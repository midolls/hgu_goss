* NGSPICE file created from hgu_cdac_half_flat.ext - technology: sky130A

.subckt hgu_cdac_half_flat d<5> db<4> d<3> db<1> db<2> d<2> db<6> db<5> db<0> d<4> d<6> d<1> d<0> db<3>
+ VSS VREF t<6> t<5> t<4> t<3> t<2> t<1> t<0> tb<6> tb<5> tb<4> tb<3> tb<2> tb<1> tb<0> VDD
X0 VREF d<3> hgu_cdac_8bit_array_3.drv<7:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1 VREF db<3> hgu_cdac_8bit_array_2.drv<7:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.35
X2 hgu_cdac_8bit_array_2.drv<31:0> db<5> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3 hgu_cdac_8bit_array_3.drv<63:0> d<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.35
X4 VREF d<5> hgu_cdac_8bit_array_3.drv<31:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X5 hgu_cdac_8bit_array_3.drv<63:0> d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X6 hgu_cdac_8bit_array_3.drv<31:0> d<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X7 VSS db<6> hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X8 VREF db<6> hgu_cdac_8bit_array_2.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X9 hgu_cdac_8bit_array_3.drv<63:0> d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X10 VREF d<4> hgu_cdac_8bit_array_3.drv<15:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X11 VSS db<5> hgu_cdac_8bit_array_2.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X12 hgu_cdac_8bit_array_3.drv<63:0> d<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X13 VREF d<6> hgu_cdac_8bit_array_3.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X14 VSS db<6> hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X15 hgu_cdac_8bit_array_3.drv<31:0> d<5> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X16 VREF d<3> hgu_cdac_8bit_array_3.drv<7:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X17 hgu_cdac_8bit_array_3.drv<1:0> d<1> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.122 ps=1.42 w=0.42 l=0.35
X18 hgu_cdac_8bit_array_3.drv<15:0> d<4> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X19 VSS db<6> hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X20 hgu_cdac_8bit_array_3.drv<31:0> d<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X21 VREF db<6> hgu_cdac_8bit_array_2.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X22 hgu_cdac_8bit_array_2.drv<15:0> db<4> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X23 hgu_cdac_8bit_array_3.drv<63:0> d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X24 VSS db<4> hgu_cdac_8bit_array_2.drv<15:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X25 VSS db<5> hgu_cdac_8bit_array_2.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X26 VREF d<6> hgu_cdac_8bit_array_3.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X27 hgu_cdac_8bit_array_3.drv<15:0> d<4> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.35
X28 hgu_cdac_8bit_array_3.drv<15:0> d<4> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X29 hgu_cdac_8bit_array_2.drv<63:0> db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X30 hgu_cdac_8bit_array_2.drv<63:0> db<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X31 hgu_cdac_8bit_array_2.drv<1:0> db<1> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.122 ps=1.42 w=0.42 l=0.35
X32 VSS d<6> hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X33 VREF db<6> hgu_cdac_8bit_array_2.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X34 hgu_cdac_8bit_array_3.drv<63:0> d<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X35 hgu_cdac_8bit_array_2.drv<7:0> db<3> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X36 hgu_cdac_8bit_array_2.drv<31:0> db<5> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X37 VSS db<6> hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X38 VREF db<6> hgu_cdac_8bit_array_2.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X39 VREF d<6> hgu_cdac_8bit_array_3.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X40 hgu_cdac_8bit_array_2.drv<63:0> db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X41 hgu_cdac_8bit_array_3.drv<63:0> d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X42 VREF d<5> hgu_cdac_8bit_array_3.drv<31:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X43 hgu_cdac_8bit_array_2.drv<7:0> db<3> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.35
X44 VREF db<2> hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X45 VSS d<6> hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X46 VSS d<5> hgu_cdac_8bit_array_3.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X47 hgu_cdac_8bit_array_3.drv<7:0> d<3> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X48 hgu_cdac_8bit_array_3.drv<63:0> d<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X49 VSS db<6> hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X50 hgu_cdac_8bit_array_3.drv<31:0> d<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X51 VREF d<6> hgu_cdac_8bit_array_3.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X52 hgu_cdac_8bit_array_3.drv<63:0> d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X53 hgu_cdac_8bit_array_3.drv<63:0> d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X54 VSS db<5> hgu_cdac_8bit_array_2.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X55 VREF db<6> hgu_cdac_8bit_array_2.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X56 VREF d<6> hgu_cdac_8bit_array_3.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X57 hgu_cdac_8bit_array_3.drv<31:0> d<5> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X58 hgu_cdac_8bit_array_2.drv<63:0> db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X59 hgu_cdac_8bit_array_2.drv<31:0> db<5> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X60 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT db<2> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X61 VREF db<6> hgu_cdac_8bit_array_2.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.35
X62 hgu_cdac_8bit_array_2.drv<0> db<0> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.35
X63 hgu_cdac_8bit_array_3.drv<63:0> d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X64 VSS db<5> hgu_cdac_8bit_array_2.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X65 VREF db<6> hgu_cdac_8bit_array_2.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X66 VREF d<6> hgu_cdac_8bit_array_3.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X67 hgu_cdac_8bit_array_3.drv<15:0> d<4> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X68 VREF d<6> hgu_cdac_8bit_array_3.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X69 VREF d<5> hgu_cdac_8bit_array_3.drv<31:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X70 VSS d<4> hgu_cdac_8bit_array_3.drv<15:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X71 hgu_cdac_8bit_array_2.drv<63:0> db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X72 VREF db<4> hgu_cdac_8bit_array_2.drv<15:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X73 VREF d<6> hgu_cdac_8bit_array_3.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X74 VREF db<5> hgu_cdac_8bit_array_2.drv<31:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X75 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT d<2> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X76 hgu_cdac_8bit_array_2.drv<63:0> db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X77 hgu_cdac_8bit_array_2.drv<63:0> db<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X78 VREF d<4> hgu_cdac_8bit_array_3.drv<15:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X79 VREF db<6> hgu_cdac_8bit_array_2.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X80 VSS d<6> hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X81 hgu_cdac_8bit_array_2.drv<15:0> db<4> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X82 VREF d<6> hgu_cdac_8bit_array_3.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X83 VSS d<4> hgu_cdac_8bit_array_3.drv<15:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X84 hgu_cdac_8bit_array_3.drv<63:0> d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X85 hgu_cdac_8bit_array_2.drv<31:0> db<5> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.35
X86 VREF d<5> hgu_cdac_8bit_array_3.drv<31:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X87 hgu_cdac_8bit_array_3.drv<31:0> d<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.122 ps=1.42 w=0.42 l=0.35
X88 VREF db<4> hgu_cdac_8bit_array_2.drv<15:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X89 VREF db<5> hgu_cdac_8bit_array_2.drv<31:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X90 VREF d<6> hgu_cdac_8bit_array_3.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X91 VSS d<6> hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X92 hgu_cdac_8bit_array_2.drv<63:0> db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X93 VSS d<5> hgu_cdac_8bit_array_3.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X94 hgu_cdac_8bit_array_3.drv<63:0> d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X95 hgu_cdac_8bit_array_2.drv<63:0> db<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X96 hgu_cdac_8bit_array_3.drv<63:0> d<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X97 VSS db<6> hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X98 hgu_cdac_8bit_array_2.drv<15:0> db<4> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.122 ps=1.42 w=0.42 l=0.35
X99 VREF d<1> hgu_cdac_8bit_array_3.drv<1:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.35
X100 hgu_cdac_8bit_array_2.drv<15:0> db<4> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X101 hgu_cdac_8bit_array_2.drv<31:0> db<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X102 VREF db<3> hgu_cdac_8bit_array_2.drv<7:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X103 hgu_cdac_8bit_array_3.drv<63:0> d<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X104 VREF d<5> hgu_cdac_8bit_array_3.drv<31:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X105 hgu_cdac_8bit_array_2.drv<63:0> db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X106 hgu_cdac_8bit_array_3.drv<63:0> d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X107 VSS db<6> hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X108 VSS d<3> hgu_cdac_8bit_array_3.drv<7:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X109 hgu_cdac_8bit_array_3.drv<31:0> d<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X110 VREF db<6> hgu_cdac_8bit_array_2.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X111 VREF d<6> hgu_cdac_8bit_array_3.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.35
X112 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT d<2> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.35
X113 VSS d<5> hgu_cdac_8bit_array_3.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X114 hgu_cdac_8bit_array_3.drv<63:0> d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.122 ps=1.42 w=0.42 l=0.35
X115 VREF d<5> hgu_cdac_8bit_array_3.drv<31:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X116 VSS db<5> hgu_cdac_8bit_array_2.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X117 hgu_cdac_8bit_array_2.drv<63:0> db<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X118 hgu_cdac_8bit_array_2.drv<15:0> db<4> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X119 VREF db<5> hgu_cdac_8bit_array_2.drv<31:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.35
X120 VSS d<4> hgu_cdac_8bit_array_3.drv<15:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X121 hgu_cdac_8bit_array_3.drv<63:0> d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X122 VSS d<6> hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X123 VSS d<3> hgu_cdac_8bit_array_3.drv<7:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X124 hgu_cdac_8bit_array_3.drv<31:0> d<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X125 VREF db<6> hgu_cdac_8bit_array_2.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X126 hgu_cdac_8bit_array_2.drv<15:0> db<4> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X127 hgu_cdac_8bit_array_2.drv<7:0> db<3> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X128 VREF d<6> hgu_cdac_8bit_array_3.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X129 VREF db<5> hgu_cdac_8bit_array_2.drv<31:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X130 hgu_cdac_8bit_array_2.drv<63:0> db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X131 VSS db<2> hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT VSS sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.35
X132 hgu_cdac_8bit_array_3.drv<15:0> d<4> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.122 ps=1.42 w=0.42 l=0.35
X133 VSS d<6> hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X134 hgu_cdac_8bit_array_2.drv<15:0> db<4> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X135 VREF d<5> hgu_cdac_8bit_array_3.drv<31:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.35
X136 hgu_cdac_8bit_array_3.drv<0> d<0> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.244 ps=2.26 w=0.84 l=0.35
X137 VSS db<6> hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X138 VREF d<6> hgu_cdac_8bit_array_3.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X139 hgu_cdac_8bit_array_2.drv<63:0> db<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X140 hgu_cdac_8bit_array_2.drv<63:0> db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X141 hgu_cdac_8bit_array_3.drv<63:0> d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X142 VSS db<5> hgu_cdac_8bit_array_2.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X143 VSS d<6> hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X144 hgu_cdac_8bit_array_2.drv<31:0> db<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X145 VSS d<5> hgu_cdac_8bit_array_3.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X146 hgu_cdac_8bit_array_2.drv<63:0> db<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X147 hgu_cdac_8bit_array_2.drv<31:0> db<5> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X148 hgu_cdac_8bit_array_3.drv<63:0> d<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X149 hgu_cdac_8bit_array_3.drv<63:0> d<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X150 VREF d<5> hgu_cdac_8bit_array_3.drv<31:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X151 hgu_cdac_8bit_array_3.drv<31:0> d<5> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X152 VSS db<6> hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X153 VREF db<6> hgu_cdac_8bit_array_2.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X154 hgu_cdac_8bit_array_3.drv<63:0> d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X155 hgu_cdac_8bit_array_2.drv<7:0> db<3> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X156 hgu_cdac_8bit_array_2.drv<31:0> db<5> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X157 VSS db<5> hgu_cdac_8bit_array_2.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X158 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT db<2> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.122 ps=1.42 w=0.42 l=0.35
X159 VREF d<6> hgu_cdac_8bit_array_3.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X160 VSS d<6> hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X161 hgu_cdac_8bit_array_3.drv<63:0> d<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X162 VSS db<6> hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X163 hgu_cdac_8bit_array_3.drv<31:0> d<5> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X164 VREF d<2> hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT VDD sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.35
X165 VSS d<6> hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X166 VSS db<6> hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X167 VSS db<6> hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X168 hgu_cdac_8bit_array_3.drv<31:0> d<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X169 VSS db<5> hgu_cdac_8bit_array_2.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X170 VREF db<6> hgu_cdac_8bit_array_2.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X171 VREF d<6> hgu_cdac_8bit_array_3.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X172 hgu_cdac_8bit_array_3.drv<15:0> d<4> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X173 VREF d<5> hgu_cdac_8bit_array_3.drv<31:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X174 hgu_cdac_8bit_array_2.drv<63:0> db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X175 VSS db<4> hgu_cdac_8bit_array_2.drv<15:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X176 hgu_cdac_8bit_array_3.drv<63:0> d<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X177 hgu_cdac_8bit_array_3.drv<15:0> d<4> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X178 VSS d<6> hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X179 VREF db<5> hgu_cdac_8bit_array_2.drv<31:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X180 hgu_cdac_8bit_array_3.drv<31:0> d<5> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X181 VSS d<5> hgu_cdac_8bit_array_3.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X182 VSS d<6> hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X183 VREF db<6> hgu_cdac_8bit_array_2.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X184 VSS db<3> hgu_cdac_8bit_array_2.drv<7:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X185 VSS d<6> hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X186 hgu_cdac_8bit_array_3.drv<15:0> d<4> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X187 VREF db<6> hgu_cdac_8bit_array_2.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X188 VSS d<4> hgu_cdac_8bit_array_3.drv<15:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X189 hgu_cdac_8bit_array_2.drv<63:0> db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X190 VSS db<4> hgu_cdac_8bit_array_2.drv<15:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X191 hgu_cdac_8bit_array_3.drv<7:0> d<3> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X192 VREF db<4> hgu_cdac_8bit_array_2.drv<15:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X193 VREF db<5> hgu_cdac_8bit_array_2.drv<31:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X194 VREF d<6> hgu_cdac_8bit_array_3.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X195 VSS d<6> hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X196 VSS d<5> hgu_cdac_8bit_array_3.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X197 hgu_cdac_8bit_array_2.drv<63:0> db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X198 hgu_cdac_8bit_array_2.drv<63:0> db<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X199 VSS d<6> hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X200 hgu_cdac_8bit_array_2.drv<1:0> db<1> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.35
X201 hgu_cdac_8bit_array_2.drv<31:0> db<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X202 hgu_cdac_8bit_array_3.drv<63:0> d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X203 hgu_cdac_8bit_array_3.drv<7:0> d<3> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X204 hgu_cdac_8bit_array_2.drv<7:0> db<3> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X205 VSS d<1> hgu_cdac_8bit_array_3.drv<1:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.35
X206 VREF db<6> hgu_cdac_8bit_array_2.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X207 hgu_cdac_8bit_array_3.drv<63:0> d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X208 hgu_cdac_8bit_array_2.drv<63:0> db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X209 VSS d<5> hgu_cdac_8bit_array_3.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X210 hgu_cdac_8bit_array_2.drv<63:0> db<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X211 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT d<2> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.122 ps=1.42 w=0.42 l=0.35
X212 VSS d<6> hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.35
X213 hgu_cdac_8bit_array_2.drv<63:0> db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X214 VSS d<5> hgu_cdac_8bit_array_3.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X215 hgu_cdac_8bit_array_2.drv<31:0> db<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X216 hgu_cdac_8bit_array_3.drv<63:0> d<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X217 VSS db<5> hgu_cdac_8bit_array_2.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X218 VSS db<6> hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X219 VREF db<6> hgu_cdac_8bit_array_2.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X220 VREF d<6> hgu_cdac_8bit_array_3.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X221 hgu_cdac_8bit_array_2.drv<31:0> db<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X222 VREF d<5> hgu_cdac_8bit_array_3.drv<31:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X223 hgu_cdac_8bit_array_2.drv<63:0> db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X224 VSS db<1> hgu_cdac_8bit_array_2.drv<1:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.35
X225 hgu_cdac_8bit_array_2.drv<63:0> db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X226 hgu_cdac_8bit_array_2.drv<63:0> db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X227 VSS db<3> hgu_cdac_8bit_array_2.drv<7:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X228 VREF db<5> hgu_cdac_8bit_array_2.drv<31:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X229 VREF d<6> hgu_cdac_8bit_array_3.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X230 hgu_cdac_8bit_array_2.drv<63:0> db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X231 hgu_cdac_8bit_array_2.drv<63:0> db<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X232 VSS d<6> hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X233 hgu_cdac_8bit_array_2.drv<31:0> db<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X234 VREF d<5> hgu_cdac_8bit_array_3.drv<31:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X235 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT db<2> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X236 hgu_cdac_8bit_array_2.drv<63:0> db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.122 ps=1.42 w=0.42 l=0.35
X237 hgu_cdac_8bit_array_2.drv<0> db<0> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.244 ps=2.26 w=0.84 l=0.35
X238 VSS db<4> hgu_cdac_8bit_array_2.drv<15:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.35
X239 VREF db<5> hgu_cdac_8bit_array_2.drv<31:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X240 VREF d<6> hgu_cdac_8bit_array_3.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X241 hgu_cdac_8bit_array_2.drv<63:0> db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X242 hgu_cdac_8bit_array_3.drv<0> d<0> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.35
X243 VSS d<5> hgu_cdac_8bit_array_3.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.35
X244 hgu_cdac_8bit_array_2.drv<63:0> db<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X245 VSS d<6> hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X246 hgu_cdac_8bit_array_2.drv<15:0> db<4> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X247 hgu_cdac_8bit_array_2.drv<31:0> db<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X248 hgu_cdac_8bit_array_2.drv<63:0> db<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X249 hgu_cdac_8bit_array_3.drv<63:0> d<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X250 VREF d<5> hgu_cdac_8bit_array_3.drv<31:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X251 VSS db<6> hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X252 VREF d<3> hgu_cdac_8bit_array_3.drv<7:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.35
X253 hgu_cdac_8bit_array_2.drv<15:0> db<4> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X254 hgu_cdac_8bit_array_3.drv<63:0> d<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X255 hgu_cdac_8bit_array_3.drv<63:0> d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X256 hgu_cdac_8bit_array_3.drv<63:0> d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X257 VSS d<5> hgu_cdac_8bit_array_3.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X258 VSS db<6> hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X259 hgu_cdac_8bit_array_3.drv<31:0> d<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X260 hgu_cdac_8bit_array_2.drv<63:0> db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X261 hgu_cdac_8bit_array_2.drv<31:0> db<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X262 hgu_cdac_8bit_array_2.drv<63:0> db<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X263 hgu_cdac_8bit_array_3.drv<63:0> d<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X264 VREF d<4> hgu_cdac_8bit_array_3.drv<15:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.35
X265 hgu_cdac_8bit_array_3.drv<31:0> d<5> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X266 VSS d<6> hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X267 VSS db<6> hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X268 VREF d<3> hgu_cdac_8bit_array_3.drv<7:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X269 VREF db<6> hgu_cdac_8bit_array_2.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X270 hgu_cdac_8bit_array_2.drv<15:0> db<4> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.35
X271 hgu_cdac_8bit_array_2.drv<31:0> db<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X272 hgu_cdac_8bit_array_3.drv<63:0> d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X273 hgu_cdac_8bit_array_2.drv<15:0> db<4> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X274 hgu_cdac_8bit_array_3.drv<63:0> d<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X275 hgu_cdac_8bit_array_2.drv<31:0> db<5> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X276 VSS d<2> hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT VSS sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.35
X277 hgu_cdac_8bit_array_3.drv<31:0> d<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X278 hgu_cdac_8bit_array_2.drv<63:0> db<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X279 VREF db<6> hgu_cdac_8bit_array_2.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X280 VREF d<6> hgu_cdac_8bit_array_3.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X281 hgu_cdac_8bit_array_3.drv<15:0> d<4> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X282 hgu_cdac_8bit_array_2.drv<63:0> db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X283 VSS db<4> hgu_cdac_8bit_array_2.drv<15:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X284 hgu_cdac_8bit_array_3.drv<31:0> d<5> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X285 hgu_cdac_8bit_array_3.drv<15:0> d<4> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X286 VSS d<6> hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X287 VREF db<5> hgu_cdac_8bit_array_2.drv<31:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X288 VSS d<5> hgu_cdac_8bit_array_3.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X289 hgu_cdac_8bit_array_2.drv<15:0> db<4> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X290 hgu_cdac_8bit_array_3.drv<63:0> d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X291 hgu_cdac_8bit_array_3.drv<31:0> d<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X292 VREF d<6> hgu_cdac_8bit_array_3.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X293 hgu_cdac_8bit_array_2.drv<63:0> db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X294 VSS db<4> hgu_cdac_8bit_array_2.drv<15:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X295 hgu_cdac_8bit_array_3.drv<15:0> d<4> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X296 hgu_cdac_8bit_array_2.drv<7:0> db<3> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X297 hgu_cdac_8bit_array_3.drv<7:0> d<3> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X298 hgu_cdac_8bit_array_2.drv<63:0> db<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X299 VREF d<2> hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X300 VREF db<2> hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT VDD sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.35
X301 VSS d<6> hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X302 hgu_cdac_8bit_array_3.drv<31:0> d<5> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X303 VSS db<6> hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X304 VREF db<6> hgu_cdac_8bit_array_2.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X305 hgu_cdac_8bit_array_3.drv<7:0> d<3> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X306 hgu_cdac_8bit_array_2.drv<63:0> db<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X307 hgu_cdac_8bit_array_3.drv<63:0> d<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X308 VSS db<5> hgu_cdac_8bit_array_2.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X309 VREF db<5> hgu_cdac_8bit_array_2.drv<31:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X310 VREF d<6> hgu_cdac_8bit_array_3.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X311 hgu_cdac_8bit_array_3.drv<31:0> d<5> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X312 hgu_cdac_8bit_array_2.drv<63:0> db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X313 hgu_cdac_8bit_array_3.drv<63:0> d<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X314 VSS db<6> hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X315 hgu_cdac_8bit_array_2.drv<31:0> db<5> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X316 VSS db<6> hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X317 VREF db<6> hgu_cdac_8bit_array_2.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X318 hgu_cdac_8bit_array_3.drv<63:0> d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X319 VSS db<5> hgu_cdac_8bit_array_2.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X320 hgu_cdac_8bit_array_2.drv<7:0> db<3> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X321 VSS d<6> hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X322 VREF db<5> hgu_cdac_8bit_array_2.drv<31:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X323 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT db<2> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.35
X324 VSS d<5> hgu_cdac_8bit_array_3.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X325 hgu_cdac_8bit_array_2.drv<63:0> db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X326 hgu_cdac_8bit_array_3.drv<63:0> d<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X327 VREF db<6> hgu_cdac_8bit_array_2.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X328 VSS db<6> hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X329 VSS d<6> hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X330 VREF db<6> hgu_cdac_8bit_array_2.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X331 hgu_cdac_8bit_array_3.drv<15:0> d<4> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X332 hgu_cdac_8bit_array_2.drv<31:0> db<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X333 VREF db<6> hgu_cdac_8bit_array_2.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X334 VREF d<4> hgu_cdac_8bit_array_3.drv<15:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X335 hgu_cdac_8bit_array_2.drv<63:0> db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X336 VREF d<5> hgu_cdac_8bit_array_3.drv<31:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X337 hgu_cdac_8bit_array_3.drv<7:0> d<3> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.35
X338 VSS db<6> hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X339 VSS db<5> hgu_cdac_8bit_array_2.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X340 VREF db<5> hgu_cdac_8bit_array_2.drv<31:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X341 VREF d<6> hgu_cdac_8bit_array_3.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X342 VREF d<6> hgu_cdac_8bit_array_3.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X343 hgu_cdac_8bit_array_3.drv<31:0> d<5> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X344 VSS d<5> hgu_cdac_8bit_array_3.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X345 hgu_cdac_8bit_array_2.drv<63:0> db<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X346 VREF db<4> hgu_cdac_8bit_array_2.drv<15:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X347 VSS d<6> hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X348 VSS db<3> hgu_cdac_8bit_array_2.drv<7:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.35
X349 hgu_cdac_8bit_array_2.drv<31:0> db<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X350 VSS db<6> hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X351 VREF db<3> hgu_cdac_8bit_array_2.drv<7:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X352 VREF d<6> hgu_cdac_8bit_array_3.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X353 hgu_cdac_8bit_array_3.drv<63:0> d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X354 VSS d<5> hgu_cdac_8bit_array_3.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X355 hgu_cdac_8bit_array_2.drv<63:0> db<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X356 VREF db<4> hgu_cdac_8bit_array_2.drv<15:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X357 VSS d<3> hgu_cdac_8bit_array_3.drv<7:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.35
X358 hgu_cdac_8bit_array_3.drv<63:0> d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X359 hgu_cdac_8bit_array_2.drv<63:0> db<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X360 hgu_cdac_8bit_array_3.drv<63:0> d<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X361 VREF d<4> hgu_cdac_8bit_array_3.drv<15:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X362 hgu_cdac_8bit_array_3.drv<31:0> d<5> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X363 VSS db<6> hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X364 hgu_cdac_8bit_array_2.drv<15:0> db<4> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X365 VSS d<4> hgu_cdac_8bit_array_3.drv<15:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.35
X366 hgu_cdac_8bit_array_3.drv<63:0> d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X367 hgu_cdac_8bit_array_2.drv<31:0> db<5> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X368 hgu_cdac_8bit_array_3.drv<31:0> d<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X369 VSS d<3> hgu_cdac_8bit_array_3.drv<7:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X370 VREF d<6> hgu_cdac_8bit_array_3.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X371 hgu_cdac_8bit_array_2.drv<63:0> db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X372 hgu_cdac_8bit_array_3.drv<63:0> d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X373 hgu_cdac_8bit_array_3.drv<63:0> d<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X374 VREF d<4> hgu_cdac_8bit_array_3.drv<15:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X375 hgu_cdac_8bit_array_2.drv<63:0> db<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X376 VREF d<6> hgu_cdac_8bit_array_3.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X377 hgu_cdac_8bit_array_3.drv<15:0> d<4> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X378 VSS db<6> hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X379 VSS d<6> hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X380 hgu_cdac_8bit_array_2.drv<31:0> db<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X381 hgu_cdac_8bit_array_2.drv<63:0> db<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X382 hgu_cdac_8bit_array_2.drv<31:0> db<5> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X383 VSS db<6> hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X384 hgu_cdac_8bit_array_3.drv<31:0> d<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X385 VREF db<6> hgu_cdac_8bit_array_2.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X386 VREF db<5> hgu_cdac_8bit_array_2.drv<31:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X387 VREF d<6> hgu_cdac_8bit_array_3.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X388 hgu_cdac_8bit_array_2.drv<7:0> db<3> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.122 ps=1.42 w=0.42 l=0.35
X389 hgu_cdac_8bit_array_2.drv<31:0> db<5> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X390 VSS db<2> hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X391 hgu_cdac_8bit_array_2.drv<63:0> db<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X392 VREF db<1> hgu_cdac_8bit_array_2.drv<1:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.35
X393 VSS d<6> hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X394 hgu_cdac_8bit_array_2.drv<63:0> db<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X395 hgu_cdac_8bit_array_2.drv<63:0> db<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X396 VREF db<3> hgu_cdac_8bit_array_2.drv<7:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X397 hgu_cdac_8bit_array_2.drv<63:0> db<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X398 hgu_cdac_8bit_array_3.drv<63:0> d<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X399 hgu_cdac_8bit_array_3.drv<63:0> d<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X400 hgu_cdac_8bit_array_2.drv<31:0> db<5> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X401 VREF d<5> hgu_cdac_8bit_array_3.drv<31:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X402 VSS d<2> hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X403 VSS db<6> hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X404 hgu_cdac_8bit_array_3.drv<31:0> d<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X405 hgu_cdac_8bit_array_2.drv<63:0> db<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.35
X406 VREF db<4> hgu_cdac_8bit_array_2.drv<15:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.35
X407 hgu_cdac_8bit_array_2.drv<31:0> db<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X408 hgu_cdac_8bit_array_2.drv<63:0> db<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X409 hgu_cdac_8bit_array_3.drv<63:0> d<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X410 hgu_cdac_8bit_array_3.drv<31:0> d<5> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X411 VSS db<6> hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.35
X412 hgu_cdac_8bit_array_2.drv<15:0> db<4> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X413 hgu_cdac_8bit_array_3.drv<63:0> d<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X414 hgu_cdac_8bit_array_3.drv<63:0> d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X415 VSS db<6> hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X416 hgu_cdac_8bit_array_2.drv<31:0> db<5> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X417 hgu_cdac_8bit_array_3.drv<31:0> d<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X418 VSS d<6> hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X419 VREF db<6> hgu_cdac_8bit_array_2.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X420 hgu_cdac_8bit_array_3.drv<1:0> d<1> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.35
X421 hgu_cdac_8bit_array_3.drv<63:0> d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X422 VSS db<4> hgu_cdac_8bit_array_2.drv<15:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X423 VSS db<5> hgu_cdac_8bit_array_2.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X424 hgu_cdac_8bit_array_3.drv<15:0> d<4> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X425 VREF db<6> hgu_cdac_8bit_array_2.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X426 hgu_cdac_8bit_array_3.drv<31:0> d<5> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X427 hgu_cdac_8bit_array_2.drv<63:0> db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X428 VSS db<6> hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X429 hgu_cdac_8bit_array_2.drv<63:0> db<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X430 hgu_cdac_8bit_array_2.drv<31:0> db<5> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X431 hgu_cdac_8bit_array_3.drv<63:0> d<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X432 hgu_cdac_8bit_array_3.drv<15:0> d<4> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X433 hgu_cdac_8bit_array_2.drv<31:0> db<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.122 ps=1.42 w=0.42 l=0.35
X434 VREF db<6> hgu_cdac_8bit_array_2.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X435 hgu_cdac_8bit_array_3.drv<63:0> d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X436 VSS db<4> hgu_cdac_8bit_array_2.drv<15:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X437 hgu_cdac_8bit_array_2.drv<31:0> db<5> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X438 VSS db<5> hgu_cdac_8bit_array_2.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X439 hgu_cdac_8bit_array_3.drv<15:0> d<4> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X440 VREF d<6> hgu_cdac_8bit_array_3.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X441 VSS d<4> hgu_cdac_8bit_array_3.drv<15:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X442 hgu_cdac_8bit_array_2.drv<63:0> db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X443 hgu_cdac_8bit_array_3.drv<7:0> d<3> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.122 ps=1.42 w=0.42 l=0.35
X444 VSS d<5> hgu_cdac_8bit_array_3.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X445 hgu_cdac_8bit_array_2.drv<63:0> db<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X446 VREF db<4> hgu_cdac_8bit_array_2.drv<15:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X447 VSS d<6> hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X448 VSS d<6> hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X449 VSS db<3> hgu_cdac_8bit_array_2.drv<7:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X450 hgu_cdac_8bit_array_3.drv<31:0> d<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X451 hgu_cdac_8bit_array_3.drv<63:0> d<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X452 VSS db<6> hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X453 VREF d<6> hgu_cdac_8bit_array_3.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X454 VREF d<5> hgu_cdac_8bit_array_3.drv<31:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X455 hgu_cdac_8bit_array_2.drv<63:0> db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X456 hgu_cdac_8bit_array_3.drv<7:0> d<3> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X457 hgu_cdac_8bit_array_2.drv<63:0> db<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X458 VREF db<4> hgu_cdac_8bit_array_2.drv<15:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X459 VSS db<5> hgu_cdac_8bit_array_2.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.35
X460 VSS d<6> hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X461 hgu_cdac_8bit_array_3.drv<31:0> d<5> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X462 hgu_cdac_8bit_array_3.drv<63:0> d<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X463 hgu_cdac_8bit_array_3.drv<63:0> d<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X464 VSS db<6> hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X465 hgu_cdac_8bit_array_2.drv<15:0> db<4> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X466 VSS d<4> hgu_cdac_8bit_array_3.drv<15:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X467 hgu_cdac_8bit_array_3.drv<63:0> d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X468 VSS db<5> hgu_cdac_8bit_array_2.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X469 hgu_cdac_8bit_array_3.drv<31:0> d<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X470 VREF db<6> hgu_cdac_8bit_array_2.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X471 hgu_cdac_8bit_array_3.drv<63:0> d<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X472 VSS d<6> hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X473 hgu_cdac_8bit_array_2.drv<15:0> db<4> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X474 VREF db<5> hgu_cdac_8bit_array_2.drv<31:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X475 VSS d<4> hgu_cdac_8bit_array_3.drv<15:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X476 hgu_cdac_8bit_array_2.drv<63:0> db<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X477 VREF d<4> hgu_cdac_8bit_array_3.drv<15:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X478 hgu_cdac_8bit_array_3.drv<63:0> d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X479 VSS d<6> hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X480 VREF db<6> hgu_cdac_8bit_array_2.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X481 hgu_cdac_8bit_array_2.drv<63:0> db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X482 VREF db<6> hgu_cdac_8bit_array_2.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X483 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT d<2> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X484 VREF d<6> hgu_cdac_8bit_array_3.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X485 VREF db<5> hgu_cdac_8bit_array_2.drv<31:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X486 VSS d<6> hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X487 hgu_cdac_8bit_array_2.drv<63:0> db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X488 hgu_cdac_8bit_array_2.drv<31:0> db<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X489 hgu_cdac_8bit_array_2.drv<63:0> db<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X490 hgu_cdac_8bit_array_3.drv<63:0> d<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X491 VREF d<4> hgu_cdac_8bit_array_3.drv<15:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X492 hgu_cdac_8bit_array_3.drv<31:0> d<5> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.35
X493 VSS db<6> hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X494 VREF db<6> hgu_cdac_8bit_array_2.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X495 VREF d<6> hgu_cdac_8bit_array_3.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X496 hgu_cdac_8bit_array_2.drv<31:0> db<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X497 hgu_cdac_8bit_array_2.drv<31:0> db<5> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X498 hgu_cdac_8bit_array_3.drv<63:0> d<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X499 VREF d<5> hgu_cdac_8bit_array_3.drv<31:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X500 hgu_cdac_8bit_array_3.drv<63:0> d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X501 hgu_cdac_8bit_array_2.drv<63:0> db<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X502 VREF db<6> hgu_cdac_8bit_array_2.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X503 VREF db<5> hgu_cdac_8bit_array_2.drv<31:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X504 VSS d<5> hgu_cdac_8bit_array_3.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X505 hgu_cdac_8bit_array_3.drv<63:0> d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X506 hgu_cdac_8bit_array_3.drv<63:0> d<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X507 hgu_cdac_8bit_array_3.drv<31:0> d<5> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
C0 t<6> hgu_cdac_8bit_array_3.drv<63:0> 0.328p
C1 tb<3> hgu_cdac_8bit_array_2.drv<7:0> 42.3f
C2 hgu_cdac_8bit_array_3.drv<15:0> d<4> 1.03f
C3 VREF hgu_cdac_8bit_array_3.drv<31:0> 5.04f
C4 hgu_cdac_8bit_array_3.drv<15:0> hgu_cdac_8bit_array_2.drv<15:0> 2.96f
C5 hgu_cdac_8bit_array_2.drv<7:0> hgu_cdac_8bit_array_2.drv<15:0> 2.27f
C6 tb<6> hgu_cdac_8bit_array_2.drv<63:0> 0.325p
C7 VREF VDD 49.1f
C8 hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_8bit_array_3.drv<63:0> 2.29f
C9 hgu_cdac_8bit_array_2.drv<7:0> hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT 1.08f
C10 hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_8bit_array_3.drv<15:0> 2.29f
C11 hgu_cdac_8bit_array_3.drv<63:0> VDD 1.5f
C12 tb<2> hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT 22.1f
C13 VREF d<6> 1.75f
C14 t<6> tb<6> 4.02f
C15 hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_8bit_array_2.drv<63:0> 2.28f
C16 VREF hgu_cdac_8bit_array_2.drv<31:0> 4.1f
C17 d<6> hgu_cdac_8bit_array_3.drv<63:0> 4.14f
C18 t<4> hgu_cdac_8bit_array_2.drv<15:0> 1.55f
C19 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT hgu_cdac_8bit_array_2.drv<1:0> 1.14f
C20 hgu_cdac_8bit_array_3.drv<7:0> hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT 1.06f
C21 hgu_cdac_8bit_array_3.drv<31:0> d<5> 2.09f
C22 hgu_cdac_8bit_array_3.drv<15:0> t<4> 83.1f
C23 tb<0> hgu_cdac_8bit_array_2.drv<0> 5.12f
C24 tb<4> hgu_cdac_8bit_array_2.drv<15:0> 82.5f
C25 t<3> hgu_cdac_8bit_array_3.drv<7:0> 42.6f
C26 hgu_cdac_8bit_array_3.drv<1:0> hgu_cdac_8bit_array_3.drv<0> 1.19f
C27 d<5> VDD 2f
C28 hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_8bit_array_2.drv<15:0> 2.28f
C29 t<0> hgu_cdac_8bit_array_3.drv<0> 5.11f
C30 d<6> VDD 4f
C31 hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_8bit_array_2.drv<31:0> 3.77f
C32 hgu_cdac_8bit_array_3.drv<1:0> hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT 1.11f
C33 hgu_cdac_8bit_array_3.drv<31:0> t<5> 0.165p
C34 db<6> hgu_cdac_8bit_array_2.drv<63:0> 3.93f
C35 VREF hgu_cdac_8bit_array_3.drv<7:0> 1.44f
C36 tb<1> hgu_cdac_8bit_array_2.drv<1:0> 11.5f
C37 VREF db<6> 1.76f
C38 t<4> tb<4> 1.12f
C39 hgu_cdac_unit_0.CBOT tb<0> 5.11f
C40 hgu_cdac_8bit_array_3.drv<7:0> hgu_cdac_8bit_array_3.drv<15:0> 2.83f
C41 hgu_cdac_8bit_array_2.drv<7:0> hgu_cdac_8bit_array_3.drv<7:0> 1.81f
C42 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT 2.13f
C43 t<2> hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT 22.2f
C44 VREF hgu_cdac_8bit_array_2.drv<63:0> 8.33f
C45 db<5> VDD 2f
C46 hgu_cdac_8bit_array_2.drv<31:0> t<5> 2.38f
C47 hgu_cdac_8bit_array_3.drv<1:0> t<1> 11.6f
C48 hgu_cdac_unit_1.CBOT t<0> 5.11f
C49 hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_8bit_array_2.drv<63:0> 7.25f
C50 t<6> hgu_cdac_8bit_array_2.drv<63:0> 4.72f
C51 VREF hgu_cdac_8bit_array_3.drv<63:0> 9.96f
C52 tb<5> hgu_cdac_8bit_array_2.drv<31:0> 0.163p
C53 db<6> VDD 4f
C54 VREF hgu_cdac_8bit_array_2.drv<15:0> 2.12f
C55 tb<5> t<5> 2.08f
C56 VREF hgu_cdac_8bit_array_3.drv<15:0> 2.69f
C57 hgu_cdac_8bit_array_2.drv<31:0> db<5> 1.88f
C58 VREF hgu_cdac_8bit_array_2.drv<7:0> 1.07f
C59 db<6> VSS 12.7f
C60 db<5> VSS 6.38f
C61 db<4> VSS 3.21f
C62 db<3> VSS 1.58f
C63 d<6> VSS 12.7f
C64 d<5> VSS 6.38f
C65 d<4> VSS 3.21f
C66 d<3> VSS 1.58f
C67 tb<6> VSS 24.1f
C68 tb<5> VSS 12.5f
C69 tb<4> VSS 6.78f
C70 tb<3> VSS 3.61f
C71 tb<2> VSS 1.91f
C72 tb<1> VSS 1.63f
C73 t<6> VSS 23.4f
C74 t<5> VSS 12.3f
C75 t<4> VSS 6.6f
C76 t<3> VSS 3.5f
C77 t<2> VSS 1.82f
C78 t<1> VSS 1.6f
C79 hgu_cdac_8bit_array_2.drv<63:0> VSS 36.4f
C80 hgu_cdac_8bit_array_2.drv<31:0> VSS 18.2f
C81 hgu_cdac_8bit_array_2.drv<15:0> VSS 9.87f
C82 hgu_cdac_8bit_array_2.drv<7:0> VSS 5.42f
C83 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT VSS 3.37f
C84 hgu_cdac_8bit_array_2.drv<1:0> VSS 1.93f
C85 hgu_cdac_8bit_array_2.drv<0> VSS 2.22f
C86 VREF VSS 13.4f
C87 hgu_cdac_8bit_array_3.drv<63:0> VSS 33f
C88 hgu_cdac_8bit_array_3.drv<31:0> VSS 16.7f
C89 hgu_cdac_8bit_array_3.drv<15:0> VSS 9f
C90 hgu_cdac_8bit_array_3.drv<7:0> VSS 5.25f
C91 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT VSS 2.8f
C92 hgu_cdac_8bit_array_3.drv<1:0> VSS 1.57f
C93 hgu_cdac_8bit_array_3.drv<0> VSS 1.83f
C94 VDD VSS 49.1f
.ends

