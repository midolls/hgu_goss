magic
tech sky130A
magscale 1 2
timestamp 1698045515
<< checkpaint >>
rect -891 2201 2051 4160
rect 3590 2201 7323 3630
rect -891 1830 7323 2201
rect -891 1034 8061 1830
rect 954 504 8061 1034
rect 954 -925 3896 504
rect 5119 -1296 8061 504
<< error_s >>
rect 405 2851 440 2864
rect 369 2830 440 2851
rect 182 2713 240 2719
rect 182 2679 194 2713
rect 182 2673 240 2679
rect 182 2519 240 2525
rect 182 2485 194 2519
rect 182 2479 240 2485
rect 369 2383 439 2830
rect 551 2762 609 2768
rect 551 2728 563 2762
rect 551 2722 609 2728
rect 551 2466 609 2472
rect 551 2432 563 2466
rect 551 2426 609 2432
rect 369 2347 422 2383
rect 4886 2321 4921 2334
rect 5677 2321 5712 2334
rect 4850 2300 4921 2321
rect 5641 2300 5712 2321
rect 4663 2183 4721 2189
rect 4663 2149 4675 2183
rect 4663 2143 4721 2149
rect 4663 1989 4721 1995
rect 4663 1955 4675 1989
rect 4663 1949 4721 1955
rect 4850 1853 4920 2300
rect 5032 2232 5090 2238
rect 5032 2198 5044 2232
rect 5032 2192 5090 2198
rect 5454 2183 5512 2189
rect 5454 2149 5466 2183
rect 5454 2143 5512 2149
rect 5454 1989 5512 1995
rect 5454 1955 5466 1989
rect 5454 1949 5512 1955
rect 5032 1936 5090 1942
rect 5032 1902 5044 1936
rect 5032 1896 5090 1902
rect 5641 1853 5711 2300
rect 5823 2232 5881 2238
rect 5823 2198 5835 2232
rect 5823 2192 5881 2198
rect 5823 1936 5881 1942
rect 5823 1902 5835 1936
rect 5823 1896 5881 1902
rect 4850 1817 4903 1853
rect 5641 1817 5694 1853
rect 1089 1251 1124 1285
rect 1090 1232 1124 1251
rect 920 1183 978 1189
rect 920 1149 932 1183
rect 920 1143 978 1149
rect 920 719 978 725
rect 920 685 932 719
rect 920 679 978 685
rect 1109 583 1124 1232
rect 1143 1198 1178 1232
rect 1143 583 1177 1198
rect 1289 1130 1347 1136
rect 1289 1096 1301 1130
rect 1289 1090 1347 1096
rect 1459 1029 1493 1047
rect 1459 993 1529 1029
rect 1476 959 1547 993
rect 1827 959 1862 993
rect 1289 666 1347 672
rect 1289 632 1301 666
rect 1289 626 1347 632
rect 1143 549 1158 583
rect 1476 530 1546 959
rect 1828 940 1862 959
rect 2214 940 2267 941
rect 1658 891 1716 897
rect 1658 857 1670 891
rect 1658 851 1716 857
rect 1658 613 1716 619
rect 1658 579 1670 613
rect 1658 573 1716 579
rect 1476 494 1529 530
rect 1847 477 1862 940
rect 1881 906 1916 940
rect 2196 906 2267 940
rect 1881 477 1915 906
rect 2197 905 2267 906
rect 2214 871 2285 905
rect 2027 838 2085 844
rect 2027 804 2039 838
rect 2027 798 2085 804
rect 2027 560 2085 566
rect 2027 526 2039 560
rect 2027 520 2085 526
rect 1881 443 1896 477
rect 2214 424 2284 871
rect 4041 827 4076 861
rect 2396 803 2454 809
rect 4042 808 4076 827
rect 2396 769 2408 803
rect 2566 786 2600 804
rect 2396 763 2454 769
rect 2566 750 2636 786
rect 2583 716 2654 750
rect 2396 507 2454 513
rect 2396 473 2408 507
rect 2396 467 2454 473
rect 2214 388 2267 424
rect 2583 371 2653 716
rect 2765 648 2823 654
rect 2765 614 2777 648
rect 2765 608 2823 614
rect 2765 454 2823 460
rect 2765 420 2777 454
rect 2765 414 2823 420
rect 2583 335 2636 371
rect 2954 318 2969 750
rect 2988 747 3023 781
rect 3303 747 3338 781
rect 3726 764 3760 782
rect 2988 318 3022 747
rect 3304 728 3338 747
rect 3134 679 3192 685
rect 3134 645 3146 679
rect 3134 639 3192 645
rect 3134 401 3192 407
rect 3134 367 3146 401
rect 3134 361 3192 367
rect 2988 284 3003 318
rect 3323 265 3338 728
rect 3357 694 3392 728
rect 3357 265 3391 694
rect 3503 626 3561 632
rect 3503 592 3515 626
rect 3503 586 3561 592
rect 3503 348 3561 354
rect 3503 314 3515 348
rect 3503 308 3561 314
rect 3357 231 3372 265
rect 3690 212 3760 764
rect 3872 759 3930 765
rect 3872 725 3884 759
rect 3872 719 3930 725
rect 3872 295 3930 301
rect 3872 261 3884 295
rect 3872 255 3930 261
rect 3690 176 3743 212
rect 4061 159 4076 808
rect 4095 774 4130 808
rect 4095 159 4129 774
rect 4241 706 4299 712
rect 4241 672 4253 706
rect 4241 666 4299 672
rect 6192 383 6250 389
rect 6192 349 6204 383
rect 6192 343 6250 349
rect 4241 242 4299 248
rect 4241 208 4253 242
rect 4241 202 4299 208
rect 6192 189 6250 195
rect 4095 125 4110 159
rect 6192 155 6204 189
rect 6192 149 6250 155
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
rect 0 -2400 200 -2200
rect 0 -2800 200 -2600
use inverter  x1
timestamp 1698045514
transform 1 0 53 0 1 1800
box -53 -1200 738 1100
use inverter  x2
timestamp 1698045514
transform 1 0 4534 0 1 1270
box -53 -1200 738 1100
use inverter  x3
timestamp 1698045514
transform 1 0 5325 0 1 1270
box -53 -1200 738 1100
use sky130_fd_pr__pfet_01v8_MQX2PY  XM1
timestamp 0
transform 1 0 2425 0 1 638
box -211 -303 211 303
use sky130_fd_pr__pfet_01v8_XY4TMQ  XM2
timestamp 0
transform 1 0 949 0 1 934
box -211 -387 211 387
use sky130_fd_pr__pfet_01v8_XY4TMQ  XM3
timestamp 0
transform 1 0 1318 0 1 881
box -211 -387 211 387
use sky130_fd_pr__nfet_01v8_L7T3GD  XM4
timestamp 0
transform 1 0 2794 0 1 534
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_9NW3WL  XM5
timestamp 0
transform 1 0 3163 0 1 523
box -211 -294 211 294
use sky130_fd_pr__nfet_01v8_9NW3WL  XM6
timestamp 0
transform 1 0 3532 0 1 470
box -211 -294 211 294
use sky130_fd_pr__pfet_01v8_XY4TMQ  XM7
timestamp 0
transform 1 0 3901 0 1 510
box -211 -387 211 387
use sky130_fd_pr__pfet_01v8_XY4TMQ  XM8
timestamp 0
transform 1 0 4270 0 1 457
box -211 -387 211 387
use sky130_fd_pr__nfet_01v8_9NW3WL  XM9
timestamp 0
transform 1 0 1687 0 1 735
box -211 -294 211 294
use sky130_fd_pr__nfet_01v8_9NW3WL  XM10
timestamp 0
transform 1 0 2056 0 1 682
box -211 -294 211 294
use sky130_fd_pr__nfet_01v8_L7T3GD  XM11
timestamp 0
transform 1 0 6221 0 1 269
box -211 -252 211 252
use sky130_fd_pr__pfet_01v8_MQX2PY  XM12
timestamp 0
transform 1 0 6590 0 1 267
box -211 -303 211 303
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 D
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 Qb
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 Q
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 CLK
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 VDD
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 VSS
port 5 nsew
flabel metal1 0 -2400 200 -2200 0 FreeSans 256 0 0 0 SET
port 6 nsew
flabel metal1 0 -2800 200 -2600 0 FreeSans 256 0 0 0 RESET
port 7 nsew
<< end >>
