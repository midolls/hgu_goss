magic
tech sky130A
magscale 1 2
timestamp 1698050879
<< error_s >>
rect 154 586 204 624
rect 230 586 292 624
rect 306 586 380 624
rect 394 586 456 624
rect 482 586 532 624
rect 322 225 364 259
rect 154 6 204 44
rect 230 6 292 44
rect 306 6 380 44
rect 394 6 456 44
rect 482 6 532 44
<< nwell >>
rect 88 279 510 665
<< nmos >>
rect 284 102 314 186
<< pmos >>
rect 284 318 314 486
<< ndiff >>
rect 226 174 284 186
rect 226 114 238 174
rect 272 114 284 174
rect 226 102 284 114
rect 314 174 372 186
rect 314 114 326 174
rect 360 114 372 174
rect 314 102 372 114
<< pdiff >>
rect 226 474 284 486
rect 226 421 238 474
rect 272 421 284 474
rect 226 383 284 421
rect 226 330 238 383
rect 272 330 284 383
rect 226 318 284 330
rect 314 474 372 486
rect 314 421 326 474
rect 360 421 372 474
rect 314 383 372 421
rect 314 330 326 383
rect 360 330 372 383
rect 314 318 372 330
<< ndiffc >>
rect 238 114 272 174
rect 326 114 360 174
<< pdiffc >>
rect 238 421 272 474
rect 238 330 272 383
rect 326 421 360 474
rect 326 330 360 383
<< psubdiff >>
rect 124 44 474 48
rect 124 6 166 44
rect 204 6 242 44
rect 280 6 318 44
rect 356 6 394 44
rect 432 6 474 44
rect 124 2 474 6
<< nsubdiff >>
rect 124 624 474 628
rect 124 586 166 624
rect 204 586 242 624
rect 280 586 318 624
rect 356 586 394 624
rect 432 586 474 624
rect 124 582 474 586
<< psubdiffcont >>
rect 166 6 204 44
rect 242 6 280 44
rect 318 6 356 44
rect 394 6 432 44
<< nsubdiffcont >>
rect 166 586 204 624
rect 242 586 280 624
rect 318 586 356 624
rect 394 586 432 624
<< poly >>
rect 284 486 314 517
rect 284 275 314 318
rect 284 259 380 275
rect 284 225 330 259
rect 364 225 380 259
rect 284 209 380 225
rect 284 186 314 209
rect 284 76 314 102
<< polycont >>
rect 330 225 364 259
<< locali >>
rect 88 624 510 628
rect 88 586 166 624
rect 204 586 242 624
rect 280 586 318 624
rect 356 586 394 624
rect 432 586 510 624
rect 88 582 510 586
rect 238 474 272 490
rect 238 383 272 421
rect 238 174 272 330
rect 326 474 360 490
rect 326 383 360 421
rect 326 314 360 330
rect 314 225 330 259
rect 364 225 380 259
rect 238 98 272 114
rect 326 174 360 190
rect 326 48 360 114
rect 88 44 510 48
rect 88 6 166 44
rect 204 6 242 44
rect 280 6 318 44
rect 356 6 394 44
rect 432 6 510 44
rect 88 2 510 6
<< viali >>
rect 166 586 204 624
rect 242 586 280 624
rect 318 586 356 624
rect 394 586 432 624
rect 238 421 272 474
rect 238 330 272 383
rect 326 421 360 474
rect 326 330 360 383
rect 330 225 364 259
rect 238 114 272 174
rect 326 114 360 174
rect 166 6 204 44
rect 242 6 280 44
rect 318 6 356 44
rect 394 6 432 44
<< metal1 >>
rect 88 624 510 630
rect 88 586 166 624
rect 204 586 242 624
rect 280 586 318 624
rect 356 586 394 624
rect 432 586 510 624
rect 88 580 510 586
rect 88 519 510 551
rect 232 474 278 486
rect 232 421 238 474
rect 272 421 278 474
rect 232 383 278 421
rect 232 330 238 383
rect 272 330 278 383
rect 232 318 278 330
rect 320 474 366 491
rect 320 421 326 474
rect 360 421 366 474
rect 320 383 366 421
rect 320 330 326 383
rect 360 330 366 383
rect 320 318 366 330
rect 314 259 380 269
rect 314 225 330 259
rect 364 225 380 259
rect 314 215 380 225
rect 232 174 278 186
rect 232 114 238 174
rect 272 114 278 174
rect 232 102 278 114
rect 320 174 366 186
rect 320 114 326 174
rect 360 114 366 174
rect 320 102 366 114
rect 88 44 510 50
rect 88 6 166 44
rect 204 6 242 44
rect 280 6 318 44
rect 356 6 394 44
rect 432 6 510 44
rect 88 0 510 6
use hgu_inverter  hgu_inverter_0
timestamp 1697875053
transform 1 0 -320 0 1 -160
box 320 160 742 825
use hgu_inverter  hgu_inverter_1
timestamp 1697875053
transform -1 0 1006 0 1 -160
box 320 160 742 825
use hgu_inverter  hgu_inverter_2
timestamp 1697875053
transform 1 0 -144 0 1 -160
box 320 160 742 825
<< labels >>
flabel metal1 470 4 496 46 0 FreeSans 160 180 0 0 VSS
port 11 nsew
flabel poly 336 213 358 269 0 FreeSans 160 180 0 0 IN
port 4 nsew
flabel locali 244 228 264 264 0 FreeSans 160 180 0 0 OUT
port 15 nsew
flabel metal1 374 529 401 544 0 FreeSans 160 180 0 0 VREF
port 19 nsew
flabel metal1 464 589 500 616 0 FreeSans 160 180 0 0 VDD
port 17 nsew
<< end >>
