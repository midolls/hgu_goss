magic
tech sky130A
magscale 1 2
timestamp 1698913229
<< nwell >>
rect -38 1236 590 1250
rect -38 1058 592 1236
rect -38 861 590 1058
<< pwell >>
rect 42 621 228 803
rect 318 621 504 803
rect 42 617 63 621
rect 318 617 339 621
rect 29 583 63 617
rect 305 583 339 617
<< scnmos >>
rect 120 647 150 777
rect 396 647 426 777
<< scpmoshvt >>
rect 120 897 150 1097
rect 396 897 426 1097
<< ndiff >>
rect 68 765 120 777
rect 68 731 76 765
rect 110 731 120 765
rect 68 697 120 731
rect 68 663 76 697
rect 110 663 120 697
rect 68 647 120 663
rect 150 765 202 777
rect 150 731 160 765
rect 194 731 202 765
rect 150 697 202 731
rect 150 663 160 697
rect 194 663 202 697
rect 150 647 202 663
rect 344 765 396 777
rect 344 731 352 765
rect 386 731 396 765
rect 344 697 396 731
rect 344 663 352 697
rect 386 663 396 697
rect 344 647 396 663
rect 426 765 478 777
rect 426 731 436 765
rect 470 731 478 765
rect 426 697 478 731
rect 426 663 436 697
rect 470 663 478 697
rect 426 647 478 663
<< pdiff >>
rect 68 1085 120 1097
rect 68 1051 76 1085
rect 110 1051 120 1085
rect 68 1017 120 1051
rect 68 983 76 1017
rect 110 983 120 1017
rect 68 949 120 983
rect 68 915 76 949
rect 110 915 120 949
rect 68 897 120 915
rect 150 1085 202 1097
rect 150 1051 160 1085
rect 194 1051 202 1085
rect 150 1017 202 1051
rect 150 983 160 1017
rect 194 983 202 1017
rect 150 949 202 983
rect 150 915 160 949
rect 194 915 202 949
rect 150 897 202 915
rect 344 1085 396 1097
rect 344 1051 352 1085
rect 386 1051 396 1085
rect 344 1017 396 1051
rect 344 983 352 1017
rect 386 983 396 1017
rect 344 949 396 983
rect 344 915 352 949
rect 386 915 396 949
rect 344 897 396 915
rect 426 1085 478 1097
rect 426 1051 436 1085
rect 470 1051 478 1085
rect 426 1017 478 1051
rect 426 983 436 1017
rect 470 983 478 1017
rect 426 949 478 983
rect 426 915 436 949
rect 470 915 478 949
rect 426 897 478 915
<< ndiffc >>
rect 76 731 110 765
rect 76 663 110 697
rect 160 731 194 765
rect 160 663 194 697
rect 352 731 386 765
rect 352 663 386 697
rect 436 731 470 765
rect 436 663 470 697
<< pdiffc >>
rect 76 1051 110 1085
rect 76 983 110 1017
rect 76 915 110 949
rect 160 1051 194 1085
rect 160 983 194 1017
rect 160 915 194 949
rect 352 1051 386 1085
rect 352 983 386 1017
rect 352 915 386 949
rect 436 1051 470 1085
rect 436 983 470 1017
rect 436 915 470 949
<< psubdiff >>
rect 2 586 554 590
rect 2 552 156 586
rect 190 552 554 586
<< nsubdiff >>
rect 0 1188 552 1190
rect 0 1154 122 1188
rect 156 1154 552 1188
rect 0 1152 552 1154
<< psubdiffcont >>
rect 156 552 190 586
<< nsubdiffcont >>
rect 122 1154 156 1188
<< poly >>
rect 120 1097 150 1123
rect 396 1097 426 1123
rect 120 865 150 897
rect 396 865 426 897
rect 64 849 150 865
rect 64 815 80 849
rect 114 815 150 849
rect 64 799 150 815
rect 340 849 426 865
rect 340 815 356 849
rect 390 815 426 849
rect 340 799 426 815
rect 120 777 150 799
rect 396 777 426 799
rect 120 621 150 647
rect 396 621 426 647
<< polycont >>
rect 80 815 114 849
rect 356 815 390 849
<< locali >>
rect 106 1188 172 1190
rect 106 1161 122 1188
rect 156 1161 172 1188
rect 0 1127 29 1161
rect 63 1127 121 1161
rect 156 1154 213 1161
rect 155 1127 213 1154
rect 247 1127 305 1161
rect 339 1127 397 1161
rect 431 1127 489 1161
rect 523 1127 552 1161
rect 68 1085 110 1127
rect 68 1051 76 1085
rect 68 1017 110 1051
rect 68 983 76 1017
rect 68 949 110 983
rect 68 915 76 949
rect 68 899 110 915
rect 144 1085 210 1093
rect 144 1051 160 1085
rect 194 1051 210 1085
rect 144 1017 210 1051
rect 144 983 160 1017
rect 194 983 210 1017
rect 144 949 210 983
rect 144 915 160 949
rect 194 915 210 949
rect 144 897 210 915
rect 344 1085 386 1127
rect 344 1051 352 1085
rect 344 1017 386 1051
rect 344 983 352 1017
rect 344 949 386 983
rect 344 915 352 949
rect 344 899 386 915
rect 420 1085 486 1093
rect 420 1051 436 1085
rect 470 1051 486 1085
rect 420 1017 486 1051
rect 420 983 436 1017
rect 470 983 486 1017
rect 420 949 486 983
rect 420 915 436 949
rect 470 915 486 949
rect 420 897 486 915
rect 64 852 130 863
rect 64 818 74 852
rect 108 849 130 852
rect 64 815 80 818
rect 114 815 130 849
rect 164 854 210 897
rect 340 854 406 863
rect 164 849 406 854
rect 164 820 356 849
rect 64 765 110 781
rect 164 777 210 820
rect 340 815 356 820
rect 390 815 406 849
rect 440 858 486 897
rect 440 824 450 858
rect 484 824 486 858
rect 64 731 76 765
rect 64 697 110 731
rect 64 663 76 697
rect 64 617 110 663
rect 144 765 210 777
rect 144 731 160 765
rect 194 731 210 765
rect 144 697 210 731
rect 144 663 160 697
rect 194 663 210 697
rect 144 651 210 663
rect 340 765 386 781
rect 440 777 486 824
rect 340 731 352 765
rect 340 697 386 731
rect 340 663 352 697
rect 340 617 386 663
rect 420 765 486 777
rect 420 731 436 765
rect 470 731 486 765
rect 420 697 486 731
rect 420 663 436 697
rect 470 663 486 697
rect 420 651 486 663
rect 0 583 29 617
rect 63 583 121 617
rect 155 586 213 617
rect 155 583 156 586
rect 138 552 156 583
rect 190 583 213 586
rect 247 583 305 617
rect 339 583 397 617
rect 431 583 489 617
rect 523 583 552 617
rect 190 552 206 583
<< viali >>
rect 29 1127 63 1161
rect 121 1154 122 1161
rect 122 1154 155 1161
rect 121 1127 155 1154
rect 213 1127 247 1161
rect 305 1127 339 1161
rect 397 1127 431 1161
rect 489 1127 523 1161
rect 74 849 108 852
rect 74 818 80 849
rect 80 818 108 849
rect 450 824 484 858
rect 29 583 63 617
rect 121 583 155 617
rect 213 583 247 617
rect 305 583 339 617
rect 397 583 431 617
rect 489 583 523 617
<< metal1 >>
rect 0 1192 550 1206
rect 0 1161 552 1192
rect 0 1127 29 1161
rect 63 1127 121 1161
rect 155 1127 213 1161
rect 247 1127 305 1161
rect 339 1127 397 1161
rect 431 1127 489 1161
rect 523 1127 552 1161
rect 0 1096 552 1127
rect 438 858 608 866
rect -54 852 124 858
rect -54 818 74 852
rect 108 818 124 852
rect -54 810 124 818
rect 438 824 450 858
rect 484 824 608 858
rect 438 816 608 824
rect -54 808 106 810
rect 0 617 552 648
rect 0 583 29 617
rect 63 583 121 617
rect 155 583 213 617
rect 247 583 305 617
rect 339 583 397 617
rect 431 583 489 617
rect 523 583 552 617
rect 0 552 552 583
rect 0 530 550 552
<< labels >>
flabel metal1 0 1108 550 1206 0 FreeSans 320 0 0 0 VDD
port 0 nsew
flabel metal1 0 530 550 628 0 FreeSans 320 0 0 0 VSS
port 1 nsew
flabel metal1 -54 808 106 858 0 FreeSans 320 0 0 0 in
port 2 nsew
flabel metal1 448 816 608 866 0 FreeSans 320 0 0 0 out
port 4 nsew
flabel locali 440 889 474 923 0 FreeSans 340 0 0 0 x2.Y
flabel locali 440 821 474 855 0 FreeSans 340 0 0 0 x2.Y
flabel locali 348 821 382 855 0 FreeSans 340 0 0 0 x2.A
flabel metal1 305 583 339 617 0 FreeSans 200 0 0 0 x2.VGND
flabel metal1 305 1127 339 1161 0 FreeSans 200 0 0 0 x2.VPWR
rlabel comment 276 600 276 600 4 x2.inv_1
rlabel metal1 276 552 552 648 1 x2.VGND
rlabel metal1 276 1096 552 1192 1 x2.VPWR
flabel pwell 305 583 339 617 0 FreeSans 200 0 0 0 x2.VNB
flabel nwell 305 1127 339 1161 0 FreeSans 200 0 0 0 x2.VPB
flabel locali 164 889 198 923 0 FreeSans 340 0 0 0 x1.Y
flabel locali 164 821 198 855 0 FreeSans 340 0 0 0 x1.Y
flabel locali 72 821 106 855 0 FreeSans 340 0 0 0 x1.A
flabel metal1 29 583 63 617 0 FreeSans 200 0 0 0 x1.VGND
flabel metal1 29 1127 63 1161 0 FreeSans 200 0 0 0 x1.VPWR
rlabel comment 0 600 0 600 4 x1.inv_1
rlabel metal1 0 552 276 648 1 x1.VGND
rlabel metal1 0 1096 276 1192 1 x1.VPWR
flabel pwell 29 583 63 617 0 FreeSans 200 0 0 0 x1.VNB
flabel nwell 29 1127 63 1161 0 FreeSans 200 0 0 0 x1.VPB
<< end >>
