magic
tech sky130A
magscale 1 2
timestamp 1701888524
<< nwell >>
rect -400 5384 -72 6034
rect 400 5768 856 6034
rect 1280 5768 1992 6034
rect 2899 5768 4123 6034
rect 400 5650 984 5768
rect 1280 5650 2504 5768
rect 2899 5650 4635 5768
rect 5392 5650 7640 6034
rect 528 5384 984 5650
rect 1792 5384 2504 5650
rect 3411 5384 4635 5650
rect 7976 5384 10224 5768
rect 10479 5650 14775 6034
rect 15740 5384 20036 5768
rect 20316 5650 28708 6034
rect 29284 5384 37676 5768
<< pwell >>
rect 17436 3572 17468 3622
rect 17436 439 17468 489
<< pmoslvt >>
rect -271 5828 -201 5996
rect 529 5828 599 5996
rect 657 5828 727 5996
rect 1409 5828 1479 5996
rect 1537 5828 1607 5996
rect 1665 5828 1735 5996
rect 1793 5828 1863 5996
rect 3028 5828 3098 5996
rect 3156 5828 3226 5996
rect 3284 5828 3354 5996
rect 3412 5828 3482 5996
rect 3540 5828 3610 5996
rect 3668 5828 3738 5996
rect 3796 5828 3866 5996
rect 3924 5828 3994 5996
rect 5521 5828 5591 5996
rect 5649 5828 5719 5996
rect 5777 5828 5847 5996
rect 5905 5828 5975 5996
rect 6033 5828 6103 5996
rect 6161 5828 6231 5996
rect 6289 5828 6359 5996
rect 6417 5828 6487 5996
rect 6545 5828 6615 5996
rect 6673 5828 6743 5996
rect 6801 5828 6871 5996
rect 6929 5828 6999 5996
rect 7057 5828 7127 5996
rect 7185 5828 7255 5996
rect 7313 5828 7383 5996
rect 7441 5828 7511 5996
rect 10608 5828 10678 5996
rect 10736 5828 10806 5996
rect 10864 5828 10934 5996
rect 10992 5828 11062 5996
rect 11120 5828 11190 5996
rect 11248 5828 11318 5996
rect 11376 5828 11446 5996
rect 11504 5828 11574 5996
rect 11632 5828 11702 5996
rect 11760 5828 11830 5996
rect 11888 5828 11958 5996
rect 12016 5828 12086 5996
rect 12144 5828 12214 5996
rect 12272 5828 12342 5996
rect 12400 5828 12470 5996
rect 12528 5828 12598 5996
rect 12656 5828 12726 5996
rect 12784 5828 12854 5996
rect 12912 5828 12982 5996
rect 13040 5828 13110 5996
rect 13168 5828 13238 5996
rect 13296 5828 13366 5996
rect 13424 5828 13494 5996
rect 13552 5828 13622 5996
rect 13680 5828 13750 5996
rect 13808 5828 13878 5996
rect 13936 5828 14006 5996
rect 14064 5828 14134 5996
rect 14192 5828 14262 5996
rect 14320 5828 14390 5996
rect 14448 5828 14518 5996
rect 14576 5828 14646 5996
rect 20445 5828 20515 5996
rect 20573 5828 20643 5996
rect 20701 5828 20771 5996
rect 20829 5828 20899 5996
rect 20957 5828 21027 5996
rect 21085 5828 21155 5996
rect 21213 5828 21283 5996
rect 21341 5828 21411 5996
rect 21469 5828 21539 5996
rect 21597 5828 21667 5996
rect 21725 5828 21795 5996
rect 21853 5828 21923 5996
rect 21981 5828 22051 5996
rect 22109 5828 22179 5996
rect 22237 5828 22307 5996
rect 22365 5828 22435 5996
rect 22493 5828 22563 5996
rect 22621 5828 22691 5996
rect 22749 5828 22819 5996
rect 22877 5828 22947 5996
rect 23005 5828 23075 5996
rect 23133 5828 23203 5996
rect 23261 5828 23331 5996
rect 23389 5828 23459 5996
rect 23517 5828 23587 5996
rect 23645 5828 23715 5996
rect 23773 5828 23843 5996
rect 23901 5828 23971 5996
rect 24029 5828 24099 5996
rect 24157 5828 24227 5996
rect 24285 5828 24355 5996
rect 24413 5828 24483 5996
rect 24541 5828 24611 5996
rect 24669 5828 24739 5996
rect 24797 5828 24867 5996
rect 24925 5828 24995 5996
rect 25053 5828 25123 5996
rect 25181 5828 25251 5996
rect 25309 5828 25379 5996
rect 25437 5828 25507 5996
rect 25565 5828 25635 5996
rect 25693 5828 25763 5996
rect 25821 5828 25891 5996
rect 25949 5828 26019 5996
rect 26077 5828 26147 5996
rect 26205 5828 26275 5996
rect 26333 5828 26403 5996
rect 26461 5828 26531 5996
rect 26589 5828 26659 5996
rect 26717 5828 26787 5996
rect 26845 5828 26915 5996
rect 26973 5828 27043 5996
rect 27101 5828 27171 5996
rect 27229 5828 27299 5996
rect 27357 5828 27427 5996
rect 27485 5828 27555 5996
rect 27613 5828 27683 5996
rect 27741 5828 27811 5996
rect 27869 5828 27939 5996
rect 27997 5828 28067 5996
rect 28125 5828 28195 5996
rect 28253 5828 28323 5996
rect 28381 5828 28451 5996
rect 28509 5828 28579 5996
rect -271 5422 -201 5590
rect 657 5422 727 5590
rect 785 5422 855 5590
rect 1921 5422 1991 5590
rect 2049 5422 2119 5590
rect 2177 5422 2247 5590
rect 2305 5422 2375 5590
rect 3540 5422 3610 5590
rect 3668 5422 3738 5590
rect 3796 5422 3866 5590
rect 3924 5422 3994 5590
rect 4052 5422 4122 5590
rect 4180 5422 4250 5590
rect 4308 5422 4378 5590
rect 4436 5422 4506 5590
rect 8105 5422 8175 5590
rect 8233 5422 8303 5590
rect 8361 5422 8431 5590
rect 8489 5422 8559 5590
rect 8617 5422 8687 5590
rect 8745 5422 8815 5590
rect 8873 5422 8943 5590
rect 9001 5422 9071 5590
rect 9129 5422 9199 5590
rect 9257 5422 9327 5590
rect 9385 5422 9455 5590
rect 9513 5422 9583 5590
rect 9641 5422 9711 5590
rect 9769 5422 9839 5590
rect 9897 5422 9967 5590
rect 10025 5422 10095 5590
rect 15869 5422 15939 5590
rect 15997 5422 16067 5590
rect 16125 5422 16195 5590
rect 16253 5422 16323 5590
rect 16381 5422 16451 5590
rect 16509 5422 16579 5590
rect 16637 5422 16707 5590
rect 16765 5422 16835 5590
rect 16893 5422 16963 5590
rect 17021 5422 17091 5590
rect 17149 5422 17219 5590
rect 17277 5422 17347 5590
rect 17405 5422 17475 5590
rect 17533 5422 17603 5590
rect 17661 5422 17731 5590
rect 17789 5422 17859 5590
rect 17917 5422 17987 5590
rect 18045 5422 18115 5590
rect 18173 5422 18243 5590
rect 18301 5422 18371 5590
rect 18429 5422 18499 5590
rect 18557 5422 18627 5590
rect 18685 5422 18755 5590
rect 18813 5422 18883 5590
rect 18941 5422 19011 5590
rect 19069 5422 19139 5590
rect 19197 5422 19267 5590
rect 19325 5422 19395 5590
rect 19453 5422 19523 5590
rect 19581 5422 19651 5590
rect 19709 5422 19779 5590
rect 19837 5422 19907 5590
rect 29413 5422 29483 5590
rect 29541 5422 29611 5590
rect 29669 5422 29739 5590
rect 29797 5422 29867 5590
rect 29925 5422 29995 5590
rect 30053 5422 30123 5590
rect 30181 5422 30251 5590
rect 30309 5422 30379 5590
rect 30437 5422 30507 5590
rect 30565 5422 30635 5590
rect 30693 5422 30763 5590
rect 30821 5422 30891 5590
rect 30949 5422 31019 5590
rect 31077 5422 31147 5590
rect 31205 5422 31275 5590
rect 31333 5422 31403 5590
rect 31461 5422 31531 5590
rect 31589 5422 31659 5590
rect 31717 5422 31787 5590
rect 31845 5422 31915 5590
rect 31973 5422 32043 5590
rect 32101 5422 32171 5590
rect 32229 5422 32299 5590
rect 32357 5422 32427 5590
rect 32485 5422 32555 5590
rect 32613 5422 32683 5590
rect 32741 5422 32811 5590
rect 32869 5422 32939 5590
rect 32997 5422 33067 5590
rect 33125 5422 33195 5590
rect 33253 5422 33323 5590
rect 33381 5422 33451 5590
rect 33509 5422 33579 5590
rect 33637 5422 33707 5590
rect 33765 5422 33835 5590
rect 33893 5422 33963 5590
rect 34021 5422 34091 5590
rect 34149 5422 34219 5590
rect 34277 5422 34347 5590
rect 34405 5422 34475 5590
rect 34533 5422 34603 5590
rect 34661 5422 34731 5590
rect 34789 5422 34859 5590
rect 34917 5422 34987 5590
rect 35045 5422 35115 5590
rect 35173 5422 35243 5590
rect 35301 5422 35371 5590
rect 35429 5422 35499 5590
rect 35557 5422 35627 5590
rect 35685 5422 35755 5590
rect 35813 5422 35883 5590
rect 35941 5422 36011 5590
rect 36069 5422 36139 5590
rect 36197 5422 36267 5590
rect 36325 5422 36395 5590
rect 36453 5422 36523 5590
rect 36581 5422 36651 5590
rect 36709 5422 36779 5590
rect 36837 5422 36907 5590
rect 36965 5422 37035 5590
rect 37093 5422 37163 5590
rect 37221 5422 37291 5590
rect 37349 5422 37419 5590
rect 37477 5422 37547 5590
<< nmoslvt >>
rect -271 6128 -201 6212
rect 529 6128 599 6212
rect 657 6128 727 6212
rect 1409 6128 1479 6212
rect 1537 6128 1607 6212
rect 1665 6128 1735 6212
rect 1793 6128 1863 6212
rect 3028 6128 3098 6212
rect 3156 6128 3226 6212
rect 3284 6128 3354 6212
rect 3412 6128 3482 6212
rect 3540 6128 3610 6212
rect 3668 6128 3738 6212
rect 3796 6128 3866 6212
rect 3924 6128 3994 6212
rect 5521 6128 5591 6212
rect 5649 6128 5719 6212
rect 5777 6128 5847 6212
rect 5905 6128 5975 6212
rect 6033 6128 6103 6212
rect 6161 6128 6231 6212
rect 6289 6128 6359 6212
rect 6417 6128 6487 6212
rect 6545 6128 6615 6212
rect 6673 6128 6743 6212
rect 6801 6128 6871 6212
rect 6929 6128 6999 6212
rect 7057 6128 7127 6212
rect 7185 6128 7255 6212
rect 7313 6128 7383 6212
rect 7441 6128 7511 6212
rect 10608 6128 10678 6212
rect 10736 6128 10806 6212
rect 10864 6128 10934 6212
rect 10992 6128 11062 6212
rect 11120 6128 11190 6212
rect 11248 6128 11318 6212
rect 11376 6128 11446 6212
rect 11504 6128 11574 6212
rect 11632 6128 11702 6212
rect 11760 6128 11830 6212
rect 11888 6128 11958 6212
rect 12016 6128 12086 6212
rect 12144 6128 12214 6212
rect 12272 6128 12342 6212
rect 12400 6128 12470 6212
rect 12528 6128 12598 6212
rect 12656 6128 12726 6212
rect 12784 6128 12854 6212
rect 12912 6128 12982 6212
rect 13040 6128 13110 6212
rect 13168 6128 13238 6212
rect 13296 6128 13366 6212
rect 13424 6128 13494 6212
rect 13552 6128 13622 6212
rect 13680 6128 13750 6212
rect 13808 6128 13878 6212
rect 13936 6128 14006 6212
rect 14064 6128 14134 6212
rect 14192 6128 14262 6212
rect 14320 6128 14390 6212
rect 14448 6128 14518 6212
rect 14576 6128 14646 6212
rect 20445 6128 20515 6212
rect 20573 6128 20643 6212
rect 20701 6128 20771 6212
rect 20829 6128 20899 6212
rect 20957 6128 21027 6212
rect 21085 6128 21155 6212
rect 21213 6128 21283 6212
rect 21341 6128 21411 6212
rect 21469 6128 21539 6212
rect 21597 6128 21667 6212
rect 21725 6128 21795 6212
rect 21853 6128 21923 6212
rect 21981 6128 22051 6212
rect 22109 6128 22179 6212
rect 22237 6128 22307 6212
rect 22365 6128 22435 6212
rect 22493 6128 22563 6212
rect 22621 6128 22691 6212
rect 22749 6128 22819 6212
rect 22877 6128 22947 6212
rect 23005 6128 23075 6212
rect 23133 6128 23203 6212
rect 23261 6128 23331 6212
rect 23389 6128 23459 6212
rect 23517 6128 23587 6212
rect 23645 6128 23715 6212
rect 23773 6128 23843 6212
rect 23901 6128 23971 6212
rect 24029 6128 24099 6212
rect 24157 6128 24227 6212
rect 24285 6128 24355 6212
rect 24413 6128 24483 6212
rect 24541 6128 24611 6212
rect 24669 6128 24739 6212
rect 24797 6128 24867 6212
rect 24925 6128 24995 6212
rect 25053 6128 25123 6212
rect 25181 6128 25251 6212
rect 25309 6128 25379 6212
rect 25437 6128 25507 6212
rect 25565 6128 25635 6212
rect 25693 6128 25763 6212
rect 25821 6128 25891 6212
rect 25949 6128 26019 6212
rect 26077 6128 26147 6212
rect 26205 6128 26275 6212
rect 26333 6128 26403 6212
rect 26461 6128 26531 6212
rect 26589 6128 26659 6212
rect 26717 6128 26787 6212
rect 26845 6128 26915 6212
rect 26973 6128 27043 6212
rect 27101 6128 27171 6212
rect 27229 6128 27299 6212
rect 27357 6128 27427 6212
rect 27485 6128 27555 6212
rect 27613 6128 27683 6212
rect 27741 6128 27811 6212
rect 27869 6128 27939 6212
rect 27997 6128 28067 6212
rect 28125 6128 28195 6212
rect 28253 6128 28323 6212
rect 28381 6128 28451 6212
rect 28509 6128 28579 6212
rect -271 5206 -201 5290
rect 657 5206 727 5290
rect 785 5206 855 5290
rect 1921 5206 1991 5290
rect 2049 5206 2119 5290
rect 2177 5206 2247 5290
rect 2305 5206 2375 5290
rect 3540 5206 3610 5290
rect 3668 5206 3738 5290
rect 3796 5206 3866 5290
rect 3924 5206 3994 5290
rect 4052 5206 4122 5290
rect 4180 5206 4250 5290
rect 4308 5206 4378 5290
rect 4436 5206 4506 5290
rect 8105 5206 8175 5290
rect 8233 5206 8303 5290
rect 8361 5206 8431 5290
rect 8489 5206 8559 5290
rect 8617 5206 8687 5290
rect 8745 5206 8815 5290
rect 8873 5206 8943 5290
rect 9001 5206 9071 5290
rect 9129 5206 9199 5290
rect 9257 5206 9327 5290
rect 9385 5206 9455 5290
rect 9513 5206 9583 5290
rect 9641 5206 9711 5290
rect 9769 5206 9839 5290
rect 9897 5206 9967 5290
rect 10025 5206 10095 5290
rect 15869 5206 15939 5290
rect 15997 5206 16067 5290
rect 16125 5206 16195 5290
rect 16253 5206 16323 5290
rect 16381 5206 16451 5290
rect 16509 5206 16579 5290
rect 16637 5206 16707 5290
rect 16765 5206 16835 5290
rect 16893 5206 16963 5290
rect 17021 5206 17091 5290
rect 17149 5206 17219 5290
rect 17277 5206 17347 5290
rect 17405 5206 17475 5290
rect 17533 5206 17603 5290
rect 17661 5206 17731 5290
rect 17789 5206 17859 5290
rect 17917 5206 17987 5290
rect 18045 5206 18115 5290
rect 18173 5206 18243 5290
rect 18301 5206 18371 5290
rect 18429 5206 18499 5290
rect 18557 5206 18627 5290
rect 18685 5206 18755 5290
rect 18813 5206 18883 5290
rect 18941 5206 19011 5290
rect 19069 5206 19139 5290
rect 19197 5206 19267 5290
rect 19325 5206 19395 5290
rect 19453 5206 19523 5290
rect 19581 5206 19651 5290
rect 19709 5206 19779 5290
rect 19837 5206 19907 5290
rect 29413 5206 29483 5290
rect 29541 5206 29611 5290
rect 29669 5206 29739 5290
rect 29797 5206 29867 5290
rect 29925 5206 29995 5290
rect 30053 5206 30123 5290
rect 30181 5206 30251 5290
rect 30309 5206 30379 5290
rect 30437 5206 30507 5290
rect 30565 5206 30635 5290
rect 30693 5206 30763 5290
rect 30821 5206 30891 5290
rect 30949 5206 31019 5290
rect 31077 5206 31147 5290
rect 31205 5206 31275 5290
rect 31333 5206 31403 5290
rect 31461 5206 31531 5290
rect 31589 5206 31659 5290
rect 31717 5206 31787 5290
rect 31845 5206 31915 5290
rect 31973 5206 32043 5290
rect 32101 5206 32171 5290
rect 32229 5206 32299 5290
rect 32357 5206 32427 5290
rect 32485 5206 32555 5290
rect 32613 5206 32683 5290
rect 32741 5206 32811 5290
rect 32869 5206 32939 5290
rect 32997 5206 33067 5290
rect 33125 5206 33195 5290
rect 33253 5206 33323 5290
rect 33381 5206 33451 5290
rect 33509 5206 33579 5290
rect 33637 5206 33707 5290
rect 33765 5206 33835 5290
rect 33893 5206 33963 5290
rect 34021 5206 34091 5290
rect 34149 5206 34219 5290
rect 34277 5206 34347 5290
rect 34405 5206 34475 5290
rect 34533 5206 34603 5290
rect 34661 5206 34731 5290
rect 34789 5206 34859 5290
rect 34917 5206 34987 5290
rect 35045 5206 35115 5290
rect 35173 5206 35243 5290
rect 35301 5206 35371 5290
rect 35429 5206 35499 5290
rect 35557 5206 35627 5290
rect 35685 5206 35755 5290
rect 35813 5206 35883 5290
rect 35941 5206 36011 5290
rect 36069 5206 36139 5290
rect 36197 5206 36267 5290
rect 36325 5206 36395 5290
rect 36453 5206 36523 5290
rect 36581 5206 36651 5290
rect 36709 5206 36779 5290
rect 36837 5206 36907 5290
rect 36965 5206 37035 5290
rect 37093 5206 37163 5290
rect 37221 5206 37291 5290
rect 37349 5206 37419 5290
rect 37477 5206 37547 5290
<< ndiff >>
rect -329 6200 -271 6212
rect -329 6140 -317 6200
rect -283 6140 -271 6200
rect -329 6128 -271 6140
rect -201 6200 -143 6212
rect -201 6140 -189 6200
rect -155 6140 -143 6200
rect -201 6128 -143 6140
rect 471 6200 529 6212
rect 471 6140 483 6200
rect 517 6140 529 6200
rect 471 6128 529 6140
rect 599 6200 657 6212
rect 599 6140 611 6200
rect 645 6140 657 6200
rect 599 6128 657 6140
rect 727 6200 785 6212
rect 727 6140 739 6200
rect 773 6140 785 6200
rect 727 6128 785 6140
rect 1351 6200 1409 6212
rect 1351 6140 1363 6200
rect 1397 6140 1409 6200
rect 1351 6128 1409 6140
rect 1479 6200 1537 6212
rect 1479 6140 1491 6200
rect 1525 6140 1537 6200
rect 1479 6128 1537 6140
rect 1607 6200 1665 6212
rect 1607 6140 1619 6200
rect 1653 6140 1665 6200
rect 1607 6128 1665 6140
rect 1735 6200 1793 6212
rect 1735 6140 1747 6200
rect 1781 6140 1793 6200
rect 1735 6128 1793 6140
rect 1863 6200 1921 6212
rect 1863 6140 1875 6200
rect 1909 6140 1921 6200
rect 1863 6128 1921 6140
rect 2970 6200 3028 6212
rect 2970 6140 2982 6200
rect 3016 6140 3028 6200
rect 2970 6128 3028 6140
rect 3098 6200 3156 6212
rect 3098 6140 3110 6200
rect 3144 6140 3156 6200
rect 3098 6128 3156 6140
rect 3226 6200 3284 6212
rect 3226 6140 3238 6200
rect 3272 6140 3284 6200
rect 3226 6128 3284 6140
rect 3354 6200 3412 6212
rect 3354 6140 3366 6200
rect 3400 6140 3412 6200
rect 3354 6128 3412 6140
rect 3482 6200 3540 6212
rect 3482 6140 3494 6200
rect 3528 6140 3540 6200
rect 3482 6128 3540 6140
rect 3610 6200 3668 6212
rect 3610 6140 3622 6200
rect 3656 6140 3668 6200
rect 3610 6128 3668 6140
rect 3738 6200 3796 6212
rect 3738 6140 3750 6200
rect 3784 6140 3796 6200
rect 3738 6128 3796 6140
rect 3866 6200 3924 6212
rect 3866 6140 3878 6200
rect 3912 6140 3924 6200
rect 3866 6128 3924 6140
rect 3994 6200 4052 6212
rect 3994 6140 4006 6200
rect 4040 6140 4052 6200
rect 5463 6200 5521 6212
rect 3994 6128 4052 6140
rect 5463 6140 5475 6200
rect 5509 6140 5521 6200
rect 5463 6128 5521 6140
rect 5591 6200 5649 6212
rect 5591 6140 5603 6200
rect 5637 6140 5649 6200
rect 5591 6128 5649 6140
rect 5719 6200 5777 6212
rect 5719 6140 5731 6200
rect 5765 6140 5777 6200
rect 5719 6128 5777 6140
rect 5847 6200 5905 6212
rect 5847 6140 5859 6200
rect 5893 6140 5905 6200
rect 5847 6128 5905 6140
rect 5975 6200 6033 6212
rect 5975 6140 5987 6200
rect 6021 6140 6033 6200
rect 5975 6128 6033 6140
rect 6103 6200 6161 6212
rect 6103 6140 6115 6200
rect 6149 6140 6161 6200
rect 6103 6128 6161 6140
rect 6231 6200 6289 6212
rect 6231 6140 6243 6200
rect 6277 6140 6289 6200
rect 6231 6128 6289 6140
rect 6359 6200 6417 6212
rect 6359 6140 6371 6200
rect 6405 6140 6417 6200
rect 6359 6128 6417 6140
rect 6487 6200 6545 6212
rect 6487 6140 6499 6200
rect 6533 6140 6545 6200
rect 6487 6128 6545 6140
rect 6615 6200 6673 6212
rect 6615 6140 6627 6200
rect 6661 6140 6673 6200
rect 6615 6128 6673 6140
rect 6743 6200 6801 6212
rect 6743 6140 6755 6200
rect 6789 6140 6801 6200
rect 6743 6128 6801 6140
rect 6871 6200 6929 6212
rect 6871 6140 6883 6200
rect 6917 6140 6929 6200
rect 6871 6128 6929 6140
rect 6999 6200 7057 6212
rect 6999 6140 7011 6200
rect 7045 6140 7057 6200
rect 6999 6128 7057 6140
rect 7127 6200 7185 6212
rect 7127 6140 7139 6200
rect 7173 6140 7185 6200
rect 7127 6128 7185 6140
rect 7255 6200 7313 6212
rect 7255 6140 7267 6200
rect 7301 6140 7313 6200
rect 7255 6128 7313 6140
rect 7383 6200 7441 6212
rect 7383 6140 7395 6200
rect 7429 6140 7441 6200
rect 7383 6128 7441 6140
rect 7511 6200 7569 6212
rect 7511 6140 7523 6200
rect 7557 6140 7569 6200
rect 10550 6200 10608 6212
rect 7511 6128 7569 6140
rect 10550 6140 10562 6200
rect 10596 6140 10608 6200
rect 10550 6128 10608 6140
rect 10678 6200 10736 6212
rect 10678 6140 10690 6200
rect 10724 6140 10736 6200
rect 10678 6128 10736 6140
rect 10806 6200 10864 6212
rect 10806 6140 10818 6200
rect 10852 6140 10864 6200
rect 10806 6128 10864 6140
rect 10934 6200 10992 6212
rect 10934 6140 10946 6200
rect 10980 6140 10992 6200
rect 10934 6128 10992 6140
rect 11062 6200 11120 6212
rect 11062 6140 11074 6200
rect 11108 6140 11120 6200
rect 11062 6128 11120 6140
rect 11190 6200 11248 6212
rect 11190 6140 11202 6200
rect 11236 6140 11248 6200
rect 11190 6128 11248 6140
rect 11318 6200 11376 6212
rect 11318 6140 11330 6200
rect 11364 6140 11376 6200
rect 11318 6128 11376 6140
rect 11446 6200 11504 6212
rect 11446 6140 11458 6200
rect 11492 6140 11504 6200
rect 11446 6128 11504 6140
rect 11574 6200 11632 6212
rect 11574 6140 11586 6200
rect 11620 6140 11632 6200
rect 11574 6128 11632 6140
rect 11702 6200 11760 6212
rect 11702 6140 11714 6200
rect 11748 6140 11760 6200
rect 11702 6128 11760 6140
rect 11830 6200 11888 6212
rect 11830 6140 11842 6200
rect 11876 6140 11888 6200
rect 11830 6128 11888 6140
rect 11958 6200 12016 6212
rect 11958 6140 11970 6200
rect 12004 6140 12016 6200
rect 11958 6128 12016 6140
rect 12086 6200 12144 6212
rect 12086 6140 12098 6200
rect 12132 6140 12144 6200
rect 12086 6128 12144 6140
rect 12214 6200 12272 6212
rect 12214 6140 12226 6200
rect 12260 6140 12272 6200
rect 12214 6128 12272 6140
rect 12342 6200 12400 6212
rect 12342 6140 12354 6200
rect 12388 6140 12400 6200
rect 12342 6128 12400 6140
rect 12470 6200 12528 6212
rect 12470 6140 12482 6200
rect 12516 6140 12528 6200
rect 12470 6128 12528 6140
rect 12598 6200 12656 6212
rect 12598 6140 12610 6200
rect 12644 6140 12656 6200
rect 12598 6128 12656 6140
rect 12726 6200 12784 6212
rect 12726 6140 12738 6200
rect 12772 6140 12784 6200
rect 12726 6128 12784 6140
rect 12854 6200 12912 6212
rect 12854 6140 12866 6200
rect 12900 6140 12912 6200
rect 12854 6128 12912 6140
rect 12982 6200 13040 6212
rect 12982 6140 12994 6200
rect 13028 6140 13040 6200
rect 12982 6128 13040 6140
rect 13110 6200 13168 6212
rect 13110 6140 13122 6200
rect 13156 6140 13168 6200
rect 13110 6128 13168 6140
rect 13238 6200 13296 6212
rect 13238 6140 13250 6200
rect 13284 6140 13296 6200
rect 13238 6128 13296 6140
rect 13366 6200 13424 6212
rect 13366 6140 13378 6200
rect 13412 6140 13424 6200
rect 13366 6128 13424 6140
rect 13494 6200 13552 6212
rect 13494 6140 13506 6200
rect 13540 6140 13552 6200
rect 13494 6128 13552 6140
rect 13622 6200 13680 6212
rect 13622 6140 13634 6200
rect 13668 6140 13680 6200
rect 13622 6128 13680 6140
rect 13750 6200 13808 6212
rect 13750 6140 13762 6200
rect 13796 6140 13808 6200
rect 13750 6128 13808 6140
rect 13878 6200 13936 6212
rect 13878 6140 13890 6200
rect 13924 6140 13936 6200
rect 13878 6128 13936 6140
rect 14006 6200 14064 6212
rect 14006 6140 14018 6200
rect 14052 6140 14064 6200
rect 14006 6128 14064 6140
rect 14134 6200 14192 6212
rect 14134 6140 14146 6200
rect 14180 6140 14192 6200
rect 14134 6128 14192 6140
rect 14262 6200 14320 6212
rect 14262 6140 14274 6200
rect 14308 6140 14320 6200
rect 14262 6128 14320 6140
rect 14390 6200 14448 6212
rect 14390 6140 14402 6200
rect 14436 6140 14448 6200
rect 14390 6128 14448 6140
rect 14518 6200 14576 6212
rect 14518 6140 14530 6200
rect 14564 6140 14576 6200
rect 14518 6128 14576 6140
rect 14646 6200 14704 6212
rect 14646 6140 14658 6200
rect 14692 6140 14704 6200
rect 14646 6128 14704 6140
rect 20387 6200 20445 6212
rect 20387 6140 20399 6200
rect 20433 6140 20445 6200
rect 20387 6128 20445 6140
rect 20515 6200 20573 6212
rect 20515 6140 20527 6200
rect 20561 6140 20573 6200
rect 20515 6128 20573 6140
rect 20643 6200 20701 6212
rect 20643 6140 20655 6200
rect 20689 6140 20701 6200
rect 20643 6128 20701 6140
rect 20771 6200 20829 6212
rect 20771 6140 20783 6200
rect 20817 6140 20829 6200
rect 20771 6128 20829 6140
rect 20899 6200 20957 6212
rect 20899 6140 20911 6200
rect 20945 6140 20957 6200
rect 20899 6128 20957 6140
rect 21027 6200 21085 6212
rect 21027 6140 21039 6200
rect 21073 6140 21085 6200
rect 21027 6128 21085 6140
rect 21155 6200 21213 6212
rect 21155 6140 21167 6200
rect 21201 6140 21213 6200
rect 21155 6128 21213 6140
rect 21283 6200 21341 6212
rect 21283 6140 21295 6200
rect 21329 6140 21341 6200
rect 21283 6128 21341 6140
rect 21411 6200 21469 6212
rect 21411 6140 21423 6200
rect 21457 6140 21469 6200
rect 21411 6128 21469 6140
rect 21539 6200 21597 6212
rect 21539 6140 21551 6200
rect 21585 6140 21597 6200
rect 21539 6128 21597 6140
rect 21667 6200 21725 6212
rect 21667 6140 21679 6200
rect 21713 6140 21725 6200
rect 21667 6128 21725 6140
rect 21795 6200 21853 6212
rect 21795 6140 21807 6200
rect 21841 6140 21853 6200
rect 21795 6128 21853 6140
rect 21923 6200 21981 6212
rect 21923 6140 21935 6200
rect 21969 6140 21981 6200
rect 21923 6128 21981 6140
rect 22051 6200 22109 6212
rect 22051 6140 22063 6200
rect 22097 6140 22109 6200
rect 22051 6128 22109 6140
rect 22179 6200 22237 6212
rect 22179 6140 22191 6200
rect 22225 6140 22237 6200
rect 22179 6128 22237 6140
rect 22307 6200 22365 6212
rect 22307 6140 22319 6200
rect 22353 6140 22365 6200
rect 22307 6128 22365 6140
rect 22435 6200 22493 6212
rect 22435 6140 22447 6200
rect 22481 6140 22493 6200
rect 22435 6128 22493 6140
rect 22563 6200 22621 6212
rect 22563 6140 22575 6200
rect 22609 6140 22621 6200
rect 22563 6128 22621 6140
rect 22691 6200 22749 6212
rect 22691 6140 22703 6200
rect 22737 6140 22749 6200
rect 22691 6128 22749 6140
rect 22819 6200 22877 6212
rect 22819 6140 22831 6200
rect 22865 6140 22877 6200
rect 22819 6128 22877 6140
rect 22947 6200 23005 6212
rect 22947 6140 22959 6200
rect 22993 6140 23005 6200
rect 22947 6128 23005 6140
rect 23075 6200 23133 6212
rect 23075 6140 23087 6200
rect 23121 6140 23133 6200
rect 23075 6128 23133 6140
rect 23203 6200 23261 6212
rect 23203 6140 23215 6200
rect 23249 6140 23261 6200
rect 23203 6128 23261 6140
rect 23331 6200 23389 6212
rect 23331 6140 23343 6200
rect 23377 6140 23389 6200
rect 23331 6128 23389 6140
rect 23459 6200 23517 6212
rect 23459 6140 23471 6200
rect 23505 6140 23517 6200
rect 23459 6128 23517 6140
rect 23587 6200 23645 6212
rect 23587 6140 23599 6200
rect 23633 6140 23645 6200
rect 23587 6128 23645 6140
rect 23715 6200 23773 6212
rect 23715 6140 23727 6200
rect 23761 6140 23773 6200
rect 23715 6128 23773 6140
rect 23843 6200 23901 6212
rect 23843 6140 23855 6200
rect 23889 6140 23901 6200
rect 23843 6128 23901 6140
rect 23971 6200 24029 6212
rect 23971 6140 23983 6200
rect 24017 6140 24029 6200
rect 23971 6128 24029 6140
rect 24099 6200 24157 6212
rect 24099 6140 24111 6200
rect 24145 6140 24157 6200
rect 24099 6128 24157 6140
rect 24227 6200 24285 6212
rect 24227 6140 24239 6200
rect 24273 6140 24285 6200
rect 24227 6128 24285 6140
rect 24355 6200 24413 6212
rect 24355 6140 24367 6200
rect 24401 6140 24413 6200
rect 24355 6128 24413 6140
rect 24483 6200 24541 6212
rect 24483 6140 24495 6200
rect 24529 6140 24541 6200
rect 24483 6128 24541 6140
rect 24611 6200 24669 6212
rect 24611 6140 24623 6200
rect 24657 6140 24669 6200
rect 24611 6128 24669 6140
rect 24739 6200 24797 6212
rect 24739 6140 24751 6200
rect 24785 6140 24797 6200
rect 24739 6128 24797 6140
rect 24867 6200 24925 6212
rect 24867 6140 24879 6200
rect 24913 6140 24925 6200
rect 24867 6128 24925 6140
rect 24995 6200 25053 6212
rect 24995 6140 25007 6200
rect 25041 6140 25053 6200
rect 24995 6128 25053 6140
rect 25123 6200 25181 6212
rect 25123 6140 25135 6200
rect 25169 6140 25181 6200
rect 25123 6128 25181 6140
rect 25251 6200 25309 6212
rect 25251 6140 25263 6200
rect 25297 6140 25309 6200
rect 25251 6128 25309 6140
rect 25379 6200 25437 6212
rect 25379 6140 25391 6200
rect 25425 6140 25437 6200
rect 25379 6128 25437 6140
rect 25507 6200 25565 6212
rect 25507 6140 25519 6200
rect 25553 6140 25565 6200
rect 25507 6128 25565 6140
rect 25635 6200 25693 6212
rect 25635 6140 25647 6200
rect 25681 6140 25693 6200
rect 25635 6128 25693 6140
rect 25763 6200 25821 6212
rect 25763 6140 25775 6200
rect 25809 6140 25821 6200
rect 25763 6128 25821 6140
rect 25891 6200 25949 6212
rect 25891 6140 25903 6200
rect 25937 6140 25949 6200
rect 25891 6128 25949 6140
rect 26019 6200 26077 6212
rect 26019 6140 26031 6200
rect 26065 6140 26077 6200
rect 26019 6128 26077 6140
rect 26147 6200 26205 6212
rect 26147 6140 26159 6200
rect 26193 6140 26205 6200
rect 26147 6128 26205 6140
rect 26275 6200 26333 6212
rect 26275 6140 26287 6200
rect 26321 6140 26333 6200
rect 26275 6128 26333 6140
rect 26403 6200 26461 6212
rect 26403 6140 26415 6200
rect 26449 6140 26461 6200
rect 26403 6128 26461 6140
rect 26531 6200 26589 6212
rect 26531 6140 26543 6200
rect 26577 6140 26589 6200
rect 26531 6128 26589 6140
rect 26659 6200 26717 6212
rect 26659 6140 26671 6200
rect 26705 6140 26717 6200
rect 26659 6128 26717 6140
rect 26787 6200 26845 6212
rect 26787 6140 26799 6200
rect 26833 6140 26845 6200
rect 26787 6128 26845 6140
rect 26915 6200 26973 6212
rect 26915 6140 26927 6200
rect 26961 6140 26973 6200
rect 26915 6128 26973 6140
rect 27043 6200 27101 6212
rect 27043 6140 27055 6200
rect 27089 6140 27101 6200
rect 27043 6128 27101 6140
rect 27171 6200 27229 6212
rect 27171 6140 27183 6200
rect 27217 6140 27229 6200
rect 27171 6128 27229 6140
rect 27299 6200 27357 6212
rect 27299 6140 27311 6200
rect 27345 6140 27357 6200
rect 27299 6128 27357 6140
rect 27427 6200 27485 6212
rect 27427 6140 27439 6200
rect 27473 6140 27485 6200
rect 27427 6128 27485 6140
rect 27555 6200 27613 6212
rect 27555 6140 27567 6200
rect 27601 6140 27613 6200
rect 27555 6128 27613 6140
rect 27683 6200 27741 6212
rect 27683 6140 27695 6200
rect 27729 6140 27741 6200
rect 27683 6128 27741 6140
rect 27811 6200 27869 6212
rect 27811 6140 27823 6200
rect 27857 6140 27869 6200
rect 27811 6128 27869 6140
rect 27939 6200 27997 6212
rect 27939 6140 27951 6200
rect 27985 6140 27997 6200
rect 27939 6128 27997 6140
rect 28067 6200 28125 6212
rect 28067 6140 28079 6200
rect 28113 6140 28125 6200
rect 28067 6128 28125 6140
rect 28195 6200 28253 6212
rect 28195 6140 28207 6200
rect 28241 6140 28253 6200
rect 28195 6128 28253 6140
rect 28323 6200 28381 6212
rect 28323 6140 28335 6200
rect 28369 6140 28381 6200
rect 28323 6128 28381 6140
rect 28451 6200 28509 6212
rect 28451 6140 28463 6200
rect 28497 6140 28509 6200
rect 28451 6128 28509 6140
rect 28579 6200 28637 6212
rect 28579 6140 28591 6200
rect 28625 6140 28637 6200
rect 28579 6128 28637 6140
rect -329 5278 -271 5290
rect -329 5218 -317 5278
rect -283 5218 -271 5278
rect -329 5206 -271 5218
rect -201 5278 -143 5290
rect -201 5218 -189 5278
rect -155 5218 -143 5278
rect -201 5206 -143 5218
rect 599 5278 657 5290
rect 599 5218 611 5278
rect 645 5218 657 5278
rect 599 5206 657 5218
rect 727 5278 785 5290
rect 727 5218 739 5278
rect 773 5218 785 5278
rect 727 5206 785 5218
rect 855 5278 913 5290
rect 855 5218 867 5278
rect 901 5218 913 5278
rect 855 5206 913 5218
rect 1863 5278 1921 5290
rect 1863 5218 1875 5278
rect 1909 5218 1921 5278
rect 1863 5206 1921 5218
rect 1991 5278 2049 5290
rect 1991 5218 2003 5278
rect 2037 5218 2049 5278
rect 1991 5206 2049 5218
rect 2119 5278 2177 5290
rect 2119 5218 2131 5278
rect 2165 5218 2177 5278
rect 2119 5206 2177 5218
rect 2247 5278 2305 5290
rect 2247 5218 2259 5278
rect 2293 5218 2305 5278
rect 2247 5206 2305 5218
rect 2375 5278 2433 5290
rect 2375 5218 2387 5278
rect 2421 5218 2433 5278
rect 2375 5206 2433 5218
rect 3482 5278 3540 5290
rect 3482 5218 3494 5278
rect 3528 5218 3540 5278
rect 3482 5206 3540 5218
rect 3610 5278 3668 5290
rect 3610 5218 3622 5278
rect 3656 5218 3668 5278
rect 3610 5206 3668 5218
rect 3738 5278 3796 5290
rect 3738 5218 3750 5278
rect 3784 5218 3796 5278
rect 3738 5206 3796 5218
rect 3866 5278 3924 5290
rect 3866 5218 3878 5278
rect 3912 5218 3924 5278
rect 3866 5206 3924 5218
rect 3994 5278 4052 5290
rect 3994 5218 4006 5278
rect 4040 5218 4052 5278
rect 3994 5206 4052 5218
rect 4122 5278 4180 5290
rect 4122 5218 4134 5278
rect 4168 5218 4180 5278
rect 4122 5206 4180 5218
rect 4250 5278 4308 5290
rect 4250 5218 4262 5278
rect 4296 5218 4308 5278
rect 4250 5206 4308 5218
rect 4378 5278 4436 5290
rect 4378 5218 4390 5278
rect 4424 5218 4436 5278
rect 4378 5206 4436 5218
rect 4506 5278 4564 5290
rect 4506 5218 4518 5278
rect 4552 5218 4564 5278
rect 4506 5206 4564 5218
rect 8047 5278 8105 5290
rect 8047 5218 8059 5278
rect 8093 5218 8105 5278
rect 8047 5206 8105 5218
rect 8175 5278 8233 5290
rect 8175 5218 8187 5278
rect 8221 5218 8233 5278
rect 8175 5206 8233 5218
rect 8303 5278 8361 5290
rect 8303 5218 8315 5278
rect 8349 5218 8361 5278
rect 8303 5206 8361 5218
rect 8431 5278 8489 5290
rect 8431 5218 8443 5278
rect 8477 5218 8489 5278
rect 8431 5206 8489 5218
rect 8559 5278 8617 5290
rect 8559 5218 8571 5278
rect 8605 5218 8617 5278
rect 8559 5206 8617 5218
rect 8687 5278 8745 5290
rect 8687 5218 8699 5278
rect 8733 5218 8745 5278
rect 8687 5206 8745 5218
rect 8815 5278 8873 5290
rect 8815 5218 8827 5278
rect 8861 5218 8873 5278
rect 8815 5206 8873 5218
rect 8943 5278 9001 5290
rect 8943 5218 8955 5278
rect 8989 5218 9001 5278
rect 8943 5206 9001 5218
rect 9071 5278 9129 5290
rect 9071 5218 9083 5278
rect 9117 5218 9129 5278
rect 9071 5206 9129 5218
rect 9199 5278 9257 5290
rect 9199 5218 9211 5278
rect 9245 5218 9257 5278
rect 9199 5206 9257 5218
rect 9327 5278 9385 5290
rect 9327 5218 9339 5278
rect 9373 5218 9385 5278
rect 9327 5206 9385 5218
rect 9455 5278 9513 5290
rect 9455 5218 9467 5278
rect 9501 5218 9513 5278
rect 9455 5206 9513 5218
rect 9583 5278 9641 5290
rect 9583 5218 9595 5278
rect 9629 5218 9641 5278
rect 9583 5206 9641 5218
rect 9711 5278 9769 5290
rect 9711 5218 9723 5278
rect 9757 5218 9769 5278
rect 9711 5206 9769 5218
rect 9839 5278 9897 5290
rect 9839 5218 9851 5278
rect 9885 5218 9897 5278
rect 9839 5206 9897 5218
rect 9967 5278 10025 5290
rect 9967 5218 9979 5278
rect 10013 5218 10025 5278
rect 9967 5206 10025 5218
rect 10095 5278 10153 5290
rect 10095 5218 10107 5278
rect 10141 5218 10153 5278
rect 10095 5206 10153 5218
rect 15811 5278 15869 5290
rect 15811 5218 15823 5278
rect 15857 5218 15869 5278
rect 15811 5206 15869 5218
rect 15939 5278 15997 5290
rect 15939 5218 15951 5278
rect 15985 5218 15997 5278
rect 15939 5206 15997 5218
rect 16067 5278 16125 5290
rect 16067 5218 16079 5278
rect 16113 5218 16125 5278
rect 16067 5206 16125 5218
rect 16195 5278 16253 5290
rect 16195 5218 16207 5278
rect 16241 5218 16253 5278
rect 16195 5206 16253 5218
rect 16323 5278 16381 5290
rect 16323 5218 16335 5278
rect 16369 5218 16381 5278
rect 16323 5206 16381 5218
rect 16451 5278 16509 5290
rect 16451 5218 16463 5278
rect 16497 5218 16509 5278
rect 16451 5206 16509 5218
rect 16579 5278 16637 5290
rect 16579 5218 16591 5278
rect 16625 5218 16637 5278
rect 16579 5206 16637 5218
rect 16707 5278 16765 5290
rect 16707 5218 16719 5278
rect 16753 5218 16765 5278
rect 16707 5206 16765 5218
rect 16835 5278 16893 5290
rect 16835 5218 16847 5278
rect 16881 5218 16893 5278
rect 16835 5206 16893 5218
rect 16963 5278 17021 5290
rect 16963 5218 16975 5278
rect 17009 5218 17021 5278
rect 16963 5206 17021 5218
rect 17091 5278 17149 5290
rect 17091 5218 17103 5278
rect 17137 5218 17149 5278
rect 17091 5206 17149 5218
rect 17219 5278 17277 5290
rect 17219 5218 17231 5278
rect 17265 5218 17277 5278
rect 17219 5206 17277 5218
rect 17347 5278 17405 5290
rect 17347 5218 17359 5278
rect 17393 5218 17405 5278
rect 17347 5206 17405 5218
rect 17475 5278 17533 5290
rect 17475 5218 17487 5278
rect 17521 5218 17533 5278
rect 17475 5206 17533 5218
rect 17603 5278 17661 5290
rect 17603 5218 17615 5278
rect 17649 5218 17661 5278
rect 17603 5206 17661 5218
rect 17731 5278 17789 5290
rect 17731 5218 17743 5278
rect 17777 5218 17789 5278
rect 17731 5206 17789 5218
rect 17859 5278 17917 5290
rect 17859 5218 17871 5278
rect 17905 5218 17917 5278
rect 17859 5206 17917 5218
rect 17987 5278 18045 5290
rect 17987 5218 17999 5278
rect 18033 5218 18045 5278
rect 17987 5206 18045 5218
rect 18115 5278 18173 5290
rect 18115 5218 18127 5278
rect 18161 5218 18173 5278
rect 18115 5206 18173 5218
rect 18243 5278 18301 5290
rect 18243 5218 18255 5278
rect 18289 5218 18301 5278
rect 18243 5206 18301 5218
rect 18371 5278 18429 5290
rect 18371 5218 18383 5278
rect 18417 5218 18429 5278
rect 18371 5206 18429 5218
rect 18499 5278 18557 5290
rect 18499 5218 18511 5278
rect 18545 5218 18557 5278
rect 18499 5206 18557 5218
rect 18627 5278 18685 5290
rect 18627 5218 18639 5278
rect 18673 5218 18685 5278
rect 18627 5206 18685 5218
rect 18755 5278 18813 5290
rect 18755 5218 18767 5278
rect 18801 5218 18813 5278
rect 18755 5206 18813 5218
rect 18883 5278 18941 5290
rect 18883 5218 18895 5278
rect 18929 5218 18941 5278
rect 18883 5206 18941 5218
rect 19011 5278 19069 5290
rect 19011 5218 19023 5278
rect 19057 5218 19069 5278
rect 19011 5206 19069 5218
rect 19139 5278 19197 5290
rect 19139 5218 19151 5278
rect 19185 5218 19197 5278
rect 19139 5206 19197 5218
rect 19267 5278 19325 5290
rect 19267 5218 19279 5278
rect 19313 5218 19325 5278
rect 19267 5206 19325 5218
rect 19395 5278 19453 5290
rect 19395 5218 19407 5278
rect 19441 5218 19453 5278
rect 19395 5206 19453 5218
rect 19523 5278 19581 5290
rect 19523 5218 19535 5278
rect 19569 5218 19581 5278
rect 19523 5206 19581 5218
rect 19651 5278 19709 5290
rect 19651 5218 19663 5278
rect 19697 5218 19709 5278
rect 19651 5206 19709 5218
rect 19779 5278 19837 5290
rect 19779 5218 19791 5278
rect 19825 5218 19837 5278
rect 19779 5206 19837 5218
rect 19907 5278 19965 5290
rect 19907 5218 19919 5278
rect 19953 5218 19965 5278
rect 19907 5206 19965 5218
rect 29355 5278 29413 5290
rect 29355 5218 29367 5278
rect 29401 5218 29413 5278
rect 29355 5206 29413 5218
rect 29483 5278 29541 5290
rect 29483 5218 29495 5278
rect 29529 5218 29541 5278
rect 29483 5206 29541 5218
rect 29611 5278 29669 5290
rect 29611 5218 29623 5278
rect 29657 5218 29669 5278
rect 29611 5206 29669 5218
rect 29739 5278 29797 5290
rect 29739 5218 29751 5278
rect 29785 5218 29797 5278
rect 29739 5206 29797 5218
rect 29867 5278 29925 5290
rect 29867 5218 29879 5278
rect 29913 5218 29925 5278
rect 29867 5206 29925 5218
rect 29995 5278 30053 5290
rect 29995 5218 30007 5278
rect 30041 5218 30053 5278
rect 29995 5206 30053 5218
rect 30123 5278 30181 5290
rect 30123 5218 30135 5278
rect 30169 5218 30181 5278
rect 30123 5206 30181 5218
rect 30251 5278 30309 5290
rect 30251 5218 30263 5278
rect 30297 5218 30309 5278
rect 30251 5206 30309 5218
rect 30379 5278 30437 5290
rect 30379 5218 30391 5278
rect 30425 5218 30437 5278
rect 30379 5206 30437 5218
rect 30507 5278 30565 5290
rect 30507 5218 30519 5278
rect 30553 5218 30565 5278
rect 30507 5206 30565 5218
rect 30635 5278 30693 5290
rect 30635 5218 30647 5278
rect 30681 5218 30693 5278
rect 30635 5206 30693 5218
rect 30763 5278 30821 5290
rect 30763 5218 30775 5278
rect 30809 5218 30821 5278
rect 30763 5206 30821 5218
rect 30891 5278 30949 5290
rect 30891 5218 30903 5278
rect 30937 5218 30949 5278
rect 30891 5206 30949 5218
rect 31019 5278 31077 5290
rect 31019 5218 31031 5278
rect 31065 5218 31077 5278
rect 31019 5206 31077 5218
rect 31147 5278 31205 5290
rect 31147 5218 31159 5278
rect 31193 5218 31205 5278
rect 31147 5206 31205 5218
rect 31275 5278 31333 5290
rect 31275 5218 31287 5278
rect 31321 5218 31333 5278
rect 31275 5206 31333 5218
rect 31403 5278 31461 5290
rect 31403 5218 31415 5278
rect 31449 5218 31461 5278
rect 31403 5206 31461 5218
rect 31531 5278 31589 5290
rect 31531 5218 31543 5278
rect 31577 5218 31589 5278
rect 31531 5206 31589 5218
rect 31659 5278 31717 5290
rect 31659 5218 31671 5278
rect 31705 5218 31717 5278
rect 31659 5206 31717 5218
rect 31787 5278 31845 5290
rect 31787 5218 31799 5278
rect 31833 5218 31845 5278
rect 31787 5206 31845 5218
rect 31915 5278 31973 5290
rect 31915 5218 31927 5278
rect 31961 5218 31973 5278
rect 31915 5206 31973 5218
rect 32043 5278 32101 5290
rect 32043 5218 32055 5278
rect 32089 5218 32101 5278
rect 32043 5206 32101 5218
rect 32171 5278 32229 5290
rect 32171 5218 32183 5278
rect 32217 5218 32229 5278
rect 32171 5206 32229 5218
rect 32299 5278 32357 5290
rect 32299 5218 32311 5278
rect 32345 5218 32357 5278
rect 32299 5206 32357 5218
rect 32427 5278 32485 5290
rect 32427 5218 32439 5278
rect 32473 5218 32485 5278
rect 32427 5206 32485 5218
rect 32555 5278 32613 5290
rect 32555 5218 32567 5278
rect 32601 5218 32613 5278
rect 32555 5206 32613 5218
rect 32683 5278 32741 5290
rect 32683 5218 32695 5278
rect 32729 5218 32741 5278
rect 32683 5206 32741 5218
rect 32811 5278 32869 5290
rect 32811 5218 32823 5278
rect 32857 5218 32869 5278
rect 32811 5206 32869 5218
rect 32939 5278 32997 5290
rect 32939 5218 32951 5278
rect 32985 5218 32997 5278
rect 32939 5206 32997 5218
rect 33067 5278 33125 5290
rect 33067 5218 33079 5278
rect 33113 5218 33125 5278
rect 33067 5206 33125 5218
rect 33195 5278 33253 5290
rect 33195 5218 33207 5278
rect 33241 5218 33253 5278
rect 33195 5206 33253 5218
rect 33323 5278 33381 5290
rect 33323 5218 33335 5278
rect 33369 5218 33381 5278
rect 33323 5206 33381 5218
rect 33451 5278 33509 5290
rect 33451 5218 33463 5278
rect 33497 5218 33509 5278
rect 33451 5206 33509 5218
rect 33579 5278 33637 5290
rect 33579 5218 33591 5278
rect 33625 5218 33637 5278
rect 33579 5206 33637 5218
rect 33707 5278 33765 5290
rect 33707 5218 33719 5278
rect 33753 5218 33765 5278
rect 33707 5206 33765 5218
rect 33835 5278 33893 5290
rect 33835 5218 33847 5278
rect 33881 5218 33893 5278
rect 33835 5206 33893 5218
rect 33963 5278 34021 5290
rect 33963 5218 33975 5278
rect 34009 5218 34021 5278
rect 33963 5206 34021 5218
rect 34091 5278 34149 5290
rect 34091 5218 34103 5278
rect 34137 5218 34149 5278
rect 34091 5206 34149 5218
rect 34219 5278 34277 5290
rect 34219 5218 34231 5278
rect 34265 5218 34277 5278
rect 34219 5206 34277 5218
rect 34347 5278 34405 5290
rect 34347 5218 34359 5278
rect 34393 5218 34405 5278
rect 34347 5206 34405 5218
rect 34475 5278 34533 5290
rect 34475 5218 34487 5278
rect 34521 5218 34533 5278
rect 34475 5206 34533 5218
rect 34603 5278 34661 5290
rect 34603 5218 34615 5278
rect 34649 5218 34661 5278
rect 34603 5206 34661 5218
rect 34731 5278 34789 5290
rect 34731 5218 34743 5278
rect 34777 5218 34789 5278
rect 34731 5206 34789 5218
rect 34859 5278 34917 5290
rect 34859 5218 34871 5278
rect 34905 5218 34917 5278
rect 34859 5206 34917 5218
rect 34987 5278 35045 5290
rect 34987 5218 34999 5278
rect 35033 5218 35045 5278
rect 34987 5206 35045 5218
rect 35115 5278 35173 5290
rect 35115 5218 35127 5278
rect 35161 5218 35173 5278
rect 35115 5206 35173 5218
rect 35243 5278 35301 5290
rect 35243 5218 35255 5278
rect 35289 5218 35301 5278
rect 35243 5206 35301 5218
rect 35371 5278 35429 5290
rect 35371 5218 35383 5278
rect 35417 5218 35429 5278
rect 35371 5206 35429 5218
rect 35499 5278 35557 5290
rect 35499 5218 35511 5278
rect 35545 5218 35557 5278
rect 35499 5206 35557 5218
rect 35627 5278 35685 5290
rect 35627 5218 35639 5278
rect 35673 5218 35685 5278
rect 35627 5206 35685 5218
rect 35755 5278 35813 5290
rect 35755 5218 35767 5278
rect 35801 5218 35813 5278
rect 35755 5206 35813 5218
rect 35883 5278 35941 5290
rect 35883 5218 35895 5278
rect 35929 5218 35941 5278
rect 35883 5206 35941 5218
rect 36011 5278 36069 5290
rect 36011 5218 36023 5278
rect 36057 5218 36069 5278
rect 36011 5206 36069 5218
rect 36139 5278 36197 5290
rect 36139 5218 36151 5278
rect 36185 5218 36197 5278
rect 36139 5206 36197 5218
rect 36267 5278 36325 5290
rect 36267 5218 36279 5278
rect 36313 5218 36325 5278
rect 36267 5206 36325 5218
rect 36395 5278 36453 5290
rect 36395 5218 36407 5278
rect 36441 5218 36453 5278
rect 36395 5206 36453 5218
rect 36523 5278 36581 5290
rect 36523 5218 36535 5278
rect 36569 5218 36581 5278
rect 36523 5206 36581 5218
rect 36651 5278 36709 5290
rect 36651 5218 36663 5278
rect 36697 5218 36709 5278
rect 36651 5206 36709 5218
rect 36779 5278 36837 5290
rect 36779 5218 36791 5278
rect 36825 5218 36837 5278
rect 36779 5206 36837 5218
rect 36907 5278 36965 5290
rect 36907 5218 36919 5278
rect 36953 5218 36965 5278
rect 36907 5206 36965 5218
rect 37035 5278 37093 5290
rect 37035 5218 37047 5278
rect 37081 5218 37093 5278
rect 37035 5206 37093 5218
rect 37163 5278 37221 5290
rect 37163 5218 37175 5278
rect 37209 5218 37221 5278
rect 37163 5206 37221 5218
rect 37291 5278 37349 5290
rect 37291 5218 37303 5278
rect 37337 5218 37349 5278
rect 37291 5206 37349 5218
rect 37419 5278 37477 5290
rect 37419 5218 37431 5278
rect 37465 5218 37477 5278
rect 37419 5206 37477 5218
rect 37547 5278 37605 5290
rect 37547 5218 37559 5278
rect 37593 5218 37605 5278
rect 37547 5206 37605 5218
<< pdiff >>
rect -329 5984 -271 5996
rect -329 5840 -317 5984
rect -283 5840 -271 5984
rect -329 5828 -271 5840
rect -201 5984 -143 5996
rect -201 5840 -189 5984
rect -155 5840 -143 5984
rect -201 5828 -143 5840
rect 471 5984 529 5996
rect 471 5840 483 5984
rect 517 5840 529 5984
rect 471 5828 529 5840
rect 599 5984 657 5996
rect 599 5840 611 5984
rect 645 5840 657 5984
rect 599 5828 657 5840
rect 727 5984 785 5996
rect 727 5840 739 5984
rect 773 5840 785 5984
rect 727 5828 785 5840
rect 1351 5984 1409 5996
rect 1351 5840 1363 5984
rect 1397 5840 1409 5984
rect 1351 5828 1409 5840
rect 1479 5984 1537 5996
rect 1479 5840 1491 5984
rect 1525 5840 1537 5984
rect 1479 5828 1537 5840
rect 1607 5984 1665 5996
rect 1607 5840 1619 5984
rect 1653 5840 1665 5984
rect 1607 5828 1665 5840
rect 1735 5984 1793 5996
rect 1735 5840 1747 5984
rect 1781 5840 1793 5984
rect 1735 5828 1793 5840
rect 1863 5984 1921 5996
rect 1863 5840 1875 5984
rect 1909 5840 1921 5984
rect 1863 5828 1921 5840
rect 2970 5984 3028 5996
rect 2970 5840 2982 5984
rect 3016 5840 3028 5984
rect 2970 5828 3028 5840
rect 3098 5984 3156 5996
rect 3098 5840 3110 5984
rect 3144 5840 3156 5984
rect 3098 5828 3156 5840
rect 3226 5984 3284 5996
rect 3226 5840 3238 5984
rect 3272 5840 3284 5984
rect 3226 5828 3284 5840
rect 3354 5984 3412 5996
rect 3354 5840 3366 5984
rect 3400 5840 3412 5984
rect 3354 5828 3412 5840
rect 3482 5984 3540 5996
rect 3482 5840 3494 5984
rect 3528 5840 3540 5984
rect 3482 5828 3540 5840
rect 3610 5984 3668 5996
rect 3610 5840 3622 5984
rect 3656 5840 3668 5984
rect 3610 5828 3668 5840
rect 3738 5984 3796 5996
rect 3738 5840 3750 5984
rect 3784 5840 3796 5984
rect 3738 5828 3796 5840
rect 3866 5984 3924 5996
rect 3866 5840 3878 5984
rect 3912 5840 3924 5984
rect 3866 5828 3924 5840
rect 3994 5984 4052 5996
rect 3994 5840 4006 5984
rect 4040 5840 4052 5984
rect 3994 5828 4052 5840
rect 5463 5984 5521 5996
rect 5463 5840 5475 5984
rect 5509 5840 5521 5984
rect 5463 5828 5521 5840
rect 5591 5984 5649 5996
rect 5591 5840 5603 5984
rect 5637 5840 5649 5984
rect 5591 5828 5649 5840
rect 5719 5984 5777 5996
rect 5719 5840 5731 5984
rect 5765 5840 5777 5984
rect 5719 5828 5777 5840
rect 5847 5984 5905 5996
rect 5847 5840 5859 5984
rect 5893 5840 5905 5984
rect 5847 5828 5905 5840
rect 5975 5984 6033 5996
rect 5975 5840 5987 5984
rect 6021 5840 6033 5984
rect 5975 5828 6033 5840
rect 6103 5984 6161 5996
rect 6103 5840 6115 5984
rect 6149 5840 6161 5984
rect 6103 5828 6161 5840
rect 6231 5984 6289 5996
rect 6231 5840 6243 5984
rect 6277 5840 6289 5984
rect 6231 5828 6289 5840
rect 6359 5984 6417 5996
rect 6359 5840 6371 5984
rect 6405 5840 6417 5984
rect 6359 5828 6417 5840
rect 6487 5984 6545 5996
rect 6487 5840 6499 5984
rect 6533 5840 6545 5984
rect 6487 5828 6545 5840
rect 6615 5984 6673 5996
rect 6615 5840 6627 5984
rect 6661 5840 6673 5984
rect 6615 5828 6673 5840
rect 6743 5984 6801 5996
rect 6743 5840 6755 5984
rect 6789 5840 6801 5984
rect 6743 5828 6801 5840
rect 6871 5984 6929 5996
rect 6871 5840 6883 5984
rect 6917 5840 6929 5984
rect 6871 5828 6929 5840
rect 6999 5984 7057 5996
rect 6999 5840 7011 5984
rect 7045 5840 7057 5984
rect 6999 5828 7057 5840
rect 7127 5984 7185 5996
rect 7127 5840 7139 5984
rect 7173 5840 7185 5984
rect 7127 5828 7185 5840
rect 7255 5984 7313 5996
rect 7255 5840 7267 5984
rect 7301 5840 7313 5984
rect 7255 5828 7313 5840
rect 7383 5984 7441 5996
rect 7383 5840 7395 5984
rect 7429 5840 7441 5984
rect 7383 5828 7441 5840
rect 7511 5984 7569 5996
rect 7511 5840 7523 5984
rect 7557 5840 7569 5984
rect 7511 5828 7569 5840
rect 10550 5984 10608 5996
rect 10550 5840 10562 5984
rect 10596 5840 10608 5984
rect 10550 5828 10608 5840
rect 10678 5984 10736 5996
rect 10678 5840 10690 5984
rect 10724 5840 10736 5984
rect 10678 5828 10736 5840
rect 10806 5984 10864 5996
rect 10806 5840 10818 5984
rect 10852 5840 10864 5984
rect 10806 5828 10864 5840
rect 10934 5984 10992 5996
rect 10934 5840 10946 5984
rect 10980 5840 10992 5984
rect 10934 5828 10992 5840
rect 11062 5984 11120 5996
rect 11062 5840 11074 5984
rect 11108 5840 11120 5984
rect 11062 5828 11120 5840
rect 11190 5984 11248 5996
rect 11190 5840 11202 5984
rect 11236 5840 11248 5984
rect 11190 5828 11248 5840
rect 11318 5984 11376 5996
rect 11318 5840 11330 5984
rect 11364 5840 11376 5984
rect 11318 5828 11376 5840
rect 11446 5984 11504 5996
rect 11446 5840 11458 5984
rect 11492 5840 11504 5984
rect 11446 5828 11504 5840
rect 11574 5984 11632 5996
rect 11574 5840 11586 5984
rect 11620 5840 11632 5984
rect 11574 5828 11632 5840
rect 11702 5984 11760 5996
rect 11702 5840 11714 5984
rect 11748 5840 11760 5984
rect 11702 5828 11760 5840
rect 11830 5984 11888 5996
rect 11830 5840 11842 5984
rect 11876 5840 11888 5984
rect 11830 5828 11888 5840
rect 11958 5984 12016 5996
rect 11958 5840 11970 5984
rect 12004 5840 12016 5984
rect 11958 5828 12016 5840
rect 12086 5984 12144 5996
rect 12086 5840 12098 5984
rect 12132 5840 12144 5984
rect 12086 5828 12144 5840
rect 12214 5984 12272 5996
rect 12214 5840 12226 5984
rect 12260 5840 12272 5984
rect 12214 5828 12272 5840
rect 12342 5984 12400 5996
rect 12342 5840 12354 5984
rect 12388 5840 12400 5984
rect 12342 5828 12400 5840
rect 12470 5984 12528 5996
rect 12470 5840 12482 5984
rect 12516 5840 12528 5984
rect 12470 5828 12528 5840
rect 12598 5984 12656 5996
rect 12598 5840 12610 5984
rect 12644 5840 12656 5984
rect 12598 5828 12656 5840
rect 12726 5984 12784 5996
rect 12726 5840 12738 5984
rect 12772 5840 12784 5984
rect 12726 5828 12784 5840
rect 12854 5984 12912 5996
rect 12854 5840 12866 5984
rect 12900 5840 12912 5984
rect 12854 5828 12912 5840
rect 12982 5984 13040 5996
rect 12982 5840 12994 5984
rect 13028 5840 13040 5984
rect 12982 5828 13040 5840
rect 13110 5984 13168 5996
rect 13110 5840 13122 5984
rect 13156 5840 13168 5984
rect 13110 5828 13168 5840
rect 13238 5984 13296 5996
rect 13238 5840 13250 5984
rect 13284 5840 13296 5984
rect 13238 5828 13296 5840
rect 13366 5984 13424 5996
rect 13366 5840 13378 5984
rect 13412 5840 13424 5984
rect 13366 5828 13424 5840
rect 13494 5984 13552 5996
rect 13494 5840 13506 5984
rect 13540 5840 13552 5984
rect 13494 5828 13552 5840
rect 13622 5984 13680 5996
rect 13622 5840 13634 5984
rect 13668 5840 13680 5984
rect 13622 5828 13680 5840
rect 13750 5984 13808 5996
rect 13750 5840 13762 5984
rect 13796 5840 13808 5984
rect 13750 5828 13808 5840
rect 13878 5984 13936 5996
rect 13878 5840 13890 5984
rect 13924 5840 13936 5984
rect 13878 5828 13936 5840
rect 14006 5984 14064 5996
rect 14006 5840 14018 5984
rect 14052 5840 14064 5984
rect 14006 5828 14064 5840
rect 14134 5984 14192 5996
rect 14134 5840 14146 5984
rect 14180 5840 14192 5984
rect 14134 5828 14192 5840
rect 14262 5984 14320 5996
rect 14262 5840 14274 5984
rect 14308 5840 14320 5984
rect 14262 5828 14320 5840
rect 14390 5984 14448 5996
rect 14390 5840 14402 5984
rect 14436 5840 14448 5984
rect 14390 5828 14448 5840
rect 14518 5984 14576 5996
rect 14518 5840 14530 5984
rect 14564 5840 14576 5984
rect 14518 5828 14576 5840
rect 14646 5984 14704 5996
rect 14646 5840 14658 5984
rect 14692 5840 14704 5984
rect 14646 5828 14704 5840
rect 20387 5984 20445 5996
rect 20387 5840 20399 5984
rect 20433 5840 20445 5984
rect 20387 5828 20445 5840
rect 20515 5984 20573 5996
rect 20515 5840 20527 5984
rect 20561 5840 20573 5984
rect 20515 5828 20573 5840
rect 20643 5984 20701 5996
rect 20643 5840 20655 5984
rect 20689 5840 20701 5984
rect 20643 5828 20701 5840
rect 20771 5984 20829 5996
rect 20771 5840 20783 5984
rect 20817 5840 20829 5984
rect 20771 5828 20829 5840
rect 20899 5984 20957 5996
rect 20899 5840 20911 5984
rect 20945 5840 20957 5984
rect 20899 5828 20957 5840
rect 21027 5984 21085 5996
rect 21027 5840 21039 5984
rect 21073 5840 21085 5984
rect 21027 5828 21085 5840
rect 21155 5984 21213 5996
rect 21155 5840 21167 5984
rect 21201 5840 21213 5984
rect 21155 5828 21213 5840
rect 21283 5984 21341 5996
rect 21283 5840 21295 5984
rect 21329 5840 21341 5984
rect 21283 5828 21341 5840
rect 21411 5984 21469 5996
rect 21411 5840 21423 5984
rect 21457 5840 21469 5984
rect 21411 5828 21469 5840
rect 21539 5984 21597 5996
rect 21539 5840 21551 5984
rect 21585 5840 21597 5984
rect 21539 5828 21597 5840
rect 21667 5984 21725 5996
rect 21667 5840 21679 5984
rect 21713 5840 21725 5984
rect 21667 5828 21725 5840
rect 21795 5984 21853 5996
rect 21795 5840 21807 5984
rect 21841 5840 21853 5984
rect 21795 5828 21853 5840
rect 21923 5984 21981 5996
rect 21923 5840 21935 5984
rect 21969 5840 21981 5984
rect 21923 5828 21981 5840
rect 22051 5984 22109 5996
rect 22051 5840 22063 5984
rect 22097 5840 22109 5984
rect 22051 5828 22109 5840
rect 22179 5984 22237 5996
rect 22179 5840 22191 5984
rect 22225 5840 22237 5984
rect 22179 5828 22237 5840
rect 22307 5984 22365 5996
rect 22307 5840 22319 5984
rect 22353 5840 22365 5984
rect 22307 5828 22365 5840
rect 22435 5984 22493 5996
rect 22435 5840 22447 5984
rect 22481 5840 22493 5984
rect 22435 5828 22493 5840
rect 22563 5984 22621 5996
rect 22563 5840 22575 5984
rect 22609 5840 22621 5984
rect 22563 5828 22621 5840
rect 22691 5984 22749 5996
rect 22691 5840 22703 5984
rect 22737 5840 22749 5984
rect 22691 5828 22749 5840
rect 22819 5984 22877 5996
rect 22819 5840 22831 5984
rect 22865 5840 22877 5984
rect 22819 5828 22877 5840
rect 22947 5984 23005 5996
rect 22947 5840 22959 5984
rect 22993 5840 23005 5984
rect 22947 5828 23005 5840
rect 23075 5984 23133 5996
rect 23075 5840 23087 5984
rect 23121 5840 23133 5984
rect 23075 5828 23133 5840
rect 23203 5984 23261 5996
rect 23203 5840 23215 5984
rect 23249 5840 23261 5984
rect 23203 5828 23261 5840
rect 23331 5984 23389 5996
rect 23331 5840 23343 5984
rect 23377 5840 23389 5984
rect 23331 5828 23389 5840
rect 23459 5984 23517 5996
rect 23459 5840 23471 5984
rect 23505 5840 23517 5984
rect 23459 5828 23517 5840
rect 23587 5984 23645 5996
rect 23587 5840 23599 5984
rect 23633 5840 23645 5984
rect 23587 5828 23645 5840
rect 23715 5984 23773 5996
rect 23715 5840 23727 5984
rect 23761 5840 23773 5984
rect 23715 5828 23773 5840
rect 23843 5984 23901 5996
rect 23843 5840 23855 5984
rect 23889 5840 23901 5984
rect 23843 5828 23901 5840
rect 23971 5984 24029 5996
rect 23971 5840 23983 5984
rect 24017 5840 24029 5984
rect 23971 5828 24029 5840
rect 24099 5984 24157 5996
rect 24099 5840 24111 5984
rect 24145 5840 24157 5984
rect 24099 5828 24157 5840
rect 24227 5984 24285 5996
rect 24227 5840 24239 5984
rect 24273 5840 24285 5984
rect 24227 5828 24285 5840
rect 24355 5984 24413 5996
rect 24355 5840 24367 5984
rect 24401 5840 24413 5984
rect 24355 5828 24413 5840
rect 24483 5984 24541 5996
rect 24483 5840 24495 5984
rect 24529 5840 24541 5984
rect 24483 5828 24541 5840
rect 24611 5984 24669 5996
rect 24611 5840 24623 5984
rect 24657 5840 24669 5984
rect 24611 5828 24669 5840
rect 24739 5984 24797 5996
rect 24739 5840 24751 5984
rect 24785 5840 24797 5984
rect 24739 5828 24797 5840
rect 24867 5984 24925 5996
rect 24867 5840 24879 5984
rect 24913 5840 24925 5984
rect 24867 5828 24925 5840
rect 24995 5984 25053 5996
rect 24995 5840 25007 5984
rect 25041 5840 25053 5984
rect 24995 5828 25053 5840
rect 25123 5984 25181 5996
rect 25123 5840 25135 5984
rect 25169 5840 25181 5984
rect 25123 5828 25181 5840
rect 25251 5984 25309 5996
rect 25251 5840 25263 5984
rect 25297 5840 25309 5984
rect 25251 5828 25309 5840
rect 25379 5984 25437 5996
rect 25379 5840 25391 5984
rect 25425 5840 25437 5984
rect 25379 5828 25437 5840
rect 25507 5984 25565 5996
rect 25507 5840 25519 5984
rect 25553 5840 25565 5984
rect 25507 5828 25565 5840
rect 25635 5984 25693 5996
rect 25635 5840 25647 5984
rect 25681 5840 25693 5984
rect 25635 5828 25693 5840
rect 25763 5984 25821 5996
rect 25763 5840 25775 5984
rect 25809 5840 25821 5984
rect 25763 5828 25821 5840
rect 25891 5984 25949 5996
rect 25891 5840 25903 5984
rect 25937 5840 25949 5984
rect 25891 5828 25949 5840
rect 26019 5984 26077 5996
rect 26019 5840 26031 5984
rect 26065 5840 26077 5984
rect 26019 5828 26077 5840
rect 26147 5984 26205 5996
rect 26147 5840 26159 5984
rect 26193 5840 26205 5984
rect 26147 5828 26205 5840
rect 26275 5984 26333 5996
rect 26275 5840 26287 5984
rect 26321 5840 26333 5984
rect 26275 5828 26333 5840
rect 26403 5984 26461 5996
rect 26403 5840 26415 5984
rect 26449 5840 26461 5984
rect 26403 5828 26461 5840
rect 26531 5984 26589 5996
rect 26531 5840 26543 5984
rect 26577 5840 26589 5984
rect 26531 5828 26589 5840
rect 26659 5984 26717 5996
rect 26659 5840 26671 5984
rect 26705 5840 26717 5984
rect 26659 5828 26717 5840
rect 26787 5984 26845 5996
rect 26787 5840 26799 5984
rect 26833 5840 26845 5984
rect 26787 5828 26845 5840
rect 26915 5984 26973 5996
rect 26915 5840 26927 5984
rect 26961 5840 26973 5984
rect 26915 5828 26973 5840
rect 27043 5984 27101 5996
rect 27043 5840 27055 5984
rect 27089 5840 27101 5984
rect 27043 5828 27101 5840
rect 27171 5984 27229 5996
rect 27171 5840 27183 5984
rect 27217 5840 27229 5984
rect 27171 5828 27229 5840
rect 27299 5984 27357 5996
rect 27299 5840 27311 5984
rect 27345 5840 27357 5984
rect 27299 5828 27357 5840
rect 27427 5984 27485 5996
rect 27427 5840 27439 5984
rect 27473 5840 27485 5984
rect 27427 5828 27485 5840
rect 27555 5984 27613 5996
rect 27555 5840 27567 5984
rect 27601 5840 27613 5984
rect 27555 5828 27613 5840
rect 27683 5984 27741 5996
rect 27683 5840 27695 5984
rect 27729 5840 27741 5984
rect 27683 5828 27741 5840
rect 27811 5984 27869 5996
rect 27811 5840 27823 5984
rect 27857 5840 27869 5984
rect 27811 5828 27869 5840
rect 27939 5984 27997 5996
rect 27939 5840 27951 5984
rect 27985 5840 27997 5984
rect 27939 5828 27997 5840
rect 28067 5984 28125 5996
rect 28067 5840 28079 5984
rect 28113 5840 28125 5984
rect 28067 5828 28125 5840
rect 28195 5984 28253 5996
rect 28195 5840 28207 5984
rect 28241 5840 28253 5984
rect 28195 5828 28253 5840
rect 28323 5984 28381 5996
rect 28323 5840 28335 5984
rect 28369 5840 28381 5984
rect 28323 5828 28381 5840
rect 28451 5984 28509 5996
rect 28451 5840 28463 5984
rect 28497 5840 28509 5984
rect 28451 5828 28509 5840
rect 28579 5984 28637 5996
rect 28579 5840 28591 5984
rect 28625 5840 28637 5984
rect 28579 5828 28637 5840
rect -329 5578 -271 5590
rect -329 5434 -317 5578
rect -283 5434 -271 5578
rect -329 5422 -271 5434
rect -201 5578 -143 5590
rect -201 5434 -189 5578
rect -155 5434 -143 5578
rect -201 5422 -143 5434
rect 599 5578 657 5590
rect 599 5434 611 5578
rect 645 5434 657 5578
rect 599 5422 657 5434
rect 727 5578 785 5590
rect 727 5434 739 5578
rect 773 5434 785 5578
rect 727 5422 785 5434
rect 855 5578 913 5590
rect 855 5434 867 5578
rect 901 5434 913 5578
rect 1863 5578 1921 5590
rect 855 5422 913 5434
rect 1863 5434 1875 5578
rect 1909 5434 1921 5578
rect 1863 5422 1921 5434
rect 1991 5578 2049 5590
rect 1991 5434 2003 5578
rect 2037 5434 2049 5578
rect 1991 5422 2049 5434
rect 2119 5578 2177 5590
rect 2119 5434 2131 5578
rect 2165 5434 2177 5578
rect 2119 5422 2177 5434
rect 2247 5578 2305 5590
rect 2247 5434 2259 5578
rect 2293 5434 2305 5578
rect 2247 5422 2305 5434
rect 2375 5578 2433 5590
rect 2375 5434 2387 5578
rect 2421 5434 2433 5578
rect 3482 5578 3540 5590
rect 2375 5422 2433 5434
rect 3482 5434 3494 5578
rect 3528 5434 3540 5578
rect 3482 5422 3540 5434
rect 3610 5578 3668 5590
rect 3610 5434 3622 5578
rect 3656 5434 3668 5578
rect 3610 5422 3668 5434
rect 3738 5578 3796 5590
rect 3738 5434 3750 5578
rect 3784 5434 3796 5578
rect 3738 5422 3796 5434
rect 3866 5578 3924 5590
rect 3866 5434 3878 5578
rect 3912 5434 3924 5578
rect 3866 5422 3924 5434
rect 3994 5578 4052 5590
rect 3994 5434 4006 5578
rect 4040 5434 4052 5578
rect 3994 5422 4052 5434
rect 4122 5578 4180 5590
rect 4122 5434 4134 5578
rect 4168 5434 4180 5578
rect 4122 5422 4180 5434
rect 4250 5578 4308 5590
rect 4250 5434 4262 5578
rect 4296 5434 4308 5578
rect 4250 5422 4308 5434
rect 4378 5578 4436 5590
rect 4378 5434 4390 5578
rect 4424 5434 4436 5578
rect 4378 5422 4436 5434
rect 4506 5578 4564 5590
rect 4506 5434 4518 5578
rect 4552 5434 4564 5578
rect 8047 5578 8105 5590
rect 4506 5422 4564 5434
rect 8047 5434 8059 5578
rect 8093 5434 8105 5578
rect 8047 5422 8105 5434
rect 8175 5578 8233 5590
rect 8175 5434 8187 5578
rect 8221 5434 8233 5578
rect 8175 5422 8233 5434
rect 8303 5578 8361 5590
rect 8303 5434 8315 5578
rect 8349 5434 8361 5578
rect 8303 5422 8361 5434
rect 8431 5578 8489 5590
rect 8431 5434 8443 5578
rect 8477 5434 8489 5578
rect 8431 5422 8489 5434
rect 8559 5578 8617 5590
rect 8559 5434 8571 5578
rect 8605 5434 8617 5578
rect 8559 5422 8617 5434
rect 8687 5578 8745 5590
rect 8687 5434 8699 5578
rect 8733 5434 8745 5578
rect 8687 5422 8745 5434
rect 8815 5578 8873 5590
rect 8815 5434 8827 5578
rect 8861 5434 8873 5578
rect 8815 5422 8873 5434
rect 8943 5578 9001 5590
rect 8943 5434 8955 5578
rect 8989 5434 9001 5578
rect 8943 5422 9001 5434
rect 9071 5578 9129 5590
rect 9071 5434 9083 5578
rect 9117 5434 9129 5578
rect 9071 5422 9129 5434
rect 9199 5578 9257 5590
rect 9199 5434 9211 5578
rect 9245 5434 9257 5578
rect 9199 5422 9257 5434
rect 9327 5578 9385 5590
rect 9327 5434 9339 5578
rect 9373 5434 9385 5578
rect 9327 5422 9385 5434
rect 9455 5578 9513 5590
rect 9455 5434 9467 5578
rect 9501 5434 9513 5578
rect 9455 5422 9513 5434
rect 9583 5578 9641 5590
rect 9583 5434 9595 5578
rect 9629 5434 9641 5578
rect 9583 5422 9641 5434
rect 9711 5578 9769 5590
rect 9711 5434 9723 5578
rect 9757 5434 9769 5578
rect 9711 5422 9769 5434
rect 9839 5578 9897 5590
rect 9839 5434 9851 5578
rect 9885 5434 9897 5578
rect 9839 5422 9897 5434
rect 9967 5578 10025 5590
rect 9967 5434 9979 5578
rect 10013 5434 10025 5578
rect 9967 5422 10025 5434
rect 10095 5578 10153 5590
rect 10095 5434 10107 5578
rect 10141 5434 10153 5578
rect 10095 5422 10153 5434
rect 15811 5578 15869 5590
rect 15811 5434 15823 5578
rect 15857 5434 15869 5578
rect 15811 5422 15869 5434
rect 15939 5578 15997 5590
rect 15939 5434 15951 5578
rect 15985 5434 15997 5578
rect 15939 5422 15997 5434
rect 16067 5578 16125 5590
rect 16067 5434 16079 5578
rect 16113 5434 16125 5578
rect 16067 5422 16125 5434
rect 16195 5578 16253 5590
rect 16195 5434 16207 5578
rect 16241 5434 16253 5578
rect 16195 5422 16253 5434
rect 16323 5578 16381 5590
rect 16323 5434 16335 5578
rect 16369 5434 16381 5578
rect 16323 5422 16381 5434
rect 16451 5578 16509 5590
rect 16451 5434 16463 5578
rect 16497 5434 16509 5578
rect 16451 5422 16509 5434
rect 16579 5578 16637 5590
rect 16579 5434 16591 5578
rect 16625 5434 16637 5578
rect 16579 5422 16637 5434
rect 16707 5578 16765 5590
rect 16707 5434 16719 5578
rect 16753 5434 16765 5578
rect 16707 5422 16765 5434
rect 16835 5578 16893 5590
rect 16835 5434 16847 5578
rect 16881 5434 16893 5578
rect 16835 5422 16893 5434
rect 16963 5578 17021 5590
rect 16963 5434 16975 5578
rect 17009 5434 17021 5578
rect 16963 5422 17021 5434
rect 17091 5578 17149 5590
rect 17091 5434 17103 5578
rect 17137 5434 17149 5578
rect 17091 5422 17149 5434
rect 17219 5578 17277 5590
rect 17219 5434 17231 5578
rect 17265 5434 17277 5578
rect 17219 5422 17277 5434
rect 17347 5578 17405 5590
rect 17347 5434 17359 5578
rect 17393 5434 17405 5578
rect 17347 5422 17405 5434
rect 17475 5578 17533 5590
rect 17475 5434 17487 5578
rect 17521 5434 17533 5578
rect 17475 5422 17533 5434
rect 17603 5578 17661 5590
rect 17603 5434 17615 5578
rect 17649 5434 17661 5578
rect 17603 5422 17661 5434
rect 17731 5578 17789 5590
rect 17731 5434 17743 5578
rect 17777 5434 17789 5578
rect 17731 5422 17789 5434
rect 17859 5578 17917 5590
rect 17859 5434 17871 5578
rect 17905 5434 17917 5578
rect 17859 5422 17917 5434
rect 17987 5578 18045 5590
rect 17987 5434 17999 5578
rect 18033 5434 18045 5578
rect 17987 5422 18045 5434
rect 18115 5578 18173 5590
rect 18115 5434 18127 5578
rect 18161 5434 18173 5578
rect 18115 5422 18173 5434
rect 18243 5578 18301 5590
rect 18243 5434 18255 5578
rect 18289 5434 18301 5578
rect 18243 5422 18301 5434
rect 18371 5578 18429 5590
rect 18371 5434 18383 5578
rect 18417 5434 18429 5578
rect 18371 5422 18429 5434
rect 18499 5578 18557 5590
rect 18499 5434 18511 5578
rect 18545 5434 18557 5578
rect 18499 5422 18557 5434
rect 18627 5578 18685 5590
rect 18627 5434 18639 5578
rect 18673 5434 18685 5578
rect 18627 5422 18685 5434
rect 18755 5578 18813 5590
rect 18755 5434 18767 5578
rect 18801 5434 18813 5578
rect 18755 5422 18813 5434
rect 18883 5578 18941 5590
rect 18883 5434 18895 5578
rect 18929 5434 18941 5578
rect 18883 5422 18941 5434
rect 19011 5578 19069 5590
rect 19011 5434 19023 5578
rect 19057 5434 19069 5578
rect 19011 5422 19069 5434
rect 19139 5578 19197 5590
rect 19139 5434 19151 5578
rect 19185 5434 19197 5578
rect 19139 5422 19197 5434
rect 19267 5578 19325 5590
rect 19267 5434 19279 5578
rect 19313 5434 19325 5578
rect 19267 5422 19325 5434
rect 19395 5578 19453 5590
rect 19395 5434 19407 5578
rect 19441 5434 19453 5578
rect 19395 5422 19453 5434
rect 19523 5578 19581 5590
rect 19523 5434 19535 5578
rect 19569 5434 19581 5578
rect 19523 5422 19581 5434
rect 19651 5578 19709 5590
rect 19651 5434 19663 5578
rect 19697 5434 19709 5578
rect 19651 5422 19709 5434
rect 19779 5578 19837 5590
rect 19779 5434 19791 5578
rect 19825 5434 19837 5578
rect 19779 5422 19837 5434
rect 19907 5578 19965 5590
rect 19907 5434 19919 5578
rect 19953 5434 19965 5578
rect 19907 5422 19965 5434
rect 29355 5578 29413 5590
rect 29355 5434 29367 5578
rect 29401 5434 29413 5578
rect 29355 5422 29413 5434
rect 29483 5578 29541 5590
rect 29483 5434 29495 5578
rect 29529 5434 29541 5578
rect 29483 5422 29541 5434
rect 29611 5578 29669 5590
rect 29611 5434 29623 5578
rect 29657 5434 29669 5578
rect 29611 5422 29669 5434
rect 29739 5578 29797 5590
rect 29739 5434 29751 5578
rect 29785 5434 29797 5578
rect 29739 5422 29797 5434
rect 29867 5578 29925 5590
rect 29867 5434 29879 5578
rect 29913 5434 29925 5578
rect 29867 5422 29925 5434
rect 29995 5578 30053 5590
rect 29995 5434 30007 5578
rect 30041 5434 30053 5578
rect 29995 5422 30053 5434
rect 30123 5578 30181 5590
rect 30123 5434 30135 5578
rect 30169 5434 30181 5578
rect 30123 5422 30181 5434
rect 30251 5578 30309 5590
rect 30251 5434 30263 5578
rect 30297 5434 30309 5578
rect 30251 5422 30309 5434
rect 30379 5578 30437 5590
rect 30379 5434 30391 5578
rect 30425 5434 30437 5578
rect 30379 5422 30437 5434
rect 30507 5578 30565 5590
rect 30507 5434 30519 5578
rect 30553 5434 30565 5578
rect 30507 5422 30565 5434
rect 30635 5578 30693 5590
rect 30635 5434 30647 5578
rect 30681 5434 30693 5578
rect 30635 5422 30693 5434
rect 30763 5578 30821 5590
rect 30763 5434 30775 5578
rect 30809 5434 30821 5578
rect 30763 5422 30821 5434
rect 30891 5578 30949 5590
rect 30891 5434 30903 5578
rect 30937 5434 30949 5578
rect 30891 5422 30949 5434
rect 31019 5578 31077 5590
rect 31019 5434 31031 5578
rect 31065 5434 31077 5578
rect 31019 5422 31077 5434
rect 31147 5578 31205 5590
rect 31147 5434 31159 5578
rect 31193 5434 31205 5578
rect 31147 5422 31205 5434
rect 31275 5578 31333 5590
rect 31275 5434 31287 5578
rect 31321 5434 31333 5578
rect 31275 5422 31333 5434
rect 31403 5578 31461 5590
rect 31403 5434 31415 5578
rect 31449 5434 31461 5578
rect 31403 5422 31461 5434
rect 31531 5578 31589 5590
rect 31531 5434 31543 5578
rect 31577 5434 31589 5578
rect 31531 5422 31589 5434
rect 31659 5578 31717 5590
rect 31659 5434 31671 5578
rect 31705 5434 31717 5578
rect 31659 5422 31717 5434
rect 31787 5578 31845 5590
rect 31787 5434 31799 5578
rect 31833 5434 31845 5578
rect 31787 5422 31845 5434
rect 31915 5578 31973 5590
rect 31915 5434 31927 5578
rect 31961 5434 31973 5578
rect 31915 5422 31973 5434
rect 32043 5578 32101 5590
rect 32043 5434 32055 5578
rect 32089 5434 32101 5578
rect 32043 5422 32101 5434
rect 32171 5578 32229 5590
rect 32171 5434 32183 5578
rect 32217 5434 32229 5578
rect 32171 5422 32229 5434
rect 32299 5578 32357 5590
rect 32299 5434 32311 5578
rect 32345 5434 32357 5578
rect 32299 5422 32357 5434
rect 32427 5578 32485 5590
rect 32427 5434 32439 5578
rect 32473 5434 32485 5578
rect 32427 5422 32485 5434
rect 32555 5578 32613 5590
rect 32555 5434 32567 5578
rect 32601 5434 32613 5578
rect 32555 5422 32613 5434
rect 32683 5578 32741 5590
rect 32683 5434 32695 5578
rect 32729 5434 32741 5578
rect 32683 5422 32741 5434
rect 32811 5578 32869 5590
rect 32811 5434 32823 5578
rect 32857 5434 32869 5578
rect 32811 5422 32869 5434
rect 32939 5578 32997 5590
rect 32939 5434 32951 5578
rect 32985 5434 32997 5578
rect 32939 5422 32997 5434
rect 33067 5578 33125 5590
rect 33067 5434 33079 5578
rect 33113 5434 33125 5578
rect 33067 5422 33125 5434
rect 33195 5578 33253 5590
rect 33195 5434 33207 5578
rect 33241 5434 33253 5578
rect 33195 5422 33253 5434
rect 33323 5578 33381 5590
rect 33323 5434 33335 5578
rect 33369 5434 33381 5578
rect 33323 5422 33381 5434
rect 33451 5578 33509 5590
rect 33451 5434 33463 5578
rect 33497 5434 33509 5578
rect 33451 5422 33509 5434
rect 33579 5578 33637 5590
rect 33579 5434 33591 5578
rect 33625 5434 33637 5578
rect 33579 5422 33637 5434
rect 33707 5578 33765 5590
rect 33707 5434 33719 5578
rect 33753 5434 33765 5578
rect 33707 5422 33765 5434
rect 33835 5578 33893 5590
rect 33835 5434 33847 5578
rect 33881 5434 33893 5578
rect 33835 5422 33893 5434
rect 33963 5578 34021 5590
rect 33963 5434 33975 5578
rect 34009 5434 34021 5578
rect 33963 5422 34021 5434
rect 34091 5578 34149 5590
rect 34091 5434 34103 5578
rect 34137 5434 34149 5578
rect 34091 5422 34149 5434
rect 34219 5578 34277 5590
rect 34219 5434 34231 5578
rect 34265 5434 34277 5578
rect 34219 5422 34277 5434
rect 34347 5578 34405 5590
rect 34347 5434 34359 5578
rect 34393 5434 34405 5578
rect 34347 5422 34405 5434
rect 34475 5578 34533 5590
rect 34475 5434 34487 5578
rect 34521 5434 34533 5578
rect 34475 5422 34533 5434
rect 34603 5578 34661 5590
rect 34603 5434 34615 5578
rect 34649 5434 34661 5578
rect 34603 5422 34661 5434
rect 34731 5578 34789 5590
rect 34731 5434 34743 5578
rect 34777 5434 34789 5578
rect 34731 5422 34789 5434
rect 34859 5578 34917 5590
rect 34859 5434 34871 5578
rect 34905 5434 34917 5578
rect 34859 5422 34917 5434
rect 34987 5578 35045 5590
rect 34987 5434 34999 5578
rect 35033 5434 35045 5578
rect 34987 5422 35045 5434
rect 35115 5578 35173 5590
rect 35115 5434 35127 5578
rect 35161 5434 35173 5578
rect 35115 5422 35173 5434
rect 35243 5578 35301 5590
rect 35243 5434 35255 5578
rect 35289 5434 35301 5578
rect 35243 5422 35301 5434
rect 35371 5578 35429 5590
rect 35371 5434 35383 5578
rect 35417 5434 35429 5578
rect 35371 5422 35429 5434
rect 35499 5578 35557 5590
rect 35499 5434 35511 5578
rect 35545 5434 35557 5578
rect 35499 5422 35557 5434
rect 35627 5578 35685 5590
rect 35627 5434 35639 5578
rect 35673 5434 35685 5578
rect 35627 5422 35685 5434
rect 35755 5578 35813 5590
rect 35755 5434 35767 5578
rect 35801 5434 35813 5578
rect 35755 5422 35813 5434
rect 35883 5578 35941 5590
rect 35883 5434 35895 5578
rect 35929 5434 35941 5578
rect 35883 5422 35941 5434
rect 36011 5578 36069 5590
rect 36011 5434 36023 5578
rect 36057 5434 36069 5578
rect 36011 5422 36069 5434
rect 36139 5578 36197 5590
rect 36139 5434 36151 5578
rect 36185 5434 36197 5578
rect 36139 5422 36197 5434
rect 36267 5578 36325 5590
rect 36267 5434 36279 5578
rect 36313 5434 36325 5578
rect 36267 5422 36325 5434
rect 36395 5578 36453 5590
rect 36395 5434 36407 5578
rect 36441 5434 36453 5578
rect 36395 5422 36453 5434
rect 36523 5578 36581 5590
rect 36523 5434 36535 5578
rect 36569 5434 36581 5578
rect 36523 5422 36581 5434
rect 36651 5578 36709 5590
rect 36651 5434 36663 5578
rect 36697 5434 36709 5578
rect 36651 5422 36709 5434
rect 36779 5578 36837 5590
rect 36779 5434 36791 5578
rect 36825 5434 36837 5578
rect 36779 5422 36837 5434
rect 36907 5578 36965 5590
rect 36907 5434 36919 5578
rect 36953 5434 36965 5578
rect 36907 5422 36965 5434
rect 37035 5578 37093 5590
rect 37035 5434 37047 5578
rect 37081 5434 37093 5578
rect 37035 5422 37093 5434
rect 37163 5578 37221 5590
rect 37163 5434 37175 5578
rect 37209 5434 37221 5578
rect 37163 5422 37221 5434
rect 37291 5578 37349 5590
rect 37291 5434 37303 5578
rect 37337 5434 37349 5578
rect 37291 5422 37349 5434
rect 37419 5578 37477 5590
rect 37419 5434 37431 5578
rect 37465 5434 37477 5578
rect 37419 5422 37477 5434
rect 37547 5578 37605 5590
rect 37547 5434 37559 5578
rect 37593 5434 37605 5578
rect 37547 5422 37605 5434
<< ndiffc >>
rect -317 6140 -283 6200
rect -189 6140 -155 6200
rect 483 6140 517 6200
rect 611 6140 645 6200
rect 739 6140 773 6200
rect 1363 6140 1397 6200
rect 1491 6140 1525 6200
rect 1619 6140 1653 6200
rect 1747 6140 1781 6200
rect 1875 6140 1909 6200
rect 2982 6140 3016 6200
rect 3110 6140 3144 6200
rect 3238 6140 3272 6200
rect 3366 6140 3400 6200
rect 3494 6140 3528 6200
rect 3622 6140 3656 6200
rect 3750 6140 3784 6200
rect 3878 6140 3912 6200
rect 4006 6140 4040 6200
rect 5475 6140 5509 6200
rect 5603 6140 5637 6200
rect 5731 6140 5765 6200
rect 5859 6140 5893 6200
rect 5987 6140 6021 6200
rect 6115 6140 6149 6200
rect 6243 6140 6277 6200
rect 6371 6140 6405 6200
rect 6499 6140 6533 6200
rect 6627 6140 6661 6200
rect 6755 6140 6789 6200
rect 6883 6140 6917 6200
rect 7011 6140 7045 6200
rect 7139 6140 7173 6200
rect 7267 6140 7301 6200
rect 7395 6140 7429 6200
rect 7523 6140 7557 6200
rect 10562 6140 10596 6200
rect 10690 6140 10724 6200
rect 10818 6140 10852 6200
rect 10946 6140 10980 6200
rect 11074 6140 11108 6200
rect 11202 6140 11236 6200
rect 11330 6140 11364 6200
rect 11458 6140 11492 6200
rect 11586 6140 11620 6200
rect 11714 6140 11748 6200
rect 11842 6140 11876 6200
rect 11970 6140 12004 6200
rect 12098 6140 12132 6200
rect 12226 6140 12260 6200
rect 12354 6140 12388 6200
rect 12482 6140 12516 6200
rect 12610 6140 12644 6200
rect 12738 6140 12772 6200
rect 12866 6140 12900 6200
rect 12994 6140 13028 6200
rect 13122 6140 13156 6200
rect 13250 6140 13284 6200
rect 13378 6140 13412 6200
rect 13506 6140 13540 6200
rect 13634 6140 13668 6200
rect 13762 6140 13796 6200
rect 13890 6140 13924 6200
rect 14018 6140 14052 6200
rect 14146 6140 14180 6200
rect 14274 6140 14308 6200
rect 14402 6140 14436 6200
rect 14530 6140 14564 6200
rect 14658 6140 14692 6200
rect 20399 6140 20433 6200
rect 20527 6140 20561 6200
rect 20655 6140 20689 6200
rect 20783 6140 20817 6200
rect 20911 6140 20945 6200
rect 21039 6140 21073 6200
rect 21167 6140 21201 6200
rect 21295 6140 21329 6200
rect 21423 6140 21457 6200
rect 21551 6140 21585 6200
rect 21679 6140 21713 6200
rect 21807 6140 21841 6200
rect 21935 6140 21969 6200
rect 22063 6140 22097 6200
rect 22191 6140 22225 6200
rect 22319 6140 22353 6200
rect 22447 6140 22481 6200
rect 22575 6140 22609 6200
rect 22703 6140 22737 6200
rect 22831 6140 22865 6200
rect 22959 6140 22993 6200
rect 23087 6140 23121 6200
rect 23215 6140 23249 6200
rect 23343 6140 23377 6200
rect 23471 6140 23505 6200
rect 23599 6140 23633 6200
rect 23727 6140 23761 6200
rect 23855 6140 23889 6200
rect 23983 6140 24017 6200
rect 24111 6140 24145 6200
rect 24239 6140 24273 6200
rect 24367 6140 24401 6200
rect 24495 6140 24529 6200
rect 24623 6140 24657 6200
rect 24751 6140 24785 6200
rect 24879 6140 24913 6200
rect 25007 6140 25041 6200
rect 25135 6140 25169 6200
rect 25263 6140 25297 6200
rect 25391 6140 25425 6200
rect 25519 6140 25553 6200
rect 25647 6140 25681 6200
rect 25775 6140 25809 6200
rect 25903 6140 25937 6200
rect 26031 6140 26065 6200
rect 26159 6140 26193 6200
rect 26287 6140 26321 6200
rect 26415 6140 26449 6200
rect 26543 6140 26577 6200
rect 26671 6140 26705 6200
rect 26799 6140 26833 6200
rect 26927 6140 26961 6200
rect 27055 6140 27089 6200
rect 27183 6140 27217 6200
rect 27311 6140 27345 6200
rect 27439 6140 27473 6200
rect 27567 6140 27601 6200
rect 27695 6140 27729 6200
rect 27823 6140 27857 6200
rect 27951 6140 27985 6200
rect 28079 6140 28113 6200
rect 28207 6140 28241 6200
rect 28335 6140 28369 6200
rect 28463 6140 28497 6200
rect 28591 6140 28625 6200
rect -317 5218 -283 5278
rect -189 5218 -155 5278
rect 611 5218 645 5278
rect 739 5218 773 5278
rect 867 5218 901 5278
rect 1875 5218 1909 5278
rect 2003 5218 2037 5278
rect 2131 5218 2165 5278
rect 2259 5218 2293 5278
rect 2387 5218 2421 5278
rect 3494 5218 3528 5278
rect 3622 5218 3656 5278
rect 3750 5218 3784 5278
rect 3878 5218 3912 5278
rect 4006 5218 4040 5278
rect 4134 5218 4168 5278
rect 4262 5218 4296 5278
rect 4390 5218 4424 5278
rect 4518 5218 4552 5278
rect 8059 5218 8093 5278
rect 8187 5218 8221 5278
rect 8315 5218 8349 5278
rect 8443 5218 8477 5278
rect 8571 5218 8605 5278
rect 8699 5218 8733 5278
rect 8827 5218 8861 5278
rect 8955 5218 8989 5278
rect 9083 5218 9117 5278
rect 9211 5218 9245 5278
rect 9339 5218 9373 5278
rect 9467 5218 9501 5278
rect 9595 5218 9629 5278
rect 9723 5218 9757 5278
rect 9851 5218 9885 5278
rect 9979 5218 10013 5278
rect 10107 5218 10141 5278
rect 15823 5218 15857 5278
rect 15951 5218 15985 5278
rect 16079 5218 16113 5278
rect 16207 5218 16241 5278
rect 16335 5218 16369 5278
rect 16463 5218 16497 5278
rect 16591 5218 16625 5278
rect 16719 5218 16753 5278
rect 16847 5218 16881 5278
rect 16975 5218 17009 5278
rect 17103 5218 17137 5278
rect 17231 5218 17265 5278
rect 17359 5218 17393 5278
rect 17487 5218 17521 5278
rect 17615 5218 17649 5278
rect 17743 5218 17777 5278
rect 17871 5218 17905 5278
rect 17999 5218 18033 5278
rect 18127 5218 18161 5278
rect 18255 5218 18289 5278
rect 18383 5218 18417 5278
rect 18511 5218 18545 5278
rect 18639 5218 18673 5278
rect 18767 5218 18801 5278
rect 18895 5218 18929 5278
rect 19023 5218 19057 5278
rect 19151 5218 19185 5278
rect 19279 5218 19313 5278
rect 19407 5218 19441 5278
rect 19535 5218 19569 5278
rect 19663 5218 19697 5278
rect 19791 5218 19825 5278
rect 19919 5218 19953 5278
rect 29367 5218 29401 5278
rect 29495 5218 29529 5278
rect 29623 5218 29657 5278
rect 29751 5218 29785 5278
rect 29879 5218 29913 5278
rect 30007 5218 30041 5278
rect 30135 5218 30169 5278
rect 30263 5218 30297 5278
rect 30391 5218 30425 5278
rect 30519 5218 30553 5278
rect 30647 5218 30681 5278
rect 30775 5218 30809 5278
rect 30903 5218 30937 5278
rect 31031 5218 31065 5278
rect 31159 5218 31193 5278
rect 31287 5218 31321 5278
rect 31415 5218 31449 5278
rect 31543 5218 31577 5278
rect 31671 5218 31705 5278
rect 31799 5218 31833 5278
rect 31927 5218 31961 5278
rect 32055 5218 32089 5278
rect 32183 5218 32217 5278
rect 32311 5218 32345 5278
rect 32439 5218 32473 5278
rect 32567 5218 32601 5278
rect 32695 5218 32729 5278
rect 32823 5218 32857 5278
rect 32951 5218 32985 5278
rect 33079 5218 33113 5278
rect 33207 5218 33241 5278
rect 33335 5218 33369 5278
rect 33463 5218 33497 5278
rect 33591 5218 33625 5278
rect 33719 5218 33753 5278
rect 33847 5218 33881 5278
rect 33975 5218 34009 5278
rect 34103 5218 34137 5278
rect 34231 5218 34265 5278
rect 34359 5218 34393 5278
rect 34487 5218 34521 5278
rect 34615 5218 34649 5278
rect 34743 5218 34777 5278
rect 34871 5218 34905 5278
rect 34999 5218 35033 5278
rect 35127 5218 35161 5278
rect 35255 5218 35289 5278
rect 35383 5218 35417 5278
rect 35511 5218 35545 5278
rect 35639 5218 35673 5278
rect 35767 5218 35801 5278
rect 35895 5218 35929 5278
rect 36023 5218 36057 5278
rect 36151 5218 36185 5278
rect 36279 5218 36313 5278
rect 36407 5218 36441 5278
rect 36535 5218 36569 5278
rect 36663 5218 36697 5278
rect 36791 5218 36825 5278
rect 36919 5218 36953 5278
rect 37047 5218 37081 5278
rect 37175 5218 37209 5278
rect 37303 5218 37337 5278
rect 37431 5218 37465 5278
rect 37559 5218 37593 5278
<< pdiffc >>
rect -317 5840 -283 5984
rect -189 5840 -155 5984
rect 483 5840 517 5984
rect 611 5840 645 5984
rect 739 5840 773 5984
rect 1363 5840 1397 5984
rect 1491 5840 1525 5984
rect 1619 5840 1653 5984
rect 1747 5840 1781 5984
rect 1875 5840 1909 5984
rect 2982 5840 3016 5984
rect 3110 5840 3144 5984
rect 3238 5840 3272 5984
rect 3366 5840 3400 5984
rect 3494 5840 3528 5984
rect 3622 5840 3656 5984
rect 3750 5840 3784 5984
rect 3878 5840 3912 5984
rect 4006 5840 4040 5984
rect 5475 5840 5509 5984
rect 5603 5840 5637 5984
rect 5731 5840 5765 5984
rect 5859 5840 5893 5984
rect 5987 5840 6021 5984
rect 6115 5840 6149 5984
rect 6243 5840 6277 5984
rect 6371 5840 6405 5984
rect 6499 5840 6533 5984
rect 6627 5840 6661 5984
rect 6755 5840 6789 5984
rect 6883 5840 6917 5984
rect 7011 5840 7045 5984
rect 7139 5840 7173 5984
rect 7267 5840 7301 5984
rect 7395 5840 7429 5984
rect 7523 5840 7557 5984
rect 10562 5840 10596 5984
rect 10690 5840 10724 5984
rect 10818 5840 10852 5984
rect 10946 5840 10980 5984
rect 11074 5840 11108 5984
rect 11202 5840 11236 5984
rect 11330 5840 11364 5984
rect 11458 5840 11492 5984
rect 11586 5840 11620 5984
rect 11714 5840 11748 5984
rect 11842 5840 11876 5984
rect 11970 5840 12004 5984
rect 12098 5840 12132 5984
rect 12226 5840 12260 5984
rect 12354 5840 12388 5984
rect 12482 5840 12516 5984
rect 12610 5840 12644 5984
rect 12738 5840 12772 5984
rect 12866 5840 12900 5984
rect 12994 5840 13028 5984
rect 13122 5840 13156 5984
rect 13250 5840 13284 5984
rect 13378 5840 13412 5984
rect 13506 5840 13540 5984
rect 13634 5840 13668 5984
rect 13762 5840 13796 5984
rect 13890 5840 13924 5984
rect 14018 5840 14052 5984
rect 14146 5840 14180 5984
rect 14274 5840 14308 5984
rect 14402 5840 14436 5984
rect 14530 5840 14564 5984
rect 14658 5840 14692 5984
rect 20399 5840 20433 5984
rect 20527 5840 20561 5984
rect 20655 5840 20689 5984
rect 20783 5840 20817 5984
rect 20911 5840 20945 5984
rect 21039 5840 21073 5984
rect 21167 5840 21201 5984
rect 21295 5840 21329 5984
rect 21423 5840 21457 5984
rect 21551 5840 21585 5984
rect 21679 5840 21713 5984
rect 21807 5840 21841 5984
rect 21935 5840 21969 5984
rect 22063 5840 22097 5984
rect 22191 5840 22225 5984
rect 22319 5840 22353 5984
rect 22447 5840 22481 5984
rect 22575 5840 22609 5984
rect 22703 5840 22737 5984
rect 22831 5840 22865 5984
rect 22959 5840 22993 5984
rect 23087 5840 23121 5984
rect 23215 5840 23249 5984
rect 23343 5840 23377 5984
rect 23471 5840 23505 5984
rect 23599 5840 23633 5984
rect 23727 5840 23761 5984
rect 23855 5840 23889 5984
rect 23983 5840 24017 5984
rect 24111 5840 24145 5984
rect 24239 5840 24273 5984
rect 24367 5840 24401 5984
rect 24495 5840 24529 5984
rect 24623 5840 24657 5984
rect 24751 5840 24785 5984
rect 24879 5840 24913 5984
rect 25007 5840 25041 5984
rect 25135 5840 25169 5984
rect 25263 5840 25297 5984
rect 25391 5840 25425 5984
rect 25519 5840 25553 5984
rect 25647 5840 25681 5984
rect 25775 5840 25809 5984
rect 25903 5840 25937 5984
rect 26031 5840 26065 5984
rect 26159 5840 26193 5984
rect 26287 5840 26321 5984
rect 26415 5840 26449 5984
rect 26543 5840 26577 5984
rect 26671 5840 26705 5984
rect 26799 5840 26833 5984
rect 26927 5840 26961 5984
rect 27055 5840 27089 5984
rect 27183 5840 27217 5984
rect 27311 5840 27345 5984
rect 27439 5840 27473 5984
rect 27567 5840 27601 5984
rect 27695 5840 27729 5984
rect 27823 5840 27857 5984
rect 27951 5840 27985 5984
rect 28079 5840 28113 5984
rect 28207 5840 28241 5984
rect 28335 5840 28369 5984
rect 28463 5840 28497 5984
rect 28591 5840 28625 5984
rect -317 5434 -283 5578
rect -189 5434 -155 5578
rect 611 5434 645 5578
rect 739 5434 773 5578
rect 867 5434 901 5578
rect 1875 5434 1909 5578
rect 2003 5434 2037 5578
rect 2131 5434 2165 5578
rect 2259 5434 2293 5578
rect 2387 5434 2421 5578
rect 3494 5434 3528 5578
rect 3622 5434 3656 5578
rect 3750 5434 3784 5578
rect 3878 5434 3912 5578
rect 4006 5434 4040 5578
rect 4134 5434 4168 5578
rect 4262 5434 4296 5578
rect 4390 5434 4424 5578
rect 4518 5434 4552 5578
rect 8059 5434 8093 5578
rect 8187 5434 8221 5578
rect 8315 5434 8349 5578
rect 8443 5434 8477 5578
rect 8571 5434 8605 5578
rect 8699 5434 8733 5578
rect 8827 5434 8861 5578
rect 8955 5434 8989 5578
rect 9083 5434 9117 5578
rect 9211 5434 9245 5578
rect 9339 5434 9373 5578
rect 9467 5434 9501 5578
rect 9595 5434 9629 5578
rect 9723 5434 9757 5578
rect 9851 5434 9885 5578
rect 9979 5434 10013 5578
rect 10107 5434 10141 5578
rect 15823 5434 15857 5578
rect 15951 5434 15985 5578
rect 16079 5434 16113 5578
rect 16207 5434 16241 5578
rect 16335 5434 16369 5578
rect 16463 5434 16497 5578
rect 16591 5434 16625 5578
rect 16719 5434 16753 5578
rect 16847 5434 16881 5578
rect 16975 5434 17009 5578
rect 17103 5434 17137 5578
rect 17231 5434 17265 5578
rect 17359 5434 17393 5578
rect 17487 5434 17521 5578
rect 17615 5434 17649 5578
rect 17743 5434 17777 5578
rect 17871 5434 17905 5578
rect 17999 5434 18033 5578
rect 18127 5434 18161 5578
rect 18255 5434 18289 5578
rect 18383 5434 18417 5578
rect 18511 5434 18545 5578
rect 18639 5434 18673 5578
rect 18767 5434 18801 5578
rect 18895 5434 18929 5578
rect 19023 5434 19057 5578
rect 19151 5434 19185 5578
rect 19279 5434 19313 5578
rect 19407 5434 19441 5578
rect 19535 5434 19569 5578
rect 19663 5434 19697 5578
rect 19791 5434 19825 5578
rect 19919 5434 19953 5578
rect 29367 5434 29401 5578
rect 29495 5434 29529 5578
rect 29623 5434 29657 5578
rect 29751 5434 29785 5578
rect 29879 5434 29913 5578
rect 30007 5434 30041 5578
rect 30135 5434 30169 5578
rect 30263 5434 30297 5578
rect 30391 5434 30425 5578
rect 30519 5434 30553 5578
rect 30647 5434 30681 5578
rect 30775 5434 30809 5578
rect 30903 5434 30937 5578
rect 31031 5434 31065 5578
rect 31159 5434 31193 5578
rect 31287 5434 31321 5578
rect 31415 5434 31449 5578
rect 31543 5434 31577 5578
rect 31671 5434 31705 5578
rect 31799 5434 31833 5578
rect 31927 5434 31961 5578
rect 32055 5434 32089 5578
rect 32183 5434 32217 5578
rect 32311 5434 32345 5578
rect 32439 5434 32473 5578
rect 32567 5434 32601 5578
rect 32695 5434 32729 5578
rect 32823 5434 32857 5578
rect 32951 5434 32985 5578
rect 33079 5434 33113 5578
rect 33207 5434 33241 5578
rect 33335 5434 33369 5578
rect 33463 5434 33497 5578
rect 33591 5434 33625 5578
rect 33719 5434 33753 5578
rect 33847 5434 33881 5578
rect 33975 5434 34009 5578
rect 34103 5434 34137 5578
rect 34231 5434 34265 5578
rect 34359 5434 34393 5578
rect 34487 5434 34521 5578
rect 34615 5434 34649 5578
rect 34743 5434 34777 5578
rect 34871 5434 34905 5578
rect 34999 5434 35033 5578
rect 35127 5434 35161 5578
rect 35255 5434 35289 5578
rect 35383 5434 35417 5578
rect 35511 5434 35545 5578
rect 35639 5434 35673 5578
rect 35767 5434 35801 5578
rect 35895 5434 35929 5578
rect 36023 5434 36057 5578
rect 36151 5434 36185 5578
rect 36279 5434 36313 5578
rect 36407 5434 36441 5578
rect 36535 5434 36569 5578
rect 36663 5434 36697 5578
rect 36791 5434 36825 5578
rect 36919 5434 36953 5578
rect 37047 5434 37081 5578
rect 37175 5434 37209 5578
rect 37303 5434 37337 5578
rect 37431 5434 37465 5578
rect 37559 5434 37593 5578
<< psubdiff >>
rect -363 6308 -109 6312
rect -363 6270 -319 6308
rect -281 6270 -191 6308
rect -153 6270 -109 6308
rect -363 6266 -109 6270
rect 437 6308 819 6312
rect 437 6270 481 6308
rect 519 6270 609 6308
rect 647 6270 737 6308
rect 775 6270 819 6308
rect 437 6266 819 6270
rect 1317 6308 1955 6312
rect 1317 6270 1361 6308
rect 1399 6270 1489 6308
rect 1527 6270 1617 6308
rect 1655 6270 1745 6308
rect 1783 6270 1873 6308
rect 1911 6270 1955 6308
rect 1317 6266 1955 6270
rect 2878 6308 4086 6312
rect 2878 6270 2980 6308
rect 3018 6270 3108 6308
rect 3146 6270 3236 6308
rect 3274 6270 3364 6308
rect 3402 6270 3492 6308
rect 3530 6270 3620 6308
rect 3658 6270 3748 6308
rect 3786 6270 3876 6308
rect 3914 6270 4004 6308
rect 4042 6270 4086 6308
rect 2878 6266 4086 6270
rect 5397 6308 7603 6312
rect 5397 6270 5473 6308
rect 5511 6270 5601 6308
rect 5639 6270 5729 6308
rect 5767 6270 5857 6308
rect 5895 6270 5985 6308
rect 6023 6270 6113 6308
rect 6151 6270 6241 6308
rect 6279 6270 6369 6308
rect 6407 6270 6497 6308
rect 6535 6270 6625 6308
rect 6663 6270 6753 6308
rect 6791 6270 6881 6308
rect 6919 6270 7009 6308
rect 7047 6270 7137 6308
rect 7175 6270 7265 6308
rect 7303 6270 7393 6308
rect 7431 6270 7521 6308
rect 7559 6270 7603 6308
rect 5397 6266 7603 6270
rect 10516 6308 14738 6312
rect 10516 6270 10560 6308
rect 10598 6270 10688 6308
rect 10726 6270 10816 6308
rect 10854 6270 10944 6308
rect 10982 6270 11072 6308
rect 11110 6270 11200 6308
rect 11238 6270 11328 6308
rect 11366 6270 11456 6308
rect 11494 6270 11584 6308
rect 11622 6270 11712 6308
rect 11750 6270 11840 6308
rect 11878 6270 11968 6308
rect 12006 6270 12096 6308
rect 12134 6270 12224 6308
rect 12262 6270 12352 6308
rect 12390 6270 12480 6308
rect 12518 6270 12608 6308
rect 12646 6270 12736 6308
rect 12774 6270 12864 6308
rect 12902 6270 12992 6308
rect 13030 6270 13120 6308
rect 13158 6270 13248 6308
rect 13286 6270 13376 6308
rect 13414 6270 13504 6308
rect 13542 6270 13632 6308
rect 13670 6270 13760 6308
rect 13798 6270 13888 6308
rect 13926 6270 14016 6308
rect 14054 6270 14144 6308
rect 14182 6270 14272 6308
rect 14310 6270 14400 6308
rect 14438 6270 14528 6308
rect 14566 6270 14656 6308
rect 14694 6270 14738 6308
rect 10516 6266 14738 6270
rect 20353 6308 28671 6312
rect 20353 6270 20397 6308
rect 20435 6270 20525 6308
rect 20563 6270 20653 6308
rect 20691 6270 20781 6308
rect 20819 6270 20909 6308
rect 20947 6270 21037 6308
rect 21075 6270 21165 6308
rect 21203 6270 21293 6308
rect 21331 6270 21421 6308
rect 21459 6270 21549 6308
rect 21587 6270 21677 6308
rect 21715 6270 21805 6308
rect 21843 6270 21933 6308
rect 21971 6270 22061 6308
rect 22099 6270 22189 6308
rect 22227 6270 22317 6308
rect 22355 6270 22445 6308
rect 22483 6270 22573 6308
rect 22611 6270 22701 6308
rect 22739 6270 22829 6308
rect 22867 6270 22957 6308
rect 22995 6270 23085 6308
rect 23123 6270 23213 6308
rect 23251 6270 23341 6308
rect 23379 6270 23469 6308
rect 23507 6270 23597 6308
rect 23635 6270 23725 6308
rect 23763 6270 23853 6308
rect 23891 6270 23981 6308
rect 24019 6270 24109 6308
rect 24147 6270 24237 6308
rect 24275 6270 24365 6308
rect 24403 6270 24493 6308
rect 24531 6270 24621 6308
rect 24659 6270 24749 6308
rect 24787 6270 24877 6308
rect 24915 6270 25005 6308
rect 25043 6270 25133 6308
rect 25171 6270 25261 6308
rect 25299 6270 25389 6308
rect 25427 6270 25517 6308
rect 25555 6270 25645 6308
rect 25683 6270 25773 6308
rect 25811 6270 25901 6308
rect 25939 6270 26029 6308
rect 26067 6270 26157 6308
rect 26195 6270 26285 6308
rect 26323 6270 26413 6308
rect 26451 6270 26541 6308
rect 26579 6270 26669 6308
rect 26707 6270 26797 6308
rect 26835 6270 26925 6308
rect 26963 6270 27053 6308
rect 27091 6270 27181 6308
rect 27219 6270 27309 6308
rect 27347 6270 27437 6308
rect 27475 6270 27565 6308
rect 27603 6270 27693 6308
rect 27731 6270 27821 6308
rect 27859 6270 27949 6308
rect 27987 6270 28077 6308
rect 28115 6270 28205 6308
rect 28243 6270 28333 6308
rect 28371 6270 28461 6308
rect 28499 6270 28589 6308
rect 28627 6270 28671 6308
rect 20353 6266 28671 6270
rect -363 5148 947 5152
rect -363 5110 -319 5148
rect -281 5110 -191 5148
rect -153 5110 609 5148
rect 647 5110 737 5148
rect 775 5110 865 5148
rect 903 5110 947 5148
rect -363 5106 947 5110
rect 1829 5148 2467 5152
rect 1829 5110 1873 5148
rect 1911 5110 2001 5148
rect 2039 5110 2129 5148
rect 2167 5110 2257 5148
rect 2295 5110 2385 5148
rect 2423 5110 2467 5148
rect 1829 5106 2467 5110
rect 3448 5148 37639 5152
rect 3448 5110 3492 5148
rect 3530 5110 3620 5148
rect 3658 5110 3748 5148
rect 3786 5110 3876 5148
rect 3914 5110 4004 5148
rect 4042 5110 4132 5148
rect 4170 5110 4260 5148
rect 4298 5110 4388 5148
rect 4426 5110 4516 5148
rect 4554 5110 8057 5148
rect 8095 5110 8185 5148
rect 8223 5110 8313 5148
rect 8351 5110 8441 5148
rect 8479 5110 8569 5148
rect 8607 5110 8697 5148
rect 8735 5110 8825 5148
rect 8863 5110 8953 5148
rect 8991 5110 9081 5148
rect 9119 5110 9209 5148
rect 9247 5110 9337 5148
rect 9375 5110 9465 5148
rect 9503 5110 9593 5148
rect 9631 5110 9721 5148
rect 9759 5110 9849 5148
rect 9887 5110 9977 5148
rect 10015 5110 10105 5148
rect 10143 5110 15821 5148
rect 15859 5110 15949 5148
rect 15987 5110 16077 5148
rect 16115 5110 16205 5148
rect 16243 5110 16333 5148
rect 16371 5110 16461 5148
rect 16499 5110 16589 5148
rect 16627 5110 16717 5148
rect 16755 5110 16845 5148
rect 16883 5110 16973 5148
rect 17011 5110 17101 5148
rect 17139 5110 17229 5148
rect 17267 5110 17357 5148
rect 17395 5110 17485 5148
rect 17523 5110 17613 5148
rect 17651 5110 17741 5148
rect 17779 5110 17869 5148
rect 17907 5110 17997 5148
rect 18035 5110 18125 5148
rect 18163 5110 18253 5148
rect 18291 5110 18381 5148
rect 18419 5110 18509 5148
rect 18547 5110 18637 5148
rect 18675 5110 18765 5148
rect 18803 5110 18893 5148
rect 18931 5110 19021 5148
rect 19059 5110 19149 5148
rect 19187 5110 19277 5148
rect 19315 5110 19405 5148
rect 19443 5110 19533 5148
rect 19571 5110 19661 5148
rect 19699 5110 19789 5148
rect 19827 5110 19917 5148
rect 19955 5110 29365 5148
rect 29403 5110 29493 5148
rect 29531 5110 29621 5148
rect 29659 5110 29749 5148
rect 29787 5110 29877 5148
rect 29915 5110 30005 5148
rect 30043 5110 30133 5148
rect 30171 5110 30261 5148
rect 30299 5110 30389 5148
rect 30427 5110 30517 5148
rect 30555 5110 30645 5148
rect 30683 5110 30773 5148
rect 30811 5110 30901 5148
rect 30939 5110 31029 5148
rect 31067 5110 31157 5148
rect 31195 5110 31285 5148
rect 31323 5110 31413 5148
rect 31451 5110 31541 5148
rect 31579 5110 31669 5148
rect 31707 5110 31797 5148
rect 31835 5110 31925 5148
rect 31963 5110 32053 5148
rect 32091 5110 32181 5148
rect 32219 5110 32309 5148
rect 32347 5110 32437 5148
rect 32475 5110 32565 5148
rect 32603 5110 32693 5148
rect 32731 5110 32821 5148
rect 32859 5110 32949 5148
rect 32987 5110 33077 5148
rect 33115 5110 33205 5148
rect 33243 5110 33333 5148
rect 33371 5110 33461 5148
rect 33499 5110 33589 5148
rect 33627 5110 33717 5148
rect 33755 5110 33845 5148
rect 33883 5110 33973 5148
rect 34011 5110 34101 5148
rect 34139 5110 34229 5148
rect 34267 5110 34357 5148
rect 34395 5110 34485 5148
rect 34523 5110 34613 5148
rect 34651 5110 34741 5148
rect 34779 5110 34869 5148
rect 34907 5110 34997 5148
rect 35035 5110 35125 5148
rect 35163 5110 35253 5148
rect 35291 5110 35381 5148
rect 35419 5110 35509 5148
rect 35547 5110 35637 5148
rect 35675 5110 35765 5148
rect 35803 5110 35893 5148
rect 35931 5110 36021 5148
rect 36059 5110 36149 5148
rect 36187 5110 36277 5148
rect 36315 5110 36405 5148
rect 36443 5110 36533 5148
rect 36571 5110 36661 5148
rect 36699 5110 36789 5148
rect 36827 5110 36917 5148
rect 36955 5110 37045 5148
rect 37083 5110 37173 5148
rect 37211 5110 37301 5148
rect 37339 5110 37429 5148
rect 37467 5110 37557 5148
rect 37595 5110 37639 5148
rect 3448 5106 37639 5110
rect 675 4600 713 4678
rect 1587 4600 1625 4678
rect 2193 4600 2231 4678
rect 3121 4600 3159 4678
rect 3727 4600 3765 4678
rect 4333 4600 4371 4678
rect 4939 4600 4977 4678
rect 5672 4600 5710 4678
rect 6278 4600 6316 4678
rect 6884 4600 6922 4678
rect 7490 4600 7528 4678
rect 8096 4600 8134 4678
rect 8702 4600 8740 4678
rect 9308 4600 9346 4678
rect 9914 4600 9952 4678
rect 10646 4600 10684 4678
rect 11252 4600 11290 4678
rect 11858 4600 11896 4678
rect 12464 4600 12502 4678
rect 13070 4600 13108 4678
rect 13676 4600 13714 4678
rect 14282 4600 14320 4678
rect 14888 4600 14926 4678
rect 15494 4600 15532 4678
rect 16100 4600 16138 4678
rect 16706 4600 16744 4678
rect 17312 4600 17350 4678
rect 17918 4600 17956 4678
rect 18524 4600 18562 4678
rect 19130 4600 19168 4678
rect 19736 4600 19774 4678
rect 20468 4600 20506 4678
rect 21074 4600 21112 4678
rect 21680 4600 21718 4678
rect 22286 4600 22324 4678
rect 22892 4600 22930 4678
rect 23498 4600 23536 4678
rect 24104 4600 24142 4678
rect 24710 4600 24748 4678
rect 25316 4600 25354 4678
rect 25922 4600 25960 4678
rect 26528 4600 26566 4678
rect 27134 4600 27172 4678
rect 27740 4600 27778 4678
rect 28346 4600 28384 4678
rect 28952 4600 28990 4678
rect 29558 4600 29596 4678
rect 30164 4600 30202 4678
rect 30770 4600 30808 4678
rect 31376 4600 31414 4678
rect 31982 4600 32020 4678
rect 32588 4600 32626 4678
rect 33194 4600 33232 4678
rect 33800 4600 33838 4678
rect 34406 4600 34444 4678
rect 35012 4600 35050 4678
rect 35618 4600 35656 4678
rect 36224 4600 36262 4678
rect 36830 4600 36868 4678
rect 37436 4600 37474 4678
rect 38042 4600 38080 4678
rect 38648 4600 38686 4678
rect 39254 4600 39292 4678
rect -145 4282 -107 4360
rect 7850 3958 7894 4040
rect 669 3615 717 3729
rect 2069 3708 2109 3818
rect 4207 3754 4251 3854
rect 14766 3754 14810 3846
rect 29070 3542 29112 3632
rect -139 3440 -101 3518
rect 669 3122 707 3200
rect 1581 3122 1619 3200
rect 2187 3122 2225 3200
rect 3115 3122 3153 3200
rect 3721 3122 3759 3200
rect 4327 3122 4365 3200
rect 4933 3122 4971 3200
rect 5666 3122 5704 3200
rect 6272 3122 6310 3200
rect 6878 3122 6916 3200
rect 7484 3122 7522 3200
rect 8090 3122 8128 3200
rect 8696 3122 8734 3200
rect 9302 3122 9340 3200
rect 9908 3122 9946 3200
rect 10640 3122 10678 3200
rect 11246 3122 11284 3200
rect 11852 3122 11890 3200
rect 12458 3122 12496 3200
rect 13064 3122 13102 3200
rect 13670 3122 13708 3200
rect 14276 3122 14314 3200
rect 14882 3122 14920 3200
rect 15488 3122 15526 3200
rect 16094 3122 16132 3200
rect 16700 3122 16738 3200
rect 17306 3122 17344 3200
rect 17912 3122 17950 3200
rect 18518 3122 18556 3200
rect 19124 3122 19162 3200
rect 19730 3122 19768 3200
rect 20462 3122 20500 3200
rect 21068 3122 21106 3200
rect 21674 3122 21712 3200
rect 22280 3122 22318 3200
rect 22886 3122 22924 3200
rect 23492 3122 23530 3200
rect 24098 3122 24136 3200
rect 24704 3122 24742 3200
rect 25310 3122 25348 3200
rect 25916 3122 25954 3200
rect 26522 3122 26560 3200
rect 27128 3122 27166 3200
rect 27734 3122 27772 3200
rect 28340 3122 28378 3200
rect 28946 3122 28984 3200
rect 29552 3122 29590 3200
rect 30158 3122 30196 3200
rect 30764 3122 30802 3200
rect 31370 3122 31408 3200
rect 31976 3122 32014 3200
rect 32582 3122 32620 3200
rect 33188 3122 33226 3200
rect 33794 3122 33832 3200
rect 34400 3122 34438 3200
rect 35006 3122 35044 3200
rect 35612 3122 35650 3200
rect 36218 3122 36256 3200
rect 36824 3122 36862 3200
rect 37430 3122 37468 3200
rect 38036 3122 38074 3200
rect 38642 3122 38680 3200
rect 39248 3122 39286 3200
rect 675 1467 713 1545
rect 1587 1467 1625 1545
rect 2193 1467 2231 1545
rect 3121 1467 3159 1545
rect 3727 1467 3765 1545
rect 4333 1467 4371 1545
rect 4939 1467 4977 1545
rect 5672 1467 5710 1545
rect 6278 1467 6316 1545
rect 6884 1467 6922 1545
rect 7490 1467 7528 1545
rect 8096 1467 8134 1545
rect 8702 1467 8740 1545
rect 9308 1467 9346 1545
rect 9914 1467 9952 1545
rect 10646 1467 10684 1545
rect 11252 1467 11290 1545
rect 11858 1467 11896 1545
rect 12464 1467 12502 1545
rect 13070 1467 13108 1545
rect 13676 1467 13714 1545
rect 14282 1467 14320 1545
rect 14888 1467 14926 1545
rect 15494 1467 15532 1545
rect 16100 1467 16138 1545
rect 16706 1467 16744 1545
rect 17312 1467 17350 1545
rect 17918 1467 17956 1545
rect 18524 1467 18562 1545
rect 19130 1467 19168 1545
rect 19736 1467 19774 1545
rect 20468 1467 20506 1545
rect 21074 1467 21112 1545
rect 21680 1467 21718 1545
rect 22286 1467 22324 1545
rect 22892 1467 22930 1545
rect 23498 1467 23536 1545
rect 24104 1467 24142 1545
rect 24710 1467 24748 1545
rect 25316 1467 25354 1545
rect 25922 1467 25960 1545
rect 26528 1467 26566 1545
rect 27134 1467 27172 1545
rect 27740 1467 27778 1545
rect 28346 1467 28384 1545
rect 28952 1467 28990 1545
rect 29558 1467 29596 1545
rect 30164 1467 30202 1545
rect 30770 1467 30808 1545
rect 31376 1467 31414 1545
rect 31982 1467 32020 1545
rect 32588 1467 32626 1545
rect 33194 1467 33232 1545
rect 33800 1467 33838 1545
rect 34406 1467 34444 1545
rect 35012 1467 35050 1545
rect 35618 1467 35656 1545
rect 36224 1467 36262 1545
rect 36830 1467 36868 1545
rect 37436 1467 37474 1545
rect 38042 1467 38080 1545
rect 38648 1467 38686 1545
rect 39254 1467 39292 1545
rect -145 1149 -107 1227
rect 7850 825 7894 907
rect 669 482 717 596
rect 2069 575 2109 685
rect 4207 621 4251 721
rect 14766 621 14810 713
rect 29070 409 29112 499
rect -139 307 -101 385
rect 669 -11 707 67
rect 1581 -11 1619 67
rect 2187 -11 2225 67
rect 3115 -11 3153 67
rect 3721 -11 3759 67
rect 4327 -11 4365 67
rect 4933 -11 4971 67
rect 5666 -11 5704 67
rect 6272 -11 6310 67
rect 6878 -11 6916 67
rect 7484 -11 7522 67
rect 8090 -11 8128 67
rect 8696 -11 8734 67
rect 9302 -11 9340 67
rect 9908 -11 9946 67
rect 10640 -11 10678 67
rect 11246 -11 11284 67
rect 11852 -11 11890 67
rect 12458 -11 12496 67
rect 13064 -11 13102 67
rect 13670 -11 13708 67
rect 14276 -11 14314 67
rect 14882 -11 14920 67
rect 15488 -11 15526 67
rect 16094 -11 16132 67
rect 16700 -11 16738 67
rect 17306 -11 17344 67
rect 17912 -11 17950 67
rect 18518 -11 18556 67
rect 19124 -11 19162 67
rect 19730 -11 19768 67
rect 20462 -11 20500 67
rect 21068 -11 21106 67
rect 21674 -11 21712 67
rect 22280 -11 22318 67
rect 22886 -11 22924 67
rect 23492 -11 23530 67
rect 24098 -11 24136 67
rect 24704 -11 24742 67
rect 25310 -11 25348 67
rect 25916 -11 25954 67
rect 26522 -11 26560 67
rect 27128 -11 27166 67
rect 27734 -11 27772 67
rect 28340 -11 28378 67
rect 28946 -11 28984 67
rect 29552 -11 29590 67
rect 30158 -11 30196 67
rect 30764 -11 30802 67
rect 31370 -11 31408 67
rect 31976 -11 32014 67
rect 32582 -11 32620 67
rect 33188 -11 33226 67
rect 33794 -11 33832 67
rect 34400 -11 34438 67
rect 35006 -11 35044 67
rect 35612 -11 35650 67
rect 36218 -11 36256 67
rect 36824 -11 36862 67
rect 37430 -11 37468 67
rect 38036 -11 38074 67
rect 38642 -11 38680 67
rect 39248 -11 39286 67
<< nsubdiff >>
rect -363 5728 -109 5732
rect -363 5690 -319 5728
rect -281 5690 -191 5728
rect -153 5690 -109 5728
rect -363 5686 -109 5690
rect 437 5728 947 5732
rect 437 5690 481 5728
rect 519 5690 609 5728
rect 647 5690 737 5728
rect 775 5690 865 5728
rect 903 5690 947 5728
rect 437 5686 947 5690
rect 1317 5728 2467 5732
rect 1317 5690 1361 5728
rect 1399 5690 1489 5728
rect 1527 5690 1617 5728
rect 1655 5690 1745 5728
rect 1783 5690 1873 5728
rect 1911 5690 2001 5728
rect 2039 5690 2129 5728
rect 2167 5690 2257 5728
rect 2295 5690 2385 5728
rect 2423 5690 2467 5728
rect 1317 5686 2467 5690
rect 2936 5728 4598 5732
rect 2936 5690 2980 5728
rect 3018 5690 3108 5728
rect 3146 5690 3236 5728
rect 3274 5690 3364 5728
rect 3402 5690 3492 5728
rect 3530 5690 3620 5728
rect 3658 5690 3748 5728
rect 3786 5690 3876 5728
rect 3914 5690 4004 5728
rect 4042 5690 4132 5728
rect 4170 5690 4260 5728
rect 4298 5690 4388 5728
rect 4426 5690 4516 5728
rect 4554 5690 4598 5728
rect 2936 5686 4598 5690
rect 5429 5728 7603 5732
rect 5429 5690 5473 5728
rect 5511 5690 5601 5728
rect 5639 5690 5729 5728
rect 5767 5690 5857 5728
rect 5895 5690 5985 5728
rect 6023 5690 6113 5728
rect 6151 5690 6241 5728
rect 6279 5690 6369 5728
rect 6407 5690 6497 5728
rect 6535 5690 6625 5728
rect 6663 5690 6753 5728
rect 6791 5690 6881 5728
rect 6919 5690 7009 5728
rect 7047 5690 7137 5728
rect 7175 5690 7265 5728
rect 7303 5690 7393 5728
rect 7431 5690 7521 5728
rect 7559 5690 7603 5728
rect 5429 5686 7603 5690
rect 8013 5728 10187 5732
rect 8013 5690 8057 5728
rect 8095 5690 8185 5728
rect 8223 5690 8313 5728
rect 8351 5690 8441 5728
rect 8479 5690 8569 5728
rect 8607 5690 8697 5728
rect 8735 5690 8825 5728
rect 8863 5690 8953 5728
rect 8991 5690 9081 5728
rect 9119 5690 9209 5728
rect 9247 5690 9337 5728
rect 9375 5690 9465 5728
rect 9503 5690 9593 5728
rect 9631 5690 9721 5728
rect 9759 5690 9849 5728
rect 9887 5690 9977 5728
rect 10015 5690 10105 5728
rect 10143 5690 10187 5728
rect 8013 5686 10187 5690
rect 10516 5728 14738 5732
rect 10516 5690 10560 5728
rect 10598 5690 10688 5728
rect 10726 5690 10816 5728
rect 10854 5690 10944 5728
rect 10982 5690 11072 5728
rect 11110 5690 11200 5728
rect 11238 5690 11328 5728
rect 11366 5690 11456 5728
rect 11494 5690 11584 5728
rect 11622 5690 11712 5728
rect 11750 5690 11840 5728
rect 11878 5690 11968 5728
rect 12006 5690 12096 5728
rect 12134 5690 12224 5728
rect 12262 5690 12352 5728
rect 12390 5690 12480 5728
rect 12518 5690 12608 5728
rect 12646 5690 12736 5728
rect 12774 5690 12864 5728
rect 12902 5690 12992 5728
rect 13030 5690 13120 5728
rect 13158 5690 13248 5728
rect 13286 5690 13376 5728
rect 13414 5690 13504 5728
rect 13542 5690 13632 5728
rect 13670 5690 13760 5728
rect 13798 5690 13888 5728
rect 13926 5690 14016 5728
rect 14054 5690 14144 5728
rect 14182 5690 14272 5728
rect 14310 5690 14400 5728
rect 14438 5690 14528 5728
rect 14566 5690 14656 5728
rect 14694 5690 14738 5728
rect 10516 5686 14738 5690
rect 15777 5728 19999 5732
rect 15777 5690 15821 5728
rect 15859 5690 15949 5728
rect 15987 5690 16077 5728
rect 16115 5690 16205 5728
rect 16243 5690 16333 5728
rect 16371 5690 16461 5728
rect 16499 5690 16589 5728
rect 16627 5690 16717 5728
rect 16755 5690 16845 5728
rect 16883 5690 16973 5728
rect 17011 5690 17101 5728
rect 17139 5690 17229 5728
rect 17267 5690 17357 5728
rect 17395 5690 17485 5728
rect 17523 5690 17613 5728
rect 17651 5690 17741 5728
rect 17779 5690 17869 5728
rect 17907 5690 17997 5728
rect 18035 5690 18125 5728
rect 18163 5690 18253 5728
rect 18291 5690 18381 5728
rect 18419 5690 18509 5728
rect 18547 5690 18637 5728
rect 18675 5690 18765 5728
rect 18803 5690 18893 5728
rect 18931 5690 19021 5728
rect 19059 5690 19149 5728
rect 19187 5690 19277 5728
rect 19315 5690 19405 5728
rect 19443 5690 19533 5728
rect 19571 5690 19661 5728
rect 19699 5690 19789 5728
rect 19827 5690 19917 5728
rect 19955 5690 19999 5728
rect 15777 5686 19999 5690
rect 20353 5728 28671 5732
rect 20353 5690 20397 5728
rect 20435 5690 20525 5728
rect 20563 5690 20653 5728
rect 20691 5690 20781 5728
rect 20819 5690 20909 5728
rect 20947 5690 21037 5728
rect 21075 5690 21165 5728
rect 21203 5690 21293 5728
rect 21331 5690 21421 5728
rect 21459 5690 21549 5728
rect 21587 5690 21677 5728
rect 21715 5690 21805 5728
rect 21843 5690 21933 5728
rect 21971 5690 22061 5728
rect 22099 5690 22189 5728
rect 22227 5690 22317 5728
rect 22355 5690 22445 5728
rect 22483 5690 22573 5728
rect 22611 5690 22701 5728
rect 22739 5690 22829 5728
rect 22867 5690 22957 5728
rect 22995 5690 23085 5728
rect 23123 5690 23213 5728
rect 23251 5690 23341 5728
rect 23379 5690 23469 5728
rect 23507 5690 23597 5728
rect 23635 5690 23725 5728
rect 23763 5690 23853 5728
rect 23891 5690 23981 5728
rect 24019 5690 24109 5728
rect 24147 5690 24237 5728
rect 24275 5690 24365 5728
rect 24403 5690 24493 5728
rect 24531 5690 24621 5728
rect 24659 5690 24749 5728
rect 24787 5690 24877 5728
rect 24915 5690 25005 5728
rect 25043 5690 25133 5728
rect 25171 5690 25261 5728
rect 25299 5690 25389 5728
rect 25427 5690 25517 5728
rect 25555 5690 25645 5728
rect 25683 5690 25773 5728
rect 25811 5690 25901 5728
rect 25939 5690 26029 5728
rect 26067 5690 26157 5728
rect 26195 5690 26285 5728
rect 26323 5690 26413 5728
rect 26451 5690 26541 5728
rect 26579 5690 26669 5728
rect 26707 5690 26797 5728
rect 26835 5690 26925 5728
rect 26963 5690 27053 5728
rect 27091 5690 27181 5728
rect 27219 5690 27309 5728
rect 27347 5690 27437 5728
rect 27475 5690 27565 5728
rect 27603 5690 27693 5728
rect 27731 5690 27821 5728
rect 27859 5690 27949 5728
rect 27987 5690 28077 5728
rect 28115 5690 28205 5728
rect 28243 5690 28333 5728
rect 28371 5690 28461 5728
rect 28499 5690 28589 5728
rect 28627 5690 28671 5728
rect 20353 5686 28671 5690
rect 29321 5728 37639 5732
rect 29321 5690 29365 5728
rect 29403 5690 29493 5728
rect 29531 5690 29621 5728
rect 29659 5690 29749 5728
rect 29787 5690 29877 5728
rect 29915 5690 30005 5728
rect 30043 5690 30133 5728
rect 30171 5690 30261 5728
rect 30299 5690 30389 5728
rect 30427 5690 30517 5728
rect 30555 5690 30645 5728
rect 30683 5690 30773 5728
rect 30811 5690 30901 5728
rect 30939 5690 31029 5728
rect 31067 5690 31157 5728
rect 31195 5690 31285 5728
rect 31323 5690 31413 5728
rect 31451 5690 31541 5728
rect 31579 5690 31669 5728
rect 31707 5690 31797 5728
rect 31835 5690 31925 5728
rect 31963 5690 32053 5728
rect 32091 5690 32181 5728
rect 32219 5690 32309 5728
rect 32347 5690 32437 5728
rect 32475 5690 32565 5728
rect 32603 5690 32693 5728
rect 32731 5690 32821 5728
rect 32859 5690 32949 5728
rect 32987 5690 33077 5728
rect 33115 5690 33205 5728
rect 33243 5690 33333 5728
rect 33371 5690 33461 5728
rect 33499 5690 33589 5728
rect 33627 5690 33717 5728
rect 33755 5690 33845 5728
rect 33883 5690 33973 5728
rect 34011 5690 34101 5728
rect 34139 5690 34229 5728
rect 34267 5690 34357 5728
rect 34395 5690 34485 5728
rect 34523 5690 34613 5728
rect 34651 5690 34741 5728
rect 34779 5690 34869 5728
rect 34907 5690 34997 5728
rect 35035 5690 35125 5728
rect 35163 5690 35253 5728
rect 35291 5690 35381 5728
rect 35419 5690 35509 5728
rect 35547 5690 35637 5728
rect 35675 5690 35765 5728
rect 35803 5690 35893 5728
rect 35931 5690 36021 5728
rect 36059 5690 36149 5728
rect 36187 5690 36277 5728
rect 36315 5690 36405 5728
rect 36443 5690 36533 5728
rect 36571 5690 36661 5728
rect 36699 5690 36789 5728
rect 36827 5690 36917 5728
rect 36955 5690 37045 5728
rect 37083 5690 37173 5728
rect 37211 5690 37301 5728
rect 37339 5690 37429 5728
rect 37467 5690 37557 5728
rect 37595 5690 37639 5728
rect 29321 5686 37639 5690
<< psubdiffcont >>
rect -319 6270 -281 6308
rect -191 6270 -153 6308
rect 481 6270 519 6308
rect 609 6270 647 6308
rect 737 6270 775 6308
rect 1361 6270 1399 6308
rect 1489 6270 1527 6308
rect 1617 6270 1655 6308
rect 1745 6270 1783 6308
rect 1873 6270 1911 6308
rect 2980 6270 3018 6308
rect 3108 6270 3146 6308
rect 3236 6270 3274 6308
rect 3364 6270 3402 6308
rect 3492 6270 3530 6308
rect 3620 6270 3658 6308
rect 3748 6270 3786 6308
rect 3876 6270 3914 6308
rect 4004 6270 4042 6308
rect 5473 6270 5511 6308
rect 5601 6270 5639 6308
rect 5729 6270 5767 6308
rect 5857 6270 5895 6308
rect 5985 6270 6023 6308
rect 6113 6270 6151 6308
rect 6241 6270 6279 6308
rect 6369 6270 6407 6308
rect 6497 6270 6535 6308
rect 6625 6270 6663 6308
rect 6753 6270 6791 6308
rect 6881 6270 6919 6308
rect 7009 6270 7047 6308
rect 7137 6270 7175 6308
rect 7265 6270 7303 6308
rect 7393 6270 7431 6308
rect 7521 6270 7559 6308
rect 10560 6270 10598 6308
rect 10688 6270 10726 6308
rect 10816 6270 10854 6308
rect 10944 6270 10982 6308
rect 11072 6270 11110 6308
rect 11200 6270 11238 6308
rect 11328 6270 11366 6308
rect 11456 6270 11494 6308
rect 11584 6270 11622 6308
rect 11712 6270 11750 6308
rect 11840 6270 11878 6308
rect 11968 6270 12006 6308
rect 12096 6270 12134 6308
rect 12224 6270 12262 6308
rect 12352 6270 12390 6308
rect 12480 6270 12518 6308
rect 12608 6270 12646 6308
rect 12736 6270 12774 6308
rect 12864 6270 12902 6308
rect 12992 6270 13030 6308
rect 13120 6270 13158 6308
rect 13248 6270 13286 6308
rect 13376 6270 13414 6308
rect 13504 6270 13542 6308
rect 13632 6270 13670 6308
rect 13760 6270 13798 6308
rect 13888 6270 13926 6308
rect 14016 6270 14054 6308
rect 14144 6270 14182 6308
rect 14272 6270 14310 6308
rect 14400 6270 14438 6308
rect 14528 6270 14566 6308
rect 14656 6270 14694 6308
rect 20397 6270 20435 6308
rect 20525 6270 20563 6308
rect 20653 6270 20691 6308
rect 20781 6270 20819 6308
rect 20909 6270 20947 6308
rect 21037 6270 21075 6308
rect 21165 6270 21203 6308
rect 21293 6270 21331 6308
rect 21421 6270 21459 6308
rect 21549 6270 21587 6308
rect 21677 6270 21715 6308
rect 21805 6270 21843 6308
rect 21933 6270 21971 6308
rect 22061 6270 22099 6308
rect 22189 6270 22227 6308
rect 22317 6270 22355 6308
rect 22445 6270 22483 6308
rect 22573 6270 22611 6308
rect 22701 6270 22739 6308
rect 22829 6270 22867 6308
rect 22957 6270 22995 6308
rect 23085 6270 23123 6308
rect 23213 6270 23251 6308
rect 23341 6270 23379 6308
rect 23469 6270 23507 6308
rect 23597 6270 23635 6308
rect 23725 6270 23763 6308
rect 23853 6270 23891 6308
rect 23981 6270 24019 6308
rect 24109 6270 24147 6308
rect 24237 6270 24275 6308
rect 24365 6270 24403 6308
rect 24493 6270 24531 6308
rect 24621 6270 24659 6308
rect 24749 6270 24787 6308
rect 24877 6270 24915 6308
rect 25005 6270 25043 6308
rect 25133 6270 25171 6308
rect 25261 6270 25299 6308
rect 25389 6270 25427 6308
rect 25517 6270 25555 6308
rect 25645 6270 25683 6308
rect 25773 6270 25811 6308
rect 25901 6270 25939 6308
rect 26029 6270 26067 6308
rect 26157 6270 26195 6308
rect 26285 6270 26323 6308
rect 26413 6270 26451 6308
rect 26541 6270 26579 6308
rect 26669 6270 26707 6308
rect 26797 6270 26835 6308
rect 26925 6270 26963 6308
rect 27053 6270 27091 6308
rect 27181 6270 27219 6308
rect 27309 6270 27347 6308
rect 27437 6270 27475 6308
rect 27565 6270 27603 6308
rect 27693 6270 27731 6308
rect 27821 6270 27859 6308
rect 27949 6270 27987 6308
rect 28077 6270 28115 6308
rect 28205 6270 28243 6308
rect 28333 6270 28371 6308
rect 28461 6270 28499 6308
rect 28589 6270 28627 6308
rect -319 5110 -281 5148
rect -191 5110 -153 5148
rect 609 5110 647 5148
rect 737 5110 775 5148
rect 865 5110 903 5148
rect 1873 5110 1911 5148
rect 2001 5110 2039 5148
rect 2129 5110 2167 5148
rect 2257 5110 2295 5148
rect 2385 5110 2423 5148
rect 3492 5110 3530 5148
rect 3620 5110 3658 5148
rect 3748 5110 3786 5148
rect 3876 5110 3914 5148
rect 4004 5110 4042 5148
rect 4132 5110 4170 5148
rect 4260 5110 4298 5148
rect 4388 5110 4426 5148
rect 4516 5110 4554 5148
rect 8057 5110 8095 5148
rect 8185 5110 8223 5148
rect 8313 5110 8351 5148
rect 8441 5110 8479 5148
rect 8569 5110 8607 5148
rect 8697 5110 8735 5148
rect 8825 5110 8863 5148
rect 8953 5110 8991 5148
rect 9081 5110 9119 5148
rect 9209 5110 9247 5148
rect 9337 5110 9375 5148
rect 9465 5110 9503 5148
rect 9593 5110 9631 5148
rect 9721 5110 9759 5148
rect 9849 5110 9887 5148
rect 9977 5110 10015 5148
rect 10105 5110 10143 5148
rect 15821 5110 15859 5148
rect 15949 5110 15987 5148
rect 16077 5110 16115 5148
rect 16205 5110 16243 5148
rect 16333 5110 16371 5148
rect 16461 5110 16499 5148
rect 16589 5110 16627 5148
rect 16717 5110 16755 5148
rect 16845 5110 16883 5148
rect 16973 5110 17011 5148
rect 17101 5110 17139 5148
rect 17229 5110 17267 5148
rect 17357 5110 17395 5148
rect 17485 5110 17523 5148
rect 17613 5110 17651 5148
rect 17741 5110 17779 5148
rect 17869 5110 17907 5148
rect 17997 5110 18035 5148
rect 18125 5110 18163 5148
rect 18253 5110 18291 5148
rect 18381 5110 18419 5148
rect 18509 5110 18547 5148
rect 18637 5110 18675 5148
rect 18765 5110 18803 5148
rect 18893 5110 18931 5148
rect 19021 5110 19059 5148
rect 19149 5110 19187 5148
rect 19277 5110 19315 5148
rect 19405 5110 19443 5148
rect 19533 5110 19571 5148
rect 19661 5110 19699 5148
rect 19789 5110 19827 5148
rect 19917 5110 19955 5148
rect 29365 5110 29403 5148
rect 29493 5110 29531 5148
rect 29621 5110 29659 5148
rect 29749 5110 29787 5148
rect 29877 5110 29915 5148
rect 30005 5110 30043 5148
rect 30133 5110 30171 5148
rect 30261 5110 30299 5148
rect 30389 5110 30427 5148
rect 30517 5110 30555 5148
rect 30645 5110 30683 5148
rect 30773 5110 30811 5148
rect 30901 5110 30939 5148
rect 31029 5110 31067 5148
rect 31157 5110 31195 5148
rect 31285 5110 31323 5148
rect 31413 5110 31451 5148
rect 31541 5110 31579 5148
rect 31669 5110 31707 5148
rect 31797 5110 31835 5148
rect 31925 5110 31963 5148
rect 32053 5110 32091 5148
rect 32181 5110 32219 5148
rect 32309 5110 32347 5148
rect 32437 5110 32475 5148
rect 32565 5110 32603 5148
rect 32693 5110 32731 5148
rect 32821 5110 32859 5148
rect 32949 5110 32987 5148
rect 33077 5110 33115 5148
rect 33205 5110 33243 5148
rect 33333 5110 33371 5148
rect 33461 5110 33499 5148
rect 33589 5110 33627 5148
rect 33717 5110 33755 5148
rect 33845 5110 33883 5148
rect 33973 5110 34011 5148
rect 34101 5110 34139 5148
rect 34229 5110 34267 5148
rect 34357 5110 34395 5148
rect 34485 5110 34523 5148
rect 34613 5110 34651 5148
rect 34741 5110 34779 5148
rect 34869 5110 34907 5148
rect 34997 5110 35035 5148
rect 35125 5110 35163 5148
rect 35253 5110 35291 5148
rect 35381 5110 35419 5148
rect 35509 5110 35547 5148
rect 35637 5110 35675 5148
rect 35765 5110 35803 5148
rect 35893 5110 35931 5148
rect 36021 5110 36059 5148
rect 36149 5110 36187 5148
rect 36277 5110 36315 5148
rect 36405 5110 36443 5148
rect 36533 5110 36571 5148
rect 36661 5110 36699 5148
rect 36789 5110 36827 5148
rect 36917 5110 36955 5148
rect 37045 5110 37083 5148
rect 37173 5110 37211 5148
rect 37301 5110 37339 5148
rect 37429 5110 37467 5148
rect 37557 5110 37595 5148
<< nsubdiffcont >>
rect -319 5690 -281 5728
rect -191 5690 -153 5728
rect 481 5690 519 5728
rect 609 5690 647 5728
rect 737 5690 775 5728
rect 865 5690 903 5728
rect 1361 5690 1399 5728
rect 1489 5690 1527 5728
rect 1617 5690 1655 5728
rect 1745 5690 1783 5728
rect 1873 5690 1911 5728
rect 2001 5690 2039 5728
rect 2129 5690 2167 5728
rect 2257 5690 2295 5728
rect 2385 5690 2423 5728
rect 2980 5690 3018 5728
rect 3108 5690 3146 5728
rect 3236 5690 3274 5728
rect 3364 5690 3402 5728
rect 3492 5690 3530 5728
rect 3620 5690 3658 5728
rect 3748 5690 3786 5728
rect 3876 5690 3914 5728
rect 4004 5690 4042 5728
rect 4132 5690 4170 5728
rect 4260 5690 4298 5728
rect 4388 5690 4426 5728
rect 4516 5690 4554 5728
rect 5473 5690 5511 5728
rect 5601 5690 5639 5728
rect 5729 5690 5767 5728
rect 5857 5690 5895 5728
rect 5985 5690 6023 5728
rect 6113 5690 6151 5728
rect 6241 5690 6279 5728
rect 6369 5690 6407 5728
rect 6497 5690 6535 5728
rect 6625 5690 6663 5728
rect 6753 5690 6791 5728
rect 6881 5690 6919 5728
rect 7009 5690 7047 5728
rect 7137 5690 7175 5728
rect 7265 5690 7303 5728
rect 7393 5690 7431 5728
rect 7521 5690 7559 5728
rect 8057 5690 8095 5728
rect 8185 5690 8223 5728
rect 8313 5690 8351 5728
rect 8441 5690 8479 5728
rect 8569 5690 8607 5728
rect 8697 5690 8735 5728
rect 8825 5690 8863 5728
rect 8953 5690 8991 5728
rect 9081 5690 9119 5728
rect 9209 5690 9247 5728
rect 9337 5690 9375 5728
rect 9465 5690 9503 5728
rect 9593 5690 9631 5728
rect 9721 5690 9759 5728
rect 9849 5690 9887 5728
rect 9977 5690 10015 5728
rect 10105 5690 10143 5728
rect 10560 5690 10598 5728
rect 10688 5690 10726 5728
rect 10816 5690 10854 5728
rect 10944 5690 10982 5728
rect 11072 5690 11110 5728
rect 11200 5690 11238 5728
rect 11328 5690 11366 5728
rect 11456 5690 11494 5728
rect 11584 5690 11622 5728
rect 11712 5690 11750 5728
rect 11840 5690 11878 5728
rect 11968 5690 12006 5728
rect 12096 5690 12134 5728
rect 12224 5690 12262 5728
rect 12352 5690 12390 5728
rect 12480 5690 12518 5728
rect 12608 5690 12646 5728
rect 12736 5690 12774 5728
rect 12864 5690 12902 5728
rect 12992 5690 13030 5728
rect 13120 5690 13158 5728
rect 13248 5690 13286 5728
rect 13376 5690 13414 5728
rect 13504 5690 13542 5728
rect 13632 5690 13670 5728
rect 13760 5690 13798 5728
rect 13888 5690 13926 5728
rect 14016 5690 14054 5728
rect 14144 5690 14182 5728
rect 14272 5690 14310 5728
rect 14400 5690 14438 5728
rect 14528 5690 14566 5728
rect 14656 5690 14694 5728
rect 15821 5690 15859 5728
rect 15949 5690 15987 5728
rect 16077 5690 16115 5728
rect 16205 5690 16243 5728
rect 16333 5690 16371 5728
rect 16461 5690 16499 5728
rect 16589 5690 16627 5728
rect 16717 5690 16755 5728
rect 16845 5690 16883 5728
rect 16973 5690 17011 5728
rect 17101 5690 17139 5728
rect 17229 5690 17267 5728
rect 17357 5690 17395 5728
rect 17485 5690 17523 5728
rect 17613 5690 17651 5728
rect 17741 5690 17779 5728
rect 17869 5690 17907 5728
rect 17997 5690 18035 5728
rect 18125 5690 18163 5728
rect 18253 5690 18291 5728
rect 18381 5690 18419 5728
rect 18509 5690 18547 5728
rect 18637 5690 18675 5728
rect 18765 5690 18803 5728
rect 18893 5690 18931 5728
rect 19021 5690 19059 5728
rect 19149 5690 19187 5728
rect 19277 5690 19315 5728
rect 19405 5690 19443 5728
rect 19533 5690 19571 5728
rect 19661 5690 19699 5728
rect 19789 5690 19827 5728
rect 19917 5690 19955 5728
rect 20397 5690 20435 5728
rect 20525 5690 20563 5728
rect 20653 5690 20691 5728
rect 20781 5690 20819 5728
rect 20909 5690 20947 5728
rect 21037 5690 21075 5728
rect 21165 5690 21203 5728
rect 21293 5690 21331 5728
rect 21421 5690 21459 5728
rect 21549 5690 21587 5728
rect 21677 5690 21715 5728
rect 21805 5690 21843 5728
rect 21933 5690 21971 5728
rect 22061 5690 22099 5728
rect 22189 5690 22227 5728
rect 22317 5690 22355 5728
rect 22445 5690 22483 5728
rect 22573 5690 22611 5728
rect 22701 5690 22739 5728
rect 22829 5690 22867 5728
rect 22957 5690 22995 5728
rect 23085 5690 23123 5728
rect 23213 5690 23251 5728
rect 23341 5690 23379 5728
rect 23469 5690 23507 5728
rect 23597 5690 23635 5728
rect 23725 5690 23763 5728
rect 23853 5690 23891 5728
rect 23981 5690 24019 5728
rect 24109 5690 24147 5728
rect 24237 5690 24275 5728
rect 24365 5690 24403 5728
rect 24493 5690 24531 5728
rect 24621 5690 24659 5728
rect 24749 5690 24787 5728
rect 24877 5690 24915 5728
rect 25005 5690 25043 5728
rect 25133 5690 25171 5728
rect 25261 5690 25299 5728
rect 25389 5690 25427 5728
rect 25517 5690 25555 5728
rect 25645 5690 25683 5728
rect 25773 5690 25811 5728
rect 25901 5690 25939 5728
rect 26029 5690 26067 5728
rect 26157 5690 26195 5728
rect 26285 5690 26323 5728
rect 26413 5690 26451 5728
rect 26541 5690 26579 5728
rect 26669 5690 26707 5728
rect 26797 5690 26835 5728
rect 26925 5690 26963 5728
rect 27053 5690 27091 5728
rect 27181 5690 27219 5728
rect 27309 5690 27347 5728
rect 27437 5690 27475 5728
rect 27565 5690 27603 5728
rect 27693 5690 27731 5728
rect 27821 5690 27859 5728
rect 27949 5690 27987 5728
rect 28077 5690 28115 5728
rect 28205 5690 28243 5728
rect 28333 5690 28371 5728
rect 28461 5690 28499 5728
rect 28589 5690 28627 5728
rect 29365 5690 29403 5728
rect 29493 5690 29531 5728
rect 29621 5690 29659 5728
rect 29749 5690 29787 5728
rect 29877 5690 29915 5728
rect 30005 5690 30043 5728
rect 30133 5690 30171 5728
rect 30261 5690 30299 5728
rect 30389 5690 30427 5728
rect 30517 5690 30555 5728
rect 30645 5690 30683 5728
rect 30773 5690 30811 5728
rect 30901 5690 30939 5728
rect 31029 5690 31067 5728
rect 31157 5690 31195 5728
rect 31285 5690 31323 5728
rect 31413 5690 31451 5728
rect 31541 5690 31579 5728
rect 31669 5690 31707 5728
rect 31797 5690 31835 5728
rect 31925 5690 31963 5728
rect 32053 5690 32091 5728
rect 32181 5690 32219 5728
rect 32309 5690 32347 5728
rect 32437 5690 32475 5728
rect 32565 5690 32603 5728
rect 32693 5690 32731 5728
rect 32821 5690 32859 5728
rect 32949 5690 32987 5728
rect 33077 5690 33115 5728
rect 33205 5690 33243 5728
rect 33333 5690 33371 5728
rect 33461 5690 33499 5728
rect 33589 5690 33627 5728
rect 33717 5690 33755 5728
rect 33845 5690 33883 5728
rect 33973 5690 34011 5728
rect 34101 5690 34139 5728
rect 34229 5690 34267 5728
rect 34357 5690 34395 5728
rect 34485 5690 34523 5728
rect 34613 5690 34651 5728
rect 34741 5690 34779 5728
rect 34869 5690 34907 5728
rect 34997 5690 35035 5728
rect 35125 5690 35163 5728
rect 35253 5690 35291 5728
rect 35381 5690 35419 5728
rect 35509 5690 35547 5728
rect 35637 5690 35675 5728
rect 35765 5690 35803 5728
rect 35893 5690 35931 5728
rect 36021 5690 36059 5728
rect 36149 5690 36187 5728
rect 36277 5690 36315 5728
rect 36405 5690 36443 5728
rect 36533 5690 36571 5728
rect 36661 5690 36699 5728
rect 36789 5690 36827 5728
rect 36917 5690 36955 5728
rect 37045 5690 37083 5728
rect 37173 5690 37211 5728
rect 37301 5690 37339 5728
rect 37429 5690 37467 5728
rect 37557 5690 37595 5728
<< poly >>
rect -271 6212 -201 6238
rect 529 6212 599 6238
rect 657 6212 727 6238
rect 1409 6212 1479 6238
rect 1537 6212 1607 6238
rect 1665 6212 1735 6238
rect 1793 6212 1863 6238
rect 3028 6212 3098 6238
rect 3156 6212 3226 6238
rect 3284 6212 3354 6238
rect 3412 6212 3482 6238
rect 3540 6212 3610 6238
rect 3668 6212 3738 6238
rect 3796 6212 3866 6238
rect 3924 6212 3994 6238
rect 5521 6212 5591 6238
rect 5649 6212 5719 6238
rect 5777 6212 5847 6238
rect 5905 6212 5975 6238
rect 6033 6212 6103 6238
rect 6161 6212 6231 6238
rect 6289 6212 6359 6238
rect 6417 6212 6487 6238
rect 6545 6212 6615 6238
rect 6673 6212 6743 6238
rect 6801 6212 6871 6238
rect 6929 6212 6999 6238
rect 7057 6212 7127 6238
rect 7185 6212 7255 6238
rect 7313 6212 7383 6238
rect 7441 6212 7511 6238
rect 10608 6212 10678 6238
rect 10736 6212 10806 6238
rect 10864 6212 10934 6238
rect 10992 6212 11062 6238
rect 11120 6212 11190 6238
rect 11248 6212 11318 6238
rect 11376 6212 11446 6238
rect 11504 6212 11574 6238
rect 11632 6212 11702 6238
rect 11760 6212 11830 6238
rect 11888 6212 11958 6238
rect 12016 6212 12086 6238
rect 12144 6212 12214 6238
rect 12272 6212 12342 6238
rect 12400 6212 12470 6238
rect 12528 6212 12598 6238
rect 12656 6212 12726 6238
rect 12784 6212 12854 6238
rect 12912 6212 12982 6238
rect 13040 6212 13110 6238
rect 13168 6212 13238 6238
rect 13296 6212 13366 6238
rect 13424 6212 13494 6238
rect 13552 6212 13622 6238
rect 13680 6212 13750 6238
rect 13808 6212 13878 6238
rect 13936 6212 14006 6238
rect 14064 6212 14134 6238
rect 14192 6212 14262 6238
rect 14320 6212 14390 6238
rect 14448 6212 14518 6238
rect 14576 6212 14646 6238
rect 20445 6212 20515 6238
rect 20573 6212 20643 6238
rect 20701 6212 20771 6238
rect 20829 6212 20899 6238
rect 20957 6212 21027 6238
rect 21085 6212 21155 6238
rect 21213 6212 21283 6238
rect 21341 6212 21411 6238
rect 21469 6212 21539 6238
rect 21597 6212 21667 6238
rect 21725 6212 21795 6238
rect 21853 6212 21923 6238
rect 21981 6212 22051 6238
rect 22109 6212 22179 6238
rect 22237 6212 22307 6238
rect 22365 6212 22435 6238
rect 22493 6212 22563 6238
rect 22621 6212 22691 6238
rect 22749 6212 22819 6238
rect 22877 6212 22947 6238
rect 23005 6212 23075 6238
rect 23133 6212 23203 6238
rect 23261 6212 23331 6238
rect 23389 6212 23459 6238
rect 23517 6212 23587 6238
rect 23645 6212 23715 6238
rect 23773 6212 23843 6238
rect 23901 6212 23971 6238
rect 24029 6212 24099 6238
rect 24157 6212 24227 6238
rect 24285 6212 24355 6238
rect 24413 6212 24483 6238
rect 24541 6212 24611 6238
rect 24669 6212 24739 6238
rect 24797 6212 24867 6238
rect 24925 6212 24995 6238
rect 25053 6212 25123 6238
rect 25181 6212 25251 6238
rect 25309 6212 25379 6238
rect 25437 6212 25507 6238
rect 25565 6212 25635 6238
rect 25693 6212 25763 6238
rect 25821 6212 25891 6238
rect 25949 6212 26019 6238
rect 26077 6212 26147 6238
rect 26205 6212 26275 6238
rect 26333 6212 26403 6238
rect 26461 6212 26531 6238
rect 26589 6212 26659 6238
rect 26717 6212 26787 6238
rect 26845 6212 26915 6238
rect 26973 6212 27043 6238
rect 27101 6212 27171 6238
rect 27229 6212 27299 6238
rect 27357 6212 27427 6238
rect 27485 6212 27555 6238
rect 27613 6212 27683 6238
rect 27741 6212 27811 6238
rect 27869 6212 27939 6238
rect 27997 6212 28067 6238
rect 28125 6212 28195 6238
rect 28253 6212 28323 6238
rect 28381 6212 28451 6238
rect 28509 6212 28579 6238
rect 4107 6157 4173 6167
rect -271 6088 -201 6128
rect -301 6078 -201 6088
rect -301 6044 -285 6078
rect -251 6044 -201 6078
rect -301 6034 -201 6044
rect -271 5996 -201 6034
rect 529 6083 599 6128
rect 657 6088 727 6128
rect 657 6083 815 6088
rect 529 6078 815 6083
rect 529 6044 765 6078
rect 799 6044 815 6078
rect 529 6031 815 6044
rect 1409 6083 1479 6128
rect 1537 6083 1607 6128
rect 1665 6083 1735 6128
rect 1793 6083 1863 6128
rect 3028 6083 3098 6128
rect 3156 6083 3226 6128
rect 3284 6083 3354 6128
rect 3412 6083 3482 6128
rect 3540 6083 3610 6128
rect 3668 6083 3738 6128
rect 3796 6083 3866 6128
rect 3924 6113 3994 6128
rect 4107 6123 4123 6157
rect 4157 6123 4173 6157
rect 7684 6154 7750 6164
rect 4107 6119 4173 6123
rect 4106 6113 4173 6119
rect 3924 6110 4173 6113
rect 3924 6108 4139 6110
rect 3924 6083 4138 6108
rect 1409 6077 1987 6083
rect 1409 6067 2035 6077
rect 1409 6033 1985 6067
rect 2019 6033 2035 6067
rect 529 6013 727 6031
rect 529 5996 599 6013
rect 657 5996 727 6013
rect 1409 6020 2035 6033
rect 3028 6075 4138 6083
rect 5521 6083 5591 6128
rect 5649 6083 5719 6128
rect 5777 6083 5847 6128
rect 5905 6083 5975 6128
rect 6033 6083 6103 6128
rect 6161 6083 6231 6128
rect 6289 6083 6359 6128
rect 6417 6083 6487 6128
rect 6545 6083 6615 6128
rect 6673 6083 6743 6128
rect 6801 6083 6871 6128
rect 6929 6083 6999 6128
rect 7057 6083 7127 6128
rect 7185 6083 7255 6128
rect 7313 6083 7383 6128
rect 7441 6113 7511 6128
rect 7684 6120 7700 6154
rect 7734 6120 7750 6154
rect 7684 6115 7750 6120
rect 7681 6113 7750 6115
rect 7441 6107 7750 6113
rect 7441 6083 7722 6107
rect 1409 6014 1987 6020
rect 1409 6013 1863 6014
rect 1409 5996 1479 6013
rect 1537 5996 1607 6013
rect 1665 5996 1735 6013
rect 1793 5996 1863 6013
rect 3028 6013 3994 6075
rect 3028 5996 3098 6013
rect 3156 5996 3226 6013
rect 3284 5996 3354 6013
rect 3412 5996 3482 6013
rect 3540 5996 3610 6013
rect 3668 5996 3738 6013
rect 3796 5996 3866 6013
rect 3924 5996 3994 6013
rect 5521 6069 7722 6083
rect 10608 6093 10678 6128
rect 10736 6093 10806 6128
rect 10864 6093 10934 6128
rect 10992 6093 11062 6128
rect 11120 6093 11190 6128
rect 11248 6093 11318 6128
rect 11376 6093 11446 6128
rect 11504 6093 11574 6128
rect 11632 6093 11702 6128
rect 11760 6093 11830 6128
rect 11888 6093 11958 6128
rect 12016 6093 12086 6128
rect 12144 6093 12214 6128
rect 12272 6093 12342 6128
rect 12400 6093 12470 6128
rect 12528 6093 12598 6128
rect 12656 6093 12726 6128
rect 12784 6093 12854 6128
rect 12912 6093 12982 6128
rect 13040 6093 13110 6128
rect 13168 6093 13238 6128
rect 13296 6093 13366 6128
rect 13424 6093 13494 6128
rect 13552 6093 13622 6128
rect 13680 6093 13750 6128
rect 13808 6093 13878 6128
rect 13936 6093 14006 6128
rect 14064 6093 14134 6128
rect 14192 6093 14262 6128
rect 14320 6093 14390 6128
rect 14448 6093 14518 6128
rect 14576 6093 14646 6128
rect 10608 6092 14646 6093
rect 10608 6082 14765 6092
rect 5521 6013 7511 6069
rect 5521 5996 5591 6013
rect 5649 5996 5719 6013
rect 5777 5996 5847 6013
rect 5905 5996 5975 6013
rect 6033 5996 6103 6013
rect 6161 5996 6231 6013
rect 6289 5996 6359 6013
rect 6417 5996 6487 6013
rect 6545 5996 6615 6013
rect 6673 5996 6743 6013
rect 6801 5996 6871 6013
rect 6929 5996 6999 6013
rect 7057 5996 7127 6013
rect 7185 5996 7255 6013
rect 7313 5996 7383 6013
rect 7441 5996 7511 6013
rect 10608 6048 14715 6082
rect 14749 6048 14765 6082
rect 10608 6035 14765 6048
rect 20445 6083 20515 6128
rect 20573 6083 20643 6128
rect 20701 6083 20771 6128
rect 20829 6083 20899 6128
rect 20957 6083 21027 6128
rect 21085 6083 21155 6128
rect 21213 6083 21283 6128
rect 21341 6083 21411 6128
rect 21469 6083 21539 6128
rect 21597 6083 21667 6128
rect 21725 6083 21795 6128
rect 21853 6083 21923 6128
rect 21981 6083 22051 6128
rect 22109 6083 22179 6128
rect 22237 6083 22307 6128
rect 22365 6083 22435 6128
rect 22493 6083 22563 6128
rect 22621 6083 22691 6128
rect 22749 6083 22819 6128
rect 22877 6083 22947 6128
rect 23005 6083 23075 6128
rect 23133 6083 23203 6128
rect 23261 6083 23331 6128
rect 23389 6083 23459 6128
rect 23517 6083 23587 6128
rect 23645 6083 23715 6128
rect 23773 6083 23843 6128
rect 23901 6083 23971 6128
rect 24029 6083 24099 6128
rect 24157 6083 24227 6128
rect 24285 6083 24355 6128
rect 24413 6083 24483 6128
rect 24541 6083 24611 6128
rect 24669 6083 24739 6128
rect 24797 6083 24867 6128
rect 24925 6083 24995 6128
rect 25053 6083 25123 6128
rect 25181 6083 25251 6128
rect 25309 6083 25379 6128
rect 25437 6083 25507 6128
rect 25565 6083 25635 6128
rect 25693 6083 25763 6128
rect 25821 6083 25891 6128
rect 25949 6083 26019 6128
rect 26077 6083 26147 6128
rect 26205 6083 26275 6128
rect 26333 6083 26403 6128
rect 26461 6083 26531 6128
rect 26589 6083 26659 6128
rect 26717 6083 26787 6128
rect 26845 6083 26915 6128
rect 26973 6083 27043 6128
rect 27101 6083 27171 6128
rect 27229 6083 27299 6128
rect 27357 6083 27427 6128
rect 27485 6083 27555 6128
rect 27613 6083 27683 6128
rect 27741 6083 27811 6128
rect 27869 6083 27939 6128
rect 27997 6083 28067 6128
rect 28125 6083 28195 6128
rect 28253 6083 28323 6128
rect 28381 6083 28451 6128
rect 28509 6108 28579 6128
rect 28724 6108 28793 6115
rect 28509 6102 28793 6108
rect 28509 6083 28743 6102
rect 20445 6068 28743 6083
rect 28777 6068 28793 6102
rect 20445 6058 28793 6068
rect 10608 6013 14646 6035
rect 10608 5996 10678 6013
rect 10736 5996 10806 6013
rect 10864 5996 10934 6013
rect 10992 5996 11062 6013
rect 11120 5996 11190 6013
rect 11248 5996 11318 6013
rect 11376 5996 11446 6013
rect 11504 5996 11574 6013
rect 11632 5996 11702 6013
rect 11760 5996 11830 6013
rect 11888 5996 11958 6013
rect 12016 5996 12086 6013
rect 12144 5996 12214 6013
rect 12272 5996 12342 6013
rect 12400 5996 12470 6013
rect 12528 5996 12598 6013
rect 12656 5996 12726 6013
rect 12784 5996 12854 6013
rect 12912 5996 12982 6013
rect 13040 5996 13110 6013
rect 13168 5996 13238 6013
rect 13296 5996 13366 6013
rect 13424 5996 13494 6013
rect 13552 5996 13622 6013
rect 13680 5996 13750 6013
rect 13808 5996 13878 6013
rect 13936 5996 14006 6013
rect 14064 5996 14134 6013
rect 14192 5996 14262 6013
rect 14320 5996 14390 6013
rect 14448 5996 14518 6013
rect 14576 5996 14646 6013
rect 20445 6013 28579 6058
rect 20445 5996 20515 6013
rect 20573 5996 20643 6013
rect 20701 5996 20771 6013
rect 20829 5996 20899 6013
rect 20957 5996 21027 6013
rect 21085 5996 21155 6013
rect 21213 5996 21283 6013
rect 21341 5996 21411 6013
rect 21469 5996 21539 6013
rect 21597 5996 21667 6013
rect 21725 5996 21795 6013
rect 21853 5996 21923 6013
rect 21981 5996 22051 6013
rect 22109 5996 22179 6013
rect 22237 5996 22307 6013
rect 22365 5996 22435 6013
rect 22493 5996 22563 6013
rect 22621 5996 22691 6013
rect 22749 5996 22819 6013
rect 22877 5996 22947 6013
rect 23005 5996 23075 6013
rect 23133 5996 23203 6013
rect 23261 5996 23331 6013
rect 23389 5996 23459 6013
rect 23517 5996 23587 6013
rect 23645 5996 23715 6013
rect 23773 5996 23843 6013
rect 23901 5996 23971 6013
rect 24029 5996 24099 6013
rect 24157 5996 24227 6013
rect 24285 5996 24355 6013
rect 24413 5996 24483 6013
rect 24541 5996 24611 6013
rect 24669 5996 24739 6013
rect 24797 5996 24867 6013
rect 24925 5996 24995 6013
rect 25053 5996 25123 6013
rect 25181 5996 25251 6013
rect 25309 5996 25379 6013
rect 25437 5996 25507 6013
rect 25565 5996 25635 6013
rect 25693 5996 25763 6013
rect 25821 5996 25891 6013
rect 25949 5996 26019 6013
rect 26077 5996 26147 6013
rect 26205 5996 26275 6013
rect 26333 5996 26403 6013
rect 26461 5996 26531 6013
rect 26589 5996 26659 6013
rect 26717 5996 26787 6013
rect 26845 5996 26915 6013
rect 26973 5996 27043 6013
rect 27101 5996 27171 6013
rect 27229 5996 27299 6013
rect 27357 5996 27427 6013
rect 27485 5996 27555 6013
rect 27613 5996 27683 6013
rect 27741 5996 27811 6013
rect 27869 5996 27939 6013
rect 27997 5996 28067 6013
rect 28125 5996 28195 6013
rect 28253 5996 28323 6013
rect 28381 5996 28451 6013
rect 28509 5996 28579 6013
rect -271 5797 -201 5828
rect 529 5797 599 5828
rect 657 5797 727 5828
rect 1409 5797 1479 5828
rect 1537 5797 1607 5828
rect 1665 5797 1735 5828
rect 1793 5797 1863 5828
rect 3028 5797 3098 5828
rect 3156 5797 3226 5828
rect 3284 5797 3354 5828
rect 3412 5797 3482 5828
rect 3540 5797 3610 5828
rect 3668 5797 3738 5828
rect 3796 5797 3866 5828
rect 3924 5797 3994 5828
rect 5521 5797 5591 5828
rect 5649 5797 5719 5828
rect 5777 5797 5847 5828
rect 5905 5797 5975 5828
rect 6033 5797 6103 5828
rect 6161 5797 6231 5828
rect 6289 5797 6359 5828
rect 6417 5797 6487 5828
rect 6545 5797 6615 5828
rect 6673 5797 6743 5828
rect 6801 5797 6871 5828
rect 6929 5797 6999 5828
rect 7057 5797 7127 5828
rect 7185 5797 7255 5828
rect 7313 5797 7383 5828
rect 7441 5797 7511 5828
rect 10608 5797 10678 5828
rect 10736 5797 10806 5828
rect 10864 5797 10934 5828
rect 10992 5797 11062 5828
rect 11120 5797 11190 5828
rect 11248 5797 11318 5828
rect 11376 5797 11446 5828
rect 11504 5797 11574 5828
rect 11632 5797 11702 5828
rect 11760 5797 11830 5828
rect 11888 5797 11958 5828
rect 12016 5797 12086 5828
rect 12144 5797 12214 5828
rect 12272 5797 12342 5828
rect 12400 5797 12470 5828
rect 12528 5797 12598 5828
rect 12656 5797 12726 5828
rect 12784 5797 12854 5828
rect 12912 5797 12982 5828
rect 13040 5797 13110 5828
rect 13168 5797 13238 5828
rect 13296 5797 13366 5828
rect 13424 5797 13494 5828
rect 13552 5797 13622 5828
rect 13680 5797 13750 5828
rect 13808 5797 13878 5828
rect 13936 5797 14006 5828
rect 14064 5797 14134 5828
rect 14192 5797 14262 5828
rect 14320 5797 14390 5828
rect 14448 5797 14518 5828
rect 14576 5797 14646 5828
rect 20445 5797 20515 5828
rect 20573 5797 20643 5828
rect 20701 5797 20771 5828
rect 20829 5797 20899 5828
rect 20957 5797 21027 5828
rect 21085 5797 21155 5828
rect 21213 5797 21283 5828
rect 21341 5797 21411 5828
rect 21469 5797 21539 5828
rect 21597 5797 21667 5828
rect 21725 5797 21795 5828
rect 21853 5797 21923 5828
rect 21981 5797 22051 5828
rect 22109 5797 22179 5828
rect 22237 5797 22307 5828
rect 22365 5797 22435 5828
rect 22493 5797 22563 5828
rect 22621 5797 22691 5828
rect 22749 5797 22819 5828
rect 22877 5797 22947 5828
rect 23005 5797 23075 5828
rect 23133 5797 23203 5828
rect 23261 5797 23331 5828
rect 23389 5797 23459 5828
rect 23517 5797 23587 5828
rect 23645 5797 23715 5828
rect 23773 5797 23843 5828
rect 23901 5797 23971 5828
rect 24029 5797 24099 5828
rect 24157 5797 24227 5828
rect 24285 5797 24355 5828
rect 24413 5797 24483 5828
rect 24541 5797 24611 5828
rect 24669 5797 24739 5828
rect 24797 5797 24867 5828
rect 24925 5797 24995 5828
rect 25053 5797 25123 5828
rect 25181 5797 25251 5828
rect 25309 5797 25379 5828
rect 25437 5797 25507 5828
rect 25565 5797 25635 5828
rect 25693 5797 25763 5828
rect 25821 5797 25891 5828
rect 25949 5797 26019 5828
rect 26077 5797 26147 5828
rect 26205 5797 26275 5828
rect 26333 5797 26403 5828
rect 26461 5797 26531 5828
rect 26589 5797 26659 5828
rect 26717 5797 26787 5828
rect 26845 5797 26915 5828
rect 26973 5797 27043 5828
rect 27101 5797 27171 5828
rect 27229 5797 27299 5828
rect 27357 5797 27427 5828
rect 27485 5797 27555 5828
rect 27613 5797 27683 5828
rect 27741 5797 27811 5828
rect 27869 5797 27939 5828
rect 27997 5797 28067 5828
rect 28125 5797 28195 5828
rect 28253 5797 28323 5828
rect 28381 5797 28451 5828
rect 28509 5797 28579 5828
rect -271 5590 -201 5621
rect 657 5590 727 5621
rect 785 5590 855 5621
rect 1921 5590 1991 5621
rect 2049 5590 2119 5621
rect 2177 5590 2247 5621
rect 2305 5590 2375 5621
rect 3540 5590 3610 5621
rect 3668 5590 3738 5621
rect 3796 5590 3866 5621
rect 3924 5590 3994 5621
rect 4052 5590 4122 5621
rect 4180 5590 4250 5621
rect 4308 5590 4378 5621
rect 4436 5590 4506 5621
rect 8105 5590 8175 5621
rect 8233 5590 8303 5621
rect 8361 5590 8431 5621
rect 8489 5590 8559 5621
rect 8617 5590 8687 5621
rect 8745 5590 8815 5621
rect 8873 5590 8943 5621
rect 9001 5590 9071 5621
rect 9129 5590 9199 5621
rect 9257 5590 9327 5621
rect 9385 5590 9455 5621
rect 9513 5590 9583 5621
rect 9641 5590 9711 5621
rect 9769 5590 9839 5621
rect 9897 5590 9967 5621
rect 10025 5590 10095 5621
rect 15869 5590 15939 5621
rect 15997 5590 16067 5621
rect 16125 5590 16195 5621
rect 16253 5590 16323 5621
rect 16381 5590 16451 5621
rect 16509 5590 16579 5621
rect 16637 5590 16707 5621
rect 16765 5590 16835 5621
rect 16893 5590 16963 5621
rect 17021 5590 17091 5621
rect 17149 5590 17219 5621
rect 17277 5590 17347 5621
rect 17405 5590 17475 5621
rect 17533 5590 17603 5621
rect 17661 5590 17731 5621
rect 17789 5590 17859 5621
rect 17917 5590 17987 5621
rect 18045 5590 18115 5621
rect 18173 5590 18243 5621
rect 18301 5590 18371 5621
rect 18429 5590 18499 5621
rect 18557 5590 18627 5621
rect 18685 5590 18755 5621
rect 18813 5590 18883 5621
rect 18941 5590 19011 5621
rect 19069 5590 19139 5621
rect 19197 5590 19267 5621
rect 19325 5590 19395 5621
rect 19453 5590 19523 5621
rect 19581 5590 19651 5621
rect 19709 5590 19779 5621
rect 19837 5590 19907 5621
rect 29413 5590 29483 5621
rect 29541 5590 29611 5621
rect 29669 5590 29739 5621
rect 29797 5590 29867 5621
rect 29925 5590 29995 5621
rect 30053 5590 30123 5621
rect 30181 5590 30251 5621
rect 30309 5590 30379 5621
rect 30437 5590 30507 5621
rect 30565 5590 30635 5621
rect 30693 5590 30763 5621
rect 30821 5590 30891 5621
rect 30949 5590 31019 5621
rect 31077 5590 31147 5621
rect 31205 5590 31275 5621
rect 31333 5590 31403 5621
rect 31461 5590 31531 5621
rect 31589 5590 31659 5621
rect 31717 5590 31787 5621
rect 31845 5590 31915 5621
rect 31973 5590 32043 5621
rect 32101 5590 32171 5621
rect 32229 5590 32299 5621
rect 32357 5590 32427 5621
rect 32485 5590 32555 5621
rect 32613 5590 32683 5621
rect 32741 5590 32811 5621
rect 32869 5590 32939 5621
rect 32997 5590 33067 5621
rect 33125 5590 33195 5621
rect 33253 5590 33323 5621
rect 33381 5590 33451 5621
rect 33509 5590 33579 5621
rect 33637 5590 33707 5621
rect 33765 5590 33835 5621
rect 33893 5590 33963 5621
rect 34021 5590 34091 5621
rect 34149 5590 34219 5621
rect 34277 5590 34347 5621
rect 34405 5590 34475 5621
rect 34533 5590 34603 5621
rect 34661 5590 34731 5621
rect 34789 5590 34859 5621
rect 34917 5590 34987 5621
rect 35045 5590 35115 5621
rect 35173 5590 35243 5621
rect 35301 5590 35371 5621
rect 35429 5590 35499 5621
rect 35557 5590 35627 5621
rect 35685 5590 35755 5621
rect 35813 5590 35883 5621
rect 35941 5590 36011 5621
rect 36069 5590 36139 5621
rect 36197 5590 36267 5621
rect 36325 5590 36395 5621
rect 36453 5590 36523 5621
rect 36581 5590 36651 5621
rect 36709 5590 36779 5621
rect 36837 5590 36907 5621
rect 36965 5590 37035 5621
rect 37093 5590 37163 5621
rect 37221 5590 37291 5621
rect 37349 5590 37419 5621
rect 37477 5590 37547 5621
rect 961 5435 1030 5445
rect -271 5382 -201 5422
rect -388 5372 -201 5382
rect -388 5338 -372 5372
rect -338 5338 -201 5372
rect -388 5328 -201 5338
rect -271 5290 -201 5328
rect 657 5405 727 5422
rect 785 5405 855 5422
rect 961 5417 977 5435
rect 657 5402 855 5405
rect 958 5402 977 5417
rect 657 5401 977 5402
rect 1011 5401 1030 5435
rect 2490 5435 2556 5445
rect 657 5391 1030 5401
rect 1921 5405 1991 5422
rect 2049 5405 2119 5422
rect 2177 5405 2247 5422
rect 2305 5406 2375 5422
rect 2490 5406 2506 5435
rect 2305 5405 2506 5406
rect 1921 5401 2506 5405
rect 2540 5401 2556 5435
rect 4661 5444 4727 5454
rect 657 5372 988 5391
rect 1921 5388 2556 5401
rect 3540 5405 3610 5422
rect 3668 5405 3738 5422
rect 3796 5405 3866 5422
rect 3924 5405 3994 5422
rect 4052 5405 4122 5422
rect 4180 5405 4250 5422
rect 4308 5405 4378 5422
rect 4436 5405 4506 5422
rect 4661 5410 4677 5444
rect 4711 5410 4727 5444
rect 4661 5405 4727 5410
rect 3540 5397 4727 5405
rect 7919 5429 7985 5439
rect 657 5335 855 5372
rect 657 5290 727 5335
rect 785 5290 855 5335
rect 1921 5361 2520 5388
rect 3540 5364 4698 5397
rect 7919 5395 7935 5429
rect 7969 5414 7985 5429
rect 7969 5407 7988 5414
rect 8105 5407 8175 5422
rect 7969 5405 8175 5407
rect 8233 5405 8303 5422
rect 8361 5405 8431 5422
rect 8489 5405 8559 5422
rect 8617 5405 8687 5422
rect 8745 5405 8815 5422
rect 8873 5405 8943 5422
rect 9001 5405 9071 5422
rect 9129 5405 9199 5422
rect 9257 5405 9327 5422
rect 9385 5405 9455 5422
rect 9513 5405 9583 5422
rect 9641 5405 9711 5422
rect 9769 5405 9839 5422
rect 9897 5405 9967 5422
rect 10025 5405 10095 5422
rect 7969 5395 10095 5405
rect 7919 5382 10095 5395
rect 1921 5335 2375 5361
rect 1921 5290 1991 5335
rect 2049 5290 2119 5335
rect 2177 5290 2247 5335
rect 2305 5290 2375 5335
rect 3540 5335 4506 5364
rect 7962 5363 10095 5382
rect 3540 5290 3610 5335
rect 3668 5290 3738 5335
rect 3796 5290 3866 5335
rect 3924 5290 3994 5335
rect 4052 5290 4122 5335
rect 4180 5290 4250 5335
rect 4308 5290 4378 5335
rect 4436 5290 4506 5335
rect 8105 5335 10095 5363
rect 15688 5407 15757 5408
rect 15869 5407 15939 5422
rect 15688 5405 15939 5407
rect 15997 5405 16067 5422
rect 16125 5405 16195 5422
rect 16253 5405 16323 5422
rect 16381 5405 16451 5422
rect 16509 5405 16579 5422
rect 16637 5405 16707 5422
rect 16765 5405 16835 5422
rect 16893 5405 16963 5422
rect 17021 5405 17091 5422
rect 17149 5405 17219 5422
rect 17277 5405 17347 5422
rect 17405 5405 17475 5422
rect 17533 5405 17603 5422
rect 17661 5405 17731 5422
rect 17789 5405 17859 5422
rect 17917 5405 17987 5422
rect 18045 5405 18115 5422
rect 18173 5405 18243 5422
rect 18301 5405 18371 5422
rect 18429 5405 18499 5422
rect 18557 5405 18627 5422
rect 18685 5405 18755 5422
rect 18813 5405 18883 5422
rect 18941 5405 19011 5422
rect 19069 5405 19139 5422
rect 19197 5405 19267 5422
rect 19325 5405 19395 5422
rect 19453 5405 19523 5422
rect 19581 5405 19651 5422
rect 19709 5405 19779 5422
rect 19837 5405 19907 5422
rect 15688 5398 19907 5405
rect 15688 5364 15704 5398
rect 15738 5364 19907 5398
rect 15688 5351 19907 5364
rect 8105 5290 8175 5335
rect 8233 5290 8303 5335
rect 8361 5290 8431 5335
rect 8489 5290 8559 5335
rect 8617 5290 8687 5335
rect 8745 5290 8815 5335
rect 8873 5290 8943 5335
rect 9001 5290 9071 5335
rect 9129 5290 9199 5335
rect 9257 5290 9327 5335
rect 9385 5290 9455 5335
rect 9513 5290 9583 5335
rect 9641 5290 9711 5335
rect 9769 5290 9839 5335
rect 9897 5290 9967 5335
rect 10025 5290 10095 5335
rect 15869 5335 19907 5351
rect 15869 5290 15939 5335
rect 15997 5290 16067 5335
rect 16125 5290 16195 5335
rect 16253 5290 16323 5335
rect 16381 5290 16451 5335
rect 16509 5290 16579 5335
rect 16637 5290 16707 5335
rect 16765 5290 16835 5335
rect 16893 5290 16963 5335
rect 17021 5290 17091 5335
rect 17149 5290 17219 5335
rect 17277 5290 17347 5335
rect 17405 5290 17475 5335
rect 17533 5290 17603 5335
rect 17661 5290 17731 5335
rect 17789 5290 17859 5335
rect 17917 5290 17987 5335
rect 18045 5290 18115 5335
rect 18173 5290 18243 5335
rect 18301 5290 18371 5335
rect 18429 5290 18499 5335
rect 18557 5290 18627 5335
rect 18685 5290 18755 5335
rect 18813 5290 18883 5335
rect 18941 5290 19011 5335
rect 19069 5290 19139 5335
rect 19197 5290 19267 5335
rect 19325 5290 19395 5335
rect 19453 5290 19523 5335
rect 19581 5290 19651 5335
rect 19709 5290 19779 5335
rect 19837 5290 19907 5335
rect 29413 5405 29483 5422
rect 29541 5405 29611 5422
rect 29669 5405 29739 5422
rect 29797 5405 29867 5422
rect 29925 5405 29995 5422
rect 30053 5405 30123 5422
rect 30181 5405 30251 5422
rect 30309 5405 30379 5422
rect 30437 5405 30507 5422
rect 30565 5405 30635 5422
rect 30693 5405 30763 5422
rect 30821 5405 30891 5422
rect 30949 5405 31019 5422
rect 31077 5405 31147 5422
rect 31205 5405 31275 5422
rect 31333 5405 31403 5422
rect 31461 5405 31531 5422
rect 31589 5405 31659 5422
rect 31717 5405 31787 5422
rect 31845 5405 31915 5422
rect 31973 5405 32043 5422
rect 32101 5405 32171 5422
rect 32229 5405 32299 5422
rect 32357 5405 32427 5422
rect 32485 5405 32555 5422
rect 32613 5405 32683 5422
rect 32741 5405 32811 5422
rect 32869 5405 32939 5422
rect 32997 5405 33067 5422
rect 33125 5405 33195 5422
rect 33253 5405 33323 5422
rect 33381 5405 33451 5422
rect 33509 5405 33579 5422
rect 33637 5405 33707 5422
rect 33765 5405 33835 5422
rect 33893 5405 33963 5422
rect 34021 5405 34091 5422
rect 34149 5405 34219 5422
rect 34277 5405 34347 5422
rect 34405 5405 34475 5422
rect 34533 5405 34603 5422
rect 34661 5405 34731 5422
rect 34789 5405 34859 5422
rect 34917 5405 34987 5422
rect 35045 5405 35115 5422
rect 35173 5405 35243 5422
rect 35301 5405 35371 5422
rect 35429 5405 35499 5422
rect 35557 5405 35627 5422
rect 35685 5405 35755 5422
rect 35813 5405 35883 5422
rect 35941 5405 36011 5422
rect 36069 5405 36139 5422
rect 36197 5405 36267 5422
rect 36325 5405 36395 5422
rect 36453 5405 36523 5422
rect 36581 5405 36651 5422
rect 36709 5405 36779 5422
rect 36837 5405 36907 5422
rect 36965 5405 37035 5422
rect 37093 5405 37163 5422
rect 37221 5405 37291 5422
rect 37349 5405 37419 5422
rect 37477 5405 37547 5422
rect 29413 5335 37547 5405
rect 29413 5290 29483 5335
rect 29541 5290 29611 5335
rect 29669 5290 29739 5335
rect 29797 5290 29867 5335
rect 29925 5290 29995 5335
rect 30053 5290 30123 5335
rect 30181 5290 30251 5335
rect 30309 5290 30379 5335
rect 30437 5290 30507 5335
rect 30565 5290 30635 5335
rect 30693 5290 30763 5335
rect 30821 5290 30891 5335
rect 30949 5290 31019 5335
rect 31077 5290 31147 5335
rect 31205 5290 31275 5335
rect 31333 5290 31403 5335
rect 31461 5290 31531 5335
rect 31589 5290 31659 5335
rect 31717 5290 31787 5335
rect 31845 5290 31915 5335
rect 31973 5290 32043 5335
rect 32101 5290 32171 5335
rect 32229 5290 32299 5335
rect 32357 5290 32427 5335
rect 32485 5290 32555 5335
rect 32613 5290 32683 5335
rect 32741 5290 32811 5335
rect 32869 5290 32939 5335
rect 32997 5290 33067 5335
rect 33125 5290 33195 5335
rect 33253 5290 33323 5335
rect 33381 5290 33451 5335
rect 33509 5290 33579 5335
rect 33637 5290 33707 5335
rect 33765 5290 33835 5335
rect 33893 5290 33963 5335
rect 34021 5290 34091 5335
rect 34149 5290 34219 5335
rect 34277 5290 34347 5335
rect 34405 5290 34475 5335
rect 34533 5290 34603 5335
rect 34661 5290 34731 5335
rect 34789 5290 34859 5335
rect 34917 5290 34987 5335
rect 35045 5290 35115 5335
rect 35173 5290 35243 5335
rect 35301 5290 35371 5335
rect 35429 5290 35499 5335
rect 35557 5290 35627 5335
rect 35685 5290 35755 5335
rect 35813 5290 35883 5335
rect 35941 5290 36011 5335
rect 36069 5290 36139 5335
rect 36197 5290 36267 5335
rect 36325 5290 36395 5335
rect 36453 5290 36523 5335
rect 36581 5290 36651 5335
rect 36709 5290 36779 5335
rect 36837 5290 36907 5335
rect 36965 5290 37035 5335
rect 37093 5290 37163 5335
rect 37221 5290 37291 5335
rect 37349 5290 37419 5335
rect 37477 5290 37547 5335
rect -271 5180 -201 5206
rect 657 5180 727 5206
rect 785 5180 855 5206
rect 1921 5180 1991 5206
rect 2049 5180 2119 5206
rect 2177 5180 2247 5206
rect 2305 5180 2375 5206
rect 3540 5180 3610 5206
rect 3668 5180 3738 5206
rect 3796 5180 3866 5206
rect 3924 5180 3994 5206
rect 4052 5180 4122 5206
rect 4180 5180 4250 5206
rect 4308 5180 4378 5206
rect 4436 5180 4506 5206
rect 8105 5180 8175 5206
rect 8233 5180 8303 5206
rect 8361 5180 8431 5206
rect 8489 5180 8559 5206
rect 8617 5180 8687 5206
rect 8745 5180 8815 5206
rect 8873 5180 8943 5206
rect 9001 5180 9071 5206
rect 9129 5180 9199 5206
rect 9257 5180 9327 5206
rect 9385 5180 9455 5206
rect 9513 5180 9583 5206
rect 9641 5180 9711 5206
rect 9769 5180 9839 5206
rect 9897 5180 9967 5206
rect 10025 5180 10095 5206
rect 15869 5180 15939 5206
rect 15997 5180 16067 5206
rect 16125 5180 16195 5206
rect 16253 5180 16323 5206
rect 16381 5180 16451 5206
rect 16509 5180 16579 5206
rect 16637 5180 16707 5206
rect 16765 5180 16835 5206
rect 16893 5180 16963 5206
rect 17021 5180 17091 5206
rect 17149 5180 17219 5206
rect 17277 5180 17347 5206
rect 17405 5180 17475 5206
rect 17533 5180 17603 5206
rect 17661 5180 17731 5206
rect 17789 5180 17859 5206
rect 17917 5180 17987 5206
rect 18045 5180 18115 5206
rect 18173 5180 18243 5206
rect 18301 5180 18371 5206
rect 18429 5180 18499 5206
rect 18557 5180 18627 5206
rect 18685 5180 18755 5206
rect 18813 5180 18883 5206
rect 18941 5180 19011 5206
rect 19069 5180 19139 5206
rect 19197 5180 19267 5206
rect 19325 5180 19395 5206
rect 19453 5180 19523 5206
rect 19581 5180 19651 5206
rect 19709 5180 19779 5206
rect 19837 5180 19907 5206
rect 29413 5180 29483 5206
rect 29541 5180 29611 5206
rect 29669 5180 29739 5206
rect 29797 5180 29867 5206
rect 29925 5180 29995 5206
rect 30053 5180 30123 5206
rect 30181 5180 30251 5206
rect 30309 5180 30379 5206
rect 30437 5180 30507 5206
rect 30565 5180 30635 5206
rect 30693 5180 30763 5206
rect 30821 5180 30891 5206
rect 30949 5180 31019 5206
rect 31077 5180 31147 5206
rect 31205 5180 31275 5206
rect 31333 5180 31403 5206
rect 31461 5180 31531 5206
rect 31589 5180 31659 5206
rect 31717 5180 31787 5206
rect 31845 5180 31915 5206
rect 31973 5180 32043 5206
rect 32101 5180 32171 5206
rect 32229 5180 32299 5206
rect 32357 5180 32427 5206
rect 32485 5180 32555 5206
rect 32613 5180 32683 5206
rect 32741 5180 32811 5206
rect 32869 5180 32939 5206
rect 32997 5180 33067 5206
rect 33125 5180 33195 5206
rect 33253 5180 33323 5206
rect 33381 5180 33451 5206
rect 33509 5180 33579 5206
rect 33637 5180 33707 5206
rect 33765 5180 33835 5206
rect 33893 5180 33963 5206
rect 34021 5180 34091 5206
rect 34149 5180 34219 5206
rect 34277 5180 34347 5206
rect 34405 5180 34475 5206
rect 34533 5180 34603 5206
rect 34661 5180 34731 5206
rect 34789 5180 34859 5206
rect 34917 5180 34987 5206
rect 35045 5180 35115 5206
rect 35173 5180 35243 5206
rect 35301 5180 35371 5206
rect 35429 5180 35499 5206
rect 35557 5180 35627 5206
rect 35685 5180 35755 5206
rect 35813 5180 35883 5206
rect 35941 5180 36011 5206
rect 36069 5180 36139 5206
rect 36197 5180 36267 5206
rect 36325 5180 36395 5206
rect 36453 5180 36523 5206
rect 36581 5180 36651 5206
rect 36709 5180 36779 5206
rect 36837 5180 36907 5206
rect 36965 5180 37035 5206
rect 37093 5180 37163 5206
rect 37221 5180 37291 5206
rect 37349 5180 37419 5206
rect 37477 5180 37547 5206
<< polycont >>
rect -285 6044 -251 6078
rect 765 6044 799 6078
rect 4123 6123 4157 6157
rect 1985 6033 2019 6067
rect 7700 6120 7734 6154
rect 14715 6048 14749 6082
rect 28743 6068 28777 6102
rect -372 5338 -338 5372
rect 977 5401 1011 5435
rect 2506 5401 2540 5435
rect 4677 5410 4711 5444
rect 7935 5395 7969 5429
rect 15704 5364 15738 5398
<< locali >>
rect -363 6308 28671 6312
rect -363 6270 -319 6308
rect -281 6270 -191 6308
rect -153 6270 481 6308
rect 519 6270 609 6308
rect 647 6270 737 6308
rect 775 6270 1361 6308
rect 1399 6270 1489 6308
rect 1527 6270 1617 6308
rect 1655 6270 1745 6308
rect 1783 6270 1873 6308
rect 1911 6270 2980 6308
rect 3018 6270 3108 6308
rect 3146 6270 3236 6308
rect 3274 6270 3364 6308
rect 3402 6270 3492 6308
rect 3530 6270 3620 6308
rect 3658 6270 3748 6308
rect 3786 6270 3876 6308
rect 3914 6270 4004 6308
rect 4042 6270 5473 6308
rect 5511 6270 5601 6308
rect 5639 6270 5729 6308
rect 5767 6270 5857 6308
rect 5895 6270 5985 6308
rect 6023 6270 6113 6308
rect 6151 6270 6241 6308
rect 6279 6270 6369 6308
rect 6407 6270 6497 6308
rect 6535 6270 6625 6308
rect 6663 6270 6753 6308
rect 6791 6270 6881 6308
rect 6919 6270 7009 6308
rect 7047 6270 7137 6308
rect 7175 6270 7265 6308
rect 7303 6270 7393 6308
rect 7431 6270 7521 6308
rect 7559 6270 10560 6308
rect 10598 6270 10688 6308
rect 10726 6270 10816 6308
rect 10854 6270 10944 6308
rect 10982 6270 11072 6308
rect 11110 6270 11200 6308
rect 11238 6270 11328 6308
rect 11366 6270 11456 6308
rect 11494 6270 11584 6308
rect 11622 6270 11712 6308
rect 11750 6270 11840 6308
rect 11878 6270 11968 6308
rect 12006 6270 12096 6308
rect 12134 6270 12224 6308
rect 12262 6270 12352 6308
rect 12390 6270 12480 6308
rect 12518 6270 12608 6308
rect 12646 6270 12736 6308
rect 12774 6270 12864 6308
rect 12902 6270 12992 6308
rect 13030 6270 13120 6308
rect 13158 6270 13248 6308
rect 13286 6270 13376 6308
rect 13414 6270 13504 6308
rect 13542 6270 13632 6308
rect 13670 6270 13760 6308
rect 13798 6270 13888 6308
rect 13926 6270 14016 6308
rect 14054 6270 14144 6308
rect 14182 6270 14272 6308
rect 14310 6270 14400 6308
rect 14438 6270 14528 6308
rect 14566 6270 14656 6308
rect 14694 6270 20397 6308
rect 20435 6270 20525 6308
rect 20563 6270 20653 6308
rect 20691 6270 20781 6308
rect 20819 6270 20909 6308
rect 20947 6270 21037 6308
rect 21075 6270 21165 6308
rect 21203 6270 21293 6308
rect 21331 6270 21421 6308
rect 21459 6270 21549 6308
rect 21587 6270 21677 6308
rect 21715 6270 21805 6308
rect 21843 6270 21933 6308
rect 21971 6270 22061 6308
rect 22099 6270 22189 6308
rect 22227 6270 22317 6308
rect 22355 6270 22445 6308
rect 22483 6270 22573 6308
rect 22611 6270 22701 6308
rect 22739 6270 22829 6308
rect 22867 6270 22957 6308
rect 22995 6270 23085 6308
rect 23123 6270 23213 6308
rect 23251 6270 23341 6308
rect 23379 6270 23469 6308
rect 23507 6270 23597 6308
rect 23635 6270 23725 6308
rect 23763 6270 23853 6308
rect 23891 6270 23981 6308
rect 24019 6270 24109 6308
rect 24147 6270 24237 6308
rect 24275 6270 24365 6308
rect 24403 6270 24493 6308
rect 24531 6270 24621 6308
rect 24659 6270 24749 6308
rect 24787 6270 24877 6308
rect 24915 6270 25005 6308
rect 25043 6270 25133 6308
rect 25171 6270 25261 6308
rect 25299 6270 25389 6308
rect 25427 6270 25517 6308
rect 25555 6270 25645 6308
rect 25683 6270 25773 6308
rect 25811 6270 25901 6308
rect 25939 6270 26029 6308
rect 26067 6270 26157 6308
rect 26195 6270 26285 6308
rect 26323 6270 26413 6308
rect 26451 6270 26541 6308
rect 26579 6270 26669 6308
rect 26707 6270 26797 6308
rect 26835 6270 26925 6308
rect 26963 6270 27053 6308
rect 27091 6270 27181 6308
rect 27219 6270 27309 6308
rect 27347 6270 27437 6308
rect 27475 6270 27565 6308
rect 27603 6270 27693 6308
rect 27731 6270 27821 6308
rect 27859 6270 27949 6308
rect 27987 6270 28077 6308
rect 28115 6270 28205 6308
rect 28243 6270 28333 6308
rect 28371 6270 28461 6308
rect 28499 6270 28589 6308
rect 28627 6270 28671 6308
rect -363 6266 28671 6270
rect -317 6200 -283 6216
rect -317 6124 -283 6140
rect -189 6200 -155 6216
rect -189 6124 -155 6140
rect 483 6200 517 6216
rect 483 6124 517 6140
rect 611 6200 645 6216
rect 611 6124 645 6140
rect 739 6200 773 6216
rect 739 6124 773 6140
rect 1363 6200 1397 6216
rect 1363 6124 1397 6140
rect 1491 6200 1525 6216
rect 1491 6124 1525 6140
rect 1619 6200 1653 6216
rect 1619 6124 1653 6140
rect 1747 6200 1781 6216
rect 1747 6124 1781 6140
rect 1875 6200 1909 6216
rect 1875 6124 1909 6140
rect 2982 6200 3016 6216
rect 2982 6124 3016 6140
rect 3110 6200 3144 6216
rect 3110 6124 3144 6140
rect 3238 6200 3272 6216
rect 3238 6124 3272 6140
rect 3366 6200 3400 6216
rect 3366 6124 3400 6140
rect 3494 6200 3528 6216
rect 3494 6124 3528 6140
rect 3622 6200 3656 6216
rect 3622 6124 3656 6140
rect 3750 6200 3784 6216
rect 3750 6124 3784 6140
rect 3878 6200 3912 6216
rect 3878 6124 3912 6140
rect 4006 6200 4040 6216
rect 5475 6200 5509 6216
rect 4006 6124 4040 6140
rect 4107 6118 4118 6161
rect 4163 6118 4173 6161
rect 5475 6124 5509 6140
rect 5603 6200 5637 6216
rect 5603 6124 5637 6140
rect 5731 6200 5765 6216
rect 5731 6124 5765 6140
rect 5859 6200 5893 6216
rect 5859 6124 5893 6140
rect 5987 6200 6021 6216
rect 5987 6124 6021 6140
rect 6115 6200 6149 6216
rect 6115 6124 6149 6140
rect 6243 6200 6277 6216
rect 6243 6124 6277 6140
rect 6371 6200 6405 6216
rect 6371 6124 6405 6140
rect 6499 6200 6533 6216
rect 6499 6124 6533 6140
rect 6627 6200 6661 6216
rect 6627 6124 6661 6140
rect 6755 6200 6789 6216
rect 6755 6124 6789 6140
rect 6883 6200 6917 6216
rect 6883 6124 6917 6140
rect 7011 6200 7045 6216
rect 7011 6124 7045 6140
rect 7139 6200 7173 6216
rect 7139 6124 7173 6140
rect 7267 6200 7301 6216
rect 7267 6124 7301 6140
rect 7395 6200 7429 6216
rect 7395 6124 7429 6140
rect 7523 6200 7557 6216
rect 10562 6200 10596 6216
rect 7523 6124 7557 6140
rect 7684 6115 7695 6158
rect 7740 6115 7750 6158
rect 10562 6124 10596 6140
rect 10690 6200 10724 6216
rect 10690 6124 10724 6140
rect 10818 6200 10852 6216
rect 10818 6124 10852 6140
rect 10946 6200 10980 6216
rect 10946 6124 10980 6140
rect 11074 6200 11108 6216
rect 11074 6124 11108 6140
rect 11202 6200 11236 6216
rect 11202 6124 11236 6140
rect 11330 6200 11364 6216
rect 11330 6124 11364 6140
rect 11458 6200 11492 6216
rect 11458 6124 11492 6140
rect 11586 6200 11620 6216
rect 11586 6124 11620 6140
rect 11714 6200 11748 6216
rect 11714 6124 11748 6140
rect 11842 6200 11876 6216
rect 11842 6124 11876 6140
rect 11970 6200 12004 6216
rect 11970 6124 12004 6140
rect 12098 6200 12132 6216
rect 12098 6124 12132 6140
rect 12226 6200 12260 6216
rect 12226 6124 12260 6140
rect 12354 6200 12388 6216
rect 12354 6124 12388 6140
rect 12482 6200 12516 6216
rect 12482 6124 12516 6140
rect 12610 6200 12644 6216
rect 12610 6124 12644 6140
rect 12738 6200 12772 6216
rect 12738 6124 12772 6140
rect 12866 6200 12900 6216
rect 12866 6124 12900 6140
rect 12994 6200 13028 6216
rect 12994 6124 13028 6140
rect 13122 6200 13156 6216
rect 13122 6124 13156 6140
rect 13250 6200 13284 6216
rect 13250 6124 13284 6140
rect 13378 6200 13412 6216
rect 13378 6124 13412 6140
rect 13506 6200 13540 6216
rect 13506 6124 13540 6140
rect 13634 6200 13668 6216
rect 13634 6124 13668 6140
rect 13762 6200 13796 6216
rect 13762 6124 13796 6140
rect 13890 6200 13924 6216
rect 13890 6124 13924 6140
rect 14018 6200 14052 6216
rect 14018 6124 14052 6140
rect 14146 6200 14180 6216
rect 14146 6124 14180 6140
rect 14274 6200 14308 6216
rect 14274 6124 14308 6140
rect 14402 6200 14436 6216
rect 14402 6124 14436 6140
rect 14530 6200 14564 6216
rect 14530 6124 14564 6140
rect 14658 6200 14692 6216
rect 14658 6124 14692 6140
rect 20399 6200 20433 6216
rect 20399 6124 20433 6140
rect 20527 6200 20561 6216
rect 20527 6124 20561 6140
rect 20655 6200 20689 6216
rect 20655 6124 20689 6140
rect 20783 6200 20817 6216
rect 20783 6124 20817 6140
rect 20911 6200 20945 6216
rect 20911 6124 20945 6140
rect 21039 6200 21073 6216
rect 21039 6124 21073 6140
rect 21167 6200 21201 6216
rect 21167 6124 21201 6140
rect 21295 6200 21329 6216
rect 21295 6124 21329 6140
rect 21423 6200 21457 6216
rect 21423 6124 21457 6140
rect 21551 6200 21585 6216
rect 21551 6124 21585 6140
rect 21679 6200 21713 6216
rect 21679 6124 21713 6140
rect 21807 6200 21841 6216
rect 21807 6124 21841 6140
rect 21935 6200 21969 6216
rect 21935 6124 21969 6140
rect 22063 6200 22097 6216
rect 22063 6124 22097 6140
rect 22191 6200 22225 6216
rect 22191 6124 22225 6140
rect 22319 6200 22353 6216
rect 22319 6124 22353 6140
rect 22447 6200 22481 6216
rect 22447 6124 22481 6140
rect 22575 6200 22609 6216
rect 22575 6124 22609 6140
rect 22703 6200 22737 6216
rect 22703 6124 22737 6140
rect 22831 6200 22865 6216
rect 22831 6124 22865 6140
rect 22959 6200 22993 6216
rect 22959 6124 22993 6140
rect 23087 6200 23121 6216
rect 23087 6124 23121 6140
rect 23215 6200 23249 6216
rect 23215 6124 23249 6140
rect 23343 6200 23377 6216
rect 23343 6124 23377 6140
rect 23471 6200 23505 6216
rect 23471 6124 23505 6140
rect 23599 6200 23633 6216
rect 23599 6124 23633 6140
rect 23727 6200 23761 6216
rect 23727 6124 23761 6140
rect 23855 6200 23889 6216
rect 23855 6124 23889 6140
rect 23983 6200 24017 6216
rect 23983 6124 24017 6140
rect 24111 6200 24145 6216
rect 24111 6124 24145 6140
rect 24239 6200 24273 6216
rect 24239 6124 24273 6140
rect 24367 6200 24401 6216
rect 24367 6124 24401 6140
rect 24495 6200 24529 6216
rect 24495 6124 24529 6140
rect 24623 6200 24657 6216
rect 24623 6124 24657 6140
rect 24751 6200 24785 6216
rect 24751 6124 24785 6140
rect 24879 6200 24913 6216
rect 24879 6124 24913 6140
rect 25007 6200 25041 6216
rect 25007 6124 25041 6140
rect 25135 6200 25169 6216
rect 25135 6124 25169 6140
rect 25263 6200 25297 6216
rect 25263 6124 25297 6140
rect 25391 6200 25425 6216
rect 25391 6124 25425 6140
rect 25519 6200 25553 6216
rect 25519 6124 25553 6140
rect 25647 6200 25681 6216
rect 25647 6124 25681 6140
rect 25775 6200 25809 6216
rect 25775 6124 25809 6140
rect 25903 6200 25937 6216
rect 25903 6124 25937 6140
rect 26031 6200 26065 6216
rect 26031 6124 26065 6140
rect 26159 6200 26193 6216
rect 26159 6124 26193 6140
rect 26287 6200 26321 6216
rect 26287 6124 26321 6140
rect 26415 6200 26449 6216
rect 26415 6124 26449 6140
rect 26543 6200 26577 6216
rect 26543 6124 26577 6140
rect 26671 6200 26705 6216
rect 26671 6124 26705 6140
rect 26799 6200 26833 6216
rect 26799 6124 26833 6140
rect 26927 6200 26961 6216
rect 26927 6124 26961 6140
rect 27055 6200 27089 6216
rect 27055 6124 27089 6140
rect 27183 6200 27217 6216
rect 27183 6124 27217 6140
rect 27311 6200 27345 6216
rect 27311 6124 27345 6140
rect 27439 6200 27473 6216
rect 27439 6124 27473 6140
rect 27567 6200 27601 6216
rect 27567 6124 27601 6140
rect 27695 6200 27729 6216
rect 27695 6124 27729 6140
rect 27823 6200 27857 6216
rect 27823 6124 27857 6140
rect 27951 6200 27985 6216
rect 27951 6124 27985 6140
rect 28079 6200 28113 6216
rect 28079 6124 28113 6140
rect 28207 6200 28241 6216
rect 28207 6124 28241 6140
rect 28335 6200 28369 6216
rect 28335 6124 28369 6140
rect 28463 6200 28497 6216
rect 28463 6124 28497 6140
rect 28591 6200 28625 6216
rect 28591 6124 28625 6140
rect -301 6039 -290 6082
rect -245 6039 -235 6082
rect 749 6039 760 6082
rect 805 6039 815 6082
rect 1969 6028 1980 6071
rect 2025 6028 2035 6071
rect 14699 6043 14710 6086
rect 14755 6043 14765 6086
rect 28727 6064 28737 6107
rect 28782 6064 28793 6107
rect -317 5984 -283 6000
rect -317 5824 -283 5840
rect -189 5984 -155 6000
rect -189 5824 -155 5840
rect 483 5984 517 6000
rect 483 5824 517 5840
rect 611 5984 645 6000
rect 611 5824 645 5840
rect 739 5984 773 6000
rect 739 5824 773 5840
rect 1363 5984 1397 6000
rect 1363 5824 1397 5840
rect 1491 5984 1525 6000
rect 1491 5824 1525 5840
rect 1619 5984 1653 6000
rect 1619 5824 1653 5840
rect 1747 5984 1781 6000
rect 1747 5824 1781 5840
rect 1875 5984 1909 6000
rect 1875 5824 1909 5840
rect 2982 5984 3016 6000
rect 2982 5824 3016 5840
rect 3110 5984 3144 6000
rect 3110 5824 3144 5840
rect 3238 5984 3272 6000
rect 3238 5824 3272 5840
rect 3366 5984 3400 6000
rect 3366 5824 3400 5840
rect 3494 5984 3528 6000
rect 3494 5824 3528 5840
rect 3622 5984 3656 6000
rect 3622 5824 3656 5840
rect 3750 5984 3784 6000
rect 3750 5824 3784 5840
rect 3878 5984 3912 6000
rect 3878 5824 3912 5840
rect 4006 5984 4040 6000
rect 4006 5824 4040 5840
rect 5475 5984 5509 6000
rect 5475 5824 5509 5840
rect 5603 5984 5637 6000
rect 5603 5824 5637 5840
rect 5731 5984 5765 6000
rect 5731 5824 5765 5840
rect 5859 5984 5893 6000
rect 5859 5824 5893 5840
rect 5987 5984 6021 6000
rect 5987 5824 6021 5840
rect 6115 5984 6149 6000
rect 6115 5824 6149 5840
rect 6243 5984 6277 6000
rect 6243 5824 6277 5840
rect 6371 5984 6405 6000
rect 6371 5824 6405 5840
rect 6499 5984 6533 6000
rect 6499 5824 6533 5840
rect 6627 5984 6661 6000
rect 6627 5824 6661 5840
rect 6755 5984 6789 6000
rect 6755 5824 6789 5840
rect 6883 5984 6917 6000
rect 6883 5824 6917 5840
rect 7011 5984 7045 6000
rect 7011 5824 7045 5840
rect 7139 5984 7173 6000
rect 7139 5824 7173 5840
rect 7267 5984 7301 6000
rect 7267 5824 7301 5840
rect 7395 5984 7429 6000
rect 7395 5824 7429 5840
rect 7523 5984 7557 6000
rect 7523 5824 7557 5840
rect 10562 5984 10596 6000
rect 10562 5824 10596 5840
rect 10690 5984 10724 6000
rect 10690 5824 10724 5840
rect 10818 5984 10852 6000
rect 10818 5824 10852 5840
rect 10946 5984 10980 6000
rect 10946 5824 10980 5840
rect 11074 5984 11108 6000
rect 11074 5824 11108 5840
rect 11202 5984 11236 6000
rect 11202 5824 11236 5840
rect 11330 5984 11364 6000
rect 11330 5824 11364 5840
rect 11458 5984 11492 6000
rect 11458 5824 11492 5840
rect 11586 5984 11620 6000
rect 11586 5824 11620 5840
rect 11714 5984 11748 6000
rect 11714 5824 11748 5840
rect 11842 5984 11876 6000
rect 11842 5824 11876 5840
rect 11970 5984 12004 6000
rect 11970 5824 12004 5840
rect 12098 5984 12132 6000
rect 12098 5824 12132 5840
rect 12226 5984 12260 6000
rect 12226 5824 12260 5840
rect 12354 5984 12388 6000
rect 12354 5824 12388 5840
rect 12482 5984 12516 6000
rect 12482 5824 12516 5840
rect 12610 5984 12644 6000
rect 12610 5824 12644 5840
rect 12738 5984 12772 6000
rect 12738 5824 12772 5840
rect 12866 5984 12900 6000
rect 12866 5824 12900 5840
rect 12994 5984 13028 6000
rect 12994 5824 13028 5840
rect 13122 5984 13156 6000
rect 13122 5824 13156 5840
rect 13250 5984 13284 6000
rect 13250 5824 13284 5840
rect 13378 5984 13412 6000
rect 13378 5824 13412 5840
rect 13506 5984 13540 6000
rect 13506 5824 13540 5840
rect 13634 5984 13668 6000
rect 13634 5824 13668 5840
rect 13762 5984 13796 6000
rect 13762 5824 13796 5840
rect 13890 5984 13924 6000
rect 13890 5824 13924 5840
rect 14018 5984 14052 6000
rect 14018 5824 14052 5840
rect 14146 5984 14180 6000
rect 14146 5824 14180 5840
rect 14274 5984 14308 6000
rect 14274 5824 14308 5840
rect 14402 5984 14436 6000
rect 14402 5824 14436 5840
rect 14530 5984 14564 6000
rect 14530 5824 14564 5840
rect 14658 5984 14692 6000
rect 14658 5824 14692 5840
rect 20399 5984 20433 6000
rect 20399 5824 20433 5840
rect 20527 5984 20561 6000
rect 20527 5824 20561 5840
rect 20655 5984 20689 6000
rect 20655 5824 20689 5840
rect 20783 5984 20817 6000
rect 20783 5824 20817 5840
rect 20911 5984 20945 6000
rect 20911 5824 20945 5840
rect 21039 5984 21073 6000
rect 21039 5824 21073 5840
rect 21167 5984 21201 6000
rect 21167 5824 21201 5840
rect 21295 5984 21329 6000
rect 21295 5824 21329 5840
rect 21423 5984 21457 6000
rect 21423 5824 21457 5840
rect 21551 5984 21585 6000
rect 21551 5824 21585 5840
rect 21679 5984 21713 6000
rect 21679 5824 21713 5840
rect 21807 5984 21841 6000
rect 21807 5824 21841 5840
rect 21935 5984 21969 6000
rect 21935 5824 21969 5840
rect 22063 5984 22097 6000
rect 22063 5824 22097 5840
rect 22191 5984 22225 6000
rect 22191 5824 22225 5840
rect 22319 5984 22353 6000
rect 22319 5824 22353 5840
rect 22447 5984 22481 6000
rect 22447 5824 22481 5840
rect 22575 5984 22609 6000
rect 22575 5824 22609 5840
rect 22703 5984 22737 6000
rect 22703 5824 22737 5840
rect 22831 5984 22865 6000
rect 22831 5824 22865 5840
rect 22959 5984 22993 6000
rect 22959 5824 22993 5840
rect 23087 5984 23121 6000
rect 23087 5824 23121 5840
rect 23215 5984 23249 6000
rect 23215 5824 23249 5840
rect 23343 5984 23377 6000
rect 23343 5824 23377 5840
rect 23471 5984 23505 6000
rect 23471 5824 23505 5840
rect 23599 5984 23633 6000
rect 23599 5824 23633 5840
rect 23727 5984 23761 6000
rect 23727 5824 23761 5840
rect 23855 5984 23889 6000
rect 23855 5824 23889 5840
rect 23983 5984 24017 6000
rect 23983 5824 24017 5840
rect 24111 5984 24145 6000
rect 24111 5824 24145 5840
rect 24239 5984 24273 6000
rect 24239 5824 24273 5840
rect 24367 5984 24401 6000
rect 24367 5824 24401 5840
rect 24495 5984 24529 6000
rect 24495 5824 24529 5840
rect 24623 5984 24657 6000
rect 24623 5824 24657 5840
rect 24751 5984 24785 6000
rect 24751 5824 24785 5840
rect 24879 5984 24913 6000
rect 24879 5824 24913 5840
rect 25007 5984 25041 6000
rect 25007 5824 25041 5840
rect 25135 5984 25169 6000
rect 25135 5824 25169 5840
rect 25263 5984 25297 6000
rect 25263 5824 25297 5840
rect 25391 5984 25425 6000
rect 25391 5824 25425 5840
rect 25519 5984 25553 6000
rect 25519 5824 25553 5840
rect 25647 5984 25681 6000
rect 25647 5824 25681 5840
rect 25775 5984 25809 6000
rect 25775 5824 25809 5840
rect 25903 5984 25937 6000
rect 25903 5824 25937 5840
rect 26031 5984 26065 6000
rect 26031 5824 26065 5840
rect 26159 5984 26193 6000
rect 26159 5824 26193 5840
rect 26287 5984 26321 6000
rect 26287 5824 26321 5840
rect 26415 5984 26449 6000
rect 26415 5824 26449 5840
rect 26543 5984 26577 6000
rect 26543 5824 26577 5840
rect 26671 5984 26705 6000
rect 26671 5824 26705 5840
rect 26799 5984 26833 6000
rect 26799 5824 26833 5840
rect 26927 5984 26961 6000
rect 26927 5824 26961 5840
rect 27055 5984 27089 6000
rect 27055 5824 27089 5840
rect 27183 5984 27217 6000
rect 27183 5824 27217 5840
rect 27311 5984 27345 6000
rect 27311 5824 27345 5840
rect 27439 5984 27473 6000
rect 27439 5824 27473 5840
rect 27567 5984 27601 6000
rect 27567 5824 27601 5840
rect 27695 5984 27729 6000
rect 27695 5824 27729 5840
rect 27823 5984 27857 6000
rect 27823 5824 27857 5840
rect 27951 5984 27985 6000
rect 27951 5824 27985 5840
rect 28079 5984 28113 6000
rect 28079 5824 28113 5840
rect 28207 5984 28241 6000
rect 28207 5824 28241 5840
rect 28335 5984 28369 6000
rect 28335 5824 28369 5840
rect 28463 5984 28497 6000
rect 28463 5824 28497 5840
rect 28591 5984 28625 6000
rect 28591 5824 28625 5840
rect -363 5728 37639 5732
rect -363 5690 -319 5728
rect -281 5690 -191 5728
rect -153 5690 481 5728
rect 519 5690 609 5728
rect 647 5690 737 5728
rect 775 5690 865 5728
rect 903 5690 1361 5728
rect 1399 5690 1489 5728
rect 1527 5690 1617 5728
rect 1655 5690 1745 5728
rect 1783 5690 1873 5728
rect 1911 5690 2001 5728
rect 2039 5690 2129 5728
rect 2167 5690 2257 5728
rect 2295 5690 2385 5728
rect 2423 5690 2980 5728
rect 3018 5690 3108 5728
rect 3146 5690 3236 5728
rect 3274 5690 3364 5728
rect 3402 5690 3492 5728
rect 3530 5690 3620 5728
rect 3658 5690 3748 5728
rect 3786 5690 3876 5728
rect 3914 5690 4004 5728
rect 4042 5690 4132 5728
rect 4170 5690 4260 5728
rect 4298 5690 4388 5728
rect 4426 5690 4516 5728
rect 4554 5690 5473 5728
rect 5511 5690 5601 5728
rect 5639 5690 5729 5728
rect 5767 5690 5857 5728
rect 5895 5690 5985 5728
rect 6023 5690 6113 5728
rect 6151 5690 6241 5728
rect 6279 5690 6369 5728
rect 6407 5690 6497 5728
rect 6535 5690 6625 5728
rect 6663 5690 6753 5728
rect 6791 5690 6881 5728
rect 6919 5690 7009 5728
rect 7047 5690 7137 5728
rect 7175 5690 7265 5728
rect 7303 5690 7393 5728
rect 7431 5690 7521 5728
rect 7559 5690 8057 5728
rect 8095 5690 8185 5728
rect 8223 5690 8313 5728
rect 8351 5690 8441 5728
rect 8479 5690 8569 5728
rect 8607 5690 8697 5728
rect 8735 5690 8825 5728
rect 8863 5690 8953 5728
rect 8991 5690 9081 5728
rect 9119 5690 9209 5728
rect 9247 5690 9337 5728
rect 9375 5690 9465 5728
rect 9503 5690 9593 5728
rect 9631 5690 9721 5728
rect 9759 5690 9849 5728
rect 9887 5690 9977 5728
rect 10015 5690 10105 5728
rect 10143 5690 10560 5728
rect 10598 5690 10688 5728
rect 10726 5690 10816 5728
rect 10854 5690 10944 5728
rect 10982 5690 11072 5728
rect 11110 5690 11200 5728
rect 11238 5690 11328 5728
rect 11366 5690 11456 5728
rect 11494 5690 11584 5728
rect 11622 5690 11712 5728
rect 11750 5690 11840 5728
rect 11878 5690 11968 5728
rect 12006 5690 12096 5728
rect 12134 5690 12224 5728
rect 12262 5690 12352 5728
rect 12390 5690 12480 5728
rect 12518 5690 12608 5728
rect 12646 5690 12736 5728
rect 12774 5690 12864 5728
rect 12902 5690 12992 5728
rect 13030 5690 13120 5728
rect 13158 5690 13248 5728
rect 13286 5690 13376 5728
rect 13414 5690 13504 5728
rect 13542 5690 13632 5728
rect 13670 5690 13760 5728
rect 13798 5690 13888 5728
rect 13926 5690 14016 5728
rect 14054 5690 14144 5728
rect 14182 5690 14272 5728
rect 14310 5690 14400 5728
rect 14438 5690 14528 5728
rect 14566 5690 14656 5728
rect 14694 5690 15821 5728
rect 15859 5690 15949 5728
rect 15987 5690 16077 5728
rect 16115 5690 16205 5728
rect 16243 5690 16333 5728
rect 16371 5690 16461 5728
rect 16499 5690 16589 5728
rect 16627 5690 16717 5728
rect 16755 5690 16845 5728
rect 16883 5690 16973 5728
rect 17011 5690 17101 5728
rect 17139 5690 17229 5728
rect 17267 5690 17357 5728
rect 17395 5690 17485 5728
rect 17523 5690 17613 5728
rect 17651 5690 17741 5728
rect 17779 5690 17869 5728
rect 17907 5690 17997 5728
rect 18035 5690 18125 5728
rect 18163 5690 18253 5728
rect 18291 5690 18381 5728
rect 18419 5690 18509 5728
rect 18547 5690 18637 5728
rect 18675 5690 18765 5728
rect 18803 5690 18893 5728
rect 18931 5690 19021 5728
rect 19059 5690 19149 5728
rect 19187 5690 19277 5728
rect 19315 5690 19405 5728
rect 19443 5690 19533 5728
rect 19571 5690 19661 5728
rect 19699 5690 19789 5728
rect 19827 5690 19917 5728
rect 19955 5690 20397 5728
rect 20435 5690 20525 5728
rect 20563 5690 20653 5728
rect 20691 5690 20781 5728
rect 20819 5690 20909 5728
rect 20947 5690 21037 5728
rect 21075 5690 21165 5728
rect 21203 5690 21293 5728
rect 21331 5690 21421 5728
rect 21459 5690 21549 5728
rect 21587 5690 21677 5728
rect 21715 5690 21805 5728
rect 21843 5690 21933 5728
rect 21971 5690 22061 5728
rect 22099 5690 22189 5728
rect 22227 5690 22317 5728
rect 22355 5690 22445 5728
rect 22483 5690 22573 5728
rect 22611 5690 22701 5728
rect 22739 5690 22829 5728
rect 22867 5690 22957 5728
rect 22995 5690 23085 5728
rect 23123 5690 23213 5728
rect 23251 5690 23341 5728
rect 23379 5690 23469 5728
rect 23507 5690 23597 5728
rect 23635 5690 23725 5728
rect 23763 5690 23853 5728
rect 23891 5690 23981 5728
rect 24019 5690 24109 5728
rect 24147 5690 24237 5728
rect 24275 5690 24365 5728
rect 24403 5690 24493 5728
rect 24531 5690 24621 5728
rect 24659 5690 24749 5728
rect 24787 5690 24877 5728
rect 24915 5690 25005 5728
rect 25043 5690 25133 5728
rect 25171 5690 25261 5728
rect 25299 5690 25389 5728
rect 25427 5690 25517 5728
rect 25555 5690 25645 5728
rect 25683 5690 25773 5728
rect 25811 5690 25901 5728
rect 25939 5690 26029 5728
rect 26067 5690 26157 5728
rect 26195 5690 26285 5728
rect 26323 5690 26413 5728
rect 26451 5690 26541 5728
rect 26579 5690 26669 5728
rect 26707 5690 26797 5728
rect 26835 5690 26925 5728
rect 26963 5690 27053 5728
rect 27091 5690 27181 5728
rect 27219 5690 27309 5728
rect 27347 5690 27437 5728
rect 27475 5690 27565 5728
rect 27603 5690 27693 5728
rect 27731 5690 27821 5728
rect 27859 5690 27949 5728
rect 27987 5690 28077 5728
rect 28115 5690 28205 5728
rect 28243 5690 28333 5728
rect 28371 5690 28461 5728
rect 28499 5690 28589 5728
rect 28627 5690 29365 5728
rect 29403 5690 29493 5728
rect 29531 5690 29621 5728
rect 29659 5690 29749 5728
rect 29787 5690 29877 5728
rect 29915 5690 30005 5728
rect 30043 5690 30133 5728
rect 30171 5690 30261 5728
rect 30299 5690 30389 5728
rect 30427 5690 30517 5728
rect 30555 5690 30645 5728
rect 30683 5690 30773 5728
rect 30811 5690 30901 5728
rect 30939 5690 31029 5728
rect 31067 5690 31157 5728
rect 31195 5690 31285 5728
rect 31323 5690 31413 5728
rect 31451 5690 31541 5728
rect 31579 5690 31669 5728
rect 31707 5690 31797 5728
rect 31835 5690 31925 5728
rect 31963 5690 32053 5728
rect 32091 5690 32181 5728
rect 32219 5690 32309 5728
rect 32347 5690 32437 5728
rect 32475 5690 32565 5728
rect 32603 5690 32693 5728
rect 32731 5690 32821 5728
rect 32859 5690 32949 5728
rect 32987 5690 33077 5728
rect 33115 5690 33205 5728
rect 33243 5690 33333 5728
rect 33371 5690 33461 5728
rect 33499 5690 33589 5728
rect 33627 5690 33717 5728
rect 33755 5690 33845 5728
rect 33883 5690 33973 5728
rect 34011 5690 34101 5728
rect 34139 5690 34229 5728
rect 34267 5690 34357 5728
rect 34395 5690 34485 5728
rect 34523 5690 34613 5728
rect 34651 5690 34741 5728
rect 34779 5690 34869 5728
rect 34907 5690 34997 5728
rect 35035 5690 35125 5728
rect 35163 5690 35253 5728
rect 35291 5690 35381 5728
rect 35419 5690 35509 5728
rect 35547 5690 35637 5728
rect 35675 5690 35765 5728
rect 35803 5690 35893 5728
rect 35931 5690 36021 5728
rect 36059 5690 36149 5728
rect 36187 5690 36277 5728
rect 36315 5690 36405 5728
rect 36443 5690 36533 5728
rect 36571 5690 36661 5728
rect 36699 5690 36789 5728
rect 36827 5690 36917 5728
rect 36955 5690 37045 5728
rect 37083 5690 37173 5728
rect 37211 5690 37301 5728
rect 37339 5690 37429 5728
rect 37467 5690 37557 5728
rect 37595 5690 37639 5728
rect -363 5686 37639 5690
rect -317 5578 -283 5594
rect -317 5418 -283 5434
rect -189 5578 -155 5594
rect -189 5418 -155 5434
rect 611 5578 645 5594
rect 611 5418 645 5434
rect 739 5578 773 5594
rect 739 5418 773 5434
rect 867 5578 901 5594
rect 1875 5578 1909 5594
rect 867 5418 901 5434
rect 961 5396 972 5439
rect 1017 5396 1027 5439
rect 1875 5418 1909 5434
rect 2003 5578 2037 5594
rect 2003 5418 2037 5434
rect 2131 5578 2165 5594
rect 2131 5418 2165 5434
rect 2259 5578 2293 5594
rect 2259 5418 2293 5434
rect 2387 5578 2421 5594
rect 3494 5578 3528 5594
rect 2387 5418 2421 5434
rect 2490 5396 2501 5439
rect 2546 5396 2556 5439
rect 3494 5418 3528 5434
rect 3622 5578 3656 5594
rect 3622 5418 3656 5434
rect 3750 5578 3784 5594
rect 3750 5418 3784 5434
rect 3878 5578 3912 5594
rect 3878 5418 3912 5434
rect 4006 5578 4040 5594
rect 4006 5418 4040 5434
rect 4134 5578 4168 5594
rect 4134 5418 4168 5434
rect 4262 5578 4296 5594
rect 4262 5418 4296 5434
rect 4390 5578 4424 5594
rect 4390 5418 4424 5434
rect 4518 5578 4552 5594
rect 8059 5578 8093 5594
rect 4518 5418 4552 5434
rect 4661 5405 4672 5448
rect 4717 5405 4727 5448
rect 7919 5390 7930 5433
rect 7975 5390 7985 5433
rect 8059 5418 8093 5434
rect 8187 5578 8221 5594
rect 8187 5418 8221 5434
rect 8315 5578 8349 5594
rect 8315 5418 8349 5434
rect 8443 5578 8477 5594
rect 8443 5418 8477 5434
rect 8571 5578 8605 5594
rect 8571 5418 8605 5434
rect 8699 5578 8733 5594
rect 8699 5418 8733 5434
rect 8827 5578 8861 5594
rect 8827 5418 8861 5434
rect 8955 5578 8989 5594
rect 8955 5418 8989 5434
rect 9083 5578 9117 5594
rect 9083 5418 9117 5434
rect 9211 5578 9245 5594
rect 9211 5418 9245 5434
rect 9339 5578 9373 5594
rect 9339 5418 9373 5434
rect 9467 5578 9501 5594
rect 9467 5418 9501 5434
rect 9595 5578 9629 5594
rect 9595 5418 9629 5434
rect 9723 5578 9757 5594
rect 9723 5418 9757 5434
rect 9851 5578 9885 5594
rect 9851 5418 9885 5434
rect 9979 5578 10013 5594
rect 9979 5418 10013 5434
rect 10107 5578 10141 5594
rect 10107 5418 10141 5434
rect 15823 5578 15857 5594
rect 15823 5418 15857 5434
rect 15951 5578 15985 5594
rect 15951 5418 15985 5434
rect 16079 5578 16113 5594
rect 16079 5418 16113 5434
rect 16207 5578 16241 5594
rect 16207 5418 16241 5434
rect 16335 5578 16369 5594
rect 16335 5418 16369 5434
rect 16463 5578 16497 5594
rect 16463 5418 16497 5434
rect 16591 5578 16625 5594
rect 16591 5418 16625 5434
rect 16719 5578 16753 5594
rect 16719 5418 16753 5434
rect 16847 5578 16881 5594
rect 16847 5418 16881 5434
rect 16975 5578 17009 5594
rect 16975 5418 17009 5434
rect 17103 5578 17137 5594
rect 17103 5418 17137 5434
rect 17231 5578 17265 5594
rect 17231 5418 17265 5434
rect 17359 5578 17393 5594
rect 17359 5418 17393 5434
rect 17487 5578 17521 5594
rect 17487 5418 17521 5434
rect 17615 5578 17649 5594
rect 17615 5418 17649 5434
rect 17743 5578 17777 5594
rect 17743 5418 17777 5434
rect 17871 5578 17905 5594
rect 17871 5418 17905 5434
rect 17999 5578 18033 5594
rect 17999 5418 18033 5434
rect 18127 5578 18161 5594
rect 18127 5418 18161 5434
rect 18255 5578 18289 5594
rect 18255 5418 18289 5434
rect 18383 5578 18417 5594
rect 18383 5418 18417 5434
rect 18511 5578 18545 5594
rect 18511 5418 18545 5434
rect 18639 5578 18673 5594
rect 18639 5418 18673 5434
rect 18767 5578 18801 5594
rect 18767 5418 18801 5434
rect 18895 5578 18929 5594
rect 18895 5418 18929 5434
rect 19023 5578 19057 5594
rect 19023 5418 19057 5434
rect 19151 5578 19185 5594
rect 19151 5418 19185 5434
rect 19279 5578 19313 5594
rect 19279 5418 19313 5434
rect 19407 5578 19441 5594
rect 19407 5418 19441 5434
rect 19535 5578 19569 5594
rect 19535 5418 19569 5434
rect 19663 5578 19697 5594
rect 19663 5418 19697 5434
rect 19791 5578 19825 5594
rect 19791 5418 19825 5434
rect 19919 5578 19953 5594
rect 19919 5418 19953 5434
rect 29367 5578 29401 5594
rect 29367 5418 29401 5434
rect 29495 5578 29529 5594
rect 29495 5418 29529 5434
rect 29623 5578 29657 5594
rect 29623 5418 29657 5434
rect 29751 5578 29785 5594
rect 29751 5418 29785 5434
rect 29879 5578 29913 5594
rect 29879 5418 29913 5434
rect 30007 5578 30041 5594
rect 30007 5418 30041 5434
rect 30135 5578 30169 5594
rect 30135 5418 30169 5434
rect 30263 5578 30297 5594
rect 30263 5418 30297 5434
rect 30391 5578 30425 5594
rect 30391 5418 30425 5434
rect 30519 5578 30553 5594
rect 30519 5418 30553 5434
rect 30647 5578 30681 5594
rect 30647 5418 30681 5434
rect 30775 5578 30809 5594
rect 30775 5418 30809 5434
rect 30903 5578 30937 5594
rect 30903 5418 30937 5434
rect 31031 5578 31065 5594
rect 31031 5418 31065 5434
rect 31159 5578 31193 5594
rect 31159 5418 31193 5434
rect 31287 5578 31321 5594
rect 31287 5418 31321 5434
rect 31415 5578 31449 5594
rect 31415 5418 31449 5434
rect 31543 5578 31577 5594
rect 31543 5418 31577 5434
rect 31671 5578 31705 5594
rect 31671 5418 31705 5434
rect 31799 5578 31833 5594
rect 31799 5418 31833 5434
rect 31927 5578 31961 5594
rect 31927 5418 31961 5434
rect 32055 5578 32089 5594
rect 32055 5418 32089 5434
rect 32183 5578 32217 5594
rect 32183 5418 32217 5434
rect 32311 5578 32345 5594
rect 32311 5418 32345 5434
rect 32439 5578 32473 5594
rect 32439 5418 32473 5434
rect 32567 5578 32601 5594
rect 32567 5418 32601 5434
rect 32695 5578 32729 5594
rect 32695 5418 32729 5434
rect 32823 5578 32857 5594
rect 32823 5418 32857 5434
rect 32951 5578 32985 5594
rect 32951 5418 32985 5434
rect 33079 5578 33113 5594
rect 33079 5418 33113 5434
rect 33207 5578 33241 5594
rect 33207 5418 33241 5434
rect 33335 5578 33369 5594
rect 33335 5418 33369 5434
rect 33463 5578 33497 5594
rect 33463 5418 33497 5434
rect 33591 5578 33625 5594
rect 33591 5418 33625 5434
rect 33719 5578 33753 5594
rect 33719 5418 33753 5434
rect 33847 5578 33881 5594
rect 33847 5418 33881 5434
rect 33975 5578 34009 5594
rect 33975 5418 34009 5434
rect 34103 5578 34137 5594
rect 34103 5418 34137 5434
rect 34231 5578 34265 5594
rect 34231 5418 34265 5434
rect 34359 5578 34393 5594
rect 34359 5418 34393 5434
rect 34487 5578 34521 5594
rect 34487 5418 34521 5434
rect 34615 5578 34649 5594
rect 34615 5418 34649 5434
rect 34743 5578 34777 5594
rect 34743 5418 34777 5434
rect 34871 5578 34905 5594
rect 34871 5418 34905 5434
rect 34999 5578 35033 5594
rect 34999 5418 35033 5434
rect 35127 5578 35161 5594
rect 35127 5418 35161 5434
rect 35255 5578 35289 5594
rect 35255 5418 35289 5434
rect 35383 5578 35417 5594
rect 35383 5418 35417 5434
rect 35511 5578 35545 5594
rect 35511 5418 35545 5434
rect 35639 5578 35673 5594
rect 35639 5418 35673 5434
rect 35767 5578 35801 5594
rect 35767 5418 35801 5434
rect 35895 5578 35929 5594
rect 35895 5418 35929 5434
rect 36023 5578 36057 5594
rect 36023 5418 36057 5434
rect 36151 5578 36185 5594
rect 36151 5418 36185 5434
rect 36279 5578 36313 5594
rect 36279 5418 36313 5434
rect 36407 5578 36441 5594
rect 36407 5418 36441 5434
rect 36535 5578 36569 5594
rect 36535 5418 36569 5434
rect 36663 5578 36697 5594
rect 36663 5418 36697 5434
rect 36791 5578 36825 5594
rect 36791 5418 36825 5434
rect 36919 5578 36953 5594
rect 36919 5418 36953 5434
rect 37047 5578 37081 5594
rect 37047 5418 37081 5434
rect 37175 5578 37209 5594
rect 37175 5418 37209 5434
rect 37303 5578 37337 5594
rect 37303 5418 37337 5434
rect 37431 5578 37465 5594
rect 37431 5418 37465 5434
rect 37559 5578 37593 5594
rect 37559 5418 37593 5434
rect -388 5333 -377 5376
rect -332 5333 -322 5376
rect 15688 5359 15699 5402
rect 15744 5359 15754 5402
rect -317 5278 -283 5294
rect -317 5202 -283 5218
rect -189 5278 -155 5294
rect -189 5202 -155 5218
rect 611 5278 645 5294
rect 611 5202 645 5218
rect 739 5278 773 5294
rect 739 5202 773 5218
rect 867 5278 901 5294
rect 867 5202 901 5218
rect 1875 5278 1909 5294
rect 1875 5202 1909 5218
rect 2003 5278 2037 5294
rect 2003 5202 2037 5218
rect 2131 5278 2165 5294
rect 2131 5202 2165 5218
rect 2259 5278 2293 5294
rect 2259 5202 2293 5218
rect 2387 5278 2421 5294
rect 2387 5202 2421 5218
rect 3494 5278 3528 5294
rect 3494 5202 3528 5218
rect 3622 5278 3656 5294
rect 3622 5202 3656 5218
rect 3750 5278 3784 5294
rect 3750 5202 3784 5218
rect 3878 5278 3912 5294
rect 3878 5202 3912 5218
rect 4006 5278 4040 5294
rect 4006 5202 4040 5218
rect 4134 5278 4168 5294
rect 4134 5202 4168 5218
rect 4262 5278 4296 5294
rect 4262 5202 4296 5218
rect 4390 5278 4424 5294
rect 4390 5202 4424 5218
rect 4518 5278 4552 5294
rect 4518 5202 4552 5218
rect 8059 5278 8093 5294
rect 8059 5202 8093 5218
rect 8187 5278 8221 5294
rect 8187 5202 8221 5218
rect 8315 5278 8349 5294
rect 8315 5202 8349 5218
rect 8443 5278 8477 5294
rect 8443 5202 8477 5218
rect 8571 5278 8605 5294
rect 8571 5202 8605 5218
rect 8699 5278 8733 5294
rect 8699 5202 8733 5218
rect 8827 5278 8861 5294
rect 8827 5202 8861 5218
rect 8955 5278 8989 5294
rect 8955 5202 8989 5218
rect 9083 5278 9117 5294
rect 9083 5202 9117 5218
rect 9211 5278 9245 5294
rect 9211 5202 9245 5218
rect 9339 5278 9373 5294
rect 9339 5202 9373 5218
rect 9467 5278 9501 5294
rect 9467 5202 9501 5218
rect 9595 5278 9629 5294
rect 9595 5202 9629 5218
rect 9723 5278 9757 5294
rect 9723 5202 9757 5218
rect 9851 5278 9885 5294
rect 9851 5202 9885 5218
rect 9979 5278 10013 5294
rect 9979 5202 10013 5218
rect 10107 5278 10141 5294
rect 10107 5202 10141 5218
rect 15823 5278 15857 5294
rect 15823 5202 15857 5218
rect 15951 5278 15985 5294
rect 15951 5202 15985 5218
rect 16079 5278 16113 5294
rect 16079 5202 16113 5218
rect 16207 5278 16241 5294
rect 16207 5202 16241 5218
rect 16335 5278 16369 5294
rect 16335 5202 16369 5218
rect 16463 5278 16497 5294
rect 16463 5202 16497 5218
rect 16591 5278 16625 5294
rect 16591 5202 16625 5218
rect 16719 5278 16753 5294
rect 16719 5202 16753 5218
rect 16847 5278 16881 5294
rect 16847 5202 16881 5218
rect 16975 5278 17009 5294
rect 16975 5202 17009 5218
rect 17103 5278 17137 5294
rect 17103 5202 17137 5218
rect 17231 5278 17265 5294
rect 17231 5202 17265 5218
rect 17359 5278 17393 5294
rect 17359 5202 17393 5218
rect 17487 5278 17521 5294
rect 17487 5202 17521 5218
rect 17615 5278 17649 5294
rect 17615 5202 17649 5218
rect 17743 5278 17777 5294
rect 17743 5202 17777 5218
rect 17871 5278 17905 5294
rect 17871 5202 17905 5218
rect 17999 5278 18033 5294
rect 17999 5202 18033 5218
rect 18127 5278 18161 5294
rect 18127 5202 18161 5218
rect 18255 5278 18289 5294
rect 18255 5202 18289 5218
rect 18383 5278 18417 5294
rect 18383 5202 18417 5218
rect 18511 5278 18545 5294
rect 18511 5202 18545 5218
rect 18639 5278 18673 5294
rect 18639 5202 18673 5218
rect 18767 5278 18801 5294
rect 18767 5202 18801 5218
rect 18895 5278 18929 5294
rect 18895 5202 18929 5218
rect 19023 5278 19057 5294
rect 19023 5202 19057 5218
rect 19151 5278 19185 5294
rect 19151 5202 19185 5218
rect 19279 5278 19313 5294
rect 19279 5202 19313 5218
rect 19407 5278 19441 5294
rect 19407 5202 19441 5218
rect 19535 5278 19569 5294
rect 19535 5202 19569 5218
rect 19663 5278 19697 5294
rect 19663 5202 19697 5218
rect 19791 5278 19825 5294
rect 19791 5202 19825 5218
rect 19919 5278 19953 5294
rect 19919 5202 19953 5218
rect 29367 5278 29401 5294
rect 29367 5202 29401 5218
rect 29495 5278 29529 5294
rect 29495 5202 29529 5218
rect 29623 5278 29657 5294
rect 29623 5202 29657 5218
rect 29751 5278 29785 5294
rect 29751 5202 29785 5218
rect 29879 5278 29913 5294
rect 29879 5202 29913 5218
rect 30007 5278 30041 5294
rect 30007 5202 30041 5218
rect 30135 5278 30169 5294
rect 30135 5202 30169 5218
rect 30263 5278 30297 5294
rect 30263 5202 30297 5218
rect 30391 5278 30425 5294
rect 30391 5202 30425 5218
rect 30519 5278 30553 5294
rect 30519 5202 30553 5218
rect 30647 5278 30681 5294
rect 30647 5202 30681 5218
rect 30775 5278 30809 5294
rect 30775 5202 30809 5218
rect 30903 5278 30937 5294
rect 30903 5202 30937 5218
rect 31031 5278 31065 5294
rect 31031 5202 31065 5218
rect 31159 5278 31193 5294
rect 31159 5202 31193 5218
rect 31287 5278 31321 5294
rect 31287 5202 31321 5218
rect 31415 5278 31449 5294
rect 31415 5202 31449 5218
rect 31543 5278 31577 5294
rect 31543 5202 31577 5218
rect 31671 5278 31705 5294
rect 31671 5202 31705 5218
rect 31799 5278 31833 5294
rect 31799 5202 31833 5218
rect 31927 5278 31961 5294
rect 31927 5202 31961 5218
rect 32055 5278 32089 5294
rect 32055 5202 32089 5218
rect 32183 5278 32217 5294
rect 32183 5202 32217 5218
rect 32311 5278 32345 5294
rect 32311 5202 32345 5218
rect 32439 5278 32473 5294
rect 32439 5202 32473 5218
rect 32567 5278 32601 5294
rect 32567 5202 32601 5218
rect 32695 5278 32729 5294
rect 32695 5202 32729 5218
rect 32823 5278 32857 5294
rect 32823 5202 32857 5218
rect 32951 5278 32985 5294
rect 32951 5202 32985 5218
rect 33079 5278 33113 5294
rect 33079 5202 33113 5218
rect 33207 5278 33241 5294
rect 33207 5202 33241 5218
rect 33335 5278 33369 5294
rect 33335 5202 33369 5218
rect 33463 5278 33497 5294
rect 33463 5202 33497 5218
rect 33591 5278 33625 5294
rect 33591 5202 33625 5218
rect 33719 5278 33753 5294
rect 33719 5202 33753 5218
rect 33847 5278 33881 5294
rect 33847 5202 33881 5218
rect 33975 5278 34009 5294
rect 33975 5202 34009 5218
rect 34103 5278 34137 5294
rect 34103 5202 34137 5218
rect 34231 5278 34265 5294
rect 34231 5202 34265 5218
rect 34359 5278 34393 5294
rect 34359 5202 34393 5218
rect 34487 5278 34521 5294
rect 34487 5202 34521 5218
rect 34615 5278 34649 5294
rect 34615 5202 34649 5218
rect 34743 5278 34777 5294
rect 34743 5202 34777 5218
rect 34871 5278 34905 5294
rect 34871 5202 34905 5218
rect 34999 5278 35033 5294
rect 34999 5202 35033 5218
rect 35127 5278 35161 5294
rect 35127 5202 35161 5218
rect 35255 5278 35289 5294
rect 35255 5202 35289 5218
rect 35383 5278 35417 5294
rect 35383 5202 35417 5218
rect 35511 5278 35545 5294
rect 35511 5202 35545 5218
rect 35639 5278 35673 5294
rect 35639 5202 35673 5218
rect 35767 5278 35801 5294
rect 35767 5202 35801 5218
rect 35895 5278 35929 5294
rect 35895 5202 35929 5218
rect 36023 5278 36057 5294
rect 36023 5202 36057 5218
rect 36151 5278 36185 5294
rect 36151 5202 36185 5218
rect 36279 5278 36313 5294
rect 36279 5202 36313 5218
rect 36407 5278 36441 5294
rect 36407 5202 36441 5218
rect 36535 5278 36569 5294
rect 36535 5202 36569 5218
rect 36663 5278 36697 5294
rect 36663 5202 36697 5218
rect 36791 5278 36825 5294
rect 36791 5202 36825 5218
rect 36919 5278 36953 5294
rect 36919 5202 36953 5218
rect 37047 5278 37081 5294
rect 37047 5202 37081 5218
rect 37175 5278 37209 5294
rect 37175 5202 37209 5218
rect 37303 5278 37337 5294
rect 37303 5202 37337 5218
rect 37431 5278 37465 5294
rect 37431 5202 37465 5218
rect 37559 5278 37593 5294
rect 37559 5202 37593 5218
rect -363 5148 37639 5152
rect -363 5110 -319 5148
rect -281 5110 -191 5148
rect -153 5110 609 5148
rect 647 5110 737 5148
rect 775 5110 865 5148
rect 903 5110 1873 5148
rect 1911 5110 2001 5148
rect 2039 5110 2129 5148
rect 2167 5110 2257 5148
rect 2295 5110 2385 5148
rect 2423 5110 3492 5148
rect 3530 5110 3620 5148
rect 3658 5110 3748 5148
rect 3786 5110 3876 5148
rect 3914 5110 4004 5148
rect 4042 5110 4132 5148
rect 4170 5110 4260 5148
rect 4298 5110 4388 5148
rect 4426 5110 4516 5148
rect 4554 5110 8057 5148
rect 8095 5110 8185 5148
rect 8223 5110 8313 5148
rect 8351 5110 8441 5148
rect 8479 5110 8569 5148
rect 8607 5110 8697 5148
rect 8735 5110 8825 5148
rect 8863 5110 8953 5148
rect 8991 5110 9081 5148
rect 9119 5110 9209 5148
rect 9247 5110 9337 5148
rect 9375 5110 9465 5148
rect 9503 5110 9593 5148
rect 9631 5110 9721 5148
rect 9759 5110 9849 5148
rect 9887 5110 9977 5148
rect 10015 5110 10105 5148
rect 10143 5110 15821 5148
rect 15859 5110 15949 5148
rect 15987 5110 16077 5148
rect 16115 5110 16205 5148
rect 16243 5110 16333 5148
rect 16371 5110 16461 5148
rect 16499 5110 16589 5148
rect 16627 5110 16717 5148
rect 16755 5110 16845 5148
rect 16883 5110 16973 5148
rect 17011 5110 17101 5148
rect 17139 5110 17229 5148
rect 17267 5110 17357 5148
rect 17395 5110 17485 5148
rect 17523 5110 17613 5148
rect 17651 5110 17741 5148
rect 17779 5110 17869 5148
rect 17907 5110 17997 5148
rect 18035 5110 18125 5148
rect 18163 5110 18253 5148
rect 18291 5110 18381 5148
rect 18419 5110 18509 5148
rect 18547 5110 18637 5148
rect 18675 5110 18765 5148
rect 18803 5110 18893 5148
rect 18931 5110 19021 5148
rect 19059 5110 19149 5148
rect 19187 5110 19277 5148
rect 19315 5110 19405 5148
rect 19443 5110 19533 5148
rect 19571 5110 19661 5148
rect 19699 5110 19789 5148
rect 19827 5110 19917 5148
rect 19955 5110 29365 5148
rect 29403 5110 29493 5148
rect 29531 5110 29621 5148
rect 29659 5110 29749 5148
rect 29787 5110 29877 5148
rect 29915 5110 30005 5148
rect 30043 5110 30133 5148
rect 30171 5110 30261 5148
rect 30299 5110 30389 5148
rect 30427 5110 30517 5148
rect 30555 5110 30645 5148
rect 30683 5110 30773 5148
rect 30811 5110 30901 5148
rect 30939 5110 31029 5148
rect 31067 5110 31157 5148
rect 31195 5110 31285 5148
rect 31323 5110 31413 5148
rect 31451 5110 31541 5148
rect 31579 5110 31669 5148
rect 31707 5110 31797 5148
rect 31835 5110 31925 5148
rect 31963 5110 32053 5148
rect 32091 5110 32181 5148
rect 32219 5110 32309 5148
rect 32347 5110 32437 5148
rect 32475 5110 32565 5148
rect 32603 5110 32693 5148
rect 32731 5110 32821 5148
rect 32859 5110 32949 5148
rect 32987 5110 33077 5148
rect 33115 5110 33205 5148
rect 33243 5110 33333 5148
rect 33371 5110 33461 5148
rect 33499 5110 33589 5148
rect 33627 5110 33717 5148
rect 33755 5110 33845 5148
rect 33883 5110 33973 5148
rect 34011 5110 34101 5148
rect 34139 5110 34229 5148
rect 34267 5110 34357 5148
rect 34395 5110 34485 5148
rect 34523 5110 34613 5148
rect 34651 5110 34741 5148
rect 34779 5110 34869 5148
rect 34907 5110 34997 5148
rect 35035 5110 35125 5148
rect 35163 5110 35253 5148
rect 35291 5110 35381 5148
rect 35419 5110 35509 5148
rect 35547 5110 35637 5148
rect 35675 5110 35765 5148
rect 35803 5110 35893 5148
rect 35931 5110 36021 5148
rect 36059 5110 36149 5148
rect 36187 5110 36277 5148
rect 36315 5110 36405 5148
rect 36443 5110 36533 5148
rect 36571 5110 36661 5148
rect 36699 5110 36789 5148
rect 36827 5110 36917 5148
rect 36955 5110 37045 5148
rect 37083 5110 37173 5148
rect 37211 5110 37301 5148
rect 37339 5110 37429 5148
rect 37467 5110 37557 5148
rect 37595 5110 37639 5148
rect -363 5106 37639 5110
<< viali >>
rect -319 6270 -281 6308
rect -191 6270 -153 6308
rect 481 6270 519 6308
rect 609 6270 647 6308
rect 737 6270 775 6308
rect 1361 6270 1399 6308
rect 1489 6270 1527 6308
rect 1617 6270 1655 6308
rect 1745 6270 1783 6308
rect 1873 6270 1911 6308
rect 2980 6270 3018 6308
rect 3108 6270 3146 6308
rect 3236 6270 3274 6308
rect 3364 6270 3402 6308
rect 3492 6270 3530 6308
rect 3620 6270 3658 6308
rect 3748 6270 3786 6308
rect 3876 6270 3914 6308
rect 4004 6270 4042 6308
rect 5473 6270 5511 6308
rect 5601 6270 5639 6308
rect 5729 6270 5767 6308
rect 5857 6270 5895 6308
rect 5985 6270 6023 6308
rect 6113 6270 6151 6308
rect 6241 6270 6279 6308
rect 6369 6270 6407 6308
rect 6497 6270 6535 6308
rect 6625 6270 6663 6308
rect 6753 6270 6791 6308
rect 6881 6270 6919 6308
rect 7009 6270 7047 6308
rect 7137 6270 7175 6308
rect 7265 6270 7303 6308
rect 7393 6270 7431 6308
rect 7521 6270 7559 6308
rect 10560 6270 10598 6308
rect 10688 6270 10726 6308
rect 10816 6270 10854 6308
rect 10944 6270 10982 6308
rect 11072 6270 11110 6308
rect 11200 6270 11238 6308
rect 11328 6270 11366 6308
rect 11456 6270 11494 6308
rect 11584 6270 11622 6308
rect 11712 6270 11750 6308
rect 11840 6270 11878 6308
rect 11968 6270 12006 6308
rect 12096 6270 12134 6308
rect 12224 6270 12262 6308
rect 12352 6270 12390 6308
rect 12480 6270 12518 6308
rect 12608 6270 12646 6308
rect 12736 6270 12774 6308
rect 12864 6270 12902 6308
rect 12992 6270 13030 6308
rect 13120 6270 13158 6308
rect 13248 6270 13286 6308
rect 13376 6270 13414 6308
rect 13504 6270 13542 6308
rect 13632 6270 13670 6308
rect 13760 6270 13798 6308
rect 13888 6270 13926 6308
rect 14016 6270 14054 6308
rect 14144 6270 14182 6308
rect 14272 6270 14310 6308
rect 14400 6270 14438 6308
rect 14528 6270 14566 6308
rect 14656 6270 14694 6308
rect 20397 6270 20435 6308
rect 20525 6270 20563 6308
rect 20653 6270 20691 6308
rect 20781 6270 20819 6308
rect 20909 6270 20947 6308
rect 21037 6270 21075 6308
rect 21165 6270 21203 6308
rect 21293 6270 21331 6308
rect 21421 6270 21459 6308
rect 21549 6270 21587 6308
rect 21677 6270 21715 6308
rect 21805 6270 21843 6308
rect 21933 6270 21971 6308
rect 22061 6270 22099 6308
rect 22189 6270 22227 6308
rect 22317 6270 22355 6308
rect 22445 6270 22483 6308
rect 22573 6270 22611 6308
rect 22701 6270 22739 6308
rect 22829 6270 22867 6308
rect 22957 6270 22995 6308
rect 23085 6270 23123 6308
rect 23213 6270 23251 6308
rect 23341 6270 23379 6308
rect 23469 6270 23507 6308
rect 23597 6270 23635 6308
rect 23725 6270 23763 6308
rect 23853 6270 23891 6308
rect 23981 6270 24019 6308
rect 24109 6270 24147 6308
rect 24237 6270 24275 6308
rect 24365 6270 24403 6308
rect 24493 6270 24531 6308
rect 24621 6270 24659 6308
rect 24749 6270 24787 6308
rect 24877 6270 24915 6308
rect 25005 6270 25043 6308
rect 25133 6270 25171 6308
rect 25261 6270 25299 6308
rect 25389 6270 25427 6308
rect 25517 6270 25555 6308
rect 25645 6270 25683 6308
rect 25773 6270 25811 6308
rect 25901 6270 25939 6308
rect 26029 6270 26067 6308
rect 26157 6270 26195 6308
rect 26285 6270 26323 6308
rect 26413 6270 26451 6308
rect 26541 6270 26579 6308
rect 26669 6270 26707 6308
rect 26797 6270 26835 6308
rect 26925 6270 26963 6308
rect 27053 6270 27091 6308
rect 27181 6270 27219 6308
rect 27309 6270 27347 6308
rect 27437 6270 27475 6308
rect 27565 6270 27603 6308
rect 27693 6270 27731 6308
rect 27821 6270 27859 6308
rect 27949 6270 27987 6308
rect 28077 6270 28115 6308
rect 28205 6270 28243 6308
rect 28333 6270 28371 6308
rect 28461 6270 28499 6308
rect 28589 6270 28627 6308
rect -317 6140 -283 6200
rect -189 6140 -155 6200
rect 483 6140 517 6200
rect 611 6140 645 6200
rect 739 6140 773 6200
rect 1363 6140 1397 6200
rect 1491 6140 1525 6200
rect 1619 6140 1653 6200
rect 1747 6140 1781 6200
rect 1875 6140 1909 6200
rect 2982 6140 3016 6200
rect 3110 6140 3144 6200
rect 3238 6140 3272 6200
rect 3366 6140 3400 6200
rect 3494 6140 3528 6200
rect 3622 6140 3656 6200
rect 3750 6140 3784 6200
rect 3878 6140 3912 6200
rect 4006 6140 4040 6200
rect 4118 6157 4163 6161
rect 4118 6123 4123 6157
rect 4123 6123 4157 6157
rect 4157 6123 4163 6157
rect 4118 6118 4163 6123
rect 5475 6140 5509 6200
rect 5603 6140 5637 6200
rect 5731 6140 5765 6200
rect 5859 6140 5893 6200
rect 5987 6140 6021 6200
rect 6115 6140 6149 6200
rect 6243 6140 6277 6200
rect 6371 6140 6405 6200
rect 6499 6140 6533 6200
rect 6627 6140 6661 6200
rect 6755 6140 6789 6200
rect 6883 6140 6917 6200
rect 7011 6140 7045 6200
rect 7139 6140 7173 6200
rect 7267 6140 7301 6200
rect 7395 6140 7429 6200
rect 7523 6140 7557 6200
rect 7695 6154 7740 6158
rect 7695 6120 7700 6154
rect 7700 6120 7734 6154
rect 7734 6120 7740 6154
rect 7695 6115 7740 6120
rect 10562 6140 10596 6200
rect 10690 6140 10724 6200
rect 10818 6140 10852 6200
rect 10946 6140 10980 6200
rect 11074 6140 11108 6200
rect 11202 6140 11236 6200
rect 11330 6140 11364 6200
rect 11458 6140 11492 6200
rect 11586 6140 11620 6200
rect 11714 6140 11748 6200
rect 11842 6140 11876 6200
rect 11970 6140 12004 6200
rect 12098 6140 12132 6200
rect 12226 6140 12260 6200
rect 12354 6140 12388 6200
rect 12482 6140 12516 6200
rect 12610 6140 12644 6200
rect 12738 6140 12772 6200
rect 12866 6140 12900 6200
rect 12994 6140 13028 6200
rect 13122 6140 13156 6200
rect 13250 6140 13284 6200
rect 13378 6140 13412 6200
rect 13506 6140 13540 6200
rect 13634 6140 13668 6200
rect 13762 6140 13796 6200
rect 13890 6140 13924 6200
rect 14018 6140 14052 6200
rect 14146 6140 14180 6200
rect 14274 6140 14308 6200
rect 14402 6140 14436 6200
rect 14530 6140 14564 6200
rect 14658 6140 14692 6200
rect 20399 6140 20433 6200
rect 20527 6140 20561 6200
rect 20655 6140 20689 6200
rect 20783 6140 20817 6200
rect 20911 6140 20945 6200
rect 21039 6140 21073 6200
rect 21167 6140 21201 6200
rect 21295 6140 21329 6200
rect 21423 6140 21457 6200
rect 21551 6140 21585 6200
rect 21679 6140 21713 6200
rect 21807 6140 21841 6200
rect 21935 6140 21969 6200
rect 22063 6140 22097 6200
rect 22191 6140 22225 6200
rect 22319 6140 22353 6200
rect 22447 6140 22481 6200
rect 22575 6140 22609 6200
rect 22703 6140 22737 6200
rect 22831 6140 22865 6200
rect 22959 6140 22993 6200
rect 23087 6140 23121 6200
rect 23215 6140 23249 6200
rect 23343 6140 23377 6200
rect 23471 6140 23505 6200
rect 23599 6140 23633 6200
rect 23727 6140 23761 6200
rect 23855 6140 23889 6200
rect 23983 6140 24017 6200
rect 24111 6140 24145 6200
rect 24239 6140 24273 6200
rect 24367 6140 24401 6200
rect 24495 6140 24529 6200
rect 24623 6140 24657 6200
rect 24751 6140 24785 6200
rect 24879 6140 24913 6200
rect 25007 6140 25041 6200
rect 25135 6140 25169 6200
rect 25263 6140 25297 6200
rect 25391 6140 25425 6200
rect 25519 6140 25553 6200
rect 25647 6140 25681 6200
rect 25775 6140 25809 6200
rect 25903 6140 25937 6200
rect 26031 6140 26065 6200
rect 26159 6140 26193 6200
rect 26287 6140 26321 6200
rect 26415 6140 26449 6200
rect 26543 6140 26577 6200
rect 26671 6140 26705 6200
rect 26799 6140 26833 6200
rect 26927 6140 26961 6200
rect 27055 6140 27089 6200
rect 27183 6140 27217 6200
rect 27311 6140 27345 6200
rect 27439 6140 27473 6200
rect 27567 6140 27601 6200
rect 27695 6140 27729 6200
rect 27823 6140 27857 6200
rect 27951 6140 27985 6200
rect 28079 6140 28113 6200
rect 28207 6140 28241 6200
rect 28335 6140 28369 6200
rect 28463 6140 28497 6200
rect 28591 6140 28625 6200
rect -290 6078 -245 6082
rect -290 6044 -285 6078
rect -285 6044 -251 6078
rect -251 6044 -245 6078
rect -290 6039 -245 6044
rect 760 6078 805 6082
rect 760 6044 765 6078
rect 765 6044 799 6078
rect 799 6044 805 6078
rect 760 6039 805 6044
rect 1980 6067 2025 6071
rect 1980 6033 1985 6067
rect 1985 6033 2019 6067
rect 2019 6033 2025 6067
rect 1980 6028 2025 6033
rect 14710 6082 14755 6086
rect 14710 6048 14715 6082
rect 14715 6048 14749 6082
rect 14749 6048 14755 6082
rect 14710 6043 14755 6048
rect 28737 6102 28782 6107
rect 28737 6068 28743 6102
rect 28743 6068 28777 6102
rect 28777 6068 28782 6102
rect 28737 6064 28782 6068
rect -317 5840 -283 5984
rect -189 5840 -155 5984
rect 483 5840 517 5984
rect 611 5840 645 5984
rect 739 5840 773 5984
rect 1363 5840 1397 5984
rect 1491 5840 1525 5984
rect 1619 5840 1653 5984
rect 1747 5840 1781 5984
rect 1875 5840 1909 5984
rect 2982 5840 3016 5984
rect 3110 5840 3144 5984
rect 3238 5840 3272 5984
rect 3366 5840 3400 5984
rect 3494 5840 3528 5984
rect 3622 5840 3656 5984
rect 3750 5840 3784 5984
rect 3878 5840 3912 5984
rect 4006 5840 4040 5984
rect 5475 5840 5509 5984
rect 5603 5840 5637 5984
rect 5731 5840 5765 5984
rect 5859 5840 5893 5984
rect 5987 5840 6021 5984
rect 6115 5840 6149 5984
rect 6243 5840 6277 5984
rect 6371 5840 6405 5984
rect 6499 5840 6533 5984
rect 6627 5840 6661 5984
rect 6755 5840 6789 5984
rect 6883 5840 6917 5984
rect 7011 5840 7045 5984
rect 7139 5840 7173 5984
rect 7267 5840 7301 5984
rect 7395 5840 7429 5984
rect 7523 5840 7557 5984
rect 10562 5840 10596 5984
rect 10690 5840 10724 5984
rect 10818 5840 10852 5984
rect 10946 5840 10980 5984
rect 11074 5840 11108 5984
rect 11202 5840 11236 5984
rect 11330 5840 11364 5984
rect 11458 5840 11492 5984
rect 11586 5840 11620 5984
rect 11714 5840 11748 5984
rect 11842 5840 11876 5984
rect 11970 5840 12004 5984
rect 12098 5840 12132 5984
rect 12226 5840 12260 5984
rect 12354 5840 12388 5984
rect 12482 5840 12516 5984
rect 12610 5840 12644 5984
rect 12738 5840 12772 5984
rect 12866 5840 12900 5984
rect 12994 5840 13028 5984
rect 13122 5840 13156 5984
rect 13250 5840 13284 5984
rect 13378 5840 13412 5984
rect 13506 5840 13540 5984
rect 13634 5840 13668 5984
rect 13762 5840 13796 5984
rect 13890 5840 13924 5984
rect 14018 5840 14052 5984
rect 14146 5840 14180 5984
rect 14274 5840 14308 5984
rect 14402 5840 14436 5984
rect 14530 5840 14564 5984
rect 14658 5840 14692 5984
rect 20399 5840 20433 5984
rect 20527 5840 20561 5984
rect 20655 5840 20689 5984
rect 20783 5840 20817 5984
rect 20911 5840 20945 5984
rect 21039 5840 21073 5984
rect 21167 5840 21201 5984
rect 21295 5840 21329 5984
rect 21423 5840 21457 5984
rect 21551 5840 21585 5984
rect 21679 5840 21713 5984
rect 21807 5840 21841 5984
rect 21935 5840 21969 5984
rect 22063 5840 22097 5984
rect 22191 5840 22225 5984
rect 22319 5840 22353 5984
rect 22447 5840 22481 5984
rect 22575 5840 22609 5984
rect 22703 5840 22737 5984
rect 22831 5840 22865 5984
rect 22959 5840 22993 5984
rect 23087 5840 23121 5984
rect 23215 5840 23249 5984
rect 23343 5840 23377 5984
rect 23471 5840 23505 5984
rect 23599 5840 23633 5984
rect 23727 5840 23761 5984
rect 23855 5840 23889 5984
rect 23983 5840 24017 5984
rect 24111 5840 24145 5984
rect 24239 5840 24273 5984
rect 24367 5840 24401 5984
rect 24495 5840 24529 5984
rect 24623 5840 24657 5984
rect 24751 5840 24785 5984
rect 24879 5840 24913 5984
rect 25007 5840 25041 5984
rect 25135 5840 25169 5984
rect 25263 5840 25297 5984
rect 25391 5840 25425 5984
rect 25519 5840 25553 5984
rect 25647 5840 25681 5984
rect 25775 5840 25809 5984
rect 25903 5840 25937 5984
rect 26031 5840 26065 5984
rect 26159 5840 26193 5984
rect 26287 5840 26321 5984
rect 26415 5840 26449 5984
rect 26543 5840 26577 5984
rect 26671 5840 26705 5984
rect 26799 5840 26833 5984
rect 26927 5840 26961 5984
rect 27055 5840 27089 5984
rect 27183 5840 27217 5984
rect 27311 5840 27345 5984
rect 27439 5840 27473 5984
rect 27567 5840 27601 5984
rect 27695 5840 27729 5984
rect 27823 5840 27857 5984
rect 27951 5840 27985 5984
rect 28079 5840 28113 5984
rect 28207 5840 28241 5984
rect 28335 5840 28369 5984
rect 28463 5840 28497 5984
rect 28591 5840 28625 5984
rect -319 5690 -281 5728
rect -191 5690 -153 5728
rect 481 5690 519 5728
rect 609 5690 647 5728
rect 737 5690 775 5728
rect 865 5690 903 5728
rect 1361 5690 1399 5728
rect 1489 5690 1527 5728
rect 1617 5690 1655 5728
rect 1745 5690 1783 5728
rect 1873 5690 1911 5728
rect 2001 5690 2039 5728
rect 2129 5690 2167 5728
rect 2257 5690 2295 5728
rect 2385 5690 2423 5728
rect 2980 5690 3018 5728
rect 3108 5690 3146 5728
rect 3236 5690 3274 5728
rect 3364 5690 3402 5728
rect 3492 5690 3530 5728
rect 3620 5690 3658 5728
rect 3748 5690 3786 5728
rect 3876 5690 3914 5728
rect 4004 5690 4042 5728
rect 4132 5690 4170 5728
rect 4260 5690 4298 5728
rect 4388 5690 4426 5728
rect 4516 5690 4554 5728
rect 5473 5690 5511 5728
rect 5601 5690 5639 5728
rect 5729 5690 5767 5728
rect 5857 5690 5895 5728
rect 5985 5690 6023 5728
rect 6113 5690 6151 5728
rect 6241 5690 6279 5728
rect 6369 5690 6407 5728
rect 6497 5690 6535 5728
rect 6625 5690 6663 5728
rect 6753 5690 6791 5728
rect 6881 5690 6919 5728
rect 7009 5690 7047 5728
rect 7137 5690 7175 5728
rect 7265 5690 7303 5728
rect 7393 5690 7431 5728
rect 7521 5690 7559 5728
rect 8057 5690 8095 5728
rect 8185 5690 8223 5728
rect 8313 5690 8351 5728
rect 8441 5690 8479 5728
rect 8569 5690 8607 5728
rect 8697 5690 8735 5728
rect 8825 5690 8863 5728
rect 8953 5690 8991 5728
rect 9081 5690 9119 5728
rect 9209 5690 9247 5728
rect 9337 5690 9375 5728
rect 9465 5690 9503 5728
rect 9593 5690 9631 5728
rect 9721 5690 9759 5728
rect 9849 5690 9887 5728
rect 9977 5690 10015 5728
rect 10105 5690 10143 5728
rect 10560 5690 10598 5728
rect 10688 5690 10726 5728
rect 10816 5690 10854 5728
rect 10944 5690 10982 5728
rect 11072 5690 11110 5728
rect 11200 5690 11238 5728
rect 11328 5690 11366 5728
rect 11456 5690 11494 5728
rect 11584 5690 11622 5728
rect 11712 5690 11750 5728
rect 11840 5690 11878 5728
rect 11968 5690 12006 5728
rect 12096 5690 12134 5728
rect 12224 5690 12262 5728
rect 12352 5690 12390 5728
rect 12480 5690 12518 5728
rect 12608 5690 12646 5728
rect 12736 5690 12774 5728
rect 12864 5690 12902 5728
rect 12992 5690 13030 5728
rect 13120 5690 13158 5728
rect 13248 5690 13286 5728
rect 13376 5690 13414 5728
rect 13504 5690 13542 5728
rect 13632 5690 13670 5728
rect 13760 5690 13798 5728
rect 13888 5690 13926 5728
rect 14016 5690 14054 5728
rect 14144 5690 14182 5728
rect 14272 5690 14310 5728
rect 14400 5690 14438 5728
rect 14528 5690 14566 5728
rect 14656 5690 14694 5728
rect 15821 5690 15859 5728
rect 15949 5690 15987 5728
rect 16077 5690 16115 5728
rect 16205 5690 16243 5728
rect 16333 5690 16371 5728
rect 16461 5690 16499 5728
rect 16589 5690 16627 5728
rect 16717 5690 16755 5728
rect 16845 5690 16883 5728
rect 16973 5690 17011 5728
rect 17101 5690 17139 5728
rect 17229 5690 17267 5728
rect 17357 5690 17395 5728
rect 17485 5690 17523 5728
rect 17613 5690 17651 5728
rect 17741 5690 17779 5728
rect 17869 5690 17907 5728
rect 17997 5690 18035 5728
rect 18125 5690 18163 5728
rect 18253 5690 18291 5728
rect 18381 5690 18419 5728
rect 18509 5690 18547 5728
rect 18637 5690 18675 5728
rect 18765 5690 18803 5728
rect 18893 5690 18931 5728
rect 19021 5690 19059 5728
rect 19149 5690 19187 5728
rect 19277 5690 19315 5728
rect 19405 5690 19443 5728
rect 19533 5690 19571 5728
rect 19661 5690 19699 5728
rect 19789 5690 19827 5728
rect 19917 5690 19955 5728
rect 20397 5690 20435 5728
rect 20525 5690 20563 5728
rect 20653 5690 20691 5728
rect 20781 5690 20819 5728
rect 20909 5690 20947 5728
rect 21037 5690 21075 5728
rect 21165 5690 21203 5728
rect 21293 5690 21331 5728
rect 21421 5690 21459 5728
rect 21549 5690 21587 5728
rect 21677 5690 21715 5728
rect 21805 5690 21843 5728
rect 21933 5690 21971 5728
rect 22061 5690 22099 5728
rect 22189 5690 22227 5728
rect 22317 5690 22355 5728
rect 22445 5690 22483 5728
rect 22573 5690 22611 5728
rect 22701 5690 22739 5728
rect 22829 5690 22867 5728
rect 22957 5690 22995 5728
rect 23085 5690 23123 5728
rect 23213 5690 23251 5728
rect 23341 5690 23379 5728
rect 23469 5690 23507 5728
rect 23597 5690 23635 5728
rect 23725 5690 23763 5728
rect 23853 5690 23891 5728
rect 23981 5690 24019 5728
rect 24109 5690 24147 5728
rect 24237 5690 24275 5728
rect 24365 5690 24403 5728
rect 24493 5690 24531 5728
rect 24621 5690 24659 5728
rect 24749 5690 24787 5728
rect 24877 5690 24915 5728
rect 25005 5690 25043 5728
rect 25133 5690 25171 5728
rect 25261 5690 25299 5728
rect 25389 5690 25427 5728
rect 25517 5690 25555 5728
rect 25645 5690 25683 5728
rect 25773 5690 25811 5728
rect 25901 5690 25939 5728
rect 26029 5690 26067 5728
rect 26157 5690 26195 5728
rect 26285 5690 26323 5728
rect 26413 5690 26451 5728
rect 26541 5690 26579 5728
rect 26669 5690 26707 5728
rect 26797 5690 26835 5728
rect 26925 5690 26963 5728
rect 27053 5690 27091 5728
rect 27181 5690 27219 5728
rect 27309 5690 27347 5728
rect 27437 5690 27475 5728
rect 27565 5690 27603 5728
rect 27693 5690 27731 5728
rect 27821 5690 27859 5728
rect 27949 5690 27987 5728
rect 28077 5690 28115 5728
rect 28205 5690 28243 5728
rect 28333 5690 28371 5728
rect 28461 5690 28499 5728
rect 28589 5690 28627 5728
rect 29365 5690 29403 5728
rect 29493 5690 29531 5728
rect 29621 5690 29659 5728
rect 29749 5690 29787 5728
rect 29877 5690 29915 5728
rect 30005 5690 30043 5728
rect 30133 5690 30171 5728
rect 30261 5690 30299 5728
rect 30389 5690 30427 5728
rect 30517 5690 30555 5728
rect 30645 5690 30683 5728
rect 30773 5690 30811 5728
rect 30901 5690 30939 5728
rect 31029 5690 31067 5728
rect 31157 5690 31195 5728
rect 31285 5690 31323 5728
rect 31413 5690 31451 5728
rect 31541 5690 31579 5728
rect 31669 5690 31707 5728
rect 31797 5690 31835 5728
rect 31925 5690 31963 5728
rect 32053 5690 32091 5728
rect 32181 5690 32219 5728
rect 32309 5690 32347 5728
rect 32437 5690 32475 5728
rect 32565 5690 32603 5728
rect 32693 5690 32731 5728
rect 32821 5690 32859 5728
rect 32949 5690 32987 5728
rect 33077 5690 33115 5728
rect 33205 5690 33243 5728
rect 33333 5690 33371 5728
rect 33461 5690 33499 5728
rect 33589 5690 33627 5728
rect 33717 5690 33755 5728
rect 33845 5690 33883 5728
rect 33973 5690 34011 5728
rect 34101 5690 34139 5728
rect 34229 5690 34267 5728
rect 34357 5690 34395 5728
rect 34485 5690 34523 5728
rect 34613 5690 34651 5728
rect 34741 5690 34779 5728
rect 34869 5690 34907 5728
rect 34997 5690 35035 5728
rect 35125 5690 35163 5728
rect 35253 5690 35291 5728
rect 35381 5690 35419 5728
rect 35509 5690 35547 5728
rect 35637 5690 35675 5728
rect 35765 5690 35803 5728
rect 35893 5690 35931 5728
rect 36021 5690 36059 5728
rect 36149 5690 36187 5728
rect 36277 5690 36315 5728
rect 36405 5690 36443 5728
rect 36533 5690 36571 5728
rect 36661 5690 36699 5728
rect 36789 5690 36827 5728
rect 36917 5690 36955 5728
rect 37045 5690 37083 5728
rect 37173 5690 37211 5728
rect 37301 5690 37339 5728
rect 37429 5690 37467 5728
rect 37557 5690 37595 5728
rect -317 5434 -283 5578
rect -189 5434 -155 5578
rect 611 5434 645 5578
rect 739 5434 773 5578
rect 867 5434 901 5578
rect 972 5435 1017 5439
rect 972 5401 977 5435
rect 977 5401 1011 5435
rect 1011 5401 1017 5435
rect 972 5396 1017 5401
rect 1875 5434 1909 5578
rect 2003 5434 2037 5578
rect 2131 5434 2165 5578
rect 2259 5434 2293 5578
rect 2387 5434 2421 5578
rect 2501 5435 2546 5439
rect 2501 5401 2506 5435
rect 2506 5401 2540 5435
rect 2540 5401 2546 5435
rect 2501 5396 2546 5401
rect 3494 5434 3528 5578
rect 3622 5434 3656 5578
rect 3750 5434 3784 5578
rect 3878 5434 3912 5578
rect 4006 5434 4040 5578
rect 4134 5434 4168 5578
rect 4262 5434 4296 5578
rect 4390 5434 4424 5578
rect 4518 5434 4552 5578
rect 4672 5444 4717 5448
rect 4672 5410 4677 5444
rect 4677 5410 4711 5444
rect 4711 5410 4717 5444
rect 4672 5405 4717 5410
rect 8059 5434 8093 5578
rect 7930 5429 7975 5433
rect 7930 5395 7935 5429
rect 7935 5395 7969 5429
rect 7969 5395 7975 5429
rect 7930 5390 7975 5395
rect 8187 5434 8221 5578
rect 8315 5434 8349 5578
rect 8443 5434 8477 5578
rect 8571 5434 8605 5578
rect 8699 5434 8733 5578
rect 8827 5434 8861 5578
rect 8955 5434 8989 5578
rect 9083 5434 9117 5578
rect 9211 5434 9245 5578
rect 9339 5434 9373 5578
rect 9467 5434 9501 5578
rect 9595 5434 9629 5578
rect 9723 5434 9757 5578
rect 9851 5434 9885 5578
rect 9979 5434 10013 5578
rect 10107 5434 10141 5578
rect 15823 5434 15857 5578
rect 15951 5434 15985 5578
rect 16079 5434 16113 5578
rect 16207 5434 16241 5578
rect 16335 5434 16369 5578
rect 16463 5434 16497 5578
rect 16591 5434 16625 5578
rect 16719 5434 16753 5578
rect 16847 5434 16881 5578
rect 16975 5434 17009 5578
rect 17103 5434 17137 5578
rect 17231 5434 17265 5578
rect 17359 5434 17393 5578
rect 17487 5434 17521 5578
rect 17615 5434 17649 5578
rect 17743 5434 17777 5578
rect 17871 5434 17905 5578
rect 17999 5434 18033 5578
rect 18127 5434 18161 5578
rect 18255 5434 18289 5578
rect 18383 5434 18417 5578
rect 18511 5434 18545 5578
rect 18639 5434 18673 5578
rect 18767 5434 18801 5578
rect 18895 5434 18929 5578
rect 19023 5434 19057 5578
rect 19151 5434 19185 5578
rect 19279 5434 19313 5578
rect 19407 5434 19441 5578
rect 19535 5434 19569 5578
rect 19663 5434 19697 5578
rect 19791 5434 19825 5578
rect 19919 5434 19953 5578
rect 29367 5434 29401 5578
rect 29495 5434 29529 5578
rect 29623 5434 29657 5578
rect 29751 5434 29785 5578
rect 29879 5434 29913 5578
rect 30007 5434 30041 5578
rect 30135 5434 30169 5578
rect 30263 5434 30297 5578
rect 30391 5434 30425 5578
rect 30519 5434 30553 5578
rect 30647 5434 30681 5578
rect 30775 5434 30809 5578
rect 30903 5434 30937 5578
rect 31031 5434 31065 5578
rect 31159 5434 31193 5578
rect 31287 5434 31321 5578
rect 31415 5434 31449 5578
rect 31543 5434 31577 5578
rect 31671 5434 31705 5578
rect 31799 5434 31833 5578
rect 31927 5434 31961 5578
rect 32055 5434 32089 5578
rect 32183 5434 32217 5578
rect 32311 5434 32345 5578
rect 32439 5434 32473 5578
rect 32567 5434 32601 5578
rect 32695 5434 32729 5578
rect 32823 5434 32857 5578
rect 32951 5434 32985 5578
rect 33079 5434 33113 5578
rect 33207 5434 33241 5578
rect 33335 5434 33369 5578
rect 33463 5434 33497 5578
rect 33591 5434 33625 5578
rect 33719 5434 33753 5578
rect 33847 5434 33881 5578
rect 33975 5434 34009 5578
rect 34103 5434 34137 5578
rect 34231 5434 34265 5578
rect 34359 5434 34393 5578
rect 34487 5434 34521 5578
rect 34615 5434 34649 5578
rect 34743 5434 34777 5578
rect 34871 5434 34905 5578
rect 34999 5434 35033 5578
rect 35127 5434 35161 5578
rect 35255 5434 35289 5578
rect 35383 5434 35417 5578
rect 35511 5434 35545 5578
rect 35639 5434 35673 5578
rect 35767 5434 35801 5578
rect 35895 5434 35929 5578
rect 36023 5434 36057 5578
rect 36151 5434 36185 5578
rect 36279 5434 36313 5578
rect 36407 5434 36441 5578
rect 36535 5434 36569 5578
rect 36663 5434 36697 5578
rect 36791 5434 36825 5578
rect 36919 5434 36953 5578
rect 37047 5434 37081 5578
rect 37175 5434 37209 5578
rect 37303 5434 37337 5578
rect 37431 5434 37465 5578
rect 37559 5434 37593 5578
rect -377 5372 -332 5376
rect -377 5338 -372 5372
rect -372 5338 -338 5372
rect -338 5338 -332 5372
rect -377 5333 -332 5338
rect 15699 5398 15744 5402
rect 15699 5364 15704 5398
rect 15704 5364 15738 5398
rect 15738 5364 15744 5398
rect 15699 5359 15744 5364
rect -317 5218 -283 5278
rect -189 5218 -155 5278
rect 611 5218 645 5278
rect 739 5218 773 5278
rect 867 5218 901 5278
rect 1875 5218 1909 5278
rect 2003 5218 2037 5278
rect 2131 5218 2165 5278
rect 2259 5218 2293 5278
rect 2387 5218 2421 5278
rect 3494 5218 3528 5278
rect 3622 5218 3656 5278
rect 3750 5218 3784 5278
rect 3878 5218 3912 5278
rect 4006 5218 4040 5278
rect 4134 5218 4168 5278
rect 4262 5218 4296 5278
rect 4390 5218 4424 5278
rect 4518 5218 4552 5278
rect 8059 5218 8093 5278
rect 8187 5218 8221 5278
rect 8315 5218 8349 5278
rect 8443 5218 8477 5278
rect 8571 5218 8605 5278
rect 8699 5218 8733 5278
rect 8827 5218 8861 5278
rect 8955 5218 8989 5278
rect 9083 5218 9117 5278
rect 9211 5218 9245 5278
rect 9339 5218 9373 5278
rect 9467 5218 9501 5278
rect 9595 5218 9629 5278
rect 9723 5218 9757 5278
rect 9851 5218 9885 5278
rect 9979 5218 10013 5278
rect 10107 5218 10141 5278
rect 15823 5218 15857 5278
rect 15951 5218 15985 5278
rect 16079 5218 16113 5278
rect 16207 5218 16241 5278
rect 16335 5218 16369 5278
rect 16463 5218 16497 5278
rect 16591 5218 16625 5278
rect 16719 5218 16753 5278
rect 16847 5218 16881 5278
rect 16975 5218 17009 5278
rect 17103 5218 17137 5278
rect 17231 5218 17265 5278
rect 17359 5218 17393 5278
rect 17487 5218 17521 5278
rect 17615 5218 17649 5278
rect 17743 5218 17777 5278
rect 17871 5218 17905 5278
rect 17999 5218 18033 5278
rect 18127 5218 18161 5278
rect 18255 5218 18289 5278
rect 18383 5218 18417 5278
rect 18511 5218 18545 5278
rect 18639 5218 18673 5278
rect 18767 5218 18801 5278
rect 18895 5218 18929 5278
rect 19023 5218 19057 5278
rect 19151 5218 19185 5278
rect 19279 5218 19313 5278
rect 19407 5218 19441 5278
rect 19535 5218 19569 5278
rect 19663 5218 19697 5278
rect 19791 5218 19825 5278
rect 19919 5218 19953 5278
rect 29367 5218 29401 5278
rect 29495 5218 29529 5278
rect 29623 5218 29657 5278
rect 29751 5218 29785 5278
rect 29879 5218 29913 5278
rect 30007 5218 30041 5278
rect 30135 5218 30169 5278
rect 30263 5218 30297 5278
rect 30391 5218 30425 5278
rect 30519 5218 30553 5278
rect 30647 5218 30681 5278
rect 30775 5218 30809 5278
rect 30903 5218 30937 5278
rect 31031 5218 31065 5278
rect 31159 5218 31193 5278
rect 31287 5218 31321 5278
rect 31415 5218 31449 5278
rect 31543 5218 31577 5278
rect 31671 5218 31705 5278
rect 31799 5218 31833 5278
rect 31927 5218 31961 5278
rect 32055 5218 32089 5278
rect 32183 5218 32217 5278
rect 32311 5218 32345 5278
rect 32439 5218 32473 5278
rect 32567 5218 32601 5278
rect 32695 5218 32729 5278
rect 32823 5218 32857 5278
rect 32951 5218 32985 5278
rect 33079 5218 33113 5278
rect 33207 5218 33241 5278
rect 33335 5218 33369 5278
rect 33463 5218 33497 5278
rect 33591 5218 33625 5278
rect 33719 5218 33753 5278
rect 33847 5218 33881 5278
rect 33975 5218 34009 5278
rect 34103 5218 34137 5278
rect 34231 5218 34265 5278
rect 34359 5218 34393 5278
rect 34487 5218 34521 5278
rect 34615 5218 34649 5278
rect 34743 5218 34777 5278
rect 34871 5218 34905 5278
rect 34999 5218 35033 5278
rect 35127 5218 35161 5278
rect 35255 5218 35289 5278
rect 35383 5218 35417 5278
rect 35511 5218 35545 5278
rect 35639 5218 35673 5278
rect 35767 5218 35801 5278
rect 35895 5218 35929 5278
rect 36023 5218 36057 5278
rect 36151 5218 36185 5278
rect 36279 5218 36313 5278
rect 36407 5218 36441 5278
rect 36535 5218 36569 5278
rect 36663 5218 36697 5278
rect 36791 5218 36825 5278
rect 36919 5218 36953 5278
rect 37047 5218 37081 5278
rect 37175 5218 37209 5278
rect 37303 5218 37337 5278
rect 37431 5218 37465 5278
rect 37559 5218 37593 5278
rect -319 5110 -281 5148
rect -191 5110 -153 5148
rect 609 5110 647 5148
rect 737 5110 775 5148
rect 865 5110 903 5148
rect 1873 5110 1911 5148
rect 2001 5110 2039 5148
rect 2129 5110 2167 5148
rect 2257 5110 2295 5148
rect 2385 5110 2423 5148
rect 3492 5110 3530 5148
rect 3620 5110 3658 5148
rect 3748 5110 3786 5148
rect 3876 5110 3914 5148
rect 4004 5110 4042 5148
rect 4132 5110 4170 5148
rect 4260 5110 4298 5148
rect 4388 5110 4426 5148
rect 4516 5110 4554 5148
rect 8057 5110 8095 5148
rect 8185 5110 8223 5148
rect 8313 5110 8351 5148
rect 8441 5110 8479 5148
rect 8569 5110 8607 5148
rect 8697 5110 8735 5148
rect 8825 5110 8863 5148
rect 8953 5110 8991 5148
rect 9081 5110 9119 5148
rect 9209 5110 9247 5148
rect 9337 5110 9375 5148
rect 9465 5110 9503 5148
rect 9593 5110 9631 5148
rect 9721 5110 9759 5148
rect 9849 5110 9887 5148
rect 9977 5110 10015 5148
rect 10105 5110 10143 5148
rect 15821 5110 15859 5148
rect 15949 5110 15987 5148
rect 16077 5110 16115 5148
rect 16205 5110 16243 5148
rect 16333 5110 16371 5148
rect 16461 5110 16499 5148
rect 16589 5110 16627 5148
rect 16717 5110 16755 5148
rect 16845 5110 16883 5148
rect 16973 5110 17011 5148
rect 17101 5110 17139 5148
rect 17229 5110 17267 5148
rect 17357 5110 17395 5148
rect 17485 5110 17523 5148
rect 17613 5110 17651 5148
rect 17741 5110 17779 5148
rect 17869 5110 17907 5148
rect 17997 5110 18035 5148
rect 18125 5110 18163 5148
rect 18253 5110 18291 5148
rect 18381 5110 18419 5148
rect 18509 5110 18547 5148
rect 18637 5110 18675 5148
rect 18765 5110 18803 5148
rect 18893 5110 18931 5148
rect 19021 5110 19059 5148
rect 19149 5110 19187 5148
rect 19277 5110 19315 5148
rect 19405 5110 19443 5148
rect 19533 5110 19571 5148
rect 19661 5110 19699 5148
rect 19789 5110 19827 5148
rect 19917 5110 19955 5148
rect 29365 5110 29403 5148
rect 29493 5110 29531 5148
rect 29621 5110 29659 5148
rect 29749 5110 29787 5148
rect 29877 5110 29915 5148
rect 30005 5110 30043 5148
rect 30133 5110 30171 5148
rect 30261 5110 30299 5148
rect 30389 5110 30427 5148
rect 30517 5110 30555 5148
rect 30645 5110 30683 5148
rect 30773 5110 30811 5148
rect 30901 5110 30939 5148
rect 31029 5110 31067 5148
rect 31157 5110 31195 5148
rect 31285 5110 31323 5148
rect 31413 5110 31451 5148
rect 31541 5110 31579 5148
rect 31669 5110 31707 5148
rect 31797 5110 31835 5148
rect 31925 5110 31963 5148
rect 32053 5110 32091 5148
rect 32181 5110 32219 5148
rect 32309 5110 32347 5148
rect 32437 5110 32475 5148
rect 32565 5110 32603 5148
rect 32693 5110 32731 5148
rect 32821 5110 32859 5148
rect 32949 5110 32987 5148
rect 33077 5110 33115 5148
rect 33205 5110 33243 5148
rect 33333 5110 33371 5148
rect 33461 5110 33499 5148
rect 33589 5110 33627 5148
rect 33717 5110 33755 5148
rect 33845 5110 33883 5148
rect 33973 5110 34011 5148
rect 34101 5110 34139 5148
rect 34229 5110 34267 5148
rect 34357 5110 34395 5148
rect 34485 5110 34523 5148
rect 34613 5110 34651 5148
rect 34741 5110 34779 5148
rect 34869 5110 34907 5148
rect 34997 5110 35035 5148
rect 35125 5110 35163 5148
rect 35253 5110 35291 5148
rect 35381 5110 35419 5148
rect 35509 5110 35547 5148
rect 35637 5110 35675 5148
rect 35765 5110 35803 5148
rect 35893 5110 35931 5148
rect 36021 5110 36059 5148
rect 36149 5110 36187 5148
rect 36277 5110 36315 5148
rect 36405 5110 36443 5148
rect 36533 5110 36571 5148
rect 36661 5110 36699 5148
rect 36789 5110 36827 5148
rect 36917 5110 36955 5148
rect 37045 5110 37083 5148
rect 37173 5110 37211 5148
rect 37301 5110 37339 5148
rect 37429 5110 37467 5148
rect 37557 5110 37595 5148
<< metal1 >>
rect -363 6308 38471 6314
rect -363 6270 -319 6308
rect -281 6270 -191 6308
rect -153 6270 481 6308
rect 519 6270 609 6308
rect 647 6270 737 6308
rect 775 6270 1361 6308
rect 1399 6270 1489 6308
rect 1527 6270 1617 6308
rect 1655 6270 1745 6308
rect 1783 6270 1873 6308
rect 1911 6270 2980 6308
rect 3018 6270 3108 6308
rect 3146 6270 3236 6308
rect 3274 6270 3364 6308
rect 3402 6270 3492 6308
rect 3530 6270 3620 6308
rect 3658 6270 3748 6308
rect 3786 6270 3876 6308
rect 3914 6270 4004 6308
rect 4042 6270 5473 6308
rect 5511 6270 5601 6308
rect 5639 6270 5729 6308
rect 5767 6270 5857 6308
rect 5895 6270 5985 6308
rect 6023 6270 6113 6308
rect 6151 6270 6241 6308
rect 6279 6270 6369 6308
rect 6407 6270 6497 6308
rect 6535 6270 6625 6308
rect 6663 6270 6753 6308
rect 6791 6270 6881 6308
rect 6919 6270 7009 6308
rect 7047 6270 7137 6308
rect 7175 6270 7265 6308
rect 7303 6270 7393 6308
rect 7431 6270 7521 6308
rect 7559 6270 10560 6308
rect 10598 6270 10688 6308
rect 10726 6270 10816 6308
rect 10854 6270 10944 6308
rect 10982 6270 11072 6308
rect 11110 6270 11200 6308
rect 11238 6270 11328 6308
rect 11366 6270 11456 6308
rect 11494 6270 11584 6308
rect 11622 6270 11712 6308
rect 11750 6270 11840 6308
rect 11878 6270 11968 6308
rect 12006 6270 12096 6308
rect 12134 6270 12224 6308
rect 12262 6270 12352 6308
rect 12390 6270 12480 6308
rect 12518 6270 12608 6308
rect 12646 6270 12736 6308
rect 12774 6270 12864 6308
rect 12902 6270 12992 6308
rect 13030 6270 13120 6308
rect 13158 6270 13248 6308
rect 13286 6270 13376 6308
rect 13414 6270 13504 6308
rect 13542 6270 13632 6308
rect 13670 6270 13760 6308
rect 13798 6270 13888 6308
rect 13926 6270 14016 6308
rect 14054 6270 14144 6308
rect 14182 6270 14272 6308
rect 14310 6270 14400 6308
rect 14438 6270 14528 6308
rect 14566 6270 14656 6308
rect 14694 6270 20397 6308
rect 20435 6270 20525 6308
rect 20563 6270 20653 6308
rect 20691 6270 20781 6308
rect 20819 6270 20909 6308
rect 20947 6270 21037 6308
rect 21075 6270 21165 6308
rect 21203 6270 21293 6308
rect 21331 6270 21421 6308
rect 21459 6270 21549 6308
rect 21587 6270 21677 6308
rect 21715 6270 21805 6308
rect 21843 6270 21933 6308
rect 21971 6270 22061 6308
rect 22099 6270 22189 6308
rect 22227 6270 22317 6308
rect 22355 6270 22445 6308
rect 22483 6270 22573 6308
rect 22611 6270 22701 6308
rect 22739 6270 22829 6308
rect 22867 6270 22957 6308
rect 22995 6270 23085 6308
rect 23123 6270 23213 6308
rect 23251 6270 23341 6308
rect 23379 6270 23469 6308
rect 23507 6270 23597 6308
rect 23635 6270 23725 6308
rect 23763 6270 23853 6308
rect 23891 6270 23981 6308
rect 24019 6270 24109 6308
rect 24147 6270 24237 6308
rect 24275 6270 24365 6308
rect 24403 6270 24493 6308
rect 24531 6270 24621 6308
rect 24659 6270 24749 6308
rect 24787 6270 24877 6308
rect 24915 6270 25005 6308
rect 25043 6270 25133 6308
rect 25171 6270 25261 6308
rect 25299 6270 25389 6308
rect 25427 6270 25517 6308
rect 25555 6270 25645 6308
rect 25683 6270 25773 6308
rect 25811 6270 25901 6308
rect 25939 6270 26029 6308
rect 26067 6270 26157 6308
rect 26195 6270 26285 6308
rect 26323 6270 26413 6308
rect 26451 6270 26541 6308
rect 26579 6270 26669 6308
rect 26707 6270 26797 6308
rect 26835 6270 26925 6308
rect 26963 6270 27053 6308
rect 27091 6270 27181 6308
rect 27219 6270 27309 6308
rect 27347 6270 27437 6308
rect 27475 6270 27565 6308
rect 27603 6270 27693 6308
rect 27731 6270 27821 6308
rect 27859 6270 27949 6308
rect 27987 6270 28077 6308
rect 28115 6270 28205 6308
rect 28243 6270 28333 6308
rect 28371 6270 28461 6308
rect 28499 6270 28589 6308
rect 28627 6270 38413 6308
rect -363 6264 38413 6270
rect -317 6212 -283 6264
rect 483 6212 517 6264
rect 739 6212 773 6264
rect 1363 6212 1397 6264
rect 1619 6212 1653 6264
rect 1875 6212 1909 6264
rect 2982 6212 3016 6264
rect 3238 6212 3272 6264
rect 3494 6212 3528 6264
rect 3750 6212 3784 6264
rect 4006 6212 4040 6264
rect 5475 6212 5509 6264
rect 5731 6212 5765 6264
rect 5987 6212 6021 6264
rect 6243 6212 6277 6264
rect 6499 6212 6533 6264
rect 6755 6212 6789 6264
rect 7011 6212 7045 6264
rect 7267 6212 7301 6264
rect 7523 6212 7557 6264
rect 10562 6212 10596 6264
rect 10818 6212 10852 6264
rect 11074 6212 11108 6264
rect 11330 6212 11364 6264
rect 11586 6212 11620 6264
rect 11842 6212 11876 6264
rect 12098 6212 12132 6264
rect 12354 6212 12388 6264
rect 12610 6212 12644 6264
rect 12866 6212 12900 6264
rect 13122 6212 13156 6264
rect 13378 6212 13412 6264
rect 13634 6212 13668 6264
rect 13890 6212 13924 6264
rect 14146 6212 14180 6264
rect 14402 6212 14436 6264
rect 14658 6212 14692 6264
rect 20399 6212 20433 6264
rect 20655 6212 20689 6264
rect 20911 6212 20945 6264
rect 21167 6212 21201 6264
rect 21423 6212 21457 6264
rect 21679 6212 21713 6264
rect 21935 6212 21969 6264
rect 22191 6212 22225 6264
rect 22447 6212 22481 6264
rect 22703 6212 22737 6264
rect 22959 6212 22993 6264
rect 23215 6212 23249 6264
rect 23471 6212 23505 6264
rect 23727 6212 23761 6264
rect 23983 6212 24017 6264
rect 24239 6212 24273 6264
rect 24495 6212 24529 6264
rect 24751 6212 24785 6264
rect 25007 6212 25041 6264
rect 25263 6212 25297 6264
rect 25519 6212 25553 6264
rect 25775 6212 25809 6264
rect 26031 6212 26065 6264
rect 26287 6212 26321 6264
rect 26543 6212 26577 6264
rect 26799 6212 26833 6264
rect 27055 6212 27089 6264
rect 27311 6212 27345 6264
rect 27567 6212 27601 6264
rect 27823 6212 27857 6264
rect 28079 6212 28113 6264
rect 28335 6212 28369 6264
rect 28591 6212 28625 6264
rect 38407 6256 38413 6264
rect 38465 6256 38471 6308
rect 38407 6250 38471 6256
rect -323 6200 -277 6212
rect -323 6140 -317 6200
rect -283 6140 -277 6200
rect -323 6128 -277 6140
rect -195 6200 -149 6212
rect -195 6140 -189 6200
rect -155 6140 -149 6200
rect -195 6128 -149 6140
rect 477 6200 523 6212
rect 477 6140 483 6200
rect 517 6140 523 6200
rect 477 6128 523 6140
rect 605 6200 651 6212
rect 605 6140 611 6200
rect 645 6140 651 6200
rect 605 6128 651 6140
rect 733 6200 779 6212
rect 733 6140 739 6200
rect 773 6140 779 6200
rect 733 6128 779 6140
rect 1357 6200 1403 6212
rect 1357 6140 1363 6200
rect 1397 6140 1403 6200
rect 1357 6128 1403 6140
rect 1485 6200 1531 6212
rect 1485 6140 1491 6200
rect 1525 6140 1531 6200
rect 1485 6128 1531 6140
rect 1613 6200 1659 6212
rect 1613 6140 1619 6200
rect 1653 6140 1659 6200
rect 1613 6128 1659 6140
rect 1741 6200 1787 6212
rect 1741 6140 1747 6200
rect 1781 6140 1787 6200
rect 1741 6128 1787 6140
rect 1869 6200 1915 6212
rect 1869 6140 1875 6200
rect 1909 6140 1915 6200
rect 1869 6128 1915 6140
rect 2976 6200 3022 6212
rect 2976 6140 2982 6200
rect 3016 6140 3022 6200
rect 2976 6128 3022 6140
rect 3104 6200 3150 6212
rect 3104 6140 3110 6200
rect 3144 6140 3150 6200
rect 3104 6128 3150 6140
rect 3232 6200 3278 6212
rect 3232 6140 3238 6200
rect 3272 6140 3278 6200
rect 3232 6128 3278 6140
rect 3360 6200 3406 6212
rect 3360 6140 3366 6200
rect 3400 6140 3406 6200
rect 3360 6128 3406 6140
rect 3488 6200 3534 6212
rect 3488 6140 3494 6200
rect 3528 6140 3534 6200
rect 3488 6128 3534 6140
rect 3616 6200 3662 6212
rect 3616 6140 3622 6200
rect 3656 6140 3662 6200
rect 3616 6128 3662 6140
rect 3744 6200 3790 6212
rect 3744 6140 3750 6200
rect 3784 6140 3790 6200
rect 3744 6128 3790 6140
rect 3872 6200 3918 6212
rect 3872 6140 3878 6200
rect 3912 6140 3918 6200
rect 3872 6128 3918 6140
rect 4000 6200 4046 6212
rect 4000 6140 4006 6200
rect 4040 6140 4046 6200
rect 5469 6200 5515 6212
rect 4000 6128 4046 6140
rect 4104 6167 4176 6173
rect -304 6088 -232 6094
rect -304 6031 -298 6088
rect -238 6031 -232 6088
rect -304 6026 -232 6031
rect -189 6073 -155 6128
rect -95 6083 -31 6089
rect -95 6073 -89 6083
rect -189 6040 -89 6073
rect -189 5996 -155 6040
rect -95 6031 -89 6040
rect -37 6031 -31 6083
rect -95 6025 -31 6031
rect 357 6066 421 6072
rect 357 6014 363 6066
rect 415 6060 421 6066
rect 611 6060 645 6128
rect 1268 6109 1332 6115
rect 415 6024 645 6060
rect 746 6088 818 6094
rect 746 6031 752 6088
rect 812 6031 818 6088
rect 1268 6057 1274 6109
rect 1326 6099 1332 6109
rect 1491 6099 1525 6128
rect 1747 6099 1781 6128
rect 2803 6112 2867 6118
rect 1326 6083 1781 6099
rect 1874 6094 1938 6100
rect 1874 6083 1880 6094
rect 1326 6070 1880 6083
rect 1326 6068 1553 6070
rect 1326 6057 1332 6068
rect 1268 6051 1332 6057
rect 746 6025 818 6031
rect 415 6014 421 6024
rect 357 6008 421 6014
rect 611 5996 645 6024
rect 1491 5996 1525 6068
rect 1747 6054 1880 6070
rect 1747 5996 1781 6054
rect 1874 6042 1880 6054
rect 1932 6042 1938 6094
rect 1874 6036 1938 6042
rect 1966 6077 2038 6083
rect 1966 6020 1972 6077
rect 2032 6020 2038 6077
rect 2803 6060 2809 6112
rect 2861 6099 2867 6112
rect 3110 6099 3144 6128
rect 3366 6099 3400 6128
rect 3622 6099 3656 6128
rect 3878 6099 3912 6128
rect 4104 6110 4110 6167
rect 4170 6110 4176 6167
rect 5469 6140 5475 6200
rect 5509 6140 5515 6200
rect 5469 6128 5515 6140
rect 5597 6200 5643 6212
rect 5597 6140 5603 6200
rect 5637 6140 5643 6200
rect 5597 6128 5643 6140
rect 5725 6200 5771 6212
rect 5725 6140 5731 6200
rect 5765 6140 5771 6200
rect 5725 6128 5771 6140
rect 5853 6200 5899 6212
rect 5853 6140 5859 6200
rect 5893 6140 5899 6200
rect 5853 6128 5899 6140
rect 5981 6200 6027 6212
rect 5981 6140 5987 6200
rect 6021 6140 6027 6200
rect 5981 6128 6027 6140
rect 6109 6200 6155 6212
rect 6109 6140 6115 6200
rect 6149 6140 6155 6200
rect 6109 6128 6155 6140
rect 6237 6200 6283 6212
rect 6237 6140 6243 6200
rect 6277 6140 6283 6200
rect 6237 6128 6283 6140
rect 6365 6200 6411 6212
rect 6365 6140 6371 6200
rect 6405 6140 6411 6200
rect 6365 6128 6411 6140
rect 6493 6200 6539 6212
rect 6493 6140 6499 6200
rect 6533 6140 6539 6200
rect 6493 6128 6539 6140
rect 6621 6200 6667 6212
rect 6621 6140 6627 6200
rect 6661 6140 6667 6200
rect 6621 6128 6667 6140
rect 6749 6200 6795 6212
rect 6749 6140 6755 6200
rect 6789 6140 6795 6200
rect 6749 6128 6795 6140
rect 6877 6200 6923 6212
rect 6877 6140 6883 6200
rect 6917 6140 6923 6200
rect 6877 6128 6923 6140
rect 7005 6200 7051 6212
rect 7005 6140 7011 6200
rect 7045 6140 7051 6200
rect 7005 6128 7051 6140
rect 7133 6200 7179 6212
rect 7133 6140 7139 6200
rect 7173 6140 7179 6200
rect 7133 6128 7179 6140
rect 7261 6200 7307 6212
rect 7261 6140 7267 6200
rect 7301 6140 7307 6200
rect 7261 6128 7307 6140
rect 7389 6200 7435 6212
rect 7389 6140 7395 6200
rect 7429 6140 7435 6200
rect 7389 6128 7435 6140
rect 7517 6200 7563 6212
rect 7517 6140 7523 6200
rect 7557 6140 7563 6200
rect 10556 6200 10602 6212
rect 7517 6128 7563 6140
rect 7681 6164 7753 6170
rect 4104 6104 4176 6110
rect 5353 6110 5417 6116
rect 2861 6086 3912 6099
rect 4015 6086 4079 6088
rect 2861 6082 4079 6086
rect 2861 6070 4021 6082
rect 2861 6060 2867 6070
rect 2803 6054 2867 6060
rect 1966 6014 2038 6020
rect 3110 5996 3144 6070
rect 3366 5996 3400 6070
rect 3622 5996 3656 6070
rect 3878 6051 4021 6070
rect 3878 5996 3912 6051
rect 4015 6030 4021 6051
rect 4073 6076 4079 6082
rect 5043 6076 5107 6081
rect 4073 6075 5107 6076
rect 4073 6030 5049 6075
rect 4015 6024 5049 6030
rect 5043 6023 5049 6024
rect 5101 6023 5107 6075
rect 5353 6058 5359 6110
rect 5411 6099 5417 6110
rect 5603 6099 5637 6128
rect 5859 6099 5893 6128
rect 5960 6099 6024 6100
rect 6115 6099 6149 6128
rect 6371 6099 6405 6128
rect 6627 6100 6661 6128
rect 6565 6099 6661 6100
rect 6883 6099 6917 6128
rect 7139 6099 7173 6128
rect 7395 6099 7429 6128
rect 7681 6107 7687 6164
rect 7747 6107 7753 6164
rect 10556 6140 10562 6200
rect 10596 6140 10602 6200
rect 10556 6128 10602 6140
rect 10684 6200 10730 6212
rect 10684 6140 10690 6200
rect 10724 6140 10730 6200
rect 10684 6128 10730 6140
rect 10812 6200 10858 6212
rect 10812 6140 10818 6200
rect 10852 6140 10858 6200
rect 10812 6128 10858 6140
rect 10940 6200 10986 6212
rect 10940 6140 10946 6200
rect 10980 6140 10986 6200
rect 10940 6128 10986 6140
rect 11068 6200 11114 6212
rect 11068 6140 11074 6200
rect 11108 6140 11114 6200
rect 11068 6128 11114 6140
rect 11196 6200 11242 6212
rect 11196 6140 11202 6200
rect 11236 6140 11242 6200
rect 11196 6128 11242 6140
rect 11324 6200 11370 6212
rect 11324 6140 11330 6200
rect 11364 6140 11370 6200
rect 11324 6128 11370 6140
rect 11452 6200 11498 6212
rect 11452 6140 11458 6200
rect 11492 6140 11498 6200
rect 11452 6128 11498 6140
rect 11580 6200 11626 6212
rect 11580 6140 11586 6200
rect 11620 6140 11626 6200
rect 11580 6128 11626 6140
rect 11708 6200 11754 6212
rect 11708 6140 11714 6200
rect 11748 6140 11754 6200
rect 11708 6128 11754 6140
rect 11836 6200 11882 6212
rect 11836 6140 11842 6200
rect 11876 6140 11882 6200
rect 11836 6128 11882 6140
rect 11964 6200 12010 6212
rect 11964 6140 11970 6200
rect 12004 6140 12010 6200
rect 11964 6128 12010 6140
rect 12092 6200 12138 6212
rect 12092 6140 12098 6200
rect 12132 6140 12138 6200
rect 12092 6128 12138 6140
rect 12220 6200 12266 6212
rect 12220 6140 12226 6200
rect 12260 6140 12266 6200
rect 12220 6128 12266 6140
rect 12348 6200 12394 6212
rect 12348 6140 12354 6200
rect 12388 6140 12394 6200
rect 12348 6128 12394 6140
rect 12476 6200 12522 6212
rect 12476 6140 12482 6200
rect 12516 6140 12522 6200
rect 12476 6128 12522 6140
rect 12604 6200 12650 6212
rect 12604 6140 12610 6200
rect 12644 6140 12650 6200
rect 12604 6128 12650 6140
rect 12732 6200 12778 6212
rect 12732 6140 12738 6200
rect 12772 6140 12778 6200
rect 12732 6128 12778 6140
rect 12860 6200 12906 6212
rect 12860 6140 12866 6200
rect 12900 6140 12906 6200
rect 12860 6128 12906 6140
rect 12988 6200 13034 6212
rect 12988 6140 12994 6200
rect 13028 6140 13034 6200
rect 12988 6128 13034 6140
rect 13116 6200 13162 6212
rect 13116 6140 13122 6200
rect 13156 6140 13162 6200
rect 13116 6128 13162 6140
rect 13244 6200 13290 6212
rect 13244 6140 13250 6200
rect 13284 6140 13290 6200
rect 13244 6128 13290 6140
rect 13372 6200 13418 6212
rect 13372 6140 13378 6200
rect 13412 6140 13418 6200
rect 13372 6128 13418 6140
rect 13500 6200 13546 6212
rect 13500 6140 13506 6200
rect 13540 6140 13546 6200
rect 13500 6128 13546 6140
rect 13628 6200 13674 6212
rect 13628 6140 13634 6200
rect 13668 6140 13674 6200
rect 13628 6128 13674 6140
rect 13756 6200 13802 6212
rect 13756 6140 13762 6200
rect 13796 6140 13802 6200
rect 13756 6128 13802 6140
rect 13884 6200 13930 6212
rect 13884 6140 13890 6200
rect 13924 6140 13930 6200
rect 13884 6128 13930 6140
rect 14012 6200 14058 6212
rect 14012 6140 14018 6200
rect 14052 6140 14058 6200
rect 14012 6128 14058 6140
rect 14140 6200 14186 6212
rect 14140 6140 14146 6200
rect 14180 6140 14186 6200
rect 14140 6128 14186 6140
rect 14268 6200 14314 6212
rect 14268 6140 14274 6200
rect 14308 6140 14314 6200
rect 14268 6128 14314 6140
rect 14396 6200 14442 6212
rect 14396 6140 14402 6200
rect 14436 6140 14442 6200
rect 14396 6128 14442 6140
rect 14524 6200 14570 6212
rect 14524 6140 14530 6200
rect 14564 6140 14570 6200
rect 14524 6128 14570 6140
rect 14652 6200 14698 6212
rect 14652 6140 14658 6200
rect 14692 6140 14698 6200
rect 14652 6128 14698 6140
rect 20393 6200 20439 6212
rect 20393 6140 20399 6200
rect 20433 6140 20439 6200
rect 20393 6128 20439 6140
rect 20521 6200 20567 6212
rect 20521 6140 20527 6200
rect 20561 6140 20567 6200
rect 20521 6128 20567 6140
rect 20649 6200 20695 6212
rect 20649 6140 20655 6200
rect 20689 6140 20695 6200
rect 20649 6128 20695 6140
rect 20777 6200 20823 6212
rect 20777 6140 20783 6200
rect 20817 6140 20823 6200
rect 20777 6128 20823 6140
rect 20905 6200 20951 6212
rect 20905 6140 20911 6200
rect 20945 6140 20951 6200
rect 20905 6128 20951 6140
rect 21033 6200 21079 6212
rect 21033 6140 21039 6200
rect 21073 6140 21079 6200
rect 21033 6128 21079 6140
rect 21161 6200 21207 6212
rect 21161 6140 21167 6200
rect 21201 6140 21207 6200
rect 21161 6128 21207 6140
rect 21289 6200 21335 6212
rect 21289 6140 21295 6200
rect 21329 6140 21335 6200
rect 21289 6128 21335 6140
rect 21417 6200 21463 6212
rect 21417 6140 21423 6200
rect 21457 6140 21463 6200
rect 21417 6128 21463 6140
rect 21545 6200 21591 6212
rect 21545 6140 21551 6200
rect 21585 6140 21591 6200
rect 21545 6128 21591 6140
rect 21673 6200 21719 6212
rect 21673 6140 21679 6200
rect 21713 6140 21719 6200
rect 21673 6128 21719 6140
rect 21801 6200 21847 6212
rect 21801 6140 21807 6200
rect 21841 6140 21847 6200
rect 21801 6128 21847 6140
rect 21929 6200 21975 6212
rect 21929 6140 21935 6200
rect 21969 6140 21975 6200
rect 21929 6128 21975 6140
rect 22057 6200 22103 6212
rect 22057 6140 22063 6200
rect 22097 6140 22103 6200
rect 22057 6128 22103 6140
rect 22185 6200 22231 6212
rect 22185 6140 22191 6200
rect 22225 6140 22231 6200
rect 22185 6128 22231 6140
rect 22313 6200 22359 6212
rect 22313 6140 22319 6200
rect 22353 6140 22359 6200
rect 22313 6128 22359 6140
rect 22441 6200 22487 6212
rect 22441 6140 22447 6200
rect 22481 6140 22487 6200
rect 22441 6128 22487 6140
rect 22569 6200 22615 6212
rect 22569 6140 22575 6200
rect 22609 6140 22615 6200
rect 22569 6128 22615 6140
rect 22697 6200 22743 6212
rect 22697 6140 22703 6200
rect 22737 6140 22743 6200
rect 22697 6128 22743 6140
rect 22825 6200 22871 6212
rect 22825 6140 22831 6200
rect 22865 6140 22871 6200
rect 22825 6128 22871 6140
rect 22953 6200 22999 6212
rect 22953 6140 22959 6200
rect 22993 6140 22999 6200
rect 22953 6128 22999 6140
rect 23081 6200 23127 6212
rect 23081 6140 23087 6200
rect 23121 6140 23127 6200
rect 23081 6128 23127 6140
rect 23209 6200 23255 6212
rect 23209 6140 23215 6200
rect 23249 6140 23255 6200
rect 23209 6128 23255 6140
rect 23337 6200 23383 6212
rect 23337 6140 23343 6200
rect 23377 6140 23383 6200
rect 23337 6128 23383 6140
rect 23465 6200 23511 6212
rect 23465 6140 23471 6200
rect 23505 6140 23511 6200
rect 23465 6128 23511 6140
rect 23593 6200 23639 6212
rect 23593 6140 23599 6200
rect 23633 6140 23639 6200
rect 23593 6128 23639 6140
rect 23721 6200 23767 6212
rect 23721 6140 23727 6200
rect 23761 6140 23767 6200
rect 23721 6128 23767 6140
rect 23849 6200 23895 6212
rect 23849 6140 23855 6200
rect 23889 6140 23895 6200
rect 23849 6128 23895 6140
rect 23977 6200 24023 6212
rect 23977 6140 23983 6200
rect 24017 6140 24023 6200
rect 23977 6128 24023 6140
rect 24105 6200 24151 6212
rect 24105 6140 24111 6200
rect 24145 6140 24151 6200
rect 24105 6128 24151 6140
rect 24233 6200 24279 6212
rect 24233 6140 24239 6200
rect 24273 6140 24279 6200
rect 24233 6128 24279 6140
rect 24361 6200 24407 6212
rect 24361 6140 24367 6200
rect 24401 6140 24407 6200
rect 24361 6128 24407 6140
rect 24489 6200 24535 6212
rect 24489 6140 24495 6200
rect 24529 6140 24535 6200
rect 24489 6128 24535 6140
rect 24617 6200 24663 6212
rect 24617 6140 24623 6200
rect 24657 6140 24663 6200
rect 24617 6128 24663 6140
rect 24745 6200 24791 6212
rect 24745 6140 24751 6200
rect 24785 6140 24791 6200
rect 24745 6128 24791 6140
rect 24873 6200 24919 6212
rect 24873 6140 24879 6200
rect 24913 6140 24919 6200
rect 24873 6128 24919 6140
rect 25001 6200 25047 6212
rect 25001 6140 25007 6200
rect 25041 6140 25047 6200
rect 25001 6128 25047 6140
rect 25129 6200 25175 6212
rect 25129 6140 25135 6200
rect 25169 6140 25175 6200
rect 25129 6128 25175 6140
rect 25257 6200 25303 6212
rect 25257 6140 25263 6200
rect 25297 6140 25303 6200
rect 25257 6128 25303 6140
rect 25385 6200 25431 6212
rect 25385 6140 25391 6200
rect 25425 6140 25431 6200
rect 25385 6128 25431 6140
rect 25513 6200 25559 6212
rect 25513 6140 25519 6200
rect 25553 6140 25559 6200
rect 25513 6128 25559 6140
rect 25641 6200 25687 6212
rect 25641 6140 25647 6200
rect 25681 6140 25687 6200
rect 25641 6128 25687 6140
rect 25769 6200 25815 6212
rect 25769 6140 25775 6200
rect 25809 6140 25815 6200
rect 25769 6128 25815 6140
rect 25897 6200 25943 6212
rect 25897 6140 25903 6200
rect 25937 6140 25943 6200
rect 25897 6128 25943 6140
rect 26025 6200 26071 6212
rect 26025 6140 26031 6200
rect 26065 6140 26071 6200
rect 26025 6128 26071 6140
rect 26153 6200 26199 6212
rect 26153 6140 26159 6200
rect 26193 6140 26199 6200
rect 26153 6128 26199 6140
rect 26281 6200 26327 6212
rect 26281 6140 26287 6200
rect 26321 6140 26327 6200
rect 26281 6128 26327 6140
rect 26409 6200 26455 6212
rect 26409 6140 26415 6200
rect 26449 6140 26455 6200
rect 26409 6128 26455 6140
rect 26537 6200 26583 6212
rect 26537 6140 26543 6200
rect 26577 6140 26583 6200
rect 26537 6128 26583 6140
rect 26665 6200 26711 6212
rect 26665 6140 26671 6200
rect 26705 6140 26711 6200
rect 26665 6128 26711 6140
rect 26793 6200 26839 6212
rect 26793 6140 26799 6200
rect 26833 6140 26839 6200
rect 26793 6128 26839 6140
rect 26921 6200 26967 6212
rect 26921 6140 26927 6200
rect 26961 6140 26967 6200
rect 26921 6128 26967 6140
rect 27049 6200 27095 6212
rect 27049 6140 27055 6200
rect 27089 6140 27095 6200
rect 27049 6128 27095 6140
rect 27177 6200 27223 6212
rect 27177 6140 27183 6200
rect 27217 6140 27223 6200
rect 27177 6128 27223 6140
rect 27305 6200 27351 6212
rect 27305 6140 27311 6200
rect 27345 6140 27351 6200
rect 27305 6128 27351 6140
rect 27433 6200 27479 6212
rect 27433 6140 27439 6200
rect 27473 6140 27479 6200
rect 27433 6128 27479 6140
rect 27561 6200 27607 6212
rect 27561 6140 27567 6200
rect 27601 6140 27607 6200
rect 27561 6128 27607 6140
rect 27689 6200 27735 6212
rect 27689 6140 27695 6200
rect 27729 6140 27735 6200
rect 27689 6128 27735 6140
rect 27817 6200 27863 6212
rect 27817 6140 27823 6200
rect 27857 6140 27863 6200
rect 27817 6128 27863 6140
rect 27945 6200 27991 6212
rect 27945 6140 27951 6200
rect 27985 6140 27991 6200
rect 27945 6128 27991 6140
rect 28073 6200 28119 6212
rect 28073 6140 28079 6200
rect 28113 6140 28119 6200
rect 28073 6128 28119 6140
rect 28201 6200 28247 6212
rect 28201 6140 28207 6200
rect 28241 6140 28247 6200
rect 28201 6128 28247 6140
rect 28329 6200 28375 6212
rect 28329 6140 28335 6200
rect 28369 6140 28375 6200
rect 28329 6128 28375 6140
rect 28457 6200 28503 6212
rect 28457 6140 28463 6200
rect 28497 6140 28503 6200
rect 28457 6128 28503 6140
rect 28585 6200 28631 6212
rect 28585 6140 28591 6200
rect 28625 6140 28631 6200
rect 28585 6128 28631 6140
rect 7681 6101 7753 6107
rect 10326 6107 10390 6113
rect 5411 6094 7429 6099
rect 5411 6070 5966 6094
rect 5411 6061 5637 6070
rect 5411 6058 5417 6061
rect 5353 6052 5417 6058
rect 5043 6017 5107 6023
rect 5603 5996 5637 6061
rect 5859 5996 5893 6070
rect 5960 6042 5966 6070
rect 6018 6070 6571 6094
rect 6018 6042 6024 6070
rect 5960 6036 6024 6042
rect 6115 5996 6149 6070
rect 6371 5996 6405 6070
rect 6565 6042 6571 6070
rect 6623 6093 7429 6094
rect 6623 6070 7177 6093
rect 6623 6042 6661 6070
rect 6565 6036 6661 6042
rect 6627 5996 6661 6036
rect 6883 5996 6917 6070
rect 7139 6041 7177 6070
rect 7229 6073 7429 6093
rect 7777 6073 7841 6076
rect 7229 6070 7841 6073
rect 7229 6041 7235 6070
rect 7139 6035 7235 6041
rect 7139 5996 7173 6035
rect 7395 6026 7783 6070
rect 7395 5996 7429 6026
rect 7777 6018 7783 6026
rect 7835 6018 7841 6070
rect 10326 6055 10332 6107
rect 10384 6097 10390 6107
rect 10690 6099 10724 6128
rect 10946 6100 10980 6128
rect 10932 6099 10996 6100
rect 11202 6099 11236 6128
rect 11458 6099 11492 6128
rect 11714 6099 11748 6128
rect 11970 6099 12004 6128
rect 12226 6099 12260 6128
rect 12482 6099 12516 6128
rect 12738 6099 12772 6128
rect 12994 6099 13028 6128
rect 13250 6099 13284 6128
rect 13506 6099 13540 6128
rect 13762 6099 13796 6128
rect 14018 6099 14052 6128
rect 14274 6099 14308 6128
rect 14530 6099 14564 6128
rect 10690 6097 14628 6099
rect 20149 6098 20213 6103
rect 20527 6099 20561 6128
rect 20783 6099 20817 6128
rect 21039 6099 21073 6128
rect 21295 6099 21329 6128
rect 21551 6099 21585 6128
rect 21807 6099 21841 6128
rect 22063 6099 22097 6128
rect 22319 6099 22353 6128
rect 22575 6099 22609 6128
rect 22831 6099 22865 6128
rect 23087 6099 23121 6128
rect 23180 6099 23244 6100
rect 23343 6099 23377 6128
rect 23599 6099 23633 6128
rect 23855 6099 23889 6128
rect 24111 6099 24145 6128
rect 24367 6099 24401 6128
rect 24623 6099 24657 6128
rect 24879 6099 24913 6128
rect 25135 6099 25169 6128
rect 25391 6099 25425 6128
rect 25647 6099 25681 6128
rect 25903 6099 25937 6128
rect 26159 6099 26193 6128
rect 26415 6099 26449 6128
rect 26671 6099 26705 6128
rect 26927 6099 26961 6128
rect 27183 6099 27217 6128
rect 27439 6099 27473 6128
rect 27695 6099 27729 6128
rect 27951 6099 27985 6128
rect 28028 6099 28092 6100
rect 28207 6099 28241 6128
rect 28463 6099 28497 6128
rect 28724 6115 28796 6121
rect 20527 6098 28696 6099
rect 10384 6094 14628 6097
rect 10384 6070 10938 6094
rect 10384 6067 10724 6070
rect 10384 6055 10390 6067
rect 10326 6049 10390 6055
rect 7777 6012 7841 6018
rect 10690 5996 10724 6067
rect 10932 6042 10938 6070
rect 10990 6093 14628 6094
rect 10990 6070 11544 6093
rect 10990 6042 10996 6070
rect 10932 6036 10996 6042
rect 10946 5996 10980 6036
rect 11202 5996 11236 6070
rect 11458 5996 11492 6070
rect 11538 6041 11544 6070
rect 11596 6070 12178 6093
rect 11596 6041 11602 6070
rect 11538 6035 11602 6041
rect 11714 5996 11748 6070
rect 11970 5996 12004 6070
rect 12172 6041 12178 6070
rect 12230 6070 12756 6093
rect 12230 6041 12260 6070
rect 12172 6035 12260 6041
rect 12226 5996 12260 6035
rect 12482 5996 12516 6070
rect 12738 6041 12756 6070
rect 12808 6087 14570 6093
rect 12808 6070 13362 6087
rect 12808 6041 12814 6070
rect 12738 6035 12814 6041
rect 12738 5996 12772 6035
rect 12994 5996 13028 6070
rect 13250 5996 13284 6070
rect 13356 6035 13362 6070
rect 13414 6070 13968 6087
rect 13414 6035 13420 6070
rect 13356 6029 13420 6035
rect 13506 5996 13540 6070
rect 13762 5996 13796 6070
rect 13962 6035 13968 6070
rect 14020 6070 14570 6087
rect 14020 6035 14052 6070
rect 13962 6029 14052 6035
rect 14018 5996 14052 6029
rect 14274 5996 14308 6070
rect 14530 6041 14570 6070
rect 14622 6041 14628 6093
rect 14530 6035 14628 6041
rect 14696 6092 14768 6098
rect 14696 6035 14702 6092
rect 14762 6035 14768 6092
rect 20149 6097 28696 6098
rect 20149 6045 20155 6097
rect 20207 6094 28696 6097
rect 20207 6093 23186 6094
rect 20207 6092 21974 6093
rect 20207 6070 20762 6092
rect 20207 6045 20213 6070
rect 20149 6039 20213 6045
rect 14530 5996 14564 6035
rect 14696 6029 14768 6035
rect 20527 5996 20561 6070
rect 20755 6052 20762 6070
rect 20756 6040 20762 6052
rect 20814 6070 21367 6092
rect 20814 6040 20820 6070
rect 20756 6034 20820 6040
rect 20783 5996 20817 6034
rect 21039 5996 21073 6070
rect 21295 5996 21329 6070
rect 21360 6052 21367 6070
rect 21361 6040 21367 6052
rect 21419 6070 21974 6092
rect 21419 6040 21425 6070
rect 21361 6034 21425 6040
rect 21551 5996 21585 6070
rect 21807 5996 21841 6070
rect 21967 6053 21974 6070
rect 21968 6041 21974 6053
rect 22026 6070 22580 6093
rect 22026 6041 22032 6070
rect 21968 6035 22032 6041
rect 22063 5996 22097 6070
rect 22319 5996 22353 6070
rect 22573 6053 22580 6070
rect 22574 6041 22580 6053
rect 22632 6070 23186 6093
rect 22632 6041 22638 6070
rect 22574 6035 22638 6041
rect 22575 5996 22609 6035
rect 22831 5996 22865 6070
rect 23087 5996 23121 6070
rect 23179 6054 23186 6070
rect 23180 6042 23186 6054
rect 23238 6093 28034 6094
rect 23238 6070 23798 6093
rect 23238 6042 23244 6070
rect 23180 6036 23244 6042
rect 23343 5996 23377 6070
rect 23599 5996 23633 6070
rect 23791 6053 23798 6070
rect 23792 6041 23798 6053
rect 23850 6070 25003 6093
rect 23850 6041 23889 6070
rect 23792 6035 23889 6041
rect 23855 5996 23889 6035
rect 24111 5996 24145 6070
rect 24367 5996 24401 6070
rect 24623 5996 24657 6070
rect 24879 5996 24913 6070
rect 24997 6041 25003 6070
rect 25055 6070 25609 6093
rect 25055 6041 25061 6070
rect 24997 6035 25061 6041
rect 25135 5996 25169 6070
rect 25391 5996 25425 6070
rect 25603 6041 25609 6070
rect 25661 6092 26822 6093
rect 25661 6070 26197 6092
rect 25661 6041 25681 6070
rect 25603 6035 25681 6041
rect 25647 5996 25681 6035
rect 25903 5996 25937 6070
rect 26159 6040 26197 6070
rect 26249 6070 26822 6092
rect 26249 6040 26255 6070
rect 26159 6034 26255 6040
rect 26159 5996 26193 6034
rect 26415 5996 26449 6070
rect 26671 5996 26705 6070
rect 26816 6041 26822 6070
rect 26874 6070 27429 6093
rect 26874 6041 26880 6070
rect 26816 6035 26880 6041
rect 26927 5996 26961 6070
rect 27183 5996 27217 6070
rect 27423 6041 27429 6070
rect 27481 6070 28034 6093
rect 27481 6041 27487 6070
rect 27423 6035 27487 6041
rect 27439 5996 27473 6035
rect 27695 5996 27729 6070
rect 27951 5996 27985 6070
rect 28028 6042 28034 6070
rect 28086 6093 28696 6094
rect 28086 6070 28638 6093
rect 28086 6042 28092 6070
rect 28028 6036 28092 6042
rect 28207 5996 28241 6070
rect 28463 5996 28497 6070
rect 28632 6041 28638 6070
rect 28690 6041 28696 6093
rect 28724 6058 28730 6115
rect 28790 6058 28796 6115
rect 28724 6052 28796 6058
rect 28632 6035 28696 6041
rect -323 5984 -277 5996
rect -323 5840 -317 5984
rect -283 5840 -277 5984
rect -323 5828 -277 5840
rect -195 5984 -149 5996
rect -195 5840 -189 5984
rect -155 5840 -149 5984
rect -195 5828 -149 5840
rect 477 5984 523 5996
rect 477 5840 483 5984
rect 517 5840 523 5984
rect 477 5828 523 5840
rect 605 5984 651 5996
rect 605 5840 611 5984
rect 645 5840 651 5984
rect 605 5828 651 5840
rect 733 5984 779 5996
rect 733 5840 739 5984
rect 773 5840 779 5984
rect 733 5828 779 5840
rect 1357 5984 1403 5996
rect 1357 5840 1363 5984
rect 1397 5840 1403 5984
rect 1357 5828 1403 5840
rect 1485 5984 1531 5996
rect 1485 5840 1491 5984
rect 1525 5840 1531 5984
rect 1485 5828 1531 5840
rect 1613 5984 1659 5996
rect 1613 5840 1619 5984
rect 1653 5840 1659 5984
rect 1613 5828 1659 5840
rect 1741 5984 1787 5996
rect 1741 5840 1747 5984
rect 1781 5840 1787 5984
rect 1741 5828 1787 5840
rect 1869 5984 1915 5996
rect 1869 5840 1875 5984
rect 1909 5840 1915 5984
rect 1869 5828 1915 5840
rect 2976 5984 3022 5996
rect 2976 5840 2982 5984
rect 3016 5840 3022 5984
rect 2976 5828 3022 5840
rect 3104 5984 3150 5996
rect 3104 5840 3110 5984
rect 3144 5840 3150 5984
rect 3104 5828 3150 5840
rect 3232 5984 3278 5996
rect 3232 5840 3238 5984
rect 3272 5840 3278 5984
rect 3232 5828 3278 5840
rect 3360 5984 3406 5996
rect 3360 5840 3366 5984
rect 3400 5840 3406 5984
rect 3360 5828 3406 5840
rect 3488 5984 3534 5996
rect 3488 5840 3494 5984
rect 3528 5840 3534 5984
rect 3488 5828 3534 5840
rect 3616 5984 3662 5996
rect 3616 5840 3622 5984
rect 3656 5840 3662 5984
rect 3616 5828 3662 5840
rect 3744 5984 3790 5996
rect 3744 5840 3750 5984
rect 3784 5840 3790 5984
rect 3744 5828 3790 5840
rect 3872 5984 3918 5996
rect 3872 5840 3878 5984
rect 3912 5840 3918 5984
rect 3872 5828 3918 5840
rect 4000 5984 4046 5996
rect 4000 5840 4006 5984
rect 4040 5840 4046 5984
rect 4000 5828 4046 5840
rect 5469 5984 5515 5996
rect 5469 5840 5475 5984
rect 5509 5840 5515 5984
rect 5469 5828 5515 5840
rect 5597 5984 5643 5996
rect 5597 5840 5603 5984
rect 5637 5840 5643 5984
rect 5597 5828 5643 5840
rect 5725 5984 5771 5996
rect 5725 5840 5731 5984
rect 5765 5840 5771 5984
rect 5725 5828 5771 5840
rect 5853 5984 5899 5996
rect 5853 5840 5859 5984
rect 5893 5840 5899 5984
rect 5853 5828 5899 5840
rect 5981 5984 6027 5996
rect 5981 5840 5987 5984
rect 6021 5840 6027 5984
rect 5981 5828 6027 5840
rect 6109 5984 6155 5996
rect 6109 5840 6115 5984
rect 6149 5840 6155 5984
rect 6109 5828 6155 5840
rect 6237 5984 6283 5996
rect 6237 5840 6243 5984
rect 6277 5840 6283 5984
rect 6237 5828 6283 5840
rect 6365 5984 6411 5996
rect 6365 5840 6371 5984
rect 6405 5840 6411 5984
rect 6365 5828 6411 5840
rect 6493 5984 6539 5996
rect 6493 5840 6499 5984
rect 6533 5840 6539 5984
rect 6493 5828 6539 5840
rect 6621 5984 6667 5996
rect 6621 5840 6627 5984
rect 6661 5840 6667 5984
rect 6621 5828 6667 5840
rect 6749 5984 6795 5996
rect 6749 5840 6755 5984
rect 6789 5840 6795 5984
rect 6749 5828 6795 5840
rect 6877 5984 6923 5996
rect 6877 5840 6883 5984
rect 6917 5840 6923 5984
rect 6877 5828 6923 5840
rect 7005 5984 7051 5996
rect 7005 5840 7011 5984
rect 7045 5840 7051 5984
rect 7005 5828 7051 5840
rect 7133 5984 7179 5996
rect 7133 5840 7139 5984
rect 7173 5840 7179 5984
rect 7133 5828 7179 5840
rect 7261 5984 7307 5996
rect 7261 5840 7267 5984
rect 7301 5840 7307 5984
rect 7261 5828 7307 5840
rect 7389 5984 7435 5996
rect 7389 5840 7395 5984
rect 7429 5840 7435 5984
rect 7389 5828 7435 5840
rect 7517 5984 7563 5996
rect 7517 5840 7523 5984
rect 7557 5840 7563 5984
rect 7517 5828 7563 5840
rect 10556 5984 10602 5996
rect 10556 5840 10562 5984
rect 10596 5840 10602 5984
rect 10556 5828 10602 5840
rect 10684 5984 10730 5996
rect 10684 5840 10690 5984
rect 10724 5840 10730 5984
rect 10684 5828 10730 5840
rect 10812 5984 10858 5996
rect 10812 5840 10818 5984
rect 10852 5840 10858 5984
rect 10812 5828 10858 5840
rect 10940 5984 10986 5996
rect 10940 5840 10946 5984
rect 10980 5840 10986 5984
rect 10940 5828 10986 5840
rect 11068 5984 11114 5996
rect 11068 5840 11074 5984
rect 11108 5840 11114 5984
rect 11068 5828 11114 5840
rect 11196 5984 11242 5996
rect 11196 5840 11202 5984
rect 11236 5840 11242 5984
rect 11196 5828 11242 5840
rect 11324 5984 11370 5996
rect 11324 5840 11330 5984
rect 11364 5840 11370 5984
rect 11324 5828 11370 5840
rect 11452 5984 11498 5996
rect 11452 5840 11458 5984
rect 11492 5840 11498 5984
rect 11452 5828 11498 5840
rect 11580 5984 11626 5996
rect 11580 5840 11586 5984
rect 11620 5840 11626 5984
rect 11580 5828 11626 5840
rect 11708 5984 11754 5996
rect 11708 5840 11714 5984
rect 11748 5840 11754 5984
rect 11708 5828 11754 5840
rect 11836 5984 11882 5996
rect 11836 5840 11842 5984
rect 11876 5840 11882 5984
rect 11836 5828 11882 5840
rect 11964 5984 12010 5996
rect 11964 5840 11970 5984
rect 12004 5840 12010 5984
rect 11964 5828 12010 5840
rect 12092 5984 12138 5996
rect 12092 5840 12098 5984
rect 12132 5840 12138 5984
rect 12092 5828 12138 5840
rect 12220 5984 12266 5996
rect 12220 5840 12226 5984
rect 12260 5840 12266 5984
rect 12220 5828 12266 5840
rect 12348 5984 12394 5996
rect 12348 5840 12354 5984
rect 12388 5840 12394 5984
rect 12348 5828 12394 5840
rect 12476 5984 12522 5996
rect 12476 5840 12482 5984
rect 12516 5840 12522 5984
rect 12476 5828 12522 5840
rect 12604 5984 12650 5996
rect 12604 5840 12610 5984
rect 12644 5840 12650 5984
rect 12604 5828 12650 5840
rect 12732 5984 12778 5996
rect 12732 5840 12738 5984
rect 12772 5840 12778 5984
rect 12732 5828 12778 5840
rect 12860 5984 12906 5996
rect 12860 5840 12866 5984
rect 12900 5840 12906 5984
rect 12860 5828 12906 5840
rect 12988 5984 13034 5996
rect 12988 5840 12994 5984
rect 13028 5840 13034 5984
rect 12988 5828 13034 5840
rect 13116 5984 13162 5996
rect 13116 5840 13122 5984
rect 13156 5840 13162 5984
rect 13116 5828 13162 5840
rect 13244 5984 13290 5996
rect 13244 5840 13250 5984
rect 13284 5840 13290 5984
rect 13244 5828 13290 5840
rect 13372 5984 13418 5996
rect 13372 5840 13378 5984
rect 13412 5840 13418 5984
rect 13372 5828 13418 5840
rect 13500 5984 13546 5996
rect 13500 5840 13506 5984
rect 13540 5840 13546 5984
rect 13500 5828 13546 5840
rect 13628 5984 13674 5996
rect 13628 5840 13634 5984
rect 13668 5840 13674 5984
rect 13628 5828 13674 5840
rect 13756 5984 13802 5996
rect 13756 5840 13762 5984
rect 13796 5840 13802 5984
rect 13756 5828 13802 5840
rect 13884 5984 13930 5996
rect 13884 5840 13890 5984
rect 13924 5840 13930 5984
rect 13884 5828 13930 5840
rect 14012 5984 14058 5996
rect 14012 5840 14018 5984
rect 14052 5840 14058 5984
rect 14012 5828 14058 5840
rect 14140 5984 14186 5996
rect 14140 5840 14146 5984
rect 14180 5840 14186 5984
rect 14140 5828 14186 5840
rect 14268 5984 14314 5996
rect 14268 5840 14274 5984
rect 14308 5840 14314 5984
rect 14268 5828 14314 5840
rect 14396 5984 14442 5996
rect 14396 5840 14402 5984
rect 14436 5840 14442 5984
rect 14396 5828 14442 5840
rect 14524 5984 14570 5996
rect 14524 5840 14530 5984
rect 14564 5840 14570 5984
rect 14524 5828 14570 5840
rect 14652 5984 14698 5996
rect 14652 5840 14658 5984
rect 14692 5840 14698 5984
rect 14652 5828 14698 5840
rect 20393 5984 20439 5996
rect 20393 5840 20399 5984
rect 20433 5840 20439 5984
rect 20393 5828 20439 5840
rect 20521 5984 20567 5996
rect 20521 5840 20527 5984
rect 20561 5840 20567 5984
rect 20521 5828 20567 5840
rect 20649 5984 20695 5996
rect 20649 5840 20655 5984
rect 20689 5840 20695 5984
rect 20649 5828 20695 5840
rect 20777 5984 20823 5996
rect 20777 5840 20783 5984
rect 20817 5840 20823 5984
rect 20777 5828 20823 5840
rect 20905 5984 20951 5996
rect 20905 5840 20911 5984
rect 20945 5840 20951 5984
rect 20905 5828 20951 5840
rect 21033 5984 21079 5996
rect 21033 5840 21039 5984
rect 21073 5840 21079 5984
rect 21033 5828 21079 5840
rect 21161 5984 21207 5996
rect 21161 5840 21167 5984
rect 21201 5840 21207 5984
rect 21161 5828 21207 5840
rect 21289 5984 21335 5996
rect 21289 5840 21295 5984
rect 21329 5840 21335 5984
rect 21289 5828 21335 5840
rect 21417 5984 21463 5996
rect 21417 5840 21423 5984
rect 21457 5840 21463 5984
rect 21417 5828 21463 5840
rect 21545 5984 21591 5996
rect 21545 5840 21551 5984
rect 21585 5840 21591 5984
rect 21545 5828 21591 5840
rect 21673 5984 21719 5996
rect 21673 5840 21679 5984
rect 21713 5840 21719 5984
rect 21673 5828 21719 5840
rect 21801 5984 21847 5996
rect 21801 5840 21807 5984
rect 21841 5840 21847 5984
rect 21801 5828 21847 5840
rect 21929 5984 21975 5996
rect 21929 5840 21935 5984
rect 21969 5840 21975 5984
rect 21929 5828 21975 5840
rect 22057 5984 22103 5996
rect 22057 5840 22063 5984
rect 22097 5840 22103 5984
rect 22057 5828 22103 5840
rect 22185 5984 22231 5996
rect 22185 5840 22191 5984
rect 22225 5840 22231 5984
rect 22185 5828 22231 5840
rect 22313 5984 22359 5996
rect 22313 5840 22319 5984
rect 22353 5840 22359 5984
rect 22313 5828 22359 5840
rect 22441 5984 22487 5996
rect 22441 5840 22447 5984
rect 22481 5840 22487 5984
rect 22441 5828 22487 5840
rect 22569 5984 22615 5996
rect 22569 5840 22575 5984
rect 22609 5840 22615 5984
rect 22569 5828 22615 5840
rect 22697 5984 22743 5996
rect 22697 5840 22703 5984
rect 22737 5840 22743 5984
rect 22697 5828 22743 5840
rect 22825 5984 22871 5996
rect 22825 5840 22831 5984
rect 22865 5840 22871 5984
rect 22825 5828 22871 5840
rect 22953 5984 22999 5996
rect 22953 5840 22959 5984
rect 22993 5840 22999 5984
rect 22953 5828 22999 5840
rect 23081 5984 23127 5996
rect 23081 5840 23087 5984
rect 23121 5840 23127 5984
rect 23081 5828 23127 5840
rect 23209 5984 23255 5996
rect 23209 5840 23215 5984
rect 23249 5840 23255 5984
rect 23209 5828 23255 5840
rect 23337 5984 23383 5996
rect 23337 5840 23343 5984
rect 23377 5840 23383 5984
rect 23337 5828 23383 5840
rect 23465 5984 23511 5996
rect 23465 5840 23471 5984
rect 23505 5840 23511 5984
rect 23465 5828 23511 5840
rect 23593 5984 23639 5996
rect 23593 5840 23599 5984
rect 23633 5840 23639 5984
rect 23593 5828 23639 5840
rect 23721 5984 23767 5996
rect 23721 5840 23727 5984
rect 23761 5840 23767 5984
rect 23721 5828 23767 5840
rect 23849 5984 23895 5996
rect 23849 5840 23855 5984
rect 23889 5840 23895 5984
rect 23849 5828 23895 5840
rect 23977 5984 24023 5996
rect 23977 5840 23983 5984
rect 24017 5840 24023 5984
rect 23977 5828 24023 5840
rect 24105 5984 24151 5996
rect 24105 5840 24111 5984
rect 24145 5840 24151 5984
rect 24105 5828 24151 5840
rect 24233 5984 24279 5996
rect 24233 5840 24239 5984
rect 24273 5840 24279 5984
rect 24233 5828 24279 5840
rect 24361 5984 24407 5996
rect 24361 5840 24367 5984
rect 24401 5840 24407 5984
rect 24361 5828 24407 5840
rect 24489 5984 24535 5996
rect 24489 5840 24495 5984
rect 24529 5840 24535 5984
rect 24489 5828 24535 5840
rect 24617 5984 24663 5996
rect 24617 5840 24623 5984
rect 24657 5840 24663 5984
rect 24617 5828 24663 5840
rect 24745 5984 24791 5996
rect 24745 5840 24751 5984
rect 24785 5840 24791 5984
rect 24745 5828 24791 5840
rect 24873 5984 24919 5996
rect 24873 5840 24879 5984
rect 24913 5840 24919 5984
rect 24873 5828 24919 5840
rect 25001 5984 25047 5996
rect 25001 5840 25007 5984
rect 25041 5840 25047 5984
rect 25001 5828 25047 5840
rect 25129 5984 25175 5996
rect 25129 5840 25135 5984
rect 25169 5840 25175 5984
rect 25129 5828 25175 5840
rect 25257 5984 25303 5996
rect 25257 5840 25263 5984
rect 25297 5840 25303 5984
rect 25257 5828 25303 5840
rect 25385 5984 25431 5996
rect 25385 5840 25391 5984
rect 25425 5840 25431 5984
rect 25385 5828 25431 5840
rect 25513 5984 25559 5996
rect 25513 5840 25519 5984
rect 25553 5840 25559 5984
rect 25513 5828 25559 5840
rect 25641 5984 25687 5996
rect 25641 5840 25647 5984
rect 25681 5840 25687 5984
rect 25641 5828 25687 5840
rect 25769 5984 25815 5996
rect 25769 5840 25775 5984
rect 25809 5840 25815 5984
rect 25769 5828 25815 5840
rect 25897 5984 25943 5996
rect 25897 5840 25903 5984
rect 25937 5840 25943 5984
rect 25897 5828 25943 5840
rect 26025 5984 26071 5996
rect 26025 5840 26031 5984
rect 26065 5840 26071 5984
rect 26025 5828 26071 5840
rect 26153 5984 26199 5996
rect 26153 5840 26159 5984
rect 26193 5840 26199 5984
rect 26153 5828 26199 5840
rect 26281 5984 26327 5996
rect 26281 5840 26287 5984
rect 26321 5840 26327 5984
rect 26281 5828 26327 5840
rect 26409 5984 26455 5996
rect 26409 5840 26415 5984
rect 26449 5840 26455 5984
rect 26409 5828 26455 5840
rect 26537 5984 26583 5996
rect 26537 5840 26543 5984
rect 26577 5840 26583 5984
rect 26537 5828 26583 5840
rect 26665 5984 26711 5996
rect 26665 5840 26671 5984
rect 26705 5840 26711 5984
rect 26665 5828 26711 5840
rect 26793 5984 26839 5996
rect 26793 5840 26799 5984
rect 26833 5840 26839 5984
rect 26793 5828 26839 5840
rect 26921 5984 26967 5996
rect 26921 5840 26927 5984
rect 26961 5840 26967 5984
rect 26921 5828 26967 5840
rect 27049 5984 27095 5996
rect 27049 5840 27055 5984
rect 27089 5840 27095 5984
rect 27049 5828 27095 5840
rect 27177 5984 27223 5996
rect 27177 5840 27183 5984
rect 27217 5840 27223 5984
rect 27177 5828 27223 5840
rect 27305 5984 27351 5996
rect 27305 5840 27311 5984
rect 27345 5840 27351 5984
rect 27305 5828 27351 5840
rect 27433 5984 27479 5996
rect 27433 5840 27439 5984
rect 27473 5840 27479 5984
rect 27433 5828 27479 5840
rect 27561 5984 27607 5996
rect 27561 5840 27567 5984
rect 27601 5840 27607 5984
rect 27561 5828 27607 5840
rect 27689 5984 27735 5996
rect 27689 5840 27695 5984
rect 27729 5840 27735 5984
rect 27689 5828 27735 5840
rect 27817 5984 27863 5996
rect 27817 5840 27823 5984
rect 27857 5840 27863 5984
rect 27817 5828 27863 5840
rect 27945 5984 27991 5996
rect 27945 5840 27951 5984
rect 27985 5840 27991 5984
rect 27945 5828 27991 5840
rect 28073 5984 28119 5996
rect 28073 5840 28079 5984
rect 28113 5840 28119 5984
rect 28073 5828 28119 5840
rect 28201 5984 28247 5996
rect 28201 5840 28207 5984
rect 28241 5840 28247 5984
rect 28201 5828 28247 5840
rect 28329 5984 28375 5996
rect 28329 5840 28335 5984
rect 28369 5840 28375 5984
rect 28329 5828 28375 5840
rect 28457 5984 28503 5996
rect 28457 5840 28463 5984
rect 28497 5840 28503 5984
rect 28457 5828 28503 5840
rect 28585 5984 28631 5996
rect 28585 5840 28591 5984
rect 28625 5840 28631 5984
rect 28585 5828 28631 5840
rect -317 5795 -283 5828
rect 483 5795 517 5828
rect 739 5795 773 5828
rect 1363 5795 1397 5828
rect 1619 5795 1653 5828
rect 1875 5795 1909 5828
rect 2982 5795 3016 5828
rect 3238 5795 3272 5828
rect 3494 5795 3528 5828
rect 3750 5795 3784 5828
rect 4006 5795 4040 5828
rect 5475 5795 5509 5828
rect 5731 5795 5765 5828
rect 5987 5795 6021 5828
rect 6243 5795 6277 5828
rect 6499 5795 6533 5828
rect 6755 5795 6789 5828
rect 7011 5795 7045 5828
rect 7267 5795 7301 5828
rect 7523 5795 7557 5828
rect 10562 5795 10596 5828
rect 10818 5795 10852 5828
rect 11074 5795 11108 5828
rect 11330 5795 11364 5828
rect 11586 5795 11620 5828
rect 11842 5795 11876 5828
rect 12098 5795 12132 5828
rect 12354 5795 12388 5828
rect 12610 5795 12644 5828
rect 12866 5795 12900 5828
rect 13122 5795 13156 5828
rect 13378 5795 13412 5828
rect 13634 5795 13668 5828
rect 13890 5795 13924 5828
rect 14146 5795 14180 5828
rect 14402 5795 14436 5828
rect 14658 5795 14692 5828
rect 20399 5795 20433 5828
rect 20655 5795 20689 5828
rect 20911 5795 20945 5828
rect 21167 5795 21201 5828
rect 21423 5795 21457 5828
rect 21679 5795 21713 5828
rect 21935 5795 21969 5828
rect 22191 5795 22225 5828
rect 22447 5795 22481 5828
rect 22703 5795 22737 5828
rect 22959 5795 22993 5828
rect 23215 5795 23249 5828
rect 23471 5795 23505 5828
rect 23727 5795 23761 5828
rect 23983 5795 24017 5828
rect 24239 5795 24273 5828
rect 24495 5795 24529 5828
rect 24751 5795 24785 5828
rect 25007 5795 25041 5828
rect 25263 5795 25297 5828
rect 25519 5795 25553 5828
rect 25775 5795 25809 5828
rect 26031 5795 26065 5828
rect 26287 5795 26321 5828
rect 26543 5795 26577 5828
rect 26799 5795 26833 5828
rect 27055 5795 27089 5828
rect 27311 5795 27345 5828
rect 27567 5795 27601 5828
rect 27823 5795 27857 5828
rect 28079 5795 28113 5828
rect 28335 5795 28369 5828
rect 28591 5795 28625 5828
rect 37698 5820 37762 5826
rect 37698 5795 37704 5820
rect -363 5768 37704 5795
rect 37756 5768 37762 5820
rect -363 5763 37762 5768
rect 37698 5762 37762 5763
rect 38683 5736 38747 5742
rect 38683 5734 38689 5736
rect -363 5732 19999 5734
rect 20353 5732 38689 5734
rect -363 5728 38689 5732
rect -363 5690 -319 5728
rect -281 5690 -191 5728
rect -153 5690 481 5728
rect 519 5690 609 5728
rect 647 5690 737 5728
rect 775 5690 865 5728
rect 903 5690 1361 5728
rect 1399 5690 1489 5728
rect 1527 5690 1617 5728
rect 1655 5690 1745 5728
rect 1783 5690 1873 5728
rect 1911 5690 2001 5728
rect 2039 5690 2129 5728
rect 2167 5690 2257 5728
rect 2295 5690 2385 5728
rect 2423 5690 2980 5728
rect 3018 5690 3108 5728
rect 3146 5690 3236 5728
rect 3274 5690 3364 5728
rect 3402 5690 3492 5728
rect 3530 5690 3620 5728
rect 3658 5690 3748 5728
rect 3786 5690 3876 5728
rect 3914 5690 4004 5728
rect 4042 5690 4132 5728
rect 4170 5690 4260 5728
rect 4298 5690 4388 5728
rect 4426 5690 4516 5728
rect 4554 5690 5473 5728
rect 5511 5690 5601 5728
rect 5639 5690 5729 5728
rect 5767 5690 5857 5728
rect 5895 5690 5985 5728
rect 6023 5690 6113 5728
rect 6151 5690 6241 5728
rect 6279 5690 6369 5728
rect 6407 5690 6497 5728
rect 6535 5690 6625 5728
rect 6663 5690 6753 5728
rect 6791 5690 6881 5728
rect 6919 5690 7009 5728
rect 7047 5690 7137 5728
rect 7175 5690 7265 5728
rect 7303 5690 7393 5728
rect 7431 5690 7521 5728
rect 7559 5690 8057 5728
rect 8095 5690 8185 5728
rect 8223 5690 8313 5728
rect 8351 5690 8441 5728
rect 8479 5690 8569 5728
rect 8607 5690 8697 5728
rect 8735 5690 8825 5728
rect 8863 5690 8953 5728
rect 8991 5690 9081 5728
rect 9119 5690 9209 5728
rect 9247 5690 9337 5728
rect 9375 5690 9465 5728
rect 9503 5690 9593 5728
rect 9631 5690 9721 5728
rect 9759 5690 9849 5728
rect 9887 5690 9977 5728
rect 10015 5690 10105 5728
rect 10143 5690 10560 5728
rect 10598 5690 10688 5728
rect 10726 5690 10816 5728
rect 10854 5690 10944 5728
rect 10982 5690 11072 5728
rect 11110 5690 11200 5728
rect 11238 5690 11328 5728
rect 11366 5690 11456 5728
rect 11494 5690 11584 5728
rect 11622 5690 11712 5728
rect 11750 5690 11840 5728
rect 11878 5690 11968 5728
rect 12006 5690 12096 5728
rect 12134 5690 12224 5728
rect 12262 5690 12352 5728
rect 12390 5690 12480 5728
rect 12518 5690 12608 5728
rect 12646 5690 12736 5728
rect 12774 5690 12864 5728
rect 12902 5690 12992 5728
rect 13030 5690 13120 5728
rect 13158 5690 13248 5728
rect 13286 5690 13376 5728
rect 13414 5690 13504 5728
rect 13542 5690 13632 5728
rect 13670 5690 13760 5728
rect 13798 5690 13888 5728
rect 13926 5690 14016 5728
rect 14054 5690 14144 5728
rect 14182 5690 14272 5728
rect 14310 5690 14400 5728
rect 14438 5690 14528 5728
rect 14566 5690 14656 5728
rect 14694 5690 15821 5728
rect 15859 5690 15949 5728
rect 15987 5690 16077 5728
rect 16115 5690 16205 5728
rect 16243 5690 16333 5728
rect 16371 5690 16461 5728
rect 16499 5690 16589 5728
rect 16627 5690 16717 5728
rect 16755 5690 16845 5728
rect 16883 5690 16973 5728
rect 17011 5690 17101 5728
rect 17139 5690 17229 5728
rect 17267 5690 17357 5728
rect 17395 5690 17485 5728
rect 17523 5690 17613 5728
rect 17651 5690 17741 5728
rect 17779 5690 17869 5728
rect 17907 5690 17997 5728
rect 18035 5690 18125 5728
rect 18163 5690 18253 5728
rect 18291 5690 18381 5728
rect 18419 5690 18509 5728
rect 18547 5690 18637 5728
rect 18675 5690 18765 5728
rect 18803 5690 18893 5728
rect 18931 5690 19021 5728
rect 19059 5690 19149 5728
rect 19187 5690 19277 5728
rect 19315 5690 19405 5728
rect 19443 5690 19533 5728
rect 19571 5690 19661 5728
rect 19699 5690 19789 5728
rect 19827 5690 19917 5728
rect 19955 5690 20397 5728
rect 20435 5690 20525 5728
rect 20563 5690 20653 5728
rect 20691 5690 20781 5728
rect 20819 5690 20909 5728
rect 20947 5690 21037 5728
rect 21075 5690 21165 5728
rect 21203 5690 21293 5728
rect 21331 5690 21421 5728
rect 21459 5690 21549 5728
rect 21587 5690 21677 5728
rect 21715 5690 21805 5728
rect 21843 5690 21933 5728
rect 21971 5690 22061 5728
rect 22099 5690 22189 5728
rect 22227 5690 22317 5728
rect 22355 5690 22445 5728
rect 22483 5690 22573 5728
rect 22611 5690 22701 5728
rect 22739 5690 22829 5728
rect 22867 5690 22957 5728
rect 22995 5690 23085 5728
rect 23123 5690 23213 5728
rect 23251 5690 23341 5728
rect 23379 5690 23469 5728
rect 23507 5690 23597 5728
rect 23635 5690 23725 5728
rect 23763 5690 23853 5728
rect 23891 5690 23981 5728
rect 24019 5690 24109 5728
rect 24147 5690 24237 5728
rect 24275 5690 24365 5728
rect 24403 5690 24493 5728
rect 24531 5690 24621 5728
rect 24659 5690 24749 5728
rect 24787 5690 24877 5728
rect 24915 5690 25005 5728
rect 25043 5690 25133 5728
rect 25171 5690 25261 5728
rect 25299 5690 25389 5728
rect 25427 5690 25517 5728
rect 25555 5690 25645 5728
rect 25683 5690 25773 5728
rect 25811 5690 25901 5728
rect 25939 5690 26029 5728
rect 26067 5690 26157 5728
rect 26195 5690 26285 5728
rect 26323 5690 26413 5728
rect 26451 5690 26541 5728
rect 26579 5690 26669 5728
rect 26707 5690 26797 5728
rect 26835 5690 26925 5728
rect 26963 5690 27053 5728
rect 27091 5690 27181 5728
rect 27219 5690 27309 5728
rect 27347 5690 27437 5728
rect 27475 5690 27565 5728
rect 27603 5690 27693 5728
rect 27731 5690 27821 5728
rect 27859 5690 27949 5728
rect 27987 5690 28077 5728
rect 28115 5690 28205 5728
rect 28243 5690 28333 5728
rect 28371 5690 28461 5728
rect 28499 5690 28589 5728
rect 28627 5690 29365 5728
rect 29403 5690 29493 5728
rect 29531 5690 29621 5728
rect 29659 5690 29749 5728
rect 29787 5690 29877 5728
rect 29915 5690 30005 5728
rect 30043 5690 30133 5728
rect 30171 5690 30261 5728
rect 30299 5690 30389 5728
rect 30427 5690 30517 5728
rect 30555 5690 30645 5728
rect 30683 5690 30773 5728
rect 30811 5690 30901 5728
rect 30939 5690 31029 5728
rect 31067 5690 31157 5728
rect 31195 5690 31285 5728
rect 31323 5690 31413 5728
rect 31451 5690 31541 5728
rect 31579 5690 31669 5728
rect 31707 5690 31797 5728
rect 31835 5690 31925 5728
rect 31963 5690 32053 5728
rect 32091 5690 32181 5728
rect 32219 5690 32309 5728
rect 32347 5690 32437 5728
rect 32475 5690 32565 5728
rect 32603 5690 32693 5728
rect 32731 5690 32821 5728
rect 32859 5690 32949 5728
rect 32987 5690 33077 5728
rect 33115 5690 33205 5728
rect 33243 5690 33333 5728
rect 33371 5690 33461 5728
rect 33499 5690 33589 5728
rect 33627 5690 33717 5728
rect 33755 5690 33845 5728
rect 33883 5690 33973 5728
rect 34011 5690 34101 5728
rect 34139 5690 34229 5728
rect 34267 5690 34357 5728
rect 34395 5690 34485 5728
rect 34523 5690 34613 5728
rect 34651 5690 34741 5728
rect 34779 5690 34869 5728
rect 34907 5690 34997 5728
rect 35035 5690 35125 5728
rect 35163 5690 35253 5728
rect 35291 5690 35381 5728
rect 35419 5690 35509 5728
rect 35547 5690 35637 5728
rect 35675 5690 35765 5728
rect 35803 5690 35893 5728
rect 35931 5690 36021 5728
rect 36059 5690 36149 5728
rect 36187 5690 36277 5728
rect 36315 5690 36405 5728
rect 36443 5690 36533 5728
rect 36571 5690 36661 5728
rect 36699 5690 36789 5728
rect 36827 5690 36917 5728
rect 36955 5690 37045 5728
rect 37083 5690 37173 5728
rect 37211 5690 37301 5728
rect 37339 5690 37429 5728
rect 37467 5690 37557 5728
rect 37595 5690 38689 5728
rect -363 5686 38689 5690
rect -363 5684 19999 5686
rect 20353 5684 38689 5686
rect 38741 5684 38747 5736
rect 38683 5678 38747 5684
rect -363 5649 37762 5655
rect -363 5623 37704 5649
rect -317 5590 -283 5623
rect 611 5590 645 5623
rect 867 5590 901 5623
rect 1875 5590 1909 5623
rect 2131 5590 2165 5623
rect 2387 5590 2421 5623
rect 3494 5590 3528 5623
rect 3750 5590 3784 5623
rect 4006 5590 4040 5623
rect 4262 5590 4296 5623
rect 4518 5590 4552 5623
rect 8059 5590 8093 5623
rect 8315 5590 8349 5623
rect 8571 5590 8605 5623
rect 8827 5590 8861 5623
rect 9083 5590 9117 5623
rect 9339 5590 9373 5623
rect 9595 5590 9629 5623
rect 9851 5590 9885 5623
rect 10107 5590 10141 5623
rect 15823 5590 15857 5623
rect 16079 5590 16113 5623
rect 16335 5590 16369 5623
rect 16591 5590 16625 5623
rect 16847 5590 16881 5623
rect 17103 5590 17137 5623
rect 17359 5590 17393 5623
rect 17615 5590 17649 5623
rect 17871 5590 17905 5623
rect 18127 5590 18161 5623
rect 18383 5590 18417 5623
rect 18639 5590 18673 5623
rect 18895 5590 18929 5623
rect 19151 5590 19185 5623
rect 19407 5590 19441 5623
rect 19663 5590 19697 5623
rect 19919 5590 19953 5623
rect 29367 5590 29401 5623
rect 29623 5590 29657 5623
rect 29879 5590 29913 5623
rect 30135 5590 30169 5623
rect 30391 5590 30425 5623
rect 30647 5590 30681 5623
rect 30903 5590 30937 5623
rect 31159 5590 31193 5623
rect 31415 5590 31449 5623
rect 31671 5590 31705 5623
rect 31927 5590 31961 5623
rect 32183 5590 32217 5623
rect 32439 5590 32473 5623
rect 32695 5590 32729 5623
rect 32951 5590 32985 5623
rect 33207 5590 33241 5623
rect 33463 5590 33497 5623
rect 33719 5590 33753 5623
rect 33975 5590 34009 5623
rect 34231 5590 34265 5623
rect 34487 5590 34521 5623
rect 34743 5590 34777 5623
rect 34999 5590 35033 5623
rect 35255 5590 35289 5623
rect 35511 5590 35545 5623
rect 35767 5590 35801 5623
rect 36023 5590 36057 5623
rect 36279 5590 36313 5623
rect 36535 5590 36569 5623
rect 36791 5590 36825 5623
rect 37047 5590 37081 5623
rect 37303 5590 37337 5623
rect 37559 5590 37593 5623
rect 37698 5597 37704 5623
rect 37756 5597 37762 5649
rect 37698 5591 37762 5597
rect -323 5578 -277 5590
rect -323 5434 -317 5578
rect -283 5434 -277 5578
rect -323 5422 -277 5434
rect -195 5578 -149 5590
rect -195 5434 -189 5578
rect -155 5434 -149 5578
rect -195 5422 -149 5434
rect 605 5578 651 5590
rect 605 5434 611 5578
rect 645 5434 651 5578
rect 605 5422 651 5434
rect 733 5578 779 5590
rect 733 5434 739 5578
rect 773 5434 779 5578
rect 733 5422 779 5434
rect 861 5578 907 5590
rect 861 5434 867 5578
rect 901 5434 907 5578
rect 1869 5578 1915 5590
rect 861 5422 907 5434
rect 958 5445 1030 5451
rect -391 5382 -319 5388
rect -391 5325 -385 5382
rect -325 5325 -319 5382
rect -391 5319 -319 5325
rect -189 5356 -155 5422
rect -95 5363 -31 5369
rect -95 5356 -89 5363
rect -189 5322 -89 5356
rect -189 5290 -155 5322
rect -95 5311 -89 5322
rect -37 5311 -31 5363
rect -95 5305 -31 5311
rect 739 5354 773 5422
rect 958 5388 964 5445
rect 1024 5388 1030 5445
rect 1869 5434 1875 5578
rect 1909 5434 1915 5578
rect 1869 5422 1915 5434
rect 1997 5578 2043 5590
rect 1997 5434 2003 5578
rect 2037 5434 2043 5578
rect 1997 5422 2043 5434
rect 2125 5578 2171 5590
rect 2125 5434 2131 5578
rect 2165 5434 2171 5578
rect 2125 5422 2171 5434
rect 2253 5578 2299 5590
rect 2253 5434 2259 5578
rect 2293 5434 2299 5578
rect 2253 5422 2299 5434
rect 2381 5578 2427 5590
rect 2381 5434 2387 5578
rect 2421 5434 2427 5578
rect 3488 5578 3534 5590
rect 2381 5422 2427 5434
rect 2487 5445 2559 5451
rect 958 5382 1030 5388
rect 1750 5358 1814 5364
rect 739 5348 1026 5354
rect 739 5318 968 5348
rect 739 5290 773 5318
rect 962 5296 968 5318
rect 1020 5296 1026 5348
rect 1750 5306 1756 5358
rect 1808 5348 1814 5358
rect 2003 5348 2037 5422
rect 2259 5354 2293 5422
rect 2487 5388 2493 5445
rect 2553 5388 2559 5445
rect 3488 5434 3494 5578
rect 3528 5434 3534 5578
rect 3488 5422 3534 5434
rect 3616 5578 3662 5590
rect 3616 5434 3622 5578
rect 3656 5434 3662 5578
rect 3616 5422 3662 5434
rect 3744 5578 3790 5590
rect 3744 5434 3750 5578
rect 3784 5434 3790 5578
rect 3744 5422 3790 5434
rect 3872 5578 3918 5590
rect 3872 5434 3878 5578
rect 3912 5434 3918 5578
rect 3872 5422 3918 5434
rect 4000 5578 4046 5590
rect 4000 5434 4006 5578
rect 4040 5434 4046 5578
rect 4000 5422 4046 5434
rect 4128 5578 4174 5590
rect 4128 5434 4134 5578
rect 4168 5434 4174 5578
rect 4128 5422 4174 5434
rect 4256 5578 4302 5590
rect 4256 5434 4262 5578
rect 4296 5434 4302 5578
rect 4256 5422 4302 5434
rect 4384 5578 4430 5590
rect 4384 5434 4390 5578
rect 4424 5434 4430 5578
rect 4384 5422 4430 5434
rect 4512 5578 4558 5590
rect 4512 5434 4518 5578
rect 4552 5434 4558 5578
rect 8053 5578 8099 5590
rect 4512 5422 4558 5434
rect 4658 5454 4730 5460
rect 2487 5382 2559 5388
rect 3408 5371 3472 5377
rect 2259 5348 2544 5354
rect 1808 5323 2486 5348
rect 1808 5319 2293 5323
rect 1808 5306 1814 5319
rect 1750 5300 1814 5306
rect 962 5290 1026 5296
rect 2003 5290 2037 5319
rect 2259 5290 2293 5319
rect 2480 5296 2486 5323
rect 2538 5296 2544 5348
rect 3408 5319 3414 5371
rect 3466 5348 3472 5371
rect 3622 5348 3656 5422
rect 3878 5348 3912 5422
rect 4134 5348 4168 5422
rect 4390 5348 4424 5422
rect 4658 5397 4664 5454
rect 4724 5397 4730 5454
rect 4658 5391 4730 5397
rect 7916 5439 7988 5445
rect 7916 5382 7922 5439
rect 7982 5382 7988 5439
rect 8053 5434 8059 5578
rect 8093 5434 8099 5578
rect 8053 5422 8099 5434
rect 8181 5578 8227 5590
rect 8181 5434 8187 5578
rect 8221 5434 8227 5578
rect 8181 5422 8227 5434
rect 8309 5578 8355 5590
rect 8309 5434 8315 5578
rect 8349 5434 8355 5578
rect 8309 5422 8355 5434
rect 8437 5578 8483 5590
rect 8437 5434 8443 5578
rect 8477 5434 8483 5578
rect 8437 5422 8483 5434
rect 8565 5578 8611 5590
rect 8565 5434 8571 5578
rect 8605 5434 8611 5578
rect 8565 5422 8611 5434
rect 8693 5578 8739 5590
rect 8693 5434 8699 5578
rect 8733 5434 8739 5578
rect 8693 5422 8739 5434
rect 8821 5578 8867 5590
rect 8821 5434 8827 5578
rect 8861 5434 8867 5578
rect 8821 5422 8867 5434
rect 8949 5578 8995 5590
rect 8949 5434 8955 5578
rect 8989 5434 8995 5578
rect 8949 5422 8995 5434
rect 9077 5578 9123 5590
rect 9077 5434 9083 5578
rect 9117 5434 9123 5578
rect 9077 5422 9123 5434
rect 9205 5578 9251 5590
rect 9205 5434 9211 5578
rect 9245 5434 9251 5578
rect 9205 5422 9251 5434
rect 9333 5578 9379 5590
rect 9333 5434 9339 5578
rect 9373 5434 9379 5578
rect 9333 5422 9379 5434
rect 9461 5578 9507 5590
rect 9461 5434 9467 5578
rect 9501 5434 9507 5578
rect 9461 5422 9507 5434
rect 9589 5578 9635 5590
rect 9589 5434 9595 5578
rect 9629 5434 9635 5578
rect 9589 5422 9635 5434
rect 9717 5578 9763 5590
rect 9717 5434 9723 5578
rect 9757 5434 9763 5578
rect 9717 5422 9763 5434
rect 9845 5578 9891 5590
rect 9845 5434 9851 5578
rect 9885 5434 9891 5578
rect 9845 5422 9891 5434
rect 9973 5578 10019 5590
rect 9973 5434 9979 5578
rect 10013 5434 10019 5578
rect 9973 5422 10019 5434
rect 10101 5578 10147 5590
rect 10101 5434 10107 5578
rect 10141 5434 10147 5578
rect 10101 5422 10147 5434
rect 15817 5578 15863 5590
rect 15817 5434 15823 5578
rect 15857 5434 15863 5578
rect 15817 5422 15863 5434
rect 15945 5578 15991 5590
rect 15945 5434 15951 5578
rect 15985 5434 15991 5578
rect 15945 5422 15991 5434
rect 16073 5578 16119 5590
rect 16073 5434 16079 5578
rect 16113 5434 16119 5578
rect 16073 5422 16119 5434
rect 16201 5578 16247 5590
rect 16201 5434 16207 5578
rect 16241 5434 16247 5578
rect 16201 5422 16247 5434
rect 16329 5578 16375 5590
rect 16329 5434 16335 5578
rect 16369 5434 16375 5578
rect 16329 5422 16375 5434
rect 16457 5578 16503 5590
rect 16457 5434 16463 5578
rect 16497 5434 16503 5578
rect 16457 5422 16503 5434
rect 16585 5578 16631 5590
rect 16585 5434 16591 5578
rect 16625 5434 16631 5578
rect 16585 5422 16631 5434
rect 16713 5578 16759 5590
rect 16713 5434 16719 5578
rect 16753 5434 16759 5578
rect 16713 5422 16759 5434
rect 16841 5578 16887 5590
rect 16841 5434 16847 5578
rect 16881 5434 16887 5578
rect 16841 5422 16887 5434
rect 16969 5578 17015 5590
rect 16969 5434 16975 5578
rect 17009 5434 17015 5578
rect 16969 5422 17015 5434
rect 17097 5578 17143 5590
rect 17097 5434 17103 5578
rect 17137 5434 17143 5578
rect 17097 5422 17143 5434
rect 17225 5578 17271 5590
rect 17225 5434 17231 5578
rect 17265 5434 17271 5578
rect 17225 5422 17271 5434
rect 17353 5578 17399 5590
rect 17353 5434 17359 5578
rect 17393 5434 17399 5578
rect 17353 5422 17399 5434
rect 17481 5578 17527 5590
rect 17481 5434 17487 5578
rect 17521 5434 17527 5578
rect 17481 5422 17527 5434
rect 17609 5578 17655 5590
rect 17609 5434 17615 5578
rect 17649 5434 17655 5578
rect 17609 5422 17655 5434
rect 17737 5578 17783 5590
rect 17737 5434 17743 5578
rect 17777 5434 17783 5578
rect 17737 5422 17783 5434
rect 17865 5578 17911 5590
rect 17865 5434 17871 5578
rect 17905 5434 17911 5578
rect 17865 5422 17911 5434
rect 17993 5578 18039 5590
rect 17993 5434 17999 5578
rect 18033 5434 18039 5578
rect 17993 5422 18039 5434
rect 18121 5578 18167 5590
rect 18121 5434 18127 5578
rect 18161 5434 18167 5578
rect 18121 5422 18167 5434
rect 18249 5578 18295 5590
rect 18249 5434 18255 5578
rect 18289 5434 18295 5578
rect 18249 5422 18295 5434
rect 18377 5578 18423 5590
rect 18377 5434 18383 5578
rect 18417 5434 18423 5578
rect 18377 5422 18423 5434
rect 18505 5578 18551 5590
rect 18505 5434 18511 5578
rect 18545 5434 18551 5578
rect 18505 5422 18551 5434
rect 18633 5578 18679 5590
rect 18633 5434 18639 5578
rect 18673 5434 18679 5578
rect 18633 5422 18679 5434
rect 18761 5578 18807 5590
rect 18761 5434 18767 5578
rect 18801 5434 18807 5578
rect 18761 5422 18807 5434
rect 18889 5578 18935 5590
rect 18889 5434 18895 5578
rect 18929 5434 18935 5578
rect 18889 5422 18935 5434
rect 19017 5578 19063 5590
rect 19017 5434 19023 5578
rect 19057 5434 19063 5578
rect 19017 5422 19063 5434
rect 19145 5578 19191 5590
rect 19145 5434 19151 5578
rect 19185 5434 19191 5578
rect 19145 5422 19191 5434
rect 19273 5578 19319 5590
rect 19273 5434 19279 5578
rect 19313 5434 19319 5578
rect 19273 5422 19319 5434
rect 19401 5578 19447 5590
rect 19401 5434 19407 5578
rect 19441 5434 19447 5578
rect 19401 5422 19447 5434
rect 19529 5578 19575 5590
rect 19529 5434 19535 5578
rect 19569 5434 19575 5578
rect 19529 5422 19575 5434
rect 19657 5578 19703 5590
rect 19657 5434 19663 5578
rect 19697 5434 19703 5578
rect 19657 5422 19703 5434
rect 19785 5578 19831 5590
rect 19785 5434 19791 5578
rect 19825 5434 19831 5578
rect 19785 5422 19831 5434
rect 19913 5578 19959 5590
rect 19913 5434 19919 5578
rect 19953 5434 19959 5578
rect 19913 5422 19959 5434
rect 29361 5578 29407 5590
rect 29361 5434 29367 5578
rect 29401 5434 29407 5578
rect 29361 5422 29407 5434
rect 29489 5578 29535 5590
rect 29489 5434 29495 5578
rect 29529 5434 29535 5578
rect 29489 5422 29535 5434
rect 29617 5578 29663 5590
rect 29617 5434 29623 5578
rect 29657 5434 29663 5578
rect 29617 5422 29663 5434
rect 29745 5578 29791 5590
rect 29745 5434 29751 5578
rect 29785 5434 29791 5578
rect 29745 5422 29791 5434
rect 29873 5578 29919 5590
rect 29873 5434 29879 5578
rect 29913 5434 29919 5578
rect 29873 5422 29919 5434
rect 30001 5578 30047 5590
rect 30001 5434 30007 5578
rect 30041 5434 30047 5578
rect 30001 5422 30047 5434
rect 30129 5578 30175 5590
rect 30129 5434 30135 5578
rect 30169 5434 30175 5578
rect 30129 5422 30175 5434
rect 30257 5578 30303 5590
rect 30257 5434 30263 5578
rect 30297 5434 30303 5578
rect 30257 5422 30303 5434
rect 30385 5578 30431 5590
rect 30385 5434 30391 5578
rect 30425 5434 30431 5578
rect 30385 5422 30431 5434
rect 30513 5578 30559 5590
rect 30513 5434 30519 5578
rect 30553 5434 30559 5578
rect 30513 5422 30559 5434
rect 30641 5578 30687 5590
rect 30641 5434 30647 5578
rect 30681 5434 30687 5578
rect 30641 5422 30687 5434
rect 30769 5578 30815 5590
rect 30769 5434 30775 5578
rect 30809 5434 30815 5578
rect 30769 5422 30815 5434
rect 30897 5578 30943 5590
rect 30897 5434 30903 5578
rect 30937 5434 30943 5578
rect 30897 5422 30943 5434
rect 31025 5578 31071 5590
rect 31025 5434 31031 5578
rect 31065 5434 31071 5578
rect 31025 5422 31071 5434
rect 31153 5578 31199 5590
rect 31153 5434 31159 5578
rect 31193 5434 31199 5578
rect 31153 5422 31199 5434
rect 31281 5578 31327 5590
rect 31281 5434 31287 5578
rect 31321 5434 31327 5578
rect 31281 5422 31327 5434
rect 31409 5578 31455 5590
rect 31409 5434 31415 5578
rect 31449 5434 31455 5578
rect 31409 5422 31455 5434
rect 31537 5578 31583 5590
rect 31537 5434 31543 5578
rect 31577 5434 31583 5578
rect 31537 5422 31583 5434
rect 31665 5578 31711 5590
rect 31665 5434 31671 5578
rect 31705 5434 31711 5578
rect 31665 5422 31711 5434
rect 31793 5578 31839 5590
rect 31793 5434 31799 5578
rect 31833 5434 31839 5578
rect 31793 5422 31839 5434
rect 31921 5578 31967 5590
rect 31921 5434 31927 5578
rect 31961 5434 31967 5578
rect 31921 5422 31967 5434
rect 32049 5578 32095 5590
rect 32049 5434 32055 5578
rect 32089 5434 32095 5578
rect 32049 5422 32095 5434
rect 32177 5578 32223 5590
rect 32177 5434 32183 5578
rect 32217 5434 32223 5578
rect 32177 5422 32223 5434
rect 32305 5578 32351 5590
rect 32305 5434 32311 5578
rect 32345 5434 32351 5578
rect 32305 5422 32351 5434
rect 32433 5578 32479 5590
rect 32433 5434 32439 5578
rect 32473 5434 32479 5578
rect 32433 5422 32479 5434
rect 32561 5578 32607 5590
rect 32561 5434 32567 5578
rect 32601 5434 32607 5578
rect 32561 5422 32607 5434
rect 32689 5578 32735 5590
rect 32689 5434 32695 5578
rect 32729 5434 32735 5578
rect 32689 5422 32735 5434
rect 32817 5578 32863 5590
rect 32817 5434 32823 5578
rect 32857 5434 32863 5578
rect 32817 5422 32863 5434
rect 32945 5578 32991 5590
rect 32945 5434 32951 5578
rect 32985 5434 32991 5578
rect 32945 5422 32991 5434
rect 33073 5578 33119 5590
rect 33073 5434 33079 5578
rect 33113 5434 33119 5578
rect 33073 5422 33119 5434
rect 33201 5578 33247 5590
rect 33201 5434 33207 5578
rect 33241 5434 33247 5578
rect 33201 5422 33247 5434
rect 33329 5578 33375 5590
rect 33329 5434 33335 5578
rect 33369 5434 33375 5578
rect 33329 5422 33375 5434
rect 33457 5578 33503 5590
rect 33457 5434 33463 5578
rect 33497 5434 33503 5578
rect 33457 5422 33503 5434
rect 33585 5578 33631 5590
rect 33585 5434 33591 5578
rect 33625 5434 33631 5578
rect 33585 5422 33631 5434
rect 33713 5578 33759 5590
rect 33713 5434 33719 5578
rect 33753 5434 33759 5578
rect 33713 5422 33759 5434
rect 33841 5578 33887 5590
rect 33841 5434 33847 5578
rect 33881 5434 33887 5578
rect 33841 5422 33887 5434
rect 33969 5578 34015 5590
rect 33969 5434 33975 5578
rect 34009 5434 34015 5578
rect 33969 5422 34015 5434
rect 34097 5578 34143 5590
rect 34097 5434 34103 5578
rect 34137 5434 34143 5578
rect 34097 5422 34143 5434
rect 34225 5578 34271 5590
rect 34225 5434 34231 5578
rect 34265 5434 34271 5578
rect 34225 5422 34271 5434
rect 34353 5578 34399 5590
rect 34353 5434 34359 5578
rect 34393 5434 34399 5578
rect 34353 5422 34399 5434
rect 34481 5578 34527 5590
rect 34481 5434 34487 5578
rect 34521 5434 34527 5578
rect 34481 5422 34527 5434
rect 34609 5578 34655 5590
rect 34609 5434 34615 5578
rect 34649 5434 34655 5578
rect 34609 5422 34655 5434
rect 34737 5578 34783 5590
rect 34737 5434 34743 5578
rect 34777 5434 34783 5578
rect 34737 5422 34783 5434
rect 34865 5578 34911 5590
rect 34865 5434 34871 5578
rect 34905 5434 34911 5578
rect 34865 5422 34911 5434
rect 34993 5578 35039 5590
rect 34993 5434 34999 5578
rect 35033 5434 35039 5578
rect 34993 5422 35039 5434
rect 35121 5578 35167 5590
rect 35121 5434 35127 5578
rect 35161 5434 35167 5578
rect 35121 5422 35167 5434
rect 35249 5578 35295 5590
rect 35249 5434 35255 5578
rect 35289 5434 35295 5578
rect 35249 5422 35295 5434
rect 35377 5578 35423 5590
rect 35377 5434 35383 5578
rect 35417 5434 35423 5578
rect 35377 5422 35423 5434
rect 35505 5578 35551 5590
rect 35505 5434 35511 5578
rect 35545 5434 35551 5578
rect 35505 5422 35551 5434
rect 35633 5578 35679 5590
rect 35633 5434 35639 5578
rect 35673 5434 35679 5578
rect 35633 5422 35679 5434
rect 35761 5578 35807 5590
rect 35761 5434 35767 5578
rect 35801 5434 35807 5578
rect 35761 5422 35807 5434
rect 35889 5578 35935 5590
rect 35889 5434 35895 5578
rect 35929 5434 35935 5578
rect 35889 5422 35935 5434
rect 36017 5578 36063 5590
rect 36017 5434 36023 5578
rect 36057 5434 36063 5578
rect 36017 5422 36063 5434
rect 36145 5578 36191 5590
rect 36145 5434 36151 5578
rect 36185 5434 36191 5578
rect 36145 5422 36191 5434
rect 36273 5578 36319 5590
rect 36273 5434 36279 5578
rect 36313 5434 36319 5578
rect 36273 5422 36319 5434
rect 36401 5578 36447 5590
rect 36401 5434 36407 5578
rect 36441 5434 36447 5578
rect 36401 5422 36447 5434
rect 36529 5578 36575 5590
rect 36529 5434 36535 5578
rect 36569 5434 36575 5578
rect 36529 5422 36575 5434
rect 36657 5578 36703 5590
rect 36657 5434 36663 5578
rect 36697 5434 36703 5578
rect 36657 5422 36703 5434
rect 36785 5578 36831 5590
rect 36785 5434 36791 5578
rect 36825 5434 36831 5578
rect 36785 5422 36831 5434
rect 36913 5578 36959 5590
rect 36913 5434 36919 5578
rect 36953 5434 36959 5578
rect 36913 5422 36959 5434
rect 37041 5578 37087 5590
rect 37041 5434 37047 5578
rect 37081 5434 37087 5578
rect 37041 5422 37087 5434
rect 37169 5578 37215 5590
rect 37169 5434 37175 5578
rect 37209 5434 37215 5578
rect 37169 5422 37215 5434
rect 37297 5578 37343 5590
rect 37297 5434 37303 5578
rect 37337 5434 37343 5578
rect 37297 5422 37343 5434
rect 37425 5578 37471 5590
rect 37425 5434 37431 5578
rect 37465 5434 37471 5578
rect 37425 5422 37471 5434
rect 37553 5578 37599 5590
rect 37553 5434 37559 5578
rect 37593 5434 37599 5578
rect 37553 5422 37599 5434
rect 7916 5376 7988 5382
rect 8187 5348 8221 5422
rect 8443 5384 8477 5422
rect 8381 5378 8477 5384
rect 8381 5348 8387 5378
rect 3466 5342 4684 5348
rect 8187 5347 8387 5348
rect 3466 5319 4626 5342
rect 3408 5313 3472 5319
rect 2480 5290 2544 5296
rect 3622 5290 3656 5319
rect 3878 5290 3912 5319
rect 4134 5290 4168 5319
rect 4390 5290 4424 5319
rect 4620 5290 4626 5319
rect 4678 5290 4684 5342
rect -323 5278 -277 5290
rect -323 5218 -317 5278
rect -283 5218 -277 5278
rect -323 5206 -277 5218
rect -195 5278 -149 5290
rect -195 5218 -189 5278
rect -155 5218 -149 5278
rect -195 5206 -149 5218
rect 605 5278 651 5290
rect 605 5218 611 5278
rect 645 5218 651 5278
rect 605 5206 651 5218
rect 733 5278 779 5290
rect 733 5218 739 5278
rect 773 5218 779 5278
rect 733 5206 779 5218
rect 861 5278 907 5290
rect 861 5218 867 5278
rect 901 5218 907 5278
rect 861 5206 907 5218
rect 1869 5278 1915 5290
rect 1869 5218 1875 5278
rect 1909 5218 1915 5278
rect 1869 5206 1915 5218
rect 1997 5278 2043 5290
rect 1997 5218 2003 5278
rect 2037 5218 2043 5278
rect 1997 5206 2043 5218
rect 2125 5278 2171 5290
rect 2125 5218 2131 5278
rect 2165 5218 2171 5278
rect 2125 5206 2171 5218
rect 2253 5278 2299 5290
rect 2253 5218 2259 5278
rect 2293 5218 2299 5278
rect 2253 5206 2299 5218
rect 2381 5278 2427 5290
rect 2381 5218 2387 5278
rect 2421 5218 2427 5278
rect 2381 5206 2427 5218
rect 3488 5278 3534 5290
rect 3488 5218 3494 5278
rect 3528 5218 3534 5278
rect 3488 5206 3534 5218
rect 3616 5278 3662 5290
rect 3616 5218 3622 5278
rect 3656 5218 3662 5278
rect 3616 5206 3662 5218
rect 3744 5278 3790 5290
rect 3744 5218 3750 5278
rect 3784 5218 3790 5278
rect 3744 5206 3790 5218
rect 3872 5278 3918 5290
rect 3872 5218 3878 5278
rect 3912 5218 3918 5278
rect 3872 5206 3918 5218
rect 4000 5278 4046 5290
rect 4000 5218 4006 5278
rect 4040 5218 4046 5278
rect 4000 5206 4046 5218
rect 4128 5278 4174 5290
rect 4128 5218 4134 5278
rect 4168 5218 4174 5278
rect 4128 5206 4174 5218
rect 4256 5278 4302 5290
rect 4256 5218 4262 5278
rect 4296 5218 4302 5278
rect 4256 5206 4302 5218
rect 4384 5278 4430 5290
rect 4384 5218 4390 5278
rect 4424 5218 4430 5278
rect 4384 5206 4430 5218
rect 4512 5278 4558 5290
rect 4620 5284 4684 5290
rect 7923 5341 8387 5347
rect 7923 5289 7929 5341
rect 7981 5326 8387 5341
rect 8439 5348 8477 5378
rect 8699 5348 8733 5422
rect 8955 5383 8989 5422
rect 8955 5377 9051 5383
rect 8955 5348 8993 5377
rect 8439 5326 8993 5348
rect 7981 5325 8993 5326
rect 9045 5348 9051 5377
rect 9211 5348 9245 5422
rect 9467 5348 9501 5422
rect 9593 5377 9657 5383
rect 9593 5348 9599 5377
rect 9045 5325 9599 5348
rect 9651 5348 9657 5377
rect 9723 5348 9757 5422
rect 9979 5353 10013 5422
rect 15685 5408 15757 5414
rect 10200 5362 10264 5368
rect 10200 5353 10206 5362
rect 9979 5348 10206 5353
rect 9651 5325 10206 5348
rect 7981 5324 10206 5325
rect 7981 5319 10013 5324
rect 7981 5318 8221 5319
rect 7981 5289 7987 5318
rect 8187 5290 8221 5318
rect 8443 5290 8477 5319
rect 8699 5290 8733 5319
rect 8955 5290 8989 5319
rect 9211 5290 9245 5319
rect 9467 5290 9501 5319
rect 9723 5290 9757 5319
rect 9979 5290 10013 5319
rect 10200 5310 10206 5324
rect 10258 5310 10264 5362
rect 15685 5351 15691 5408
rect 15751 5351 15757 5408
rect 15685 5345 15757 5351
rect 15786 5376 15850 5382
rect 15786 5324 15792 5376
rect 15844 5362 15850 5376
rect 15951 5362 15985 5422
rect 15844 5348 15985 5362
rect 16207 5348 16241 5422
rect 16463 5382 16497 5422
rect 16402 5376 16497 5382
rect 16402 5348 16408 5376
rect 15844 5329 16408 5348
rect 15844 5324 15850 5329
rect 15786 5318 15850 5324
rect 15951 5324 16408 5329
rect 16460 5348 16497 5376
rect 16719 5348 16753 5422
rect 16975 5348 17009 5422
rect 17231 5348 17265 5422
rect 17487 5348 17521 5422
rect 17743 5348 17777 5422
rect 17999 5348 18033 5422
rect 18255 5348 18289 5422
rect 18511 5348 18545 5422
rect 18767 5348 18801 5422
rect 19023 5348 19057 5422
rect 19279 5348 19313 5422
rect 19535 5348 19569 5422
rect 19791 5348 19825 5422
rect 16460 5347 19825 5348
rect 20023 5358 20087 5364
rect 20023 5347 20029 5358
rect 16460 5324 20029 5347
rect 15951 5319 20029 5324
rect 10200 5304 10264 5310
rect 15951 5290 15985 5319
rect 16207 5290 16241 5319
rect 16402 5318 16497 5319
rect 16463 5290 16497 5318
rect 16719 5290 16753 5319
rect 16975 5290 17009 5319
rect 17231 5290 17265 5319
rect 17487 5290 17521 5319
rect 17743 5290 17777 5319
rect 17999 5290 18033 5319
rect 18255 5290 18289 5319
rect 18511 5290 18545 5319
rect 18767 5290 18801 5319
rect 19023 5290 19057 5319
rect 19279 5290 19313 5319
rect 19535 5290 19569 5319
rect 19791 5318 20029 5319
rect 19791 5290 19825 5318
rect 20023 5306 20029 5318
rect 20081 5306 20087 5358
rect 29495 5349 29529 5422
rect 20023 5300 20087 5306
rect 29239 5348 29529 5349
rect 29751 5348 29785 5422
rect 29846 5378 29910 5384
rect 29846 5348 29852 5378
rect 29239 5343 29852 5348
rect 29239 5291 29245 5343
rect 29297 5326 29852 5343
rect 29904 5348 29910 5378
rect 30007 5348 30041 5422
rect 30263 5348 30297 5422
rect 30519 5383 30553 5422
rect 30455 5377 30553 5383
rect 30455 5348 30461 5377
rect 29904 5326 30461 5348
rect 29297 5325 30461 5326
rect 30513 5348 30553 5377
rect 30775 5348 30809 5422
rect 31031 5383 31065 5422
rect 31031 5377 31121 5383
rect 31031 5348 31063 5377
rect 30513 5325 31063 5348
rect 31115 5348 31121 5377
rect 31287 5348 31321 5422
rect 31543 5348 31577 5422
rect 31663 5377 31727 5383
rect 31663 5348 31669 5377
rect 31115 5325 31669 5348
rect 31721 5348 31727 5377
rect 31799 5348 31833 5422
rect 32055 5348 32089 5422
rect 32311 5383 32345 5422
rect 32269 5377 32345 5383
rect 32269 5348 32275 5377
rect 31721 5325 32275 5348
rect 32327 5348 32345 5377
rect 32567 5348 32601 5422
rect 32823 5348 32857 5422
rect 32885 5377 32949 5383
rect 32885 5348 32891 5377
rect 32327 5325 32891 5348
rect 32943 5348 32949 5377
rect 33079 5348 33113 5422
rect 33335 5348 33369 5422
rect 33481 5377 33545 5383
rect 33481 5348 33487 5377
rect 32943 5325 33487 5348
rect 33539 5348 33545 5377
rect 33591 5348 33625 5422
rect 33847 5348 33881 5422
rect 34103 5383 34137 5422
rect 34087 5377 34151 5383
rect 34087 5348 34093 5377
rect 33539 5325 34093 5348
rect 34145 5348 34151 5377
rect 34359 5348 34393 5422
rect 34615 5348 34649 5422
rect 34694 5377 34758 5383
rect 34694 5348 34700 5377
rect 34145 5325 34700 5348
rect 34752 5348 34758 5377
rect 34871 5348 34905 5422
rect 35127 5348 35161 5422
rect 35291 5376 35355 5382
rect 35291 5348 35297 5376
rect 34752 5325 35297 5348
rect 29297 5324 35297 5325
rect 35349 5348 35355 5376
rect 35383 5348 35417 5422
rect 35639 5348 35673 5422
rect 35895 5382 35929 5422
rect 35895 5376 35970 5382
rect 35895 5348 35912 5376
rect 35349 5324 35912 5348
rect 35964 5348 35970 5376
rect 36151 5348 36185 5422
rect 36407 5348 36441 5422
rect 36512 5377 36576 5383
rect 36512 5348 36518 5377
rect 35964 5325 36518 5348
rect 36570 5348 36576 5377
rect 36663 5348 36697 5422
rect 36919 5348 36953 5422
rect 37175 5383 37209 5422
rect 37118 5377 37209 5383
rect 37118 5348 37124 5377
rect 36570 5325 37124 5348
rect 37176 5348 37209 5377
rect 37431 5349 37465 5422
rect 37720 5359 37784 5365
rect 37720 5349 37726 5359
rect 37431 5348 37726 5349
rect 37176 5325 37726 5348
rect 35964 5324 37726 5325
rect 29297 5320 37726 5324
rect 29297 5291 29303 5320
rect 7923 5283 7987 5289
rect 4512 5218 4518 5278
rect 4552 5218 4558 5278
rect 4512 5206 4558 5218
rect 8053 5278 8099 5290
rect 8053 5218 8059 5278
rect 8093 5218 8099 5278
rect 8053 5206 8099 5218
rect 8181 5278 8227 5290
rect 8181 5218 8187 5278
rect 8221 5218 8227 5278
rect 8181 5206 8227 5218
rect 8309 5278 8355 5290
rect 8309 5218 8315 5278
rect 8349 5218 8355 5278
rect 8309 5206 8355 5218
rect 8437 5278 8483 5290
rect 8437 5218 8443 5278
rect 8477 5218 8483 5278
rect 8437 5206 8483 5218
rect 8565 5278 8611 5290
rect 8565 5218 8571 5278
rect 8605 5218 8611 5278
rect 8565 5206 8611 5218
rect 8693 5278 8739 5290
rect 8693 5218 8699 5278
rect 8733 5218 8739 5278
rect 8693 5206 8739 5218
rect 8821 5278 8867 5290
rect 8821 5218 8827 5278
rect 8861 5218 8867 5278
rect 8821 5206 8867 5218
rect 8949 5278 8995 5290
rect 8949 5218 8955 5278
rect 8989 5218 8995 5278
rect 8949 5206 8995 5218
rect 9077 5278 9123 5290
rect 9077 5218 9083 5278
rect 9117 5218 9123 5278
rect 9077 5206 9123 5218
rect 9205 5278 9251 5290
rect 9205 5218 9211 5278
rect 9245 5218 9251 5278
rect 9205 5206 9251 5218
rect 9333 5278 9379 5290
rect 9333 5218 9339 5278
rect 9373 5218 9379 5278
rect 9333 5206 9379 5218
rect 9461 5278 9507 5290
rect 9461 5218 9467 5278
rect 9501 5218 9507 5278
rect 9461 5206 9507 5218
rect 9589 5278 9635 5290
rect 9589 5218 9595 5278
rect 9629 5218 9635 5278
rect 9589 5206 9635 5218
rect 9717 5278 9763 5290
rect 9717 5218 9723 5278
rect 9757 5218 9763 5278
rect 9717 5206 9763 5218
rect 9845 5278 9891 5290
rect 9845 5218 9851 5278
rect 9885 5218 9891 5278
rect 9845 5206 9891 5218
rect 9973 5278 10019 5290
rect 9973 5218 9979 5278
rect 10013 5218 10019 5278
rect 9973 5206 10019 5218
rect 10101 5278 10147 5290
rect 10101 5218 10107 5278
rect 10141 5218 10147 5278
rect 10101 5206 10147 5218
rect 15817 5278 15863 5290
rect 15817 5218 15823 5278
rect 15857 5218 15863 5278
rect 15817 5206 15863 5218
rect 15945 5278 15991 5290
rect 15945 5218 15951 5278
rect 15985 5218 15991 5278
rect 15945 5206 15991 5218
rect 16073 5278 16119 5290
rect 16073 5218 16079 5278
rect 16113 5218 16119 5278
rect 16073 5206 16119 5218
rect 16201 5278 16247 5290
rect 16201 5218 16207 5278
rect 16241 5218 16247 5278
rect 16201 5206 16247 5218
rect 16329 5278 16375 5290
rect 16329 5218 16335 5278
rect 16369 5218 16375 5278
rect 16329 5206 16375 5218
rect 16457 5278 16503 5290
rect 16457 5218 16463 5278
rect 16497 5218 16503 5278
rect 16457 5206 16503 5218
rect 16585 5278 16631 5290
rect 16585 5218 16591 5278
rect 16625 5218 16631 5278
rect 16585 5206 16631 5218
rect 16713 5278 16759 5290
rect 16713 5218 16719 5278
rect 16753 5218 16759 5278
rect 16713 5206 16759 5218
rect 16841 5278 16887 5290
rect 16841 5218 16847 5278
rect 16881 5218 16887 5278
rect 16841 5206 16887 5218
rect 16969 5278 17015 5290
rect 16969 5218 16975 5278
rect 17009 5218 17015 5278
rect 16969 5206 17015 5218
rect 17097 5278 17143 5290
rect 17097 5218 17103 5278
rect 17137 5218 17143 5278
rect 17097 5206 17143 5218
rect 17225 5278 17271 5290
rect 17225 5218 17231 5278
rect 17265 5218 17271 5278
rect 17225 5206 17271 5218
rect 17353 5278 17399 5290
rect 17353 5218 17359 5278
rect 17393 5218 17399 5278
rect 17353 5206 17399 5218
rect 17481 5278 17527 5290
rect 17481 5218 17487 5278
rect 17521 5218 17527 5278
rect 17481 5206 17527 5218
rect 17609 5278 17655 5290
rect 17609 5218 17615 5278
rect 17649 5218 17655 5278
rect 17609 5206 17655 5218
rect 17737 5278 17783 5290
rect 17737 5218 17743 5278
rect 17777 5218 17783 5278
rect 17737 5206 17783 5218
rect 17865 5278 17911 5290
rect 17865 5218 17871 5278
rect 17905 5218 17911 5278
rect 17865 5206 17911 5218
rect 17993 5278 18039 5290
rect 17993 5218 17999 5278
rect 18033 5218 18039 5278
rect 17993 5206 18039 5218
rect 18121 5278 18167 5290
rect 18121 5218 18127 5278
rect 18161 5218 18167 5278
rect 18121 5206 18167 5218
rect 18249 5278 18295 5290
rect 18249 5218 18255 5278
rect 18289 5218 18295 5278
rect 18249 5206 18295 5218
rect 18377 5278 18423 5290
rect 18377 5218 18383 5278
rect 18417 5218 18423 5278
rect 18377 5206 18423 5218
rect 18505 5278 18551 5290
rect 18505 5218 18511 5278
rect 18545 5218 18551 5278
rect 18505 5206 18551 5218
rect 18633 5278 18679 5290
rect 18633 5218 18639 5278
rect 18673 5218 18679 5278
rect 18633 5206 18679 5218
rect 18761 5278 18807 5290
rect 18761 5218 18767 5278
rect 18801 5218 18807 5278
rect 18761 5206 18807 5218
rect 18889 5278 18935 5290
rect 18889 5218 18895 5278
rect 18929 5218 18935 5278
rect 18889 5206 18935 5218
rect 19017 5278 19063 5290
rect 19017 5218 19023 5278
rect 19057 5218 19063 5278
rect 19017 5206 19063 5218
rect 19145 5278 19191 5290
rect 19145 5218 19151 5278
rect 19185 5218 19191 5278
rect 19145 5206 19191 5218
rect 19273 5278 19319 5290
rect 19273 5218 19279 5278
rect 19313 5218 19319 5278
rect 19273 5206 19319 5218
rect 19401 5278 19447 5290
rect 19401 5218 19407 5278
rect 19441 5218 19447 5278
rect 19401 5206 19447 5218
rect 19529 5278 19575 5290
rect 19529 5218 19535 5278
rect 19569 5218 19575 5278
rect 19529 5206 19575 5218
rect 19657 5278 19703 5290
rect 19657 5218 19663 5278
rect 19697 5218 19703 5278
rect 19657 5206 19703 5218
rect 19785 5278 19831 5290
rect 19785 5218 19791 5278
rect 19825 5218 19831 5278
rect 19785 5206 19831 5218
rect 19913 5278 19959 5290
rect 29239 5285 29303 5291
rect 29495 5319 37465 5320
rect 29495 5290 29529 5319
rect 29751 5290 29785 5319
rect 30007 5290 30041 5319
rect 30263 5290 30297 5319
rect 30519 5290 30553 5319
rect 30775 5290 30809 5319
rect 31031 5290 31065 5319
rect 31287 5290 31321 5319
rect 31543 5290 31577 5319
rect 31799 5290 31833 5319
rect 32055 5290 32089 5319
rect 32311 5290 32345 5319
rect 32567 5290 32601 5319
rect 32823 5290 32857 5319
rect 33079 5290 33113 5319
rect 33335 5290 33369 5319
rect 33591 5290 33625 5319
rect 33847 5290 33881 5319
rect 34103 5290 34137 5319
rect 34359 5290 34393 5319
rect 34615 5290 34649 5319
rect 34871 5290 34905 5319
rect 35127 5290 35161 5319
rect 35291 5318 35355 5319
rect 35383 5290 35417 5319
rect 35639 5290 35673 5319
rect 35895 5318 35970 5319
rect 35895 5290 35929 5318
rect 36151 5290 36185 5319
rect 36407 5290 36441 5319
rect 36663 5290 36697 5319
rect 36919 5290 36953 5319
rect 37175 5290 37209 5319
rect 37431 5290 37465 5319
rect 37720 5307 37726 5320
rect 37778 5307 37784 5359
rect 37720 5301 37784 5307
rect 19913 5218 19919 5278
rect 19953 5218 19959 5278
rect 19913 5206 19959 5218
rect 29361 5278 29407 5290
rect 29361 5218 29367 5278
rect 29401 5218 29407 5278
rect 29361 5206 29407 5218
rect 29489 5278 29535 5290
rect 29489 5218 29495 5278
rect 29529 5218 29535 5278
rect 29489 5206 29535 5218
rect 29617 5278 29663 5290
rect 29617 5218 29623 5278
rect 29657 5218 29663 5278
rect 29617 5206 29663 5218
rect 29745 5278 29791 5290
rect 29745 5218 29751 5278
rect 29785 5218 29791 5278
rect 29745 5206 29791 5218
rect 29873 5278 29919 5290
rect 29873 5218 29879 5278
rect 29913 5218 29919 5278
rect 29873 5206 29919 5218
rect 30001 5278 30047 5290
rect 30001 5218 30007 5278
rect 30041 5218 30047 5278
rect 30001 5206 30047 5218
rect 30129 5278 30175 5290
rect 30129 5218 30135 5278
rect 30169 5218 30175 5278
rect 30129 5206 30175 5218
rect 30257 5278 30303 5290
rect 30257 5218 30263 5278
rect 30297 5218 30303 5278
rect 30257 5206 30303 5218
rect 30385 5278 30431 5290
rect 30385 5218 30391 5278
rect 30425 5218 30431 5278
rect 30385 5206 30431 5218
rect 30513 5278 30559 5290
rect 30513 5218 30519 5278
rect 30553 5218 30559 5278
rect 30513 5206 30559 5218
rect 30641 5278 30687 5290
rect 30641 5218 30647 5278
rect 30681 5218 30687 5278
rect 30641 5206 30687 5218
rect 30769 5278 30815 5290
rect 30769 5218 30775 5278
rect 30809 5218 30815 5278
rect 30769 5206 30815 5218
rect 30897 5278 30943 5290
rect 30897 5218 30903 5278
rect 30937 5218 30943 5278
rect 30897 5206 30943 5218
rect 31025 5278 31071 5290
rect 31025 5218 31031 5278
rect 31065 5218 31071 5278
rect 31025 5206 31071 5218
rect 31153 5278 31199 5290
rect 31153 5218 31159 5278
rect 31193 5218 31199 5278
rect 31153 5206 31199 5218
rect 31281 5278 31327 5290
rect 31281 5218 31287 5278
rect 31321 5218 31327 5278
rect 31281 5206 31327 5218
rect 31409 5278 31455 5290
rect 31409 5218 31415 5278
rect 31449 5218 31455 5278
rect 31409 5206 31455 5218
rect 31537 5278 31583 5290
rect 31537 5218 31543 5278
rect 31577 5218 31583 5278
rect 31537 5206 31583 5218
rect 31665 5278 31711 5290
rect 31665 5218 31671 5278
rect 31705 5218 31711 5278
rect 31665 5206 31711 5218
rect 31793 5278 31839 5290
rect 31793 5218 31799 5278
rect 31833 5218 31839 5278
rect 31793 5206 31839 5218
rect 31921 5278 31967 5290
rect 31921 5218 31927 5278
rect 31961 5218 31967 5278
rect 31921 5206 31967 5218
rect 32049 5278 32095 5290
rect 32049 5218 32055 5278
rect 32089 5218 32095 5278
rect 32049 5206 32095 5218
rect 32177 5278 32223 5290
rect 32177 5218 32183 5278
rect 32217 5218 32223 5278
rect 32177 5206 32223 5218
rect 32305 5278 32351 5290
rect 32305 5218 32311 5278
rect 32345 5218 32351 5278
rect 32305 5206 32351 5218
rect 32433 5278 32479 5290
rect 32433 5218 32439 5278
rect 32473 5218 32479 5278
rect 32433 5206 32479 5218
rect 32561 5278 32607 5290
rect 32561 5218 32567 5278
rect 32601 5218 32607 5278
rect 32561 5206 32607 5218
rect 32689 5278 32735 5290
rect 32689 5218 32695 5278
rect 32729 5218 32735 5278
rect 32689 5206 32735 5218
rect 32817 5278 32863 5290
rect 32817 5218 32823 5278
rect 32857 5218 32863 5278
rect 32817 5206 32863 5218
rect 32945 5278 32991 5290
rect 32945 5218 32951 5278
rect 32985 5218 32991 5278
rect 32945 5206 32991 5218
rect 33073 5278 33119 5290
rect 33073 5218 33079 5278
rect 33113 5218 33119 5278
rect 33073 5206 33119 5218
rect 33201 5278 33247 5290
rect 33201 5218 33207 5278
rect 33241 5218 33247 5278
rect 33201 5206 33247 5218
rect 33329 5278 33375 5290
rect 33329 5218 33335 5278
rect 33369 5218 33375 5278
rect 33329 5206 33375 5218
rect 33457 5278 33503 5290
rect 33457 5218 33463 5278
rect 33497 5218 33503 5278
rect 33457 5206 33503 5218
rect 33585 5278 33631 5290
rect 33585 5218 33591 5278
rect 33625 5218 33631 5278
rect 33585 5206 33631 5218
rect 33713 5278 33759 5290
rect 33713 5218 33719 5278
rect 33753 5218 33759 5278
rect 33713 5206 33759 5218
rect 33841 5278 33887 5290
rect 33841 5218 33847 5278
rect 33881 5218 33887 5278
rect 33841 5206 33887 5218
rect 33969 5278 34015 5290
rect 33969 5218 33975 5278
rect 34009 5218 34015 5278
rect 33969 5206 34015 5218
rect 34097 5278 34143 5290
rect 34097 5218 34103 5278
rect 34137 5218 34143 5278
rect 34097 5206 34143 5218
rect 34225 5278 34271 5290
rect 34225 5218 34231 5278
rect 34265 5218 34271 5278
rect 34225 5206 34271 5218
rect 34353 5278 34399 5290
rect 34353 5218 34359 5278
rect 34393 5218 34399 5278
rect 34353 5206 34399 5218
rect 34481 5278 34527 5290
rect 34481 5218 34487 5278
rect 34521 5218 34527 5278
rect 34481 5206 34527 5218
rect 34609 5278 34655 5290
rect 34609 5218 34615 5278
rect 34649 5218 34655 5278
rect 34609 5206 34655 5218
rect 34737 5278 34783 5290
rect 34737 5218 34743 5278
rect 34777 5218 34783 5278
rect 34737 5206 34783 5218
rect 34865 5278 34911 5290
rect 34865 5218 34871 5278
rect 34905 5218 34911 5278
rect 34865 5206 34911 5218
rect 34993 5278 35039 5290
rect 34993 5218 34999 5278
rect 35033 5218 35039 5278
rect 34993 5206 35039 5218
rect 35121 5278 35167 5290
rect 35121 5218 35127 5278
rect 35161 5218 35167 5278
rect 35121 5206 35167 5218
rect 35249 5278 35295 5290
rect 35249 5218 35255 5278
rect 35289 5218 35295 5278
rect 35249 5206 35295 5218
rect 35377 5278 35423 5290
rect 35377 5218 35383 5278
rect 35417 5218 35423 5278
rect 35377 5206 35423 5218
rect 35505 5278 35551 5290
rect 35505 5218 35511 5278
rect 35545 5218 35551 5278
rect 35505 5206 35551 5218
rect 35633 5278 35679 5290
rect 35633 5218 35639 5278
rect 35673 5218 35679 5278
rect 35633 5206 35679 5218
rect 35761 5278 35807 5290
rect 35761 5218 35767 5278
rect 35801 5218 35807 5278
rect 35761 5206 35807 5218
rect 35889 5278 35935 5290
rect 35889 5218 35895 5278
rect 35929 5218 35935 5278
rect 35889 5206 35935 5218
rect 36017 5278 36063 5290
rect 36017 5218 36023 5278
rect 36057 5218 36063 5278
rect 36017 5206 36063 5218
rect 36145 5278 36191 5290
rect 36145 5218 36151 5278
rect 36185 5218 36191 5278
rect 36145 5206 36191 5218
rect 36273 5278 36319 5290
rect 36273 5218 36279 5278
rect 36313 5218 36319 5278
rect 36273 5206 36319 5218
rect 36401 5278 36447 5290
rect 36401 5218 36407 5278
rect 36441 5218 36447 5278
rect 36401 5206 36447 5218
rect 36529 5278 36575 5290
rect 36529 5218 36535 5278
rect 36569 5218 36575 5278
rect 36529 5206 36575 5218
rect 36657 5278 36703 5290
rect 36657 5218 36663 5278
rect 36697 5218 36703 5278
rect 36657 5206 36703 5218
rect 36785 5278 36831 5290
rect 36785 5218 36791 5278
rect 36825 5218 36831 5278
rect 36785 5206 36831 5218
rect 36913 5278 36959 5290
rect 36913 5218 36919 5278
rect 36953 5218 36959 5278
rect 36913 5206 36959 5218
rect 37041 5278 37087 5290
rect 37041 5218 37047 5278
rect 37081 5218 37087 5278
rect 37041 5206 37087 5218
rect 37169 5278 37215 5290
rect 37169 5218 37175 5278
rect 37209 5218 37215 5278
rect 37169 5206 37215 5218
rect 37297 5278 37343 5290
rect 37297 5218 37303 5278
rect 37337 5218 37343 5278
rect 37297 5206 37343 5218
rect 37425 5278 37471 5290
rect 37425 5218 37431 5278
rect 37465 5218 37471 5278
rect 37425 5206 37471 5218
rect 37553 5278 37599 5290
rect 37553 5218 37559 5278
rect 37593 5218 37599 5278
rect 37553 5206 37599 5218
rect -317 5154 -283 5206
rect 611 5154 645 5206
rect 867 5154 901 5206
rect 1875 5154 1909 5206
rect 2131 5154 2165 5206
rect 2387 5154 2421 5206
rect 3494 5154 3528 5206
rect 3750 5154 3784 5206
rect 4006 5154 4040 5206
rect 4262 5154 4296 5206
rect 4518 5154 4552 5206
rect 8059 5154 8093 5206
rect 8315 5154 8349 5206
rect 8571 5154 8605 5206
rect 8827 5154 8861 5206
rect 9083 5154 9117 5206
rect 9339 5154 9373 5206
rect 9595 5154 9629 5206
rect 9851 5154 9885 5206
rect 10107 5154 10141 5206
rect 15823 5154 15857 5206
rect 16079 5154 16113 5206
rect 16335 5154 16369 5206
rect 16591 5154 16625 5206
rect 16847 5154 16881 5206
rect 17103 5154 17137 5206
rect 17359 5154 17393 5206
rect 17615 5154 17649 5206
rect 17871 5154 17905 5206
rect 18127 5154 18161 5206
rect 18383 5154 18417 5206
rect 18639 5154 18673 5206
rect 18895 5154 18929 5206
rect 19151 5154 19185 5206
rect 19407 5154 19441 5206
rect 19663 5154 19697 5206
rect 19919 5154 19953 5206
rect 29367 5154 29401 5206
rect 29623 5154 29657 5206
rect 29879 5154 29913 5206
rect 30135 5154 30169 5206
rect 30391 5154 30425 5206
rect 30647 5154 30681 5206
rect 30903 5154 30937 5206
rect 31159 5154 31193 5206
rect 31415 5154 31449 5206
rect 31671 5154 31705 5206
rect 31927 5154 31961 5206
rect 32183 5154 32217 5206
rect 32439 5154 32473 5206
rect 32695 5154 32729 5206
rect 32951 5154 32985 5206
rect 33207 5154 33241 5206
rect 33463 5154 33497 5206
rect 33719 5154 33753 5206
rect 33975 5154 34009 5206
rect 34231 5154 34265 5206
rect 34487 5154 34521 5206
rect 34743 5154 34777 5206
rect 34999 5154 35033 5206
rect 35255 5154 35289 5206
rect 35511 5154 35545 5206
rect 35767 5154 35801 5206
rect 36023 5154 36057 5206
rect 36279 5154 36313 5206
rect 36535 5154 36569 5206
rect 36791 5154 36825 5206
rect 37047 5154 37081 5206
rect 37303 5154 37337 5206
rect 37559 5154 37593 5206
rect 38407 5158 38471 5164
rect 38407 5154 38413 5158
rect -363 5148 38413 5154
rect -363 5110 -319 5148
rect -281 5110 -191 5148
rect -153 5110 609 5148
rect 647 5110 737 5148
rect 775 5110 865 5148
rect 903 5110 1873 5148
rect 1911 5110 2001 5148
rect 2039 5110 2129 5148
rect 2167 5110 2257 5148
rect 2295 5110 2385 5148
rect 2423 5110 3492 5148
rect 3530 5110 3620 5148
rect 3658 5110 3748 5148
rect 3786 5110 3876 5148
rect 3914 5110 4004 5148
rect 4042 5110 4132 5148
rect 4170 5110 4260 5148
rect 4298 5110 4388 5148
rect 4426 5110 4516 5148
rect 4554 5110 8057 5148
rect 8095 5110 8185 5148
rect 8223 5110 8313 5148
rect 8351 5110 8441 5148
rect 8479 5110 8569 5148
rect 8607 5110 8697 5148
rect 8735 5110 8825 5148
rect 8863 5110 8953 5148
rect 8991 5110 9081 5148
rect 9119 5110 9209 5148
rect 9247 5110 9337 5148
rect 9375 5110 9465 5148
rect 9503 5110 9593 5148
rect 9631 5110 9721 5148
rect 9759 5110 9849 5148
rect 9887 5110 9977 5148
rect 10015 5110 10105 5148
rect 10143 5110 15821 5148
rect 15859 5110 15949 5148
rect 15987 5110 16077 5148
rect 16115 5110 16205 5148
rect 16243 5110 16333 5148
rect 16371 5110 16461 5148
rect 16499 5110 16589 5148
rect 16627 5110 16717 5148
rect 16755 5110 16845 5148
rect 16883 5110 16973 5148
rect 17011 5110 17101 5148
rect 17139 5110 17229 5148
rect 17267 5110 17357 5148
rect 17395 5110 17485 5148
rect 17523 5110 17613 5148
rect 17651 5110 17741 5148
rect 17779 5110 17869 5148
rect 17907 5110 17997 5148
rect 18035 5110 18125 5148
rect 18163 5110 18253 5148
rect 18291 5110 18381 5148
rect 18419 5110 18509 5148
rect 18547 5110 18637 5148
rect 18675 5110 18765 5148
rect 18803 5110 18893 5148
rect 18931 5110 19021 5148
rect 19059 5110 19149 5148
rect 19187 5110 19277 5148
rect 19315 5110 19405 5148
rect 19443 5110 19533 5148
rect 19571 5110 19661 5148
rect 19699 5110 19789 5148
rect 19827 5110 19917 5148
rect 19955 5110 29365 5148
rect 29403 5110 29493 5148
rect 29531 5110 29621 5148
rect 29659 5110 29749 5148
rect 29787 5110 29877 5148
rect 29915 5110 30005 5148
rect 30043 5110 30133 5148
rect 30171 5110 30261 5148
rect 30299 5110 30389 5148
rect 30427 5110 30517 5148
rect 30555 5110 30645 5148
rect 30683 5110 30773 5148
rect 30811 5110 30901 5148
rect 30939 5110 31029 5148
rect 31067 5110 31157 5148
rect 31195 5110 31285 5148
rect 31323 5110 31413 5148
rect 31451 5110 31541 5148
rect 31579 5110 31669 5148
rect 31707 5110 31797 5148
rect 31835 5110 31925 5148
rect 31963 5110 32053 5148
rect 32091 5110 32181 5148
rect 32219 5110 32309 5148
rect 32347 5110 32437 5148
rect 32475 5110 32565 5148
rect 32603 5110 32693 5148
rect 32731 5110 32821 5148
rect 32859 5110 32949 5148
rect 32987 5110 33077 5148
rect 33115 5110 33205 5148
rect 33243 5110 33333 5148
rect 33371 5110 33461 5148
rect 33499 5110 33589 5148
rect 33627 5110 33717 5148
rect 33755 5110 33845 5148
rect 33883 5110 33973 5148
rect 34011 5110 34101 5148
rect 34139 5110 34229 5148
rect 34267 5110 34357 5148
rect 34395 5110 34485 5148
rect 34523 5110 34613 5148
rect 34651 5110 34741 5148
rect 34779 5110 34869 5148
rect 34907 5110 34997 5148
rect 35035 5110 35125 5148
rect 35163 5110 35253 5148
rect 35291 5110 35381 5148
rect 35419 5110 35509 5148
rect 35547 5110 35637 5148
rect 35675 5110 35765 5148
rect 35803 5110 35893 5148
rect 35931 5110 36021 5148
rect 36059 5110 36149 5148
rect 36187 5110 36277 5148
rect 36315 5110 36405 5148
rect 36443 5110 36533 5148
rect 36571 5110 36661 5148
rect 36699 5110 36789 5148
rect 36827 5110 36917 5148
rect 36955 5110 37045 5148
rect 37083 5110 37173 5148
rect 37211 5110 37301 5148
rect 37339 5110 37429 5148
rect 37467 5110 37557 5148
rect 37595 5110 38413 5148
rect -363 5106 38413 5110
rect 38465 5106 38471 5158
rect -363 5104 38471 5106
rect 38407 5102 38471 5104
rect 150 4070 210 4078
rect 150 4018 154 4070
rect 206 4018 210 4070
rect 150 4007 210 4018
rect 162 3998 196 4007
rect 5102 3925 5169 3929
rect 5102 3873 5108 3925
rect 5160 3915 5169 3925
rect 5160 3881 5175 3915
rect 5160 3873 5169 3881
rect 5102 3869 5169 3873
rect 358 3085 418 3091
rect 358 3033 362 3085
rect 414 3033 418 3085
rect 358 3024 418 3033
rect 370 3013 404 3024
rect 358 2914 418 2920
rect 358 2862 362 2914
rect 414 2862 418 2914
rect 358 2853 418 2862
rect 1270 2914 1330 2920
rect 1270 2862 1274 2914
rect 1326 2862 1330 2914
rect 1270 2853 1330 2862
rect 1876 2913 1936 2919
rect 1876 2861 1880 2913
rect 1932 2861 1936 2913
rect 370 2842 404 2853
rect 1282 2842 1316 2853
rect 1876 2852 1936 2861
rect 2804 2912 2864 2918
rect 2804 2860 2808 2912
rect 2860 2860 2864 2912
rect 1888 2841 1922 2852
rect 2804 2849 2864 2860
rect 4016 2914 4076 2920
rect 4016 2862 4020 2914
rect 4072 2862 4076 2914
rect 4016 2853 4076 2862
rect 5352 2907 5418 2918
rect 5352 2855 5358 2907
rect 5410 2855 5418 2907
rect 2816 2840 2850 2849
rect 4028 2842 4062 2853
rect 5352 2844 5418 2855
rect 5959 2905 6023 2911
rect 5959 2853 5965 2905
rect 6017 2853 6023 2905
rect 5959 2847 6023 2853
rect 6565 2905 6629 2911
rect 6565 2853 6571 2905
rect 6623 2853 6629 2905
rect 6565 2847 6629 2853
rect 7171 2905 7235 2911
rect 7171 2853 7177 2905
rect 7229 2853 7235 2905
rect 7171 2847 7235 2853
rect 7777 2905 7841 2911
rect 7777 2853 7783 2905
rect 7835 2853 7841 2905
rect 7777 2847 7841 2853
rect 10327 2910 10391 2921
rect 10327 2858 10332 2910
rect 10384 2858 10391 2910
rect 10327 2847 10391 2858
rect 10932 2901 10998 2912
rect 10932 2849 10938 2901
rect 10990 2849 10998 2901
rect 5367 2840 5401 2844
rect 5973 2839 6007 2847
rect 6579 2839 6613 2847
rect 7185 2839 7219 2847
rect 7791 2839 7825 2847
rect 10341 2843 10375 2847
rect 10932 2838 10998 2849
rect 11538 2902 11604 2913
rect 11538 2850 11544 2902
rect 11596 2850 11604 2902
rect 11538 2839 11604 2850
rect 12144 2901 12210 2912
rect 12144 2849 12150 2901
rect 12202 2849 12210 2901
rect 12144 2838 12210 2849
rect 12750 2901 12816 2912
rect 12750 2849 12756 2901
rect 12808 2849 12816 2901
rect 12750 2838 12816 2849
rect 13356 2903 13422 2914
rect 13356 2851 13362 2903
rect 13414 2851 13422 2903
rect 13356 2840 13422 2851
rect 13962 2903 14028 2914
rect 13962 2851 13968 2903
rect 14020 2851 14028 2903
rect 13962 2840 14028 2851
rect 14568 2902 14634 2913
rect 14568 2850 14574 2902
rect 14626 2850 14634 2902
rect 14568 2839 14634 2850
rect 20149 2902 20213 2908
rect 20149 2850 20155 2902
rect 20207 2850 20213 2902
rect 20149 2844 20213 2850
rect 20755 2902 20819 2908
rect 20755 2850 20761 2902
rect 20813 2850 20819 2902
rect 20755 2844 20819 2850
rect 21361 2903 21425 2909
rect 21361 2851 21367 2903
rect 21419 2851 21425 2903
rect 21361 2845 21425 2851
rect 21967 2902 22031 2908
rect 21967 2850 21973 2902
rect 22025 2850 22031 2902
rect 20163 2839 20197 2844
rect 20769 2839 20803 2844
rect 21375 2840 21409 2845
rect 21967 2844 22031 2850
rect 22573 2902 22637 2908
rect 22573 2850 22579 2902
rect 22631 2850 22637 2902
rect 22573 2844 22637 2850
rect 23179 2902 23243 2908
rect 23179 2850 23185 2902
rect 23237 2850 23243 2902
rect 23179 2844 23243 2850
rect 23785 2902 23849 2908
rect 23785 2850 23791 2902
rect 23843 2850 23849 2902
rect 23785 2844 23849 2850
rect 24391 2902 24455 2908
rect 24391 2850 24397 2902
rect 24449 2850 24455 2902
rect 24391 2844 24455 2850
rect 24997 2902 25061 2908
rect 24997 2850 25003 2902
rect 25055 2850 25061 2902
rect 24997 2844 25061 2850
rect 25603 2902 25667 2908
rect 25603 2850 25609 2902
rect 25661 2850 25667 2902
rect 25603 2844 25667 2850
rect 26209 2902 26273 2908
rect 26209 2850 26215 2902
rect 26267 2850 26273 2902
rect 26209 2844 26273 2850
rect 26815 2902 26879 2908
rect 26815 2850 26821 2902
rect 26873 2850 26879 2902
rect 26815 2844 26879 2850
rect 27421 2902 27485 2908
rect 27421 2850 27427 2902
rect 27479 2850 27485 2902
rect 27421 2844 27485 2850
rect 28027 2902 28091 2908
rect 28027 2850 28033 2902
rect 28085 2850 28091 2902
rect 28027 2844 28091 2850
rect 28633 2902 28697 2908
rect 28633 2850 28639 2902
rect 28691 2850 28697 2902
rect 28633 2844 28697 2850
rect 21981 2839 22015 2844
rect 22587 2839 22621 2844
rect 23193 2839 23227 2844
rect 23799 2839 23833 2844
rect 24405 2839 24439 2844
rect 25011 2839 25045 2844
rect 25617 2839 25651 2844
rect 26223 2839 26257 2844
rect 26829 2839 26863 2844
rect 27435 2839 27469 2844
rect 28041 2839 28075 2844
rect 28647 2839 28681 2844
rect -93 1954 -33 1960
rect -93 1902 -89 1954
rect -37 1902 -33 1954
rect -93 1896 -33 1902
rect -81 1882 -47 1896
rect 964 1815 1024 1821
rect 964 1763 968 1815
rect 1020 1763 1024 1815
rect 964 1754 1024 1763
rect 1876 1814 1936 1820
rect 1876 1762 1880 1814
rect 1932 1762 1936 1814
rect 976 1743 1010 1754
rect 1876 1753 1936 1762
rect 2482 1815 2542 1821
rect 2482 1763 2486 1815
rect 2538 1763 2542 1815
rect 7776 1818 7842 1829
rect 2482 1754 2542 1763
rect 3408 1804 3472 1810
rect 1888 1742 1922 1753
rect 2494 1743 2528 1754
rect 3408 1752 3414 1804
rect 3466 1752 3472 1804
rect 3408 1746 3472 1752
rect 4620 1805 4684 1811
rect 4620 1753 4626 1805
rect 4678 1753 4684 1805
rect 4620 1747 4684 1753
rect 5226 1805 5290 1811
rect 5226 1753 5232 1805
rect 5284 1753 5290 1805
rect 7776 1766 7782 1818
rect 7834 1766 7842 1818
rect 7776 1755 7842 1766
rect 8382 1818 8448 1829
rect 8382 1766 8388 1818
rect 8440 1766 8448 1818
rect 8382 1755 8448 1766
rect 8988 1818 9054 1829
rect 8988 1766 8994 1818
rect 9046 1766 9054 1818
rect 8988 1755 9054 1766
rect 9594 1818 9660 1829
rect 15780 1818 15846 1829
rect 9594 1766 9600 1818
rect 9652 1766 9660 1818
rect 9594 1755 9660 1766
rect 10200 1807 10266 1818
rect 10200 1755 10206 1807
rect 10258 1755 10266 1807
rect 15780 1766 15786 1818
rect 15838 1766 15846 1818
rect 15780 1755 15846 1766
rect 16386 1817 16452 1828
rect 16386 1765 16392 1817
rect 16444 1765 16452 1817
rect 5226 1747 5290 1753
rect 3422 1738 3456 1746
rect 4634 1733 4668 1747
rect 5240 1739 5274 1747
rect 10200 1744 10266 1755
rect 16386 1754 16452 1765
rect 16992 1817 17058 1828
rect 16992 1765 16998 1817
rect 17050 1765 17058 1817
rect 16992 1754 17058 1765
rect 17598 1816 17664 1827
rect 17598 1764 17604 1816
rect 17656 1764 17664 1816
rect 17598 1753 17664 1764
rect 18204 1816 18270 1827
rect 18204 1764 18210 1816
rect 18262 1764 18270 1816
rect 18204 1753 18270 1764
rect 18810 1816 18876 1827
rect 18810 1764 18816 1816
rect 18868 1764 18876 1816
rect 18810 1753 18876 1764
rect 19416 1815 19482 1826
rect 19416 1763 19422 1815
rect 19474 1763 19482 1815
rect 19416 1752 19482 1763
rect 20023 1815 20087 1821
rect 20023 1763 20029 1815
rect 20081 1763 20087 1815
rect 20023 1757 20087 1763
rect 29239 1814 29303 1820
rect 29239 1762 29245 1814
rect 29297 1762 29303 1814
rect 20037 1752 20071 1757
rect 29239 1756 29303 1762
rect 29845 1814 29909 1820
rect 29845 1762 29851 1814
rect 29903 1762 29909 1814
rect 29845 1756 29909 1762
rect 30451 1813 30515 1819
rect 30451 1761 30457 1813
rect 30509 1761 30515 1813
rect 29253 1751 29287 1756
rect 29859 1751 29893 1756
rect 30451 1755 30515 1761
rect 31057 1814 31121 1820
rect 31057 1762 31063 1814
rect 31115 1762 31121 1814
rect 31057 1756 31121 1762
rect 31663 1814 31727 1820
rect 31663 1762 31669 1814
rect 31721 1762 31727 1814
rect 31663 1756 31727 1762
rect 32269 1814 32333 1820
rect 32269 1762 32275 1814
rect 32327 1762 32333 1814
rect 32269 1756 32333 1762
rect 32875 1814 32939 1820
rect 32875 1762 32881 1814
rect 32933 1762 32939 1814
rect 32875 1756 32939 1762
rect 33481 1814 33545 1820
rect 33481 1762 33487 1814
rect 33539 1762 33545 1814
rect 33481 1756 33545 1762
rect 34087 1814 34151 1820
rect 34087 1762 34093 1814
rect 34145 1762 34151 1814
rect 34087 1756 34151 1762
rect 34693 1814 34757 1820
rect 34693 1762 34699 1814
rect 34751 1762 34757 1814
rect 34693 1756 34757 1762
rect 35299 1814 35363 1820
rect 35299 1762 35305 1814
rect 35357 1762 35363 1814
rect 35299 1756 35363 1762
rect 35905 1813 35969 1819
rect 35905 1761 35911 1813
rect 35963 1761 35969 1813
rect 30465 1750 30499 1755
rect 31071 1751 31105 1756
rect 31677 1751 31711 1756
rect 32283 1751 32317 1756
rect 32889 1751 32923 1756
rect 33495 1751 33529 1756
rect 34101 1751 34135 1756
rect 34707 1751 34741 1756
rect 35313 1751 35347 1756
rect 35905 1755 35969 1761
rect 36511 1814 36575 1820
rect 36511 1762 36517 1814
rect 36569 1762 36575 1814
rect 36511 1756 36575 1762
rect 37117 1814 37181 1820
rect 37117 1762 37123 1814
rect 37175 1762 37181 1814
rect 37117 1756 37181 1762
rect 37723 1814 37787 1820
rect 37723 1762 37729 1814
rect 37781 1762 37787 1814
rect 37723 1756 37787 1762
rect 35919 1750 35953 1755
rect 36525 1751 36559 1756
rect 37131 1751 37165 1756
rect 37737 1751 37771 1756
rect 10215 1735 10249 1744
rect 964 1669 1024 1675
rect 964 1617 968 1669
rect 1020 1617 1024 1669
rect 964 1608 1024 1617
rect 976 1597 1010 1608
<< via1 >>
rect 38413 6256 38465 6308
rect -298 6082 -238 6088
rect -298 6039 -290 6082
rect -290 6039 -245 6082
rect -245 6039 -238 6082
rect -298 6031 -238 6039
rect -89 6031 -37 6083
rect 363 6014 415 6066
rect 752 6082 812 6088
rect 752 6039 760 6082
rect 760 6039 805 6082
rect 805 6039 812 6082
rect 752 6031 812 6039
rect 1274 6057 1326 6109
rect 1880 6042 1932 6094
rect 1972 6071 2032 6077
rect 1972 6028 1980 6071
rect 1980 6028 2025 6071
rect 2025 6028 2032 6071
rect 1972 6020 2032 6028
rect 2809 6060 2861 6112
rect 4110 6161 4170 6167
rect 4110 6118 4118 6161
rect 4118 6118 4163 6161
rect 4163 6118 4170 6161
rect 4110 6110 4170 6118
rect 4021 6030 4073 6082
rect 5049 6023 5101 6075
rect 5359 6058 5411 6110
rect 7687 6158 7747 6164
rect 7687 6115 7695 6158
rect 7695 6115 7740 6158
rect 7740 6115 7747 6158
rect 7687 6107 7747 6115
rect 5966 6042 6018 6094
rect 6571 6042 6623 6094
rect 7177 6041 7229 6093
rect 7783 6018 7835 6070
rect 10332 6055 10384 6107
rect 10938 6042 10990 6094
rect 11544 6041 11596 6093
rect 12178 6041 12230 6093
rect 12756 6041 12808 6093
rect 13362 6035 13414 6087
rect 13968 6035 14020 6087
rect 14570 6041 14622 6093
rect 14702 6086 14762 6092
rect 14702 6043 14710 6086
rect 14710 6043 14755 6086
rect 14755 6043 14762 6086
rect 14702 6035 14762 6043
rect 20155 6045 20207 6097
rect 20762 6040 20814 6092
rect 21367 6040 21419 6092
rect 21974 6041 22026 6093
rect 22580 6041 22632 6093
rect 23186 6042 23238 6094
rect 23798 6041 23850 6093
rect 25003 6041 25055 6093
rect 25609 6041 25661 6093
rect 26197 6040 26249 6092
rect 26822 6041 26874 6093
rect 27429 6041 27481 6093
rect 28034 6042 28086 6094
rect 28638 6041 28690 6093
rect 28730 6107 28790 6115
rect 28730 6064 28737 6107
rect 28737 6064 28782 6107
rect 28782 6064 28790 6107
rect 28730 6058 28790 6064
rect 37704 5768 37756 5820
rect 38689 5684 38741 5736
rect 37704 5597 37756 5649
rect -385 5376 -325 5382
rect -385 5333 -377 5376
rect -377 5333 -332 5376
rect -332 5333 -325 5376
rect -385 5325 -325 5333
rect -89 5311 -37 5363
rect 964 5439 1024 5445
rect 964 5396 972 5439
rect 972 5396 1017 5439
rect 1017 5396 1024 5439
rect 964 5388 1024 5396
rect 968 5296 1020 5348
rect 1756 5306 1808 5358
rect 2493 5439 2553 5445
rect 2493 5396 2501 5439
rect 2501 5396 2546 5439
rect 2546 5396 2553 5439
rect 2493 5388 2553 5396
rect 2486 5296 2538 5348
rect 3414 5319 3466 5371
rect 4664 5448 4724 5454
rect 4664 5405 4672 5448
rect 4672 5405 4717 5448
rect 4717 5405 4724 5448
rect 4664 5397 4724 5405
rect 7922 5433 7982 5439
rect 7922 5390 7930 5433
rect 7930 5390 7975 5433
rect 7975 5390 7982 5433
rect 7922 5382 7982 5390
rect 4626 5290 4678 5342
rect 7929 5289 7981 5341
rect 8387 5326 8439 5378
rect 8993 5325 9045 5377
rect 9599 5325 9651 5377
rect 10206 5310 10258 5362
rect 15691 5402 15751 5408
rect 15691 5359 15699 5402
rect 15699 5359 15744 5402
rect 15744 5359 15751 5402
rect 15691 5351 15751 5359
rect 15792 5324 15844 5376
rect 16408 5324 16460 5376
rect 20029 5306 20081 5358
rect 29245 5291 29297 5343
rect 29852 5326 29904 5378
rect 30461 5325 30513 5377
rect 31063 5325 31115 5377
rect 31669 5325 31721 5377
rect 32275 5325 32327 5377
rect 32891 5325 32943 5377
rect 33487 5325 33539 5377
rect 34093 5325 34145 5377
rect 34700 5325 34752 5377
rect 35297 5324 35349 5376
rect 35912 5324 35964 5376
rect 36518 5325 36570 5377
rect 37124 5325 37176 5377
rect 37726 5307 37778 5359
rect 38413 5106 38465 5158
rect 154 4018 206 4070
rect 5108 3873 5160 3925
rect 362 3033 414 3085
rect 362 2862 414 2914
rect 1274 2862 1326 2914
rect 1880 2861 1932 2913
rect 2808 2860 2860 2912
rect 4020 2862 4072 2914
rect 5358 2855 5410 2907
rect 5965 2853 6017 2905
rect 6571 2853 6623 2905
rect 7177 2853 7229 2905
rect 7783 2853 7835 2905
rect 10332 2858 10384 2910
rect 10938 2849 10990 2901
rect 11544 2850 11596 2902
rect 12150 2849 12202 2901
rect 12756 2849 12808 2901
rect 13362 2851 13414 2903
rect 13968 2851 14020 2903
rect 14574 2850 14626 2902
rect 20155 2850 20207 2902
rect 20761 2850 20813 2902
rect 21367 2851 21419 2903
rect 21973 2850 22025 2902
rect 22579 2850 22631 2902
rect 23185 2850 23237 2902
rect 23791 2850 23843 2902
rect 24397 2850 24449 2902
rect 25003 2850 25055 2902
rect 25609 2850 25661 2902
rect 26215 2850 26267 2902
rect 26821 2850 26873 2902
rect 27427 2850 27479 2902
rect 28033 2850 28085 2902
rect 28639 2850 28691 2902
rect -89 1902 -37 1954
rect 968 1763 1020 1815
rect 1880 1762 1932 1814
rect 2486 1763 2538 1815
rect 3414 1752 3466 1804
rect 4626 1753 4678 1805
rect 5232 1753 5284 1805
rect 7782 1766 7834 1818
rect 8388 1766 8440 1818
rect 8994 1766 9046 1818
rect 9600 1766 9652 1818
rect 10206 1755 10258 1807
rect 15786 1766 15838 1818
rect 16392 1765 16444 1817
rect 16998 1765 17050 1817
rect 17604 1764 17656 1816
rect 18210 1764 18262 1816
rect 18816 1764 18868 1816
rect 19422 1763 19474 1815
rect 20029 1763 20081 1815
rect 29245 1762 29297 1814
rect 29851 1762 29903 1814
rect 30457 1761 30509 1813
rect 31063 1762 31115 1814
rect 31669 1762 31721 1814
rect 32275 1762 32327 1814
rect 32881 1762 32933 1814
rect 33487 1762 33539 1814
rect 34093 1762 34145 1814
rect 34699 1762 34751 1814
rect 35305 1762 35357 1814
rect 35911 1761 35963 1813
rect 36517 1762 36569 1814
rect 37123 1762 37175 1814
rect 37729 1762 37781 1814
rect 968 1617 1020 1669
<< metal2 >>
rect 38407 6308 38471 6314
rect 38407 6256 38413 6308
rect 38465 6256 38471 6308
rect -95 6198 210 6254
rect 38407 6250 38471 6256
rect -304 6088 -238 6094
rect -304 6031 -298 6088
rect -304 6026 -238 6031
rect -95 6083 -31 6198
rect -95 6031 -89 6083
rect -37 6031 -31 6083
rect -95 6025 -31 6031
rect -391 5382 -380 5388
rect -332 5382 -319 5388
rect -391 5325 -385 5382
rect -325 5325 -319 5382
rect -391 5319 -319 5325
rect -95 5363 -31 5369
rect -95 5311 -89 5363
rect -37 5311 -31 5363
rect -95 5305 -31 5311
rect -93 1960 -31 5305
rect 150 4072 210 6198
rect 4104 6167 4116 6173
rect 4164 6167 4176 6173
rect 1268 6109 1332 6115
rect 746 6088 758 6094
rect 806 6088 818 6094
rect 357 6066 421 6072
rect 357 6014 363 6066
rect 415 6014 421 6066
rect 746 6031 752 6088
rect 812 6031 818 6088
rect 1268 6057 1274 6109
rect 1326 6057 1332 6109
rect 2803 6112 2867 6118
rect 1268 6051 1332 6057
rect 1874 6094 1938 6100
rect 746 6025 818 6031
rect 357 6008 421 6014
rect 150 4016 152 4072
rect 208 4016 210 4072
rect 150 4007 210 4016
rect 363 3096 414 6008
rect 958 5445 970 5451
rect 1018 5445 1030 5451
rect 958 5388 964 5445
rect 1024 5388 1030 5445
rect 958 5382 1030 5388
rect 962 5348 1026 5354
rect 962 5296 968 5348
rect 1020 5296 1026 5348
rect 962 5290 1026 5296
rect 358 3087 418 3096
rect 358 3031 360 3087
rect 416 3031 418 3087
rect 358 3022 418 3031
rect 363 2925 414 3022
rect 358 2916 418 2925
rect 358 2860 360 2916
rect 416 2860 418 2916
rect 358 2851 418 2860
rect -93 1956 -33 1960
rect -93 1900 -91 1956
rect -35 1900 -33 1956
rect -93 1891 -33 1900
rect 968 1826 1024 5290
rect 1274 2925 1326 6051
rect 1874 6042 1880 6094
rect 1932 6042 1938 6094
rect 1874 6036 1938 6042
rect 1966 6077 1978 6083
rect 2026 6077 2038 6083
rect 1750 5358 1814 5364
rect 1750 5306 1756 5358
rect 1808 5306 1814 5358
rect 1750 5300 1814 5306
rect 1270 2916 1330 2925
rect 1270 2860 1272 2916
rect 1328 2860 1330 2916
rect 1270 2851 1330 2860
rect 964 1817 1024 1826
rect 964 1761 966 1817
rect 1022 1761 1024 1817
rect 1756 1814 1808 5300
rect 1880 2924 1932 6036
rect 1966 6020 1972 6077
rect 2032 6020 2038 6077
rect 2803 6060 2809 6112
rect 2861 6060 2867 6112
rect 4104 6110 4110 6167
rect 4170 6110 4176 6167
rect 7681 6164 7694 6170
rect 7742 6164 7753 6170
rect 4104 6104 4176 6110
rect 5353 6110 5417 6116
rect 2803 6054 2867 6060
rect 4015 6082 4079 6088
rect 1966 6014 2038 6020
rect 2487 5445 2500 5451
rect 2548 5445 2559 5451
rect 2487 5388 2493 5445
rect 2553 5388 2559 5445
rect 2487 5382 2559 5388
rect 2480 5348 2544 5354
rect 2480 5296 2486 5348
rect 2538 5296 2544 5348
rect 2480 5290 2544 5296
rect 1876 2915 1936 2924
rect 1876 2859 1878 2915
rect 1934 2859 1936 2915
rect 1876 2850 1936 2859
rect 1889 1825 1923 1829
rect 2486 1826 2538 5290
rect 2808 2923 2861 6054
rect 4015 6030 4021 6082
rect 4073 6030 4079 6082
rect 4015 6024 4079 6030
rect 5043 6076 5107 6081
rect 5043 6075 5160 6076
rect 3408 5371 3472 5377
rect 3408 5319 3414 5371
rect 3466 5319 3472 5371
rect 3408 5313 3472 5319
rect 2804 2914 2864 2923
rect 2804 2858 2806 2914
rect 2862 2858 2864 2914
rect 2804 2849 2864 2858
rect 1876 1816 1936 1825
rect 1876 1814 1878 1816
rect 1756 1762 1878 1814
rect 964 1752 1024 1761
rect 968 1680 1024 1752
rect 1876 1760 1878 1762
rect 1934 1760 1936 1816
rect 1876 1751 1936 1760
rect 2482 1817 2542 1826
rect 2482 1761 2484 1817
rect 2540 1761 2542 1817
rect 3414 1815 3466 5313
rect 4020 2925 4073 6024
rect 5043 6023 5049 6075
rect 5101 6023 5160 6075
rect 5353 6058 5359 6110
rect 5411 6058 5417 6110
rect 7681 6107 7687 6164
rect 7747 6107 7753 6164
rect 28724 6115 28796 6121
rect 7681 6101 7753 6107
rect 10326 6107 10390 6113
rect 5353 6052 5417 6058
rect 5960 6094 6024 6100
rect 5043 6017 5160 6023
rect 4658 5454 4671 5460
rect 4719 5454 4730 5460
rect 4658 5397 4664 5454
rect 4724 5397 4730 5454
rect 4658 5391 4730 5397
rect 4620 5342 4684 5348
rect 4620 5290 4626 5342
rect 4678 5290 4684 5342
rect 4620 5284 4684 5290
rect 4016 2916 4076 2925
rect 4016 2860 4018 2916
rect 4074 2860 4076 2916
rect 4016 2851 4076 2860
rect 4626 2017 4678 5284
rect 5108 3929 5160 6017
rect 5097 3927 5171 3929
rect 5097 3926 5106 3927
rect 5094 3873 5106 3926
rect 5097 3871 5106 3873
rect 5162 3871 5171 3927
rect 5097 3869 5171 3871
rect 5358 2918 5411 6052
rect 5960 6042 5966 6094
rect 6018 6042 6024 6094
rect 5960 6036 6024 6042
rect 6565 6094 6629 6100
rect 6565 6042 6571 6094
rect 6623 6042 6629 6094
rect 6565 6036 6629 6042
rect 7171 6093 7235 6099
rect 7171 6041 7177 6093
rect 7229 6041 7235 6093
rect 5352 2909 5418 2918
rect 5965 2916 6018 6036
rect 6571 2916 6624 6036
rect 7171 6035 7235 6041
rect 7777 6070 7841 6076
rect 7177 2916 7230 6035
rect 7777 6018 7783 6070
rect 7835 6018 7841 6070
rect 10326 6055 10332 6107
rect 10384 6055 10390 6107
rect 10326 6049 10390 6055
rect 10932 6094 10996 6100
rect 7777 6012 7841 6018
rect 7783 2916 7836 6012
rect 7916 5439 7918 5445
rect 7966 5439 7988 5445
rect 7916 5382 7922 5439
rect 7982 5382 7988 5439
rect 7916 5376 7988 5382
rect 8381 5378 8445 5384
rect 7923 5341 7987 5347
rect 7923 5289 7929 5341
rect 7981 5289 7987 5341
rect 8381 5326 8387 5378
rect 8439 5326 8445 5378
rect 8381 5320 8445 5326
rect 8987 5377 9051 5383
rect 8987 5325 8993 5377
rect 9045 5325 9051 5377
rect 7923 5283 7987 5289
rect 5352 2853 5357 2909
rect 5413 2853 5418 2909
rect 5352 2844 5418 2853
rect 5959 2907 6023 2916
rect 5959 2851 5963 2907
rect 6019 2851 6023 2907
rect 5959 2842 6023 2851
rect 6565 2907 6629 2916
rect 6565 2851 6569 2907
rect 6625 2851 6629 2907
rect 6565 2842 6629 2851
rect 7171 2907 7235 2916
rect 7171 2851 7175 2907
rect 7231 2851 7235 2907
rect 7171 2842 7235 2851
rect 7777 2907 7841 2916
rect 7777 2851 7781 2907
rect 7837 2851 7841 2907
rect 7777 2842 7841 2851
rect 4626 1965 5284 2017
rect 4626 1816 4678 1965
rect 5232 1816 5284 1965
rect 7776 1820 7842 1829
rect 2482 1752 2542 1761
rect 3408 1806 3472 1815
rect 3408 1750 3412 1806
rect 3468 1750 3472 1806
rect 3408 1741 3472 1750
rect 4620 1807 4684 1816
rect 4620 1751 4624 1807
rect 4680 1751 4684 1807
rect 4620 1742 4684 1751
rect 5226 1807 5290 1816
rect 5226 1751 5230 1807
rect 5286 1751 5290 1807
rect 7776 1764 7781 1820
rect 7837 1818 7842 1820
rect 7930 1818 7982 5283
rect 8388 1829 8440 5320
rect 8987 5319 9051 5325
rect 9593 5377 9657 5383
rect 9593 5325 9599 5377
rect 9651 5325 9657 5377
rect 9593 5319 9657 5325
rect 10200 5362 10264 5368
rect 8994 1829 9046 5319
rect 9600 1829 9652 5319
rect 10200 5310 10206 5362
rect 10258 5310 10264 5362
rect 10200 5304 10264 5310
rect 7837 1766 7982 1818
rect 8382 1820 8448 1829
rect 7837 1764 7842 1766
rect 7776 1755 7842 1764
rect 8382 1764 8387 1820
rect 8443 1764 8448 1820
rect 8382 1755 8448 1764
rect 8988 1820 9054 1829
rect 8988 1764 8993 1820
rect 9049 1764 9054 1820
rect 8988 1755 9054 1764
rect 9594 1820 9660 1829
rect 9594 1764 9599 1820
rect 9655 1764 9660 1820
rect 10206 1818 10258 5304
rect 10332 2921 10384 6049
rect 10932 6042 10938 6094
rect 10990 6042 10996 6094
rect 10932 6036 10996 6042
rect 11538 6093 11602 6099
rect 11538 6041 11544 6093
rect 11596 6041 11602 6093
rect 10327 2912 10391 2921
rect 10938 2912 10990 6036
rect 11538 6035 11602 6041
rect 12150 6093 12236 6099
rect 12150 6041 12178 6093
rect 12230 6041 12236 6093
rect 12150 6035 12236 6041
rect 12750 6093 12814 6099
rect 14564 6093 14628 6099
rect 12750 6041 12756 6093
rect 12808 6041 12814 6093
rect 12750 6035 12814 6041
rect 13356 6087 13420 6093
rect 13356 6035 13362 6087
rect 13414 6035 13420 6087
rect 11544 2913 11596 6035
rect 10327 2856 10331 2912
rect 10387 2856 10391 2912
rect 10327 2847 10391 2856
rect 10932 2903 10998 2912
rect 10932 2847 10937 2903
rect 10993 2847 10998 2903
rect 10932 2838 10998 2847
rect 11538 2904 11604 2913
rect 12150 2912 12202 6035
rect 12756 2912 12808 6035
rect 13356 6029 13420 6035
rect 13962 6087 14026 6093
rect 13962 6035 13968 6087
rect 14020 6035 14026 6087
rect 14564 6041 14570 6093
rect 14622 6041 14628 6093
rect 14564 6035 14628 6041
rect 14696 6092 14709 6098
rect 14757 6092 14768 6098
rect 14696 6035 14702 6092
rect 14762 6035 14768 6092
rect 20149 6097 20213 6103
rect 20149 6045 20155 6097
rect 20207 6045 20213 6097
rect 20149 6039 20213 6045
rect 20756 6092 20820 6098
rect 20756 6040 20762 6092
rect 20814 6040 20820 6092
rect 13962 6029 14026 6035
rect 13362 2914 13414 6029
rect 13968 2914 14020 6029
rect 11538 2848 11543 2904
rect 11599 2848 11604 2904
rect 11538 2839 11604 2848
rect 12144 2903 12210 2912
rect 12144 2847 12149 2903
rect 12205 2847 12210 2903
rect 12144 2838 12210 2847
rect 12750 2903 12816 2912
rect 12750 2847 12755 2903
rect 12811 2847 12816 2903
rect 12750 2838 12816 2847
rect 13356 2905 13422 2914
rect 13356 2849 13361 2905
rect 13417 2849 13422 2905
rect 13356 2840 13422 2849
rect 13962 2905 14028 2914
rect 14574 2913 14626 6035
rect 14696 6029 14768 6035
rect 15685 5408 15697 5414
rect 15745 5408 15757 5414
rect 15685 5351 15691 5408
rect 15751 5351 15757 5408
rect 15685 5345 15757 5351
rect 15786 5376 15850 5382
rect 15786 5324 15792 5376
rect 15844 5324 15850 5376
rect 16402 5376 16466 5382
rect 16402 5325 16408 5376
rect 15786 5318 15850 5324
rect 16392 5324 16408 5325
rect 16460 5324 16466 5376
rect 16392 5318 16466 5324
rect 20023 5358 20087 5364
rect 13962 2849 13967 2905
rect 14023 2849 14028 2905
rect 13962 2840 14028 2849
rect 14568 2904 14634 2913
rect 14568 2848 14573 2904
rect 14629 2848 14634 2904
rect 14568 2839 14634 2848
rect 15786 1829 15838 5318
rect 15780 1820 15846 1829
rect 16392 1828 16444 5318
rect 20023 5306 20029 5358
rect 20081 5306 20087 5358
rect 16998 1828 17050 5306
rect 9594 1755 9660 1764
rect 10200 1809 10266 1818
rect 5226 1742 5290 1751
rect 10200 1753 10205 1809
rect 10261 1753 10266 1809
rect 15780 1764 15785 1820
rect 15841 1764 15846 1820
rect 15780 1755 15846 1764
rect 16386 1819 16452 1828
rect 16386 1763 16391 1819
rect 16447 1763 16452 1819
rect 16386 1754 16452 1763
rect 16992 1819 17058 1828
rect 17604 1827 17656 5305
rect 18210 1827 18262 5305
rect 18816 1827 18868 5305
rect 16992 1763 16997 1819
rect 17053 1763 17058 1819
rect 16992 1754 17058 1763
rect 17598 1818 17664 1827
rect 17598 1762 17603 1818
rect 17659 1762 17664 1818
rect 17598 1753 17664 1762
rect 18204 1818 18270 1827
rect 18204 1762 18209 1818
rect 18265 1762 18270 1818
rect 18204 1753 18270 1762
rect 18810 1818 18876 1827
rect 19422 1826 19474 5304
rect 20023 5300 20087 5306
rect 20029 1826 20081 5300
rect 20155 2913 20208 6039
rect 20756 6034 20820 6040
rect 21361 6092 21425 6098
rect 21361 6040 21367 6092
rect 21419 6040 21425 6092
rect 21361 6034 21425 6040
rect 21968 6093 22032 6099
rect 21968 6041 21974 6093
rect 22026 6041 22032 6093
rect 21968 6035 22032 6041
rect 22574 6093 22638 6099
rect 22574 6041 22580 6093
rect 22632 6041 22638 6093
rect 22574 6035 22638 6041
rect 23180 6094 23244 6100
rect 23180 6042 23186 6094
rect 23238 6042 23244 6094
rect 23792 6093 23856 6099
rect 23792 6062 23798 6093
rect 23180 6036 23244 6042
rect 23791 6041 23798 6062
rect 23850 6041 23856 6093
rect 20761 2913 20814 6034
rect 21367 2914 21420 6034
rect 20149 2904 20213 2913
rect 20149 2848 20153 2904
rect 20209 2848 20213 2904
rect 20149 2839 20213 2848
rect 20755 2904 20819 2913
rect 20755 2848 20759 2904
rect 20815 2848 20819 2904
rect 20755 2839 20819 2848
rect 21361 2905 21425 2914
rect 21973 2913 22026 6035
rect 22579 2913 22632 6035
rect 23185 2913 23238 6036
rect 23791 6035 23856 6041
rect 24997 6093 25061 6099
rect 24997 6041 25003 6093
rect 25055 6041 25061 6093
rect 23791 6034 23850 6035
rect 23791 2913 23844 6034
rect 24397 2913 24450 6039
rect 24997 6035 25061 6041
rect 25603 6093 25667 6099
rect 25603 6041 25609 6093
rect 25661 6041 25667 6093
rect 25603 6035 25667 6041
rect 26191 6092 26268 6098
rect 26191 6040 26197 6092
rect 26249 6040 26268 6092
rect 25003 2913 25056 6035
rect 25609 2913 25662 6035
rect 26191 6034 26268 6040
rect 26816 6093 26880 6099
rect 26816 6041 26822 6093
rect 26874 6041 26880 6093
rect 26816 6035 26880 6041
rect 27423 6093 27487 6099
rect 27423 6041 27429 6093
rect 27481 6041 27487 6093
rect 27423 6035 27487 6041
rect 28028 6094 28092 6100
rect 28028 6042 28034 6094
rect 28086 6042 28092 6094
rect 28028 6036 28092 6042
rect 28632 6093 28696 6099
rect 28632 6041 28638 6093
rect 28690 6041 28696 6093
rect 28724 6058 28730 6115
rect 28790 6058 28796 6115
rect 28724 6052 28796 6058
rect 38413 6078 38465 6250
rect 38520 6078 38595 6080
rect 38413 6071 38595 6078
rect 26215 2913 26268 6034
rect 26821 2913 26874 6035
rect 27427 2913 27480 6035
rect 28033 2913 28086 6036
rect 28632 6035 28696 6041
rect 28638 2913 28691 6035
rect 38413 6015 38529 6071
rect 38585 6015 38595 6071
rect 38413 6008 38595 6015
rect 37698 5820 37762 5826
rect 37698 5768 37704 5820
rect 37756 5768 37762 5820
rect 37698 5762 37762 5768
rect 37713 5734 37747 5762
rect 37806 5744 37915 5753
rect 37806 5734 37849 5744
rect 37713 5688 37849 5734
rect 37905 5688 37915 5744
rect 37713 5683 37915 5688
rect 37713 5655 37747 5683
rect 37806 5679 37915 5683
rect 37698 5649 37762 5655
rect 37698 5597 37704 5649
rect 37756 5597 37762 5649
rect 37698 5591 37762 5597
rect 29846 5378 29910 5384
rect 29239 5343 29303 5349
rect 29239 5291 29245 5343
rect 29297 5291 29303 5343
rect 29846 5326 29852 5378
rect 29904 5326 29910 5378
rect 29846 5320 29910 5326
rect 30455 5377 30519 5383
rect 30455 5325 30461 5377
rect 30513 5325 30519 5377
rect 29239 5285 29303 5291
rect 21361 2849 21365 2905
rect 21421 2849 21425 2905
rect 21361 2840 21425 2849
rect 21967 2904 22031 2913
rect 21967 2848 21971 2904
rect 22027 2848 22031 2904
rect 21967 2839 22031 2848
rect 22573 2904 22637 2913
rect 22573 2848 22577 2904
rect 22633 2848 22637 2904
rect 22573 2839 22637 2848
rect 23179 2904 23243 2913
rect 23179 2848 23183 2904
rect 23239 2848 23243 2904
rect 23179 2839 23243 2848
rect 23785 2904 23849 2913
rect 23785 2848 23789 2904
rect 23845 2848 23849 2904
rect 23785 2839 23849 2848
rect 24391 2904 24455 2913
rect 24391 2848 24395 2904
rect 24451 2848 24455 2904
rect 24391 2839 24455 2848
rect 24997 2904 25061 2913
rect 24997 2848 25001 2904
rect 25057 2848 25061 2904
rect 24997 2839 25061 2848
rect 25603 2904 25667 2913
rect 25603 2848 25607 2904
rect 25663 2848 25667 2904
rect 25603 2839 25667 2848
rect 26209 2904 26273 2913
rect 26209 2848 26213 2904
rect 26269 2848 26273 2904
rect 26209 2839 26273 2848
rect 26815 2904 26879 2913
rect 26815 2848 26819 2904
rect 26875 2848 26879 2904
rect 26815 2839 26879 2848
rect 27421 2904 27485 2913
rect 27421 2848 27425 2904
rect 27481 2848 27485 2904
rect 27421 2839 27485 2848
rect 28027 2904 28091 2913
rect 28027 2848 28031 2904
rect 28087 2848 28091 2904
rect 28027 2839 28091 2848
rect 28633 2904 28697 2913
rect 28633 2848 28637 2904
rect 28693 2848 28697 2904
rect 28633 2839 28697 2848
rect 18810 1762 18815 1818
rect 18871 1762 18876 1818
rect 18810 1753 18876 1762
rect 19416 1817 19482 1826
rect 19416 1761 19421 1817
rect 19477 1761 19482 1817
rect 10200 1744 10266 1753
rect 19416 1752 19482 1761
rect 20023 1817 20087 1826
rect 29245 1825 29297 5285
rect 29851 1825 29903 5320
rect 30455 5319 30519 5325
rect 31057 5377 31121 5383
rect 31057 5325 31063 5377
rect 31115 5325 31121 5377
rect 31057 5319 31121 5325
rect 31663 5377 31727 5383
rect 31663 5325 31669 5377
rect 31721 5325 31727 5377
rect 31663 5319 31727 5325
rect 32269 5377 32333 5383
rect 32269 5325 32275 5377
rect 32327 5325 32333 5377
rect 32269 5319 32333 5325
rect 32885 5377 32949 5383
rect 32885 5325 32891 5377
rect 32943 5325 32949 5377
rect 32885 5320 32949 5325
rect 32881 5319 32949 5320
rect 33481 5377 33545 5383
rect 33481 5325 33487 5377
rect 33539 5325 33545 5377
rect 33481 5319 33545 5325
rect 34087 5377 34151 5383
rect 34087 5325 34093 5377
rect 34145 5325 34151 5377
rect 34087 5319 34151 5325
rect 34694 5377 34758 5383
rect 34694 5325 34700 5377
rect 34752 5325 34758 5377
rect 34694 5319 34758 5325
rect 35291 5376 35355 5382
rect 35291 5324 35297 5376
rect 35349 5324 35355 5376
rect 35291 5320 35355 5324
rect 35906 5376 35970 5382
rect 35906 5324 35912 5376
rect 35964 5324 35970 5376
rect 20023 1761 20027 1817
rect 20083 1761 20087 1817
rect 20023 1752 20087 1761
rect 29239 1816 29303 1825
rect 29239 1760 29243 1816
rect 29299 1760 29303 1816
rect 29239 1751 29303 1760
rect 29845 1816 29909 1825
rect 30457 1824 30509 5319
rect 31063 1825 31115 5319
rect 31669 1825 31721 5319
rect 32275 1825 32327 5319
rect 32881 1825 32933 5319
rect 33487 1825 33539 5319
rect 34093 1825 34145 5319
rect 34699 1825 34751 5319
rect 35291 5318 35357 5320
rect 35906 5318 35970 5324
rect 36512 5377 36576 5383
rect 36512 5325 36518 5377
rect 36570 5325 36576 5377
rect 36512 5319 36576 5325
rect 37118 5377 37182 5383
rect 37118 5325 37124 5377
rect 37176 5325 37182 5377
rect 37118 5319 37182 5325
rect 37720 5359 37784 5365
rect 35305 1825 35357 5318
rect 29845 1760 29849 1816
rect 29905 1760 29909 1816
rect 29845 1751 29909 1760
rect 30451 1815 30515 1824
rect 30451 1759 30455 1815
rect 30511 1759 30515 1815
rect 30451 1750 30515 1759
rect 31057 1816 31121 1825
rect 31057 1760 31061 1816
rect 31117 1760 31121 1816
rect 31057 1751 31121 1760
rect 31663 1816 31727 1825
rect 31663 1760 31667 1816
rect 31723 1760 31727 1816
rect 31663 1751 31727 1760
rect 32269 1816 32333 1825
rect 32269 1760 32273 1816
rect 32329 1760 32333 1816
rect 32269 1751 32333 1760
rect 32875 1816 32939 1825
rect 32875 1760 32879 1816
rect 32935 1760 32939 1816
rect 32875 1751 32939 1760
rect 33481 1816 33545 1825
rect 33481 1760 33485 1816
rect 33541 1760 33545 1816
rect 33481 1751 33545 1760
rect 34087 1816 34151 1825
rect 34087 1760 34091 1816
rect 34147 1760 34151 1816
rect 34087 1751 34151 1760
rect 34693 1816 34757 1825
rect 34693 1760 34697 1816
rect 34753 1760 34757 1816
rect 34693 1751 34757 1760
rect 35299 1816 35363 1825
rect 35911 1824 35963 5318
rect 36517 1825 36569 5319
rect 37123 1825 37175 5319
rect 37720 5307 37726 5359
rect 37778 5307 37784 5359
rect 37720 5301 37784 5307
rect 37729 1825 37781 5301
rect 38413 5164 38465 6008
rect 38520 6006 38595 6008
rect 39085 5745 39160 5747
rect 39081 5744 39160 5745
rect 38683 5738 39160 5744
rect 38683 5736 39094 5738
rect 38683 5684 38689 5736
rect 38741 5684 39094 5736
rect 38683 5682 39094 5684
rect 39150 5682 39160 5738
rect 38683 5676 39160 5682
rect 39081 5675 39160 5676
rect 39085 5673 39160 5675
rect 38407 5158 38471 5164
rect 38407 5106 38413 5158
rect 38465 5106 38471 5158
rect 38407 5102 38471 5106
rect 35299 1760 35303 1816
rect 35359 1760 35363 1816
rect 35299 1751 35363 1760
rect 35905 1815 35969 1824
rect 35905 1759 35909 1815
rect 35965 1759 35969 1815
rect 35905 1750 35969 1759
rect 36511 1816 36575 1825
rect 36511 1760 36515 1816
rect 36571 1760 36575 1816
rect 36511 1751 36575 1760
rect 37117 1816 37181 1825
rect 37117 1760 37121 1816
rect 37177 1760 37181 1816
rect 37117 1751 37181 1760
rect 37723 1816 37787 1825
rect 37723 1760 37727 1816
rect 37783 1760 37787 1816
rect 37723 1751 37787 1760
rect 964 1671 1024 1680
rect 964 1615 966 1671
rect 1022 1615 1024 1671
rect 964 1606 1024 1615
<< via2 >>
rect 152 4070 208 4072
rect 152 4018 154 4070
rect 154 4018 206 4070
rect 206 4018 208 4070
rect 152 4016 208 4018
rect 360 3085 416 3087
rect 360 3033 362 3085
rect 362 3033 414 3085
rect 414 3033 416 3085
rect 360 3031 416 3033
rect 360 2914 416 2916
rect 360 2862 362 2914
rect 362 2862 414 2914
rect 414 2862 416 2914
rect 360 2860 416 2862
rect -91 1954 -35 1956
rect -91 1902 -89 1954
rect -89 1902 -37 1954
rect -37 1902 -35 1954
rect -91 1900 -35 1902
rect 1272 2914 1328 2916
rect 1272 2862 1274 2914
rect 1274 2862 1326 2914
rect 1326 2862 1328 2914
rect 1272 2860 1328 2862
rect 966 1815 1022 1817
rect 966 1763 968 1815
rect 968 1763 1020 1815
rect 1020 1763 1022 1815
rect 966 1761 1022 1763
rect 1878 2913 1934 2915
rect 1878 2861 1880 2913
rect 1880 2861 1932 2913
rect 1932 2861 1934 2913
rect 1878 2859 1934 2861
rect 2806 2912 2862 2914
rect 2806 2860 2808 2912
rect 2808 2860 2860 2912
rect 2860 2860 2862 2912
rect 2806 2858 2862 2860
rect 1878 1814 1934 1816
rect 1878 1762 1880 1814
rect 1880 1762 1932 1814
rect 1932 1762 1934 1814
rect 1878 1760 1934 1762
rect 2484 1815 2540 1817
rect 2484 1763 2486 1815
rect 2486 1763 2538 1815
rect 2538 1763 2540 1815
rect 2484 1761 2540 1763
rect 4018 2914 4074 2916
rect 4018 2862 4020 2914
rect 4020 2862 4072 2914
rect 4072 2862 4074 2914
rect 4018 2860 4074 2862
rect 5106 3925 5162 3927
rect 5106 3873 5108 3925
rect 5108 3873 5160 3925
rect 5160 3873 5162 3925
rect 5106 3871 5162 3873
rect 5357 2907 5413 2909
rect 5357 2855 5358 2907
rect 5358 2855 5410 2907
rect 5410 2855 5413 2907
rect 5357 2853 5413 2855
rect 5963 2905 6019 2907
rect 5963 2853 5965 2905
rect 5965 2853 6017 2905
rect 6017 2853 6019 2905
rect 5963 2851 6019 2853
rect 6569 2905 6625 2907
rect 6569 2853 6571 2905
rect 6571 2853 6623 2905
rect 6623 2853 6625 2905
rect 6569 2851 6625 2853
rect 7175 2905 7231 2907
rect 7175 2853 7177 2905
rect 7177 2853 7229 2905
rect 7229 2853 7231 2905
rect 7175 2851 7231 2853
rect 7781 2905 7837 2907
rect 7781 2853 7783 2905
rect 7783 2853 7835 2905
rect 7835 2853 7837 2905
rect 7781 2851 7837 2853
rect 3412 1804 3468 1806
rect 3412 1752 3414 1804
rect 3414 1752 3466 1804
rect 3466 1752 3468 1804
rect 3412 1750 3468 1752
rect 4624 1805 4680 1807
rect 4624 1753 4626 1805
rect 4626 1753 4678 1805
rect 4678 1753 4680 1805
rect 4624 1751 4680 1753
rect 5230 1805 5286 1807
rect 5230 1753 5232 1805
rect 5232 1753 5284 1805
rect 5284 1753 5286 1805
rect 5230 1751 5286 1753
rect 7781 1818 7837 1820
rect 7781 1766 7782 1818
rect 7782 1766 7834 1818
rect 7834 1766 7837 1818
rect 7781 1764 7837 1766
rect 8387 1818 8443 1820
rect 8387 1766 8388 1818
rect 8388 1766 8440 1818
rect 8440 1766 8443 1818
rect 8387 1764 8443 1766
rect 8993 1818 9049 1820
rect 8993 1766 8994 1818
rect 8994 1766 9046 1818
rect 9046 1766 9049 1818
rect 8993 1764 9049 1766
rect 9599 1818 9655 1820
rect 9599 1766 9600 1818
rect 9600 1766 9652 1818
rect 9652 1766 9655 1818
rect 9599 1764 9655 1766
rect 10331 2910 10387 2912
rect 10331 2858 10332 2910
rect 10332 2858 10384 2910
rect 10384 2858 10387 2910
rect 10331 2856 10387 2858
rect 10937 2901 10993 2903
rect 10937 2849 10938 2901
rect 10938 2849 10990 2901
rect 10990 2849 10993 2901
rect 10937 2847 10993 2849
rect 11543 2902 11599 2904
rect 11543 2850 11544 2902
rect 11544 2850 11596 2902
rect 11596 2850 11599 2902
rect 11543 2848 11599 2850
rect 12149 2901 12205 2903
rect 12149 2849 12150 2901
rect 12150 2849 12202 2901
rect 12202 2849 12205 2901
rect 12149 2847 12205 2849
rect 12755 2901 12811 2903
rect 12755 2849 12756 2901
rect 12756 2849 12808 2901
rect 12808 2849 12811 2901
rect 12755 2847 12811 2849
rect 13361 2903 13417 2905
rect 13361 2851 13362 2903
rect 13362 2851 13414 2903
rect 13414 2851 13417 2903
rect 13361 2849 13417 2851
rect 13967 2903 14023 2905
rect 13967 2851 13968 2903
rect 13968 2851 14020 2903
rect 14020 2851 14023 2903
rect 13967 2849 14023 2851
rect 14573 2902 14629 2904
rect 14573 2850 14574 2902
rect 14574 2850 14626 2902
rect 14626 2850 14629 2902
rect 14573 2848 14629 2850
rect 10205 1807 10261 1809
rect 10205 1755 10206 1807
rect 10206 1755 10258 1807
rect 10258 1755 10261 1807
rect 10205 1753 10261 1755
rect 15785 1818 15841 1820
rect 15785 1766 15786 1818
rect 15786 1766 15838 1818
rect 15838 1766 15841 1818
rect 15785 1764 15841 1766
rect 16391 1817 16447 1819
rect 16391 1765 16392 1817
rect 16392 1765 16444 1817
rect 16444 1765 16447 1817
rect 16391 1763 16447 1765
rect 16997 1817 17053 1819
rect 16997 1765 16998 1817
rect 16998 1765 17050 1817
rect 17050 1765 17053 1817
rect 16997 1763 17053 1765
rect 17603 1816 17659 1818
rect 17603 1764 17604 1816
rect 17604 1764 17656 1816
rect 17656 1764 17659 1816
rect 17603 1762 17659 1764
rect 18209 1816 18265 1818
rect 18209 1764 18210 1816
rect 18210 1764 18262 1816
rect 18262 1764 18265 1816
rect 18209 1762 18265 1764
rect 20153 2902 20209 2904
rect 20153 2850 20155 2902
rect 20155 2850 20207 2902
rect 20207 2850 20209 2902
rect 20153 2848 20209 2850
rect 20759 2902 20815 2904
rect 20759 2850 20761 2902
rect 20761 2850 20813 2902
rect 20813 2850 20815 2902
rect 20759 2848 20815 2850
rect 38529 6015 38585 6071
rect 37849 5688 37905 5744
rect 21365 2903 21421 2905
rect 21365 2851 21367 2903
rect 21367 2851 21419 2903
rect 21419 2851 21421 2903
rect 21365 2849 21421 2851
rect 21971 2902 22027 2904
rect 21971 2850 21973 2902
rect 21973 2850 22025 2902
rect 22025 2850 22027 2902
rect 21971 2848 22027 2850
rect 22577 2902 22633 2904
rect 22577 2850 22579 2902
rect 22579 2850 22631 2902
rect 22631 2850 22633 2902
rect 22577 2848 22633 2850
rect 23183 2902 23239 2904
rect 23183 2850 23185 2902
rect 23185 2850 23237 2902
rect 23237 2850 23239 2902
rect 23183 2848 23239 2850
rect 23789 2902 23845 2904
rect 23789 2850 23791 2902
rect 23791 2850 23843 2902
rect 23843 2850 23845 2902
rect 23789 2848 23845 2850
rect 24395 2902 24451 2904
rect 24395 2850 24397 2902
rect 24397 2850 24449 2902
rect 24449 2850 24451 2902
rect 24395 2848 24451 2850
rect 25001 2902 25057 2904
rect 25001 2850 25003 2902
rect 25003 2850 25055 2902
rect 25055 2850 25057 2902
rect 25001 2848 25057 2850
rect 25607 2902 25663 2904
rect 25607 2850 25609 2902
rect 25609 2850 25661 2902
rect 25661 2850 25663 2902
rect 25607 2848 25663 2850
rect 26213 2902 26269 2904
rect 26213 2850 26215 2902
rect 26215 2850 26267 2902
rect 26267 2850 26269 2902
rect 26213 2848 26269 2850
rect 26819 2902 26875 2904
rect 26819 2850 26821 2902
rect 26821 2850 26873 2902
rect 26873 2850 26875 2902
rect 26819 2848 26875 2850
rect 27425 2902 27481 2904
rect 27425 2850 27427 2902
rect 27427 2850 27479 2902
rect 27479 2850 27481 2902
rect 27425 2848 27481 2850
rect 28031 2902 28087 2904
rect 28031 2850 28033 2902
rect 28033 2850 28085 2902
rect 28085 2850 28087 2902
rect 28031 2848 28087 2850
rect 28637 2902 28693 2904
rect 28637 2850 28639 2902
rect 28639 2850 28691 2902
rect 28691 2850 28693 2902
rect 28637 2848 28693 2850
rect 18815 1816 18871 1818
rect 18815 1764 18816 1816
rect 18816 1764 18868 1816
rect 18868 1764 18871 1816
rect 18815 1762 18871 1764
rect 19421 1815 19477 1817
rect 19421 1763 19422 1815
rect 19422 1763 19474 1815
rect 19474 1763 19477 1815
rect 19421 1761 19477 1763
rect 20027 1815 20083 1817
rect 20027 1763 20029 1815
rect 20029 1763 20081 1815
rect 20081 1763 20083 1815
rect 20027 1761 20083 1763
rect 29243 1814 29299 1816
rect 29243 1762 29245 1814
rect 29245 1762 29297 1814
rect 29297 1762 29299 1814
rect 29243 1760 29299 1762
rect 29849 1814 29905 1816
rect 29849 1762 29851 1814
rect 29851 1762 29903 1814
rect 29903 1762 29905 1814
rect 29849 1760 29905 1762
rect 30455 1813 30511 1815
rect 30455 1761 30457 1813
rect 30457 1761 30509 1813
rect 30509 1761 30511 1813
rect 30455 1759 30511 1761
rect 31061 1814 31117 1816
rect 31061 1762 31063 1814
rect 31063 1762 31115 1814
rect 31115 1762 31117 1814
rect 31061 1760 31117 1762
rect 31667 1814 31723 1816
rect 31667 1762 31669 1814
rect 31669 1762 31721 1814
rect 31721 1762 31723 1814
rect 31667 1760 31723 1762
rect 32273 1814 32329 1816
rect 32273 1762 32275 1814
rect 32275 1762 32327 1814
rect 32327 1762 32329 1814
rect 32273 1760 32329 1762
rect 32879 1814 32935 1816
rect 32879 1762 32881 1814
rect 32881 1762 32933 1814
rect 32933 1762 32935 1814
rect 32879 1760 32935 1762
rect 33485 1814 33541 1816
rect 33485 1762 33487 1814
rect 33487 1762 33539 1814
rect 33539 1762 33541 1814
rect 33485 1760 33541 1762
rect 34091 1814 34147 1816
rect 34091 1762 34093 1814
rect 34093 1762 34145 1814
rect 34145 1762 34147 1814
rect 34091 1760 34147 1762
rect 34697 1814 34753 1816
rect 34697 1762 34699 1814
rect 34699 1762 34751 1814
rect 34751 1762 34753 1814
rect 34697 1760 34753 1762
rect 39094 5682 39150 5738
rect 35303 1814 35359 1816
rect 35303 1762 35305 1814
rect 35305 1762 35357 1814
rect 35357 1762 35359 1814
rect 35303 1760 35359 1762
rect 35909 1813 35965 1815
rect 35909 1761 35911 1813
rect 35911 1761 35963 1813
rect 35963 1761 35965 1813
rect 35909 1759 35965 1761
rect 36515 1814 36571 1816
rect 36515 1762 36517 1814
rect 36517 1762 36569 1814
rect 36569 1762 36571 1814
rect 36515 1760 36571 1762
rect 37121 1814 37177 1816
rect 37121 1762 37123 1814
rect 37123 1762 37175 1814
rect 37175 1762 37177 1814
rect 37121 1760 37177 1762
rect 37727 1814 37783 1816
rect 37727 1762 37729 1814
rect 37729 1762 37781 1814
rect 37781 1762 37783 1814
rect 37727 1760 37783 1762
rect 966 1669 1022 1671
rect 966 1617 968 1669
rect 968 1617 1020 1669
rect 1020 1617 1022 1669
rect 966 1615 1022 1617
<< metal3 >>
rect 38516 6075 38613 6095
rect 38516 6011 38525 6075
rect 38589 6011 38613 6075
rect 38516 5991 38613 6011
rect 37836 5748 37933 5768
rect 37836 5684 37845 5748
rect 37909 5684 37933 5748
rect 37836 5664 37933 5684
rect 39081 5742 39178 5762
rect 39081 5678 39090 5742
rect 39154 5678 39178 5742
rect 39081 5658 39178 5678
rect -459 5092 213 5094
rect -459 5028 -355 5092
rect -291 5028 -275 5092
rect -211 5028 -195 5092
rect -131 5028 -115 5092
rect -51 5028 -35 5092
rect 29 5028 45 5092
rect 109 5028 213 5092
rect -459 5026 213 5028
rect 355 5092 1027 5094
rect 355 5028 459 5092
rect 523 5028 539 5092
rect 603 5028 619 5092
rect 683 5028 699 5092
rect 763 5028 779 5092
rect 843 5028 859 5092
rect 923 5028 1027 5092
rect 355 5026 1027 5028
rect 1267 5092 2545 5094
rect 1267 5028 1371 5092
rect 1435 5028 1451 5092
rect 1515 5028 1531 5092
rect 1595 5028 1611 5092
rect 1675 5028 1691 5092
rect 1755 5028 1771 5092
rect 1835 5028 1977 5092
rect 2041 5028 2057 5092
rect 2121 5028 2137 5092
rect 2201 5028 2217 5092
rect 2281 5028 2297 5092
rect 2361 5028 2377 5092
rect 2441 5028 2545 5092
rect 1267 5026 2545 5028
rect 2801 5092 5291 5094
rect 2801 5028 2905 5092
rect 2969 5028 2985 5092
rect 3049 5028 3065 5092
rect 3129 5028 3145 5092
rect 3209 5028 3225 5092
rect 3289 5028 3305 5092
rect 3369 5028 3511 5092
rect 3575 5028 3591 5092
rect 3655 5028 3671 5092
rect 3735 5028 3751 5092
rect 3815 5028 3831 5092
rect 3895 5028 3911 5092
rect 3975 5028 4117 5092
rect 4181 5028 4197 5092
rect 4261 5028 4277 5092
rect 4341 5028 4357 5092
rect 4421 5028 4437 5092
rect 4501 5028 4517 5092
rect 4581 5028 4723 5092
rect 4787 5028 4803 5092
rect 4867 5028 4883 5092
rect 4947 5028 4963 5092
rect 5027 5028 5043 5092
rect 5107 5028 5123 5092
rect 5187 5028 5291 5092
rect 2801 5026 5291 5028
rect 5352 5092 10266 5094
rect 5352 5028 5456 5092
rect 5520 5028 5536 5092
rect 5600 5028 5616 5092
rect 5680 5028 5696 5092
rect 5760 5028 5776 5092
rect 5840 5028 5856 5092
rect 5920 5028 6062 5092
rect 6126 5028 6142 5092
rect 6206 5028 6222 5092
rect 6286 5028 6302 5092
rect 6366 5028 6382 5092
rect 6446 5028 6462 5092
rect 6526 5028 6668 5092
rect 6732 5028 6748 5092
rect 6812 5028 6828 5092
rect 6892 5028 6908 5092
rect 6972 5028 6988 5092
rect 7052 5028 7068 5092
rect 7132 5028 7274 5092
rect 7338 5028 7354 5092
rect 7418 5028 7434 5092
rect 7498 5028 7514 5092
rect 7578 5028 7594 5092
rect 7658 5028 7674 5092
rect 7738 5028 7880 5092
rect 7944 5028 7960 5092
rect 8024 5028 8040 5092
rect 8104 5028 8120 5092
rect 8184 5028 8200 5092
rect 8264 5028 8280 5092
rect 8344 5028 8486 5092
rect 8550 5028 8566 5092
rect 8630 5028 8646 5092
rect 8710 5028 8726 5092
rect 8790 5028 8806 5092
rect 8870 5028 8886 5092
rect 8950 5028 9092 5092
rect 9156 5028 9172 5092
rect 9236 5028 9252 5092
rect 9316 5028 9332 5092
rect 9396 5028 9412 5092
rect 9476 5028 9492 5092
rect 9556 5028 9698 5092
rect 9762 5028 9778 5092
rect 9842 5028 9858 5092
rect 9922 5028 9938 5092
rect 10002 5028 10018 5092
rect 10082 5028 10098 5092
rect 10162 5028 10266 5092
rect 5352 5026 10266 5028
rect 10326 5092 20088 5094
rect 10326 5028 10430 5092
rect 10494 5028 10510 5092
rect 10574 5028 10590 5092
rect 10654 5028 10670 5092
rect 10734 5028 10750 5092
rect 10814 5028 10830 5092
rect 10894 5028 11036 5092
rect 11100 5028 11116 5092
rect 11180 5028 11196 5092
rect 11260 5028 11276 5092
rect 11340 5028 11356 5092
rect 11420 5028 11436 5092
rect 11500 5028 11642 5092
rect 11706 5028 11722 5092
rect 11786 5028 11802 5092
rect 11866 5028 11882 5092
rect 11946 5028 11962 5092
rect 12026 5028 12042 5092
rect 12106 5028 12248 5092
rect 12312 5028 12328 5092
rect 12392 5028 12408 5092
rect 12472 5028 12488 5092
rect 12552 5028 12568 5092
rect 12632 5028 12648 5092
rect 12712 5028 12854 5092
rect 12918 5028 12934 5092
rect 12998 5028 13014 5092
rect 13078 5028 13094 5092
rect 13158 5028 13174 5092
rect 13238 5028 13254 5092
rect 13318 5028 13460 5092
rect 13524 5028 13540 5092
rect 13604 5028 13620 5092
rect 13684 5028 13700 5092
rect 13764 5028 13780 5092
rect 13844 5028 13860 5092
rect 13924 5028 14066 5092
rect 14130 5028 14146 5092
rect 14210 5028 14226 5092
rect 14290 5028 14306 5092
rect 14370 5028 14386 5092
rect 14450 5028 14466 5092
rect 14530 5028 14672 5092
rect 14736 5028 14752 5092
rect 14816 5028 14832 5092
rect 14896 5028 14912 5092
rect 14976 5028 14992 5092
rect 15056 5028 15072 5092
rect 15136 5028 15278 5092
rect 15342 5028 15358 5092
rect 15422 5028 15438 5092
rect 15502 5028 15518 5092
rect 15582 5028 15598 5092
rect 15662 5028 15678 5092
rect 15742 5028 15884 5092
rect 15948 5028 15964 5092
rect 16028 5028 16044 5092
rect 16108 5028 16124 5092
rect 16188 5028 16204 5092
rect 16268 5028 16284 5092
rect 16348 5028 16490 5092
rect 16554 5028 16570 5092
rect 16634 5028 16650 5092
rect 16714 5028 16730 5092
rect 16794 5028 16810 5092
rect 16874 5028 16890 5092
rect 16954 5028 17096 5092
rect 17160 5028 17176 5092
rect 17240 5028 17256 5092
rect 17320 5028 17336 5092
rect 17400 5028 17416 5092
rect 17480 5028 17496 5092
rect 17560 5028 17702 5092
rect 17766 5028 17782 5092
rect 17846 5028 17862 5092
rect 17926 5028 17942 5092
rect 18006 5028 18022 5092
rect 18086 5028 18102 5092
rect 18166 5028 18308 5092
rect 18372 5028 18388 5092
rect 18452 5028 18468 5092
rect 18532 5028 18548 5092
rect 18612 5028 18628 5092
rect 18692 5028 18708 5092
rect 18772 5028 18914 5092
rect 18978 5028 18994 5092
rect 19058 5028 19074 5092
rect 19138 5028 19154 5092
rect 19218 5028 19234 5092
rect 19298 5028 19314 5092
rect 19378 5028 19520 5092
rect 19584 5028 19600 5092
rect 19664 5028 19680 5092
rect 19744 5028 19760 5092
rect 19824 5028 19840 5092
rect 19904 5028 19920 5092
rect 19984 5028 20088 5092
rect 10326 5026 20088 5028
rect 20148 5092 39606 5094
rect 20148 5028 20252 5092
rect 20316 5028 20332 5092
rect 20396 5028 20412 5092
rect 20476 5028 20492 5092
rect 20556 5028 20572 5092
rect 20636 5028 20652 5092
rect 20716 5028 20858 5092
rect 20922 5028 20938 5092
rect 21002 5028 21018 5092
rect 21082 5028 21098 5092
rect 21162 5028 21178 5092
rect 21242 5028 21258 5092
rect 21322 5028 21464 5092
rect 21528 5028 21544 5092
rect 21608 5028 21624 5092
rect 21688 5028 21704 5092
rect 21768 5028 21784 5092
rect 21848 5028 21864 5092
rect 21928 5028 22070 5092
rect 22134 5028 22150 5092
rect 22214 5028 22230 5092
rect 22294 5028 22310 5092
rect 22374 5028 22390 5092
rect 22454 5028 22470 5092
rect 22534 5028 22676 5092
rect 22740 5028 22756 5092
rect 22820 5028 22836 5092
rect 22900 5028 22916 5092
rect 22980 5028 22996 5092
rect 23060 5028 23076 5092
rect 23140 5028 23282 5092
rect 23346 5028 23362 5092
rect 23426 5028 23442 5092
rect 23506 5028 23522 5092
rect 23586 5028 23602 5092
rect 23666 5028 23682 5092
rect 23746 5028 23888 5092
rect 23952 5028 23968 5092
rect 24032 5028 24048 5092
rect 24112 5028 24128 5092
rect 24192 5028 24208 5092
rect 24272 5028 24288 5092
rect 24352 5028 24494 5092
rect 24558 5028 24574 5092
rect 24638 5028 24654 5092
rect 24718 5028 24734 5092
rect 24798 5028 24814 5092
rect 24878 5028 24894 5092
rect 24958 5028 25100 5092
rect 25164 5028 25180 5092
rect 25244 5028 25260 5092
rect 25324 5028 25340 5092
rect 25404 5028 25420 5092
rect 25484 5028 25500 5092
rect 25564 5028 25706 5092
rect 25770 5028 25786 5092
rect 25850 5028 25866 5092
rect 25930 5028 25946 5092
rect 26010 5028 26026 5092
rect 26090 5028 26106 5092
rect 26170 5028 26312 5092
rect 26376 5028 26392 5092
rect 26456 5028 26472 5092
rect 26536 5028 26552 5092
rect 26616 5028 26632 5092
rect 26696 5028 26712 5092
rect 26776 5028 26918 5092
rect 26982 5028 26998 5092
rect 27062 5028 27078 5092
rect 27142 5028 27158 5092
rect 27222 5028 27238 5092
rect 27302 5028 27318 5092
rect 27382 5028 27524 5092
rect 27588 5028 27604 5092
rect 27668 5028 27684 5092
rect 27748 5028 27764 5092
rect 27828 5028 27844 5092
rect 27908 5028 27924 5092
rect 27988 5028 28130 5092
rect 28194 5028 28210 5092
rect 28274 5028 28290 5092
rect 28354 5028 28370 5092
rect 28434 5028 28450 5092
rect 28514 5028 28530 5092
rect 28594 5028 28736 5092
rect 28800 5028 28816 5092
rect 28880 5028 28896 5092
rect 28960 5028 28976 5092
rect 29040 5028 29056 5092
rect 29120 5028 29136 5092
rect 29200 5028 29342 5092
rect 29406 5028 29422 5092
rect 29486 5028 29502 5092
rect 29566 5028 29582 5092
rect 29646 5028 29662 5092
rect 29726 5028 29742 5092
rect 29806 5028 29948 5092
rect 30012 5028 30028 5092
rect 30092 5028 30108 5092
rect 30172 5028 30188 5092
rect 30252 5028 30268 5092
rect 30332 5028 30348 5092
rect 30412 5028 30554 5092
rect 30618 5028 30634 5092
rect 30698 5028 30714 5092
rect 30778 5028 30794 5092
rect 30858 5028 30874 5092
rect 30938 5028 30954 5092
rect 31018 5028 31160 5092
rect 31224 5028 31240 5092
rect 31304 5028 31320 5092
rect 31384 5028 31400 5092
rect 31464 5028 31480 5092
rect 31544 5028 31560 5092
rect 31624 5028 31766 5092
rect 31830 5028 31846 5092
rect 31910 5028 31926 5092
rect 31990 5028 32006 5092
rect 32070 5028 32086 5092
rect 32150 5028 32166 5092
rect 32230 5028 32372 5092
rect 32436 5028 32452 5092
rect 32516 5028 32532 5092
rect 32596 5028 32612 5092
rect 32676 5028 32692 5092
rect 32756 5028 32772 5092
rect 32836 5028 32978 5092
rect 33042 5028 33058 5092
rect 33122 5028 33138 5092
rect 33202 5028 33218 5092
rect 33282 5028 33298 5092
rect 33362 5028 33378 5092
rect 33442 5028 33584 5092
rect 33648 5028 33664 5092
rect 33728 5028 33744 5092
rect 33808 5028 33824 5092
rect 33888 5028 33904 5092
rect 33968 5028 33984 5092
rect 34048 5028 34190 5092
rect 34254 5028 34270 5092
rect 34334 5028 34350 5092
rect 34414 5028 34430 5092
rect 34494 5028 34510 5092
rect 34574 5028 34590 5092
rect 34654 5028 34796 5092
rect 34860 5028 34876 5092
rect 34940 5028 34956 5092
rect 35020 5028 35036 5092
rect 35100 5028 35116 5092
rect 35180 5028 35196 5092
rect 35260 5028 35402 5092
rect 35466 5028 35482 5092
rect 35546 5028 35562 5092
rect 35626 5028 35642 5092
rect 35706 5028 35722 5092
rect 35786 5028 35802 5092
rect 35866 5028 36008 5092
rect 36072 5028 36088 5092
rect 36152 5028 36168 5092
rect 36232 5028 36248 5092
rect 36312 5028 36328 5092
rect 36392 5028 36408 5092
rect 36472 5028 36614 5092
rect 36678 5028 36694 5092
rect 36758 5028 36774 5092
rect 36838 5028 36854 5092
rect 36918 5028 36934 5092
rect 36998 5028 37014 5092
rect 37078 5028 37220 5092
rect 37284 5028 37300 5092
rect 37364 5028 37380 5092
rect 37444 5028 37460 5092
rect 37524 5028 37540 5092
rect 37604 5028 37620 5092
rect 37684 5028 37826 5092
rect 37890 5028 37906 5092
rect 37970 5028 37986 5092
rect 38050 5028 38066 5092
rect 38130 5028 38146 5092
rect 38210 5028 38226 5092
rect 38290 5028 38432 5092
rect 38496 5028 38512 5092
rect 38576 5028 38592 5092
rect 38656 5028 38672 5092
rect 38736 5028 38752 5092
rect 38816 5028 38832 5092
rect 38896 5028 39038 5092
rect 39102 5028 39118 5092
rect 39182 5028 39198 5092
rect 39262 5028 39278 5092
rect 39342 5028 39358 5092
rect 39422 5028 39438 5092
rect 39502 5028 39606 5092
rect 20148 5026 39606 5028
rect -459 4872 -393 5026
rect -459 4808 -458 4872
rect -394 4808 -393 4872
rect -459 4792 -393 4808
rect -459 4728 -458 4792
rect -394 4728 -393 4792
rect -459 4712 -393 4728
rect -459 4648 -458 4712
rect -394 4648 -393 4712
rect -459 4632 -393 4648
rect -459 4568 -458 4632
rect -394 4568 -393 4632
rect -459 4552 -393 4568
rect -459 4488 -458 4552
rect -394 4488 -393 4552
rect -459 4472 -393 4488
rect -459 4408 -458 4472
rect -394 4408 -393 4472
rect -459 4392 -393 4408
rect -459 4328 -458 4392
rect -394 4328 -393 4392
rect -459 4312 -393 4328
rect -459 4248 -458 4312
rect -394 4248 -393 4312
rect -459 4232 -393 4248
rect -459 4168 -458 4232
rect -394 4168 -393 4232
rect -459 4152 -393 4168
rect -459 4088 -458 4152
rect -394 4088 -393 4152
rect -459 3998 -393 4088
rect -333 3934 -273 4964
rect -213 3994 -153 5026
rect -93 3934 -33 4964
rect 27 3994 87 5026
rect 147 4872 213 5026
rect 147 4808 148 4872
rect 212 4808 213 4872
rect 147 4792 213 4808
rect 147 4728 148 4792
rect 212 4728 213 4792
rect 147 4712 213 4728
rect 147 4648 148 4712
rect 212 4648 213 4712
rect 147 4632 213 4648
rect 147 4568 148 4632
rect 212 4568 213 4632
rect 147 4552 213 4568
rect 147 4488 148 4552
rect 212 4488 213 4552
rect 147 4472 213 4488
rect 147 4408 148 4472
rect 212 4408 213 4472
rect 147 4392 213 4408
rect 147 4328 148 4392
rect 212 4328 213 4392
rect 147 4312 213 4328
rect 147 4248 148 4312
rect 212 4248 213 4312
rect 147 4232 213 4248
rect 147 4168 148 4232
rect 212 4168 213 4232
rect 147 4152 213 4168
rect 147 4088 148 4152
rect 212 4088 213 4152
rect 147 4072 213 4088
rect 147 4016 152 4072
rect 208 4016 213 4072
rect 147 3998 213 4016
rect 355 4872 421 4962
rect 355 4808 356 4872
rect 420 4808 421 4872
rect 355 4792 421 4808
rect 355 4728 356 4792
rect 420 4728 421 4792
rect 355 4712 421 4728
rect 355 4648 356 4712
rect 420 4648 421 4712
rect 355 4632 421 4648
rect 355 4568 356 4632
rect 420 4568 421 4632
rect 355 4552 421 4568
rect 355 4488 356 4552
rect 420 4488 421 4552
rect 355 4472 421 4488
rect 355 4408 356 4472
rect 420 4408 421 4472
rect 355 4392 421 4408
rect 355 4328 356 4392
rect 420 4328 421 4392
rect 355 4312 421 4328
rect 355 4248 356 4312
rect 420 4248 421 4312
rect 355 4232 421 4248
rect 355 4168 356 4232
rect 420 4168 421 4232
rect 355 4152 421 4168
rect 355 4088 356 4152
rect 420 4088 421 4152
rect 355 3934 421 4088
rect 481 3934 541 4966
rect 601 3996 661 5026
rect 721 3934 781 4966
rect 841 3996 901 5026
rect 961 4872 1027 4962
rect 961 4808 962 4872
rect 1026 4808 1027 4872
rect 961 4792 1027 4808
rect 961 4728 962 4792
rect 1026 4728 1027 4792
rect 961 4712 1027 4728
rect 961 4648 962 4712
rect 1026 4648 1027 4712
rect 961 4632 1027 4648
rect 961 4568 962 4632
rect 1026 4568 1027 4632
rect 961 4552 1027 4568
rect 961 4488 962 4552
rect 1026 4488 1027 4552
rect 961 4472 1027 4488
rect 961 4408 962 4472
rect 1026 4408 1027 4472
rect 961 4392 1027 4408
rect 961 4328 962 4392
rect 1026 4328 1027 4392
rect 961 4312 1027 4328
rect 961 4248 962 4312
rect 1026 4248 1027 4312
rect 961 4232 1027 4248
rect 961 4168 962 4232
rect 1026 4168 1027 4232
rect 961 4152 1027 4168
rect 961 4088 962 4152
rect 1026 4088 1027 4152
rect 961 3934 1027 4088
rect -459 3932 213 3934
rect -459 3868 -355 3932
rect -291 3868 -275 3932
rect -211 3868 -195 3932
rect -131 3868 -115 3932
rect -51 3868 -35 3932
rect 29 3868 45 3932
rect 109 3868 213 3932
rect -459 3866 213 3868
rect 355 3932 1027 3934
rect 355 3868 459 3932
rect 523 3868 539 3932
rect 603 3868 619 3932
rect 683 3868 699 3932
rect 763 3868 779 3932
rect 843 3868 859 3932
rect 923 3868 1027 3932
rect 355 3866 1027 3868
rect -459 3712 -393 3802
rect -459 3648 -458 3712
rect -394 3648 -393 3712
rect -459 3632 -393 3648
rect -459 3568 -458 3632
rect -394 3568 -393 3632
rect -459 3552 -393 3568
rect -459 3488 -458 3552
rect -394 3488 -393 3552
rect -459 3472 -393 3488
rect -459 3408 -458 3472
rect -394 3408 -393 3472
rect -459 3392 -393 3408
rect -459 3328 -458 3392
rect -394 3328 -393 3392
rect -459 3312 -393 3328
rect -459 3248 -458 3312
rect -394 3248 -393 3312
rect -459 3232 -393 3248
rect -459 3168 -458 3232
rect -394 3168 -393 3232
rect -459 3152 -393 3168
rect -459 3088 -458 3152
rect -394 3088 -393 3152
rect -459 3072 -393 3088
rect -459 3008 -458 3072
rect -394 3008 -393 3072
rect -459 2992 -393 3008
rect -459 2928 -458 2992
rect -394 2928 -393 2992
rect -459 2774 -393 2928
rect -333 2774 -273 3806
rect -213 2836 -153 3866
rect -93 2774 -33 3806
rect 27 2836 87 3866
rect 147 3712 213 3802
rect 147 3648 148 3712
rect 212 3648 213 3712
rect 147 3632 213 3648
rect 147 3568 148 3632
rect 212 3568 213 3632
rect 147 3552 213 3568
rect 147 3488 148 3552
rect 212 3488 213 3552
rect 147 3472 213 3488
rect 147 3408 148 3472
rect 212 3408 213 3472
rect 147 3392 213 3408
rect 147 3328 148 3392
rect 212 3328 213 3392
rect 147 3312 213 3328
rect 147 3248 148 3312
rect 212 3248 213 3312
rect 147 3232 213 3248
rect 147 3168 148 3232
rect 212 3168 213 3232
rect 147 3152 213 3168
rect 147 3088 148 3152
rect 212 3088 213 3152
rect 147 3072 213 3088
rect 147 3008 148 3072
rect 212 3008 213 3072
rect 147 2992 213 3008
rect 147 2928 148 2992
rect 212 2928 213 2992
rect 147 2774 213 2928
rect 355 3712 421 3866
rect 355 3648 356 3712
rect 420 3648 421 3712
rect 355 3632 421 3648
rect 355 3568 356 3632
rect 420 3568 421 3632
rect 355 3552 421 3568
rect 355 3488 356 3552
rect 420 3488 421 3552
rect 355 3472 421 3488
rect 355 3408 356 3472
rect 420 3408 421 3472
rect 355 3392 421 3408
rect 355 3328 356 3392
rect 420 3328 421 3392
rect 355 3312 421 3328
rect 355 3248 356 3312
rect 420 3248 421 3312
rect 355 3232 421 3248
rect 355 3168 356 3232
rect 420 3168 421 3232
rect 355 3152 421 3168
rect 355 3088 356 3152
rect 420 3088 421 3152
rect 355 3087 421 3088
rect 355 3072 360 3087
rect 416 3072 421 3087
rect 355 3008 356 3072
rect 420 3008 421 3072
rect 355 2992 421 3008
rect 355 2928 356 2992
rect 420 2928 421 2992
rect 355 2916 421 2928
rect 355 2860 360 2916
rect 416 2860 421 2916
rect 355 2838 421 2860
rect 481 2774 541 3804
rect 601 2834 661 3866
rect 721 2774 781 3804
rect 841 2834 901 3866
rect 961 3712 1027 3866
rect 961 3648 962 3712
rect 1026 3648 1027 3712
rect 961 3632 1027 3648
rect 961 3568 962 3632
rect 1026 3568 1027 3632
rect 961 3552 1027 3568
rect 961 3488 962 3552
rect 1026 3488 1027 3552
rect 961 3472 1027 3488
rect 961 3408 962 3472
rect 1026 3408 1027 3472
rect 961 3392 1027 3408
rect 961 3328 962 3392
rect 1026 3328 1027 3392
rect 961 3312 1027 3328
rect 961 3248 962 3312
rect 1026 3248 1027 3312
rect 961 3232 1027 3248
rect 961 3168 962 3232
rect 1026 3168 1027 3232
rect 961 3152 1027 3168
rect 961 3088 962 3152
rect 1026 3088 1027 3152
rect 961 3072 1027 3088
rect 961 3008 962 3072
rect 1026 3008 1027 3072
rect 961 2992 1027 3008
rect 961 2928 962 2992
rect 1026 2928 1027 2992
rect 961 2838 1027 2928
rect 1267 4872 1333 4962
rect 1267 4808 1268 4872
rect 1332 4808 1333 4872
rect 1267 4792 1333 4808
rect 1267 4728 1268 4792
rect 1332 4728 1333 4792
rect 1267 4712 1333 4728
rect 1267 4648 1268 4712
rect 1332 4648 1333 4712
rect 1267 4632 1333 4648
rect 1267 4568 1268 4632
rect 1332 4568 1333 4632
rect 1267 4552 1333 4568
rect 1267 4488 1268 4552
rect 1332 4488 1333 4552
rect 1267 4472 1333 4488
rect 1267 4408 1268 4472
rect 1332 4408 1333 4472
rect 1267 4392 1333 4408
rect 1267 4328 1268 4392
rect 1332 4328 1333 4392
rect 1267 4312 1333 4328
rect 1267 4248 1268 4312
rect 1332 4248 1333 4312
rect 1267 4232 1333 4248
rect 1267 4168 1268 4232
rect 1332 4168 1333 4232
rect 1267 4152 1333 4168
rect 1267 4088 1268 4152
rect 1332 4088 1333 4152
rect 1267 3934 1333 4088
rect 1393 3934 1453 4966
rect 1513 3996 1573 5026
rect 1633 3934 1693 4966
rect 1753 3996 1813 5026
rect 1873 4872 1939 4962
rect 1873 4808 1874 4872
rect 1938 4808 1939 4872
rect 1873 4792 1939 4808
rect 1873 4728 1874 4792
rect 1938 4728 1939 4792
rect 1873 4712 1939 4728
rect 1873 4648 1874 4712
rect 1938 4648 1939 4712
rect 1873 4632 1939 4648
rect 1873 4568 1874 4632
rect 1938 4568 1939 4632
rect 1873 4552 1939 4568
rect 1873 4488 1874 4552
rect 1938 4488 1939 4552
rect 1873 4472 1939 4488
rect 1873 4408 1874 4472
rect 1938 4408 1939 4472
rect 1873 4392 1939 4408
rect 1873 4328 1874 4392
rect 1938 4328 1939 4392
rect 1873 4312 1939 4328
rect 1873 4248 1874 4312
rect 1938 4248 1939 4312
rect 1873 4232 1939 4248
rect 1873 4168 1874 4232
rect 1938 4168 1939 4232
rect 1873 4152 1939 4168
rect 1873 4088 1874 4152
rect 1938 4088 1939 4152
rect 1873 3934 1939 4088
rect 1999 3934 2059 4966
rect 2119 3996 2179 5026
rect 2239 3934 2299 4966
rect 2359 3996 2419 5026
rect 2479 4872 2545 4962
rect 2479 4808 2480 4872
rect 2544 4808 2545 4872
rect 2479 4792 2545 4808
rect 2479 4728 2480 4792
rect 2544 4728 2545 4792
rect 2479 4712 2545 4728
rect 2479 4648 2480 4712
rect 2544 4648 2545 4712
rect 2479 4632 2545 4648
rect 2479 4568 2480 4632
rect 2544 4568 2545 4632
rect 2479 4552 2545 4568
rect 2479 4488 2480 4552
rect 2544 4488 2545 4552
rect 2479 4472 2545 4488
rect 2479 4408 2480 4472
rect 2544 4408 2545 4472
rect 2479 4392 2545 4408
rect 2479 4328 2480 4392
rect 2544 4328 2545 4392
rect 2479 4312 2545 4328
rect 2479 4248 2480 4312
rect 2544 4248 2545 4312
rect 2479 4232 2545 4248
rect 2479 4168 2480 4232
rect 2544 4168 2545 4232
rect 2479 4152 2545 4168
rect 2479 4088 2480 4152
rect 2544 4088 2545 4152
rect 2479 3934 2545 4088
rect 1267 3932 2545 3934
rect 1267 3868 1371 3932
rect 1435 3868 1451 3932
rect 1515 3868 1531 3932
rect 1595 3868 1611 3932
rect 1675 3868 1691 3932
rect 1755 3868 1771 3932
rect 1835 3868 1977 3932
rect 2041 3868 2057 3932
rect 2121 3868 2137 3932
rect 2201 3868 2217 3932
rect 2281 3868 2297 3932
rect 2361 3868 2377 3932
rect 2441 3868 2545 3932
rect 1267 3866 2545 3868
rect 1267 3712 1333 3866
rect 1267 3648 1268 3712
rect 1332 3648 1333 3712
rect 1267 3632 1333 3648
rect 1267 3568 1268 3632
rect 1332 3568 1333 3632
rect 1267 3552 1333 3568
rect 1267 3488 1268 3552
rect 1332 3488 1333 3552
rect 1267 3472 1333 3488
rect 1267 3408 1268 3472
rect 1332 3408 1333 3472
rect 1267 3392 1333 3408
rect 1267 3328 1268 3392
rect 1332 3328 1333 3392
rect 1267 3312 1333 3328
rect 1267 3248 1268 3312
rect 1332 3248 1333 3312
rect 1267 3232 1333 3248
rect 1267 3168 1268 3232
rect 1332 3168 1333 3232
rect 1267 3152 1333 3168
rect 1267 3088 1268 3152
rect 1332 3088 1333 3152
rect 1267 3072 1333 3088
rect 1267 3008 1268 3072
rect 1332 3008 1333 3072
rect 1267 2992 1333 3008
rect 1267 2928 1268 2992
rect 1332 2928 1333 2992
rect 1267 2916 1333 2928
rect 1267 2860 1272 2916
rect 1328 2860 1333 2916
rect 1267 2838 1333 2860
rect 1393 2774 1453 3804
rect 1513 2834 1573 3866
rect 1633 2774 1693 3804
rect 1753 2834 1813 3866
rect 1873 3712 1939 3866
rect 1873 3648 1874 3712
rect 1938 3648 1939 3712
rect 1873 3632 1939 3648
rect 1873 3568 1874 3632
rect 1938 3568 1939 3632
rect 1873 3552 1939 3568
rect 1873 3488 1874 3552
rect 1938 3488 1939 3552
rect 1873 3472 1939 3488
rect 1873 3408 1874 3472
rect 1938 3408 1939 3472
rect 1873 3392 1939 3408
rect 1873 3328 1874 3392
rect 1938 3328 1939 3392
rect 1873 3312 1939 3328
rect 1873 3248 1874 3312
rect 1938 3248 1939 3312
rect 1873 3232 1939 3248
rect 1873 3168 1874 3232
rect 1938 3168 1939 3232
rect 1873 3152 1939 3168
rect 1873 3088 1874 3152
rect 1938 3088 1939 3152
rect 1873 3072 1939 3088
rect 1873 3008 1874 3072
rect 1938 3008 1939 3072
rect 1873 2992 1939 3008
rect 1873 2928 1874 2992
rect 1938 2928 1939 2992
rect 1873 2915 1939 2928
rect 1873 2859 1878 2915
rect 1934 2859 1939 2915
rect 1873 2838 1939 2859
rect 1999 2774 2059 3804
rect 2119 2834 2179 3866
rect 2239 2774 2299 3804
rect 2359 2834 2419 3866
rect 2479 3712 2545 3866
rect 2479 3648 2480 3712
rect 2544 3648 2545 3712
rect 2479 3632 2545 3648
rect 2479 3568 2480 3632
rect 2544 3568 2545 3632
rect 2479 3552 2545 3568
rect 2479 3488 2480 3552
rect 2544 3488 2545 3552
rect 2479 3472 2545 3488
rect 2479 3408 2480 3472
rect 2544 3408 2545 3472
rect 2479 3392 2545 3408
rect 2479 3328 2480 3392
rect 2544 3328 2545 3392
rect 2479 3312 2545 3328
rect 2479 3248 2480 3312
rect 2544 3248 2545 3312
rect 2479 3232 2545 3248
rect 2479 3168 2480 3232
rect 2544 3168 2545 3232
rect 2479 3152 2545 3168
rect 2479 3088 2480 3152
rect 2544 3088 2545 3152
rect 2479 3072 2545 3088
rect 2479 3008 2480 3072
rect 2544 3008 2545 3072
rect 2479 2992 2545 3008
rect 2479 2928 2480 2992
rect 2544 2928 2545 2992
rect 2479 2838 2545 2928
rect 2801 4872 2867 4962
rect 2801 4808 2802 4872
rect 2866 4808 2867 4872
rect 2801 4792 2867 4808
rect 2801 4728 2802 4792
rect 2866 4728 2867 4792
rect 2801 4712 2867 4728
rect 2801 4648 2802 4712
rect 2866 4648 2867 4712
rect 2801 4632 2867 4648
rect 2801 4568 2802 4632
rect 2866 4568 2867 4632
rect 2801 4552 2867 4568
rect 2801 4488 2802 4552
rect 2866 4488 2867 4552
rect 2801 4472 2867 4488
rect 2801 4408 2802 4472
rect 2866 4408 2867 4472
rect 2801 4392 2867 4408
rect 2801 4328 2802 4392
rect 2866 4328 2867 4392
rect 2801 4312 2867 4328
rect 2801 4248 2802 4312
rect 2866 4248 2867 4312
rect 2801 4232 2867 4248
rect 2801 4168 2802 4232
rect 2866 4168 2867 4232
rect 2801 4152 2867 4168
rect 2801 4088 2802 4152
rect 2866 4088 2867 4152
rect 2801 3934 2867 4088
rect 2927 3934 2987 4966
rect 3047 3996 3107 5026
rect 3167 3934 3227 4966
rect 3287 3996 3347 5026
rect 3407 4872 3473 4962
rect 3407 4808 3408 4872
rect 3472 4808 3473 4872
rect 3407 4792 3473 4808
rect 3407 4728 3408 4792
rect 3472 4728 3473 4792
rect 3407 4712 3473 4728
rect 3407 4648 3408 4712
rect 3472 4648 3473 4712
rect 3407 4632 3473 4648
rect 3407 4568 3408 4632
rect 3472 4568 3473 4632
rect 3407 4552 3473 4568
rect 3407 4488 3408 4552
rect 3472 4488 3473 4552
rect 3407 4472 3473 4488
rect 3407 4408 3408 4472
rect 3472 4408 3473 4472
rect 3407 4392 3473 4408
rect 3407 4328 3408 4392
rect 3472 4328 3473 4392
rect 3407 4312 3473 4328
rect 3407 4248 3408 4312
rect 3472 4248 3473 4312
rect 3407 4232 3473 4248
rect 3407 4168 3408 4232
rect 3472 4168 3473 4232
rect 3407 4152 3473 4168
rect 3407 4088 3408 4152
rect 3472 4088 3473 4152
rect 3407 3934 3473 4088
rect 3533 3934 3593 4966
rect 3653 3996 3713 5026
rect 3773 3934 3833 4966
rect 3893 3996 3953 5026
rect 4013 4872 4079 4962
rect 4013 4808 4014 4872
rect 4078 4808 4079 4872
rect 4013 4792 4079 4808
rect 4013 4728 4014 4792
rect 4078 4728 4079 4792
rect 4013 4712 4079 4728
rect 4013 4648 4014 4712
rect 4078 4648 4079 4712
rect 4013 4632 4079 4648
rect 4013 4568 4014 4632
rect 4078 4568 4079 4632
rect 4013 4552 4079 4568
rect 4013 4488 4014 4552
rect 4078 4488 4079 4552
rect 4013 4472 4079 4488
rect 4013 4408 4014 4472
rect 4078 4408 4079 4472
rect 4013 4392 4079 4408
rect 4013 4328 4014 4392
rect 4078 4328 4079 4392
rect 4013 4312 4079 4328
rect 4013 4248 4014 4312
rect 4078 4248 4079 4312
rect 4013 4232 4079 4248
rect 4013 4168 4014 4232
rect 4078 4168 4079 4232
rect 4013 4152 4079 4168
rect 4013 4088 4014 4152
rect 4078 4088 4079 4152
rect 4013 3934 4079 4088
rect 4139 3934 4199 4966
rect 4259 3996 4319 5026
rect 4379 3934 4439 4966
rect 4499 3996 4559 5026
rect 4619 4872 4685 4962
rect 4619 4808 4620 4872
rect 4684 4808 4685 4872
rect 4619 4792 4685 4808
rect 4619 4728 4620 4792
rect 4684 4728 4685 4792
rect 4619 4712 4685 4728
rect 4619 4648 4620 4712
rect 4684 4648 4685 4712
rect 4619 4632 4685 4648
rect 4619 4568 4620 4632
rect 4684 4568 4685 4632
rect 4619 4552 4685 4568
rect 4619 4488 4620 4552
rect 4684 4488 4685 4552
rect 4619 4472 4685 4488
rect 4619 4408 4620 4472
rect 4684 4408 4685 4472
rect 4619 4392 4685 4408
rect 4619 4328 4620 4392
rect 4684 4328 4685 4392
rect 4619 4312 4685 4328
rect 4619 4248 4620 4312
rect 4684 4248 4685 4312
rect 4619 4232 4685 4248
rect 4619 4168 4620 4232
rect 4684 4168 4685 4232
rect 4619 4152 4685 4168
rect 4619 4088 4620 4152
rect 4684 4088 4685 4152
rect 4619 3934 4685 4088
rect 4745 3934 4805 4966
rect 4865 3996 4925 5026
rect 4985 3934 5045 4966
rect 5105 3996 5165 5026
rect 5225 4872 5291 4962
rect 5225 4808 5226 4872
rect 5290 4808 5291 4872
rect 5225 4792 5291 4808
rect 5225 4728 5226 4792
rect 5290 4728 5291 4792
rect 5225 4712 5291 4728
rect 5225 4648 5226 4712
rect 5290 4648 5291 4712
rect 5225 4632 5291 4648
rect 5225 4568 5226 4632
rect 5290 4568 5291 4632
rect 5225 4552 5291 4568
rect 5225 4488 5226 4552
rect 5290 4488 5291 4552
rect 5225 4472 5291 4488
rect 5225 4408 5226 4472
rect 5290 4408 5291 4472
rect 5225 4392 5291 4408
rect 5225 4328 5226 4392
rect 5290 4328 5291 4392
rect 5225 4312 5291 4328
rect 5225 4248 5226 4312
rect 5290 4248 5291 4312
rect 5225 4232 5291 4248
rect 5225 4168 5226 4232
rect 5290 4168 5291 4232
rect 5225 4152 5291 4168
rect 5225 4088 5226 4152
rect 5290 4088 5291 4152
rect 5225 3934 5291 4088
rect 2801 3932 5291 3934
rect 2801 3868 2905 3932
rect 2969 3868 2985 3932
rect 3049 3868 3065 3932
rect 3129 3868 3145 3932
rect 3209 3868 3225 3932
rect 3289 3868 3305 3932
rect 3369 3868 3511 3932
rect 3575 3868 3591 3932
rect 3655 3868 3671 3932
rect 3735 3868 3751 3932
rect 3815 3868 3831 3932
rect 3895 3868 3911 3932
rect 3975 3868 4117 3932
rect 4181 3868 4197 3932
rect 4261 3868 4277 3932
rect 4341 3868 4357 3932
rect 4421 3868 4437 3932
rect 4501 3868 4517 3932
rect 4581 3868 4723 3932
rect 4787 3868 4803 3932
rect 4867 3868 4883 3932
rect 4947 3868 4963 3932
rect 5027 3868 5043 3932
rect 5107 3927 5123 3932
rect 5107 3868 5123 3871
rect 5187 3868 5291 3932
rect 2801 3866 5291 3868
rect 2801 3712 2867 3866
rect 2801 3648 2802 3712
rect 2866 3648 2867 3712
rect 2801 3632 2867 3648
rect 2801 3568 2802 3632
rect 2866 3568 2867 3632
rect 2801 3552 2867 3568
rect 2801 3488 2802 3552
rect 2866 3488 2867 3552
rect 2801 3472 2867 3488
rect 2801 3408 2802 3472
rect 2866 3408 2867 3472
rect 2801 3392 2867 3408
rect 2801 3328 2802 3392
rect 2866 3328 2867 3392
rect 2801 3312 2867 3328
rect 2801 3248 2802 3312
rect 2866 3248 2867 3312
rect 2801 3232 2867 3248
rect 2801 3168 2802 3232
rect 2866 3168 2867 3232
rect 2801 3152 2867 3168
rect 2801 3088 2802 3152
rect 2866 3088 2867 3152
rect 2801 3072 2867 3088
rect 2801 3008 2802 3072
rect 2866 3008 2867 3072
rect 2801 2992 2867 3008
rect 2801 2928 2802 2992
rect 2866 2928 2867 2992
rect 2801 2914 2867 2928
rect 2801 2858 2806 2914
rect 2862 2858 2867 2914
rect 2801 2838 2867 2858
rect 2927 2774 2987 3804
rect 3047 2834 3107 3866
rect 3167 2774 3227 3804
rect 3287 2834 3347 3866
rect 3407 3712 3473 3866
rect 3407 3648 3408 3712
rect 3472 3648 3473 3712
rect 3407 3632 3473 3648
rect 3407 3568 3408 3632
rect 3472 3568 3473 3632
rect 3407 3552 3473 3568
rect 3407 3488 3408 3552
rect 3472 3488 3473 3552
rect 3407 3472 3473 3488
rect 3407 3408 3408 3472
rect 3472 3408 3473 3472
rect 3407 3392 3473 3408
rect 3407 3328 3408 3392
rect 3472 3328 3473 3392
rect 3407 3312 3473 3328
rect 3407 3248 3408 3312
rect 3472 3248 3473 3312
rect 3407 3232 3473 3248
rect 3407 3168 3408 3232
rect 3472 3168 3473 3232
rect 3407 3152 3473 3168
rect 3407 3088 3408 3152
rect 3472 3088 3473 3152
rect 3407 3072 3473 3088
rect 3407 3008 3408 3072
rect 3472 3008 3473 3072
rect 3407 2992 3473 3008
rect 3407 2928 3408 2992
rect 3472 2928 3473 2992
rect 3407 2838 3473 2928
rect 3533 2774 3593 3804
rect 3653 2834 3713 3866
rect 3773 2774 3833 3804
rect 3893 2834 3953 3866
rect 4013 3712 4079 3866
rect 4013 3648 4014 3712
rect 4078 3648 4079 3712
rect 4013 3632 4079 3648
rect 4013 3568 4014 3632
rect 4078 3568 4079 3632
rect 4013 3552 4079 3568
rect 4013 3488 4014 3552
rect 4078 3488 4079 3552
rect 4013 3472 4079 3488
rect 4013 3408 4014 3472
rect 4078 3408 4079 3472
rect 4013 3392 4079 3408
rect 4013 3328 4014 3392
rect 4078 3328 4079 3392
rect 4013 3312 4079 3328
rect 4013 3248 4014 3312
rect 4078 3248 4079 3312
rect 4013 3232 4079 3248
rect 4013 3168 4014 3232
rect 4078 3168 4079 3232
rect 4013 3152 4079 3168
rect 4013 3088 4014 3152
rect 4078 3088 4079 3152
rect 4013 3072 4079 3088
rect 4013 3008 4014 3072
rect 4078 3008 4079 3072
rect 4013 2992 4079 3008
rect 4013 2928 4014 2992
rect 4078 2928 4079 2992
rect 4013 2916 4079 2928
rect 4013 2860 4018 2916
rect 4074 2860 4079 2916
rect 4013 2838 4079 2860
rect 4139 2774 4199 3804
rect 4259 2834 4319 3866
rect 4379 2774 4439 3804
rect 4499 2834 4559 3866
rect 4619 3712 4685 3866
rect 4619 3648 4620 3712
rect 4684 3648 4685 3712
rect 4619 3632 4685 3648
rect 4619 3568 4620 3632
rect 4684 3568 4685 3632
rect 4619 3552 4685 3568
rect 4619 3488 4620 3552
rect 4684 3488 4685 3552
rect 4619 3472 4685 3488
rect 4619 3408 4620 3472
rect 4684 3408 4685 3472
rect 4619 3392 4685 3408
rect 4619 3328 4620 3392
rect 4684 3328 4685 3392
rect 4619 3312 4685 3328
rect 4619 3248 4620 3312
rect 4684 3248 4685 3312
rect 4619 3232 4685 3248
rect 4619 3168 4620 3232
rect 4684 3168 4685 3232
rect 4619 3152 4685 3168
rect 4619 3088 4620 3152
rect 4684 3088 4685 3152
rect 4619 3072 4685 3088
rect 4619 3008 4620 3072
rect 4684 3008 4685 3072
rect 4619 2992 4685 3008
rect 4619 2928 4620 2992
rect 4684 2928 4685 2992
rect 4619 2838 4685 2928
rect 4745 2774 4805 3804
rect 4865 2834 4925 3866
rect 4985 2774 5045 3804
rect 5105 2834 5165 3866
rect 5225 3712 5291 3866
rect 5225 3648 5226 3712
rect 5290 3648 5291 3712
rect 5225 3632 5291 3648
rect 5225 3568 5226 3632
rect 5290 3568 5291 3632
rect 5225 3552 5291 3568
rect 5225 3488 5226 3552
rect 5290 3488 5291 3552
rect 5225 3472 5291 3488
rect 5225 3408 5226 3472
rect 5290 3408 5291 3472
rect 5225 3392 5291 3408
rect 5225 3328 5226 3392
rect 5290 3328 5291 3392
rect 5225 3312 5291 3328
rect 5225 3248 5226 3312
rect 5290 3248 5291 3312
rect 5225 3232 5291 3248
rect 5225 3168 5226 3232
rect 5290 3168 5291 3232
rect 5225 3152 5291 3168
rect 5225 3088 5226 3152
rect 5290 3088 5291 3152
rect 5225 3072 5291 3088
rect 5225 3008 5226 3072
rect 5290 3008 5291 3072
rect 5225 2992 5291 3008
rect 5225 2928 5226 2992
rect 5290 2928 5291 2992
rect 5225 2838 5291 2928
rect 5352 4872 5418 4962
rect 5352 4808 5353 4872
rect 5417 4808 5418 4872
rect 5352 4792 5418 4808
rect 5352 4728 5353 4792
rect 5417 4728 5418 4792
rect 5352 4712 5418 4728
rect 5352 4648 5353 4712
rect 5417 4648 5418 4712
rect 5352 4632 5418 4648
rect 5352 4568 5353 4632
rect 5417 4568 5418 4632
rect 5352 4552 5418 4568
rect 5352 4488 5353 4552
rect 5417 4488 5418 4552
rect 5352 4472 5418 4488
rect 5352 4408 5353 4472
rect 5417 4408 5418 4472
rect 5352 4392 5418 4408
rect 5352 4328 5353 4392
rect 5417 4328 5418 4392
rect 5352 4312 5418 4328
rect 5352 4248 5353 4312
rect 5417 4248 5418 4312
rect 5352 4232 5418 4248
rect 5352 4168 5353 4232
rect 5417 4168 5418 4232
rect 5352 4152 5418 4168
rect 5352 4088 5353 4152
rect 5417 4088 5418 4152
rect 5352 3934 5418 4088
rect 5478 3934 5538 4966
rect 5598 3996 5658 5026
rect 5718 3934 5778 4966
rect 5838 3996 5898 5026
rect 5958 4872 6024 4962
rect 5958 4808 5959 4872
rect 6023 4808 6024 4872
rect 5958 4792 6024 4808
rect 5958 4728 5959 4792
rect 6023 4728 6024 4792
rect 5958 4712 6024 4728
rect 5958 4648 5959 4712
rect 6023 4648 6024 4712
rect 5958 4632 6024 4648
rect 5958 4568 5959 4632
rect 6023 4568 6024 4632
rect 5958 4552 6024 4568
rect 5958 4488 5959 4552
rect 6023 4488 6024 4552
rect 5958 4472 6024 4488
rect 5958 4408 5959 4472
rect 6023 4408 6024 4472
rect 5958 4392 6024 4408
rect 5958 4328 5959 4392
rect 6023 4328 6024 4392
rect 5958 4312 6024 4328
rect 5958 4248 5959 4312
rect 6023 4248 6024 4312
rect 5958 4232 6024 4248
rect 5958 4168 5959 4232
rect 6023 4168 6024 4232
rect 5958 4152 6024 4168
rect 5958 4088 5959 4152
rect 6023 4088 6024 4152
rect 5958 3934 6024 4088
rect 6084 3934 6144 4966
rect 6204 3996 6264 5026
rect 6324 3934 6384 4966
rect 6444 3996 6504 5026
rect 6564 4872 6630 4962
rect 6564 4808 6565 4872
rect 6629 4808 6630 4872
rect 6564 4792 6630 4808
rect 6564 4728 6565 4792
rect 6629 4728 6630 4792
rect 6564 4712 6630 4728
rect 6564 4648 6565 4712
rect 6629 4648 6630 4712
rect 6564 4632 6630 4648
rect 6564 4568 6565 4632
rect 6629 4568 6630 4632
rect 6564 4552 6630 4568
rect 6564 4488 6565 4552
rect 6629 4488 6630 4552
rect 6564 4472 6630 4488
rect 6564 4408 6565 4472
rect 6629 4408 6630 4472
rect 6564 4392 6630 4408
rect 6564 4328 6565 4392
rect 6629 4328 6630 4392
rect 6564 4312 6630 4328
rect 6564 4248 6565 4312
rect 6629 4248 6630 4312
rect 6564 4232 6630 4248
rect 6564 4168 6565 4232
rect 6629 4168 6630 4232
rect 6564 4152 6630 4168
rect 6564 4088 6565 4152
rect 6629 4088 6630 4152
rect 6564 3934 6630 4088
rect 6690 3934 6750 4966
rect 6810 3996 6870 5026
rect 6930 3934 6990 4966
rect 7050 3996 7110 5026
rect 7170 4872 7236 4962
rect 7170 4808 7171 4872
rect 7235 4808 7236 4872
rect 7170 4792 7236 4808
rect 7170 4728 7171 4792
rect 7235 4728 7236 4792
rect 7170 4712 7236 4728
rect 7170 4648 7171 4712
rect 7235 4648 7236 4712
rect 7170 4632 7236 4648
rect 7170 4568 7171 4632
rect 7235 4568 7236 4632
rect 7170 4552 7236 4568
rect 7170 4488 7171 4552
rect 7235 4488 7236 4552
rect 7170 4472 7236 4488
rect 7170 4408 7171 4472
rect 7235 4408 7236 4472
rect 7170 4392 7236 4408
rect 7170 4328 7171 4392
rect 7235 4328 7236 4392
rect 7170 4312 7236 4328
rect 7170 4248 7171 4312
rect 7235 4248 7236 4312
rect 7170 4232 7236 4248
rect 7170 4168 7171 4232
rect 7235 4168 7236 4232
rect 7170 4152 7236 4168
rect 7170 4088 7171 4152
rect 7235 4088 7236 4152
rect 7170 3934 7236 4088
rect 7296 3934 7356 4966
rect 7416 3996 7476 5026
rect 7536 3934 7596 4966
rect 7656 3996 7716 5026
rect 7776 4872 7842 4962
rect 7776 4808 7777 4872
rect 7841 4808 7842 4872
rect 7776 4792 7842 4808
rect 7776 4728 7777 4792
rect 7841 4728 7842 4792
rect 7776 4712 7842 4728
rect 7776 4648 7777 4712
rect 7841 4648 7842 4712
rect 7776 4632 7842 4648
rect 7776 4568 7777 4632
rect 7841 4568 7842 4632
rect 7776 4552 7842 4568
rect 7776 4488 7777 4552
rect 7841 4488 7842 4552
rect 7776 4472 7842 4488
rect 7776 4408 7777 4472
rect 7841 4408 7842 4472
rect 7776 4392 7842 4408
rect 7776 4328 7777 4392
rect 7841 4328 7842 4392
rect 7776 4312 7842 4328
rect 7776 4248 7777 4312
rect 7841 4248 7842 4312
rect 7776 4232 7842 4248
rect 7776 4168 7777 4232
rect 7841 4168 7842 4232
rect 7776 4152 7842 4168
rect 7776 4088 7777 4152
rect 7841 4088 7842 4152
rect 7776 3934 7842 4088
rect 7902 3934 7962 4966
rect 8022 3996 8082 5026
rect 8142 3934 8202 4966
rect 8262 3996 8322 5026
rect 8382 4872 8448 4962
rect 8382 4808 8383 4872
rect 8447 4808 8448 4872
rect 8382 4792 8448 4808
rect 8382 4728 8383 4792
rect 8447 4728 8448 4792
rect 8382 4712 8448 4728
rect 8382 4648 8383 4712
rect 8447 4648 8448 4712
rect 8382 4632 8448 4648
rect 8382 4568 8383 4632
rect 8447 4568 8448 4632
rect 8382 4552 8448 4568
rect 8382 4488 8383 4552
rect 8447 4488 8448 4552
rect 8382 4472 8448 4488
rect 8382 4408 8383 4472
rect 8447 4408 8448 4472
rect 8382 4392 8448 4408
rect 8382 4328 8383 4392
rect 8447 4328 8448 4392
rect 8382 4312 8448 4328
rect 8382 4248 8383 4312
rect 8447 4248 8448 4312
rect 8382 4232 8448 4248
rect 8382 4168 8383 4232
rect 8447 4168 8448 4232
rect 8382 4152 8448 4168
rect 8382 4088 8383 4152
rect 8447 4088 8448 4152
rect 8382 3934 8448 4088
rect 8508 3934 8568 4966
rect 8628 3996 8688 5026
rect 8748 3934 8808 4966
rect 8868 3996 8928 5026
rect 8988 4872 9054 4962
rect 8988 4808 8989 4872
rect 9053 4808 9054 4872
rect 8988 4792 9054 4808
rect 8988 4728 8989 4792
rect 9053 4728 9054 4792
rect 8988 4712 9054 4728
rect 8988 4648 8989 4712
rect 9053 4648 9054 4712
rect 8988 4632 9054 4648
rect 8988 4568 8989 4632
rect 9053 4568 9054 4632
rect 8988 4552 9054 4568
rect 8988 4488 8989 4552
rect 9053 4488 9054 4552
rect 8988 4472 9054 4488
rect 8988 4408 8989 4472
rect 9053 4408 9054 4472
rect 8988 4392 9054 4408
rect 8988 4328 8989 4392
rect 9053 4328 9054 4392
rect 8988 4312 9054 4328
rect 8988 4248 8989 4312
rect 9053 4248 9054 4312
rect 8988 4232 9054 4248
rect 8988 4168 8989 4232
rect 9053 4168 9054 4232
rect 8988 4152 9054 4168
rect 8988 4088 8989 4152
rect 9053 4088 9054 4152
rect 8988 3934 9054 4088
rect 9114 3934 9174 4966
rect 9234 3996 9294 5026
rect 9354 3934 9414 4966
rect 9474 3996 9534 5026
rect 9594 4872 9660 4962
rect 9594 4808 9595 4872
rect 9659 4808 9660 4872
rect 9594 4792 9660 4808
rect 9594 4728 9595 4792
rect 9659 4728 9660 4792
rect 9594 4712 9660 4728
rect 9594 4648 9595 4712
rect 9659 4648 9660 4712
rect 9594 4632 9660 4648
rect 9594 4568 9595 4632
rect 9659 4568 9660 4632
rect 9594 4552 9660 4568
rect 9594 4488 9595 4552
rect 9659 4488 9660 4552
rect 9594 4472 9660 4488
rect 9594 4408 9595 4472
rect 9659 4408 9660 4472
rect 9594 4392 9660 4408
rect 9594 4328 9595 4392
rect 9659 4328 9660 4392
rect 9594 4312 9660 4328
rect 9594 4248 9595 4312
rect 9659 4248 9660 4312
rect 9594 4232 9660 4248
rect 9594 4168 9595 4232
rect 9659 4168 9660 4232
rect 9594 4152 9660 4168
rect 9594 4088 9595 4152
rect 9659 4088 9660 4152
rect 9594 3934 9660 4088
rect 9720 3934 9780 4966
rect 9840 3996 9900 5026
rect 9960 3934 10020 4966
rect 10080 3996 10140 5026
rect 10200 4872 10266 4962
rect 10200 4808 10201 4872
rect 10265 4808 10266 4872
rect 10200 4792 10266 4808
rect 10200 4728 10201 4792
rect 10265 4728 10266 4792
rect 10200 4712 10266 4728
rect 10200 4648 10201 4712
rect 10265 4648 10266 4712
rect 10200 4632 10266 4648
rect 10200 4568 10201 4632
rect 10265 4568 10266 4632
rect 10200 4552 10266 4568
rect 10200 4488 10201 4552
rect 10265 4488 10266 4552
rect 10200 4472 10266 4488
rect 10200 4408 10201 4472
rect 10265 4408 10266 4472
rect 10200 4392 10266 4408
rect 10200 4328 10201 4392
rect 10265 4328 10266 4392
rect 10200 4312 10266 4328
rect 10200 4248 10201 4312
rect 10265 4248 10266 4312
rect 10200 4232 10266 4248
rect 10200 4168 10201 4232
rect 10265 4168 10266 4232
rect 10200 4152 10266 4168
rect 10200 4088 10201 4152
rect 10265 4088 10266 4152
rect 10200 3934 10266 4088
rect 5352 3932 10266 3934
rect 5352 3868 5456 3932
rect 5520 3868 5536 3932
rect 5600 3868 5616 3932
rect 5680 3868 5696 3932
rect 5760 3868 5776 3932
rect 5840 3868 5856 3932
rect 5920 3868 6062 3932
rect 6126 3868 6142 3932
rect 6206 3868 6222 3932
rect 6286 3868 6302 3932
rect 6366 3868 6382 3932
rect 6446 3868 6462 3932
rect 6526 3868 6668 3932
rect 6732 3868 6748 3932
rect 6812 3868 6828 3932
rect 6892 3868 6908 3932
rect 6972 3868 6988 3932
rect 7052 3868 7068 3932
rect 7132 3868 7274 3932
rect 7338 3868 7354 3932
rect 7418 3868 7434 3932
rect 7498 3868 7514 3932
rect 7578 3868 7594 3932
rect 7658 3868 7674 3932
rect 7738 3868 7880 3932
rect 7944 3868 7960 3932
rect 8024 3868 8040 3932
rect 8104 3868 8120 3932
rect 8184 3868 8200 3932
rect 8264 3868 8280 3932
rect 8344 3868 8486 3932
rect 8550 3868 8566 3932
rect 8630 3868 8646 3932
rect 8710 3868 8726 3932
rect 8790 3868 8806 3932
rect 8870 3868 8886 3932
rect 8950 3868 9092 3932
rect 9156 3868 9172 3932
rect 9236 3868 9252 3932
rect 9316 3868 9332 3932
rect 9396 3868 9412 3932
rect 9476 3868 9492 3932
rect 9556 3868 9698 3932
rect 9762 3868 9778 3932
rect 9842 3868 9858 3932
rect 9922 3868 9938 3932
rect 10002 3868 10018 3932
rect 10082 3868 10098 3932
rect 10162 3868 10266 3932
rect 5352 3866 10266 3868
rect 5352 3712 5418 3866
rect 5352 3648 5353 3712
rect 5417 3648 5418 3712
rect 5352 3632 5418 3648
rect 5352 3568 5353 3632
rect 5417 3568 5418 3632
rect 5352 3552 5418 3568
rect 5352 3488 5353 3552
rect 5417 3488 5418 3552
rect 5352 3472 5418 3488
rect 5352 3408 5353 3472
rect 5417 3408 5418 3472
rect 5352 3392 5418 3408
rect 5352 3328 5353 3392
rect 5417 3328 5418 3392
rect 5352 3312 5418 3328
rect 5352 3248 5353 3312
rect 5417 3248 5418 3312
rect 5352 3232 5418 3248
rect 5352 3168 5353 3232
rect 5417 3168 5418 3232
rect 5352 3152 5418 3168
rect 5352 3088 5353 3152
rect 5417 3088 5418 3152
rect 5352 3072 5418 3088
rect 5352 3008 5353 3072
rect 5417 3008 5418 3072
rect 5352 2992 5418 3008
rect 5352 2928 5353 2992
rect 5417 2928 5418 2992
rect 5352 2909 5418 2928
rect 5352 2853 5357 2909
rect 5413 2853 5418 2909
rect 5352 2838 5418 2853
rect 5478 2774 5538 3804
rect 5598 2834 5658 3866
rect 5718 2774 5778 3804
rect 5838 2834 5898 3866
rect 5958 3712 6024 3866
rect 5958 3648 5959 3712
rect 6023 3648 6024 3712
rect 5958 3632 6024 3648
rect 5958 3568 5959 3632
rect 6023 3568 6024 3632
rect 5958 3552 6024 3568
rect 5958 3488 5959 3552
rect 6023 3488 6024 3552
rect 5958 3472 6024 3488
rect 5958 3408 5959 3472
rect 6023 3408 6024 3472
rect 5958 3392 6024 3408
rect 5958 3328 5959 3392
rect 6023 3328 6024 3392
rect 5958 3312 6024 3328
rect 5958 3248 5959 3312
rect 6023 3248 6024 3312
rect 5958 3232 6024 3248
rect 5958 3168 5959 3232
rect 6023 3168 6024 3232
rect 5958 3152 6024 3168
rect 5958 3088 5959 3152
rect 6023 3088 6024 3152
rect 5958 3072 6024 3088
rect 5958 3008 5959 3072
rect 6023 3008 6024 3072
rect 5958 2992 6024 3008
rect 5958 2928 5959 2992
rect 6023 2928 6024 2992
rect 5958 2907 6024 2928
rect 5958 2851 5963 2907
rect 6019 2851 6024 2907
rect 5958 2838 6024 2851
rect 6084 2774 6144 3804
rect 6204 2834 6264 3866
rect 6324 2774 6384 3804
rect 6444 2834 6504 3866
rect 6564 3712 6630 3866
rect 6564 3648 6565 3712
rect 6629 3648 6630 3712
rect 6564 3632 6630 3648
rect 6564 3568 6565 3632
rect 6629 3568 6630 3632
rect 6564 3552 6630 3568
rect 6564 3488 6565 3552
rect 6629 3488 6630 3552
rect 6564 3472 6630 3488
rect 6564 3408 6565 3472
rect 6629 3408 6630 3472
rect 6564 3392 6630 3408
rect 6564 3328 6565 3392
rect 6629 3328 6630 3392
rect 6564 3312 6630 3328
rect 6564 3248 6565 3312
rect 6629 3248 6630 3312
rect 6564 3232 6630 3248
rect 6564 3168 6565 3232
rect 6629 3168 6630 3232
rect 6564 3152 6630 3168
rect 6564 3088 6565 3152
rect 6629 3088 6630 3152
rect 6564 3072 6630 3088
rect 6564 3008 6565 3072
rect 6629 3008 6630 3072
rect 6564 2992 6630 3008
rect 6564 2928 6565 2992
rect 6629 2928 6630 2992
rect 6564 2907 6630 2928
rect 6564 2851 6569 2907
rect 6625 2851 6630 2907
rect 6564 2838 6630 2851
rect 6690 2774 6750 3804
rect 6810 2834 6870 3866
rect 6930 2774 6990 3804
rect 7050 2834 7110 3866
rect 7170 3712 7236 3866
rect 7170 3648 7171 3712
rect 7235 3648 7236 3712
rect 7170 3632 7236 3648
rect 7170 3568 7171 3632
rect 7235 3568 7236 3632
rect 7170 3552 7236 3568
rect 7170 3488 7171 3552
rect 7235 3488 7236 3552
rect 7170 3472 7236 3488
rect 7170 3408 7171 3472
rect 7235 3408 7236 3472
rect 7170 3392 7236 3408
rect 7170 3328 7171 3392
rect 7235 3328 7236 3392
rect 7170 3312 7236 3328
rect 7170 3248 7171 3312
rect 7235 3248 7236 3312
rect 7170 3232 7236 3248
rect 7170 3168 7171 3232
rect 7235 3168 7236 3232
rect 7170 3152 7236 3168
rect 7170 3088 7171 3152
rect 7235 3088 7236 3152
rect 7170 3072 7236 3088
rect 7170 3008 7171 3072
rect 7235 3008 7236 3072
rect 7170 2992 7236 3008
rect 7170 2928 7171 2992
rect 7235 2928 7236 2992
rect 7170 2907 7236 2928
rect 7170 2851 7175 2907
rect 7231 2851 7236 2907
rect 7170 2838 7236 2851
rect 7296 2774 7356 3804
rect 7416 2834 7476 3866
rect 7536 2774 7596 3804
rect 7656 2834 7716 3866
rect 7776 3712 7842 3866
rect 7776 3648 7777 3712
rect 7841 3648 7842 3712
rect 7776 3632 7842 3648
rect 7776 3568 7777 3632
rect 7841 3568 7842 3632
rect 7776 3552 7842 3568
rect 7776 3488 7777 3552
rect 7841 3488 7842 3552
rect 7776 3472 7842 3488
rect 7776 3408 7777 3472
rect 7841 3408 7842 3472
rect 7776 3392 7842 3408
rect 7776 3328 7777 3392
rect 7841 3328 7842 3392
rect 7776 3312 7842 3328
rect 7776 3248 7777 3312
rect 7841 3248 7842 3312
rect 7776 3232 7842 3248
rect 7776 3168 7777 3232
rect 7841 3168 7842 3232
rect 7776 3152 7842 3168
rect 7776 3088 7777 3152
rect 7841 3088 7842 3152
rect 7776 3072 7842 3088
rect 7776 3008 7777 3072
rect 7841 3008 7842 3072
rect 7776 2992 7842 3008
rect 7776 2928 7777 2992
rect 7841 2928 7842 2992
rect 7776 2907 7842 2928
rect 7776 2851 7781 2907
rect 7837 2851 7842 2907
rect 7776 2838 7842 2851
rect 7902 2774 7962 3804
rect 8022 2834 8082 3866
rect 8142 2774 8202 3804
rect 8262 2834 8322 3866
rect 8382 3712 8448 3866
rect 8382 3648 8383 3712
rect 8447 3648 8448 3712
rect 8382 3632 8448 3648
rect 8382 3568 8383 3632
rect 8447 3568 8448 3632
rect 8382 3552 8448 3568
rect 8382 3488 8383 3552
rect 8447 3488 8448 3552
rect 8382 3472 8448 3488
rect 8382 3408 8383 3472
rect 8447 3408 8448 3472
rect 8382 3392 8448 3408
rect 8382 3328 8383 3392
rect 8447 3328 8448 3392
rect 8382 3312 8448 3328
rect 8382 3248 8383 3312
rect 8447 3248 8448 3312
rect 8382 3232 8448 3248
rect 8382 3168 8383 3232
rect 8447 3168 8448 3232
rect 8382 3152 8448 3168
rect 8382 3088 8383 3152
rect 8447 3088 8448 3152
rect 8382 3072 8448 3088
rect 8382 3008 8383 3072
rect 8447 3008 8448 3072
rect 8382 2992 8448 3008
rect 8382 2928 8383 2992
rect 8447 2928 8448 2992
rect 8382 2838 8448 2928
rect 8508 2774 8568 3804
rect 8628 2834 8688 3866
rect 8748 2774 8808 3804
rect 8868 2834 8928 3866
rect 8988 3712 9054 3866
rect 8988 3648 8989 3712
rect 9053 3648 9054 3712
rect 8988 3632 9054 3648
rect 8988 3568 8989 3632
rect 9053 3568 9054 3632
rect 8988 3552 9054 3568
rect 8988 3488 8989 3552
rect 9053 3488 9054 3552
rect 8988 3472 9054 3488
rect 8988 3408 8989 3472
rect 9053 3408 9054 3472
rect 8988 3392 9054 3408
rect 8988 3328 8989 3392
rect 9053 3328 9054 3392
rect 8988 3312 9054 3328
rect 8988 3248 8989 3312
rect 9053 3248 9054 3312
rect 8988 3232 9054 3248
rect 8988 3168 8989 3232
rect 9053 3168 9054 3232
rect 8988 3152 9054 3168
rect 8988 3088 8989 3152
rect 9053 3088 9054 3152
rect 8988 3072 9054 3088
rect 8988 3008 8989 3072
rect 9053 3008 9054 3072
rect 8988 2992 9054 3008
rect 8988 2928 8989 2992
rect 9053 2928 9054 2992
rect 8988 2838 9054 2928
rect 9114 2774 9174 3804
rect 9234 2834 9294 3866
rect 9354 2774 9414 3804
rect 9474 2834 9534 3866
rect 9594 3712 9660 3866
rect 9594 3648 9595 3712
rect 9659 3648 9660 3712
rect 9594 3632 9660 3648
rect 9594 3568 9595 3632
rect 9659 3568 9660 3632
rect 9594 3552 9660 3568
rect 9594 3488 9595 3552
rect 9659 3488 9660 3552
rect 9594 3472 9660 3488
rect 9594 3408 9595 3472
rect 9659 3408 9660 3472
rect 9594 3392 9660 3408
rect 9594 3328 9595 3392
rect 9659 3328 9660 3392
rect 9594 3312 9660 3328
rect 9594 3248 9595 3312
rect 9659 3248 9660 3312
rect 9594 3232 9660 3248
rect 9594 3168 9595 3232
rect 9659 3168 9660 3232
rect 9594 3152 9660 3168
rect 9594 3088 9595 3152
rect 9659 3088 9660 3152
rect 9594 3072 9660 3088
rect 9594 3008 9595 3072
rect 9659 3008 9660 3072
rect 9594 2992 9660 3008
rect 9594 2928 9595 2992
rect 9659 2928 9660 2992
rect 9594 2838 9660 2928
rect 9720 2774 9780 3804
rect 9840 2834 9900 3866
rect 9960 2774 10020 3804
rect 10080 2834 10140 3866
rect 10200 3712 10266 3866
rect 10200 3648 10201 3712
rect 10265 3648 10266 3712
rect 10200 3632 10266 3648
rect 10200 3568 10201 3632
rect 10265 3568 10266 3632
rect 10200 3552 10266 3568
rect 10200 3488 10201 3552
rect 10265 3488 10266 3552
rect 10200 3472 10266 3488
rect 10200 3408 10201 3472
rect 10265 3408 10266 3472
rect 10200 3392 10266 3408
rect 10200 3328 10201 3392
rect 10265 3328 10266 3392
rect 10200 3312 10266 3328
rect 10200 3248 10201 3312
rect 10265 3248 10266 3312
rect 10200 3232 10266 3248
rect 10200 3168 10201 3232
rect 10265 3168 10266 3232
rect 10200 3152 10266 3168
rect 10200 3088 10201 3152
rect 10265 3088 10266 3152
rect 10200 3072 10266 3088
rect 10200 3008 10201 3072
rect 10265 3008 10266 3072
rect 10200 2992 10266 3008
rect 10200 2928 10201 2992
rect 10265 2928 10266 2992
rect 10200 2838 10266 2928
rect 10326 4872 10392 4962
rect 10326 4808 10327 4872
rect 10391 4808 10392 4872
rect 10326 4792 10392 4808
rect 10326 4728 10327 4792
rect 10391 4728 10392 4792
rect 10326 4712 10392 4728
rect 10326 4648 10327 4712
rect 10391 4648 10392 4712
rect 10326 4632 10392 4648
rect 10326 4568 10327 4632
rect 10391 4568 10392 4632
rect 10326 4552 10392 4568
rect 10326 4488 10327 4552
rect 10391 4488 10392 4552
rect 10326 4472 10392 4488
rect 10326 4408 10327 4472
rect 10391 4408 10392 4472
rect 10326 4392 10392 4408
rect 10326 4328 10327 4392
rect 10391 4328 10392 4392
rect 10326 4312 10392 4328
rect 10326 4248 10327 4312
rect 10391 4248 10392 4312
rect 10326 4232 10392 4248
rect 10326 4168 10327 4232
rect 10391 4168 10392 4232
rect 10326 4152 10392 4168
rect 10326 4088 10327 4152
rect 10391 4088 10392 4152
rect 10326 3934 10392 4088
rect 10452 3934 10512 4966
rect 10572 3996 10632 5026
rect 10692 3934 10752 4966
rect 10812 3996 10872 5026
rect 10932 4872 10998 4962
rect 10932 4808 10933 4872
rect 10997 4808 10998 4872
rect 10932 4792 10998 4808
rect 10932 4728 10933 4792
rect 10997 4728 10998 4792
rect 10932 4712 10998 4728
rect 10932 4648 10933 4712
rect 10997 4648 10998 4712
rect 10932 4632 10998 4648
rect 10932 4568 10933 4632
rect 10997 4568 10998 4632
rect 10932 4552 10998 4568
rect 10932 4488 10933 4552
rect 10997 4488 10998 4552
rect 10932 4472 10998 4488
rect 10932 4408 10933 4472
rect 10997 4408 10998 4472
rect 10932 4392 10998 4408
rect 10932 4328 10933 4392
rect 10997 4328 10998 4392
rect 10932 4312 10998 4328
rect 10932 4248 10933 4312
rect 10997 4248 10998 4312
rect 10932 4232 10998 4248
rect 10932 4168 10933 4232
rect 10997 4168 10998 4232
rect 10932 4152 10998 4168
rect 10932 4088 10933 4152
rect 10997 4088 10998 4152
rect 10932 3934 10998 4088
rect 11058 3934 11118 4966
rect 11178 3996 11238 5026
rect 11298 3934 11358 4966
rect 11418 3996 11478 5026
rect 11538 4872 11604 4962
rect 11538 4808 11539 4872
rect 11603 4808 11604 4872
rect 11538 4792 11604 4808
rect 11538 4728 11539 4792
rect 11603 4728 11604 4792
rect 11538 4712 11604 4728
rect 11538 4648 11539 4712
rect 11603 4648 11604 4712
rect 11538 4632 11604 4648
rect 11538 4568 11539 4632
rect 11603 4568 11604 4632
rect 11538 4552 11604 4568
rect 11538 4488 11539 4552
rect 11603 4488 11604 4552
rect 11538 4472 11604 4488
rect 11538 4408 11539 4472
rect 11603 4408 11604 4472
rect 11538 4392 11604 4408
rect 11538 4328 11539 4392
rect 11603 4328 11604 4392
rect 11538 4312 11604 4328
rect 11538 4248 11539 4312
rect 11603 4248 11604 4312
rect 11538 4232 11604 4248
rect 11538 4168 11539 4232
rect 11603 4168 11604 4232
rect 11538 4152 11604 4168
rect 11538 4088 11539 4152
rect 11603 4088 11604 4152
rect 11538 3934 11604 4088
rect 11664 3934 11724 4966
rect 11784 3996 11844 5026
rect 11904 3934 11964 4966
rect 12024 3996 12084 5026
rect 12144 4872 12210 4962
rect 12144 4808 12145 4872
rect 12209 4808 12210 4872
rect 12144 4792 12210 4808
rect 12144 4728 12145 4792
rect 12209 4728 12210 4792
rect 12144 4712 12210 4728
rect 12144 4648 12145 4712
rect 12209 4648 12210 4712
rect 12144 4632 12210 4648
rect 12144 4568 12145 4632
rect 12209 4568 12210 4632
rect 12144 4552 12210 4568
rect 12144 4488 12145 4552
rect 12209 4488 12210 4552
rect 12144 4472 12210 4488
rect 12144 4408 12145 4472
rect 12209 4408 12210 4472
rect 12144 4392 12210 4408
rect 12144 4328 12145 4392
rect 12209 4328 12210 4392
rect 12144 4312 12210 4328
rect 12144 4248 12145 4312
rect 12209 4248 12210 4312
rect 12144 4232 12210 4248
rect 12144 4168 12145 4232
rect 12209 4168 12210 4232
rect 12144 4152 12210 4168
rect 12144 4088 12145 4152
rect 12209 4088 12210 4152
rect 12144 3934 12210 4088
rect 12270 3934 12330 4966
rect 12390 3996 12450 5026
rect 12510 3934 12570 4966
rect 12630 3996 12690 5026
rect 12750 4872 12816 4962
rect 12750 4808 12751 4872
rect 12815 4808 12816 4872
rect 12750 4792 12816 4808
rect 12750 4728 12751 4792
rect 12815 4728 12816 4792
rect 12750 4712 12816 4728
rect 12750 4648 12751 4712
rect 12815 4648 12816 4712
rect 12750 4632 12816 4648
rect 12750 4568 12751 4632
rect 12815 4568 12816 4632
rect 12750 4552 12816 4568
rect 12750 4488 12751 4552
rect 12815 4488 12816 4552
rect 12750 4472 12816 4488
rect 12750 4408 12751 4472
rect 12815 4408 12816 4472
rect 12750 4392 12816 4408
rect 12750 4328 12751 4392
rect 12815 4328 12816 4392
rect 12750 4312 12816 4328
rect 12750 4248 12751 4312
rect 12815 4248 12816 4312
rect 12750 4232 12816 4248
rect 12750 4168 12751 4232
rect 12815 4168 12816 4232
rect 12750 4152 12816 4168
rect 12750 4088 12751 4152
rect 12815 4088 12816 4152
rect 12750 3934 12816 4088
rect 12876 3934 12936 4966
rect 12996 3996 13056 5026
rect 13116 3934 13176 4966
rect 13236 3996 13296 5026
rect 13356 4872 13422 4962
rect 13356 4808 13357 4872
rect 13421 4808 13422 4872
rect 13356 4792 13422 4808
rect 13356 4728 13357 4792
rect 13421 4728 13422 4792
rect 13356 4712 13422 4728
rect 13356 4648 13357 4712
rect 13421 4648 13422 4712
rect 13356 4632 13422 4648
rect 13356 4568 13357 4632
rect 13421 4568 13422 4632
rect 13356 4552 13422 4568
rect 13356 4488 13357 4552
rect 13421 4488 13422 4552
rect 13356 4472 13422 4488
rect 13356 4408 13357 4472
rect 13421 4408 13422 4472
rect 13356 4392 13422 4408
rect 13356 4328 13357 4392
rect 13421 4328 13422 4392
rect 13356 4312 13422 4328
rect 13356 4248 13357 4312
rect 13421 4248 13422 4312
rect 13356 4232 13422 4248
rect 13356 4168 13357 4232
rect 13421 4168 13422 4232
rect 13356 4152 13422 4168
rect 13356 4088 13357 4152
rect 13421 4088 13422 4152
rect 13356 3934 13422 4088
rect 13482 3934 13542 4966
rect 13602 3996 13662 5026
rect 13722 3934 13782 4966
rect 13842 3996 13902 5026
rect 13962 4872 14028 4962
rect 13962 4808 13963 4872
rect 14027 4808 14028 4872
rect 13962 4792 14028 4808
rect 13962 4728 13963 4792
rect 14027 4728 14028 4792
rect 13962 4712 14028 4728
rect 13962 4648 13963 4712
rect 14027 4648 14028 4712
rect 13962 4632 14028 4648
rect 13962 4568 13963 4632
rect 14027 4568 14028 4632
rect 13962 4552 14028 4568
rect 13962 4488 13963 4552
rect 14027 4488 14028 4552
rect 13962 4472 14028 4488
rect 13962 4408 13963 4472
rect 14027 4408 14028 4472
rect 13962 4392 14028 4408
rect 13962 4328 13963 4392
rect 14027 4328 14028 4392
rect 13962 4312 14028 4328
rect 13962 4248 13963 4312
rect 14027 4248 14028 4312
rect 13962 4232 14028 4248
rect 13962 4168 13963 4232
rect 14027 4168 14028 4232
rect 13962 4152 14028 4168
rect 13962 4088 13963 4152
rect 14027 4088 14028 4152
rect 13962 3934 14028 4088
rect 14088 3934 14148 4966
rect 14208 3996 14268 5026
rect 14328 3934 14388 4966
rect 14448 3996 14508 5026
rect 14568 4872 14634 4962
rect 14568 4808 14569 4872
rect 14633 4808 14634 4872
rect 14568 4792 14634 4808
rect 14568 4728 14569 4792
rect 14633 4728 14634 4792
rect 14568 4712 14634 4728
rect 14568 4648 14569 4712
rect 14633 4648 14634 4712
rect 14568 4632 14634 4648
rect 14568 4568 14569 4632
rect 14633 4568 14634 4632
rect 14568 4552 14634 4568
rect 14568 4488 14569 4552
rect 14633 4488 14634 4552
rect 14568 4472 14634 4488
rect 14568 4408 14569 4472
rect 14633 4408 14634 4472
rect 14568 4392 14634 4408
rect 14568 4328 14569 4392
rect 14633 4328 14634 4392
rect 14568 4312 14634 4328
rect 14568 4248 14569 4312
rect 14633 4248 14634 4312
rect 14568 4232 14634 4248
rect 14568 4168 14569 4232
rect 14633 4168 14634 4232
rect 14568 4152 14634 4168
rect 14568 4088 14569 4152
rect 14633 4088 14634 4152
rect 14568 3934 14634 4088
rect 14694 3934 14754 4966
rect 14814 3996 14874 5026
rect 14934 3934 14994 4966
rect 15054 3996 15114 5026
rect 15174 4872 15240 4962
rect 15174 4808 15175 4872
rect 15239 4808 15240 4872
rect 15174 4792 15240 4808
rect 15174 4728 15175 4792
rect 15239 4728 15240 4792
rect 15174 4712 15240 4728
rect 15174 4648 15175 4712
rect 15239 4648 15240 4712
rect 15174 4632 15240 4648
rect 15174 4568 15175 4632
rect 15239 4568 15240 4632
rect 15174 4552 15240 4568
rect 15174 4488 15175 4552
rect 15239 4488 15240 4552
rect 15174 4472 15240 4488
rect 15174 4408 15175 4472
rect 15239 4408 15240 4472
rect 15174 4392 15240 4408
rect 15174 4328 15175 4392
rect 15239 4328 15240 4392
rect 15174 4312 15240 4328
rect 15174 4248 15175 4312
rect 15239 4248 15240 4312
rect 15174 4232 15240 4248
rect 15174 4168 15175 4232
rect 15239 4168 15240 4232
rect 15174 4152 15240 4168
rect 15174 4088 15175 4152
rect 15239 4088 15240 4152
rect 15174 3934 15240 4088
rect 15300 3934 15360 4966
rect 15420 3996 15480 5026
rect 15540 3934 15600 4966
rect 15660 3996 15720 5026
rect 15780 4872 15846 4962
rect 15780 4808 15781 4872
rect 15845 4808 15846 4872
rect 15780 4792 15846 4808
rect 15780 4728 15781 4792
rect 15845 4728 15846 4792
rect 15780 4712 15846 4728
rect 15780 4648 15781 4712
rect 15845 4648 15846 4712
rect 15780 4632 15846 4648
rect 15780 4568 15781 4632
rect 15845 4568 15846 4632
rect 15780 4552 15846 4568
rect 15780 4488 15781 4552
rect 15845 4488 15846 4552
rect 15780 4472 15846 4488
rect 15780 4408 15781 4472
rect 15845 4408 15846 4472
rect 15780 4392 15846 4408
rect 15780 4328 15781 4392
rect 15845 4328 15846 4392
rect 15780 4312 15846 4328
rect 15780 4248 15781 4312
rect 15845 4248 15846 4312
rect 15780 4232 15846 4248
rect 15780 4168 15781 4232
rect 15845 4168 15846 4232
rect 15780 4152 15846 4168
rect 15780 4088 15781 4152
rect 15845 4088 15846 4152
rect 15780 3934 15846 4088
rect 15906 3934 15966 4966
rect 16026 3996 16086 5026
rect 16146 3934 16206 4966
rect 16266 3996 16326 5026
rect 16386 4872 16452 4962
rect 16386 4808 16387 4872
rect 16451 4808 16452 4872
rect 16386 4792 16452 4808
rect 16386 4728 16387 4792
rect 16451 4728 16452 4792
rect 16386 4712 16452 4728
rect 16386 4648 16387 4712
rect 16451 4648 16452 4712
rect 16386 4632 16452 4648
rect 16386 4568 16387 4632
rect 16451 4568 16452 4632
rect 16386 4552 16452 4568
rect 16386 4488 16387 4552
rect 16451 4488 16452 4552
rect 16386 4472 16452 4488
rect 16386 4408 16387 4472
rect 16451 4408 16452 4472
rect 16386 4392 16452 4408
rect 16386 4328 16387 4392
rect 16451 4328 16452 4392
rect 16386 4312 16452 4328
rect 16386 4248 16387 4312
rect 16451 4248 16452 4312
rect 16386 4232 16452 4248
rect 16386 4168 16387 4232
rect 16451 4168 16452 4232
rect 16386 4152 16452 4168
rect 16386 4088 16387 4152
rect 16451 4088 16452 4152
rect 16386 3934 16452 4088
rect 16512 3934 16572 4966
rect 16632 3996 16692 5026
rect 16752 3934 16812 4966
rect 16872 3996 16932 5026
rect 16992 4872 17058 4962
rect 16992 4808 16993 4872
rect 17057 4808 17058 4872
rect 16992 4792 17058 4808
rect 16992 4728 16993 4792
rect 17057 4728 17058 4792
rect 16992 4712 17058 4728
rect 16992 4648 16993 4712
rect 17057 4648 17058 4712
rect 16992 4632 17058 4648
rect 16992 4568 16993 4632
rect 17057 4568 17058 4632
rect 16992 4552 17058 4568
rect 16992 4488 16993 4552
rect 17057 4488 17058 4552
rect 16992 4472 17058 4488
rect 16992 4408 16993 4472
rect 17057 4408 17058 4472
rect 16992 4392 17058 4408
rect 16992 4328 16993 4392
rect 17057 4328 17058 4392
rect 16992 4312 17058 4328
rect 16992 4248 16993 4312
rect 17057 4248 17058 4312
rect 16992 4232 17058 4248
rect 16992 4168 16993 4232
rect 17057 4168 17058 4232
rect 16992 4152 17058 4168
rect 16992 4088 16993 4152
rect 17057 4088 17058 4152
rect 16992 3934 17058 4088
rect 17118 3934 17178 4966
rect 17238 3996 17298 5026
rect 17358 3934 17418 4966
rect 17478 3996 17538 5026
rect 17598 4872 17664 4962
rect 17598 4808 17599 4872
rect 17663 4808 17664 4872
rect 17598 4792 17664 4808
rect 17598 4728 17599 4792
rect 17663 4728 17664 4792
rect 17598 4712 17664 4728
rect 17598 4648 17599 4712
rect 17663 4648 17664 4712
rect 17598 4632 17664 4648
rect 17598 4568 17599 4632
rect 17663 4568 17664 4632
rect 17598 4552 17664 4568
rect 17598 4488 17599 4552
rect 17663 4488 17664 4552
rect 17598 4472 17664 4488
rect 17598 4408 17599 4472
rect 17663 4408 17664 4472
rect 17598 4392 17664 4408
rect 17598 4328 17599 4392
rect 17663 4328 17664 4392
rect 17598 4312 17664 4328
rect 17598 4248 17599 4312
rect 17663 4248 17664 4312
rect 17598 4232 17664 4248
rect 17598 4168 17599 4232
rect 17663 4168 17664 4232
rect 17598 4152 17664 4168
rect 17598 4088 17599 4152
rect 17663 4088 17664 4152
rect 17598 3934 17664 4088
rect 17724 3934 17784 4966
rect 17844 3996 17904 5026
rect 17964 3934 18024 4966
rect 18084 3996 18144 5026
rect 18204 4872 18270 4962
rect 18204 4808 18205 4872
rect 18269 4808 18270 4872
rect 18204 4792 18270 4808
rect 18204 4728 18205 4792
rect 18269 4728 18270 4792
rect 18204 4712 18270 4728
rect 18204 4648 18205 4712
rect 18269 4648 18270 4712
rect 18204 4632 18270 4648
rect 18204 4568 18205 4632
rect 18269 4568 18270 4632
rect 18204 4552 18270 4568
rect 18204 4488 18205 4552
rect 18269 4488 18270 4552
rect 18204 4472 18270 4488
rect 18204 4408 18205 4472
rect 18269 4408 18270 4472
rect 18204 4392 18270 4408
rect 18204 4328 18205 4392
rect 18269 4328 18270 4392
rect 18204 4312 18270 4328
rect 18204 4248 18205 4312
rect 18269 4248 18270 4312
rect 18204 4232 18270 4248
rect 18204 4168 18205 4232
rect 18269 4168 18270 4232
rect 18204 4152 18270 4168
rect 18204 4088 18205 4152
rect 18269 4088 18270 4152
rect 18204 3934 18270 4088
rect 18330 3934 18390 4966
rect 18450 3996 18510 5026
rect 18570 3934 18630 4966
rect 18690 3996 18750 5026
rect 18810 4872 18876 4962
rect 18810 4808 18811 4872
rect 18875 4808 18876 4872
rect 18810 4792 18876 4808
rect 18810 4728 18811 4792
rect 18875 4728 18876 4792
rect 18810 4712 18876 4728
rect 18810 4648 18811 4712
rect 18875 4648 18876 4712
rect 18810 4632 18876 4648
rect 18810 4568 18811 4632
rect 18875 4568 18876 4632
rect 18810 4552 18876 4568
rect 18810 4488 18811 4552
rect 18875 4488 18876 4552
rect 18810 4472 18876 4488
rect 18810 4408 18811 4472
rect 18875 4408 18876 4472
rect 18810 4392 18876 4408
rect 18810 4328 18811 4392
rect 18875 4328 18876 4392
rect 18810 4312 18876 4328
rect 18810 4248 18811 4312
rect 18875 4248 18876 4312
rect 18810 4232 18876 4248
rect 18810 4168 18811 4232
rect 18875 4168 18876 4232
rect 18810 4152 18876 4168
rect 18810 4088 18811 4152
rect 18875 4088 18876 4152
rect 18810 3934 18876 4088
rect 18936 3934 18996 4966
rect 19056 3996 19116 5026
rect 19176 3934 19236 4966
rect 19296 3996 19356 5026
rect 19416 4872 19482 4962
rect 19416 4808 19417 4872
rect 19481 4808 19482 4872
rect 19416 4792 19482 4808
rect 19416 4728 19417 4792
rect 19481 4728 19482 4792
rect 19416 4712 19482 4728
rect 19416 4648 19417 4712
rect 19481 4648 19482 4712
rect 19416 4632 19482 4648
rect 19416 4568 19417 4632
rect 19481 4568 19482 4632
rect 19416 4552 19482 4568
rect 19416 4488 19417 4552
rect 19481 4488 19482 4552
rect 19416 4472 19482 4488
rect 19416 4408 19417 4472
rect 19481 4408 19482 4472
rect 19416 4392 19482 4408
rect 19416 4328 19417 4392
rect 19481 4328 19482 4392
rect 19416 4312 19482 4328
rect 19416 4248 19417 4312
rect 19481 4248 19482 4312
rect 19416 4232 19482 4248
rect 19416 4168 19417 4232
rect 19481 4168 19482 4232
rect 19416 4152 19482 4168
rect 19416 4088 19417 4152
rect 19481 4088 19482 4152
rect 19416 3934 19482 4088
rect 19542 3934 19602 4966
rect 19662 3996 19722 5026
rect 19782 3934 19842 4966
rect 19902 3996 19962 5026
rect 20022 4872 20088 4962
rect 20022 4808 20023 4872
rect 20087 4808 20088 4872
rect 20022 4792 20088 4808
rect 20022 4728 20023 4792
rect 20087 4728 20088 4792
rect 20022 4712 20088 4728
rect 20022 4648 20023 4712
rect 20087 4648 20088 4712
rect 20022 4632 20088 4648
rect 20022 4568 20023 4632
rect 20087 4568 20088 4632
rect 20022 4552 20088 4568
rect 20022 4488 20023 4552
rect 20087 4488 20088 4552
rect 20022 4472 20088 4488
rect 20022 4408 20023 4472
rect 20087 4408 20088 4472
rect 20022 4392 20088 4408
rect 20022 4328 20023 4392
rect 20087 4328 20088 4392
rect 20022 4312 20088 4328
rect 20022 4248 20023 4312
rect 20087 4248 20088 4312
rect 20022 4232 20088 4248
rect 20022 4168 20023 4232
rect 20087 4168 20088 4232
rect 20022 4152 20088 4168
rect 20022 4088 20023 4152
rect 20087 4088 20088 4152
rect 20022 3934 20088 4088
rect 10326 3932 20088 3934
rect 10326 3868 10430 3932
rect 10494 3868 10510 3932
rect 10574 3868 10590 3932
rect 10654 3868 10670 3932
rect 10734 3868 10750 3932
rect 10814 3868 10830 3932
rect 10894 3868 11036 3932
rect 11100 3868 11116 3932
rect 11180 3868 11196 3932
rect 11260 3868 11276 3932
rect 11340 3868 11356 3932
rect 11420 3868 11436 3932
rect 11500 3868 11642 3932
rect 11706 3868 11722 3932
rect 11786 3868 11802 3932
rect 11866 3868 11882 3932
rect 11946 3868 11962 3932
rect 12026 3868 12042 3932
rect 12106 3868 12248 3932
rect 12312 3868 12328 3932
rect 12392 3868 12408 3932
rect 12472 3868 12488 3932
rect 12552 3868 12568 3932
rect 12632 3868 12648 3932
rect 12712 3868 12854 3932
rect 12918 3868 12934 3932
rect 12998 3868 13014 3932
rect 13078 3868 13094 3932
rect 13158 3868 13174 3932
rect 13238 3868 13254 3932
rect 13318 3868 13460 3932
rect 13524 3868 13540 3932
rect 13604 3868 13620 3932
rect 13684 3868 13700 3932
rect 13764 3868 13780 3932
rect 13844 3868 13860 3932
rect 13924 3868 14066 3932
rect 14130 3868 14146 3932
rect 14210 3868 14226 3932
rect 14290 3868 14306 3932
rect 14370 3868 14386 3932
rect 14450 3868 14466 3932
rect 14530 3868 14672 3932
rect 14736 3868 14752 3932
rect 14816 3868 14832 3932
rect 14896 3868 14912 3932
rect 14976 3868 14992 3932
rect 15056 3868 15072 3932
rect 15136 3868 15278 3932
rect 15342 3868 15358 3932
rect 15422 3868 15438 3932
rect 15502 3868 15518 3932
rect 15582 3868 15598 3932
rect 15662 3868 15678 3932
rect 15742 3868 15884 3932
rect 15948 3868 15964 3932
rect 16028 3868 16044 3932
rect 16108 3868 16124 3932
rect 16188 3868 16204 3932
rect 16268 3868 16284 3932
rect 16348 3868 16490 3932
rect 16554 3868 16570 3932
rect 16634 3868 16650 3932
rect 16714 3868 16730 3932
rect 16794 3868 16810 3932
rect 16874 3868 16890 3932
rect 16954 3868 17096 3932
rect 17160 3868 17176 3932
rect 17240 3868 17256 3932
rect 17320 3868 17336 3932
rect 17400 3868 17416 3932
rect 17480 3868 17496 3932
rect 17560 3868 17702 3932
rect 17766 3868 17782 3932
rect 17846 3868 17862 3932
rect 17926 3868 17942 3932
rect 18006 3868 18022 3932
rect 18086 3868 18102 3932
rect 18166 3868 18308 3932
rect 18372 3868 18388 3932
rect 18452 3868 18468 3932
rect 18532 3868 18548 3932
rect 18612 3868 18628 3932
rect 18692 3868 18708 3932
rect 18772 3868 18914 3932
rect 18978 3868 18994 3932
rect 19058 3868 19074 3932
rect 19138 3868 19154 3932
rect 19218 3868 19234 3932
rect 19298 3868 19314 3932
rect 19378 3868 19520 3932
rect 19584 3868 19600 3932
rect 19664 3868 19680 3932
rect 19744 3868 19760 3932
rect 19824 3868 19840 3932
rect 19904 3868 19920 3932
rect 19984 3868 20088 3932
rect 10326 3866 20088 3868
rect 10326 3712 10392 3866
rect 10326 3648 10327 3712
rect 10391 3648 10392 3712
rect 10326 3632 10392 3648
rect 10326 3568 10327 3632
rect 10391 3568 10392 3632
rect 10326 3552 10392 3568
rect 10326 3488 10327 3552
rect 10391 3488 10392 3552
rect 10326 3472 10392 3488
rect 10326 3408 10327 3472
rect 10391 3408 10392 3472
rect 10326 3392 10392 3408
rect 10326 3328 10327 3392
rect 10391 3328 10392 3392
rect 10326 3312 10392 3328
rect 10326 3248 10327 3312
rect 10391 3248 10392 3312
rect 10326 3232 10392 3248
rect 10326 3168 10327 3232
rect 10391 3168 10392 3232
rect 10326 3152 10392 3168
rect 10326 3088 10327 3152
rect 10391 3088 10392 3152
rect 10326 3072 10392 3088
rect 10326 3008 10327 3072
rect 10391 3008 10392 3072
rect 10326 2992 10392 3008
rect 10326 2928 10327 2992
rect 10391 2928 10392 2992
rect 10326 2912 10392 2928
rect 10326 2856 10331 2912
rect 10387 2856 10392 2912
rect 10326 2838 10392 2856
rect 10452 2774 10512 3804
rect 10572 2834 10632 3866
rect 10692 2774 10752 3804
rect 10812 2834 10872 3866
rect 10932 3712 10998 3866
rect 10932 3648 10933 3712
rect 10997 3648 10998 3712
rect 10932 3632 10998 3648
rect 10932 3568 10933 3632
rect 10997 3568 10998 3632
rect 10932 3552 10998 3568
rect 10932 3488 10933 3552
rect 10997 3488 10998 3552
rect 10932 3472 10998 3488
rect 10932 3408 10933 3472
rect 10997 3408 10998 3472
rect 10932 3392 10998 3408
rect 10932 3328 10933 3392
rect 10997 3328 10998 3392
rect 10932 3312 10998 3328
rect 10932 3248 10933 3312
rect 10997 3248 10998 3312
rect 10932 3232 10998 3248
rect 10932 3168 10933 3232
rect 10997 3168 10998 3232
rect 10932 3152 10998 3168
rect 10932 3088 10933 3152
rect 10997 3088 10998 3152
rect 10932 3072 10998 3088
rect 10932 3008 10933 3072
rect 10997 3008 10998 3072
rect 10932 2992 10998 3008
rect 10932 2928 10933 2992
rect 10997 2928 10998 2992
rect 10932 2903 10998 2928
rect 10932 2847 10937 2903
rect 10993 2847 10998 2903
rect 10932 2838 10998 2847
rect 11058 2774 11118 3804
rect 11178 2834 11238 3866
rect 11298 2774 11358 3804
rect 11418 2834 11478 3866
rect 11538 3712 11604 3866
rect 11538 3648 11539 3712
rect 11603 3648 11604 3712
rect 11538 3632 11604 3648
rect 11538 3568 11539 3632
rect 11603 3568 11604 3632
rect 11538 3552 11604 3568
rect 11538 3488 11539 3552
rect 11603 3488 11604 3552
rect 11538 3472 11604 3488
rect 11538 3408 11539 3472
rect 11603 3408 11604 3472
rect 11538 3392 11604 3408
rect 11538 3328 11539 3392
rect 11603 3328 11604 3392
rect 11538 3312 11604 3328
rect 11538 3248 11539 3312
rect 11603 3248 11604 3312
rect 11538 3232 11604 3248
rect 11538 3168 11539 3232
rect 11603 3168 11604 3232
rect 11538 3152 11604 3168
rect 11538 3088 11539 3152
rect 11603 3088 11604 3152
rect 11538 3072 11604 3088
rect 11538 3008 11539 3072
rect 11603 3008 11604 3072
rect 11538 2992 11604 3008
rect 11538 2928 11539 2992
rect 11603 2928 11604 2992
rect 11538 2904 11604 2928
rect 11538 2848 11543 2904
rect 11599 2848 11604 2904
rect 11538 2838 11604 2848
rect 11664 2774 11724 3804
rect 11784 2834 11844 3866
rect 11904 2774 11964 3804
rect 12024 2834 12084 3866
rect 12144 3712 12210 3866
rect 12144 3648 12145 3712
rect 12209 3648 12210 3712
rect 12144 3632 12210 3648
rect 12144 3568 12145 3632
rect 12209 3568 12210 3632
rect 12144 3552 12210 3568
rect 12144 3488 12145 3552
rect 12209 3488 12210 3552
rect 12144 3472 12210 3488
rect 12144 3408 12145 3472
rect 12209 3408 12210 3472
rect 12144 3392 12210 3408
rect 12144 3328 12145 3392
rect 12209 3328 12210 3392
rect 12144 3312 12210 3328
rect 12144 3248 12145 3312
rect 12209 3248 12210 3312
rect 12144 3232 12210 3248
rect 12144 3168 12145 3232
rect 12209 3168 12210 3232
rect 12144 3152 12210 3168
rect 12144 3088 12145 3152
rect 12209 3088 12210 3152
rect 12144 3072 12210 3088
rect 12144 3008 12145 3072
rect 12209 3008 12210 3072
rect 12144 2992 12210 3008
rect 12144 2928 12145 2992
rect 12209 2928 12210 2992
rect 12144 2903 12210 2928
rect 12144 2847 12149 2903
rect 12205 2847 12210 2903
rect 12144 2838 12210 2847
rect 12270 2774 12330 3804
rect 12390 2834 12450 3866
rect 12510 2774 12570 3804
rect 12630 2834 12690 3866
rect 12750 3712 12816 3866
rect 12750 3648 12751 3712
rect 12815 3648 12816 3712
rect 12750 3632 12816 3648
rect 12750 3568 12751 3632
rect 12815 3568 12816 3632
rect 12750 3552 12816 3568
rect 12750 3488 12751 3552
rect 12815 3488 12816 3552
rect 12750 3472 12816 3488
rect 12750 3408 12751 3472
rect 12815 3408 12816 3472
rect 12750 3392 12816 3408
rect 12750 3328 12751 3392
rect 12815 3328 12816 3392
rect 12750 3312 12816 3328
rect 12750 3248 12751 3312
rect 12815 3248 12816 3312
rect 12750 3232 12816 3248
rect 12750 3168 12751 3232
rect 12815 3168 12816 3232
rect 12750 3152 12816 3168
rect 12750 3088 12751 3152
rect 12815 3088 12816 3152
rect 12750 3072 12816 3088
rect 12750 3008 12751 3072
rect 12815 3008 12816 3072
rect 12750 2992 12816 3008
rect 12750 2928 12751 2992
rect 12815 2928 12816 2992
rect 12750 2903 12816 2928
rect 12750 2847 12755 2903
rect 12811 2847 12816 2903
rect 12750 2838 12816 2847
rect 12876 2774 12936 3804
rect 12996 2834 13056 3866
rect 13116 2774 13176 3804
rect 13236 2834 13296 3866
rect 13356 3712 13422 3866
rect 13356 3648 13357 3712
rect 13421 3648 13422 3712
rect 13356 3632 13422 3648
rect 13356 3568 13357 3632
rect 13421 3568 13422 3632
rect 13356 3552 13422 3568
rect 13356 3488 13357 3552
rect 13421 3488 13422 3552
rect 13356 3472 13422 3488
rect 13356 3408 13357 3472
rect 13421 3408 13422 3472
rect 13356 3392 13422 3408
rect 13356 3328 13357 3392
rect 13421 3328 13422 3392
rect 13356 3312 13422 3328
rect 13356 3248 13357 3312
rect 13421 3248 13422 3312
rect 13356 3232 13422 3248
rect 13356 3168 13357 3232
rect 13421 3168 13422 3232
rect 13356 3152 13422 3168
rect 13356 3088 13357 3152
rect 13421 3088 13422 3152
rect 13356 3072 13422 3088
rect 13356 3008 13357 3072
rect 13421 3008 13422 3072
rect 13356 2992 13422 3008
rect 13356 2928 13357 2992
rect 13421 2928 13422 2992
rect 13356 2905 13422 2928
rect 13356 2849 13361 2905
rect 13417 2849 13422 2905
rect 13356 2838 13422 2849
rect 13482 2774 13542 3804
rect 13602 2834 13662 3866
rect 13722 2774 13782 3804
rect 13842 2834 13902 3866
rect 13962 3712 14028 3866
rect 13962 3648 13963 3712
rect 14027 3648 14028 3712
rect 13962 3632 14028 3648
rect 13962 3568 13963 3632
rect 14027 3568 14028 3632
rect 13962 3552 14028 3568
rect 13962 3488 13963 3552
rect 14027 3488 14028 3552
rect 13962 3472 14028 3488
rect 13962 3408 13963 3472
rect 14027 3408 14028 3472
rect 13962 3392 14028 3408
rect 13962 3328 13963 3392
rect 14027 3328 14028 3392
rect 13962 3312 14028 3328
rect 13962 3248 13963 3312
rect 14027 3248 14028 3312
rect 13962 3232 14028 3248
rect 13962 3168 13963 3232
rect 14027 3168 14028 3232
rect 13962 3152 14028 3168
rect 13962 3088 13963 3152
rect 14027 3088 14028 3152
rect 13962 3072 14028 3088
rect 13962 3008 13963 3072
rect 14027 3008 14028 3072
rect 13962 2992 14028 3008
rect 13962 2928 13963 2992
rect 14027 2928 14028 2992
rect 13962 2905 14028 2928
rect 13962 2849 13967 2905
rect 14023 2849 14028 2905
rect 13962 2838 14028 2849
rect 14088 2774 14148 3804
rect 14208 2834 14268 3866
rect 14328 2774 14388 3804
rect 14448 2834 14508 3866
rect 14568 3712 14634 3866
rect 14568 3648 14569 3712
rect 14633 3648 14634 3712
rect 14568 3632 14634 3648
rect 14568 3568 14569 3632
rect 14633 3568 14634 3632
rect 14568 3552 14634 3568
rect 14568 3488 14569 3552
rect 14633 3488 14634 3552
rect 14568 3472 14634 3488
rect 14568 3408 14569 3472
rect 14633 3408 14634 3472
rect 14568 3392 14634 3408
rect 14568 3328 14569 3392
rect 14633 3328 14634 3392
rect 14568 3312 14634 3328
rect 14568 3248 14569 3312
rect 14633 3248 14634 3312
rect 14568 3232 14634 3248
rect 14568 3168 14569 3232
rect 14633 3168 14634 3232
rect 14568 3152 14634 3168
rect 14568 3088 14569 3152
rect 14633 3088 14634 3152
rect 14568 3072 14634 3088
rect 14568 3008 14569 3072
rect 14633 3008 14634 3072
rect 14568 2992 14634 3008
rect 14568 2928 14569 2992
rect 14633 2928 14634 2992
rect 14568 2904 14634 2928
rect 14568 2848 14573 2904
rect 14629 2848 14634 2904
rect 14568 2838 14634 2848
rect 14694 2774 14754 3804
rect 14814 2834 14874 3866
rect 14934 2774 14994 3804
rect 15054 2834 15114 3866
rect 15174 3712 15240 3866
rect 15174 3648 15175 3712
rect 15239 3648 15240 3712
rect 15174 3632 15240 3648
rect 15174 3568 15175 3632
rect 15239 3568 15240 3632
rect 15174 3552 15240 3568
rect 15174 3488 15175 3552
rect 15239 3488 15240 3552
rect 15174 3472 15240 3488
rect 15174 3408 15175 3472
rect 15239 3408 15240 3472
rect 15174 3392 15240 3408
rect 15174 3328 15175 3392
rect 15239 3328 15240 3392
rect 15174 3312 15240 3328
rect 15174 3248 15175 3312
rect 15239 3248 15240 3312
rect 15174 3232 15240 3248
rect 15174 3168 15175 3232
rect 15239 3168 15240 3232
rect 15174 3152 15240 3168
rect 15174 3088 15175 3152
rect 15239 3088 15240 3152
rect 15174 3072 15240 3088
rect 15174 3008 15175 3072
rect 15239 3008 15240 3072
rect 15174 2992 15240 3008
rect 15174 2928 15175 2992
rect 15239 2928 15240 2992
rect 15174 2838 15240 2928
rect 15300 2774 15360 3804
rect 15420 2834 15480 3866
rect 15540 2774 15600 3804
rect 15660 2834 15720 3866
rect 15780 3712 15846 3866
rect 15780 3648 15781 3712
rect 15845 3648 15846 3712
rect 15780 3632 15846 3648
rect 15780 3568 15781 3632
rect 15845 3568 15846 3632
rect 15780 3552 15846 3568
rect 15780 3488 15781 3552
rect 15845 3488 15846 3552
rect 15780 3472 15846 3488
rect 15780 3408 15781 3472
rect 15845 3408 15846 3472
rect 15780 3392 15846 3408
rect 15780 3328 15781 3392
rect 15845 3328 15846 3392
rect 15780 3312 15846 3328
rect 15780 3248 15781 3312
rect 15845 3248 15846 3312
rect 15780 3232 15846 3248
rect 15780 3168 15781 3232
rect 15845 3168 15846 3232
rect 15780 3152 15846 3168
rect 15780 3088 15781 3152
rect 15845 3088 15846 3152
rect 15780 3072 15846 3088
rect 15780 3008 15781 3072
rect 15845 3008 15846 3072
rect 15780 2992 15846 3008
rect 15780 2928 15781 2992
rect 15845 2928 15846 2992
rect 15780 2838 15846 2928
rect 15906 2774 15966 3804
rect 16026 2834 16086 3866
rect 16146 2774 16206 3804
rect 16266 2834 16326 3866
rect 16386 3712 16452 3866
rect 16386 3648 16387 3712
rect 16451 3648 16452 3712
rect 16386 3632 16452 3648
rect 16386 3568 16387 3632
rect 16451 3568 16452 3632
rect 16386 3552 16452 3568
rect 16386 3488 16387 3552
rect 16451 3488 16452 3552
rect 16386 3472 16452 3488
rect 16386 3408 16387 3472
rect 16451 3408 16452 3472
rect 16386 3392 16452 3408
rect 16386 3328 16387 3392
rect 16451 3328 16452 3392
rect 16386 3312 16452 3328
rect 16386 3248 16387 3312
rect 16451 3248 16452 3312
rect 16386 3232 16452 3248
rect 16386 3168 16387 3232
rect 16451 3168 16452 3232
rect 16386 3152 16452 3168
rect 16386 3088 16387 3152
rect 16451 3088 16452 3152
rect 16386 3072 16452 3088
rect 16386 3008 16387 3072
rect 16451 3008 16452 3072
rect 16386 2992 16452 3008
rect 16386 2928 16387 2992
rect 16451 2928 16452 2992
rect 16386 2838 16452 2928
rect 16512 2774 16572 3804
rect 16632 2834 16692 3866
rect 16752 2774 16812 3804
rect 16872 2834 16932 3866
rect 16992 3712 17058 3866
rect 16992 3648 16993 3712
rect 17057 3648 17058 3712
rect 16992 3632 17058 3648
rect 16992 3568 16993 3632
rect 17057 3568 17058 3632
rect 16992 3552 17058 3568
rect 16992 3488 16993 3552
rect 17057 3488 17058 3552
rect 16992 3472 17058 3488
rect 16992 3408 16993 3472
rect 17057 3408 17058 3472
rect 16992 3392 17058 3408
rect 16992 3328 16993 3392
rect 17057 3328 17058 3392
rect 16992 3312 17058 3328
rect 16992 3248 16993 3312
rect 17057 3248 17058 3312
rect 16992 3232 17058 3248
rect 16992 3168 16993 3232
rect 17057 3168 17058 3232
rect 16992 3152 17058 3168
rect 16992 3088 16993 3152
rect 17057 3088 17058 3152
rect 16992 3072 17058 3088
rect 16992 3008 16993 3072
rect 17057 3008 17058 3072
rect 16992 2992 17058 3008
rect 16992 2928 16993 2992
rect 17057 2928 17058 2992
rect 16992 2838 17058 2928
rect 17118 2774 17178 3804
rect 17238 2834 17298 3866
rect 17358 2774 17418 3804
rect 17478 2834 17538 3866
rect 17598 3712 17664 3866
rect 17598 3648 17599 3712
rect 17663 3648 17664 3712
rect 17598 3632 17664 3648
rect 17598 3568 17599 3632
rect 17663 3568 17664 3632
rect 17598 3552 17664 3568
rect 17598 3488 17599 3552
rect 17663 3488 17664 3552
rect 17598 3472 17664 3488
rect 17598 3408 17599 3472
rect 17663 3408 17664 3472
rect 17598 3392 17664 3408
rect 17598 3328 17599 3392
rect 17663 3328 17664 3392
rect 17598 3312 17664 3328
rect 17598 3248 17599 3312
rect 17663 3248 17664 3312
rect 17598 3232 17664 3248
rect 17598 3168 17599 3232
rect 17663 3168 17664 3232
rect 17598 3152 17664 3168
rect 17598 3088 17599 3152
rect 17663 3088 17664 3152
rect 17598 3072 17664 3088
rect 17598 3008 17599 3072
rect 17663 3008 17664 3072
rect 17598 2992 17664 3008
rect 17598 2928 17599 2992
rect 17663 2928 17664 2992
rect 17598 2838 17664 2928
rect 17724 2774 17784 3804
rect 17844 2834 17904 3866
rect 17964 2774 18024 3804
rect 18084 2834 18144 3866
rect 18204 3712 18270 3866
rect 18204 3648 18205 3712
rect 18269 3648 18270 3712
rect 18204 3632 18270 3648
rect 18204 3568 18205 3632
rect 18269 3568 18270 3632
rect 18204 3552 18270 3568
rect 18204 3488 18205 3552
rect 18269 3488 18270 3552
rect 18204 3472 18270 3488
rect 18204 3408 18205 3472
rect 18269 3408 18270 3472
rect 18204 3392 18270 3408
rect 18204 3328 18205 3392
rect 18269 3328 18270 3392
rect 18204 3312 18270 3328
rect 18204 3248 18205 3312
rect 18269 3248 18270 3312
rect 18204 3232 18270 3248
rect 18204 3168 18205 3232
rect 18269 3168 18270 3232
rect 18204 3152 18270 3168
rect 18204 3088 18205 3152
rect 18269 3088 18270 3152
rect 18204 3072 18270 3088
rect 18204 3008 18205 3072
rect 18269 3008 18270 3072
rect 18204 2992 18270 3008
rect 18204 2928 18205 2992
rect 18269 2928 18270 2992
rect 18204 2838 18270 2928
rect 18330 2774 18390 3804
rect 18450 2834 18510 3866
rect 18570 2774 18630 3804
rect 18690 2834 18750 3866
rect 18810 3712 18876 3866
rect 18810 3648 18811 3712
rect 18875 3648 18876 3712
rect 18810 3632 18876 3648
rect 18810 3568 18811 3632
rect 18875 3568 18876 3632
rect 18810 3552 18876 3568
rect 18810 3488 18811 3552
rect 18875 3488 18876 3552
rect 18810 3472 18876 3488
rect 18810 3408 18811 3472
rect 18875 3408 18876 3472
rect 18810 3392 18876 3408
rect 18810 3328 18811 3392
rect 18875 3328 18876 3392
rect 18810 3312 18876 3328
rect 18810 3248 18811 3312
rect 18875 3248 18876 3312
rect 18810 3232 18876 3248
rect 18810 3168 18811 3232
rect 18875 3168 18876 3232
rect 18810 3152 18876 3168
rect 18810 3088 18811 3152
rect 18875 3088 18876 3152
rect 18810 3072 18876 3088
rect 18810 3008 18811 3072
rect 18875 3008 18876 3072
rect 18810 2992 18876 3008
rect 18810 2928 18811 2992
rect 18875 2928 18876 2992
rect 18810 2838 18876 2928
rect 18936 2774 18996 3804
rect 19056 2834 19116 3866
rect 19176 2774 19236 3804
rect 19296 2834 19356 3866
rect 19416 3712 19482 3866
rect 19416 3648 19417 3712
rect 19481 3648 19482 3712
rect 19416 3632 19482 3648
rect 19416 3568 19417 3632
rect 19481 3568 19482 3632
rect 19416 3552 19482 3568
rect 19416 3488 19417 3552
rect 19481 3488 19482 3552
rect 19416 3472 19482 3488
rect 19416 3408 19417 3472
rect 19481 3408 19482 3472
rect 19416 3392 19482 3408
rect 19416 3328 19417 3392
rect 19481 3328 19482 3392
rect 19416 3312 19482 3328
rect 19416 3248 19417 3312
rect 19481 3248 19482 3312
rect 19416 3232 19482 3248
rect 19416 3168 19417 3232
rect 19481 3168 19482 3232
rect 19416 3152 19482 3168
rect 19416 3088 19417 3152
rect 19481 3088 19482 3152
rect 19416 3072 19482 3088
rect 19416 3008 19417 3072
rect 19481 3008 19482 3072
rect 19416 2992 19482 3008
rect 19416 2928 19417 2992
rect 19481 2928 19482 2992
rect 19416 2838 19482 2928
rect 19542 2774 19602 3804
rect 19662 2834 19722 3866
rect 19782 2774 19842 3804
rect 19902 2834 19962 3866
rect 20022 3712 20088 3866
rect 20022 3648 20023 3712
rect 20087 3648 20088 3712
rect 20022 3632 20088 3648
rect 20022 3568 20023 3632
rect 20087 3568 20088 3632
rect 20022 3552 20088 3568
rect 20022 3488 20023 3552
rect 20087 3488 20088 3552
rect 20022 3472 20088 3488
rect 20022 3408 20023 3472
rect 20087 3408 20088 3472
rect 20022 3392 20088 3408
rect 20022 3328 20023 3392
rect 20087 3328 20088 3392
rect 20022 3312 20088 3328
rect 20022 3248 20023 3312
rect 20087 3248 20088 3312
rect 20022 3232 20088 3248
rect 20022 3168 20023 3232
rect 20087 3168 20088 3232
rect 20022 3152 20088 3168
rect 20022 3088 20023 3152
rect 20087 3088 20088 3152
rect 20022 3072 20088 3088
rect 20022 3008 20023 3072
rect 20087 3008 20088 3072
rect 20022 2992 20088 3008
rect 20022 2928 20023 2992
rect 20087 2928 20088 2992
rect 20022 2838 20088 2928
rect 20148 4872 20214 4962
rect 20148 4808 20149 4872
rect 20213 4808 20214 4872
rect 20148 4792 20214 4808
rect 20148 4728 20149 4792
rect 20213 4728 20214 4792
rect 20148 4712 20214 4728
rect 20148 4648 20149 4712
rect 20213 4648 20214 4712
rect 20148 4632 20214 4648
rect 20148 4568 20149 4632
rect 20213 4568 20214 4632
rect 20148 4552 20214 4568
rect 20148 4488 20149 4552
rect 20213 4488 20214 4552
rect 20148 4472 20214 4488
rect 20148 4408 20149 4472
rect 20213 4408 20214 4472
rect 20148 4392 20214 4408
rect 20148 4328 20149 4392
rect 20213 4328 20214 4392
rect 20148 4312 20214 4328
rect 20148 4248 20149 4312
rect 20213 4248 20214 4312
rect 20148 4232 20214 4248
rect 20148 4168 20149 4232
rect 20213 4168 20214 4232
rect 20148 4152 20214 4168
rect 20148 4088 20149 4152
rect 20213 4088 20214 4152
rect 20148 3934 20214 4088
rect 20274 3934 20334 4966
rect 20394 3996 20454 5026
rect 20514 3934 20574 4966
rect 20634 3996 20694 5026
rect 20754 4872 20820 4962
rect 20754 4808 20755 4872
rect 20819 4808 20820 4872
rect 20754 4792 20820 4808
rect 20754 4728 20755 4792
rect 20819 4728 20820 4792
rect 20754 4712 20820 4728
rect 20754 4648 20755 4712
rect 20819 4648 20820 4712
rect 20754 4632 20820 4648
rect 20754 4568 20755 4632
rect 20819 4568 20820 4632
rect 20754 4552 20820 4568
rect 20754 4488 20755 4552
rect 20819 4488 20820 4552
rect 20754 4472 20820 4488
rect 20754 4408 20755 4472
rect 20819 4408 20820 4472
rect 20754 4392 20820 4408
rect 20754 4328 20755 4392
rect 20819 4328 20820 4392
rect 20754 4312 20820 4328
rect 20754 4248 20755 4312
rect 20819 4248 20820 4312
rect 20754 4232 20820 4248
rect 20754 4168 20755 4232
rect 20819 4168 20820 4232
rect 20754 4152 20820 4168
rect 20754 4088 20755 4152
rect 20819 4088 20820 4152
rect 20754 3934 20820 4088
rect 20880 3934 20940 4966
rect 21000 3996 21060 5026
rect 21120 3934 21180 4966
rect 21240 3996 21300 5026
rect 21360 4872 21426 4962
rect 21360 4808 21361 4872
rect 21425 4808 21426 4872
rect 21360 4792 21426 4808
rect 21360 4728 21361 4792
rect 21425 4728 21426 4792
rect 21360 4712 21426 4728
rect 21360 4648 21361 4712
rect 21425 4648 21426 4712
rect 21360 4632 21426 4648
rect 21360 4568 21361 4632
rect 21425 4568 21426 4632
rect 21360 4552 21426 4568
rect 21360 4488 21361 4552
rect 21425 4488 21426 4552
rect 21360 4472 21426 4488
rect 21360 4408 21361 4472
rect 21425 4408 21426 4472
rect 21360 4392 21426 4408
rect 21360 4328 21361 4392
rect 21425 4328 21426 4392
rect 21360 4312 21426 4328
rect 21360 4248 21361 4312
rect 21425 4248 21426 4312
rect 21360 4232 21426 4248
rect 21360 4168 21361 4232
rect 21425 4168 21426 4232
rect 21360 4152 21426 4168
rect 21360 4088 21361 4152
rect 21425 4088 21426 4152
rect 21360 3934 21426 4088
rect 21486 3934 21546 4966
rect 21606 3996 21666 5026
rect 21726 3934 21786 4966
rect 21846 3996 21906 5026
rect 21966 4872 22032 4962
rect 21966 4808 21967 4872
rect 22031 4808 22032 4872
rect 21966 4792 22032 4808
rect 21966 4728 21967 4792
rect 22031 4728 22032 4792
rect 21966 4712 22032 4728
rect 21966 4648 21967 4712
rect 22031 4648 22032 4712
rect 21966 4632 22032 4648
rect 21966 4568 21967 4632
rect 22031 4568 22032 4632
rect 21966 4552 22032 4568
rect 21966 4488 21967 4552
rect 22031 4488 22032 4552
rect 21966 4472 22032 4488
rect 21966 4408 21967 4472
rect 22031 4408 22032 4472
rect 21966 4392 22032 4408
rect 21966 4328 21967 4392
rect 22031 4328 22032 4392
rect 21966 4312 22032 4328
rect 21966 4248 21967 4312
rect 22031 4248 22032 4312
rect 21966 4232 22032 4248
rect 21966 4168 21967 4232
rect 22031 4168 22032 4232
rect 21966 4152 22032 4168
rect 21966 4088 21967 4152
rect 22031 4088 22032 4152
rect 21966 3934 22032 4088
rect 22092 3934 22152 4966
rect 22212 3996 22272 5026
rect 22332 3934 22392 4966
rect 22452 3996 22512 5026
rect 22572 4872 22638 4962
rect 22572 4808 22573 4872
rect 22637 4808 22638 4872
rect 22572 4792 22638 4808
rect 22572 4728 22573 4792
rect 22637 4728 22638 4792
rect 22572 4712 22638 4728
rect 22572 4648 22573 4712
rect 22637 4648 22638 4712
rect 22572 4632 22638 4648
rect 22572 4568 22573 4632
rect 22637 4568 22638 4632
rect 22572 4552 22638 4568
rect 22572 4488 22573 4552
rect 22637 4488 22638 4552
rect 22572 4472 22638 4488
rect 22572 4408 22573 4472
rect 22637 4408 22638 4472
rect 22572 4392 22638 4408
rect 22572 4328 22573 4392
rect 22637 4328 22638 4392
rect 22572 4312 22638 4328
rect 22572 4248 22573 4312
rect 22637 4248 22638 4312
rect 22572 4232 22638 4248
rect 22572 4168 22573 4232
rect 22637 4168 22638 4232
rect 22572 4152 22638 4168
rect 22572 4088 22573 4152
rect 22637 4088 22638 4152
rect 22572 3934 22638 4088
rect 22698 3934 22758 4966
rect 22818 3996 22878 5026
rect 22938 3934 22998 4966
rect 23058 3996 23118 5026
rect 23178 4872 23244 4962
rect 23178 4808 23179 4872
rect 23243 4808 23244 4872
rect 23178 4792 23244 4808
rect 23178 4728 23179 4792
rect 23243 4728 23244 4792
rect 23178 4712 23244 4728
rect 23178 4648 23179 4712
rect 23243 4648 23244 4712
rect 23178 4632 23244 4648
rect 23178 4568 23179 4632
rect 23243 4568 23244 4632
rect 23178 4552 23244 4568
rect 23178 4488 23179 4552
rect 23243 4488 23244 4552
rect 23178 4472 23244 4488
rect 23178 4408 23179 4472
rect 23243 4408 23244 4472
rect 23178 4392 23244 4408
rect 23178 4328 23179 4392
rect 23243 4328 23244 4392
rect 23178 4312 23244 4328
rect 23178 4248 23179 4312
rect 23243 4248 23244 4312
rect 23178 4232 23244 4248
rect 23178 4168 23179 4232
rect 23243 4168 23244 4232
rect 23178 4152 23244 4168
rect 23178 4088 23179 4152
rect 23243 4088 23244 4152
rect 23178 3934 23244 4088
rect 23304 3934 23364 4966
rect 23424 3996 23484 5026
rect 23544 3934 23604 4966
rect 23664 3996 23724 5026
rect 23784 4872 23850 4962
rect 23784 4808 23785 4872
rect 23849 4808 23850 4872
rect 23784 4792 23850 4808
rect 23784 4728 23785 4792
rect 23849 4728 23850 4792
rect 23784 4712 23850 4728
rect 23784 4648 23785 4712
rect 23849 4648 23850 4712
rect 23784 4632 23850 4648
rect 23784 4568 23785 4632
rect 23849 4568 23850 4632
rect 23784 4552 23850 4568
rect 23784 4488 23785 4552
rect 23849 4488 23850 4552
rect 23784 4472 23850 4488
rect 23784 4408 23785 4472
rect 23849 4408 23850 4472
rect 23784 4392 23850 4408
rect 23784 4328 23785 4392
rect 23849 4328 23850 4392
rect 23784 4312 23850 4328
rect 23784 4248 23785 4312
rect 23849 4248 23850 4312
rect 23784 4232 23850 4248
rect 23784 4168 23785 4232
rect 23849 4168 23850 4232
rect 23784 4152 23850 4168
rect 23784 4088 23785 4152
rect 23849 4088 23850 4152
rect 23784 3934 23850 4088
rect 23910 3934 23970 4966
rect 24030 3996 24090 5026
rect 24150 3934 24210 4966
rect 24270 3996 24330 5026
rect 24390 4872 24456 4962
rect 24390 4808 24391 4872
rect 24455 4808 24456 4872
rect 24390 4792 24456 4808
rect 24390 4728 24391 4792
rect 24455 4728 24456 4792
rect 24390 4712 24456 4728
rect 24390 4648 24391 4712
rect 24455 4648 24456 4712
rect 24390 4632 24456 4648
rect 24390 4568 24391 4632
rect 24455 4568 24456 4632
rect 24390 4552 24456 4568
rect 24390 4488 24391 4552
rect 24455 4488 24456 4552
rect 24390 4472 24456 4488
rect 24390 4408 24391 4472
rect 24455 4408 24456 4472
rect 24390 4392 24456 4408
rect 24390 4328 24391 4392
rect 24455 4328 24456 4392
rect 24390 4312 24456 4328
rect 24390 4248 24391 4312
rect 24455 4248 24456 4312
rect 24390 4232 24456 4248
rect 24390 4168 24391 4232
rect 24455 4168 24456 4232
rect 24390 4152 24456 4168
rect 24390 4088 24391 4152
rect 24455 4088 24456 4152
rect 24390 3934 24456 4088
rect 24516 3934 24576 4966
rect 24636 3996 24696 5026
rect 24756 3934 24816 4966
rect 24876 3996 24936 5026
rect 24996 4872 25062 4962
rect 24996 4808 24997 4872
rect 25061 4808 25062 4872
rect 24996 4792 25062 4808
rect 24996 4728 24997 4792
rect 25061 4728 25062 4792
rect 24996 4712 25062 4728
rect 24996 4648 24997 4712
rect 25061 4648 25062 4712
rect 24996 4632 25062 4648
rect 24996 4568 24997 4632
rect 25061 4568 25062 4632
rect 24996 4552 25062 4568
rect 24996 4488 24997 4552
rect 25061 4488 25062 4552
rect 24996 4472 25062 4488
rect 24996 4408 24997 4472
rect 25061 4408 25062 4472
rect 24996 4392 25062 4408
rect 24996 4328 24997 4392
rect 25061 4328 25062 4392
rect 24996 4312 25062 4328
rect 24996 4248 24997 4312
rect 25061 4248 25062 4312
rect 24996 4232 25062 4248
rect 24996 4168 24997 4232
rect 25061 4168 25062 4232
rect 24996 4152 25062 4168
rect 24996 4088 24997 4152
rect 25061 4088 25062 4152
rect 24996 3934 25062 4088
rect 25122 3934 25182 4966
rect 25242 3996 25302 5026
rect 25362 3934 25422 4966
rect 25482 3996 25542 5026
rect 25602 4872 25668 4962
rect 25602 4808 25603 4872
rect 25667 4808 25668 4872
rect 25602 4792 25668 4808
rect 25602 4728 25603 4792
rect 25667 4728 25668 4792
rect 25602 4712 25668 4728
rect 25602 4648 25603 4712
rect 25667 4648 25668 4712
rect 25602 4632 25668 4648
rect 25602 4568 25603 4632
rect 25667 4568 25668 4632
rect 25602 4552 25668 4568
rect 25602 4488 25603 4552
rect 25667 4488 25668 4552
rect 25602 4472 25668 4488
rect 25602 4408 25603 4472
rect 25667 4408 25668 4472
rect 25602 4392 25668 4408
rect 25602 4328 25603 4392
rect 25667 4328 25668 4392
rect 25602 4312 25668 4328
rect 25602 4248 25603 4312
rect 25667 4248 25668 4312
rect 25602 4232 25668 4248
rect 25602 4168 25603 4232
rect 25667 4168 25668 4232
rect 25602 4152 25668 4168
rect 25602 4088 25603 4152
rect 25667 4088 25668 4152
rect 25602 3934 25668 4088
rect 25728 3934 25788 4966
rect 25848 3996 25908 5026
rect 25968 3934 26028 4966
rect 26088 3996 26148 5026
rect 26208 4872 26274 4962
rect 26208 4808 26209 4872
rect 26273 4808 26274 4872
rect 26208 4792 26274 4808
rect 26208 4728 26209 4792
rect 26273 4728 26274 4792
rect 26208 4712 26274 4728
rect 26208 4648 26209 4712
rect 26273 4648 26274 4712
rect 26208 4632 26274 4648
rect 26208 4568 26209 4632
rect 26273 4568 26274 4632
rect 26208 4552 26274 4568
rect 26208 4488 26209 4552
rect 26273 4488 26274 4552
rect 26208 4472 26274 4488
rect 26208 4408 26209 4472
rect 26273 4408 26274 4472
rect 26208 4392 26274 4408
rect 26208 4328 26209 4392
rect 26273 4328 26274 4392
rect 26208 4312 26274 4328
rect 26208 4248 26209 4312
rect 26273 4248 26274 4312
rect 26208 4232 26274 4248
rect 26208 4168 26209 4232
rect 26273 4168 26274 4232
rect 26208 4152 26274 4168
rect 26208 4088 26209 4152
rect 26273 4088 26274 4152
rect 26208 3934 26274 4088
rect 26334 3934 26394 4966
rect 26454 3996 26514 5026
rect 26574 3934 26634 4966
rect 26694 3996 26754 5026
rect 26814 4872 26880 4962
rect 26814 4808 26815 4872
rect 26879 4808 26880 4872
rect 26814 4792 26880 4808
rect 26814 4728 26815 4792
rect 26879 4728 26880 4792
rect 26814 4712 26880 4728
rect 26814 4648 26815 4712
rect 26879 4648 26880 4712
rect 26814 4632 26880 4648
rect 26814 4568 26815 4632
rect 26879 4568 26880 4632
rect 26814 4552 26880 4568
rect 26814 4488 26815 4552
rect 26879 4488 26880 4552
rect 26814 4472 26880 4488
rect 26814 4408 26815 4472
rect 26879 4408 26880 4472
rect 26814 4392 26880 4408
rect 26814 4328 26815 4392
rect 26879 4328 26880 4392
rect 26814 4312 26880 4328
rect 26814 4248 26815 4312
rect 26879 4248 26880 4312
rect 26814 4232 26880 4248
rect 26814 4168 26815 4232
rect 26879 4168 26880 4232
rect 26814 4152 26880 4168
rect 26814 4088 26815 4152
rect 26879 4088 26880 4152
rect 26814 3934 26880 4088
rect 26940 3934 27000 4966
rect 27060 3996 27120 5026
rect 27180 3934 27240 4966
rect 27300 3996 27360 5026
rect 27420 4872 27486 4962
rect 27420 4808 27421 4872
rect 27485 4808 27486 4872
rect 27420 4792 27486 4808
rect 27420 4728 27421 4792
rect 27485 4728 27486 4792
rect 27420 4712 27486 4728
rect 27420 4648 27421 4712
rect 27485 4648 27486 4712
rect 27420 4632 27486 4648
rect 27420 4568 27421 4632
rect 27485 4568 27486 4632
rect 27420 4552 27486 4568
rect 27420 4488 27421 4552
rect 27485 4488 27486 4552
rect 27420 4472 27486 4488
rect 27420 4408 27421 4472
rect 27485 4408 27486 4472
rect 27420 4392 27486 4408
rect 27420 4328 27421 4392
rect 27485 4328 27486 4392
rect 27420 4312 27486 4328
rect 27420 4248 27421 4312
rect 27485 4248 27486 4312
rect 27420 4232 27486 4248
rect 27420 4168 27421 4232
rect 27485 4168 27486 4232
rect 27420 4152 27486 4168
rect 27420 4088 27421 4152
rect 27485 4088 27486 4152
rect 27420 3934 27486 4088
rect 27546 3934 27606 4966
rect 27666 3996 27726 5026
rect 27786 3934 27846 4966
rect 27906 3996 27966 5026
rect 28026 4872 28092 4962
rect 28026 4808 28027 4872
rect 28091 4808 28092 4872
rect 28026 4792 28092 4808
rect 28026 4728 28027 4792
rect 28091 4728 28092 4792
rect 28026 4712 28092 4728
rect 28026 4648 28027 4712
rect 28091 4648 28092 4712
rect 28026 4632 28092 4648
rect 28026 4568 28027 4632
rect 28091 4568 28092 4632
rect 28026 4552 28092 4568
rect 28026 4488 28027 4552
rect 28091 4488 28092 4552
rect 28026 4472 28092 4488
rect 28026 4408 28027 4472
rect 28091 4408 28092 4472
rect 28026 4392 28092 4408
rect 28026 4328 28027 4392
rect 28091 4328 28092 4392
rect 28026 4312 28092 4328
rect 28026 4248 28027 4312
rect 28091 4248 28092 4312
rect 28026 4232 28092 4248
rect 28026 4168 28027 4232
rect 28091 4168 28092 4232
rect 28026 4152 28092 4168
rect 28026 4088 28027 4152
rect 28091 4088 28092 4152
rect 28026 3934 28092 4088
rect 28152 3934 28212 4966
rect 28272 3996 28332 5026
rect 28392 3934 28452 4966
rect 28512 3996 28572 5026
rect 28632 4872 28698 4962
rect 28632 4808 28633 4872
rect 28697 4808 28698 4872
rect 28632 4792 28698 4808
rect 28632 4728 28633 4792
rect 28697 4728 28698 4792
rect 28632 4712 28698 4728
rect 28632 4648 28633 4712
rect 28697 4648 28698 4712
rect 28632 4632 28698 4648
rect 28632 4568 28633 4632
rect 28697 4568 28698 4632
rect 28632 4552 28698 4568
rect 28632 4488 28633 4552
rect 28697 4488 28698 4552
rect 28632 4472 28698 4488
rect 28632 4408 28633 4472
rect 28697 4408 28698 4472
rect 28632 4392 28698 4408
rect 28632 4328 28633 4392
rect 28697 4328 28698 4392
rect 28632 4312 28698 4328
rect 28632 4248 28633 4312
rect 28697 4248 28698 4312
rect 28632 4232 28698 4248
rect 28632 4168 28633 4232
rect 28697 4168 28698 4232
rect 28632 4152 28698 4168
rect 28632 4088 28633 4152
rect 28697 4088 28698 4152
rect 28632 3934 28698 4088
rect 28758 3934 28818 4966
rect 28878 3996 28938 5026
rect 28998 3934 29058 4966
rect 29118 3996 29178 5026
rect 29238 4872 29304 4962
rect 29238 4808 29239 4872
rect 29303 4808 29304 4872
rect 29238 4792 29304 4808
rect 29238 4728 29239 4792
rect 29303 4728 29304 4792
rect 29238 4712 29304 4728
rect 29238 4648 29239 4712
rect 29303 4648 29304 4712
rect 29238 4632 29304 4648
rect 29238 4568 29239 4632
rect 29303 4568 29304 4632
rect 29238 4552 29304 4568
rect 29238 4488 29239 4552
rect 29303 4488 29304 4552
rect 29238 4472 29304 4488
rect 29238 4408 29239 4472
rect 29303 4408 29304 4472
rect 29238 4392 29304 4408
rect 29238 4328 29239 4392
rect 29303 4328 29304 4392
rect 29238 4312 29304 4328
rect 29238 4248 29239 4312
rect 29303 4248 29304 4312
rect 29238 4232 29304 4248
rect 29238 4168 29239 4232
rect 29303 4168 29304 4232
rect 29238 4152 29304 4168
rect 29238 4088 29239 4152
rect 29303 4088 29304 4152
rect 29238 3934 29304 4088
rect 29364 3934 29424 4966
rect 29484 3996 29544 5026
rect 29604 3934 29664 4966
rect 29724 3996 29784 5026
rect 29844 4872 29910 4962
rect 29844 4808 29845 4872
rect 29909 4808 29910 4872
rect 29844 4792 29910 4808
rect 29844 4728 29845 4792
rect 29909 4728 29910 4792
rect 29844 4712 29910 4728
rect 29844 4648 29845 4712
rect 29909 4648 29910 4712
rect 29844 4632 29910 4648
rect 29844 4568 29845 4632
rect 29909 4568 29910 4632
rect 29844 4552 29910 4568
rect 29844 4488 29845 4552
rect 29909 4488 29910 4552
rect 29844 4472 29910 4488
rect 29844 4408 29845 4472
rect 29909 4408 29910 4472
rect 29844 4392 29910 4408
rect 29844 4328 29845 4392
rect 29909 4328 29910 4392
rect 29844 4312 29910 4328
rect 29844 4248 29845 4312
rect 29909 4248 29910 4312
rect 29844 4232 29910 4248
rect 29844 4168 29845 4232
rect 29909 4168 29910 4232
rect 29844 4152 29910 4168
rect 29844 4088 29845 4152
rect 29909 4088 29910 4152
rect 29844 3934 29910 4088
rect 29970 3934 30030 4966
rect 30090 3996 30150 5026
rect 30210 3934 30270 4966
rect 30330 3996 30390 5026
rect 30450 4872 30516 4962
rect 30450 4808 30451 4872
rect 30515 4808 30516 4872
rect 30450 4792 30516 4808
rect 30450 4728 30451 4792
rect 30515 4728 30516 4792
rect 30450 4712 30516 4728
rect 30450 4648 30451 4712
rect 30515 4648 30516 4712
rect 30450 4632 30516 4648
rect 30450 4568 30451 4632
rect 30515 4568 30516 4632
rect 30450 4552 30516 4568
rect 30450 4488 30451 4552
rect 30515 4488 30516 4552
rect 30450 4472 30516 4488
rect 30450 4408 30451 4472
rect 30515 4408 30516 4472
rect 30450 4392 30516 4408
rect 30450 4328 30451 4392
rect 30515 4328 30516 4392
rect 30450 4312 30516 4328
rect 30450 4248 30451 4312
rect 30515 4248 30516 4312
rect 30450 4232 30516 4248
rect 30450 4168 30451 4232
rect 30515 4168 30516 4232
rect 30450 4152 30516 4168
rect 30450 4088 30451 4152
rect 30515 4088 30516 4152
rect 30450 3934 30516 4088
rect 30576 3934 30636 4966
rect 30696 3996 30756 5026
rect 30816 3934 30876 4966
rect 30936 3996 30996 5026
rect 31056 4872 31122 4962
rect 31056 4808 31057 4872
rect 31121 4808 31122 4872
rect 31056 4792 31122 4808
rect 31056 4728 31057 4792
rect 31121 4728 31122 4792
rect 31056 4712 31122 4728
rect 31056 4648 31057 4712
rect 31121 4648 31122 4712
rect 31056 4632 31122 4648
rect 31056 4568 31057 4632
rect 31121 4568 31122 4632
rect 31056 4552 31122 4568
rect 31056 4488 31057 4552
rect 31121 4488 31122 4552
rect 31056 4472 31122 4488
rect 31056 4408 31057 4472
rect 31121 4408 31122 4472
rect 31056 4392 31122 4408
rect 31056 4328 31057 4392
rect 31121 4328 31122 4392
rect 31056 4312 31122 4328
rect 31056 4248 31057 4312
rect 31121 4248 31122 4312
rect 31056 4232 31122 4248
rect 31056 4168 31057 4232
rect 31121 4168 31122 4232
rect 31056 4152 31122 4168
rect 31056 4088 31057 4152
rect 31121 4088 31122 4152
rect 31056 3934 31122 4088
rect 31182 3934 31242 4966
rect 31302 3996 31362 5026
rect 31422 3934 31482 4966
rect 31542 3996 31602 5026
rect 31662 4872 31728 4962
rect 31662 4808 31663 4872
rect 31727 4808 31728 4872
rect 31662 4792 31728 4808
rect 31662 4728 31663 4792
rect 31727 4728 31728 4792
rect 31662 4712 31728 4728
rect 31662 4648 31663 4712
rect 31727 4648 31728 4712
rect 31662 4632 31728 4648
rect 31662 4568 31663 4632
rect 31727 4568 31728 4632
rect 31662 4552 31728 4568
rect 31662 4488 31663 4552
rect 31727 4488 31728 4552
rect 31662 4472 31728 4488
rect 31662 4408 31663 4472
rect 31727 4408 31728 4472
rect 31662 4392 31728 4408
rect 31662 4328 31663 4392
rect 31727 4328 31728 4392
rect 31662 4312 31728 4328
rect 31662 4248 31663 4312
rect 31727 4248 31728 4312
rect 31662 4232 31728 4248
rect 31662 4168 31663 4232
rect 31727 4168 31728 4232
rect 31662 4152 31728 4168
rect 31662 4088 31663 4152
rect 31727 4088 31728 4152
rect 31662 3934 31728 4088
rect 31788 3934 31848 4966
rect 31908 3996 31968 5026
rect 32028 3934 32088 4966
rect 32148 3996 32208 5026
rect 32268 4872 32334 4962
rect 32268 4808 32269 4872
rect 32333 4808 32334 4872
rect 32268 4792 32334 4808
rect 32268 4728 32269 4792
rect 32333 4728 32334 4792
rect 32268 4712 32334 4728
rect 32268 4648 32269 4712
rect 32333 4648 32334 4712
rect 32268 4632 32334 4648
rect 32268 4568 32269 4632
rect 32333 4568 32334 4632
rect 32268 4552 32334 4568
rect 32268 4488 32269 4552
rect 32333 4488 32334 4552
rect 32268 4472 32334 4488
rect 32268 4408 32269 4472
rect 32333 4408 32334 4472
rect 32268 4392 32334 4408
rect 32268 4328 32269 4392
rect 32333 4328 32334 4392
rect 32268 4312 32334 4328
rect 32268 4248 32269 4312
rect 32333 4248 32334 4312
rect 32268 4232 32334 4248
rect 32268 4168 32269 4232
rect 32333 4168 32334 4232
rect 32268 4152 32334 4168
rect 32268 4088 32269 4152
rect 32333 4088 32334 4152
rect 32268 3934 32334 4088
rect 32394 3934 32454 4966
rect 32514 3996 32574 5026
rect 32634 3934 32694 4966
rect 32754 3996 32814 5026
rect 32874 4872 32940 4962
rect 32874 4808 32875 4872
rect 32939 4808 32940 4872
rect 32874 4792 32940 4808
rect 32874 4728 32875 4792
rect 32939 4728 32940 4792
rect 32874 4712 32940 4728
rect 32874 4648 32875 4712
rect 32939 4648 32940 4712
rect 32874 4632 32940 4648
rect 32874 4568 32875 4632
rect 32939 4568 32940 4632
rect 32874 4552 32940 4568
rect 32874 4488 32875 4552
rect 32939 4488 32940 4552
rect 32874 4472 32940 4488
rect 32874 4408 32875 4472
rect 32939 4408 32940 4472
rect 32874 4392 32940 4408
rect 32874 4328 32875 4392
rect 32939 4328 32940 4392
rect 32874 4312 32940 4328
rect 32874 4248 32875 4312
rect 32939 4248 32940 4312
rect 32874 4232 32940 4248
rect 32874 4168 32875 4232
rect 32939 4168 32940 4232
rect 32874 4152 32940 4168
rect 32874 4088 32875 4152
rect 32939 4088 32940 4152
rect 32874 3934 32940 4088
rect 33000 3934 33060 4966
rect 33120 3996 33180 5026
rect 33240 3934 33300 4966
rect 33360 3996 33420 5026
rect 33480 4872 33546 4962
rect 33480 4808 33481 4872
rect 33545 4808 33546 4872
rect 33480 4792 33546 4808
rect 33480 4728 33481 4792
rect 33545 4728 33546 4792
rect 33480 4712 33546 4728
rect 33480 4648 33481 4712
rect 33545 4648 33546 4712
rect 33480 4632 33546 4648
rect 33480 4568 33481 4632
rect 33545 4568 33546 4632
rect 33480 4552 33546 4568
rect 33480 4488 33481 4552
rect 33545 4488 33546 4552
rect 33480 4472 33546 4488
rect 33480 4408 33481 4472
rect 33545 4408 33546 4472
rect 33480 4392 33546 4408
rect 33480 4328 33481 4392
rect 33545 4328 33546 4392
rect 33480 4312 33546 4328
rect 33480 4248 33481 4312
rect 33545 4248 33546 4312
rect 33480 4232 33546 4248
rect 33480 4168 33481 4232
rect 33545 4168 33546 4232
rect 33480 4152 33546 4168
rect 33480 4088 33481 4152
rect 33545 4088 33546 4152
rect 33480 3934 33546 4088
rect 33606 3934 33666 4966
rect 33726 3996 33786 5026
rect 33846 3934 33906 4966
rect 33966 3996 34026 5026
rect 34086 4872 34152 4962
rect 34086 4808 34087 4872
rect 34151 4808 34152 4872
rect 34086 4792 34152 4808
rect 34086 4728 34087 4792
rect 34151 4728 34152 4792
rect 34086 4712 34152 4728
rect 34086 4648 34087 4712
rect 34151 4648 34152 4712
rect 34086 4632 34152 4648
rect 34086 4568 34087 4632
rect 34151 4568 34152 4632
rect 34086 4552 34152 4568
rect 34086 4488 34087 4552
rect 34151 4488 34152 4552
rect 34086 4472 34152 4488
rect 34086 4408 34087 4472
rect 34151 4408 34152 4472
rect 34086 4392 34152 4408
rect 34086 4328 34087 4392
rect 34151 4328 34152 4392
rect 34086 4312 34152 4328
rect 34086 4248 34087 4312
rect 34151 4248 34152 4312
rect 34086 4232 34152 4248
rect 34086 4168 34087 4232
rect 34151 4168 34152 4232
rect 34086 4152 34152 4168
rect 34086 4088 34087 4152
rect 34151 4088 34152 4152
rect 34086 3934 34152 4088
rect 34212 3934 34272 4966
rect 34332 3996 34392 5026
rect 34452 3934 34512 4966
rect 34572 3996 34632 5026
rect 34692 4872 34758 4962
rect 34692 4808 34693 4872
rect 34757 4808 34758 4872
rect 34692 4792 34758 4808
rect 34692 4728 34693 4792
rect 34757 4728 34758 4792
rect 34692 4712 34758 4728
rect 34692 4648 34693 4712
rect 34757 4648 34758 4712
rect 34692 4632 34758 4648
rect 34692 4568 34693 4632
rect 34757 4568 34758 4632
rect 34692 4552 34758 4568
rect 34692 4488 34693 4552
rect 34757 4488 34758 4552
rect 34692 4472 34758 4488
rect 34692 4408 34693 4472
rect 34757 4408 34758 4472
rect 34692 4392 34758 4408
rect 34692 4328 34693 4392
rect 34757 4328 34758 4392
rect 34692 4312 34758 4328
rect 34692 4248 34693 4312
rect 34757 4248 34758 4312
rect 34692 4232 34758 4248
rect 34692 4168 34693 4232
rect 34757 4168 34758 4232
rect 34692 4152 34758 4168
rect 34692 4088 34693 4152
rect 34757 4088 34758 4152
rect 34692 3934 34758 4088
rect 34818 3934 34878 4966
rect 34938 3996 34998 5026
rect 35058 3934 35118 4966
rect 35178 3996 35238 5026
rect 35298 4872 35364 4962
rect 35298 4808 35299 4872
rect 35363 4808 35364 4872
rect 35298 4792 35364 4808
rect 35298 4728 35299 4792
rect 35363 4728 35364 4792
rect 35298 4712 35364 4728
rect 35298 4648 35299 4712
rect 35363 4648 35364 4712
rect 35298 4632 35364 4648
rect 35298 4568 35299 4632
rect 35363 4568 35364 4632
rect 35298 4552 35364 4568
rect 35298 4488 35299 4552
rect 35363 4488 35364 4552
rect 35298 4472 35364 4488
rect 35298 4408 35299 4472
rect 35363 4408 35364 4472
rect 35298 4392 35364 4408
rect 35298 4328 35299 4392
rect 35363 4328 35364 4392
rect 35298 4312 35364 4328
rect 35298 4248 35299 4312
rect 35363 4248 35364 4312
rect 35298 4232 35364 4248
rect 35298 4168 35299 4232
rect 35363 4168 35364 4232
rect 35298 4152 35364 4168
rect 35298 4088 35299 4152
rect 35363 4088 35364 4152
rect 35298 3934 35364 4088
rect 35424 3934 35484 4966
rect 35544 3996 35604 5026
rect 35664 3934 35724 4966
rect 35784 3996 35844 5026
rect 35904 4872 35970 4962
rect 35904 4808 35905 4872
rect 35969 4808 35970 4872
rect 35904 4792 35970 4808
rect 35904 4728 35905 4792
rect 35969 4728 35970 4792
rect 35904 4712 35970 4728
rect 35904 4648 35905 4712
rect 35969 4648 35970 4712
rect 35904 4632 35970 4648
rect 35904 4568 35905 4632
rect 35969 4568 35970 4632
rect 35904 4552 35970 4568
rect 35904 4488 35905 4552
rect 35969 4488 35970 4552
rect 35904 4472 35970 4488
rect 35904 4408 35905 4472
rect 35969 4408 35970 4472
rect 35904 4392 35970 4408
rect 35904 4328 35905 4392
rect 35969 4328 35970 4392
rect 35904 4312 35970 4328
rect 35904 4248 35905 4312
rect 35969 4248 35970 4312
rect 35904 4232 35970 4248
rect 35904 4168 35905 4232
rect 35969 4168 35970 4232
rect 35904 4152 35970 4168
rect 35904 4088 35905 4152
rect 35969 4088 35970 4152
rect 35904 3934 35970 4088
rect 36030 3934 36090 4966
rect 36150 3996 36210 5026
rect 36270 3934 36330 4966
rect 36390 3996 36450 5026
rect 36510 4872 36576 4962
rect 36510 4808 36511 4872
rect 36575 4808 36576 4872
rect 36510 4792 36576 4808
rect 36510 4728 36511 4792
rect 36575 4728 36576 4792
rect 36510 4712 36576 4728
rect 36510 4648 36511 4712
rect 36575 4648 36576 4712
rect 36510 4632 36576 4648
rect 36510 4568 36511 4632
rect 36575 4568 36576 4632
rect 36510 4552 36576 4568
rect 36510 4488 36511 4552
rect 36575 4488 36576 4552
rect 36510 4472 36576 4488
rect 36510 4408 36511 4472
rect 36575 4408 36576 4472
rect 36510 4392 36576 4408
rect 36510 4328 36511 4392
rect 36575 4328 36576 4392
rect 36510 4312 36576 4328
rect 36510 4248 36511 4312
rect 36575 4248 36576 4312
rect 36510 4232 36576 4248
rect 36510 4168 36511 4232
rect 36575 4168 36576 4232
rect 36510 4152 36576 4168
rect 36510 4088 36511 4152
rect 36575 4088 36576 4152
rect 36510 3934 36576 4088
rect 36636 3934 36696 4966
rect 36756 3996 36816 5026
rect 36876 3934 36936 4966
rect 36996 3996 37056 5026
rect 37116 4872 37182 4962
rect 37116 4808 37117 4872
rect 37181 4808 37182 4872
rect 37116 4792 37182 4808
rect 37116 4728 37117 4792
rect 37181 4728 37182 4792
rect 37116 4712 37182 4728
rect 37116 4648 37117 4712
rect 37181 4648 37182 4712
rect 37116 4632 37182 4648
rect 37116 4568 37117 4632
rect 37181 4568 37182 4632
rect 37116 4552 37182 4568
rect 37116 4488 37117 4552
rect 37181 4488 37182 4552
rect 37116 4472 37182 4488
rect 37116 4408 37117 4472
rect 37181 4408 37182 4472
rect 37116 4392 37182 4408
rect 37116 4328 37117 4392
rect 37181 4328 37182 4392
rect 37116 4312 37182 4328
rect 37116 4248 37117 4312
rect 37181 4248 37182 4312
rect 37116 4232 37182 4248
rect 37116 4168 37117 4232
rect 37181 4168 37182 4232
rect 37116 4152 37182 4168
rect 37116 4088 37117 4152
rect 37181 4088 37182 4152
rect 37116 3934 37182 4088
rect 37242 3934 37302 4966
rect 37362 3996 37422 5026
rect 37482 3934 37542 4966
rect 37602 3996 37662 5026
rect 37722 4872 37788 4962
rect 37722 4808 37723 4872
rect 37787 4808 37788 4872
rect 37722 4792 37788 4808
rect 37722 4728 37723 4792
rect 37787 4728 37788 4792
rect 37722 4712 37788 4728
rect 37722 4648 37723 4712
rect 37787 4648 37788 4712
rect 37722 4632 37788 4648
rect 37722 4568 37723 4632
rect 37787 4568 37788 4632
rect 37722 4552 37788 4568
rect 37722 4488 37723 4552
rect 37787 4488 37788 4552
rect 37722 4472 37788 4488
rect 37722 4408 37723 4472
rect 37787 4408 37788 4472
rect 37722 4392 37788 4408
rect 37722 4328 37723 4392
rect 37787 4328 37788 4392
rect 37722 4312 37788 4328
rect 37722 4248 37723 4312
rect 37787 4248 37788 4312
rect 37722 4232 37788 4248
rect 37722 4168 37723 4232
rect 37787 4168 37788 4232
rect 37722 4152 37788 4168
rect 37722 4088 37723 4152
rect 37787 4088 37788 4152
rect 37722 3934 37788 4088
rect 37848 3934 37908 4966
rect 37968 3996 38028 5026
rect 38088 3934 38148 4966
rect 38208 3996 38268 5026
rect 38328 4872 38394 4962
rect 38328 4808 38329 4872
rect 38393 4808 38394 4872
rect 38328 4792 38394 4808
rect 38328 4728 38329 4792
rect 38393 4728 38394 4792
rect 38328 4712 38394 4728
rect 38328 4648 38329 4712
rect 38393 4648 38394 4712
rect 38328 4632 38394 4648
rect 38328 4568 38329 4632
rect 38393 4568 38394 4632
rect 38328 4552 38394 4568
rect 38328 4488 38329 4552
rect 38393 4488 38394 4552
rect 38328 4472 38394 4488
rect 38328 4408 38329 4472
rect 38393 4408 38394 4472
rect 38328 4392 38394 4408
rect 38328 4328 38329 4392
rect 38393 4328 38394 4392
rect 38328 4312 38394 4328
rect 38328 4248 38329 4312
rect 38393 4248 38394 4312
rect 38328 4232 38394 4248
rect 38328 4168 38329 4232
rect 38393 4168 38394 4232
rect 38328 4152 38394 4168
rect 38328 4088 38329 4152
rect 38393 4088 38394 4152
rect 38328 3934 38394 4088
rect 38454 3934 38514 4966
rect 38574 3996 38634 5026
rect 38694 3934 38754 4966
rect 38814 3996 38874 5026
rect 38934 4872 39000 4962
rect 38934 4808 38935 4872
rect 38999 4808 39000 4872
rect 38934 4792 39000 4808
rect 38934 4728 38935 4792
rect 38999 4728 39000 4792
rect 38934 4712 39000 4728
rect 38934 4648 38935 4712
rect 38999 4648 39000 4712
rect 38934 4632 39000 4648
rect 38934 4568 38935 4632
rect 38999 4568 39000 4632
rect 38934 4552 39000 4568
rect 38934 4488 38935 4552
rect 38999 4488 39000 4552
rect 38934 4472 39000 4488
rect 38934 4408 38935 4472
rect 38999 4408 39000 4472
rect 38934 4392 39000 4408
rect 38934 4328 38935 4392
rect 38999 4328 39000 4392
rect 38934 4312 39000 4328
rect 38934 4248 38935 4312
rect 38999 4248 39000 4312
rect 38934 4232 39000 4248
rect 38934 4168 38935 4232
rect 38999 4168 39000 4232
rect 38934 4152 39000 4168
rect 38934 4088 38935 4152
rect 38999 4088 39000 4152
rect 38934 3934 39000 4088
rect 39060 3934 39120 4966
rect 39180 3996 39240 5026
rect 39300 3934 39360 4966
rect 39420 3996 39480 5026
rect 39540 4872 39606 4962
rect 39540 4808 39541 4872
rect 39605 4808 39606 4872
rect 39540 4792 39606 4808
rect 39540 4728 39541 4792
rect 39605 4728 39606 4792
rect 39540 4712 39606 4728
rect 39540 4648 39541 4712
rect 39605 4648 39606 4712
rect 39540 4632 39606 4648
rect 39540 4568 39541 4632
rect 39605 4568 39606 4632
rect 39540 4552 39606 4568
rect 39540 4488 39541 4552
rect 39605 4488 39606 4552
rect 39540 4472 39606 4488
rect 39540 4408 39541 4472
rect 39605 4408 39606 4472
rect 39540 4392 39606 4408
rect 39540 4328 39541 4392
rect 39605 4328 39606 4392
rect 39540 4312 39606 4328
rect 39540 4248 39541 4312
rect 39605 4248 39606 4312
rect 39540 4232 39606 4248
rect 39540 4168 39541 4232
rect 39605 4168 39606 4232
rect 39540 4152 39606 4168
rect 39540 4088 39541 4152
rect 39605 4088 39606 4152
rect 39540 3934 39606 4088
rect 20148 3932 39606 3934
rect 20148 3868 20252 3932
rect 20316 3868 20332 3932
rect 20396 3868 20412 3932
rect 20476 3868 20492 3932
rect 20556 3868 20572 3932
rect 20636 3868 20652 3932
rect 20716 3868 20858 3932
rect 20922 3868 20938 3932
rect 21002 3868 21018 3932
rect 21082 3868 21098 3932
rect 21162 3868 21178 3932
rect 21242 3868 21258 3932
rect 21322 3868 21464 3932
rect 21528 3868 21544 3932
rect 21608 3868 21624 3932
rect 21688 3868 21704 3932
rect 21768 3868 21784 3932
rect 21848 3868 21864 3932
rect 21928 3868 22070 3932
rect 22134 3868 22150 3932
rect 22214 3868 22230 3932
rect 22294 3868 22310 3932
rect 22374 3868 22390 3932
rect 22454 3868 22470 3932
rect 22534 3868 22676 3932
rect 22740 3868 22756 3932
rect 22820 3868 22836 3932
rect 22900 3868 22916 3932
rect 22980 3868 22996 3932
rect 23060 3868 23076 3932
rect 23140 3868 23282 3932
rect 23346 3868 23362 3932
rect 23426 3868 23442 3932
rect 23506 3868 23522 3932
rect 23586 3868 23602 3932
rect 23666 3868 23682 3932
rect 23746 3868 23888 3932
rect 23952 3868 23968 3932
rect 24032 3868 24048 3932
rect 24112 3868 24128 3932
rect 24192 3868 24208 3932
rect 24272 3868 24288 3932
rect 24352 3868 24494 3932
rect 24558 3868 24574 3932
rect 24638 3868 24654 3932
rect 24718 3868 24734 3932
rect 24798 3868 24814 3932
rect 24878 3868 24894 3932
rect 24958 3868 25100 3932
rect 25164 3868 25180 3932
rect 25244 3868 25260 3932
rect 25324 3868 25340 3932
rect 25404 3868 25420 3932
rect 25484 3868 25500 3932
rect 25564 3868 25706 3932
rect 25770 3868 25786 3932
rect 25850 3868 25866 3932
rect 25930 3868 25946 3932
rect 26010 3868 26026 3932
rect 26090 3868 26106 3932
rect 26170 3868 26312 3932
rect 26376 3868 26392 3932
rect 26456 3868 26472 3932
rect 26536 3868 26552 3932
rect 26616 3868 26632 3932
rect 26696 3868 26712 3932
rect 26776 3868 26918 3932
rect 26982 3868 26998 3932
rect 27062 3868 27078 3932
rect 27142 3868 27158 3932
rect 27222 3868 27238 3932
rect 27302 3868 27318 3932
rect 27382 3868 27524 3932
rect 27588 3868 27604 3932
rect 27668 3868 27684 3932
rect 27748 3868 27764 3932
rect 27828 3868 27844 3932
rect 27908 3868 27924 3932
rect 27988 3868 28130 3932
rect 28194 3868 28210 3932
rect 28274 3868 28290 3932
rect 28354 3868 28370 3932
rect 28434 3868 28450 3932
rect 28514 3868 28530 3932
rect 28594 3868 28736 3932
rect 28800 3868 28816 3932
rect 28880 3868 28896 3932
rect 28960 3868 28976 3932
rect 29040 3868 29056 3932
rect 29120 3868 29136 3932
rect 29200 3868 29342 3932
rect 29406 3868 29422 3932
rect 29486 3868 29502 3932
rect 29566 3868 29582 3932
rect 29646 3868 29662 3932
rect 29726 3868 29742 3932
rect 29806 3868 29948 3932
rect 30012 3868 30028 3932
rect 30092 3868 30108 3932
rect 30172 3868 30188 3932
rect 30252 3868 30268 3932
rect 30332 3868 30348 3932
rect 30412 3868 30554 3932
rect 30618 3868 30634 3932
rect 30698 3868 30714 3932
rect 30778 3868 30794 3932
rect 30858 3868 30874 3932
rect 30938 3868 30954 3932
rect 31018 3868 31160 3932
rect 31224 3868 31240 3932
rect 31304 3868 31320 3932
rect 31384 3868 31400 3932
rect 31464 3868 31480 3932
rect 31544 3868 31560 3932
rect 31624 3868 31766 3932
rect 31830 3868 31846 3932
rect 31910 3868 31926 3932
rect 31990 3868 32006 3932
rect 32070 3868 32086 3932
rect 32150 3868 32166 3932
rect 32230 3868 32372 3932
rect 32436 3868 32452 3932
rect 32516 3868 32532 3932
rect 32596 3868 32612 3932
rect 32676 3868 32692 3932
rect 32756 3868 32772 3932
rect 32836 3868 32978 3932
rect 33042 3868 33058 3932
rect 33122 3868 33138 3932
rect 33202 3868 33218 3932
rect 33282 3868 33298 3932
rect 33362 3868 33378 3932
rect 33442 3868 33584 3932
rect 33648 3868 33664 3932
rect 33728 3868 33744 3932
rect 33808 3868 33824 3932
rect 33888 3868 33904 3932
rect 33968 3868 33984 3932
rect 34048 3868 34190 3932
rect 34254 3868 34270 3932
rect 34334 3868 34350 3932
rect 34414 3868 34430 3932
rect 34494 3868 34510 3932
rect 34574 3868 34590 3932
rect 34654 3868 34796 3932
rect 34860 3868 34876 3932
rect 34940 3868 34956 3932
rect 35020 3868 35036 3932
rect 35100 3868 35116 3932
rect 35180 3868 35196 3932
rect 35260 3868 35402 3932
rect 35466 3868 35482 3932
rect 35546 3868 35562 3932
rect 35626 3868 35642 3932
rect 35706 3868 35722 3932
rect 35786 3868 35802 3932
rect 35866 3868 36008 3932
rect 36072 3868 36088 3932
rect 36152 3868 36168 3932
rect 36232 3868 36248 3932
rect 36312 3868 36328 3932
rect 36392 3868 36408 3932
rect 36472 3868 36614 3932
rect 36678 3868 36694 3932
rect 36758 3868 36774 3932
rect 36838 3868 36854 3932
rect 36918 3868 36934 3932
rect 36998 3868 37014 3932
rect 37078 3868 37220 3932
rect 37284 3868 37300 3932
rect 37364 3868 37380 3932
rect 37444 3868 37460 3932
rect 37524 3868 37540 3932
rect 37604 3868 37620 3932
rect 37684 3868 37826 3932
rect 37890 3868 37906 3932
rect 37970 3868 37986 3932
rect 38050 3868 38066 3932
rect 38130 3868 38146 3932
rect 38210 3868 38226 3932
rect 38290 3868 38432 3932
rect 38496 3868 38512 3932
rect 38576 3868 38592 3932
rect 38656 3868 38672 3932
rect 38736 3868 38752 3932
rect 38816 3868 38832 3932
rect 38896 3868 39038 3932
rect 39102 3868 39118 3932
rect 39182 3868 39198 3932
rect 39262 3868 39278 3932
rect 39342 3868 39358 3932
rect 39422 3868 39438 3932
rect 39502 3868 39606 3932
rect 20148 3866 39606 3868
rect 20148 3712 20214 3866
rect 20148 3648 20149 3712
rect 20213 3648 20214 3712
rect 20148 3632 20214 3648
rect 20148 3568 20149 3632
rect 20213 3568 20214 3632
rect 20148 3552 20214 3568
rect 20148 3488 20149 3552
rect 20213 3488 20214 3552
rect 20148 3472 20214 3488
rect 20148 3408 20149 3472
rect 20213 3408 20214 3472
rect 20148 3392 20214 3408
rect 20148 3328 20149 3392
rect 20213 3328 20214 3392
rect 20148 3312 20214 3328
rect 20148 3248 20149 3312
rect 20213 3248 20214 3312
rect 20148 3232 20214 3248
rect 20148 3168 20149 3232
rect 20213 3168 20214 3232
rect 20148 3152 20214 3168
rect 20148 3088 20149 3152
rect 20213 3088 20214 3152
rect 20148 3072 20214 3088
rect 20148 3008 20149 3072
rect 20213 3008 20214 3072
rect 20148 2992 20214 3008
rect 20148 2928 20149 2992
rect 20213 2928 20214 2992
rect 20148 2904 20214 2928
rect 20148 2848 20153 2904
rect 20209 2848 20214 2904
rect 20148 2838 20214 2848
rect 20274 2774 20334 3804
rect 20394 2834 20454 3866
rect 20514 2774 20574 3804
rect 20634 2834 20694 3866
rect 20754 3712 20820 3866
rect 20754 3648 20755 3712
rect 20819 3648 20820 3712
rect 20754 3632 20820 3648
rect 20754 3568 20755 3632
rect 20819 3568 20820 3632
rect 20754 3552 20820 3568
rect 20754 3488 20755 3552
rect 20819 3488 20820 3552
rect 20754 3472 20820 3488
rect 20754 3408 20755 3472
rect 20819 3408 20820 3472
rect 20754 3392 20820 3408
rect 20754 3328 20755 3392
rect 20819 3328 20820 3392
rect 20754 3312 20820 3328
rect 20754 3248 20755 3312
rect 20819 3248 20820 3312
rect 20754 3232 20820 3248
rect 20754 3168 20755 3232
rect 20819 3168 20820 3232
rect 20754 3152 20820 3168
rect 20754 3088 20755 3152
rect 20819 3088 20820 3152
rect 20754 3072 20820 3088
rect 20754 3008 20755 3072
rect 20819 3008 20820 3072
rect 20754 2992 20820 3008
rect 20754 2928 20755 2992
rect 20819 2928 20820 2992
rect 20754 2904 20820 2928
rect 20754 2848 20759 2904
rect 20815 2848 20820 2904
rect 20754 2838 20820 2848
rect 20880 2774 20940 3804
rect 21000 2834 21060 3866
rect 21120 2774 21180 3804
rect 21240 2834 21300 3866
rect 21360 3712 21426 3866
rect 21360 3648 21361 3712
rect 21425 3648 21426 3712
rect 21360 3632 21426 3648
rect 21360 3568 21361 3632
rect 21425 3568 21426 3632
rect 21360 3552 21426 3568
rect 21360 3488 21361 3552
rect 21425 3488 21426 3552
rect 21360 3472 21426 3488
rect 21360 3408 21361 3472
rect 21425 3408 21426 3472
rect 21360 3392 21426 3408
rect 21360 3328 21361 3392
rect 21425 3328 21426 3392
rect 21360 3312 21426 3328
rect 21360 3248 21361 3312
rect 21425 3248 21426 3312
rect 21360 3232 21426 3248
rect 21360 3168 21361 3232
rect 21425 3168 21426 3232
rect 21360 3152 21426 3168
rect 21360 3088 21361 3152
rect 21425 3088 21426 3152
rect 21360 3072 21426 3088
rect 21360 3008 21361 3072
rect 21425 3008 21426 3072
rect 21360 2992 21426 3008
rect 21360 2928 21361 2992
rect 21425 2928 21426 2992
rect 21360 2905 21426 2928
rect 21360 2849 21365 2905
rect 21421 2849 21426 2905
rect 21360 2838 21426 2849
rect 21486 2774 21546 3804
rect 21606 2834 21666 3866
rect 21726 2774 21786 3804
rect 21846 2834 21906 3866
rect 21966 3712 22032 3866
rect 21966 3648 21967 3712
rect 22031 3648 22032 3712
rect 21966 3632 22032 3648
rect 21966 3568 21967 3632
rect 22031 3568 22032 3632
rect 21966 3552 22032 3568
rect 21966 3488 21967 3552
rect 22031 3488 22032 3552
rect 21966 3472 22032 3488
rect 21966 3408 21967 3472
rect 22031 3408 22032 3472
rect 21966 3392 22032 3408
rect 21966 3328 21967 3392
rect 22031 3328 22032 3392
rect 21966 3312 22032 3328
rect 21966 3248 21967 3312
rect 22031 3248 22032 3312
rect 21966 3232 22032 3248
rect 21966 3168 21967 3232
rect 22031 3168 22032 3232
rect 21966 3152 22032 3168
rect 21966 3088 21967 3152
rect 22031 3088 22032 3152
rect 21966 3072 22032 3088
rect 21966 3008 21967 3072
rect 22031 3008 22032 3072
rect 21966 2992 22032 3008
rect 21966 2928 21967 2992
rect 22031 2928 22032 2992
rect 21966 2904 22032 2928
rect 21966 2848 21971 2904
rect 22027 2848 22032 2904
rect 21966 2838 22032 2848
rect 22092 2774 22152 3804
rect 22212 2834 22272 3866
rect 22332 2774 22392 3804
rect 22452 2834 22512 3866
rect 22572 3712 22638 3866
rect 22572 3648 22573 3712
rect 22637 3648 22638 3712
rect 22572 3632 22638 3648
rect 22572 3568 22573 3632
rect 22637 3568 22638 3632
rect 22572 3552 22638 3568
rect 22572 3488 22573 3552
rect 22637 3488 22638 3552
rect 22572 3472 22638 3488
rect 22572 3408 22573 3472
rect 22637 3408 22638 3472
rect 22572 3392 22638 3408
rect 22572 3328 22573 3392
rect 22637 3328 22638 3392
rect 22572 3312 22638 3328
rect 22572 3248 22573 3312
rect 22637 3248 22638 3312
rect 22572 3232 22638 3248
rect 22572 3168 22573 3232
rect 22637 3168 22638 3232
rect 22572 3152 22638 3168
rect 22572 3088 22573 3152
rect 22637 3088 22638 3152
rect 22572 3072 22638 3088
rect 22572 3008 22573 3072
rect 22637 3008 22638 3072
rect 22572 2992 22638 3008
rect 22572 2928 22573 2992
rect 22637 2928 22638 2992
rect 22572 2904 22638 2928
rect 22572 2848 22577 2904
rect 22633 2848 22638 2904
rect 22572 2838 22638 2848
rect 22698 2774 22758 3804
rect 22818 2834 22878 3866
rect 22938 2774 22998 3804
rect 23058 2834 23118 3866
rect 23178 3712 23244 3866
rect 23178 3648 23179 3712
rect 23243 3648 23244 3712
rect 23178 3632 23244 3648
rect 23178 3568 23179 3632
rect 23243 3568 23244 3632
rect 23178 3552 23244 3568
rect 23178 3488 23179 3552
rect 23243 3488 23244 3552
rect 23178 3472 23244 3488
rect 23178 3408 23179 3472
rect 23243 3408 23244 3472
rect 23178 3392 23244 3408
rect 23178 3328 23179 3392
rect 23243 3328 23244 3392
rect 23178 3312 23244 3328
rect 23178 3248 23179 3312
rect 23243 3248 23244 3312
rect 23178 3232 23244 3248
rect 23178 3168 23179 3232
rect 23243 3168 23244 3232
rect 23178 3152 23244 3168
rect 23178 3088 23179 3152
rect 23243 3088 23244 3152
rect 23178 3072 23244 3088
rect 23178 3008 23179 3072
rect 23243 3008 23244 3072
rect 23178 2992 23244 3008
rect 23178 2928 23179 2992
rect 23243 2928 23244 2992
rect 23178 2904 23244 2928
rect 23178 2848 23183 2904
rect 23239 2848 23244 2904
rect 23178 2838 23244 2848
rect 23304 2774 23364 3804
rect 23424 2834 23484 3866
rect 23544 2774 23604 3804
rect 23664 2834 23724 3866
rect 23784 3712 23850 3866
rect 23784 3648 23785 3712
rect 23849 3648 23850 3712
rect 23784 3632 23850 3648
rect 23784 3568 23785 3632
rect 23849 3568 23850 3632
rect 23784 3552 23850 3568
rect 23784 3488 23785 3552
rect 23849 3488 23850 3552
rect 23784 3472 23850 3488
rect 23784 3408 23785 3472
rect 23849 3408 23850 3472
rect 23784 3392 23850 3408
rect 23784 3328 23785 3392
rect 23849 3328 23850 3392
rect 23784 3312 23850 3328
rect 23784 3248 23785 3312
rect 23849 3248 23850 3312
rect 23784 3232 23850 3248
rect 23784 3168 23785 3232
rect 23849 3168 23850 3232
rect 23784 3152 23850 3168
rect 23784 3088 23785 3152
rect 23849 3088 23850 3152
rect 23784 3072 23850 3088
rect 23784 3008 23785 3072
rect 23849 3008 23850 3072
rect 23784 2992 23850 3008
rect 23784 2928 23785 2992
rect 23849 2928 23850 2992
rect 23784 2904 23850 2928
rect 23784 2848 23789 2904
rect 23845 2848 23850 2904
rect 23784 2838 23850 2848
rect 23910 2774 23970 3804
rect 24030 2834 24090 3866
rect 24150 2774 24210 3804
rect 24270 2834 24330 3866
rect 24390 3712 24456 3866
rect 24390 3648 24391 3712
rect 24455 3648 24456 3712
rect 24390 3632 24456 3648
rect 24390 3568 24391 3632
rect 24455 3568 24456 3632
rect 24390 3552 24456 3568
rect 24390 3488 24391 3552
rect 24455 3488 24456 3552
rect 24390 3472 24456 3488
rect 24390 3408 24391 3472
rect 24455 3408 24456 3472
rect 24390 3392 24456 3408
rect 24390 3328 24391 3392
rect 24455 3328 24456 3392
rect 24390 3312 24456 3328
rect 24390 3248 24391 3312
rect 24455 3248 24456 3312
rect 24390 3232 24456 3248
rect 24390 3168 24391 3232
rect 24455 3168 24456 3232
rect 24390 3152 24456 3168
rect 24390 3088 24391 3152
rect 24455 3088 24456 3152
rect 24390 3072 24456 3088
rect 24390 3008 24391 3072
rect 24455 3008 24456 3072
rect 24390 2992 24456 3008
rect 24390 2928 24391 2992
rect 24455 2928 24456 2992
rect 24390 2904 24456 2928
rect 24390 2848 24395 2904
rect 24451 2848 24456 2904
rect 24390 2838 24456 2848
rect 24516 2774 24576 3804
rect 24636 2834 24696 3866
rect 24756 2774 24816 3804
rect 24876 2834 24936 3866
rect 24996 3712 25062 3866
rect 24996 3648 24997 3712
rect 25061 3648 25062 3712
rect 24996 3632 25062 3648
rect 24996 3568 24997 3632
rect 25061 3568 25062 3632
rect 24996 3552 25062 3568
rect 24996 3488 24997 3552
rect 25061 3488 25062 3552
rect 24996 3472 25062 3488
rect 24996 3408 24997 3472
rect 25061 3408 25062 3472
rect 24996 3392 25062 3408
rect 24996 3328 24997 3392
rect 25061 3328 25062 3392
rect 24996 3312 25062 3328
rect 24996 3248 24997 3312
rect 25061 3248 25062 3312
rect 24996 3232 25062 3248
rect 24996 3168 24997 3232
rect 25061 3168 25062 3232
rect 24996 3152 25062 3168
rect 24996 3088 24997 3152
rect 25061 3088 25062 3152
rect 24996 3072 25062 3088
rect 24996 3008 24997 3072
rect 25061 3008 25062 3072
rect 24996 2992 25062 3008
rect 24996 2928 24997 2992
rect 25061 2928 25062 2992
rect 24996 2904 25062 2928
rect 24996 2848 25001 2904
rect 25057 2848 25062 2904
rect 24996 2838 25062 2848
rect 25122 2774 25182 3804
rect 25242 2834 25302 3866
rect 25362 2774 25422 3804
rect 25482 2834 25542 3866
rect 25602 3712 25668 3866
rect 25602 3648 25603 3712
rect 25667 3648 25668 3712
rect 25602 3632 25668 3648
rect 25602 3568 25603 3632
rect 25667 3568 25668 3632
rect 25602 3552 25668 3568
rect 25602 3488 25603 3552
rect 25667 3488 25668 3552
rect 25602 3472 25668 3488
rect 25602 3408 25603 3472
rect 25667 3408 25668 3472
rect 25602 3392 25668 3408
rect 25602 3328 25603 3392
rect 25667 3328 25668 3392
rect 25602 3312 25668 3328
rect 25602 3248 25603 3312
rect 25667 3248 25668 3312
rect 25602 3232 25668 3248
rect 25602 3168 25603 3232
rect 25667 3168 25668 3232
rect 25602 3152 25668 3168
rect 25602 3088 25603 3152
rect 25667 3088 25668 3152
rect 25602 3072 25668 3088
rect 25602 3008 25603 3072
rect 25667 3008 25668 3072
rect 25602 2992 25668 3008
rect 25602 2928 25603 2992
rect 25667 2928 25668 2992
rect 25602 2904 25668 2928
rect 25602 2848 25607 2904
rect 25663 2848 25668 2904
rect 25602 2838 25668 2848
rect 25728 2774 25788 3804
rect 25848 2834 25908 3866
rect 25968 2774 26028 3804
rect 26088 2834 26148 3866
rect 26208 3712 26274 3866
rect 26208 3648 26209 3712
rect 26273 3648 26274 3712
rect 26208 3632 26274 3648
rect 26208 3568 26209 3632
rect 26273 3568 26274 3632
rect 26208 3552 26274 3568
rect 26208 3488 26209 3552
rect 26273 3488 26274 3552
rect 26208 3472 26274 3488
rect 26208 3408 26209 3472
rect 26273 3408 26274 3472
rect 26208 3392 26274 3408
rect 26208 3328 26209 3392
rect 26273 3328 26274 3392
rect 26208 3312 26274 3328
rect 26208 3248 26209 3312
rect 26273 3248 26274 3312
rect 26208 3232 26274 3248
rect 26208 3168 26209 3232
rect 26273 3168 26274 3232
rect 26208 3152 26274 3168
rect 26208 3088 26209 3152
rect 26273 3088 26274 3152
rect 26208 3072 26274 3088
rect 26208 3008 26209 3072
rect 26273 3008 26274 3072
rect 26208 2992 26274 3008
rect 26208 2928 26209 2992
rect 26273 2928 26274 2992
rect 26208 2904 26274 2928
rect 26208 2848 26213 2904
rect 26269 2848 26274 2904
rect 26208 2838 26274 2848
rect 26334 2774 26394 3804
rect 26454 2834 26514 3866
rect 26574 2774 26634 3804
rect 26694 2834 26754 3866
rect 26814 3712 26880 3866
rect 26814 3648 26815 3712
rect 26879 3648 26880 3712
rect 26814 3632 26880 3648
rect 26814 3568 26815 3632
rect 26879 3568 26880 3632
rect 26814 3552 26880 3568
rect 26814 3488 26815 3552
rect 26879 3488 26880 3552
rect 26814 3472 26880 3488
rect 26814 3408 26815 3472
rect 26879 3408 26880 3472
rect 26814 3392 26880 3408
rect 26814 3328 26815 3392
rect 26879 3328 26880 3392
rect 26814 3312 26880 3328
rect 26814 3248 26815 3312
rect 26879 3248 26880 3312
rect 26814 3232 26880 3248
rect 26814 3168 26815 3232
rect 26879 3168 26880 3232
rect 26814 3152 26880 3168
rect 26814 3088 26815 3152
rect 26879 3088 26880 3152
rect 26814 3072 26880 3088
rect 26814 3008 26815 3072
rect 26879 3008 26880 3072
rect 26814 2992 26880 3008
rect 26814 2928 26815 2992
rect 26879 2928 26880 2992
rect 26814 2904 26880 2928
rect 26814 2848 26819 2904
rect 26875 2848 26880 2904
rect 26814 2838 26880 2848
rect 26940 2774 27000 3804
rect 27060 2834 27120 3866
rect 27180 2774 27240 3804
rect 27300 2834 27360 3866
rect 27420 3712 27486 3866
rect 27420 3648 27421 3712
rect 27485 3648 27486 3712
rect 27420 3632 27486 3648
rect 27420 3568 27421 3632
rect 27485 3568 27486 3632
rect 27420 3552 27486 3568
rect 27420 3488 27421 3552
rect 27485 3488 27486 3552
rect 27420 3472 27486 3488
rect 27420 3408 27421 3472
rect 27485 3408 27486 3472
rect 27420 3392 27486 3408
rect 27420 3328 27421 3392
rect 27485 3328 27486 3392
rect 27420 3312 27486 3328
rect 27420 3248 27421 3312
rect 27485 3248 27486 3312
rect 27420 3232 27486 3248
rect 27420 3168 27421 3232
rect 27485 3168 27486 3232
rect 27420 3152 27486 3168
rect 27420 3088 27421 3152
rect 27485 3088 27486 3152
rect 27420 3072 27486 3088
rect 27420 3008 27421 3072
rect 27485 3008 27486 3072
rect 27420 2992 27486 3008
rect 27420 2928 27421 2992
rect 27485 2928 27486 2992
rect 27420 2904 27486 2928
rect 27420 2848 27425 2904
rect 27481 2848 27486 2904
rect 27420 2838 27486 2848
rect 27546 2774 27606 3804
rect 27666 2834 27726 3866
rect 27786 2774 27846 3804
rect 27906 2834 27966 3866
rect 28026 3712 28092 3866
rect 28026 3648 28027 3712
rect 28091 3648 28092 3712
rect 28026 3632 28092 3648
rect 28026 3568 28027 3632
rect 28091 3568 28092 3632
rect 28026 3552 28092 3568
rect 28026 3488 28027 3552
rect 28091 3488 28092 3552
rect 28026 3472 28092 3488
rect 28026 3408 28027 3472
rect 28091 3408 28092 3472
rect 28026 3392 28092 3408
rect 28026 3328 28027 3392
rect 28091 3328 28092 3392
rect 28026 3312 28092 3328
rect 28026 3248 28027 3312
rect 28091 3248 28092 3312
rect 28026 3232 28092 3248
rect 28026 3168 28027 3232
rect 28091 3168 28092 3232
rect 28026 3152 28092 3168
rect 28026 3088 28027 3152
rect 28091 3088 28092 3152
rect 28026 3072 28092 3088
rect 28026 3008 28027 3072
rect 28091 3008 28092 3072
rect 28026 2992 28092 3008
rect 28026 2928 28027 2992
rect 28091 2928 28092 2992
rect 28026 2904 28092 2928
rect 28026 2848 28031 2904
rect 28087 2848 28092 2904
rect 28026 2838 28092 2848
rect 28152 2774 28212 3804
rect 28272 2834 28332 3866
rect 28392 2774 28452 3804
rect 28512 2834 28572 3866
rect 28632 3712 28698 3866
rect 28632 3648 28633 3712
rect 28697 3648 28698 3712
rect 28632 3632 28698 3648
rect 28632 3568 28633 3632
rect 28697 3568 28698 3632
rect 28632 3552 28698 3568
rect 28632 3488 28633 3552
rect 28697 3488 28698 3552
rect 28632 3472 28698 3488
rect 28632 3408 28633 3472
rect 28697 3408 28698 3472
rect 28632 3392 28698 3408
rect 28632 3328 28633 3392
rect 28697 3328 28698 3392
rect 28632 3312 28698 3328
rect 28632 3248 28633 3312
rect 28697 3248 28698 3312
rect 28632 3232 28698 3248
rect 28632 3168 28633 3232
rect 28697 3168 28698 3232
rect 28632 3152 28698 3168
rect 28632 3088 28633 3152
rect 28697 3088 28698 3152
rect 28632 3072 28698 3088
rect 28632 3008 28633 3072
rect 28697 3008 28698 3072
rect 28632 2992 28698 3008
rect 28632 2928 28633 2992
rect 28697 2928 28698 2992
rect 28632 2904 28698 2928
rect 28632 2848 28637 2904
rect 28693 2848 28698 2904
rect 28632 2838 28698 2848
rect 28758 2774 28818 3804
rect 28878 2834 28938 3866
rect 28998 2774 29058 3804
rect 29118 2834 29178 3866
rect 29238 3712 29304 3866
rect 29238 3648 29239 3712
rect 29303 3648 29304 3712
rect 29238 3632 29304 3648
rect 29238 3568 29239 3632
rect 29303 3568 29304 3632
rect 29238 3552 29304 3568
rect 29238 3488 29239 3552
rect 29303 3488 29304 3552
rect 29238 3472 29304 3488
rect 29238 3408 29239 3472
rect 29303 3408 29304 3472
rect 29238 3392 29304 3408
rect 29238 3328 29239 3392
rect 29303 3328 29304 3392
rect 29238 3312 29304 3328
rect 29238 3248 29239 3312
rect 29303 3248 29304 3312
rect 29238 3232 29304 3248
rect 29238 3168 29239 3232
rect 29303 3168 29304 3232
rect 29238 3152 29304 3168
rect 29238 3088 29239 3152
rect 29303 3088 29304 3152
rect 29238 3072 29304 3088
rect 29238 3008 29239 3072
rect 29303 3008 29304 3072
rect 29238 2992 29304 3008
rect 29238 2928 29239 2992
rect 29303 2928 29304 2992
rect 29238 2838 29304 2928
rect 29364 2774 29424 3804
rect 29484 2834 29544 3866
rect 29604 2774 29664 3804
rect 29724 2834 29784 3866
rect 29844 3712 29910 3866
rect 29844 3648 29845 3712
rect 29909 3648 29910 3712
rect 29844 3632 29910 3648
rect 29844 3568 29845 3632
rect 29909 3568 29910 3632
rect 29844 3552 29910 3568
rect 29844 3488 29845 3552
rect 29909 3488 29910 3552
rect 29844 3472 29910 3488
rect 29844 3408 29845 3472
rect 29909 3408 29910 3472
rect 29844 3392 29910 3408
rect 29844 3328 29845 3392
rect 29909 3328 29910 3392
rect 29844 3312 29910 3328
rect 29844 3248 29845 3312
rect 29909 3248 29910 3312
rect 29844 3232 29910 3248
rect 29844 3168 29845 3232
rect 29909 3168 29910 3232
rect 29844 3152 29910 3168
rect 29844 3088 29845 3152
rect 29909 3088 29910 3152
rect 29844 3072 29910 3088
rect 29844 3008 29845 3072
rect 29909 3008 29910 3072
rect 29844 2992 29910 3008
rect 29844 2928 29845 2992
rect 29909 2928 29910 2992
rect 29844 2838 29910 2928
rect 29970 2774 30030 3804
rect 30090 2834 30150 3866
rect 30210 2774 30270 3804
rect 30330 2834 30390 3866
rect 30450 3712 30516 3866
rect 30450 3648 30451 3712
rect 30515 3648 30516 3712
rect 30450 3632 30516 3648
rect 30450 3568 30451 3632
rect 30515 3568 30516 3632
rect 30450 3552 30516 3568
rect 30450 3488 30451 3552
rect 30515 3488 30516 3552
rect 30450 3472 30516 3488
rect 30450 3408 30451 3472
rect 30515 3408 30516 3472
rect 30450 3392 30516 3408
rect 30450 3328 30451 3392
rect 30515 3328 30516 3392
rect 30450 3312 30516 3328
rect 30450 3248 30451 3312
rect 30515 3248 30516 3312
rect 30450 3232 30516 3248
rect 30450 3168 30451 3232
rect 30515 3168 30516 3232
rect 30450 3152 30516 3168
rect 30450 3088 30451 3152
rect 30515 3088 30516 3152
rect 30450 3072 30516 3088
rect 30450 3008 30451 3072
rect 30515 3008 30516 3072
rect 30450 2992 30516 3008
rect 30450 2928 30451 2992
rect 30515 2928 30516 2992
rect 30450 2838 30516 2928
rect 30576 2774 30636 3804
rect 30696 2834 30756 3866
rect 30816 2774 30876 3804
rect 30936 2834 30996 3866
rect 31056 3712 31122 3866
rect 31056 3648 31057 3712
rect 31121 3648 31122 3712
rect 31056 3632 31122 3648
rect 31056 3568 31057 3632
rect 31121 3568 31122 3632
rect 31056 3552 31122 3568
rect 31056 3488 31057 3552
rect 31121 3488 31122 3552
rect 31056 3472 31122 3488
rect 31056 3408 31057 3472
rect 31121 3408 31122 3472
rect 31056 3392 31122 3408
rect 31056 3328 31057 3392
rect 31121 3328 31122 3392
rect 31056 3312 31122 3328
rect 31056 3248 31057 3312
rect 31121 3248 31122 3312
rect 31056 3232 31122 3248
rect 31056 3168 31057 3232
rect 31121 3168 31122 3232
rect 31056 3152 31122 3168
rect 31056 3088 31057 3152
rect 31121 3088 31122 3152
rect 31056 3072 31122 3088
rect 31056 3008 31057 3072
rect 31121 3008 31122 3072
rect 31056 2992 31122 3008
rect 31056 2928 31057 2992
rect 31121 2928 31122 2992
rect 31056 2838 31122 2928
rect 31182 2774 31242 3804
rect 31302 2834 31362 3866
rect 31422 2774 31482 3804
rect 31542 2834 31602 3866
rect 31662 3712 31728 3866
rect 31662 3648 31663 3712
rect 31727 3648 31728 3712
rect 31662 3632 31728 3648
rect 31662 3568 31663 3632
rect 31727 3568 31728 3632
rect 31662 3552 31728 3568
rect 31662 3488 31663 3552
rect 31727 3488 31728 3552
rect 31662 3472 31728 3488
rect 31662 3408 31663 3472
rect 31727 3408 31728 3472
rect 31662 3392 31728 3408
rect 31662 3328 31663 3392
rect 31727 3328 31728 3392
rect 31662 3312 31728 3328
rect 31662 3248 31663 3312
rect 31727 3248 31728 3312
rect 31662 3232 31728 3248
rect 31662 3168 31663 3232
rect 31727 3168 31728 3232
rect 31662 3152 31728 3168
rect 31662 3088 31663 3152
rect 31727 3088 31728 3152
rect 31662 3072 31728 3088
rect 31662 3008 31663 3072
rect 31727 3008 31728 3072
rect 31662 2992 31728 3008
rect 31662 2928 31663 2992
rect 31727 2928 31728 2992
rect 31662 2838 31728 2928
rect 31788 2774 31848 3804
rect 31908 2834 31968 3866
rect 32028 2774 32088 3804
rect 32148 2834 32208 3866
rect 32268 3712 32334 3866
rect 32268 3648 32269 3712
rect 32333 3648 32334 3712
rect 32268 3632 32334 3648
rect 32268 3568 32269 3632
rect 32333 3568 32334 3632
rect 32268 3552 32334 3568
rect 32268 3488 32269 3552
rect 32333 3488 32334 3552
rect 32268 3472 32334 3488
rect 32268 3408 32269 3472
rect 32333 3408 32334 3472
rect 32268 3392 32334 3408
rect 32268 3328 32269 3392
rect 32333 3328 32334 3392
rect 32268 3312 32334 3328
rect 32268 3248 32269 3312
rect 32333 3248 32334 3312
rect 32268 3232 32334 3248
rect 32268 3168 32269 3232
rect 32333 3168 32334 3232
rect 32268 3152 32334 3168
rect 32268 3088 32269 3152
rect 32333 3088 32334 3152
rect 32268 3072 32334 3088
rect 32268 3008 32269 3072
rect 32333 3008 32334 3072
rect 32268 2992 32334 3008
rect 32268 2928 32269 2992
rect 32333 2928 32334 2992
rect 32268 2838 32334 2928
rect 32394 2774 32454 3804
rect 32514 2834 32574 3866
rect 32634 2774 32694 3804
rect 32754 2834 32814 3866
rect 32874 3712 32940 3866
rect 32874 3648 32875 3712
rect 32939 3648 32940 3712
rect 32874 3632 32940 3648
rect 32874 3568 32875 3632
rect 32939 3568 32940 3632
rect 32874 3552 32940 3568
rect 32874 3488 32875 3552
rect 32939 3488 32940 3552
rect 32874 3472 32940 3488
rect 32874 3408 32875 3472
rect 32939 3408 32940 3472
rect 32874 3392 32940 3408
rect 32874 3328 32875 3392
rect 32939 3328 32940 3392
rect 32874 3312 32940 3328
rect 32874 3248 32875 3312
rect 32939 3248 32940 3312
rect 32874 3232 32940 3248
rect 32874 3168 32875 3232
rect 32939 3168 32940 3232
rect 32874 3152 32940 3168
rect 32874 3088 32875 3152
rect 32939 3088 32940 3152
rect 32874 3072 32940 3088
rect 32874 3008 32875 3072
rect 32939 3008 32940 3072
rect 32874 2992 32940 3008
rect 32874 2928 32875 2992
rect 32939 2928 32940 2992
rect 32874 2838 32940 2928
rect 33000 2774 33060 3804
rect 33120 2834 33180 3866
rect 33240 2774 33300 3804
rect 33360 2834 33420 3866
rect 33480 3712 33546 3866
rect 33480 3648 33481 3712
rect 33545 3648 33546 3712
rect 33480 3632 33546 3648
rect 33480 3568 33481 3632
rect 33545 3568 33546 3632
rect 33480 3552 33546 3568
rect 33480 3488 33481 3552
rect 33545 3488 33546 3552
rect 33480 3472 33546 3488
rect 33480 3408 33481 3472
rect 33545 3408 33546 3472
rect 33480 3392 33546 3408
rect 33480 3328 33481 3392
rect 33545 3328 33546 3392
rect 33480 3312 33546 3328
rect 33480 3248 33481 3312
rect 33545 3248 33546 3312
rect 33480 3232 33546 3248
rect 33480 3168 33481 3232
rect 33545 3168 33546 3232
rect 33480 3152 33546 3168
rect 33480 3088 33481 3152
rect 33545 3088 33546 3152
rect 33480 3072 33546 3088
rect 33480 3008 33481 3072
rect 33545 3008 33546 3072
rect 33480 2992 33546 3008
rect 33480 2928 33481 2992
rect 33545 2928 33546 2992
rect 33480 2838 33546 2928
rect 33606 2774 33666 3804
rect 33726 2834 33786 3866
rect 33846 2774 33906 3804
rect 33966 2834 34026 3866
rect 34086 3712 34152 3866
rect 34086 3648 34087 3712
rect 34151 3648 34152 3712
rect 34086 3632 34152 3648
rect 34086 3568 34087 3632
rect 34151 3568 34152 3632
rect 34086 3552 34152 3568
rect 34086 3488 34087 3552
rect 34151 3488 34152 3552
rect 34086 3472 34152 3488
rect 34086 3408 34087 3472
rect 34151 3408 34152 3472
rect 34086 3392 34152 3408
rect 34086 3328 34087 3392
rect 34151 3328 34152 3392
rect 34086 3312 34152 3328
rect 34086 3248 34087 3312
rect 34151 3248 34152 3312
rect 34086 3232 34152 3248
rect 34086 3168 34087 3232
rect 34151 3168 34152 3232
rect 34086 3152 34152 3168
rect 34086 3088 34087 3152
rect 34151 3088 34152 3152
rect 34086 3072 34152 3088
rect 34086 3008 34087 3072
rect 34151 3008 34152 3072
rect 34086 2992 34152 3008
rect 34086 2928 34087 2992
rect 34151 2928 34152 2992
rect 34086 2838 34152 2928
rect 34212 2774 34272 3804
rect 34332 2834 34392 3866
rect 34452 2774 34512 3804
rect 34572 2834 34632 3866
rect 34692 3712 34758 3866
rect 34692 3648 34693 3712
rect 34757 3648 34758 3712
rect 34692 3632 34758 3648
rect 34692 3568 34693 3632
rect 34757 3568 34758 3632
rect 34692 3552 34758 3568
rect 34692 3488 34693 3552
rect 34757 3488 34758 3552
rect 34692 3472 34758 3488
rect 34692 3408 34693 3472
rect 34757 3408 34758 3472
rect 34692 3392 34758 3408
rect 34692 3328 34693 3392
rect 34757 3328 34758 3392
rect 34692 3312 34758 3328
rect 34692 3248 34693 3312
rect 34757 3248 34758 3312
rect 34692 3232 34758 3248
rect 34692 3168 34693 3232
rect 34757 3168 34758 3232
rect 34692 3152 34758 3168
rect 34692 3088 34693 3152
rect 34757 3088 34758 3152
rect 34692 3072 34758 3088
rect 34692 3008 34693 3072
rect 34757 3008 34758 3072
rect 34692 2992 34758 3008
rect 34692 2928 34693 2992
rect 34757 2928 34758 2992
rect 34692 2838 34758 2928
rect 34818 2774 34878 3804
rect 34938 2834 34998 3866
rect 35058 2774 35118 3804
rect 35178 2834 35238 3866
rect 35298 3712 35364 3866
rect 35298 3648 35299 3712
rect 35363 3648 35364 3712
rect 35298 3632 35364 3648
rect 35298 3568 35299 3632
rect 35363 3568 35364 3632
rect 35298 3552 35364 3568
rect 35298 3488 35299 3552
rect 35363 3488 35364 3552
rect 35298 3472 35364 3488
rect 35298 3408 35299 3472
rect 35363 3408 35364 3472
rect 35298 3392 35364 3408
rect 35298 3328 35299 3392
rect 35363 3328 35364 3392
rect 35298 3312 35364 3328
rect 35298 3248 35299 3312
rect 35363 3248 35364 3312
rect 35298 3232 35364 3248
rect 35298 3168 35299 3232
rect 35363 3168 35364 3232
rect 35298 3152 35364 3168
rect 35298 3088 35299 3152
rect 35363 3088 35364 3152
rect 35298 3072 35364 3088
rect 35298 3008 35299 3072
rect 35363 3008 35364 3072
rect 35298 2992 35364 3008
rect 35298 2928 35299 2992
rect 35363 2928 35364 2992
rect 35298 2838 35364 2928
rect 35424 2774 35484 3804
rect 35544 2834 35604 3866
rect 35664 2774 35724 3804
rect 35784 2834 35844 3866
rect 35904 3712 35970 3866
rect 35904 3648 35905 3712
rect 35969 3648 35970 3712
rect 35904 3632 35970 3648
rect 35904 3568 35905 3632
rect 35969 3568 35970 3632
rect 35904 3552 35970 3568
rect 35904 3488 35905 3552
rect 35969 3488 35970 3552
rect 35904 3472 35970 3488
rect 35904 3408 35905 3472
rect 35969 3408 35970 3472
rect 35904 3392 35970 3408
rect 35904 3328 35905 3392
rect 35969 3328 35970 3392
rect 35904 3312 35970 3328
rect 35904 3248 35905 3312
rect 35969 3248 35970 3312
rect 35904 3232 35970 3248
rect 35904 3168 35905 3232
rect 35969 3168 35970 3232
rect 35904 3152 35970 3168
rect 35904 3088 35905 3152
rect 35969 3088 35970 3152
rect 35904 3072 35970 3088
rect 35904 3008 35905 3072
rect 35969 3008 35970 3072
rect 35904 2992 35970 3008
rect 35904 2928 35905 2992
rect 35969 2928 35970 2992
rect 35904 2838 35970 2928
rect 36030 2774 36090 3804
rect 36150 2834 36210 3866
rect 36270 2774 36330 3804
rect 36390 2834 36450 3866
rect 36510 3712 36576 3866
rect 36510 3648 36511 3712
rect 36575 3648 36576 3712
rect 36510 3632 36576 3648
rect 36510 3568 36511 3632
rect 36575 3568 36576 3632
rect 36510 3552 36576 3568
rect 36510 3488 36511 3552
rect 36575 3488 36576 3552
rect 36510 3472 36576 3488
rect 36510 3408 36511 3472
rect 36575 3408 36576 3472
rect 36510 3392 36576 3408
rect 36510 3328 36511 3392
rect 36575 3328 36576 3392
rect 36510 3312 36576 3328
rect 36510 3248 36511 3312
rect 36575 3248 36576 3312
rect 36510 3232 36576 3248
rect 36510 3168 36511 3232
rect 36575 3168 36576 3232
rect 36510 3152 36576 3168
rect 36510 3088 36511 3152
rect 36575 3088 36576 3152
rect 36510 3072 36576 3088
rect 36510 3008 36511 3072
rect 36575 3008 36576 3072
rect 36510 2992 36576 3008
rect 36510 2928 36511 2992
rect 36575 2928 36576 2992
rect 36510 2838 36576 2928
rect 36636 2774 36696 3804
rect 36756 2834 36816 3866
rect 36876 2774 36936 3804
rect 36996 2834 37056 3866
rect 37116 3712 37182 3866
rect 37116 3648 37117 3712
rect 37181 3648 37182 3712
rect 37116 3632 37182 3648
rect 37116 3568 37117 3632
rect 37181 3568 37182 3632
rect 37116 3552 37182 3568
rect 37116 3488 37117 3552
rect 37181 3488 37182 3552
rect 37116 3472 37182 3488
rect 37116 3408 37117 3472
rect 37181 3408 37182 3472
rect 37116 3392 37182 3408
rect 37116 3328 37117 3392
rect 37181 3328 37182 3392
rect 37116 3312 37182 3328
rect 37116 3248 37117 3312
rect 37181 3248 37182 3312
rect 37116 3232 37182 3248
rect 37116 3168 37117 3232
rect 37181 3168 37182 3232
rect 37116 3152 37182 3168
rect 37116 3088 37117 3152
rect 37181 3088 37182 3152
rect 37116 3072 37182 3088
rect 37116 3008 37117 3072
rect 37181 3008 37182 3072
rect 37116 2992 37182 3008
rect 37116 2928 37117 2992
rect 37181 2928 37182 2992
rect 37116 2838 37182 2928
rect 37242 2774 37302 3804
rect 37362 2834 37422 3866
rect 37482 2774 37542 3804
rect 37602 2834 37662 3866
rect 37722 3712 37788 3866
rect 37722 3648 37723 3712
rect 37787 3648 37788 3712
rect 37722 3632 37788 3648
rect 37722 3568 37723 3632
rect 37787 3568 37788 3632
rect 37722 3552 37788 3568
rect 37722 3488 37723 3552
rect 37787 3488 37788 3552
rect 37722 3472 37788 3488
rect 37722 3408 37723 3472
rect 37787 3408 37788 3472
rect 37722 3392 37788 3408
rect 37722 3328 37723 3392
rect 37787 3328 37788 3392
rect 37722 3312 37788 3328
rect 37722 3248 37723 3312
rect 37787 3248 37788 3312
rect 37722 3232 37788 3248
rect 37722 3168 37723 3232
rect 37787 3168 37788 3232
rect 37722 3152 37788 3168
rect 37722 3088 37723 3152
rect 37787 3088 37788 3152
rect 37722 3072 37788 3088
rect 37722 3008 37723 3072
rect 37787 3008 37788 3072
rect 37722 2992 37788 3008
rect 37722 2928 37723 2992
rect 37787 2928 37788 2992
rect 37722 2838 37788 2928
rect 37848 2774 37908 3804
rect 37968 2834 38028 3866
rect 38088 2774 38148 3804
rect 38208 2834 38268 3866
rect 38328 3712 38394 3866
rect 38328 3648 38329 3712
rect 38393 3648 38394 3712
rect 38328 3632 38394 3648
rect 38328 3568 38329 3632
rect 38393 3568 38394 3632
rect 38328 3552 38394 3568
rect 38328 3488 38329 3552
rect 38393 3488 38394 3552
rect 38328 3472 38394 3488
rect 38328 3408 38329 3472
rect 38393 3408 38394 3472
rect 38328 3392 38394 3408
rect 38328 3328 38329 3392
rect 38393 3328 38394 3392
rect 38328 3312 38394 3328
rect 38328 3248 38329 3312
rect 38393 3248 38394 3312
rect 38328 3232 38394 3248
rect 38328 3168 38329 3232
rect 38393 3168 38394 3232
rect 38328 3152 38394 3168
rect 38328 3088 38329 3152
rect 38393 3088 38394 3152
rect 38328 3072 38394 3088
rect 38328 3008 38329 3072
rect 38393 3008 38394 3072
rect 38328 2992 38394 3008
rect 38328 2928 38329 2992
rect 38393 2928 38394 2992
rect 38328 2838 38394 2928
rect 38454 2774 38514 3804
rect 38574 2834 38634 3866
rect 38694 2774 38754 3804
rect 38814 2834 38874 3866
rect 38934 3712 39000 3866
rect 38934 3648 38935 3712
rect 38999 3648 39000 3712
rect 38934 3632 39000 3648
rect 38934 3568 38935 3632
rect 38999 3568 39000 3632
rect 38934 3552 39000 3568
rect 38934 3488 38935 3552
rect 38999 3488 39000 3552
rect 38934 3472 39000 3488
rect 38934 3408 38935 3472
rect 38999 3408 39000 3472
rect 38934 3392 39000 3408
rect 38934 3328 38935 3392
rect 38999 3328 39000 3392
rect 38934 3312 39000 3328
rect 38934 3248 38935 3312
rect 38999 3248 39000 3312
rect 38934 3232 39000 3248
rect 38934 3168 38935 3232
rect 38999 3168 39000 3232
rect 38934 3152 39000 3168
rect 38934 3088 38935 3152
rect 38999 3088 39000 3152
rect 38934 3072 39000 3088
rect 38934 3008 38935 3072
rect 38999 3008 39000 3072
rect 38934 2992 39000 3008
rect 38934 2928 38935 2992
rect 38999 2928 39000 2992
rect 38934 2838 39000 2928
rect 39060 2774 39120 3804
rect 39180 2834 39240 3866
rect 39300 2774 39360 3804
rect 39420 2834 39480 3866
rect 39540 3712 39606 3866
rect 39540 3648 39541 3712
rect 39605 3648 39606 3712
rect 39540 3632 39606 3648
rect 39540 3568 39541 3632
rect 39605 3568 39606 3632
rect 39540 3552 39606 3568
rect 39540 3488 39541 3552
rect 39605 3488 39606 3552
rect 39540 3472 39606 3488
rect 39540 3408 39541 3472
rect 39605 3408 39606 3472
rect 39540 3392 39606 3408
rect 39540 3328 39541 3392
rect 39605 3328 39606 3392
rect 39540 3312 39606 3328
rect 39540 3248 39541 3312
rect 39605 3248 39606 3312
rect 39540 3232 39606 3248
rect 39540 3168 39541 3232
rect 39605 3168 39606 3232
rect 39540 3152 39606 3168
rect 39540 3088 39541 3152
rect 39605 3088 39606 3152
rect 39540 3072 39606 3088
rect 39540 3008 39541 3072
rect 39605 3008 39606 3072
rect 39540 2992 39606 3008
rect 39540 2928 39541 2992
rect 39605 2928 39606 2992
rect 39540 2838 39606 2928
rect -459 2772 213 2774
rect -459 2708 -355 2772
rect -291 2708 -275 2772
rect -211 2708 -195 2772
rect -131 2708 -115 2772
rect -51 2708 -35 2772
rect 29 2708 45 2772
rect 109 2708 213 2772
rect -459 2706 213 2708
rect 355 2772 1027 2774
rect 355 2708 459 2772
rect 523 2708 539 2772
rect 603 2708 619 2772
rect 683 2708 699 2772
rect 763 2708 779 2772
rect 843 2708 859 2772
rect 923 2708 1027 2772
rect 355 2706 1027 2708
rect 1267 2772 2545 2774
rect 1267 2708 1371 2772
rect 1435 2708 1451 2772
rect 1515 2708 1531 2772
rect 1595 2708 1611 2772
rect 1675 2708 1691 2772
rect 1755 2708 1771 2772
rect 1835 2708 1977 2772
rect 2041 2708 2057 2772
rect 2121 2708 2137 2772
rect 2201 2708 2217 2772
rect 2281 2708 2297 2772
rect 2361 2708 2377 2772
rect 2441 2708 2545 2772
rect 1267 2706 2545 2708
rect 2801 2772 5291 2774
rect 2801 2708 2905 2772
rect 2969 2708 2985 2772
rect 3049 2708 3065 2772
rect 3129 2708 3145 2772
rect 3209 2708 3225 2772
rect 3289 2708 3305 2772
rect 3369 2708 3511 2772
rect 3575 2708 3591 2772
rect 3655 2708 3671 2772
rect 3735 2708 3751 2772
rect 3815 2708 3831 2772
rect 3895 2708 3911 2772
rect 3975 2708 4117 2772
rect 4181 2708 4197 2772
rect 4261 2708 4277 2772
rect 4341 2708 4357 2772
rect 4421 2708 4437 2772
rect 4501 2708 4517 2772
rect 4581 2708 4723 2772
rect 4787 2708 4803 2772
rect 4867 2708 4883 2772
rect 4947 2708 4963 2772
rect 5027 2708 5043 2772
rect 5107 2708 5123 2772
rect 5187 2708 5291 2772
rect 2801 2706 5291 2708
rect 5352 2772 10266 2774
rect 5352 2708 5456 2772
rect 5520 2708 5536 2772
rect 5600 2708 5616 2772
rect 5680 2708 5696 2772
rect 5760 2708 5776 2772
rect 5840 2708 5856 2772
rect 5920 2708 6062 2772
rect 6126 2708 6142 2772
rect 6206 2708 6222 2772
rect 6286 2708 6302 2772
rect 6366 2708 6382 2772
rect 6446 2708 6462 2772
rect 6526 2708 6668 2772
rect 6732 2708 6748 2772
rect 6812 2708 6828 2772
rect 6892 2708 6908 2772
rect 6972 2708 6988 2772
rect 7052 2708 7068 2772
rect 7132 2708 7274 2772
rect 7338 2708 7354 2772
rect 7418 2708 7434 2772
rect 7498 2708 7514 2772
rect 7578 2708 7594 2772
rect 7658 2708 7674 2772
rect 7738 2708 7880 2772
rect 7944 2708 7960 2772
rect 8024 2708 8040 2772
rect 8104 2708 8120 2772
rect 8184 2708 8200 2772
rect 8264 2708 8280 2772
rect 8344 2708 8486 2772
rect 8550 2708 8566 2772
rect 8630 2708 8646 2772
rect 8710 2708 8726 2772
rect 8790 2708 8806 2772
rect 8870 2708 8886 2772
rect 8950 2708 9092 2772
rect 9156 2708 9172 2772
rect 9236 2708 9252 2772
rect 9316 2708 9332 2772
rect 9396 2708 9412 2772
rect 9476 2708 9492 2772
rect 9556 2708 9698 2772
rect 9762 2708 9778 2772
rect 9842 2708 9858 2772
rect 9922 2708 9938 2772
rect 10002 2708 10018 2772
rect 10082 2708 10098 2772
rect 10162 2708 10266 2772
rect 5352 2706 10266 2708
rect 10326 2772 20088 2774
rect 10326 2708 10430 2772
rect 10494 2708 10510 2772
rect 10574 2708 10590 2772
rect 10654 2708 10670 2772
rect 10734 2708 10750 2772
rect 10814 2708 10830 2772
rect 10894 2708 11036 2772
rect 11100 2708 11116 2772
rect 11180 2708 11196 2772
rect 11260 2708 11276 2772
rect 11340 2708 11356 2772
rect 11420 2708 11436 2772
rect 11500 2708 11642 2772
rect 11706 2708 11722 2772
rect 11786 2708 11802 2772
rect 11866 2708 11882 2772
rect 11946 2708 11962 2772
rect 12026 2708 12042 2772
rect 12106 2708 12248 2772
rect 12312 2708 12328 2772
rect 12392 2708 12408 2772
rect 12472 2708 12488 2772
rect 12552 2708 12568 2772
rect 12632 2708 12648 2772
rect 12712 2708 12854 2772
rect 12918 2708 12934 2772
rect 12998 2708 13014 2772
rect 13078 2708 13094 2772
rect 13158 2708 13174 2772
rect 13238 2708 13254 2772
rect 13318 2708 13460 2772
rect 13524 2708 13540 2772
rect 13604 2708 13620 2772
rect 13684 2708 13700 2772
rect 13764 2708 13780 2772
rect 13844 2708 13860 2772
rect 13924 2708 14066 2772
rect 14130 2708 14146 2772
rect 14210 2708 14226 2772
rect 14290 2708 14306 2772
rect 14370 2708 14386 2772
rect 14450 2708 14466 2772
rect 14530 2708 14672 2772
rect 14736 2708 14752 2772
rect 14816 2708 14832 2772
rect 14896 2708 14912 2772
rect 14976 2708 14992 2772
rect 15056 2708 15072 2772
rect 15136 2708 15278 2772
rect 15342 2708 15358 2772
rect 15422 2708 15438 2772
rect 15502 2708 15518 2772
rect 15582 2708 15598 2772
rect 15662 2708 15678 2772
rect 15742 2708 15884 2772
rect 15948 2708 15964 2772
rect 16028 2708 16044 2772
rect 16108 2708 16124 2772
rect 16188 2708 16204 2772
rect 16268 2708 16284 2772
rect 16348 2708 16490 2772
rect 16554 2708 16570 2772
rect 16634 2708 16650 2772
rect 16714 2708 16730 2772
rect 16794 2708 16810 2772
rect 16874 2708 16890 2772
rect 16954 2708 17096 2772
rect 17160 2708 17176 2772
rect 17240 2708 17256 2772
rect 17320 2708 17336 2772
rect 17400 2708 17416 2772
rect 17480 2708 17496 2772
rect 17560 2708 17702 2772
rect 17766 2708 17782 2772
rect 17846 2708 17862 2772
rect 17926 2708 17942 2772
rect 18006 2708 18022 2772
rect 18086 2708 18102 2772
rect 18166 2708 18308 2772
rect 18372 2708 18388 2772
rect 18452 2708 18468 2772
rect 18532 2708 18548 2772
rect 18612 2708 18628 2772
rect 18692 2708 18708 2772
rect 18772 2708 18914 2772
rect 18978 2708 18994 2772
rect 19058 2708 19074 2772
rect 19138 2708 19154 2772
rect 19218 2708 19234 2772
rect 19298 2708 19314 2772
rect 19378 2708 19520 2772
rect 19584 2708 19600 2772
rect 19664 2708 19680 2772
rect 19744 2708 19760 2772
rect 19824 2708 19840 2772
rect 19904 2708 19920 2772
rect 19984 2708 20088 2772
rect 10326 2706 20088 2708
rect 20148 2772 39606 2774
rect 20148 2708 20252 2772
rect 20316 2708 20332 2772
rect 20396 2708 20412 2772
rect 20476 2708 20492 2772
rect 20556 2708 20572 2772
rect 20636 2708 20652 2772
rect 20716 2708 20858 2772
rect 20922 2708 20938 2772
rect 21002 2708 21018 2772
rect 21082 2708 21098 2772
rect 21162 2708 21178 2772
rect 21242 2708 21258 2772
rect 21322 2708 21464 2772
rect 21528 2708 21544 2772
rect 21608 2708 21624 2772
rect 21688 2708 21704 2772
rect 21768 2708 21784 2772
rect 21848 2708 21864 2772
rect 21928 2708 22070 2772
rect 22134 2708 22150 2772
rect 22214 2708 22230 2772
rect 22294 2708 22310 2772
rect 22374 2708 22390 2772
rect 22454 2708 22470 2772
rect 22534 2708 22676 2772
rect 22740 2708 22756 2772
rect 22820 2708 22836 2772
rect 22900 2708 22916 2772
rect 22980 2708 22996 2772
rect 23060 2708 23076 2772
rect 23140 2708 23282 2772
rect 23346 2708 23362 2772
rect 23426 2708 23442 2772
rect 23506 2708 23522 2772
rect 23586 2708 23602 2772
rect 23666 2708 23682 2772
rect 23746 2708 23888 2772
rect 23952 2708 23968 2772
rect 24032 2708 24048 2772
rect 24112 2708 24128 2772
rect 24192 2708 24208 2772
rect 24272 2708 24288 2772
rect 24352 2708 24494 2772
rect 24558 2708 24574 2772
rect 24638 2708 24654 2772
rect 24718 2708 24734 2772
rect 24798 2708 24814 2772
rect 24878 2708 24894 2772
rect 24958 2708 25100 2772
rect 25164 2708 25180 2772
rect 25244 2708 25260 2772
rect 25324 2708 25340 2772
rect 25404 2708 25420 2772
rect 25484 2708 25500 2772
rect 25564 2708 25706 2772
rect 25770 2708 25786 2772
rect 25850 2708 25866 2772
rect 25930 2708 25946 2772
rect 26010 2708 26026 2772
rect 26090 2708 26106 2772
rect 26170 2708 26312 2772
rect 26376 2708 26392 2772
rect 26456 2708 26472 2772
rect 26536 2708 26552 2772
rect 26616 2708 26632 2772
rect 26696 2708 26712 2772
rect 26776 2708 26918 2772
rect 26982 2708 26998 2772
rect 27062 2708 27078 2772
rect 27142 2708 27158 2772
rect 27222 2708 27238 2772
rect 27302 2708 27318 2772
rect 27382 2708 27524 2772
rect 27588 2708 27604 2772
rect 27668 2708 27684 2772
rect 27748 2708 27764 2772
rect 27828 2708 27844 2772
rect 27908 2708 27924 2772
rect 27988 2708 28130 2772
rect 28194 2708 28210 2772
rect 28274 2708 28290 2772
rect 28354 2708 28370 2772
rect 28434 2708 28450 2772
rect 28514 2708 28530 2772
rect 28594 2708 28736 2772
rect 28800 2708 28816 2772
rect 28880 2708 28896 2772
rect 28960 2708 28976 2772
rect 29040 2708 29056 2772
rect 29120 2708 29136 2772
rect 29200 2708 29342 2772
rect 29406 2708 29422 2772
rect 29486 2708 29502 2772
rect 29566 2708 29582 2772
rect 29646 2708 29662 2772
rect 29726 2708 29742 2772
rect 29806 2708 29948 2772
rect 30012 2708 30028 2772
rect 30092 2708 30108 2772
rect 30172 2708 30188 2772
rect 30252 2708 30268 2772
rect 30332 2708 30348 2772
rect 30412 2708 30554 2772
rect 30618 2708 30634 2772
rect 30698 2708 30714 2772
rect 30778 2708 30794 2772
rect 30858 2708 30874 2772
rect 30938 2708 30954 2772
rect 31018 2708 31160 2772
rect 31224 2708 31240 2772
rect 31304 2708 31320 2772
rect 31384 2708 31400 2772
rect 31464 2708 31480 2772
rect 31544 2708 31560 2772
rect 31624 2708 31766 2772
rect 31830 2708 31846 2772
rect 31910 2708 31926 2772
rect 31990 2708 32006 2772
rect 32070 2708 32086 2772
rect 32150 2708 32166 2772
rect 32230 2708 32372 2772
rect 32436 2708 32452 2772
rect 32516 2708 32532 2772
rect 32596 2708 32612 2772
rect 32676 2708 32692 2772
rect 32756 2708 32772 2772
rect 32836 2708 32978 2772
rect 33042 2708 33058 2772
rect 33122 2708 33138 2772
rect 33202 2708 33218 2772
rect 33282 2708 33298 2772
rect 33362 2708 33378 2772
rect 33442 2708 33584 2772
rect 33648 2708 33664 2772
rect 33728 2708 33744 2772
rect 33808 2708 33824 2772
rect 33888 2708 33904 2772
rect 33968 2708 33984 2772
rect 34048 2708 34190 2772
rect 34254 2708 34270 2772
rect 34334 2708 34350 2772
rect 34414 2708 34430 2772
rect 34494 2708 34510 2772
rect 34574 2708 34590 2772
rect 34654 2708 34796 2772
rect 34860 2708 34876 2772
rect 34940 2708 34956 2772
rect 35020 2708 35036 2772
rect 35100 2708 35116 2772
rect 35180 2708 35196 2772
rect 35260 2708 35402 2772
rect 35466 2708 35482 2772
rect 35546 2708 35562 2772
rect 35626 2708 35642 2772
rect 35706 2708 35722 2772
rect 35786 2708 35802 2772
rect 35866 2708 36008 2772
rect 36072 2708 36088 2772
rect 36152 2708 36168 2772
rect 36232 2708 36248 2772
rect 36312 2708 36328 2772
rect 36392 2708 36408 2772
rect 36472 2708 36614 2772
rect 36678 2708 36694 2772
rect 36758 2708 36774 2772
rect 36838 2708 36854 2772
rect 36918 2708 36934 2772
rect 36998 2708 37014 2772
rect 37078 2708 37220 2772
rect 37284 2708 37300 2772
rect 37364 2708 37380 2772
rect 37444 2708 37460 2772
rect 37524 2708 37540 2772
rect 37604 2708 37620 2772
rect 37684 2708 37826 2772
rect 37890 2708 37906 2772
rect 37970 2708 37986 2772
rect 38050 2708 38066 2772
rect 38130 2708 38146 2772
rect 38210 2708 38226 2772
rect 38290 2708 38432 2772
rect 38496 2708 38512 2772
rect 38576 2708 38592 2772
rect 38656 2708 38672 2772
rect 38736 2708 38752 2772
rect 38816 2708 38832 2772
rect 38896 2708 39038 2772
rect 39102 2708 39118 2772
rect 39182 2708 39198 2772
rect 39262 2708 39278 2772
rect 39342 2708 39358 2772
rect 39422 2708 39438 2772
rect 39502 2708 39606 2772
rect 20148 2706 39606 2708
rect -459 1959 213 1961
rect -459 1895 -355 1959
rect -291 1895 -275 1959
rect -211 1895 -195 1959
rect -131 1895 -115 1959
rect -51 1956 -35 1959
rect -51 1895 -35 1900
rect 29 1895 45 1959
rect 109 1895 213 1959
rect -459 1893 213 1895
rect 355 1959 1027 1961
rect 355 1895 459 1959
rect 523 1895 539 1959
rect 603 1895 619 1959
rect 683 1895 699 1959
rect 763 1895 779 1959
rect 843 1895 859 1959
rect 923 1895 1027 1959
rect 355 1893 1027 1895
rect 1267 1959 2545 1961
rect 1267 1895 1371 1959
rect 1435 1895 1451 1959
rect 1515 1895 1531 1959
rect 1595 1895 1611 1959
rect 1675 1895 1691 1959
rect 1755 1895 1771 1959
rect 1835 1895 1977 1959
rect 2041 1895 2057 1959
rect 2121 1895 2137 1959
rect 2201 1895 2217 1959
rect 2281 1895 2297 1959
rect 2361 1895 2377 1959
rect 2441 1895 2545 1959
rect 1267 1893 2545 1895
rect 2801 1959 5291 1961
rect 2801 1895 2905 1959
rect 2969 1895 2985 1959
rect 3049 1895 3065 1959
rect 3129 1895 3145 1959
rect 3209 1895 3225 1959
rect 3289 1895 3305 1959
rect 3369 1895 3511 1959
rect 3575 1895 3591 1959
rect 3655 1895 3671 1959
rect 3735 1895 3751 1959
rect 3815 1895 3831 1959
rect 3895 1895 3911 1959
rect 3975 1895 4117 1959
rect 4181 1895 4197 1959
rect 4261 1895 4277 1959
rect 4341 1895 4357 1959
rect 4421 1895 4437 1959
rect 4501 1895 4517 1959
rect 4581 1895 4723 1959
rect 4787 1895 4803 1959
rect 4867 1895 4883 1959
rect 4947 1895 4963 1959
rect 5027 1895 5043 1959
rect 5107 1895 5123 1959
rect 5187 1895 5291 1959
rect 2801 1893 5291 1895
rect 5352 1959 10266 1961
rect 5352 1895 5456 1959
rect 5520 1895 5536 1959
rect 5600 1895 5616 1959
rect 5680 1895 5696 1959
rect 5760 1895 5776 1959
rect 5840 1895 5856 1959
rect 5920 1895 6062 1959
rect 6126 1895 6142 1959
rect 6206 1895 6222 1959
rect 6286 1895 6302 1959
rect 6366 1895 6382 1959
rect 6446 1895 6462 1959
rect 6526 1895 6668 1959
rect 6732 1895 6748 1959
rect 6812 1895 6828 1959
rect 6892 1895 6908 1959
rect 6972 1895 6988 1959
rect 7052 1895 7068 1959
rect 7132 1895 7274 1959
rect 7338 1895 7354 1959
rect 7418 1895 7434 1959
rect 7498 1895 7514 1959
rect 7578 1895 7594 1959
rect 7658 1895 7674 1959
rect 7738 1895 7880 1959
rect 7944 1895 7960 1959
rect 8024 1895 8040 1959
rect 8104 1895 8120 1959
rect 8184 1895 8200 1959
rect 8264 1895 8280 1959
rect 8344 1895 8486 1959
rect 8550 1895 8566 1959
rect 8630 1895 8646 1959
rect 8710 1895 8726 1959
rect 8790 1895 8806 1959
rect 8870 1895 8886 1959
rect 8950 1895 9092 1959
rect 9156 1895 9172 1959
rect 9236 1895 9252 1959
rect 9316 1895 9332 1959
rect 9396 1895 9412 1959
rect 9476 1895 9492 1959
rect 9556 1895 9698 1959
rect 9762 1895 9778 1959
rect 9842 1895 9858 1959
rect 9922 1895 9938 1959
rect 10002 1895 10018 1959
rect 10082 1895 10098 1959
rect 10162 1895 10266 1959
rect 5352 1893 10266 1895
rect 10326 1959 20088 1961
rect 10326 1895 10430 1959
rect 10494 1895 10510 1959
rect 10574 1895 10590 1959
rect 10654 1895 10670 1959
rect 10734 1895 10750 1959
rect 10814 1895 10830 1959
rect 10894 1895 11036 1959
rect 11100 1895 11116 1959
rect 11180 1895 11196 1959
rect 11260 1895 11276 1959
rect 11340 1895 11356 1959
rect 11420 1895 11436 1959
rect 11500 1895 11642 1959
rect 11706 1895 11722 1959
rect 11786 1895 11802 1959
rect 11866 1895 11882 1959
rect 11946 1895 11962 1959
rect 12026 1895 12042 1959
rect 12106 1895 12248 1959
rect 12312 1895 12328 1959
rect 12392 1895 12408 1959
rect 12472 1895 12488 1959
rect 12552 1895 12568 1959
rect 12632 1895 12648 1959
rect 12712 1895 12854 1959
rect 12918 1895 12934 1959
rect 12998 1895 13014 1959
rect 13078 1895 13094 1959
rect 13158 1895 13174 1959
rect 13238 1895 13254 1959
rect 13318 1895 13460 1959
rect 13524 1895 13540 1959
rect 13604 1895 13620 1959
rect 13684 1895 13700 1959
rect 13764 1895 13780 1959
rect 13844 1895 13860 1959
rect 13924 1895 14066 1959
rect 14130 1895 14146 1959
rect 14210 1895 14226 1959
rect 14290 1895 14306 1959
rect 14370 1895 14386 1959
rect 14450 1895 14466 1959
rect 14530 1895 14672 1959
rect 14736 1895 14752 1959
rect 14816 1895 14832 1959
rect 14896 1895 14912 1959
rect 14976 1895 14992 1959
rect 15056 1895 15072 1959
rect 15136 1895 15278 1959
rect 15342 1895 15358 1959
rect 15422 1895 15438 1959
rect 15502 1895 15518 1959
rect 15582 1895 15598 1959
rect 15662 1895 15678 1959
rect 15742 1895 15884 1959
rect 15948 1895 15964 1959
rect 16028 1895 16044 1959
rect 16108 1895 16124 1959
rect 16188 1895 16204 1959
rect 16268 1895 16284 1959
rect 16348 1895 16490 1959
rect 16554 1895 16570 1959
rect 16634 1895 16650 1959
rect 16714 1895 16730 1959
rect 16794 1895 16810 1959
rect 16874 1895 16890 1959
rect 16954 1895 17096 1959
rect 17160 1895 17176 1959
rect 17240 1895 17256 1959
rect 17320 1895 17336 1959
rect 17400 1895 17416 1959
rect 17480 1895 17496 1959
rect 17560 1895 17702 1959
rect 17766 1895 17782 1959
rect 17846 1895 17862 1959
rect 17926 1895 17942 1959
rect 18006 1895 18022 1959
rect 18086 1895 18102 1959
rect 18166 1895 18308 1959
rect 18372 1895 18388 1959
rect 18452 1895 18468 1959
rect 18532 1895 18548 1959
rect 18612 1895 18628 1959
rect 18692 1895 18708 1959
rect 18772 1895 18914 1959
rect 18978 1895 18994 1959
rect 19058 1895 19074 1959
rect 19138 1895 19154 1959
rect 19218 1895 19234 1959
rect 19298 1895 19314 1959
rect 19378 1895 19520 1959
rect 19584 1895 19600 1959
rect 19664 1895 19680 1959
rect 19744 1895 19760 1959
rect 19824 1895 19840 1959
rect 19904 1895 19920 1959
rect 19984 1895 20088 1959
rect 10326 1893 20088 1895
rect 20148 1959 39606 1961
rect 20148 1895 20252 1959
rect 20316 1895 20332 1959
rect 20396 1895 20412 1959
rect 20476 1895 20492 1959
rect 20556 1895 20572 1959
rect 20636 1895 20652 1959
rect 20716 1895 20858 1959
rect 20922 1895 20938 1959
rect 21002 1895 21018 1959
rect 21082 1895 21098 1959
rect 21162 1895 21178 1959
rect 21242 1895 21258 1959
rect 21322 1895 21464 1959
rect 21528 1895 21544 1959
rect 21608 1895 21624 1959
rect 21688 1895 21704 1959
rect 21768 1895 21784 1959
rect 21848 1895 21864 1959
rect 21928 1895 22070 1959
rect 22134 1895 22150 1959
rect 22214 1895 22230 1959
rect 22294 1895 22310 1959
rect 22374 1895 22390 1959
rect 22454 1895 22470 1959
rect 22534 1895 22676 1959
rect 22740 1895 22756 1959
rect 22820 1895 22836 1959
rect 22900 1895 22916 1959
rect 22980 1895 22996 1959
rect 23060 1895 23076 1959
rect 23140 1895 23282 1959
rect 23346 1895 23362 1959
rect 23426 1895 23442 1959
rect 23506 1895 23522 1959
rect 23586 1895 23602 1959
rect 23666 1895 23682 1959
rect 23746 1895 23888 1959
rect 23952 1895 23968 1959
rect 24032 1895 24048 1959
rect 24112 1895 24128 1959
rect 24192 1895 24208 1959
rect 24272 1895 24288 1959
rect 24352 1895 24494 1959
rect 24558 1895 24574 1959
rect 24638 1895 24654 1959
rect 24718 1895 24734 1959
rect 24798 1895 24814 1959
rect 24878 1895 24894 1959
rect 24958 1895 25100 1959
rect 25164 1895 25180 1959
rect 25244 1895 25260 1959
rect 25324 1895 25340 1959
rect 25404 1895 25420 1959
rect 25484 1895 25500 1959
rect 25564 1895 25706 1959
rect 25770 1895 25786 1959
rect 25850 1895 25866 1959
rect 25930 1895 25946 1959
rect 26010 1895 26026 1959
rect 26090 1895 26106 1959
rect 26170 1895 26312 1959
rect 26376 1895 26392 1959
rect 26456 1895 26472 1959
rect 26536 1895 26552 1959
rect 26616 1895 26632 1959
rect 26696 1895 26712 1959
rect 26776 1895 26918 1959
rect 26982 1895 26998 1959
rect 27062 1895 27078 1959
rect 27142 1895 27158 1959
rect 27222 1895 27238 1959
rect 27302 1895 27318 1959
rect 27382 1895 27524 1959
rect 27588 1895 27604 1959
rect 27668 1895 27684 1959
rect 27748 1895 27764 1959
rect 27828 1895 27844 1959
rect 27908 1895 27924 1959
rect 27988 1895 28130 1959
rect 28194 1895 28210 1959
rect 28274 1895 28290 1959
rect 28354 1895 28370 1959
rect 28434 1895 28450 1959
rect 28514 1895 28530 1959
rect 28594 1895 28736 1959
rect 28800 1895 28816 1959
rect 28880 1895 28896 1959
rect 28960 1895 28976 1959
rect 29040 1895 29056 1959
rect 29120 1895 29136 1959
rect 29200 1895 29342 1959
rect 29406 1895 29422 1959
rect 29486 1895 29502 1959
rect 29566 1895 29582 1959
rect 29646 1895 29662 1959
rect 29726 1895 29742 1959
rect 29806 1895 29948 1959
rect 30012 1895 30028 1959
rect 30092 1895 30108 1959
rect 30172 1895 30188 1959
rect 30252 1895 30268 1959
rect 30332 1895 30348 1959
rect 30412 1895 30554 1959
rect 30618 1895 30634 1959
rect 30698 1895 30714 1959
rect 30778 1895 30794 1959
rect 30858 1895 30874 1959
rect 30938 1895 30954 1959
rect 31018 1895 31160 1959
rect 31224 1895 31240 1959
rect 31304 1895 31320 1959
rect 31384 1895 31400 1959
rect 31464 1895 31480 1959
rect 31544 1895 31560 1959
rect 31624 1895 31766 1959
rect 31830 1895 31846 1959
rect 31910 1895 31926 1959
rect 31990 1895 32006 1959
rect 32070 1895 32086 1959
rect 32150 1895 32166 1959
rect 32230 1895 32372 1959
rect 32436 1895 32452 1959
rect 32516 1895 32532 1959
rect 32596 1895 32612 1959
rect 32676 1895 32692 1959
rect 32756 1895 32772 1959
rect 32836 1895 32978 1959
rect 33042 1895 33058 1959
rect 33122 1895 33138 1959
rect 33202 1895 33218 1959
rect 33282 1895 33298 1959
rect 33362 1895 33378 1959
rect 33442 1895 33584 1959
rect 33648 1895 33664 1959
rect 33728 1895 33744 1959
rect 33808 1895 33824 1959
rect 33888 1895 33904 1959
rect 33968 1895 33984 1959
rect 34048 1895 34190 1959
rect 34254 1895 34270 1959
rect 34334 1895 34350 1959
rect 34414 1895 34430 1959
rect 34494 1895 34510 1959
rect 34574 1895 34590 1959
rect 34654 1895 34796 1959
rect 34860 1895 34876 1959
rect 34940 1895 34956 1959
rect 35020 1895 35036 1959
rect 35100 1895 35116 1959
rect 35180 1895 35196 1959
rect 35260 1895 35402 1959
rect 35466 1895 35482 1959
rect 35546 1895 35562 1959
rect 35626 1895 35642 1959
rect 35706 1895 35722 1959
rect 35786 1895 35802 1959
rect 35866 1895 36008 1959
rect 36072 1895 36088 1959
rect 36152 1895 36168 1959
rect 36232 1895 36248 1959
rect 36312 1895 36328 1959
rect 36392 1895 36408 1959
rect 36472 1895 36614 1959
rect 36678 1895 36694 1959
rect 36758 1895 36774 1959
rect 36838 1895 36854 1959
rect 36918 1895 36934 1959
rect 36998 1895 37014 1959
rect 37078 1895 37220 1959
rect 37284 1895 37300 1959
rect 37364 1895 37380 1959
rect 37444 1895 37460 1959
rect 37524 1895 37540 1959
rect 37604 1895 37620 1959
rect 37684 1895 37826 1959
rect 37890 1895 37906 1959
rect 37970 1895 37986 1959
rect 38050 1895 38066 1959
rect 38130 1895 38146 1959
rect 38210 1895 38226 1959
rect 38290 1895 38432 1959
rect 38496 1895 38512 1959
rect 38576 1895 38592 1959
rect 38656 1895 38672 1959
rect 38736 1895 38752 1959
rect 38816 1895 38832 1959
rect 38896 1895 39038 1959
rect 39102 1895 39118 1959
rect 39182 1895 39198 1959
rect 39262 1895 39278 1959
rect 39342 1895 39358 1959
rect 39422 1895 39438 1959
rect 39502 1895 39606 1959
rect 20148 1893 39606 1895
rect -459 1739 -393 1893
rect -459 1675 -458 1739
rect -394 1675 -393 1739
rect -459 1659 -393 1675
rect -459 1595 -458 1659
rect -394 1595 -393 1659
rect -459 1579 -393 1595
rect -459 1515 -458 1579
rect -394 1515 -393 1579
rect -459 1499 -393 1515
rect -459 1435 -458 1499
rect -394 1435 -393 1499
rect -459 1419 -393 1435
rect -459 1355 -458 1419
rect -394 1355 -393 1419
rect -459 1339 -393 1355
rect -459 1275 -458 1339
rect -394 1275 -393 1339
rect -459 1259 -393 1275
rect -459 1195 -458 1259
rect -394 1195 -393 1259
rect -459 1179 -393 1195
rect -459 1115 -458 1179
rect -394 1115 -393 1179
rect -459 1099 -393 1115
rect -459 1035 -458 1099
rect -394 1035 -393 1099
rect -459 1019 -393 1035
rect -459 955 -458 1019
rect -394 955 -393 1019
rect -459 865 -393 955
rect -333 801 -273 1831
rect -213 861 -153 1893
rect -93 801 -33 1831
rect 27 861 87 1893
rect 147 1739 213 1893
rect 147 1675 148 1739
rect 212 1675 213 1739
rect 147 1659 213 1675
rect 147 1595 148 1659
rect 212 1595 213 1659
rect 147 1579 213 1595
rect 147 1515 148 1579
rect 212 1515 213 1579
rect 147 1499 213 1515
rect 147 1435 148 1499
rect 212 1435 213 1499
rect 147 1419 213 1435
rect 147 1355 148 1419
rect 212 1355 213 1419
rect 147 1339 213 1355
rect 147 1275 148 1339
rect 212 1275 213 1339
rect 147 1259 213 1275
rect 147 1195 148 1259
rect 212 1195 213 1259
rect 147 1179 213 1195
rect 147 1115 148 1179
rect 212 1115 213 1179
rect 147 1099 213 1115
rect 147 1035 148 1099
rect 212 1035 213 1099
rect 147 1019 213 1035
rect 147 955 148 1019
rect 212 955 213 1019
rect 147 865 213 955
rect 355 1739 421 1829
rect 355 1675 356 1739
rect 420 1675 421 1739
rect 355 1659 421 1675
rect 355 1595 356 1659
rect 420 1595 421 1659
rect 355 1579 421 1595
rect 355 1515 356 1579
rect 420 1515 421 1579
rect 355 1499 421 1515
rect 355 1435 356 1499
rect 420 1435 421 1499
rect 355 1419 421 1435
rect 355 1355 356 1419
rect 420 1355 421 1419
rect 355 1339 421 1355
rect 355 1275 356 1339
rect 420 1275 421 1339
rect 355 1259 421 1275
rect 355 1195 356 1259
rect 420 1195 421 1259
rect 355 1179 421 1195
rect 355 1115 356 1179
rect 420 1115 421 1179
rect 355 1099 421 1115
rect 355 1035 356 1099
rect 420 1035 421 1099
rect 355 1019 421 1035
rect 355 955 356 1019
rect 420 955 421 1019
rect 355 801 421 955
rect 481 801 541 1833
rect 601 863 661 1893
rect 721 801 781 1833
rect 841 863 901 1893
rect 964 1829 1024 1832
rect 961 1821 1027 1829
rect 961 1757 962 1821
rect 1026 1757 1027 1821
rect 961 1739 1027 1757
rect 961 1675 962 1739
rect 1026 1675 1027 1739
rect 961 1671 1027 1675
rect 961 1659 966 1671
rect 1022 1659 1027 1671
rect 961 1595 962 1659
rect 1026 1595 1027 1659
rect 961 1579 1027 1595
rect 961 1515 962 1579
rect 1026 1515 1027 1579
rect 961 1499 1027 1515
rect 961 1435 962 1499
rect 1026 1435 1027 1499
rect 961 1419 1027 1435
rect 961 1355 962 1419
rect 1026 1355 1027 1419
rect 961 1339 1027 1355
rect 961 1275 962 1339
rect 1026 1275 1027 1339
rect 961 1259 1027 1275
rect 961 1195 962 1259
rect 1026 1195 1027 1259
rect 961 1179 1027 1195
rect 961 1115 962 1179
rect 1026 1115 1027 1179
rect 961 1099 1027 1115
rect 961 1035 962 1099
rect 1026 1035 1027 1099
rect 961 1019 1027 1035
rect 961 955 962 1019
rect 1026 955 1027 1019
rect 961 801 1027 955
rect -459 799 213 801
rect -459 735 -355 799
rect -291 735 -275 799
rect -211 735 -195 799
rect -131 735 -115 799
rect -51 735 -35 799
rect 29 735 45 799
rect 109 735 213 799
rect -459 733 213 735
rect 355 799 1027 801
rect 355 735 459 799
rect 523 735 539 799
rect 603 735 619 799
rect 683 735 699 799
rect 763 735 779 799
rect 843 735 859 799
rect 923 735 1027 799
rect 355 733 1027 735
rect -459 579 -393 669
rect -459 515 -458 579
rect -394 515 -393 579
rect -459 499 -393 515
rect -459 435 -458 499
rect -394 435 -393 499
rect -459 419 -393 435
rect -459 355 -458 419
rect -394 355 -393 419
rect -459 339 -393 355
rect -459 275 -458 339
rect -394 275 -393 339
rect -459 259 -393 275
rect -459 195 -458 259
rect -394 195 -393 259
rect -459 179 -393 195
rect -459 115 -458 179
rect -394 115 -393 179
rect -459 99 -393 115
rect -459 35 -458 99
rect -394 35 -393 99
rect -459 19 -393 35
rect -459 -45 -458 19
rect -394 -45 -393 19
rect -459 -61 -393 -45
rect -459 -125 -458 -61
rect -394 -125 -393 -61
rect -459 -141 -393 -125
rect -459 -205 -458 -141
rect -394 -205 -393 -141
rect -459 -359 -393 -205
rect -333 -359 -273 673
rect -213 -297 -153 733
rect -93 -359 -33 673
rect 27 -297 87 733
rect 147 579 213 669
rect 147 515 148 579
rect 212 515 213 579
rect 147 499 213 515
rect 147 435 148 499
rect 212 435 213 499
rect 147 419 213 435
rect 147 355 148 419
rect 212 355 213 419
rect 147 339 213 355
rect 147 275 148 339
rect 212 275 213 339
rect 147 259 213 275
rect 147 195 148 259
rect 212 195 213 259
rect 147 179 213 195
rect 147 115 148 179
rect 212 115 213 179
rect 147 99 213 115
rect 147 35 148 99
rect 212 35 213 99
rect 147 19 213 35
rect 147 -45 148 19
rect 212 -45 213 19
rect 147 -61 213 -45
rect 147 -125 148 -61
rect 212 -125 213 -61
rect 147 -141 213 -125
rect 147 -205 148 -141
rect 212 -205 213 -141
rect 147 -359 213 -205
rect 355 579 421 733
rect 355 515 356 579
rect 420 515 421 579
rect 355 499 421 515
rect 355 435 356 499
rect 420 435 421 499
rect 355 419 421 435
rect 355 355 356 419
rect 420 355 421 419
rect 355 339 421 355
rect 355 275 356 339
rect 420 275 421 339
rect 355 259 421 275
rect 355 195 356 259
rect 420 195 421 259
rect 355 179 421 195
rect 355 115 356 179
rect 420 115 421 179
rect 355 99 421 115
rect 355 35 356 99
rect 420 35 421 99
rect 355 19 421 35
rect 355 -45 356 19
rect 420 -45 421 19
rect 355 -61 421 -45
rect 355 -125 356 -61
rect 420 -125 421 -61
rect 355 -141 421 -125
rect 355 -205 356 -141
rect 420 -205 421 -141
rect 355 -295 421 -205
rect 481 -359 541 671
rect 601 -299 661 733
rect 721 -359 781 671
rect 841 -299 901 733
rect 961 579 1027 733
rect 961 515 962 579
rect 1026 515 1027 579
rect 961 499 1027 515
rect 961 435 962 499
rect 1026 435 1027 499
rect 961 419 1027 435
rect 961 355 962 419
rect 1026 355 1027 419
rect 961 339 1027 355
rect 961 275 962 339
rect 1026 275 1027 339
rect 961 259 1027 275
rect 961 195 962 259
rect 1026 195 1027 259
rect 961 179 1027 195
rect 961 115 962 179
rect 1026 115 1027 179
rect 961 99 1027 115
rect 961 35 962 99
rect 1026 35 1027 99
rect 961 19 1027 35
rect 961 -45 962 19
rect 1026 -45 1027 19
rect 961 -61 1027 -45
rect 961 -125 962 -61
rect 1026 -125 1027 -61
rect 961 -141 1027 -125
rect 961 -205 962 -141
rect 1026 -205 1027 -141
rect 961 -295 1027 -205
rect 1267 1739 1333 1829
rect 1267 1675 1268 1739
rect 1332 1675 1333 1739
rect 1267 1659 1333 1675
rect 1267 1595 1268 1659
rect 1332 1595 1333 1659
rect 1267 1579 1333 1595
rect 1267 1515 1268 1579
rect 1332 1515 1333 1579
rect 1267 1499 1333 1515
rect 1267 1435 1268 1499
rect 1332 1435 1333 1499
rect 1267 1419 1333 1435
rect 1267 1355 1268 1419
rect 1332 1355 1333 1419
rect 1267 1339 1333 1355
rect 1267 1275 1268 1339
rect 1332 1275 1333 1339
rect 1267 1259 1333 1275
rect 1267 1195 1268 1259
rect 1332 1195 1333 1259
rect 1267 1179 1333 1195
rect 1267 1115 1268 1179
rect 1332 1115 1333 1179
rect 1267 1099 1333 1115
rect 1267 1035 1268 1099
rect 1332 1035 1333 1099
rect 1267 1019 1333 1035
rect 1267 955 1268 1019
rect 1332 955 1333 1019
rect 1267 801 1333 955
rect 1393 801 1453 1833
rect 1513 863 1573 1893
rect 1633 801 1693 1833
rect 1753 863 1813 1893
rect 1873 1820 1939 1829
rect 1873 1756 1874 1820
rect 1938 1756 1939 1820
rect 1873 1739 1939 1756
rect 1873 1675 1874 1739
rect 1938 1675 1939 1739
rect 1873 1659 1939 1675
rect 1873 1595 1874 1659
rect 1938 1595 1939 1659
rect 1873 1579 1939 1595
rect 1873 1515 1874 1579
rect 1938 1515 1939 1579
rect 1873 1499 1939 1515
rect 1873 1435 1874 1499
rect 1938 1435 1939 1499
rect 1873 1419 1939 1435
rect 1873 1355 1874 1419
rect 1938 1355 1939 1419
rect 1873 1339 1939 1355
rect 1873 1275 1874 1339
rect 1938 1275 1939 1339
rect 1873 1259 1939 1275
rect 1873 1195 1874 1259
rect 1938 1195 1939 1259
rect 1873 1179 1939 1195
rect 1873 1115 1874 1179
rect 1938 1115 1939 1179
rect 1873 1099 1939 1115
rect 1873 1035 1874 1099
rect 1938 1035 1939 1099
rect 1873 1019 1939 1035
rect 1873 955 1874 1019
rect 1938 955 1939 1019
rect 1873 801 1939 955
rect 1999 801 2059 1833
rect 2119 863 2179 1893
rect 2239 801 2299 1833
rect 2359 863 2419 1893
rect 2482 1830 2542 1832
rect 2479 1821 2545 1830
rect 2479 1757 2480 1821
rect 2544 1757 2545 1821
rect 2479 1739 2545 1757
rect 2479 1675 2480 1739
rect 2544 1675 2545 1739
rect 2479 1659 2545 1675
rect 2479 1595 2480 1659
rect 2544 1595 2545 1659
rect 2479 1579 2545 1595
rect 2479 1515 2480 1579
rect 2544 1515 2545 1579
rect 2479 1499 2545 1515
rect 2479 1435 2480 1499
rect 2544 1435 2545 1499
rect 2479 1419 2545 1435
rect 2479 1355 2480 1419
rect 2544 1355 2545 1419
rect 2479 1339 2545 1355
rect 2479 1275 2480 1339
rect 2544 1275 2545 1339
rect 2479 1259 2545 1275
rect 2479 1195 2480 1259
rect 2544 1195 2545 1259
rect 2479 1179 2545 1195
rect 2479 1115 2480 1179
rect 2544 1115 2545 1179
rect 2479 1099 2545 1115
rect 2479 1035 2480 1099
rect 2544 1035 2545 1099
rect 2479 1019 2545 1035
rect 2479 955 2480 1019
rect 2544 955 2545 1019
rect 2479 801 2545 955
rect 1267 799 2545 801
rect 1267 735 1371 799
rect 1435 735 1451 799
rect 1515 735 1531 799
rect 1595 735 1611 799
rect 1675 735 1691 799
rect 1755 735 1771 799
rect 1835 735 1977 799
rect 2041 735 2057 799
rect 2121 735 2137 799
rect 2201 735 2217 799
rect 2281 735 2297 799
rect 2361 735 2377 799
rect 2441 735 2545 799
rect 1267 733 2545 735
rect 1267 579 1333 733
rect 1267 515 1268 579
rect 1332 515 1333 579
rect 1267 499 1333 515
rect 1267 435 1268 499
rect 1332 435 1333 499
rect 1267 419 1333 435
rect 1267 355 1268 419
rect 1332 355 1333 419
rect 1267 339 1333 355
rect 1267 275 1268 339
rect 1332 275 1333 339
rect 1267 259 1333 275
rect 1267 195 1268 259
rect 1332 195 1333 259
rect 1267 179 1333 195
rect 1267 115 1268 179
rect 1332 115 1333 179
rect 1267 99 1333 115
rect 1267 35 1268 99
rect 1332 35 1333 99
rect 1267 19 1333 35
rect 1267 -45 1268 19
rect 1332 -45 1333 19
rect 1267 -61 1333 -45
rect 1267 -125 1268 -61
rect 1332 -125 1333 -61
rect 1267 -141 1333 -125
rect 1267 -205 1268 -141
rect 1332 -205 1333 -141
rect 1267 -295 1333 -205
rect 1393 -359 1453 671
rect 1513 -299 1573 733
rect 1633 -359 1693 671
rect 1753 -299 1813 733
rect 1873 579 1939 733
rect 1873 515 1874 579
rect 1938 515 1939 579
rect 1873 499 1939 515
rect 1873 435 1874 499
rect 1938 435 1939 499
rect 1873 419 1939 435
rect 1873 355 1874 419
rect 1938 355 1939 419
rect 1873 339 1939 355
rect 1873 275 1874 339
rect 1938 275 1939 339
rect 1873 259 1939 275
rect 1873 195 1874 259
rect 1938 195 1939 259
rect 1873 179 1939 195
rect 1873 115 1874 179
rect 1938 115 1939 179
rect 1873 99 1939 115
rect 1873 35 1874 99
rect 1938 35 1939 99
rect 1873 19 1939 35
rect 1873 -45 1874 19
rect 1938 -45 1939 19
rect 1873 -61 1939 -45
rect 1873 -125 1874 -61
rect 1938 -125 1939 -61
rect 1873 -141 1939 -125
rect 1873 -205 1874 -141
rect 1938 -205 1939 -141
rect 1873 -295 1939 -205
rect 1999 -359 2059 671
rect 2119 -299 2179 733
rect 2239 -359 2299 671
rect 2359 -299 2419 733
rect 2479 579 2545 733
rect 2479 515 2480 579
rect 2544 515 2545 579
rect 2479 499 2545 515
rect 2479 435 2480 499
rect 2544 435 2545 499
rect 2479 419 2545 435
rect 2479 355 2480 419
rect 2544 355 2545 419
rect 2479 339 2545 355
rect 2479 275 2480 339
rect 2544 275 2545 339
rect 2479 259 2545 275
rect 2479 195 2480 259
rect 2544 195 2545 259
rect 2479 179 2545 195
rect 2479 115 2480 179
rect 2544 115 2545 179
rect 2479 99 2545 115
rect 2479 35 2480 99
rect 2544 35 2545 99
rect 2479 19 2545 35
rect 2479 -45 2480 19
rect 2544 -45 2545 19
rect 2479 -61 2545 -45
rect 2479 -125 2480 -61
rect 2544 -125 2545 -61
rect 2479 -141 2545 -125
rect 2479 -205 2480 -141
rect 2544 -205 2545 -141
rect 2479 -295 2545 -205
rect 2801 1739 2867 1829
rect 2801 1675 2802 1739
rect 2866 1675 2867 1739
rect 2801 1659 2867 1675
rect 2801 1595 2802 1659
rect 2866 1595 2867 1659
rect 2801 1579 2867 1595
rect 2801 1515 2802 1579
rect 2866 1515 2867 1579
rect 2801 1499 2867 1515
rect 2801 1435 2802 1499
rect 2866 1435 2867 1499
rect 2801 1419 2867 1435
rect 2801 1355 2802 1419
rect 2866 1355 2867 1419
rect 2801 1339 2867 1355
rect 2801 1275 2802 1339
rect 2866 1275 2867 1339
rect 2801 1259 2867 1275
rect 2801 1195 2802 1259
rect 2866 1195 2867 1259
rect 2801 1179 2867 1195
rect 2801 1115 2802 1179
rect 2866 1115 2867 1179
rect 2801 1099 2867 1115
rect 2801 1035 2802 1099
rect 2866 1035 2867 1099
rect 2801 1019 2867 1035
rect 2801 955 2802 1019
rect 2866 955 2867 1019
rect 2801 801 2867 955
rect 2927 801 2987 1833
rect 3047 863 3107 1893
rect 3167 801 3227 1833
rect 3287 863 3347 1893
rect 3407 1806 3473 1829
rect 3407 1750 3412 1806
rect 3468 1750 3473 1806
rect 3407 1739 3473 1750
rect 3407 1675 3408 1739
rect 3472 1675 3473 1739
rect 3407 1659 3473 1675
rect 3407 1595 3408 1659
rect 3472 1595 3473 1659
rect 3407 1579 3473 1595
rect 3407 1515 3408 1579
rect 3472 1515 3473 1579
rect 3407 1499 3473 1515
rect 3407 1435 3408 1499
rect 3472 1435 3473 1499
rect 3407 1419 3473 1435
rect 3407 1355 3408 1419
rect 3472 1355 3473 1419
rect 3407 1339 3473 1355
rect 3407 1275 3408 1339
rect 3472 1275 3473 1339
rect 3407 1259 3473 1275
rect 3407 1195 3408 1259
rect 3472 1195 3473 1259
rect 3407 1179 3473 1195
rect 3407 1115 3408 1179
rect 3472 1115 3473 1179
rect 3407 1099 3473 1115
rect 3407 1035 3408 1099
rect 3472 1035 3473 1099
rect 3407 1019 3473 1035
rect 3407 955 3408 1019
rect 3472 955 3473 1019
rect 3407 801 3473 955
rect 3533 801 3593 1833
rect 3653 863 3713 1893
rect 3773 801 3833 1833
rect 3893 863 3953 1893
rect 4013 1739 4079 1829
rect 4013 1675 4014 1739
rect 4078 1675 4079 1739
rect 4013 1659 4079 1675
rect 4013 1595 4014 1659
rect 4078 1595 4079 1659
rect 4013 1579 4079 1595
rect 4013 1515 4014 1579
rect 4078 1515 4079 1579
rect 4013 1499 4079 1515
rect 4013 1435 4014 1499
rect 4078 1435 4079 1499
rect 4013 1419 4079 1435
rect 4013 1355 4014 1419
rect 4078 1355 4079 1419
rect 4013 1339 4079 1355
rect 4013 1275 4014 1339
rect 4078 1275 4079 1339
rect 4013 1259 4079 1275
rect 4013 1195 4014 1259
rect 4078 1195 4079 1259
rect 4013 1179 4079 1195
rect 4013 1115 4014 1179
rect 4078 1115 4079 1179
rect 4013 1099 4079 1115
rect 4013 1035 4014 1099
rect 4078 1035 4079 1099
rect 4013 1019 4079 1035
rect 4013 955 4014 1019
rect 4078 955 4079 1019
rect 4013 801 4079 955
rect 4139 801 4199 1833
rect 4259 863 4319 1893
rect 4379 801 4439 1833
rect 4499 863 4559 1893
rect 4619 1807 4685 1829
rect 4619 1751 4624 1807
rect 4680 1751 4685 1807
rect 4619 1739 4685 1751
rect 4619 1675 4620 1739
rect 4684 1675 4685 1739
rect 4619 1659 4685 1675
rect 4619 1595 4620 1659
rect 4684 1595 4685 1659
rect 4619 1579 4685 1595
rect 4619 1515 4620 1579
rect 4684 1515 4685 1579
rect 4619 1499 4685 1515
rect 4619 1435 4620 1499
rect 4684 1435 4685 1499
rect 4619 1419 4685 1435
rect 4619 1355 4620 1419
rect 4684 1355 4685 1419
rect 4619 1339 4685 1355
rect 4619 1275 4620 1339
rect 4684 1275 4685 1339
rect 4619 1259 4685 1275
rect 4619 1195 4620 1259
rect 4684 1195 4685 1259
rect 4619 1179 4685 1195
rect 4619 1115 4620 1179
rect 4684 1115 4685 1179
rect 4619 1099 4685 1115
rect 4619 1035 4620 1099
rect 4684 1035 4685 1099
rect 4619 1019 4685 1035
rect 4619 955 4620 1019
rect 4684 955 4685 1019
rect 4619 801 4685 955
rect 4745 801 4805 1833
rect 4865 863 4925 1893
rect 4985 801 5045 1833
rect 5105 863 5165 1893
rect 5225 1807 5291 1829
rect 5225 1751 5230 1807
rect 5286 1751 5291 1807
rect 5225 1739 5291 1751
rect 5225 1675 5226 1739
rect 5290 1675 5291 1739
rect 5225 1659 5291 1675
rect 5225 1595 5226 1659
rect 5290 1595 5291 1659
rect 5225 1579 5291 1595
rect 5225 1515 5226 1579
rect 5290 1515 5291 1579
rect 5225 1499 5291 1515
rect 5225 1435 5226 1499
rect 5290 1435 5291 1499
rect 5225 1419 5291 1435
rect 5225 1355 5226 1419
rect 5290 1355 5291 1419
rect 5225 1339 5291 1355
rect 5225 1275 5226 1339
rect 5290 1275 5291 1339
rect 5225 1259 5291 1275
rect 5225 1195 5226 1259
rect 5290 1195 5291 1259
rect 5225 1179 5291 1195
rect 5225 1115 5226 1179
rect 5290 1115 5291 1179
rect 5225 1099 5291 1115
rect 5225 1035 5226 1099
rect 5290 1035 5291 1099
rect 5225 1019 5291 1035
rect 5225 955 5226 1019
rect 5290 955 5291 1019
rect 5225 801 5291 955
rect 2801 799 5291 801
rect 2801 735 2905 799
rect 2969 735 2985 799
rect 3049 735 3065 799
rect 3129 735 3145 799
rect 3209 735 3225 799
rect 3289 735 3305 799
rect 3369 735 3511 799
rect 3575 735 3591 799
rect 3655 735 3671 799
rect 3735 735 3751 799
rect 3815 735 3831 799
rect 3895 735 3911 799
rect 3975 735 4117 799
rect 4181 735 4197 799
rect 4261 735 4277 799
rect 4341 735 4357 799
rect 4421 735 4437 799
rect 4501 735 4517 799
rect 4581 735 4723 799
rect 4787 735 4803 799
rect 4867 735 4883 799
rect 4947 735 4963 799
rect 5027 735 5043 799
rect 5107 735 5123 799
rect 5187 735 5291 799
rect 2801 733 5291 735
rect 2801 579 2867 733
rect 2801 515 2802 579
rect 2866 515 2867 579
rect 2801 499 2867 515
rect 2801 435 2802 499
rect 2866 435 2867 499
rect 2801 419 2867 435
rect 2801 355 2802 419
rect 2866 355 2867 419
rect 2801 339 2867 355
rect 2801 275 2802 339
rect 2866 275 2867 339
rect 2801 259 2867 275
rect 2801 195 2802 259
rect 2866 195 2867 259
rect 2801 179 2867 195
rect 2801 115 2802 179
rect 2866 115 2867 179
rect 2801 99 2867 115
rect 2801 35 2802 99
rect 2866 35 2867 99
rect 2801 19 2867 35
rect 2801 -45 2802 19
rect 2866 -45 2867 19
rect 2801 -61 2867 -45
rect 2801 -125 2802 -61
rect 2866 -125 2867 -61
rect 2801 -141 2867 -125
rect 2801 -205 2802 -141
rect 2866 -205 2867 -141
rect 2801 -295 2867 -205
rect 2927 -359 2987 671
rect 3047 -299 3107 733
rect 3167 -359 3227 671
rect 3287 -299 3347 733
rect 3407 579 3473 733
rect 3407 515 3408 579
rect 3472 515 3473 579
rect 3407 499 3473 515
rect 3407 435 3408 499
rect 3472 435 3473 499
rect 3407 419 3473 435
rect 3407 355 3408 419
rect 3472 355 3473 419
rect 3407 339 3473 355
rect 3407 275 3408 339
rect 3472 275 3473 339
rect 3407 259 3473 275
rect 3407 195 3408 259
rect 3472 195 3473 259
rect 3407 179 3473 195
rect 3407 115 3408 179
rect 3472 115 3473 179
rect 3407 99 3473 115
rect 3407 35 3408 99
rect 3472 35 3473 99
rect 3407 19 3473 35
rect 3407 -45 3408 19
rect 3472 -45 3473 19
rect 3407 -61 3473 -45
rect 3407 -125 3408 -61
rect 3472 -125 3473 -61
rect 3407 -141 3473 -125
rect 3407 -205 3408 -141
rect 3472 -205 3473 -141
rect 3407 -295 3473 -205
rect 3533 -359 3593 671
rect 3653 -299 3713 733
rect 3773 -359 3833 671
rect 3893 -299 3953 733
rect 4013 579 4079 733
rect 4013 515 4014 579
rect 4078 515 4079 579
rect 4013 499 4079 515
rect 4013 435 4014 499
rect 4078 435 4079 499
rect 4013 419 4079 435
rect 4013 355 4014 419
rect 4078 355 4079 419
rect 4013 339 4079 355
rect 4013 275 4014 339
rect 4078 275 4079 339
rect 4013 259 4079 275
rect 4013 195 4014 259
rect 4078 195 4079 259
rect 4013 179 4079 195
rect 4013 115 4014 179
rect 4078 115 4079 179
rect 4013 99 4079 115
rect 4013 35 4014 99
rect 4078 35 4079 99
rect 4013 19 4079 35
rect 4013 -45 4014 19
rect 4078 -45 4079 19
rect 4013 -61 4079 -45
rect 4013 -125 4014 -61
rect 4078 -125 4079 -61
rect 4013 -141 4079 -125
rect 4013 -205 4014 -141
rect 4078 -205 4079 -141
rect 4013 -295 4079 -205
rect 4139 -359 4199 671
rect 4259 -299 4319 733
rect 4379 -359 4439 671
rect 4499 -299 4559 733
rect 4619 579 4685 733
rect 4619 515 4620 579
rect 4684 515 4685 579
rect 4619 499 4685 515
rect 4619 435 4620 499
rect 4684 435 4685 499
rect 4619 419 4685 435
rect 4619 355 4620 419
rect 4684 355 4685 419
rect 4619 339 4685 355
rect 4619 275 4620 339
rect 4684 275 4685 339
rect 4619 259 4685 275
rect 4619 195 4620 259
rect 4684 195 4685 259
rect 4619 179 4685 195
rect 4619 115 4620 179
rect 4684 115 4685 179
rect 4619 99 4685 115
rect 4619 35 4620 99
rect 4684 35 4685 99
rect 4619 19 4685 35
rect 4619 -45 4620 19
rect 4684 -45 4685 19
rect 4619 -61 4685 -45
rect 4619 -125 4620 -61
rect 4684 -125 4685 -61
rect 4619 -141 4685 -125
rect 4619 -205 4620 -141
rect 4684 -205 4685 -141
rect 4619 -295 4685 -205
rect 4745 -359 4805 671
rect 4865 -299 4925 733
rect 4985 -359 5045 671
rect 5105 -299 5165 733
rect 5225 579 5291 733
rect 5225 515 5226 579
rect 5290 515 5291 579
rect 5225 499 5291 515
rect 5225 435 5226 499
rect 5290 435 5291 499
rect 5225 419 5291 435
rect 5225 355 5226 419
rect 5290 355 5291 419
rect 5225 339 5291 355
rect 5225 275 5226 339
rect 5290 275 5291 339
rect 5225 259 5291 275
rect 5225 195 5226 259
rect 5290 195 5291 259
rect 5225 179 5291 195
rect 5225 115 5226 179
rect 5290 115 5291 179
rect 5225 99 5291 115
rect 5225 35 5226 99
rect 5290 35 5291 99
rect 5225 19 5291 35
rect 5225 -45 5226 19
rect 5290 -45 5291 19
rect 5225 -61 5291 -45
rect 5225 -125 5226 -61
rect 5290 -125 5291 -61
rect 5225 -141 5291 -125
rect 5225 -205 5226 -141
rect 5290 -205 5291 -141
rect 5225 -295 5291 -205
rect 5352 1739 5418 1829
rect 5352 1675 5353 1739
rect 5417 1675 5418 1739
rect 5352 1659 5418 1675
rect 5352 1595 5353 1659
rect 5417 1595 5418 1659
rect 5352 1579 5418 1595
rect 5352 1515 5353 1579
rect 5417 1515 5418 1579
rect 5352 1499 5418 1515
rect 5352 1435 5353 1499
rect 5417 1435 5418 1499
rect 5352 1419 5418 1435
rect 5352 1355 5353 1419
rect 5417 1355 5418 1419
rect 5352 1339 5418 1355
rect 5352 1275 5353 1339
rect 5417 1275 5418 1339
rect 5352 1259 5418 1275
rect 5352 1195 5353 1259
rect 5417 1195 5418 1259
rect 5352 1179 5418 1195
rect 5352 1115 5353 1179
rect 5417 1115 5418 1179
rect 5352 1099 5418 1115
rect 5352 1035 5353 1099
rect 5417 1035 5418 1099
rect 5352 1019 5418 1035
rect 5352 955 5353 1019
rect 5417 955 5418 1019
rect 5352 801 5418 955
rect 5478 801 5538 1833
rect 5598 863 5658 1893
rect 5718 801 5778 1833
rect 5838 863 5898 1893
rect 5958 1739 6024 1829
rect 5958 1675 5959 1739
rect 6023 1675 6024 1739
rect 5958 1659 6024 1675
rect 5958 1595 5959 1659
rect 6023 1595 6024 1659
rect 5958 1579 6024 1595
rect 5958 1515 5959 1579
rect 6023 1515 6024 1579
rect 5958 1499 6024 1515
rect 5958 1435 5959 1499
rect 6023 1435 6024 1499
rect 5958 1419 6024 1435
rect 5958 1355 5959 1419
rect 6023 1355 6024 1419
rect 5958 1339 6024 1355
rect 5958 1275 5959 1339
rect 6023 1275 6024 1339
rect 5958 1259 6024 1275
rect 5958 1195 5959 1259
rect 6023 1195 6024 1259
rect 5958 1179 6024 1195
rect 5958 1115 5959 1179
rect 6023 1115 6024 1179
rect 5958 1099 6024 1115
rect 5958 1035 5959 1099
rect 6023 1035 6024 1099
rect 5958 1019 6024 1035
rect 5958 955 5959 1019
rect 6023 955 6024 1019
rect 5958 801 6024 955
rect 6084 801 6144 1833
rect 6204 863 6264 1893
rect 6324 801 6384 1833
rect 6444 863 6504 1893
rect 6564 1739 6630 1829
rect 6564 1675 6565 1739
rect 6629 1675 6630 1739
rect 6564 1659 6630 1675
rect 6564 1595 6565 1659
rect 6629 1595 6630 1659
rect 6564 1579 6630 1595
rect 6564 1515 6565 1579
rect 6629 1515 6630 1579
rect 6564 1499 6630 1515
rect 6564 1435 6565 1499
rect 6629 1435 6630 1499
rect 6564 1419 6630 1435
rect 6564 1355 6565 1419
rect 6629 1355 6630 1419
rect 6564 1339 6630 1355
rect 6564 1275 6565 1339
rect 6629 1275 6630 1339
rect 6564 1259 6630 1275
rect 6564 1195 6565 1259
rect 6629 1195 6630 1259
rect 6564 1179 6630 1195
rect 6564 1115 6565 1179
rect 6629 1115 6630 1179
rect 6564 1099 6630 1115
rect 6564 1035 6565 1099
rect 6629 1035 6630 1099
rect 6564 1019 6630 1035
rect 6564 955 6565 1019
rect 6629 955 6630 1019
rect 6564 801 6630 955
rect 6690 801 6750 1833
rect 6810 863 6870 1893
rect 6930 801 6990 1833
rect 7050 863 7110 1893
rect 7170 1739 7236 1829
rect 7170 1675 7171 1739
rect 7235 1675 7236 1739
rect 7170 1659 7236 1675
rect 7170 1595 7171 1659
rect 7235 1595 7236 1659
rect 7170 1579 7236 1595
rect 7170 1515 7171 1579
rect 7235 1515 7236 1579
rect 7170 1499 7236 1515
rect 7170 1435 7171 1499
rect 7235 1435 7236 1499
rect 7170 1419 7236 1435
rect 7170 1355 7171 1419
rect 7235 1355 7236 1419
rect 7170 1339 7236 1355
rect 7170 1275 7171 1339
rect 7235 1275 7236 1339
rect 7170 1259 7236 1275
rect 7170 1195 7171 1259
rect 7235 1195 7236 1259
rect 7170 1179 7236 1195
rect 7170 1115 7171 1179
rect 7235 1115 7236 1179
rect 7170 1099 7236 1115
rect 7170 1035 7171 1099
rect 7235 1035 7236 1099
rect 7170 1019 7236 1035
rect 7170 955 7171 1019
rect 7235 955 7236 1019
rect 7170 801 7236 955
rect 7296 801 7356 1833
rect 7416 863 7476 1893
rect 7536 801 7596 1833
rect 7656 863 7716 1893
rect 7776 1820 7842 1829
rect 7776 1764 7781 1820
rect 7837 1764 7842 1820
rect 7776 1739 7842 1764
rect 7776 1675 7777 1739
rect 7841 1675 7842 1739
rect 7776 1659 7842 1675
rect 7776 1595 7777 1659
rect 7841 1595 7842 1659
rect 7776 1579 7842 1595
rect 7776 1515 7777 1579
rect 7841 1515 7842 1579
rect 7776 1499 7842 1515
rect 7776 1435 7777 1499
rect 7841 1435 7842 1499
rect 7776 1419 7842 1435
rect 7776 1355 7777 1419
rect 7841 1355 7842 1419
rect 7776 1339 7842 1355
rect 7776 1275 7777 1339
rect 7841 1275 7842 1339
rect 7776 1259 7842 1275
rect 7776 1195 7777 1259
rect 7841 1195 7842 1259
rect 7776 1179 7842 1195
rect 7776 1115 7777 1179
rect 7841 1115 7842 1179
rect 7776 1099 7842 1115
rect 7776 1035 7777 1099
rect 7841 1035 7842 1099
rect 7776 1019 7842 1035
rect 7776 955 7777 1019
rect 7841 955 7842 1019
rect 7776 801 7842 955
rect 7902 801 7962 1833
rect 8022 863 8082 1893
rect 8142 801 8202 1833
rect 8262 863 8322 1893
rect 8382 1820 8448 1829
rect 8382 1764 8387 1820
rect 8443 1764 8448 1820
rect 8382 1739 8448 1764
rect 8382 1675 8383 1739
rect 8447 1675 8448 1739
rect 8382 1659 8448 1675
rect 8382 1595 8383 1659
rect 8447 1595 8448 1659
rect 8382 1579 8448 1595
rect 8382 1515 8383 1579
rect 8447 1515 8448 1579
rect 8382 1499 8448 1515
rect 8382 1435 8383 1499
rect 8447 1435 8448 1499
rect 8382 1419 8448 1435
rect 8382 1355 8383 1419
rect 8447 1355 8448 1419
rect 8382 1339 8448 1355
rect 8382 1275 8383 1339
rect 8447 1275 8448 1339
rect 8382 1259 8448 1275
rect 8382 1195 8383 1259
rect 8447 1195 8448 1259
rect 8382 1179 8448 1195
rect 8382 1115 8383 1179
rect 8447 1115 8448 1179
rect 8382 1099 8448 1115
rect 8382 1035 8383 1099
rect 8447 1035 8448 1099
rect 8382 1019 8448 1035
rect 8382 955 8383 1019
rect 8447 955 8448 1019
rect 8382 801 8448 955
rect 8508 801 8568 1833
rect 8628 863 8688 1893
rect 8748 801 8808 1833
rect 8868 863 8928 1893
rect 8988 1820 9054 1829
rect 8988 1764 8993 1820
rect 9049 1764 9054 1820
rect 8988 1739 9054 1764
rect 8988 1675 8989 1739
rect 9053 1675 9054 1739
rect 8988 1659 9054 1675
rect 8988 1595 8989 1659
rect 9053 1595 9054 1659
rect 8988 1579 9054 1595
rect 8988 1515 8989 1579
rect 9053 1515 9054 1579
rect 8988 1499 9054 1515
rect 8988 1435 8989 1499
rect 9053 1435 9054 1499
rect 8988 1419 9054 1435
rect 8988 1355 8989 1419
rect 9053 1355 9054 1419
rect 8988 1339 9054 1355
rect 8988 1275 8989 1339
rect 9053 1275 9054 1339
rect 8988 1259 9054 1275
rect 8988 1195 8989 1259
rect 9053 1195 9054 1259
rect 8988 1179 9054 1195
rect 8988 1115 8989 1179
rect 9053 1115 9054 1179
rect 8988 1099 9054 1115
rect 8988 1035 8989 1099
rect 9053 1035 9054 1099
rect 8988 1019 9054 1035
rect 8988 955 8989 1019
rect 9053 955 9054 1019
rect 8988 801 9054 955
rect 9114 801 9174 1833
rect 9234 863 9294 1893
rect 9354 801 9414 1833
rect 9474 863 9534 1893
rect 9594 1820 9660 1829
rect 9594 1764 9599 1820
rect 9655 1764 9660 1820
rect 9594 1739 9660 1764
rect 9594 1675 9595 1739
rect 9659 1675 9660 1739
rect 9594 1659 9660 1675
rect 9594 1595 9595 1659
rect 9659 1595 9660 1659
rect 9594 1579 9660 1595
rect 9594 1515 9595 1579
rect 9659 1515 9660 1579
rect 9594 1499 9660 1515
rect 9594 1435 9595 1499
rect 9659 1435 9660 1499
rect 9594 1419 9660 1435
rect 9594 1355 9595 1419
rect 9659 1355 9660 1419
rect 9594 1339 9660 1355
rect 9594 1275 9595 1339
rect 9659 1275 9660 1339
rect 9594 1259 9660 1275
rect 9594 1195 9595 1259
rect 9659 1195 9660 1259
rect 9594 1179 9660 1195
rect 9594 1115 9595 1179
rect 9659 1115 9660 1179
rect 9594 1099 9660 1115
rect 9594 1035 9595 1099
rect 9659 1035 9660 1099
rect 9594 1019 9660 1035
rect 9594 955 9595 1019
rect 9659 955 9660 1019
rect 9594 801 9660 955
rect 9720 801 9780 1833
rect 9840 863 9900 1893
rect 9960 801 10020 1833
rect 10080 863 10140 1893
rect 10200 1809 10266 1829
rect 10200 1753 10205 1809
rect 10261 1753 10266 1809
rect 10200 1739 10266 1753
rect 10200 1675 10201 1739
rect 10265 1675 10266 1739
rect 10200 1659 10266 1675
rect 10200 1595 10201 1659
rect 10265 1595 10266 1659
rect 10200 1579 10266 1595
rect 10200 1515 10201 1579
rect 10265 1515 10266 1579
rect 10200 1499 10266 1515
rect 10200 1435 10201 1499
rect 10265 1435 10266 1499
rect 10200 1419 10266 1435
rect 10200 1355 10201 1419
rect 10265 1355 10266 1419
rect 10200 1339 10266 1355
rect 10200 1275 10201 1339
rect 10265 1275 10266 1339
rect 10200 1259 10266 1275
rect 10200 1195 10201 1259
rect 10265 1195 10266 1259
rect 10200 1179 10266 1195
rect 10200 1115 10201 1179
rect 10265 1115 10266 1179
rect 10200 1099 10266 1115
rect 10200 1035 10201 1099
rect 10265 1035 10266 1099
rect 10200 1019 10266 1035
rect 10200 955 10201 1019
rect 10265 955 10266 1019
rect 10200 801 10266 955
rect 5352 799 10266 801
rect 5352 735 5456 799
rect 5520 735 5536 799
rect 5600 735 5616 799
rect 5680 735 5696 799
rect 5760 735 5776 799
rect 5840 735 5856 799
rect 5920 735 6062 799
rect 6126 735 6142 799
rect 6206 735 6222 799
rect 6286 735 6302 799
rect 6366 735 6382 799
rect 6446 735 6462 799
rect 6526 735 6668 799
rect 6732 735 6748 799
rect 6812 735 6828 799
rect 6892 735 6908 799
rect 6972 735 6988 799
rect 7052 735 7068 799
rect 7132 735 7274 799
rect 7338 735 7354 799
rect 7418 735 7434 799
rect 7498 735 7514 799
rect 7578 735 7594 799
rect 7658 735 7674 799
rect 7738 735 7880 799
rect 7944 735 7960 799
rect 8024 735 8040 799
rect 8104 735 8120 799
rect 8184 735 8200 799
rect 8264 735 8280 799
rect 8344 735 8486 799
rect 8550 735 8566 799
rect 8630 735 8646 799
rect 8710 735 8726 799
rect 8790 735 8806 799
rect 8870 735 8886 799
rect 8950 735 9092 799
rect 9156 735 9172 799
rect 9236 735 9252 799
rect 9316 735 9332 799
rect 9396 735 9412 799
rect 9476 735 9492 799
rect 9556 735 9698 799
rect 9762 735 9778 799
rect 9842 735 9858 799
rect 9922 735 9938 799
rect 10002 735 10018 799
rect 10082 735 10098 799
rect 10162 735 10266 799
rect 5352 733 10266 735
rect 5352 579 5418 733
rect 5352 515 5353 579
rect 5417 515 5418 579
rect 5352 499 5418 515
rect 5352 435 5353 499
rect 5417 435 5418 499
rect 5352 419 5418 435
rect 5352 355 5353 419
rect 5417 355 5418 419
rect 5352 339 5418 355
rect 5352 275 5353 339
rect 5417 275 5418 339
rect 5352 259 5418 275
rect 5352 195 5353 259
rect 5417 195 5418 259
rect 5352 179 5418 195
rect 5352 115 5353 179
rect 5417 115 5418 179
rect 5352 99 5418 115
rect 5352 35 5353 99
rect 5417 35 5418 99
rect 5352 19 5418 35
rect 5352 -45 5353 19
rect 5417 -45 5418 19
rect 5352 -61 5418 -45
rect 5352 -125 5353 -61
rect 5417 -125 5418 -61
rect 5352 -141 5418 -125
rect 5352 -205 5353 -141
rect 5417 -205 5418 -141
rect 5352 -295 5418 -205
rect 5478 -359 5538 671
rect 5598 -299 5658 733
rect 5718 -359 5778 671
rect 5838 -299 5898 733
rect 5958 579 6024 733
rect 5958 515 5959 579
rect 6023 515 6024 579
rect 5958 499 6024 515
rect 5958 435 5959 499
rect 6023 435 6024 499
rect 5958 419 6024 435
rect 5958 355 5959 419
rect 6023 355 6024 419
rect 5958 339 6024 355
rect 5958 275 5959 339
rect 6023 275 6024 339
rect 5958 259 6024 275
rect 5958 195 5959 259
rect 6023 195 6024 259
rect 5958 179 6024 195
rect 5958 115 5959 179
rect 6023 115 6024 179
rect 5958 99 6024 115
rect 5958 35 5959 99
rect 6023 35 6024 99
rect 5958 19 6024 35
rect 5958 -45 5959 19
rect 6023 -45 6024 19
rect 5958 -61 6024 -45
rect 5958 -125 5959 -61
rect 6023 -125 6024 -61
rect 5958 -141 6024 -125
rect 5958 -205 5959 -141
rect 6023 -205 6024 -141
rect 5958 -295 6024 -205
rect 6084 -359 6144 671
rect 6204 -299 6264 733
rect 6324 -359 6384 671
rect 6444 -299 6504 733
rect 6564 579 6630 733
rect 6564 515 6565 579
rect 6629 515 6630 579
rect 6564 499 6630 515
rect 6564 435 6565 499
rect 6629 435 6630 499
rect 6564 419 6630 435
rect 6564 355 6565 419
rect 6629 355 6630 419
rect 6564 339 6630 355
rect 6564 275 6565 339
rect 6629 275 6630 339
rect 6564 259 6630 275
rect 6564 195 6565 259
rect 6629 195 6630 259
rect 6564 179 6630 195
rect 6564 115 6565 179
rect 6629 115 6630 179
rect 6564 99 6630 115
rect 6564 35 6565 99
rect 6629 35 6630 99
rect 6564 19 6630 35
rect 6564 -45 6565 19
rect 6629 -45 6630 19
rect 6564 -61 6630 -45
rect 6564 -125 6565 -61
rect 6629 -125 6630 -61
rect 6564 -141 6630 -125
rect 6564 -205 6565 -141
rect 6629 -205 6630 -141
rect 6564 -295 6630 -205
rect 6690 -359 6750 671
rect 6810 -299 6870 733
rect 6930 -359 6990 671
rect 7050 -299 7110 733
rect 7170 579 7236 733
rect 7170 515 7171 579
rect 7235 515 7236 579
rect 7170 499 7236 515
rect 7170 435 7171 499
rect 7235 435 7236 499
rect 7170 419 7236 435
rect 7170 355 7171 419
rect 7235 355 7236 419
rect 7170 339 7236 355
rect 7170 275 7171 339
rect 7235 275 7236 339
rect 7170 259 7236 275
rect 7170 195 7171 259
rect 7235 195 7236 259
rect 7170 179 7236 195
rect 7170 115 7171 179
rect 7235 115 7236 179
rect 7170 99 7236 115
rect 7170 35 7171 99
rect 7235 35 7236 99
rect 7170 19 7236 35
rect 7170 -45 7171 19
rect 7235 -45 7236 19
rect 7170 -61 7236 -45
rect 7170 -125 7171 -61
rect 7235 -125 7236 -61
rect 7170 -141 7236 -125
rect 7170 -205 7171 -141
rect 7235 -205 7236 -141
rect 7170 -295 7236 -205
rect 7296 -359 7356 671
rect 7416 -299 7476 733
rect 7536 -359 7596 671
rect 7656 -299 7716 733
rect 7776 579 7842 733
rect 7776 515 7777 579
rect 7841 515 7842 579
rect 7776 499 7842 515
rect 7776 435 7777 499
rect 7841 435 7842 499
rect 7776 419 7842 435
rect 7776 355 7777 419
rect 7841 355 7842 419
rect 7776 339 7842 355
rect 7776 275 7777 339
rect 7841 275 7842 339
rect 7776 259 7842 275
rect 7776 195 7777 259
rect 7841 195 7842 259
rect 7776 179 7842 195
rect 7776 115 7777 179
rect 7841 115 7842 179
rect 7776 99 7842 115
rect 7776 35 7777 99
rect 7841 35 7842 99
rect 7776 19 7842 35
rect 7776 -45 7777 19
rect 7841 -45 7842 19
rect 7776 -61 7842 -45
rect 7776 -125 7777 -61
rect 7841 -125 7842 -61
rect 7776 -141 7842 -125
rect 7776 -205 7777 -141
rect 7841 -205 7842 -141
rect 7776 -295 7842 -205
rect 7902 -359 7962 671
rect 8022 -299 8082 733
rect 8142 -359 8202 671
rect 8262 -299 8322 733
rect 8382 579 8448 733
rect 8382 515 8383 579
rect 8447 515 8448 579
rect 8382 499 8448 515
rect 8382 435 8383 499
rect 8447 435 8448 499
rect 8382 419 8448 435
rect 8382 355 8383 419
rect 8447 355 8448 419
rect 8382 339 8448 355
rect 8382 275 8383 339
rect 8447 275 8448 339
rect 8382 259 8448 275
rect 8382 195 8383 259
rect 8447 195 8448 259
rect 8382 179 8448 195
rect 8382 115 8383 179
rect 8447 115 8448 179
rect 8382 99 8448 115
rect 8382 35 8383 99
rect 8447 35 8448 99
rect 8382 19 8448 35
rect 8382 -45 8383 19
rect 8447 -45 8448 19
rect 8382 -61 8448 -45
rect 8382 -125 8383 -61
rect 8447 -125 8448 -61
rect 8382 -141 8448 -125
rect 8382 -205 8383 -141
rect 8447 -205 8448 -141
rect 8382 -295 8448 -205
rect 8508 -359 8568 671
rect 8628 -299 8688 733
rect 8748 -359 8808 671
rect 8868 -299 8928 733
rect 8988 579 9054 733
rect 8988 515 8989 579
rect 9053 515 9054 579
rect 8988 499 9054 515
rect 8988 435 8989 499
rect 9053 435 9054 499
rect 8988 419 9054 435
rect 8988 355 8989 419
rect 9053 355 9054 419
rect 8988 339 9054 355
rect 8988 275 8989 339
rect 9053 275 9054 339
rect 8988 259 9054 275
rect 8988 195 8989 259
rect 9053 195 9054 259
rect 8988 179 9054 195
rect 8988 115 8989 179
rect 9053 115 9054 179
rect 8988 99 9054 115
rect 8988 35 8989 99
rect 9053 35 9054 99
rect 8988 19 9054 35
rect 8988 -45 8989 19
rect 9053 -45 9054 19
rect 8988 -61 9054 -45
rect 8988 -125 8989 -61
rect 9053 -125 9054 -61
rect 8988 -141 9054 -125
rect 8988 -205 8989 -141
rect 9053 -205 9054 -141
rect 8988 -295 9054 -205
rect 9114 -359 9174 671
rect 9234 -299 9294 733
rect 9354 -359 9414 671
rect 9474 -299 9534 733
rect 9594 579 9660 733
rect 9594 515 9595 579
rect 9659 515 9660 579
rect 9594 499 9660 515
rect 9594 435 9595 499
rect 9659 435 9660 499
rect 9594 419 9660 435
rect 9594 355 9595 419
rect 9659 355 9660 419
rect 9594 339 9660 355
rect 9594 275 9595 339
rect 9659 275 9660 339
rect 9594 259 9660 275
rect 9594 195 9595 259
rect 9659 195 9660 259
rect 9594 179 9660 195
rect 9594 115 9595 179
rect 9659 115 9660 179
rect 9594 99 9660 115
rect 9594 35 9595 99
rect 9659 35 9660 99
rect 9594 19 9660 35
rect 9594 -45 9595 19
rect 9659 -45 9660 19
rect 9594 -61 9660 -45
rect 9594 -125 9595 -61
rect 9659 -125 9660 -61
rect 9594 -141 9660 -125
rect 9594 -205 9595 -141
rect 9659 -205 9660 -141
rect 9594 -295 9660 -205
rect 9720 -359 9780 671
rect 9840 -299 9900 733
rect 9960 -359 10020 671
rect 10080 -299 10140 733
rect 10200 579 10266 733
rect 10200 515 10201 579
rect 10265 515 10266 579
rect 10200 499 10266 515
rect 10200 435 10201 499
rect 10265 435 10266 499
rect 10200 419 10266 435
rect 10200 355 10201 419
rect 10265 355 10266 419
rect 10200 339 10266 355
rect 10200 275 10201 339
rect 10265 275 10266 339
rect 10200 259 10266 275
rect 10200 195 10201 259
rect 10265 195 10266 259
rect 10200 179 10266 195
rect 10200 115 10201 179
rect 10265 115 10266 179
rect 10200 99 10266 115
rect 10200 35 10201 99
rect 10265 35 10266 99
rect 10200 19 10266 35
rect 10200 -45 10201 19
rect 10265 -45 10266 19
rect 10200 -61 10266 -45
rect 10200 -125 10201 -61
rect 10265 -125 10266 -61
rect 10200 -141 10266 -125
rect 10200 -205 10201 -141
rect 10265 -205 10266 -141
rect 10200 -295 10266 -205
rect 10326 1739 10392 1829
rect 10326 1675 10327 1739
rect 10391 1675 10392 1739
rect 10326 1659 10392 1675
rect 10326 1595 10327 1659
rect 10391 1595 10392 1659
rect 10326 1579 10392 1595
rect 10326 1515 10327 1579
rect 10391 1515 10392 1579
rect 10326 1499 10392 1515
rect 10326 1435 10327 1499
rect 10391 1435 10392 1499
rect 10326 1419 10392 1435
rect 10326 1355 10327 1419
rect 10391 1355 10392 1419
rect 10326 1339 10392 1355
rect 10326 1275 10327 1339
rect 10391 1275 10392 1339
rect 10326 1259 10392 1275
rect 10326 1195 10327 1259
rect 10391 1195 10392 1259
rect 10326 1179 10392 1195
rect 10326 1115 10327 1179
rect 10391 1115 10392 1179
rect 10326 1099 10392 1115
rect 10326 1035 10327 1099
rect 10391 1035 10392 1099
rect 10326 1019 10392 1035
rect 10326 955 10327 1019
rect 10391 955 10392 1019
rect 10326 801 10392 955
rect 10452 801 10512 1833
rect 10572 863 10632 1893
rect 10692 801 10752 1833
rect 10812 863 10872 1893
rect 10932 1739 10998 1829
rect 10932 1675 10933 1739
rect 10997 1675 10998 1739
rect 10932 1659 10998 1675
rect 10932 1595 10933 1659
rect 10997 1595 10998 1659
rect 10932 1579 10998 1595
rect 10932 1515 10933 1579
rect 10997 1515 10998 1579
rect 10932 1499 10998 1515
rect 10932 1435 10933 1499
rect 10997 1435 10998 1499
rect 10932 1419 10998 1435
rect 10932 1355 10933 1419
rect 10997 1355 10998 1419
rect 10932 1339 10998 1355
rect 10932 1275 10933 1339
rect 10997 1275 10998 1339
rect 10932 1259 10998 1275
rect 10932 1195 10933 1259
rect 10997 1195 10998 1259
rect 10932 1179 10998 1195
rect 10932 1115 10933 1179
rect 10997 1115 10998 1179
rect 10932 1099 10998 1115
rect 10932 1035 10933 1099
rect 10997 1035 10998 1099
rect 10932 1019 10998 1035
rect 10932 955 10933 1019
rect 10997 955 10998 1019
rect 10932 801 10998 955
rect 11058 801 11118 1833
rect 11178 863 11238 1893
rect 11298 801 11358 1833
rect 11418 863 11478 1893
rect 11538 1739 11604 1829
rect 11538 1675 11539 1739
rect 11603 1675 11604 1739
rect 11538 1659 11604 1675
rect 11538 1595 11539 1659
rect 11603 1595 11604 1659
rect 11538 1579 11604 1595
rect 11538 1515 11539 1579
rect 11603 1515 11604 1579
rect 11538 1499 11604 1515
rect 11538 1435 11539 1499
rect 11603 1435 11604 1499
rect 11538 1419 11604 1435
rect 11538 1355 11539 1419
rect 11603 1355 11604 1419
rect 11538 1339 11604 1355
rect 11538 1275 11539 1339
rect 11603 1275 11604 1339
rect 11538 1259 11604 1275
rect 11538 1195 11539 1259
rect 11603 1195 11604 1259
rect 11538 1179 11604 1195
rect 11538 1115 11539 1179
rect 11603 1115 11604 1179
rect 11538 1099 11604 1115
rect 11538 1035 11539 1099
rect 11603 1035 11604 1099
rect 11538 1019 11604 1035
rect 11538 955 11539 1019
rect 11603 955 11604 1019
rect 11538 801 11604 955
rect 11664 801 11724 1833
rect 11784 863 11844 1893
rect 11904 801 11964 1833
rect 12024 863 12084 1893
rect 12144 1739 12210 1829
rect 12144 1675 12145 1739
rect 12209 1675 12210 1739
rect 12144 1659 12210 1675
rect 12144 1595 12145 1659
rect 12209 1595 12210 1659
rect 12144 1579 12210 1595
rect 12144 1515 12145 1579
rect 12209 1515 12210 1579
rect 12144 1499 12210 1515
rect 12144 1435 12145 1499
rect 12209 1435 12210 1499
rect 12144 1419 12210 1435
rect 12144 1355 12145 1419
rect 12209 1355 12210 1419
rect 12144 1339 12210 1355
rect 12144 1275 12145 1339
rect 12209 1275 12210 1339
rect 12144 1259 12210 1275
rect 12144 1195 12145 1259
rect 12209 1195 12210 1259
rect 12144 1179 12210 1195
rect 12144 1115 12145 1179
rect 12209 1115 12210 1179
rect 12144 1099 12210 1115
rect 12144 1035 12145 1099
rect 12209 1035 12210 1099
rect 12144 1019 12210 1035
rect 12144 955 12145 1019
rect 12209 955 12210 1019
rect 12144 801 12210 955
rect 12270 801 12330 1833
rect 12390 863 12450 1893
rect 12510 801 12570 1833
rect 12630 863 12690 1893
rect 12750 1739 12816 1829
rect 12750 1675 12751 1739
rect 12815 1675 12816 1739
rect 12750 1659 12816 1675
rect 12750 1595 12751 1659
rect 12815 1595 12816 1659
rect 12750 1579 12816 1595
rect 12750 1515 12751 1579
rect 12815 1515 12816 1579
rect 12750 1499 12816 1515
rect 12750 1435 12751 1499
rect 12815 1435 12816 1499
rect 12750 1419 12816 1435
rect 12750 1355 12751 1419
rect 12815 1355 12816 1419
rect 12750 1339 12816 1355
rect 12750 1275 12751 1339
rect 12815 1275 12816 1339
rect 12750 1259 12816 1275
rect 12750 1195 12751 1259
rect 12815 1195 12816 1259
rect 12750 1179 12816 1195
rect 12750 1115 12751 1179
rect 12815 1115 12816 1179
rect 12750 1099 12816 1115
rect 12750 1035 12751 1099
rect 12815 1035 12816 1099
rect 12750 1019 12816 1035
rect 12750 955 12751 1019
rect 12815 955 12816 1019
rect 12750 801 12816 955
rect 12876 801 12936 1833
rect 12996 863 13056 1893
rect 13116 801 13176 1833
rect 13236 863 13296 1893
rect 13356 1739 13422 1829
rect 13356 1675 13357 1739
rect 13421 1675 13422 1739
rect 13356 1659 13422 1675
rect 13356 1595 13357 1659
rect 13421 1595 13422 1659
rect 13356 1579 13422 1595
rect 13356 1515 13357 1579
rect 13421 1515 13422 1579
rect 13356 1499 13422 1515
rect 13356 1435 13357 1499
rect 13421 1435 13422 1499
rect 13356 1419 13422 1435
rect 13356 1355 13357 1419
rect 13421 1355 13422 1419
rect 13356 1339 13422 1355
rect 13356 1275 13357 1339
rect 13421 1275 13422 1339
rect 13356 1259 13422 1275
rect 13356 1195 13357 1259
rect 13421 1195 13422 1259
rect 13356 1179 13422 1195
rect 13356 1115 13357 1179
rect 13421 1115 13422 1179
rect 13356 1099 13422 1115
rect 13356 1035 13357 1099
rect 13421 1035 13422 1099
rect 13356 1019 13422 1035
rect 13356 955 13357 1019
rect 13421 955 13422 1019
rect 13356 801 13422 955
rect 13482 801 13542 1833
rect 13602 863 13662 1893
rect 13722 801 13782 1833
rect 13842 863 13902 1893
rect 13962 1739 14028 1829
rect 13962 1675 13963 1739
rect 14027 1675 14028 1739
rect 13962 1659 14028 1675
rect 13962 1595 13963 1659
rect 14027 1595 14028 1659
rect 13962 1579 14028 1595
rect 13962 1515 13963 1579
rect 14027 1515 14028 1579
rect 13962 1499 14028 1515
rect 13962 1435 13963 1499
rect 14027 1435 14028 1499
rect 13962 1419 14028 1435
rect 13962 1355 13963 1419
rect 14027 1355 14028 1419
rect 13962 1339 14028 1355
rect 13962 1275 13963 1339
rect 14027 1275 14028 1339
rect 13962 1259 14028 1275
rect 13962 1195 13963 1259
rect 14027 1195 14028 1259
rect 13962 1179 14028 1195
rect 13962 1115 13963 1179
rect 14027 1115 14028 1179
rect 13962 1099 14028 1115
rect 13962 1035 13963 1099
rect 14027 1035 14028 1099
rect 13962 1019 14028 1035
rect 13962 955 13963 1019
rect 14027 955 14028 1019
rect 13962 801 14028 955
rect 14088 801 14148 1833
rect 14208 863 14268 1893
rect 14328 801 14388 1833
rect 14448 863 14508 1893
rect 14568 1739 14634 1829
rect 14568 1675 14569 1739
rect 14633 1675 14634 1739
rect 14568 1659 14634 1675
rect 14568 1595 14569 1659
rect 14633 1595 14634 1659
rect 14568 1579 14634 1595
rect 14568 1515 14569 1579
rect 14633 1515 14634 1579
rect 14568 1499 14634 1515
rect 14568 1435 14569 1499
rect 14633 1435 14634 1499
rect 14568 1419 14634 1435
rect 14568 1355 14569 1419
rect 14633 1355 14634 1419
rect 14568 1339 14634 1355
rect 14568 1275 14569 1339
rect 14633 1275 14634 1339
rect 14568 1259 14634 1275
rect 14568 1195 14569 1259
rect 14633 1195 14634 1259
rect 14568 1179 14634 1195
rect 14568 1115 14569 1179
rect 14633 1115 14634 1179
rect 14568 1099 14634 1115
rect 14568 1035 14569 1099
rect 14633 1035 14634 1099
rect 14568 1019 14634 1035
rect 14568 955 14569 1019
rect 14633 955 14634 1019
rect 14568 801 14634 955
rect 14694 801 14754 1833
rect 14814 863 14874 1893
rect 14934 801 14994 1833
rect 15054 863 15114 1893
rect 15174 1739 15240 1829
rect 15174 1675 15175 1739
rect 15239 1675 15240 1739
rect 15174 1659 15240 1675
rect 15174 1595 15175 1659
rect 15239 1595 15240 1659
rect 15174 1579 15240 1595
rect 15174 1515 15175 1579
rect 15239 1515 15240 1579
rect 15174 1499 15240 1515
rect 15174 1435 15175 1499
rect 15239 1435 15240 1499
rect 15174 1419 15240 1435
rect 15174 1355 15175 1419
rect 15239 1355 15240 1419
rect 15174 1339 15240 1355
rect 15174 1275 15175 1339
rect 15239 1275 15240 1339
rect 15174 1259 15240 1275
rect 15174 1195 15175 1259
rect 15239 1195 15240 1259
rect 15174 1179 15240 1195
rect 15174 1115 15175 1179
rect 15239 1115 15240 1179
rect 15174 1099 15240 1115
rect 15174 1035 15175 1099
rect 15239 1035 15240 1099
rect 15174 1019 15240 1035
rect 15174 955 15175 1019
rect 15239 955 15240 1019
rect 15174 801 15240 955
rect 15300 801 15360 1833
rect 15420 863 15480 1893
rect 15540 801 15600 1833
rect 15660 863 15720 1893
rect 15780 1820 15846 1829
rect 15780 1764 15785 1820
rect 15841 1764 15846 1820
rect 15780 1739 15846 1764
rect 15780 1675 15781 1739
rect 15845 1675 15846 1739
rect 15780 1659 15846 1675
rect 15780 1595 15781 1659
rect 15845 1595 15846 1659
rect 15780 1579 15846 1595
rect 15780 1515 15781 1579
rect 15845 1515 15846 1579
rect 15780 1499 15846 1515
rect 15780 1435 15781 1499
rect 15845 1435 15846 1499
rect 15780 1419 15846 1435
rect 15780 1355 15781 1419
rect 15845 1355 15846 1419
rect 15780 1339 15846 1355
rect 15780 1275 15781 1339
rect 15845 1275 15846 1339
rect 15780 1259 15846 1275
rect 15780 1195 15781 1259
rect 15845 1195 15846 1259
rect 15780 1179 15846 1195
rect 15780 1115 15781 1179
rect 15845 1115 15846 1179
rect 15780 1099 15846 1115
rect 15780 1035 15781 1099
rect 15845 1035 15846 1099
rect 15780 1019 15846 1035
rect 15780 955 15781 1019
rect 15845 955 15846 1019
rect 15780 801 15846 955
rect 15906 801 15966 1833
rect 16026 863 16086 1893
rect 16146 801 16206 1833
rect 16266 863 16326 1893
rect 16386 1819 16452 1829
rect 16386 1763 16391 1819
rect 16447 1763 16452 1819
rect 16386 1739 16452 1763
rect 16386 1675 16387 1739
rect 16451 1675 16452 1739
rect 16386 1659 16452 1675
rect 16386 1595 16387 1659
rect 16451 1595 16452 1659
rect 16386 1579 16452 1595
rect 16386 1515 16387 1579
rect 16451 1515 16452 1579
rect 16386 1499 16452 1515
rect 16386 1435 16387 1499
rect 16451 1435 16452 1499
rect 16386 1419 16452 1435
rect 16386 1355 16387 1419
rect 16451 1355 16452 1419
rect 16386 1339 16452 1355
rect 16386 1275 16387 1339
rect 16451 1275 16452 1339
rect 16386 1259 16452 1275
rect 16386 1195 16387 1259
rect 16451 1195 16452 1259
rect 16386 1179 16452 1195
rect 16386 1115 16387 1179
rect 16451 1115 16452 1179
rect 16386 1099 16452 1115
rect 16386 1035 16387 1099
rect 16451 1035 16452 1099
rect 16386 1019 16452 1035
rect 16386 955 16387 1019
rect 16451 955 16452 1019
rect 16386 801 16452 955
rect 16512 801 16572 1833
rect 16632 863 16692 1893
rect 16752 801 16812 1833
rect 16872 863 16932 1893
rect 16992 1819 17058 1829
rect 16992 1763 16997 1819
rect 17053 1763 17058 1819
rect 16992 1739 17058 1763
rect 16992 1675 16993 1739
rect 17057 1675 17058 1739
rect 16992 1659 17058 1675
rect 16992 1595 16993 1659
rect 17057 1595 17058 1659
rect 16992 1579 17058 1595
rect 16992 1515 16993 1579
rect 17057 1515 17058 1579
rect 16992 1499 17058 1515
rect 16992 1435 16993 1499
rect 17057 1435 17058 1499
rect 16992 1419 17058 1435
rect 16992 1355 16993 1419
rect 17057 1355 17058 1419
rect 16992 1339 17058 1355
rect 16992 1275 16993 1339
rect 17057 1275 17058 1339
rect 16992 1259 17058 1275
rect 16992 1195 16993 1259
rect 17057 1195 17058 1259
rect 16992 1179 17058 1195
rect 16992 1115 16993 1179
rect 17057 1115 17058 1179
rect 16992 1099 17058 1115
rect 16992 1035 16993 1099
rect 17057 1035 17058 1099
rect 16992 1019 17058 1035
rect 16992 955 16993 1019
rect 17057 955 17058 1019
rect 16992 801 17058 955
rect 17118 801 17178 1833
rect 17238 863 17298 1893
rect 17358 801 17418 1833
rect 17478 863 17538 1893
rect 17598 1818 17664 1829
rect 17598 1762 17603 1818
rect 17659 1762 17664 1818
rect 17598 1739 17664 1762
rect 17598 1675 17599 1739
rect 17663 1675 17664 1739
rect 17598 1659 17664 1675
rect 17598 1595 17599 1659
rect 17663 1595 17664 1659
rect 17598 1579 17664 1595
rect 17598 1515 17599 1579
rect 17663 1515 17664 1579
rect 17598 1499 17664 1515
rect 17598 1435 17599 1499
rect 17663 1435 17664 1499
rect 17598 1419 17664 1435
rect 17598 1355 17599 1419
rect 17663 1355 17664 1419
rect 17598 1339 17664 1355
rect 17598 1275 17599 1339
rect 17663 1275 17664 1339
rect 17598 1259 17664 1275
rect 17598 1195 17599 1259
rect 17663 1195 17664 1259
rect 17598 1179 17664 1195
rect 17598 1115 17599 1179
rect 17663 1115 17664 1179
rect 17598 1099 17664 1115
rect 17598 1035 17599 1099
rect 17663 1035 17664 1099
rect 17598 1019 17664 1035
rect 17598 955 17599 1019
rect 17663 955 17664 1019
rect 17598 801 17664 955
rect 17724 801 17784 1833
rect 17844 863 17904 1893
rect 17964 801 18024 1833
rect 18084 863 18144 1893
rect 18204 1818 18270 1829
rect 18204 1762 18209 1818
rect 18265 1762 18270 1818
rect 18204 1739 18270 1762
rect 18204 1675 18205 1739
rect 18269 1675 18270 1739
rect 18204 1659 18270 1675
rect 18204 1595 18205 1659
rect 18269 1595 18270 1659
rect 18204 1579 18270 1595
rect 18204 1515 18205 1579
rect 18269 1515 18270 1579
rect 18204 1499 18270 1515
rect 18204 1435 18205 1499
rect 18269 1435 18270 1499
rect 18204 1419 18270 1435
rect 18204 1355 18205 1419
rect 18269 1355 18270 1419
rect 18204 1339 18270 1355
rect 18204 1275 18205 1339
rect 18269 1275 18270 1339
rect 18204 1259 18270 1275
rect 18204 1195 18205 1259
rect 18269 1195 18270 1259
rect 18204 1179 18270 1195
rect 18204 1115 18205 1179
rect 18269 1115 18270 1179
rect 18204 1099 18270 1115
rect 18204 1035 18205 1099
rect 18269 1035 18270 1099
rect 18204 1019 18270 1035
rect 18204 955 18205 1019
rect 18269 955 18270 1019
rect 18204 801 18270 955
rect 18330 801 18390 1833
rect 18450 863 18510 1893
rect 18570 801 18630 1833
rect 18690 863 18750 1893
rect 18810 1818 18876 1829
rect 18810 1762 18815 1818
rect 18871 1762 18876 1818
rect 18810 1739 18876 1762
rect 18810 1675 18811 1739
rect 18875 1675 18876 1739
rect 18810 1659 18876 1675
rect 18810 1595 18811 1659
rect 18875 1595 18876 1659
rect 18810 1579 18876 1595
rect 18810 1515 18811 1579
rect 18875 1515 18876 1579
rect 18810 1499 18876 1515
rect 18810 1435 18811 1499
rect 18875 1435 18876 1499
rect 18810 1419 18876 1435
rect 18810 1355 18811 1419
rect 18875 1355 18876 1419
rect 18810 1339 18876 1355
rect 18810 1275 18811 1339
rect 18875 1275 18876 1339
rect 18810 1259 18876 1275
rect 18810 1195 18811 1259
rect 18875 1195 18876 1259
rect 18810 1179 18876 1195
rect 18810 1115 18811 1179
rect 18875 1115 18876 1179
rect 18810 1099 18876 1115
rect 18810 1035 18811 1099
rect 18875 1035 18876 1099
rect 18810 1019 18876 1035
rect 18810 955 18811 1019
rect 18875 955 18876 1019
rect 18810 801 18876 955
rect 18936 801 18996 1833
rect 19056 863 19116 1893
rect 19176 801 19236 1833
rect 19296 863 19356 1893
rect 19416 1817 19482 1829
rect 19416 1761 19421 1817
rect 19477 1761 19482 1817
rect 19416 1739 19482 1761
rect 19416 1675 19417 1739
rect 19481 1675 19482 1739
rect 19416 1659 19482 1675
rect 19416 1595 19417 1659
rect 19481 1595 19482 1659
rect 19416 1579 19482 1595
rect 19416 1515 19417 1579
rect 19481 1515 19482 1579
rect 19416 1499 19482 1515
rect 19416 1435 19417 1499
rect 19481 1435 19482 1499
rect 19416 1419 19482 1435
rect 19416 1355 19417 1419
rect 19481 1355 19482 1419
rect 19416 1339 19482 1355
rect 19416 1275 19417 1339
rect 19481 1275 19482 1339
rect 19416 1259 19482 1275
rect 19416 1195 19417 1259
rect 19481 1195 19482 1259
rect 19416 1179 19482 1195
rect 19416 1115 19417 1179
rect 19481 1115 19482 1179
rect 19416 1099 19482 1115
rect 19416 1035 19417 1099
rect 19481 1035 19482 1099
rect 19416 1019 19482 1035
rect 19416 955 19417 1019
rect 19481 955 19482 1019
rect 19416 801 19482 955
rect 19542 801 19602 1833
rect 19662 863 19722 1893
rect 19782 801 19842 1833
rect 19902 863 19962 1893
rect 20022 1817 20088 1829
rect 20022 1761 20027 1817
rect 20083 1761 20088 1817
rect 20022 1739 20088 1761
rect 20022 1675 20023 1739
rect 20087 1675 20088 1739
rect 20022 1659 20088 1675
rect 20022 1595 20023 1659
rect 20087 1595 20088 1659
rect 20022 1579 20088 1595
rect 20022 1515 20023 1579
rect 20087 1515 20088 1579
rect 20022 1499 20088 1515
rect 20022 1435 20023 1499
rect 20087 1435 20088 1499
rect 20022 1419 20088 1435
rect 20022 1355 20023 1419
rect 20087 1355 20088 1419
rect 20022 1339 20088 1355
rect 20022 1275 20023 1339
rect 20087 1275 20088 1339
rect 20022 1259 20088 1275
rect 20022 1195 20023 1259
rect 20087 1195 20088 1259
rect 20022 1179 20088 1195
rect 20022 1115 20023 1179
rect 20087 1115 20088 1179
rect 20022 1099 20088 1115
rect 20022 1035 20023 1099
rect 20087 1035 20088 1099
rect 20022 1019 20088 1035
rect 20022 955 20023 1019
rect 20087 955 20088 1019
rect 20022 801 20088 955
rect 10326 799 20088 801
rect 10326 735 10430 799
rect 10494 735 10510 799
rect 10574 735 10590 799
rect 10654 735 10670 799
rect 10734 735 10750 799
rect 10814 735 10830 799
rect 10894 735 11036 799
rect 11100 735 11116 799
rect 11180 735 11196 799
rect 11260 735 11276 799
rect 11340 735 11356 799
rect 11420 735 11436 799
rect 11500 735 11642 799
rect 11706 735 11722 799
rect 11786 735 11802 799
rect 11866 735 11882 799
rect 11946 735 11962 799
rect 12026 735 12042 799
rect 12106 735 12248 799
rect 12312 735 12328 799
rect 12392 735 12408 799
rect 12472 735 12488 799
rect 12552 735 12568 799
rect 12632 735 12648 799
rect 12712 735 12854 799
rect 12918 735 12934 799
rect 12998 735 13014 799
rect 13078 735 13094 799
rect 13158 735 13174 799
rect 13238 735 13254 799
rect 13318 735 13460 799
rect 13524 735 13540 799
rect 13604 735 13620 799
rect 13684 735 13700 799
rect 13764 735 13780 799
rect 13844 735 13860 799
rect 13924 735 14066 799
rect 14130 735 14146 799
rect 14210 735 14226 799
rect 14290 735 14306 799
rect 14370 735 14386 799
rect 14450 735 14466 799
rect 14530 735 14672 799
rect 14736 735 14752 799
rect 14816 735 14832 799
rect 14896 735 14912 799
rect 14976 735 14992 799
rect 15056 735 15072 799
rect 15136 735 15278 799
rect 15342 735 15358 799
rect 15422 735 15438 799
rect 15502 735 15518 799
rect 15582 735 15598 799
rect 15662 735 15678 799
rect 15742 735 15884 799
rect 15948 735 15964 799
rect 16028 735 16044 799
rect 16108 735 16124 799
rect 16188 735 16204 799
rect 16268 735 16284 799
rect 16348 735 16490 799
rect 16554 735 16570 799
rect 16634 735 16650 799
rect 16714 735 16730 799
rect 16794 735 16810 799
rect 16874 735 16890 799
rect 16954 735 17096 799
rect 17160 735 17176 799
rect 17240 735 17256 799
rect 17320 735 17336 799
rect 17400 735 17416 799
rect 17480 735 17496 799
rect 17560 735 17702 799
rect 17766 735 17782 799
rect 17846 735 17862 799
rect 17926 735 17942 799
rect 18006 735 18022 799
rect 18086 735 18102 799
rect 18166 735 18308 799
rect 18372 735 18388 799
rect 18452 735 18468 799
rect 18532 735 18548 799
rect 18612 735 18628 799
rect 18692 735 18708 799
rect 18772 735 18914 799
rect 18978 735 18994 799
rect 19058 735 19074 799
rect 19138 735 19154 799
rect 19218 735 19234 799
rect 19298 735 19314 799
rect 19378 735 19520 799
rect 19584 735 19600 799
rect 19664 735 19680 799
rect 19744 735 19760 799
rect 19824 735 19840 799
rect 19904 735 19920 799
rect 19984 735 20088 799
rect 10326 733 20088 735
rect 10326 579 10392 733
rect 10326 515 10327 579
rect 10391 515 10392 579
rect 10326 499 10392 515
rect 10326 435 10327 499
rect 10391 435 10392 499
rect 10326 419 10392 435
rect 10326 355 10327 419
rect 10391 355 10392 419
rect 10326 339 10392 355
rect 10326 275 10327 339
rect 10391 275 10392 339
rect 10326 259 10392 275
rect 10326 195 10327 259
rect 10391 195 10392 259
rect 10326 179 10392 195
rect 10326 115 10327 179
rect 10391 115 10392 179
rect 10326 99 10392 115
rect 10326 35 10327 99
rect 10391 35 10392 99
rect 10326 19 10392 35
rect 10326 -45 10327 19
rect 10391 -45 10392 19
rect 10326 -61 10392 -45
rect 10326 -125 10327 -61
rect 10391 -125 10392 -61
rect 10326 -141 10392 -125
rect 10326 -205 10327 -141
rect 10391 -205 10392 -141
rect 10326 -295 10392 -205
rect 10452 -359 10512 671
rect 10572 -299 10632 733
rect 10692 -359 10752 671
rect 10812 -299 10872 733
rect 10932 579 10998 733
rect 10932 515 10933 579
rect 10997 515 10998 579
rect 10932 499 10998 515
rect 10932 435 10933 499
rect 10997 435 10998 499
rect 10932 419 10998 435
rect 10932 355 10933 419
rect 10997 355 10998 419
rect 10932 339 10998 355
rect 10932 275 10933 339
rect 10997 275 10998 339
rect 10932 259 10998 275
rect 10932 195 10933 259
rect 10997 195 10998 259
rect 10932 179 10998 195
rect 10932 115 10933 179
rect 10997 115 10998 179
rect 10932 99 10998 115
rect 10932 35 10933 99
rect 10997 35 10998 99
rect 10932 19 10998 35
rect 10932 -45 10933 19
rect 10997 -45 10998 19
rect 10932 -61 10998 -45
rect 10932 -125 10933 -61
rect 10997 -125 10998 -61
rect 10932 -141 10998 -125
rect 10932 -205 10933 -141
rect 10997 -205 10998 -141
rect 10932 -295 10998 -205
rect 11058 -359 11118 671
rect 11178 -299 11238 733
rect 11298 -359 11358 671
rect 11418 -299 11478 733
rect 11538 579 11604 733
rect 11538 515 11539 579
rect 11603 515 11604 579
rect 11538 499 11604 515
rect 11538 435 11539 499
rect 11603 435 11604 499
rect 11538 419 11604 435
rect 11538 355 11539 419
rect 11603 355 11604 419
rect 11538 339 11604 355
rect 11538 275 11539 339
rect 11603 275 11604 339
rect 11538 259 11604 275
rect 11538 195 11539 259
rect 11603 195 11604 259
rect 11538 179 11604 195
rect 11538 115 11539 179
rect 11603 115 11604 179
rect 11538 99 11604 115
rect 11538 35 11539 99
rect 11603 35 11604 99
rect 11538 19 11604 35
rect 11538 -45 11539 19
rect 11603 -45 11604 19
rect 11538 -61 11604 -45
rect 11538 -125 11539 -61
rect 11603 -125 11604 -61
rect 11538 -141 11604 -125
rect 11538 -205 11539 -141
rect 11603 -205 11604 -141
rect 11538 -295 11604 -205
rect 11664 -359 11724 671
rect 11784 -299 11844 733
rect 11904 -359 11964 671
rect 12024 -299 12084 733
rect 12144 579 12210 733
rect 12144 515 12145 579
rect 12209 515 12210 579
rect 12144 499 12210 515
rect 12144 435 12145 499
rect 12209 435 12210 499
rect 12144 419 12210 435
rect 12144 355 12145 419
rect 12209 355 12210 419
rect 12144 339 12210 355
rect 12144 275 12145 339
rect 12209 275 12210 339
rect 12144 259 12210 275
rect 12144 195 12145 259
rect 12209 195 12210 259
rect 12144 179 12210 195
rect 12144 115 12145 179
rect 12209 115 12210 179
rect 12144 99 12210 115
rect 12144 35 12145 99
rect 12209 35 12210 99
rect 12144 19 12210 35
rect 12144 -45 12145 19
rect 12209 -45 12210 19
rect 12144 -61 12210 -45
rect 12144 -125 12145 -61
rect 12209 -125 12210 -61
rect 12144 -141 12210 -125
rect 12144 -205 12145 -141
rect 12209 -205 12210 -141
rect 12144 -295 12210 -205
rect 12270 -359 12330 671
rect 12390 -299 12450 733
rect 12510 -359 12570 671
rect 12630 -299 12690 733
rect 12750 579 12816 733
rect 12750 515 12751 579
rect 12815 515 12816 579
rect 12750 499 12816 515
rect 12750 435 12751 499
rect 12815 435 12816 499
rect 12750 419 12816 435
rect 12750 355 12751 419
rect 12815 355 12816 419
rect 12750 339 12816 355
rect 12750 275 12751 339
rect 12815 275 12816 339
rect 12750 259 12816 275
rect 12750 195 12751 259
rect 12815 195 12816 259
rect 12750 179 12816 195
rect 12750 115 12751 179
rect 12815 115 12816 179
rect 12750 99 12816 115
rect 12750 35 12751 99
rect 12815 35 12816 99
rect 12750 19 12816 35
rect 12750 -45 12751 19
rect 12815 -45 12816 19
rect 12750 -61 12816 -45
rect 12750 -125 12751 -61
rect 12815 -125 12816 -61
rect 12750 -141 12816 -125
rect 12750 -205 12751 -141
rect 12815 -205 12816 -141
rect 12750 -295 12816 -205
rect 12876 -359 12936 671
rect 12996 -299 13056 733
rect 13116 -359 13176 671
rect 13236 -299 13296 733
rect 13356 579 13422 733
rect 13356 515 13357 579
rect 13421 515 13422 579
rect 13356 499 13422 515
rect 13356 435 13357 499
rect 13421 435 13422 499
rect 13356 419 13422 435
rect 13356 355 13357 419
rect 13421 355 13422 419
rect 13356 339 13422 355
rect 13356 275 13357 339
rect 13421 275 13422 339
rect 13356 259 13422 275
rect 13356 195 13357 259
rect 13421 195 13422 259
rect 13356 179 13422 195
rect 13356 115 13357 179
rect 13421 115 13422 179
rect 13356 99 13422 115
rect 13356 35 13357 99
rect 13421 35 13422 99
rect 13356 19 13422 35
rect 13356 -45 13357 19
rect 13421 -45 13422 19
rect 13356 -61 13422 -45
rect 13356 -125 13357 -61
rect 13421 -125 13422 -61
rect 13356 -141 13422 -125
rect 13356 -205 13357 -141
rect 13421 -205 13422 -141
rect 13356 -295 13422 -205
rect 13482 -359 13542 671
rect 13602 -299 13662 733
rect 13722 -359 13782 671
rect 13842 -299 13902 733
rect 13962 579 14028 733
rect 13962 515 13963 579
rect 14027 515 14028 579
rect 13962 499 14028 515
rect 13962 435 13963 499
rect 14027 435 14028 499
rect 13962 419 14028 435
rect 13962 355 13963 419
rect 14027 355 14028 419
rect 13962 339 14028 355
rect 13962 275 13963 339
rect 14027 275 14028 339
rect 13962 259 14028 275
rect 13962 195 13963 259
rect 14027 195 14028 259
rect 13962 179 14028 195
rect 13962 115 13963 179
rect 14027 115 14028 179
rect 13962 99 14028 115
rect 13962 35 13963 99
rect 14027 35 14028 99
rect 13962 19 14028 35
rect 13962 -45 13963 19
rect 14027 -45 14028 19
rect 13962 -61 14028 -45
rect 13962 -125 13963 -61
rect 14027 -125 14028 -61
rect 13962 -141 14028 -125
rect 13962 -205 13963 -141
rect 14027 -205 14028 -141
rect 13962 -295 14028 -205
rect 14088 -359 14148 671
rect 14208 -299 14268 733
rect 14328 -359 14388 671
rect 14448 -299 14508 733
rect 14568 579 14634 733
rect 14568 515 14569 579
rect 14633 515 14634 579
rect 14568 499 14634 515
rect 14568 435 14569 499
rect 14633 435 14634 499
rect 14568 419 14634 435
rect 14568 355 14569 419
rect 14633 355 14634 419
rect 14568 339 14634 355
rect 14568 275 14569 339
rect 14633 275 14634 339
rect 14568 259 14634 275
rect 14568 195 14569 259
rect 14633 195 14634 259
rect 14568 179 14634 195
rect 14568 115 14569 179
rect 14633 115 14634 179
rect 14568 99 14634 115
rect 14568 35 14569 99
rect 14633 35 14634 99
rect 14568 19 14634 35
rect 14568 -45 14569 19
rect 14633 -45 14634 19
rect 14568 -61 14634 -45
rect 14568 -125 14569 -61
rect 14633 -125 14634 -61
rect 14568 -141 14634 -125
rect 14568 -205 14569 -141
rect 14633 -205 14634 -141
rect 14568 -295 14634 -205
rect 14694 -359 14754 671
rect 14814 -299 14874 733
rect 14934 -359 14994 671
rect 15054 -299 15114 733
rect 15174 579 15240 733
rect 15174 515 15175 579
rect 15239 515 15240 579
rect 15174 499 15240 515
rect 15174 435 15175 499
rect 15239 435 15240 499
rect 15174 419 15240 435
rect 15174 355 15175 419
rect 15239 355 15240 419
rect 15174 339 15240 355
rect 15174 275 15175 339
rect 15239 275 15240 339
rect 15174 259 15240 275
rect 15174 195 15175 259
rect 15239 195 15240 259
rect 15174 179 15240 195
rect 15174 115 15175 179
rect 15239 115 15240 179
rect 15174 99 15240 115
rect 15174 35 15175 99
rect 15239 35 15240 99
rect 15174 19 15240 35
rect 15174 -45 15175 19
rect 15239 -45 15240 19
rect 15174 -61 15240 -45
rect 15174 -125 15175 -61
rect 15239 -125 15240 -61
rect 15174 -141 15240 -125
rect 15174 -205 15175 -141
rect 15239 -205 15240 -141
rect 15174 -295 15240 -205
rect 15300 -359 15360 671
rect 15420 -299 15480 733
rect 15540 -359 15600 671
rect 15660 -299 15720 733
rect 15780 579 15846 733
rect 15780 515 15781 579
rect 15845 515 15846 579
rect 15780 499 15846 515
rect 15780 435 15781 499
rect 15845 435 15846 499
rect 15780 419 15846 435
rect 15780 355 15781 419
rect 15845 355 15846 419
rect 15780 339 15846 355
rect 15780 275 15781 339
rect 15845 275 15846 339
rect 15780 259 15846 275
rect 15780 195 15781 259
rect 15845 195 15846 259
rect 15780 179 15846 195
rect 15780 115 15781 179
rect 15845 115 15846 179
rect 15780 99 15846 115
rect 15780 35 15781 99
rect 15845 35 15846 99
rect 15780 19 15846 35
rect 15780 -45 15781 19
rect 15845 -45 15846 19
rect 15780 -61 15846 -45
rect 15780 -125 15781 -61
rect 15845 -125 15846 -61
rect 15780 -141 15846 -125
rect 15780 -205 15781 -141
rect 15845 -205 15846 -141
rect 15780 -295 15846 -205
rect 15906 -359 15966 671
rect 16026 -299 16086 733
rect 16146 -359 16206 671
rect 16266 -299 16326 733
rect 16386 579 16452 733
rect 16386 515 16387 579
rect 16451 515 16452 579
rect 16386 499 16452 515
rect 16386 435 16387 499
rect 16451 435 16452 499
rect 16386 419 16452 435
rect 16386 355 16387 419
rect 16451 355 16452 419
rect 16386 339 16452 355
rect 16386 275 16387 339
rect 16451 275 16452 339
rect 16386 259 16452 275
rect 16386 195 16387 259
rect 16451 195 16452 259
rect 16386 179 16452 195
rect 16386 115 16387 179
rect 16451 115 16452 179
rect 16386 99 16452 115
rect 16386 35 16387 99
rect 16451 35 16452 99
rect 16386 19 16452 35
rect 16386 -45 16387 19
rect 16451 -45 16452 19
rect 16386 -61 16452 -45
rect 16386 -125 16387 -61
rect 16451 -125 16452 -61
rect 16386 -141 16452 -125
rect 16386 -205 16387 -141
rect 16451 -205 16452 -141
rect 16386 -295 16452 -205
rect 16512 -359 16572 671
rect 16632 -299 16692 733
rect 16752 -359 16812 671
rect 16872 -299 16932 733
rect 16992 579 17058 733
rect 16992 515 16993 579
rect 17057 515 17058 579
rect 16992 499 17058 515
rect 16992 435 16993 499
rect 17057 435 17058 499
rect 16992 419 17058 435
rect 16992 355 16993 419
rect 17057 355 17058 419
rect 16992 339 17058 355
rect 16992 275 16993 339
rect 17057 275 17058 339
rect 16992 259 17058 275
rect 16992 195 16993 259
rect 17057 195 17058 259
rect 16992 179 17058 195
rect 16992 115 16993 179
rect 17057 115 17058 179
rect 16992 99 17058 115
rect 16992 35 16993 99
rect 17057 35 17058 99
rect 16992 19 17058 35
rect 16992 -45 16993 19
rect 17057 -45 17058 19
rect 16992 -61 17058 -45
rect 16992 -125 16993 -61
rect 17057 -125 17058 -61
rect 16992 -141 17058 -125
rect 16992 -205 16993 -141
rect 17057 -205 17058 -141
rect 16992 -295 17058 -205
rect 17118 -359 17178 671
rect 17238 -299 17298 733
rect 17358 -359 17418 671
rect 17478 -299 17538 733
rect 17598 579 17664 733
rect 17598 515 17599 579
rect 17663 515 17664 579
rect 17598 499 17664 515
rect 17598 435 17599 499
rect 17663 435 17664 499
rect 17598 419 17664 435
rect 17598 355 17599 419
rect 17663 355 17664 419
rect 17598 339 17664 355
rect 17598 275 17599 339
rect 17663 275 17664 339
rect 17598 259 17664 275
rect 17598 195 17599 259
rect 17663 195 17664 259
rect 17598 179 17664 195
rect 17598 115 17599 179
rect 17663 115 17664 179
rect 17598 99 17664 115
rect 17598 35 17599 99
rect 17663 35 17664 99
rect 17598 19 17664 35
rect 17598 -45 17599 19
rect 17663 -45 17664 19
rect 17598 -61 17664 -45
rect 17598 -125 17599 -61
rect 17663 -125 17664 -61
rect 17598 -141 17664 -125
rect 17598 -205 17599 -141
rect 17663 -205 17664 -141
rect 17598 -295 17664 -205
rect 17724 -359 17784 671
rect 17844 -299 17904 733
rect 17964 -359 18024 671
rect 18084 -299 18144 733
rect 18204 579 18270 733
rect 18204 515 18205 579
rect 18269 515 18270 579
rect 18204 499 18270 515
rect 18204 435 18205 499
rect 18269 435 18270 499
rect 18204 419 18270 435
rect 18204 355 18205 419
rect 18269 355 18270 419
rect 18204 339 18270 355
rect 18204 275 18205 339
rect 18269 275 18270 339
rect 18204 259 18270 275
rect 18204 195 18205 259
rect 18269 195 18270 259
rect 18204 179 18270 195
rect 18204 115 18205 179
rect 18269 115 18270 179
rect 18204 99 18270 115
rect 18204 35 18205 99
rect 18269 35 18270 99
rect 18204 19 18270 35
rect 18204 -45 18205 19
rect 18269 -45 18270 19
rect 18204 -61 18270 -45
rect 18204 -125 18205 -61
rect 18269 -125 18270 -61
rect 18204 -141 18270 -125
rect 18204 -205 18205 -141
rect 18269 -205 18270 -141
rect 18204 -295 18270 -205
rect 18330 -359 18390 671
rect 18450 -299 18510 733
rect 18570 -359 18630 671
rect 18690 -299 18750 733
rect 18810 579 18876 733
rect 18810 515 18811 579
rect 18875 515 18876 579
rect 18810 499 18876 515
rect 18810 435 18811 499
rect 18875 435 18876 499
rect 18810 419 18876 435
rect 18810 355 18811 419
rect 18875 355 18876 419
rect 18810 339 18876 355
rect 18810 275 18811 339
rect 18875 275 18876 339
rect 18810 259 18876 275
rect 18810 195 18811 259
rect 18875 195 18876 259
rect 18810 179 18876 195
rect 18810 115 18811 179
rect 18875 115 18876 179
rect 18810 99 18876 115
rect 18810 35 18811 99
rect 18875 35 18876 99
rect 18810 19 18876 35
rect 18810 -45 18811 19
rect 18875 -45 18876 19
rect 18810 -61 18876 -45
rect 18810 -125 18811 -61
rect 18875 -125 18876 -61
rect 18810 -141 18876 -125
rect 18810 -205 18811 -141
rect 18875 -205 18876 -141
rect 18810 -295 18876 -205
rect 18936 -359 18996 671
rect 19056 -299 19116 733
rect 19176 -359 19236 671
rect 19296 -299 19356 733
rect 19416 579 19482 733
rect 19416 515 19417 579
rect 19481 515 19482 579
rect 19416 499 19482 515
rect 19416 435 19417 499
rect 19481 435 19482 499
rect 19416 419 19482 435
rect 19416 355 19417 419
rect 19481 355 19482 419
rect 19416 339 19482 355
rect 19416 275 19417 339
rect 19481 275 19482 339
rect 19416 259 19482 275
rect 19416 195 19417 259
rect 19481 195 19482 259
rect 19416 179 19482 195
rect 19416 115 19417 179
rect 19481 115 19482 179
rect 19416 99 19482 115
rect 19416 35 19417 99
rect 19481 35 19482 99
rect 19416 19 19482 35
rect 19416 -45 19417 19
rect 19481 -45 19482 19
rect 19416 -61 19482 -45
rect 19416 -125 19417 -61
rect 19481 -125 19482 -61
rect 19416 -141 19482 -125
rect 19416 -205 19417 -141
rect 19481 -205 19482 -141
rect 19416 -295 19482 -205
rect 19542 -359 19602 671
rect 19662 -299 19722 733
rect 19782 -359 19842 671
rect 19902 -299 19962 733
rect 20022 579 20088 733
rect 20022 515 20023 579
rect 20087 515 20088 579
rect 20022 499 20088 515
rect 20022 435 20023 499
rect 20087 435 20088 499
rect 20022 419 20088 435
rect 20022 355 20023 419
rect 20087 355 20088 419
rect 20022 339 20088 355
rect 20022 275 20023 339
rect 20087 275 20088 339
rect 20022 259 20088 275
rect 20022 195 20023 259
rect 20087 195 20088 259
rect 20022 179 20088 195
rect 20022 115 20023 179
rect 20087 115 20088 179
rect 20022 99 20088 115
rect 20022 35 20023 99
rect 20087 35 20088 99
rect 20022 19 20088 35
rect 20022 -45 20023 19
rect 20087 -45 20088 19
rect 20022 -61 20088 -45
rect 20022 -125 20023 -61
rect 20087 -125 20088 -61
rect 20022 -141 20088 -125
rect 20022 -205 20023 -141
rect 20087 -205 20088 -141
rect 20022 -295 20088 -205
rect 20148 1739 20214 1829
rect 20148 1675 20149 1739
rect 20213 1675 20214 1739
rect 20148 1659 20214 1675
rect 20148 1595 20149 1659
rect 20213 1595 20214 1659
rect 20148 1579 20214 1595
rect 20148 1515 20149 1579
rect 20213 1515 20214 1579
rect 20148 1499 20214 1515
rect 20148 1435 20149 1499
rect 20213 1435 20214 1499
rect 20148 1419 20214 1435
rect 20148 1355 20149 1419
rect 20213 1355 20214 1419
rect 20148 1339 20214 1355
rect 20148 1275 20149 1339
rect 20213 1275 20214 1339
rect 20148 1259 20214 1275
rect 20148 1195 20149 1259
rect 20213 1195 20214 1259
rect 20148 1179 20214 1195
rect 20148 1115 20149 1179
rect 20213 1115 20214 1179
rect 20148 1099 20214 1115
rect 20148 1035 20149 1099
rect 20213 1035 20214 1099
rect 20148 1019 20214 1035
rect 20148 955 20149 1019
rect 20213 955 20214 1019
rect 20148 801 20214 955
rect 20274 801 20334 1833
rect 20394 863 20454 1893
rect 20514 801 20574 1833
rect 20634 863 20694 1893
rect 20754 1739 20820 1829
rect 20754 1675 20755 1739
rect 20819 1675 20820 1739
rect 20754 1659 20820 1675
rect 20754 1595 20755 1659
rect 20819 1595 20820 1659
rect 20754 1579 20820 1595
rect 20754 1515 20755 1579
rect 20819 1515 20820 1579
rect 20754 1499 20820 1515
rect 20754 1435 20755 1499
rect 20819 1435 20820 1499
rect 20754 1419 20820 1435
rect 20754 1355 20755 1419
rect 20819 1355 20820 1419
rect 20754 1339 20820 1355
rect 20754 1275 20755 1339
rect 20819 1275 20820 1339
rect 20754 1259 20820 1275
rect 20754 1195 20755 1259
rect 20819 1195 20820 1259
rect 20754 1179 20820 1195
rect 20754 1115 20755 1179
rect 20819 1115 20820 1179
rect 20754 1099 20820 1115
rect 20754 1035 20755 1099
rect 20819 1035 20820 1099
rect 20754 1019 20820 1035
rect 20754 955 20755 1019
rect 20819 955 20820 1019
rect 20754 801 20820 955
rect 20880 801 20940 1833
rect 21000 863 21060 1893
rect 21120 801 21180 1833
rect 21240 863 21300 1893
rect 21360 1739 21426 1829
rect 21360 1675 21361 1739
rect 21425 1675 21426 1739
rect 21360 1659 21426 1675
rect 21360 1595 21361 1659
rect 21425 1595 21426 1659
rect 21360 1579 21426 1595
rect 21360 1515 21361 1579
rect 21425 1515 21426 1579
rect 21360 1499 21426 1515
rect 21360 1435 21361 1499
rect 21425 1435 21426 1499
rect 21360 1419 21426 1435
rect 21360 1355 21361 1419
rect 21425 1355 21426 1419
rect 21360 1339 21426 1355
rect 21360 1275 21361 1339
rect 21425 1275 21426 1339
rect 21360 1259 21426 1275
rect 21360 1195 21361 1259
rect 21425 1195 21426 1259
rect 21360 1179 21426 1195
rect 21360 1115 21361 1179
rect 21425 1115 21426 1179
rect 21360 1099 21426 1115
rect 21360 1035 21361 1099
rect 21425 1035 21426 1099
rect 21360 1019 21426 1035
rect 21360 955 21361 1019
rect 21425 955 21426 1019
rect 21360 801 21426 955
rect 21486 801 21546 1833
rect 21606 863 21666 1893
rect 21726 801 21786 1833
rect 21846 863 21906 1893
rect 21966 1739 22032 1829
rect 21966 1675 21967 1739
rect 22031 1675 22032 1739
rect 21966 1659 22032 1675
rect 21966 1595 21967 1659
rect 22031 1595 22032 1659
rect 21966 1579 22032 1595
rect 21966 1515 21967 1579
rect 22031 1515 22032 1579
rect 21966 1499 22032 1515
rect 21966 1435 21967 1499
rect 22031 1435 22032 1499
rect 21966 1419 22032 1435
rect 21966 1355 21967 1419
rect 22031 1355 22032 1419
rect 21966 1339 22032 1355
rect 21966 1275 21967 1339
rect 22031 1275 22032 1339
rect 21966 1259 22032 1275
rect 21966 1195 21967 1259
rect 22031 1195 22032 1259
rect 21966 1179 22032 1195
rect 21966 1115 21967 1179
rect 22031 1115 22032 1179
rect 21966 1099 22032 1115
rect 21966 1035 21967 1099
rect 22031 1035 22032 1099
rect 21966 1019 22032 1035
rect 21966 955 21967 1019
rect 22031 955 22032 1019
rect 21966 801 22032 955
rect 22092 801 22152 1833
rect 22212 863 22272 1893
rect 22332 801 22392 1833
rect 22452 863 22512 1893
rect 22572 1739 22638 1829
rect 22572 1675 22573 1739
rect 22637 1675 22638 1739
rect 22572 1659 22638 1675
rect 22572 1595 22573 1659
rect 22637 1595 22638 1659
rect 22572 1579 22638 1595
rect 22572 1515 22573 1579
rect 22637 1515 22638 1579
rect 22572 1499 22638 1515
rect 22572 1435 22573 1499
rect 22637 1435 22638 1499
rect 22572 1419 22638 1435
rect 22572 1355 22573 1419
rect 22637 1355 22638 1419
rect 22572 1339 22638 1355
rect 22572 1275 22573 1339
rect 22637 1275 22638 1339
rect 22572 1259 22638 1275
rect 22572 1195 22573 1259
rect 22637 1195 22638 1259
rect 22572 1179 22638 1195
rect 22572 1115 22573 1179
rect 22637 1115 22638 1179
rect 22572 1099 22638 1115
rect 22572 1035 22573 1099
rect 22637 1035 22638 1099
rect 22572 1019 22638 1035
rect 22572 955 22573 1019
rect 22637 955 22638 1019
rect 22572 801 22638 955
rect 22698 801 22758 1833
rect 22818 863 22878 1893
rect 22938 801 22998 1833
rect 23058 863 23118 1893
rect 23178 1739 23244 1829
rect 23178 1675 23179 1739
rect 23243 1675 23244 1739
rect 23178 1659 23244 1675
rect 23178 1595 23179 1659
rect 23243 1595 23244 1659
rect 23178 1579 23244 1595
rect 23178 1515 23179 1579
rect 23243 1515 23244 1579
rect 23178 1499 23244 1515
rect 23178 1435 23179 1499
rect 23243 1435 23244 1499
rect 23178 1419 23244 1435
rect 23178 1355 23179 1419
rect 23243 1355 23244 1419
rect 23178 1339 23244 1355
rect 23178 1275 23179 1339
rect 23243 1275 23244 1339
rect 23178 1259 23244 1275
rect 23178 1195 23179 1259
rect 23243 1195 23244 1259
rect 23178 1179 23244 1195
rect 23178 1115 23179 1179
rect 23243 1115 23244 1179
rect 23178 1099 23244 1115
rect 23178 1035 23179 1099
rect 23243 1035 23244 1099
rect 23178 1019 23244 1035
rect 23178 955 23179 1019
rect 23243 955 23244 1019
rect 23178 801 23244 955
rect 23304 801 23364 1833
rect 23424 863 23484 1893
rect 23544 801 23604 1833
rect 23664 863 23724 1893
rect 23784 1739 23850 1829
rect 23784 1675 23785 1739
rect 23849 1675 23850 1739
rect 23784 1659 23850 1675
rect 23784 1595 23785 1659
rect 23849 1595 23850 1659
rect 23784 1579 23850 1595
rect 23784 1515 23785 1579
rect 23849 1515 23850 1579
rect 23784 1499 23850 1515
rect 23784 1435 23785 1499
rect 23849 1435 23850 1499
rect 23784 1419 23850 1435
rect 23784 1355 23785 1419
rect 23849 1355 23850 1419
rect 23784 1339 23850 1355
rect 23784 1275 23785 1339
rect 23849 1275 23850 1339
rect 23784 1259 23850 1275
rect 23784 1195 23785 1259
rect 23849 1195 23850 1259
rect 23784 1179 23850 1195
rect 23784 1115 23785 1179
rect 23849 1115 23850 1179
rect 23784 1099 23850 1115
rect 23784 1035 23785 1099
rect 23849 1035 23850 1099
rect 23784 1019 23850 1035
rect 23784 955 23785 1019
rect 23849 955 23850 1019
rect 23784 801 23850 955
rect 23910 801 23970 1833
rect 24030 863 24090 1893
rect 24150 801 24210 1833
rect 24270 863 24330 1893
rect 24390 1739 24456 1829
rect 24390 1675 24391 1739
rect 24455 1675 24456 1739
rect 24390 1659 24456 1675
rect 24390 1595 24391 1659
rect 24455 1595 24456 1659
rect 24390 1579 24456 1595
rect 24390 1515 24391 1579
rect 24455 1515 24456 1579
rect 24390 1499 24456 1515
rect 24390 1435 24391 1499
rect 24455 1435 24456 1499
rect 24390 1419 24456 1435
rect 24390 1355 24391 1419
rect 24455 1355 24456 1419
rect 24390 1339 24456 1355
rect 24390 1275 24391 1339
rect 24455 1275 24456 1339
rect 24390 1259 24456 1275
rect 24390 1195 24391 1259
rect 24455 1195 24456 1259
rect 24390 1179 24456 1195
rect 24390 1115 24391 1179
rect 24455 1115 24456 1179
rect 24390 1099 24456 1115
rect 24390 1035 24391 1099
rect 24455 1035 24456 1099
rect 24390 1019 24456 1035
rect 24390 955 24391 1019
rect 24455 955 24456 1019
rect 24390 801 24456 955
rect 24516 801 24576 1833
rect 24636 863 24696 1893
rect 24756 801 24816 1833
rect 24876 863 24936 1893
rect 24996 1739 25062 1829
rect 24996 1675 24997 1739
rect 25061 1675 25062 1739
rect 24996 1659 25062 1675
rect 24996 1595 24997 1659
rect 25061 1595 25062 1659
rect 24996 1579 25062 1595
rect 24996 1515 24997 1579
rect 25061 1515 25062 1579
rect 24996 1499 25062 1515
rect 24996 1435 24997 1499
rect 25061 1435 25062 1499
rect 24996 1419 25062 1435
rect 24996 1355 24997 1419
rect 25061 1355 25062 1419
rect 24996 1339 25062 1355
rect 24996 1275 24997 1339
rect 25061 1275 25062 1339
rect 24996 1259 25062 1275
rect 24996 1195 24997 1259
rect 25061 1195 25062 1259
rect 24996 1179 25062 1195
rect 24996 1115 24997 1179
rect 25061 1115 25062 1179
rect 24996 1099 25062 1115
rect 24996 1035 24997 1099
rect 25061 1035 25062 1099
rect 24996 1019 25062 1035
rect 24996 955 24997 1019
rect 25061 955 25062 1019
rect 24996 801 25062 955
rect 25122 801 25182 1833
rect 25242 863 25302 1893
rect 25362 801 25422 1833
rect 25482 863 25542 1893
rect 25602 1739 25668 1829
rect 25602 1675 25603 1739
rect 25667 1675 25668 1739
rect 25602 1659 25668 1675
rect 25602 1595 25603 1659
rect 25667 1595 25668 1659
rect 25602 1579 25668 1595
rect 25602 1515 25603 1579
rect 25667 1515 25668 1579
rect 25602 1499 25668 1515
rect 25602 1435 25603 1499
rect 25667 1435 25668 1499
rect 25602 1419 25668 1435
rect 25602 1355 25603 1419
rect 25667 1355 25668 1419
rect 25602 1339 25668 1355
rect 25602 1275 25603 1339
rect 25667 1275 25668 1339
rect 25602 1259 25668 1275
rect 25602 1195 25603 1259
rect 25667 1195 25668 1259
rect 25602 1179 25668 1195
rect 25602 1115 25603 1179
rect 25667 1115 25668 1179
rect 25602 1099 25668 1115
rect 25602 1035 25603 1099
rect 25667 1035 25668 1099
rect 25602 1019 25668 1035
rect 25602 955 25603 1019
rect 25667 955 25668 1019
rect 25602 801 25668 955
rect 25728 801 25788 1833
rect 25848 863 25908 1893
rect 25968 801 26028 1833
rect 26088 863 26148 1893
rect 26208 1739 26274 1829
rect 26208 1675 26209 1739
rect 26273 1675 26274 1739
rect 26208 1659 26274 1675
rect 26208 1595 26209 1659
rect 26273 1595 26274 1659
rect 26208 1579 26274 1595
rect 26208 1515 26209 1579
rect 26273 1515 26274 1579
rect 26208 1499 26274 1515
rect 26208 1435 26209 1499
rect 26273 1435 26274 1499
rect 26208 1419 26274 1435
rect 26208 1355 26209 1419
rect 26273 1355 26274 1419
rect 26208 1339 26274 1355
rect 26208 1275 26209 1339
rect 26273 1275 26274 1339
rect 26208 1259 26274 1275
rect 26208 1195 26209 1259
rect 26273 1195 26274 1259
rect 26208 1179 26274 1195
rect 26208 1115 26209 1179
rect 26273 1115 26274 1179
rect 26208 1099 26274 1115
rect 26208 1035 26209 1099
rect 26273 1035 26274 1099
rect 26208 1019 26274 1035
rect 26208 955 26209 1019
rect 26273 955 26274 1019
rect 26208 801 26274 955
rect 26334 801 26394 1833
rect 26454 863 26514 1893
rect 26574 801 26634 1833
rect 26694 863 26754 1893
rect 26814 1739 26880 1829
rect 26814 1675 26815 1739
rect 26879 1675 26880 1739
rect 26814 1659 26880 1675
rect 26814 1595 26815 1659
rect 26879 1595 26880 1659
rect 26814 1579 26880 1595
rect 26814 1515 26815 1579
rect 26879 1515 26880 1579
rect 26814 1499 26880 1515
rect 26814 1435 26815 1499
rect 26879 1435 26880 1499
rect 26814 1419 26880 1435
rect 26814 1355 26815 1419
rect 26879 1355 26880 1419
rect 26814 1339 26880 1355
rect 26814 1275 26815 1339
rect 26879 1275 26880 1339
rect 26814 1259 26880 1275
rect 26814 1195 26815 1259
rect 26879 1195 26880 1259
rect 26814 1179 26880 1195
rect 26814 1115 26815 1179
rect 26879 1115 26880 1179
rect 26814 1099 26880 1115
rect 26814 1035 26815 1099
rect 26879 1035 26880 1099
rect 26814 1019 26880 1035
rect 26814 955 26815 1019
rect 26879 955 26880 1019
rect 26814 801 26880 955
rect 26940 801 27000 1833
rect 27060 863 27120 1893
rect 27180 801 27240 1833
rect 27300 863 27360 1893
rect 27420 1739 27486 1829
rect 27420 1675 27421 1739
rect 27485 1675 27486 1739
rect 27420 1659 27486 1675
rect 27420 1595 27421 1659
rect 27485 1595 27486 1659
rect 27420 1579 27486 1595
rect 27420 1515 27421 1579
rect 27485 1515 27486 1579
rect 27420 1499 27486 1515
rect 27420 1435 27421 1499
rect 27485 1435 27486 1499
rect 27420 1419 27486 1435
rect 27420 1355 27421 1419
rect 27485 1355 27486 1419
rect 27420 1339 27486 1355
rect 27420 1275 27421 1339
rect 27485 1275 27486 1339
rect 27420 1259 27486 1275
rect 27420 1195 27421 1259
rect 27485 1195 27486 1259
rect 27420 1179 27486 1195
rect 27420 1115 27421 1179
rect 27485 1115 27486 1179
rect 27420 1099 27486 1115
rect 27420 1035 27421 1099
rect 27485 1035 27486 1099
rect 27420 1019 27486 1035
rect 27420 955 27421 1019
rect 27485 955 27486 1019
rect 27420 801 27486 955
rect 27546 801 27606 1833
rect 27666 863 27726 1893
rect 27786 801 27846 1833
rect 27906 863 27966 1893
rect 28026 1739 28092 1829
rect 28026 1675 28027 1739
rect 28091 1675 28092 1739
rect 28026 1659 28092 1675
rect 28026 1595 28027 1659
rect 28091 1595 28092 1659
rect 28026 1579 28092 1595
rect 28026 1515 28027 1579
rect 28091 1515 28092 1579
rect 28026 1499 28092 1515
rect 28026 1435 28027 1499
rect 28091 1435 28092 1499
rect 28026 1419 28092 1435
rect 28026 1355 28027 1419
rect 28091 1355 28092 1419
rect 28026 1339 28092 1355
rect 28026 1275 28027 1339
rect 28091 1275 28092 1339
rect 28026 1259 28092 1275
rect 28026 1195 28027 1259
rect 28091 1195 28092 1259
rect 28026 1179 28092 1195
rect 28026 1115 28027 1179
rect 28091 1115 28092 1179
rect 28026 1099 28092 1115
rect 28026 1035 28027 1099
rect 28091 1035 28092 1099
rect 28026 1019 28092 1035
rect 28026 955 28027 1019
rect 28091 955 28092 1019
rect 28026 801 28092 955
rect 28152 801 28212 1833
rect 28272 863 28332 1893
rect 28392 801 28452 1833
rect 28512 863 28572 1893
rect 28632 1739 28698 1829
rect 28632 1675 28633 1739
rect 28697 1675 28698 1739
rect 28632 1659 28698 1675
rect 28632 1595 28633 1659
rect 28697 1595 28698 1659
rect 28632 1579 28698 1595
rect 28632 1515 28633 1579
rect 28697 1515 28698 1579
rect 28632 1499 28698 1515
rect 28632 1435 28633 1499
rect 28697 1435 28698 1499
rect 28632 1419 28698 1435
rect 28632 1355 28633 1419
rect 28697 1355 28698 1419
rect 28632 1339 28698 1355
rect 28632 1275 28633 1339
rect 28697 1275 28698 1339
rect 28632 1259 28698 1275
rect 28632 1195 28633 1259
rect 28697 1195 28698 1259
rect 28632 1179 28698 1195
rect 28632 1115 28633 1179
rect 28697 1115 28698 1179
rect 28632 1099 28698 1115
rect 28632 1035 28633 1099
rect 28697 1035 28698 1099
rect 28632 1019 28698 1035
rect 28632 955 28633 1019
rect 28697 955 28698 1019
rect 28632 801 28698 955
rect 28758 801 28818 1833
rect 28878 863 28938 1893
rect 28998 801 29058 1833
rect 29118 863 29178 1893
rect 29238 1816 29304 1829
rect 29238 1760 29243 1816
rect 29299 1760 29304 1816
rect 29238 1739 29304 1760
rect 29238 1675 29239 1739
rect 29303 1675 29304 1739
rect 29238 1659 29304 1675
rect 29238 1595 29239 1659
rect 29303 1595 29304 1659
rect 29238 1579 29304 1595
rect 29238 1515 29239 1579
rect 29303 1515 29304 1579
rect 29238 1499 29304 1515
rect 29238 1435 29239 1499
rect 29303 1435 29304 1499
rect 29238 1419 29304 1435
rect 29238 1355 29239 1419
rect 29303 1355 29304 1419
rect 29238 1339 29304 1355
rect 29238 1275 29239 1339
rect 29303 1275 29304 1339
rect 29238 1259 29304 1275
rect 29238 1195 29239 1259
rect 29303 1195 29304 1259
rect 29238 1179 29304 1195
rect 29238 1115 29239 1179
rect 29303 1115 29304 1179
rect 29238 1099 29304 1115
rect 29238 1035 29239 1099
rect 29303 1035 29304 1099
rect 29238 1019 29304 1035
rect 29238 955 29239 1019
rect 29303 955 29304 1019
rect 29238 801 29304 955
rect 29364 801 29424 1833
rect 29484 863 29544 1893
rect 29604 801 29664 1833
rect 29724 863 29784 1893
rect 29844 1816 29910 1829
rect 29844 1760 29849 1816
rect 29905 1760 29910 1816
rect 29844 1739 29910 1760
rect 29844 1675 29845 1739
rect 29909 1675 29910 1739
rect 29844 1659 29910 1675
rect 29844 1595 29845 1659
rect 29909 1595 29910 1659
rect 29844 1579 29910 1595
rect 29844 1515 29845 1579
rect 29909 1515 29910 1579
rect 29844 1499 29910 1515
rect 29844 1435 29845 1499
rect 29909 1435 29910 1499
rect 29844 1419 29910 1435
rect 29844 1355 29845 1419
rect 29909 1355 29910 1419
rect 29844 1339 29910 1355
rect 29844 1275 29845 1339
rect 29909 1275 29910 1339
rect 29844 1259 29910 1275
rect 29844 1195 29845 1259
rect 29909 1195 29910 1259
rect 29844 1179 29910 1195
rect 29844 1115 29845 1179
rect 29909 1115 29910 1179
rect 29844 1099 29910 1115
rect 29844 1035 29845 1099
rect 29909 1035 29910 1099
rect 29844 1019 29910 1035
rect 29844 955 29845 1019
rect 29909 955 29910 1019
rect 29844 801 29910 955
rect 29970 801 30030 1833
rect 30090 863 30150 1893
rect 30210 801 30270 1833
rect 30330 863 30390 1893
rect 30450 1815 30516 1829
rect 30450 1759 30455 1815
rect 30511 1759 30516 1815
rect 30450 1739 30516 1759
rect 30450 1675 30451 1739
rect 30515 1675 30516 1739
rect 30450 1659 30516 1675
rect 30450 1595 30451 1659
rect 30515 1595 30516 1659
rect 30450 1579 30516 1595
rect 30450 1515 30451 1579
rect 30515 1515 30516 1579
rect 30450 1499 30516 1515
rect 30450 1435 30451 1499
rect 30515 1435 30516 1499
rect 30450 1419 30516 1435
rect 30450 1355 30451 1419
rect 30515 1355 30516 1419
rect 30450 1339 30516 1355
rect 30450 1275 30451 1339
rect 30515 1275 30516 1339
rect 30450 1259 30516 1275
rect 30450 1195 30451 1259
rect 30515 1195 30516 1259
rect 30450 1179 30516 1195
rect 30450 1115 30451 1179
rect 30515 1115 30516 1179
rect 30450 1099 30516 1115
rect 30450 1035 30451 1099
rect 30515 1035 30516 1099
rect 30450 1019 30516 1035
rect 30450 955 30451 1019
rect 30515 955 30516 1019
rect 30450 801 30516 955
rect 30576 801 30636 1833
rect 30696 863 30756 1893
rect 30816 801 30876 1833
rect 30936 863 30996 1893
rect 31056 1816 31122 1829
rect 31056 1760 31061 1816
rect 31117 1760 31122 1816
rect 31056 1739 31122 1760
rect 31056 1675 31057 1739
rect 31121 1675 31122 1739
rect 31056 1659 31122 1675
rect 31056 1595 31057 1659
rect 31121 1595 31122 1659
rect 31056 1579 31122 1595
rect 31056 1515 31057 1579
rect 31121 1515 31122 1579
rect 31056 1499 31122 1515
rect 31056 1435 31057 1499
rect 31121 1435 31122 1499
rect 31056 1419 31122 1435
rect 31056 1355 31057 1419
rect 31121 1355 31122 1419
rect 31056 1339 31122 1355
rect 31056 1275 31057 1339
rect 31121 1275 31122 1339
rect 31056 1259 31122 1275
rect 31056 1195 31057 1259
rect 31121 1195 31122 1259
rect 31056 1179 31122 1195
rect 31056 1115 31057 1179
rect 31121 1115 31122 1179
rect 31056 1099 31122 1115
rect 31056 1035 31057 1099
rect 31121 1035 31122 1099
rect 31056 1019 31122 1035
rect 31056 955 31057 1019
rect 31121 955 31122 1019
rect 31056 801 31122 955
rect 31182 801 31242 1833
rect 31302 863 31362 1893
rect 31422 801 31482 1833
rect 31542 863 31602 1893
rect 31662 1816 31728 1829
rect 31662 1760 31667 1816
rect 31723 1760 31728 1816
rect 31662 1739 31728 1760
rect 31662 1675 31663 1739
rect 31727 1675 31728 1739
rect 31662 1659 31728 1675
rect 31662 1595 31663 1659
rect 31727 1595 31728 1659
rect 31662 1579 31728 1595
rect 31662 1515 31663 1579
rect 31727 1515 31728 1579
rect 31662 1499 31728 1515
rect 31662 1435 31663 1499
rect 31727 1435 31728 1499
rect 31662 1419 31728 1435
rect 31662 1355 31663 1419
rect 31727 1355 31728 1419
rect 31662 1339 31728 1355
rect 31662 1275 31663 1339
rect 31727 1275 31728 1339
rect 31662 1259 31728 1275
rect 31662 1195 31663 1259
rect 31727 1195 31728 1259
rect 31662 1179 31728 1195
rect 31662 1115 31663 1179
rect 31727 1115 31728 1179
rect 31662 1099 31728 1115
rect 31662 1035 31663 1099
rect 31727 1035 31728 1099
rect 31662 1019 31728 1035
rect 31662 955 31663 1019
rect 31727 955 31728 1019
rect 31662 801 31728 955
rect 31788 801 31848 1833
rect 31908 863 31968 1893
rect 32028 801 32088 1833
rect 32148 863 32208 1893
rect 32268 1816 32334 1829
rect 32268 1760 32273 1816
rect 32329 1760 32334 1816
rect 32268 1739 32334 1760
rect 32268 1675 32269 1739
rect 32333 1675 32334 1739
rect 32268 1659 32334 1675
rect 32268 1595 32269 1659
rect 32333 1595 32334 1659
rect 32268 1579 32334 1595
rect 32268 1515 32269 1579
rect 32333 1515 32334 1579
rect 32268 1499 32334 1515
rect 32268 1435 32269 1499
rect 32333 1435 32334 1499
rect 32268 1419 32334 1435
rect 32268 1355 32269 1419
rect 32333 1355 32334 1419
rect 32268 1339 32334 1355
rect 32268 1275 32269 1339
rect 32333 1275 32334 1339
rect 32268 1259 32334 1275
rect 32268 1195 32269 1259
rect 32333 1195 32334 1259
rect 32268 1179 32334 1195
rect 32268 1115 32269 1179
rect 32333 1115 32334 1179
rect 32268 1099 32334 1115
rect 32268 1035 32269 1099
rect 32333 1035 32334 1099
rect 32268 1019 32334 1035
rect 32268 955 32269 1019
rect 32333 955 32334 1019
rect 32268 801 32334 955
rect 32394 801 32454 1833
rect 32514 863 32574 1893
rect 32634 801 32694 1833
rect 32754 863 32814 1893
rect 32874 1816 32940 1829
rect 32874 1760 32879 1816
rect 32935 1760 32940 1816
rect 32874 1739 32940 1760
rect 32874 1675 32875 1739
rect 32939 1675 32940 1739
rect 32874 1659 32940 1675
rect 32874 1595 32875 1659
rect 32939 1595 32940 1659
rect 32874 1579 32940 1595
rect 32874 1515 32875 1579
rect 32939 1515 32940 1579
rect 32874 1499 32940 1515
rect 32874 1435 32875 1499
rect 32939 1435 32940 1499
rect 32874 1419 32940 1435
rect 32874 1355 32875 1419
rect 32939 1355 32940 1419
rect 32874 1339 32940 1355
rect 32874 1275 32875 1339
rect 32939 1275 32940 1339
rect 32874 1259 32940 1275
rect 32874 1195 32875 1259
rect 32939 1195 32940 1259
rect 32874 1179 32940 1195
rect 32874 1115 32875 1179
rect 32939 1115 32940 1179
rect 32874 1099 32940 1115
rect 32874 1035 32875 1099
rect 32939 1035 32940 1099
rect 32874 1019 32940 1035
rect 32874 955 32875 1019
rect 32939 955 32940 1019
rect 32874 801 32940 955
rect 33000 801 33060 1833
rect 33120 863 33180 1893
rect 33240 801 33300 1833
rect 33360 863 33420 1893
rect 33480 1816 33546 1829
rect 33480 1760 33485 1816
rect 33541 1760 33546 1816
rect 33480 1739 33546 1760
rect 33480 1675 33481 1739
rect 33545 1675 33546 1739
rect 33480 1659 33546 1675
rect 33480 1595 33481 1659
rect 33545 1595 33546 1659
rect 33480 1579 33546 1595
rect 33480 1515 33481 1579
rect 33545 1515 33546 1579
rect 33480 1499 33546 1515
rect 33480 1435 33481 1499
rect 33545 1435 33546 1499
rect 33480 1419 33546 1435
rect 33480 1355 33481 1419
rect 33545 1355 33546 1419
rect 33480 1339 33546 1355
rect 33480 1275 33481 1339
rect 33545 1275 33546 1339
rect 33480 1259 33546 1275
rect 33480 1195 33481 1259
rect 33545 1195 33546 1259
rect 33480 1179 33546 1195
rect 33480 1115 33481 1179
rect 33545 1115 33546 1179
rect 33480 1099 33546 1115
rect 33480 1035 33481 1099
rect 33545 1035 33546 1099
rect 33480 1019 33546 1035
rect 33480 955 33481 1019
rect 33545 955 33546 1019
rect 33480 801 33546 955
rect 33606 801 33666 1833
rect 33726 863 33786 1893
rect 33846 801 33906 1833
rect 33966 863 34026 1893
rect 34086 1816 34152 1829
rect 34086 1760 34091 1816
rect 34147 1760 34152 1816
rect 34086 1739 34152 1760
rect 34086 1675 34087 1739
rect 34151 1675 34152 1739
rect 34086 1659 34152 1675
rect 34086 1595 34087 1659
rect 34151 1595 34152 1659
rect 34086 1579 34152 1595
rect 34086 1515 34087 1579
rect 34151 1515 34152 1579
rect 34086 1499 34152 1515
rect 34086 1435 34087 1499
rect 34151 1435 34152 1499
rect 34086 1419 34152 1435
rect 34086 1355 34087 1419
rect 34151 1355 34152 1419
rect 34086 1339 34152 1355
rect 34086 1275 34087 1339
rect 34151 1275 34152 1339
rect 34086 1259 34152 1275
rect 34086 1195 34087 1259
rect 34151 1195 34152 1259
rect 34086 1179 34152 1195
rect 34086 1115 34087 1179
rect 34151 1115 34152 1179
rect 34086 1099 34152 1115
rect 34086 1035 34087 1099
rect 34151 1035 34152 1099
rect 34086 1019 34152 1035
rect 34086 955 34087 1019
rect 34151 955 34152 1019
rect 34086 801 34152 955
rect 34212 801 34272 1833
rect 34332 863 34392 1893
rect 34452 801 34512 1833
rect 34572 863 34632 1893
rect 34692 1816 34758 1829
rect 34692 1760 34697 1816
rect 34753 1760 34758 1816
rect 34692 1739 34758 1760
rect 34692 1675 34693 1739
rect 34757 1675 34758 1739
rect 34692 1659 34758 1675
rect 34692 1595 34693 1659
rect 34757 1595 34758 1659
rect 34692 1579 34758 1595
rect 34692 1515 34693 1579
rect 34757 1515 34758 1579
rect 34692 1499 34758 1515
rect 34692 1435 34693 1499
rect 34757 1435 34758 1499
rect 34692 1419 34758 1435
rect 34692 1355 34693 1419
rect 34757 1355 34758 1419
rect 34692 1339 34758 1355
rect 34692 1275 34693 1339
rect 34757 1275 34758 1339
rect 34692 1259 34758 1275
rect 34692 1195 34693 1259
rect 34757 1195 34758 1259
rect 34692 1179 34758 1195
rect 34692 1115 34693 1179
rect 34757 1115 34758 1179
rect 34692 1099 34758 1115
rect 34692 1035 34693 1099
rect 34757 1035 34758 1099
rect 34692 1019 34758 1035
rect 34692 955 34693 1019
rect 34757 955 34758 1019
rect 34692 801 34758 955
rect 34818 801 34878 1833
rect 34938 863 34998 1893
rect 35058 801 35118 1833
rect 35178 863 35238 1893
rect 35298 1816 35364 1829
rect 35298 1760 35303 1816
rect 35359 1760 35364 1816
rect 35298 1739 35364 1760
rect 35298 1675 35299 1739
rect 35363 1675 35364 1739
rect 35298 1659 35364 1675
rect 35298 1595 35299 1659
rect 35363 1595 35364 1659
rect 35298 1579 35364 1595
rect 35298 1515 35299 1579
rect 35363 1515 35364 1579
rect 35298 1499 35364 1515
rect 35298 1435 35299 1499
rect 35363 1435 35364 1499
rect 35298 1419 35364 1435
rect 35298 1355 35299 1419
rect 35363 1355 35364 1419
rect 35298 1339 35364 1355
rect 35298 1275 35299 1339
rect 35363 1275 35364 1339
rect 35298 1259 35364 1275
rect 35298 1195 35299 1259
rect 35363 1195 35364 1259
rect 35298 1179 35364 1195
rect 35298 1115 35299 1179
rect 35363 1115 35364 1179
rect 35298 1099 35364 1115
rect 35298 1035 35299 1099
rect 35363 1035 35364 1099
rect 35298 1019 35364 1035
rect 35298 955 35299 1019
rect 35363 955 35364 1019
rect 35298 801 35364 955
rect 35424 801 35484 1833
rect 35544 863 35604 1893
rect 35664 801 35724 1833
rect 35784 863 35844 1893
rect 35904 1815 35970 1829
rect 35904 1759 35909 1815
rect 35965 1759 35970 1815
rect 35904 1739 35970 1759
rect 35904 1675 35905 1739
rect 35969 1675 35970 1739
rect 35904 1659 35970 1675
rect 35904 1595 35905 1659
rect 35969 1595 35970 1659
rect 35904 1579 35970 1595
rect 35904 1515 35905 1579
rect 35969 1515 35970 1579
rect 35904 1499 35970 1515
rect 35904 1435 35905 1499
rect 35969 1435 35970 1499
rect 35904 1419 35970 1435
rect 35904 1355 35905 1419
rect 35969 1355 35970 1419
rect 35904 1339 35970 1355
rect 35904 1275 35905 1339
rect 35969 1275 35970 1339
rect 35904 1259 35970 1275
rect 35904 1195 35905 1259
rect 35969 1195 35970 1259
rect 35904 1179 35970 1195
rect 35904 1115 35905 1179
rect 35969 1115 35970 1179
rect 35904 1099 35970 1115
rect 35904 1035 35905 1099
rect 35969 1035 35970 1099
rect 35904 1019 35970 1035
rect 35904 955 35905 1019
rect 35969 955 35970 1019
rect 35904 801 35970 955
rect 36030 801 36090 1833
rect 36150 863 36210 1893
rect 36270 801 36330 1833
rect 36390 863 36450 1893
rect 36510 1816 36576 1829
rect 36510 1760 36515 1816
rect 36571 1760 36576 1816
rect 36510 1739 36576 1760
rect 36510 1675 36511 1739
rect 36575 1675 36576 1739
rect 36510 1659 36576 1675
rect 36510 1595 36511 1659
rect 36575 1595 36576 1659
rect 36510 1579 36576 1595
rect 36510 1515 36511 1579
rect 36575 1515 36576 1579
rect 36510 1499 36576 1515
rect 36510 1435 36511 1499
rect 36575 1435 36576 1499
rect 36510 1419 36576 1435
rect 36510 1355 36511 1419
rect 36575 1355 36576 1419
rect 36510 1339 36576 1355
rect 36510 1275 36511 1339
rect 36575 1275 36576 1339
rect 36510 1259 36576 1275
rect 36510 1195 36511 1259
rect 36575 1195 36576 1259
rect 36510 1179 36576 1195
rect 36510 1115 36511 1179
rect 36575 1115 36576 1179
rect 36510 1099 36576 1115
rect 36510 1035 36511 1099
rect 36575 1035 36576 1099
rect 36510 1019 36576 1035
rect 36510 955 36511 1019
rect 36575 955 36576 1019
rect 36510 801 36576 955
rect 36636 801 36696 1833
rect 36756 863 36816 1893
rect 36876 801 36936 1833
rect 36996 863 37056 1893
rect 37116 1816 37182 1829
rect 37116 1760 37121 1816
rect 37177 1760 37182 1816
rect 37116 1739 37182 1760
rect 37116 1675 37117 1739
rect 37181 1675 37182 1739
rect 37116 1659 37182 1675
rect 37116 1595 37117 1659
rect 37181 1595 37182 1659
rect 37116 1579 37182 1595
rect 37116 1515 37117 1579
rect 37181 1515 37182 1579
rect 37116 1499 37182 1515
rect 37116 1435 37117 1499
rect 37181 1435 37182 1499
rect 37116 1419 37182 1435
rect 37116 1355 37117 1419
rect 37181 1355 37182 1419
rect 37116 1339 37182 1355
rect 37116 1275 37117 1339
rect 37181 1275 37182 1339
rect 37116 1259 37182 1275
rect 37116 1195 37117 1259
rect 37181 1195 37182 1259
rect 37116 1179 37182 1195
rect 37116 1115 37117 1179
rect 37181 1115 37182 1179
rect 37116 1099 37182 1115
rect 37116 1035 37117 1099
rect 37181 1035 37182 1099
rect 37116 1019 37182 1035
rect 37116 955 37117 1019
rect 37181 955 37182 1019
rect 37116 801 37182 955
rect 37242 801 37302 1833
rect 37362 863 37422 1893
rect 37482 801 37542 1833
rect 37602 863 37662 1893
rect 37722 1816 37788 1829
rect 37722 1760 37727 1816
rect 37783 1760 37788 1816
rect 37722 1739 37788 1760
rect 37722 1675 37723 1739
rect 37787 1675 37788 1739
rect 37722 1659 37788 1675
rect 37722 1595 37723 1659
rect 37787 1595 37788 1659
rect 37722 1579 37788 1595
rect 37722 1515 37723 1579
rect 37787 1515 37788 1579
rect 37722 1499 37788 1515
rect 37722 1435 37723 1499
rect 37787 1435 37788 1499
rect 37722 1419 37788 1435
rect 37722 1355 37723 1419
rect 37787 1355 37788 1419
rect 37722 1339 37788 1355
rect 37722 1275 37723 1339
rect 37787 1275 37788 1339
rect 37722 1259 37788 1275
rect 37722 1195 37723 1259
rect 37787 1195 37788 1259
rect 37722 1179 37788 1195
rect 37722 1115 37723 1179
rect 37787 1115 37788 1179
rect 37722 1099 37788 1115
rect 37722 1035 37723 1099
rect 37787 1035 37788 1099
rect 37722 1019 37788 1035
rect 37722 955 37723 1019
rect 37787 955 37788 1019
rect 37722 801 37788 955
rect 37848 801 37908 1833
rect 37968 863 38028 1893
rect 38088 801 38148 1833
rect 38208 863 38268 1893
rect 38328 1739 38394 1829
rect 38328 1675 38329 1739
rect 38393 1675 38394 1739
rect 38328 1659 38394 1675
rect 38328 1595 38329 1659
rect 38393 1595 38394 1659
rect 38328 1579 38394 1595
rect 38328 1515 38329 1579
rect 38393 1515 38394 1579
rect 38328 1499 38394 1515
rect 38328 1435 38329 1499
rect 38393 1435 38394 1499
rect 38328 1419 38394 1435
rect 38328 1355 38329 1419
rect 38393 1355 38394 1419
rect 38328 1339 38394 1355
rect 38328 1275 38329 1339
rect 38393 1275 38394 1339
rect 38328 1259 38394 1275
rect 38328 1195 38329 1259
rect 38393 1195 38394 1259
rect 38328 1179 38394 1195
rect 38328 1115 38329 1179
rect 38393 1115 38394 1179
rect 38328 1099 38394 1115
rect 38328 1035 38329 1099
rect 38393 1035 38394 1099
rect 38328 1019 38394 1035
rect 38328 955 38329 1019
rect 38393 955 38394 1019
rect 38328 801 38394 955
rect 38454 801 38514 1833
rect 38574 863 38634 1893
rect 38694 801 38754 1833
rect 38814 863 38874 1893
rect 38934 1739 39000 1829
rect 38934 1675 38935 1739
rect 38999 1675 39000 1739
rect 38934 1659 39000 1675
rect 38934 1595 38935 1659
rect 38999 1595 39000 1659
rect 38934 1579 39000 1595
rect 38934 1515 38935 1579
rect 38999 1515 39000 1579
rect 38934 1499 39000 1515
rect 38934 1435 38935 1499
rect 38999 1435 39000 1499
rect 38934 1419 39000 1435
rect 38934 1355 38935 1419
rect 38999 1355 39000 1419
rect 38934 1339 39000 1355
rect 38934 1275 38935 1339
rect 38999 1275 39000 1339
rect 38934 1259 39000 1275
rect 38934 1195 38935 1259
rect 38999 1195 39000 1259
rect 38934 1179 39000 1195
rect 38934 1115 38935 1179
rect 38999 1115 39000 1179
rect 38934 1099 39000 1115
rect 38934 1035 38935 1099
rect 38999 1035 39000 1099
rect 38934 1019 39000 1035
rect 38934 955 38935 1019
rect 38999 955 39000 1019
rect 38934 801 39000 955
rect 39060 801 39120 1833
rect 39180 863 39240 1893
rect 39300 801 39360 1833
rect 39420 863 39480 1893
rect 39540 1739 39606 1829
rect 39540 1675 39541 1739
rect 39605 1675 39606 1739
rect 39540 1659 39606 1675
rect 39540 1595 39541 1659
rect 39605 1595 39606 1659
rect 39540 1579 39606 1595
rect 39540 1515 39541 1579
rect 39605 1515 39606 1579
rect 39540 1499 39606 1515
rect 39540 1435 39541 1499
rect 39605 1435 39606 1499
rect 39540 1419 39606 1435
rect 39540 1355 39541 1419
rect 39605 1355 39606 1419
rect 39540 1339 39606 1355
rect 39540 1275 39541 1339
rect 39605 1275 39606 1339
rect 39540 1259 39606 1275
rect 39540 1195 39541 1259
rect 39605 1195 39606 1259
rect 39540 1179 39606 1195
rect 39540 1115 39541 1179
rect 39605 1115 39606 1179
rect 39540 1099 39606 1115
rect 39540 1035 39541 1099
rect 39605 1035 39606 1099
rect 39540 1019 39606 1035
rect 39540 955 39541 1019
rect 39605 955 39606 1019
rect 39540 801 39606 955
rect 20148 799 39606 801
rect 20148 735 20252 799
rect 20316 735 20332 799
rect 20396 735 20412 799
rect 20476 735 20492 799
rect 20556 735 20572 799
rect 20636 735 20652 799
rect 20716 735 20858 799
rect 20922 735 20938 799
rect 21002 735 21018 799
rect 21082 735 21098 799
rect 21162 735 21178 799
rect 21242 735 21258 799
rect 21322 735 21464 799
rect 21528 735 21544 799
rect 21608 735 21624 799
rect 21688 735 21704 799
rect 21768 735 21784 799
rect 21848 735 21864 799
rect 21928 735 22070 799
rect 22134 735 22150 799
rect 22214 735 22230 799
rect 22294 735 22310 799
rect 22374 735 22390 799
rect 22454 735 22470 799
rect 22534 735 22676 799
rect 22740 735 22756 799
rect 22820 735 22836 799
rect 22900 735 22916 799
rect 22980 735 22996 799
rect 23060 735 23076 799
rect 23140 735 23282 799
rect 23346 735 23362 799
rect 23426 735 23442 799
rect 23506 735 23522 799
rect 23586 735 23602 799
rect 23666 735 23682 799
rect 23746 735 23888 799
rect 23952 735 23968 799
rect 24032 735 24048 799
rect 24112 735 24128 799
rect 24192 735 24208 799
rect 24272 735 24288 799
rect 24352 735 24494 799
rect 24558 735 24574 799
rect 24638 735 24654 799
rect 24718 735 24734 799
rect 24798 735 24814 799
rect 24878 735 24894 799
rect 24958 735 25100 799
rect 25164 735 25180 799
rect 25244 735 25260 799
rect 25324 735 25340 799
rect 25404 735 25420 799
rect 25484 735 25500 799
rect 25564 735 25706 799
rect 25770 735 25786 799
rect 25850 735 25866 799
rect 25930 735 25946 799
rect 26010 735 26026 799
rect 26090 735 26106 799
rect 26170 735 26312 799
rect 26376 735 26392 799
rect 26456 735 26472 799
rect 26536 735 26552 799
rect 26616 735 26632 799
rect 26696 735 26712 799
rect 26776 735 26918 799
rect 26982 735 26998 799
rect 27062 735 27078 799
rect 27142 735 27158 799
rect 27222 735 27238 799
rect 27302 735 27318 799
rect 27382 735 27524 799
rect 27588 735 27604 799
rect 27668 735 27684 799
rect 27748 735 27764 799
rect 27828 735 27844 799
rect 27908 735 27924 799
rect 27988 735 28130 799
rect 28194 735 28210 799
rect 28274 735 28290 799
rect 28354 735 28370 799
rect 28434 735 28450 799
rect 28514 735 28530 799
rect 28594 735 28736 799
rect 28800 735 28816 799
rect 28880 735 28896 799
rect 28960 735 28976 799
rect 29040 735 29056 799
rect 29120 735 29136 799
rect 29200 735 29342 799
rect 29406 735 29422 799
rect 29486 735 29502 799
rect 29566 735 29582 799
rect 29646 735 29662 799
rect 29726 735 29742 799
rect 29806 735 29948 799
rect 30012 735 30028 799
rect 30092 735 30108 799
rect 30172 735 30188 799
rect 30252 735 30268 799
rect 30332 735 30348 799
rect 30412 735 30554 799
rect 30618 735 30634 799
rect 30698 735 30714 799
rect 30778 735 30794 799
rect 30858 735 30874 799
rect 30938 735 30954 799
rect 31018 735 31160 799
rect 31224 735 31240 799
rect 31304 735 31320 799
rect 31384 735 31400 799
rect 31464 735 31480 799
rect 31544 735 31560 799
rect 31624 735 31766 799
rect 31830 735 31846 799
rect 31910 735 31926 799
rect 31990 735 32006 799
rect 32070 735 32086 799
rect 32150 735 32166 799
rect 32230 735 32372 799
rect 32436 735 32452 799
rect 32516 735 32532 799
rect 32596 735 32612 799
rect 32676 735 32692 799
rect 32756 735 32772 799
rect 32836 735 32978 799
rect 33042 735 33058 799
rect 33122 735 33138 799
rect 33202 735 33218 799
rect 33282 735 33298 799
rect 33362 735 33378 799
rect 33442 735 33584 799
rect 33648 735 33664 799
rect 33728 735 33744 799
rect 33808 735 33824 799
rect 33888 735 33904 799
rect 33968 735 33984 799
rect 34048 735 34190 799
rect 34254 735 34270 799
rect 34334 735 34350 799
rect 34414 735 34430 799
rect 34494 735 34510 799
rect 34574 735 34590 799
rect 34654 735 34796 799
rect 34860 735 34876 799
rect 34940 735 34956 799
rect 35020 735 35036 799
rect 35100 735 35116 799
rect 35180 735 35196 799
rect 35260 735 35402 799
rect 35466 735 35482 799
rect 35546 735 35562 799
rect 35626 735 35642 799
rect 35706 735 35722 799
rect 35786 735 35802 799
rect 35866 735 36008 799
rect 36072 735 36088 799
rect 36152 735 36168 799
rect 36232 735 36248 799
rect 36312 735 36328 799
rect 36392 735 36408 799
rect 36472 735 36614 799
rect 36678 735 36694 799
rect 36758 735 36774 799
rect 36838 735 36854 799
rect 36918 735 36934 799
rect 36998 735 37014 799
rect 37078 735 37220 799
rect 37284 735 37300 799
rect 37364 735 37380 799
rect 37444 735 37460 799
rect 37524 735 37540 799
rect 37604 735 37620 799
rect 37684 735 37826 799
rect 37890 735 37906 799
rect 37970 735 37986 799
rect 38050 735 38066 799
rect 38130 735 38146 799
rect 38210 735 38226 799
rect 38290 735 38432 799
rect 38496 735 38512 799
rect 38576 735 38592 799
rect 38656 735 38672 799
rect 38736 735 38752 799
rect 38816 735 38832 799
rect 38896 735 39038 799
rect 39102 735 39118 799
rect 39182 735 39198 799
rect 39262 735 39278 799
rect 39342 735 39358 799
rect 39422 735 39438 799
rect 39502 735 39606 799
rect 20148 733 39606 735
rect 20148 579 20214 733
rect 20148 515 20149 579
rect 20213 515 20214 579
rect 20148 499 20214 515
rect 20148 435 20149 499
rect 20213 435 20214 499
rect 20148 419 20214 435
rect 20148 355 20149 419
rect 20213 355 20214 419
rect 20148 339 20214 355
rect 20148 275 20149 339
rect 20213 275 20214 339
rect 20148 259 20214 275
rect 20148 195 20149 259
rect 20213 195 20214 259
rect 20148 179 20214 195
rect 20148 115 20149 179
rect 20213 115 20214 179
rect 20148 99 20214 115
rect 20148 35 20149 99
rect 20213 35 20214 99
rect 20148 19 20214 35
rect 20148 -45 20149 19
rect 20213 -45 20214 19
rect 20148 -61 20214 -45
rect 20148 -125 20149 -61
rect 20213 -125 20214 -61
rect 20148 -141 20214 -125
rect 20148 -205 20149 -141
rect 20213 -205 20214 -141
rect 20148 -295 20214 -205
rect 20274 -359 20334 671
rect 20394 -299 20454 733
rect 20514 -359 20574 671
rect 20634 -299 20694 733
rect 20754 579 20820 733
rect 20754 515 20755 579
rect 20819 515 20820 579
rect 20754 499 20820 515
rect 20754 435 20755 499
rect 20819 435 20820 499
rect 20754 419 20820 435
rect 20754 355 20755 419
rect 20819 355 20820 419
rect 20754 339 20820 355
rect 20754 275 20755 339
rect 20819 275 20820 339
rect 20754 259 20820 275
rect 20754 195 20755 259
rect 20819 195 20820 259
rect 20754 179 20820 195
rect 20754 115 20755 179
rect 20819 115 20820 179
rect 20754 99 20820 115
rect 20754 35 20755 99
rect 20819 35 20820 99
rect 20754 19 20820 35
rect 20754 -45 20755 19
rect 20819 -45 20820 19
rect 20754 -61 20820 -45
rect 20754 -125 20755 -61
rect 20819 -125 20820 -61
rect 20754 -141 20820 -125
rect 20754 -205 20755 -141
rect 20819 -205 20820 -141
rect 20754 -295 20820 -205
rect 20880 -359 20940 671
rect 21000 -299 21060 733
rect 21120 -359 21180 671
rect 21240 -299 21300 733
rect 21360 579 21426 733
rect 21360 515 21361 579
rect 21425 515 21426 579
rect 21360 499 21426 515
rect 21360 435 21361 499
rect 21425 435 21426 499
rect 21360 419 21426 435
rect 21360 355 21361 419
rect 21425 355 21426 419
rect 21360 339 21426 355
rect 21360 275 21361 339
rect 21425 275 21426 339
rect 21360 259 21426 275
rect 21360 195 21361 259
rect 21425 195 21426 259
rect 21360 179 21426 195
rect 21360 115 21361 179
rect 21425 115 21426 179
rect 21360 99 21426 115
rect 21360 35 21361 99
rect 21425 35 21426 99
rect 21360 19 21426 35
rect 21360 -45 21361 19
rect 21425 -45 21426 19
rect 21360 -61 21426 -45
rect 21360 -125 21361 -61
rect 21425 -125 21426 -61
rect 21360 -141 21426 -125
rect 21360 -205 21361 -141
rect 21425 -205 21426 -141
rect 21360 -295 21426 -205
rect 21486 -359 21546 671
rect 21606 -299 21666 733
rect 21726 -359 21786 671
rect 21846 -299 21906 733
rect 21966 579 22032 733
rect 21966 515 21967 579
rect 22031 515 22032 579
rect 21966 499 22032 515
rect 21966 435 21967 499
rect 22031 435 22032 499
rect 21966 419 22032 435
rect 21966 355 21967 419
rect 22031 355 22032 419
rect 21966 339 22032 355
rect 21966 275 21967 339
rect 22031 275 22032 339
rect 21966 259 22032 275
rect 21966 195 21967 259
rect 22031 195 22032 259
rect 21966 179 22032 195
rect 21966 115 21967 179
rect 22031 115 22032 179
rect 21966 99 22032 115
rect 21966 35 21967 99
rect 22031 35 22032 99
rect 21966 19 22032 35
rect 21966 -45 21967 19
rect 22031 -45 22032 19
rect 21966 -61 22032 -45
rect 21966 -125 21967 -61
rect 22031 -125 22032 -61
rect 21966 -141 22032 -125
rect 21966 -205 21967 -141
rect 22031 -205 22032 -141
rect 21966 -295 22032 -205
rect 22092 -359 22152 671
rect 22212 -299 22272 733
rect 22332 -359 22392 671
rect 22452 -299 22512 733
rect 22572 579 22638 733
rect 22572 515 22573 579
rect 22637 515 22638 579
rect 22572 499 22638 515
rect 22572 435 22573 499
rect 22637 435 22638 499
rect 22572 419 22638 435
rect 22572 355 22573 419
rect 22637 355 22638 419
rect 22572 339 22638 355
rect 22572 275 22573 339
rect 22637 275 22638 339
rect 22572 259 22638 275
rect 22572 195 22573 259
rect 22637 195 22638 259
rect 22572 179 22638 195
rect 22572 115 22573 179
rect 22637 115 22638 179
rect 22572 99 22638 115
rect 22572 35 22573 99
rect 22637 35 22638 99
rect 22572 19 22638 35
rect 22572 -45 22573 19
rect 22637 -45 22638 19
rect 22572 -61 22638 -45
rect 22572 -125 22573 -61
rect 22637 -125 22638 -61
rect 22572 -141 22638 -125
rect 22572 -205 22573 -141
rect 22637 -205 22638 -141
rect 22572 -295 22638 -205
rect 22698 -359 22758 671
rect 22818 -299 22878 733
rect 22938 -359 22998 671
rect 23058 -299 23118 733
rect 23178 579 23244 733
rect 23178 515 23179 579
rect 23243 515 23244 579
rect 23178 499 23244 515
rect 23178 435 23179 499
rect 23243 435 23244 499
rect 23178 419 23244 435
rect 23178 355 23179 419
rect 23243 355 23244 419
rect 23178 339 23244 355
rect 23178 275 23179 339
rect 23243 275 23244 339
rect 23178 259 23244 275
rect 23178 195 23179 259
rect 23243 195 23244 259
rect 23178 179 23244 195
rect 23178 115 23179 179
rect 23243 115 23244 179
rect 23178 99 23244 115
rect 23178 35 23179 99
rect 23243 35 23244 99
rect 23178 19 23244 35
rect 23178 -45 23179 19
rect 23243 -45 23244 19
rect 23178 -61 23244 -45
rect 23178 -125 23179 -61
rect 23243 -125 23244 -61
rect 23178 -141 23244 -125
rect 23178 -205 23179 -141
rect 23243 -205 23244 -141
rect 23178 -295 23244 -205
rect 23304 -359 23364 671
rect 23424 -299 23484 733
rect 23544 -359 23604 671
rect 23664 -299 23724 733
rect 23784 579 23850 733
rect 23784 515 23785 579
rect 23849 515 23850 579
rect 23784 499 23850 515
rect 23784 435 23785 499
rect 23849 435 23850 499
rect 23784 419 23850 435
rect 23784 355 23785 419
rect 23849 355 23850 419
rect 23784 339 23850 355
rect 23784 275 23785 339
rect 23849 275 23850 339
rect 23784 259 23850 275
rect 23784 195 23785 259
rect 23849 195 23850 259
rect 23784 179 23850 195
rect 23784 115 23785 179
rect 23849 115 23850 179
rect 23784 99 23850 115
rect 23784 35 23785 99
rect 23849 35 23850 99
rect 23784 19 23850 35
rect 23784 -45 23785 19
rect 23849 -45 23850 19
rect 23784 -61 23850 -45
rect 23784 -125 23785 -61
rect 23849 -125 23850 -61
rect 23784 -141 23850 -125
rect 23784 -205 23785 -141
rect 23849 -205 23850 -141
rect 23784 -295 23850 -205
rect 23910 -359 23970 671
rect 24030 -299 24090 733
rect 24150 -359 24210 671
rect 24270 -299 24330 733
rect 24390 579 24456 733
rect 24390 515 24391 579
rect 24455 515 24456 579
rect 24390 499 24456 515
rect 24390 435 24391 499
rect 24455 435 24456 499
rect 24390 419 24456 435
rect 24390 355 24391 419
rect 24455 355 24456 419
rect 24390 339 24456 355
rect 24390 275 24391 339
rect 24455 275 24456 339
rect 24390 259 24456 275
rect 24390 195 24391 259
rect 24455 195 24456 259
rect 24390 179 24456 195
rect 24390 115 24391 179
rect 24455 115 24456 179
rect 24390 99 24456 115
rect 24390 35 24391 99
rect 24455 35 24456 99
rect 24390 19 24456 35
rect 24390 -45 24391 19
rect 24455 -45 24456 19
rect 24390 -61 24456 -45
rect 24390 -125 24391 -61
rect 24455 -125 24456 -61
rect 24390 -141 24456 -125
rect 24390 -205 24391 -141
rect 24455 -205 24456 -141
rect 24390 -295 24456 -205
rect 24516 -359 24576 671
rect 24636 -299 24696 733
rect 24756 -359 24816 671
rect 24876 -299 24936 733
rect 24996 579 25062 733
rect 24996 515 24997 579
rect 25061 515 25062 579
rect 24996 499 25062 515
rect 24996 435 24997 499
rect 25061 435 25062 499
rect 24996 419 25062 435
rect 24996 355 24997 419
rect 25061 355 25062 419
rect 24996 339 25062 355
rect 24996 275 24997 339
rect 25061 275 25062 339
rect 24996 259 25062 275
rect 24996 195 24997 259
rect 25061 195 25062 259
rect 24996 179 25062 195
rect 24996 115 24997 179
rect 25061 115 25062 179
rect 24996 99 25062 115
rect 24996 35 24997 99
rect 25061 35 25062 99
rect 24996 19 25062 35
rect 24996 -45 24997 19
rect 25061 -45 25062 19
rect 24996 -61 25062 -45
rect 24996 -125 24997 -61
rect 25061 -125 25062 -61
rect 24996 -141 25062 -125
rect 24996 -205 24997 -141
rect 25061 -205 25062 -141
rect 24996 -295 25062 -205
rect 25122 -359 25182 671
rect 25242 -299 25302 733
rect 25362 -359 25422 671
rect 25482 -299 25542 733
rect 25602 579 25668 733
rect 25602 515 25603 579
rect 25667 515 25668 579
rect 25602 499 25668 515
rect 25602 435 25603 499
rect 25667 435 25668 499
rect 25602 419 25668 435
rect 25602 355 25603 419
rect 25667 355 25668 419
rect 25602 339 25668 355
rect 25602 275 25603 339
rect 25667 275 25668 339
rect 25602 259 25668 275
rect 25602 195 25603 259
rect 25667 195 25668 259
rect 25602 179 25668 195
rect 25602 115 25603 179
rect 25667 115 25668 179
rect 25602 99 25668 115
rect 25602 35 25603 99
rect 25667 35 25668 99
rect 25602 19 25668 35
rect 25602 -45 25603 19
rect 25667 -45 25668 19
rect 25602 -61 25668 -45
rect 25602 -125 25603 -61
rect 25667 -125 25668 -61
rect 25602 -141 25668 -125
rect 25602 -205 25603 -141
rect 25667 -205 25668 -141
rect 25602 -295 25668 -205
rect 25728 -359 25788 671
rect 25848 -299 25908 733
rect 25968 -359 26028 671
rect 26088 -299 26148 733
rect 26208 579 26274 733
rect 26208 515 26209 579
rect 26273 515 26274 579
rect 26208 499 26274 515
rect 26208 435 26209 499
rect 26273 435 26274 499
rect 26208 419 26274 435
rect 26208 355 26209 419
rect 26273 355 26274 419
rect 26208 339 26274 355
rect 26208 275 26209 339
rect 26273 275 26274 339
rect 26208 259 26274 275
rect 26208 195 26209 259
rect 26273 195 26274 259
rect 26208 179 26274 195
rect 26208 115 26209 179
rect 26273 115 26274 179
rect 26208 99 26274 115
rect 26208 35 26209 99
rect 26273 35 26274 99
rect 26208 19 26274 35
rect 26208 -45 26209 19
rect 26273 -45 26274 19
rect 26208 -61 26274 -45
rect 26208 -125 26209 -61
rect 26273 -125 26274 -61
rect 26208 -141 26274 -125
rect 26208 -205 26209 -141
rect 26273 -205 26274 -141
rect 26208 -295 26274 -205
rect 26334 -359 26394 671
rect 26454 -299 26514 733
rect 26574 -359 26634 671
rect 26694 -299 26754 733
rect 26814 579 26880 733
rect 26814 515 26815 579
rect 26879 515 26880 579
rect 26814 499 26880 515
rect 26814 435 26815 499
rect 26879 435 26880 499
rect 26814 419 26880 435
rect 26814 355 26815 419
rect 26879 355 26880 419
rect 26814 339 26880 355
rect 26814 275 26815 339
rect 26879 275 26880 339
rect 26814 259 26880 275
rect 26814 195 26815 259
rect 26879 195 26880 259
rect 26814 179 26880 195
rect 26814 115 26815 179
rect 26879 115 26880 179
rect 26814 99 26880 115
rect 26814 35 26815 99
rect 26879 35 26880 99
rect 26814 19 26880 35
rect 26814 -45 26815 19
rect 26879 -45 26880 19
rect 26814 -61 26880 -45
rect 26814 -125 26815 -61
rect 26879 -125 26880 -61
rect 26814 -141 26880 -125
rect 26814 -205 26815 -141
rect 26879 -205 26880 -141
rect 26814 -295 26880 -205
rect 26940 -359 27000 671
rect 27060 -299 27120 733
rect 27180 -359 27240 671
rect 27300 -299 27360 733
rect 27420 579 27486 733
rect 27420 515 27421 579
rect 27485 515 27486 579
rect 27420 499 27486 515
rect 27420 435 27421 499
rect 27485 435 27486 499
rect 27420 419 27486 435
rect 27420 355 27421 419
rect 27485 355 27486 419
rect 27420 339 27486 355
rect 27420 275 27421 339
rect 27485 275 27486 339
rect 27420 259 27486 275
rect 27420 195 27421 259
rect 27485 195 27486 259
rect 27420 179 27486 195
rect 27420 115 27421 179
rect 27485 115 27486 179
rect 27420 99 27486 115
rect 27420 35 27421 99
rect 27485 35 27486 99
rect 27420 19 27486 35
rect 27420 -45 27421 19
rect 27485 -45 27486 19
rect 27420 -61 27486 -45
rect 27420 -125 27421 -61
rect 27485 -125 27486 -61
rect 27420 -141 27486 -125
rect 27420 -205 27421 -141
rect 27485 -205 27486 -141
rect 27420 -295 27486 -205
rect 27546 -359 27606 671
rect 27666 -299 27726 733
rect 27786 -359 27846 671
rect 27906 -299 27966 733
rect 28026 579 28092 733
rect 28026 515 28027 579
rect 28091 515 28092 579
rect 28026 499 28092 515
rect 28026 435 28027 499
rect 28091 435 28092 499
rect 28026 419 28092 435
rect 28026 355 28027 419
rect 28091 355 28092 419
rect 28026 339 28092 355
rect 28026 275 28027 339
rect 28091 275 28092 339
rect 28026 259 28092 275
rect 28026 195 28027 259
rect 28091 195 28092 259
rect 28026 179 28092 195
rect 28026 115 28027 179
rect 28091 115 28092 179
rect 28026 99 28092 115
rect 28026 35 28027 99
rect 28091 35 28092 99
rect 28026 19 28092 35
rect 28026 -45 28027 19
rect 28091 -45 28092 19
rect 28026 -61 28092 -45
rect 28026 -125 28027 -61
rect 28091 -125 28092 -61
rect 28026 -141 28092 -125
rect 28026 -205 28027 -141
rect 28091 -205 28092 -141
rect 28026 -295 28092 -205
rect 28152 -359 28212 671
rect 28272 -299 28332 733
rect 28392 -359 28452 671
rect 28512 -299 28572 733
rect 28632 579 28698 733
rect 28632 515 28633 579
rect 28697 515 28698 579
rect 28632 499 28698 515
rect 28632 435 28633 499
rect 28697 435 28698 499
rect 28632 419 28698 435
rect 28632 355 28633 419
rect 28697 355 28698 419
rect 28632 339 28698 355
rect 28632 275 28633 339
rect 28697 275 28698 339
rect 28632 259 28698 275
rect 28632 195 28633 259
rect 28697 195 28698 259
rect 28632 179 28698 195
rect 28632 115 28633 179
rect 28697 115 28698 179
rect 28632 99 28698 115
rect 28632 35 28633 99
rect 28697 35 28698 99
rect 28632 19 28698 35
rect 28632 -45 28633 19
rect 28697 -45 28698 19
rect 28632 -61 28698 -45
rect 28632 -125 28633 -61
rect 28697 -125 28698 -61
rect 28632 -141 28698 -125
rect 28632 -205 28633 -141
rect 28697 -205 28698 -141
rect 28632 -295 28698 -205
rect 28758 -359 28818 671
rect 28878 -299 28938 733
rect 28998 -359 29058 671
rect 29118 -299 29178 733
rect 29238 579 29304 733
rect 29238 515 29239 579
rect 29303 515 29304 579
rect 29238 499 29304 515
rect 29238 435 29239 499
rect 29303 435 29304 499
rect 29238 419 29304 435
rect 29238 355 29239 419
rect 29303 355 29304 419
rect 29238 339 29304 355
rect 29238 275 29239 339
rect 29303 275 29304 339
rect 29238 259 29304 275
rect 29238 195 29239 259
rect 29303 195 29304 259
rect 29238 179 29304 195
rect 29238 115 29239 179
rect 29303 115 29304 179
rect 29238 99 29304 115
rect 29238 35 29239 99
rect 29303 35 29304 99
rect 29238 19 29304 35
rect 29238 -45 29239 19
rect 29303 -45 29304 19
rect 29238 -61 29304 -45
rect 29238 -125 29239 -61
rect 29303 -125 29304 -61
rect 29238 -141 29304 -125
rect 29238 -205 29239 -141
rect 29303 -205 29304 -141
rect 29238 -295 29304 -205
rect 29364 -359 29424 671
rect 29484 -299 29544 733
rect 29604 -359 29664 671
rect 29724 -299 29784 733
rect 29844 579 29910 733
rect 29844 515 29845 579
rect 29909 515 29910 579
rect 29844 499 29910 515
rect 29844 435 29845 499
rect 29909 435 29910 499
rect 29844 419 29910 435
rect 29844 355 29845 419
rect 29909 355 29910 419
rect 29844 339 29910 355
rect 29844 275 29845 339
rect 29909 275 29910 339
rect 29844 259 29910 275
rect 29844 195 29845 259
rect 29909 195 29910 259
rect 29844 179 29910 195
rect 29844 115 29845 179
rect 29909 115 29910 179
rect 29844 99 29910 115
rect 29844 35 29845 99
rect 29909 35 29910 99
rect 29844 19 29910 35
rect 29844 -45 29845 19
rect 29909 -45 29910 19
rect 29844 -61 29910 -45
rect 29844 -125 29845 -61
rect 29909 -125 29910 -61
rect 29844 -141 29910 -125
rect 29844 -205 29845 -141
rect 29909 -205 29910 -141
rect 29844 -295 29910 -205
rect 29970 -359 30030 671
rect 30090 -299 30150 733
rect 30210 -359 30270 671
rect 30330 -299 30390 733
rect 30450 579 30516 733
rect 30450 515 30451 579
rect 30515 515 30516 579
rect 30450 499 30516 515
rect 30450 435 30451 499
rect 30515 435 30516 499
rect 30450 419 30516 435
rect 30450 355 30451 419
rect 30515 355 30516 419
rect 30450 339 30516 355
rect 30450 275 30451 339
rect 30515 275 30516 339
rect 30450 259 30516 275
rect 30450 195 30451 259
rect 30515 195 30516 259
rect 30450 179 30516 195
rect 30450 115 30451 179
rect 30515 115 30516 179
rect 30450 99 30516 115
rect 30450 35 30451 99
rect 30515 35 30516 99
rect 30450 19 30516 35
rect 30450 -45 30451 19
rect 30515 -45 30516 19
rect 30450 -61 30516 -45
rect 30450 -125 30451 -61
rect 30515 -125 30516 -61
rect 30450 -141 30516 -125
rect 30450 -205 30451 -141
rect 30515 -205 30516 -141
rect 30450 -295 30516 -205
rect 30576 -359 30636 671
rect 30696 -299 30756 733
rect 30816 -359 30876 671
rect 30936 -299 30996 733
rect 31056 579 31122 733
rect 31056 515 31057 579
rect 31121 515 31122 579
rect 31056 499 31122 515
rect 31056 435 31057 499
rect 31121 435 31122 499
rect 31056 419 31122 435
rect 31056 355 31057 419
rect 31121 355 31122 419
rect 31056 339 31122 355
rect 31056 275 31057 339
rect 31121 275 31122 339
rect 31056 259 31122 275
rect 31056 195 31057 259
rect 31121 195 31122 259
rect 31056 179 31122 195
rect 31056 115 31057 179
rect 31121 115 31122 179
rect 31056 99 31122 115
rect 31056 35 31057 99
rect 31121 35 31122 99
rect 31056 19 31122 35
rect 31056 -45 31057 19
rect 31121 -45 31122 19
rect 31056 -61 31122 -45
rect 31056 -125 31057 -61
rect 31121 -125 31122 -61
rect 31056 -141 31122 -125
rect 31056 -205 31057 -141
rect 31121 -205 31122 -141
rect 31056 -295 31122 -205
rect 31182 -359 31242 671
rect 31302 -299 31362 733
rect 31422 -359 31482 671
rect 31542 -299 31602 733
rect 31662 579 31728 733
rect 31662 515 31663 579
rect 31727 515 31728 579
rect 31662 499 31728 515
rect 31662 435 31663 499
rect 31727 435 31728 499
rect 31662 419 31728 435
rect 31662 355 31663 419
rect 31727 355 31728 419
rect 31662 339 31728 355
rect 31662 275 31663 339
rect 31727 275 31728 339
rect 31662 259 31728 275
rect 31662 195 31663 259
rect 31727 195 31728 259
rect 31662 179 31728 195
rect 31662 115 31663 179
rect 31727 115 31728 179
rect 31662 99 31728 115
rect 31662 35 31663 99
rect 31727 35 31728 99
rect 31662 19 31728 35
rect 31662 -45 31663 19
rect 31727 -45 31728 19
rect 31662 -61 31728 -45
rect 31662 -125 31663 -61
rect 31727 -125 31728 -61
rect 31662 -141 31728 -125
rect 31662 -205 31663 -141
rect 31727 -205 31728 -141
rect 31662 -295 31728 -205
rect 31788 -359 31848 671
rect 31908 -299 31968 733
rect 32028 -359 32088 671
rect 32148 -299 32208 733
rect 32268 579 32334 733
rect 32268 515 32269 579
rect 32333 515 32334 579
rect 32268 499 32334 515
rect 32268 435 32269 499
rect 32333 435 32334 499
rect 32268 419 32334 435
rect 32268 355 32269 419
rect 32333 355 32334 419
rect 32268 339 32334 355
rect 32268 275 32269 339
rect 32333 275 32334 339
rect 32268 259 32334 275
rect 32268 195 32269 259
rect 32333 195 32334 259
rect 32268 179 32334 195
rect 32268 115 32269 179
rect 32333 115 32334 179
rect 32268 99 32334 115
rect 32268 35 32269 99
rect 32333 35 32334 99
rect 32268 19 32334 35
rect 32268 -45 32269 19
rect 32333 -45 32334 19
rect 32268 -61 32334 -45
rect 32268 -125 32269 -61
rect 32333 -125 32334 -61
rect 32268 -141 32334 -125
rect 32268 -205 32269 -141
rect 32333 -205 32334 -141
rect 32268 -295 32334 -205
rect 32394 -359 32454 671
rect 32514 -299 32574 733
rect 32634 -359 32694 671
rect 32754 -299 32814 733
rect 32874 579 32940 733
rect 32874 515 32875 579
rect 32939 515 32940 579
rect 32874 499 32940 515
rect 32874 435 32875 499
rect 32939 435 32940 499
rect 32874 419 32940 435
rect 32874 355 32875 419
rect 32939 355 32940 419
rect 32874 339 32940 355
rect 32874 275 32875 339
rect 32939 275 32940 339
rect 32874 259 32940 275
rect 32874 195 32875 259
rect 32939 195 32940 259
rect 32874 179 32940 195
rect 32874 115 32875 179
rect 32939 115 32940 179
rect 32874 99 32940 115
rect 32874 35 32875 99
rect 32939 35 32940 99
rect 32874 19 32940 35
rect 32874 -45 32875 19
rect 32939 -45 32940 19
rect 32874 -61 32940 -45
rect 32874 -125 32875 -61
rect 32939 -125 32940 -61
rect 32874 -141 32940 -125
rect 32874 -205 32875 -141
rect 32939 -205 32940 -141
rect 32874 -295 32940 -205
rect 33000 -359 33060 671
rect 33120 -299 33180 733
rect 33240 -359 33300 671
rect 33360 -299 33420 733
rect 33480 579 33546 733
rect 33480 515 33481 579
rect 33545 515 33546 579
rect 33480 499 33546 515
rect 33480 435 33481 499
rect 33545 435 33546 499
rect 33480 419 33546 435
rect 33480 355 33481 419
rect 33545 355 33546 419
rect 33480 339 33546 355
rect 33480 275 33481 339
rect 33545 275 33546 339
rect 33480 259 33546 275
rect 33480 195 33481 259
rect 33545 195 33546 259
rect 33480 179 33546 195
rect 33480 115 33481 179
rect 33545 115 33546 179
rect 33480 99 33546 115
rect 33480 35 33481 99
rect 33545 35 33546 99
rect 33480 19 33546 35
rect 33480 -45 33481 19
rect 33545 -45 33546 19
rect 33480 -61 33546 -45
rect 33480 -125 33481 -61
rect 33545 -125 33546 -61
rect 33480 -141 33546 -125
rect 33480 -205 33481 -141
rect 33545 -205 33546 -141
rect 33480 -295 33546 -205
rect 33606 -359 33666 671
rect 33726 -299 33786 733
rect 33846 -359 33906 671
rect 33966 -299 34026 733
rect 34086 579 34152 733
rect 34086 515 34087 579
rect 34151 515 34152 579
rect 34086 499 34152 515
rect 34086 435 34087 499
rect 34151 435 34152 499
rect 34086 419 34152 435
rect 34086 355 34087 419
rect 34151 355 34152 419
rect 34086 339 34152 355
rect 34086 275 34087 339
rect 34151 275 34152 339
rect 34086 259 34152 275
rect 34086 195 34087 259
rect 34151 195 34152 259
rect 34086 179 34152 195
rect 34086 115 34087 179
rect 34151 115 34152 179
rect 34086 99 34152 115
rect 34086 35 34087 99
rect 34151 35 34152 99
rect 34086 19 34152 35
rect 34086 -45 34087 19
rect 34151 -45 34152 19
rect 34086 -61 34152 -45
rect 34086 -125 34087 -61
rect 34151 -125 34152 -61
rect 34086 -141 34152 -125
rect 34086 -205 34087 -141
rect 34151 -205 34152 -141
rect 34086 -295 34152 -205
rect 34212 -359 34272 671
rect 34332 -299 34392 733
rect 34452 -359 34512 671
rect 34572 -299 34632 733
rect 34692 579 34758 733
rect 34692 515 34693 579
rect 34757 515 34758 579
rect 34692 499 34758 515
rect 34692 435 34693 499
rect 34757 435 34758 499
rect 34692 419 34758 435
rect 34692 355 34693 419
rect 34757 355 34758 419
rect 34692 339 34758 355
rect 34692 275 34693 339
rect 34757 275 34758 339
rect 34692 259 34758 275
rect 34692 195 34693 259
rect 34757 195 34758 259
rect 34692 179 34758 195
rect 34692 115 34693 179
rect 34757 115 34758 179
rect 34692 99 34758 115
rect 34692 35 34693 99
rect 34757 35 34758 99
rect 34692 19 34758 35
rect 34692 -45 34693 19
rect 34757 -45 34758 19
rect 34692 -61 34758 -45
rect 34692 -125 34693 -61
rect 34757 -125 34758 -61
rect 34692 -141 34758 -125
rect 34692 -205 34693 -141
rect 34757 -205 34758 -141
rect 34692 -295 34758 -205
rect 34818 -359 34878 671
rect 34938 -299 34998 733
rect 35058 -359 35118 671
rect 35178 -299 35238 733
rect 35298 579 35364 733
rect 35298 515 35299 579
rect 35363 515 35364 579
rect 35298 499 35364 515
rect 35298 435 35299 499
rect 35363 435 35364 499
rect 35298 419 35364 435
rect 35298 355 35299 419
rect 35363 355 35364 419
rect 35298 339 35364 355
rect 35298 275 35299 339
rect 35363 275 35364 339
rect 35298 259 35364 275
rect 35298 195 35299 259
rect 35363 195 35364 259
rect 35298 179 35364 195
rect 35298 115 35299 179
rect 35363 115 35364 179
rect 35298 99 35364 115
rect 35298 35 35299 99
rect 35363 35 35364 99
rect 35298 19 35364 35
rect 35298 -45 35299 19
rect 35363 -45 35364 19
rect 35298 -61 35364 -45
rect 35298 -125 35299 -61
rect 35363 -125 35364 -61
rect 35298 -141 35364 -125
rect 35298 -205 35299 -141
rect 35363 -205 35364 -141
rect 35298 -295 35364 -205
rect 35424 -359 35484 671
rect 35544 -299 35604 733
rect 35664 -359 35724 671
rect 35784 -299 35844 733
rect 35904 579 35970 733
rect 35904 515 35905 579
rect 35969 515 35970 579
rect 35904 499 35970 515
rect 35904 435 35905 499
rect 35969 435 35970 499
rect 35904 419 35970 435
rect 35904 355 35905 419
rect 35969 355 35970 419
rect 35904 339 35970 355
rect 35904 275 35905 339
rect 35969 275 35970 339
rect 35904 259 35970 275
rect 35904 195 35905 259
rect 35969 195 35970 259
rect 35904 179 35970 195
rect 35904 115 35905 179
rect 35969 115 35970 179
rect 35904 99 35970 115
rect 35904 35 35905 99
rect 35969 35 35970 99
rect 35904 19 35970 35
rect 35904 -45 35905 19
rect 35969 -45 35970 19
rect 35904 -61 35970 -45
rect 35904 -125 35905 -61
rect 35969 -125 35970 -61
rect 35904 -141 35970 -125
rect 35904 -205 35905 -141
rect 35969 -205 35970 -141
rect 35904 -295 35970 -205
rect 36030 -359 36090 671
rect 36150 -299 36210 733
rect 36270 -359 36330 671
rect 36390 -299 36450 733
rect 36510 579 36576 733
rect 36510 515 36511 579
rect 36575 515 36576 579
rect 36510 499 36576 515
rect 36510 435 36511 499
rect 36575 435 36576 499
rect 36510 419 36576 435
rect 36510 355 36511 419
rect 36575 355 36576 419
rect 36510 339 36576 355
rect 36510 275 36511 339
rect 36575 275 36576 339
rect 36510 259 36576 275
rect 36510 195 36511 259
rect 36575 195 36576 259
rect 36510 179 36576 195
rect 36510 115 36511 179
rect 36575 115 36576 179
rect 36510 99 36576 115
rect 36510 35 36511 99
rect 36575 35 36576 99
rect 36510 19 36576 35
rect 36510 -45 36511 19
rect 36575 -45 36576 19
rect 36510 -61 36576 -45
rect 36510 -125 36511 -61
rect 36575 -125 36576 -61
rect 36510 -141 36576 -125
rect 36510 -205 36511 -141
rect 36575 -205 36576 -141
rect 36510 -295 36576 -205
rect 36636 -359 36696 671
rect 36756 -299 36816 733
rect 36876 -359 36936 671
rect 36996 -299 37056 733
rect 37116 579 37182 733
rect 37116 515 37117 579
rect 37181 515 37182 579
rect 37116 499 37182 515
rect 37116 435 37117 499
rect 37181 435 37182 499
rect 37116 419 37182 435
rect 37116 355 37117 419
rect 37181 355 37182 419
rect 37116 339 37182 355
rect 37116 275 37117 339
rect 37181 275 37182 339
rect 37116 259 37182 275
rect 37116 195 37117 259
rect 37181 195 37182 259
rect 37116 179 37182 195
rect 37116 115 37117 179
rect 37181 115 37182 179
rect 37116 99 37182 115
rect 37116 35 37117 99
rect 37181 35 37182 99
rect 37116 19 37182 35
rect 37116 -45 37117 19
rect 37181 -45 37182 19
rect 37116 -61 37182 -45
rect 37116 -125 37117 -61
rect 37181 -125 37182 -61
rect 37116 -141 37182 -125
rect 37116 -205 37117 -141
rect 37181 -205 37182 -141
rect 37116 -295 37182 -205
rect 37242 -359 37302 671
rect 37362 -299 37422 733
rect 37482 -359 37542 671
rect 37602 -299 37662 733
rect 37722 579 37788 733
rect 37722 515 37723 579
rect 37787 515 37788 579
rect 37722 499 37788 515
rect 37722 435 37723 499
rect 37787 435 37788 499
rect 37722 419 37788 435
rect 37722 355 37723 419
rect 37787 355 37788 419
rect 37722 339 37788 355
rect 37722 275 37723 339
rect 37787 275 37788 339
rect 37722 259 37788 275
rect 37722 195 37723 259
rect 37787 195 37788 259
rect 37722 179 37788 195
rect 37722 115 37723 179
rect 37787 115 37788 179
rect 37722 99 37788 115
rect 37722 35 37723 99
rect 37787 35 37788 99
rect 37722 19 37788 35
rect 37722 -45 37723 19
rect 37787 -45 37788 19
rect 37722 -61 37788 -45
rect 37722 -125 37723 -61
rect 37787 -125 37788 -61
rect 37722 -141 37788 -125
rect 37722 -205 37723 -141
rect 37787 -205 37788 -141
rect 37722 -295 37788 -205
rect 37848 -359 37908 671
rect 37968 -299 38028 733
rect 38088 -359 38148 671
rect 38208 -299 38268 733
rect 38328 579 38394 733
rect 38328 515 38329 579
rect 38393 515 38394 579
rect 38328 499 38394 515
rect 38328 435 38329 499
rect 38393 435 38394 499
rect 38328 419 38394 435
rect 38328 355 38329 419
rect 38393 355 38394 419
rect 38328 339 38394 355
rect 38328 275 38329 339
rect 38393 275 38394 339
rect 38328 259 38394 275
rect 38328 195 38329 259
rect 38393 195 38394 259
rect 38328 179 38394 195
rect 38328 115 38329 179
rect 38393 115 38394 179
rect 38328 99 38394 115
rect 38328 35 38329 99
rect 38393 35 38394 99
rect 38328 19 38394 35
rect 38328 -45 38329 19
rect 38393 -45 38394 19
rect 38328 -61 38394 -45
rect 38328 -125 38329 -61
rect 38393 -125 38394 -61
rect 38328 -141 38394 -125
rect 38328 -205 38329 -141
rect 38393 -205 38394 -141
rect 38328 -295 38394 -205
rect 38454 -359 38514 671
rect 38574 -299 38634 733
rect 38694 -359 38754 671
rect 38814 -299 38874 733
rect 38934 579 39000 733
rect 38934 515 38935 579
rect 38999 515 39000 579
rect 38934 499 39000 515
rect 38934 435 38935 499
rect 38999 435 39000 499
rect 38934 419 39000 435
rect 38934 355 38935 419
rect 38999 355 39000 419
rect 38934 339 39000 355
rect 38934 275 38935 339
rect 38999 275 39000 339
rect 38934 259 39000 275
rect 38934 195 38935 259
rect 38999 195 39000 259
rect 38934 179 39000 195
rect 38934 115 38935 179
rect 38999 115 39000 179
rect 38934 99 39000 115
rect 38934 35 38935 99
rect 38999 35 39000 99
rect 38934 19 39000 35
rect 38934 -45 38935 19
rect 38999 -45 39000 19
rect 38934 -61 39000 -45
rect 38934 -125 38935 -61
rect 38999 -125 39000 -61
rect 38934 -141 39000 -125
rect 38934 -205 38935 -141
rect 38999 -205 39000 -141
rect 38934 -295 39000 -205
rect 39060 -359 39120 671
rect 39180 -299 39240 733
rect 39300 -359 39360 671
rect 39420 -299 39480 733
rect 39540 579 39606 733
rect 39540 515 39541 579
rect 39605 515 39606 579
rect 39540 499 39606 515
rect 39540 435 39541 499
rect 39605 435 39606 499
rect 39540 419 39606 435
rect 39540 355 39541 419
rect 39605 355 39606 419
rect 39540 339 39606 355
rect 39540 275 39541 339
rect 39605 275 39606 339
rect 39540 259 39606 275
rect 39540 195 39541 259
rect 39605 195 39606 259
rect 39540 179 39606 195
rect 39540 115 39541 179
rect 39605 115 39606 179
rect 39540 99 39606 115
rect 39540 35 39541 99
rect 39605 35 39606 99
rect 39540 19 39606 35
rect 39540 -45 39541 19
rect 39605 -45 39606 19
rect 39540 -61 39606 -45
rect 39540 -125 39541 -61
rect 39605 -125 39606 -61
rect 39540 -141 39606 -125
rect 39540 -205 39541 -141
rect 39605 -205 39606 -141
rect 39540 -295 39606 -205
rect -459 -361 213 -359
rect -459 -425 -355 -361
rect -291 -425 -275 -361
rect -211 -425 -195 -361
rect -131 -425 -115 -361
rect -51 -425 -35 -361
rect 29 -425 45 -361
rect 109 -425 213 -361
rect -459 -427 213 -425
rect 355 -361 1027 -359
rect 355 -425 459 -361
rect 523 -425 539 -361
rect 603 -425 619 -361
rect 683 -425 699 -361
rect 763 -425 779 -361
rect 843 -425 859 -361
rect 923 -425 1027 -361
rect 355 -427 1027 -425
rect 1267 -361 2545 -359
rect 1267 -425 1371 -361
rect 1435 -425 1451 -361
rect 1515 -425 1531 -361
rect 1595 -425 1611 -361
rect 1675 -425 1691 -361
rect 1755 -425 1771 -361
rect 1835 -425 1977 -361
rect 2041 -425 2057 -361
rect 2121 -425 2137 -361
rect 2201 -425 2217 -361
rect 2281 -425 2297 -361
rect 2361 -425 2377 -361
rect 2441 -425 2545 -361
rect 1267 -427 2545 -425
rect 2801 -361 5291 -359
rect 2801 -425 2905 -361
rect 2969 -425 2985 -361
rect 3049 -425 3065 -361
rect 3129 -425 3145 -361
rect 3209 -425 3225 -361
rect 3289 -425 3305 -361
rect 3369 -425 3511 -361
rect 3575 -425 3591 -361
rect 3655 -425 3671 -361
rect 3735 -425 3751 -361
rect 3815 -425 3831 -361
rect 3895 -425 3911 -361
rect 3975 -425 4117 -361
rect 4181 -425 4197 -361
rect 4261 -425 4277 -361
rect 4341 -425 4357 -361
rect 4421 -425 4437 -361
rect 4501 -425 4517 -361
rect 4581 -425 4723 -361
rect 4787 -425 4803 -361
rect 4867 -425 4883 -361
rect 4947 -425 4963 -361
rect 5027 -425 5043 -361
rect 5107 -425 5123 -361
rect 5187 -425 5291 -361
rect 2801 -427 5291 -425
rect 5352 -361 10266 -359
rect 5352 -425 5456 -361
rect 5520 -425 5536 -361
rect 5600 -425 5616 -361
rect 5680 -425 5696 -361
rect 5760 -425 5776 -361
rect 5840 -425 5856 -361
rect 5920 -425 6062 -361
rect 6126 -425 6142 -361
rect 6206 -425 6222 -361
rect 6286 -425 6302 -361
rect 6366 -425 6382 -361
rect 6446 -425 6462 -361
rect 6526 -425 6668 -361
rect 6732 -425 6748 -361
rect 6812 -425 6828 -361
rect 6892 -425 6908 -361
rect 6972 -425 6988 -361
rect 7052 -425 7068 -361
rect 7132 -425 7274 -361
rect 7338 -425 7354 -361
rect 7418 -425 7434 -361
rect 7498 -425 7514 -361
rect 7578 -425 7594 -361
rect 7658 -425 7674 -361
rect 7738 -425 7880 -361
rect 7944 -425 7960 -361
rect 8024 -425 8040 -361
rect 8104 -425 8120 -361
rect 8184 -425 8200 -361
rect 8264 -425 8280 -361
rect 8344 -425 8486 -361
rect 8550 -425 8566 -361
rect 8630 -425 8646 -361
rect 8710 -425 8726 -361
rect 8790 -425 8806 -361
rect 8870 -425 8886 -361
rect 8950 -425 9092 -361
rect 9156 -425 9172 -361
rect 9236 -425 9252 -361
rect 9316 -425 9332 -361
rect 9396 -425 9412 -361
rect 9476 -425 9492 -361
rect 9556 -425 9698 -361
rect 9762 -425 9778 -361
rect 9842 -425 9858 -361
rect 9922 -425 9938 -361
rect 10002 -425 10018 -361
rect 10082 -425 10098 -361
rect 10162 -425 10266 -361
rect 5352 -427 10266 -425
rect 10326 -361 20088 -359
rect 10326 -425 10430 -361
rect 10494 -425 10510 -361
rect 10574 -425 10590 -361
rect 10654 -425 10670 -361
rect 10734 -425 10750 -361
rect 10814 -425 10830 -361
rect 10894 -425 11036 -361
rect 11100 -425 11116 -361
rect 11180 -425 11196 -361
rect 11260 -425 11276 -361
rect 11340 -425 11356 -361
rect 11420 -425 11436 -361
rect 11500 -425 11642 -361
rect 11706 -425 11722 -361
rect 11786 -425 11802 -361
rect 11866 -425 11882 -361
rect 11946 -425 11962 -361
rect 12026 -425 12042 -361
rect 12106 -425 12248 -361
rect 12312 -425 12328 -361
rect 12392 -425 12408 -361
rect 12472 -425 12488 -361
rect 12552 -425 12568 -361
rect 12632 -425 12648 -361
rect 12712 -425 12854 -361
rect 12918 -425 12934 -361
rect 12998 -425 13014 -361
rect 13078 -425 13094 -361
rect 13158 -425 13174 -361
rect 13238 -425 13254 -361
rect 13318 -425 13460 -361
rect 13524 -425 13540 -361
rect 13604 -425 13620 -361
rect 13684 -425 13700 -361
rect 13764 -425 13780 -361
rect 13844 -425 13860 -361
rect 13924 -425 14066 -361
rect 14130 -425 14146 -361
rect 14210 -425 14226 -361
rect 14290 -425 14306 -361
rect 14370 -425 14386 -361
rect 14450 -425 14466 -361
rect 14530 -425 14672 -361
rect 14736 -425 14752 -361
rect 14816 -425 14832 -361
rect 14896 -425 14912 -361
rect 14976 -425 14992 -361
rect 15056 -425 15072 -361
rect 15136 -425 15278 -361
rect 15342 -425 15358 -361
rect 15422 -425 15438 -361
rect 15502 -425 15518 -361
rect 15582 -425 15598 -361
rect 15662 -425 15678 -361
rect 15742 -425 15884 -361
rect 15948 -425 15964 -361
rect 16028 -425 16044 -361
rect 16108 -425 16124 -361
rect 16188 -425 16204 -361
rect 16268 -425 16284 -361
rect 16348 -425 16490 -361
rect 16554 -425 16570 -361
rect 16634 -425 16650 -361
rect 16714 -425 16730 -361
rect 16794 -425 16810 -361
rect 16874 -425 16890 -361
rect 16954 -425 17096 -361
rect 17160 -425 17176 -361
rect 17240 -425 17256 -361
rect 17320 -425 17336 -361
rect 17400 -425 17416 -361
rect 17480 -425 17496 -361
rect 17560 -425 17702 -361
rect 17766 -425 17782 -361
rect 17846 -425 17862 -361
rect 17926 -425 17942 -361
rect 18006 -425 18022 -361
rect 18086 -425 18102 -361
rect 18166 -425 18308 -361
rect 18372 -425 18388 -361
rect 18452 -425 18468 -361
rect 18532 -425 18548 -361
rect 18612 -425 18628 -361
rect 18692 -425 18708 -361
rect 18772 -425 18914 -361
rect 18978 -425 18994 -361
rect 19058 -425 19074 -361
rect 19138 -425 19154 -361
rect 19218 -425 19234 -361
rect 19298 -425 19314 -361
rect 19378 -425 19520 -361
rect 19584 -425 19600 -361
rect 19664 -425 19680 -361
rect 19744 -425 19760 -361
rect 19824 -425 19840 -361
rect 19904 -425 19920 -361
rect 19984 -425 20088 -361
rect 10326 -427 20088 -425
rect 20148 -361 39606 -359
rect 20148 -425 20252 -361
rect 20316 -425 20332 -361
rect 20396 -425 20412 -361
rect 20476 -425 20492 -361
rect 20556 -425 20572 -361
rect 20636 -425 20652 -361
rect 20716 -425 20858 -361
rect 20922 -425 20938 -361
rect 21002 -425 21018 -361
rect 21082 -425 21098 -361
rect 21162 -425 21178 -361
rect 21242 -425 21258 -361
rect 21322 -425 21464 -361
rect 21528 -425 21544 -361
rect 21608 -425 21624 -361
rect 21688 -425 21704 -361
rect 21768 -425 21784 -361
rect 21848 -425 21864 -361
rect 21928 -425 22070 -361
rect 22134 -425 22150 -361
rect 22214 -425 22230 -361
rect 22294 -425 22310 -361
rect 22374 -425 22390 -361
rect 22454 -425 22470 -361
rect 22534 -425 22676 -361
rect 22740 -425 22756 -361
rect 22820 -425 22836 -361
rect 22900 -425 22916 -361
rect 22980 -425 22996 -361
rect 23060 -425 23076 -361
rect 23140 -425 23282 -361
rect 23346 -425 23362 -361
rect 23426 -425 23442 -361
rect 23506 -425 23522 -361
rect 23586 -425 23602 -361
rect 23666 -425 23682 -361
rect 23746 -425 23888 -361
rect 23952 -425 23968 -361
rect 24032 -425 24048 -361
rect 24112 -425 24128 -361
rect 24192 -425 24208 -361
rect 24272 -425 24288 -361
rect 24352 -425 24494 -361
rect 24558 -425 24574 -361
rect 24638 -425 24654 -361
rect 24718 -425 24734 -361
rect 24798 -425 24814 -361
rect 24878 -425 24894 -361
rect 24958 -425 25100 -361
rect 25164 -425 25180 -361
rect 25244 -425 25260 -361
rect 25324 -425 25340 -361
rect 25404 -425 25420 -361
rect 25484 -425 25500 -361
rect 25564 -425 25706 -361
rect 25770 -425 25786 -361
rect 25850 -425 25866 -361
rect 25930 -425 25946 -361
rect 26010 -425 26026 -361
rect 26090 -425 26106 -361
rect 26170 -425 26312 -361
rect 26376 -425 26392 -361
rect 26456 -425 26472 -361
rect 26536 -425 26552 -361
rect 26616 -425 26632 -361
rect 26696 -425 26712 -361
rect 26776 -425 26918 -361
rect 26982 -425 26998 -361
rect 27062 -425 27078 -361
rect 27142 -425 27158 -361
rect 27222 -425 27238 -361
rect 27302 -425 27318 -361
rect 27382 -425 27524 -361
rect 27588 -425 27604 -361
rect 27668 -425 27684 -361
rect 27748 -425 27764 -361
rect 27828 -425 27844 -361
rect 27908 -425 27924 -361
rect 27988 -425 28130 -361
rect 28194 -425 28210 -361
rect 28274 -425 28290 -361
rect 28354 -425 28370 -361
rect 28434 -425 28450 -361
rect 28514 -425 28530 -361
rect 28594 -425 28736 -361
rect 28800 -425 28816 -361
rect 28880 -425 28896 -361
rect 28960 -425 28976 -361
rect 29040 -425 29056 -361
rect 29120 -425 29136 -361
rect 29200 -425 29342 -361
rect 29406 -425 29422 -361
rect 29486 -425 29502 -361
rect 29566 -425 29582 -361
rect 29646 -425 29662 -361
rect 29726 -425 29742 -361
rect 29806 -425 29948 -361
rect 30012 -425 30028 -361
rect 30092 -425 30108 -361
rect 30172 -425 30188 -361
rect 30252 -425 30268 -361
rect 30332 -425 30348 -361
rect 30412 -425 30554 -361
rect 30618 -425 30634 -361
rect 30698 -425 30714 -361
rect 30778 -425 30794 -361
rect 30858 -425 30874 -361
rect 30938 -425 30954 -361
rect 31018 -425 31160 -361
rect 31224 -425 31240 -361
rect 31304 -425 31320 -361
rect 31384 -425 31400 -361
rect 31464 -425 31480 -361
rect 31544 -425 31560 -361
rect 31624 -425 31766 -361
rect 31830 -425 31846 -361
rect 31910 -425 31926 -361
rect 31990 -425 32006 -361
rect 32070 -425 32086 -361
rect 32150 -425 32166 -361
rect 32230 -425 32372 -361
rect 32436 -425 32452 -361
rect 32516 -425 32532 -361
rect 32596 -425 32612 -361
rect 32676 -425 32692 -361
rect 32756 -425 32772 -361
rect 32836 -425 32978 -361
rect 33042 -425 33058 -361
rect 33122 -425 33138 -361
rect 33202 -425 33218 -361
rect 33282 -425 33298 -361
rect 33362 -425 33378 -361
rect 33442 -425 33584 -361
rect 33648 -425 33664 -361
rect 33728 -425 33744 -361
rect 33808 -425 33824 -361
rect 33888 -425 33904 -361
rect 33968 -425 33984 -361
rect 34048 -425 34190 -361
rect 34254 -425 34270 -361
rect 34334 -425 34350 -361
rect 34414 -425 34430 -361
rect 34494 -425 34510 -361
rect 34574 -425 34590 -361
rect 34654 -425 34796 -361
rect 34860 -425 34876 -361
rect 34940 -425 34956 -361
rect 35020 -425 35036 -361
rect 35100 -425 35116 -361
rect 35180 -425 35196 -361
rect 35260 -425 35402 -361
rect 35466 -425 35482 -361
rect 35546 -425 35562 -361
rect 35626 -425 35642 -361
rect 35706 -425 35722 -361
rect 35786 -425 35802 -361
rect 35866 -425 36008 -361
rect 36072 -425 36088 -361
rect 36152 -425 36168 -361
rect 36232 -425 36248 -361
rect 36312 -425 36328 -361
rect 36392 -425 36408 -361
rect 36472 -425 36614 -361
rect 36678 -425 36694 -361
rect 36758 -425 36774 -361
rect 36838 -425 36854 -361
rect 36918 -425 36934 -361
rect 36998 -425 37014 -361
rect 37078 -425 37220 -361
rect 37284 -425 37300 -361
rect 37364 -425 37380 -361
rect 37444 -425 37460 -361
rect 37524 -425 37540 -361
rect 37604 -425 37620 -361
rect 37684 -425 37826 -361
rect 37890 -425 37906 -361
rect 37970 -425 37986 -361
rect 38050 -425 38066 -361
rect 38130 -425 38146 -361
rect 38210 -425 38226 -361
rect 38290 -425 38432 -361
rect 38496 -425 38512 -361
rect 38576 -425 38592 -361
rect 38656 -425 38672 -361
rect 38736 -425 38752 -361
rect 38816 -425 38832 -361
rect 38896 -425 39038 -361
rect 39102 -425 39118 -361
rect 39182 -425 39198 -361
rect 39262 -425 39278 -361
rect 39342 -425 39358 -361
rect 39422 -425 39438 -361
rect 39502 -425 39606 -361
rect 20148 -427 39606 -425
<< via3 >>
rect 38525 6071 38589 6075
rect 38525 6015 38529 6071
rect 38529 6015 38585 6071
rect 38585 6015 38589 6071
rect 38525 6011 38589 6015
rect 37845 5744 37909 5748
rect 37845 5688 37849 5744
rect 37849 5688 37905 5744
rect 37905 5688 37909 5744
rect 37845 5684 37909 5688
rect 39090 5738 39154 5742
rect 39090 5682 39094 5738
rect 39094 5682 39150 5738
rect 39150 5682 39154 5738
rect 39090 5678 39154 5682
rect -355 5028 -291 5092
rect -275 5028 -211 5092
rect -195 5028 -131 5092
rect -115 5028 -51 5092
rect -35 5028 29 5092
rect 45 5028 109 5092
rect 459 5028 523 5092
rect 539 5028 603 5092
rect 619 5028 683 5092
rect 699 5028 763 5092
rect 779 5028 843 5092
rect 859 5028 923 5092
rect 1371 5028 1435 5092
rect 1451 5028 1515 5092
rect 1531 5028 1595 5092
rect 1611 5028 1675 5092
rect 1691 5028 1755 5092
rect 1771 5028 1835 5092
rect 1977 5028 2041 5092
rect 2057 5028 2121 5092
rect 2137 5028 2201 5092
rect 2217 5028 2281 5092
rect 2297 5028 2361 5092
rect 2377 5028 2441 5092
rect 2905 5028 2969 5092
rect 2985 5028 3049 5092
rect 3065 5028 3129 5092
rect 3145 5028 3209 5092
rect 3225 5028 3289 5092
rect 3305 5028 3369 5092
rect 3511 5028 3575 5092
rect 3591 5028 3655 5092
rect 3671 5028 3735 5092
rect 3751 5028 3815 5092
rect 3831 5028 3895 5092
rect 3911 5028 3975 5092
rect 4117 5028 4181 5092
rect 4197 5028 4261 5092
rect 4277 5028 4341 5092
rect 4357 5028 4421 5092
rect 4437 5028 4501 5092
rect 4517 5028 4581 5092
rect 4723 5028 4787 5092
rect 4803 5028 4867 5092
rect 4883 5028 4947 5092
rect 4963 5028 5027 5092
rect 5043 5028 5107 5092
rect 5123 5028 5187 5092
rect 5456 5028 5520 5092
rect 5536 5028 5600 5092
rect 5616 5028 5680 5092
rect 5696 5028 5760 5092
rect 5776 5028 5840 5092
rect 5856 5028 5920 5092
rect 6062 5028 6126 5092
rect 6142 5028 6206 5092
rect 6222 5028 6286 5092
rect 6302 5028 6366 5092
rect 6382 5028 6446 5092
rect 6462 5028 6526 5092
rect 6668 5028 6732 5092
rect 6748 5028 6812 5092
rect 6828 5028 6892 5092
rect 6908 5028 6972 5092
rect 6988 5028 7052 5092
rect 7068 5028 7132 5092
rect 7274 5028 7338 5092
rect 7354 5028 7418 5092
rect 7434 5028 7498 5092
rect 7514 5028 7578 5092
rect 7594 5028 7658 5092
rect 7674 5028 7738 5092
rect 7880 5028 7944 5092
rect 7960 5028 8024 5092
rect 8040 5028 8104 5092
rect 8120 5028 8184 5092
rect 8200 5028 8264 5092
rect 8280 5028 8344 5092
rect 8486 5028 8550 5092
rect 8566 5028 8630 5092
rect 8646 5028 8710 5092
rect 8726 5028 8790 5092
rect 8806 5028 8870 5092
rect 8886 5028 8950 5092
rect 9092 5028 9156 5092
rect 9172 5028 9236 5092
rect 9252 5028 9316 5092
rect 9332 5028 9396 5092
rect 9412 5028 9476 5092
rect 9492 5028 9556 5092
rect 9698 5028 9762 5092
rect 9778 5028 9842 5092
rect 9858 5028 9922 5092
rect 9938 5028 10002 5092
rect 10018 5028 10082 5092
rect 10098 5028 10162 5092
rect 10430 5028 10494 5092
rect 10510 5028 10574 5092
rect 10590 5028 10654 5092
rect 10670 5028 10734 5092
rect 10750 5028 10814 5092
rect 10830 5028 10894 5092
rect 11036 5028 11100 5092
rect 11116 5028 11180 5092
rect 11196 5028 11260 5092
rect 11276 5028 11340 5092
rect 11356 5028 11420 5092
rect 11436 5028 11500 5092
rect 11642 5028 11706 5092
rect 11722 5028 11786 5092
rect 11802 5028 11866 5092
rect 11882 5028 11946 5092
rect 11962 5028 12026 5092
rect 12042 5028 12106 5092
rect 12248 5028 12312 5092
rect 12328 5028 12392 5092
rect 12408 5028 12472 5092
rect 12488 5028 12552 5092
rect 12568 5028 12632 5092
rect 12648 5028 12712 5092
rect 12854 5028 12918 5092
rect 12934 5028 12998 5092
rect 13014 5028 13078 5092
rect 13094 5028 13158 5092
rect 13174 5028 13238 5092
rect 13254 5028 13318 5092
rect 13460 5028 13524 5092
rect 13540 5028 13604 5092
rect 13620 5028 13684 5092
rect 13700 5028 13764 5092
rect 13780 5028 13844 5092
rect 13860 5028 13924 5092
rect 14066 5028 14130 5092
rect 14146 5028 14210 5092
rect 14226 5028 14290 5092
rect 14306 5028 14370 5092
rect 14386 5028 14450 5092
rect 14466 5028 14530 5092
rect 14672 5028 14736 5092
rect 14752 5028 14816 5092
rect 14832 5028 14896 5092
rect 14912 5028 14976 5092
rect 14992 5028 15056 5092
rect 15072 5028 15136 5092
rect 15278 5028 15342 5092
rect 15358 5028 15422 5092
rect 15438 5028 15502 5092
rect 15518 5028 15582 5092
rect 15598 5028 15662 5092
rect 15678 5028 15742 5092
rect 15884 5028 15948 5092
rect 15964 5028 16028 5092
rect 16044 5028 16108 5092
rect 16124 5028 16188 5092
rect 16204 5028 16268 5092
rect 16284 5028 16348 5092
rect 16490 5028 16554 5092
rect 16570 5028 16634 5092
rect 16650 5028 16714 5092
rect 16730 5028 16794 5092
rect 16810 5028 16874 5092
rect 16890 5028 16954 5092
rect 17096 5028 17160 5092
rect 17176 5028 17240 5092
rect 17256 5028 17320 5092
rect 17336 5028 17400 5092
rect 17416 5028 17480 5092
rect 17496 5028 17560 5092
rect 17702 5028 17766 5092
rect 17782 5028 17846 5092
rect 17862 5028 17926 5092
rect 17942 5028 18006 5092
rect 18022 5028 18086 5092
rect 18102 5028 18166 5092
rect 18308 5028 18372 5092
rect 18388 5028 18452 5092
rect 18468 5028 18532 5092
rect 18548 5028 18612 5092
rect 18628 5028 18692 5092
rect 18708 5028 18772 5092
rect 18914 5028 18978 5092
rect 18994 5028 19058 5092
rect 19074 5028 19138 5092
rect 19154 5028 19218 5092
rect 19234 5028 19298 5092
rect 19314 5028 19378 5092
rect 19520 5028 19584 5092
rect 19600 5028 19664 5092
rect 19680 5028 19744 5092
rect 19760 5028 19824 5092
rect 19840 5028 19904 5092
rect 19920 5028 19984 5092
rect 20252 5028 20316 5092
rect 20332 5028 20396 5092
rect 20412 5028 20476 5092
rect 20492 5028 20556 5092
rect 20572 5028 20636 5092
rect 20652 5028 20716 5092
rect 20858 5028 20922 5092
rect 20938 5028 21002 5092
rect 21018 5028 21082 5092
rect 21098 5028 21162 5092
rect 21178 5028 21242 5092
rect 21258 5028 21322 5092
rect 21464 5028 21528 5092
rect 21544 5028 21608 5092
rect 21624 5028 21688 5092
rect 21704 5028 21768 5092
rect 21784 5028 21848 5092
rect 21864 5028 21928 5092
rect 22070 5028 22134 5092
rect 22150 5028 22214 5092
rect 22230 5028 22294 5092
rect 22310 5028 22374 5092
rect 22390 5028 22454 5092
rect 22470 5028 22534 5092
rect 22676 5028 22740 5092
rect 22756 5028 22820 5092
rect 22836 5028 22900 5092
rect 22916 5028 22980 5092
rect 22996 5028 23060 5092
rect 23076 5028 23140 5092
rect 23282 5028 23346 5092
rect 23362 5028 23426 5092
rect 23442 5028 23506 5092
rect 23522 5028 23586 5092
rect 23602 5028 23666 5092
rect 23682 5028 23746 5092
rect 23888 5028 23952 5092
rect 23968 5028 24032 5092
rect 24048 5028 24112 5092
rect 24128 5028 24192 5092
rect 24208 5028 24272 5092
rect 24288 5028 24352 5092
rect 24494 5028 24558 5092
rect 24574 5028 24638 5092
rect 24654 5028 24718 5092
rect 24734 5028 24798 5092
rect 24814 5028 24878 5092
rect 24894 5028 24958 5092
rect 25100 5028 25164 5092
rect 25180 5028 25244 5092
rect 25260 5028 25324 5092
rect 25340 5028 25404 5092
rect 25420 5028 25484 5092
rect 25500 5028 25564 5092
rect 25706 5028 25770 5092
rect 25786 5028 25850 5092
rect 25866 5028 25930 5092
rect 25946 5028 26010 5092
rect 26026 5028 26090 5092
rect 26106 5028 26170 5092
rect 26312 5028 26376 5092
rect 26392 5028 26456 5092
rect 26472 5028 26536 5092
rect 26552 5028 26616 5092
rect 26632 5028 26696 5092
rect 26712 5028 26776 5092
rect 26918 5028 26982 5092
rect 26998 5028 27062 5092
rect 27078 5028 27142 5092
rect 27158 5028 27222 5092
rect 27238 5028 27302 5092
rect 27318 5028 27382 5092
rect 27524 5028 27588 5092
rect 27604 5028 27668 5092
rect 27684 5028 27748 5092
rect 27764 5028 27828 5092
rect 27844 5028 27908 5092
rect 27924 5028 27988 5092
rect 28130 5028 28194 5092
rect 28210 5028 28274 5092
rect 28290 5028 28354 5092
rect 28370 5028 28434 5092
rect 28450 5028 28514 5092
rect 28530 5028 28594 5092
rect 28736 5028 28800 5092
rect 28816 5028 28880 5092
rect 28896 5028 28960 5092
rect 28976 5028 29040 5092
rect 29056 5028 29120 5092
rect 29136 5028 29200 5092
rect 29342 5028 29406 5092
rect 29422 5028 29486 5092
rect 29502 5028 29566 5092
rect 29582 5028 29646 5092
rect 29662 5028 29726 5092
rect 29742 5028 29806 5092
rect 29948 5028 30012 5092
rect 30028 5028 30092 5092
rect 30108 5028 30172 5092
rect 30188 5028 30252 5092
rect 30268 5028 30332 5092
rect 30348 5028 30412 5092
rect 30554 5028 30618 5092
rect 30634 5028 30698 5092
rect 30714 5028 30778 5092
rect 30794 5028 30858 5092
rect 30874 5028 30938 5092
rect 30954 5028 31018 5092
rect 31160 5028 31224 5092
rect 31240 5028 31304 5092
rect 31320 5028 31384 5092
rect 31400 5028 31464 5092
rect 31480 5028 31544 5092
rect 31560 5028 31624 5092
rect 31766 5028 31830 5092
rect 31846 5028 31910 5092
rect 31926 5028 31990 5092
rect 32006 5028 32070 5092
rect 32086 5028 32150 5092
rect 32166 5028 32230 5092
rect 32372 5028 32436 5092
rect 32452 5028 32516 5092
rect 32532 5028 32596 5092
rect 32612 5028 32676 5092
rect 32692 5028 32756 5092
rect 32772 5028 32836 5092
rect 32978 5028 33042 5092
rect 33058 5028 33122 5092
rect 33138 5028 33202 5092
rect 33218 5028 33282 5092
rect 33298 5028 33362 5092
rect 33378 5028 33442 5092
rect 33584 5028 33648 5092
rect 33664 5028 33728 5092
rect 33744 5028 33808 5092
rect 33824 5028 33888 5092
rect 33904 5028 33968 5092
rect 33984 5028 34048 5092
rect 34190 5028 34254 5092
rect 34270 5028 34334 5092
rect 34350 5028 34414 5092
rect 34430 5028 34494 5092
rect 34510 5028 34574 5092
rect 34590 5028 34654 5092
rect 34796 5028 34860 5092
rect 34876 5028 34940 5092
rect 34956 5028 35020 5092
rect 35036 5028 35100 5092
rect 35116 5028 35180 5092
rect 35196 5028 35260 5092
rect 35402 5028 35466 5092
rect 35482 5028 35546 5092
rect 35562 5028 35626 5092
rect 35642 5028 35706 5092
rect 35722 5028 35786 5092
rect 35802 5028 35866 5092
rect 36008 5028 36072 5092
rect 36088 5028 36152 5092
rect 36168 5028 36232 5092
rect 36248 5028 36312 5092
rect 36328 5028 36392 5092
rect 36408 5028 36472 5092
rect 36614 5028 36678 5092
rect 36694 5028 36758 5092
rect 36774 5028 36838 5092
rect 36854 5028 36918 5092
rect 36934 5028 36998 5092
rect 37014 5028 37078 5092
rect 37220 5028 37284 5092
rect 37300 5028 37364 5092
rect 37380 5028 37444 5092
rect 37460 5028 37524 5092
rect 37540 5028 37604 5092
rect 37620 5028 37684 5092
rect 37826 5028 37890 5092
rect 37906 5028 37970 5092
rect 37986 5028 38050 5092
rect 38066 5028 38130 5092
rect 38146 5028 38210 5092
rect 38226 5028 38290 5092
rect 38432 5028 38496 5092
rect 38512 5028 38576 5092
rect 38592 5028 38656 5092
rect 38672 5028 38736 5092
rect 38752 5028 38816 5092
rect 38832 5028 38896 5092
rect 39038 5028 39102 5092
rect 39118 5028 39182 5092
rect 39198 5028 39262 5092
rect 39278 5028 39342 5092
rect 39358 5028 39422 5092
rect 39438 5028 39502 5092
rect -458 4808 -394 4872
rect -458 4728 -394 4792
rect -458 4648 -394 4712
rect -458 4568 -394 4632
rect -458 4488 -394 4552
rect -458 4408 -394 4472
rect -458 4328 -394 4392
rect -458 4248 -394 4312
rect -458 4168 -394 4232
rect -458 4088 -394 4152
rect 148 4808 212 4872
rect 148 4728 212 4792
rect 148 4648 212 4712
rect 148 4568 212 4632
rect 148 4488 212 4552
rect 148 4408 212 4472
rect 148 4328 212 4392
rect 148 4248 212 4312
rect 148 4168 212 4232
rect 148 4088 212 4152
rect 356 4808 420 4872
rect 356 4728 420 4792
rect 356 4648 420 4712
rect 356 4568 420 4632
rect 356 4488 420 4552
rect 356 4408 420 4472
rect 356 4328 420 4392
rect 356 4248 420 4312
rect 356 4168 420 4232
rect 356 4088 420 4152
rect 962 4808 1026 4872
rect 962 4728 1026 4792
rect 962 4648 1026 4712
rect 962 4568 1026 4632
rect 962 4488 1026 4552
rect 962 4408 1026 4472
rect 962 4328 1026 4392
rect 962 4248 1026 4312
rect 962 4168 1026 4232
rect 962 4088 1026 4152
rect -355 3868 -291 3932
rect -275 3868 -211 3932
rect -195 3868 -131 3932
rect -115 3868 -51 3932
rect -35 3868 29 3932
rect 45 3868 109 3932
rect 459 3868 523 3932
rect 539 3868 603 3932
rect 619 3868 683 3932
rect 699 3868 763 3932
rect 779 3868 843 3932
rect 859 3868 923 3932
rect -458 3648 -394 3712
rect -458 3568 -394 3632
rect -458 3488 -394 3552
rect -458 3408 -394 3472
rect -458 3328 -394 3392
rect -458 3248 -394 3312
rect -458 3168 -394 3232
rect -458 3088 -394 3152
rect -458 3008 -394 3072
rect -458 2928 -394 2992
rect 148 3648 212 3712
rect 148 3568 212 3632
rect 148 3488 212 3552
rect 148 3408 212 3472
rect 148 3328 212 3392
rect 148 3248 212 3312
rect 148 3168 212 3232
rect 148 3088 212 3152
rect 148 3008 212 3072
rect 148 2928 212 2992
rect 356 3648 420 3712
rect 356 3568 420 3632
rect 356 3488 420 3552
rect 356 3408 420 3472
rect 356 3328 420 3392
rect 356 3248 420 3312
rect 356 3168 420 3232
rect 356 3088 420 3152
rect 356 3031 360 3072
rect 360 3031 416 3072
rect 416 3031 420 3072
rect 356 3008 420 3031
rect 356 2928 420 2992
rect 962 3648 1026 3712
rect 962 3568 1026 3632
rect 962 3488 1026 3552
rect 962 3408 1026 3472
rect 962 3328 1026 3392
rect 962 3248 1026 3312
rect 962 3168 1026 3232
rect 962 3088 1026 3152
rect 962 3008 1026 3072
rect 962 2928 1026 2992
rect 1268 4808 1332 4872
rect 1268 4728 1332 4792
rect 1268 4648 1332 4712
rect 1268 4568 1332 4632
rect 1268 4488 1332 4552
rect 1268 4408 1332 4472
rect 1268 4328 1332 4392
rect 1268 4248 1332 4312
rect 1268 4168 1332 4232
rect 1268 4088 1332 4152
rect 1874 4808 1938 4872
rect 1874 4728 1938 4792
rect 1874 4648 1938 4712
rect 1874 4568 1938 4632
rect 1874 4488 1938 4552
rect 1874 4408 1938 4472
rect 1874 4328 1938 4392
rect 1874 4248 1938 4312
rect 1874 4168 1938 4232
rect 1874 4088 1938 4152
rect 2480 4808 2544 4872
rect 2480 4728 2544 4792
rect 2480 4648 2544 4712
rect 2480 4568 2544 4632
rect 2480 4488 2544 4552
rect 2480 4408 2544 4472
rect 2480 4328 2544 4392
rect 2480 4248 2544 4312
rect 2480 4168 2544 4232
rect 2480 4088 2544 4152
rect 1371 3868 1435 3932
rect 1451 3868 1515 3932
rect 1531 3868 1595 3932
rect 1611 3868 1675 3932
rect 1691 3868 1755 3932
rect 1771 3868 1835 3932
rect 1977 3868 2041 3932
rect 2057 3868 2121 3932
rect 2137 3868 2201 3932
rect 2217 3868 2281 3932
rect 2297 3868 2361 3932
rect 2377 3868 2441 3932
rect 1268 3648 1332 3712
rect 1268 3568 1332 3632
rect 1268 3488 1332 3552
rect 1268 3408 1332 3472
rect 1268 3328 1332 3392
rect 1268 3248 1332 3312
rect 1268 3168 1332 3232
rect 1268 3088 1332 3152
rect 1268 3008 1332 3072
rect 1268 2928 1332 2992
rect 1874 3648 1938 3712
rect 1874 3568 1938 3632
rect 1874 3488 1938 3552
rect 1874 3408 1938 3472
rect 1874 3328 1938 3392
rect 1874 3248 1938 3312
rect 1874 3168 1938 3232
rect 1874 3088 1938 3152
rect 1874 3008 1938 3072
rect 1874 2928 1938 2992
rect 2480 3648 2544 3712
rect 2480 3568 2544 3632
rect 2480 3488 2544 3552
rect 2480 3408 2544 3472
rect 2480 3328 2544 3392
rect 2480 3248 2544 3312
rect 2480 3168 2544 3232
rect 2480 3088 2544 3152
rect 2480 3008 2544 3072
rect 2480 2928 2544 2992
rect 2802 4808 2866 4872
rect 2802 4728 2866 4792
rect 2802 4648 2866 4712
rect 2802 4568 2866 4632
rect 2802 4488 2866 4552
rect 2802 4408 2866 4472
rect 2802 4328 2866 4392
rect 2802 4248 2866 4312
rect 2802 4168 2866 4232
rect 2802 4088 2866 4152
rect 3408 4808 3472 4872
rect 3408 4728 3472 4792
rect 3408 4648 3472 4712
rect 3408 4568 3472 4632
rect 3408 4488 3472 4552
rect 3408 4408 3472 4472
rect 3408 4328 3472 4392
rect 3408 4248 3472 4312
rect 3408 4168 3472 4232
rect 3408 4088 3472 4152
rect 4014 4808 4078 4872
rect 4014 4728 4078 4792
rect 4014 4648 4078 4712
rect 4014 4568 4078 4632
rect 4014 4488 4078 4552
rect 4014 4408 4078 4472
rect 4014 4328 4078 4392
rect 4014 4248 4078 4312
rect 4014 4168 4078 4232
rect 4014 4088 4078 4152
rect 4620 4808 4684 4872
rect 4620 4728 4684 4792
rect 4620 4648 4684 4712
rect 4620 4568 4684 4632
rect 4620 4488 4684 4552
rect 4620 4408 4684 4472
rect 4620 4328 4684 4392
rect 4620 4248 4684 4312
rect 4620 4168 4684 4232
rect 4620 4088 4684 4152
rect 5226 4808 5290 4872
rect 5226 4728 5290 4792
rect 5226 4648 5290 4712
rect 5226 4568 5290 4632
rect 5226 4488 5290 4552
rect 5226 4408 5290 4472
rect 5226 4328 5290 4392
rect 5226 4248 5290 4312
rect 5226 4168 5290 4232
rect 5226 4088 5290 4152
rect 2905 3868 2969 3932
rect 2985 3868 3049 3932
rect 3065 3868 3129 3932
rect 3145 3868 3209 3932
rect 3225 3868 3289 3932
rect 3305 3868 3369 3932
rect 3511 3868 3575 3932
rect 3591 3868 3655 3932
rect 3671 3868 3735 3932
rect 3751 3868 3815 3932
rect 3831 3868 3895 3932
rect 3911 3868 3975 3932
rect 4117 3868 4181 3932
rect 4197 3868 4261 3932
rect 4277 3868 4341 3932
rect 4357 3868 4421 3932
rect 4437 3868 4501 3932
rect 4517 3868 4581 3932
rect 4723 3868 4787 3932
rect 4803 3868 4867 3932
rect 4883 3868 4947 3932
rect 4963 3868 5027 3932
rect 5043 3927 5107 3932
rect 5123 3927 5187 3932
rect 5043 3871 5106 3927
rect 5106 3871 5107 3927
rect 5123 3871 5162 3927
rect 5162 3871 5187 3927
rect 5043 3868 5107 3871
rect 5123 3868 5187 3871
rect 2802 3648 2866 3712
rect 2802 3568 2866 3632
rect 2802 3488 2866 3552
rect 2802 3408 2866 3472
rect 2802 3328 2866 3392
rect 2802 3248 2866 3312
rect 2802 3168 2866 3232
rect 2802 3088 2866 3152
rect 2802 3008 2866 3072
rect 2802 2928 2866 2992
rect 3408 3648 3472 3712
rect 3408 3568 3472 3632
rect 3408 3488 3472 3552
rect 3408 3408 3472 3472
rect 3408 3328 3472 3392
rect 3408 3248 3472 3312
rect 3408 3168 3472 3232
rect 3408 3088 3472 3152
rect 3408 3008 3472 3072
rect 3408 2928 3472 2992
rect 4014 3648 4078 3712
rect 4014 3568 4078 3632
rect 4014 3488 4078 3552
rect 4014 3408 4078 3472
rect 4014 3328 4078 3392
rect 4014 3248 4078 3312
rect 4014 3168 4078 3232
rect 4014 3088 4078 3152
rect 4014 3008 4078 3072
rect 4014 2928 4078 2992
rect 4620 3648 4684 3712
rect 4620 3568 4684 3632
rect 4620 3488 4684 3552
rect 4620 3408 4684 3472
rect 4620 3328 4684 3392
rect 4620 3248 4684 3312
rect 4620 3168 4684 3232
rect 4620 3088 4684 3152
rect 4620 3008 4684 3072
rect 4620 2928 4684 2992
rect 5226 3648 5290 3712
rect 5226 3568 5290 3632
rect 5226 3488 5290 3552
rect 5226 3408 5290 3472
rect 5226 3328 5290 3392
rect 5226 3248 5290 3312
rect 5226 3168 5290 3232
rect 5226 3088 5290 3152
rect 5226 3008 5290 3072
rect 5226 2928 5290 2992
rect 5353 4808 5417 4872
rect 5353 4728 5417 4792
rect 5353 4648 5417 4712
rect 5353 4568 5417 4632
rect 5353 4488 5417 4552
rect 5353 4408 5417 4472
rect 5353 4328 5417 4392
rect 5353 4248 5417 4312
rect 5353 4168 5417 4232
rect 5353 4088 5417 4152
rect 5959 4808 6023 4872
rect 5959 4728 6023 4792
rect 5959 4648 6023 4712
rect 5959 4568 6023 4632
rect 5959 4488 6023 4552
rect 5959 4408 6023 4472
rect 5959 4328 6023 4392
rect 5959 4248 6023 4312
rect 5959 4168 6023 4232
rect 5959 4088 6023 4152
rect 6565 4808 6629 4872
rect 6565 4728 6629 4792
rect 6565 4648 6629 4712
rect 6565 4568 6629 4632
rect 6565 4488 6629 4552
rect 6565 4408 6629 4472
rect 6565 4328 6629 4392
rect 6565 4248 6629 4312
rect 6565 4168 6629 4232
rect 6565 4088 6629 4152
rect 7171 4808 7235 4872
rect 7171 4728 7235 4792
rect 7171 4648 7235 4712
rect 7171 4568 7235 4632
rect 7171 4488 7235 4552
rect 7171 4408 7235 4472
rect 7171 4328 7235 4392
rect 7171 4248 7235 4312
rect 7171 4168 7235 4232
rect 7171 4088 7235 4152
rect 7777 4808 7841 4872
rect 7777 4728 7841 4792
rect 7777 4648 7841 4712
rect 7777 4568 7841 4632
rect 7777 4488 7841 4552
rect 7777 4408 7841 4472
rect 7777 4328 7841 4392
rect 7777 4248 7841 4312
rect 7777 4168 7841 4232
rect 7777 4088 7841 4152
rect 8383 4808 8447 4872
rect 8383 4728 8447 4792
rect 8383 4648 8447 4712
rect 8383 4568 8447 4632
rect 8383 4488 8447 4552
rect 8383 4408 8447 4472
rect 8383 4328 8447 4392
rect 8383 4248 8447 4312
rect 8383 4168 8447 4232
rect 8383 4088 8447 4152
rect 8989 4808 9053 4872
rect 8989 4728 9053 4792
rect 8989 4648 9053 4712
rect 8989 4568 9053 4632
rect 8989 4488 9053 4552
rect 8989 4408 9053 4472
rect 8989 4328 9053 4392
rect 8989 4248 9053 4312
rect 8989 4168 9053 4232
rect 8989 4088 9053 4152
rect 9595 4808 9659 4872
rect 9595 4728 9659 4792
rect 9595 4648 9659 4712
rect 9595 4568 9659 4632
rect 9595 4488 9659 4552
rect 9595 4408 9659 4472
rect 9595 4328 9659 4392
rect 9595 4248 9659 4312
rect 9595 4168 9659 4232
rect 9595 4088 9659 4152
rect 10201 4808 10265 4872
rect 10201 4728 10265 4792
rect 10201 4648 10265 4712
rect 10201 4568 10265 4632
rect 10201 4488 10265 4552
rect 10201 4408 10265 4472
rect 10201 4328 10265 4392
rect 10201 4248 10265 4312
rect 10201 4168 10265 4232
rect 10201 4088 10265 4152
rect 5456 3868 5520 3932
rect 5536 3868 5600 3932
rect 5616 3868 5680 3932
rect 5696 3868 5760 3932
rect 5776 3868 5840 3932
rect 5856 3868 5920 3932
rect 6062 3868 6126 3932
rect 6142 3868 6206 3932
rect 6222 3868 6286 3932
rect 6302 3868 6366 3932
rect 6382 3868 6446 3932
rect 6462 3868 6526 3932
rect 6668 3868 6732 3932
rect 6748 3868 6812 3932
rect 6828 3868 6892 3932
rect 6908 3868 6972 3932
rect 6988 3868 7052 3932
rect 7068 3868 7132 3932
rect 7274 3868 7338 3932
rect 7354 3868 7418 3932
rect 7434 3868 7498 3932
rect 7514 3868 7578 3932
rect 7594 3868 7658 3932
rect 7674 3868 7738 3932
rect 7880 3868 7944 3932
rect 7960 3868 8024 3932
rect 8040 3868 8104 3932
rect 8120 3868 8184 3932
rect 8200 3868 8264 3932
rect 8280 3868 8344 3932
rect 8486 3868 8550 3932
rect 8566 3868 8630 3932
rect 8646 3868 8710 3932
rect 8726 3868 8790 3932
rect 8806 3868 8870 3932
rect 8886 3868 8950 3932
rect 9092 3868 9156 3932
rect 9172 3868 9236 3932
rect 9252 3868 9316 3932
rect 9332 3868 9396 3932
rect 9412 3868 9476 3932
rect 9492 3868 9556 3932
rect 9698 3868 9762 3932
rect 9778 3868 9842 3932
rect 9858 3868 9922 3932
rect 9938 3868 10002 3932
rect 10018 3868 10082 3932
rect 10098 3868 10162 3932
rect 5353 3648 5417 3712
rect 5353 3568 5417 3632
rect 5353 3488 5417 3552
rect 5353 3408 5417 3472
rect 5353 3328 5417 3392
rect 5353 3248 5417 3312
rect 5353 3168 5417 3232
rect 5353 3088 5417 3152
rect 5353 3008 5417 3072
rect 5353 2928 5417 2992
rect 5959 3648 6023 3712
rect 5959 3568 6023 3632
rect 5959 3488 6023 3552
rect 5959 3408 6023 3472
rect 5959 3328 6023 3392
rect 5959 3248 6023 3312
rect 5959 3168 6023 3232
rect 5959 3088 6023 3152
rect 5959 3008 6023 3072
rect 5959 2928 6023 2992
rect 6565 3648 6629 3712
rect 6565 3568 6629 3632
rect 6565 3488 6629 3552
rect 6565 3408 6629 3472
rect 6565 3328 6629 3392
rect 6565 3248 6629 3312
rect 6565 3168 6629 3232
rect 6565 3088 6629 3152
rect 6565 3008 6629 3072
rect 6565 2928 6629 2992
rect 7171 3648 7235 3712
rect 7171 3568 7235 3632
rect 7171 3488 7235 3552
rect 7171 3408 7235 3472
rect 7171 3328 7235 3392
rect 7171 3248 7235 3312
rect 7171 3168 7235 3232
rect 7171 3088 7235 3152
rect 7171 3008 7235 3072
rect 7171 2928 7235 2992
rect 7777 3648 7841 3712
rect 7777 3568 7841 3632
rect 7777 3488 7841 3552
rect 7777 3408 7841 3472
rect 7777 3328 7841 3392
rect 7777 3248 7841 3312
rect 7777 3168 7841 3232
rect 7777 3088 7841 3152
rect 7777 3008 7841 3072
rect 7777 2928 7841 2992
rect 8383 3648 8447 3712
rect 8383 3568 8447 3632
rect 8383 3488 8447 3552
rect 8383 3408 8447 3472
rect 8383 3328 8447 3392
rect 8383 3248 8447 3312
rect 8383 3168 8447 3232
rect 8383 3088 8447 3152
rect 8383 3008 8447 3072
rect 8383 2928 8447 2992
rect 8989 3648 9053 3712
rect 8989 3568 9053 3632
rect 8989 3488 9053 3552
rect 8989 3408 9053 3472
rect 8989 3328 9053 3392
rect 8989 3248 9053 3312
rect 8989 3168 9053 3232
rect 8989 3088 9053 3152
rect 8989 3008 9053 3072
rect 8989 2928 9053 2992
rect 9595 3648 9659 3712
rect 9595 3568 9659 3632
rect 9595 3488 9659 3552
rect 9595 3408 9659 3472
rect 9595 3328 9659 3392
rect 9595 3248 9659 3312
rect 9595 3168 9659 3232
rect 9595 3088 9659 3152
rect 9595 3008 9659 3072
rect 9595 2928 9659 2992
rect 10201 3648 10265 3712
rect 10201 3568 10265 3632
rect 10201 3488 10265 3552
rect 10201 3408 10265 3472
rect 10201 3328 10265 3392
rect 10201 3248 10265 3312
rect 10201 3168 10265 3232
rect 10201 3088 10265 3152
rect 10201 3008 10265 3072
rect 10201 2928 10265 2992
rect 10327 4808 10391 4872
rect 10327 4728 10391 4792
rect 10327 4648 10391 4712
rect 10327 4568 10391 4632
rect 10327 4488 10391 4552
rect 10327 4408 10391 4472
rect 10327 4328 10391 4392
rect 10327 4248 10391 4312
rect 10327 4168 10391 4232
rect 10327 4088 10391 4152
rect 10933 4808 10997 4872
rect 10933 4728 10997 4792
rect 10933 4648 10997 4712
rect 10933 4568 10997 4632
rect 10933 4488 10997 4552
rect 10933 4408 10997 4472
rect 10933 4328 10997 4392
rect 10933 4248 10997 4312
rect 10933 4168 10997 4232
rect 10933 4088 10997 4152
rect 11539 4808 11603 4872
rect 11539 4728 11603 4792
rect 11539 4648 11603 4712
rect 11539 4568 11603 4632
rect 11539 4488 11603 4552
rect 11539 4408 11603 4472
rect 11539 4328 11603 4392
rect 11539 4248 11603 4312
rect 11539 4168 11603 4232
rect 11539 4088 11603 4152
rect 12145 4808 12209 4872
rect 12145 4728 12209 4792
rect 12145 4648 12209 4712
rect 12145 4568 12209 4632
rect 12145 4488 12209 4552
rect 12145 4408 12209 4472
rect 12145 4328 12209 4392
rect 12145 4248 12209 4312
rect 12145 4168 12209 4232
rect 12145 4088 12209 4152
rect 12751 4808 12815 4872
rect 12751 4728 12815 4792
rect 12751 4648 12815 4712
rect 12751 4568 12815 4632
rect 12751 4488 12815 4552
rect 12751 4408 12815 4472
rect 12751 4328 12815 4392
rect 12751 4248 12815 4312
rect 12751 4168 12815 4232
rect 12751 4088 12815 4152
rect 13357 4808 13421 4872
rect 13357 4728 13421 4792
rect 13357 4648 13421 4712
rect 13357 4568 13421 4632
rect 13357 4488 13421 4552
rect 13357 4408 13421 4472
rect 13357 4328 13421 4392
rect 13357 4248 13421 4312
rect 13357 4168 13421 4232
rect 13357 4088 13421 4152
rect 13963 4808 14027 4872
rect 13963 4728 14027 4792
rect 13963 4648 14027 4712
rect 13963 4568 14027 4632
rect 13963 4488 14027 4552
rect 13963 4408 14027 4472
rect 13963 4328 14027 4392
rect 13963 4248 14027 4312
rect 13963 4168 14027 4232
rect 13963 4088 14027 4152
rect 14569 4808 14633 4872
rect 14569 4728 14633 4792
rect 14569 4648 14633 4712
rect 14569 4568 14633 4632
rect 14569 4488 14633 4552
rect 14569 4408 14633 4472
rect 14569 4328 14633 4392
rect 14569 4248 14633 4312
rect 14569 4168 14633 4232
rect 14569 4088 14633 4152
rect 15175 4808 15239 4872
rect 15175 4728 15239 4792
rect 15175 4648 15239 4712
rect 15175 4568 15239 4632
rect 15175 4488 15239 4552
rect 15175 4408 15239 4472
rect 15175 4328 15239 4392
rect 15175 4248 15239 4312
rect 15175 4168 15239 4232
rect 15175 4088 15239 4152
rect 15781 4808 15845 4872
rect 15781 4728 15845 4792
rect 15781 4648 15845 4712
rect 15781 4568 15845 4632
rect 15781 4488 15845 4552
rect 15781 4408 15845 4472
rect 15781 4328 15845 4392
rect 15781 4248 15845 4312
rect 15781 4168 15845 4232
rect 15781 4088 15845 4152
rect 16387 4808 16451 4872
rect 16387 4728 16451 4792
rect 16387 4648 16451 4712
rect 16387 4568 16451 4632
rect 16387 4488 16451 4552
rect 16387 4408 16451 4472
rect 16387 4328 16451 4392
rect 16387 4248 16451 4312
rect 16387 4168 16451 4232
rect 16387 4088 16451 4152
rect 16993 4808 17057 4872
rect 16993 4728 17057 4792
rect 16993 4648 17057 4712
rect 16993 4568 17057 4632
rect 16993 4488 17057 4552
rect 16993 4408 17057 4472
rect 16993 4328 17057 4392
rect 16993 4248 17057 4312
rect 16993 4168 17057 4232
rect 16993 4088 17057 4152
rect 17599 4808 17663 4872
rect 17599 4728 17663 4792
rect 17599 4648 17663 4712
rect 17599 4568 17663 4632
rect 17599 4488 17663 4552
rect 17599 4408 17663 4472
rect 17599 4328 17663 4392
rect 17599 4248 17663 4312
rect 17599 4168 17663 4232
rect 17599 4088 17663 4152
rect 18205 4808 18269 4872
rect 18205 4728 18269 4792
rect 18205 4648 18269 4712
rect 18205 4568 18269 4632
rect 18205 4488 18269 4552
rect 18205 4408 18269 4472
rect 18205 4328 18269 4392
rect 18205 4248 18269 4312
rect 18205 4168 18269 4232
rect 18205 4088 18269 4152
rect 18811 4808 18875 4872
rect 18811 4728 18875 4792
rect 18811 4648 18875 4712
rect 18811 4568 18875 4632
rect 18811 4488 18875 4552
rect 18811 4408 18875 4472
rect 18811 4328 18875 4392
rect 18811 4248 18875 4312
rect 18811 4168 18875 4232
rect 18811 4088 18875 4152
rect 19417 4808 19481 4872
rect 19417 4728 19481 4792
rect 19417 4648 19481 4712
rect 19417 4568 19481 4632
rect 19417 4488 19481 4552
rect 19417 4408 19481 4472
rect 19417 4328 19481 4392
rect 19417 4248 19481 4312
rect 19417 4168 19481 4232
rect 19417 4088 19481 4152
rect 20023 4808 20087 4872
rect 20023 4728 20087 4792
rect 20023 4648 20087 4712
rect 20023 4568 20087 4632
rect 20023 4488 20087 4552
rect 20023 4408 20087 4472
rect 20023 4328 20087 4392
rect 20023 4248 20087 4312
rect 20023 4168 20087 4232
rect 20023 4088 20087 4152
rect 10430 3868 10494 3932
rect 10510 3868 10574 3932
rect 10590 3868 10654 3932
rect 10670 3868 10734 3932
rect 10750 3868 10814 3932
rect 10830 3868 10894 3932
rect 11036 3868 11100 3932
rect 11116 3868 11180 3932
rect 11196 3868 11260 3932
rect 11276 3868 11340 3932
rect 11356 3868 11420 3932
rect 11436 3868 11500 3932
rect 11642 3868 11706 3932
rect 11722 3868 11786 3932
rect 11802 3868 11866 3932
rect 11882 3868 11946 3932
rect 11962 3868 12026 3932
rect 12042 3868 12106 3932
rect 12248 3868 12312 3932
rect 12328 3868 12392 3932
rect 12408 3868 12472 3932
rect 12488 3868 12552 3932
rect 12568 3868 12632 3932
rect 12648 3868 12712 3932
rect 12854 3868 12918 3932
rect 12934 3868 12998 3932
rect 13014 3868 13078 3932
rect 13094 3868 13158 3932
rect 13174 3868 13238 3932
rect 13254 3868 13318 3932
rect 13460 3868 13524 3932
rect 13540 3868 13604 3932
rect 13620 3868 13684 3932
rect 13700 3868 13764 3932
rect 13780 3868 13844 3932
rect 13860 3868 13924 3932
rect 14066 3868 14130 3932
rect 14146 3868 14210 3932
rect 14226 3868 14290 3932
rect 14306 3868 14370 3932
rect 14386 3868 14450 3932
rect 14466 3868 14530 3932
rect 14672 3868 14736 3932
rect 14752 3868 14816 3932
rect 14832 3868 14896 3932
rect 14912 3868 14976 3932
rect 14992 3868 15056 3932
rect 15072 3868 15136 3932
rect 15278 3868 15342 3932
rect 15358 3868 15422 3932
rect 15438 3868 15502 3932
rect 15518 3868 15582 3932
rect 15598 3868 15662 3932
rect 15678 3868 15742 3932
rect 15884 3868 15948 3932
rect 15964 3868 16028 3932
rect 16044 3868 16108 3932
rect 16124 3868 16188 3932
rect 16204 3868 16268 3932
rect 16284 3868 16348 3932
rect 16490 3868 16554 3932
rect 16570 3868 16634 3932
rect 16650 3868 16714 3932
rect 16730 3868 16794 3932
rect 16810 3868 16874 3932
rect 16890 3868 16954 3932
rect 17096 3868 17160 3932
rect 17176 3868 17240 3932
rect 17256 3868 17320 3932
rect 17336 3868 17400 3932
rect 17416 3868 17480 3932
rect 17496 3868 17560 3932
rect 17702 3868 17766 3932
rect 17782 3868 17846 3932
rect 17862 3868 17926 3932
rect 17942 3868 18006 3932
rect 18022 3868 18086 3932
rect 18102 3868 18166 3932
rect 18308 3868 18372 3932
rect 18388 3868 18452 3932
rect 18468 3868 18532 3932
rect 18548 3868 18612 3932
rect 18628 3868 18692 3932
rect 18708 3868 18772 3932
rect 18914 3868 18978 3932
rect 18994 3868 19058 3932
rect 19074 3868 19138 3932
rect 19154 3868 19218 3932
rect 19234 3868 19298 3932
rect 19314 3868 19378 3932
rect 19520 3868 19584 3932
rect 19600 3868 19664 3932
rect 19680 3868 19744 3932
rect 19760 3868 19824 3932
rect 19840 3868 19904 3932
rect 19920 3868 19984 3932
rect 10327 3648 10391 3712
rect 10327 3568 10391 3632
rect 10327 3488 10391 3552
rect 10327 3408 10391 3472
rect 10327 3328 10391 3392
rect 10327 3248 10391 3312
rect 10327 3168 10391 3232
rect 10327 3088 10391 3152
rect 10327 3008 10391 3072
rect 10327 2928 10391 2992
rect 10933 3648 10997 3712
rect 10933 3568 10997 3632
rect 10933 3488 10997 3552
rect 10933 3408 10997 3472
rect 10933 3328 10997 3392
rect 10933 3248 10997 3312
rect 10933 3168 10997 3232
rect 10933 3088 10997 3152
rect 10933 3008 10997 3072
rect 10933 2928 10997 2992
rect 11539 3648 11603 3712
rect 11539 3568 11603 3632
rect 11539 3488 11603 3552
rect 11539 3408 11603 3472
rect 11539 3328 11603 3392
rect 11539 3248 11603 3312
rect 11539 3168 11603 3232
rect 11539 3088 11603 3152
rect 11539 3008 11603 3072
rect 11539 2928 11603 2992
rect 12145 3648 12209 3712
rect 12145 3568 12209 3632
rect 12145 3488 12209 3552
rect 12145 3408 12209 3472
rect 12145 3328 12209 3392
rect 12145 3248 12209 3312
rect 12145 3168 12209 3232
rect 12145 3088 12209 3152
rect 12145 3008 12209 3072
rect 12145 2928 12209 2992
rect 12751 3648 12815 3712
rect 12751 3568 12815 3632
rect 12751 3488 12815 3552
rect 12751 3408 12815 3472
rect 12751 3328 12815 3392
rect 12751 3248 12815 3312
rect 12751 3168 12815 3232
rect 12751 3088 12815 3152
rect 12751 3008 12815 3072
rect 12751 2928 12815 2992
rect 13357 3648 13421 3712
rect 13357 3568 13421 3632
rect 13357 3488 13421 3552
rect 13357 3408 13421 3472
rect 13357 3328 13421 3392
rect 13357 3248 13421 3312
rect 13357 3168 13421 3232
rect 13357 3088 13421 3152
rect 13357 3008 13421 3072
rect 13357 2928 13421 2992
rect 13963 3648 14027 3712
rect 13963 3568 14027 3632
rect 13963 3488 14027 3552
rect 13963 3408 14027 3472
rect 13963 3328 14027 3392
rect 13963 3248 14027 3312
rect 13963 3168 14027 3232
rect 13963 3088 14027 3152
rect 13963 3008 14027 3072
rect 13963 2928 14027 2992
rect 14569 3648 14633 3712
rect 14569 3568 14633 3632
rect 14569 3488 14633 3552
rect 14569 3408 14633 3472
rect 14569 3328 14633 3392
rect 14569 3248 14633 3312
rect 14569 3168 14633 3232
rect 14569 3088 14633 3152
rect 14569 3008 14633 3072
rect 14569 2928 14633 2992
rect 15175 3648 15239 3712
rect 15175 3568 15239 3632
rect 15175 3488 15239 3552
rect 15175 3408 15239 3472
rect 15175 3328 15239 3392
rect 15175 3248 15239 3312
rect 15175 3168 15239 3232
rect 15175 3088 15239 3152
rect 15175 3008 15239 3072
rect 15175 2928 15239 2992
rect 15781 3648 15845 3712
rect 15781 3568 15845 3632
rect 15781 3488 15845 3552
rect 15781 3408 15845 3472
rect 15781 3328 15845 3392
rect 15781 3248 15845 3312
rect 15781 3168 15845 3232
rect 15781 3088 15845 3152
rect 15781 3008 15845 3072
rect 15781 2928 15845 2992
rect 16387 3648 16451 3712
rect 16387 3568 16451 3632
rect 16387 3488 16451 3552
rect 16387 3408 16451 3472
rect 16387 3328 16451 3392
rect 16387 3248 16451 3312
rect 16387 3168 16451 3232
rect 16387 3088 16451 3152
rect 16387 3008 16451 3072
rect 16387 2928 16451 2992
rect 16993 3648 17057 3712
rect 16993 3568 17057 3632
rect 16993 3488 17057 3552
rect 16993 3408 17057 3472
rect 16993 3328 17057 3392
rect 16993 3248 17057 3312
rect 16993 3168 17057 3232
rect 16993 3088 17057 3152
rect 16993 3008 17057 3072
rect 16993 2928 17057 2992
rect 17599 3648 17663 3712
rect 17599 3568 17663 3632
rect 17599 3488 17663 3552
rect 17599 3408 17663 3472
rect 17599 3328 17663 3392
rect 17599 3248 17663 3312
rect 17599 3168 17663 3232
rect 17599 3088 17663 3152
rect 17599 3008 17663 3072
rect 17599 2928 17663 2992
rect 18205 3648 18269 3712
rect 18205 3568 18269 3632
rect 18205 3488 18269 3552
rect 18205 3408 18269 3472
rect 18205 3328 18269 3392
rect 18205 3248 18269 3312
rect 18205 3168 18269 3232
rect 18205 3088 18269 3152
rect 18205 3008 18269 3072
rect 18205 2928 18269 2992
rect 18811 3648 18875 3712
rect 18811 3568 18875 3632
rect 18811 3488 18875 3552
rect 18811 3408 18875 3472
rect 18811 3328 18875 3392
rect 18811 3248 18875 3312
rect 18811 3168 18875 3232
rect 18811 3088 18875 3152
rect 18811 3008 18875 3072
rect 18811 2928 18875 2992
rect 19417 3648 19481 3712
rect 19417 3568 19481 3632
rect 19417 3488 19481 3552
rect 19417 3408 19481 3472
rect 19417 3328 19481 3392
rect 19417 3248 19481 3312
rect 19417 3168 19481 3232
rect 19417 3088 19481 3152
rect 19417 3008 19481 3072
rect 19417 2928 19481 2992
rect 20023 3648 20087 3712
rect 20023 3568 20087 3632
rect 20023 3488 20087 3552
rect 20023 3408 20087 3472
rect 20023 3328 20087 3392
rect 20023 3248 20087 3312
rect 20023 3168 20087 3232
rect 20023 3088 20087 3152
rect 20023 3008 20087 3072
rect 20023 2928 20087 2992
rect 20149 4808 20213 4872
rect 20149 4728 20213 4792
rect 20149 4648 20213 4712
rect 20149 4568 20213 4632
rect 20149 4488 20213 4552
rect 20149 4408 20213 4472
rect 20149 4328 20213 4392
rect 20149 4248 20213 4312
rect 20149 4168 20213 4232
rect 20149 4088 20213 4152
rect 20755 4808 20819 4872
rect 20755 4728 20819 4792
rect 20755 4648 20819 4712
rect 20755 4568 20819 4632
rect 20755 4488 20819 4552
rect 20755 4408 20819 4472
rect 20755 4328 20819 4392
rect 20755 4248 20819 4312
rect 20755 4168 20819 4232
rect 20755 4088 20819 4152
rect 21361 4808 21425 4872
rect 21361 4728 21425 4792
rect 21361 4648 21425 4712
rect 21361 4568 21425 4632
rect 21361 4488 21425 4552
rect 21361 4408 21425 4472
rect 21361 4328 21425 4392
rect 21361 4248 21425 4312
rect 21361 4168 21425 4232
rect 21361 4088 21425 4152
rect 21967 4808 22031 4872
rect 21967 4728 22031 4792
rect 21967 4648 22031 4712
rect 21967 4568 22031 4632
rect 21967 4488 22031 4552
rect 21967 4408 22031 4472
rect 21967 4328 22031 4392
rect 21967 4248 22031 4312
rect 21967 4168 22031 4232
rect 21967 4088 22031 4152
rect 22573 4808 22637 4872
rect 22573 4728 22637 4792
rect 22573 4648 22637 4712
rect 22573 4568 22637 4632
rect 22573 4488 22637 4552
rect 22573 4408 22637 4472
rect 22573 4328 22637 4392
rect 22573 4248 22637 4312
rect 22573 4168 22637 4232
rect 22573 4088 22637 4152
rect 23179 4808 23243 4872
rect 23179 4728 23243 4792
rect 23179 4648 23243 4712
rect 23179 4568 23243 4632
rect 23179 4488 23243 4552
rect 23179 4408 23243 4472
rect 23179 4328 23243 4392
rect 23179 4248 23243 4312
rect 23179 4168 23243 4232
rect 23179 4088 23243 4152
rect 23785 4808 23849 4872
rect 23785 4728 23849 4792
rect 23785 4648 23849 4712
rect 23785 4568 23849 4632
rect 23785 4488 23849 4552
rect 23785 4408 23849 4472
rect 23785 4328 23849 4392
rect 23785 4248 23849 4312
rect 23785 4168 23849 4232
rect 23785 4088 23849 4152
rect 24391 4808 24455 4872
rect 24391 4728 24455 4792
rect 24391 4648 24455 4712
rect 24391 4568 24455 4632
rect 24391 4488 24455 4552
rect 24391 4408 24455 4472
rect 24391 4328 24455 4392
rect 24391 4248 24455 4312
rect 24391 4168 24455 4232
rect 24391 4088 24455 4152
rect 24997 4808 25061 4872
rect 24997 4728 25061 4792
rect 24997 4648 25061 4712
rect 24997 4568 25061 4632
rect 24997 4488 25061 4552
rect 24997 4408 25061 4472
rect 24997 4328 25061 4392
rect 24997 4248 25061 4312
rect 24997 4168 25061 4232
rect 24997 4088 25061 4152
rect 25603 4808 25667 4872
rect 25603 4728 25667 4792
rect 25603 4648 25667 4712
rect 25603 4568 25667 4632
rect 25603 4488 25667 4552
rect 25603 4408 25667 4472
rect 25603 4328 25667 4392
rect 25603 4248 25667 4312
rect 25603 4168 25667 4232
rect 25603 4088 25667 4152
rect 26209 4808 26273 4872
rect 26209 4728 26273 4792
rect 26209 4648 26273 4712
rect 26209 4568 26273 4632
rect 26209 4488 26273 4552
rect 26209 4408 26273 4472
rect 26209 4328 26273 4392
rect 26209 4248 26273 4312
rect 26209 4168 26273 4232
rect 26209 4088 26273 4152
rect 26815 4808 26879 4872
rect 26815 4728 26879 4792
rect 26815 4648 26879 4712
rect 26815 4568 26879 4632
rect 26815 4488 26879 4552
rect 26815 4408 26879 4472
rect 26815 4328 26879 4392
rect 26815 4248 26879 4312
rect 26815 4168 26879 4232
rect 26815 4088 26879 4152
rect 27421 4808 27485 4872
rect 27421 4728 27485 4792
rect 27421 4648 27485 4712
rect 27421 4568 27485 4632
rect 27421 4488 27485 4552
rect 27421 4408 27485 4472
rect 27421 4328 27485 4392
rect 27421 4248 27485 4312
rect 27421 4168 27485 4232
rect 27421 4088 27485 4152
rect 28027 4808 28091 4872
rect 28027 4728 28091 4792
rect 28027 4648 28091 4712
rect 28027 4568 28091 4632
rect 28027 4488 28091 4552
rect 28027 4408 28091 4472
rect 28027 4328 28091 4392
rect 28027 4248 28091 4312
rect 28027 4168 28091 4232
rect 28027 4088 28091 4152
rect 28633 4808 28697 4872
rect 28633 4728 28697 4792
rect 28633 4648 28697 4712
rect 28633 4568 28697 4632
rect 28633 4488 28697 4552
rect 28633 4408 28697 4472
rect 28633 4328 28697 4392
rect 28633 4248 28697 4312
rect 28633 4168 28697 4232
rect 28633 4088 28697 4152
rect 29239 4808 29303 4872
rect 29239 4728 29303 4792
rect 29239 4648 29303 4712
rect 29239 4568 29303 4632
rect 29239 4488 29303 4552
rect 29239 4408 29303 4472
rect 29239 4328 29303 4392
rect 29239 4248 29303 4312
rect 29239 4168 29303 4232
rect 29239 4088 29303 4152
rect 29845 4808 29909 4872
rect 29845 4728 29909 4792
rect 29845 4648 29909 4712
rect 29845 4568 29909 4632
rect 29845 4488 29909 4552
rect 29845 4408 29909 4472
rect 29845 4328 29909 4392
rect 29845 4248 29909 4312
rect 29845 4168 29909 4232
rect 29845 4088 29909 4152
rect 30451 4808 30515 4872
rect 30451 4728 30515 4792
rect 30451 4648 30515 4712
rect 30451 4568 30515 4632
rect 30451 4488 30515 4552
rect 30451 4408 30515 4472
rect 30451 4328 30515 4392
rect 30451 4248 30515 4312
rect 30451 4168 30515 4232
rect 30451 4088 30515 4152
rect 31057 4808 31121 4872
rect 31057 4728 31121 4792
rect 31057 4648 31121 4712
rect 31057 4568 31121 4632
rect 31057 4488 31121 4552
rect 31057 4408 31121 4472
rect 31057 4328 31121 4392
rect 31057 4248 31121 4312
rect 31057 4168 31121 4232
rect 31057 4088 31121 4152
rect 31663 4808 31727 4872
rect 31663 4728 31727 4792
rect 31663 4648 31727 4712
rect 31663 4568 31727 4632
rect 31663 4488 31727 4552
rect 31663 4408 31727 4472
rect 31663 4328 31727 4392
rect 31663 4248 31727 4312
rect 31663 4168 31727 4232
rect 31663 4088 31727 4152
rect 32269 4808 32333 4872
rect 32269 4728 32333 4792
rect 32269 4648 32333 4712
rect 32269 4568 32333 4632
rect 32269 4488 32333 4552
rect 32269 4408 32333 4472
rect 32269 4328 32333 4392
rect 32269 4248 32333 4312
rect 32269 4168 32333 4232
rect 32269 4088 32333 4152
rect 32875 4808 32939 4872
rect 32875 4728 32939 4792
rect 32875 4648 32939 4712
rect 32875 4568 32939 4632
rect 32875 4488 32939 4552
rect 32875 4408 32939 4472
rect 32875 4328 32939 4392
rect 32875 4248 32939 4312
rect 32875 4168 32939 4232
rect 32875 4088 32939 4152
rect 33481 4808 33545 4872
rect 33481 4728 33545 4792
rect 33481 4648 33545 4712
rect 33481 4568 33545 4632
rect 33481 4488 33545 4552
rect 33481 4408 33545 4472
rect 33481 4328 33545 4392
rect 33481 4248 33545 4312
rect 33481 4168 33545 4232
rect 33481 4088 33545 4152
rect 34087 4808 34151 4872
rect 34087 4728 34151 4792
rect 34087 4648 34151 4712
rect 34087 4568 34151 4632
rect 34087 4488 34151 4552
rect 34087 4408 34151 4472
rect 34087 4328 34151 4392
rect 34087 4248 34151 4312
rect 34087 4168 34151 4232
rect 34087 4088 34151 4152
rect 34693 4808 34757 4872
rect 34693 4728 34757 4792
rect 34693 4648 34757 4712
rect 34693 4568 34757 4632
rect 34693 4488 34757 4552
rect 34693 4408 34757 4472
rect 34693 4328 34757 4392
rect 34693 4248 34757 4312
rect 34693 4168 34757 4232
rect 34693 4088 34757 4152
rect 35299 4808 35363 4872
rect 35299 4728 35363 4792
rect 35299 4648 35363 4712
rect 35299 4568 35363 4632
rect 35299 4488 35363 4552
rect 35299 4408 35363 4472
rect 35299 4328 35363 4392
rect 35299 4248 35363 4312
rect 35299 4168 35363 4232
rect 35299 4088 35363 4152
rect 35905 4808 35969 4872
rect 35905 4728 35969 4792
rect 35905 4648 35969 4712
rect 35905 4568 35969 4632
rect 35905 4488 35969 4552
rect 35905 4408 35969 4472
rect 35905 4328 35969 4392
rect 35905 4248 35969 4312
rect 35905 4168 35969 4232
rect 35905 4088 35969 4152
rect 36511 4808 36575 4872
rect 36511 4728 36575 4792
rect 36511 4648 36575 4712
rect 36511 4568 36575 4632
rect 36511 4488 36575 4552
rect 36511 4408 36575 4472
rect 36511 4328 36575 4392
rect 36511 4248 36575 4312
rect 36511 4168 36575 4232
rect 36511 4088 36575 4152
rect 37117 4808 37181 4872
rect 37117 4728 37181 4792
rect 37117 4648 37181 4712
rect 37117 4568 37181 4632
rect 37117 4488 37181 4552
rect 37117 4408 37181 4472
rect 37117 4328 37181 4392
rect 37117 4248 37181 4312
rect 37117 4168 37181 4232
rect 37117 4088 37181 4152
rect 37723 4808 37787 4872
rect 37723 4728 37787 4792
rect 37723 4648 37787 4712
rect 37723 4568 37787 4632
rect 37723 4488 37787 4552
rect 37723 4408 37787 4472
rect 37723 4328 37787 4392
rect 37723 4248 37787 4312
rect 37723 4168 37787 4232
rect 37723 4088 37787 4152
rect 38329 4808 38393 4872
rect 38329 4728 38393 4792
rect 38329 4648 38393 4712
rect 38329 4568 38393 4632
rect 38329 4488 38393 4552
rect 38329 4408 38393 4472
rect 38329 4328 38393 4392
rect 38329 4248 38393 4312
rect 38329 4168 38393 4232
rect 38329 4088 38393 4152
rect 38935 4808 38999 4872
rect 38935 4728 38999 4792
rect 38935 4648 38999 4712
rect 38935 4568 38999 4632
rect 38935 4488 38999 4552
rect 38935 4408 38999 4472
rect 38935 4328 38999 4392
rect 38935 4248 38999 4312
rect 38935 4168 38999 4232
rect 38935 4088 38999 4152
rect 39541 4808 39605 4872
rect 39541 4728 39605 4792
rect 39541 4648 39605 4712
rect 39541 4568 39605 4632
rect 39541 4488 39605 4552
rect 39541 4408 39605 4472
rect 39541 4328 39605 4392
rect 39541 4248 39605 4312
rect 39541 4168 39605 4232
rect 39541 4088 39605 4152
rect 20252 3868 20316 3932
rect 20332 3868 20396 3932
rect 20412 3868 20476 3932
rect 20492 3868 20556 3932
rect 20572 3868 20636 3932
rect 20652 3868 20716 3932
rect 20858 3868 20922 3932
rect 20938 3868 21002 3932
rect 21018 3868 21082 3932
rect 21098 3868 21162 3932
rect 21178 3868 21242 3932
rect 21258 3868 21322 3932
rect 21464 3868 21528 3932
rect 21544 3868 21608 3932
rect 21624 3868 21688 3932
rect 21704 3868 21768 3932
rect 21784 3868 21848 3932
rect 21864 3868 21928 3932
rect 22070 3868 22134 3932
rect 22150 3868 22214 3932
rect 22230 3868 22294 3932
rect 22310 3868 22374 3932
rect 22390 3868 22454 3932
rect 22470 3868 22534 3932
rect 22676 3868 22740 3932
rect 22756 3868 22820 3932
rect 22836 3868 22900 3932
rect 22916 3868 22980 3932
rect 22996 3868 23060 3932
rect 23076 3868 23140 3932
rect 23282 3868 23346 3932
rect 23362 3868 23426 3932
rect 23442 3868 23506 3932
rect 23522 3868 23586 3932
rect 23602 3868 23666 3932
rect 23682 3868 23746 3932
rect 23888 3868 23952 3932
rect 23968 3868 24032 3932
rect 24048 3868 24112 3932
rect 24128 3868 24192 3932
rect 24208 3868 24272 3932
rect 24288 3868 24352 3932
rect 24494 3868 24558 3932
rect 24574 3868 24638 3932
rect 24654 3868 24718 3932
rect 24734 3868 24798 3932
rect 24814 3868 24878 3932
rect 24894 3868 24958 3932
rect 25100 3868 25164 3932
rect 25180 3868 25244 3932
rect 25260 3868 25324 3932
rect 25340 3868 25404 3932
rect 25420 3868 25484 3932
rect 25500 3868 25564 3932
rect 25706 3868 25770 3932
rect 25786 3868 25850 3932
rect 25866 3868 25930 3932
rect 25946 3868 26010 3932
rect 26026 3868 26090 3932
rect 26106 3868 26170 3932
rect 26312 3868 26376 3932
rect 26392 3868 26456 3932
rect 26472 3868 26536 3932
rect 26552 3868 26616 3932
rect 26632 3868 26696 3932
rect 26712 3868 26776 3932
rect 26918 3868 26982 3932
rect 26998 3868 27062 3932
rect 27078 3868 27142 3932
rect 27158 3868 27222 3932
rect 27238 3868 27302 3932
rect 27318 3868 27382 3932
rect 27524 3868 27588 3932
rect 27604 3868 27668 3932
rect 27684 3868 27748 3932
rect 27764 3868 27828 3932
rect 27844 3868 27908 3932
rect 27924 3868 27988 3932
rect 28130 3868 28194 3932
rect 28210 3868 28274 3932
rect 28290 3868 28354 3932
rect 28370 3868 28434 3932
rect 28450 3868 28514 3932
rect 28530 3868 28594 3932
rect 28736 3868 28800 3932
rect 28816 3868 28880 3932
rect 28896 3868 28960 3932
rect 28976 3868 29040 3932
rect 29056 3868 29120 3932
rect 29136 3868 29200 3932
rect 29342 3868 29406 3932
rect 29422 3868 29486 3932
rect 29502 3868 29566 3932
rect 29582 3868 29646 3932
rect 29662 3868 29726 3932
rect 29742 3868 29806 3932
rect 29948 3868 30012 3932
rect 30028 3868 30092 3932
rect 30108 3868 30172 3932
rect 30188 3868 30252 3932
rect 30268 3868 30332 3932
rect 30348 3868 30412 3932
rect 30554 3868 30618 3932
rect 30634 3868 30698 3932
rect 30714 3868 30778 3932
rect 30794 3868 30858 3932
rect 30874 3868 30938 3932
rect 30954 3868 31018 3932
rect 31160 3868 31224 3932
rect 31240 3868 31304 3932
rect 31320 3868 31384 3932
rect 31400 3868 31464 3932
rect 31480 3868 31544 3932
rect 31560 3868 31624 3932
rect 31766 3868 31830 3932
rect 31846 3868 31910 3932
rect 31926 3868 31990 3932
rect 32006 3868 32070 3932
rect 32086 3868 32150 3932
rect 32166 3868 32230 3932
rect 32372 3868 32436 3932
rect 32452 3868 32516 3932
rect 32532 3868 32596 3932
rect 32612 3868 32676 3932
rect 32692 3868 32756 3932
rect 32772 3868 32836 3932
rect 32978 3868 33042 3932
rect 33058 3868 33122 3932
rect 33138 3868 33202 3932
rect 33218 3868 33282 3932
rect 33298 3868 33362 3932
rect 33378 3868 33442 3932
rect 33584 3868 33648 3932
rect 33664 3868 33728 3932
rect 33744 3868 33808 3932
rect 33824 3868 33888 3932
rect 33904 3868 33968 3932
rect 33984 3868 34048 3932
rect 34190 3868 34254 3932
rect 34270 3868 34334 3932
rect 34350 3868 34414 3932
rect 34430 3868 34494 3932
rect 34510 3868 34574 3932
rect 34590 3868 34654 3932
rect 34796 3868 34860 3932
rect 34876 3868 34940 3932
rect 34956 3868 35020 3932
rect 35036 3868 35100 3932
rect 35116 3868 35180 3932
rect 35196 3868 35260 3932
rect 35402 3868 35466 3932
rect 35482 3868 35546 3932
rect 35562 3868 35626 3932
rect 35642 3868 35706 3932
rect 35722 3868 35786 3932
rect 35802 3868 35866 3932
rect 36008 3868 36072 3932
rect 36088 3868 36152 3932
rect 36168 3868 36232 3932
rect 36248 3868 36312 3932
rect 36328 3868 36392 3932
rect 36408 3868 36472 3932
rect 36614 3868 36678 3932
rect 36694 3868 36758 3932
rect 36774 3868 36838 3932
rect 36854 3868 36918 3932
rect 36934 3868 36998 3932
rect 37014 3868 37078 3932
rect 37220 3868 37284 3932
rect 37300 3868 37364 3932
rect 37380 3868 37444 3932
rect 37460 3868 37524 3932
rect 37540 3868 37604 3932
rect 37620 3868 37684 3932
rect 37826 3868 37890 3932
rect 37906 3868 37970 3932
rect 37986 3868 38050 3932
rect 38066 3868 38130 3932
rect 38146 3868 38210 3932
rect 38226 3868 38290 3932
rect 38432 3868 38496 3932
rect 38512 3868 38576 3932
rect 38592 3868 38656 3932
rect 38672 3868 38736 3932
rect 38752 3868 38816 3932
rect 38832 3868 38896 3932
rect 39038 3868 39102 3932
rect 39118 3868 39182 3932
rect 39198 3868 39262 3932
rect 39278 3868 39342 3932
rect 39358 3868 39422 3932
rect 39438 3868 39502 3932
rect 20149 3648 20213 3712
rect 20149 3568 20213 3632
rect 20149 3488 20213 3552
rect 20149 3408 20213 3472
rect 20149 3328 20213 3392
rect 20149 3248 20213 3312
rect 20149 3168 20213 3232
rect 20149 3088 20213 3152
rect 20149 3008 20213 3072
rect 20149 2928 20213 2992
rect 20755 3648 20819 3712
rect 20755 3568 20819 3632
rect 20755 3488 20819 3552
rect 20755 3408 20819 3472
rect 20755 3328 20819 3392
rect 20755 3248 20819 3312
rect 20755 3168 20819 3232
rect 20755 3088 20819 3152
rect 20755 3008 20819 3072
rect 20755 2928 20819 2992
rect 21361 3648 21425 3712
rect 21361 3568 21425 3632
rect 21361 3488 21425 3552
rect 21361 3408 21425 3472
rect 21361 3328 21425 3392
rect 21361 3248 21425 3312
rect 21361 3168 21425 3232
rect 21361 3088 21425 3152
rect 21361 3008 21425 3072
rect 21361 2928 21425 2992
rect 21967 3648 22031 3712
rect 21967 3568 22031 3632
rect 21967 3488 22031 3552
rect 21967 3408 22031 3472
rect 21967 3328 22031 3392
rect 21967 3248 22031 3312
rect 21967 3168 22031 3232
rect 21967 3088 22031 3152
rect 21967 3008 22031 3072
rect 21967 2928 22031 2992
rect 22573 3648 22637 3712
rect 22573 3568 22637 3632
rect 22573 3488 22637 3552
rect 22573 3408 22637 3472
rect 22573 3328 22637 3392
rect 22573 3248 22637 3312
rect 22573 3168 22637 3232
rect 22573 3088 22637 3152
rect 22573 3008 22637 3072
rect 22573 2928 22637 2992
rect 23179 3648 23243 3712
rect 23179 3568 23243 3632
rect 23179 3488 23243 3552
rect 23179 3408 23243 3472
rect 23179 3328 23243 3392
rect 23179 3248 23243 3312
rect 23179 3168 23243 3232
rect 23179 3088 23243 3152
rect 23179 3008 23243 3072
rect 23179 2928 23243 2992
rect 23785 3648 23849 3712
rect 23785 3568 23849 3632
rect 23785 3488 23849 3552
rect 23785 3408 23849 3472
rect 23785 3328 23849 3392
rect 23785 3248 23849 3312
rect 23785 3168 23849 3232
rect 23785 3088 23849 3152
rect 23785 3008 23849 3072
rect 23785 2928 23849 2992
rect 24391 3648 24455 3712
rect 24391 3568 24455 3632
rect 24391 3488 24455 3552
rect 24391 3408 24455 3472
rect 24391 3328 24455 3392
rect 24391 3248 24455 3312
rect 24391 3168 24455 3232
rect 24391 3088 24455 3152
rect 24391 3008 24455 3072
rect 24391 2928 24455 2992
rect 24997 3648 25061 3712
rect 24997 3568 25061 3632
rect 24997 3488 25061 3552
rect 24997 3408 25061 3472
rect 24997 3328 25061 3392
rect 24997 3248 25061 3312
rect 24997 3168 25061 3232
rect 24997 3088 25061 3152
rect 24997 3008 25061 3072
rect 24997 2928 25061 2992
rect 25603 3648 25667 3712
rect 25603 3568 25667 3632
rect 25603 3488 25667 3552
rect 25603 3408 25667 3472
rect 25603 3328 25667 3392
rect 25603 3248 25667 3312
rect 25603 3168 25667 3232
rect 25603 3088 25667 3152
rect 25603 3008 25667 3072
rect 25603 2928 25667 2992
rect 26209 3648 26273 3712
rect 26209 3568 26273 3632
rect 26209 3488 26273 3552
rect 26209 3408 26273 3472
rect 26209 3328 26273 3392
rect 26209 3248 26273 3312
rect 26209 3168 26273 3232
rect 26209 3088 26273 3152
rect 26209 3008 26273 3072
rect 26209 2928 26273 2992
rect 26815 3648 26879 3712
rect 26815 3568 26879 3632
rect 26815 3488 26879 3552
rect 26815 3408 26879 3472
rect 26815 3328 26879 3392
rect 26815 3248 26879 3312
rect 26815 3168 26879 3232
rect 26815 3088 26879 3152
rect 26815 3008 26879 3072
rect 26815 2928 26879 2992
rect 27421 3648 27485 3712
rect 27421 3568 27485 3632
rect 27421 3488 27485 3552
rect 27421 3408 27485 3472
rect 27421 3328 27485 3392
rect 27421 3248 27485 3312
rect 27421 3168 27485 3232
rect 27421 3088 27485 3152
rect 27421 3008 27485 3072
rect 27421 2928 27485 2992
rect 28027 3648 28091 3712
rect 28027 3568 28091 3632
rect 28027 3488 28091 3552
rect 28027 3408 28091 3472
rect 28027 3328 28091 3392
rect 28027 3248 28091 3312
rect 28027 3168 28091 3232
rect 28027 3088 28091 3152
rect 28027 3008 28091 3072
rect 28027 2928 28091 2992
rect 28633 3648 28697 3712
rect 28633 3568 28697 3632
rect 28633 3488 28697 3552
rect 28633 3408 28697 3472
rect 28633 3328 28697 3392
rect 28633 3248 28697 3312
rect 28633 3168 28697 3232
rect 28633 3088 28697 3152
rect 28633 3008 28697 3072
rect 28633 2928 28697 2992
rect 29239 3648 29303 3712
rect 29239 3568 29303 3632
rect 29239 3488 29303 3552
rect 29239 3408 29303 3472
rect 29239 3328 29303 3392
rect 29239 3248 29303 3312
rect 29239 3168 29303 3232
rect 29239 3088 29303 3152
rect 29239 3008 29303 3072
rect 29239 2928 29303 2992
rect 29845 3648 29909 3712
rect 29845 3568 29909 3632
rect 29845 3488 29909 3552
rect 29845 3408 29909 3472
rect 29845 3328 29909 3392
rect 29845 3248 29909 3312
rect 29845 3168 29909 3232
rect 29845 3088 29909 3152
rect 29845 3008 29909 3072
rect 29845 2928 29909 2992
rect 30451 3648 30515 3712
rect 30451 3568 30515 3632
rect 30451 3488 30515 3552
rect 30451 3408 30515 3472
rect 30451 3328 30515 3392
rect 30451 3248 30515 3312
rect 30451 3168 30515 3232
rect 30451 3088 30515 3152
rect 30451 3008 30515 3072
rect 30451 2928 30515 2992
rect 31057 3648 31121 3712
rect 31057 3568 31121 3632
rect 31057 3488 31121 3552
rect 31057 3408 31121 3472
rect 31057 3328 31121 3392
rect 31057 3248 31121 3312
rect 31057 3168 31121 3232
rect 31057 3088 31121 3152
rect 31057 3008 31121 3072
rect 31057 2928 31121 2992
rect 31663 3648 31727 3712
rect 31663 3568 31727 3632
rect 31663 3488 31727 3552
rect 31663 3408 31727 3472
rect 31663 3328 31727 3392
rect 31663 3248 31727 3312
rect 31663 3168 31727 3232
rect 31663 3088 31727 3152
rect 31663 3008 31727 3072
rect 31663 2928 31727 2992
rect 32269 3648 32333 3712
rect 32269 3568 32333 3632
rect 32269 3488 32333 3552
rect 32269 3408 32333 3472
rect 32269 3328 32333 3392
rect 32269 3248 32333 3312
rect 32269 3168 32333 3232
rect 32269 3088 32333 3152
rect 32269 3008 32333 3072
rect 32269 2928 32333 2992
rect 32875 3648 32939 3712
rect 32875 3568 32939 3632
rect 32875 3488 32939 3552
rect 32875 3408 32939 3472
rect 32875 3328 32939 3392
rect 32875 3248 32939 3312
rect 32875 3168 32939 3232
rect 32875 3088 32939 3152
rect 32875 3008 32939 3072
rect 32875 2928 32939 2992
rect 33481 3648 33545 3712
rect 33481 3568 33545 3632
rect 33481 3488 33545 3552
rect 33481 3408 33545 3472
rect 33481 3328 33545 3392
rect 33481 3248 33545 3312
rect 33481 3168 33545 3232
rect 33481 3088 33545 3152
rect 33481 3008 33545 3072
rect 33481 2928 33545 2992
rect 34087 3648 34151 3712
rect 34087 3568 34151 3632
rect 34087 3488 34151 3552
rect 34087 3408 34151 3472
rect 34087 3328 34151 3392
rect 34087 3248 34151 3312
rect 34087 3168 34151 3232
rect 34087 3088 34151 3152
rect 34087 3008 34151 3072
rect 34087 2928 34151 2992
rect 34693 3648 34757 3712
rect 34693 3568 34757 3632
rect 34693 3488 34757 3552
rect 34693 3408 34757 3472
rect 34693 3328 34757 3392
rect 34693 3248 34757 3312
rect 34693 3168 34757 3232
rect 34693 3088 34757 3152
rect 34693 3008 34757 3072
rect 34693 2928 34757 2992
rect 35299 3648 35363 3712
rect 35299 3568 35363 3632
rect 35299 3488 35363 3552
rect 35299 3408 35363 3472
rect 35299 3328 35363 3392
rect 35299 3248 35363 3312
rect 35299 3168 35363 3232
rect 35299 3088 35363 3152
rect 35299 3008 35363 3072
rect 35299 2928 35363 2992
rect 35905 3648 35969 3712
rect 35905 3568 35969 3632
rect 35905 3488 35969 3552
rect 35905 3408 35969 3472
rect 35905 3328 35969 3392
rect 35905 3248 35969 3312
rect 35905 3168 35969 3232
rect 35905 3088 35969 3152
rect 35905 3008 35969 3072
rect 35905 2928 35969 2992
rect 36511 3648 36575 3712
rect 36511 3568 36575 3632
rect 36511 3488 36575 3552
rect 36511 3408 36575 3472
rect 36511 3328 36575 3392
rect 36511 3248 36575 3312
rect 36511 3168 36575 3232
rect 36511 3088 36575 3152
rect 36511 3008 36575 3072
rect 36511 2928 36575 2992
rect 37117 3648 37181 3712
rect 37117 3568 37181 3632
rect 37117 3488 37181 3552
rect 37117 3408 37181 3472
rect 37117 3328 37181 3392
rect 37117 3248 37181 3312
rect 37117 3168 37181 3232
rect 37117 3088 37181 3152
rect 37117 3008 37181 3072
rect 37117 2928 37181 2992
rect 37723 3648 37787 3712
rect 37723 3568 37787 3632
rect 37723 3488 37787 3552
rect 37723 3408 37787 3472
rect 37723 3328 37787 3392
rect 37723 3248 37787 3312
rect 37723 3168 37787 3232
rect 37723 3088 37787 3152
rect 37723 3008 37787 3072
rect 37723 2928 37787 2992
rect 38329 3648 38393 3712
rect 38329 3568 38393 3632
rect 38329 3488 38393 3552
rect 38329 3408 38393 3472
rect 38329 3328 38393 3392
rect 38329 3248 38393 3312
rect 38329 3168 38393 3232
rect 38329 3088 38393 3152
rect 38329 3008 38393 3072
rect 38329 2928 38393 2992
rect 38935 3648 38999 3712
rect 38935 3568 38999 3632
rect 38935 3488 38999 3552
rect 38935 3408 38999 3472
rect 38935 3328 38999 3392
rect 38935 3248 38999 3312
rect 38935 3168 38999 3232
rect 38935 3088 38999 3152
rect 38935 3008 38999 3072
rect 38935 2928 38999 2992
rect 39541 3648 39605 3712
rect 39541 3568 39605 3632
rect 39541 3488 39605 3552
rect 39541 3408 39605 3472
rect 39541 3328 39605 3392
rect 39541 3248 39605 3312
rect 39541 3168 39605 3232
rect 39541 3088 39605 3152
rect 39541 3008 39605 3072
rect 39541 2928 39605 2992
rect -355 2708 -291 2772
rect -275 2708 -211 2772
rect -195 2708 -131 2772
rect -115 2708 -51 2772
rect -35 2708 29 2772
rect 45 2708 109 2772
rect 459 2708 523 2772
rect 539 2708 603 2772
rect 619 2708 683 2772
rect 699 2708 763 2772
rect 779 2708 843 2772
rect 859 2708 923 2772
rect 1371 2708 1435 2772
rect 1451 2708 1515 2772
rect 1531 2708 1595 2772
rect 1611 2708 1675 2772
rect 1691 2708 1755 2772
rect 1771 2708 1835 2772
rect 1977 2708 2041 2772
rect 2057 2708 2121 2772
rect 2137 2708 2201 2772
rect 2217 2708 2281 2772
rect 2297 2708 2361 2772
rect 2377 2708 2441 2772
rect 2905 2708 2969 2772
rect 2985 2708 3049 2772
rect 3065 2708 3129 2772
rect 3145 2708 3209 2772
rect 3225 2708 3289 2772
rect 3305 2708 3369 2772
rect 3511 2708 3575 2772
rect 3591 2708 3655 2772
rect 3671 2708 3735 2772
rect 3751 2708 3815 2772
rect 3831 2708 3895 2772
rect 3911 2708 3975 2772
rect 4117 2708 4181 2772
rect 4197 2708 4261 2772
rect 4277 2708 4341 2772
rect 4357 2708 4421 2772
rect 4437 2708 4501 2772
rect 4517 2708 4581 2772
rect 4723 2708 4787 2772
rect 4803 2708 4867 2772
rect 4883 2708 4947 2772
rect 4963 2708 5027 2772
rect 5043 2708 5107 2772
rect 5123 2708 5187 2772
rect 5456 2708 5520 2772
rect 5536 2708 5600 2772
rect 5616 2708 5680 2772
rect 5696 2708 5760 2772
rect 5776 2708 5840 2772
rect 5856 2708 5920 2772
rect 6062 2708 6126 2772
rect 6142 2708 6206 2772
rect 6222 2708 6286 2772
rect 6302 2708 6366 2772
rect 6382 2708 6446 2772
rect 6462 2708 6526 2772
rect 6668 2708 6732 2772
rect 6748 2708 6812 2772
rect 6828 2708 6892 2772
rect 6908 2708 6972 2772
rect 6988 2708 7052 2772
rect 7068 2708 7132 2772
rect 7274 2708 7338 2772
rect 7354 2708 7418 2772
rect 7434 2708 7498 2772
rect 7514 2708 7578 2772
rect 7594 2708 7658 2772
rect 7674 2708 7738 2772
rect 7880 2708 7944 2772
rect 7960 2708 8024 2772
rect 8040 2708 8104 2772
rect 8120 2708 8184 2772
rect 8200 2708 8264 2772
rect 8280 2708 8344 2772
rect 8486 2708 8550 2772
rect 8566 2708 8630 2772
rect 8646 2708 8710 2772
rect 8726 2708 8790 2772
rect 8806 2708 8870 2772
rect 8886 2708 8950 2772
rect 9092 2708 9156 2772
rect 9172 2708 9236 2772
rect 9252 2708 9316 2772
rect 9332 2708 9396 2772
rect 9412 2708 9476 2772
rect 9492 2708 9556 2772
rect 9698 2708 9762 2772
rect 9778 2708 9842 2772
rect 9858 2708 9922 2772
rect 9938 2708 10002 2772
rect 10018 2708 10082 2772
rect 10098 2708 10162 2772
rect 10430 2708 10494 2772
rect 10510 2708 10574 2772
rect 10590 2708 10654 2772
rect 10670 2708 10734 2772
rect 10750 2708 10814 2772
rect 10830 2708 10894 2772
rect 11036 2708 11100 2772
rect 11116 2708 11180 2772
rect 11196 2708 11260 2772
rect 11276 2708 11340 2772
rect 11356 2708 11420 2772
rect 11436 2708 11500 2772
rect 11642 2708 11706 2772
rect 11722 2708 11786 2772
rect 11802 2708 11866 2772
rect 11882 2708 11946 2772
rect 11962 2708 12026 2772
rect 12042 2708 12106 2772
rect 12248 2708 12312 2772
rect 12328 2708 12392 2772
rect 12408 2708 12472 2772
rect 12488 2708 12552 2772
rect 12568 2708 12632 2772
rect 12648 2708 12712 2772
rect 12854 2708 12918 2772
rect 12934 2708 12998 2772
rect 13014 2708 13078 2772
rect 13094 2708 13158 2772
rect 13174 2708 13238 2772
rect 13254 2708 13318 2772
rect 13460 2708 13524 2772
rect 13540 2708 13604 2772
rect 13620 2708 13684 2772
rect 13700 2708 13764 2772
rect 13780 2708 13844 2772
rect 13860 2708 13924 2772
rect 14066 2708 14130 2772
rect 14146 2708 14210 2772
rect 14226 2708 14290 2772
rect 14306 2708 14370 2772
rect 14386 2708 14450 2772
rect 14466 2708 14530 2772
rect 14672 2708 14736 2772
rect 14752 2708 14816 2772
rect 14832 2708 14896 2772
rect 14912 2708 14976 2772
rect 14992 2708 15056 2772
rect 15072 2708 15136 2772
rect 15278 2708 15342 2772
rect 15358 2708 15422 2772
rect 15438 2708 15502 2772
rect 15518 2708 15582 2772
rect 15598 2708 15662 2772
rect 15678 2708 15742 2772
rect 15884 2708 15948 2772
rect 15964 2708 16028 2772
rect 16044 2708 16108 2772
rect 16124 2708 16188 2772
rect 16204 2708 16268 2772
rect 16284 2708 16348 2772
rect 16490 2708 16554 2772
rect 16570 2708 16634 2772
rect 16650 2708 16714 2772
rect 16730 2708 16794 2772
rect 16810 2708 16874 2772
rect 16890 2708 16954 2772
rect 17096 2708 17160 2772
rect 17176 2708 17240 2772
rect 17256 2708 17320 2772
rect 17336 2708 17400 2772
rect 17416 2708 17480 2772
rect 17496 2708 17560 2772
rect 17702 2708 17766 2772
rect 17782 2708 17846 2772
rect 17862 2708 17926 2772
rect 17942 2708 18006 2772
rect 18022 2708 18086 2772
rect 18102 2708 18166 2772
rect 18308 2708 18372 2772
rect 18388 2708 18452 2772
rect 18468 2708 18532 2772
rect 18548 2708 18612 2772
rect 18628 2708 18692 2772
rect 18708 2708 18772 2772
rect 18914 2708 18978 2772
rect 18994 2708 19058 2772
rect 19074 2708 19138 2772
rect 19154 2708 19218 2772
rect 19234 2708 19298 2772
rect 19314 2708 19378 2772
rect 19520 2708 19584 2772
rect 19600 2708 19664 2772
rect 19680 2708 19744 2772
rect 19760 2708 19824 2772
rect 19840 2708 19904 2772
rect 19920 2708 19984 2772
rect 20252 2708 20316 2772
rect 20332 2708 20396 2772
rect 20412 2708 20476 2772
rect 20492 2708 20556 2772
rect 20572 2708 20636 2772
rect 20652 2708 20716 2772
rect 20858 2708 20922 2772
rect 20938 2708 21002 2772
rect 21018 2708 21082 2772
rect 21098 2708 21162 2772
rect 21178 2708 21242 2772
rect 21258 2708 21322 2772
rect 21464 2708 21528 2772
rect 21544 2708 21608 2772
rect 21624 2708 21688 2772
rect 21704 2708 21768 2772
rect 21784 2708 21848 2772
rect 21864 2708 21928 2772
rect 22070 2708 22134 2772
rect 22150 2708 22214 2772
rect 22230 2708 22294 2772
rect 22310 2708 22374 2772
rect 22390 2708 22454 2772
rect 22470 2708 22534 2772
rect 22676 2708 22740 2772
rect 22756 2708 22820 2772
rect 22836 2708 22900 2772
rect 22916 2708 22980 2772
rect 22996 2708 23060 2772
rect 23076 2708 23140 2772
rect 23282 2708 23346 2772
rect 23362 2708 23426 2772
rect 23442 2708 23506 2772
rect 23522 2708 23586 2772
rect 23602 2708 23666 2772
rect 23682 2708 23746 2772
rect 23888 2708 23952 2772
rect 23968 2708 24032 2772
rect 24048 2708 24112 2772
rect 24128 2708 24192 2772
rect 24208 2708 24272 2772
rect 24288 2708 24352 2772
rect 24494 2708 24558 2772
rect 24574 2708 24638 2772
rect 24654 2708 24718 2772
rect 24734 2708 24798 2772
rect 24814 2708 24878 2772
rect 24894 2708 24958 2772
rect 25100 2708 25164 2772
rect 25180 2708 25244 2772
rect 25260 2708 25324 2772
rect 25340 2708 25404 2772
rect 25420 2708 25484 2772
rect 25500 2708 25564 2772
rect 25706 2708 25770 2772
rect 25786 2708 25850 2772
rect 25866 2708 25930 2772
rect 25946 2708 26010 2772
rect 26026 2708 26090 2772
rect 26106 2708 26170 2772
rect 26312 2708 26376 2772
rect 26392 2708 26456 2772
rect 26472 2708 26536 2772
rect 26552 2708 26616 2772
rect 26632 2708 26696 2772
rect 26712 2708 26776 2772
rect 26918 2708 26982 2772
rect 26998 2708 27062 2772
rect 27078 2708 27142 2772
rect 27158 2708 27222 2772
rect 27238 2708 27302 2772
rect 27318 2708 27382 2772
rect 27524 2708 27588 2772
rect 27604 2708 27668 2772
rect 27684 2708 27748 2772
rect 27764 2708 27828 2772
rect 27844 2708 27908 2772
rect 27924 2708 27988 2772
rect 28130 2708 28194 2772
rect 28210 2708 28274 2772
rect 28290 2708 28354 2772
rect 28370 2708 28434 2772
rect 28450 2708 28514 2772
rect 28530 2708 28594 2772
rect 28736 2708 28800 2772
rect 28816 2708 28880 2772
rect 28896 2708 28960 2772
rect 28976 2708 29040 2772
rect 29056 2708 29120 2772
rect 29136 2708 29200 2772
rect 29342 2708 29406 2772
rect 29422 2708 29486 2772
rect 29502 2708 29566 2772
rect 29582 2708 29646 2772
rect 29662 2708 29726 2772
rect 29742 2708 29806 2772
rect 29948 2708 30012 2772
rect 30028 2708 30092 2772
rect 30108 2708 30172 2772
rect 30188 2708 30252 2772
rect 30268 2708 30332 2772
rect 30348 2708 30412 2772
rect 30554 2708 30618 2772
rect 30634 2708 30698 2772
rect 30714 2708 30778 2772
rect 30794 2708 30858 2772
rect 30874 2708 30938 2772
rect 30954 2708 31018 2772
rect 31160 2708 31224 2772
rect 31240 2708 31304 2772
rect 31320 2708 31384 2772
rect 31400 2708 31464 2772
rect 31480 2708 31544 2772
rect 31560 2708 31624 2772
rect 31766 2708 31830 2772
rect 31846 2708 31910 2772
rect 31926 2708 31990 2772
rect 32006 2708 32070 2772
rect 32086 2708 32150 2772
rect 32166 2708 32230 2772
rect 32372 2708 32436 2772
rect 32452 2708 32516 2772
rect 32532 2708 32596 2772
rect 32612 2708 32676 2772
rect 32692 2708 32756 2772
rect 32772 2708 32836 2772
rect 32978 2708 33042 2772
rect 33058 2708 33122 2772
rect 33138 2708 33202 2772
rect 33218 2708 33282 2772
rect 33298 2708 33362 2772
rect 33378 2708 33442 2772
rect 33584 2708 33648 2772
rect 33664 2708 33728 2772
rect 33744 2708 33808 2772
rect 33824 2708 33888 2772
rect 33904 2708 33968 2772
rect 33984 2708 34048 2772
rect 34190 2708 34254 2772
rect 34270 2708 34334 2772
rect 34350 2708 34414 2772
rect 34430 2708 34494 2772
rect 34510 2708 34574 2772
rect 34590 2708 34654 2772
rect 34796 2708 34860 2772
rect 34876 2708 34940 2772
rect 34956 2708 35020 2772
rect 35036 2708 35100 2772
rect 35116 2708 35180 2772
rect 35196 2708 35260 2772
rect 35402 2708 35466 2772
rect 35482 2708 35546 2772
rect 35562 2708 35626 2772
rect 35642 2708 35706 2772
rect 35722 2708 35786 2772
rect 35802 2708 35866 2772
rect 36008 2708 36072 2772
rect 36088 2708 36152 2772
rect 36168 2708 36232 2772
rect 36248 2708 36312 2772
rect 36328 2708 36392 2772
rect 36408 2708 36472 2772
rect 36614 2708 36678 2772
rect 36694 2708 36758 2772
rect 36774 2708 36838 2772
rect 36854 2708 36918 2772
rect 36934 2708 36998 2772
rect 37014 2708 37078 2772
rect 37220 2708 37284 2772
rect 37300 2708 37364 2772
rect 37380 2708 37444 2772
rect 37460 2708 37524 2772
rect 37540 2708 37604 2772
rect 37620 2708 37684 2772
rect 37826 2708 37890 2772
rect 37906 2708 37970 2772
rect 37986 2708 38050 2772
rect 38066 2708 38130 2772
rect 38146 2708 38210 2772
rect 38226 2708 38290 2772
rect 38432 2708 38496 2772
rect 38512 2708 38576 2772
rect 38592 2708 38656 2772
rect 38672 2708 38736 2772
rect 38752 2708 38816 2772
rect 38832 2708 38896 2772
rect 39038 2708 39102 2772
rect 39118 2708 39182 2772
rect 39198 2708 39262 2772
rect 39278 2708 39342 2772
rect 39358 2708 39422 2772
rect 39438 2708 39502 2772
rect -355 1895 -291 1959
rect -275 1895 -211 1959
rect -195 1895 -131 1959
rect -115 1956 -51 1959
rect -115 1900 -91 1956
rect -91 1900 -51 1956
rect -115 1895 -51 1900
rect -35 1895 29 1959
rect 45 1895 109 1959
rect 459 1895 523 1959
rect 539 1895 603 1959
rect 619 1895 683 1959
rect 699 1895 763 1959
rect 779 1895 843 1959
rect 859 1895 923 1959
rect 1371 1895 1435 1959
rect 1451 1895 1515 1959
rect 1531 1895 1595 1959
rect 1611 1895 1675 1959
rect 1691 1895 1755 1959
rect 1771 1895 1835 1959
rect 1977 1895 2041 1959
rect 2057 1895 2121 1959
rect 2137 1895 2201 1959
rect 2217 1895 2281 1959
rect 2297 1895 2361 1959
rect 2377 1895 2441 1959
rect 2905 1895 2969 1959
rect 2985 1895 3049 1959
rect 3065 1895 3129 1959
rect 3145 1895 3209 1959
rect 3225 1895 3289 1959
rect 3305 1895 3369 1959
rect 3511 1895 3575 1959
rect 3591 1895 3655 1959
rect 3671 1895 3735 1959
rect 3751 1895 3815 1959
rect 3831 1895 3895 1959
rect 3911 1895 3975 1959
rect 4117 1895 4181 1959
rect 4197 1895 4261 1959
rect 4277 1895 4341 1959
rect 4357 1895 4421 1959
rect 4437 1895 4501 1959
rect 4517 1895 4581 1959
rect 4723 1895 4787 1959
rect 4803 1895 4867 1959
rect 4883 1895 4947 1959
rect 4963 1895 5027 1959
rect 5043 1895 5107 1959
rect 5123 1895 5187 1959
rect 5456 1895 5520 1959
rect 5536 1895 5600 1959
rect 5616 1895 5680 1959
rect 5696 1895 5760 1959
rect 5776 1895 5840 1959
rect 5856 1895 5920 1959
rect 6062 1895 6126 1959
rect 6142 1895 6206 1959
rect 6222 1895 6286 1959
rect 6302 1895 6366 1959
rect 6382 1895 6446 1959
rect 6462 1895 6526 1959
rect 6668 1895 6732 1959
rect 6748 1895 6812 1959
rect 6828 1895 6892 1959
rect 6908 1895 6972 1959
rect 6988 1895 7052 1959
rect 7068 1895 7132 1959
rect 7274 1895 7338 1959
rect 7354 1895 7418 1959
rect 7434 1895 7498 1959
rect 7514 1895 7578 1959
rect 7594 1895 7658 1959
rect 7674 1895 7738 1959
rect 7880 1895 7944 1959
rect 7960 1895 8024 1959
rect 8040 1895 8104 1959
rect 8120 1895 8184 1959
rect 8200 1895 8264 1959
rect 8280 1895 8344 1959
rect 8486 1895 8550 1959
rect 8566 1895 8630 1959
rect 8646 1895 8710 1959
rect 8726 1895 8790 1959
rect 8806 1895 8870 1959
rect 8886 1895 8950 1959
rect 9092 1895 9156 1959
rect 9172 1895 9236 1959
rect 9252 1895 9316 1959
rect 9332 1895 9396 1959
rect 9412 1895 9476 1959
rect 9492 1895 9556 1959
rect 9698 1895 9762 1959
rect 9778 1895 9842 1959
rect 9858 1895 9922 1959
rect 9938 1895 10002 1959
rect 10018 1895 10082 1959
rect 10098 1895 10162 1959
rect 10430 1895 10494 1959
rect 10510 1895 10574 1959
rect 10590 1895 10654 1959
rect 10670 1895 10734 1959
rect 10750 1895 10814 1959
rect 10830 1895 10894 1959
rect 11036 1895 11100 1959
rect 11116 1895 11180 1959
rect 11196 1895 11260 1959
rect 11276 1895 11340 1959
rect 11356 1895 11420 1959
rect 11436 1895 11500 1959
rect 11642 1895 11706 1959
rect 11722 1895 11786 1959
rect 11802 1895 11866 1959
rect 11882 1895 11946 1959
rect 11962 1895 12026 1959
rect 12042 1895 12106 1959
rect 12248 1895 12312 1959
rect 12328 1895 12392 1959
rect 12408 1895 12472 1959
rect 12488 1895 12552 1959
rect 12568 1895 12632 1959
rect 12648 1895 12712 1959
rect 12854 1895 12918 1959
rect 12934 1895 12998 1959
rect 13014 1895 13078 1959
rect 13094 1895 13158 1959
rect 13174 1895 13238 1959
rect 13254 1895 13318 1959
rect 13460 1895 13524 1959
rect 13540 1895 13604 1959
rect 13620 1895 13684 1959
rect 13700 1895 13764 1959
rect 13780 1895 13844 1959
rect 13860 1895 13924 1959
rect 14066 1895 14130 1959
rect 14146 1895 14210 1959
rect 14226 1895 14290 1959
rect 14306 1895 14370 1959
rect 14386 1895 14450 1959
rect 14466 1895 14530 1959
rect 14672 1895 14736 1959
rect 14752 1895 14816 1959
rect 14832 1895 14896 1959
rect 14912 1895 14976 1959
rect 14992 1895 15056 1959
rect 15072 1895 15136 1959
rect 15278 1895 15342 1959
rect 15358 1895 15422 1959
rect 15438 1895 15502 1959
rect 15518 1895 15582 1959
rect 15598 1895 15662 1959
rect 15678 1895 15742 1959
rect 15884 1895 15948 1959
rect 15964 1895 16028 1959
rect 16044 1895 16108 1959
rect 16124 1895 16188 1959
rect 16204 1895 16268 1959
rect 16284 1895 16348 1959
rect 16490 1895 16554 1959
rect 16570 1895 16634 1959
rect 16650 1895 16714 1959
rect 16730 1895 16794 1959
rect 16810 1895 16874 1959
rect 16890 1895 16954 1959
rect 17096 1895 17160 1959
rect 17176 1895 17240 1959
rect 17256 1895 17320 1959
rect 17336 1895 17400 1959
rect 17416 1895 17480 1959
rect 17496 1895 17560 1959
rect 17702 1895 17766 1959
rect 17782 1895 17846 1959
rect 17862 1895 17926 1959
rect 17942 1895 18006 1959
rect 18022 1895 18086 1959
rect 18102 1895 18166 1959
rect 18308 1895 18372 1959
rect 18388 1895 18452 1959
rect 18468 1895 18532 1959
rect 18548 1895 18612 1959
rect 18628 1895 18692 1959
rect 18708 1895 18772 1959
rect 18914 1895 18978 1959
rect 18994 1895 19058 1959
rect 19074 1895 19138 1959
rect 19154 1895 19218 1959
rect 19234 1895 19298 1959
rect 19314 1895 19378 1959
rect 19520 1895 19584 1959
rect 19600 1895 19664 1959
rect 19680 1895 19744 1959
rect 19760 1895 19824 1959
rect 19840 1895 19904 1959
rect 19920 1895 19984 1959
rect 20252 1895 20316 1959
rect 20332 1895 20396 1959
rect 20412 1895 20476 1959
rect 20492 1895 20556 1959
rect 20572 1895 20636 1959
rect 20652 1895 20716 1959
rect 20858 1895 20922 1959
rect 20938 1895 21002 1959
rect 21018 1895 21082 1959
rect 21098 1895 21162 1959
rect 21178 1895 21242 1959
rect 21258 1895 21322 1959
rect 21464 1895 21528 1959
rect 21544 1895 21608 1959
rect 21624 1895 21688 1959
rect 21704 1895 21768 1959
rect 21784 1895 21848 1959
rect 21864 1895 21928 1959
rect 22070 1895 22134 1959
rect 22150 1895 22214 1959
rect 22230 1895 22294 1959
rect 22310 1895 22374 1959
rect 22390 1895 22454 1959
rect 22470 1895 22534 1959
rect 22676 1895 22740 1959
rect 22756 1895 22820 1959
rect 22836 1895 22900 1959
rect 22916 1895 22980 1959
rect 22996 1895 23060 1959
rect 23076 1895 23140 1959
rect 23282 1895 23346 1959
rect 23362 1895 23426 1959
rect 23442 1895 23506 1959
rect 23522 1895 23586 1959
rect 23602 1895 23666 1959
rect 23682 1895 23746 1959
rect 23888 1895 23952 1959
rect 23968 1895 24032 1959
rect 24048 1895 24112 1959
rect 24128 1895 24192 1959
rect 24208 1895 24272 1959
rect 24288 1895 24352 1959
rect 24494 1895 24558 1959
rect 24574 1895 24638 1959
rect 24654 1895 24718 1959
rect 24734 1895 24798 1959
rect 24814 1895 24878 1959
rect 24894 1895 24958 1959
rect 25100 1895 25164 1959
rect 25180 1895 25244 1959
rect 25260 1895 25324 1959
rect 25340 1895 25404 1959
rect 25420 1895 25484 1959
rect 25500 1895 25564 1959
rect 25706 1895 25770 1959
rect 25786 1895 25850 1959
rect 25866 1895 25930 1959
rect 25946 1895 26010 1959
rect 26026 1895 26090 1959
rect 26106 1895 26170 1959
rect 26312 1895 26376 1959
rect 26392 1895 26456 1959
rect 26472 1895 26536 1959
rect 26552 1895 26616 1959
rect 26632 1895 26696 1959
rect 26712 1895 26776 1959
rect 26918 1895 26982 1959
rect 26998 1895 27062 1959
rect 27078 1895 27142 1959
rect 27158 1895 27222 1959
rect 27238 1895 27302 1959
rect 27318 1895 27382 1959
rect 27524 1895 27588 1959
rect 27604 1895 27668 1959
rect 27684 1895 27748 1959
rect 27764 1895 27828 1959
rect 27844 1895 27908 1959
rect 27924 1895 27988 1959
rect 28130 1895 28194 1959
rect 28210 1895 28274 1959
rect 28290 1895 28354 1959
rect 28370 1895 28434 1959
rect 28450 1895 28514 1959
rect 28530 1895 28594 1959
rect 28736 1895 28800 1959
rect 28816 1895 28880 1959
rect 28896 1895 28960 1959
rect 28976 1895 29040 1959
rect 29056 1895 29120 1959
rect 29136 1895 29200 1959
rect 29342 1895 29406 1959
rect 29422 1895 29486 1959
rect 29502 1895 29566 1959
rect 29582 1895 29646 1959
rect 29662 1895 29726 1959
rect 29742 1895 29806 1959
rect 29948 1895 30012 1959
rect 30028 1895 30092 1959
rect 30108 1895 30172 1959
rect 30188 1895 30252 1959
rect 30268 1895 30332 1959
rect 30348 1895 30412 1959
rect 30554 1895 30618 1959
rect 30634 1895 30698 1959
rect 30714 1895 30778 1959
rect 30794 1895 30858 1959
rect 30874 1895 30938 1959
rect 30954 1895 31018 1959
rect 31160 1895 31224 1959
rect 31240 1895 31304 1959
rect 31320 1895 31384 1959
rect 31400 1895 31464 1959
rect 31480 1895 31544 1959
rect 31560 1895 31624 1959
rect 31766 1895 31830 1959
rect 31846 1895 31910 1959
rect 31926 1895 31990 1959
rect 32006 1895 32070 1959
rect 32086 1895 32150 1959
rect 32166 1895 32230 1959
rect 32372 1895 32436 1959
rect 32452 1895 32516 1959
rect 32532 1895 32596 1959
rect 32612 1895 32676 1959
rect 32692 1895 32756 1959
rect 32772 1895 32836 1959
rect 32978 1895 33042 1959
rect 33058 1895 33122 1959
rect 33138 1895 33202 1959
rect 33218 1895 33282 1959
rect 33298 1895 33362 1959
rect 33378 1895 33442 1959
rect 33584 1895 33648 1959
rect 33664 1895 33728 1959
rect 33744 1895 33808 1959
rect 33824 1895 33888 1959
rect 33904 1895 33968 1959
rect 33984 1895 34048 1959
rect 34190 1895 34254 1959
rect 34270 1895 34334 1959
rect 34350 1895 34414 1959
rect 34430 1895 34494 1959
rect 34510 1895 34574 1959
rect 34590 1895 34654 1959
rect 34796 1895 34860 1959
rect 34876 1895 34940 1959
rect 34956 1895 35020 1959
rect 35036 1895 35100 1959
rect 35116 1895 35180 1959
rect 35196 1895 35260 1959
rect 35402 1895 35466 1959
rect 35482 1895 35546 1959
rect 35562 1895 35626 1959
rect 35642 1895 35706 1959
rect 35722 1895 35786 1959
rect 35802 1895 35866 1959
rect 36008 1895 36072 1959
rect 36088 1895 36152 1959
rect 36168 1895 36232 1959
rect 36248 1895 36312 1959
rect 36328 1895 36392 1959
rect 36408 1895 36472 1959
rect 36614 1895 36678 1959
rect 36694 1895 36758 1959
rect 36774 1895 36838 1959
rect 36854 1895 36918 1959
rect 36934 1895 36998 1959
rect 37014 1895 37078 1959
rect 37220 1895 37284 1959
rect 37300 1895 37364 1959
rect 37380 1895 37444 1959
rect 37460 1895 37524 1959
rect 37540 1895 37604 1959
rect 37620 1895 37684 1959
rect 37826 1895 37890 1959
rect 37906 1895 37970 1959
rect 37986 1895 38050 1959
rect 38066 1895 38130 1959
rect 38146 1895 38210 1959
rect 38226 1895 38290 1959
rect 38432 1895 38496 1959
rect 38512 1895 38576 1959
rect 38592 1895 38656 1959
rect 38672 1895 38736 1959
rect 38752 1895 38816 1959
rect 38832 1895 38896 1959
rect 39038 1895 39102 1959
rect 39118 1895 39182 1959
rect 39198 1895 39262 1959
rect 39278 1895 39342 1959
rect 39358 1895 39422 1959
rect 39438 1895 39502 1959
rect -458 1675 -394 1739
rect -458 1595 -394 1659
rect -458 1515 -394 1579
rect -458 1435 -394 1499
rect -458 1355 -394 1419
rect -458 1275 -394 1339
rect -458 1195 -394 1259
rect -458 1115 -394 1179
rect -458 1035 -394 1099
rect -458 955 -394 1019
rect 148 1675 212 1739
rect 148 1595 212 1659
rect 148 1515 212 1579
rect 148 1435 212 1499
rect 148 1355 212 1419
rect 148 1275 212 1339
rect 148 1195 212 1259
rect 148 1115 212 1179
rect 148 1035 212 1099
rect 148 955 212 1019
rect 356 1675 420 1739
rect 356 1595 420 1659
rect 356 1515 420 1579
rect 356 1435 420 1499
rect 356 1355 420 1419
rect 356 1275 420 1339
rect 356 1195 420 1259
rect 356 1115 420 1179
rect 356 1035 420 1099
rect 356 955 420 1019
rect 962 1817 1026 1821
rect 962 1761 966 1817
rect 966 1761 1022 1817
rect 1022 1761 1026 1817
rect 962 1757 1026 1761
rect 962 1675 1026 1739
rect 962 1615 966 1659
rect 966 1615 1022 1659
rect 1022 1615 1026 1659
rect 962 1595 1026 1615
rect 962 1515 1026 1579
rect 962 1435 1026 1499
rect 962 1355 1026 1419
rect 962 1275 1026 1339
rect 962 1195 1026 1259
rect 962 1115 1026 1179
rect 962 1035 1026 1099
rect 962 955 1026 1019
rect -355 735 -291 799
rect -275 735 -211 799
rect -195 735 -131 799
rect -115 735 -51 799
rect -35 735 29 799
rect 45 735 109 799
rect 459 735 523 799
rect 539 735 603 799
rect 619 735 683 799
rect 699 735 763 799
rect 779 735 843 799
rect 859 735 923 799
rect -458 515 -394 579
rect -458 435 -394 499
rect -458 355 -394 419
rect -458 275 -394 339
rect -458 195 -394 259
rect -458 115 -394 179
rect -458 35 -394 99
rect -458 -45 -394 19
rect -458 -125 -394 -61
rect -458 -205 -394 -141
rect 148 515 212 579
rect 148 435 212 499
rect 148 355 212 419
rect 148 275 212 339
rect 148 195 212 259
rect 148 115 212 179
rect 148 35 212 99
rect 148 -45 212 19
rect 148 -125 212 -61
rect 148 -205 212 -141
rect 356 515 420 579
rect 356 435 420 499
rect 356 355 420 419
rect 356 275 420 339
rect 356 195 420 259
rect 356 115 420 179
rect 356 35 420 99
rect 356 -45 420 19
rect 356 -125 420 -61
rect 356 -205 420 -141
rect 962 515 1026 579
rect 962 435 1026 499
rect 962 355 1026 419
rect 962 275 1026 339
rect 962 195 1026 259
rect 962 115 1026 179
rect 962 35 1026 99
rect 962 -45 1026 19
rect 962 -125 1026 -61
rect 962 -205 1026 -141
rect 1268 1675 1332 1739
rect 1268 1595 1332 1659
rect 1268 1515 1332 1579
rect 1268 1435 1332 1499
rect 1268 1355 1332 1419
rect 1268 1275 1332 1339
rect 1268 1195 1332 1259
rect 1268 1115 1332 1179
rect 1268 1035 1332 1099
rect 1268 955 1332 1019
rect 1874 1816 1938 1820
rect 1874 1760 1878 1816
rect 1878 1760 1934 1816
rect 1934 1760 1938 1816
rect 1874 1756 1938 1760
rect 1874 1675 1938 1739
rect 1874 1595 1938 1659
rect 1874 1515 1938 1579
rect 1874 1435 1938 1499
rect 1874 1355 1938 1419
rect 1874 1275 1938 1339
rect 1874 1195 1938 1259
rect 1874 1115 1938 1179
rect 1874 1035 1938 1099
rect 1874 955 1938 1019
rect 2480 1817 2544 1821
rect 2480 1761 2484 1817
rect 2484 1761 2540 1817
rect 2540 1761 2544 1817
rect 2480 1757 2544 1761
rect 2480 1675 2544 1739
rect 2480 1595 2544 1659
rect 2480 1515 2544 1579
rect 2480 1435 2544 1499
rect 2480 1355 2544 1419
rect 2480 1275 2544 1339
rect 2480 1195 2544 1259
rect 2480 1115 2544 1179
rect 2480 1035 2544 1099
rect 2480 955 2544 1019
rect 1371 735 1435 799
rect 1451 735 1515 799
rect 1531 735 1595 799
rect 1611 735 1675 799
rect 1691 735 1755 799
rect 1771 735 1835 799
rect 1977 735 2041 799
rect 2057 735 2121 799
rect 2137 735 2201 799
rect 2217 735 2281 799
rect 2297 735 2361 799
rect 2377 735 2441 799
rect 1268 515 1332 579
rect 1268 435 1332 499
rect 1268 355 1332 419
rect 1268 275 1332 339
rect 1268 195 1332 259
rect 1268 115 1332 179
rect 1268 35 1332 99
rect 1268 -45 1332 19
rect 1268 -125 1332 -61
rect 1268 -205 1332 -141
rect 1874 515 1938 579
rect 1874 435 1938 499
rect 1874 355 1938 419
rect 1874 275 1938 339
rect 1874 195 1938 259
rect 1874 115 1938 179
rect 1874 35 1938 99
rect 1874 -45 1938 19
rect 1874 -125 1938 -61
rect 1874 -205 1938 -141
rect 2480 515 2544 579
rect 2480 435 2544 499
rect 2480 355 2544 419
rect 2480 275 2544 339
rect 2480 195 2544 259
rect 2480 115 2544 179
rect 2480 35 2544 99
rect 2480 -45 2544 19
rect 2480 -125 2544 -61
rect 2480 -205 2544 -141
rect 2802 1675 2866 1739
rect 2802 1595 2866 1659
rect 2802 1515 2866 1579
rect 2802 1435 2866 1499
rect 2802 1355 2866 1419
rect 2802 1275 2866 1339
rect 2802 1195 2866 1259
rect 2802 1115 2866 1179
rect 2802 1035 2866 1099
rect 2802 955 2866 1019
rect 3408 1675 3472 1739
rect 3408 1595 3472 1659
rect 3408 1515 3472 1579
rect 3408 1435 3472 1499
rect 3408 1355 3472 1419
rect 3408 1275 3472 1339
rect 3408 1195 3472 1259
rect 3408 1115 3472 1179
rect 3408 1035 3472 1099
rect 3408 955 3472 1019
rect 4014 1675 4078 1739
rect 4014 1595 4078 1659
rect 4014 1515 4078 1579
rect 4014 1435 4078 1499
rect 4014 1355 4078 1419
rect 4014 1275 4078 1339
rect 4014 1195 4078 1259
rect 4014 1115 4078 1179
rect 4014 1035 4078 1099
rect 4014 955 4078 1019
rect 4620 1675 4684 1739
rect 4620 1595 4684 1659
rect 4620 1515 4684 1579
rect 4620 1435 4684 1499
rect 4620 1355 4684 1419
rect 4620 1275 4684 1339
rect 4620 1195 4684 1259
rect 4620 1115 4684 1179
rect 4620 1035 4684 1099
rect 4620 955 4684 1019
rect 5226 1675 5290 1739
rect 5226 1595 5290 1659
rect 5226 1515 5290 1579
rect 5226 1435 5290 1499
rect 5226 1355 5290 1419
rect 5226 1275 5290 1339
rect 5226 1195 5290 1259
rect 5226 1115 5290 1179
rect 5226 1035 5290 1099
rect 5226 955 5290 1019
rect 2905 735 2969 799
rect 2985 735 3049 799
rect 3065 735 3129 799
rect 3145 735 3209 799
rect 3225 735 3289 799
rect 3305 735 3369 799
rect 3511 735 3575 799
rect 3591 735 3655 799
rect 3671 735 3735 799
rect 3751 735 3815 799
rect 3831 735 3895 799
rect 3911 735 3975 799
rect 4117 735 4181 799
rect 4197 735 4261 799
rect 4277 735 4341 799
rect 4357 735 4421 799
rect 4437 735 4501 799
rect 4517 735 4581 799
rect 4723 735 4787 799
rect 4803 735 4867 799
rect 4883 735 4947 799
rect 4963 735 5027 799
rect 5043 735 5107 799
rect 5123 735 5187 799
rect 2802 515 2866 579
rect 2802 435 2866 499
rect 2802 355 2866 419
rect 2802 275 2866 339
rect 2802 195 2866 259
rect 2802 115 2866 179
rect 2802 35 2866 99
rect 2802 -45 2866 19
rect 2802 -125 2866 -61
rect 2802 -205 2866 -141
rect 3408 515 3472 579
rect 3408 435 3472 499
rect 3408 355 3472 419
rect 3408 275 3472 339
rect 3408 195 3472 259
rect 3408 115 3472 179
rect 3408 35 3472 99
rect 3408 -45 3472 19
rect 3408 -125 3472 -61
rect 3408 -205 3472 -141
rect 4014 515 4078 579
rect 4014 435 4078 499
rect 4014 355 4078 419
rect 4014 275 4078 339
rect 4014 195 4078 259
rect 4014 115 4078 179
rect 4014 35 4078 99
rect 4014 -45 4078 19
rect 4014 -125 4078 -61
rect 4014 -205 4078 -141
rect 4620 515 4684 579
rect 4620 435 4684 499
rect 4620 355 4684 419
rect 4620 275 4684 339
rect 4620 195 4684 259
rect 4620 115 4684 179
rect 4620 35 4684 99
rect 4620 -45 4684 19
rect 4620 -125 4684 -61
rect 4620 -205 4684 -141
rect 5226 515 5290 579
rect 5226 435 5290 499
rect 5226 355 5290 419
rect 5226 275 5290 339
rect 5226 195 5290 259
rect 5226 115 5290 179
rect 5226 35 5290 99
rect 5226 -45 5290 19
rect 5226 -125 5290 -61
rect 5226 -205 5290 -141
rect 5353 1675 5417 1739
rect 5353 1595 5417 1659
rect 5353 1515 5417 1579
rect 5353 1435 5417 1499
rect 5353 1355 5417 1419
rect 5353 1275 5417 1339
rect 5353 1195 5417 1259
rect 5353 1115 5417 1179
rect 5353 1035 5417 1099
rect 5353 955 5417 1019
rect 5959 1675 6023 1739
rect 5959 1595 6023 1659
rect 5959 1515 6023 1579
rect 5959 1435 6023 1499
rect 5959 1355 6023 1419
rect 5959 1275 6023 1339
rect 5959 1195 6023 1259
rect 5959 1115 6023 1179
rect 5959 1035 6023 1099
rect 5959 955 6023 1019
rect 6565 1675 6629 1739
rect 6565 1595 6629 1659
rect 6565 1515 6629 1579
rect 6565 1435 6629 1499
rect 6565 1355 6629 1419
rect 6565 1275 6629 1339
rect 6565 1195 6629 1259
rect 6565 1115 6629 1179
rect 6565 1035 6629 1099
rect 6565 955 6629 1019
rect 7171 1675 7235 1739
rect 7171 1595 7235 1659
rect 7171 1515 7235 1579
rect 7171 1435 7235 1499
rect 7171 1355 7235 1419
rect 7171 1275 7235 1339
rect 7171 1195 7235 1259
rect 7171 1115 7235 1179
rect 7171 1035 7235 1099
rect 7171 955 7235 1019
rect 7777 1675 7841 1739
rect 7777 1595 7841 1659
rect 7777 1515 7841 1579
rect 7777 1435 7841 1499
rect 7777 1355 7841 1419
rect 7777 1275 7841 1339
rect 7777 1195 7841 1259
rect 7777 1115 7841 1179
rect 7777 1035 7841 1099
rect 7777 955 7841 1019
rect 8383 1675 8447 1739
rect 8383 1595 8447 1659
rect 8383 1515 8447 1579
rect 8383 1435 8447 1499
rect 8383 1355 8447 1419
rect 8383 1275 8447 1339
rect 8383 1195 8447 1259
rect 8383 1115 8447 1179
rect 8383 1035 8447 1099
rect 8383 955 8447 1019
rect 8989 1675 9053 1739
rect 8989 1595 9053 1659
rect 8989 1515 9053 1579
rect 8989 1435 9053 1499
rect 8989 1355 9053 1419
rect 8989 1275 9053 1339
rect 8989 1195 9053 1259
rect 8989 1115 9053 1179
rect 8989 1035 9053 1099
rect 8989 955 9053 1019
rect 9595 1675 9659 1739
rect 9595 1595 9659 1659
rect 9595 1515 9659 1579
rect 9595 1435 9659 1499
rect 9595 1355 9659 1419
rect 9595 1275 9659 1339
rect 9595 1195 9659 1259
rect 9595 1115 9659 1179
rect 9595 1035 9659 1099
rect 9595 955 9659 1019
rect 10201 1675 10265 1739
rect 10201 1595 10265 1659
rect 10201 1515 10265 1579
rect 10201 1435 10265 1499
rect 10201 1355 10265 1419
rect 10201 1275 10265 1339
rect 10201 1195 10265 1259
rect 10201 1115 10265 1179
rect 10201 1035 10265 1099
rect 10201 955 10265 1019
rect 5456 735 5520 799
rect 5536 735 5600 799
rect 5616 735 5680 799
rect 5696 735 5760 799
rect 5776 735 5840 799
rect 5856 735 5920 799
rect 6062 735 6126 799
rect 6142 735 6206 799
rect 6222 735 6286 799
rect 6302 735 6366 799
rect 6382 735 6446 799
rect 6462 735 6526 799
rect 6668 735 6732 799
rect 6748 735 6812 799
rect 6828 735 6892 799
rect 6908 735 6972 799
rect 6988 735 7052 799
rect 7068 735 7132 799
rect 7274 735 7338 799
rect 7354 735 7418 799
rect 7434 735 7498 799
rect 7514 735 7578 799
rect 7594 735 7658 799
rect 7674 735 7738 799
rect 7880 735 7944 799
rect 7960 735 8024 799
rect 8040 735 8104 799
rect 8120 735 8184 799
rect 8200 735 8264 799
rect 8280 735 8344 799
rect 8486 735 8550 799
rect 8566 735 8630 799
rect 8646 735 8710 799
rect 8726 735 8790 799
rect 8806 735 8870 799
rect 8886 735 8950 799
rect 9092 735 9156 799
rect 9172 735 9236 799
rect 9252 735 9316 799
rect 9332 735 9396 799
rect 9412 735 9476 799
rect 9492 735 9556 799
rect 9698 735 9762 799
rect 9778 735 9842 799
rect 9858 735 9922 799
rect 9938 735 10002 799
rect 10018 735 10082 799
rect 10098 735 10162 799
rect 5353 515 5417 579
rect 5353 435 5417 499
rect 5353 355 5417 419
rect 5353 275 5417 339
rect 5353 195 5417 259
rect 5353 115 5417 179
rect 5353 35 5417 99
rect 5353 -45 5417 19
rect 5353 -125 5417 -61
rect 5353 -205 5417 -141
rect 5959 515 6023 579
rect 5959 435 6023 499
rect 5959 355 6023 419
rect 5959 275 6023 339
rect 5959 195 6023 259
rect 5959 115 6023 179
rect 5959 35 6023 99
rect 5959 -45 6023 19
rect 5959 -125 6023 -61
rect 5959 -205 6023 -141
rect 6565 515 6629 579
rect 6565 435 6629 499
rect 6565 355 6629 419
rect 6565 275 6629 339
rect 6565 195 6629 259
rect 6565 115 6629 179
rect 6565 35 6629 99
rect 6565 -45 6629 19
rect 6565 -125 6629 -61
rect 6565 -205 6629 -141
rect 7171 515 7235 579
rect 7171 435 7235 499
rect 7171 355 7235 419
rect 7171 275 7235 339
rect 7171 195 7235 259
rect 7171 115 7235 179
rect 7171 35 7235 99
rect 7171 -45 7235 19
rect 7171 -125 7235 -61
rect 7171 -205 7235 -141
rect 7777 515 7841 579
rect 7777 435 7841 499
rect 7777 355 7841 419
rect 7777 275 7841 339
rect 7777 195 7841 259
rect 7777 115 7841 179
rect 7777 35 7841 99
rect 7777 -45 7841 19
rect 7777 -125 7841 -61
rect 7777 -205 7841 -141
rect 8383 515 8447 579
rect 8383 435 8447 499
rect 8383 355 8447 419
rect 8383 275 8447 339
rect 8383 195 8447 259
rect 8383 115 8447 179
rect 8383 35 8447 99
rect 8383 -45 8447 19
rect 8383 -125 8447 -61
rect 8383 -205 8447 -141
rect 8989 515 9053 579
rect 8989 435 9053 499
rect 8989 355 9053 419
rect 8989 275 9053 339
rect 8989 195 9053 259
rect 8989 115 9053 179
rect 8989 35 9053 99
rect 8989 -45 9053 19
rect 8989 -125 9053 -61
rect 8989 -205 9053 -141
rect 9595 515 9659 579
rect 9595 435 9659 499
rect 9595 355 9659 419
rect 9595 275 9659 339
rect 9595 195 9659 259
rect 9595 115 9659 179
rect 9595 35 9659 99
rect 9595 -45 9659 19
rect 9595 -125 9659 -61
rect 9595 -205 9659 -141
rect 10201 515 10265 579
rect 10201 435 10265 499
rect 10201 355 10265 419
rect 10201 275 10265 339
rect 10201 195 10265 259
rect 10201 115 10265 179
rect 10201 35 10265 99
rect 10201 -45 10265 19
rect 10201 -125 10265 -61
rect 10201 -205 10265 -141
rect 10327 1675 10391 1739
rect 10327 1595 10391 1659
rect 10327 1515 10391 1579
rect 10327 1435 10391 1499
rect 10327 1355 10391 1419
rect 10327 1275 10391 1339
rect 10327 1195 10391 1259
rect 10327 1115 10391 1179
rect 10327 1035 10391 1099
rect 10327 955 10391 1019
rect 10933 1675 10997 1739
rect 10933 1595 10997 1659
rect 10933 1515 10997 1579
rect 10933 1435 10997 1499
rect 10933 1355 10997 1419
rect 10933 1275 10997 1339
rect 10933 1195 10997 1259
rect 10933 1115 10997 1179
rect 10933 1035 10997 1099
rect 10933 955 10997 1019
rect 11539 1675 11603 1739
rect 11539 1595 11603 1659
rect 11539 1515 11603 1579
rect 11539 1435 11603 1499
rect 11539 1355 11603 1419
rect 11539 1275 11603 1339
rect 11539 1195 11603 1259
rect 11539 1115 11603 1179
rect 11539 1035 11603 1099
rect 11539 955 11603 1019
rect 12145 1675 12209 1739
rect 12145 1595 12209 1659
rect 12145 1515 12209 1579
rect 12145 1435 12209 1499
rect 12145 1355 12209 1419
rect 12145 1275 12209 1339
rect 12145 1195 12209 1259
rect 12145 1115 12209 1179
rect 12145 1035 12209 1099
rect 12145 955 12209 1019
rect 12751 1675 12815 1739
rect 12751 1595 12815 1659
rect 12751 1515 12815 1579
rect 12751 1435 12815 1499
rect 12751 1355 12815 1419
rect 12751 1275 12815 1339
rect 12751 1195 12815 1259
rect 12751 1115 12815 1179
rect 12751 1035 12815 1099
rect 12751 955 12815 1019
rect 13357 1675 13421 1739
rect 13357 1595 13421 1659
rect 13357 1515 13421 1579
rect 13357 1435 13421 1499
rect 13357 1355 13421 1419
rect 13357 1275 13421 1339
rect 13357 1195 13421 1259
rect 13357 1115 13421 1179
rect 13357 1035 13421 1099
rect 13357 955 13421 1019
rect 13963 1675 14027 1739
rect 13963 1595 14027 1659
rect 13963 1515 14027 1579
rect 13963 1435 14027 1499
rect 13963 1355 14027 1419
rect 13963 1275 14027 1339
rect 13963 1195 14027 1259
rect 13963 1115 14027 1179
rect 13963 1035 14027 1099
rect 13963 955 14027 1019
rect 14569 1675 14633 1739
rect 14569 1595 14633 1659
rect 14569 1515 14633 1579
rect 14569 1435 14633 1499
rect 14569 1355 14633 1419
rect 14569 1275 14633 1339
rect 14569 1195 14633 1259
rect 14569 1115 14633 1179
rect 14569 1035 14633 1099
rect 14569 955 14633 1019
rect 15175 1675 15239 1739
rect 15175 1595 15239 1659
rect 15175 1515 15239 1579
rect 15175 1435 15239 1499
rect 15175 1355 15239 1419
rect 15175 1275 15239 1339
rect 15175 1195 15239 1259
rect 15175 1115 15239 1179
rect 15175 1035 15239 1099
rect 15175 955 15239 1019
rect 15781 1675 15845 1739
rect 15781 1595 15845 1659
rect 15781 1515 15845 1579
rect 15781 1435 15845 1499
rect 15781 1355 15845 1419
rect 15781 1275 15845 1339
rect 15781 1195 15845 1259
rect 15781 1115 15845 1179
rect 15781 1035 15845 1099
rect 15781 955 15845 1019
rect 16387 1675 16451 1739
rect 16387 1595 16451 1659
rect 16387 1515 16451 1579
rect 16387 1435 16451 1499
rect 16387 1355 16451 1419
rect 16387 1275 16451 1339
rect 16387 1195 16451 1259
rect 16387 1115 16451 1179
rect 16387 1035 16451 1099
rect 16387 955 16451 1019
rect 16993 1675 17057 1739
rect 16993 1595 17057 1659
rect 16993 1515 17057 1579
rect 16993 1435 17057 1499
rect 16993 1355 17057 1419
rect 16993 1275 17057 1339
rect 16993 1195 17057 1259
rect 16993 1115 17057 1179
rect 16993 1035 17057 1099
rect 16993 955 17057 1019
rect 17599 1675 17663 1739
rect 17599 1595 17663 1659
rect 17599 1515 17663 1579
rect 17599 1435 17663 1499
rect 17599 1355 17663 1419
rect 17599 1275 17663 1339
rect 17599 1195 17663 1259
rect 17599 1115 17663 1179
rect 17599 1035 17663 1099
rect 17599 955 17663 1019
rect 18205 1675 18269 1739
rect 18205 1595 18269 1659
rect 18205 1515 18269 1579
rect 18205 1435 18269 1499
rect 18205 1355 18269 1419
rect 18205 1275 18269 1339
rect 18205 1195 18269 1259
rect 18205 1115 18269 1179
rect 18205 1035 18269 1099
rect 18205 955 18269 1019
rect 18811 1675 18875 1739
rect 18811 1595 18875 1659
rect 18811 1515 18875 1579
rect 18811 1435 18875 1499
rect 18811 1355 18875 1419
rect 18811 1275 18875 1339
rect 18811 1195 18875 1259
rect 18811 1115 18875 1179
rect 18811 1035 18875 1099
rect 18811 955 18875 1019
rect 19417 1675 19481 1739
rect 19417 1595 19481 1659
rect 19417 1515 19481 1579
rect 19417 1435 19481 1499
rect 19417 1355 19481 1419
rect 19417 1275 19481 1339
rect 19417 1195 19481 1259
rect 19417 1115 19481 1179
rect 19417 1035 19481 1099
rect 19417 955 19481 1019
rect 20023 1675 20087 1739
rect 20023 1595 20087 1659
rect 20023 1515 20087 1579
rect 20023 1435 20087 1499
rect 20023 1355 20087 1419
rect 20023 1275 20087 1339
rect 20023 1195 20087 1259
rect 20023 1115 20087 1179
rect 20023 1035 20087 1099
rect 20023 955 20087 1019
rect 10430 735 10494 799
rect 10510 735 10574 799
rect 10590 735 10654 799
rect 10670 735 10734 799
rect 10750 735 10814 799
rect 10830 735 10894 799
rect 11036 735 11100 799
rect 11116 735 11180 799
rect 11196 735 11260 799
rect 11276 735 11340 799
rect 11356 735 11420 799
rect 11436 735 11500 799
rect 11642 735 11706 799
rect 11722 735 11786 799
rect 11802 735 11866 799
rect 11882 735 11946 799
rect 11962 735 12026 799
rect 12042 735 12106 799
rect 12248 735 12312 799
rect 12328 735 12392 799
rect 12408 735 12472 799
rect 12488 735 12552 799
rect 12568 735 12632 799
rect 12648 735 12712 799
rect 12854 735 12918 799
rect 12934 735 12998 799
rect 13014 735 13078 799
rect 13094 735 13158 799
rect 13174 735 13238 799
rect 13254 735 13318 799
rect 13460 735 13524 799
rect 13540 735 13604 799
rect 13620 735 13684 799
rect 13700 735 13764 799
rect 13780 735 13844 799
rect 13860 735 13924 799
rect 14066 735 14130 799
rect 14146 735 14210 799
rect 14226 735 14290 799
rect 14306 735 14370 799
rect 14386 735 14450 799
rect 14466 735 14530 799
rect 14672 735 14736 799
rect 14752 735 14816 799
rect 14832 735 14896 799
rect 14912 735 14976 799
rect 14992 735 15056 799
rect 15072 735 15136 799
rect 15278 735 15342 799
rect 15358 735 15422 799
rect 15438 735 15502 799
rect 15518 735 15582 799
rect 15598 735 15662 799
rect 15678 735 15742 799
rect 15884 735 15948 799
rect 15964 735 16028 799
rect 16044 735 16108 799
rect 16124 735 16188 799
rect 16204 735 16268 799
rect 16284 735 16348 799
rect 16490 735 16554 799
rect 16570 735 16634 799
rect 16650 735 16714 799
rect 16730 735 16794 799
rect 16810 735 16874 799
rect 16890 735 16954 799
rect 17096 735 17160 799
rect 17176 735 17240 799
rect 17256 735 17320 799
rect 17336 735 17400 799
rect 17416 735 17480 799
rect 17496 735 17560 799
rect 17702 735 17766 799
rect 17782 735 17846 799
rect 17862 735 17926 799
rect 17942 735 18006 799
rect 18022 735 18086 799
rect 18102 735 18166 799
rect 18308 735 18372 799
rect 18388 735 18452 799
rect 18468 735 18532 799
rect 18548 735 18612 799
rect 18628 735 18692 799
rect 18708 735 18772 799
rect 18914 735 18978 799
rect 18994 735 19058 799
rect 19074 735 19138 799
rect 19154 735 19218 799
rect 19234 735 19298 799
rect 19314 735 19378 799
rect 19520 735 19584 799
rect 19600 735 19664 799
rect 19680 735 19744 799
rect 19760 735 19824 799
rect 19840 735 19904 799
rect 19920 735 19984 799
rect 10327 515 10391 579
rect 10327 435 10391 499
rect 10327 355 10391 419
rect 10327 275 10391 339
rect 10327 195 10391 259
rect 10327 115 10391 179
rect 10327 35 10391 99
rect 10327 -45 10391 19
rect 10327 -125 10391 -61
rect 10327 -205 10391 -141
rect 10933 515 10997 579
rect 10933 435 10997 499
rect 10933 355 10997 419
rect 10933 275 10997 339
rect 10933 195 10997 259
rect 10933 115 10997 179
rect 10933 35 10997 99
rect 10933 -45 10997 19
rect 10933 -125 10997 -61
rect 10933 -205 10997 -141
rect 11539 515 11603 579
rect 11539 435 11603 499
rect 11539 355 11603 419
rect 11539 275 11603 339
rect 11539 195 11603 259
rect 11539 115 11603 179
rect 11539 35 11603 99
rect 11539 -45 11603 19
rect 11539 -125 11603 -61
rect 11539 -205 11603 -141
rect 12145 515 12209 579
rect 12145 435 12209 499
rect 12145 355 12209 419
rect 12145 275 12209 339
rect 12145 195 12209 259
rect 12145 115 12209 179
rect 12145 35 12209 99
rect 12145 -45 12209 19
rect 12145 -125 12209 -61
rect 12145 -205 12209 -141
rect 12751 515 12815 579
rect 12751 435 12815 499
rect 12751 355 12815 419
rect 12751 275 12815 339
rect 12751 195 12815 259
rect 12751 115 12815 179
rect 12751 35 12815 99
rect 12751 -45 12815 19
rect 12751 -125 12815 -61
rect 12751 -205 12815 -141
rect 13357 515 13421 579
rect 13357 435 13421 499
rect 13357 355 13421 419
rect 13357 275 13421 339
rect 13357 195 13421 259
rect 13357 115 13421 179
rect 13357 35 13421 99
rect 13357 -45 13421 19
rect 13357 -125 13421 -61
rect 13357 -205 13421 -141
rect 13963 515 14027 579
rect 13963 435 14027 499
rect 13963 355 14027 419
rect 13963 275 14027 339
rect 13963 195 14027 259
rect 13963 115 14027 179
rect 13963 35 14027 99
rect 13963 -45 14027 19
rect 13963 -125 14027 -61
rect 13963 -205 14027 -141
rect 14569 515 14633 579
rect 14569 435 14633 499
rect 14569 355 14633 419
rect 14569 275 14633 339
rect 14569 195 14633 259
rect 14569 115 14633 179
rect 14569 35 14633 99
rect 14569 -45 14633 19
rect 14569 -125 14633 -61
rect 14569 -205 14633 -141
rect 15175 515 15239 579
rect 15175 435 15239 499
rect 15175 355 15239 419
rect 15175 275 15239 339
rect 15175 195 15239 259
rect 15175 115 15239 179
rect 15175 35 15239 99
rect 15175 -45 15239 19
rect 15175 -125 15239 -61
rect 15175 -205 15239 -141
rect 15781 515 15845 579
rect 15781 435 15845 499
rect 15781 355 15845 419
rect 15781 275 15845 339
rect 15781 195 15845 259
rect 15781 115 15845 179
rect 15781 35 15845 99
rect 15781 -45 15845 19
rect 15781 -125 15845 -61
rect 15781 -205 15845 -141
rect 16387 515 16451 579
rect 16387 435 16451 499
rect 16387 355 16451 419
rect 16387 275 16451 339
rect 16387 195 16451 259
rect 16387 115 16451 179
rect 16387 35 16451 99
rect 16387 -45 16451 19
rect 16387 -125 16451 -61
rect 16387 -205 16451 -141
rect 16993 515 17057 579
rect 16993 435 17057 499
rect 16993 355 17057 419
rect 16993 275 17057 339
rect 16993 195 17057 259
rect 16993 115 17057 179
rect 16993 35 17057 99
rect 16993 -45 17057 19
rect 16993 -125 17057 -61
rect 16993 -205 17057 -141
rect 17599 515 17663 579
rect 17599 435 17663 499
rect 17599 355 17663 419
rect 17599 275 17663 339
rect 17599 195 17663 259
rect 17599 115 17663 179
rect 17599 35 17663 99
rect 17599 -45 17663 19
rect 17599 -125 17663 -61
rect 17599 -205 17663 -141
rect 18205 515 18269 579
rect 18205 435 18269 499
rect 18205 355 18269 419
rect 18205 275 18269 339
rect 18205 195 18269 259
rect 18205 115 18269 179
rect 18205 35 18269 99
rect 18205 -45 18269 19
rect 18205 -125 18269 -61
rect 18205 -205 18269 -141
rect 18811 515 18875 579
rect 18811 435 18875 499
rect 18811 355 18875 419
rect 18811 275 18875 339
rect 18811 195 18875 259
rect 18811 115 18875 179
rect 18811 35 18875 99
rect 18811 -45 18875 19
rect 18811 -125 18875 -61
rect 18811 -205 18875 -141
rect 19417 515 19481 579
rect 19417 435 19481 499
rect 19417 355 19481 419
rect 19417 275 19481 339
rect 19417 195 19481 259
rect 19417 115 19481 179
rect 19417 35 19481 99
rect 19417 -45 19481 19
rect 19417 -125 19481 -61
rect 19417 -205 19481 -141
rect 20023 515 20087 579
rect 20023 435 20087 499
rect 20023 355 20087 419
rect 20023 275 20087 339
rect 20023 195 20087 259
rect 20023 115 20087 179
rect 20023 35 20087 99
rect 20023 -45 20087 19
rect 20023 -125 20087 -61
rect 20023 -205 20087 -141
rect 20149 1675 20213 1739
rect 20149 1595 20213 1659
rect 20149 1515 20213 1579
rect 20149 1435 20213 1499
rect 20149 1355 20213 1419
rect 20149 1275 20213 1339
rect 20149 1195 20213 1259
rect 20149 1115 20213 1179
rect 20149 1035 20213 1099
rect 20149 955 20213 1019
rect 20755 1675 20819 1739
rect 20755 1595 20819 1659
rect 20755 1515 20819 1579
rect 20755 1435 20819 1499
rect 20755 1355 20819 1419
rect 20755 1275 20819 1339
rect 20755 1195 20819 1259
rect 20755 1115 20819 1179
rect 20755 1035 20819 1099
rect 20755 955 20819 1019
rect 21361 1675 21425 1739
rect 21361 1595 21425 1659
rect 21361 1515 21425 1579
rect 21361 1435 21425 1499
rect 21361 1355 21425 1419
rect 21361 1275 21425 1339
rect 21361 1195 21425 1259
rect 21361 1115 21425 1179
rect 21361 1035 21425 1099
rect 21361 955 21425 1019
rect 21967 1675 22031 1739
rect 21967 1595 22031 1659
rect 21967 1515 22031 1579
rect 21967 1435 22031 1499
rect 21967 1355 22031 1419
rect 21967 1275 22031 1339
rect 21967 1195 22031 1259
rect 21967 1115 22031 1179
rect 21967 1035 22031 1099
rect 21967 955 22031 1019
rect 22573 1675 22637 1739
rect 22573 1595 22637 1659
rect 22573 1515 22637 1579
rect 22573 1435 22637 1499
rect 22573 1355 22637 1419
rect 22573 1275 22637 1339
rect 22573 1195 22637 1259
rect 22573 1115 22637 1179
rect 22573 1035 22637 1099
rect 22573 955 22637 1019
rect 23179 1675 23243 1739
rect 23179 1595 23243 1659
rect 23179 1515 23243 1579
rect 23179 1435 23243 1499
rect 23179 1355 23243 1419
rect 23179 1275 23243 1339
rect 23179 1195 23243 1259
rect 23179 1115 23243 1179
rect 23179 1035 23243 1099
rect 23179 955 23243 1019
rect 23785 1675 23849 1739
rect 23785 1595 23849 1659
rect 23785 1515 23849 1579
rect 23785 1435 23849 1499
rect 23785 1355 23849 1419
rect 23785 1275 23849 1339
rect 23785 1195 23849 1259
rect 23785 1115 23849 1179
rect 23785 1035 23849 1099
rect 23785 955 23849 1019
rect 24391 1675 24455 1739
rect 24391 1595 24455 1659
rect 24391 1515 24455 1579
rect 24391 1435 24455 1499
rect 24391 1355 24455 1419
rect 24391 1275 24455 1339
rect 24391 1195 24455 1259
rect 24391 1115 24455 1179
rect 24391 1035 24455 1099
rect 24391 955 24455 1019
rect 24997 1675 25061 1739
rect 24997 1595 25061 1659
rect 24997 1515 25061 1579
rect 24997 1435 25061 1499
rect 24997 1355 25061 1419
rect 24997 1275 25061 1339
rect 24997 1195 25061 1259
rect 24997 1115 25061 1179
rect 24997 1035 25061 1099
rect 24997 955 25061 1019
rect 25603 1675 25667 1739
rect 25603 1595 25667 1659
rect 25603 1515 25667 1579
rect 25603 1435 25667 1499
rect 25603 1355 25667 1419
rect 25603 1275 25667 1339
rect 25603 1195 25667 1259
rect 25603 1115 25667 1179
rect 25603 1035 25667 1099
rect 25603 955 25667 1019
rect 26209 1675 26273 1739
rect 26209 1595 26273 1659
rect 26209 1515 26273 1579
rect 26209 1435 26273 1499
rect 26209 1355 26273 1419
rect 26209 1275 26273 1339
rect 26209 1195 26273 1259
rect 26209 1115 26273 1179
rect 26209 1035 26273 1099
rect 26209 955 26273 1019
rect 26815 1675 26879 1739
rect 26815 1595 26879 1659
rect 26815 1515 26879 1579
rect 26815 1435 26879 1499
rect 26815 1355 26879 1419
rect 26815 1275 26879 1339
rect 26815 1195 26879 1259
rect 26815 1115 26879 1179
rect 26815 1035 26879 1099
rect 26815 955 26879 1019
rect 27421 1675 27485 1739
rect 27421 1595 27485 1659
rect 27421 1515 27485 1579
rect 27421 1435 27485 1499
rect 27421 1355 27485 1419
rect 27421 1275 27485 1339
rect 27421 1195 27485 1259
rect 27421 1115 27485 1179
rect 27421 1035 27485 1099
rect 27421 955 27485 1019
rect 28027 1675 28091 1739
rect 28027 1595 28091 1659
rect 28027 1515 28091 1579
rect 28027 1435 28091 1499
rect 28027 1355 28091 1419
rect 28027 1275 28091 1339
rect 28027 1195 28091 1259
rect 28027 1115 28091 1179
rect 28027 1035 28091 1099
rect 28027 955 28091 1019
rect 28633 1675 28697 1739
rect 28633 1595 28697 1659
rect 28633 1515 28697 1579
rect 28633 1435 28697 1499
rect 28633 1355 28697 1419
rect 28633 1275 28697 1339
rect 28633 1195 28697 1259
rect 28633 1115 28697 1179
rect 28633 1035 28697 1099
rect 28633 955 28697 1019
rect 29239 1675 29303 1739
rect 29239 1595 29303 1659
rect 29239 1515 29303 1579
rect 29239 1435 29303 1499
rect 29239 1355 29303 1419
rect 29239 1275 29303 1339
rect 29239 1195 29303 1259
rect 29239 1115 29303 1179
rect 29239 1035 29303 1099
rect 29239 955 29303 1019
rect 29845 1675 29909 1739
rect 29845 1595 29909 1659
rect 29845 1515 29909 1579
rect 29845 1435 29909 1499
rect 29845 1355 29909 1419
rect 29845 1275 29909 1339
rect 29845 1195 29909 1259
rect 29845 1115 29909 1179
rect 29845 1035 29909 1099
rect 29845 955 29909 1019
rect 30451 1675 30515 1739
rect 30451 1595 30515 1659
rect 30451 1515 30515 1579
rect 30451 1435 30515 1499
rect 30451 1355 30515 1419
rect 30451 1275 30515 1339
rect 30451 1195 30515 1259
rect 30451 1115 30515 1179
rect 30451 1035 30515 1099
rect 30451 955 30515 1019
rect 31057 1675 31121 1739
rect 31057 1595 31121 1659
rect 31057 1515 31121 1579
rect 31057 1435 31121 1499
rect 31057 1355 31121 1419
rect 31057 1275 31121 1339
rect 31057 1195 31121 1259
rect 31057 1115 31121 1179
rect 31057 1035 31121 1099
rect 31057 955 31121 1019
rect 31663 1675 31727 1739
rect 31663 1595 31727 1659
rect 31663 1515 31727 1579
rect 31663 1435 31727 1499
rect 31663 1355 31727 1419
rect 31663 1275 31727 1339
rect 31663 1195 31727 1259
rect 31663 1115 31727 1179
rect 31663 1035 31727 1099
rect 31663 955 31727 1019
rect 32269 1675 32333 1739
rect 32269 1595 32333 1659
rect 32269 1515 32333 1579
rect 32269 1435 32333 1499
rect 32269 1355 32333 1419
rect 32269 1275 32333 1339
rect 32269 1195 32333 1259
rect 32269 1115 32333 1179
rect 32269 1035 32333 1099
rect 32269 955 32333 1019
rect 32875 1675 32939 1739
rect 32875 1595 32939 1659
rect 32875 1515 32939 1579
rect 32875 1435 32939 1499
rect 32875 1355 32939 1419
rect 32875 1275 32939 1339
rect 32875 1195 32939 1259
rect 32875 1115 32939 1179
rect 32875 1035 32939 1099
rect 32875 955 32939 1019
rect 33481 1675 33545 1739
rect 33481 1595 33545 1659
rect 33481 1515 33545 1579
rect 33481 1435 33545 1499
rect 33481 1355 33545 1419
rect 33481 1275 33545 1339
rect 33481 1195 33545 1259
rect 33481 1115 33545 1179
rect 33481 1035 33545 1099
rect 33481 955 33545 1019
rect 34087 1675 34151 1739
rect 34087 1595 34151 1659
rect 34087 1515 34151 1579
rect 34087 1435 34151 1499
rect 34087 1355 34151 1419
rect 34087 1275 34151 1339
rect 34087 1195 34151 1259
rect 34087 1115 34151 1179
rect 34087 1035 34151 1099
rect 34087 955 34151 1019
rect 34693 1675 34757 1739
rect 34693 1595 34757 1659
rect 34693 1515 34757 1579
rect 34693 1435 34757 1499
rect 34693 1355 34757 1419
rect 34693 1275 34757 1339
rect 34693 1195 34757 1259
rect 34693 1115 34757 1179
rect 34693 1035 34757 1099
rect 34693 955 34757 1019
rect 35299 1675 35363 1739
rect 35299 1595 35363 1659
rect 35299 1515 35363 1579
rect 35299 1435 35363 1499
rect 35299 1355 35363 1419
rect 35299 1275 35363 1339
rect 35299 1195 35363 1259
rect 35299 1115 35363 1179
rect 35299 1035 35363 1099
rect 35299 955 35363 1019
rect 35905 1675 35969 1739
rect 35905 1595 35969 1659
rect 35905 1515 35969 1579
rect 35905 1435 35969 1499
rect 35905 1355 35969 1419
rect 35905 1275 35969 1339
rect 35905 1195 35969 1259
rect 35905 1115 35969 1179
rect 35905 1035 35969 1099
rect 35905 955 35969 1019
rect 36511 1675 36575 1739
rect 36511 1595 36575 1659
rect 36511 1515 36575 1579
rect 36511 1435 36575 1499
rect 36511 1355 36575 1419
rect 36511 1275 36575 1339
rect 36511 1195 36575 1259
rect 36511 1115 36575 1179
rect 36511 1035 36575 1099
rect 36511 955 36575 1019
rect 37117 1675 37181 1739
rect 37117 1595 37181 1659
rect 37117 1515 37181 1579
rect 37117 1435 37181 1499
rect 37117 1355 37181 1419
rect 37117 1275 37181 1339
rect 37117 1195 37181 1259
rect 37117 1115 37181 1179
rect 37117 1035 37181 1099
rect 37117 955 37181 1019
rect 37723 1675 37787 1739
rect 37723 1595 37787 1659
rect 37723 1515 37787 1579
rect 37723 1435 37787 1499
rect 37723 1355 37787 1419
rect 37723 1275 37787 1339
rect 37723 1195 37787 1259
rect 37723 1115 37787 1179
rect 37723 1035 37787 1099
rect 37723 955 37787 1019
rect 38329 1675 38393 1739
rect 38329 1595 38393 1659
rect 38329 1515 38393 1579
rect 38329 1435 38393 1499
rect 38329 1355 38393 1419
rect 38329 1275 38393 1339
rect 38329 1195 38393 1259
rect 38329 1115 38393 1179
rect 38329 1035 38393 1099
rect 38329 955 38393 1019
rect 38935 1675 38999 1739
rect 38935 1595 38999 1659
rect 38935 1515 38999 1579
rect 38935 1435 38999 1499
rect 38935 1355 38999 1419
rect 38935 1275 38999 1339
rect 38935 1195 38999 1259
rect 38935 1115 38999 1179
rect 38935 1035 38999 1099
rect 38935 955 38999 1019
rect 39541 1675 39605 1739
rect 39541 1595 39605 1659
rect 39541 1515 39605 1579
rect 39541 1435 39605 1499
rect 39541 1355 39605 1419
rect 39541 1275 39605 1339
rect 39541 1195 39605 1259
rect 39541 1115 39605 1179
rect 39541 1035 39605 1099
rect 39541 955 39605 1019
rect 20252 735 20316 799
rect 20332 735 20396 799
rect 20412 735 20476 799
rect 20492 735 20556 799
rect 20572 735 20636 799
rect 20652 735 20716 799
rect 20858 735 20922 799
rect 20938 735 21002 799
rect 21018 735 21082 799
rect 21098 735 21162 799
rect 21178 735 21242 799
rect 21258 735 21322 799
rect 21464 735 21528 799
rect 21544 735 21608 799
rect 21624 735 21688 799
rect 21704 735 21768 799
rect 21784 735 21848 799
rect 21864 735 21928 799
rect 22070 735 22134 799
rect 22150 735 22214 799
rect 22230 735 22294 799
rect 22310 735 22374 799
rect 22390 735 22454 799
rect 22470 735 22534 799
rect 22676 735 22740 799
rect 22756 735 22820 799
rect 22836 735 22900 799
rect 22916 735 22980 799
rect 22996 735 23060 799
rect 23076 735 23140 799
rect 23282 735 23346 799
rect 23362 735 23426 799
rect 23442 735 23506 799
rect 23522 735 23586 799
rect 23602 735 23666 799
rect 23682 735 23746 799
rect 23888 735 23952 799
rect 23968 735 24032 799
rect 24048 735 24112 799
rect 24128 735 24192 799
rect 24208 735 24272 799
rect 24288 735 24352 799
rect 24494 735 24558 799
rect 24574 735 24638 799
rect 24654 735 24718 799
rect 24734 735 24798 799
rect 24814 735 24878 799
rect 24894 735 24958 799
rect 25100 735 25164 799
rect 25180 735 25244 799
rect 25260 735 25324 799
rect 25340 735 25404 799
rect 25420 735 25484 799
rect 25500 735 25564 799
rect 25706 735 25770 799
rect 25786 735 25850 799
rect 25866 735 25930 799
rect 25946 735 26010 799
rect 26026 735 26090 799
rect 26106 735 26170 799
rect 26312 735 26376 799
rect 26392 735 26456 799
rect 26472 735 26536 799
rect 26552 735 26616 799
rect 26632 735 26696 799
rect 26712 735 26776 799
rect 26918 735 26982 799
rect 26998 735 27062 799
rect 27078 735 27142 799
rect 27158 735 27222 799
rect 27238 735 27302 799
rect 27318 735 27382 799
rect 27524 735 27588 799
rect 27604 735 27668 799
rect 27684 735 27748 799
rect 27764 735 27828 799
rect 27844 735 27908 799
rect 27924 735 27988 799
rect 28130 735 28194 799
rect 28210 735 28274 799
rect 28290 735 28354 799
rect 28370 735 28434 799
rect 28450 735 28514 799
rect 28530 735 28594 799
rect 28736 735 28800 799
rect 28816 735 28880 799
rect 28896 735 28960 799
rect 28976 735 29040 799
rect 29056 735 29120 799
rect 29136 735 29200 799
rect 29342 735 29406 799
rect 29422 735 29486 799
rect 29502 735 29566 799
rect 29582 735 29646 799
rect 29662 735 29726 799
rect 29742 735 29806 799
rect 29948 735 30012 799
rect 30028 735 30092 799
rect 30108 735 30172 799
rect 30188 735 30252 799
rect 30268 735 30332 799
rect 30348 735 30412 799
rect 30554 735 30618 799
rect 30634 735 30698 799
rect 30714 735 30778 799
rect 30794 735 30858 799
rect 30874 735 30938 799
rect 30954 735 31018 799
rect 31160 735 31224 799
rect 31240 735 31304 799
rect 31320 735 31384 799
rect 31400 735 31464 799
rect 31480 735 31544 799
rect 31560 735 31624 799
rect 31766 735 31830 799
rect 31846 735 31910 799
rect 31926 735 31990 799
rect 32006 735 32070 799
rect 32086 735 32150 799
rect 32166 735 32230 799
rect 32372 735 32436 799
rect 32452 735 32516 799
rect 32532 735 32596 799
rect 32612 735 32676 799
rect 32692 735 32756 799
rect 32772 735 32836 799
rect 32978 735 33042 799
rect 33058 735 33122 799
rect 33138 735 33202 799
rect 33218 735 33282 799
rect 33298 735 33362 799
rect 33378 735 33442 799
rect 33584 735 33648 799
rect 33664 735 33728 799
rect 33744 735 33808 799
rect 33824 735 33888 799
rect 33904 735 33968 799
rect 33984 735 34048 799
rect 34190 735 34254 799
rect 34270 735 34334 799
rect 34350 735 34414 799
rect 34430 735 34494 799
rect 34510 735 34574 799
rect 34590 735 34654 799
rect 34796 735 34860 799
rect 34876 735 34940 799
rect 34956 735 35020 799
rect 35036 735 35100 799
rect 35116 735 35180 799
rect 35196 735 35260 799
rect 35402 735 35466 799
rect 35482 735 35546 799
rect 35562 735 35626 799
rect 35642 735 35706 799
rect 35722 735 35786 799
rect 35802 735 35866 799
rect 36008 735 36072 799
rect 36088 735 36152 799
rect 36168 735 36232 799
rect 36248 735 36312 799
rect 36328 735 36392 799
rect 36408 735 36472 799
rect 36614 735 36678 799
rect 36694 735 36758 799
rect 36774 735 36838 799
rect 36854 735 36918 799
rect 36934 735 36998 799
rect 37014 735 37078 799
rect 37220 735 37284 799
rect 37300 735 37364 799
rect 37380 735 37444 799
rect 37460 735 37524 799
rect 37540 735 37604 799
rect 37620 735 37684 799
rect 37826 735 37890 799
rect 37906 735 37970 799
rect 37986 735 38050 799
rect 38066 735 38130 799
rect 38146 735 38210 799
rect 38226 735 38290 799
rect 38432 735 38496 799
rect 38512 735 38576 799
rect 38592 735 38656 799
rect 38672 735 38736 799
rect 38752 735 38816 799
rect 38832 735 38896 799
rect 39038 735 39102 799
rect 39118 735 39182 799
rect 39198 735 39262 799
rect 39278 735 39342 799
rect 39358 735 39422 799
rect 39438 735 39502 799
rect 20149 515 20213 579
rect 20149 435 20213 499
rect 20149 355 20213 419
rect 20149 275 20213 339
rect 20149 195 20213 259
rect 20149 115 20213 179
rect 20149 35 20213 99
rect 20149 -45 20213 19
rect 20149 -125 20213 -61
rect 20149 -205 20213 -141
rect 20755 515 20819 579
rect 20755 435 20819 499
rect 20755 355 20819 419
rect 20755 275 20819 339
rect 20755 195 20819 259
rect 20755 115 20819 179
rect 20755 35 20819 99
rect 20755 -45 20819 19
rect 20755 -125 20819 -61
rect 20755 -205 20819 -141
rect 21361 515 21425 579
rect 21361 435 21425 499
rect 21361 355 21425 419
rect 21361 275 21425 339
rect 21361 195 21425 259
rect 21361 115 21425 179
rect 21361 35 21425 99
rect 21361 -45 21425 19
rect 21361 -125 21425 -61
rect 21361 -205 21425 -141
rect 21967 515 22031 579
rect 21967 435 22031 499
rect 21967 355 22031 419
rect 21967 275 22031 339
rect 21967 195 22031 259
rect 21967 115 22031 179
rect 21967 35 22031 99
rect 21967 -45 22031 19
rect 21967 -125 22031 -61
rect 21967 -205 22031 -141
rect 22573 515 22637 579
rect 22573 435 22637 499
rect 22573 355 22637 419
rect 22573 275 22637 339
rect 22573 195 22637 259
rect 22573 115 22637 179
rect 22573 35 22637 99
rect 22573 -45 22637 19
rect 22573 -125 22637 -61
rect 22573 -205 22637 -141
rect 23179 515 23243 579
rect 23179 435 23243 499
rect 23179 355 23243 419
rect 23179 275 23243 339
rect 23179 195 23243 259
rect 23179 115 23243 179
rect 23179 35 23243 99
rect 23179 -45 23243 19
rect 23179 -125 23243 -61
rect 23179 -205 23243 -141
rect 23785 515 23849 579
rect 23785 435 23849 499
rect 23785 355 23849 419
rect 23785 275 23849 339
rect 23785 195 23849 259
rect 23785 115 23849 179
rect 23785 35 23849 99
rect 23785 -45 23849 19
rect 23785 -125 23849 -61
rect 23785 -205 23849 -141
rect 24391 515 24455 579
rect 24391 435 24455 499
rect 24391 355 24455 419
rect 24391 275 24455 339
rect 24391 195 24455 259
rect 24391 115 24455 179
rect 24391 35 24455 99
rect 24391 -45 24455 19
rect 24391 -125 24455 -61
rect 24391 -205 24455 -141
rect 24997 515 25061 579
rect 24997 435 25061 499
rect 24997 355 25061 419
rect 24997 275 25061 339
rect 24997 195 25061 259
rect 24997 115 25061 179
rect 24997 35 25061 99
rect 24997 -45 25061 19
rect 24997 -125 25061 -61
rect 24997 -205 25061 -141
rect 25603 515 25667 579
rect 25603 435 25667 499
rect 25603 355 25667 419
rect 25603 275 25667 339
rect 25603 195 25667 259
rect 25603 115 25667 179
rect 25603 35 25667 99
rect 25603 -45 25667 19
rect 25603 -125 25667 -61
rect 25603 -205 25667 -141
rect 26209 515 26273 579
rect 26209 435 26273 499
rect 26209 355 26273 419
rect 26209 275 26273 339
rect 26209 195 26273 259
rect 26209 115 26273 179
rect 26209 35 26273 99
rect 26209 -45 26273 19
rect 26209 -125 26273 -61
rect 26209 -205 26273 -141
rect 26815 515 26879 579
rect 26815 435 26879 499
rect 26815 355 26879 419
rect 26815 275 26879 339
rect 26815 195 26879 259
rect 26815 115 26879 179
rect 26815 35 26879 99
rect 26815 -45 26879 19
rect 26815 -125 26879 -61
rect 26815 -205 26879 -141
rect 27421 515 27485 579
rect 27421 435 27485 499
rect 27421 355 27485 419
rect 27421 275 27485 339
rect 27421 195 27485 259
rect 27421 115 27485 179
rect 27421 35 27485 99
rect 27421 -45 27485 19
rect 27421 -125 27485 -61
rect 27421 -205 27485 -141
rect 28027 515 28091 579
rect 28027 435 28091 499
rect 28027 355 28091 419
rect 28027 275 28091 339
rect 28027 195 28091 259
rect 28027 115 28091 179
rect 28027 35 28091 99
rect 28027 -45 28091 19
rect 28027 -125 28091 -61
rect 28027 -205 28091 -141
rect 28633 515 28697 579
rect 28633 435 28697 499
rect 28633 355 28697 419
rect 28633 275 28697 339
rect 28633 195 28697 259
rect 28633 115 28697 179
rect 28633 35 28697 99
rect 28633 -45 28697 19
rect 28633 -125 28697 -61
rect 28633 -205 28697 -141
rect 29239 515 29303 579
rect 29239 435 29303 499
rect 29239 355 29303 419
rect 29239 275 29303 339
rect 29239 195 29303 259
rect 29239 115 29303 179
rect 29239 35 29303 99
rect 29239 -45 29303 19
rect 29239 -125 29303 -61
rect 29239 -205 29303 -141
rect 29845 515 29909 579
rect 29845 435 29909 499
rect 29845 355 29909 419
rect 29845 275 29909 339
rect 29845 195 29909 259
rect 29845 115 29909 179
rect 29845 35 29909 99
rect 29845 -45 29909 19
rect 29845 -125 29909 -61
rect 29845 -205 29909 -141
rect 30451 515 30515 579
rect 30451 435 30515 499
rect 30451 355 30515 419
rect 30451 275 30515 339
rect 30451 195 30515 259
rect 30451 115 30515 179
rect 30451 35 30515 99
rect 30451 -45 30515 19
rect 30451 -125 30515 -61
rect 30451 -205 30515 -141
rect 31057 515 31121 579
rect 31057 435 31121 499
rect 31057 355 31121 419
rect 31057 275 31121 339
rect 31057 195 31121 259
rect 31057 115 31121 179
rect 31057 35 31121 99
rect 31057 -45 31121 19
rect 31057 -125 31121 -61
rect 31057 -205 31121 -141
rect 31663 515 31727 579
rect 31663 435 31727 499
rect 31663 355 31727 419
rect 31663 275 31727 339
rect 31663 195 31727 259
rect 31663 115 31727 179
rect 31663 35 31727 99
rect 31663 -45 31727 19
rect 31663 -125 31727 -61
rect 31663 -205 31727 -141
rect 32269 515 32333 579
rect 32269 435 32333 499
rect 32269 355 32333 419
rect 32269 275 32333 339
rect 32269 195 32333 259
rect 32269 115 32333 179
rect 32269 35 32333 99
rect 32269 -45 32333 19
rect 32269 -125 32333 -61
rect 32269 -205 32333 -141
rect 32875 515 32939 579
rect 32875 435 32939 499
rect 32875 355 32939 419
rect 32875 275 32939 339
rect 32875 195 32939 259
rect 32875 115 32939 179
rect 32875 35 32939 99
rect 32875 -45 32939 19
rect 32875 -125 32939 -61
rect 32875 -205 32939 -141
rect 33481 515 33545 579
rect 33481 435 33545 499
rect 33481 355 33545 419
rect 33481 275 33545 339
rect 33481 195 33545 259
rect 33481 115 33545 179
rect 33481 35 33545 99
rect 33481 -45 33545 19
rect 33481 -125 33545 -61
rect 33481 -205 33545 -141
rect 34087 515 34151 579
rect 34087 435 34151 499
rect 34087 355 34151 419
rect 34087 275 34151 339
rect 34087 195 34151 259
rect 34087 115 34151 179
rect 34087 35 34151 99
rect 34087 -45 34151 19
rect 34087 -125 34151 -61
rect 34087 -205 34151 -141
rect 34693 515 34757 579
rect 34693 435 34757 499
rect 34693 355 34757 419
rect 34693 275 34757 339
rect 34693 195 34757 259
rect 34693 115 34757 179
rect 34693 35 34757 99
rect 34693 -45 34757 19
rect 34693 -125 34757 -61
rect 34693 -205 34757 -141
rect 35299 515 35363 579
rect 35299 435 35363 499
rect 35299 355 35363 419
rect 35299 275 35363 339
rect 35299 195 35363 259
rect 35299 115 35363 179
rect 35299 35 35363 99
rect 35299 -45 35363 19
rect 35299 -125 35363 -61
rect 35299 -205 35363 -141
rect 35905 515 35969 579
rect 35905 435 35969 499
rect 35905 355 35969 419
rect 35905 275 35969 339
rect 35905 195 35969 259
rect 35905 115 35969 179
rect 35905 35 35969 99
rect 35905 -45 35969 19
rect 35905 -125 35969 -61
rect 35905 -205 35969 -141
rect 36511 515 36575 579
rect 36511 435 36575 499
rect 36511 355 36575 419
rect 36511 275 36575 339
rect 36511 195 36575 259
rect 36511 115 36575 179
rect 36511 35 36575 99
rect 36511 -45 36575 19
rect 36511 -125 36575 -61
rect 36511 -205 36575 -141
rect 37117 515 37181 579
rect 37117 435 37181 499
rect 37117 355 37181 419
rect 37117 275 37181 339
rect 37117 195 37181 259
rect 37117 115 37181 179
rect 37117 35 37181 99
rect 37117 -45 37181 19
rect 37117 -125 37181 -61
rect 37117 -205 37181 -141
rect 37723 515 37787 579
rect 37723 435 37787 499
rect 37723 355 37787 419
rect 37723 275 37787 339
rect 37723 195 37787 259
rect 37723 115 37787 179
rect 37723 35 37787 99
rect 37723 -45 37787 19
rect 37723 -125 37787 -61
rect 37723 -205 37787 -141
rect 38329 515 38393 579
rect 38329 435 38393 499
rect 38329 355 38393 419
rect 38329 275 38393 339
rect 38329 195 38393 259
rect 38329 115 38393 179
rect 38329 35 38393 99
rect 38329 -45 38393 19
rect 38329 -125 38393 -61
rect 38329 -205 38393 -141
rect 38935 515 38999 579
rect 38935 435 38999 499
rect 38935 355 38999 419
rect 38935 275 38999 339
rect 38935 195 38999 259
rect 38935 115 38999 179
rect 38935 35 38999 99
rect 38935 -45 38999 19
rect 38935 -125 38999 -61
rect 38935 -205 38999 -141
rect 39541 515 39605 579
rect 39541 435 39605 499
rect 39541 355 39605 419
rect 39541 275 39605 339
rect 39541 195 39605 259
rect 39541 115 39605 179
rect 39541 35 39605 99
rect 39541 -45 39605 19
rect 39541 -125 39605 -61
rect 39541 -205 39605 -141
rect -355 -425 -291 -361
rect -275 -425 -211 -361
rect -195 -425 -131 -361
rect -115 -425 -51 -361
rect -35 -425 29 -361
rect 45 -425 109 -361
rect 459 -425 523 -361
rect 539 -425 603 -361
rect 619 -425 683 -361
rect 699 -425 763 -361
rect 779 -425 843 -361
rect 859 -425 923 -361
rect 1371 -425 1435 -361
rect 1451 -425 1515 -361
rect 1531 -425 1595 -361
rect 1611 -425 1675 -361
rect 1691 -425 1755 -361
rect 1771 -425 1835 -361
rect 1977 -425 2041 -361
rect 2057 -425 2121 -361
rect 2137 -425 2201 -361
rect 2217 -425 2281 -361
rect 2297 -425 2361 -361
rect 2377 -425 2441 -361
rect 2905 -425 2969 -361
rect 2985 -425 3049 -361
rect 3065 -425 3129 -361
rect 3145 -425 3209 -361
rect 3225 -425 3289 -361
rect 3305 -425 3369 -361
rect 3511 -425 3575 -361
rect 3591 -425 3655 -361
rect 3671 -425 3735 -361
rect 3751 -425 3815 -361
rect 3831 -425 3895 -361
rect 3911 -425 3975 -361
rect 4117 -425 4181 -361
rect 4197 -425 4261 -361
rect 4277 -425 4341 -361
rect 4357 -425 4421 -361
rect 4437 -425 4501 -361
rect 4517 -425 4581 -361
rect 4723 -425 4787 -361
rect 4803 -425 4867 -361
rect 4883 -425 4947 -361
rect 4963 -425 5027 -361
rect 5043 -425 5107 -361
rect 5123 -425 5187 -361
rect 5456 -425 5520 -361
rect 5536 -425 5600 -361
rect 5616 -425 5680 -361
rect 5696 -425 5760 -361
rect 5776 -425 5840 -361
rect 5856 -425 5920 -361
rect 6062 -425 6126 -361
rect 6142 -425 6206 -361
rect 6222 -425 6286 -361
rect 6302 -425 6366 -361
rect 6382 -425 6446 -361
rect 6462 -425 6526 -361
rect 6668 -425 6732 -361
rect 6748 -425 6812 -361
rect 6828 -425 6892 -361
rect 6908 -425 6972 -361
rect 6988 -425 7052 -361
rect 7068 -425 7132 -361
rect 7274 -425 7338 -361
rect 7354 -425 7418 -361
rect 7434 -425 7498 -361
rect 7514 -425 7578 -361
rect 7594 -425 7658 -361
rect 7674 -425 7738 -361
rect 7880 -425 7944 -361
rect 7960 -425 8024 -361
rect 8040 -425 8104 -361
rect 8120 -425 8184 -361
rect 8200 -425 8264 -361
rect 8280 -425 8344 -361
rect 8486 -425 8550 -361
rect 8566 -425 8630 -361
rect 8646 -425 8710 -361
rect 8726 -425 8790 -361
rect 8806 -425 8870 -361
rect 8886 -425 8950 -361
rect 9092 -425 9156 -361
rect 9172 -425 9236 -361
rect 9252 -425 9316 -361
rect 9332 -425 9396 -361
rect 9412 -425 9476 -361
rect 9492 -425 9556 -361
rect 9698 -425 9762 -361
rect 9778 -425 9842 -361
rect 9858 -425 9922 -361
rect 9938 -425 10002 -361
rect 10018 -425 10082 -361
rect 10098 -425 10162 -361
rect 10430 -425 10494 -361
rect 10510 -425 10574 -361
rect 10590 -425 10654 -361
rect 10670 -425 10734 -361
rect 10750 -425 10814 -361
rect 10830 -425 10894 -361
rect 11036 -425 11100 -361
rect 11116 -425 11180 -361
rect 11196 -425 11260 -361
rect 11276 -425 11340 -361
rect 11356 -425 11420 -361
rect 11436 -425 11500 -361
rect 11642 -425 11706 -361
rect 11722 -425 11786 -361
rect 11802 -425 11866 -361
rect 11882 -425 11946 -361
rect 11962 -425 12026 -361
rect 12042 -425 12106 -361
rect 12248 -425 12312 -361
rect 12328 -425 12392 -361
rect 12408 -425 12472 -361
rect 12488 -425 12552 -361
rect 12568 -425 12632 -361
rect 12648 -425 12712 -361
rect 12854 -425 12918 -361
rect 12934 -425 12998 -361
rect 13014 -425 13078 -361
rect 13094 -425 13158 -361
rect 13174 -425 13238 -361
rect 13254 -425 13318 -361
rect 13460 -425 13524 -361
rect 13540 -425 13604 -361
rect 13620 -425 13684 -361
rect 13700 -425 13764 -361
rect 13780 -425 13844 -361
rect 13860 -425 13924 -361
rect 14066 -425 14130 -361
rect 14146 -425 14210 -361
rect 14226 -425 14290 -361
rect 14306 -425 14370 -361
rect 14386 -425 14450 -361
rect 14466 -425 14530 -361
rect 14672 -425 14736 -361
rect 14752 -425 14816 -361
rect 14832 -425 14896 -361
rect 14912 -425 14976 -361
rect 14992 -425 15056 -361
rect 15072 -425 15136 -361
rect 15278 -425 15342 -361
rect 15358 -425 15422 -361
rect 15438 -425 15502 -361
rect 15518 -425 15582 -361
rect 15598 -425 15662 -361
rect 15678 -425 15742 -361
rect 15884 -425 15948 -361
rect 15964 -425 16028 -361
rect 16044 -425 16108 -361
rect 16124 -425 16188 -361
rect 16204 -425 16268 -361
rect 16284 -425 16348 -361
rect 16490 -425 16554 -361
rect 16570 -425 16634 -361
rect 16650 -425 16714 -361
rect 16730 -425 16794 -361
rect 16810 -425 16874 -361
rect 16890 -425 16954 -361
rect 17096 -425 17160 -361
rect 17176 -425 17240 -361
rect 17256 -425 17320 -361
rect 17336 -425 17400 -361
rect 17416 -425 17480 -361
rect 17496 -425 17560 -361
rect 17702 -425 17766 -361
rect 17782 -425 17846 -361
rect 17862 -425 17926 -361
rect 17942 -425 18006 -361
rect 18022 -425 18086 -361
rect 18102 -425 18166 -361
rect 18308 -425 18372 -361
rect 18388 -425 18452 -361
rect 18468 -425 18532 -361
rect 18548 -425 18612 -361
rect 18628 -425 18692 -361
rect 18708 -425 18772 -361
rect 18914 -425 18978 -361
rect 18994 -425 19058 -361
rect 19074 -425 19138 -361
rect 19154 -425 19218 -361
rect 19234 -425 19298 -361
rect 19314 -425 19378 -361
rect 19520 -425 19584 -361
rect 19600 -425 19664 -361
rect 19680 -425 19744 -361
rect 19760 -425 19824 -361
rect 19840 -425 19904 -361
rect 19920 -425 19984 -361
rect 20252 -425 20316 -361
rect 20332 -425 20396 -361
rect 20412 -425 20476 -361
rect 20492 -425 20556 -361
rect 20572 -425 20636 -361
rect 20652 -425 20716 -361
rect 20858 -425 20922 -361
rect 20938 -425 21002 -361
rect 21018 -425 21082 -361
rect 21098 -425 21162 -361
rect 21178 -425 21242 -361
rect 21258 -425 21322 -361
rect 21464 -425 21528 -361
rect 21544 -425 21608 -361
rect 21624 -425 21688 -361
rect 21704 -425 21768 -361
rect 21784 -425 21848 -361
rect 21864 -425 21928 -361
rect 22070 -425 22134 -361
rect 22150 -425 22214 -361
rect 22230 -425 22294 -361
rect 22310 -425 22374 -361
rect 22390 -425 22454 -361
rect 22470 -425 22534 -361
rect 22676 -425 22740 -361
rect 22756 -425 22820 -361
rect 22836 -425 22900 -361
rect 22916 -425 22980 -361
rect 22996 -425 23060 -361
rect 23076 -425 23140 -361
rect 23282 -425 23346 -361
rect 23362 -425 23426 -361
rect 23442 -425 23506 -361
rect 23522 -425 23586 -361
rect 23602 -425 23666 -361
rect 23682 -425 23746 -361
rect 23888 -425 23952 -361
rect 23968 -425 24032 -361
rect 24048 -425 24112 -361
rect 24128 -425 24192 -361
rect 24208 -425 24272 -361
rect 24288 -425 24352 -361
rect 24494 -425 24558 -361
rect 24574 -425 24638 -361
rect 24654 -425 24718 -361
rect 24734 -425 24798 -361
rect 24814 -425 24878 -361
rect 24894 -425 24958 -361
rect 25100 -425 25164 -361
rect 25180 -425 25244 -361
rect 25260 -425 25324 -361
rect 25340 -425 25404 -361
rect 25420 -425 25484 -361
rect 25500 -425 25564 -361
rect 25706 -425 25770 -361
rect 25786 -425 25850 -361
rect 25866 -425 25930 -361
rect 25946 -425 26010 -361
rect 26026 -425 26090 -361
rect 26106 -425 26170 -361
rect 26312 -425 26376 -361
rect 26392 -425 26456 -361
rect 26472 -425 26536 -361
rect 26552 -425 26616 -361
rect 26632 -425 26696 -361
rect 26712 -425 26776 -361
rect 26918 -425 26982 -361
rect 26998 -425 27062 -361
rect 27078 -425 27142 -361
rect 27158 -425 27222 -361
rect 27238 -425 27302 -361
rect 27318 -425 27382 -361
rect 27524 -425 27588 -361
rect 27604 -425 27668 -361
rect 27684 -425 27748 -361
rect 27764 -425 27828 -361
rect 27844 -425 27908 -361
rect 27924 -425 27988 -361
rect 28130 -425 28194 -361
rect 28210 -425 28274 -361
rect 28290 -425 28354 -361
rect 28370 -425 28434 -361
rect 28450 -425 28514 -361
rect 28530 -425 28594 -361
rect 28736 -425 28800 -361
rect 28816 -425 28880 -361
rect 28896 -425 28960 -361
rect 28976 -425 29040 -361
rect 29056 -425 29120 -361
rect 29136 -425 29200 -361
rect 29342 -425 29406 -361
rect 29422 -425 29486 -361
rect 29502 -425 29566 -361
rect 29582 -425 29646 -361
rect 29662 -425 29726 -361
rect 29742 -425 29806 -361
rect 29948 -425 30012 -361
rect 30028 -425 30092 -361
rect 30108 -425 30172 -361
rect 30188 -425 30252 -361
rect 30268 -425 30332 -361
rect 30348 -425 30412 -361
rect 30554 -425 30618 -361
rect 30634 -425 30698 -361
rect 30714 -425 30778 -361
rect 30794 -425 30858 -361
rect 30874 -425 30938 -361
rect 30954 -425 31018 -361
rect 31160 -425 31224 -361
rect 31240 -425 31304 -361
rect 31320 -425 31384 -361
rect 31400 -425 31464 -361
rect 31480 -425 31544 -361
rect 31560 -425 31624 -361
rect 31766 -425 31830 -361
rect 31846 -425 31910 -361
rect 31926 -425 31990 -361
rect 32006 -425 32070 -361
rect 32086 -425 32150 -361
rect 32166 -425 32230 -361
rect 32372 -425 32436 -361
rect 32452 -425 32516 -361
rect 32532 -425 32596 -361
rect 32612 -425 32676 -361
rect 32692 -425 32756 -361
rect 32772 -425 32836 -361
rect 32978 -425 33042 -361
rect 33058 -425 33122 -361
rect 33138 -425 33202 -361
rect 33218 -425 33282 -361
rect 33298 -425 33362 -361
rect 33378 -425 33442 -361
rect 33584 -425 33648 -361
rect 33664 -425 33728 -361
rect 33744 -425 33808 -361
rect 33824 -425 33888 -361
rect 33904 -425 33968 -361
rect 33984 -425 34048 -361
rect 34190 -425 34254 -361
rect 34270 -425 34334 -361
rect 34350 -425 34414 -361
rect 34430 -425 34494 -361
rect 34510 -425 34574 -361
rect 34590 -425 34654 -361
rect 34796 -425 34860 -361
rect 34876 -425 34940 -361
rect 34956 -425 35020 -361
rect 35036 -425 35100 -361
rect 35116 -425 35180 -361
rect 35196 -425 35260 -361
rect 35402 -425 35466 -361
rect 35482 -425 35546 -361
rect 35562 -425 35626 -361
rect 35642 -425 35706 -361
rect 35722 -425 35786 -361
rect 35802 -425 35866 -361
rect 36008 -425 36072 -361
rect 36088 -425 36152 -361
rect 36168 -425 36232 -361
rect 36248 -425 36312 -361
rect 36328 -425 36392 -361
rect 36408 -425 36472 -361
rect 36614 -425 36678 -361
rect 36694 -425 36758 -361
rect 36774 -425 36838 -361
rect 36854 -425 36918 -361
rect 36934 -425 36998 -361
rect 37014 -425 37078 -361
rect 37220 -425 37284 -361
rect 37300 -425 37364 -361
rect 37380 -425 37444 -361
rect 37460 -425 37524 -361
rect 37540 -425 37604 -361
rect 37620 -425 37684 -361
rect 37826 -425 37890 -361
rect 37906 -425 37970 -361
rect 37986 -425 38050 -361
rect 38066 -425 38130 -361
rect 38146 -425 38210 -361
rect 38226 -425 38290 -361
rect 38432 -425 38496 -361
rect 38512 -425 38576 -361
rect 38592 -425 38656 -361
rect 38672 -425 38736 -361
rect 38752 -425 38816 -361
rect 38832 -425 38896 -361
rect 39038 -425 39102 -361
rect 39118 -425 39182 -361
rect 39198 -425 39262 -361
rect 39278 -425 39342 -361
rect 39358 -425 39422 -361
rect 39438 -425 39502 -361
<< metal4 >>
rect 38511 6075 38950 6291
rect 38065 6013 38298 6014
rect 37836 5748 38298 6013
rect 38511 6011 38525 6075
rect 38589 6011 38950 6075
rect 38511 5806 38950 6011
rect 37836 5684 37845 5748
rect 37909 5684 38298 5748
rect 37836 5449 38298 5684
rect 38065 5448 38298 5449
rect 39077 5742 39565 6049
rect 39077 5678 39090 5742
rect 39154 5678 39565 5742
rect 39077 5415 39565 5678
rect -459 5092 213 5094
rect -459 5028 -355 5092
rect -291 5028 -275 5092
rect -211 5028 -195 5092
rect -131 5028 -115 5092
rect -51 5028 -35 5092
rect 29 5028 45 5092
rect 109 5028 213 5092
rect -459 5026 213 5028
rect 524 5092 1027 5094
rect 524 5028 539 5092
rect 603 5028 619 5092
rect 683 5028 699 5092
rect 763 5028 779 5092
rect 843 5028 859 5092
rect 923 5028 1027 5092
rect 524 5026 1027 5028
rect 1267 5092 1717 5094
rect 1954 5092 2545 5094
rect 1267 5028 1371 5092
rect 1435 5028 1451 5092
rect 1515 5028 1531 5092
rect 1595 5028 1611 5092
rect 1675 5028 1691 5092
rect 1954 5028 1977 5092
rect 2041 5028 2057 5092
rect 2121 5028 2137 5092
rect 2201 5028 2217 5092
rect 2281 5028 2297 5092
rect 2361 5028 2377 5092
rect 2441 5028 2545 5092
rect 1267 5026 1717 5028
rect 1954 5026 2545 5028
rect 2801 5092 3301 5094
rect 3538 5092 5291 5094
rect 2801 5028 2905 5092
rect 2969 5028 2985 5092
rect 3049 5028 3065 5092
rect 3129 5028 3145 5092
rect 3209 5028 3225 5092
rect 3289 5028 3301 5092
rect 3575 5028 3591 5092
rect 3655 5028 3671 5092
rect 3735 5028 3751 5092
rect 3815 5028 3831 5092
rect 3895 5028 3911 5092
rect 3975 5028 4117 5092
rect 4181 5028 4197 5092
rect 4261 5028 4277 5092
rect 4341 5028 4357 5092
rect 4421 5028 4437 5092
rect 4501 5028 4517 5092
rect 4581 5028 4723 5092
rect 4787 5028 4803 5092
rect 4867 5028 4883 5092
rect 4947 5028 4963 5092
rect 5027 5028 5043 5092
rect 5107 5028 5123 5092
rect 5187 5028 5291 5092
rect 2801 5026 3301 5028
rect 3538 5026 5291 5028
rect 5352 5026 5394 5094
rect 5631 5092 10266 5094
rect 5680 5028 5696 5092
rect 5760 5028 5776 5092
rect 5840 5028 5856 5092
rect 5920 5028 6062 5092
rect 6126 5028 6142 5092
rect 6206 5028 6222 5092
rect 6286 5028 6302 5092
rect 6366 5028 6382 5092
rect 6446 5028 6462 5092
rect 6526 5028 6668 5092
rect 6732 5028 6748 5092
rect 6812 5028 6828 5092
rect 6892 5028 6908 5092
rect 6972 5028 6988 5092
rect 7052 5028 7068 5092
rect 7132 5028 7274 5092
rect 7338 5028 7354 5092
rect 7418 5028 7434 5092
rect 7498 5028 7514 5092
rect 7578 5028 7594 5092
rect 7658 5028 7674 5092
rect 7738 5028 7880 5092
rect 7944 5028 7960 5092
rect 8024 5028 8040 5092
rect 8104 5028 8120 5092
rect 8184 5028 8200 5092
rect 8264 5028 8280 5092
rect 8344 5028 8486 5092
rect 8550 5028 8566 5092
rect 8630 5028 8646 5092
rect 8710 5028 8726 5092
rect 8790 5028 8806 5092
rect 8870 5028 8886 5092
rect 8950 5028 9092 5092
rect 9156 5028 9172 5092
rect 9236 5028 9252 5092
rect 9316 5028 9332 5092
rect 9396 5028 9412 5092
rect 9476 5028 9492 5092
rect 9556 5028 9698 5092
rect 9762 5028 9778 5092
rect 9842 5028 9858 5092
rect 9922 5028 9938 5092
rect 10002 5028 10018 5092
rect 10082 5028 10098 5092
rect 10162 5028 10266 5092
rect 5631 5026 10266 5028
rect 10326 5026 10368 5094
rect 10605 5092 20088 5094
rect 10654 5028 10670 5092
rect 10734 5028 10750 5092
rect 10814 5028 10830 5092
rect 10894 5028 11036 5092
rect 11100 5028 11116 5092
rect 11180 5028 11196 5092
rect 11260 5028 11276 5092
rect 11340 5028 11356 5092
rect 11420 5028 11436 5092
rect 11500 5028 11642 5092
rect 11706 5028 11722 5092
rect 11786 5028 11802 5092
rect 11866 5028 11882 5092
rect 11946 5028 11962 5092
rect 12026 5028 12042 5092
rect 12106 5028 12248 5092
rect 12312 5028 12328 5092
rect 12392 5028 12408 5092
rect 12472 5028 12488 5092
rect 12552 5028 12568 5092
rect 12632 5028 12648 5092
rect 12712 5028 12854 5092
rect 12918 5028 12934 5092
rect 12998 5028 13014 5092
rect 13078 5028 13094 5092
rect 13158 5028 13174 5092
rect 13238 5028 13254 5092
rect 13318 5028 13460 5092
rect 13524 5028 13540 5092
rect 13604 5028 13620 5092
rect 13684 5028 13700 5092
rect 13764 5028 13780 5092
rect 13844 5028 13860 5092
rect 13924 5028 14066 5092
rect 14130 5028 14146 5092
rect 14210 5028 14226 5092
rect 14290 5028 14306 5092
rect 14370 5028 14386 5092
rect 14450 5028 14466 5092
rect 14530 5028 14672 5092
rect 14736 5028 14752 5092
rect 14816 5028 14832 5092
rect 14896 5028 14912 5092
rect 14976 5028 14992 5092
rect 15056 5028 15072 5092
rect 15136 5028 15278 5092
rect 15342 5028 15358 5092
rect 15422 5028 15438 5092
rect 15502 5028 15518 5092
rect 15582 5028 15598 5092
rect 15662 5028 15678 5092
rect 15742 5028 15884 5092
rect 15948 5028 15964 5092
rect 16028 5028 16044 5092
rect 16108 5028 16124 5092
rect 16188 5028 16204 5092
rect 16268 5028 16284 5092
rect 16348 5028 16490 5092
rect 16554 5028 16570 5092
rect 16634 5028 16650 5092
rect 16714 5028 16730 5092
rect 16794 5028 16810 5092
rect 16874 5028 16890 5092
rect 16954 5028 17096 5092
rect 17160 5028 17176 5092
rect 17240 5028 17256 5092
rect 17320 5028 17336 5092
rect 17400 5028 17416 5092
rect 17480 5028 17496 5092
rect 17560 5028 17702 5092
rect 17766 5028 17782 5092
rect 17846 5028 17862 5092
rect 17926 5028 17942 5092
rect 18006 5028 18022 5092
rect 18086 5028 18102 5092
rect 18166 5028 18308 5092
rect 18372 5028 18388 5092
rect 18452 5028 18468 5092
rect 18532 5028 18548 5092
rect 18612 5028 18628 5092
rect 18692 5028 18708 5092
rect 18772 5028 18914 5092
rect 18978 5028 18994 5092
rect 19058 5028 19074 5092
rect 19138 5028 19154 5092
rect 19218 5028 19234 5092
rect 19298 5028 19314 5092
rect 19378 5028 19520 5092
rect 19584 5028 19600 5092
rect 19664 5028 19680 5092
rect 19744 5028 19760 5092
rect 19824 5028 19840 5092
rect 19904 5028 19920 5092
rect 19984 5028 20088 5092
rect 10605 5026 20088 5028
rect 20148 5092 39298 5094
rect 20148 5028 20252 5092
rect 20316 5028 20332 5092
rect 20396 5028 20412 5092
rect 20476 5028 20492 5092
rect 20556 5028 20572 5092
rect 20636 5028 20652 5092
rect 20716 5028 20858 5092
rect 20922 5028 20938 5092
rect 21002 5028 21018 5092
rect 21082 5028 21098 5092
rect 21162 5028 21178 5092
rect 21242 5028 21258 5092
rect 21322 5028 21464 5092
rect 21528 5028 21544 5092
rect 21608 5028 21624 5092
rect 21688 5028 21704 5092
rect 21768 5028 21784 5092
rect 21848 5028 21864 5092
rect 21928 5028 22070 5092
rect 22134 5028 22150 5092
rect 22214 5028 22230 5092
rect 22294 5028 22310 5092
rect 22374 5028 22390 5092
rect 22454 5028 22470 5092
rect 22534 5028 22676 5092
rect 22740 5028 22756 5092
rect 22820 5028 22836 5092
rect 22900 5028 22916 5092
rect 22980 5028 22996 5092
rect 23060 5028 23076 5092
rect 23140 5028 23282 5092
rect 23346 5028 23362 5092
rect 23426 5028 23442 5092
rect 23506 5028 23522 5092
rect 23586 5028 23602 5092
rect 23666 5028 23682 5092
rect 23746 5028 23888 5092
rect 23952 5028 23968 5092
rect 24032 5028 24048 5092
rect 24112 5028 24128 5092
rect 24192 5028 24208 5092
rect 24272 5028 24288 5092
rect 24352 5028 24494 5092
rect 24558 5028 24574 5092
rect 24638 5028 24654 5092
rect 24718 5028 24734 5092
rect 24798 5028 24814 5092
rect 24878 5028 24894 5092
rect 24958 5028 25100 5092
rect 25164 5028 25180 5092
rect 25244 5028 25260 5092
rect 25324 5028 25340 5092
rect 25404 5028 25420 5092
rect 25484 5028 25500 5092
rect 25564 5028 25706 5092
rect 25770 5028 25786 5092
rect 25850 5028 25866 5092
rect 25930 5028 25946 5092
rect 26010 5028 26026 5092
rect 26090 5028 26106 5092
rect 26170 5028 26312 5092
rect 26376 5028 26392 5092
rect 26456 5028 26472 5092
rect 26536 5028 26552 5092
rect 26616 5028 26632 5092
rect 26696 5028 26712 5092
rect 26776 5028 26918 5092
rect 26982 5028 26998 5092
rect 27062 5028 27078 5092
rect 27142 5028 27158 5092
rect 27222 5028 27238 5092
rect 27302 5028 27318 5092
rect 27382 5028 27524 5092
rect 27588 5028 27604 5092
rect 27668 5028 27684 5092
rect 27748 5028 27764 5092
rect 27828 5028 27844 5092
rect 27908 5028 27924 5092
rect 27988 5028 28130 5092
rect 28194 5028 28210 5092
rect 28274 5028 28290 5092
rect 28354 5028 28370 5092
rect 28434 5028 28450 5092
rect 28514 5028 28530 5092
rect 28594 5028 28736 5092
rect 28800 5028 28816 5092
rect 28880 5028 28896 5092
rect 28960 5028 28976 5092
rect 29040 5028 29056 5092
rect 29120 5028 29136 5092
rect 29200 5028 29342 5092
rect 29406 5028 29422 5092
rect 29486 5028 29502 5092
rect 29566 5028 29582 5092
rect 29646 5028 29662 5092
rect 29726 5028 29742 5092
rect 29806 5028 29948 5092
rect 30012 5028 30028 5092
rect 30092 5028 30108 5092
rect 30172 5028 30188 5092
rect 30252 5028 30268 5092
rect 30332 5028 30348 5092
rect 30412 5028 30554 5092
rect 30618 5028 30634 5092
rect 30698 5028 30714 5092
rect 30778 5028 30794 5092
rect 30858 5028 30874 5092
rect 30938 5028 30954 5092
rect 31018 5028 31160 5092
rect 31224 5028 31240 5092
rect 31304 5028 31320 5092
rect 31384 5028 31400 5092
rect 31464 5028 31480 5092
rect 31544 5028 31560 5092
rect 31624 5028 31766 5092
rect 31830 5028 31846 5092
rect 31910 5028 31926 5092
rect 31990 5028 32006 5092
rect 32070 5028 32086 5092
rect 32150 5028 32166 5092
rect 32230 5028 32372 5092
rect 32436 5028 32452 5092
rect 32516 5028 32532 5092
rect 32596 5028 32612 5092
rect 32676 5028 32692 5092
rect 32756 5028 32772 5092
rect 32836 5028 32978 5092
rect 33042 5028 33058 5092
rect 33122 5028 33138 5092
rect 33202 5028 33218 5092
rect 33282 5028 33298 5092
rect 33362 5028 33378 5092
rect 33442 5028 33584 5092
rect 33648 5028 33664 5092
rect 33728 5028 33744 5092
rect 33808 5028 33824 5092
rect 33888 5028 33904 5092
rect 33968 5028 33984 5092
rect 34048 5028 34190 5092
rect 34254 5028 34270 5092
rect 34334 5028 34350 5092
rect 34414 5028 34430 5092
rect 34494 5028 34510 5092
rect 34574 5028 34590 5092
rect 34654 5028 34796 5092
rect 34860 5028 34876 5092
rect 34940 5028 34956 5092
rect 35020 5028 35036 5092
rect 35100 5028 35116 5092
rect 35180 5028 35196 5092
rect 35260 5028 35402 5092
rect 35466 5028 35482 5092
rect 35546 5028 35562 5092
rect 35626 5028 35642 5092
rect 35706 5028 35722 5092
rect 35786 5028 35802 5092
rect 35866 5028 36008 5092
rect 36072 5028 36088 5092
rect 36152 5028 36168 5092
rect 36232 5028 36248 5092
rect 36312 5028 36328 5092
rect 36392 5028 36408 5092
rect 36472 5028 36614 5092
rect 36678 5028 36694 5092
rect 36758 5028 36774 5092
rect 36838 5028 36854 5092
rect 36918 5028 36934 5092
rect 36998 5028 37014 5092
rect 37078 5028 37220 5092
rect 37284 5028 37300 5092
rect 37364 5028 37380 5092
rect 37444 5028 37460 5092
rect 37524 5028 37540 5092
rect 37604 5028 37620 5092
rect 37684 5028 37826 5092
rect 37890 5028 37906 5092
rect 37970 5028 37986 5092
rect 38050 5028 38066 5092
rect 38130 5028 38146 5092
rect 38210 5028 38226 5092
rect 38290 5028 38432 5092
rect 38496 5028 38512 5092
rect 38576 5028 38592 5092
rect 38656 5028 38672 5092
rect 38736 5028 38752 5092
rect 38816 5028 38832 5092
rect 38896 5028 39038 5092
rect 39102 5028 39118 5092
rect 39182 5028 39198 5092
rect 39262 5028 39278 5092
rect 20148 5026 39298 5028
rect 39534 5026 39606 5094
rect -459 4872 -393 5026
rect -459 4808 -458 4872
rect -394 4808 -393 4872
rect -459 4792 -393 4808
rect -459 4728 -458 4792
rect -394 4728 -393 4792
rect -459 4712 -393 4728
rect -459 4648 -458 4712
rect -394 4648 -393 4712
rect -459 4632 -393 4648
rect -459 4568 -458 4632
rect -394 4568 -393 4632
rect -459 4552 -393 4568
rect -459 4488 -458 4552
rect -394 4488 -393 4552
rect -459 4472 -393 4488
rect -459 4408 -458 4472
rect -394 4408 -393 4472
rect -459 4392 -393 4408
rect -459 4328 -458 4392
rect -394 4328 -393 4392
rect -459 4312 -393 4328
rect -459 4248 -458 4312
rect -394 4248 -393 4312
rect -459 4232 -393 4248
rect -459 4168 -458 4232
rect -394 4168 -393 4232
rect -459 4152 -393 4168
rect -459 4088 -458 4152
rect -394 4088 -393 4152
rect -459 3998 -393 4088
rect -333 3994 -273 5026
rect -213 3934 -153 4964
rect -93 3994 -33 5026
rect 27 3934 87 4964
rect 147 4872 213 5026
rect 147 4808 148 4872
rect 212 4808 213 4872
rect 147 4792 213 4808
rect 147 4728 148 4792
rect 212 4728 213 4792
rect 147 4712 213 4728
rect 147 4648 148 4712
rect 212 4648 213 4712
rect 147 4632 213 4648
rect 147 4568 148 4632
rect 212 4568 213 4632
rect 147 4552 213 4568
rect 147 4488 148 4552
rect 212 4488 213 4552
rect 147 4472 213 4488
rect 147 4408 148 4472
rect 212 4408 213 4472
rect 147 4392 213 4408
rect 147 4328 148 4392
rect 212 4328 213 4392
rect 147 4312 213 4328
rect 147 4248 148 4312
rect 212 4248 213 4312
rect 147 4232 213 4248
rect 147 4168 148 4232
rect 212 4168 213 4232
rect 147 4152 213 4168
rect 147 4088 148 4152
rect 212 4088 213 4152
rect 147 3998 213 4088
rect 355 4872 421 4962
rect 355 4808 356 4872
rect 420 4808 421 4872
rect 355 4792 421 4808
rect 355 4728 356 4792
rect 420 4728 421 4792
rect 355 4712 421 4728
rect 355 4648 356 4712
rect 420 4648 421 4712
rect 355 4632 421 4648
rect 355 4568 356 4632
rect 420 4568 421 4632
rect 355 4552 421 4568
rect 355 4488 356 4552
rect 420 4488 421 4552
rect 355 4472 421 4488
rect 355 4408 356 4472
rect 420 4408 421 4472
rect 355 4392 421 4408
rect 355 4328 356 4392
rect 420 4328 421 4392
rect 355 4312 421 4328
rect 355 4248 356 4312
rect 420 4248 421 4312
rect 355 4232 421 4248
rect 355 4168 356 4232
rect 420 4168 421 4232
rect 355 4152 421 4168
rect 355 4088 356 4152
rect 420 4088 421 4152
rect 150 3994 210 3998
rect 355 3934 421 4088
rect 481 3996 541 5026
rect 601 3934 661 4966
rect 721 3996 781 5026
rect 841 3934 901 4966
rect 961 4872 1027 4962
rect 961 4808 962 4872
rect 1026 4808 1027 4872
rect 961 4792 1027 4808
rect 961 4728 962 4792
rect 1026 4728 1027 4792
rect 961 4712 1027 4728
rect 961 4648 962 4712
rect 1026 4648 1027 4712
rect 961 4632 1027 4648
rect 961 4568 962 4632
rect 1026 4568 1027 4632
rect 961 4552 1027 4568
rect 961 4488 962 4552
rect 1026 4488 1027 4552
rect 961 4472 1027 4488
rect 961 4408 962 4472
rect 1026 4408 1027 4472
rect 961 4392 1027 4408
rect 961 4328 962 4392
rect 1026 4328 1027 4392
rect 961 4312 1027 4328
rect 961 4248 962 4312
rect 1026 4248 1027 4312
rect 961 4232 1027 4248
rect 961 4168 962 4232
rect 1026 4168 1027 4232
rect 961 4152 1027 4168
rect 961 4088 962 4152
rect 1026 4088 1027 4152
rect 961 3934 1027 4088
rect -459 3932 213 3934
rect -459 3868 -355 3932
rect -291 3868 -275 3932
rect -211 3868 -195 3932
rect -131 3868 -115 3932
rect -51 3868 -35 3932
rect 29 3868 45 3932
rect 109 3868 213 3932
rect -459 3866 213 3868
rect 355 3932 1027 3934
rect 355 3868 459 3932
rect 523 3868 539 3932
rect 603 3868 619 3932
rect 683 3868 699 3932
rect 763 3868 779 3932
rect 843 3868 859 3932
rect 923 3868 1027 3932
rect 355 3866 1027 3868
rect -459 3712 -393 3802
rect -459 3648 -458 3712
rect -394 3648 -393 3712
rect -459 3632 -393 3648
rect -459 3568 -458 3632
rect -394 3568 -393 3632
rect -459 3552 -393 3568
rect -459 3488 -458 3552
rect -394 3488 -393 3552
rect -459 3472 -393 3488
rect -459 3408 -458 3472
rect -394 3408 -393 3472
rect -459 3392 -393 3408
rect -459 3328 -458 3392
rect -394 3328 -393 3392
rect -459 3312 -393 3328
rect -459 3248 -458 3312
rect -394 3248 -393 3312
rect -459 3232 -393 3248
rect -459 3168 -458 3232
rect -394 3168 -393 3232
rect -459 3152 -393 3168
rect -459 3088 -458 3152
rect -394 3088 -393 3152
rect -459 3072 -393 3088
rect -459 3008 -458 3072
rect -394 3008 -393 3072
rect -459 2992 -393 3008
rect -459 2928 -458 2992
rect -394 2928 -393 2992
rect -459 2774 -393 2928
rect -333 2836 -273 3866
rect -213 2774 -153 3806
rect -93 2836 -33 3866
rect 27 2774 87 3806
rect 147 3712 213 3802
rect 147 3648 148 3712
rect 212 3648 213 3712
rect 147 3632 213 3648
rect 147 3568 148 3632
rect 212 3568 213 3632
rect 147 3552 213 3568
rect 147 3488 148 3552
rect 212 3488 213 3552
rect 147 3472 213 3488
rect 147 3408 148 3472
rect 212 3408 213 3472
rect 147 3392 213 3408
rect 147 3328 148 3392
rect 212 3328 213 3392
rect 147 3312 213 3328
rect 147 3248 148 3312
rect 212 3248 213 3312
rect 147 3232 213 3248
rect 147 3168 148 3232
rect 212 3168 213 3232
rect 147 3152 213 3168
rect 147 3088 148 3152
rect 212 3088 213 3152
rect 147 3072 213 3088
rect 147 3008 148 3072
rect 212 3008 213 3072
rect 147 2992 213 3008
rect 147 2928 148 2992
rect 212 2928 213 2992
rect 147 2774 213 2928
rect 355 3712 421 3866
rect 355 3648 356 3712
rect 420 3648 421 3712
rect 355 3632 421 3648
rect 355 3568 356 3632
rect 420 3568 421 3632
rect 355 3552 421 3568
rect 355 3488 356 3552
rect 420 3488 421 3552
rect 355 3472 421 3488
rect 355 3408 356 3472
rect 420 3408 421 3472
rect 355 3392 421 3408
rect 355 3328 356 3392
rect 420 3328 421 3392
rect 355 3312 421 3328
rect 355 3248 356 3312
rect 420 3248 421 3312
rect 355 3232 421 3248
rect 355 3168 356 3232
rect 420 3168 421 3232
rect 355 3152 421 3168
rect 355 3088 356 3152
rect 420 3088 421 3152
rect 355 3072 421 3088
rect 355 3008 356 3072
rect 420 3008 421 3072
rect 355 2992 421 3008
rect 355 2928 356 2992
rect 420 2928 421 2992
rect 355 2838 421 2928
rect 481 2834 541 3866
rect 601 2774 661 3804
rect 721 2834 781 3866
rect 841 2774 901 3804
rect 961 3712 1027 3866
rect 961 3648 962 3712
rect 1026 3648 1027 3712
rect 961 3632 1027 3648
rect 961 3568 962 3632
rect 1026 3568 1027 3632
rect 961 3552 1027 3568
rect 961 3488 962 3552
rect 1026 3488 1027 3552
rect 961 3472 1027 3488
rect 961 3408 962 3472
rect 1026 3408 1027 3472
rect 961 3392 1027 3408
rect 961 3328 962 3392
rect 1026 3328 1027 3392
rect 961 3312 1027 3328
rect 961 3248 962 3312
rect 1026 3248 1027 3312
rect 961 3232 1027 3248
rect 961 3168 962 3232
rect 1026 3168 1027 3232
rect 961 3152 1027 3168
rect 961 3088 962 3152
rect 1026 3088 1027 3152
rect 961 3072 1027 3088
rect 961 3008 962 3072
rect 1026 3008 1027 3072
rect 961 2992 1027 3008
rect 961 2928 962 2992
rect 1026 2928 1027 2992
rect 961 2838 1027 2928
rect 1267 4872 1333 4962
rect 1267 4808 1268 4872
rect 1332 4808 1333 4872
rect 1267 4792 1333 4808
rect 1267 4728 1268 4792
rect 1332 4728 1333 4792
rect 1267 4712 1333 4728
rect 1267 4648 1268 4712
rect 1332 4648 1333 4712
rect 1267 4632 1333 4648
rect 1267 4568 1268 4632
rect 1332 4568 1333 4632
rect 1267 4552 1333 4568
rect 1267 4488 1268 4552
rect 1332 4488 1333 4552
rect 1267 4472 1333 4488
rect 1267 4408 1268 4472
rect 1332 4408 1333 4472
rect 1267 4392 1333 4408
rect 1267 4328 1268 4392
rect 1332 4328 1333 4392
rect 1267 4312 1333 4328
rect 1267 4248 1268 4312
rect 1332 4248 1333 4312
rect 1267 4232 1333 4248
rect 1267 4168 1268 4232
rect 1332 4168 1333 4232
rect 1267 4152 1333 4168
rect 1267 4088 1268 4152
rect 1332 4088 1333 4152
rect 1267 3934 1333 4088
rect 1393 3996 1453 5026
rect 1513 3934 1573 4966
rect 1633 3996 1693 5026
rect 1753 3934 1813 4966
rect 1873 4872 1939 4962
rect 1873 4808 1874 4872
rect 1938 4808 1939 4872
rect 1873 4792 1939 4808
rect 1873 4728 1874 4792
rect 1938 4728 1939 4792
rect 1873 4712 1939 4728
rect 1873 4648 1874 4712
rect 1938 4648 1939 4712
rect 1873 4632 1939 4648
rect 1873 4568 1874 4632
rect 1938 4568 1939 4632
rect 1873 4552 1939 4568
rect 1873 4488 1874 4552
rect 1938 4488 1939 4552
rect 1873 4472 1939 4488
rect 1873 4408 1874 4472
rect 1938 4408 1939 4472
rect 1873 4392 1939 4408
rect 1873 4328 1874 4392
rect 1938 4328 1939 4392
rect 1873 4312 1939 4328
rect 1873 4248 1874 4312
rect 1938 4248 1939 4312
rect 1873 4232 1939 4248
rect 1873 4168 1874 4232
rect 1938 4168 1939 4232
rect 1873 4152 1939 4168
rect 1873 4088 1874 4152
rect 1938 4088 1939 4152
rect 1873 3934 1939 4088
rect 1999 3996 2059 5026
rect 2119 3934 2179 4966
rect 2239 3996 2299 5026
rect 2359 3934 2419 4966
rect 2479 4872 2545 4962
rect 2479 4808 2480 4872
rect 2544 4808 2545 4872
rect 2479 4792 2545 4808
rect 2479 4728 2480 4792
rect 2544 4728 2545 4792
rect 2479 4712 2545 4728
rect 2479 4648 2480 4712
rect 2544 4648 2545 4712
rect 2479 4632 2545 4648
rect 2479 4568 2480 4632
rect 2544 4568 2545 4632
rect 2479 4552 2545 4568
rect 2479 4488 2480 4552
rect 2544 4488 2545 4552
rect 2479 4472 2545 4488
rect 2479 4408 2480 4472
rect 2544 4408 2545 4472
rect 2479 4392 2545 4408
rect 2479 4328 2480 4392
rect 2544 4328 2545 4392
rect 2479 4312 2545 4328
rect 2479 4248 2480 4312
rect 2544 4248 2545 4312
rect 2479 4232 2545 4248
rect 2479 4168 2480 4232
rect 2544 4168 2545 4232
rect 2479 4152 2545 4168
rect 2479 4088 2480 4152
rect 2544 4088 2545 4152
rect 2479 3934 2545 4088
rect 1267 3932 2545 3934
rect 1267 3868 1371 3932
rect 1435 3868 1451 3932
rect 1515 3868 1531 3932
rect 1595 3868 1611 3932
rect 1675 3868 1691 3932
rect 1755 3868 1771 3932
rect 1835 3868 1977 3932
rect 2041 3868 2057 3932
rect 2121 3868 2137 3932
rect 2201 3868 2217 3932
rect 2281 3868 2297 3932
rect 2361 3868 2377 3932
rect 2441 3868 2545 3932
rect 1267 3866 2545 3868
rect 1267 3712 1333 3866
rect 1267 3648 1268 3712
rect 1332 3648 1333 3712
rect 1267 3632 1333 3648
rect 1267 3568 1268 3632
rect 1332 3568 1333 3632
rect 1267 3552 1333 3568
rect 1267 3488 1268 3552
rect 1332 3488 1333 3552
rect 1267 3472 1333 3488
rect 1267 3408 1268 3472
rect 1332 3408 1333 3472
rect 1267 3392 1333 3408
rect 1267 3328 1268 3392
rect 1332 3328 1333 3392
rect 1267 3312 1333 3328
rect 1267 3248 1268 3312
rect 1332 3248 1333 3312
rect 1267 3232 1333 3248
rect 1267 3168 1268 3232
rect 1332 3168 1333 3232
rect 1267 3152 1333 3168
rect 1267 3088 1268 3152
rect 1332 3088 1333 3152
rect 1267 3072 1333 3088
rect 1267 3008 1268 3072
rect 1332 3008 1333 3072
rect 1267 2992 1333 3008
rect 1267 2928 1268 2992
rect 1332 2928 1333 2992
rect 1267 2838 1333 2928
rect 1393 2834 1453 3866
rect 1513 2774 1573 3804
rect 1633 2834 1693 3866
rect 1753 2774 1813 3804
rect 1873 3712 1939 3866
rect 1873 3648 1874 3712
rect 1938 3648 1939 3712
rect 1873 3632 1939 3648
rect 1873 3568 1874 3632
rect 1938 3568 1939 3632
rect 1873 3552 1939 3568
rect 1873 3488 1874 3552
rect 1938 3488 1939 3552
rect 1873 3472 1939 3488
rect 1873 3408 1874 3472
rect 1938 3408 1939 3472
rect 1873 3392 1939 3408
rect 1873 3328 1874 3392
rect 1938 3328 1939 3392
rect 1873 3312 1939 3328
rect 1873 3248 1874 3312
rect 1938 3248 1939 3312
rect 1873 3232 1939 3248
rect 1873 3168 1874 3232
rect 1938 3168 1939 3232
rect 1873 3152 1939 3168
rect 1873 3088 1874 3152
rect 1938 3088 1939 3152
rect 1873 3072 1939 3088
rect 1873 3008 1874 3072
rect 1938 3008 1939 3072
rect 1873 2992 1939 3008
rect 1873 2928 1874 2992
rect 1938 2928 1939 2992
rect 1873 2838 1939 2928
rect 1999 2834 2059 3866
rect 2119 2774 2179 3804
rect 2239 2834 2299 3866
rect 2359 2774 2419 3804
rect 2479 3712 2545 3866
rect 2479 3648 2480 3712
rect 2544 3648 2545 3712
rect 2479 3632 2545 3648
rect 2479 3568 2480 3632
rect 2544 3568 2545 3632
rect 2479 3552 2545 3568
rect 2479 3488 2480 3552
rect 2544 3488 2545 3552
rect 2479 3472 2545 3488
rect 2479 3408 2480 3472
rect 2544 3408 2545 3472
rect 2479 3392 2545 3408
rect 2479 3328 2480 3392
rect 2544 3328 2545 3392
rect 2479 3312 2545 3328
rect 2479 3248 2480 3312
rect 2544 3248 2545 3312
rect 2479 3232 2545 3248
rect 2479 3168 2480 3232
rect 2544 3168 2545 3232
rect 2479 3152 2545 3168
rect 2479 3088 2480 3152
rect 2544 3088 2545 3152
rect 2479 3072 2545 3088
rect 2479 3008 2480 3072
rect 2544 3008 2545 3072
rect 2479 2992 2545 3008
rect 2479 2928 2480 2992
rect 2544 2928 2545 2992
rect 2479 2838 2545 2928
rect 2801 4872 2867 4962
rect 2801 4808 2802 4872
rect 2866 4808 2867 4872
rect 2801 4792 2867 4808
rect 2801 4728 2802 4792
rect 2866 4728 2867 4792
rect 2801 4712 2867 4728
rect 2801 4648 2802 4712
rect 2866 4648 2867 4712
rect 2801 4632 2867 4648
rect 2801 4568 2802 4632
rect 2866 4568 2867 4632
rect 2801 4552 2867 4568
rect 2801 4488 2802 4552
rect 2866 4488 2867 4552
rect 2801 4472 2867 4488
rect 2801 4408 2802 4472
rect 2866 4408 2867 4472
rect 2801 4392 2867 4408
rect 2801 4328 2802 4392
rect 2866 4328 2867 4392
rect 2801 4312 2867 4328
rect 2801 4248 2802 4312
rect 2866 4248 2867 4312
rect 2801 4232 2867 4248
rect 2801 4168 2802 4232
rect 2866 4168 2867 4232
rect 2801 4152 2867 4168
rect 2801 4088 2802 4152
rect 2866 4088 2867 4152
rect 2801 3934 2867 4088
rect 2927 3996 2987 5026
rect 3047 3934 3107 4966
rect 3167 3996 3227 5026
rect 3287 3934 3347 4966
rect 3407 4872 3473 4962
rect 3407 4808 3408 4872
rect 3472 4808 3473 4872
rect 3407 4792 3473 4808
rect 3407 4728 3408 4792
rect 3472 4728 3473 4792
rect 3407 4712 3473 4728
rect 3407 4648 3408 4712
rect 3472 4648 3473 4712
rect 3407 4632 3473 4648
rect 3407 4568 3408 4632
rect 3472 4568 3473 4632
rect 3407 4552 3473 4568
rect 3407 4488 3408 4552
rect 3472 4488 3473 4552
rect 3407 4472 3473 4488
rect 3407 4408 3408 4472
rect 3472 4408 3473 4472
rect 3407 4392 3473 4408
rect 3407 4328 3408 4392
rect 3472 4328 3473 4392
rect 3407 4312 3473 4328
rect 3407 4248 3408 4312
rect 3472 4248 3473 4312
rect 3407 4232 3473 4248
rect 3407 4168 3408 4232
rect 3472 4168 3473 4232
rect 3407 4152 3473 4168
rect 3407 4088 3408 4152
rect 3472 4088 3473 4152
rect 3407 3934 3473 4088
rect 3533 3996 3593 5026
rect 3653 3934 3713 4966
rect 3773 3996 3833 5026
rect 3893 3934 3953 4966
rect 4013 4872 4079 4962
rect 4013 4808 4014 4872
rect 4078 4808 4079 4872
rect 4013 4792 4079 4808
rect 4013 4728 4014 4792
rect 4078 4728 4079 4792
rect 4013 4712 4079 4728
rect 4013 4648 4014 4712
rect 4078 4648 4079 4712
rect 4013 4632 4079 4648
rect 4013 4568 4014 4632
rect 4078 4568 4079 4632
rect 4013 4552 4079 4568
rect 4013 4488 4014 4552
rect 4078 4488 4079 4552
rect 4013 4472 4079 4488
rect 4013 4408 4014 4472
rect 4078 4408 4079 4472
rect 4013 4392 4079 4408
rect 4013 4328 4014 4392
rect 4078 4328 4079 4392
rect 4013 4312 4079 4328
rect 4013 4248 4014 4312
rect 4078 4248 4079 4312
rect 4013 4232 4079 4248
rect 4013 4168 4014 4232
rect 4078 4168 4079 4232
rect 4013 4152 4079 4168
rect 4013 4088 4014 4152
rect 4078 4088 4079 4152
rect 4013 3934 4079 4088
rect 4139 3996 4199 5026
rect 4259 3934 4319 4966
rect 4379 3996 4439 5026
rect 4499 3934 4559 4966
rect 4619 4872 4685 4962
rect 4619 4808 4620 4872
rect 4684 4808 4685 4872
rect 4619 4792 4685 4808
rect 4619 4728 4620 4792
rect 4684 4728 4685 4792
rect 4619 4712 4685 4728
rect 4619 4648 4620 4712
rect 4684 4648 4685 4712
rect 4619 4632 4685 4648
rect 4619 4568 4620 4632
rect 4684 4568 4685 4632
rect 4619 4552 4685 4568
rect 4619 4488 4620 4552
rect 4684 4488 4685 4552
rect 4619 4472 4685 4488
rect 4619 4408 4620 4472
rect 4684 4408 4685 4472
rect 4619 4392 4685 4408
rect 4619 4328 4620 4392
rect 4684 4328 4685 4392
rect 4619 4312 4685 4328
rect 4619 4248 4620 4312
rect 4684 4248 4685 4312
rect 4619 4232 4685 4248
rect 4619 4168 4620 4232
rect 4684 4168 4685 4232
rect 4619 4152 4685 4168
rect 4619 4088 4620 4152
rect 4684 4088 4685 4152
rect 4619 3934 4685 4088
rect 4745 3996 4805 5026
rect 4865 3934 4925 4966
rect 4985 3996 5045 5026
rect 5105 3934 5165 4966
rect 5225 4872 5291 4962
rect 5225 4808 5226 4872
rect 5290 4808 5291 4872
rect 5225 4792 5291 4808
rect 5225 4728 5226 4792
rect 5290 4728 5291 4792
rect 5225 4712 5291 4728
rect 5225 4648 5226 4712
rect 5290 4648 5291 4712
rect 5225 4632 5291 4648
rect 5225 4568 5226 4632
rect 5290 4568 5291 4632
rect 5225 4552 5291 4568
rect 5225 4488 5226 4552
rect 5290 4488 5291 4552
rect 5225 4472 5291 4488
rect 5225 4408 5226 4472
rect 5290 4408 5291 4472
rect 5225 4392 5291 4408
rect 5225 4328 5226 4392
rect 5290 4328 5291 4392
rect 5225 4312 5291 4328
rect 5225 4248 5226 4312
rect 5290 4248 5291 4312
rect 5225 4232 5291 4248
rect 5225 4168 5226 4232
rect 5290 4168 5291 4232
rect 5225 4152 5291 4168
rect 5225 4088 5226 4152
rect 5290 4088 5291 4152
rect 5225 3934 5291 4088
rect 2801 3932 5291 3934
rect 2801 3868 2905 3932
rect 2969 3868 2985 3932
rect 3049 3868 3065 3932
rect 3129 3868 3145 3932
rect 3209 3868 3225 3932
rect 3289 3868 3305 3932
rect 3369 3868 3511 3932
rect 3575 3868 3591 3932
rect 3655 3868 3671 3932
rect 3735 3868 3751 3932
rect 3815 3868 3831 3932
rect 3895 3868 3911 3932
rect 3975 3868 4117 3932
rect 4181 3868 4197 3932
rect 4261 3868 4277 3932
rect 4341 3868 4357 3932
rect 4421 3868 4437 3932
rect 4501 3868 4517 3932
rect 4581 3868 4723 3932
rect 4787 3868 4803 3932
rect 4867 3868 4883 3932
rect 4947 3868 4963 3932
rect 5027 3868 5043 3932
rect 5107 3868 5123 3932
rect 5187 3868 5291 3932
rect 2801 3866 5291 3868
rect 2801 3712 2867 3866
rect 2801 3648 2802 3712
rect 2866 3648 2867 3712
rect 2801 3632 2867 3648
rect 2801 3568 2802 3632
rect 2866 3568 2867 3632
rect 2801 3552 2867 3568
rect 2801 3488 2802 3552
rect 2866 3488 2867 3552
rect 2801 3472 2867 3488
rect 2801 3408 2802 3472
rect 2866 3408 2867 3472
rect 2801 3392 2867 3408
rect 2801 3328 2802 3392
rect 2866 3328 2867 3392
rect 2801 3312 2867 3328
rect 2801 3248 2802 3312
rect 2866 3248 2867 3312
rect 2801 3232 2867 3248
rect 2801 3168 2802 3232
rect 2866 3168 2867 3232
rect 2801 3152 2867 3168
rect 2801 3088 2802 3152
rect 2866 3088 2867 3152
rect 2801 3072 2867 3088
rect 2801 3008 2802 3072
rect 2866 3008 2867 3072
rect 2801 2992 2867 3008
rect 2801 2928 2802 2992
rect 2866 2928 2867 2992
rect 2801 2838 2867 2928
rect 2927 2834 2987 3866
rect 3047 2774 3107 3804
rect 3167 2834 3227 3866
rect 3287 2774 3347 3804
rect 3407 3712 3473 3866
rect 3407 3648 3408 3712
rect 3472 3648 3473 3712
rect 3407 3632 3473 3648
rect 3407 3568 3408 3632
rect 3472 3568 3473 3632
rect 3407 3552 3473 3568
rect 3407 3488 3408 3552
rect 3472 3488 3473 3552
rect 3407 3472 3473 3488
rect 3407 3408 3408 3472
rect 3472 3408 3473 3472
rect 3407 3392 3473 3408
rect 3407 3328 3408 3392
rect 3472 3328 3473 3392
rect 3407 3312 3473 3328
rect 3407 3248 3408 3312
rect 3472 3248 3473 3312
rect 3407 3232 3473 3248
rect 3407 3168 3408 3232
rect 3472 3168 3473 3232
rect 3407 3152 3473 3168
rect 3407 3088 3408 3152
rect 3472 3088 3473 3152
rect 3407 3072 3473 3088
rect 3407 3008 3408 3072
rect 3472 3008 3473 3072
rect 3407 2992 3473 3008
rect 3407 2928 3408 2992
rect 3472 2928 3473 2992
rect 3407 2838 3473 2928
rect 3533 2834 3593 3866
rect 3653 2774 3713 3804
rect 3773 2834 3833 3866
rect 3893 2774 3953 3804
rect 4013 3712 4079 3866
rect 4013 3648 4014 3712
rect 4078 3648 4079 3712
rect 4013 3632 4079 3648
rect 4013 3568 4014 3632
rect 4078 3568 4079 3632
rect 4013 3552 4079 3568
rect 4013 3488 4014 3552
rect 4078 3488 4079 3552
rect 4013 3472 4079 3488
rect 4013 3408 4014 3472
rect 4078 3408 4079 3472
rect 4013 3392 4079 3408
rect 4013 3328 4014 3392
rect 4078 3328 4079 3392
rect 4013 3312 4079 3328
rect 4013 3248 4014 3312
rect 4078 3248 4079 3312
rect 4013 3232 4079 3248
rect 4013 3168 4014 3232
rect 4078 3168 4079 3232
rect 4013 3152 4079 3168
rect 4013 3088 4014 3152
rect 4078 3088 4079 3152
rect 4013 3072 4079 3088
rect 4013 3008 4014 3072
rect 4078 3008 4079 3072
rect 4013 2992 4079 3008
rect 4013 2928 4014 2992
rect 4078 2928 4079 2992
rect 4013 2838 4079 2928
rect 4139 2834 4199 3866
rect 4259 2774 4319 3804
rect 4379 2834 4439 3866
rect 4499 2774 4559 3804
rect 4619 3712 4685 3866
rect 4619 3648 4620 3712
rect 4684 3648 4685 3712
rect 4619 3632 4685 3648
rect 4619 3568 4620 3632
rect 4684 3568 4685 3632
rect 4619 3552 4685 3568
rect 4619 3488 4620 3552
rect 4684 3488 4685 3552
rect 4619 3472 4685 3488
rect 4619 3408 4620 3472
rect 4684 3408 4685 3472
rect 4619 3392 4685 3408
rect 4619 3328 4620 3392
rect 4684 3328 4685 3392
rect 4619 3312 4685 3328
rect 4619 3248 4620 3312
rect 4684 3248 4685 3312
rect 4619 3232 4685 3248
rect 4619 3168 4620 3232
rect 4684 3168 4685 3232
rect 4619 3152 4685 3168
rect 4619 3088 4620 3152
rect 4684 3088 4685 3152
rect 4619 3072 4685 3088
rect 4619 3008 4620 3072
rect 4684 3008 4685 3072
rect 4619 2992 4685 3008
rect 4619 2928 4620 2992
rect 4684 2928 4685 2992
rect 4619 2838 4685 2928
rect 4745 2834 4805 3866
rect 4865 2774 4925 3804
rect 4985 2834 5045 3866
rect 5105 2774 5165 3804
rect 5225 3712 5291 3866
rect 5225 3648 5226 3712
rect 5290 3648 5291 3712
rect 5225 3632 5291 3648
rect 5225 3568 5226 3632
rect 5290 3568 5291 3632
rect 5225 3552 5291 3568
rect 5225 3488 5226 3552
rect 5290 3488 5291 3552
rect 5225 3472 5291 3488
rect 5225 3408 5226 3472
rect 5290 3408 5291 3472
rect 5225 3392 5291 3408
rect 5225 3328 5226 3392
rect 5290 3328 5291 3392
rect 5225 3312 5291 3328
rect 5225 3248 5226 3312
rect 5290 3248 5291 3312
rect 5225 3232 5291 3248
rect 5225 3168 5226 3232
rect 5290 3168 5291 3232
rect 5225 3152 5291 3168
rect 5225 3088 5226 3152
rect 5290 3088 5291 3152
rect 5225 3072 5291 3088
rect 5225 3008 5226 3072
rect 5290 3008 5291 3072
rect 5225 2992 5291 3008
rect 5225 2928 5226 2992
rect 5290 2928 5291 2992
rect 5225 2838 5291 2928
rect 5352 4872 5418 4962
rect 5352 4808 5353 4872
rect 5417 4808 5418 4872
rect 5352 4792 5418 4808
rect 5352 4728 5353 4792
rect 5417 4728 5418 4792
rect 5352 4712 5418 4728
rect 5352 4648 5353 4712
rect 5417 4648 5418 4712
rect 5352 4632 5418 4648
rect 5352 4568 5353 4632
rect 5417 4568 5418 4632
rect 5352 4552 5418 4568
rect 5352 4488 5353 4552
rect 5417 4488 5418 4552
rect 5352 4472 5418 4488
rect 5352 4408 5353 4472
rect 5417 4408 5418 4472
rect 5352 4392 5418 4408
rect 5352 4328 5353 4392
rect 5417 4328 5418 4392
rect 5352 4312 5418 4328
rect 5352 4248 5353 4312
rect 5417 4248 5418 4312
rect 5352 4232 5418 4248
rect 5352 4168 5353 4232
rect 5417 4168 5418 4232
rect 5352 4152 5418 4168
rect 5352 4088 5353 4152
rect 5417 4088 5418 4152
rect 5352 3934 5418 4088
rect 5478 3996 5538 5026
rect 5598 3934 5658 4966
rect 5718 3996 5778 5026
rect 5838 3934 5898 4966
rect 5958 4872 6024 4962
rect 5958 4808 5959 4872
rect 6023 4808 6024 4872
rect 5958 4792 6024 4808
rect 5958 4728 5959 4792
rect 6023 4728 6024 4792
rect 5958 4712 6024 4728
rect 5958 4648 5959 4712
rect 6023 4648 6024 4712
rect 5958 4632 6024 4648
rect 5958 4568 5959 4632
rect 6023 4568 6024 4632
rect 5958 4552 6024 4568
rect 5958 4488 5959 4552
rect 6023 4488 6024 4552
rect 5958 4472 6024 4488
rect 5958 4408 5959 4472
rect 6023 4408 6024 4472
rect 5958 4392 6024 4408
rect 5958 4328 5959 4392
rect 6023 4328 6024 4392
rect 5958 4312 6024 4328
rect 5958 4248 5959 4312
rect 6023 4248 6024 4312
rect 5958 4232 6024 4248
rect 5958 4168 5959 4232
rect 6023 4168 6024 4232
rect 5958 4152 6024 4168
rect 5958 4088 5959 4152
rect 6023 4088 6024 4152
rect 5958 3934 6024 4088
rect 6084 3996 6144 5026
rect 6204 3934 6264 4966
rect 6324 3996 6384 5026
rect 6444 3934 6504 4966
rect 6564 4872 6630 4962
rect 6564 4808 6565 4872
rect 6629 4808 6630 4872
rect 6564 4792 6630 4808
rect 6564 4728 6565 4792
rect 6629 4728 6630 4792
rect 6564 4712 6630 4728
rect 6564 4648 6565 4712
rect 6629 4648 6630 4712
rect 6564 4632 6630 4648
rect 6564 4568 6565 4632
rect 6629 4568 6630 4632
rect 6564 4552 6630 4568
rect 6564 4488 6565 4552
rect 6629 4488 6630 4552
rect 6564 4472 6630 4488
rect 6564 4408 6565 4472
rect 6629 4408 6630 4472
rect 6564 4392 6630 4408
rect 6564 4328 6565 4392
rect 6629 4328 6630 4392
rect 6564 4312 6630 4328
rect 6564 4248 6565 4312
rect 6629 4248 6630 4312
rect 6564 4232 6630 4248
rect 6564 4168 6565 4232
rect 6629 4168 6630 4232
rect 6564 4152 6630 4168
rect 6564 4088 6565 4152
rect 6629 4088 6630 4152
rect 6564 3934 6630 4088
rect 6690 3996 6750 5026
rect 6810 3934 6870 4966
rect 6930 3996 6990 5026
rect 7050 3934 7110 4966
rect 7170 4872 7236 4962
rect 7170 4808 7171 4872
rect 7235 4808 7236 4872
rect 7170 4792 7236 4808
rect 7170 4728 7171 4792
rect 7235 4728 7236 4792
rect 7170 4712 7236 4728
rect 7170 4648 7171 4712
rect 7235 4648 7236 4712
rect 7170 4632 7236 4648
rect 7170 4568 7171 4632
rect 7235 4568 7236 4632
rect 7170 4552 7236 4568
rect 7170 4488 7171 4552
rect 7235 4488 7236 4552
rect 7170 4472 7236 4488
rect 7170 4408 7171 4472
rect 7235 4408 7236 4472
rect 7170 4392 7236 4408
rect 7170 4328 7171 4392
rect 7235 4328 7236 4392
rect 7170 4312 7236 4328
rect 7170 4248 7171 4312
rect 7235 4248 7236 4312
rect 7170 4232 7236 4248
rect 7170 4168 7171 4232
rect 7235 4168 7236 4232
rect 7170 4152 7236 4168
rect 7170 4088 7171 4152
rect 7235 4088 7236 4152
rect 7170 3934 7236 4088
rect 7296 3996 7356 5026
rect 7416 3934 7476 4966
rect 7536 3996 7596 5026
rect 7656 3934 7716 4966
rect 7776 4872 7842 4962
rect 7776 4808 7777 4872
rect 7841 4808 7842 4872
rect 7776 4792 7842 4808
rect 7776 4728 7777 4792
rect 7841 4728 7842 4792
rect 7776 4712 7842 4728
rect 7776 4648 7777 4712
rect 7841 4648 7842 4712
rect 7776 4632 7842 4648
rect 7776 4568 7777 4632
rect 7841 4568 7842 4632
rect 7776 4552 7842 4568
rect 7776 4488 7777 4552
rect 7841 4488 7842 4552
rect 7776 4472 7842 4488
rect 7776 4408 7777 4472
rect 7841 4408 7842 4472
rect 7776 4392 7842 4408
rect 7776 4328 7777 4392
rect 7841 4328 7842 4392
rect 7776 4312 7842 4328
rect 7776 4248 7777 4312
rect 7841 4248 7842 4312
rect 7776 4232 7842 4248
rect 7776 4168 7777 4232
rect 7841 4168 7842 4232
rect 7776 4152 7842 4168
rect 7776 4088 7777 4152
rect 7841 4088 7842 4152
rect 7776 3934 7842 4088
rect 7902 3996 7962 5026
rect 8022 3934 8082 4966
rect 8142 3996 8202 5026
rect 8262 3934 8322 4966
rect 8382 4872 8448 4962
rect 8382 4808 8383 4872
rect 8447 4808 8448 4872
rect 8382 4792 8448 4808
rect 8382 4728 8383 4792
rect 8447 4728 8448 4792
rect 8382 4712 8448 4728
rect 8382 4648 8383 4712
rect 8447 4648 8448 4712
rect 8382 4632 8448 4648
rect 8382 4568 8383 4632
rect 8447 4568 8448 4632
rect 8382 4552 8448 4568
rect 8382 4488 8383 4552
rect 8447 4488 8448 4552
rect 8382 4472 8448 4488
rect 8382 4408 8383 4472
rect 8447 4408 8448 4472
rect 8382 4392 8448 4408
rect 8382 4328 8383 4392
rect 8447 4328 8448 4392
rect 8382 4312 8448 4328
rect 8382 4248 8383 4312
rect 8447 4248 8448 4312
rect 8382 4232 8448 4248
rect 8382 4168 8383 4232
rect 8447 4168 8448 4232
rect 8382 4152 8448 4168
rect 8382 4088 8383 4152
rect 8447 4088 8448 4152
rect 8382 3934 8448 4088
rect 8508 3996 8568 5026
rect 8628 3934 8688 4966
rect 8748 3996 8808 5026
rect 8868 3934 8928 4966
rect 8988 4872 9054 4962
rect 8988 4808 8989 4872
rect 9053 4808 9054 4872
rect 8988 4792 9054 4808
rect 8988 4728 8989 4792
rect 9053 4728 9054 4792
rect 8988 4712 9054 4728
rect 8988 4648 8989 4712
rect 9053 4648 9054 4712
rect 8988 4632 9054 4648
rect 8988 4568 8989 4632
rect 9053 4568 9054 4632
rect 8988 4552 9054 4568
rect 8988 4488 8989 4552
rect 9053 4488 9054 4552
rect 8988 4472 9054 4488
rect 8988 4408 8989 4472
rect 9053 4408 9054 4472
rect 8988 4392 9054 4408
rect 8988 4328 8989 4392
rect 9053 4328 9054 4392
rect 8988 4312 9054 4328
rect 8988 4248 8989 4312
rect 9053 4248 9054 4312
rect 8988 4232 9054 4248
rect 8988 4168 8989 4232
rect 9053 4168 9054 4232
rect 8988 4152 9054 4168
rect 8988 4088 8989 4152
rect 9053 4088 9054 4152
rect 8988 3934 9054 4088
rect 9114 3996 9174 5026
rect 9234 3934 9294 4966
rect 9354 3996 9414 5026
rect 9474 3934 9534 4966
rect 9594 4872 9660 4962
rect 9594 4808 9595 4872
rect 9659 4808 9660 4872
rect 9594 4792 9660 4808
rect 9594 4728 9595 4792
rect 9659 4728 9660 4792
rect 9594 4712 9660 4728
rect 9594 4648 9595 4712
rect 9659 4648 9660 4712
rect 9594 4632 9660 4648
rect 9594 4568 9595 4632
rect 9659 4568 9660 4632
rect 9594 4552 9660 4568
rect 9594 4488 9595 4552
rect 9659 4488 9660 4552
rect 9594 4472 9660 4488
rect 9594 4408 9595 4472
rect 9659 4408 9660 4472
rect 9594 4392 9660 4408
rect 9594 4328 9595 4392
rect 9659 4328 9660 4392
rect 9594 4312 9660 4328
rect 9594 4248 9595 4312
rect 9659 4248 9660 4312
rect 9594 4232 9660 4248
rect 9594 4168 9595 4232
rect 9659 4168 9660 4232
rect 9594 4152 9660 4168
rect 9594 4088 9595 4152
rect 9659 4088 9660 4152
rect 9594 3934 9660 4088
rect 9720 3996 9780 5026
rect 9840 3934 9900 4966
rect 9960 3996 10020 5026
rect 10080 3934 10140 4966
rect 10200 4872 10266 4962
rect 10200 4808 10201 4872
rect 10265 4808 10266 4872
rect 10200 4792 10266 4808
rect 10200 4728 10201 4792
rect 10265 4728 10266 4792
rect 10200 4712 10266 4728
rect 10200 4648 10201 4712
rect 10265 4648 10266 4712
rect 10200 4632 10266 4648
rect 10200 4568 10201 4632
rect 10265 4568 10266 4632
rect 10200 4552 10266 4568
rect 10200 4488 10201 4552
rect 10265 4488 10266 4552
rect 10200 4472 10266 4488
rect 10200 4408 10201 4472
rect 10265 4408 10266 4472
rect 10200 4392 10266 4408
rect 10200 4328 10201 4392
rect 10265 4328 10266 4392
rect 10200 4312 10266 4328
rect 10200 4248 10201 4312
rect 10265 4248 10266 4312
rect 10200 4232 10266 4248
rect 10200 4168 10201 4232
rect 10265 4168 10266 4232
rect 10200 4152 10266 4168
rect 10200 4088 10201 4152
rect 10265 4088 10266 4152
rect 10200 3934 10266 4088
rect 5352 3932 10266 3934
rect 5352 3868 5456 3932
rect 5520 3868 5536 3932
rect 5600 3868 5616 3932
rect 5680 3868 5696 3932
rect 5760 3868 5776 3932
rect 5840 3868 5856 3932
rect 5920 3868 6062 3932
rect 6126 3868 6142 3932
rect 6206 3868 6222 3932
rect 6286 3868 6302 3932
rect 6366 3868 6382 3932
rect 6446 3868 6462 3932
rect 6526 3868 6668 3932
rect 6732 3868 6748 3932
rect 6812 3868 6828 3932
rect 6892 3868 6908 3932
rect 6972 3868 6988 3932
rect 7052 3868 7068 3932
rect 7132 3868 7274 3932
rect 7338 3868 7354 3932
rect 7418 3868 7434 3932
rect 7498 3868 7514 3932
rect 7578 3868 7594 3932
rect 7658 3868 7674 3932
rect 7738 3868 7880 3932
rect 7944 3868 7960 3932
rect 8024 3868 8040 3932
rect 8104 3868 8120 3932
rect 8184 3868 8200 3932
rect 8264 3868 8280 3932
rect 8344 3868 8486 3932
rect 8550 3868 8566 3932
rect 8630 3868 8646 3932
rect 8710 3868 8726 3932
rect 8790 3868 8806 3932
rect 8870 3868 8886 3932
rect 8950 3868 9092 3932
rect 9156 3868 9172 3932
rect 9236 3868 9252 3932
rect 9316 3868 9332 3932
rect 9396 3868 9412 3932
rect 9476 3868 9492 3932
rect 9556 3868 9698 3932
rect 9762 3868 9778 3932
rect 9842 3868 9858 3932
rect 9922 3868 9938 3932
rect 10002 3868 10018 3932
rect 10082 3868 10098 3932
rect 10162 3868 10266 3932
rect 5352 3866 10266 3868
rect 5352 3712 5418 3866
rect 5352 3648 5353 3712
rect 5417 3648 5418 3712
rect 5352 3632 5418 3648
rect 5352 3568 5353 3632
rect 5417 3568 5418 3632
rect 5352 3552 5418 3568
rect 5352 3488 5353 3552
rect 5417 3488 5418 3552
rect 5352 3472 5418 3488
rect 5352 3408 5353 3472
rect 5417 3408 5418 3472
rect 5352 3392 5418 3408
rect 5352 3328 5353 3392
rect 5417 3328 5418 3392
rect 5352 3312 5418 3328
rect 5352 3248 5353 3312
rect 5417 3248 5418 3312
rect 5352 3232 5418 3248
rect 5352 3168 5353 3232
rect 5417 3168 5418 3232
rect 5352 3152 5418 3168
rect 5352 3088 5353 3152
rect 5417 3088 5418 3152
rect 5352 3072 5418 3088
rect 5352 3008 5353 3072
rect 5417 3008 5418 3072
rect 5352 2992 5418 3008
rect 5352 2928 5353 2992
rect 5417 2928 5418 2992
rect 5352 2838 5418 2928
rect 5478 2834 5538 3866
rect 5598 2774 5658 3804
rect 5718 2834 5778 3866
rect 5838 2774 5898 3804
rect 5958 3712 6024 3866
rect 5958 3648 5959 3712
rect 6023 3648 6024 3712
rect 5958 3632 6024 3648
rect 5958 3568 5959 3632
rect 6023 3568 6024 3632
rect 5958 3552 6024 3568
rect 5958 3488 5959 3552
rect 6023 3488 6024 3552
rect 5958 3472 6024 3488
rect 5958 3408 5959 3472
rect 6023 3408 6024 3472
rect 5958 3392 6024 3408
rect 5958 3328 5959 3392
rect 6023 3328 6024 3392
rect 5958 3312 6024 3328
rect 5958 3248 5959 3312
rect 6023 3248 6024 3312
rect 5958 3232 6024 3248
rect 5958 3168 5959 3232
rect 6023 3168 6024 3232
rect 5958 3152 6024 3168
rect 5958 3088 5959 3152
rect 6023 3088 6024 3152
rect 5958 3072 6024 3088
rect 5958 3008 5959 3072
rect 6023 3008 6024 3072
rect 5958 2992 6024 3008
rect 5958 2928 5959 2992
rect 6023 2928 6024 2992
rect 5958 2838 6024 2928
rect 6084 2834 6144 3866
rect 6204 2774 6264 3804
rect 6324 2834 6384 3866
rect 6444 2774 6504 3804
rect 6564 3712 6630 3866
rect 6564 3648 6565 3712
rect 6629 3648 6630 3712
rect 6564 3632 6630 3648
rect 6564 3568 6565 3632
rect 6629 3568 6630 3632
rect 6564 3552 6630 3568
rect 6564 3488 6565 3552
rect 6629 3488 6630 3552
rect 6564 3472 6630 3488
rect 6564 3408 6565 3472
rect 6629 3408 6630 3472
rect 6564 3392 6630 3408
rect 6564 3328 6565 3392
rect 6629 3328 6630 3392
rect 6564 3312 6630 3328
rect 6564 3248 6565 3312
rect 6629 3248 6630 3312
rect 6564 3232 6630 3248
rect 6564 3168 6565 3232
rect 6629 3168 6630 3232
rect 6564 3152 6630 3168
rect 6564 3088 6565 3152
rect 6629 3088 6630 3152
rect 6564 3072 6630 3088
rect 6564 3008 6565 3072
rect 6629 3008 6630 3072
rect 6564 2992 6630 3008
rect 6564 2928 6565 2992
rect 6629 2928 6630 2992
rect 6564 2838 6630 2928
rect 6690 2834 6750 3866
rect 6810 2774 6870 3804
rect 6930 2834 6990 3866
rect 7050 2774 7110 3804
rect 7170 3712 7236 3866
rect 7170 3648 7171 3712
rect 7235 3648 7236 3712
rect 7170 3632 7236 3648
rect 7170 3568 7171 3632
rect 7235 3568 7236 3632
rect 7170 3552 7236 3568
rect 7170 3488 7171 3552
rect 7235 3488 7236 3552
rect 7170 3472 7236 3488
rect 7170 3408 7171 3472
rect 7235 3408 7236 3472
rect 7170 3392 7236 3408
rect 7170 3328 7171 3392
rect 7235 3328 7236 3392
rect 7170 3312 7236 3328
rect 7170 3248 7171 3312
rect 7235 3248 7236 3312
rect 7170 3232 7236 3248
rect 7170 3168 7171 3232
rect 7235 3168 7236 3232
rect 7170 3152 7236 3168
rect 7170 3088 7171 3152
rect 7235 3088 7236 3152
rect 7170 3072 7236 3088
rect 7170 3008 7171 3072
rect 7235 3008 7236 3072
rect 7170 2992 7236 3008
rect 7170 2928 7171 2992
rect 7235 2928 7236 2992
rect 7170 2838 7236 2928
rect 7296 2834 7356 3866
rect 7416 2774 7476 3804
rect 7536 2834 7596 3866
rect 7656 2774 7716 3804
rect 7776 3712 7842 3866
rect 7776 3648 7777 3712
rect 7841 3648 7842 3712
rect 7776 3632 7842 3648
rect 7776 3568 7777 3632
rect 7841 3568 7842 3632
rect 7776 3552 7842 3568
rect 7776 3488 7777 3552
rect 7841 3488 7842 3552
rect 7776 3472 7842 3488
rect 7776 3408 7777 3472
rect 7841 3408 7842 3472
rect 7776 3392 7842 3408
rect 7776 3328 7777 3392
rect 7841 3328 7842 3392
rect 7776 3312 7842 3328
rect 7776 3248 7777 3312
rect 7841 3248 7842 3312
rect 7776 3232 7842 3248
rect 7776 3168 7777 3232
rect 7841 3168 7842 3232
rect 7776 3152 7842 3168
rect 7776 3088 7777 3152
rect 7841 3088 7842 3152
rect 7776 3072 7842 3088
rect 7776 3008 7777 3072
rect 7841 3008 7842 3072
rect 7776 2992 7842 3008
rect 7776 2928 7777 2992
rect 7841 2928 7842 2992
rect 7776 2838 7842 2928
rect 7902 2834 7962 3866
rect 8022 2774 8082 3804
rect 8142 2834 8202 3866
rect 8262 2774 8322 3804
rect 8382 3712 8448 3866
rect 8382 3648 8383 3712
rect 8447 3648 8448 3712
rect 8382 3632 8448 3648
rect 8382 3568 8383 3632
rect 8447 3568 8448 3632
rect 8382 3552 8448 3568
rect 8382 3488 8383 3552
rect 8447 3488 8448 3552
rect 8382 3472 8448 3488
rect 8382 3408 8383 3472
rect 8447 3408 8448 3472
rect 8382 3392 8448 3408
rect 8382 3328 8383 3392
rect 8447 3328 8448 3392
rect 8382 3312 8448 3328
rect 8382 3248 8383 3312
rect 8447 3248 8448 3312
rect 8382 3232 8448 3248
rect 8382 3168 8383 3232
rect 8447 3168 8448 3232
rect 8382 3152 8448 3168
rect 8382 3088 8383 3152
rect 8447 3088 8448 3152
rect 8382 3072 8448 3088
rect 8382 3008 8383 3072
rect 8447 3008 8448 3072
rect 8382 2992 8448 3008
rect 8382 2928 8383 2992
rect 8447 2928 8448 2992
rect 8382 2838 8448 2928
rect 8508 2834 8568 3866
rect 8628 2774 8688 3804
rect 8748 2834 8808 3866
rect 8868 2774 8928 3804
rect 8988 3712 9054 3866
rect 8988 3648 8989 3712
rect 9053 3648 9054 3712
rect 8988 3632 9054 3648
rect 8988 3568 8989 3632
rect 9053 3568 9054 3632
rect 8988 3552 9054 3568
rect 8988 3488 8989 3552
rect 9053 3488 9054 3552
rect 8988 3472 9054 3488
rect 8988 3408 8989 3472
rect 9053 3408 9054 3472
rect 8988 3392 9054 3408
rect 8988 3328 8989 3392
rect 9053 3328 9054 3392
rect 8988 3312 9054 3328
rect 8988 3248 8989 3312
rect 9053 3248 9054 3312
rect 8988 3232 9054 3248
rect 8988 3168 8989 3232
rect 9053 3168 9054 3232
rect 8988 3152 9054 3168
rect 8988 3088 8989 3152
rect 9053 3088 9054 3152
rect 8988 3072 9054 3088
rect 8988 3008 8989 3072
rect 9053 3008 9054 3072
rect 8988 2992 9054 3008
rect 8988 2928 8989 2992
rect 9053 2928 9054 2992
rect 8988 2838 9054 2928
rect 9114 2834 9174 3866
rect 9234 2774 9294 3804
rect 9354 2834 9414 3866
rect 9474 2774 9534 3804
rect 9594 3712 9660 3866
rect 9594 3648 9595 3712
rect 9659 3648 9660 3712
rect 9594 3632 9660 3648
rect 9594 3568 9595 3632
rect 9659 3568 9660 3632
rect 9594 3552 9660 3568
rect 9594 3488 9595 3552
rect 9659 3488 9660 3552
rect 9594 3472 9660 3488
rect 9594 3408 9595 3472
rect 9659 3408 9660 3472
rect 9594 3392 9660 3408
rect 9594 3328 9595 3392
rect 9659 3328 9660 3392
rect 9594 3312 9660 3328
rect 9594 3248 9595 3312
rect 9659 3248 9660 3312
rect 9594 3232 9660 3248
rect 9594 3168 9595 3232
rect 9659 3168 9660 3232
rect 9594 3152 9660 3168
rect 9594 3088 9595 3152
rect 9659 3088 9660 3152
rect 9594 3072 9660 3088
rect 9594 3008 9595 3072
rect 9659 3008 9660 3072
rect 9594 2992 9660 3008
rect 9594 2928 9595 2992
rect 9659 2928 9660 2992
rect 9594 2838 9660 2928
rect 9720 2834 9780 3866
rect 9840 2774 9900 3804
rect 9960 2834 10020 3866
rect 10080 2774 10140 3804
rect 10200 3712 10266 3866
rect 10200 3648 10201 3712
rect 10265 3648 10266 3712
rect 10200 3632 10266 3648
rect 10200 3568 10201 3632
rect 10265 3568 10266 3632
rect 10200 3552 10266 3568
rect 10200 3488 10201 3552
rect 10265 3488 10266 3552
rect 10200 3472 10266 3488
rect 10200 3408 10201 3472
rect 10265 3408 10266 3472
rect 10200 3392 10266 3408
rect 10200 3328 10201 3392
rect 10265 3328 10266 3392
rect 10200 3312 10266 3328
rect 10200 3248 10201 3312
rect 10265 3248 10266 3312
rect 10200 3232 10266 3248
rect 10200 3168 10201 3232
rect 10265 3168 10266 3232
rect 10200 3152 10266 3168
rect 10200 3088 10201 3152
rect 10265 3088 10266 3152
rect 10200 3072 10266 3088
rect 10200 3008 10201 3072
rect 10265 3008 10266 3072
rect 10200 2992 10266 3008
rect 10200 2928 10201 2992
rect 10265 2928 10266 2992
rect 10200 2838 10266 2928
rect 10326 4872 10392 4962
rect 10326 4808 10327 4872
rect 10391 4808 10392 4872
rect 10326 4792 10392 4808
rect 10326 4728 10327 4792
rect 10391 4728 10392 4792
rect 10326 4712 10392 4728
rect 10326 4648 10327 4712
rect 10391 4648 10392 4712
rect 10326 4632 10392 4648
rect 10326 4568 10327 4632
rect 10391 4568 10392 4632
rect 10326 4552 10392 4568
rect 10326 4488 10327 4552
rect 10391 4488 10392 4552
rect 10326 4472 10392 4488
rect 10326 4408 10327 4472
rect 10391 4408 10392 4472
rect 10326 4392 10392 4408
rect 10326 4328 10327 4392
rect 10391 4328 10392 4392
rect 10326 4312 10392 4328
rect 10326 4248 10327 4312
rect 10391 4248 10392 4312
rect 10326 4232 10392 4248
rect 10326 4168 10327 4232
rect 10391 4168 10392 4232
rect 10326 4152 10392 4168
rect 10326 4088 10327 4152
rect 10391 4088 10392 4152
rect 10326 3934 10392 4088
rect 10452 3996 10512 5026
rect 10572 3934 10632 4966
rect 10692 3996 10752 5026
rect 10812 3934 10872 4966
rect 10932 4872 10998 4962
rect 10932 4808 10933 4872
rect 10997 4808 10998 4872
rect 10932 4792 10998 4808
rect 10932 4728 10933 4792
rect 10997 4728 10998 4792
rect 10932 4712 10998 4728
rect 10932 4648 10933 4712
rect 10997 4648 10998 4712
rect 10932 4632 10998 4648
rect 10932 4568 10933 4632
rect 10997 4568 10998 4632
rect 10932 4552 10998 4568
rect 10932 4488 10933 4552
rect 10997 4488 10998 4552
rect 10932 4472 10998 4488
rect 10932 4408 10933 4472
rect 10997 4408 10998 4472
rect 10932 4392 10998 4408
rect 10932 4328 10933 4392
rect 10997 4328 10998 4392
rect 10932 4312 10998 4328
rect 10932 4248 10933 4312
rect 10997 4248 10998 4312
rect 10932 4232 10998 4248
rect 10932 4168 10933 4232
rect 10997 4168 10998 4232
rect 10932 4152 10998 4168
rect 10932 4088 10933 4152
rect 10997 4088 10998 4152
rect 10932 3934 10998 4088
rect 11058 3996 11118 5026
rect 11178 3934 11238 4966
rect 11298 3996 11358 5026
rect 11418 3934 11478 4966
rect 11538 4872 11604 4962
rect 11538 4808 11539 4872
rect 11603 4808 11604 4872
rect 11538 4792 11604 4808
rect 11538 4728 11539 4792
rect 11603 4728 11604 4792
rect 11538 4712 11604 4728
rect 11538 4648 11539 4712
rect 11603 4648 11604 4712
rect 11538 4632 11604 4648
rect 11538 4568 11539 4632
rect 11603 4568 11604 4632
rect 11538 4552 11604 4568
rect 11538 4488 11539 4552
rect 11603 4488 11604 4552
rect 11538 4472 11604 4488
rect 11538 4408 11539 4472
rect 11603 4408 11604 4472
rect 11538 4392 11604 4408
rect 11538 4328 11539 4392
rect 11603 4328 11604 4392
rect 11538 4312 11604 4328
rect 11538 4248 11539 4312
rect 11603 4248 11604 4312
rect 11538 4232 11604 4248
rect 11538 4168 11539 4232
rect 11603 4168 11604 4232
rect 11538 4152 11604 4168
rect 11538 4088 11539 4152
rect 11603 4088 11604 4152
rect 11538 3934 11604 4088
rect 11664 3996 11724 5026
rect 11784 3934 11844 4966
rect 11904 3996 11964 5026
rect 12024 3934 12084 4966
rect 12144 4872 12210 4962
rect 12144 4808 12145 4872
rect 12209 4808 12210 4872
rect 12144 4792 12210 4808
rect 12144 4728 12145 4792
rect 12209 4728 12210 4792
rect 12144 4712 12210 4728
rect 12144 4648 12145 4712
rect 12209 4648 12210 4712
rect 12144 4632 12210 4648
rect 12144 4568 12145 4632
rect 12209 4568 12210 4632
rect 12144 4552 12210 4568
rect 12144 4488 12145 4552
rect 12209 4488 12210 4552
rect 12144 4472 12210 4488
rect 12144 4408 12145 4472
rect 12209 4408 12210 4472
rect 12144 4392 12210 4408
rect 12144 4328 12145 4392
rect 12209 4328 12210 4392
rect 12144 4312 12210 4328
rect 12144 4248 12145 4312
rect 12209 4248 12210 4312
rect 12144 4232 12210 4248
rect 12144 4168 12145 4232
rect 12209 4168 12210 4232
rect 12144 4152 12210 4168
rect 12144 4088 12145 4152
rect 12209 4088 12210 4152
rect 12144 3934 12210 4088
rect 12270 3996 12330 5026
rect 12390 3934 12450 4966
rect 12510 3996 12570 5026
rect 12630 3934 12690 4966
rect 12750 4872 12816 4962
rect 12750 4808 12751 4872
rect 12815 4808 12816 4872
rect 12750 4792 12816 4808
rect 12750 4728 12751 4792
rect 12815 4728 12816 4792
rect 12750 4712 12816 4728
rect 12750 4648 12751 4712
rect 12815 4648 12816 4712
rect 12750 4632 12816 4648
rect 12750 4568 12751 4632
rect 12815 4568 12816 4632
rect 12750 4552 12816 4568
rect 12750 4488 12751 4552
rect 12815 4488 12816 4552
rect 12750 4472 12816 4488
rect 12750 4408 12751 4472
rect 12815 4408 12816 4472
rect 12750 4392 12816 4408
rect 12750 4328 12751 4392
rect 12815 4328 12816 4392
rect 12750 4312 12816 4328
rect 12750 4248 12751 4312
rect 12815 4248 12816 4312
rect 12750 4232 12816 4248
rect 12750 4168 12751 4232
rect 12815 4168 12816 4232
rect 12750 4152 12816 4168
rect 12750 4088 12751 4152
rect 12815 4088 12816 4152
rect 12750 3934 12816 4088
rect 12876 3996 12936 5026
rect 12996 3934 13056 4966
rect 13116 3996 13176 5026
rect 13236 3934 13296 4966
rect 13356 4872 13422 4962
rect 13356 4808 13357 4872
rect 13421 4808 13422 4872
rect 13356 4792 13422 4808
rect 13356 4728 13357 4792
rect 13421 4728 13422 4792
rect 13356 4712 13422 4728
rect 13356 4648 13357 4712
rect 13421 4648 13422 4712
rect 13356 4632 13422 4648
rect 13356 4568 13357 4632
rect 13421 4568 13422 4632
rect 13356 4552 13422 4568
rect 13356 4488 13357 4552
rect 13421 4488 13422 4552
rect 13356 4472 13422 4488
rect 13356 4408 13357 4472
rect 13421 4408 13422 4472
rect 13356 4392 13422 4408
rect 13356 4328 13357 4392
rect 13421 4328 13422 4392
rect 13356 4312 13422 4328
rect 13356 4248 13357 4312
rect 13421 4248 13422 4312
rect 13356 4232 13422 4248
rect 13356 4168 13357 4232
rect 13421 4168 13422 4232
rect 13356 4152 13422 4168
rect 13356 4088 13357 4152
rect 13421 4088 13422 4152
rect 13356 3934 13422 4088
rect 13482 3996 13542 5026
rect 13602 3934 13662 4966
rect 13722 3996 13782 5026
rect 13842 3934 13902 4966
rect 13962 4872 14028 4962
rect 13962 4808 13963 4872
rect 14027 4808 14028 4872
rect 13962 4792 14028 4808
rect 13962 4728 13963 4792
rect 14027 4728 14028 4792
rect 13962 4712 14028 4728
rect 13962 4648 13963 4712
rect 14027 4648 14028 4712
rect 13962 4632 14028 4648
rect 13962 4568 13963 4632
rect 14027 4568 14028 4632
rect 13962 4552 14028 4568
rect 13962 4488 13963 4552
rect 14027 4488 14028 4552
rect 13962 4472 14028 4488
rect 13962 4408 13963 4472
rect 14027 4408 14028 4472
rect 13962 4392 14028 4408
rect 13962 4328 13963 4392
rect 14027 4328 14028 4392
rect 13962 4312 14028 4328
rect 13962 4248 13963 4312
rect 14027 4248 14028 4312
rect 13962 4232 14028 4248
rect 13962 4168 13963 4232
rect 14027 4168 14028 4232
rect 13962 4152 14028 4168
rect 13962 4088 13963 4152
rect 14027 4088 14028 4152
rect 13962 3934 14028 4088
rect 14088 3996 14148 5026
rect 14208 3934 14268 4966
rect 14328 3996 14388 5026
rect 14448 3934 14508 4966
rect 14568 4872 14634 4962
rect 14568 4808 14569 4872
rect 14633 4808 14634 4872
rect 14568 4792 14634 4808
rect 14568 4728 14569 4792
rect 14633 4728 14634 4792
rect 14568 4712 14634 4728
rect 14568 4648 14569 4712
rect 14633 4648 14634 4712
rect 14568 4632 14634 4648
rect 14568 4568 14569 4632
rect 14633 4568 14634 4632
rect 14568 4552 14634 4568
rect 14568 4488 14569 4552
rect 14633 4488 14634 4552
rect 14568 4472 14634 4488
rect 14568 4408 14569 4472
rect 14633 4408 14634 4472
rect 14568 4392 14634 4408
rect 14568 4328 14569 4392
rect 14633 4328 14634 4392
rect 14568 4312 14634 4328
rect 14568 4248 14569 4312
rect 14633 4248 14634 4312
rect 14568 4232 14634 4248
rect 14568 4168 14569 4232
rect 14633 4168 14634 4232
rect 14568 4152 14634 4168
rect 14568 4088 14569 4152
rect 14633 4088 14634 4152
rect 14568 3934 14634 4088
rect 14694 3996 14754 5026
rect 14814 3934 14874 4966
rect 14934 3996 14994 5026
rect 15054 3934 15114 4966
rect 15174 4872 15240 4962
rect 15174 4808 15175 4872
rect 15239 4808 15240 4872
rect 15174 4792 15240 4808
rect 15174 4728 15175 4792
rect 15239 4728 15240 4792
rect 15174 4712 15240 4728
rect 15174 4648 15175 4712
rect 15239 4648 15240 4712
rect 15174 4632 15240 4648
rect 15174 4568 15175 4632
rect 15239 4568 15240 4632
rect 15174 4552 15240 4568
rect 15174 4488 15175 4552
rect 15239 4488 15240 4552
rect 15174 4472 15240 4488
rect 15174 4408 15175 4472
rect 15239 4408 15240 4472
rect 15174 4392 15240 4408
rect 15174 4328 15175 4392
rect 15239 4328 15240 4392
rect 15174 4312 15240 4328
rect 15174 4248 15175 4312
rect 15239 4248 15240 4312
rect 15174 4232 15240 4248
rect 15174 4168 15175 4232
rect 15239 4168 15240 4232
rect 15174 4152 15240 4168
rect 15174 4088 15175 4152
rect 15239 4088 15240 4152
rect 15174 3934 15240 4088
rect 15300 3996 15360 5026
rect 15420 3934 15480 4966
rect 15540 3996 15600 5026
rect 15660 3934 15720 4966
rect 15780 4872 15846 4962
rect 15780 4808 15781 4872
rect 15845 4808 15846 4872
rect 15780 4792 15846 4808
rect 15780 4728 15781 4792
rect 15845 4728 15846 4792
rect 15780 4712 15846 4728
rect 15780 4648 15781 4712
rect 15845 4648 15846 4712
rect 15780 4632 15846 4648
rect 15780 4568 15781 4632
rect 15845 4568 15846 4632
rect 15780 4552 15846 4568
rect 15780 4488 15781 4552
rect 15845 4488 15846 4552
rect 15780 4472 15846 4488
rect 15780 4408 15781 4472
rect 15845 4408 15846 4472
rect 15780 4392 15846 4408
rect 15780 4328 15781 4392
rect 15845 4328 15846 4392
rect 15780 4312 15846 4328
rect 15780 4248 15781 4312
rect 15845 4248 15846 4312
rect 15780 4232 15846 4248
rect 15780 4168 15781 4232
rect 15845 4168 15846 4232
rect 15780 4152 15846 4168
rect 15780 4088 15781 4152
rect 15845 4088 15846 4152
rect 15780 3934 15846 4088
rect 15906 3996 15966 5026
rect 16026 3934 16086 4966
rect 16146 3996 16206 5026
rect 16266 3934 16326 4966
rect 16386 4872 16452 4962
rect 16386 4808 16387 4872
rect 16451 4808 16452 4872
rect 16386 4792 16452 4808
rect 16386 4728 16387 4792
rect 16451 4728 16452 4792
rect 16386 4712 16452 4728
rect 16386 4648 16387 4712
rect 16451 4648 16452 4712
rect 16386 4632 16452 4648
rect 16386 4568 16387 4632
rect 16451 4568 16452 4632
rect 16386 4552 16452 4568
rect 16386 4488 16387 4552
rect 16451 4488 16452 4552
rect 16386 4472 16452 4488
rect 16386 4408 16387 4472
rect 16451 4408 16452 4472
rect 16386 4392 16452 4408
rect 16386 4328 16387 4392
rect 16451 4328 16452 4392
rect 16386 4312 16452 4328
rect 16386 4248 16387 4312
rect 16451 4248 16452 4312
rect 16386 4232 16452 4248
rect 16386 4168 16387 4232
rect 16451 4168 16452 4232
rect 16386 4152 16452 4168
rect 16386 4088 16387 4152
rect 16451 4088 16452 4152
rect 16386 3934 16452 4088
rect 16512 3996 16572 5026
rect 16632 3934 16692 4966
rect 16752 3996 16812 5026
rect 16872 3934 16932 4966
rect 16992 4872 17058 4962
rect 16992 4808 16993 4872
rect 17057 4808 17058 4872
rect 16992 4792 17058 4808
rect 16992 4728 16993 4792
rect 17057 4728 17058 4792
rect 16992 4712 17058 4728
rect 16992 4648 16993 4712
rect 17057 4648 17058 4712
rect 16992 4632 17058 4648
rect 16992 4568 16993 4632
rect 17057 4568 17058 4632
rect 16992 4552 17058 4568
rect 16992 4488 16993 4552
rect 17057 4488 17058 4552
rect 16992 4472 17058 4488
rect 16992 4408 16993 4472
rect 17057 4408 17058 4472
rect 16992 4392 17058 4408
rect 16992 4328 16993 4392
rect 17057 4328 17058 4392
rect 16992 4312 17058 4328
rect 16992 4248 16993 4312
rect 17057 4248 17058 4312
rect 16992 4232 17058 4248
rect 16992 4168 16993 4232
rect 17057 4168 17058 4232
rect 16992 4152 17058 4168
rect 16992 4088 16993 4152
rect 17057 4088 17058 4152
rect 16992 3934 17058 4088
rect 17118 3996 17178 5026
rect 17238 3934 17298 4966
rect 17358 3996 17418 5026
rect 17478 3934 17538 4966
rect 17598 4872 17664 4962
rect 17598 4808 17599 4872
rect 17663 4808 17664 4872
rect 17598 4792 17664 4808
rect 17598 4728 17599 4792
rect 17663 4728 17664 4792
rect 17598 4712 17664 4728
rect 17598 4648 17599 4712
rect 17663 4648 17664 4712
rect 17598 4632 17664 4648
rect 17598 4568 17599 4632
rect 17663 4568 17664 4632
rect 17598 4552 17664 4568
rect 17598 4488 17599 4552
rect 17663 4488 17664 4552
rect 17598 4472 17664 4488
rect 17598 4408 17599 4472
rect 17663 4408 17664 4472
rect 17598 4392 17664 4408
rect 17598 4328 17599 4392
rect 17663 4328 17664 4392
rect 17598 4312 17664 4328
rect 17598 4248 17599 4312
rect 17663 4248 17664 4312
rect 17598 4232 17664 4248
rect 17598 4168 17599 4232
rect 17663 4168 17664 4232
rect 17598 4152 17664 4168
rect 17598 4088 17599 4152
rect 17663 4088 17664 4152
rect 17598 3934 17664 4088
rect 17724 3996 17784 5026
rect 17844 3934 17904 4966
rect 17964 3996 18024 5026
rect 18084 3934 18144 4966
rect 18204 4872 18270 4962
rect 18204 4808 18205 4872
rect 18269 4808 18270 4872
rect 18204 4792 18270 4808
rect 18204 4728 18205 4792
rect 18269 4728 18270 4792
rect 18204 4712 18270 4728
rect 18204 4648 18205 4712
rect 18269 4648 18270 4712
rect 18204 4632 18270 4648
rect 18204 4568 18205 4632
rect 18269 4568 18270 4632
rect 18204 4552 18270 4568
rect 18204 4488 18205 4552
rect 18269 4488 18270 4552
rect 18204 4472 18270 4488
rect 18204 4408 18205 4472
rect 18269 4408 18270 4472
rect 18204 4392 18270 4408
rect 18204 4328 18205 4392
rect 18269 4328 18270 4392
rect 18204 4312 18270 4328
rect 18204 4248 18205 4312
rect 18269 4248 18270 4312
rect 18204 4232 18270 4248
rect 18204 4168 18205 4232
rect 18269 4168 18270 4232
rect 18204 4152 18270 4168
rect 18204 4088 18205 4152
rect 18269 4088 18270 4152
rect 18204 3934 18270 4088
rect 18330 3996 18390 5026
rect 18450 3934 18510 4966
rect 18570 3996 18630 5026
rect 18690 3934 18750 4966
rect 18810 4872 18876 4962
rect 18810 4808 18811 4872
rect 18875 4808 18876 4872
rect 18810 4792 18876 4808
rect 18810 4728 18811 4792
rect 18875 4728 18876 4792
rect 18810 4712 18876 4728
rect 18810 4648 18811 4712
rect 18875 4648 18876 4712
rect 18810 4632 18876 4648
rect 18810 4568 18811 4632
rect 18875 4568 18876 4632
rect 18810 4552 18876 4568
rect 18810 4488 18811 4552
rect 18875 4488 18876 4552
rect 18810 4472 18876 4488
rect 18810 4408 18811 4472
rect 18875 4408 18876 4472
rect 18810 4392 18876 4408
rect 18810 4328 18811 4392
rect 18875 4328 18876 4392
rect 18810 4312 18876 4328
rect 18810 4248 18811 4312
rect 18875 4248 18876 4312
rect 18810 4232 18876 4248
rect 18810 4168 18811 4232
rect 18875 4168 18876 4232
rect 18810 4152 18876 4168
rect 18810 4088 18811 4152
rect 18875 4088 18876 4152
rect 18810 3934 18876 4088
rect 18936 3996 18996 5026
rect 19056 3934 19116 4966
rect 19176 3996 19236 5026
rect 19296 3934 19356 4966
rect 19416 4872 19482 4962
rect 19416 4808 19417 4872
rect 19481 4808 19482 4872
rect 19416 4792 19482 4808
rect 19416 4728 19417 4792
rect 19481 4728 19482 4792
rect 19416 4712 19482 4728
rect 19416 4648 19417 4712
rect 19481 4648 19482 4712
rect 19416 4632 19482 4648
rect 19416 4568 19417 4632
rect 19481 4568 19482 4632
rect 19416 4552 19482 4568
rect 19416 4488 19417 4552
rect 19481 4488 19482 4552
rect 19416 4472 19482 4488
rect 19416 4408 19417 4472
rect 19481 4408 19482 4472
rect 19416 4392 19482 4408
rect 19416 4328 19417 4392
rect 19481 4328 19482 4392
rect 19416 4312 19482 4328
rect 19416 4248 19417 4312
rect 19481 4248 19482 4312
rect 19416 4232 19482 4248
rect 19416 4168 19417 4232
rect 19481 4168 19482 4232
rect 19416 4152 19482 4168
rect 19416 4088 19417 4152
rect 19481 4088 19482 4152
rect 19416 3934 19482 4088
rect 19542 3996 19602 5026
rect 19662 3934 19722 4966
rect 19782 3996 19842 5026
rect 19902 3934 19962 4966
rect 20022 4872 20088 4962
rect 20022 4808 20023 4872
rect 20087 4808 20088 4872
rect 20022 4792 20088 4808
rect 20022 4728 20023 4792
rect 20087 4728 20088 4792
rect 20022 4712 20088 4728
rect 20022 4648 20023 4712
rect 20087 4648 20088 4712
rect 20022 4632 20088 4648
rect 20022 4568 20023 4632
rect 20087 4568 20088 4632
rect 20022 4552 20088 4568
rect 20022 4488 20023 4552
rect 20087 4488 20088 4552
rect 20022 4472 20088 4488
rect 20022 4408 20023 4472
rect 20087 4408 20088 4472
rect 20022 4392 20088 4408
rect 20022 4328 20023 4392
rect 20087 4328 20088 4392
rect 20022 4312 20088 4328
rect 20022 4248 20023 4312
rect 20087 4248 20088 4312
rect 20022 4232 20088 4248
rect 20022 4168 20023 4232
rect 20087 4168 20088 4232
rect 20022 4152 20088 4168
rect 20022 4088 20023 4152
rect 20087 4088 20088 4152
rect 20022 3934 20088 4088
rect 10326 3932 20088 3934
rect 10326 3868 10430 3932
rect 10494 3868 10510 3932
rect 10574 3868 10590 3932
rect 10654 3868 10670 3932
rect 10734 3868 10750 3932
rect 10814 3868 10830 3932
rect 10894 3868 11036 3932
rect 11100 3868 11116 3932
rect 11180 3868 11196 3932
rect 11260 3868 11276 3932
rect 11340 3868 11356 3932
rect 11420 3868 11436 3932
rect 11500 3868 11642 3932
rect 11706 3868 11722 3932
rect 11786 3868 11802 3932
rect 11866 3868 11882 3932
rect 11946 3868 11962 3932
rect 12026 3868 12042 3932
rect 12106 3868 12248 3932
rect 12312 3868 12328 3932
rect 12392 3868 12408 3932
rect 12472 3868 12488 3932
rect 12552 3868 12568 3932
rect 12632 3868 12648 3932
rect 12712 3868 12854 3932
rect 12918 3868 12934 3932
rect 12998 3868 13014 3932
rect 13078 3868 13094 3932
rect 13158 3868 13174 3932
rect 13238 3868 13254 3932
rect 13318 3868 13460 3932
rect 13524 3868 13540 3932
rect 13604 3868 13620 3932
rect 13684 3868 13700 3932
rect 13764 3868 13780 3932
rect 13844 3868 13860 3932
rect 13924 3868 14066 3932
rect 14130 3868 14146 3932
rect 14210 3868 14226 3932
rect 14290 3868 14306 3932
rect 14370 3868 14386 3932
rect 14450 3868 14466 3932
rect 14530 3868 14672 3932
rect 14736 3868 14752 3932
rect 14816 3868 14832 3932
rect 14896 3868 14912 3932
rect 14976 3868 14992 3932
rect 15056 3868 15072 3932
rect 15136 3868 15278 3932
rect 15342 3868 15358 3932
rect 15422 3868 15438 3932
rect 15502 3868 15518 3932
rect 15582 3868 15598 3932
rect 15662 3868 15678 3932
rect 15742 3868 15884 3932
rect 15948 3868 15964 3932
rect 16028 3868 16044 3932
rect 16108 3868 16124 3932
rect 16188 3868 16204 3932
rect 16268 3868 16284 3932
rect 16348 3868 16490 3932
rect 16554 3868 16570 3932
rect 16634 3868 16650 3932
rect 16714 3868 16730 3932
rect 16794 3868 16810 3932
rect 16874 3868 16890 3932
rect 16954 3868 17096 3932
rect 17160 3868 17176 3932
rect 17240 3868 17256 3932
rect 17320 3868 17336 3932
rect 17400 3868 17416 3932
rect 17480 3868 17496 3932
rect 17560 3868 17702 3932
rect 17766 3868 17782 3932
rect 17846 3868 17862 3932
rect 17926 3868 17942 3932
rect 18006 3868 18022 3932
rect 18086 3868 18102 3932
rect 18166 3868 18308 3932
rect 18372 3868 18388 3932
rect 18452 3868 18468 3932
rect 18532 3868 18548 3932
rect 18612 3868 18628 3932
rect 18692 3868 18708 3932
rect 18772 3868 18914 3932
rect 18978 3868 18994 3932
rect 19058 3868 19074 3932
rect 19138 3868 19154 3932
rect 19218 3868 19234 3932
rect 19298 3868 19314 3932
rect 19378 3868 19520 3932
rect 19584 3868 19600 3932
rect 19664 3868 19680 3932
rect 19744 3868 19760 3932
rect 19824 3868 19840 3932
rect 19904 3868 19920 3932
rect 19984 3868 20088 3932
rect 10326 3866 20088 3868
rect 10326 3712 10392 3866
rect 10326 3648 10327 3712
rect 10391 3648 10392 3712
rect 10326 3632 10392 3648
rect 10326 3568 10327 3632
rect 10391 3568 10392 3632
rect 10326 3552 10392 3568
rect 10326 3488 10327 3552
rect 10391 3488 10392 3552
rect 10326 3472 10392 3488
rect 10326 3408 10327 3472
rect 10391 3408 10392 3472
rect 10326 3392 10392 3408
rect 10326 3328 10327 3392
rect 10391 3328 10392 3392
rect 10326 3312 10392 3328
rect 10326 3248 10327 3312
rect 10391 3248 10392 3312
rect 10326 3232 10392 3248
rect 10326 3168 10327 3232
rect 10391 3168 10392 3232
rect 10326 3152 10392 3168
rect 10326 3088 10327 3152
rect 10391 3088 10392 3152
rect 10326 3072 10392 3088
rect 10326 3008 10327 3072
rect 10391 3008 10392 3072
rect 10326 2992 10392 3008
rect 10326 2928 10327 2992
rect 10391 2928 10392 2992
rect 10326 2838 10392 2928
rect 10452 2834 10512 3866
rect 10572 2774 10632 3804
rect 10692 2834 10752 3866
rect 10812 2774 10872 3804
rect 10932 3712 10998 3866
rect 10932 3648 10933 3712
rect 10997 3648 10998 3712
rect 10932 3632 10998 3648
rect 10932 3568 10933 3632
rect 10997 3568 10998 3632
rect 10932 3552 10998 3568
rect 10932 3488 10933 3552
rect 10997 3488 10998 3552
rect 10932 3472 10998 3488
rect 10932 3408 10933 3472
rect 10997 3408 10998 3472
rect 10932 3392 10998 3408
rect 10932 3328 10933 3392
rect 10997 3328 10998 3392
rect 10932 3312 10998 3328
rect 10932 3248 10933 3312
rect 10997 3248 10998 3312
rect 10932 3232 10998 3248
rect 10932 3168 10933 3232
rect 10997 3168 10998 3232
rect 10932 3152 10998 3168
rect 10932 3088 10933 3152
rect 10997 3088 10998 3152
rect 10932 3072 10998 3088
rect 10932 3008 10933 3072
rect 10997 3008 10998 3072
rect 10932 2992 10998 3008
rect 10932 2928 10933 2992
rect 10997 2928 10998 2992
rect 10932 2838 10998 2928
rect 11058 2834 11118 3866
rect 11178 2774 11238 3804
rect 11298 2834 11358 3866
rect 11418 2774 11478 3804
rect 11538 3712 11604 3866
rect 11538 3648 11539 3712
rect 11603 3648 11604 3712
rect 11538 3632 11604 3648
rect 11538 3568 11539 3632
rect 11603 3568 11604 3632
rect 11538 3552 11604 3568
rect 11538 3488 11539 3552
rect 11603 3488 11604 3552
rect 11538 3472 11604 3488
rect 11538 3408 11539 3472
rect 11603 3408 11604 3472
rect 11538 3392 11604 3408
rect 11538 3328 11539 3392
rect 11603 3328 11604 3392
rect 11538 3312 11604 3328
rect 11538 3248 11539 3312
rect 11603 3248 11604 3312
rect 11538 3232 11604 3248
rect 11538 3168 11539 3232
rect 11603 3168 11604 3232
rect 11538 3152 11604 3168
rect 11538 3088 11539 3152
rect 11603 3088 11604 3152
rect 11538 3072 11604 3088
rect 11538 3008 11539 3072
rect 11603 3008 11604 3072
rect 11538 2992 11604 3008
rect 11538 2928 11539 2992
rect 11603 2928 11604 2992
rect 11538 2838 11604 2928
rect 11664 2834 11724 3866
rect 11784 2774 11844 3804
rect 11904 2834 11964 3866
rect 12024 2774 12084 3804
rect 12144 3712 12210 3866
rect 12144 3648 12145 3712
rect 12209 3648 12210 3712
rect 12144 3632 12210 3648
rect 12144 3568 12145 3632
rect 12209 3568 12210 3632
rect 12144 3552 12210 3568
rect 12144 3488 12145 3552
rect 12209 3488 12210 3552
rect 12144 3472 12210 3488
rect 12144 3408 12145 3472
rect 12209 3408 12210 3472
rect 12144 3392 12210 3408
rect 12144 3328 12145 3392
rect 12209 3328 12210 3392
rect 12144 3312 12210 3328
rect 12144 3248 12145 3312
rect 12209 3248 12210 3312
rect 12144 3232 12210 3248
rect 12144 3168 12145 3232
rect 12209 3168 12210 3232
rect 12144 3152 12210 3168
rect 12144 3088 12145 3152
rect 12209 3088 12210 3152
rect 12144 3072 12210 3088
rect 12144 3008 12145 3072
rect 12209 3008 12210 3072
rect 12144 2992 12210 3008
rect 12144 2928 12145 2992
rect 12209 2928 12210 2992
rect 12144 2838 12210 2928
rect 12270 2834 12330 3866
rect 12390 2774 12450 3804
rect 12510 2834 12570 3866
rect 12630 2774 12690 3804
rect 12750 3712 12816 3866
rect 12750 3648 12751 3712
rect 12815 3648 12816 3712
rect 12750 3632 12816 3648
rect 12750 3568 12751 3632
rect 12815 3568 12816 3632
rect 12750 3552 12816 3568
rect 12750 3488 12751 3552
rect 12815 3488 12816 3552
rect 12750 3472 12816 3488
rect 12750 3408 12751 3472
rect 12815 3408 12816 3472
rect 12750 3392 12816 3408
rect 12750 3328 12751 3392
rect 12815 3328 12816 3392
rect 12750 3312 12816 3328
rect 12750 3248 12751 3312
rect 12815 3248 12816 3312
rect 12750 3232 12816 3248
rect 12750 3168 12751 3232
rect 12815 3168 12816 3232
rect 12750 3152 12816 3168
rect 12750 3088 12751 3152
rect 12815 3088 12816 3152
rect 12750 3072 12816 3088
rect 12750 3008 12751 3072
rect 12815 3008 12816 3072
rect 12750 2992 12816 3008
rect 12750 2928 12751 2992
rect 12815 2928 12816 2992
rect 12750 2838 12816 2928
rect 12876 2834 12936 3866
rect 12996 2774 13056 3804
rect 13116 2834 13176 3866
rect 13236 2774 13296 3804
rect 13356 3712 13422 3866
rect 13356 3648 13357 3712
rect 13421 3648 13422 3712
rect 13356 3632 13422 3648
rect 13356 3568 13357 3632
rect 13421 3568 13422 3632
rect 13356 3552 13422 3568
rect 13356 3488 13357 3552
rect 13421 3488 13422 3552
rect 13356 3472 13422 3488
rect 13356 3408 13357 3472
rect 13421 3408 13422 3472
rect 13356 3392 13422 3408
rect 13356 3328 13357 3392
rect 13421 3328 13422 3392
rect 13356 3312 13422 3328
rect 13356 3248 13357 3312
rect 13421 3248 13422 3312
rect 13356 3232 13422 3248
rect 13356 3168 13357 3232
rect 13421 3168 13422 3232
rect 13356 3152 13422 3168
rect 13356 3088 13357 3152
rect 13421 3088 13422 3152
rect 13356 3072 13422 3088
rect 13356 3008 13357 3072
rect 13421 3008 13422 3072
rect 13356 2992 13422 3008
rect 13356 2928 13357 2992
rect 13421 2928 13422 2992
rect 13356 2838 13422 2928
rect 13482 2834 13542 3866
rect 13602 2774 13662 3804
rect 13722 2834 13782 3866
rect 13842 2774 13902 3804
rect 13962 3712 14028 3866
rect 13962 3648 13963 3712
rect 14027 3648 14028 3712
rect 13962 3632 14028 3648
rect 13962 3568 13963 3632
rect 14027 3568 14028 3632
rect 13962 3552 14028 3568
rect 13962 3488 13963 3552
rect 14027 3488 14028 3552
rect 13962 3472 14028 3488
rect 13962 3408 13963 3472
rect 14027 3408 14028 3472
rect 13962 3392 14028 3408
rect 13962 3328 13963 3392
rect 14027 3328 14028 3392
rect 13962 3312 14028 3328
rect 13962 3248 13963 3312
rect 14027 3248 14028 3312
rect 13962 3232 14028 3248
rect 13962 3168 13963 3232
rect 14027 3168 14028 3232
rect 13962 3152 14028 3168
rect 13962 3088 13963 3152
rect 14027 3088 14028 3152
rect 13962 3072 14028 3088
rect 13962 3008 13963 3072
rect 14027 3008 14028 3072
rect 13962 2992 14028 3008
rect 13962 2928 13963 2992
rect 14027 2928 14028 2992
rect 13962 2838 14028 2928
rect 14088 2834 14148 3866
rect 14208 2774 14268 3804
rect 14328 2834 14388 3866
rect 14448 2774 14508 3804
rect 14568 3712 14634 3866
rect 14568 3648 14569 3712
rect 14633 3648 14634 3712
rect 14568 3632 14634 3648
rect 14568 3568 14569 3632
rect 14633 3568 14634 3632
rect 14568 3552 14634 3568
rect 14568 3488 14569 3552
rect 14633 3488 14634 3552
rect 14568 3472 14634 3488
rect 14568 3408 14569 3472
rect 14633 3408 14634 3472
rect 14568 3392 14634 3408
rect 14568 3328 14569 3392
rect 14633 3328 14634 3392
rect 14568 3312 14634 3328
rect 14568 3248 14569 3312
rect 14633 3248 14634 3312
rect 14568 3232 14634 3248
rect 14568 3168 14569 3232
rect 14633 3168 14634 3232
rect 14568 3152 14634 3168
rect 14568 3088 14569 3152
rect 14633 3088 14634 3152
rect 14568 3072 14634 3088
rect 14568 3008 14569 3072
rect 14633 3008 14634 3072
rect 14568 2992 14634 3008
rect 14568 2928 14569 2992
rect 14633 2928 14634 2992
rect 14568 2838 14634 2928
rect 14694 2834 14754 3866
rect 14814 2774 14874 3804
rect 14934 2834 14994 3866
rect 15054 2774 15114 3804
rect 15174 3712 15240 3866
rect 15174 3648 15175 3712
rect 15239 3648 15240 3712
rect 15174 3632 15240 3648
rect 15174 3568 15175 3632
rect 15239 3568 15240 3632
rect 15174 3552 15240 3568
rect 15174 3488 15175 3552
rect 15239 3488 15240 3552
rect 15174 3472 15240 3488
rect 15174 3408 15175 3472
rect 15239 3408 15240 3472
rect 15174 3392 15240 3408
rect 15174 3328 15175 3392
rect 15239 3328 15240 3392
rect 15174 3312 15240 3328
rect 15174 3248 15175 3312
rect 15239 3248 15240 3312
rect 15174 3232 15240 3248
rect 15174 3168 15175 3232
rect 15239 3168 15240 3232
rect 15174 3152 15240 3168
rect 15174 3088 15175 3152
rect 15239 3088 15240 3152
rect 15174 3072 15240 3088
rect 15174 3008 15175 3072
rect 15239 3008 15240 3072
rect 15174 2992 15240 3008
rect 15174 2928 15175 2992
rect 15239 2928 15240 2992
rect 15174 2838 15240 2928
rect 15300 2834 15360 3866
rect 15420 2774 15480 3804
rect 15540 2834 15600 3866
rect 15660 2774 15720 3804
rect 15780 3712 15846 3866
rect 15780 3648 15781 3712
rect 15845 3648 15846 3712
rect 15780 3632 15846 3648
rect 15780 3568 15781 3632
rect 15845 3568 15846 3632
rect 15780 3552 15846 3568
rect 15780 3488 15781 3552
rect 15845 3488 15846 3552
rect 15780 3472 15846 3488
rect 15780 3408 15781 3472
rect 15845 3408 15846 3472
rect 15780 3392 15846 3408
rect 15780 3328 15781 3392
rect 15845 3328 15846 3392
rect 15780 3312 15846 3328
rect 15780 3248 15781 3312
rect 15845 3248 15846 3312
rect 15780 3232 15846 3248
rect 15780 3168 15781 3232
rect 15845 3168 15846 3232
rect 15780 3152 15846 3168
rect 15780 3088 15781 3152
rect 15845 3088 15846 3152
rect 15780 3072 15846 3088
rect 15780 3008 15781 3072
rect 15845 3008 15846 3072
rect 15780 2992 15846 3008
rect 15780 2928 15781 2992
rect 15845 2928 15846 2992
rect 15780 2838 15846 2928
rect 15906 2834 15966 3866
rect 16026 2774 16086 3804
rect 16146 2834 16206 3866
rect 16266 2774 16326 3804
rect 16386 3712 16452 3866
rect 16386 3648 16387 3712
rect 16451 3648 16452 3712
rect 16386 3632 16452 3648
rect 16386 3568 16387 3632
rect 16451 3568 16452 3632
rect 16386 3552 16452 3568
rect 16386 3488 16387 3552
rect 16451 3488 16452 3552
rect 16386 3472 16452 3488
rect 16386 3408 16387 3472
rect 16451 3408 16452 3472
rect 16386 3392 16452 3408
rect 16386 3328 16387 3392
rect 16451 3328 16452 3392
rect 16386 3312 16452 3328
rect 16386 3248 16387 3312
rect 16451 3248 16452 3312
rect 16386 3232 16452 3248
rect 16386 3168 16387 3232
rect 16451 3168 16452 3232
rect 16386 3152 16452 3168
rect 16386 3088 16387 3152
rect 16451 3088 16452 3152
rect 16386 3072 16452 3088
rect 16386 3008 16387 3072
rect 16451 3008 16452 3072
rect 16386 2992 16452 3008
rect 16386 2928 16387 2992
rect 16451 2928 16452 2992
rect 16386 2838 16452 2928
rect 16512 2834 16572 3866
rect 16632 2774 16692 3804
rect 16752 2834 16812 3866
rect 16872 2774 16932 3804
rect 16992 3712 17058 3866
rect 16992 3648 16993 3712
rect 17057 3648 17058 3712
rect 16992 3632 17058 3648
rect 16992 3568 16993 3632
rect 17057 3568 17058 3632
rect 16992 3552 17058 3568
rect 16992 3488 16993 3552
rect 17057 3488 17058 3552
rect 16992 3472 17058 3488
rect 16992 3408 16993 3472
rect 17057 3408 17058 3472
rect 16992 3392 17058 3408
rect 16992 3328 16993 3392
rect 17057 3328 17058 3392
rect 16992 3312 17058 3328
rect 16992 3248 16993 3312
rect 17057 3248 17058 3312
rect 16992 3232 17058 3248
rect 16992 3168 16993 3232
rect 17057 3168 17058 3232
rect 16992 3152 17058 3168
rect 16992 3088 16993 3152
rect 17057 3088 17058 3152
rect 16992 3072 17058 3088
rect 16992 3008 16993 3072
rect 17057 3008 17058 3072
rect 16992 2992 17058 3008
rect 16992 2928 16993 2992
rect 17057 2928 17058 2992
rect 16992 2838 17058 2928
rect 17118 2834 17178 3866
rect 17238 2774 17298 3804
rect 17358 2834 17418 3866
rect 17478 2774 17538 3804
rect 17598 3712 17664 3866
rect 17598 3648 17599 3712
rect 17663 3648 17664 3712
rect 17598 3632 17664 3648
rect 17598 3568 17599 3632
rect 17663 3568 17664 3632
rect 17598 3552 17664 3568
rect 17598 3488 17599 3552
rect 17663 3488 17664 3552
rect 17598 3472 17664 3488
rect 17598 3408 17599 3472
rect 17663 3408 17664 3472
rect 17598 3392 17664 3408
rect 17598 3328 17599 3392
rect 17663 3328 17664 3392
rect 17598 3312 17664 3328
rect 17598 3248 17599 3312
rect 17663 3248 17664 3312
rect 17598 3232 17664 3248
rect 17598 3168 17599 3232
rect 17663 3168 17664 3232
rect 17598 3152 17664 3168
rect 17598 3088 17599 3152
rect 17663 3088 17664 3152
rect 17598 3072 17664 3088
rect 17598 3008 17599 3072
rect 17663 3008 17664 3072
rect 17598 2992 17664 3008
rect 17598 2928 17599 2992
rect 17663 2928 17664 2992
rect 17598 2838 17664 2928
rect 17724 2834 17784 3866
rect 17844 2774 17904 3804
rect 17964 2834 18024 3866
rect 18084 2774 18144 3804
rect 18204 3712 18270 3866
rect 18204 3648 18205 3712
rect 18269 3648 18270 3712
rect 18204 3632 18270 3648
rect 18204 3568 18205 3632
rect 18269 3568 18270 3632
rect 18204 3552 18270 3568
rect 18204 3488 18205 3552
rect 18269 3488 18270 3552
rect 18204 3472 18270 3488
rect 18204 3408 18205 3472
rect 18269 3408 18270 3472
rect 18204 3392 18270 3408
rect 18204 3328 18205 3392
rect 18269 3328 18270 3392
rect 18204 3312 18270 3328
rect 18204 3248 18205 3312
rect 18269 3248 18270 3312
rect 18204 3232 18270 3248
rect 18204 3168 18205 3232
rect 18269 3168 18270 3232
rect 18204 3152 18270 3168
rect 18204 3088 18205 3152
rect 18269 3088 18270 3152
rect 18204 3072 18270 3088
rect 18204 3008 18205 3072
rect 18269 3008 18270 3072
rect 18204 2992 18270 3008
rect 18204 2928 18205 2992
rect 18269 2928 18270 2992
rect 18204 2838 18270 2928
rect 18330 2834 18390 3866
rect 18450 2774 18510 3804
rect 18570 2834 18630 3866
rect 18690 2774 18750 3804
rect 18810 3712 18876 3866
rect 18810 3648 18811 3712
rect 18875 3648 18876 3712
rect 18810 3632 18876 3648
rect 18810 3568 18811 3632
rect 18875 3568 18876 3632
rect 18810 3552 18876 3568
rect 18810 3488 18811 3552
rect 18875 3488 18876 3552
rect 18810 3472 18876 3488
rect 18810 3408 18811 3472
rect 18875 3408 18876 3472
rect 18810 3392 18876 3408
rect 18810 3328 18811 3392
rect 18875 3328 18876 3392
rect 18810 3312 18876 3328
rect 18810 3248 18811 3312
rect 18875 3248 18876 3312
rect 18810 3232 18876 3248
rect 18810 3168 18811 3232
rect 18875 3168 18876 3232
rect 18810 3152 18876 3168
rect 18810 3088 18811 3152
rect 18875 3088 18876 3152
rect 18810 3072 18876 3088
rect 18810 3008 18811 3072
rect 18875 3008 18876 3072
rect 18810 2992 18876 3008
rect 18810 2928 18811 2992
rect 18875 2928 18876 2992
rect 18810 2838 18876 2928
rect 18936 2834 18996 3866
rect 19056 2774 19116 3804
rect 19176 2834 19236 3866
rect 19296 2774 19356 3804
rect 19416 3712 19482 3866
rect 19416 3648 19417 3712
rect 19481 3648 19482 3712
rect 19416 3632 19482 3648
rect 19416 3568 19417 3632
rect 19481 3568 19482 3632
rect 19416 3552 19482 3568
rect 19416 3488 19417 3552
rect 19481 3488 19482 3552
rect 19416 3472 19482 3488
rect 19416 3408 19417 3472
rect 19481 3408 19482 3472
rect 19416 3392 19482 3408
rect 19416 3328 19417 3392
rect 19481 3328 19482 3392
rect 19416 3312 19482 3328
rect 19416 3248 19417 3312
rect 19481 3248 19482 3312
rect 19416 3232 19482 3248
rect 19416 3168 19417 3232
rect 19481 3168 19482 3232
rect 19416 3152 19482 3168
rect 19416 3088 19417 3152
rect 19481 3088 19482 3152
rect 19416 3072 19482 3088
rect 19416 3008 19417 3072
rect 19481 3008 19482 3072
rect 19416 2992 19482 3008
rect 19416 2928 19417 2992
rect 19481 2928 19482 2992
rect 19416 2838 19482 2928
rect 19542 2834 19602 3866
rect 19662 2774 19722 3804
rect 19782 2834 19842 3866
rect 19902 2774 19962 3804
rect 20022 3712 20088 3866
rect 20022 3648 20023 3712
rect 20087 3648 20088 3712
rect 20022 3632 20088 3648
rect 20022 3568 20023 3632
rect 20087 3568 20088 3632
rect 20022 3552 20088 3568
rect 20022 3488 20023 3552
rect 20087 3488 20088 3552
rect 20022 3472 20088 3488
rect 20022 3408 20023 3472
rect 20087 3408 20088 3472
rect 20022 3392 20088 3408
rect 20022 3328 20023 3392
rect 20087 3328 20088 3392
rect 20022 3312 20088 3328
rect 20022 3248 20023 3312
rect 20087 3248 20088 3312
rect 20022 3232 20088 3248
rect 20022 3168 20023 3232
rect 20087 3168 20088 3232
rect 20022 3152 20088 3168
rect 20022 3088 20023 3152
rect 20087 3088 20088 3152
rect 20022 3072 20088 3088
rect 20022 3008 20023 3072
rect 20087 3008 20088 3072
rect 20022 2992 20088 3008
rect 20022 2928 20023 2992
rect 20087 2928 20088 2992
rect 20022 2838 20088 2928
rect 20148 4872 20214 4962
rect 20148 4808 20149 4872
rect 20213 4808 20214 4872
rect 20148 4792 20214 4808
rect 20148 4728 20149 4792
rect 20213 4728 20214 4792
rect 20148 4712 20214 4728
rect 20148 4648 20149 4712
rect 20213 4648 20214 4712
rect 20148 4632 20214 4648
rect 20148 4568 20149 4632
rect 20213 4568 20214 4632
rect 20148 4552 20214 4568
rect 20148 4488 20149 4552
rect 20213 4488 20214 4552
rect 20148 4472 20214 4488
rect 20148 4408 20149 4472
rect 20213 4408 20214 4472
rect 20148 4392 20214 4408
rect 20148 4328 20149 4392
rect 20213 4328 20214 4392
rect 20148 4312 20214 4328
rect 20148 4248 20149 4312
rect 20213 4248 20214 4312
rect 20148 4232 20214 4248
rect 20148 4168 20149 4232
rect 20213 4168 20214 4232
rect 20148 4152 20214 4168
rect 20148 4088 20149 4152
rect 20213 4088 20214 4152
rect 20148 3934 20214 4088
rect 20274 3996 20334 5026
rect 20394 3934 20454 4966
rect 20514 3996 20574 5026
rect 20634 3934 20694 4966
rect 20754 4872 20820 4962
rect 20754 4808 20755 4872
rect 20819 4808 20820 4872
rect 20754 4792 20820 4808
rect 20754 4728 20755 4792
rect 20819 4728 20820 4792
rect 20754 4712 20820 4728
rect 20754 4648 20755 4712
rect 20819 4648 20820 4712
rect 20754 4632 20820 4648
rect 20754 4568 20755 4632
rect 20819 4568 20820 4632
rect 20754 4552 20820 4568
rect 20754 4488 20755 4552
rect 20819 4488 20820 4552
rect 20754 4472 20820 4488
rect 20754 4408 20755 4472
rect 20819 4408 20820 4472
rect 20754 4392 20820 4408
rect 20754 4328 20755 4392
rect 20819 4328 20820 4392
rect 20754 4312 20820 4328
rect 20754 4248 20755 4312
rect 20819 4248 20820 4312
rect 20754 4232 20820 4248
rect 20754 4168 20755 4232
rect 20819 4168 20820 4232
rect 20754 4152 20820 4168
rect 20754 4088 20755 4152
rect 20819 4088 20820 4152
rect 20754 3934 20820 4088
rect 20880 3996 20940 5026
rect 21000 3934 21060 4966
rect 21120 3996 21180 5026
rect 21240 3934 21300 4966
rect 21360 4872 21426 4962
rect 21360 4808 21361 4872
rect 21425 4808 21426 4872
rect 21360 4792 21426 4808
rect 21360 4728 21361 4792
rect 21425 4728 21426 4792
rect 21360 4712 21426 4728
rect 21360 4648 21361 4712
rect 21425 4648 21426 4712
rect 21360 4632 21426 4648
rect 21360 4568 21361 4632
rect 21425 4568 21426 4632
rect 21360 4552 21426 4568
rect 21360 4488 21361 4552
rect 21425 4488 21426 4552
rect 21360 4472 21426 4488
rect 21360 4408 21361 4472
rect 21425 4408 21426 4472
rect 21360 4392 21426 4408
rect 21360 4328 21361 4392
rect 21425 4328 21426 4392
rect 21360 4312 21426 4328
rect 21360 4248 21361 4312
rect 21425 4248 21426 4312
rect 21360 4232 21426 4248
rect 21360 4168 21361 4232
rect 21425 4168 21426 4232
rect 21360 4152 21426 4168
rect 21360 4088 21361 4152
rect 21425 4088 21426 4152
rect 21360 3934 21426 4088
rect 21486 3996 21546 5026
rect 21606 3934 21666 4966
rect 21726 3996 21786 5026
rect 21846 3934 21906 4966
rect 21966 4872 22032 4962
rect 21966 4808 21967 4872
rect 22031 4808 22032 4872
rect 21966 4792 22032 4808
rect 21966 4728 21967 4792
rect 22031 4728 22032 4792
rect 21966 4712 22032 4728
rect 21966 4648 21967 4712
rect 22031 4648 22032 4712
rect 21966 4632 22032 4648
rect 21966 4568 21967 4632
rect 22031 4568 22032 4632
rect 21966 4552 22032 4568
rect 21966 4488 21967 4552
rect 22031 4488 22032 4552
rect 21966 4472 22032 4488
rect 21966 4408 21967 4472
rect 22031 4408 22032 4472
rect 21966 4392 22032 4408
rect 21966 4328 21967 4392
rect 22031 4328 22032 4392
rect 21966 4312 22032 4328
rect 21966 4248 21967 4312
rect 22031 4248 22032 4312
rect 21966 4232 22032 4248
rect 21966 4168 21967 4232
rect 22031 4168 22032 4232
rect 21966 4152 22032 4168
rect 21966 4088 21967 4152
rect 22031 4088 22032 4152
rect 21966 3934 22032 4088
rect 22092 3996 22152 5026
rect 22212 3934 22272 4966
rect 22332 3996 22392 5026
rect 22452 3934 22512 4966
rect 22572 4872 22638 4962
rect 22572 4808 22573 4872
rect 22637 4808 22638 4872
rect 22572 4792 22638 4808
rect 22572 4728 22573 4792
rect 22637 4728 22638 4792
rect 22572 4712 22638 4728
rect 22572 4648 22573 4712
rect 22637 4648 22638 4712
rect 22572 4632 22638 4648
rect 22572 4568 22573 4632
rect 22637 4568 22638 4632
rect 22572 4552 22638 4568
rect 22572 4488 22573 4552
rect 22637 4488 22638 4552
rect 22572 4472 22638 4488
rect 22572 4408 22573 4472
rect 22637 4408 22638 4472
rect 22572 4392 22638 4408
rect 22572 4328 22573 4392
rect 22637 4328 22638 4392
rect 22572 4312 22638 4328
rect 22572 4248 22573 4312
rect 22637 4248 22638 4312
rect 22572 4232 22638 4248
rect 22572 4168 22573 4232
rect 22637 4168 22638 4232
rect 22572 4152 22638 4168
rect 22572 4088 22573 4152
rect 22637 4088 22638 4152
rect 22572 3934 22638 4088
rect 22698 3996 22758 5026
rect 22818 3934 22878 4966
rect 22938 3996 22998 5026
rect 23058 3934 23118 4966
rect 23178 4872 23244 4962
rect 23178 4808 23179 4872
rect 23243 4808 23244 4872
rect 23178 4792 23244 4808
rect 23178 4728 23179 4792
rect 23243 4728 23244 4792
rect 23178 4712 23244 4728
rect 23178 4648 23179 4712
rect 23243 4648 23244 4712
rect 23178 4632 23244 4648
rect 23178 4568 23179 4632
rect 23243 4568 23244 4632
rect 23178 4552 23244 4568
rect 23178 4488 23179 4552
rect 23243 4488 23244 4552
rect 23178 4472 23244 4488
rect 23178 4408 23179 4472
rect 23243 4408 23244 4472
rect 23178 4392 23244 4408
rect 23178 4328 23179 4392
rect 23243 4328 23244 4392
rect 23178 4312 23244 4328
rect 23178 4248 23179 4312
rect 23243 4248 23244 4312
rect 23178 4232 23244 4248
rect 23178 4168 23179 4232
rect 23243 4168 23244 4232
rect 23178 4152 23244 4168
rect 23178 4088 23179 4152
rect 23243 4088 23244 4152
rect 23178 3934 23244 4088
rect 23304 3996 23364 5026
rect 23424 3934 23484 4966
rect 23544 3996 23604 5026
rect 23664 3934 23724 4966
rect 23784 4872 23850 4962
rect 23784 4808 23785 4872
rect 23849 4808 23850 4872
rect 23784 4792 23850 4808
rect 23784 4728 23785 4792
rect 23849 4728 23850 4792
rect 23784 4712 23850 4728
rect 23784 4648 23785 4712
rect 23849 4648 23850 4712
rect 23784 4632 23850 4648
rect 23784 4568 23785 4632
rect 23849 4568 23850 4632
rect 23784 4552 23850 4568
rect 23784 4488 23785 4552
rect 23849 4488 23850 4552
rect 23784 4472 23850 4488
rect 23784 4408 23785 4472
rect 23849 4408 23850 4472
rect 23784 4392 23850 4408
rect 23784 4328 23785 4392
rect 23849 4328 23850 4392
rect 23784 4312 23850 4328
rect 23784 4248 23785 4312
rect 23849 4248 23850 4312
rect 23784 4232 23850 4248
rect 23784 4168 23785 4232
rect 23849 4168 23850 4232
rect 23784 4152 23850 4168
rect 23784 4088 23785 4152
rect 23849 4088 23850 4152
rect 23784 3934 23850 4088
rect 23910 3996 23970 5026
rect 24030 3934 24090 4966
rect 24150 3996 24210 5026
rect 24270 3934 24330 4966
rect 24390 4872 24456 4962
rect 24390 4808 24391 4872
rect 24455 4808 24456 4872
rect 24390 4792 24456 4808
rect 24390 4728 24391 4792
rect 24455 4728 24456 4792
rect 24390 4712 24456 4728
rect 24390 4648 24391 4712
rect 24455 4648 24456 4712
rect 24390 4632 24456 4648
rect 24390 4568 24391 4632
rect 24455 4568 24456 4632
rect 24390 4552 24456 4568
rect 24390 4488 24391 4552
rect 24455 4488 24456 4552
rect 24390 4472 24456 4488
rect 24390 4408 24391 4472
rect 24455 4408 24456 4472
rect 24390 4392 24456 4408
rect 24390 4328 24391 4392
rect 24455 4328 24456 4392
rect 24390 4312 24456 4328
rect 24390 4248 24391 4312
rect 24455 4248 24456 4312
rect 24390 4232 24456 4248
rect 24390 4168 24391 4232
rect 24455 4168 24456 4232
rect 24390 4152 24456 4168
rect 24390 4088 24391 4152
rect 24455 4088 24456 4152
rect 24390 3934 24456 4088
rect 24516 3996 24576 5026
rect 24636 3934 24696 4966
rect 24756 3996 24816 5026
rect 24876 3934 24936 4966
rect 24996 4872 25062 4962
rect 24996 4808 24997 4872
rect 25061 4808 25062 4872
rect 24996 4792 25062 4808
rect 24996 4728 24997 4792
rect 25061 4728 25062 4792
rect 24996 4712 25062 4728
rect 24996 4648 24997 4712
rect 25061 4648 25062 4712
rect 24996 4632 25062 4648
rect 24996 4568 24997 4632
rect 25061 4568 25062 4632
rect 24996 4552 25062 4568
rect 24996 4488 24997 4552
rect 25061 4488 25062 4552
rect 24996 4472 25062 4488
rect 24996 4408 24997 4472
rect 25061 4408 25062 4472
rect 24996 4392 25062 4408
rect 24996 4328 24997 4392
rect 25061 4328 25062 4392
rect 24996 4312 25062 4328
rect 24996 4248 24997 4312
rect 25061 4248 25062 4312
rect 24996 4232 25062 4248
rect 24996 4168 24997 4232
rect 25061 4168 25062 4232
rect 24996 4152 25062 4168
rect 24996 4088 24997 4152
rect 25061 4088 25062 4152
rect 24996 3934 25062 4088
rect 25122 3996 25182 5026
rect 25242 3934 25302 4966
rect 25362 3996 25422 5026
rect 25482 3934 25542 4966
rect 25602 4872 25668 4962
rect 25602 4808 25603 4872
rect 25667 4808 25668 4872
rect 25602 4792 25668 4808
rect 25602 4728 25603 4792
rect 25667 4728 25668 4792
rect 25602 4712 25668 4728
rect 25602 4648 25603 4712
rect 25667 4648 25668 4712
rect 25602 4632 25668 4648
rect 25602 4568 25603 4632
rect 25667 4568 25668 4632
rect 25602 4552 25668 4568
rect 25602 4488 25603 4552
rect 25667 4488 25668 4552
rect 25602 4472 25668 4488
rect 25602 4408 25603 4472
rect 25667 4408 25668 4472
rect 25602 4392 25668 4408
rect 25602 4328 25603 4392
rect 25667 4328 25668 4392
rect 25602 4312 25668 4328
rect 25602 4248 25603 4312
rect 25667 4248 25668 4312
rect 25602 4232 25668 4248
rect 25602 4168 25603 4232
rect 25667 4168 25668 4232
rect 25602 4152 25668 4168
rect 25602 4088 25603 4152
rect 25667 4088 25668 4152
rect 25602 3934 25668 4088
rect 25728 3996 25788 5026
rect 25848 3934 25908 4966
rect 25968 3996 26028 5026
rect 26088 3934 26148 4966
rect 26208 4872 26274 4962
rect 26208 4808 26209 4872
rect 26273 4808 26274 4872
rect 26208 4792 26274 4808
rect 26208 4728 26209 4792
rect 26273 4728 26274 4792
rect 26208 4712 26274 4728
rect 26208 4648 26209 4712
rect 26273 4648 26274 4712
rect 26208 4632 26274 4648
rect 26208 4568 26209 4632
rect 26273 4568 26274 4632
rect 26208 4552 26274 4568
rect 26208 4488 26209 4552
rect 26273 4488 26274 4552
rect 26208 4472 26274 4488
rect 26208 4408 26209 4472
rect 26273 4408 26274 4472
rect 26208 4392 26274 4408
rect 26208 4328 26209 4392
rect 26273 4328 26274 4392
rect 26208 4312 26274 4328
rect 26208 4248 26209 4312
rect 26273 4248 26274 4312
rect 26208 4232 26274 4248
rect 26208 4168 26209 4232
rect 26273 4168 26274 4232
rect 26208 4152 26274 4168
rect 26208 4088 26209 4152
rect 26273 4088 26274 4152
rect 26208 3934 26274 4088
rect 26334 3996 26394 5026
rect 26454 3934 26514 4966
rect 26574 3996 26634 5026
rect 26694 3934 26754 4966
rect 26814 4872 26880 4962
rect 26814 4808 26815 4872
rect 26879 4808 26880 4872
rect 26814 4792 26880 4808
rect 26814 4728 26815 4792
rect 26879 4728 26880 4792
rect 26814 4712 26880 4728
rect 26814 4648 26815 4712
rect 26879 4648 26880 4712
rect 26814 4632 26880 4648
rect 26814 4568 26815 4632
rect 26879 4568 26880 4632
rect 26814 4552 26880 4568
rect 26814 4488 26815 4552
rect 26879 4488 26880 4552
rect 26814 4472 26880 4488
rect 26814 4408 26815 4472
rect 26879 4408 26880 4472
rect 26814 4392 26880 4408
rect 26814 4328 26815 4392
rect 26879 4328 26880 4392
rect 26814 4312 26880 4328
rect 26814 4248 26815 4312
rect 26879 4248 26880 4312
rect 26814 4232 26880 4248
rect 26814 4168 26815 4232
rect 26879 4168 26880 4232
rect 26814 4152 26880 4168
rect 26814 4088 26815 4152
rect 26879 4088 26880 4152
rect 26814 3934 26880 4088
rect 26940 3996 27000 5026
rect 27060 3934 27120 4966
rect 27180 3996 27240 5026
rect 27300 3934 27360 4966
rect 27420 4872 27486 4962
rect 27420 4808 27421 4872
rect 27485 4808 27486 4872
rect 27420 4792 27486 4808
rect 27420 4728 27421 4792
rect 27485 4728 27486 4792
rect 27420 4712 27486 4728
rect 27420 4648 27421 4712
rect 27485 4648 27486 4712
rect 27420 4632 27486 4648
rect 27420 4568 27421 4632
rect 27485 4568 27486 4632
rect 27420 4552 27486 4568
rect 27420 4488 27421 4552
rect 27485 4488 27486 4552
rect 27420 4472 27486 4488
rect 27420 4408 27421 4472
rect 27485 4408 27486 4472
rect 27420 4392 27486 4408
rect 27420 4328 27421 4392
rect 27485 4328 27486 4392
rect 27420 4312 27486 4328
rect 27420 4248 27421 4312
rect 27485 4248 27486 4312
rect 27420 4232 27486 4248
rect 27420 4168 27421 4232
rect 27485 4168 27486 4232
rect 27420 4152 27486 4168
rect 27420 4088 27421 4152
rect 27485 4088 27486 4152
rect 27420 3934 27486 4088
rect 27546 3996 27606 5026
rect 27666 3934 27726 4966
rect 27786 3996 27846 5026
rect 27906 3934 27966 4966
rect 28026 4872 28092 4962
rect 28026 4808 28027 4872
rect 28091 4808 28092 4872
rect 28026 4792 28092 4808
rect 28026 4728 28027 4792
rect 28091 4728 28092 4792
rect 28026 4712 28092 4728
rect 28026 4648 28027 4712
rect 28091 4648 28092 4712
rect 28026 4632 28092 4648
rect 28026 4568 28027 4632
rect 28091 4568 28092 4632
rect 28026 4552 28092 4568
rect 28026 4488 28027 4552
rect 28091 4488 28092 4552
rect 28026 4472 28092 4488
rect 28026 4408 28027 4472
rect 28091 4408 28092 4472
rect 28026 4392 28092 4408
rect 28026 4328 28027 4392
rect 28091 4328 28092 4392
rect 28026 4312 28092 4328
rect 28026 4248 28027 4312
rect 28091 4248 28092 4312
rect 28026 4232 28092 4248
rect 28026 4168 28027 4232
rect 28091 4168 28092 4232
rect 28026 4152 28092 4168
rect 28026 4088 28027 4152
rect 28091 4088 28092 4152
rect 28026 3934 28092 4088
rect 28152 3996 28212 5026
rect 28272 3934 28332 4966
rect 28392 3996 28452 5026
rect 28512 3934 28572 4966
rect 28632 4872 28698 4962
rect 28632 4808 28633 4872
rect 28697 4808 28698 4872
rect 28632 4792 28698 4808
rect 28632 4728 28633 4792
rect 28697 4728 28698 4792
rect 28632 4712 28698 4728
rect 28632 4648 28633 4712
rect 28697 4648 28698 4712
rect 28632 4632 28698 4648
rect 28632 4568 28633 4632
rect 28697 4568 28698 4632
rect 28632 4552 28698 4568
rect 28632 4488 28633 4552
rect 28697 4488 28698 4552
rect 28632 4472 28698 4488
rect 28632 4408 28633 4472
rect 28697 4408 28698 4472
rect 28632 4392 28698 4408
rect 28632 4328 28633 4392
rect 28697 4328 28698 4392
rect 28632 4312 28698 4328
rect 28632 4248 28633 4312
rect 28697 4248 28698 4312
rect 28632 4232 28698 4248
rect 28632 4168 28633 4232
rect 28697 4168 28698 4232
rect 28632 4152 28698 4168
rect 28632 4088 28633 4152
rect 28697 4088 28698 4152
rect 28632 3934 28698 4088
rect 28758 3996 28818 5026
rect 28878 3934 28938 4966
rect 28998 3996 29058 5026
rect 29118 3934 29178 4966
rect 29238 4872 29304 4962
rect 29238 4808 29239 4872
rect 29303 4808 29304 4872
rect 29238 4792 29304 4808
rect 29238 4728 29239 4792
rect 29303 4728 29304 4792
rect 29238 4712 29304 4728
rect 29238 4648 29239 4712
rect 29303 4648 29304 4712
rect 29238 4632 29304 4648
rect 29238 4568 29239 4632
rect 29303 4568 29304 4632
rect 29238 4552 29304 4568
rect 29238 4488 29239 4552
rect 29303 4488 29304 4552
rect 29238 4472 29304 4488
rect 29238 4408 29239 4472
rect 29303 4408 29304 4472
rect 29238 4392 29304 4408
rect 29238 4328 29239 4392
rect 29303 4328 29304 4392
rect 29238 4312 29304 4328
rect 29238 4248 29239 4312
rect 29303 4248 29304 4312
rect 29238 4232 29304 4248
rect 29238 4168 29239 4232
rect 29303 4168 29304 4232
rect 29238 4152 29304 4168
rect 29238 4088 29239 4152
rect 29303 4088 29304 4152
rect 29238 3934 29304 4088
rect 29364 3996 29424 5026
rect 29484 3934 29544 4966
rect 29604 3996 29664 5026
rect 29724 3934 29784 4966
rect 29844 4872 29910 4962
rect 29844 4808 29845 4872
rect 29909 4808 29910 4872
rect 29844 4792 29910 4808
rect 29844 4728 29845 4792
rect 29909 4728 29910 4792
rect 29844 4712 29910 4728
rect 29844 4648 29845 4712
rect 29909 4648 29910 4712
rect 29844 4632 29910 4648
rect 29844 4568 29845 4632
rect 29909 4568 29910 4632
rect 29844 4552 29910 4568
rect 29844 4488 29845 4552
rect 29909 4488 29910 4552
rect 29844 4472 29910 4488
rect 29844 4408 29845 4472
rect 29909 4408 29910 4472
rect 29844 4392 29910 4408
rect 29844 4328 29845 4392
rect 29909 4328 29910 4392
rect 29844 4312 29910 4328
rect 29844 4248 29845 4312
rect 29909 4248 29910 4312
rect 29844 4232 29910 4248
rect 29844 4168 29845 4232
rect 29909 4168 29910 4232
rect 29844 4152 29910 4168
rect 29844 4088 29845 4152
rect 29909 4088 29910 4152
rect 29844 3934 29910 4088
rect 29970 3996 30030 5026
rect 30090 3934 30150 4966
rect 30210 3996 30270 5026
rect 30330 3934 30390 4966
rect 30450 4872 30516 4962
rect 30450 4808 30451 4872
rect 30515 4808 30516 4872
rect 30450 4792 30516 4808
rect 30450 4728 30451 4792
rect 30515 4728 30516 4792
rect 30450 4712 30516 4728
rect 30450 4648 30451 4712
rect 30515 4648 30516 4712
rect 30450 4632 30516 4648
rect 30450 4568 30451 4632
rect 30515 4568 30516 4632
rect 30450 4552 30516 4568
rect 30450 4488 30451 4552
rect 30515 4488 30516 4552
rect 30450 4472 30516 4488
rect 30450 4408 30451 4472
rect 30515 4408 30516 4472
rect 30450 4392 30516 4408
rect 30450 4328 30451 4392
rect 30515 4328 30516 4392
rect 30450 4312 30516 4328
rect 30450 4248 30451 4312
rect 30515 4248 30516 4312
rect 30450 4232 30516 4248
rect 30450 4168 30451 4232
rect 30515 4168 30516 4232
rect 30450 4152 30516 4168
rect 30450 4088 30451 4152
rect 30515 4088 30516 4152
rect 30450 3934 30516 4088
rect 30576 3996 30636 5026
rect 30696 3934 30756 4966
rect 30816 3996 30876 5026
rect 30936 3934 30996 4966
rect 31056 4872 31122 4962
rect 31056 4808 31057 4872
rect 31121 4808 31122 4872
rect 31056 4792 31122 4808
rect 31056 4728 31057 4792
rect 31121 4728 31122 4792
rect 31056 4712 31122 4728
rect 31056 4648 31057 4712
rect 31121 4648 31122 4712
rect 31056 4632 31122 4648
rect 31056 4568 31057 4632
rect 31121 4568 31122 4632
rect 31056 4552 31122 4568
rect 31056 4488 31057 4552
rect 31121 4488 31122 4552
rect 31056 4472 31122 4488
rect 31056 4408 31057 4472
rect 31121 4408 31122 4472
rect 31056 4392 31122 4408
rect 31056 4328 31057 4392
rect 31121 4328 31122 4392
rect 31056 4312 31122 4328
rect 31056 4248 31057 4312
rect 31121 4248 31122 4312
rect 31056 4232 31122 4248
rect 31056 4168 31057 4232
rect 31121 4168 31122 4232
rect 31056 4152 31122 4168
rect 31056 4088 31057 4152
rect 31121 4088 31122 4152
rect 31056 3934 31122 4088
rect 31182 3996 31242 5026
rect 31302 3934 31362 4966
rect 31422 3996 31482 5026
rect 31542 3934 31602 4966
rect 31662 4872 31728 4962
rect 31662 4808 31663 4872
rect 31727 4808 31728 4872
rect 31662 4792 31728 4808
rect 31662 4728 31663 4792
rect 31727 4728 31728 4792
rect 31662 4712 31728 4728
rect 31662 4648 31663 4712
rect 31727 4648 31728 4712
rect 31662 4632 31728 4648
rect 31662 4568 31663 4632
rect 31727 4568 31728 4632
rect 31662 4552 31728 4568
rect 31662 4488 31663 4552
rect 31727 4488 31728 4552
rect 31662 4472 31728 4488
rect 31662 4408 31663 4472
rect 31727 4408 31728 4472
rect 31662 4392 31728 4408
rect 31662 4328 31663 4392
rect 31727 4328 31728 4392
rect 31662 4312 31728 4328
rect 31662 4248 31663 4312
rect 31727 4248 31728 4312
rect 31662 4232 31728 4248
rect 31662 4168 31663 4232
rect 31727 4168 31728 4232
rect 31662 4152 31728 4168
rect 31662 4088 31663 4152
rect 31727 4088 31728 4152
rect 31662 3934 31728 4088
rect 31788 3996 31848 5026
rect 31908 3934 31968 4966
rect 32028 3996 32088 5026
rect 32148 3934 32208 4966
rect 32268 4872 32334 4962
rect 32268 4808 32269 4872
rect 32333 4808 32334 4872
rect 32268 4792 32334 4808
rect 32268 4728 32269 4792
rect 32333 4728 32334 4792
rect 32268 4712 32334 4728
rect 32268 4648 32269 4712
rect 32333 4648 32334 4712
rect 32268 4632 32334 4648
rect 32268 4568 32269 4632
rect 32333 4568 32334 4632
rect 32268 4552 32334 4568
rect 32268 4488 32269 4552
rect 32333 4488 32334 4552
rect 32268 4472 32334 4488
rect 32268 4408 32269 4472
rect 32333 4408 32334 4472
rect 32268 4392 32334 4408
rect 32268 4328 32269 4392
rect 32333 4328 32334 4392
rect 32268 4312 32334 4328
rect 32268 4248 32269 4312
rect 32333 4248 32334 4312
rect 32268 4232 32334 4248
rect 32268 4168 32269 4232
rect 32333 4168 32334 4232
rect 32268 4152 32334 4168
rect 32268 4088 32269 4152
rect 32333 4088 32334 4152
rect 32268 3934 32334 4088
rect 32394 3996 32454 5026
rect 32514 3934 32574 4966
rect 32634 3996 32694 5026
rect 32754 3934 32814 4966
rect 32874 4872 32940 4962
rect 32874 4808 32875 4872
rect 32939 4808 32940 4872
rect 32874 4792 32940 4808
rect 32874 4728 32875 4792
rect 32939 4728 32940 4792
rect 32874 4712 32940 4728
rect 32874 4648 32875 4712
rect 32939 4648 32940 4712
rect 32874 4632 32940 4648
rect 32874 4568 32875 4632
rect 32939 4568 32940 4632
rect 32874 4552 32940 4568
rect 32874 4488 32875 4552
rect 32939 4488 32940 4552
rect 32874 4472 32940 4488
rect 32874 4408 32875 4472
rect 32939 4408 32940 4472
rect 32874 4392 32940 4408
rect 32874 4328 32875 4392
rect 32939 4328 32940 4392
rect 32874 4312 32940 4328
rect 32874 4248 32875 4312
rect 32939 4248 32940 4312
rect 32874 4232 32940 4248
rect 32874 4168 32875 4232
rect 32939 4168 32940 4232
rect 32874 4152 32940 4168
rect 32874 4088 32875 4152
rect 32939 4088 32940 4152
rect 32874 3934 32940 4088
rect 33000 3996 33060 5026
rect 33120 3934 33180 4966
rect 33240 3996 33300 5026
rect 33360 3934 33420 4966
rect 33480 4872 33546 4962
rect 33480 4808 33481 4872
rect 33545 4808 33546 4872
rect 33480 4792 33546 4808
rect 33480 4728 33481 4792
rect 33545 4728 33546 4792
rect 33480 4712 33546 4728
rect 33480 4648 33481 4712
rect 33545 4648 33546 4712
rect 33480 4632 33546 4648
rect 33480 4568 33481 4632
rect 33545 4568 33546 4632
rect 33480 4552 33546 4568
rect 33480 4488 33481 4552
rect 33545 4488 33546 4552
rect 33480 4472 33546 4488
rect 33480 4408 33481 4472
rect 33545 4408 33546 4472
rect 33480 4392 33546 4408
rect 33480 4328 33481 4392
rect 33545 4328 33546 4392
rect 33480 4312 33546 4328
rect 33480 4248 33481 4312
rect 33545 4248 33546 4312
rect 33480 4232 33546 4248
rect 33480 4168 33481 4232
rect 33545 4168 33546 4232
rect 33480 4152 33546 4168
rect 33480 4088 33481 4152
rect 33545 4088 33546 4152
rect 33480 3934 33546 4088
rect 33606 3996 33666 5026
rect 33726 3934 33786 4966
rect 33846 3996 33906 5026
rect 33966 3934 34026 4966
rect 34086 4872 34152 4962
rect 34086 4808 34087 4872
rect 34151 4808 34152 4872
rect 34086 4792 34152 4808
rect 34086 4728 34087 4792
rect 34151 4728 34152 4792
rect 34086 4712 34152 4728
rect 34086 4648 34087 4712
rect 34151 4648 34152 4712
rect 34086 4632 34152 4648
rect 34086 4568 34087 4632
rect 34151 4568 34152 4632
rect 34086 4552 34152 4568
rect 34086 4488 34087 4552
rect 34151 4488 34152 4552
rect 34086 4472 34152 4488
rect 34086 4408 34087 4472
rect 34151 4408 34152 4472
rect 34086 4392 34152 4408
rect 34086 4328 34087 4392
rect 34151 4328 34152 4392
rect 34086 4312 34152 4328
rect 34086 4248 34087 4312
rect 34151 4248 34152 4312
rect 34086 4232 34152 4248
rect 34086 4168 34087 4232
rect 34151 4168 34152 4232
rect 34086 4152 34152 4168
rect 34086 4088 34087 4152
rect 34151 4088 34152 4152
rect 34086 3934 34152 4088
rect 34212 3996 34272 5026
rect 34332 3934 34392 4966
rect 34452 3996 34512 5026
rect 34572 3934 34632 4966
rect 34692 4872 34758 4962
rect 34692 4808 34693 4872
rect 34757 4808 34758 4872
rect 34692 4792 34758 4808
rect 34692 4728 34693 4792
rect 34757 4728 34758 4792
rect 34692 4712 34758 4728
rect 34692 4648 34693 4712
rect 34757 4648 34758 4712
rect 34692 4632 34758 4648
rect 34692 4568 34693 4632
rect 34757 4568 34758 4632
rect 34692 4552 34758 4568
rect 34692 4488 34693 4552
rect 34757 4488 34758 4552
rect 34692 4472 34758 4488
rect 34692 4408 34693 4472
rect 34757 4408 34758 4472
rect 34692 4392 34758 4408
rect 34692 4328 34693 4392
rect 34757 4328 34758 4392
rect 34692 4312 34758 4328
rect 34692 4248 34693 4312
rect 34757 4248 34758 4312
rect 34692 4232 34758 4248
rect 34692 4168 34693 4232
rect 34757 4168 34758 4232
rect 34692 4152 34758 4168
rect 34692 4088 34693 4152
rect 34757 4088 34758 4152
rect 34692 3934 34758 4088
rect 34818 3996 34878 5026
rect 34938 3934 34998 4966
rect 35058 3996 35118 5026
rect 35178 3934 35238 4966
rect 35298 4872 35364 4962
rect 35298 4808 35299 4872
rect 35363 4808 35364 4872
rect 35298 4792 35364 4808
rect 35298 4728 35299 4792
rect 35363 4728 35364 4792
rect 35298 4712 35364 4728
rect 35298 4648 35299 4712
rect 35363 4648 35364 4712
rect 35298 4632 35364 4648
rect 35298 4568 35299 4632
rect 35363 4568 35364 4632
rect 35298 4552 35364 4568
rect 35298 4488 35299 4552
rect 35363 4488 35364 4552
rect 35298 4472 35364 4488
rect 35298 4408 35299 4472
rect 35363 4408 35364 4472
rect 35298 4392 35364 4408
rect 35298 4328 35299 4392
rect 35363 4328 35364 4392
rect 35298 4312 35364 4328
rect 35298 4248 35299 4312
rect 35363 4248 35364 4312
rect 35298 4232 35364 4248
rect 35298 4168 35299 4232
rect 35363 4168 35364 4232
rect 35298 4152 35364 4168
rect 35298 4088 35299 4152
rect 35363 4088 35364 4152
rect 35298 3934 35364 4088
rect 35424 3996 35484 5026
rect 35544 3934 35604 4966
rect 35664 3996 35724 5026
rect 35784 3934 35844 4966
rect 35904 4872 35970 4962
rect 35904 4808 35905 4872
rect 35969 4808 35970 4872
rect 35904 4792 35970 4808
rect 35904 4728 35905 4792
rect 35969 4728 35970 4792
rect 35904 4712 35970 4728
rect 35904 4648 35905 4712
rect 35969 4648 35970 4712
rect 35904 4632 35970 4648
rect 35904 4568 35905 4632
rect 35969 4568 35970 4632
rect 35904 4552 35970 4568
rect 35904 4488 35905 4552
rect 35969 4488 35970 4552
rect 35904 4472 35970 4488
rect 35904 4408 35905 4472
rect 35969 4408 35970 4472
rect 35904 4392 35970 4408
rect 35904 4328 35905 4392
rect 35969 4328 35970 4392
rect 35904 4312 35970 4328
rect 35904 4248 35905 4312
rect 35969 4248 35970 4312
rect 35904 4232 35970 4248
rect 35904 4168 35905 4232
rect 35969 4168 35970 4232
rect 35904 4152 35970 4168
rect 35904 4088 35905 4152
rect 35969 4088 35970 4152
rect 35904 3934 35970 4088
rect 36030 3996 36090 5026
rect 36150 3934 36210 4966
rect 36270 3996 36330 5026
rect 36390 3934 36450 4966
rect 36510 4872 36576 4962
rect 36510 4808 36511 4872
rect 36575 4808 36576 4872
rect 36510 4792 36576 4808
rect 36510 4728 36511 4792
rect 36575 4728 36576 4792
rect 36510 4712 36576 4728
rect 36510 4648 36511 4712
rect 36575 4648 36576 4712
rect 36510 4632 36576 4648
rect 36510 4568 36511 4632
rect 36575 4568 36576 4632
rect 36510 4552 36576 4568
rect 36510 4488 36511 4552
rect 36575 4488 36576 4552
rect 36510 4472 36576 4488
rect 36510 4408 36511 4472
rect 36575 4408 36576 4472
rect 36510 4392 36576 4408
rect 36510 4328 36511 4392
rect 36575 4328 36576 4392
rect 36510 4312 36576 4328
rect 36510 4248 36511 4312
rect 36575 4248 36576 4312
rect 36510 4232 36576 4248
rect 36510 4168 36511 4232
rect 36575 4168 36576 4232
rect 36510 4152 36576 4168
rect 36510 4088 36511 4152
rect 36575 4088 36576 4152
rect 36510 3934 36576 4088
rect 36636 3996 36696 5026
rect 36756 3934 36816 4966
rect 36876 3996 36936 5026
rect 36996 3934 37056 4966
rect 37116 4872 37182 4962
rect 37116 4808 37117 4872
rect 37181 4808 37182 4872
rect 37116 4792 37182 4808
rect 37116 4728 37117 4792
rect 37181 4728 37182 4792
rect 37116 4712 37182 4728
rect 37116 4648 37117 4712
rect 37181 4648 37182 4712
rect 37116 4632 37182 4648
rect 37116 4568 37117 4632
rect 37181 4568 37182 4632
rect 37116 4552 37182 4568
rect 37116 4488 37117 4552
rect 37181 4488 37182 4552
rect 37116 4472 37182 4488
rect 37116 4408 37117 4472
rect 37181 4408 37182 4472
rect 37116 4392 37182 4408
rect 37116 4328 37117 4392
rect 37181 4328 37182 4392
rect 37116 4312 37182 4328
rect 37116 4248 37117 4312
rect 37181 4248 37182 4312
rect 37116 4232 37182 4248
rect 37116 4168 37117 4232
rect 37181 4168 37182 4232
rect 37116 4152 37182 4168
rect 37116 4088 37117 4152
rect 37181 4088 37182 4152
rect 37116 3934 37182 4088
rect 37242 3996 37302 5026
rect 37362 3934 37422 4966
rect 37482 3996 37542 5026
rect 37602 3934 37662 4966
rect 37722 4872 37788 4962
rect 37722 4808 37723 4872
rect 37787 4808 37788 4872
rect 37722 4792 37788 4808
rect 37722 4728 37723 4792
rect 37787 4728 37788 4792
rect 37722 4712 37788 4728
rect 37722 4648 37723 4712
rect 37787 4648 37788 4712
rect 37722 4632 37788 4648
rect 37722 4568 37723 4632
rect 37787 4568 37788 4632
rect 37722 4552 37788 4568
rect 37722 4488 37723 4552
rect 37787 4488 37788 4552
rect 37722 4472 37788 4488
rect 37722 4408 37723 4472
rect 37787 4408 37788 4472
rect 37722 4392 37788 4408
rect 37722 4328 37723 4392
rect 37787 4328 37788 4392
rect 37722 4312 37788 4328
rect 37722 4248 37723 4312
rect 37787 4248 37788 4312
rect 37722 4232 37788 4248
rect 37722 4168 37723 4232
rect 37787 4168 37788 4232
rect 37722 4152 37788 4168
rect 37722 4088 37723 4152
rect 37787 4088 37788 4152
rect 37722 3934 37788 4088
rect 37848 3996 37908 5026
rect 37968 3934 38028 4966
rect 38088 3996 38148 5026
rect 38208 3934 38268 4966
rect 38328 4872 38394 4962
rect 38328 4808 38329 4872
rect 38393 4808 38394 4872
rect 38328 4792 38394 4808
rect 38328 4728 38329 4792
rect 38393 4728 38394 4792
rect 38328 4712 38394 4728
rect 38328 4648 38329 4712
rect 38393 4648 38394 4712
rect 38328 4632 38394 4648
rect 38328 4568 38329 4632
rect 38393 4568 38394 4632
rect 38328 4552 38394 4568
rect 38328 4488 38329 4552
rect 38393 4488 38394 4552
rect 38328 4472 38394 4488
rect 38328 4408 38329 4472
rect 38393 4408 38394 4472
rect 38328 4392 38394 4408
rect 38328 4328 38329 4392
rect 38393 4328 38394 4392
rect 38328 4312 38394 4328
rect 38328 4248 38329 4312
rect 38393 4248 38394 4312
rect 38328 4232 38394 4248
rect 38328 4168 38329 4232
rect 38393 4168 38394 4232
rect 38328 4152 38394 4168
rect 38328 4088 38329 4152
rect 38393 4088 38394 4152
rect 38328 3934 38394 4088
rect 38454 3996 38514 5026
rect 38574 3934 38634 4966
rect 38694 3996 38754 5026
rect 38814 3934 38874 4966
rect 38934 4872 39000 4962
rect 38934 4808 38935 4872
rect 38999 4808 39000 4872
rect 38934 4792 39000 4808
rect 38934 4728 38935 4792
rect 38999 4728 39000 4792
rect 38934 4712 39000 4728
rect 38934 4648 38935 4712
rect 38999 4648 39000 4712
rect 38934 4632 39000 4648
rect 38934 4568 38935 4632
rect 38999 4568 39000 4632
rect 38934 4552 39000 4568
rect 38934 4488 38935 4552
rect 38999 4488 39000 4552
rect 38934 4472 39000 4488
rect 38934 4408 38935 4472
rect 38999 4408 39000 4472
rect 38934 4392 39000 4408
rect 38934 4328 38935 4392
rect 38999 4328 39000 4392
rect 38934 4312 39000 4328
rect 38934 4248 38935 4312
rect 38999 4248 39000 4312
rect 38934 4232 39000 4248
rect 38934 4168 38935 4232
rect 38999 4168 39000 4232
rect 38934 4152 39000 4168
rect 38934 4088 38935 4152
rect 38999 4088 39000 4152
rect 38934 3934 39000 4088
rect 39060 3996 39120 5026
rect 39180 3934 39240 4966
rect 39300 3996 39360 5026
rect 39420 3934 39480 4966
rect 39540 4872 39606 4962
rect 39540 4808 39541 4872
rect 39605 4808 39606 4872
rect 39540 4792 39606 4808
rect 39540 4728 39541 4792
rect 39605 4728 39606 4792
rect 39540 4712 39606 4728
rect 39540 4648 39541 4712
rect 39605 4648 39606 4712
rect 39540 4632 39606 4648
rect 39540 4568 39541 4632
rect 39605 4568 39606 4632
rect 39540 4552 39606 4568
rect 39540 4488 39541 4552
rect 39605 4488 39606 4552
rect 39540 4472 39606 4488
rect 39540 4408 39541 4472
rect 39605 4408 39606 4472
rect 39540 4392 39606 4408
rect 39540 4328 39541 4392
rect 39605 4328 39606 4392
rect 39540 4312 39606 4328
rect 39540 4248 39541 4312
rect 39605 4248 39606 4312
rect 39540 4232 39606 4248
rect 39540 4168 39541 4232
rect 39605 4168 39606 4232
rect 39540 4152 39606 4168
rect 39540 4088 39541 4152
rect 39605 4088 39606 4152
rect 39540 3934 39606 4088
rect 20148 3932 39606 3934
rect 20148 3868 20252 3932
rect 20316 3868 20332 3932
rect 20396 3868 20412 3932
rect 20476 3868 20492 3932
rect 20556 3868 20572 3932
rect 20636 3868 20652 3932
rect 20716 3868 20858 3932
rect 20922 3868 20938 3932
rect 21002 3868 21018 3932
rect 21082 3868 21098 3932
rect 21162 3868 21178 3932
rect 21242 3868 21258 3932
rect 21322 3868 21464 3932
rect 21528 3868 21544 3932
rect 21608 3868 21624 3932
rect 21688 3868 21704 3932
rect 21768 3868 21784 3932
rect 21848 3868 21864 3932
rect 21928 3868 22070 3932
rect 22134 3868 22150 3932
rect 22214 3868 22230 3932
rect 22294 3868 22310 3932
rect 22374 3868 22390 3932
rect 22454 3868 22470 3932
rect 22534 3868 22676 3932
rect 22740 3868 22756 3932
rect 22820 3868 22836 3932
rect 22900 3868 22916 3932
rect 22980 3868 22996 3932
rect 23060 3868 23076 3932
rect 23140 3868 23282 3932
rect 23346 3868 23362 3932
rect 23426 3868 23442 3932
rect 23506 3868 23522 3932
rect 23586 3868 23602 3932
rect 23666 3868 23682 3932
rect 23746 3868 23888 3932
rect 23952 3868 23968 3932
rect 24032 3868 24048 3932
rect 24112 3868 24128 3932
rect 24192 3868 24208 3932
rect 24272 3868 24288 3932
rect 24352 3868 24494 3932
rect 24558 3868 24574 3932
rect 24638 3868 24654 3932
rect 24718 3868 24734 3932
rect 24798 3868 24814 3932
rect 24878 3868 24894 3932
rect 24958 3868 25100 3932
rect 25164 3868 25180 3932
rect 25244 3868 25260 3932
rect 25324 3868 25340 3932
rect 25404 3868 25420 3932
rect 25484 3868 25500 3932
rect 25564 3868 25706 3932
rect 25770 3868 25786 3932
rect 25850 3868 25866 3932
rect 25930 3868 25946 3932
rect 26010 3868 26026 3932
rect 26090 3868 26106 3932
rect 26170 3868 26312 3932
rect 26376 3868 26392 3932
rect 26456 3868 26472 3932
rect 26536 3868 26552 3932
rect 26616 3868 26632 3932
rect 26696 3868 26712 3932
rect 26776 3868 26918 3932
rect 26982 3868 26998 3932
rect 27062 3868 27078 3932
rect 27142 3868 27158 3932
rect 27222 3868 27238 3932
rect 27302 3868 27318 3932
rect 27382 3868 27524 3932
rect 27588 3868 27604 3932
rect 27668 3868 27684 3932
rect 27748 3868 27764 3932
rect 27828 3868 27844 3932
rect 27908 3868 27924 3932
rect 27988 3868 28130 3932
rect 28194 3868 28210 3932
rect 28274 3868 28290 3932
rect 28354 3868 28370 3932
rect 28434 3868 28450 3932
rect 28514 3868 28530 3932
rect 28594 3868 28736 3932
rect 28800 3868 28816 3932
rect 28880 3868 28896 3932
rect 28960 3868 28976 3932
rect 29040 3868 29056 3932
rect 29120 3868 29136 3932
rect 29200 3868 29342 3932
rect 29406 3868 29422 3932
rect 29486 3868 29502 3932
rect 29566 3868 29582 3932
rect 29646 3868 29662 3932
rect 29726 3868 29742 3932
rect 29806 3868 29948 3932
rect 30012 3868 30028 3932
rect 30092 3868 30108 3932
rect 30172 3868 30188 3932
rect 30252 3868 30268 3932
rect 30332 3868 30348 3932
rect 30412 3868 30554 3932
rect 30618 3868 30634 3932
rect 30698 3868 30714 3932
rect 30778 3868 30794 3932
rect 30858 3868 30874 3932
rect 30938 3868 30954 3932
rect 31018 3868 31160 3932
rect 31224 3868 31240 3932
rect 31304 3868 31320 3932
rect 31384 3868 31400 3932
rect 31464 3868 31480 3932
rect 31544 3868 31560 3932
rect 31624 3868 31766 3932
rect 31830 3868 31846 3932
rect 31910 3868 31926 3932
rect 31990 3868 32006 3932
rect 32070 3868 32086 3932
rect 32150 3868 32166 3932
rect 32230 3868 32372 3932
rect 32436 3868 32452 3932
rect 32516 3868 32532 3932
rect 32596 3868 32612 3932
rect 32676 3868 32692 3932
rect 32756 3868 32772 3932
rect 32836 3868 32978 3932
rect 33042 3868 33058 3932
rect 33122 3868 33138 3932
rect 33202 3868 33218 3932
rect 33282 3868 33298 3932
rect 33362 3868 33378 3932
rect 33442 3868 33584 3932
rect 33648 3868 33664 3932
rect 33728 3868 33744 3932
rect 33808 3868 33824 3932
rect 33888 3868 33904 3932
rect 33968 3868 33984 3932
rect 34048 3868 34190 3932
rect 34254 3868 34270 3932
rect 34334 3868 34350 3932
rect 34414 3868 34430 3932
rect 34494 3868 34510 3932
rect 34574 3868 34590 3932
rect 34654 3868 34796 3932
rect 34860 3868 34876 3932
rect 34940 3868 34956 3932
rect 35020 3868 35036 3932
rect 35100 3868 35116 3932
rect 35180 3868 35196 3932
rect 35260 3868 35402 3932
rect 35466 3868 35482 3932
rect 35546 3868 35562 3932
rect 35626 3868 35642 3932
rect 35706 3868 35722 3932
rect 35786 3868 35802 3932
rect 35866 3868 36008 3932
rect 36072 3868 36088 3932
rect 36152 3868 36168 3932
rect 36232 3868 36248 3932
rect 36312 3868 36328 3932
rect 36392 3868 36408 3932
rect 36472 3868 36614 3932
rect 36678 3868 36694 3932
rect 36758 3868 36774 3932
rect 36838 3868 36854 3932
rect 36918 3868 36934 3932
rect 36998 3868 37014 3932
rect 37078 3868 37220 3932
rect 37284 3868 37300 3932
rect 37364 3868 37380 3932
rect 37444 3868 37460 3932
rect 37524 3868 37540 3932
rect 37604 3868 37620 3932
rect 37684 3868 37826 3932
rect 37890 3868 37906 3932
rect 37970 3868 37986 3932
rect 38050 3868 38066 3932
rect 38130 3868 38146 3932
rect 38210 3868 38226 3932
rect 38290 3868 38432 3932
rect 38496 3868 38512 3932
rect 38576 3868 38592 3932
rect 38656 3868 38672 3932
rect 38736 3868 38752 3932
rect 38816 3868 38832 3932
rect 38896 3868 39038 3932
rect 39102 3868 39118 3932
rect 39182 3868 39198 3932
rect 39262 3868 39278 3932
rect 39342 3868 39358 3932
rect 39422 3868 39438 3932
rect 39502 3868 39606 3932
rect 20148 3866 39606 3868
rect 20148 3712 20214 3866
rect 20148 3648 20149 3712
rect 20213 3648 20214 3712
rect 20148 3632 20214 3648
rect 20148 3568 20149 3632
rect 20213 3568 20214 3632
rect 20148 3552 20214 3568
rect 20148 3488 20149 3552
rect 20213 3488 20214 3552
rect 20148 3472 20214 3488
rect 20148 3408 20149 3472
rect 20213 3408 20214 3472
rect 20148 3392 20214 3408
rect 20148 3328 20149 3392
rect 20213 3328 20214 3392
rect 20148 3312 20214 3328
rect 20148 3248 20149 3312
rect 20213 3248 20214 3312
rect 20148 3232 20214 3248
rect 20148 3168 20149 3232
rect 20213 3168 20214 3232
rect 20148 3152 20214 3168
rect 20148 3088 20149 3152
rect 20213 3088 20214 3152
rect 20148 3072 20214 3088
rect 20148 3008 20149 3072
rect 20213 3008 20214 3072
rect 20148 2992 20214 3008
rect 20148 2928 20149 2992
rect 20213 2928 20214 2992
rect 20148 2838 20214 2928
rect 20274 2834 20334 3866
rect 20394 2774 20454 3804
rect 20514 2834 20574 3866
rect 20634 2774 20694 3804
rect 20754 3712 20820 3866
rect 20754 3648 20755 3712
rect 20819 3648 20820 3712
rect 20754 3632 20820 3648
rect 20754 3568 20755 3632
rect 20819 3568 20820 3632
rect 20754 3552 20820 3568
rect 20754 3488 20755 3552
rect 20819 3488 20820 3552
rect 20754 3472 20820 3488
rect 20754 3408 20755 3472
rect 20819 3408 20820 3472
rect 20754 3392 20820 3408
rect 20754 3328 20755 3392
rect 20819 3328 20820 3392
rect 20754 3312 20820 3328
rect 20754 3248 20755 3312
rect 20819 3248 20820 3312
rect 20754 3232 20820 3248
rect 20754 3168 20755 3232
rect 20819 3168 20820 3232
rect 20754 3152 20820 3168
rect 20754 3088 20755 3152
rect 20819 3088 20820 3152
rect 20754 3072 20820 3088
rect 20754 3008 20755 3072
rect 20819 3008 20820 3072
rect 20754 2992 20820 3008
rect 20754 2928 20755 2992
rect 20819 2928 20820 2992
rect 20754 2838 20820 2928
rect 20880 2834 20940 3866
rect 21000 2774 21060 3804
rect 21120 2834 21180 3866
rect 21240 2774 21300 3804
rect 21360 3712 21426 3866
rect 21360 3648 21361 3712
rect 21425 3648 21426 3712
rect 21360 3632 21426 3648
rect 21360 3568 21361 3632
rect 21425 3568 21426 3632
rect 21360 3552 21426 3568
rect 21360 3488 21361 3552
rect 21425 3488 21426 3552
rect 21360 3472 21426 3488
rect 21360 3408 21361 3472
rect 21425 3408 21426 3472
rect 21360 3392 21426 3408
rect 21360 3328 21361 3392
rect 21425 3328 21426 3392
rect 21360 3312 21426 3328
rect 21360 3248 21361 3312
rect 21425 3248 21426 3312
rect 21360 3232 21426 3248
rect 21360 3168 21361 3232
rect 21425 3168 21426 3232
rect 21360 3152 21426 3168
rect 21360 3088 21361 3152
rect 21425 3088 21426 3152
rect 21360 3072 21426 3088
rect 21360 3008 21361 3072
rect 21425 3008 21426 3072
rect 21360 2992 21426 3008
rect 21360 2928 21361 2992
rect 21425 2928 21426 2992
rect 21360 2838 21426 2928
rect 21486 2834 21546 3866
rect 21606 2774 21666 3804
rect 21726 2834 21786 3866
rect 21846 2774 21906 3804
rect 21966 3712 22032 3866
rect 21966 3648 21967 3712
rect 22031 3648 22032 3712
rect 21966 3632 22032 3648
rect 21966 3568 21967 3632
rect 22031 3568 22032 3632
rect 21966 3552 22032 3568
rect 21966 3488 21967 3552
rect 22031 3488 22032 3552
rect 21966 3472 22032 3488
rect 21966 3408 21967 3472
rect 22031 3408 22032 3472
rect 21966 3392 22032 3408
rect 21966 3328 21967 3392
rect 22031 3328 22032 3392
rect 21966 3312 22032 3328
rect 21966 3248 21967 3312
rect 22031 3248 22032 3312
rect 21966 3232 22032 3248
rect 21966 3168 21967 3232
rect 22031 3168 22032 3232
rect 21966 3152 22032 3168
rect 21966 3088 21967 3152
rect 22031 3088 22032 3152
rect 21966 3072 22032 3088
rect 21966 3008 21967 3072
rect 22031 3008 22032 3072
rect 21966 2992 22032 3008
rect 21966 2928 21967 2992
rect 22031 2928 22032 2992
rect 21966 2838 22032 2928
rect 22092 2834 22152 3866
rect 22212 2774 22272 3804
rect 22332 2834 22392 3866
rect 22452 2774 22512 3804
rect 22572 3712 22638 3866
rect 22572 3648 22573 3712
rect 22637 3648 22638 3712
rect 22572 3632 22638 3648
rect 22572 3568 22573 3632
rect 22637 3568 22638 3632
rect 22572 3552 22638 3568
rect 22572 3488 22573 3552
rect 22637 3488 22638 3552
rect 22572 3472 22638 3488
rect 22572 3408 22573 3472
rect 22637 3408 22638 3472
rect 22572 3392 22638 3408
rect 22572 3328 22573 3392
rect 22637 3328 22638 3392
rect 22572 3312 22638 3328
rect 22572 3248 22573 3312
rect 22637 3248 22638 3312
rect 22572 3232 22638 3248
rect 22572 3168 22573 3232
rect 22637 3168 22638 3232
rect 22572 3152 22638 3168
rect 22572 3088 22573 3152
rect 22637 3088 22638 3152
rect 22572 3072 22638 3088
rect 22572 3008 22573 3072
rect 22637 3008 22638 3072
rect 22572 2992 22638 3008
rect 22572 2928 22573 2992
rect 22637 2928 22638 2992
rect 22572 2838 22638 2928
rect 22698 2834 22758 3866
rect 22818 2774 22878 3804
rect 22938 2834 22998 3866
rect 23058 2774 23118 3804
rect 23178 3712 23244 3866
rect 23178 3648 23179 3712
rect 23243 3648 23244 3712
rect 23178 3632 23244 3648
rect 23178 3568 23179 3632
rect 23243 3568 23244 3632
rect 23178 3552 23244 3568
rect 23178 3488 23179 3552
rect 23243 3488 23244 3552
rect 23178 3472 23244 3488
rect 23178 3408 23179 3472
rect 23243 3408 23244 3472
rect 23178 3392 23244 3408
rect 23178 3328 23179 3392
rect 23243 3328 23244 3392
rect 23178 3312 23244 3328
rect 23178 3248 23179 3312
rect 23243 3248 23244 3312
rect 23178 3232 23244 3248
rect 23178 3168 23179 3232
rect 23243 3168 23244 3232
rect 23178 3152 23244 3168
rect 23178 3088 23179 3152
rect 23243 3088 23244 3152
rect 23178 3072 23244 3088
rect 23178 3008 23179 3072
rect 23243 3008 23244 3072
rect 23178 2992 23244 3008
rect 23178 2928 23179 2992
rect 23243 2928 23244 2992
rect 23178 2838 23244 2928
rect 23304 2834 23364 3866
rect 23424 2774 23484 3804
rect 23544 2834 23604 3866
rect 23664 2774 23724 3804
rect 23784 3712 23850 3866
rect 23784 3648 23785 3712
rect 23849 3648 23850 3712
rect 23784 3632 23850 3648
rect 23784 3568 23785 3632
rect 23849 3568 23850 3632
rect 23784 3552 23850 3568
rect 23784 3488 23785 3552
rect 23849 3488 23850 3552
rect 23784 3472 23850 3488
rect 23784 3408 23785 3472
rect 23849 3408 23850 3472
rect 23784 3392 23850 3408
rect 23784 3328 23785 3392
rect 23849 3328 23850 3392
rect 23784 3312 23850 3328
rect 23784 3248 23785 3312
rect 23849 3248 23850 3312
rect 23784 3232 23850 3248
rect 23784 3168 23785 3232
rect 23849 3168 23850 3232
rect 23784 3152 23850 3168
rect 23784 3088 23785 3152
rect 23849 3088 23850 3152
rect 23784 3072 23850 3088
rect 23784 3008 23785 3072
rect 23849 3008 23850 3072
rect 23784 2992 23850 3008
rect 23784 2928 23785 2992
rect 23849 2928 23850 2992
rect 23784 2838 23850 2928
rect 23910 2834 23970 3866
rect 24030 2774 24090 3804
rect 24150 2834 24210 3866
rect 24270 2774 24330 3804
rect 24390 3712 24456 3866
rect 24390 3648 24391 3712
rect 24455 3648 24456 3712
rect 24390 3632 24456 3648
rect 24390 3568 24391 3632
rect 24455 3568 24456 3632
rect 24390 3552 24456 3568
rect 24390 3488 24391 3552
rect 24455 3488 24456 3552
rect 24390 3472 24456 3488
rect 24390 3408 24391 3472
rect 24455 3408 24456 3472
rect 24390 3392 24456 3408
rect 24390 3328 24391 3392
rect 24455 3328 24456 3392
rect 24390 3312 24456 3328
rect 24390 3248 24391 3312
rect 24455 3248 24456 3312
rect 24390 3232 24456 3248
rect 24390 3168 24391 3232
rect 24455 3168 24456 3232
rect 24390 3152 24456 3168
rect 24390 3088 24391 3152
rect 24455 3088 24456 3152
rect 24390 3072 24456 3088
rect 24390 3008 24391 3072
rect 24455 3008 24456 3072
rect 24390 2992 24456 3008
rect 24390 2928 24391 2992
rect 24455 2928 24456 2992
rect 24390 2838 24456 2928
rect 24516 2834 24576 3866
rect 24636 2774 24696 3804
rect 24756 2834 24816 3866
rect 24876 2774 24936 3804
rect 24996 3712 25062 3866
rect 24996 3648 24997 3712
rect 25061 3648 25062 3712
rect 24996 3632 25062 3648
rect 24996 3568 24997 3632
rect 25061 3568 25062 3632
rect 24996 3552 25062 3568
rect 24996 3488 24997 3552
rect 25061 3488 25062 3552
rect 24996 3472 25062 3488
rect 24996 3408 24997 3472
rect 25061 3408 25062 3472
rect 24996 3392 25062 3408
rect 24996 3328 24997 3392
rect 25061 3328 25062 3392
rect 24996 3312 25062 3328
rect 24996 3248 24997 3312
rect 25061 3248 25062 3312
rect 24996 3232 25062 3248
rect 24996 3168 24997 3232
rect 25061 3168 25062 3232
rect 24996 3152 25062 3168
rect 24996 3088 24997 3152
rect 25061 3088 25062 3152
rect 24996 3072 25062 3088
rect 24996 3008 24997 3072
rect 25061 3008 25062 3072
rect 24996 2992 25062 3008
rect 24996 2928 24997 2992
rect 25061 2928 25062 2992
rect 24996 2838 25062 2928
rect 25122 2834 25182 3866
rect 25242 2774 25302 3804
rect 25362 2834 25422 3866
rect 25482 2774 25542 3804
rect 25602 3712 25668 3866
rect 25602 3648 25603 3712
rect 25667 3648 25668 3712
rect 25602 3632 25668 3648
rect 25602 3568 25603 3632
rect 25667 3568 25668 3632
rect 25602 3552 25668 3568
rect 25602 3488 25603 3552
rect 25667 3488 25668 3552
rect 25602 3472 25668 3488
rect 25602 3408 25603 3472
rect 25667 3408 25668 3472
rect 25602 3392 25668 3408
rect 25602 3328 25603 3392
rect 25667 3328 25668 3392
rect 25602 3312 25668 3328
rect 25602 3248 25603 3312
rect 25667 3248 25668 3312
rect 25602 3232 25668 3248
rect 25602 3168 25603 3232
rect 25667 3168 25668 3232
rect 25602 3152 25668 3168
rect 25602 3088 25603 3152
rect 25667 3088 25668 3152
rect 25602 3072 25668 3088
rect 25602 3008 25603 3072
rect 25667 3008 25668 3072
rect 25602 2992 25668 3008
rect 25602 2928 25603 2992
rect 25667 2928 25668 2992
rect 25602 2838 25668 2928
rect 25728 2834 25788 3866
rect 25848 2774 25908 3804
rect 25968 2834 26028 3866
rect 26088 2774 26148 3804
rect 26208 3712 26274 3866
rect 26208 3648 26209 3712
rect 26273 3648 26274 3712
rect 26208 3632 26274 3648
rect 26208 3568 26209 3632
rect 26273 3568 26274 3632
rect 26208 3552 26274 3568
rect 26208 3488 26209 3552
rect 26273 3488 26274 3552
rect 26208 3472 26274 3488
rect 26208 3408 26209 3472
rect 26273 3408 26274 3472
rect 26208 3392 26274 3408
rect 26208 3328 26209 3392
rect 26273 3328 26274 3392
rect 26208 3312 26274 3328
rect 26208 3248 26209 3312
rect 26273 3248 26274 3312
rect 26208 3232 26274 3248
rect 26208 3168 26209 3232
rect 26273 3168 26274 3232
rect 26208 3152 26274 3168
rect 26208 3088 26209 3152
rect 26273 3088 26274 3152
rect 26208 3072 26274 3088
rect 26208 3008 26209 3072
rect 26273 3008 26274 3072
rect 26208 2992 26274 3008
rect 26208 2928 26209 2992
rect 26273 2928 26274 2992
rect 26208 2838 26274 2928
rect 26334 2834 26394 3866
rect 26454 2774 26514 3804
rect 26574 2834 26634 3866
rect 26694 2774 26754 3804
rect 26814 3712 26880 3866
rect 26814 3648 26815 3712
rect 26879 3648 26880 3712
rect 26814 3632 26880 3648
rect 26814 3568 26815 3632
rect 26879 3568 26880 3632
rect 26814 3552 26880 3568
rect 26814 3488 26815 3552
rect 26879 3488 26880 3552
rect 26814 3472 26880 3488
rect 26814 3408 26815 3472
rect 26879 3408 26880 3472
rect 26814 3392 26880 3408
rect 26814 3328 26815 3392
rect 26879 3328 26880 3392
rect 26814 3312 26880 3328
rect 26814 3248 26815 3312
rect 26879 3248 26880 3312
rect 26814 3232 26880 3248
rect 26814 3168 26815 3232
rect 26879 3168 26880 3232
rect 26814 3152 26880 3168
rect 26814 3088 26815 3152
rect 26879 3088 26880 3152
rect 26814 3072 26880 3088
rect 26814 3008 26815 3072
rect 26879 3008 26880 3072
rect 26814 2992 26880 3008
rect 26814 2928 26815 2992
rect 26879 2928 26880 2992
rect 26814 2838 26880 2928
rect 26940 2834 27000 3866
rect 27060 2774 27120 3804
rect 27180 2834 27240 3866
rect 27300 2774 27360 3804
rect 27420 3712 27486 3866
rect 27420 3648 27421 3712
rect 27485 3648 27486 3712
rect 27420 3632 27486 3648
rect 27420 3568 27421 3632
rect 27485 3568 27486 3632
rect 27420 3552 27486 3568
rect 27420 3488 27421 3552
rect 27485 3488 27486 3552
rect 27420 3472 27486 3488
rect 27420 3408 27421 3472
rect 27485 3408 27486 3472
rect 27420 3392 27486 3408
rect 27420 3328 27421 3392
rect 27485 3328 27486 3392
rect 27420 3312 27486 3328
rect 27420 3248 27421 3312
rect 27485 3248 27486 3312
rect 27420 3232 27486 3248
rect 27420 3168 27421 3232
rect 27485 3168 27486 3232
rect 27420 3152 27486 3168
rect 27420 3088 27421 3152
rect 27485 3088 27486 3152
rect 27420 3072 27486 3088
rect 27420 3008 27421 3072
rect 27485 3008 27486 3072
rect 27420 2992 27486 3008
rect 27420 2928 27421 2992
rect 27485 2928 27486 2992
rect 27420 2838 27486 2928
rect 27546 2834 27606 3866
rect 27666 2774 27726 3804
rect 27786 2834 27846 3866
rect 27906 2774 27966 3804
rect 28026 3712 28092 3866
rect 28026 3648 28027 3712
rect 28091 3648 28092 3712
rect 28026 3632 28092 3648
rect 28026 3568 28027 3632
rect 28091 3568 28092 3632
rect 28026 3552 28092 3568
rect 28026 3488 28027 3552
rect 28091 3488 28092 3552
rect 28026 3472 28092 3488
rect 28026 3408 28027 3472
rect 28091 3408 28092 3472
rect 28026 3392 28092 3408
rect 28026 3328 28027 3392
rect 28091 3328 28092 3392
rect 28026 3312 28092 3328
rect 28026 3248 28027 3312
rect 28091 3248 28092 3312
rect 28026 3232 28092 3248
rect 28026 3168 28027 3232
rect 28091 3168 28092 3232
rect 28026 3152 28092 3168
rect 28026 3088 28027 3152
rect 28091 3088 28092 3152
rect 28026 3072 28092 3088
rect 28026 3008 28027 3072
rect 28091 3008 28092 3072
rect 28026 2992 28092 3008
rect 28026 2928 28027 2992
rect 28091 2928 28092 2992
rect 28026 2838 28092 2928
rect 28152 2834 28212 3866
rect 28272 2774 28332 3804
rect 28392 2834 28452 3866
rect 28512 2774 28572 3804
rect 28632 3712 28698 3866
rect 28632 3648 28633 3712
rect 28697 3648 28698 3712
rect 28632 3632 28698 3648
rect 28632 3568 28633 3632
rect 28697 3568 28698 3632
rect 28632 3552 28698 3568
rect 28632 3488 28633 3552
rect 28697 3488 28698 3552
rect 28632 3472 28698 3488
rect 28632 3408 28633 3472
rect 28697 3408 28698 3472
rect 28632 3392 28698 3408
rect 28632 3328 28633 3392
rect 28697 3328 28698 3392
rect 28632 3312 28698 3328
rect 28632 3248 28633 3312
rect 28697 3248 28698 3312
rect 28632 3232 28698 3248
rect 28632 3168 28633 3232
rect 28697 3168 28698 3232
rect 28632 3152 28698 3168
rect 28632 3088 28633 3152
rect 28697 3088 28698 3152
rect 28632 3072 28698 3088
rect 28632 3008 28633 3072
rect 28697 3008 28698 3072
rect 28632 2992 28698 3008
rect 28632 2928 28633 2992
rect 28697 2928 28698 2992
rect 28632 2838 28698 2928
rect 28758 2834 28818 3866
rect 28878 2774 28938 3804
rect 28998 2834 29058 3866
rect 29118 2774 29178 3804
rect 29238 3712 29304 3866
rect 29238 3648 29239 3712
rect 29303 3648 29304 3712
rect 29238 3632 29304 3648
rect 29238 3568 29239 3632
rect 29303 3568 29304 3632
rect 29238 3552 29304 3568
rect 29238 3488 29239 3552
rect 29303 3488 29304 3552
rect 29238 3472 29304 3488
rect 29238 3408 29239 3472
rect 29303 3408 29304 3472
rect 29238 3392 29304 3408
rect 29238 3328 29239 3392
rect 29303 3328 29304 3392
rect 29238 3312 29304 3328
rect 29238 3248 29239 3312
rect 29303 3248 29304 3312
rect 29238 3232 29304 3248
rect 29238 3168 29239 3232
rect 29303 3168 29304 3232
rect 29238 3152 29304 3168
rect 29238 3088 29239 3152
rect 29303 3088 29304 3152
rect 29238 3072 29304 3088
rect 29238 3008 29239 3072
rect 29303 3008 29304 3072
rect 29238 2992 29304 3008
rect 29238 2928 29239 2992
rect 29303 2928 29304 2992
rect 29238 2838 29304 2928
rect 29364 2834 29424 3866
rect 29484 2774 29544 3804
rect 29604 2834 29664 3866
rect 29724 2774 29784 3804
rect 29844 3712 29910 3866
rect 29844 3648 29845 3712
rect 29909 3648 29910 3712
rect 29844 3632 29910 3648
rect 29844 3568 29845 3632
rect 29909 3568 29910 3632
rect 29844 3552 29910 3568
rect 29844 3488 29845 3552
rect 29909 3488 29910 3552
rect 29844 3472 29910 3488
rect 29844 3408 29845 3472
rect 29909 3408 29910 3472
rect 29844 3392 29910 3408
rect 29844 3328 29845 3392
rect 29909 3328 29910 3392
rect 29844 3312 29910 3328
rect 29844 3248 29845 3312
rect 29909 3248 29910 3312
rect 29844 3232 29910 3248
rect 29844 3168 29845 3232
rect 29909 3168 29910 3232
rect 29844 3152 29910 3168
rect 29844 3088 29845 3152
rect 29909 3088 29910 3152
rect 29844 3072 29910 3088
rect 29844 3008 29845 3072
rect 29909 3008 29910 3072
rect 29844 2992 29910 3008
rect 29844 2928 29845 2992
rect 29909 2928 29910 2992
rect 29844 2838 29910 2928
rect 29970 2834 30030 3866
rect 30090 2774 30150 3804
rect 30210 2834 30270 3866
rect 30330 2774 30390 3804
rect 30450 3712 30516 3866
rect 30450 3648 30451 3712
rect 30515 3648 30516 3712
rect 30450 3632 30516 3648
rect 30450 3568 30451 3632
rect 30515 3568 30516 3632
rect 30450 3552 30516 3568
rect 30450 3488 30451 3552
rect 30515 3488 30516 3552
rect 30450 3472 30516 3488
rect 30450 3408 30451 3472
rect 30515 3408 30516 3472
rect 30450 3392 30516 3408
rect 30450 3328 30451 3392
rect 30515 3328 30516 3392
rect 30450 3312 30516 3328
rect 30450 3248 30451 3312
rect 30515 3248 30516 3312
rect 30450 3232 30516 3248
rect 30450 3168 30451 3232
rect 30515 3168 30516 3232
rect 30450 3152 30516 3168
rect 30450 3088 30451 3152
rect 30515 3088 30516 3152
rect 30450 3072 30516 3088
rect 30450 3008 30451 3072
rect 30515 3008 30516 3072
rect 30450 2992 30516 3008
rect 30450 2928 30451 2992
rect 30515 2928 30516 2992
rect 30450 2838 30516 2928
rect 30576 2834 30636 3866
rect 30696 2774 30756 3804
rect 30816 2834 30876 3866
rect 30936 2774 30996 3804
rect 31056 3712 31122 3866
rect 31056 3648 31057 3712
rect 31121 3648 31122 3712
rect 31056 3632 31122 3648
rect 31056 3568 31057 3632
rect 31121 3568 31122 3632
rect 31056 3552 31122 3568
rect 31056 3488 31057 3552
rect 31121 3488 31122 3552
rect 31056 3472 31122 3488
rect 31056 3408 31057 3472
rect 31121 3408 31122 3472
rect 31056 3392 31122 3408
rect 31056 3328 31057 3392
rect 31121 3328 31122 3392
rect 31056 3312 31122 3328
rect 31056 3248 31057 3312
rect 31121 3248 31122 3312
rect 31056 3232 31122 3248
rect 31056 3168 31057 3232
rect 31121 3168 31122 3232
rect 31056 3152 31122 3168
rect 31056 3088 31057 3152
rect 31121 3088 31122 3152
rect 31056 3072 31122 3088
rect 31056 3008 31057 3072
rect 31121 3008 31122 3072
rect 31056 2992 31122 3008
rect 31056 2928 31057 2992
rect 31121 2928 31122 2992
rect 31056 2838 31122 2928
rect 31182 2834 31242 3866
rect 31302 2774 31362 3804
rect 31422 2834 31482 3866
rect 31542 2774 31602 3804
rect 31662 3712 31728 3866
rect 31662 3648 31663 3712
rect 31727 3648 31728 3712
rect 31662 3632 31728 3648
rect 31662 3568 31663 3632
rect 31727 3568 31728 3632
rect 31662 3552 31728 3568
rect 31662 3488 31663 3552
rect 31727 3488 31728 3552
rect 31662 3472 31728 3488
rect 31662 3408 31663 3472
rect 31727 3408 31728 3472
rect 31662 3392 31728 3408
rect 31662 3328 31663 3392
rect 31727 3328 31728 3392
rect 31662 3312 31728 3328
rect 31662 3248 31663 3312
rect 31727 3248 31728 3312
rect 31662 3232 31728 3248
rect 31662 3168 31663 3232
rect 31727 3168 31728 3232
rect 31662 3152 31728 3168
rect 31662 3088 31663 3152
rect 31727 3088 31728 3152
rect 31662 3072 31728 3088
rect 31662 3008 31663 3072
rect 31727 3008 31728 3072
rect 31662 2992 31728 3008
rect 31662 2928 31663 2992
rect 31727 2928 31728 2992
rect 31662 2838 31728 2928
rect 31788 2834 31848 3866
rect 31908 2774 31968 3804
rect 32028 2834 32088 3866
rect 32148 2774 32208 3804
rect 32268 3712 32334 3866
rect 32268 3648 32269 3712
rect 32333 3648 32334 3712
rect 32268 3632 32334 3648
rect 32268 3568 32269 3632
rect 32333 3568 32334 3632
rect 32268 3552 32334 3568
rect 32268 3488 32269 3552
rect 32333 3488 32334 3552
rect 32268 3472 32334 3488
rect 32268 3408 32269 3472
rect 32333 3408 32334 3472
rect 32268 3392 32334 3408
rect 32268 3328 32269 3392
rect 32333 3328 32334 3392
rect 32268 3312 32334 3328
rect 32268 3248 32269 3312
rect 32333 3248 32334 3312
rect 32268 3232 32334 3248
rect 32268 3168 32269 3232
rect 32333 3168 32334 3232
rect 32268 3152 32334 3168
rect 32268 3088 32269 3152
rect 32333 3088 32334 3152
rect 32268 3072 32334 3088
rect 32268 3008 32269 3072
rect 32333 3008 32334 3072
rect 32268 2992 32334 3008
rect 32268 2928 32269 2992
rect 32333 2928 32334 2992
rect 32268 2838 32334 2928
rect 32394 2834 32454 3866
rect 32514 2774 32574 3804
rect 32634 2834 32694 3866
rect 32754 2774 32814 3804
rect 32874 3712 32940 3866
rect 32874 3648 32875 3712
rect 32939 3648 32940 3712
rect 32874 3632 32940 3648
rect 32874 3568 32875 3632
rect 32939 3568 32940 3632
rect 32874 3552 32940 3568
rect 32874 3488 32875 3552
rect 32939 3488 32940 3552
rect 32874 3472 32940 3488
rect 32874 3408 32875 3472
rect 32939 3408 32940 3472
rect 32874 3392 32940 3408
rect 32874 3328 32875 3392
rect 32939 3328 32940 3392
rect 32874 3312 32940 3328
rect 32874 3248 32875 3312
rect 32939 3248 32940 3312
rect 32874 3232 32940 3248
rect 32874 3168 32875 3232
rect 32939 3168 32940 3232
rect 32874 3152 32940 3168
rect 32874 3088 32875 3152
rect 32939 3088 32940 3152
rect 32874 3072 32940 3088
rect 32874 3008 32875 3072
rect 32939 3008 32940 3072
rect 32874 2992 32940 3008
rect 32874 2928 32875 2992
rect 32939 2928 32940 2992
rect 32874 2838 32940 2928
rect 33000 2834 33060 3866
rect 33120 2774 33180 3804
rect 33240 2834 33300 3866
rect 33360 2774 33420 3804
rect 33480 3712 33546 3866
rect 33480 3648 33481 3712
rect 33545 3648 33546 3712
rect 33480 3632 33546 3648
rect 33480 3568 33481 3632
rect 33545 3568 33546 3632
rect 33480 3552 33546 3568
rect 33480 3488 33481 3552
rect 33545 3488 33546 3552
rect 33480 3472 33546 3488
rect 33480 3408 33481 3472
rect 33545 3408 33546 3472
rect 33480 3392 33546 3408
rect 33480 3328 33481 3392
rect 33545 3328 33546 3392
rect 33480 3312 33546 3328
rect 33480 3248 33481 3312
rect 33545 3248 33546 3312
rect 33480 3232 33546 3248
rect 33480 3168 33481 3232
rect 33545 3168 33546 3232
rect 33480 3152 33546 3168
rect 33480 3088 33481 3152
rect 33545 3088 33546 3152
rect 33480 3072 33546 3088
rect 33480 3008 33481 3072
rect 33545 3008 33546 3072
rect 33480 2992 33546 3008
rect 33480 2928 33481 2992
rect 33545 2928 33546 2992
rect 33480 2838 33546 2928
rect 33606 2834 33666 3866
rect 33726 2774 33786 3804
rect 33846 2834 33906 3866
rect 33966 2774 34026 3804
rect 34086 3712 34152 3866
rect 34086 3648 34087 3712
rect 34151 3648 34152 3712
rect 34086 3632 34152 3648
rect 34086 3568 34087 3632
rect 34151 3568 34152 3632
rect 34086 3552 34152 3568
rect 34086 3488 34087 3552
rect 34151 3488 34152 3552
rect 34086 3472 34152 3488
rect 34086 3408 34087 3472
rect 34151 3408 34152 3472
rect 34086 3392 34152 3408
rect 34086 3328 34087 3392
rect 34151 3328 34152 3392
rect 34086 3312 34152 3328
rect 34086 3248 34087 3312
rect 34151 3248 34152 3312
rect 34086 3232 34152 3248
rect 34086 3168 34087 3232
rect 34151 3168 34152 3232
rect 34086 3152 34152 3168
rect 34086 3088 34087 3152
rect 34151 3088 34152 3152
rect 34086 3072 34152 3088
rect 34086 3008 34087 3072
rect 34151 3008 34152 3072
rect 34086 2992 34152 3008
rect 34086 2928 34087 2992
rect 34151 2928 34152 2992
rect 34086 2838 34152 2928
rect 34212 2834 34272 3866
rect 34332 2774 34392 3804
rect 34452 2834 34512 3866
rect 34572 2774 34632 3804
rect 34692 3712 34758 3866
rect 34692 3648 34693 3712
rect 34757 3648 34758 3712
rect 34692 3632 34758 3648
rect 34692 3568 34693 3632
rect 34757 3568 34758 3632
rect 34692 3552 34758 3568
rect 34692 3488 34693 3552
rect 34757 3488 34758 3552
rect 34692 3472 34758 3488
rect 34692 3408 34693 3472
rect 34757 3408 34758 3472
rect 34692 3392 34758 3408
rect 34692 3328 34693 3392
rect 34757 3328 34758 3392
rect 34692 3312 34758 3328
rect 34692 3248 34693 3312
rect 34757 3248 34758 3312
rect 34692 3232 34758 3248
rect 34692 3168 34693 3232
rect 34757 3168 34758 3232
rect 34692 3152 34758 3168
rect 34692 3088 34693 3152
rect 34757 3088 34758 3152
rect 34692 3072 34758 3088
rect 34692 3008 34693 3072
rect 34757 3008 34758 3072
rect 34692 2992 34758 3008
rect 34692 2928 34693 2992
rect 34757 2928 34758 2992
rect 34692 2838 34758 2928
rect 34818 2834 34878 3866
rect 34938 2774 34998 3804
rect 35058 2834 35118 3866
rect 35178 2774 35238 3804
rect 35298 3712 35364 3866
rect 35298 3648 35299 3712
rect 35363 3648 35364 3712
rect 35298 3632 35364 3648
rect 35298 3568 35299 3632
rect 35363 3568 35364 3632
rect 35298 3552 35364 3568
rect 35298 3488 35299 3552
rect 35363 3488 35364 3552
rect 35298 3472 35364 3488
rect 35298 3408 35299 3472
rect 35363 3408 35364 3472
rect 35298 3392 35364 3408
rect 35298 3328 35299 3392
rect 35363 3328 35364 3392
rect 35298 3312 35364 3328
rect 35298 3248 35299 3312
rect 35363 3248 35364 3312
rect 35298 3232 35364 3248
rect 35298 3168 35299 3232
rect 35363 3168 35364 3232
rect 35298 3152 35364 3168
rect 35298 3088 35299 3152
rect 35363 3088 35364 3152
rect 35298 3072 35364 3088
rect 35298 3008 35299 3072
rect 35363 3008 35364 3072
rect 35298 2992 35364 3008
rect 35298 2928 35299 2992
rect 35363 2928 35364 2992
rect 35298 2838 35364 2928
rect 35424 2834 35484 3866
rect 35544 2774 35604 3804
rect 35664 2834 35724 3866
rect 35784 2774 35844 3804
rect 35904 3712 35970 3866
rect 35904 3648 35905 3712
rect 35969 3648 35970 3712
rect 35904 3632 35970 3648
rect 35904 3568 35905 3632
rect 35969 3568 35970 3632
rect 35904 3552 35970 3568
rect 35904 3488 35905 3552
rect 35969 3488 35970 3552
rect 35904 3472 35970 3488
rect 35904 3408 35905 3472
rect 35969 3408 35970 3472
rect 35904 3392 35970 3408
rect 35904 3328 35905 3392
rect 35969 3328 35970 3392
rect 35904 3312 35970 3328
rect 35904 3248 35905 3312
rect 35969 3248 35970 3312
rect 35904 3232 35970 3248
rect 35904 3168 35905 3232
rect 35969 3168 35970 3232
rect 35904 3152 35970 3168
rect 35904 3088 35905 3152
rect 35969 3088 35970 3152
rect 35904 3072 35970 3088
rect 35904 3008 35905 3072
rect 35969 3008 35970 3072
rect 35904 2992 35970 3008
rect 35904 2928 35905 2992
rect 35969 2928 35970 2992
rect 35904 2838 35970 2928
rect 36030 2834 36090 3866
rect 36150 2774 36210 3804
rect 36270 2834 36330 3866
rect 36390 2774 36450 3804
rect 36510 3712 36576 3866
rect 36510 3648 36511 3712
rect 36575 3648 36576 3712
rect 36510 3632 36576 3648
rect 36510 3568 36511 3632
rect 36575 3568 36576 3632
rect 36510 3552 36576 3568
rect 36510 3488 36511 3552
rect 36575 3488 36576 3552
rect 36510 3472 36576 3488
rect 36510 3408 36511 3472
rect 36575 3408 36576 3472
rect 36510 3392 36576 3408
rect 36510 3328 36511 3392
rect 36575 3328 36576 3392
rect 36510 3312 36576 3328
rect 36510 3248 36511 3312
rect 36575 3248 36576 3312
rect 36510 3232 36576 3248
rect 36510 3168 36511 3232
rect 36575 3168 36576 3232
rect 36510 3152 36576 3168
rect 36510 3088 36511 3152
rect 36575 3088 36576 3152
rect 36510 3072 36576 3088
rect 36510 3008 36511 3072
rect 36575 3008 36576 3072
rect 36510 2992 36576 3008
rect 36510 2928 36511 2992
rect 36575 2928 36576 2992
rect 36510 2838 36576 2928
rect 36636 2834 36696 3866
rect 36756 2774 36816 3804
rect 36876 2834 36936 3866
rect 36996 2774 37056 3804
rect 37116 3712 37182 3866
rect 37116 3648 37117 3712
rect 37181 3648 37182 3712
rect 37116 3632 37182 3648
rect 37116 3568 37117 3632
rect 37181 3568 37182 3632
rect 37116 3552 37182 3568
rect 37116 3488 37117 3552
rect 37181 3488 37182 3552
rect 37116 3472 37182 3488
rect 37116 3408 37117 3472
rect 37181 3408 37182 3472
rect 37116 3392 37182 3408
rect 37116 3328 37117 3392
rect 37181 3328 37182 3392
rect 37116 3312 37182 3328
rect 37116 3248 37117 3312
rect 37181 3248 37182 3312
rect 37116 3232 37182 3248
rect 37116 3168 37117 3232
rect 37181 3168 37182 3232
rect 37116 3152 37182 3168
rect 37116 3088 37117 3152
rect 37181 3088 37182 3152
rect 37116 3072 37182 3088
rect 37116 3008 37117 3072
rect 37181 3008 37182 3072
rect 37116 2992 37182 3008
rect 37116 2928 37117 2992
rect 37181 2928 37182 2992
rect 37116 2838 37182 2928
rect 37242 2834 37302 3866
rect 37362 2774 37422 3804
rect 37482 2834 37542 3866
rect 37602 2774 37662 3804
rect 37722 3712 37788 3866
rect 37722 3648 37723 3712
rect 37787 3648 37788 3712
rect 37722 3632 37788 3648
rect 37722 3568 37723 3632
rect 37787 3568 37788 3632
rect 37722 3552 37788 3568
rect 37722 3488 37723 3552
rect 37787 3488 37788 3552
rect 37722 3472 37788 3488
rect 37722 3408 37723 3472
rect 37787 3408 37788 3472
rect 37722 3392 37788 3408
rect 37722 3328 37723 3392
rect 37787 3328 37788 3392
rect 37722 3312 37788 3328
rect 37722 3248 37723 3312
rect 37787 3248 37788 3312
rect 37722 3232 37788 3248
rect 37722 3168 37723 3232
rect 37787 3168 37788 3232
rect 37722 3152 37788 3168
rect 37722 3088 37723 3152
rect 37787 3088 37788 3152
rect 37722 3072 37788 3088
rect 37722 3008 37723 3072
rect 37787 3008 37788 3072
rect 37722 2992 37788 3008
rect 37722 2928 37723 2992
rect 37787 2928 37788 2992
rect 37722 2838 37788 2928
rect 37848 2834 37908 3866
rect 37968 2774 38028 3804
rect 38088 2834 38148 3866
rect 38208 2774 38268 3804
rect 38328 3712 38394 3866
rect 38328 3648 38329 3712
rect 38393 3648 38394 3712
rect 38328 3632 38394 3648
rect 38328 3568 38329 3632
rect 38393 3568 38394 3632
rect 38328 3552 38394 3568
rect 38328 3488 38329 3552
rect 38393 3488 38394 3552
rect 38328 3472 38394 3488
rect 38328 3408 38329 3472
rect 38393 3408 38394 3472
rect 38328 3392 38394 3408
rect 38328 3328 38329 3392
rect 38393 3328 38394 3392
rect 38328 3312 38394 3328
rect 38328 3248 38329 3312
rect 38393 3248 38394 3312
rect 38328 3232 38394 3248
rect 38328 3168 38329 3232
rect 38393 3168 38394 3232
rect 38328 3152 38394 3168
rect 38328 3088 38329 3152
rect 38393 3088 38394 3152
rect 38328 3072 38394 3088
rect 38328 3008 38329 3072
rect 38393 3008 38394 3072
rect 38328 2992 38394 3008
rect 38328 2928 38329 2992
rect 38393 2928 38394 2992
rect 38328 2838 38394 2928
rect 38454 2834 38514 3866
rect 38574 2774 38634 3804
rect 38694 2834 38754 3866
rect 38814 2774 38874 3804
rect 38934 3712 39000 3866
rect 38934 3648 38935 3712
rect 38999 3648 39000 3712
rect 38934 3632 39000 3648
rect 38934 3568 38935 3632
rect 38999 3568 39000 3632
rect 38934 3552 39000 3568
rect 38934 3488 38935 3552
rect 38999 3488 39000 3552
rect 38934 3472 39000 3488
rect 38934 3408 38935 3472
rect 38999 3408 39000 3472
rect 38934 3392 39000 3408
rect 38934 3328 38935 3392
rect 38999 3328 39000 3392
rect 38934 3312 39000 3328
rect 38934 3248 38935 3312
rect 38999 3248 39000 3312
rect 38934 3232 39000 3248
rect 38934 3168 38935 3232
rect 38999 3168 39000 3232
rect 38934 3152 39000 3168
rect 38934 3088 38935 3152
rect 38999 3088 39000 3152
rect 38934 3072 39000 3088
rect 38934 3008 38935 3072
rect 38999 3008 39000 3072
rect 38934 2992 39000 3008
rect 38934 2928 38935 2992
rect 38999 2928 39000 2992
rect 38934 2838 39000 2928
rect 39060 2834 39120 3866
rect 39180 2774 39240 3804
rect 39300 2834 39360 3866
rect 39420 2774 39480 3804
rect 39540 3712 39606 3866
rect 39540 3648 39541 3712
rect 39605 3648 39606 3712
rect 39540 3632 39606 3648
rect 39540 3568 39541 3632
rect 39605 3568 39606 3632
rect 39540 3552 39606 3568
rect 39540 3488 39541 3552
rect 39605 3488 39606 3552
rect 39540 3472 39606 3488
rect 39540 3408 39541 3472
rect 39605 3408 39606 3472
rect 39540 3392 39606 3408
rect 39540 3328 39541 3392
rect 39605 3328 39606 3392
rect 39540 3312 39606 3328
rect 39540 3248 39541 3312
rect 39605 3248 39606 3312
rect 39540 3232 39606 3248
rect 39540 3168 39541 3232
rect 39605 3168 39606 3232
rect 39540 3152 39606 3168
rect 39540 3088 39541 3152
rect 39605 3088 39606 3152
rect 39540 3072 39606 3088
rect 39540 3008 39541 3072
rect 39605 3008 39606 3072
rect 39540 2992 39606 3008
rect 39540 2928 39541 2992
rect 39605 2928 39606 2992
rect 39540 2838 39606 2928
rect -459 2772 213 2774
rect -459 2708 -355 2772
rect -291 2708 -275 2772
rect -211 2708 -195 2772
rect -131 2708 -115 2772
rect -51 2708 -35 2772
rect 29 2708 45 2772
rect 109 2708 213 2772
rect -459 2706 213 2708
rect 524 2772 1027 2774
rect 524 2708 539 2772
rect 603 2708 619 2772
rect 683 2708 699 2772
rect 763 2708 779 2772
rect 843 2708 859 2772
rect 923 2708 1027 2772
rect 524 2706 1027 2708
rect 1267 2772 1717 2774
rect 1954 2772 2545 2774
rect 1267 2708 1371 2772
rect 1435 2708 1451 2772
rect 1515 2708 1531 2772
rect 1595 2708 1611 2772
rect 1675 2708 1691 2772
rect 1954 2708 1977 2772
rect 2041 2708 2057 2772
rect 2121 2708 2137 2772
rect 2201 2708 2217 2772
rect 2281 2708 2297 2772
rect 2361 2708 2377 2772
rect 2441 2708 2545 2772
rect 1267 2706 1717 2708
rect 1954 2706 2545 2708
rect 2801 2772 3301 2774
rect 3538 2772 5291 2774
rect 2801 2708 2905 2772
rect 2969 2708 2985 2772
rect 3049 2708 3065 2772
rect 3129 2708 3145 2772
rect 3209 2708 3225 2772
rect 3289 2708 3301 2772
rect 3575 2708 3591 2772
rect 3655 2708 3671 2772
rect 3735 2708 3751 2772
rect 3815 2708 3831 2772
rect 3895 2708 3911 2772
rect 3975 2708 4117 2772
rect 4181 2708 4197 2772
rect 4261 2708 4277 2772
rect 4341 2708 4357 2772
rect 4421 2708 4437 2772
rect 4501 2708 4517 2772
rect 4581 2708 4723 2772
rect 4787 2708 4803 2772
rect 4867 2708 4883 2772
rect 4947 2708 4963 2772
rect 5027 2708 5043 2772
rect 5107 2708 5123 2772
rect 5187 2708 5291 2772
rect 2801 2706 3301 2708
rect 3538 2706 5291 2708
rect 5352 2706 5394 2774
rect 5631 2772 10266 2774
rect 5680 2708 5696 2772
rect 5760 2708 5776 2772
rect 5840 2708 5856 2772
rect 5920 2708 6062 2772
rect 6126 2708 6142 2772
rect 6206 2708 6222 2772
rect 6286 2708 6302 2772
rect 6366 2708 6382 2772
rect 6446 2708 6462 2772
rect 6526 2708 6668 2772
rect 6732 2708 6748 2772
rect 6812 2708 6828 2772
rect 6892 2708 6908 2772
rect 6972 2708 6988 2772
rect 7052 2708 7068 2772
rect 7132 2708 7274 2772
rect 7338 2708 7354 2772
rect 7418 2708 7434 2772
rect 7498 2708 7514 2772
rect 7578 2708 7594 2772
rect 7658 2708 7674 2772
rect 7738 2708 7880 2772
rect 7944 2708 7960 2772
rect 8024 2708 8040 2772
rect 8104 2708 8120 2772
rect 8184 2708 8200 2772
rect 8264 2708 8280 2772
rect 8344 2708 8486 2772
rect 8550 2708 8566 2772
rect 8630 2708 8646 2772
rect 8710 2708 8726 2772
rect 8790 2708 8806 2772
rect 8870 2708 8886 2772
rect 8950 2708 9092 2772
rect 9156 2708 9172 2772
rect 9236 2708 9252 2772
rect 9316 2708 9332 2772
rect 9396 2708 9412 2772
rect 9476 2708 9492 2772
rect 9556 2708 9698 2772
rect 9762 2708 9778 2772
rect 9842 2708 9858 2772
rect 9922 2708 9938 2772
rect 10002 2708 10018 2772
rect 10082 2708 10098 2772
rect 10162 2708 10266 2772
rect 5631 2706 10266 2708
rect 10326 2706 10368 2774
rect 10605 2772 20088 2774
rect 10654 2708 10670 2772
rect 10734 2708 10750 2772
rect 10814 2708 10830 2772
rect 10894 2708 11036 2772
rect 11100 2708 11116 2772
rect 11180 2708 11196 2772
rect 11260 2708 11276 2772
rect 11340 2708 11356 2772
rect 11420 2708 11436 2772
rect 11500 2708 11642 2772
rect 11706 2708 11722 2772
rect 11786 2708 11802 2772
rect 11866 2708 11882 2772
rect 11946 2708 11962 2772
rect 12026 2708 12042 2772
rect 12106 2708 12248 2772
rect 12312 2708 12328 2772
rect 12392 2708 12408 2772
rect 12472 2708 12488 2772
rect 12552 2708 12568 2772
rect 12632 2708 12648 2772
rect 12712 2708 12854 2772
rect 12918 2708 12934 2772
rect 12998 2708 13014 2772
rect 13078 2708 13094 2772
rect 13158 2708 13174 2772
rect 13238 2708 13254 2772
rect 13318 2708 13460 2772
rect 13524 2708 13540 2772
rect 13604 2708 13620 2772
rect 13684 2708 13700 2772
rect 13764 2708 13780 2772
rect 13844 2708 13860 2772
rect 13924 2708 14066 2772
rect 14130 2708 14146 2772
rect 14210 2708 14226 2772
rect 14290 2708 14306 2772
rect 14370 2708 14386 2772
rect 14450 2708 14466 2772
rect 14530 2708 14672 2772
rect 14736 2708 14752 2772
rect 14816 2708 14832 2772
rect 14896 2708 14912 2772
rect 14976 2708 14992 2772
rect 15056 2708 15072 2772
rect 15136 2708 15278 2772
rect 15342 2708 15358 2772
rect 15422 2708 15438 2772
rect 15502 2708 15518 2772
rect 15582 2708 15598 2772
rect 15662 2708 15678 2772
rect 15742 2708 15884 2772
rect 15948 2708 15964 2772
rect 16028 2708 16044 2772
rect 16108 2708 16124 2772
rect 16188 2708 16204 2772
rect 16268 2708 16284 2772
rect 16348 2708 16490 2772
rect 16554 2708 16570 2772
rect 16634 2708 16650 2772
rect 16714 2708 16730 2772
rect 16794 2708 16810 2772
rect 16874 2708 16890 2772
rect 16954 2708 17096 2772
rect 17160 2708 17176 2772
rect 17240 2708 17256 2772
rect 17320 2708 17336 2772
rect 17400 2708 17416 2772
rect 17480 2708 17496 2772
rect 17560 2708 17702 2772
rect 17766 2708 17782 2772
rect 17846 2708 17862 2772
rect 17926 2708 17942 2772
rect 18006 2708 18022 2772
rect 18086 2708 18102 2772
rect 18166 2708 18308 2772
rect 18372 2708 18388 2772
rect 18452 2708 18468 2772
rect 18532 2708 18548 2772
rect 18612 2708 18628 2772
rect 18692 2708 18708 2772
rect 18772 2708 18914 2772
rect 18978 2708 18994 2772
rect 19058 2708 19074 2772
rect 19138 2708 19154 2772
rect 19218 2708 19234 2772
rect 19298 2708 19314 2772
rect 19378 2708 19520 2772
rect 19584 2708 19600 2772
rect 19664 2708 19680 2772
rect 19744 2708 19760 2772
rect 19824 2708 19840 2772
rect 19904 2708 19920 2772
rect 19984 2708 20088 2772
rect 10605 2706 20088 2708
rect 20148 2772 39298 2774
rect 20148 2708 20252 2772
rect 20316 2708 20332 2772
rect 20396 2708 20412 2772
rect 20476 2708 20492 2772
rect 20556 2708 20572 2772
rect 20636 2708 20652 2772
rect 20716 2708 20858 2772
rect 20922 2708 20938 2772
rect 21002 2708 21018 2772
rect 21082 2708 21098 2772
rect 21162 2708 21178 2772
rect 21242 2708 21258 2772
rect 21322 2708 21464 2772
rect 21528 2708 21544 2772
rect 21608 2708 21624 2772
rect 21688 2708 21704 2772
rect 21768 2708 21784 2772
rect 21848 2708 21864 2772
rect 21928 2708 22070 2772
rect 22134 2708 22150 2772
rect 22214 2708 22230 2772
rect 22294 2708 22310 2772
rect 22374 2708 22390 2772
rect 22454 2708 22470 2772
rect 22534 2708 22676 2772
rect 22740 2708 22756 2772
rect 22820 2708 22836 2772
rect 22900 2708 22916 2772
rect 22980 2708 22996 2772
rect 23060 2708 23076 2772
rect 23140 2708 23282 2772
rect 23346 2708 23362 2772
rect 23426 2708 23442 2772
rect 23506 2708 23522 2772
rect 23586 2708 23602 2772
rect 23666 2708 23682 2772
rect 23746 2708 23888 2772
rect 23952 2708 23968 2772
rect 24032 2708 24048 2772
rect 24112 2708 24128 2772
rect 24192 2708 24208 2772
rect 24272 2708 24288 2772
rect 24352 2708 24494 2772
rect 24558 2708 24574 2772
rect 24638 2708 24654 2772
rect 24718 2708 24734 2772
rect 24798 2708 24814 2772
rect 24878 2708 24894 2772
rect 24958 2708 25100 2772
rect 25164 2708 25180 2772
rect 25244 2708 25260 2772
rect 25324 2708 25340 2772
rect 25404 2708 25420 2772
rect 25484 2708 25500 2772
rect 25564 2708 25706 2772
rect 25770 2708 25786 2772
rect 25850 2708 25866 2772
rect 25930 2708 25946 2772
rect 26010 2708 26026 2772
rect 26090 2708 26106 2772
rect 26170 2708 26312 2772
rect 26376 2708 26392 2772
rect 26456 2708 26472 2772
rect 26536 2708 26552 2772
rect 26616 2708 26632 2772
rect 26696 2708 26712 2772
rect 26776 2708 26918 2772
rect 26982 2708 26998 2772
rect 27062 2708 27078 2772
rect 27142 2708 27158 2772
rect 27222 2708 27238 2772
rect 27302 2708 27318 2772
rect 27382 2708 27524 2772
rect 27588 2708 27604 2772
rect 27668 2708 27684 2772
rect 27748 2708 27764 2772
rect 27828 2708 27844 2772
rect 27908 2708 27924 2772
rect 27988 2708 28130 2772
rect 28194 2708 28210 2772
rect 28274 2708 28290 2772
rect 28354 2708 28370 2772
rect 28434 2708 28450 2772
rect 28514 2708 28530 2772
rect 28594 2708 28736 2772
rect 28800 2708 28816 2772
rect 28880 2708 28896 2772
rect 28960 2708 28976 2772
rect 29040 2708 29056 2772
rect 29120 2708 29136 2772
rect 29200 2708 29342 2772
rect 29406 2708 29422 2772
rect 29486 2708 29502 2772
rect 29566 2708 29582 2772
rect 29646 2708 29662 2772
rect 29726 2708 29742 2772
rect 29806 2708 29948 2772
rect 30012 2708 30028 2772
rect 30092 2708 30108 2772
rect 30172 2708 30188 2772
rect 30252 2708 30268 2772
rect 30332 2708 30348 2772
rect 30412 2708 30554 2772
rect 30618 2708 30634 2772
rect 30698 2708 30714 2772
rect 30778 2708 30794 2772
rect 30858 2708 30874 2772
rect 30938 2708 30954 2772
rect 31018 2708 31160 2772
rect 31224 2708 31240 2772
rect 31304 2708 31320 2772
rect 31384 2708 31400 2772
rect 31464 2708 31480 2772
rect 31544 2708 31560 2772
rect 31624 2708 31766 2772
rect 31830 2708 31846 2772
rect 31910 2708 31926 2772
rect 31990 2708 32006 2772
rect 32070 2708 32086 2772
rect 32150 2708 32166 2772
rect 32230 2708 32372 2772
rect 32436 2708 32452 2772
rect 32516 2708 32532 2772
rect 32596 2708 32612 2772
rect 32676 2708 32692 2772
rect 32756 2708 32772 2772
rect 32836 2708 32978 2772
rect 33042 2708 33058 2772
rect 33122 2708 33138 2772
rect 33202 2708 33218 2772
rect 33282 2708 33298 2772
rect 33362 2708 33378 2772
rect 33442 2708 33584 2772
rect 33648 2708 33664 2772
rect 33728 2708 33744 2772
rect 33808 2708 33824 2772
rect 33888 2708 33904 2772
rect 33968 2708 33984 2772
rect 34048 2708 34190 2772
rect 34254 2708 34270 2772
rect 34334 2708 34350 2772
rect 34414 2708 34430 2772
rect 34494 2708 34510 2772
rect 34574 2708 34590 2772
rect 34654 2708 34796 2772
rect 34860 2708 34876 2772
rect 34940 2708 34956 2772
rect 35020 2708 35036 2772
rect 35100 2708 35116 2772
rect 35180 2708 35196 2772
rect 35260 2708 35402 2772
rect 35466 2708 35482 2772
rect 35546 2708 35562 2772
rect 35626 2708 35642 2772
rect 35706 2708 35722 2772
rect 35786 2708 35802 2772
rect 35866 2708 36008 2772
rect 36072 2708 36088 2772
rect 36152 2708 36168 2772
rect 36232 2708 36248 2772
rect 36312 2708 36328 2772
rect 36392 2708 36408 2772
rect 36472 2708 36614 2772
rect 36678 2708 36694 2772
rect 36758 2708 36774 2772
rect 36838 2708 36854 2772
rect 36918 2708 36934 2772
rect 36998 2708 37014 2772
rect 37078 2708 37220 2772
rect 37284 2708 37300 2772
rect 37364 2708 37380 2772
rect 37444 2708 37460 2772
rect 37524 2708 37540 2772
rect 37604 2708 37620 2772
rect 37684 2708 37826 2772
rect 37890 2708 37906 2772
rect 37970 2708 37986 2772
rect 38050 2708 38066 2772
rect 38130 2708 38146 2772
rect 38210 2708 38226 2772
rect 38290 2708 38432 2772
rect 38496 2708 38512 2772
rect 38576 2708 38592 2772
rect 38656 2708 38672 2772
rect 38736 2708 38752 2772
rect 38816 2708 38832 2772
rect 38896 2708 39038 2772
rect 39102 2708 39118 2772
rect 39182 2708 39198 2772
rect 39262 2708 39278 2772
rect 20148 2706 39298 2708
rect 39534 2706 39606 2774
rect -459 1959 213 1961
rect -459 1895 -355 1959
rect -291 1895 -275 1959
rect -211 1895 -195 1959
rect -131 1895 -115 1959
rect -51 1895 -35 1959
rect 29 1895 45 1959
rect 109 1895 213 1959
rect -459 1893 213 1895
rect 524 1959 1027 1961
rect 524 1895 539 1959
rect 603 1895 619 1959
rect 683 1895 699 1959
rect 763 1895 779 1959
rect 843 1895 859 1959
rect 923 1895 1027 1959
rect 524 1893 1027 1895
rect 1267 1959 1717 1961
rect 1954 1959 2545 1961
rect 1267 1895 1371 1959
rect 1435 1895 1451 1959
rect 1515 1895 1531 1959
rect 1595 1895 1611 1959
rect 1675 1895 1691 1959
rect 1954 1895 1977 1959
rect 2041 1895 2057 1959
rect 2121 1895 2137 1959
rect 2201 1895 2217 1959
rect 2281 1895 2297 1959
rect 2361 1895 2377 1959
rect 2441 1895 2545 1959
rect 1267 1893 1717 1895
rect 1954 1893 2545 1895
rect 2801 1959 3301 1961
rect 3538 1959 5291 1961
rect 2801 1895 2905 1959
rect 2969 1895 2985 1959
rect 3049 1895 3065 1959
rect 3129 1895 3145 1959
rect 3209 1895 3225 1959
rect 3289 1895 3301 1959
rect 3575 1895 3591 1959
rect 3655 1895 3671 1959
rect 3735 1895 3751 1959
rect 3815 1895 3831 1959
rect 3895 1895 3911 1959
rect 3975 1895 4117 1959
rect 4181 1895 4197 1959
rect 4261 1895 4277 1959
rect 4341 1895 4357 1959
rect 4421 1895 4437 1959
rect 4501 1895 4517 1959
rect 4581 1895 4723 1959
rect 4787 1895 4803 1959
rect 4867 1895 4883 1959
rect 4947 1895 4963 1959
rect 5027 1895 5043 1959
rect 5107 1895 5123 1959
rect 5187 1895 5291 1959
rect 2801 1893 3301 1895
rect 3538 1893 5291 1895
rect 5352 1893 5394 1961
rect 5631 1959 10266 1961
rect 5680 1895 5696 1959
rect 5760 1895 5776 1959
rect 5840 1895 5856 1959
rect 5920 1895 6062 1959
rect 6126 1895 6142 1959
rect 6206 1895 6222 1959
rect 6286 1895 6302 1959
rect 6366 1895 6382 1959
rect 6446 1895 6462 1959
rect 6526 1895 6668 1959
rect 6732 1895 6748 1959
rect 6812 1895 6828 1959
rect 6892 1895 6908 1959
rect 6972 1895 6988 1959
rect 7052 1895 7068 1959
rect 7132 1895 7274 1959
rect 7338 1895 7354 1959
rect 7418 1895 7434 1959
rect 7498 1895 7514 1959
rect 7578 1895 7594 1959
rect 7658 1895 7674 1959
rect 7738 1895 7880 1959
rect 7944 1895 7960 1959
rect 8024 1895 8040 1959
rect 8104 1895 8120 1959
rect 8184 1895 8200 1959
rect 8264 1895 8280 1959
rect 8344 1895 8486 1959
rect 8550 1895 8566 1959
rect 8630 1895 8646 1959
rect 8710 1895 8726 1959
rect 8790 1895 8806 1959
rect 8870 1895 8886 1959
rect 8950 1895 9092 1959
rect 9156 1895 9172 1959
rect 9236 1895 9252 1959
rect 9316 1895 9332 1959
rect 9396 1895 9412 1959
rect 9476 1895 9492 1959
rect 9556 1895 9698 1959
rect 9762 1895 9778 1959
rect 9842 1895 9858 1959
rect 9922 1895 9938 1959
rect 10002 1895 10018 1959
rect 10082 1895 10098 1959
rect 10162 1895 10266 1959
rect 5631 1893 10266 1895
rect 10326 1893 10368 1961
rect 10605 1959 20088 1961
rect 10654 1895 10670 1959
rect 10734 1895 10750 1959
rect 10814 1895 10830 1959
rect 10894 1895 11036 1959
rect 11100 1895 11116 1959
rect 11180 1895 11196 1959
rect 11260 1895 11276 1959
rect 11340 1895 11356 1959
rect 11420 1895 11436 1959
rect 11500 1895 11642 1959
rect 11706 1895 11722 1959
rect 11786 1895 11802 1959
rect 11866 1895 11882 1959
rect 11946 1895 11962 1959
rect 12026 1895 12042 1959
rect 12106 1895 12248 1959
rect 12312 1895 12328 1959
rect 12392 1895 12408 1959
rect 12472 1895 12488 1959
rect 12552 1895 12568 1959
rect 12632 1895 12648 1959
rect 12712 1895 12854 1959
rect 12918 1895 12934 1959
rect 12998 1895 13014 1959
rect 13078 1895 13094 1959
rect 13158 1895 13174 1959
rect 13238 1895 13254 1959
rect 13318 1895 13460 1959
rect 13524 1895 13540 1959
rect 13604 1895 13620 1959
rect 13684 1895 13700 1959
rect 13764 1895 13780 1959
rect 13844 1895 13860 1959
rect 13924 1895 14066 1959
rect 14130 1895 14146 1959
rect 14210 1895 14226 1959
rect 14290 1895 14306 1959
rect 14370 1895 14386 1959
rect 14450 1895 14466 1959
rect 14530 1895 14672 1959
rect 14736 1895 14752 1959
rect 14816 1895 14832 1959
rect 14896 1895 14912 1959
rect 14976 1895 14992 1959
rect 15056 1895 15072 1959
rect 15136 1895 15278 1959
rect 15342 1895 15358 1959
rect 15422 1895 15438 1959
rect 15502 1895 15518 1959
rect 15582 1895 15598 1959
rect 15662 1895 15678 1959
rect 15742 1895 15884 1959
rect 15948 1895 15964 1959
rect 16028 1895 16044 1959
rect 16108 1895 16124 1959
rect 16188 1895 16204 1959
rect 16268 1895 16284 1959
rect 16348 1895 16490 1959
rect 16554 1895 16570 1959
rect 16634 1895 16650 1959
rect 16714 1895 16730 1959
rect 16794 1895 16810 1959
rect 16874 1895 16890 1959
rect 16954 1895 17096 1959
rect 17160 1895 17176 1959
rect 17240 1895 17256 1959
rect 17320 1895 17336 1959
rect 17400 1895 17416 1959
rect 17480 1895 17496 1959
rect 17560 1895 17702 1959
rect 17766 1895 17782 1959
rect 17846 1895 17862 1959
rect 17926 1895 17942 1959
rect 18006 1895 18022 1959
rect 18086 1895 18102 1959
rect 18166 1895 18308 1959
rect 18372 1895 18388 1959
rect 18452 1895 18468 1959
rect 18532 1895 18548 1959
rect 18612 1895 18628 1959
rect 18692 1895 18708 1959
rect 18772 1895 18914 1959
rect 18978 1895 18994 1959
rect 19058 1895 19074 1959
rect 19138 1895 19154 1959
rect 19218 1895 19234 1959
rect 19298 1895 19314 1959
rect 19378 1895 19520 1959
rect 19584 1895 19600 1959
rect 19664 1895 19680 1959
rect 19744 1895 19760 1959
rect 19824 1895 19840 1959
rect 19904 1895 19920 1959
rect 19984 1895 20088 1959
rect 10605 1893 20088 1895
rect 20148 1959 39298 1961
rect 20148 1895 20252 1959
rect 20316 1895 20332 1959
rect 20396 1895 20412 1959
rect 20476 1895 20492 1959
rect 20556 1895 20572 1959
rect 20636 1895 20652 1959
rect 20716 1895 20858 1959
rect 20922 1895 20938 1959
rect 21002 1895 21018 1959
rect 21082 1895 21098 1959
rect 21162 1895 21178 1959
rect 21242 1895 21258 1959
rect 21322 1895 21464 1959
rect 21528 1895 21544 1959
rect 21608 1895 21624 1959
rect 21688 1895 21704 1959
rect 21768 1895 21784 1959
rect 21848 1895 21864 1959
rect 21928 1895 22070 1959
rect 22134 1895 22150 1959
rect 22214 1895 22230 1959
rect 22294 1895 22310 1959
rect 22374 1895 22390 1959
rect 22454 1895 22470 1959
rect 22534 1895 22676 1959
rect 22740 1895 22756 1959
rect 22820 1895 22836 1959
rect 22900 1895 22916 1959
rect 22980 1895 22996 1959
rect 23060 1895 23076 1959
rect 23140 1895 23282 1959
rect 23346 1895 23362 1959
rect 23426 1895 23442 1959
rect 23506 1895 23522 1959
rect 23586 1895 23602 1959
rect 23666 1895 23682 1959
rect 23746 1895 23888 1959
rect 23952 1895 23968 1959
rect 24032 1895 24048 1959
rect 24112 1895 24128 1959
rect 24192 1895 24208 1959
rect 24272 1895 24288 1959
rect 24352 1895 24494 1959
rect 24558 1895 24574 1959
rect 24638 1895 24654 1959
rect 24718 1895 24734 1959
rect 24798 1895 24814 1959
rect 24878 1895 24894 1959
rect 24958 1895 25100 1959
rect 25164 1895 25180 1959
rect 25244 1895 25260 1959
rect 25324 1895 25340 1959
rect 25404 1895 25420 1959
rect 25484 1895 25500 1959
rect 25564 1895 25706 1959
rect 25770 1895 25786 1959
rect 25850 1895 25866 1959
rect 25930 1895 25946 1959
rect 26010 1895 26026 1959
rect 26090 1895 26106 1959
rect 26170 1895 26312 1959
rect 26376 1895 26392 1959
rect 26456 1895 26472 1959
rect 26536 1895 26552 1959
rect 26616 1895 26632 1959
rect 26696 1895 26712 1959
rect 26776 1895 26918 1959
rect 26982 1895 26998 1959
rect 27062 1895 27078 1959
rect 27142 1895 27158 1959
rect 27222 1895 27238 1959
rect 27302 1895 27318 1959
rect 27382 1895 27524 1959
rect 27588 1895 27604 1959
rect 27668 1895 27684 1959
rect 27748 1895 27764 1959
rect 27828 1895 27844 1959
rect 27908 1895 27924 1959
rect 27988 1895 28130 1959
rect 28194 1895 28210 1959
rect 28274 1895 28290 1959
rect 28354 1895 28370 1959
rect 28434 1895 28450 1959
rect 28514 1895 28530 1959
rect 28594 1895 28736 1959
rect 28800 1895 28816 1959
rect 28880 1895 28896 1959
rect 28960 1895 28976 1959
rect 29040 1895 29056 1959
rect 29120 1895 29136 1959
rect 29200 1895 29342 1959
rect 29406 1895 29422 1959
rect 29486 1895 29502 1959
rect 29566 1895 29582 1959
rect 29646 1895 29662 1959
rect 29726 1895 29742 1959
rect 29806 1895 29948 1959
rect 30012 1895 30028 1959
rect 30092 1895 30108 1959
rect 30172 1895 30188 1959
rect 30252 1895 30268 1959
rect 30332 1895 30348 1959
rect 30412 1895 30554 1959
rect 30618 1895 30634 1959
rect 30698 1895 30714 1959
rect 30778 1895 30794 1959
rect 30858 1895 30874 1959
rect 30938 1895 30954 1959
rect 31018 1895 31160 1959
rect 31224 1895 31240 1959
rect 31304 1895 31320 1959
rect 31384 1895 31400 1959
rect 31464 1895 31480 1959
rect 31544 1895 31560 1959
rect 31624 1895 31766 1959
rect 31830 1895 31846 1959
rect 31910 1895 31926 1959
rect 31990 1895 32006 1959
rect 32070 1895 32086 1959
rect 32150 1895 32166 1959
rect 32230 1895 32372 1959
rect 32436 1895 32452 1959
rect 32516 1895 32532 1959
rect 32596 1895 32612 1959
rect 32676 1895 32692 1959
rect 32756 1895 32772 1959
rect 32836 1895 32978 1959
rect 33042 1895 33058 1959
rect 33122 1895 33138 1959
rect 33202 1895 33218 1959
rect 33282 1895 33298 1959
rect 33362 1895 33378 1959
rect 33442 1895 33584 1959
rect 33648 1895 33664 1959
rect 33728 1895 33744 1959
rect 33808 1895 33824 1959
rect 33888 1895 33904 1959
rect 33968 1895 33984 1959
rect 34048 1895 34190 1959
rect 34254 1895 34270 1959
rect 34334 1895 34350 1959
rect 34414 1895 34430 1959
rect 34494 1895 34510 1959
rect 34574 1895 34590 1959
rect 34654 1895 34796 1959
rect 34860 1895 34876 1959
rect 34940 1895 34956 1959
rect 35020 1895 35036 1959
rect 35100 1895 35116 1959
rect 35180 1895 35196 1959
rect 35260 1895 35402 1959
rect 35466 1895 35482 1959
rect 35546 1895 35562 1959
rect 35626 1895 35642 1959
rect 35706 1895 35722 1959
rect 35786 1895 35802 1959
rect 35866 1895 36008 1959
rect 36072 1895 36088 1959
rect 36152 1895 36168 1959
rect 36232 1895 36248 1959
rect 36312 1895 36328 1959
rect 36392 1895 36408 1959
rect 36472 1895 36614 1959
rect 36678 1895 36694 1959
rect 36758 1895 36774 1959
rect 36838 1895 36854 1959
rect 36918 1895 36934 1959
rect 36998 1895 37014 1959
rect 37078 1895 37220 1959
rect 37284 1895 37300 1959
rect 37364 1895 37380 1959
rect 37444 1895 37460 1959
rect 37524 1895 37540 1959
rect 37604 1895 37620 1959
rect 37684 1895 37826 1959
rect 37890 1895 37906 1959
rect 37970 1895 37986 1959
rect 38050 1895 38066 1959
rect 38130 1895 38146 1959
rect 38210 1895 38226 1959
rect 38290 1895 38432 1959
rect 38496 1895 38512 1959
rect 38576 1895 38592 1959
rect 38656 1895 38672 1959
rect 38736 1895 38752 1959
rect 38816 1895 38832 1959
rect 38896 1895 39038 1959
rect 39102 1895 39118 1959
rect 39182 1895 39198 1959
rect 39262 1895 39278 1959
rect 20148 1893 39298 1895
rect 39534 1893 39606 1961
rect -459 1739 -393 1893
rect -459 1675 -458 1739
rect -394 1675 -393 1739
rect -459 1659 -393 1675
rect -459 1595 -458 1659
rect -394 1595 -393 1659
rect -459 1579 -393 1595
rect -459 1515 -458 1579
rect -394 1515 -393 1579
rect -459 1499 -393 1515
rect -459 1435 -458 1499
rect -394 1435 -393 1499
rect -459 1419 -393 1435
rect -459 1355 -458 1419
rect -394 1355 -393 1419
rect -459 1339 -393 1355
rect -459 1275 -458 1339
rect -394 1275 -393 1339
rect -459 1259 -393 1275
rect -459 1195 -458 1259
rect -394 1195 -393 1259
rect -459 1179 -393 1195
rect -459 1115 -458 1179
rect -394 1115 -393 1179
rect -459 1099 -393 1115
rect -459 1035 -458 1099
rect -394 1035 -393 1099
rect -459 1019 -393 1035
rect -459 955 -458 1019
rect -394 955 -393 1019
rect -459 865 -393 955
rect -333 861 -273 1893
rect -213 801 -153 1831
rect -93 861 -33 1893
rect 27 801 87 1831
rect 147 1739 213 1893
rect 147 1675 148 1739
rect 212 1675 213 1739
rect 147 1659 213 1675
rect 147 1595 148 1659
rect 212 1595 213 1659
rect 147 1579 213 1595
rect 147 1515 148 1579
rect 212 1515 213 1579
rect 147 1499 213 1515
rect 147 1435 148 1499
rect 212 1435 213 1499
rect 147 1419 213 1435
rect 147 1355 148 1419
rect 212 1355 213 1419
rect 147 1339 213 1355
rect 147 1275 148 1339
rect 212 1275 213 1339
rect 147 1259 213 1275
rect 147 1195 148 1259
rect 212 1195 213 1259
rect 147 1179 213 1195
rect 147 1115 148 1179
rect 212 1115 213 1179
rect 147 1099 213 1115
rect 147 1035 148 1099
rect 212 1035 213 1099
rect 147 1019 213 1035
rect 147 955 148 1019
rect 212 955 213 1019
rect 147 865 213 955
rect 355 1739 421 1829
rect 355 1675 356 1739
rect 420 1675 421 1739
rect 355 1659 421 1675
rect 355 1595 356 1659
rect 420 1595 421 1659
rect 355 1579 421 1595
rect 355 1515 356 1579
rect 420 1515 421 1579
rect 355 1499 421 1515
rect 355 1435 356 1499
rect 420 1435 421 1499
rect 355 1419 421 1435
rect 355 1355 356 1419
rect 420 1355 421 1419
rect 355 1339 421 1355
rect 355 1275 356 1339
rect 420 1275 421 1339
rect 355 1259 421 1275
rect 355 1195 356 1259
rect 420 1195 421 1259
rect 355 1179 421 1195
rect 355 1115 356 1179
rect 420 1115 421 1179
rect 355 1099 421 1115
rect 355 1035 356 1099
rect 420 1035 421 1099
rect 355 1019 421 1035
rect 355 955 356 1019
rect 420 955 421 1019
rect 355 801 421 955
rect 481 863 541 1893
rect 601 801 661 1833
rect 721 863 781 1893
rect 841 801 901 1833
rect 964 1829 1024 1830
rect 961 1821 1027 1829
rect 961 1757 962 1821
rect 1026 1757 1027 1821
rect 961 1739 1027 1757
rect 961 1675 962 1739
rect 1026 1675 1027 1739
rect 961 1659 1027 1675
rect 961 1595 962 1659
rect 1026 1595 1027 1659
rect 961 1579 1027 1595
rect 961 1515 962 1579
rect 1026 1515 1027 1579
rect 961 1499 1027 1515
rect 961 1435 962 1499
rect 1026 1435 1027 1499
rect 961 1419 1027 1435
rect 961 1355 962 1419
rect 1026 1355 1027 1419
rect 961 1339 1027 1355
rect 961 1275 962 1339
rect 1026 1275 1027 1339
rect 961 1259 1027 1275
rect 961 1195 962 1259
rect 1026 1195 1027 1259
rect 961 1179 1027 1195
rect 961 1115 962 1179
rect 1026 1115 1027 1179
rect 961 1099 1027 1115
rect 961 1035 962 1099
rect 1026 1035 1027 1099
rect 961 1019 1027 1035
rect 961 955 962 1019
rect 1026 955 1027 1019
rect 961 801 1027 955
rect -459 799 213 801
rect -459 735 -355 799
rect -291 735 -275 799
rect -211 735 -195 799
rect -131 735 -115 799
rect -51 735 -35 799
rect 29 735 45 799
rect 109 735 213 799
rect -459 733 213 735
rect 355 799 1027 801
rect 355 735 459 799
rect 523 735 539 799
rect 603 735 619 799
rect 683 735 699 799
rect 763 735 779 799
rect 843 735 859 799
rect 923 735 1027 799
rect 355 733 1027 735
rect -459 579 -393 669
rect -459 515 -458 579
rect -394 515 -393 579
rect -459 499 -393 515
rect -459 435 -458 499
rect -394 435 -393 499
rect -459 419 -393 435
rect -459 355 -458 419
rect -394 355 -393 419
rect -459 339 -393 355
rect -459 275 -458 339
rect -394 275 -393 339
rect -459 259 -393 275
rect -459 195 -458 259
rect -394 195 -393 259
rect -459 179 -393 195
rect -459 115 -458 179
rect -394 115 -393 179
rect -459 99 -393 115
rect -459 35 -458 99
rect -394 35 -393 99
rect -459 19 -393 35
rect -459 -45 -458 19
rect -394 -45 -393 19
rect -459 -61 -393 -45
rect -459 -125 -458 -61
rect -394 -125 -393 -61
rect -459 -141 -393 -125
rect -459 -205 -458 -141
rect -394 -205 -393 -141
rect -459 -359 -393 -205
rect -333 -297 -273 733
rect -213 -359 -153 673
rect -93 -297 -33 733
rect 27 -359 87 673
rect 147 579 213 669
rect 147 515 148 579
rect 212 515 213 579
rect 147 499 213 515
rect 147 435 148 499
rect 212 435 213 499
rect 147 419 213 435
rect 147 355 148 419
rect 212 355 213 419
rect 147 339 213 355
rect 147 275 148 339
rect 212 275 213 339
rect 147 259 213 275
rect 147 195 148 259
rect 212 195 213 259
rect 147 179 213 195
rect 147 115 148 179
rect 212 115 213 179
rect 147 99 213 115
rect 147 35 148 99
rect 212 35 213 99
rect 147 19 213 35
rect 147 -45 148 19
rect 212 -45 213 19
rect 147 -61 213 -45
rect 147 -125 148 -61
rect 212 -125 213 -61
rect 147 -141 213 -125
rect 147 -205 148 -141
rect 212 -205 213 -141
rect 147 -359 213 -205
rect 355 579 421 733
rect 355 515 356 579
rect 420 515 421 579
rect 355 499 421 515
rect 355 435 356 499
rect 420 435 421 499
rect 355 419 421 435
rect 355 355 356 419
rect 420 355 421 419
rect 355 339 421 355
rect 355 275 356 339
rect 420 275 421 339
rect 355 259 421 275
rect 355 195 356 259
rect 420 195 421 259
rect 355 179 421 195
rect 355 115 356 179
rect 420 115 421 179
rect 355 99 421 115
rect 355 35 356 99
rect 420 35 421 99
rect 355 19 421 35
rect 355 -45 356 19
rect 420 -45 421 19
rect 355 -61 421 -45
rect 355 -125 356 -61
rect 420 -125 421 -61
rect 355 -141 421 -125
rect 355 -205 356 -141
rect 420 -205 421 -141
rect 355 -295 421 -205
rect 481 -299 541 733
rect 601 -359 661 671
rect 721 -299 781 733
rect 841 -359 901 671
rect 961 579 1027 733
rect 961 515 962 579
rect 1026 515 1027 579
rect 961 499 1027 515
rect 961 435 962 499
rect 1026 435 1027 499
rect 961 419 1027 435
rect 961 355 962 419
rect 1026 355 1027 419
rect 961 339 1027 355
rect 961 275 962 339
rect 1026 275 1027 339
rect 961 259 1027 275
rect 961 195 962 259
rect 1026 195 1027 259
rect 961 179 1027 195
rect 961 115 962 179
rect 1026 115 1027 179
rect 961 99 1027 115
rect 961 35 962 99
rect 1026 35 1027 99
rect 961 19 1027 35
rect 961 -45 962 19
rect 1026 -45 1027 19
rect 961 -61 1027 -45
rect 961 -125 962 -61
rect 1026 -125 1027 -61
rect 961 -141 1027 -125
rect 961 -205 962 -141
rect 1026 -205 1027 -141
rect 961 -295 1027 -205
rect 1267 1739 1333 1829
rect 1267 1675 1268 1739
rect 1332 1675 1333 1739
rect 1267 1659 1333 1675
rect 1267 1595 1268 1659
rect 1332 1595 1333 1659
rect 1267 1579 1333 1595
rect 1267 1515 1268 1579
rect 1332 1515 1333 1579
rect 1267 1499 1333 1515
rect 1267 1435 1268 1499
rect 1332 1435 1333 1499
rect 1267 1419 1333 1435
rect 1267 1355 1268 1419
rect 1332 1355 1333 1419
rect 1267 1339 1333 1355
rect 1267 1275 1268 1339
rect 1332 1275 1333 1339
rect 1267 1259 1333 1275
rect 1267 1195 1268 1259
rect 1332 1195 1333 1259
rect 1267 1179 1333 1195
rect 1267 1115 1268 1179
rect 1332 1115 1333 1179
rect 1267 1099 1333 1115
rect 1267 1035 1268 1099
rect 1332 1035 1333 1099
rect 1267 1019 1333 1035
rect 1267 955 1268 1019
rect 1332 955 1333 1019
rect 1267 801 1333 955
rect 1393 863 1453 1893
rect 1513 801 1573 1833
rect 1633 863 1693 1893
rect 1753 801 1813 1833
rect 1873 1820 1939 1829
rect 1873 1756 1874 1820
rect 1938 1756 1939 1820
rect 1873 1739 1939 1756
rect 1873 1675 1874 1739
rect 1938 1675 1939 1739
rect 1873 1659 1939 1675
rect 1873 1595 1874 1659
rect 1938 1595 1939 1659
rect 1873 1579 1939 1595
rect 1873 1515 1874 1579
rect 1938 1515 1939 1579
rect 1873 1499 1939 1515
rect 1873 1435 1874 1499
rect 1938 1435 1939 1499
rect 1873 1419 1939 1435
rect 1873 1355 1874 1419
rect 1938 1355 1939 1419
rect 1873 1339 1939 1355
rect 1873 1275 1874 1339
rect 1938 1275 1939 1339
rect 1873 1259 1939 1275
rect 1873 1195 1874 1259
rect 1938 1195 1939 1259
rect 1873 1179 1939 1195
rect 1873 1115 1874 1179
rect 1938 1115 1939 1179
rect 1873 1099 1939 1115
rect 1873 1035 1874 1099
rect 1938 1035 1939 1099
rect 1873 1019 1939 1035
rect 1873 955 1874 1019
rect 1938 955 1939 1019
rect 1873 801 1939 955
rect 1999 863 2059 1893
rect 2119 801 2179 1833
rect 2239 863 2299 1893
rect 2359 801 2419 1833
rect 2479 1821 2545 1830
rect 2479 1757 2480 1821
rect 2544 1757 2545 1821
rect 2479 1739 2545 1757
rect 2479 1675 2480 1739
rect 2544 1675 2545 1739
rect 2479 1659 2545 1675
rect 2479 1595 2480 1659
rect 2544 1595 2545 1659
rect 2479 1579 2545 1595
rect 2479 1515 2480 1579
rect 2544 1515 2545 1579
rect 2479 1499 2545 1515
rect 2479 1435 2480 1499
rect 2544 1435 2545 1499
rect 2479 1419 2545 1435
rect 2479 1355 2480 1419
rect 2544 1355 2545 1419
rect 2479 1339 2545 1355
rect 2479 1275 2480 1339
rect 2544 1275 2545 1339
rect 2479 1259 2545 1275
rect 2479 1195 2480 1259
rect 2544 1195 2545 1259
rect 2479 1179 2545 1195
rect 2479 1115 2480 1179
rect 2544 1115 2545 1179
rect 2479 1099 2545 1115
rect 2479 1035 2480 1099
rect 2544 1035 2545 1099
rect 2479 1019 2545 1035
rect 2479 955 2480 1019
rect 2544 955 2545 1019
rect 2479 801 2545 955
rect 1267 799 2545 801
rect 1267 735 1371 799
rect 1435 735 1451 799
rect 1515 735 1531 799
rect 1595 735 1611 799
rect 1675 735 1691 799
rect 1755 735 1771 799
rect 1835 735 1977 799
rect 2041 735 2057 799
rect 2121 735 2137 799
rect 2201 735 2217 799
rect 2281 735 2297 799
rect 2361 735 2377 799
rect 2441 735 2545 799
rect 1267 733 2545 735
rect 1267 579 1333 733
rect 1267 515 1268 579
rect 1332 515 1333 579
rect 1267 499 1333 515
rect 1267 435 1268 499
rect 1332 435 1333 499
rect 1267 419 1333 435
rect 1267 355 1268 419
rect 1332 355 1333 419
rect 1267 339 1333 355
rect 1267 275 1268 339
rect 1332 275 1333 339
rect 1267 259 1333 275
rect 1267 195 1268 259
rect 1332 195 1333 259
rect 1267 179 1333 195
rect 1267 115 1268 179
rect 1332 115 1333 179
rect 1267 99 1333 115
rect 1267 35 1268 99
rect 1332 35 1333 99
rect 1267 19 1333 35
rect 1267 -45 1268 19
rect 1332 -45 1333 19
rect 1267 -61 1333 -45
rect 1267 -125 1268 -61
rect 1332 -125 1333 -61
rect 1267 -141 1333 -125
rect 1267 -205 1268 -141
rect 1332 -205 1333 -141
rect 1267 -295 1333 -205
rect 1393 -299 1453 733
rect 1513 -359 1573 671
rect 1633 -299 1693 733
rect 1753 -359 1813 671
rect 1873 579 1939 733
rect 1873 515 1874 579
rect 1938 515 1939 579
rect 1873 499 1939 515
rect 1873 435 1874 499
rect 1938 435 1939 499
rect 1873 419 1939 435
rect 1873 355 1874 419
rect 1938 355 1939 419
rect 1873 339 1939 355
rect 1873 275 1874 339
rect 1938 275 1939 339
rect 1873 259 1939 275
rect 1873 195 1874 259
rect 1938 195 1939 259
rect 1873 179 1939 195
rect 1873 115 1874 179
rect 1938 115 1939 179
rect 1873 99 1939 115
rect 1873 35 1874 99
rect 1938 35 1939 99
rect 1873 19 1939 35
rect 1873 -45 1874 19
rect 1938 -45 1939 19
rect 1873 -61 1939 -45
rect 1873 -125 1874 -61
rect 1938 -125 1939 -61
rect 1873 -141 1939 -125
rect 1873 -205 1874 -141
rect 1938 -205 1939 -141
rect 1873 -295 1939 -205
rect 1999 -299 2059 733
rect 2119 -359 2179 671
rect 2239 -299 2299 733
rect 2359 -359 2419 671
rect 2479 579 2545 733
rect 2479 515 2480 579
rect 2544 515 2545 579
rect 2479 499 2545 515
rect 2479 435 2480 499
rect 2544 435 2545 499
rect 2479 419 2545 435
rect 2479 355 2480 419
rect 2544 355 2545 419
rect 2479 339 2545 355
rect 2479 275 2480 339
rect 2544 275 2545 339
rect 2479 259 2545 275
rect 2479 195 2480 259
rect 2544 195 2545 259
rect 2479 179 2545 195
rect 2479 115 2480 179
rect 2544 115 2545 179
rect 2479 99 2545 115
rect 2479 35 2480 99
rect 2544 35 2545 99
rect 2479 19 2545 35
rect 2479 -45 2480 19
rect 2544 -45 2545 19
rect 2479 -61 2545 -45
rect 2479 -125 2480 -61
rect 2544 -125 2545 -61
rect 2479 -141 2545 -125
rect 2479 -205 2480 -141
rect 2544 -205 2545 -141
rect 2479 -295 2545 -205
rect 2801 1739 2867 1829
rect 2801 1675 2802 1739
rect 2866 1675 2867 1739
rect 2801 1659 2867 1675
rect 2801 1595 2802 1659
rect 2866 1595 2867 1659
rect 2801 1579 2867 1595
rect 2801 1515 2802 1579
rect 2866 1515 2867 1579
rect 2801 1499 2867 1515
rect 2801 1435 2802 1499
rect 2866 1435 2867 1499
rect 2801 1419 2867 1435
rect 2801 1355 2802 1419
rect 2866 1355 2867 1419
rect 2801 1339 2867 1355
rect 2801 1275 2802 1339
rect 2866 1275 2867 1339
rect 2801 1259 2867 1275
rect 2801 1195 2802 1259
rect 2866 1195 2867 1259
rect 2801 1179 2867 1195
rect 2801 1115 2802 1179
rect 2866 1115 2867 1179
rect 2801 1099 2867 1115
rect 2801 1035 2802 1099
rect 2866 1035 2867 1099
rect 2801 1019 2867 1035
rect 2801 955 2802 1019
rect 2866 955 2867 1019
rect 2801 801 2867 955
rect 2927 863 2987 1893
rect 3047 801 3107 1833
rect 3167 863 3227 1893
rect 3287 801 3347 1833
rect 3407 1739 3473 1829
rect 3407 1675 3408 1739
rect 3472 1675 3473 1739
rect 3407 1659 3473 1675
rect 3407 1595 3408 1659
rect 3472 1595 3473 1659
rect 3407 1579 3473 1595
rect 3407 1515 3408 1579
rect 3472 1515 3473 1579
rect 3407 1499 3473 1515
rect 3407 1435 3408 1499
rect 3472 1435 3473 1499
rect 3407 1419 3473 1435
rect 3407 1355 3408 1419
rect 3472 1355 3473 1419
rect 3407 1339 3473 1355
rect 3407 1275 3408 1339
rect 3472 1275 3473 1339
rect 3407 1259 3473 1275
rect 3407 1195 3408 1259
rect 3472 1195 3473 1259
rect 3407 1179 3473 1195
rect 3407 1115 3408 1179
rect 3472 1115 3473 1179
rect 3407 1099 3473 1115
rect 3407 1035 3408 1099
rect 3472 1035 3473 1099
rect 3407 1019 3473 1035
rect 3407 955 3408 1019
rect 3472 955 3473 1019
rect 3407 801 3473 955
rect 3533 863 3593 1893
rect 3653 801 3713 1833
rect 3773 863 3833 1893
rect 3893 801 3953 1833
rect 4013 1739 4079 1829
rect 4013 1675 4014 1739
rect 4078 1675 4079 1739
rect 4013 1659 4079 1675
rect 4013 1595 4014 1659
rect 4078 1595 4079 1659
rect 4013 1579 4079 1595
rect 4013 1515 4014 1579
rect 4078 1515 4079 1579
rect 4013 1499 4079 1515
rect 4013 1435 4014 1499
rect 4078 1435 4079 1499
rect 4013 1419 4079 1435
rect 4013 1355 4014 1419
rect 4078 1355 4079 1419
rect 4013 1339 4079 1355
rect 4013 1275 4014 1339
rect 4078 1275 4079 1339
rect 4013 1259 4079 1275
rect 4013 1195 4014 1259
rect 4078 1195 4079 1259
rect 4013 1179 4079 1195
rect 4013 1115 4014 1179
rect 4078 1115 4079 1179
rect 4013 1099 4079 1115
rect 4013 1035 4014 1099
rect 4078 1035 4079 1099
rect 4013 1019 4079 1035
rect 4013 955 4014 1019
rect 4078 955 4079 1019
rect 4013 801 4079 955
rect 4139 863 4199 1893
rect 4259 801 4319 1833
rect 4379 863 4439 1893
rect 4499 801 4559 1833
rect 4619 1739 4685 1829
rect 4619 1675 4620 1739
rect 4684 1675 4685 1739
rect 4619 1659 4685 1675
rect 4619 1595 4620 1659
rect 4684 1595 4685 1659
rect 4619 1579 4685 1595
rect 4619 1515 4620 1579
rect 4684 1515 4685 1579
rect 4619 1499 4685 1515
rect 4619 1435 4620 1499
rect 4684 1435 4685 1499
rect 4619 1419 4685 1435
rect 4619 1355 4620 1419
rect 4684 1355 4685 1419
rect 4619 1339 4685 1355
rect 4619 1275 4620 1339
rect 4684 1275 4685 1339
rect 4619 1259 4685 1275
rect 4619 1195 4620 1259
rect 4684 1195 4685 1259
rect 4619 1179 4685 1195
rect 4619 1115 4620 1179
rect 4684 1115 4685 1179
rect 4619 1099 4685 1115
rect 4619 1035 4620 1099
rect 4684 1035 4685 1099
rect 4619 1019 4685 1035
rect 4619 955 4620 1019
rect 4684 955 4685 1019
rect 4619 801 4685 955
rect 4745 863 4805 1893
rect 4865 801 4925 1833
rect 4985 863 5045 1893
rect 5105 801 5165 1833
rect 5225 1739 5291 1829
rect 5225 1675 5226 1739
rect 5290 1675 5291 1739
rect 5225 1659 5291 1675
rect 5225 1595 5226 1659
rect 5290 1595 5291 1659
rect 5225 1579 5291 1595
rect 5225 1515 5226 1579
rect 5290 1515 5291 1579
rect 5225 1499 5291 1515
rect 5225 1435 5226 1499
rect 5290 1435 5291 1499
rect 5225 1419 5291 1435
rect 5225 1355 5226 1419
rect 5290 1355 5291 1419
rect 5225 1339 5291 1355
rect 5225 1275 5226 1339
rect 5290 1275 5291 1339
rect 5225 1259 5291 1275
rect 5225 1195 5226 1259
rect 5290 1195 5291 1259
rect 5225 1179 5291 1195
rect 5225 1115 5226 1179
rect 5290 1115 5291 1179
rect 5225 1099 5291 1115
rect 5225 1035 5226 1099
rect 5290 1035 5291 1099
rect 5225 1019 5291 1035
rect 5225 955 5226 1019
rect 5290 955 5291 1019
rect 5225 801 5291 955
rect 2801 799 5291 801
rect 2801 735 2905 799
rect 2969 735 2985 799
rect 3049 735 3065 799
rect 3129 735 3145 799
rect 3209 735 3225 799
rect 3289 735 3305 799
rect 3369 735 3511 799
rect 3575 735 3591 799
rect 3655 735 3671 799
rect 3735 735 3751 799
rect 3815 735 3831 799
rect 3895 735 3911 799
rect 3975 735 4117 799
rect 4181 735 4197 799
rect 4261 735 4277 799
rect 4341 735 4357 799
rect 4421 735 4437 799
rect 4501 735 4517 799
rect 4581 735 4723 799
rect 4787 735 4803 799
rect 4867 735 4883 799
rect 4947 735 4963 799
rect 5027 735 5043 799
rect 5107 735 5123 799
rect 5187 735 5291 799
rect 2801 733 5291 735
rect 2801 579 2867 733
rect 2801 515 2802 579
rect 2866 515 2867 579
rect 2801 499 2867 515
rect 2801 435 2802 499
rect 2866 435 2867 499
rect 2801 419 2867 435
rect 2801 355 2802 419
rect 2866 355 2867 419
rect 2801 339 2867 355
rect 2801 275 2802 339
rect 2866 275 2867 339
rect 2801 259 2867 275
rect 2801 195 2802 259
rect 2866 195 2867 259
rect 2801 179 2867 195
rect 2801 115 2802 179
rect 2866 115 2867 179
rect 2801 99 2867 115
rect 2801 35 2802 99
rect 2866 35 2867 99
rect 2801 19 2867 35
rect 2801 -45 2802 19
rect 2866 -45 2867 19
rect 2801 -61 2867 -45
rect 2801 -125 2802 -61
rect 2866 -125 2867 -61
rect 2801 -141 2867 -125
rect 2801 -205 2802 -141
rect 2866 -205 2867 -141
rect 2801 -295 2867 -205
rect 2927 -299 2987 733
rect 3047 -359 3107 671
rect 3167 -299 3227 733
rect 3287 -359 3347 671
rect 3407 579 3473 733
rect 3407 515 3408 579
rect 3472 515 3473 579
rect 3407 499 3473 515
rect 3407 435 3408 499
rect 3472 435 3473 499
rect 3407 419 3473 435
rect 3407 355 3408 419
rect 3472 355 3473 419
rect 3407 339 3473 355
rect 3407 275 3408 339
rect 3472 275 3473 339
rect 3407 259 3473 275
rect 3407 195 3408 259
rect 3472 195 3473 259
rect 3407 179 3473 195
rect 3407 115 3408 179
rect 3472 115 3473 179
rect 3407 99 3473 115
rect 3407 35 3408 99
rect 3472 35 3473 99
rect 3407 19 3473 35
rect 3407 -45 3408 19
rect 3472 -45 3473 19
rect 3407 -61 3473 -45
rect 3407 -125 3408 -61
rect 3472 -125 3473 -61
rect 3407 -141 3473 -125
rect 3407 -205 3408 -141
rect 3472 -205 3473 -141
rect 3407 -295 3473 -205
rect 3533 -299 3593 733
rect 3653 -359 3713 671
rect 3773 -299 3833 733
rect 3893 -359 3953 671
rect 4013 579 4079 733
rect 4013 515 4014 579
rect 4078 515 4079 579
rect 4013 499 4079 515
rect 4013 435 4014 499
rect 4078 435 4079 499
rect 4013 419 4079 435
rect 4013 355 4014 419
rect 4078 355 4079 419
rect 4013 339 4079 355
rect 4013 275 4014 339
rect 4078 275 4079 339
rect 4013 259 4079 275
rect 4013 195 4014 259
rect 4078 195 4079 259
rect 4013 179 4079 195
rect 4013 115 4014 179
rect 4078 115 4079 179
rect 4013 99 4079 115
rect 4013 35 4014 99
rect 4078 35 4079 99
rect 4013 19 4079 35
rect 4013 -45 4014 19
rect 4078 -45 4079 19
rect 4013 -61 4079 -45
rect 4013 -125 4014 -61
rect 4078 -125 4079 -61
rect 4013 -141 4079 -125
rect 4013 -205 4014 -141
rect 4078 -205 4079 -141
rect 4013 -295 4079 -205
rect 4139 -299 4199 733
rect 4259 -359 4319 671
rect 4379 -299 4439 733
rect 4499 -359 4559 671
rect 4619 579 4685 733
rect 4619 515 4620 579
rect 4684 515 4685 579
rect 4619 499 4685 515
rect 4619 435 4620 499
rect 4684 435 4685 499
rect 4619 419 4685 435
rect 4619 355 4620 419
rect 4684 355 4685 419
rect 4619 339 4685 355
rect 4619 275 4620 339
rect 4684 275 4685 339
rect 4619 259 4685 275
rect 4619 195 4620 259
rect 4684 195 4685 259
rect 4619 179 4685 195
rect 4619 115 4620 179
rect 4684 115 4685 179
rect 4619 99 4685 115
rect 4619 35 4620 99
rect 4684 35 4685 99
rect 4619 19 4685 35
rect 4619 -45 4620 19
rect 4684 -45 4685 19
rect 4619 -61 4685 -45
rect 4619 -125 4620 -61
rect 4684 -125 4685 -61
rect 4619 -141 4685 -125
rect 4619 -205 4620 -141
rect 4684 -205 4685 -141
rect 4619 -295 4685 -205
rect 4745 -299 4805 733
rect 4865 -359 4925 671
rect 4985 -299 5045 733
rect 5105 -359 5165 671
rect 5225 579 5291 733
rect 5225 515 5226 579
rect 5290 515 5291 579
rect 5225 499 5291 515
rect 5225 435 5226 499
rect 5290 435 5291 499
rect 5225 419 5291 435
rect 5225 355 5226 419
rect 5290 355 5291 419
rect 5225 339 5291 355
rect 5225 275 5226 339
rect 5290 275 5291 339
rect 5225 259 5291 275
rect 5225 195 5226 259
rect 5290 195 5291 259
rect 5225 179 5291 195
rect 5225 115 5226 179
rect 5290 115 5291 179
rect 5225 99 5291 115
rect 5225 35 5226 99
rect 5290 35 5291 99
rect 5225 19 5291 35
rect 5225 -45 5226 19
rect 5290 -45 5291 19
rect 5225 -61 5291 -45
rect 5225 -125 5226 -61
rect 5290 -125 5291 -61
rect 5225 -141 5291 -125
rect 5225 -205 5226 -141
rect 5290 -205 5291 -141
rect 5225 -295 5291 -205
rect 5352 1739 5418 1829
rect 5352 1675 5353 1739
rect 5417 1675 5418 1739
rect 5352 1659 5418 1675
rect 5352 1595 5353 1659
rect 5417 1595 5418 1659
rect 5352 1579 5418 1595
rect 5352 1515 5353 1579
rect 5417 1515 5418 1579
rect 5352 1499 5418 1515
rect 5352 1435 5353 1499
rect 5417 1435 5418 1499
rect 5352 1419 5418 1435
rect 5352 1355 5353 1419
rect 5417 1355 5418 1419
rect 5352 1339 5418 1355
rect 5352 1275 5353 1339
rect 5417 1275 5418 1339
rect 5352 1259 5418 1275
rect 5352 1195 5353 1259
rect 5417 1195 5418 1259
rect 5352 1179 5418 1195
rect 5352 1115 5353 1179
rect 5417 1115 5418 1179
rect 5352 1099 5418 1115
rect 5352 1035 5353 1099
rect 5417 1035 5418 1099
rect 5352 1019 5418 1035
rect 5352 955 5353 1019
rect 5417 955 5418 1019
rect 5352 801 5418 955
rect 5478 863 5538 1893
rect 5598 801 5658 1833
rect 5718 863 5778 1893
rect 5838 801 5898 1833
rect 5958 1739 6024 1829
rect 5958 1675 5959 1739
rect 6023 1675 6024 1739
rect 5958 1659 6024 1675
rect 5958 1595 5959 1659
rect 6023 1595 6024 1659
rect 5958 1579 6024 1595
rect 5958 1515 5959 1579
rect 6023 1515 6024 1579
rect 5958 1499 6024 1515
rect 5958 1435 5959 1499
rect 6023 1435 6024 1499
rect 5958 1419 6024 1435
rect 5958 1355 5959 1419
rect 6023 1355 6024 1419
rect 5958 1339 6024 1355
rect 5958 1275 5959 1339
rect 6023 1275 6024 1339
rect 5958 1259 6024 1275
rect 5958 1195 5959 1259
rect 6023 1195 6024 1259
rect 5958 1179 6024 1195
rect 5958 1115 5959 1179
rect 6023 1115 6024 1179
rect 5958 1099 6024 1115
rect 5958 1035 5959 1099
rect 6023 1035 6024 1099
rect 5958 1019 6024 1035
rect 5958 955 5959 1019
rect 6023 955 6024 1019
rect 5958 801 6024 955
rect 6084 863 6144 1893
rect 6204 801 6264 1833
rect 6324 863 6384 1893
rect 6444 801 6504 1833
rect 6564 1739 6630 1829
rect 6564 1675 6565 1739
rect 6629 1675 6630 1739
rect 6564 1659 6630 1675
rect 6564 1595 6565 1659
rect 6629 1595 6630 1659
rect 6564 1579 6630 1595
rect 6564 1515 6565 1579
rect 6629 1515 6630 1579
rect 6564 1499 6630 1515
rect 6564 1435 6565 1499
rect 6629 1435 6630 1499
rect 6564 1419 6630 1435
rect 6564 1355 6565 1419
rect 6629 1355 6630 1419
rect 6564 1339 6630 1355
rect 6564 1275 6565 1339
rect 6629 1275 6630 1339
rect 6564 1259 6630 1275
rect 6564 1195 6565 1259
rect 6629 1195 6630 1259
rect 6564 1179 6630 1195
rect 6564 1115 6565 1179
rect 6629 1115 6630 1179
rect 6564 1099 6630 1115
rect 6564 1035 6565 1099
rect 6629 1035 6630 1099
rect 6564 1019 6630 1035
rect 6564 955 6565 1019
rect 6629 955 6630 1019
rect 6564 801 6630 955
rect 6690 863 6750 1893
rect 6810 801 6870 1833
rect 6930 863 6990 1893
rect 7050 801 7110 1833
rect 7170 1739 7236 1829
rect 7170 1675 7171 1739
rect 7235 1675 7236 1739
rect 7170 1659 7236 1675
rect 7170 1595 7171 1659
rect 7235 1595 7236 1659
rect 7170 1579 7236 1595
rect 7170 1515 7171 1579
rect 7235 1515 7236 1579
rect 7170 1499 7236 1515
rect 7170 1435 7171 1499
rect 7235 1435 7236 1499
rect 7170 1419 7236 1435
rect 7170 1355 7171 1419
rect 7235 1355 7236 1419
rect 7170 1339 7236 1355
rect 7170 1275 7171 1339
rect 7235 1275 7236 1339
rect 7170 1259 7236 1275
rect 7170 1195 7171 1259
rect 7235 1195 7236 1259
rect 7170 1179 7236 1195
rect 7170 1115 7171 1179
rect 7235 1115 7236 1179
rect 7170 1099 7236 1115
rect 7170 1035 7171 1099
rect 7235 1035 7236 1099
rect 7170 1019 7236 1035
rect 7170 955 7171 1019
rect 7235 955 7236 1019
rect 7170 801 7236 955
rect 7296 863 7356 1893
rect 7416 801 7476 1833
rect 7536 863 7596 1893
rect 7656 801 7716 1833
rect 7776 1739 7842 1829
rect 7776 1675 7777 1739
rect 7841 1675 7842 1739
rect 7776 1659 7842 1675
rect 7776 1595 7777 1659
rect 7841 1595 7842 1659
rect 7776 1579 7842 1595
rect 7776 1515 7777 1579
rect 7841 1515 7842 1579
rect 7776 1499 7842 1515
rect 7776 1435 7777 1499
rect 7841 1435 7842 1499
rect 7776 1419 7842 1435
rect 7776 1355 7777 1419
rect 7841 1355 7842 1419
rect 7776 1339 7842 1355
rect 7776 1275 7777 1339
rect 7841 1275 7842 1339
rect 7776 1259 7842 1275
rect 7776 1195 7777 1259
rect 7841 1195 7842 1259
rect 7776 1179 7842 1195
rect 7776 1115 7777 1179
rect 7841 1115 7842 1179
rect 7776 1099 7842 1115
rect 7776 1035 7777 1099
rect 7841 1035 7842 1099
rect 7776 1019 7842 1035
rect 7776 955 7777 1019
rect 7841 955 7842 1019
rect 7776 801 7842 955
rect 7902 863 7962 1893
rect 8022 801 8082 1833
rect 8142 863 8202 1893
rect 8262 801 8322 1833
rect 8382 1739 8448 1829
rect 8382 1675 8383 1739
rect 8447 1675 8448 1739
rect 8382 1659 8448 1675
rect 8382 1595 8383 1659
rect 8447 1595 8448 1659
rect 8382 1579 8448 1595
rect 8382 1515 8383 1579
rect 8447 1515 8448 1579
rect 8382 1499 8448 1515
rect 8382 1435 8383 1499
rect 8447 1435 8448 1499
rect 8382 1419 8448 1435
rect 8382 1355 8383 1419
rect 8447 1355 8448 1419
rect 8382 1339 8448 1355
rect 8382 1275 8383 1339
rect 8447 1275 8448 1339
rect 8382 1259 8448 1275
rect 8382 1195 8383 1259
rect 8447 1195 8448 1259
rect 8382 1179 8448 1195
rect 8382 1115 8383 1179
rect 8447 1115 8448 1179
rect 8382 1099 8448 1115
rect 8382 1035 8383 1099
rect 8447 1035 8448 1099
rect 8382 1019 8448 1035
rect 8382 955 8383 1019
rect 8447 955 8448 1019
rect 8382 801 8448 955
rect 8508 863 8568 1893
rect 8628 801 8688 1833
rect 8748 863 8808 1893
rect 8868 801 8928 1833
rect 8988 1739 9054 1829
rect 8988 1675 8989 1739
rect 9053 1675 9054 1739
rect 8988 1659 9054 1675
rect 8988 1595 8989 1659
rect 9053 1595 9054 1659
rect 8988 1579 9054 1595
rect 8988 1515 8989 1579
rect 9053 1515 9054 1579
rect 8988 1499 9054 1515
rect 8988 1435 8989 1499
rect 9053 1435 9054 1499
rect 8988 1419 9054 1435
rect 8988 1355 8989 1419
rect 9053 1355 9054 1419
rect 8988 1339 9054 1355
rect 8988 1275 8989 1339
rect 9053 1275 9054 1339
rect 8988 1259 9054 1275
rect 8988 1195 8989 1259
rect 9053 1195 9054 1259
rect 8988 1179 9054 1195
rect 8988 1115 8989 1179
rect 9053 1115 9054 1179
rect 8988 1099 9054 1115
rect 8988 1035 8989 1099
rect 9053 1035 9054 1099
rect 8988 1019 9054 1035
rect 8988 955 8989 1019
rect 9053 955 9054 1019
rect 8988 801 9054 955
rect 9114 863 9174 1893
rect 9234 801 9294 1833
rect 9354 863 9414 1893
rect 9474 801 9534 1833
rect 9594 1739 9660 1829
rect 9594 1675 9595 1739
rect 9659 1675 9660 1739
rect 9594 1659 9660 1675
rect 9594 1595 9595 1659
rect 9659 1595 9660 1659
rect 9594 1579 9660 1595
rect 9594 1515 9595 1579
rect 9659 1515 9660 1579
rect 9594 1499 9660 1515
rect 9594 1435 9595 1499
rect 9659 1435 9660 1499
rect 9594 1419 9660 1435
rect 9594 1355 9595 1419
rect 9659 1355 9660 1419
rect 9594 1339 9660 1355
rect 9594 1275 9595 1339
rect 9659 1275 9660 1339
rect 9594 1259 9660 1275
rect 9594 1195 9595 1259
rect 9659 1195 9660 1259
rect 9594 1179 9660 1195
rect 9594 1115 9595 1179
rect 9659 1115 9660 1179
rect 9594 1099 9660 1115
rect 9594 1035 9595 1099
rect 9659 1035 9660 1099
rect 9594 1019 9660 1035
rect 9594 955 9595 1019
rect 9659 955 9660 1019
rect 9594 801 9660 955
rect 9720 863 9780 1893
rect 9840 801 9900 1833
rect 9960 863 10020 1893
rect 10080 801 10140 1833
rect 10200 1739 10266 1829
rect 10200 1675 10201 1739
rect 10265 1675 10266 1739
rect 10200 1659 10266 1675
rect 10200 1595 10201 1659
rect 10265 1595 10266 1659
rect 10200 1579 10266 1595
rect 10200 1515 10201 1579
rect 10265 1515 10266 1579
rect 10200 1499 10266 1515
rect 10200 1435 10201 1499
rect 10265 1435 10266 1499
rect 10200 1419 10266 1435
rect 10200 1355 10201 1419
rect 10265 1355 10266 1419
rect 10200 1339 10266 1355
rect 10200 1275 10201 1339
rect 10265 1275 10266 1339
rect 10200 1259 10266 1275
rect 10200 1195 10201 1259
rect 10265 1195 10266 1259
rect 10200 1179 10266 1195
rect 10200 1115 10201 1179
rect 10265 1115 10266 1179
rect 10200 1099 10266 1115
rect 10200 1035 10201 1099
rect 10265 1035 10266 1099
rect 10200 1019 10266 1035
rect 10200 955 10201 1019
rect 10265 955 10266 1019
rect 10200 801 10266 955
rect 5352 799 10266 801
rect 5352 735 5456 799
rect 5520 735 5536 799
rect 5600 735 5616 799
rect 5680 735 5696 799
rect 5760 735 5776 799
rect 5840 735 5856 799
rect 5920 735 6062 799
rect 6126 735 6142 799
rect 6206 735 6222 799
rect 6286 735 6302 799
rect 6366 735 6382 799
rect 6446 735 6462 799
rect 6526 735 6668 799
rect 6732 735 6748 799
rect 6812 735 6828 799
rect 6892 735 6908 799
rect 6972 735 6988 799
rect 7052 735 7068 799
rect 7132 735 7274 799
rect 7338 735 7354 799
rect 7418 735 7434 799
rect 7498 735 7514 799
rect 7578 735 7594 799
rect 7658 735 7674 799
rect 7738 735 7880 799
rect 7944 735 7960 799
rect 8024 735 8040 799
rect 8104 735 8120 799
rect 8184 735 8200 799
rect 8264 735 8280 799
rect 8344 735 8486 799
rect 8550 735 8566 799
rect 8630 735 8646 799
rect 8710 735 8726 799
rect 8790 735 8806 799
rect 8870 735 8886 799
rect 8950 735 9092 799
rect 9156 735 9172 799
rect 9236 735 9252 799
rect 9316 735 9332 799
rect 9396 735 9412 799
rect 9476 735 9492 799
rect 9556 735 9698 799
rect 9762 735 9778 799
rect 9842 735 9858 799
rect 9922 735 9938 799
rect 10002 735 10018 799
rect 10082 735 10098 799
rect 10162 735 10266 799
rect 5352 733 10266 735
rect 5352 579 5418 733
rect 5352 515 5353 579
rect 5417 515 5418 579
rect 5352 499 5418 515
rect 5352 435 5353 499
rect 5417 435 5418 499
rect 5352 419 5418 435
rect 5352 355 5353 419
rect 5417 355 5418 419
rect 5352 339 5418 355
rect 5352 275 5353 339
rect 5417 275 5418 339
rect 5352 259 5418 275
rect 5352 195 5353 259
rect 5417 195 5418 259
rect 5352 179 5418 195
rect 5352 115 5353 179
rect 5417 115 5418 179
rect 5352 99 5418 115
rect 5352 35 5353 99
rect 5417 35 5418 99
rect 5352 19 5418 35
rect 5352 -45 5353 19
rect 5417 -45 5418 19
rect 5352 -61 5418 -45
rect 5352 -125 5353 -61
rect 5417 -125 5418 -61
rect 5352 -141 5418 -125
rect 5352 -205 5353 -141
rect 5417 -205 5418 -141
rect 5352 -295 5418 -205
rect 5478 -299 5538 733
rect 5598 -359 5658 671
rect 5718 -299 5778 733
rect 5838 -359 5898 671
rect 5958 579 6024 733
rect 5958 515 5959 579
rect 6023 515 6024 579
rect 5958 499 6024 515
rect 5958 435 5959 499
rect 6023 435 6024 499
rect 5958 419 6024 435
rect 5958 355 5959 419
rect 6023 355 6024 419
rect 5958 339 6024 355
rect 5958 275 5959 339
rect 6023 275 6024 339
rect 5958 259 6024 275
rect 5958 195 5959 259
rect 6023 195 6024 259
rect 5958 179 6024 195
rect 5958 115 5959 179
rect 6023 115 6024 179
rect 5958 99 6024 115
rect 5958 35 5959 99
rect 6023 35 6024 99
rect 5958 19 6024 35
rect 5958 -45 5959 19
rect 6023 -45 6024 19
rect 5958 -61 6024 -45
rect 5958 -125 5959 -61
rect 6023 -125 6024 -61
rect 5958 -141 6024 -125
rect 5958 -205 5959 -141
rect 6023 -205 6024 -141
rect 5958 -295 6024 -205
rect 6084 -299 6144 733
rect 6204 -359 6264 671
rect 6324 -299 6384 733
rect 6444 -359 6504 671
rect 6564 579 6630 733
rect 6564 515 6565 579
rect 6629 515 6630 579
rect 6564 499 6630 515
rect 6564 435 6565 499
rect 6629 435 6630 499
rect 6564 419 6630 435
rect 6564 355 6565 419
rect 6629 355 6630 419
rect 6564 339 6630 355
rect 6564 275 6565 339
rect 6629 275 6630 339
rect 6564 259 6630 275
rect 6564 195 6565 259
rect 6629 195 6630 259
rect 6564 179 6630 195
rect 6564 115 6565 179
rect 6629 115 6630 179
rect 6564 99 6630 115
rect 6564 35 6565 99
rect 6629 35 6630 99
rect 6564 19 6630 35
rect 6564 -45 6565 19
rect 6629 -45 6630 19
rect 6564 -61 6630 -45
rect 6564 -125 6565 -61
rect 6629 -125 6630 -61
rect 6564 -141 6630 -125
rect 6564 -205 6565 -141
rect 6629 -205 6630 -141
rect 6564 -295 6630 -205
rect 6690 -299 6750 733
rect 6810 -359 6870 671
rect 6930 -299 6990 733
rect 7050 -359 7110 671
rect 7170 579 7236 733
rect 7170 515 7171 579
rect 7235 515 7236 579
rect 7170 499 7236 515
rect 7170 435 7171 499
rect 7235 435 7236 499
rect 7170 419 7236 435
rect 7170 355 7171 419
rect 7235 355 7236 419
rect 7170 339 7236 355
rect 7170 275 7171 339
rect 7235 275 7236 339
rect 7170 259 7236 275
rect 7170 195 7171 259
rect 7235 195 7236 259
rect 7170 179 7236 195
rect 7170 115 7171 179
rect 7235 115 7236 179
rect 7170 99 7236 115
rect 7170 35 7171 99
rect 7235 35 7236 99
rect 7170 19 7236 35
rect 7170 -45 7171 19
rect 7235 -45 7236 19
rect 7170 -61 7236 -45
rect 7170 -125 7171 -61
rect 7235 -125 7236 -61
rect 7170 -141 7236 -125
rect 7170 -205 7171 -141
rect 7235 -205 7236 -141
rect 7170 -295 7236 -205
rect 7296 -299 7356 733
rect 7416 -359 7476 671
rect 7536 -299 7596 733
rect 7656 -359 7716 671
rect 7776 579 7842 733
rect 7776 515 7777 579
rect 7841 515 7842 579
rect 7776 499 7842 515
rect 7776 435 7777 499
rect 7841 435 7842 499
rect 7776 419 7842 435
rect 7776 355 7777 419
rect 7841 355 7842 419
rect 7776 339 7842 355
rect 7776 275 7777 339
rect 7841 275 7842 339
rect 7776 259 7842 275
rect 7776 195 7777 259
rect 7841 195 7842 259
rect 7776 179 7842 195
rect 7776 115 7777 179
rect 7841 115 7842 179
rect 7776 99 7842 115
rect 7776 35 7777 99
rect 7841 35 7842 99
rect 7776 19 7842 35
rect 7776 -45 7777 19
rect 7841 -45 7842 19
rect 7776 -61 7842 -45
rect 7776 -125 7777 -61
rect 7841 -125 7842 -61
rect 7776 -141 7842 -125
rect 7776 -205 7777 -141
rect 7841 -205 7842 -141
rect 7776 -295 7842 -205
rect 7902 -299 7962 733
rect 8022 -359 8082 671
rect 8142 -299 8202 733
rect 8262 -359 8322 671
rect 8382 579 8448 733
rect 8382 515 8383 579
rect 8447 515 8448 579
rect 8382 499 8448 515
rect 8382 435 8383 499
rect 8447 435 8448 499
rect 8382 419 8448 435
rect 8382 355 8383 419
rect 8447 355 8448 419
rect 8382 339 8448 355
rect 8382 275 8383 339
rect 8447 275 8448 339
rect 8382 259 8448 275
rect 8382 195 8383 259
rect 8447 195 8448 259
rect 8382 179 8448 195
rect 8382 115 8383 179
rect 8447 115 8448 179
rect 8382 99 8448 115
rect 8382 35 8383 99
rect 8447 35 8448 99
rect 8382 19 8448 35
rect 8382 -45 8383 19
rect 8447 -45 8448 19
rect 8382 -61 8448 -45
rect 8382 -125 8383 -61
rect 8447 -125 8448 -61
rect 8382 -141 8448 -125
rect 8382 -205 8383 -141
rect 8447 -205 8448 -141
rect 8382 -295 8448 -205
rect 8508 -299 8568 733
rect 8628 -359 8688 671
rect 8748 -299 8808 733
rect 8868 -359 8928 671
rect 8988 579 9054 733
rect 8988 515 8989 579
rect 9053 515 9054 579
rect 8988 499 9054 515
rect 8988 435 8989 499
rect 9053 435 9054 499
rect 8988 419 9054 435
rect 8988 355 8989 419
rect 9053 355 9054 419
rect 8988 339 9054 355
rect 8988 275 8989 339
rect 9053 275 9054 339
rect 8988 259 9054 275
rect 8988 195 8989 259
rect 9053 195 9054 259
rect 8988 179 9054 195
rect 8988 115 8989 179
rect 9053 115 9054 179
rect 8988 99 9054 115
rect 8988 35 8989 99
rect 9053 35 9054 99
rect 8988 19 9054 35
rect 8988 -45 8989 19
rect 9053 -45 9054 19
rect 8988 -61 9054 -45
rect 8988 -125 8989 -61
rect 9053 -125 9054 -61
rect 8988 -141 9054 -125
rect 8988 -205 8989 -141
rect 9053 -205 9054 -141
rect 8988 -295 9054 -205
rect 9114 -299 9174 733
rect 9234 -359 9294 671
rect 9354 -299 9414 733
rect 9474 -359 9534 671
rect 9594 579 9660 733
rect 9594 515 9595 579
rect 9659 515 9660 579
rect 9594 499 9660 515
rect 9594 435 9595 499
rect 9659 435 9660 499
rect 9594 419 9660 435
rect 9594 355 9595 419
rect 9659 355 9660 419
rect 9594 339 9660 355
rect 9594 275 9595 339
rect 9659 275 9660 339
rect 9594 259 9660 275
rect 9594 195 9595 259
rect 9659 195 9660 259
rect 9594 179 9660 195
rect 9594 115 9595 179
rect 9659 115 9660 179
rect 9594 99 9660 115
rect 9594 35 9595 99
rect 9659 35 9660 99
rect 9594 19 9660 35
rect 9594 -45 9595 19
rect 9659 -45 9660 19
rect 9594 -61 9660 -45
rect 9594 -125 9595 -61
rect 9659 -125 9660 -61
rect 9594 -141 9660 -125
rect 9594 -205 9595 -141
rect 9659 -205 9660 -141
rect 9594 -295 9660 -205
rect 9720 -299 9780 733
rect 9840 -359 9900 671
rect 9960 -299 10020 733
rect 10080 -359 10140 671
rect 10200 579 10266 733
rect 10200 515 10201 579
rect 10265 515 10266 579
rect 10200 499 10266 515
rect 10200 435 10201 499
rect 10265 435 10266 499
rect 10200 419 10266 435
rect 10200 355 10201 419
rect 10265 355 10266 419
rect 10200 339 10266 355
rect 10200 275 10201 339
rect 10265 275 10266 339
rect 10200 259 10266 275
rect 10200 195 10201 259
rect 10265 195 10266 259
rect 10200 179 10266 195
rect 10200 115 10201 179
rect 10265 115 10266 179
rect 10200 99 10266 115
rect 10200 35 10201 99
rect 10265 35 10266 99
rect 10200 19 10266 35
rect 10200 -45 10201 19
rect 10265 -45 10266 19
rect 10200 -61 10266 -45
rect 10200 -125 10201 -61
rect 10265 -125 10266 -61
rect 10200 -141 10266 -125
rect 10200 -205 10201 -141
rect 10265 -205 10266 -141
rect 10200 -295 10266 -205
rect 10326 1739 10392 1829
rect 10326 1675 10327 1739
rect 10391 1675 10392 1739
rect 10326 1659 10392 1675
rect 10326 1595 10327 1659
rect 10391 1595 10392 1659
rect 10326 1579 10392 1595
rect 10326 1515 10327 1579
rect 10391 1515 10392 1579
rect 10326 1499 10392 1515
rect 10326 1435 10327 1499
rect 10391 1435 10392 1499
rect 10326 1419 10392 1435
rect 10326 1355 10327 1419
rect 10391 1355 10392 1419
rect 10326 1339 10392 1355
rect 10326 1275 10327 1339
rect 10391 1275 10392 1339
rect 10326 1259 10392 1275
rect 10326 1195 10327 1259
rect 10391 1195 10392 1259
rect 10326 1179 10392 1195
rect 10326 1115 10327 1179
rect 10391 1115 10392 1179
rect 10326 1099 10392 1115
rect 10326 1035 10327 1099
rect 10391 1035 10392 1099
rect 10326 1019 10392 1035
rect 10326 955 10327 1019
rect 10391 955 10392 1019
rect 10326 801 10392 955
rect 10452 863 10512 1893
rect 10572 801 10632 1833
rect 10692 863 10752 1893
rect 10812 801 10872 1833
rect 10932 1739 10998 1829
rect 10932 1675 10933 1739
rect 10997 1675 10998 1739
rect 10932 1659 10998 1675
rect 10932 1595 10933 1659
rect 10997 1595 10998 1659
rect 10932 1579 10998 1595
rect 10932 1515 10933 1579
rect 10997 1515 10998 1579
rect 10932 1499 10998 1515
rect 10932 1435 10933 1499
rect 10997 1435 10998 1499
rect 10932 1419 10998 1435
rect 10932 1355 10933 1419
rect 10997 1355 10998 1419
rect 10932 1339 10998 1355
rect 10932 1275 10933 1339
rect 10997 1275 10998 1339
rect 10932 1259 10998 1275
rect 10932 1195 10933 1259
rect 10997 1195 10998 1259
rect 10932 1179 10998 1195
rect 10932 1115 10933 1179
rect 10997 1115 10998 1179
rect 10932 1099 10998 1115
rect 10932 1035 10933 1099
rect 10997 1035 10998 1099
rect 10932 1019 10998 1035
rect 10932 955 10933 1019
rect 10997 955 10998 1019
rect 10932 801 10998 955
rect 11058 863 11118 1893
rect 11178 801 11238 1833
rect 11298 863 11358 1893
rect 11418 801 11478 1833
rect 11538 1739 11604 1829
rect 11538 1675 11539 1739
rect 11603 1675 11604 1739
rect 11538 1659 11604 1675
rect 11538 1595 11539 1659
rect 11603 1595 11604 1659
rect 11538 1579 11604 1595
rect 11538 1515 11539 1579
rect 11603 1515 11604 1579
rect 11538 1499 11604 1515
rect 11538 1435 11539 1499
rect 11603 1435 11604 1499
rect 11538 1419 11604 1435
rect 11538 1355 11539 1419
rect 11603 1355 11604 1419
rect 11538 1339 11604 1355
rect 11538 1275 11539 1339
rect 11603 1275 11604 1339
rect 11538 1259 11604 1275
rect 11538 1195 11539 1259
rect 11603 1195 11604 1259
rect 11538 1179 11604 1195
rect 11538 1115 11539 1179
rect 11603 1115 11604 1179
rect 11538 1099 11604 1115
rect 11538 1035 11539 1099
rect 11603 1035 11604 1099
rect 11538 1019 11604 1035
rect 11538 955 11539 1019
rect 11603 955 11604 1019
rect 11538 801 11604 955
rect 11664 863 11724 1893
rect 11784 801 11844 1833
rect 11904 863 11964 1893
rect 12024 801 12084 1833
rect 12144 1739 12210 1829
rect 12144 1675 12145 1739
rect 12209 1675 12210 1739
rect 12144 1659 12210 1675
rect 12144 1595 12145 1659
rect 12209 1595 12210 1659
rect 12144 1579 12210 1595
rect 12144 1515 12145 1579
rect 12209 1515 12210 1579
rect 12144 1499 12210 1515
rect 12144 1435 12145 1499
rect 12209 1435 12210 1499
rect 12144 1419 12210 1435
rect 12144 1355 12145 1419
rect 12209 1355 12210 1419
rect 12144 1339 12210 1355
rect 12144 1275 12145 1339
rect 12209 1275 12210 1339
rect 12144 1259 12210 1275
rect 12144 1195 12145 1259
rect 12209 1195 12210 1259
rect 12144 1179 12210 1195
rect 12144 1115 12145 1179
rect 12209 1115 12210 1179
rect 12144 1099 12210 1115
rect 12144 1035 12145 1099
rect 12209 1035 12210 1099
rect 12144 1019 12210 1035
rect 12144 955 12145 1019
rect 12209 955 12210 1019
rect 12144 801 12210 955
rect 12270 863 12330 1893
rect 12390 801 12450 1833
rect 12510 863 12570 1893
rect 12630 801 12690 1833
rect 12750 1739 12816 1829
rect 12750 1675 12751 1739
rect 12815 1675 12816 1739
rect 12750 1659 12816 1675
rect 12750 1595 12751 1659
rect 12815 1595 12816 1659
rect 12750 1579 12816 1595
rect 12750 1515 12751 1579
rect 12815 1515 12816 1579
rect 12750 1499 12816 1515
rect 12750 1435 12751 1499
rect 12815 1435 12816 1499
rect 12750 1419 12816 1435
rect 12750 1355 12751 1419
rect 12815 1355 12816 1419
rect 12750 1339 12816 1355
rect 12750 1275 12751 1339
rect 12815 1275 12816 1339
rect 12750 1259 12816 1275
rect 12750 1195 12751 1259
rect 12815 1195 12816 1259
rect 12750 1179 12816 1195
rect 12750 1115 12751 1179
rect 12815 1115 12816 1179
rect 12750 1099 12816 1115
rect 12750 1035 12751 1099
rect 12815 1035 12816 1099
rect 12750 1019 12816 1035
rect 12750 955 12751 1019
rect 12815 955 12816 1019
rect 12750 801 12816 955
rect 12876 863 12936 1893
rect 12996 801 13056 1833
rect 13116 863 13176 1893
rect 13236 801 13296 1833
rect 13356 1739 13422 1829
rect 13356 1675 13357 1739
rect 13421 1675 13422 1739
rect 13356 1659 13422 1675
rect 13356 1595 13357 1659
rect 13421 1595 13422 1659
rect 13356 1579 13422 1595
rect 13356 1515 13357 1579
rect 13421 1515 13422 1579
rect 13356 1499 13422 1515
rect 13356 1435 13357 1499
rect 13421 1435 13422 1499
rect 13356 1419 13422 1435
rect 13356 1355 13357 1419
rect 13421 1355 13422 1419
rect 13356 1339 13422 1355
rect 13356 1275 13357 1339
rect 13421 1275 13422 1339
rect 13356 1259 13422 1275
rect 13356 1195 13357 1259
rect 13421 1195 13422 1259
rect 13356 1179 13422 1195
rect 13356 1115 13357 1179
rect 13421 1115 13422 1179
rect 13356 1099 13422 1115
rect 13356 1035 13357 1099
rect 13421 1035 13422 1099
rect 13356 1019 13422 1035
rect 13356 955 13357 1019
rect 13421 955 13422 1019
rect 13356 801 13422 955
rect 13482 863 13542 1893
rect 13602 801 13662 1833
rect 13722 863 13782 1893
rect 13842 801 13902 1833
rect 13962 1739 14028 1829
rect 13962 1675 13963 1739
rect 14027 1675 14028 1739
rect 13962 1659 14028 1675
rect 13962 1595 13963 1659
rect 14027 1595 14028 1659
rect 13962 1579 14028 1595
rect 13962 1515 13963 1579
rect 14027 1515 14028 1579
rect 13962 1499 14028 1515
rect 13962 1435 13963 1499
rect 14027 1435 14028 1499
rect 13962 1419 14028 1435
rect 13962 1355 13963 1419
rect 14027 1355 14028 1419
rect 13962 1339 14028 1355
rect 13962 1275 13963 1339
rect 14027 1275 14028 1339
rect 13962 1259 14028 1275
rect 13962 1195 13963 1259
rect 14027 1195 14028 1259
rect 13962 1179 14028 1195
rect 13962 1115 13963 1179
rect 14027 1115 14028 1179
rect 13962 1099 14028 1115
rect 13962 1035 13963 1099
rect 14027 1035 14028 1099
rect 13962 1019 14028 1035
rect 13962 955 13963 1019
rect 14027 955 14028 1019
rect 13962 801 14028 955
rect 14088 863 14148 1893
rect 14208 801 14268 1833
rect 14328 863 14388 1893
rect 14448 801 14508 1833
rect 14568 1739 14634 1829
rect 14568 1675 14569 1739
rect 14633 1675 14634 1739
rect 14568 1659 14634 1675
rect 14568 1595 14569 1659
rect 14633 1595 14634 1659
rect 14568 1579 14634 1595
rect 14568 1515 14569 1579
rect 14633 1515 14634 1579
rect 14568 1499 14634 1515
rect 14568 1435 14569 1499
rect 14633 1435 14634 1499
rect 14568 1419 14634 1435
rect 14568 1355 14569 1419
rect 14633 1355 14634 1419
rect 14568 1339 14634 1355
rect 14568 1275 14569 1339
rect 14633 1275 14634 1339
rect 14568 1259 14634 1275
rect 14568 1195 14569 1259
rect 14633 1195 14634 1259
rect 14568 1179 14634 1195
rect 14568 1115 14569 1179
rect 14633 1115 14634 1179
rect 14568 1099 14634 1115
rect 14568 1035 14569 1099
rect 14633 1035 14634 1099
rect 14568 1019 14634 1035
rect 14568 955 14569 1019
rect 14633 955 14634 1019
rect 14568 801 14634 955
rect 14694 863 14754 1893
rect 14814 801 14874 1833
rect 14934 863 14994 1893
rect 15054 801 15114 1833
rect 15174 1739 15240 1829
rect 15174 1675 15175 1739
rect 15239 1675 15240 1739
rect 15174 1659 15240 1675
rect 15174 1595 15175 1659
rect 15239 1595 15240 1659
rect 15174 1579 15240 1595
rect 15174 1515 15175 1579
rect 15239 1515 15240 1579
rect 15174 1499 15240 1515
rect 15174 1435 15175 1499
rect 15239 1435 15240 1499
rect 15174 1419 15240 1435
rect 15174 1355 15175 1419
rect 15239 1355 15240 1419
rect 15174 1339 15240 1355
rect 15174 1275 15175 1339
rect 15239 1275 15240 1339
rect 15174 1259 15240 1275
rect 15174 1195 15175 1259
rect 15239 1195 15240 1259
rect 15174 1179 15240 1195
rect 15174 1115 15175 1179
rect 15239 1115 15240 1179
rect 15174 1099 15240 1115
rect 15174 1035 15175 1099
rect 15239 1035 15240 1099
rect 15174 1019 15240 1035
rect 15174 955 15175 1019
rect 15239 955 15240 1019
rect 15174 801 15240 955
rect 15300 863 15360 1893
rect 15420 801 15480 1833
rect 15540 863 15600 1893
rect 15660 801 15720 1833
rect 15780 1739 15846 1829
rect 15780 1675 15781 1739
rect 15845 1675 15846 1739
rect 15780 1659 15846 1675
rect 15780 1595 15781 1659
rect 15845 1595 15846 1659
rect 15780 1579 15846 1595
rect 15780 1515 15781 1579
rect 15845 1515 15846 1579
rect 15780 1499 15846 1515
rect 15780 1435 15781 1499
rect 15845 1435 15846 1499
rect 15780 1419 15846 1435
rect 15780 1355 15781 1419
rect 15845 1355 15846 1419
rect 15780 1339 15846 1355
rect 15780 1275 15781 1339
rect 15845 1275 15846 1339
rect 15780 1259 15846 1275
rect 15780 1195 15781 1259
rect 15845 1195 15846 1259
rect 15780 1179 15846 1195
rect 15780 1115 15781 1179
rect 15845 1115 15846 1179
rect 15780 1099 15846 1115
rect 15780 1035 15781 1099
rect 15845 1035 15846 1099
rect 15780 1019 15846 1035
rect 15780 955 15781 1019
rect 15845 955 15846 1019
rect 15780 801 15846 955
rect 15906 863 15966 1893
rect 16026 801 16086 1833
rect 16146 863 16206 1893
rect 16266 801 16326 1833
rect 16386 1739 16452 1829
rect 16386 1675 16387 1739
rect 16451 1675 16452 1739
rect 16386 1659 16452 1675
rect 16386 1595 16387 1659
rect 16451 1595 16452 1659
rect 16386 1579 16452 1595
rect 16386 1515 16387 1579
rect 16451 1515 16452 1579
rect 16386 1499 16452 1515
rect 16386 1435 16387 1499
rect 16451 1435 16452 1499
rect 16386 1419 16452 1435
rect 16386 1355 16387 1419
rect 16451 1355 16452 1419
rect 16386 1339 16452 1355
rect 16386 1275 16387 1339
rect 16451 1275 16452 1339
rect 16386 1259 16452 1275
rect 16386 1195 16387 1259
rect 16451 1195 16452 1259
rect 16386 1179 16452 1195
rect 16386 1115 16387 1179
rect 16451 1115 16452 1179
rect 16386 1099 16452 1115
rect 16386 1035 16387 1099
rect 16451 1035 16452 1099
rect 16386 1019 16452 1035
rect 16386 955 16387 1019
rect 16451 955 16452 1019
rect 16386 801 16452 955
rect 16512 863 16572 1893
rect 16632 801 16692 1833
rect 16752 863 16812 1893
rect 16872 801 16932 1833
rect 16992 1739 17058 1829
rect 16992 1675 16993 1739
rect 17057 1675 17058 1739
rect 16992 1659 17058 1675
rect 16992 1595 16993 1659
rect 17057 1595 17058 1659
rect 16992 1579 17058 1595
rect 16992 1515 16993 1579
rect 17057 1515 17058 1579
rect 16992 1499 17058 1515
rect 16992 1435 16993 1499
rect 17057 1435 17058 1499
rect 16992 1419 17058 1435
rect 16992 1355 16993 1419
rect 17057 1355 17058 1419
rect 16992 1339 17058 1355
rect 16992 1275 16993 1339
rect 17057 1275 17058 1339
rect 16992 1259 17058 1275
rect 16992 1195 16993 1259
rect 17057 1195 17058 1259
rect 16992 1179 17058 1195
rect 16992 1115 16993 1179
rect 17057 1115 17058 1179
rect 16992 1099 17058 1115
rect 16992 1035 16993 1099
rect 17057 1035 17058 1099
rect 16992 1019 17058 1035
rect 16992 955 16993 1019
rect 17057 955 17058 1019
rect 16992 801 17058 955
rect 17118 863 17178 1893
rect 17238 801 17298 1833
rect 17358 863 17418 1893
rect 17478 801 17538 1833
rect 17598 1739 17664 1829
rect 17598 1675 17599 1739
rect 17663 1675 17664 1739
rect 17598 1659 17664 1675
rect 17598 1595 17599 1659
rect 17663 1595 17664 1659
rect 17598 1579 17664 1595
rect 17598 1515 17599 1579
rect 17663 1515 17664 1579
rect 17598 1499 17664 1515
rect 17598 1435 17599 1499
rect 17663 1435 17664 1499
rect 17598 1419 17664 1435
rect 17598 1355 17599 1419
rect 17663 1355 17664 1419
rect 17598 1339 17664 1355
rect 17598 1275 17599 1339
rect 17663 1275 17664 1339
rect 17598 1259 17664 1275
rect 17598 1195 17599 1259
rect 17663 1195 17664 1259
rect 17598 1179 17664 1195
rect 17598 1115 17599 1179
rect 17663 1115 17664 1179
rect 17598 1099 17664 1115
rect 17598 1035 17599 1099
rect 17663 1035 17664 1099
rect 17598 1019 17664 1035
rect 17598 955 17599 1019
rect 17663 955 17664 1019
rect 17598 801 17664 955
rect 17724 863 17784 1893
rect 17844 801 17904 1833
rect 17964 863 18024 1893
rect 18084 801 18144 1833
rect 18204 1739 18270 1829
rect 18204 1675 18205 1739
rect 18269 1675 18270 1739
rect 18204 1659 18270 1675
rect 18204 1595 18205 1659
rect 18269 1595 18270 1659
rect 18204 1579 18270 1595
rect 18204 1515 18205 1579
rect 18269 1515 18270 1579
rect 18204 1499 18270 1515
rect 18204 1435 18205 1499
rect 18269 1435 18270 1499
rect 18204 1419 18270 1435
rect 18204 1355 18205 1419
rect 18269 1355 18270 1419
rect 18204 1339 18270 1355
rect 18204 1275 18205 1339
rect 18269 1275 18270 1339
rect 18204 1259 18270 1275
rect 18204 1195 18205 1259
rect 18269 1195 18270 1259
rect 18204 1179 18270 1195
rect 18204 1115 18205 1179
rect 18269 1115 18270 1179
rect 18204 1099 18270 1115
rect 18204 1035 18205 1099
rect 18269 1035 18270 1099
rect 18204 1019 18270 1035
rect 18204 955 18205 1019
rect 18269 955 18270 1019
rect 18204 801 18270 955
rect 18330 863 18390 1893
rect 18450 801 18510 1833
rect 18570 863 18630 1893
rect 18690 801 18750 1833
rect 18810 1739 18876 1829
rect 18810 1675 18811 1739
rect 18875 1675 18876 1739
rect 18810 1659 18876 1675
rect 18810 1595 18811 1659
rect 18875 1595 18876 1659
rect 18810 1579 18876 1595
rect 18810 1515 18811 1579
rect 18875 1515 18876 1579
rect 18810 1499 18876 1515
rect 18810 1435 18811 1499
rect 18875 1435 18876 1499
rect 18810 1419 18876 1435
rect 18810 1355 18811 1419
rect 18875 1355 18876 1419
rect 18810 1339 18876 1355
rect 18810 1275 18811 1339
rect 18875 1275 18876 1339
rect 18810 1259 18876 1275
rect 18810 1195 18811 1259
rect 18875 1195 18876 1259
rect 18810 1179 18876 1195
rect 18810 1115 18811 1179
rect 18875 1115 18876 1179
rect 18810 1099 18876 1115
rect 18810 1035 18811 1099
rect 18875 1035 18876 1099
rect 18810 1019 18876 1035
rect 18810 955 18811 1019
rect 18875 955 18876 1019
rect 18810 801 18876 955
rect 18936 863 18996 1893
rect 19056 801 19116 1833
rect 19176 863 19236 1893
rect 19296 801 19356 1833
rect 19416 1739 19482 1829
rect 19416 1675 19417 1739
rect 19481 1675 19482 1739
rect 19416 1659 19482 1675
rect 19416 1595 19417 1659
rect 19481 1595 19482 1659
rect 19416 1579 19482 1595
rect 19416 1515 19417 1579
rect 19481 1515 19482 1579
rect 19416 1499 19482 1515
rect 19416 1435 19417 1499
rect 19481 1435 19482 1499
rect 19416 1419 19482 1435
rect 19416 1355 19417 1419
rect 19481 1355 19482 1419
rect 19416 1339 19482 1355
rect 19416 1275 19417 1339
rect 19481 1275 19482 1339
rect 19416 1259 19482 1275
rect 19416 1195 19417 1259
rect 19481 1195 19482 1259
rect 19416 1179 19482 1195
rect 19416 1115 19417 1179
rect 19481 1115 19482 1179
rect 19416 1099 19482 1115
rect 19416 1035 19417 1099
rect 19481 1035 19482 1099
rect 19416 1019 19482 1035
rect 19416 955 19417 1019
rect 19481 955 19482 1019
rect 19416 801 19482 955
rect 19542 863 19602 1893
rect 19662 801 19722 1833
rect 19782 863 19842 1893
rect 19902 801 19962 1833
rect 20022 1739 20088 1829
rect 20022 1675 20023 1739
rect 20087 1675 20088 1739
rect 20022 1659 20088 1675
rect 20022 1595 20023 1659
rect 20087 1595 20088 1659
rect 20022 1579 20088 1595
rect 20022 1515 20023 1579
rect 20087 1515 20088 1579
rect 20022 1499 20088 1515
rect 20022 1435 20023 1499
rect 20087 1435 20088 1499
rect 20022 1419 20088 1435
rect 20022 1355 20023 1419
rect 20087 1355 20088 1419
rect 20022 1339 20088 1355
rect 20022 1275 20023 1339
rect 20087 1275 20088 1339
rect 20022 1259 20088 1275
rect 20022 1195 20023 1259
rect 20087 1195 20088 1259
rect 20022 1179 20088 1195
rect 20022 1115 20023 1179
rect 20087 1115 20088 1179
rect 20022 1099 20088 1115
rect 20022 1035 20023 1099
rect 20087 1035 20088 1099
rect 20022 1019 20088 1035
rect 20022 955 20023 1019
rect 20087 955 20088 1019
rect 20022 801 20088 955
rect 10326 799 20088 801
rect 10326 735 10430 799
rect 10494 735 10510 799
rect 10574 735 10590 799
rect 10654 735 10670 799
rect 10734 735 10750 799
rect 10814 735 10830 799
rect 10894 735 11036 799
rect 11100 735 11116 799
rect 11180 735 11196 799
rect 11260 735 11276 799
rect 11340 735 11356 799
rect 11420 735 11436 799
rect 11500 735 11642 799
rect 11706 735 11722 799
rect 11786 735 11802 799
rect 11866 735 11882 799
rect 11946 735 11962 799
rect 12026 735 12042 799
rect 12106 735 12248 799
rect 12312 735 12328 799
rect 12392 735 12408 799
rect 12472 735 12488 799
rect 12552 735 12568 799
rect 12632 735 12648 799
rect 12712 735 12854 799
rect 12918 735 12934 799
rect 12998 735 13014 799
rect 13078 735 13094 799
rect 13158 735 13174 799
rect 13238 735 13254 799
rect 13318 735 13460 799
rect 13524 735 13540 799
rect 13604 735 13620 799
rect 13684 735 13700 799
rect 13764 735 13780 799
rect 13844 735 13860 799
rect 13924 735 14066 799
rect 14130 735 14146 799
rect 14210 735 14226 799
rect 14290 735 14306 799
rect 14370 735 14386 799
rect 14450 735 14466 799
rect 14530 735 14672 799
rect 14736 735 14752 799
rect 14816 735 14832 799
rect 14896 735 14912 799
rect 14976 735 14992 799
rect 15056 735 15072 799
rect 15136 735 15278 799
rect 15342 735 15358 799
rect 15422 735 15438 799
rect 15502 735 15518 799
rect 15582 735 15598 799
rect 15662 735 15678 799
rect 15742 735 15884 799
rect 15948 735 15964 799
rect 16028 735 16044 799
rect 16108 735 16124 799
rect 16188 735 16204 799
rect 16268 735 16284 799
rect 16348 735 16490 799
rect 16554 735 16570 799
rect 16634 735 16650 799
rect 16714 735 16730 799
rect 16794 735 16810 799
rect 16874 735 16890 799
rect 16954 735 17096 799
rect 17160 735 17176 799
rect 17240 735 17256 799
rect 17320 735 17336 799
rect 17400 735 17416 799
rect 17480 735 17496 799
rect 17560 735 17702 799
rect 17766 735 17782 799
rect 17846 735 17862 799
rect 17926 735 17942 799
rect 18006 735 18022 799
rect 18086 735 18102 799
rect 18166 735 18308 799
rect 18372 735 18388 799
rect 18452 735 18468 799
rect 18532 735 18548 799
rect 18612 735 18628 799
rect 18692 735 18708 799
rect 18772 735 18914 799
rect 18978 735 18994 799
rect 19058 735 19074 799
rect 19138 735 19154 799
rect 19218 735 19234 799
rect 19298 735 19314 799
rect 19378 735 19520 799
rect 19584 735 19600 799
rect 19664 735 19680 799
rect 19744 735 19760 799
rect 19824 735 19840 799
rect 19904 735 19920 799
rect 19984 735 20088 799
rect 10326 733 20088 735
rect 10326 579 10392 733
rect 10326 515 10327 579
rect 10391 515 10392 579
rect 10326 499 10392 515
rect 10326 435 10327 499
rect 10391 435 10392 499
rect 10326 419 10392 435
rect 10326 355 10327 419
rect 10391 355 10392 419
rect 10326 339 10392 355
rect 10326 275 10327 339
rect 10391 275 10392 339
rect 10326 259 10392 275
rect 10326 195 10327 259
rect 10391 195 10392 259
rect 10326 179 10392 195
rect 10326 115 10327 179
rect 10391 115 10392 179
rect 10326 99 10392 115
rect 10326 35 10327 99
rect 10391 35 10392 99
rect 10326 19 10392 35
rect 10326 -45 10327 19
rect 10391 -45 10392 19
rect 10326 -61 10392 -45
rect 10326 -125 10327 -61
rect 10391 -125 10392 -61
rect 10326 -141 10392 -125
rect 10326 -205 10327 -141
rect 10391 -205 10392 -141
rect 10326 -295 10392 -205
rect 10452 -299 10512 733
rect 10572 -359 10632 671
rect 10692 -299 10752 733
rect 10812 -359 10872 671
rect 10932 579 10998 733
rect 10932 515 10933 579
rect 10997 515 10998 579
rect 10932 499 10998 515
rect 10932 435 10933 499
rect 10997 435 10998 499
rect 10932 419 10998 435
rect 10932 355 10933 419
rect 10997 355 10998 419
rect 10932 339 10998 355
rect 10932 275 10933 339
rect 10997 275 10998 339
rect 10932 259 10998 275
rect 10932 195 10933 259
rect 10997 195 10998 259
rect 10932 179 10998 195
rect 10932 115 10933 179
rect 10997 115 10998 179
rect 10932 99 10998 115
rect 10932 35 10933 99
rect 10997 35 10998 99
rect 10932 19 10998 35
rect 10932 -45 10933 19
rect 10997 -45 10998 19
rect 10932 -61 10998 -45
rect 10932 -125 10933 -61
rect 10997 -125 10998 -61
rect 10932 -141 10998 -125
rect 10932 -205 10933 -141
rect 10997 -205 10998 -141
rect 10932 -295 10998 -205
rect 11058 -299 11118 733
rect 11178 -359 11238 671
rect 11298 -299 11358 733
rect 11418 -359 11478 671
rect 11538 579 11604 733
rect 11538 515 11539 579
rect 11603 515 11604 579
rect 11538 499 11604 515
rect 11538 435 11539 499
rect 11603 435 11604 499
rect 11538 419 11604 435
rect 11538 355 11539 419
rect 11603 355 11604 419
rect 11538 339 11604 355
rect 11538 275 11539 339
rect 11603 275 11604 339
rect 11538 259 11604 275
rect 11538 195 11539 259
rect 11603 195 11604 259
rect 11538 179 11604 195
rect 11538 115 11539 179
rect 11603 115 11604 179
rect 11538 99 11604 115
rect 11538 35 11539 99
rect 11603 35 11604 99
rect 11538 19 11604 35
rect 11538 -45 11539 19
rect 11603 -45 11604 19
rect 11538 -61 11604 -45
rect 11538 -125 11539 -61
rect 11603 -125 11604 -61
rect 11538 -141 11604 -125
rect 11538 -205 11539 -141
rect 11603 -205 11604 -141
rect 11538 -295 11604 -205
rect 11664 -299 11724 733
rect 11784 -359 11844 671
rect 11904 -299 11964 733
rect 12024 -359 12084 671
rect 12144 579 12210 733
rect 12144 515 12145 579
rect 12209 515 12210 579
rect 12144 499 12210 515
rect 12144 435 12145 499
rect 12209 435 12210 499
rect 12144 419 12210 435
rect 12144 355 12145 419
rect 12209 355 12210 419
rect 12144 339 12210 355
rect 12144 275 12145 339
rect 12209 275 12210 339
rect 12144 259 12210 275
rect 12144 195 12145 259
rect 12209 195 12210 259
rect 12144 179 12210 195
rect 12144 115 12145 179
rect 12209 115 12210 179
rect 12144 99 12210 115
rect 12144 35 12145 99
rect 12209 35 12210 99
rect 12144 19 12210 35
rect 12144 -45 12145 19
rect 12209 -45 12210 19
rect 12144 -61 12210 -45
rect 12144 -125 12145 -61
rect 12209 -125 12210 -61
rect 12144 -141 12210 -125
rect 12144 -205 12145 -141
rect 12209 -205 12210 -141
rect 12144 -295 12210 -205
rect 12270 -299 12330 733
rect 12390 -359 12450 671
rect 12510 -299 12570 733
rect 12630 -359 12690 671
rect 12750 579 12816 733
rect 12750 515 12751 579
rect 12815 515 12816 579
rect 12750 499 12816 515
rect 12750 435 12751 499
rect 12815 435 12816 499
rect 12750 419 12816 435
rect 12750 355 12751 419
rect 12815 355 12816 419
rect 12750 339 12816 355
rect 12750 275 12751 339
rect 12815 275 12816 339
rect 12750 259 12816 275
rect 12750 195 12751 259
rect 12815 195 12816 259
rect 12750 179 12816 195
rect 12750 115 12751 179
rect 12815 115 12816 179
rect 12750 99 12816 115
rect 12750 35 12751 99
rect 12815 35 12816 99
rect 12750 19 12816 35
rect 12750 -45 12751 19
rect 12815 -45 12816 19
rect 12750 -61 12816 -45
rect 12750 -125 12751 -61
rect 12815 -125 12816 -61
rect 12750 -141 12816 -125
rect 12750 -205 12751 -141
rect 12815 -205 12816 -141
rect 12750 -295 12816 -205
rect 12876 -299 12936 733
rect 12996 -359 13056 671
rect 13116 -299 13176 733
rect 13236 -359 13296 671
rect 13356 579 13422 733
rect 13356 515 13357 579
rect 13421 515 13422 579
rect 13356 499 13422 515
rect 13356 435 13357 499
rect 13421 435 13422 499
rect 13356 419 13422 435
rect 13356 355 13357 419
rect 13421 355 13422 419
rect 13356 339 13422 355
rect 13356 275 13357 339
rect 13421 275 13422 339
rect 13356 259 13422 275
rect 13356 195 13357 259
rect 13421 195 13422 259
rect 13356 179 13422 195
rect 13356 115 13357 179
rect 13421 115 13422 179
rect 13356 99 13422 115
rect 13356 35 13357 99
rect 13421 35 13422 99
rect 13356 19 13422 35
rect 13356 -45 13357 19
rect 13421 -45 13422 19
rect 13356 -61 13422 -45
rect 13356 -125 13357 -61
rect 13421 -125 13422 -61
rect 13356 -141 13422 -125
rect 13356 -205 13357 -141
rect 13421 -205 13422 -141
rect 13356 -295 13422 -205
rect 13482 -299 13542 733
rect 13602 -359 13662 671
rect 13722 -299 13782 733
rect 13842 -359 13902 671
rect 13962 579 14028 733
rect 13962 515 13963 579
rect 14027 515 14028 579
rect 13962 499 14028 515
rect 13962 435 13963 499
rect 14027 435 14028 499
rect 13962 419 14028 435
rect 13962 355 13963 419
rect 14027 355 14028 419
rect 13962 339 14028 355
rect 13962 275 13963 339
rect 14027 275 14028 339
rect 13962 259 14028 275
rect 13962 195 13963 259
rect 14027 195 14028 259
rect 13962 179 14028 195
rect 13962 115 13963 179
rect 14027 115 14028 179
rect 13962 99 14028 115
rect 13962 35 13963 99
rect 14027 35 14028 99
rect 13962 19 14028 35
rect 13962 -45 13963 19
rect 14027 -45 14028 19
rect 13962 -61 14028 -45
rect 13962 -125 13963 -61
rect 14027 -125 14028 -61
rect 13962 -141 14028 -125
rect 13962 -205 13963 -141
rect 14027 -205 14028 -141
rect 13962 -295 14028 -205
rect 14088 -299 14148 733
rect 14208 -359 14268 671
rect 14328 -299 14388 733
rect 14448 -359 14508 671
rect 14568 579 14634 733
rect 14568 515 14569 579
rect 14633 515 14634 579
rect 14568 499 14634 515
rect 14568 435 14569 499
rect 14633 435 14634 499
rect 14568 419 14634 435
rect 14568 355 14569 419
rect 14633 355 14634 419
rect 14568 339 14634 355
rect 14568 275 14569 339
rect 14633 275 14634 339
rect 14568 259 14634 275
rect 14568 195 14569 259
rect 14633 195 14634 259
rect 14568 179 14634 195
rect 14568 115 14569 179
rect 14633 115 14634 179
rect 14568 99 14634 115
rect 14568 35 14569 99
rect 14633 35 14634 99
rect 14568 19 14634 35
rect 14568 -45 14569 19
rect 14633 -45 14634 19
rect 14568 -61 14634 -45
rect 14568 -125 14569 -61
rect 14633 -125 14634 -61
rect 14568 -141 14634 -125
rect 14568 -205 14569 -141
rect 14633 -205 14634 -141
rect 14568 -295 14634 -205
rect 14694 -299 14754 733
rect 14814 -359 14874 671
rect 14934 -299 14994 733
rect 15054 -359 15114 671
rect 15174 579 15240 733
rect 15174 515 15175 579
rect 15239 515 15240 579
rect 15174 499 15240 515
rect 15174 435 15175 499
rect 15239 435 15240 499
rect 15174 419 15240 435
rect 15174 355 15175 419
rect 15239 355 15240 419
rect 15174 339 15240 355
rect 15174 275 15175 339
rect 15239 275 15240 339
rect 15174 259 15240 275
rect 15174 195 15175 259
rect 15239 195 15240 259
rect 15174 179 15240 195
rect 15174 115 15175 179
rect 15239 115 15240 179
rect 15174 99 15240 115
rect 15174 35 15175 99
rect 15239 35 15240 99
rect 15174 19 15240 35
rect 15174 -45 15175 19
rect 15239 -45 15240 19
rect 15174 -61 15240 -45
rect 15174 -125 15175 -61
rect 15239 -125 15240 -61
rect 15174 -141 15240 -125
rect 15174 -205 15175 -141
rect 15239 -205 15240 -141
rect 15174 -295 15240 -205
rect 15300 -299 15360 733
rect 15420 -359 15480 671
rect 15540 -299 15600 733
rect 15660 -359 15720 671
rect 15780 579 15846 733
rect 15780 515 15781 579
rect 15845 515 15846 579
rect 15780 499 15846 515
rect 15780 435 15781 499
rect 15845 435 15846 499
rect 15780 419 15846 435
rect 15780 355 15781 419
rect 15845 355 15846 419
rect 15780 339 15846 355
rect 15780 275 15781 339
rect 15845 275 15846 339
rect 15780 259 15846 275
rect 15780 195 15781 259
rect 15845 195 15846 259
rect 15780 179 15846 195
rect 15780 115 15781 179
rect 15845 115 15846 179
rect 15780 99 15846 115
rect 15780 35 15781 99
rect 15845 35 15846 99
rect 15780 19 15846 35
rect 15780 -45 15781 19
rect 15845 -45 15846 19
rect 15780 -61 15846 -45
rect 15780 -125 15781 -61
rect 15845 -125 15846 -61
rect 15780 -141 15846 -125
rect 15780 -205 15781 -141
rect 15845 -205 15846 -141
rect 15780 -295 15846 -205
rect 15906 -299 15966 733
rect 16026 -359 16086 671
rect 16146 -299 16206 733
rect 16266 -359 16326 671
rect 16386 579 16452 733
rect 16386 515 16387 579
rect 16451 515 16452 579
rect 16386 499 16452 515
rect 16386 435 16387 499
rect 16451 435 16452 499
rect 16386 419 16452 435
rect 16386 355 16387 419
rect 16451 355 16452 419
rect 16386 339 16452 355
rect 16386 275 16387 339
rect 16451 275 16452 339
rect 16386 259 16452 275
rect 16386 195 16387 259
rect 16451 195 16452 259
rect 16386 179 16452 195
rect 16386 115 16387 179
rect 16451 115 16452 179
rect 16386 99 16452 115
rect 16386 35 16387 99
rect 16451 35 16452 99
rect 16386 19 16452 35
rect 16386 -45 16387 19
rect 16451 -45 16452 19
rect 16386 -61 16452 -45
rect 16386 -125 16387 -61
rect 16451 -125 16452 -61
rect 16386 -141 16452 -125
rect 16386 -205 16387 -141
rect 16451 -205 16452 -141
rect 16386 -295 16452 -205
rect 16512 -299 16572 733
rect 16632 -359 16692 671
rect 16752 -299 16812 733
rect 16872 -359 16932 671
rect 16992 579 17058 733
rect 16992 515 16993 579
rect 17057 515 17058 579
rect 16992 499 17058 515
rect 16992 435 16993 499
rect 17057 435 17058 499
rect 16992 419 17058 435
rect 16992 355 16993 419
rect 17057 355 17058 419
rect 16992 339 17058 355
rect 16992 275 16993 339
rect 17057 275 17058 339
rect 16992 259 17058 275
rect 16992 195 16993 259
rect 17057 195 17058 259
rect 16992 179 17058 195
rect 16992 115 16993 179
rect 17057 115 17058 179
rect 16992 99 17058 115
rect 16992 35 16993 99
rect 17057 35 17058 99
rect 16992 19 17058 35
rect 16992 -45 16993 19
rect 17057 -45 17058 19
rect 16992 -61 17058 -45
rect 16992 -125 16993 -61
rect 17057 -125 17058 -61
rect 16992 -141 17058 -125
rect 16992 -205 16993 -141
rect 17057 -205 17058 -141
rect 16992 -295 17058 -205
rect 17118 -299 17178 733
rect 17238 -359 17298 671
rect 17358 -299 17418 733
rect 17478 -359 17538 671
rect 17598 579 17664 733
rect 17598 515 17599 579
rect 17663 515 17664 579
rect 17598 499 17664 515
rect 17598 435 17599 499
rect 17663 435 17664 499
rect 17598 419 17664 435
rect 17598 355 17599 419
rect 17663 355 17664 419
rect 17598 339 17664 355
rect 17598 275 17599 339
rect 17663 275 17664 339
rect 17598 259 17664 275
rect 17598 195 17599 259
rect 17663 195 17664 259
rect 17598 179 17664 195
rect 17598 115 17599 179
rect 17663 115 17664 179
rect 17598 99 17664 115
rect 17598 35 17599 99
rect 17663 35 17664 99
rect 17598 19 17664 35
rect 17598 -45 17599 19
rect 17663 -45 17664 19
rect 17598 -61 17664 -45
rect 17598 -125 17599 -61
rect 17663 -125 17664 -61
rect 17598 -141 17664 -125
rect 17598 -205 17599 -141
rect 17663 -205 17664 -141
rect 17598 -295 17664 -205
rect 17724 -299 17784 733
rect 17844 -359 17904 671
rect 17964 -299 18024 733
rect 18084 -359 18144 671
rect 18204 579 18270 733
rect 18204 515 18205 579
rect 18269 515 18270 579
rect 18204 499 18270 515
rect 18204 435 18205 499
rect 18269 435 18270 499
rect 18204 419 18270 435
rect 18204 355 18205 419
rect 18269 355 18270 419
rect 18204 339 18270 355
rect 18204 275 18205 339
rect 18269 275 18270 339
rect 18204 259 18270 275
rect 18204 195 18205 259
rect 18269 195 18270 259
rect 18204 179 18270 195
rect 18204 115 18205 179
rect 18269 115 18270 179
rect 18204 99 18270 115
rect 18204 35 18205 99
rect 18269 35 18270 99
rect 18204 19 18270 35
rect 18204 -45 18205 19
rect 18269 -45 18270 19
rect 18204 -61 18270 -45
rect 18204 -125 18205 -61
rect 18269 -125 18270 -61
rect 18204 -141 18270 -125
rect 18204 -205 18205 -141
rect 18269 -205 18270 -141
rect 18204 -295 18270 -205
rect 18330 -299 18390 733
rect 18450 -359 18510 671
rect 18570 -299 18630 733
rect 18690 -359 18750 671
rect 18810 579 18876 733
rect 18810 515 18811 579
rect 18875 515 18876 579
rect 18810 499 18876 515
rect 18810 435 18811 499
rect 18875 435 18876 499
rect 18810 419 18876 435
rect 18810 355 18811 419
rect 18875 355 18876 419
rect 18810 339 18876 355
rect 18810 275 18811 339
rect 18875 275 18876 339
rect 18810 259 18876 275
rect 18810 195 18811 259
rect 18875 195 18876 259
rect 18810 179 18876 195
rect 18810 115 18811 179
rect 18875 115 18876 179
rect 18810 99 18876 115
rect 18810 35 18811 99
rect 18875 35 18876 99
rect 18810 19 18876 35
rect 18810 -45 18811 19
rect 18875 -45 18876 19
rect 18810 -61 18876 -45
rect 18810 -125 18811 -61
rect 18875 -125 18876 -61
rect 18810 -141 18876 -125
rect 18810 -205 18811 -141
rect 18875 -205 18876 -141
rect 18810 -295 18876 -205
rect 18936 -299 18996 733
rect 19056 -359 19116 671
rect 19176 -299 19236 733
rect 19296 -359 19356 671
rect 19416 579 19482 733
rect 19416 515 19417 579
rect 19481 515 19482 579
rect 19416 499 19482 515
rect 19416 435 19417 499
rect 19481 435 19482 499
rect 19416 419 19482 435
rect 19416 355 19417 419
rect 19481 355 19482 419
rect 19416 339 19482 355
rect 19416 275 19417 339
rect 19481 275 19482 339
rect 19416 259 19482 275
rect 19416 195 19417 259
rect 19481 195 19482 259
rect 19416 179 19482 195
rect 19416 115 19417 179
rect 19481 115 19482 179
rect 19416 99 19482 115
rect 19416 35 19417 99
rect 19481 35 19482 99
rect 19416 19 19482 35
rect 19416 -45 19417 19
rect 19481 -45 19482 19
rect 19416 -61 19482 -45
rect 19416 -125 19417 -61
rect 19481 -125 19482 -61
rect 19416 -141 19482 -125
rect 19416 -205 19417 -141
rect 19481 -205 19482 -141
rect 19416 -295 19482 -205
rect 19542 -299 19602 733
rect 19662 -359 19722 671
rect 19782 -299 19842 733
rect 19902 -359 19962 671
rect 20022 579 20088 733
rect 20022 515 20023 579
rect 20087 515 20088 579
rect 20022 499 20088 515
rect 20022 435 20023 499
rect 20087 435 20088 499
rect 20022 419 20088 435
rect 20022 355 20023 419
rect 20087 355 20088 419
rect 20022 339 20088 355
rect 20022 275 20023 339
rect 20087 275 20088 339
rect 20022 259 20088 275
rect 20022 195 20023 259
rect 20087 195 20088 259
rect 20022 179 20088 195
rect 20022 115 20023 179
rect 20087 115 20088 179
rect 20022 99 20088 115
rect 20022 35 20023 99
rect 20087 35 20088 99
rect 20022 19 20088 35
rect 20022 -45 20023 19
rect 20087 -45 20088 19
rect 20022 -61 20088 -45
rect 20022 -125 20023 -61
rect 20087 -125 20088 -61
rect 20022 -141 20088 -125
rect 20022 -205 20023 -141
rect 20087 -205 20088 -141
rect 20022 -295 20088 -205
rect 20148 1739 20214 1829
rect 20148 1675 20149 1739
rect 20213 1675 20214 1739
rect 20148 1659 20214 1675
rect 20148 1595 20149 1659
rect 20213 1595 20214 1659
rect 20148 1579 20214 1595
rect 20148 1515 20149 1579
rect 20213 1515 20214 1579
rect 20148 1499 20214 1515
rect 20148 1435 20149 1499
rect 20213 1435 20214 1499
rect 20148 1419 20214 1435
rect 20148 1355 20149 1419
rect 20213 1355 20214 1419
rect 20148 1339 20214 1355
rect 20148 1275 20149 1339
rect 20213 1275 20214 1339
rect 20148 1259 20214 1275
rect 20148 1195 20149 1259
rect 20213 1195 20214 1259
rect 20148 1179 20214 1195
rect 20148 1115 20149 1179
rect 20213 1115 20214 1179
rect 20148 1099 20214 1115
rect 20148 1035 20149 1099
rect 20213 1035 20214 1099
rect 20148 1019 20214 1035
rect 20148 955 20149 1019
rect 20213 955 20214 1019
rect 20148 801 20214 955
rect 20274 863 20334 1893
rect 20394 801 20454 1833
rect 20514 863 20574 1893
rect 20634 801 20694 1833
rect 20754 1739 20820 1829
rect 20754 1675 20755 1739
rect 20819 1675 20820 1739
rect 20754 1659 20820 1675
rect 20754 1595 20755 1659
rect 20819 1595 20820 1659
rect 20754 1579 20820 1595
rect 20754 1515 20755 1579
rect 20819 1515 20820 1579
rect 20754 1499 20820 1515
rect 20754 1435 20755 1499
rect 20819 1435 20820 1499
rect 20754 1419 20820 1435
rect 20754 1355 20755 1419
rect 20819 1355 20820 1419
rect 20754 1339 20820 1355
rect 20754 1275 20755 1339
rect 20819 1275 20820 1339
rect 20754 1259 20820 1275
rect 20754 1195 20755 1259
rect 20819 1195 20820 1259
rect 20754 1179 20820 1195
rect 20754 1115 20755 1179
rect 20819 1115 20820 1179
rect 20754 1099 20820 1115
rect 20754 1035 20755 1099
rect 20819 1035 20820 1099
rect 20754 1019 20820 1035
rect 20754 955 20755 1019
rect 20819 955 20820 1019
rect 20754 801 20820 955
rect 20880 863 20940 1893
rect 21000 801 21060 1833
rect 21120 863 21180 1893
rect 21240 801 21300 1833
rect 21360 1739 21426 1829
rect 21360 1675 21361 1739
rect 21425 1675 21426 1739
rect 21360 1659 21426 1675
rect 21360 1595 21361 1659
rect 21425 1595 21426 1659
rect 21360 1579 21426 1595
rect 21360 1515 21361 1579
rect 21425 1515 21426 1579
rect 21360 1499 21426 1515
rect 21360 1435 21361 1499
rect 21425 1435 21426 1499
rect 21360 1419 21426 1435
rect 21360 1355 21361 1419
rect 21425 1355 21426 1419
rect 21360 1339 21426 1355
rect 21360 1275 21361 1339
rect 21425 1275 21426 1339
rect 21360 1259 21426 1275
rect 21360 1195 21361 1259
rect 21425 1195 21426 1259
rect 21360 1179 21426 1195
rect 21360 1115 21361 1179
rect 21425 1115 21426 1179
rect 21360 1099 21426 1115
rect 21360 1035 21361 1099
rect 21425 1035 21426 1099
rect 21360 1019 21426 1035
rect 21360 955 21361 1019
rect 21425 955 21426 1019
rect 21360 801 21426 955
rect 21486 863 21546 1893
rect 21606 801 21666 1833
rect 21726 863 21786 1893
rect 21846 801 21906 1833
rect 21966 1739 22032 1829
rect 21966 1675 21967 1739
rect 22031 1675 22032 1739
rect 21966 1659 22032 1675
rect 21966 1595 21967 1659
rect 22031 1595 22032 1659
rect 21966 1579 22032 1595
rect 21966 1515 21967 1579
rect 22031 1515 22032 1579
rect 21966 1499 22032 1515
rect 21966 1435 21967 1499
rect 22031 1435 22032 1499
rect 21966 1419 22032 1435
rect 21966 1355 21967 1419
rect 22031 1355 22032 1419
rect 21966 1339 22032 1355
rect 21966 1275 21967 1339
rect 22031 1275 22032 1339
rect 21966 1259 22032 1275
rect 21966 1195 21967 1259
rect 22031 1195 22032 1259
rect 21966 1179 22032 1195
rect 21966 1115 21967 1179
rect 22031 1115 22032 1179
rect 21966 1099 22032 1115
rect 21966 1035 21967 1099
rect 22031 1035 22032 1099
rect 21966 1019 22032 1035
rect 21966 955 21967 1019
rect 22031 955 22032 1019
rect 21966 801 22032 955
rect 22092 863 22152 1893
rect 22212 801 22272 1833
rect 22332 863 22392 1893
rect 22452 801 22512 1833
rect 22572 1739 22638 1829
rect 22572 1675 22573 1739
rect 22637 1675 22638 1739
rect 22572 1659 22638 1675
rect 22572 1595 22573 1659
rect 22637 1595 22638 1659
rect 22572 1579 22638 1595
rect 22572 1515 22573 1579
rect 22637 1515 22638 1579
rect 22572 1499 22638 1515
rect 22572 1435 22573 1499
rect 22637 1435 22638 1499
rect 22572 1419 22638 1435
rect 22572 1355 22573 1419
rect 22637 1355 22638 1419
rect 22572 1339 22638 1355
rect 22572 1275 22573 1339
rect 22637 1275 22638 1339
rect 22572 1259 22638 1275
rect 22572 1195 22573 1259
rect 22637 1195 22638 1259
rect 22572 1179 22638 1195
rect 22572 1115 22573 1179
rect 22637 1115 22638 1179
rect 22572 1099 22638 1115
rect 22572 1035 22573 1099
rect 22637 1035 22638 1099
rect 22572 1019 22638 1035
rect 22572 955 22573 1019
rect 22637 955 22638 1019
rect 22572 801 22638 955
rect 22698 863 22758 1893
rect 22818 801 22878 1833
rect 22938 863 22998 1893
rect 23058 801 23118 1833
rect 23178 1739 23244 1829
rect 23178 1675 23179 1739
rect 23243 1675 23244 1739
rect 23178 1659 23244 1675
rect 23178 1595 23179 1659
rect 23243 1595 23244 1659
rect 23178 1579 23244 1595
rect 23178 1515 23179 1579
rect 23243 1515 23244 1579
rect 23178 1499 23244 1515
rect 23178 1435 23179 1499
rect 23243 1435 23244 1499
rect 23178 1419 23244 1435
rect 23178 1355 23179 1419
rect 23243 1355 23244 1419
rect 23178 1339 23244 1355
rect 23178 1275 23179 1339
rect 23243 1275 23244 1339
rect 23178 1259 23244 1275
rect 23178 1195 23179 1259
rect 23243 1195 23244 1259
rect 23178 1179 23244 1195
rect 23178 1115 23179 1179
rect 23243 1115 23244 1179
rect 23178 1099 23244 1115
rect 23178 1035 23179 1099
rect 23243 1035 23244 1099
rect 23178 1019 23244 1035
rect 23178 955 23179 1019
rect 23243 955 23244 1019
rect 23178 801 23244 955
rect 23304 863 23364 1893
rect 23424 801 23484 1833
rect 23544 863 23604 1893
rect 23664 801 23724 1833
rect 23784 1739 23850 1829
rect 23784 1675 23785 1739
rect 23849 1675 23850 1739
rect 23784 1659 23850 1675
rect 23784 1595 23785 1659
rect 23849 1595 23850 1659
rect 23784 1579 23850 1595
rect 23784 1515 23785 1579
rect 23849 1515 23850 1579
rect 23784 1499 23850 1515
rect 23784 1435 23785 1499
rect 23849 1435 23850 1499
rect 23784 1419 23850 1435
rect 23784 1355 23785 1419
rect 23849 1355 23850 1419
rect 23784 1339 23850 1355
rect 23784 1275 23785 1339
rect 23849 1275 23850 1339
rect 23784 1259 23850 1275
rect 23784 1195 23785 1259
rect 23849 1195 23850 1259
rect 23784 1179 23850 1195
rect 23784 1115 23785 1179
rect 23849 1115 23850 1179
rect 23784 1099 23850 1115
rect 23784 1035 23785 1099
rect 23849 1035 23850 1099
rect 23784 1019 23850 1035
rect 23784 955 23785 1019
rect 23849 955 23850 1019
rect 23784 801 23850 955
rect 23910 863 23970 1893
rect 24030 801 24090 1833
rect 24150 863 24210 1893
rect 24270 801 24330 1833
rect 24390 1739 24456 1829
rect 24390 1675 24391 1739
rect 24455 1675 24456 1739
rect 24390 1659 24456 1675
rect 24390 1595 24391 1659
rect 24455 1595 24456 1659
rect 24390 1579 24456 1595
rect 24390 1515 24391 1579
rect 24455 1515 24456 1579
rect 24390 1499 24456 1515
rect 24390 1435 24391 1499
rect 24455 1435 24456 1499
rect 24390 1419 24456 1435
rect 24390 1355 24391 1419
rect 24455 1355 24456 1419
rect 24390 1339 24456 1355
rect 24390 1275 24391 1339
rect 24455 1275 24456 1339
rect 24390 1259 24456 1275
rect 24390 1195 24391 1259
rect 24455 1195 24456 1259
rect 24390 1179 24456 1195
rect 24390 1115 24391 1179
rect 24455 1115 24456 1179
rect 24390 1099 24456 1115
rect 24390 1035 24391 1099
rect 24455 1035 24456 1099
rect 24390 1019 24456 1035
rect 24390 955 24391 1019
rect 24455 955 24456 1019
rect 24390 801 24456 955
rect 24516 863 24576 1893
rect 24636 801 24696 1833
rect 24756 863 24816 1893
rect 24876 801 24936 1833
rect 24996 1739 25062 1829
rect 24996 1675 24997 1739
rect 25061 1675 25062 1739
rect 24996 1659 25062 1675
rect 24996 1595 24997 1659
rect 25061 1595 25062 1659
rect 24996 1579 25062 1595
rect 24996 1515 24997 1579
rect 25061 1515 25062 1579
rect 24996 1499 25062 1515
rect 24996 1435 24997 1499
rect 25061 1435 25062 1499
rect 24996 1419 25062 1435
rect 24996 1355 24997 1419
rect 25061 1355 25062 1419
rect 24996 1339 25062 1355
rect 24996 1275 24997 1339
rect 25061 1275 25062 1339
rect 24996 1259 25062 1275
rect 24996 1195 24997 1259
rect 25061 1195 25062 1259
rect 24996 1179 25062 1195
rect 24996 1115 24997 1179
rect 25061 1115 25062 1179
rect 24996 1099 25062 1115
rect 24996 1035 24997 1099
rect 25061 1035 25062 1099
rect 24996 1019 25062 1035
rect 24996 955 24997 1019
rect 25061 955 25062 1019
rect 24996 801 25062 955
rect 25122 863 25182 1893
rect 25242 801 25302 1833
rect 25362 863 25422 1893
rect 25482 801 25542 1833
rect 25602 1739 25668 1829
rect 25602 1675 25603 1739
rect 25667 1675 25668 1739
rect 25602 1659 25668 1675
rect 25602 1595 25603 1659
rect 25667 1595 25668 1659
rect 25602 1579 25668 1595
rect 25602 1515 25603 1579
rect 25667 1515 25668 1579
rect 25602 1499 25668 1515
rect 25602 1435 25603 1499
rect 25667 1435 25668 1499
rect 25602 1419 25668 1435
rect 25602 1355 25603 1419
rect 25667 1355 25668 1419
rect 25602 1339 25668 1355
rect 25602 1275 25603 1339
rect 25667 1275 25668 1339
rect 25602 1259 25668 1275
rect 25602 1195 25603 1259
rect 25667 1195 25668 1259
rect 25602 1179 25668 1195
rect 25602 1115 25603 1179
rect 25667 1115 25668 1179
rect 25602 1099 25668 1115
rect 25602 1035 25603 1099
rect 25667 1035 25668 1099
rect 25602 1019 25668 1035
rect 25602 955 25603 1019
rect 25667 955 25668 1019
rect 25602 801 25668 955
rect 25728 863 25788 1893
rect 25848 801 25908 1833
rect 25968 863 26028 1893
rect 26088 801 26148 1833
rect 26208 1739 26274 1829
rect 26208 1675 26209 1739
rect 26273 1675 26274 1739
rect 26208 1659 26274 1675
rect 26208 1595 26209 1659
rect 26273 1595 26274 1659
rect 26208 1579 26274 1595
rect 26208 1515 26209 1579
rect 26273 1515 26274 1579
rect 26208 1499 26274 1515
rect 26208 1435 26209 1499
rect 26273 1435 26274 1499
rect 26208 1419 26274 1435
rect 26208 1355 26209 1419
rect 26273 1355 26274 1419
rect 26208 1339 26274 1355
rect 26208 1275 26209 1339
rect 26273 1275 26274 1339
rect 26208 1259 26274 1275
rect 26208 1195 26209 1259
rect 26273 1195 26274 1259
rect 26208 1179 26274 1195
rect 26208 1115 26209 1179
rect 26273 1115 26274 1179
rect 26208 1099 26274 1115
rect 26208 1035 26209 1099
rect 26273 1035 26274 1099
rect 26208 1019 26274 1035
rect 26208 955 26209 1019
rect 26273 955 26274 1019
rect 26208 801 26274 955
rect 26334 863 26394 1893
rect 26454 801 26514 1833
rect 26574 863 26634 1893
rect 26694 801 26754 1833
rect 26814 1739 26880 1829
rect 26814 1675 26815 1739
rect 26879 1675 26880 1739
rect 26814 1659 26880 1675
rect 26814 1595 26815 1659
rect 26879 1595 26880 1659
rect 26814 1579 26880 1595
rect 26814 1515 26815 1579
rect 26879 1515 26880 1579
rect 26814 1499 26880 1515
rect 26814 1435 26815 1499
rect 26879 1435 26880 1499
rect 26814 1419 26880 1435
rect 26814 1355 26815 1419
rect 26879 1355 26880 1419
rect 26814 1339 26880 1355
rect 26814 1275 26815 1339
rect 26879 1275 26880 1339
rect 26814 1259 26880 1275
rect 26814 1195 26815 1259
rect 26879 1195 26880 1259
rect 26814 1179 26880 1195
rect 26814 1115 26815 1179
rect 26879 1115 26880 1179
rect 26814 1099 26880 1115
rect 26814 1035 26815 1099
rect 26879 1035 26880 1099
rect 26814 1019 26880 1035
rect 26814 955 26815 1019
rect 26879 955 26880 1019
rect 26814 801 26880 955
rect 26940 863 27000 1893
rect 27060 801 27120 1833
rect 27180 863 27240 1893
rect 27300 801 27360 1833
rect 27420 1739 27486 1829
rect 27420 1675 27421 1739
rect 27485 1675 27486 1739
rect 27420 1659 27486 1675
rect 27420 1595 27421 1659
rect 27485 1595 27486 1659
rect 27420 1579 27486 1595
rect 27420 1515 27421 1579
rect 27485 1515 27486 1579
rect 27420 1499 27486 1515
rect 27420 1435 27421 1499
rect 27485 1435 27486 1499
rect 27420 1419 27486 1435
rect 27420 1355 27421 1419
rect 27485 1355 27486 1419
rect 27420 1339 27486 1355
rect 27420 1275 27421 1339
rect 27485 1275 27486 1339
rect 27420 1259 27486 1275
rect 27420 1195 27421 1259
rect 27485 1195 27486 1259
rect 27420 1179 27486 1195
rect 27420 1115 27421 1179
rect 27485 1115 27486 1179
rect 27420 1099 27486 1115
rect 27420 1035 27421 1099
rect 27485 1035 27486 1099
rect 27420 1019 27486 1035
rect 27420 955 27421 1019
rect 27485 955 27486 1019
rect 27420 801 27486 955
rect 27546 863 27606 1893
rect 27666 801 27726 1833
rect 27786 863 27846 1893
rect 27906 801 27966 1833
rect 28026 1739 28092 1829
rect 28026 1675 28027 1739
rect 28091 1675 28092 1739
rect 28026 1659 28092 1675
rect 28026 1595 28027 1659
rect 28091 1595 28092 1659
rect 28026 1579 28092 1595
rect 28026 1515 28027 1579
rect 28091 1515 28092 1579
rect 28026 1499 28092 1515
rect 28026 1435 28027 1499
rect 28091 1435 28092 1499
rect 28026 1419 28092 1435
rect 28026 1355 28027 1419
rect 28091 1355 28092 1419
rect 28026 1339 28092 1355
rect 28026 1275 28027 1339
rect 28091 1275 28092 1339
rect 28026 1259 28092 1275
rect 28026 1195 28027 1259
rect 28091 1195 28092 1259
rect 28026 1179 28092 1195
rect 28026 1115 28027 1179
rect 28091 1115 28092 1179
rect 28026 1099 28092 1115
rect 28026 1035 28027 1099
rect 28091 1035 28092 1099
rect 28026 1019 28092 1035
rect 28026 955 28027 1019
rect 28091 955 28092 1019
rect 28026 801 28092 955
rect 28152 863 28212 1893
rect 28272 801 28332 1833
rect 28392 863 28452 1893
rect 28512 801 28572 1833
rect 28632 1739 28698 1829
rect 28632 1675 28633 1739
rect 28697 1675 28698 1739
rect 28632 1659 28698 1675
rect 28632 1595 28633 1659
rect 28697 1595 28698 1659
rect 28632 1579 28698 1595
rect 28632 1515 28633 1579
rect 28697 1515 28698 1579
rect 28632 1499 28698 1515
rect 28632 1435 28633 1499
rect 28697 1435 28698 1499
rect 28632 1419 28698 1435
rect 28632 1355 28633 1419
rect 28697 1355 28698 1419
rect 28632 1339 28698 1355
rect 28632 1275 28633 1339
rect 28697 1275 28698 1339
rect 28632 1259 28698 1275
rect 28632 1195 28633 1259
rect 28697 1195 28698 1259
rect 28632 1179 28698 1195
rect 28632 1115 28633 1179
rect 28697 1115 28698 1179
rect 28632 1099 28698 1115
rect 28632 1035 28633 1099
rect 28697 1035 28698 1099
rect 28632 1019 28698 1035
rect 28632 955 28633 1019
rect 28697 955 28698 1019
rect 28632 801 28698 955
rect 28758 863 28818 1893
rect 28878 801 28938 1833
rect 28998 863 29058 1893
rect 29118 801 29178 1833
rect 29238 1739 29304 1829
rect 29238 1675 29239 1739
rect 29303 1675 29304 1739
rect 29238 1659 29304 1675
rect 29238 1595 29239 1659
rect 29303 1595 29304 1659
rect 29238 1579 29304 1595
rect 29238 1515 29239 1579
rect 29303 1515 29304 1579
rect 29238 1499 29304 1515
rect 29238 1435 29239 1499
rect 29303 1435 29304 1499
rect 29238 1419 29304 1435
rect 29238 1355 29239 1419
rect 29303 1355 29304 1419
rect 29238 1339 29304 1355
rect 29238 1275 29239 1339
rect 29303 1275 29304 1339
rect 29238 1259 29304 1275
rect 29238 1195 29239 1259
rect 29303 1195 29304 1259
rect 29238 1179 29304 1195
rect 29238 1115 29239 1179
rect 29303 1115 29304 1179
rect 29238 1099 29304 1115
rect 29238 1035 29239 1099
rect 29303 1035 29304 1099
rect 29238 1019 29304 1035
rect 29238 955 29239 1019
rect 29303 955 29304 1019
rect 29238 801 29304 955
rect 29364 863 29424 1893
rect 29484 801 29544 1833
rect 29604 863 29664 1893
rect 29724 801 29784 1833
rect 29844 1739 29910 1829
rect 29844 1675 29845 1739
rect 29909 1675 29910 1739
rect 29844 1659 29910 1675
rect 29844 1595 29845 1659
rect 29909 1595 29910 1659
rect 29844 1579 29910 1595
rect 29844 1515 29845 1579
rect 29909 1515 29910 1579
rect 29844 1499 29910 1515
rect 29844 1435 29845 1499
rect 29909 1435 29910 1499
rect 29844 1419 29910 1435
rect 29844 1355 29845 1419
rect 29909 1355 29910 1419
rect 29844 1339 29910 1355
rect 29844 1275 29845 1339
rect 29909 1275 29910 1339
rect 29844 1259 29910 1275
rect 29844 1195 29845 1259
rect 29909 1195 29910 1259
rect 29844 1179 29910 1195
rect 29844 1115 29845 1179
rect 29909 1115 29910 1179
rect 29844 1099 29910 1115
rect 29844 1035 29845 1099
rect 29909 1035 29910 1099
rect 29844 1019 29910 1035
rect 29844 955 29845 1019
rect 29909 955 29910 1019
rect 29844 801 29910 955
rect 29970 863 30030 1893
rect 30090 801 30150 1833
rect 30210 863 30270 1893
rect 30330 801 30390 1833
rect 30450 1739 30516 1829
rect 30450 1675 30451 1739
rect 30515 1675 30516 1739
rect 30450 1659 30516 1675
rect 30450 1595 30451 1659
rect 30515 1595 30516 1659
rect 30450 1579 30516 1595
rect 30450 1515 30451 1579
rect 30515 1515 30516 1579
rect 30450 1499 30516 1515
rect 30450 1435 30451 1499
rect 30515 1435 30516 1499
rect 30450 1419 30516 1435
rect 30450 1355 30451 1419
rect 30515 1355 30516 1419
rect 30450 1339 30516 1355
rect 30450 1275 30451 1339
rect 30515 1275 30516 1339
rect 30450 1259 30516 1275
rect 30450 1195 30451 1259
rect 30515 1195 30516 1259
rect 30450 1179 30516 1195
rect 30450 1115 30451 1179
rect 30515 1115 30516 1179
rect 30450 1099 30516 1115
rect 30450 1035 30451 1099
rect 30515 1035 30516 1099
rect 30450 1019 30516 1035
rect 30450 955 30451 1019
rect 30515 955 30516 1019
rect 30450 801 30516 955
rect 30576 863 30636 1893
rect 30696 801 30756 1833
rect 30816 863 30876 1893
rect 30936 801 30996 1833
rect 31056 1739 31122 1829
rect 31056 1675 31057 1739
rect 31121 1675 31122 1739
rect 31056 1659 31122 1675
rect 31056 1595 31057 1659
rect 31121 1595 31122 1659
rect 31056 1579 31122 1595
rect 31056 1515 31057 1579
rect 31121 1515 31122 1579
rect 31056 1499 31122 1515
rect 31056 1435 31057 1499
rect 31121 1435 31122 1499
rect 31056 1419 31122 1435
rect 31056 1355 31057 1419
rect 31121 1355 31122 1419
rect 31056 1339 31122 1355
rect 31056 1275 31057 1339
rect 31121 1275 31122 1339
rect 31056 1259 31122 1275
rect 31056 1195 31057 1259
rect 31121 1195 31122 1259
rect 31056 1179 31122 1195
rect 31056 1115 31057 1179
rect 31121 1115 31122 1179
rect 31056 1099 31122 1115
rect 31056 1035 31057 1099
rect 31121 1035 31122 1099
rect 31056 1019 31122 1035
rect 31056 955 31057 1019
rect 31121 955 31122 1019
rect 31056 801 31122 955
rect 31182 863 31242 1893
rect 31302 801 31362 1833
rect 31422 863 31482 1893
rect 31542 801 31602 1833
rect 31662 1739 31728 1829
rect 31662 1675 31663 1739
rect 31727 1675 31728 1739
rect 31662 1659 31728 1675
rect 31662 1595 31663 1659
rect 31727 1595 31728 1659
rect 31662 1579 31728 1595
rect 31662 1515 31663 1579
rect 31727 1515 31728 1579
rect 31662 1499 31728 1515
rect 31662 1435 31663 1499
rect 31727 1435 31728 1499
rect 31662 1419 31728 1435
rect 31662 1355 31663 1419
rect 31727 1355 31728 1419
rect 31662 1339 31728 1355
rect 31662 1275 31663 1339
rect 31727 1275 31728 1339
rect 31662 1259 31728 1275
rect 31662 1195 31663 1259
rect 31727 1195 31728 1259
rect 31662 1179 31728 1195
rect 31662 1115 31663 1179
rect 31727 1115 31728 1179
rect 31662 1099 31728 1115
rect 31662 1035 31663 1099
rect 31727 1035 31728 1099
rect 31662 1019 31728 1035
rect 31662 955 31663 1019
rect 31727 955 31728 1019
rect 31662 801 31728 955
rect 31788 863 31848 1893
rect 31908 801 31968 1833
rect 32028 863 32088 1893
rect 32148 801 32208 1833
rect 32268 1739 32334 1829
rect 32268 1675 32269 1739
rect 32333 1675 32334 1739
rect 32268 1659 32334 1675
rect 32268 1595 32269 1659
rect 32333 1595 32334 1659
rect 32268 1579 32334 1595
rect 32268 1515 32269 1579
rect 32333 1515 32334 1579
rect 32268 1499 32334 1515
rect 32268 1435 32269 1499
rect 32333 1435 32334 1499
rect 32268 1419 32334 1435
rect 32268 1355 32269 1419
rect 32333 1355 32334 1419
rect 32268 1339 32334 1355
rect 32268 1275 32269 1339
rect 32333 1275 32334 1339
rect 32268 1259 32334 1275
rect 32268 1195 32269 1259
rect 32333 1195 32334 1259
rect 32268 1179 32334 1195
rect 32268 1115 32269 1179
rect 32333 1115 32334 1179
rect 32268 1099 32334 1115
rect 32268 1035 32269 1099
rect 32333 1035 32334 1099
rect 32268 1019 32334 1035
rect 32268 955 32269 1019
rect 32333 955 32334 1019
rect 32268 801 32334 955
rect 32394 863 32454 1893
rect 32514 801 32574 1833
rect 32634 863 32694 1893
rect 32754 801 32814 1833
rect 32874 1739 32940 1829
rect 32874 1675 32875 1739
rect 32939 1675 32940 1739
rect 32874 1659 32940 1675
rect 32874 1595 32875 1659
rect 32939 1595 32940 1659
rect 32874 1579 32940 1595
rect 32874 1515 32875 1579
rect 32939 1515 32940 1579
rect 32874 1499 32940 1515
rect 32874 1435 32875 1499
rect 32939 1435 32940 1499
rect 32874 1419 32940 1435
rect 32874 1355 32875 1419
rect 32939 1355 32940 1419
rect 32874 1339 32940 1355
rect 32874 1275 32875 1339
rect 32939 1275 32940 1339
rect 32874 1259 32940 1275
rect 32874 1195 32875 1259
rect 32939 1195 32940 1259
rect 32874 1179 32940 1195
rect 32874 1115 32875 1179
rect 32939 1115 32940 1179
rect 32874 1099 32940 1115
rect 32874 1035 32875 1099
rect 32939 1035 32940 1099
rect 32874 1019 32940 1035
rect 32874 955 32875 1019
rect 32939 955 32940 1019
rect 32874 801 32940 955
rect 33000 863 33060 1893
rect 33120 801 33180 1833
rect 33240 863 33300 1893
rect 33360 801 33420 1833
rect 33480 1739 33546 1829
rect 33480 1675 33481 1739
rect 33545 1675 33546 1739
rect 33480 1659 33546 1675
rect 33480 1595 33481 1659
rect 33545 1595 33546 1659
rect 33480 1579 33546 1595
rect 33480 1515 33481 1579
rect 33545 1515 33546 1579
rect 33480 1499 33546 1515
rect 33480 1435 33481 1499
rect 33545 1435 33546 1499
rect 33480 1419 33546 1435
rect 33480 1355 33481 1419
rect 33545 1355 33546 1419
rect 33480 1339 33546 1355
rect 33480 1275 33481 1339
rect 33545 1275 33546 1339
rect 33480 1259 33546 1275
rect 33480 1195 33481 1259
rect 33545 1195 33546 1259
rect 33480 1179 33546 1195
rect 33480 1115 33481 1179
rect 33545 1115 33546 1179
rect 33480 1099 33546 1115
rect 33480 1035 33481 1099
rect 33545 1035 33546 1099
rect 33480 1019 33546 1035
rect 33480 955 33481 1019
rect 33545 955 33546 1019
rect 33480 801 33546 955
rect 33606 863 33666 1893
rect 33726 801 33786 1833
rect 33846 863 33906 1893
rect 33966 801 34026 1833
rect 34086 1739 34152 1829
rect 34086 1675 34087 1739
rect 34151 1675 34152 1739
rect 34086 1659 34152 1675
rect 34086 1595 34087 1659
rect 34151 1595 34152 1659
rect 34086 1579 34152 1595
rect 34086 1515 34087 1579
rect 34151 1515 34152 1579
rect 34086 1499 34152 1515
rect 34086 1435 34087 1499
rect 34151 1435 34152 1499
rect 34086 1419 34152 1435
rect 34086 1355 34087 1419
rect 34151 1355 34152 1419
rect 34086 1339 34152 1355
rect 34086 1275 34087 1339
rect 34151 1275 34152 1339
rect 34086 1259 34152 1275
rect 34086 1195 34087 1259
rect 34151 1195 34152 1259
rect 34086 1179 34152 1195
rect 34086 1115 34087 1179
rect 34151 1115 34152 1179
rect 34086 1099 34152 1115
rect 34086 1035 34087 1099
rect 34151 1035 34152 1099
rect 34086 1019 34152 1035
rect 34086 955 34087 1019
rect 34151 955 34152 1019
rect 34086 801 34152 955
rect 34212 863 34272 1893
rect 34332 801 34392 1833
rect 34452 863 34512 1893
rect 34572 801 34632 1833
rect 34692 1739 34758 1829
rect 34692 1675 34693 1739
rect 34757 1675 34758 1739
rect 34692 1659 34758 1675
rect 34692 1595 34693 1659
rect 34757 1595 34758 1659
rect 34692 1579 34758 1595
rect 34692 1515 34693 1579
rect 34757 1515 34758 1579
rect 34692 1499 34758 1515
rect 34692 1435 34693 1499
rect 34757 1435 34758 1499
rect 34692 1419 34758 1435
rect 34692 1355 34693 1419
rect 34757 1355 34758 1419
rect 34692 1339 34758 1355
rect 34692 1275 34693 1339
rect 34757 1275 34758 1339
rect 34692 1259 34758 1275
rect 34692 1195 34693 1259
rect 34757 1195 34758 1259
rect 34692 1179 34758 1195
rect 34692 1115 34693 1179
rect 34757 1115 34758 1179
rect 34692 1099 34758 1115
rect 34692 1035 34693 1099
rect 34757 1035 34758 1099
rect 34692 1019 34758 1035
rect 34692 955 34693 1019
rect 34757 955 34758 1019
rect 34692 801 34758 955
rect 34818 863 34878 1893
rect 34938 801 34998 1833
rect 35058 863 35118 1893
rect 35178 801 35238 1833
rect 35298 1739 35364 1829
rect 35298 1675 35299 1739
rect 35363 1675 35364 1739
rect 35298 1659 35364 1675
rect 35298 1595 35299 1659
rect 35363 1595 35364 1659
rect 35298 1579 35364 1595
rect 35298 1515 35299 1579
rect 35363 1515 35364 1579
rect 35298 1499 35364 1515
rect 35298 1435 35299 1499
rect 35363 1435 35364 1499
rect 35298 1419 35364 1435
rect 35298 1355 35299 1419
rect 35363 1355 35364 1419
rect 35298 1339 35364 1355
rect 35298 1275 35299 1339
rect 35363 1275 35364 1339
rect 35298 1259 35364 1275
rect 35298 1195 35299 1259
rect 35363 1195 35364 1259
rect 35298 1179 35364 1195
rect 35298 1115 35299 1179
rect 35363 1115 35364 1179
rect 35298 1099 35364 1115
rect 35298 1035 35299 1099
rect 35363 1035 35364 1099
rect 35298 1019 35364 1035
rect 35298 955 35299 1019
rect 35363 955 35364 1019
rect 35298 801 35364 955
rect 35424 863 35484 1893
rect 35544 801 35604 1833
rect 35664 863 35724 1893
rect 35784 801 35844 1833
rect 35904 1739 35970 1829
rect 35904 1675 35905 1739
rect 35969 1675 35970 1739
rect 35904 1659 35970 1675
rect 35904 1595 35905 1659
rect 35969 1595 35970 1659
rect 35904 1579 35970 1595
rect 35904 1515 35905 1579
rect 35969 1515 35970 1579
rect 35904 1499 35970 1515
rect 35904 1435 35905 1499
rect 35969 1435 35970 1499
rect 35904 1419 35970 1435
rect 35904 1355 35905 1419
rect 35969 1355 35970 1419
rect 35904 1339 35970 1355
rect 35904 1275 35905 1339
rect 35969 1275 35970 1339
rect 35904 1259 35970 1275
rect 35904 1195 35905 1259
rect 35969 1195 35970 1259
rect 35904 1179 35970 1195
rect 35904 1115 35905 1179
rect 35969 1115 35970 1179
rect 35904 1099 35970 1115
rect 35904 1035 35905 1099
rect 35969 1035 35970 1099
rect 35904 1019 35970 1035
rect 35904 955 35905 1019
rect 35969 955 35970 1019
rect 35904 801 35970 955
rect 36030 863 36090 1893
rect 36150 801 36210 1833
rect 36270 863 36330 1893
rect 36390 801 36450 1833
rect 36510 1739 36576 1829
rect 36510 1675 36511 1739
rect 36575 1675 36576 1739
rect 36510 1659 36576 1675
rect 36510 1595 36511 1659
rect 36575 1595 36576 1659
rect 36510 1579 36576 1595
rect 36510 1515 36511 1579
rect 36575 1515 36576 1579
rect 36510 1499 36576 1515
rect 36510 1435 36511 1499
rect 36575 1435 36576 1499
rect 36510 1419 36576 1435
rect 36510 1355 36511 1419
rect 36575 1355 36576 1419
rect 36510 1339 36576 1355
rect 36510 1275 36511 1339
rect 36575 1275 36576 1339
rect 36510 1259 36576 1275
rect 36510 1195 36511 1259
rect 36575 1195 36576 1259
rect 36510 1179 36576 1195
rect 36510 1115 36511 1179
rect 36575 1115 36576 1179
rect 36510 1099 36576 1115
rect 36510 1035 36511 1099
rect 36575 1035 36576 1099
rect 36510 1019 36576 1035
rect 36510 955 36511 1019
rect 36575 955 36576 1019
rect 36510 801 36576 955
rect 36636 863 36696 1893
rect 36756 801 36816 1833
rect 36876 863 36936 1893
rect 36996 801 37056 1833
rect 37116 1739 37182 1829
rect 37116 1675 37117 1739
rect 37181 1675 37182 1739
rect 37116 1659 37182 1675
rect 37116 1595 37117 1659
rect 37181 1595 37182 1659
rect 37116 1579 37182 1595
rect 37116 1515 37117 1579
rect 37181 1515 37182 1579
rect 37116 1499 37182 1515
rect 37116 1435 37117 1499
rect 37181 1435 37182 1499
rect 37116 1419 37182 1435
rect 37116 1355 37117 1419
rect 37181 1355 37182 1419
rect 37116 1339 37182 1355
rect 37116 1275 37117 1339
rect 37181 1275 37182 1339
rect 37116 1259 37182 1275
rect 37116 1195 37117 1259
rect 37181 1195 37182 1259
rect 37116 1179 37182 1195
rect 37116 1115 37117 1179
rect 37181 1115 37182 1179
rect 37116 1099 37182 1115
rect 37116 1035 37117 1099
rect 37181 1035 37182 1099
rect 37116 1019 37182 1035
rect 37116 955 37117 1019
rect 37181 955 37182 1019
rect 37116 801 37182 955
rect 37242 863 37302 1893
rect 37362 801 37422 1833
rect 37482 863 37542 1893
rect 37602 801 37662 1833
rect 37722 1739 37788 1829
rect 37722 1675 37723 1739
rect 37787 1675 37788 1739
rect 37722 1659 37788 1675
rect 37722 1595 37723 1659
rect 37787 1595 37788 1659
rect 37722 1579 37788 1595
rect 37722 1515 37723 1579
rect 37787 1515 37788 1579
rect 37722 1499 37788 1515
rect 37722 1435 37723 1499
rect 37787 1435 37788 1499
rect 37722 1419 37788 1435
rect 37722 1355 37723 1419
rect 37787 1355 37788 1419
rect 37722 1339 37788 1355
rect 37722 1275 37723 1339
rect 37787 1275 37788 1339
rect 37722 1259 37788 1275
rect 37722 1195 37723 1259
rect 37787 1195 37788 1259
rect 37722 1179 37788 1195
rect 37722 1115 37723 1179
rect 37787 1115 37788 1179
rect 37722 1099 37788 1115
rect 37722 1035 37723 1099
rect 37787 1035 37788 1099
rect 37722 1019 37788 1035
rect 37722 955 37723 1019
rect 37787 955 37788 1019
rect 37722 801 37788 955
rect 37848 863 37908 1893
rect 37968 801 38028 1833
rect 38088 863 38148 1893
rect 38208 801 38268 1833
rect 38328 1739 38394 1829
rect 38328 1675 38329 1739
rect 38393 1675 38394 1739
rect 38328 1659 38394 1675
rect 38328 1595 38329 1659
rect 38393 1595 38394 1659
rect 38328 1579 38394 1595
rect 38328 1515 38329 1579
rect 38393 1515 38394 1579
rect 38328 1499 38394 1515
rect 38328 1435 38329 1499
rect 38393 1435 38394 1499
rect 38328 1419 38394 1435
rect 38328 1355 38329 1419
rect 38393 1355 38394 1419
rect 38328 1339 38394 1355
rect 38328 1275 38329 1339
rect 38393 1275 38394 1339
rect 38328 1259 38394 1275
rect 38328 1195 38329 1259
rect 38393 1195 38394 1259
rect 38328 1179 38394 1195
rect 38328 1115 38329 1179
rect 38393 1115 38394 1179
rect 38328 1099 38394 1115
rect 38328 1035 38329 1099
rect 38393 1035 38394 1099
rect 38328 1019 38394 1035
rect 38328 955 38329 1019
rect 38393 955 38394 1019
rect 38328 801 38394 955
rect 38454 863 38514 1893
rect 38574 801 38634 1833
rect 38694 863 38754 1893
rect 38814 801 38874 1833
rect 38934 1739 39000 1829
rect 38934 1675 38935 1739
rect 38999 1675 39000 1739
rect 38934 1659 39000 1675
rect 38934 1595 38935 1659
rect 38999 1595 39000 1659
rect 38934 1579 39000 1595
rect 38934 1515 38935 1579
rect 38999 1515 39000 1579
rect 38934 1499 39000 1515
rect 38934 1435 38935 1499
rect 38999 1435 39000 1499
rect 38934 1419 39000 1435
rect 38934 1355 38935 1419
rect 38999 1355 39000 1419
rect 38934 1339 39000 1355
rect 38934 1275 38935 1339
rect 38999 1275 39000 1339
rect 38934 1259 39000 1275
rect 38934 1195 38935 1259
rect 38999 1195 39000 1259
rect 38934 1179 39000 1195
rect 38934 1115 38935 1179
rect 38999 1115 39000 1179
rect 38934 1099 39000 1115
rect 38934 1035 38935 1099
rect 38999 1035 39000 1099
rect 38934 1019 39000 1035
rect 38934 955 38935 1019
rect 38999 955 39000 1019
rect 38934 801 39000 955
rect 39060 863 39120 1893
rect 39180 801 39240 1833
rect 39300 863 39360 1893
rect 39420 801 39480 1833
rect 39540 1739 39606 1829
rect 39540 1675 39541 1739
rect 39605 1675 39606 1739
rect 39540 1659 39606 1675
rect 39540 1595 39541 1659
rect 39605 1595 39606 1659
rect 39540 1579 39606 1595
rect 39540 1515 39541 1579
rect 39605 1515 39606 1579
rect 39540 1499 39606 1515
rect 39540 1435 39541 1499
rect 39605 1435 39606 1499
rect 39540 1419 39606 1435
rect 39540 1355 39541 1419
rect 39605 1355 39606 1419
rect 39540 1339 39606 1355
rect 39540 1275 39541 1339
rect 39605 1275 39606 1339
rect 39540 1259 39606 1275
rect 39540 1195 39541 1259
rect 39605 1195 39606 1259
rect 39540 1179 39606 1195
rect 39540 1115 39541 1179
rect 39605 1115 39606 1179
rect 39540 1099 39606 1115
rect 39540 1035 39541 1099
rect 39605 1035 39606 1099
rect 39540 1019 39606 1035
rect 39540 955 39541 1019
rect 39605 955 39606 1019
rect 39540 801 39606 955
rect 20148 799 39606 801
rect 20148 735 20252 799
rect 20316 735 20332 799
rect 20396 735 20412 799
rect 20476 735 20492 799
rect 20556 735 20572 799
rect 20636 735 20652 799
rect 20716 735 20858 799
rect 20922 735 20938 799
rect 21002 735 21018 799
rect 21082 735 21098 799
rect 21162 735 21178 799
rect 21242 735 21258 799
rect 21322 735 21464 799
rect 21528 735 21544 799
rect 21608 735 21624 799
rect 21688 735 21704 799
rect 21768 735 21784 799
rect 21848 735 21864 799
rect 21928 735 22070 799
rect 22134 735 22150 799
rect 22214 735 22230 799
rect 22294 735 22310 799
rect 22374 735 22390 799
rect 22454 735 22470 799
rect 22534 735 22676 799
rect 22740 735 22756 799
rect 22820 735 22836 799
rect 22900 735 22916 799
rect 22980 735 22996 799
rect 23060 735 23076 799
rect 23140 735 23282 799
rect 23346 735 23362 799
rect 23426 735 23442 799
rect 23506 735 23522 799
rect 23586 735 23602 799
rect 23666 735 23682 799
rect 23746 735 23888 799
rect 23952 735 23968 799
rect 24032 735 24048 799
rect 24112 735 24128 799
rect 24192 735 24208 799
rect 24272 735 24288 799
rect 24352 735 24494 799
rect 24558 735 24574 799
rect 24638 735 24654 799
rect 24718 735 24734 799
rect 24798 735 24814 799
rect 24878 735 24894 799
rect 24958 735 25100 799
rect 25164 735 25180 799
rect 25244 735 25260 799
rect 25324 735 25340 799
rect 25404 735 25420 799
rect 25484 735 25500 799
rect 25564 735 25706 799
rect 25770 735 25786 799
rect 25850 735 25866 799
rect 25930 735 25946 799
rect 26010 735 26026 799
rect 26090 735 26106 799
rect 26170 735 26312 799
rect 26376 735 26392 799
rect 26456 735 26472 799
rect 26536 735 26552 799
rect 26616 735 26632 799
rect 26696 735 26712 799
rect 26776 735 26918 799
rect 26982 735 26998 799
rect 27062 735 27078 799
rect 27142 735 27158 799
rect 27222 735 27238 799
rect 27302 735 27318 799
rect 27382 735 27524 799
rect 27588 735 27604 799
rect 27668 735 27684 799
rect 27748 735 27764 799
rect 27828 735 27844 799
rect 27908 735 27924 799
rect 27988 735 28130 799
rect 28194 735 28210 799
rect 28274 735 28290 799
rect 28354 735 28370 799
rect 28434 735 28450 799
rect 28514 735 28530 799
rect 28594 735 28736 799
rect 28800 735 28816 799
rect 28880 735 28896 799
rect 28960 735 28976 799
rect 29040 735 29056 799
rect 29120 735 29136 799
rect 29200 735 29342 799
rect 29406 735 29422 799
rect 29486 735 29502 799
rect 29566 735 29582 799
rect 29646 735 29662 799
rect 29726 735 29742 799
rect 29806 735 29948 799
rect 30012 735 30028 799
rect 30092 735 30108 799
rect 30172 735 30188 799
rect 30252 735 30268 799
rect 30332 735 30348 799
rect 30412 735 30554 799
rect 30618 735 30634 799
rect 30698 735 30714 799
rect 30778 735 30794 799
rect 30858 735 30874 799
rect 30938 735 30954 799
rect 31018 735 31160 799
rect 31224 735 31240 799
rect 31304 735 31320 799
rect 31384 735 31400 799
rect 31464 735 31480 799
rect 31544 735 31560 799
rect 31624 735 31766 799
rect 31830 735 31846 799
rect 31910 735 31926 799
rect 31990 735 32006 799
rect 32070 735 32086 799
rect 32150 735 32166 799
rect 32230 735 32372 799
rect 32436 735 32452 799
rect 32516 735 32532 799
rect 32596 735 32612 799
rect 32676 735 32692 799
rect 32756 735 32772 799
rect 32836 735 32978 799
rect 33042 735 33058 799
rect 33122 735 33138 799
rect 33202 735 33218 799
rect 33282 735 33298 799
rect 33362 735 33378 799
rect 33442 735 33584 799
rect 33648 735 33664 799
rect 33728 735 33744 799
rect 33808 735 33824 799
rect 33888 735 33904 799
rect 33968 735 33984 799
rect 34048 735 34190 799
rect 34254 735 34270 799
rect 34334 735 34350 799
rect 34414 735 34430 799
rect 34494 735 34510 799
rect 34574 735 34590 799
rect 34654 735 34796 799
rect 34860 735 34876 799
rect 34940 735 34956 799
rect 35020 735 35036 799
rect 35100 735 35116 799
rect 35180 735 35196 799
rect 35260 735 35402 799
rect 35466 735 35482 799
rect 35546 735 35562 799
rect 35626 735 35642 799
rect 35706 735 35722 799
rect 35786 735 35802 799
rect 35866 735 36008 799
rect 36072 735 36088 799
rect 36152 735 36168 799
rect 36232 735 36248 799
rect 36312 735 36328 799
rect 36392 735 36408 799
rect 36472 735 36614 799
rect 36678 735 36694 799
rect 36758 735 36774 799
rect 36838 735 36854 799
rect 36918 735 36934 799
rect 36998 735 37014 799
rect 37078 735 37220 799
rect 37284 735 37300 799
rect 37364 735 37380 799
rect 37444 735 37460 799
rect 37524 735 37540 799
rect 37604 735 37620 799
rect 37684 735 37826 799
rect 37890 735 37906 799
rect 37970 735 37986 799
rect 38050 735 38066 799
rect 38130 735 38146 799
rect 38210 735 38226 799
rect 38290 735 38432 799
rect 38496 735 38512 799
rect 38576 735 38592 799
rect 38656 735 38672 799
rect 38736 735 38752 799
rect 38816 735 38832 799
rect 38896 735 39038 799
rect 39102 735 39118 799
rect 39182 735 39198 799
rect 39262 735 39278 799
rect 39342 735 39358 799
rect 39422 735 39438 799
rect 39502 735 39606 799
rect 20148 733 39606 735
rect 20148 579 20214 733
rect 20148 515 20149 579
rect 20213 515 20214 579
rect 20148 499 20214 515
rect 20148 435 20149 499
rect 20213 435 20214 499
rect 20148 419 20214 435
rect 20148 355 20149 419
rect 20213 355 20214 419
rect 20148 339 20214 355
rect 20148 275 20149 339
rect 20213 275 20214 339
rect 20148 259 20214 275
rect 20148 195 20149 259
rect 20213 195 20214 259
rect 20148 179 20214 195
rect 20148 115 20149 179
rect 20213 115 20214 179
rect 20148 99 20214 115
rect 20148 35 20149 99
rect 20213 35 20214 99
rect 20148 19 20214 35
rect 20148 -45 20149 19
rect 20213 -45 20214 19
rect 20148 -61 20214 -45
rect 20148 -125 20149 -61
rect 20213 -125 20214 -61
rect 20148 -141 20214 -125
rect 20148 -205 20149 -141
rect 20213 -205 20214 -141
rect 20148 -295 20214 -205
rect 20274 -299 20334 733
rect 20394 -359 20454 671
rect 20514 -299 20574 733
rect 20634 -359 20694 671
rect 20754 579 20820 733
rect 20754 515 20755 579
rect 20819 515 20820 579
rect 20754 499 20820 515
rect 20754 435 20755 499
rect 20819 435 20820 499
rect 20754 419 20820 435
rect 20754 355 20755 419
rect 20819 355 20820 419
rect 20754 339 20820 355
rect 20754 275 20755 339
rect 20819 275 20820 339
rect 20754 259 20820 275
rect 20754 195 20755 259
rect 20819 195 20820 259
rect 20754 179 20820 195
rect 20754 115 20755 179
rect 20819 115 20820 179
rect 20754 99 20820 115
rect 20754 35 20755 99
rect 20819 35 20820 99
rect 20754 19 20820 35
rect 20754 -45 20755 19
rect 20819 -45 20820 19
rect 20754 -61 20820 -45
rect 20754 -125 20755 -61
rect 20819 -125 20820 -61
rect 20754 -141 20820 -125
rect 20754 -205 20755 -141
rect 20819 -205 20820 -141
rect 20754 -295 20820 -205
rect 20880 -299 20940 733
rect 21000 -359 21060 671
rect 21120 -299 21180 733
rect 21240 -359 21300 671
rect 21360 579 21426 733
rect 21360 515 21361 579
rect 21425 515 21426 579
rect 21360 499 21426 515
rect 21360 435 21361 499
rect 21425 435 21426 499
rect 21360 419 21426 435
rect 21360 355 21361 419
rect 21425 355 21426 419
rect 21360 339 21426 355
rect 21360 275 21361 339
rect 21425 275 21426 339
rect 21360 259 21426 275
rect 21360 195 21361 259
rect 21425 195 21426 259
rect 21360 179 21426 195
rect 21360 115 21361 179
rect 21425 115 21426 179
rect 21360 99 21426 115
rect 21360 35 21361 99
rect 21425 35 21426 99
rect 21360 19 21426 35
rect 21360 -45 21361 19
rect 21425 -45 21426 19
rect 21360 -61 21426 -45
rect 21360 -125 21361 -61
rect 21425 -125 21426 -61
rect 21360 -141 21426 -125
rect 21360 -205 21361 -141
rect 21425 -205 21426 -141
rect 21360 -295 21426 -205
rect 21486 -299 21546 733
rect 21606 -359 21666 671
rect 21726 -299 21786 733
rect 21846 -359 21906 671
rect 21966 579 22032 733
rect 21966 515 21967 579
rect 22031 515 22032 579
rect 21966 499 22032 515
rect 21966 435 21967 499
rect 22031 435 22032 499
rect 21966 419 22032 435
rect 21966 355 21967 419
rect 22031 355 22032 419
rect 21966 339 22032 355
rect 21966 275 21967 339
rect 22031 275 22032 339
rect 21966 259 22032 275
rect 21966 195 21967 259
rect 22031 195 22032 259
rect 21966 179 22032 195
rect 21966 115 21967 179
rect 22031 115 22032 179
rect 21966 99 22032 115
rect 21966 35 21967 99
rect 22031 35 22032 99
rect 21966 19 22032 35
rect 21966 -45 21967 19
rect 22031 -45 22032 19
rect 21966 -61 22032 -45
rect 21966 -125 21967 -61
rect 22031 -125 22032 -61
rect 21966 -141 22032 -125
rect 21966 -205 21967 -141
rect 22031 -205 22032 -141
rect 21966 -295 22032 -205
rect 22092 -299 22152 733
rect 22212 -359 22272 671
rect 22332 -299 22392 733
rect 22452 -359 22512 671
rect 22572 579 22638 733
rect 22572 515 22573 579
rect 22637 515 22638 579
rect 22572 499 22638 515
rect 22572 435 22573 499
rect 22637 435 22638 499
rect 22572 419 22638 435
rect 22572 355 22573 419
rect 22637 355 22638 419
rect 22572 339 22638 355
rect 22572 275 22573 339
rect 22637 275 22638 339
rect 22572 259 22638 275
rect 22572 195 22573 259
rect 22637 195 22638 259
rect 22572 179 22638 195
rect 22572 115 22573 179
rect 22637 115 22638 179
rect 22572 99 22638 115
rect 22572 35 22573 99
rect 22637 35 22638 99
rect 22572 19 22638 35
rect 22572 -45 22573 19
rect 22637 -45 22638 19
rect 22572 -61 22638 -45
rect 22572 -125 22573 -61
rect 22637 -125 22638 -61
rect 22572 -141 22638 -125
rect 22572 -205 22573 -141
rect 22637 -205 22638 -141
rect 22572 -295 22638 -205
rect 22698 -299 22758 733
rect 22818 -359 22878 671
rect 22938 -299 22998 733
rect 23058 -359 23118 671
rect 23178 579 23244 733
rect 23178 515 23179 579
rect 23243 515 23244 579
rect 23178 499 23244 515
rect 23178 435 23179 499
rect 23243 435 23244 499
rect 23178 419 23244 435
rect 23178 355 23179 419
rect 23243 355 23244 419
rect 23178 339 23244 355
rect 23178 275 23179 339
rect 23243 275 23244 339
rect 23178 259 23244 275
rect 23178 195 23179 259
rect 23243 195 23244 259
rect 23178 179 23244 195
rect 23178 115 23179 179
rect 23243 115 23244 179
rect 23178 99 23244 115
rect 23178 35 23179 99
rect 23243 35 23244 99
rect 23178 19 23244 35
rect 23178 -45 23179 19
rect 23243 -45 23244 19
rect 23178 -61 23244 -45
rect 23178 -125 23179 -61
rect 23243 -125 23244 -61
rect 23178 -141 23244 -125
rect 23178 -205 23179 -141
rect 23243 -205 23244 -141
rect 23178 -295 23244 -205
rect 23304 -299 23364 733
rect 23424 -359 23484 671
rect 23544 -299 23604 733
rect 23664 -359 23724 671
rect 23784 579 23850 733
rect 23784 515 23785 579
rect 23849 515 23850 579
rect 23784 499 23850 515
rect 23784 435 23785 499
rect 23849 435 23850 499
rect 23784 419 23850 435
rect 23784 355 23785 419
rect 23849 355 23850 419
rect 23784 339 23850 355
rect 23784 275 23785 339
rect 23849 275 23850 339
rect 23784 259 23850 275
rect 23784 195 23785 259
rect 23849 195 23850 259
rect 23784 179 23850 195
rect 23784 115 23785 179
rect 23849 115 23850 179
rect 23784 99 23850 115
rect 23784 35 23785 99
rect 23849 35 23850 99
rect 23784 19 23850 35
rect 23784 -45 23785 19
rect 23849 -45 23850 19
rect 23784 -61 23850 -45
rect 23784 -125 23785 -61
rect 23849 -125 23850 -61
rect 23784 -141 23850 -125
rect 23784 -205 23785 -141
rect 23849 -205 23850 -141
rect 23784 -295 23850 -205
rect 23910 -299 23970 733
rect 24030 -359 24090 671
rect 24150 -299 24210 733
rect 24270 -359 24330 671
rect 24390 579 24456 733
rect 24390 515 24391 579
rect 24455 515 24456 579
rect 24390 499 24456 515
rect 24390 435 24391 499
rect 24455 435 24456 499
rect 24390 419 24456 435
rect 24390 355 24391 419
rect 24455 355 24456 419
rect 24390 339 24456 355
rect 24390 275 24391 339
rect 24455 275 24456 339
rect 24390 259 24456 275
rect 24390 195 24391 259
rect 24455 195 24456 259
rect 24390 179 24456 195
rect 24390 115 24391 179
rect 24455 115 24456 179
rect 24390 99 24456 115
rect 24390 35 24391 99
rect 24455 35 24456 99
rect 24390 19 24456 35
rect 24390 -45 24391 19
rect 24455 -45 24456 19
rect 24390 -61 24456 -45
rect 24390 -125 24391 -61
rect 24455 -125 24456 -61
rect 24390 -141 24456 -125
rect 24390 -205 24391 -141
rect 24455 -205 24456 -141
rect 24390 -295 24456 -205
rect 24516 -299 24576 733
rect 24636 -359 24696 671
rect 24756 -299 24816 733
rect 24876 -359 24936 671
rect 24996 579 25062 733
rect 24996 515 24997 579
rect 25061 515 25062 579
rect 24996 499 25062 515
rect 24996 435 24997 499
rect 25061 435 25062 499
rect 24996 419 25062 435
rect 24996 355 24997 419
rect 25061 355 25062 419
rect 24996 339 25062 355
rect 24996 275 24997 339
rect 25061 275 25062 339
rect 24996 259 25062 275
rect 24996 195 24997 259
rect 25061 195 25062 259
rect 24996 179 25062 195
rect 24996 115 24997 179
rect 25061 115 25062 179
rect 24996 99 25062 115
rect 24996 35 24997 99
rect 25061 35 25062 99
rect 24996 19 25062 35
rect 24996 -45 24997 19
rect 25061 -45 25062 19
rect 24996 -61 25062 -45
rect 24996 -125 24997 -61
rect 25061 -125 25062 -61
rect 24996 -141 25062 -125
rect 24996 -205 24997 -141
rect 25061 -205 25062 -141
rect 24996 -295 25062 -205
rect 25122 -299 25182 733
rect 25242 -359 25302 671
rect 25362 -299 25422 733
rect 25482 -359 25542 671
rect 25602 579 25668 733
rect 25602 515 25603 579
rect 25667 515 25668 579
rect 25602 499 25668 515
rect 25602 435 25603 499
rect 25667 435 25668 499
rect 25602 419 25668 435
rect 25602 355 25603 419
rect 25667 355 25668 419
rect 25602 339 25668 355
rect 25602 275 25603 339
rect 25667 275 25668 339
rect 25602 259 25668 275
rect 25602 195 25603 259
rect 25667 195 25668 259
rect 25602 179 25668 195
rect 25602 115 25603 179
rect 25667 115 25668 179
rect 25602 99 25668 115
rect 25602 35 25603 99
rect 25667 35 25668 99
rect 25602 19 25668 35
rect 25602 -45 25603 19
rect 25667 -45 25668 19
rect 25602 -61 25668 -45
rect 25602 -125 25603 -61
rect 25667 -125 25668 -61
rect 25602 -141 25668 -125
rect 25602 -205 25603 -141
rect 25667 -205 25668 -141
rect 25602 -295 25668 -205
rect 25728 -299 25788 733
rect 25848 -359 25908 671
rect 25968 -299 26028 733
rect 26088 -359 26148 671
rect 26208 579 26274 733
rect 26208 515 26209 579
rect 26273 515 26274 579
rect 26208 499 26274 515
rect 26208 435 26209 499
rect 26273 435 26274 499
rect 26208 419 26274 435
rect 26208 355 26209 419
rect 26273 355 26274 419
rect 26208 339 26274 355
rect 26208 275 26209 339
rect 26273 275 26274 339
rect 26208 259 26274 275
rect 26208 195 26209 259
rect 26273 195 26274 259
rect 26208 179 26274 195
rect 26208 115 26209 179
rect 26273 115 26274 179
rect 26208 99 26274 115
rect 26208 35 26209 99
rect 26273 35 26274 99
rect 26208 19 26274 35
rect 26208 -45 26209 19
rect 26273 -45 26274 19
rect 26208 -61 26274 -45
rect 26208 -125 26209 -61
rect 26273 -125 26274 -61
rect 26208 -141 26274 -125
rect 26208 -205 26209 -141
rect 26273 -205 26274 -141
rect 26208 -295 26274 -205
rect 26334 -299 26394 733
rect 26454 -359 26514 671
rect 26574 -299 26634 733
rect 26694 -359 26754 671
rect 26814 579 26880 733
rect 26814 515 26815 579
rect 26879 515 26880 579
rect 26814 499 26880 515
rect 26814 435 26815 499
rect 26879 435 26880 499
rect 26814 419 26880 435
rect 26814 355 26815 419
rect 26879 355 26880 419
rect 26814 339 26880 355
rect 26814 275 26815 339
rect 26879 275 26880 339
rect 26814 259 26880 275
rect 26814 195 26815 259
rect 26879 195 26880 259
rect 26814 179 26880 195
rect 26814 115 26815 179
rect 26879 115 26880 179
rect 26814 99 26880 115
rect 26814 35 26815 99
rect 26879 35 26880 99
rect 26814 19 26880 35
rect 26814 -45 26815 19
rect 26879 -45 26880 19
rect 26814 -61 26880 -45
rect 26814 -125 26815 -61
rect 26879 -125 26880 -61
rect 26814 -141 26880 -125
rect 26814 -205 26815 -141
rect 26879 -205 26880 -141
rect 26814 -295 26880 -205
rect 26940 -299 27000 733
rect 27060 -359 27120 671
rect 27180 -299 27240 733
rect 27300 -359 27360 671
rect 27420 579 27486 733
rect 27420 515 27421 579
rect 27485 515 27486 579
rect 27420 499 27486 515
rect 27420 435 27421 499
rect 27485 435 27486 499
rect 27420 419 27486 435
rect 27420 355 27421 419
rect 27485 355 27486 419
rect 27420 339 27486 355
rect 27420 275 27421 339
rect 27485 275 27486 339
rect 27420 259 27486 275
rect 27420 195 27421 259
rect 27485 195 27486 259
rect 27420 179 27486 195
rect 27420 115 27421 179
rect 27485 115 27486 179
rect 27420 99 27486 115
rect 27420 35 27421 99
rect 27485 35 27486 99
rect 27420 19 27486 35
rect 27420 -45 27421 19
rect 27485 -45 27486 19
rect 27420 -61 27486 -45
rect 27420 -125 27421 -61
rect 27485 -125 27486 -61
rect 27420 -141 27486 -125
rect 27420 -205 27421 -141
rect 27485 -205 27486 -141
rect 27420 -295 27486 -205
rect 27546 -299 27606 733
rect 27666 -359 27726 671
rect 27786 -299 27846 733
rect 27906 -359 27966 671
rect 28026 579 28092 733
rect 28026 515 28027 579
rect 28091 515 28092 579
rect 28026 499 28092 515
rect 28026 435 28027 499
rect 28091 435 28092 499
rect 28026 419 28092 435
rect 28026 355 28027 419
rect 28091 355 28092 419
rect 28026 339 28092 355
rect 28026 275 28027 339
rect 28091 275 28092 339
rect 28026 259 28092 275
rect 28026 195 28027 259
rect 28091 195 28092 259
rect 28026 179 28092 195
rect 28026 115 28027 179
rect 28091 115 28092 179
rect 28026 99 28092 115
rect 28026 35 28027 99
rect 28091 35 28092 99
rect 28026 19 28092 35
rect 28026 -45 28027 19
rect 28091 -45 28092 19
rect 28026 -61 28092 -45
rect 28026 -125 28027 -61
rect 28091 -125 28092 -61
rect 28026 -141 28092 -125
rect 28026 -205 28027 -141
rect 28091 -205 28092 -141
rect 28026 -295 28092 -205
rect 28152 -299 28212 733
rect 28272 -359 28332 671
rect 28392 -299 28452 733
rect 28512 -359 28572 671
rect 28632 579 28698 733
rect 28632 515 28633 579
rect 28697 515 28698 579
rect 28632 499 28698 515
rect 28632 435 28633 499
rect 28697 435 28698 499
rect 28632 419 28698 435
rect 28632 355 28633 419
rect 28697 355 28698 419
rect 28632 339 28698 355
rect 28632 275 28633 339
rect 28697 275 28698 339
rect 28632 259 28698 275
rect 28632 195 28633 259
rect 28697 195 28698 259
rect 28632 179 28698 195
rect 28632 115 28633 179
rect 28697 115 28698 179
rect 28632 99 28698 115
rect 28632 35 28633 99
rect 28697 35 28698 99
rect 28632 19 28698 35
rect 28632 -45 28633 19
rect 28697 -45 28698 19
rect 28632 -61 28698 -45
rect 28632 -125 28633 -61
rect 28697 -125 28698 -61
rect 28632 -141 28698 -125
rect 28632 -205 28633 -141
rect 28697 -205 28698 -141
rect 28632 -295 28698 -205
rect 28758 -299 28818 733
rect 28878 -359 28938 671
rect 28998 -299 29058 733
rect 29118 -359 29178 671
rect 29238 579 29304 733
rect 29238 515 29239 579
rect 29303 515 29304 579
rect 29238 499 29304 515
rect 29238 435 29239 499
rect 29303 435 29304 499
rect 29238 419 29304 435
rect 29238 355 29239 419
rect 29303 355 29304 419
rect 29238 339 29304 355
rect 29238 275 29239 339
rect 29303 275 29304 339
rect 29238 259 29304 275
rect 29238 195 29239 259
rect 29303 195 29304 259
rect 29238 179 29304 195
rect 29238 115 29239 179
rect 29303 115 29304 179
rect 29238 99 29304 115
rect 29238 35 29239 99
rect 29303 35 29304 99
rect 29238 19 29304 35
rect 29238 -45 29239 19
rect 29303 -45 29304 19
rect 29238 -61 29304 -45
rect 29238 -125 29239 -61
rect 29303 -125 29304 -61
rect 29238 -141 29304 -125
rect 29238 -205 29239 -141
rect 29303 -205 29304 -141
rect 29238 -295 29304 -205
rect 29364 -299 29424 733
rect 29484 -359 29544 671
rect 29604 -299 29664 733
rect 29724 -359 29784 671
rect 29844 579 29910 733
rect 29844 515 29845 579
rect 29909 515 29910 579
rect 29844 499 29910 515
rect 29844 435 29845 499
rect 29909 435 29910 499
rect 29844 419 29910 435
rect 29844 355 29845 419
rect 29909 355 29910 419
rect 29844 339 29910 355
rect 29844 275 29845 339
rect 29909 275 29910 339
rect 29844 259 29910 275
rect 29844 195 29845 259
rect 29909 195 29910 259
rect 29844 179 29910 195
rect 29844 115 29845 179
rect 29909 115 29910 179
rect 29844 99 29910 115
rect 29844 35 29845 99
rect 29909 35 29910 99
rect 29844 19 29910 35
rect 29844 -45 29845 19
rect 29909 -45 29910 19
rect 29844 -61 29910 -45
rect 29844 -125 29845 -61
rect 29909 -125 29910 -61
rect 29844 -141 29910 -125
rect 29844 -205 29845 -141
rect 29909 -205 29910 -141
rect 29844 -295 29910 -205
rect 29970 -299 30030 733
rect 30090 -359 30150 671
rect 30210 -299 30270 733
rect 30330 -359 30390 671
rect 30450 579 30516 733
rect 30450 515 30451 579
rect 30515 515 30516 579
rect 30450 499 30516 515
rect 30450 435 30451 499
rect 30515 435 30516 499
rect 30450 419 30516 435
rect 30450 355 30451 419
rect 30515 355 30516 419
rect 30450 339 30516 355
rect 30450 275 30451 339
rect 30515 275 30516 339
rect 30450 259 30516 275
rect 30450 195 30451 259
rect 30515 195 30516 259
rect 30450 179 30516 195
rect 30450 115 30451 179
rect 30515 115 30516 179
rect 30450 99 30516 115
rect 30450 35 30451 99
rect 30515 35 30516 99
rect 30450 19 30516 35
rect 30450 -45 30451 19
rect 30515 -45 30516 19
rect 30450 -61 30516 -45
rect 30450 -125 30451 -61
rect 30515 -125 30516 -61
rect 30450 -141 30516 -125
rect 30450 -205 30451 -141
rect 30515 -205 30516 -141
rect 30450 -295 30516 -205
rect 30576 -299 30636 733
rect 30696 -359 30756 671
rect 30816 -299 30876 733
rect 30936 -359 30996 671
rect 31056 579 31122 733
rect 31056 515 31057 579
rect 31121 515 31122 579
rect 31056 499 31122 515
rect 31056 435 31057 499
rect 31121 435 31122 499
rect 31056 419 31122 435
rect 31056 355 31057 419
rect 31121 355 31122 419
rect 31056 339 31122 355
rect 31056 275 31057 339
rect 31121 275 31122 339
rect 31056 259 31122 275
rect 31056 195 31057 259
rect 31121 195 31122 259
rect 31056 179 31122 195
rect 31056 115 31057 179
rect 31121 115 31122 179
rect 31056 99 31122 115
rect 31056 35 31057 99
rect 31121 35 31122 99
rect 31056 19 31122 35
rect 31056 -45 31057 19
rect 31121 -45 31122 19
rect 31056 -61 31122 -45
rect 31056 -125 31057 -61
rect 31121 -125 31122 -61
rect 31056 -141 31122 -125
rect 31056 -205 31057 -141
rect 31121 -205 31122 -141
rect 31056 -295 31122 -205
rect 31182 -299 31242 733
rect 31302 -359 31362 671
rect 31422 -299 31482 733
rect 31542 -359 31602 671
rect 31662 579 31728 733
rect 31662 515 31663 579
rect 31727 515 31728 579
rect 31662 499 31728 515
rect 31662 435 31663 499
rect 31727 435 31728 499
rect 31662 419 31728 435
rect 31662 355 31663 419
rect 31727 355 31728 419
rect 31662 339 31728 355
rect 31662 275 31663 339
rect 31727 275 31728 339
rect 31662 259 31728 275
rect 31662 195 31663 259
rect 31727 195 31728 259
rect 31662 179 31728 195
rect 31662 115 31663 179
rect 31727 115 31728 179
rect 31662 99 31728 115
rect 31662 35 31663 99
rect 31727 35 31728 99
rect 31662 19 31728 35
rect 31662 -45 31663 19
rect 31727 -45 31728 19
rect 31662 -61 31728 -45
rect 31662 -125 31663 -61
rect 31727 -125 31728 -61
rect 31662 -141 31728 -125
rect 31662 -205 31663 -141
rect 31727 -205 31728 -141
rect 31662 -295 31728 -205
rect 31788 -299 31848 733
rect 31908 -359 31968 671
rect 32028 -299 32088 733
rect 32148 -359 32208 671
rect 32268 579 32334 733
rect 32268 515 32269 579
rect 32333 515 32334 579
rect 32268 499 32334 515
rect 32268 435 32269 499
rect 32333 435 32334 499
rect 32268 419 32334 435
rect 32268 355 32269 419
rect 32333 355 32334 419
rect 32268 339 32334 355
rect 32268 275 32269 339
rect 32333 275 32334 339
rect 32268 259 32334 275
rect 32268 195 32269 259
rect 32333 195 32334 259
rect 32268 179 32334 195
rect 32268 115 32269 179
rect 32333 115 32334 179
rect 32268 99 32334 115
rect 32268 35 32269 99
rect 32333 35 32334 99
rect 32268 19 32334 35
rect 32268 -45 32269 19
rect 32333 -45 32334 19
rect 32268 -61 32334 -45
rect 32268 -125 32269 -61
rect 32333 -125 32334 -61
rect 32268 -141 32334 -125
rect 32268 -205 32269 -141
rect 32333 -205 32334 -141
rect 32268 -295 32334 -205
rect 32394 -299 32454 733
rect 32514 -359 32574 671
rect 32634 -299 32694 733
rect 32754 -359 32814 671
rect 32874 579 32940 733
rect 32874 515 32875 579
rect 32939 515 32940 579
rect 32874 499 32940 515
rect 32874 435 32875 499
rect 32939 435 32940 499
rect 32874 419 32940 435
rect 32874 355 32875 419
rect 32939 355 32940 419
rect 32874 339 32940 355
rect 32874 275 32875 339
rect 32939 275 32940 339
rect 32874 259 32940 275
rect 32874 195 32875 259
rect 32939 195 32940 259
rect 32874 179 32940 195
rect 32874 115 32875 179
rect 32939 115 32940 179
rect 32874 99 32940 115
rect 32874 35 32875 99
rect 32939 35 32940 99
rect 32874 19 32940 35
rect 32874 -45 32875 19
rect 32939 -45 32940 19
rect 32874 -61 32940 -45
rect 32874 -125 32875 -61
rect 32939 -125 32940 -61
rect 32874 -141 32940 -125
rect 32874 -205 32875 -141
rect 32939 -205 32940 -141
rect 32874 -295 32940 -205
rect 33000 -299 33060 733
rect 33120 -359 33180 671
rect 33240 -299 33300 733
rect 33360 -359 33420 671
rect 33480 579 33546 733
rect 33480 515 33481 579
rect 33545 515 33546 579
rect 33480 499 33546 515
rect 33480 435 33481 499
rect 33545 435 33546 499
rect 33480 419 33546 435
rect 33480 355 33481 419
rect 33545 355 33546 419
rect 33480 339 33546 355
rect 33480 275 33481 339
rect 33545 275 33546 339
rect 33480 259 33546 275
rect 33480 195 33481 259
rect 33545 195 33546 259
rect 33480 179 33546 195
rect 33480 115 33481 179
rect 33545 115 33546 179
rect 33480 99 33546 115
rect 33480 35 33481 99
rect 33545 35 33546 99
rect 33480 19 33546 35
rect 33480 -45 33481 19
rect 33545 -45 33546 19
rect 33480 -61 33546 -45
rect 33480 -125 33481 -61
rect 33545 -125 33546 -61
rect 33480 -141 33546 -125
rect 33480 -205 33481 -141
rect 33545 -205 33546 -141
rect 33480 -295 33546 -205
rect 33606 -299 33666 733
rect 33726 -359 33786 671
rect 33846 -299 33906 733
rect 33966 -359 34026 671
rect 34086 579 34152 733
rect 34086 515 34087 579
rect 34151 515 34152 579
rect 34086 499 34152 515
rect 34086 435 34087 499
rect 34151 435 34152 499
rect 34086 419 34152 435
rect 34086 355 34087 419
rect 34151 355 34152 419
rect 34086 339 34152 355
rect 34086 275 34087 339
rect 34151 275 34152 339
rect 34086 259 34152 275
rect 34086 195 34087 259
rect 34151 195 34152 259
rect 34086 179 34152 195
rect 34086 115 34087 179
rect 34151 115 34152 179
rect 34086 99 34152 115
rect 34086 35 34087 99
rect 34151 35 34152 99
rect 34086 19 34152 35
rect 34086 -45 34087 19
rect 34151 -45 34152 19
rect 34086 -61 34152 -45
rect 34086 -125 34087 -61
rect 34151 -125 34152 -61
rect 34086 -141 34152 -125
rect 34086 -205 34087 -141
rect 34151 -205 34152 -141
rect 34086 -295 34152 -205
rect 34212 -299 34272 733
rect 34332 -359 34392 671
rect 34452 -299 34512 733
rect 34572 -359 34632 671
rect 34692 579 34758 733
rect 34692 515 34693 579
rect 34757 515 34758 579
rect 34692 499 34758 515
rect 34692 435 34693 499
rect 34757 435 34758 499
rect 34692 419 34758 435
rect 34692 355 34693 419
rect 34757 355 34758 419
rect 34692 339 34758 355
rect 34692 275 34693 339
rect 34757 275 34758 339
rect 34692 259 34758 275
rect 34692 195 34693 259
rect 34757 195 34758 259
rect 34692 179 34758 195
rect 34692 115 34693 179
rect 34757 115 34758 179
rect 34692 99 34758 115
rect 34692 35 34693 99
rect 34757 35 34758 99
rect 34692 19 34758 35
rect 34692 -45 34693 19
rect 34757 -45 34758 19
rect 34692 -61 34758 -45
rect 34692 -125 34693 -61
rect 34757 -125 34758 -61
rect 34692 -141 34758 -125
rect 34692 -205 34693 -141
rect 34757 -205 34758 -141
rect 34692 -295 34758 -205
rect 34818 -299 34878 733
rect 34938 -359 34998 671
rect 35058 -299 35118 733
rect 35178 -359 35238 671
rect 35298 579 35364 733
rect 35298 515 35299 579
rect 35363 515 35364 579
rect 35298 499 35364 515
rect 35298 435 35299 499
rect 35363 435 35364 499
rect 35298 419 35364 435
rect 35298 355 35299 419
rect 35363 355 35364 419
rect 35298 339 35364 355
rect 35298 275 35299 339
rect 35363 275 35364 339
rect 35298 259 35364 275
rect 35298 195 35299 259
rect 35363 195 35364 259
rect 35298 179 35364 195
rect 35298 115 35299 179
rect 35363 115 35364 179
rect 35298 99 35364 115
rect 35298 35 35299 99
rect 35363 35 35364 99
rect 35298 19 35364 35
rect 35298 -45 35299 19
rect 35363 -45 35364 19
rect 35298 -61 35364 -45
rect 35298 -125 35299 -61
rect 35363 -125 35364 -61
rect 35298 -141 35364 -125
rect 35298 -205 35299 -141
rect 35363 -205 35364 -141
rect 35298 -295 35364 -205
rect 35424 -299 35484 733
rect 35544 -359 35604 671
rect 35664 -299 35724 733
rect 35784 -359 35844 671
rect 35904 579 35970 733
rect 35904 515 35905 579
rect 35969 515 35970 579
rect 35904 499 35970 515
rect 35904 435 35905 499
rect 35969 435 35970 499
rect 35904 419 35970 435
rect 35904 355 35905 419
rect 35969 355 35970 419
rect 35904 339 35970 355
rect 35904 275 35905 339
rect 35969 275 35970 339
rect 35904 259 35970 275
rect 35904 195 35905 259
rect 35969 195 35970 259
rect 35904 179 35970 195
rect 35904 115 35905 179
rect 35969 115 35970 179
rect 35904 99 35970 115
rect 35904 35 35905 99
rect 35969 35 35970 99
rect 35904 19 35970 35
rect 35904 -45 35905 19
rect 35969 -45 35970 19
rect 35904 -61 35970 -45
rect 35904 -125 35905 -61
rect 35969 -125 35970 -61
rect 35904 -141 35970 -125
rect 35904 -205 35905 -141
rect 35969 -205 35970 -141
rect 35904 -295 35970 -205
rect 36030 -299 36090 733
rect 36150 -359 36210 671
rect 36270 -299 36330 733
rect 36390 -359 36450 671
rect 36510 579 36576 733
rect 36510 515 36511 579
rect 36575 515 36576 579
rect 36510 499 36576 515
rect 36510 435 36511 499
rect 36575 435 36576 499
rect 36510 419 36576 435
rect 36510 355 36511 419
rect 36575 355 36576 419
rect 36510 339 36576 355
rect 36510 275 36511 339
rect 36575 275 36576 339
rect 36510 259 36576 275
rect 36510 195 36511 259
rect 36575 195 36576 259
rect 36510 179 36576 195
rect 36510 115 36511 179
rect 36575 115 36576 179
rect 36510 99 36576 115
rect 36510 35 36511 99
rect 36575 35 36576 99
rect 36510 19 36576 35
rect 36510 -45 36511 19
rect 36575 -45 36576 19
rect 36510 -61 36576 -45
rect 36510 -125 36511 -61
rect 36575 -125 36576 -61
rect 36510 -141 36576 -125
rect 36510 -205 36511 -141
rect 36575 -205 36576 -141
rect 36510 -295 36576 -205
rect 36636 -299 36696 733
rect 36756 -359 36816 671
rect 36876 -299 36936 733
rect 36996 -359 37056 671
rect 37116 579 37182 733
rect 37116 515 37117 579
rect 37181 515 37182 579
rect 37116 499 37182 515
rect 37116 435 37117 499
rect 37181 435 37182 499
rect 37116 419 37182 435
rect 37116 355 37117 419
rect 37181 355 37182 419
rect 37116 339 37182 355
rect 37116 275 37117 339
rect 37181 275 37182 339
rect 37116 259 37182 275
rect 37116 195 37117 259
rect 37181 195 37182 259
rect 37116 179 37182 195
rect 37116 115 37117 179
rect 37181 115 37182 179
rect 37116 99 37182 115
rect 37116 35 37117 99
rect 37181 35 37182 99
rect 37116 19 37182 35
rect 37116 -45 37117 19
rect 37181 -45 37182 19
rect 37116 -61 37182 -45
rect 37116 -125 37117 -61
rect 37181 -125 37182 -61
rect 37116 -141 37182 -125
rect 37116 -205 37117 -141
rect 37181 -205 37182 -141
rect 37116 -295 37182 -205
rect 37242 -299 37302 733
rect 37362 -359 37422 671
rect 37482 -299 37542 733
rect 37602 -359 37662 671
rect 37722 579 37788 733
rect 37722 515 37723 579
rect 37787 515 37788 579
rect 37722 499 37788 515
rect 37722 435 37723 499
rect 37787 435 37788 499
rect 37722 419 37788 435
rect 37722 355 37723 419
rect 37787 355 37788 419
rect 37722 339 37788 355
rect 37722 275 37723 339
rect 37787 275 37788 339
rect 37722 259 37788 275
rect 37722 195 37723 259
rect 37787 195 37788 259
rect 37722 179 37788 195
rect 37722 115 37723 179
rect 37787 115 37788 179
rect 37722 99 37788 115
rect 37722 35 37723 99
rect 37787 35 37788 99
rect 37722 19 37788 35
rect 37722 -45 37723 19
rect 37787 -45 37788 19
rect 37722 -61 37788 -45
rect 37722 -125 37723 -61
rect 37787 -125 37788 -61
rect 37722 -141 37788 -125
rect 37722 -205 37723 -141
rect 37787 -205 37788 -141
rect 37722 -295 37788 -205
rect 37848 -299 37908 733
rect 37968 -359 38028 671
rect 38088 -299 38148 733
rect 38208 -359 38268 671
rect 38328 579 38394 733
rect 38328 515 38329 579
rect 38393 515 38394 579
rect 38328 499 38394 515
rect 38328 435 38329 499
rect 38393 435 38394 499
rect 38328 419 38394 435
rect 38328 355 38329 419
rect 38393 355 38394 419
rect 38328 339 38394 355
rect 38328 275 38329 339
rect 38393 275 38394 339
rect 38328 259 38394 275
rect 38328 195 38329 259
rect 38393 195 38394 259
rect 38328 179 38394 195
rect 38328 115 38329 179
rect 38393 115 38394 179
rect 38328 99 38394 115
rect 38328 35 38329 99
rect 38393 35 38394 99
rect 38328 19 38394 35
rect 38328 -45 38329 19
rect 38393 -45 38394 19
rect 38328 -61 38394 -45
rect 38328 -125 38329 -61
rect 38393 -125 38394 -61
rect 38328 -141 38394 -125
rect 38328 -205 38329 -141
rect 38393 -205 38394 -141
rect 38328 -295 38394 -205
rect 38454 -299 38514 733
rect 38574 -359 38634 671
rect 38694 -299 38754 733
rect 38814 -359 38874 671
rect 38934 579 39000 733
rect 38934 515 38935 579
rect 38999 515 39000 579
rect 38934 499 39000 515
rect 38934 435 38935 499
rect 38999 435 39000 499
rect 38934 419 39000 435
rect 38934 355 38935 419
rect 38999 355 39000 419
rect 38934 339 39000 355
rect 38934 275 38935 339
rect 38999 275 39000 339
rect 38934 259 39000 275
rect 38934 195 38935 259
rect 38999 195 39000 259
rect 38934 179 39000 195
rect 38934 115 38935 179
rect 38999 115 39000 179
rect 38934 99 39000 115
rect 38934 35 38935 99
rect 38999 35 39000 99
rect 38934 19 39000 35
rect 38934 -45 38935 19
rect 38999 -45 39000 19
rect 38934 -61 39000 -45
rect 38934 -125 38935 -61
rect 38999 -125 39000 -61
rect 38934 -141 39000 -125
rect 38934 -205 38935 -141
rect 38999 -205 39000 -141
rect 38934 -295 39000 -205
rect 39060 -299 39120 733
rect 39180 -359 39240 671
rect 39300 -299 39360 733
rect 39420 -359 39480 671
rect 39540 579 39606 733
rect 39540 515 39541 579
rect 39605 515 39606 579
rect 39540 499 39606 515
rect 39540 435 39541 499
rect 39605 435 39606 499
rect 39540 419 39606 435
rect 39540 355 39541 419
rect 39605 355 39606 419
rect 39540 339 39606 355
rect 39540 275 39541 339
rect 39605 275 39606 339
rect 39540 259 39606 275
rect 39540 195 39541 259
rect 39605 195 39606 259
rect 39540 179 39606 195
rect 39540 115 39541 179
rect 39605 115 39606 179
rect 39540 99 39606 115
rect 39540 35 39541 99
rect 39605 35 39606 99
rect 39540 19 39606 35
rect 39540 -45 39541 19
rect 39605 -45 39606 19
rect 39540 -61 39606 -45
rect 39540 -125 39541 -61
rect 39605 -125 39606 -61
rect 39540 -141 39606 -125
rect 39540 -205 39541 -141
rect 39605 -205 39606 -141
rect 39540 -295 39606 -205
rect -459 -361 213 -359
rect -459 -425 -355 -361
rect -291 -425 -275 -361
rect -211 -425 -195 -361
rect -131 -425 -115 -361
rect -51 -425 -35 -361
rect 29 -425 45 -361
rect 109 -425 213 -361
rect -459 -427 213 -425
rect 524 -361 1027 -359
rect 524 -425 539 -361
rect 603 -425 619 -361
rect 683 -425 699 -361
rect 763 -425 779 -361
rect 843 -425 859 -361
rect 923 -425 1027 -361
rect 524 -427 1027 -425
rect 1267 -361 1717 -359
rect 1954 -361 2545 -359
rect 1267 -425 1371 -361
rect 1435 -425 1451 -361
rect 1515 -425 1531 -361
rect 1595 -425 1611 -361
rect 1675 -425 1691 -361
rect 1954 -425 1977 -361
rect 2041 -425 2057 -361
rect 2121 -425 2137 -361
rect 2201 -425 2217 -361
rect 2281 -425 2297 -361
rect 2361 -425 2377 -361
rect 2441 -425 2545 -361
rect 1267 -427 1717 -425
rect 1954 -427 2545 -425
rect 2801 -361 3301 -359
rect 3538 -361 5291 -359
rect 2801 -425 2905 -361
rect 2969 -425 2985 -361
rect 3049 -425 3065 -361
rect 3129 -425 3145 -361
rect 3209 -425 3225 -361
rect 3289 -425 3301 -361
rect 3575 -425 3591 -361
rect 3655 -425 3671 -361
rect 3735 -425 3751 -361
rect 3815 -425 3831 -361
rect 3895 -425 3911 -361
rect 3975 -425 4117 -361
rect 4181 -425 4197 -361
rect 4261 -425 4277 -361
rect 4341 -425 4357 -361
rect 4421 -425 4437 -361
rect 4501 -425 4517 -361
rect 4581 -425 4723 -361
rect 4787 -425 4803 -361
rect 4867 -425 4883 -361
rect 4947 -425 4963 -361
rect 5027 -425 5043 -361
rect 5107 -425 5123 -361
rect 5187 -425 5291 -361
rect 2801 -427 3301 -425
rect 3538 -427 5291 -425
rect 5352 -427 5394 -359
rect 5631 -361 10266 -359
rect 5680 -425 5696 -361
rect 5760 -425 5776 -361
rect 5840 -425 5856 -361
rect 5920 -425 6062 -361
rect 6126 -425 6142 -361
rect 6206 -425 6222 -361
rect 6286 -425 6302 -361
rect 6366 -425 6382 -361
rect 6446 -425 6462 -361
rect 6526 -425 6668 -361
rect 6732 -425 6748 -361
rect 6812 -425 6828 -361
rect 6892 -425 6908 -361
rect 6972 -425 6988 -361
rect 7052 -425 7068 -361
rect 7132 -425 7274 -361
rect 7338 -425 7354 -361
rect 7418 -425 7434 -361
rect 7498 -425 7514 -361
rect 7578 -425 7594 -361
rect 7658 -425 7674 -361
rect 7738 -425 7880 -361
rect 7944 -425 7960 -361
rect 8024 -425 8040 -361
rect 8104 -425 8120 -361
rect 8184 -425 8200 -361
rect 8264 -425 8280 -361
rect 8344 -425 8486 -361
rect 8550 -425 8566 -361
rect 8630 -425 8646 -361
rect 8710 -425 8726 -361
rect 8790 -425 8806 -361
rect 8870 -425 8886 -361
rect 8950 -425 9092 -361
rect 9156 -425 9172 -361
rect 9236 -425 9252 -361
rect 9316 -425 9332 -361
rect 9396 -425 9412 -361
rect 9476 -425 9492 -361
rect 9556 -425 9698 -361
rect 9762 -425 9778 -361
rect 9842 -425 9858 -361
rect 9922 -425 9938 -361
rect 10002 -425 10018 -361
rect 10082 -425 10098 -361
rect 10162 -425 10266 -361
rect 5631 -427 10266 -425
rect 10326 -427 10368 -359
rect 10605 -361 20088 -359
rect 10654 -425 10670 -361
rect 10734 -425 10750 -361
rect 10814 -425 10830 -361
rect 10894 -425 11036 -361
rect 11100 -425 11116 -361
rect 11180 -425 11196 -361
rect 11260 -425 11276 -361
rect 11340 -425 11356 -361
rect 11420 -425 11436 -361
rect 11500 -425 11642 -361
rect 11706 -425 11722 -361
rect 11786 -425 11802 -361
rect 11866 -425 11882 -361
rect 11946 -425 11962 -361
rect 12026 -425 12042 -361
rect 12106 -425 12248 -361
rect 12312 -425 12328 -361
rect 12392 -425 12408 -361
rect 12472 -425 12488 -361
rect 12552 -425 12568 -361
rect 12632 -425 12648 -361
rect 12712 -425 12854 -361
rect 12918 -425 12934 -361
rect 12998 -425 13014 -361
rect 13078 -425 13094 -361
rect 13158 -425 13174 -361
rect 13238 -425 13254 -361
rect 13318 -425 13460 -361
rect 13524 -425 13540 -361
rect 13604 -425 13620 -361
rect 13684 -425 13700 -361
rect 13764 -425 13780 -361
rect 13844 -425 13860 -361
rect 13924 -425 14066 -361
rect 14130 -425 14146 -361
rect 14210 -425 14226 -361
rect 14290 -425 14306 -361
rect 14370 -425 14386 -361
rect 14450 -425 14466 -361
rect 14530 -425 14672 -361
rect 14736 -425 14752 -361
rect 14816 -425 14832 -361
rect 14896 -425 14912 -361
rect 14976 -425 14992 -361
rect 15056 -425 15072 -361
rect 15136 -425 15278 -361
rect 15342 -425 15358 -361
rect 15422 -425 15438 -361
rect 15502 -425 15518 -361
rect 15582 -425 15598 -361
rect 15662 -425 15678 -361
rect 15742 -425 15884 -361
rect 15948 -425 15964 -361
rect 16028 -425 16044 -361
rect 16108 -425 16124 -361
rect 16188 -425 16204 -361
rect 16268 -425 16284 -361
rect 16348 -425 16490 -361
rect 16554 -425 16570 -361
rect 16634 -425 16650 -361
rect 16714 -425 16730 -361
rect 16794 -425 16810 -361
rect 16874 -425 16890 -361
rect 16954 -425 17096 -361
rect 17160 -425 17176 -361
rect 17240 -425 17256 -361
rect 17320 -425 17336 -361
rect 17400 -425 17416 -361
rect 17480 -425 17496 -361
rect 17560 -425 17702 -361
rect 17766 -425 17782 -361
rect 17846 -425 17862 -361
rect 17926 -425 17942 -361
rect 18006 -425 18022 -361
rect 18086 -425 18102 -361
rect 18166 -425 18308 -361
rect 18372 -425 18388 -361
rect 18452 -425 18468 -361
rect 18532 -425 18548 -361
rect 18612 -425 18628 -361
rect 18692 -425 18708 -361
rect 18772 -425 18914 -361
rect 18978 -425 18994 -361
rect 19058 -425 19074 -361
rect 19138 -425 19154 -361
rect 19218 -425 19234 -361
rect 19298 -425 19314 -361
rect 19378 -425 19520 -361
rect 19584 -425 19600 -361
rect 19664 -425 19680 -361
rect 19744 -425 19760 -361
rect 19824 -425 19840 -361
rect 19904 -425 19920 -361
rect 19984 -425 20088 -361
rect 10605 -427 20088 -425
rect 20148 -361 39298 -359
rect 20148 -425 20252 -361
rect 20316 -425 20332 -361
rect 20396 -425 20412 -361
rect 20476 -425 20492 -361
rect 20556 -425 20572 -361
rect 20636 -425 20652 -361
rect 20716 -425 20858 -361
rect 20922 -425 20938 -361
rect 21002 -425 21018 -361
rect 21082 -425 21098 -361
rect 21162 -425 21178 -361
rect 21242 -425 21258 -361
rect 21322 -425 21464 -361
rect 21528 -425 21544 -361
rect 21608 -425 21624 -361
rect 21688 -425 21704 -361
rect 21768 -425 21784 -361
rect 21848 -425 21864 -361
rect 21928 -425 22070 -361
rect 22134 -425 22150 -361
rect 22214 -425 22230 -361
rect 22294 -425 22310 -361
rect 22374 -425 22390 -361
rect 22454 -425 22470 -361
rect 22534 -425 22676 -361
rect 22740 -425 22756 -361
rect 22820 -425 22836 -361
rect 22900 -425 22916 -361
rect 22980 -425 22996 -361
rect 23060 -425 23076 -361
rect 23140 -425 23282 -361
rect 23346 -425 23362 -361
rect 23426 -425 23442 -361
rect 23506 -425 23522 -361
rect 23586 -425 23602 -361
rect 23666 -425 23682 -361
rect 23746 -425 23888 -361
rect 23952 -425 23968 -361
rect 24032 -425 24048 -361
rect 24112 -425 24128 -361
rect 24192 -425 24208 -361
rect 24272 -425 24288 -361
rect 24352 -425 24494 -361
rect 24558 -425 24574 -361
rect 24638 -425 24654 -361
rect 24718 -425 24734 -361
rect 24798 -425 24814 -361
rect 24878 -425 24894 -361
rect 24958 -425 25100 -361
rect 25164 -425 25180 -361
rect 25244 -425 25260 -361
rect 25324 -425 25340 -361
rect 25404 -425 25420 -361
rect 25484 -425 25500 -361
rect 25564 -425 25706 -361
rect 25770 -425 25786 -361
rect 25850 -425 25866 -361
rect 25930 -425 25946 -361
rect 26010 -425 26026 -361
rect 26090 -425 26106 -361
rect 26170 -425 26312 -361
rect 26376 -425 26392 -361
rect 26456 -425 26472 -361
rect 26536 -425 26552 -361
rect 26616 -425 26632 -361
rect 26696 -425 26712 -361
rect 26776 -425 26918 -361
rect 26982 -425 26998 -361
rect 27062 -425 27078 -361
rect 27142 -425 27158 -361
rect 27222 -425 27238 -361
rect 27302 -425 27318 -361
rect 27382 -425 27524 -361
rect 27588 -425 27604 -361
rect 27668 -425 27684 -361
rect 27748 -425 27764 -361
rect 27828 -425 27844 -361
rect 27908 -425 27924 -361
rect 27988 -425 28130 -361
rect 28194 -425 28210 -361
rect 28274 -425 28290 -361
rect 28354 -425 28370 -361
rect 28434 -425 28450 -361
rect 28514 -425 28530 -361
rect 28594 -425 28736 -361
rect 28800 -425 28816 -361
rect 28880 -425 28896 -361
rect 28960 -425 28976 -361
rect 29040 -425 29056 -361
rect 29120 -425 29136 -361
rect 29200 -425 29342 -361
rect 29406 -425 29422 -361
rect 29486 -425 29502 -361
rect 29566 -425 29582 -361
rect 29646 -425 29662 -361
rect 29726 -425 29742 -361
rect 29806 -425 29948 -361
rect 30012 -425 30028 -361
rect 30092 -425 30108 -361
rect 30172 -425 30188 -361
rect 30252 -425 30268 -361
rect 30332 -425 30348 -361
rect 30412 -425 30554 -361
rect 30618 -425 30634 -361
rect 30698 -425 30714 -361
rect 30778 -425 30794 -361
rect 30858 -425 30874 -361
rect 30938 -425 30954 -361
rect 31018 -425 31160 -361
rect 31224 -425 31240 -361
rect 31304 -425 31320 -361
rect 31384 -425 31400 -361
rect 31464 -425 31480 -361
rect 31544 -425 31560 -361
rect 31624 -425 31766 -361
rect 31830 -425 31846 -361
rect 31910 -425 31926 -361
rect 31990 -425 32006 -361
rect 32070 -425 32086 -361
rect 32150 -425 32166 -361
rect 32230 -425 32372 -361
rect 32436 -425 32452 -361
rect 32516 -425 32532 -361
rect 32596 -425 32612 -361
rect 32676 -425 32692 -361
rect 32756 -425 32772 -361
rect 32836 -425 32978 -361
rect 33042 -425 33058 -361
rect 33122 -425 33138 -361
rect 33202 -425 33218 -361
rect 33282 -425 33298 -361
rect 33362 -425 33378 -361
rect 33442 -425 33584 -361
rect 33648 -425 33664 -361
rect 33728 -425 33744 -361
rect 33808 -425 33824 -361
rect 33888 -425 33904 -361
rect 33968 -425 33984 -361
rect 34048 -425 34190 -361
rect 34254 -425 34270 -361
rect 34334 -425 34350 -361
rect 34414 -425 34430 -361
rect 34494 -425 34510 -361
rect 34574 -425 34590 -361
rect 34654 -425 34796 -361
rect 34860 -425 34876 -361
rect 34940 -425 34956 -361
rect 35020 -425 35036 -361
rect 35100 -425 35116 -361
rect 35180 -425 35196 -361
rect 35260 -425 35402 -361
rect 35466 -425 35482 -361
rect 35546 -425 35562 -361
rect 35626 -425 35642 -361
rect 35706 -425 35722 -361
rect 35786 -425 35802 -361
rect 35866 -425 36008 -361
rect 36072 -425 36088 -361
rect 36152 -425 36168 -361
rect 36232 -425 36248 -361
rect 36312 -425 36328 -361
rect 36392 -425 36408 -361
rect 36472 -425 36614 -361
rect 36678 -425 36694 -361
rect 36758 -425 36774 -361
rect 36838 -425 36854 -361
rect 36918 -425 36934 -361
rect 36998 -425 37014 -361
rect 37078 -425 37220 -361
rect 37284 -425 37300 -361
rect 37364 -425 37380 -361
rect 37444 -425 37460 -361
rect 37524 -425 37540 -361
rect 37604 -425 37620 -361
rect 37684 -425 37826 -361
rect 37890 -425 37906 -361
rect 37970 -425 37986 -361
rect 38050 -425 38066 -361
rect 38130 -425 38146 -361
rect 38210 -425 38226 -361
rect 38290 -425 38432 -361
rect 38496 -425 38512 -361
rect 38576 -425 38592 -361
rect 38656 -425 38672 -361
rect 38736 -425 38752 -361
rect 38816 -425 38832 -361
rect 38896 -425 39038 -361
rect 39102 -425 39118 -361
rect 39182 -425 39198 -361
rect 39262 -425 39278 -361
rect 20148 -427 39298 -425
rect 39534 -427 39606 -359
<< via4 >>
rect 287 5092 524 5262
rect 287 5028 459 5092
rect 459 5028 523 5092
rect 523 5028 524 5092
rect 287 5026 524 5028
rect 1717 5092 1954 5262
rect 1717 5028 1755 5092
rect 1755 5028 1771 5092
rect 1771 5028 1835 5092
rect 1835 5028 1954 5092
rect 1717 5026 1954 5028
rect 3301 5092 3538 5262
rect 3301 5028 3305 5092
rect 3305 5028 3369 5092
rect 3369 5028 3511 5092
rect 3511 5028 3538 5092
rect 3301 5026 3538 5028
rect 5394 5092 5631 5262
rect 5394 5028 5456 5092
rect 5456 5028 5520 5092
rect 5520 5028 5536 5092
rect 5536 5028 5600 5092
rect 5600 5028 5616 5092
rect 5616 5028 5631 5092
rect 5394 5026 5631 5028
rect 10368 5092 10605 5262
rect 10368 5028 10430 5092
rect 10430 5028 10494 5092
rect 10494 5028 10510 5092
rect 10510 5028 10574 5092
rect 10574 5028 10590 5092
rect 10590 5028 10605 5092
rect 10368 5026 10605 5028
rect 39298 5092 39534 5262
rect 39298 5028 39342 5092
rect 39342 5028 39358 5092
rect 39358 5028 39422 5092
rect 39422 5028 39438 5092
rect 39438 5028 39502 5092
rect 39502 5028 39534 5092
rect 39298 5026 39534 5028
rect 287 2772 524 2774
rect 287 2708 459 2772
rect 459 2708 523 2772
rect 523 2708 524 2772
rect 287 2538 524 2708
rect 1717 2772 1954 2774
rect 1717 2708 1755 2772
rect 1755 2708 1771 2772
rect 1771 2708 1835 2772
rect 1835 2708 1954 2772
rect 1717 2538 1954 2708
rect 3301 2772 3538 2774
rect 3301 2708 3305 2772
rect 3305 2708 3369 2772
rect 3369 2708 3511 2772
rect 3511 2708 3538 2772
rect 3301 2538 3538 2708
rect 5394 2772 5631 2774
rect 5394 2708 5456 2772
rect 5456 2708 5520 2772
rect 5520 2708 5536 2772
rect 5536 2708 5600 2772
rect 5600 2708 5616 2772
rect 5616 2708 5631 2772
rect 5394 2538 5631 2708
rect 10368 2772 10605 2774
rect 10368 2708 10430 2772
rect 10430 2708 10494 2772
rect 10494 2708 10510 2772
rect 10510 2708 10574 2772
rect 10574 2708 10590 2772
rect 10590 2708 10605 2772
rect 10368 2538 10605 2708
rect 39298 2772 39534 2774
rect 39298 2708 39342 2772
rect 39342 2708 39358 2772
rect 39358 2708 39422 2772
rect 39422 2708 39438 2772
rect 39438 2708 39502 2772
rect 39502 2708 39534 2772
rect 39298 2538 39534 2708
rect 287 1959 524 2129
rect 287 1895 459 1959
rect 459 1895 523 1959
rect 523 1895 524 1959
rect 287 1893 524 1895
rect 1717 1959 1954 2129
rect 1717 1895 1755 1959
rect 1755 1895 1771 1959
rect 1771 1895 1835 1959
rect 1835 1895 1954 1959
rect 1717 1893 1954 1895
rect 3301 1959 3538 2129
rect 3301 1895 3305 1959
rect 3305 1895 3369 1959
rect 3369 1895 3511 1959
rect 3511 1895 3538 1959
rect 3301 1893 3538 1895
rect 5394 1959 5631 2129
rect 5394 1895 5456 1959
rect 5456 1895 5520 1959
rect 5520 1895 5536 1959
rect 5536 1895 5600 1959
rect 5600 1895 5616 1959
rect 5616 1895 5631 1959
rect 5394 1893 5631 1895
rect 10368 1959 10605 2129
rect 10368 1895 10430 1959
rect 10430 1895 10494 1959
rect 10494 1895 10510 1959
rect 10510 1895 10574 1959
rect 10574 1895 10590 1959
rect 10590 1895 10605 1959
rect 10368 1893 10605 1895
rect 39298 1959 39534 2129
rect 39298 1895 39342 1959
rect 39342 1895 39358 1959
rect 39358 1895 39422 1959
rect 39422 1895 39438 1959
rect 39438 1895 39502 1959
rect 39502 1895 39534 1959
rect 39298 1893 39534 1895
rect 287 -361 524 -359
rect 287 -425 459 -361
rect 459 -425 523 -361
rect 523 -425 524 -361
rect 287 -595 524 -425
rect 1717 -361 1954 -359
rect 1717 -425 1755 -361
rect 1755 -425 1771 -361
rect 1771 -425 1835 -361
rect 1835 -425 1954 -361
rect 1717 -595 1954 -425
rect 3301 -361 3538 -359
rect 3301 -425 3305 -361
rect 3305 -425 3369 -361
rect 3369 -425 3511 -361
rect 3511 -425 3538 -361
rect 3301 -595 3538 -425
rect 5394 -361 5631 -359
rect 5394 -425 5456 -361
rect 5456 -425 5520 -361
rect 5520 -425 5536 -361
rect 5536 -425 5600 -361
rect 5600 -425 5616 -361
rect 5616 -425 5631 -361
rect 5394 -595 5631 -425
rect 10368 -361 10605 -359
rect 10368 -425 10430 -361
rect 10430 -425 10494 -361
rect 10494 -425 10510 -361
rect 10510 -425 10574 -361
rect 10574 -425 10590 -361
rect 10590 -425 10605 -361
rect 10368 -595 10605 -425
rect 39298 -361 39534 -359
rect 39298 -425 39342 -361
rect 39342 -425 39358 -361
rect 39358 -425 39422 -361
rect 39422 -425 39438 -361
rect 39438 -425 39502 -361
rect 39502 -425 39534 -361
rect 39298 -595 39534 -425
<< metal5 >>
rect 245 5262 565 5300
rect 245 5026 287 5262
rect 524 5026 565 5262
rect 245 2774 565 5026
rect 245 2538 287 2774
rect 524 2538 565 2774
rect 245 2499 565 2538
rect 1675 5262 1995 5300
rect 1675 5026 1717 5262
rect 1954 5026 1995 5262
rect 1675 2774 1995 5026
rect 1675 2538 1717 2774
rect 1954 2538 1995 2774
rect 1675 2499 1995 2538
rect 3259 5262 3579 5300
rect 3259 5026 3301 5262
rect 3538 5026 3579 5262
rect 3259 2774 3579 5026
rect 3259 2538 3301 2774
rect 3538 2538 3579 2774
rect 3259 2499 3579 2538
rect 5352 5262 5672 5300
rect 5352 5026 5394 5262
rect 5631 5026 5672 5262
rect 5352 2774 5672 5026
rect 5352 2538 5394 2774
rect 5631 2538 5672 2774
rect 5352 2499 5672 2538
rect 10326 5262 10646 5300
rect 10326 5026 10368 5262
rect 10605 5026 10646 5262
rect 10326 2774 10646 5026
rect 10326 2538 10368 2774
rect 10605 2538 10646 2774
rect 10326 2499 10646 2538
rect 39256 5262 39576 5300
rect 39256 5026 39298 5262
rect 39534 5026 39576 5262
rect 39256 2808 39576 5026
rect 39256 2774 39578 2808
rect 39256 2538 39298 2774
rect 39534 2538 39578 2774
rect 39256 2488 39578 2538
rect 245 2129 565 2167
rect 245 1893 287 2129
rect 524 1893 565 2129
rect 245 -359 565 1893
rect 245 -595 287 -359
rect 524 -595 565 -359
rect 245 -634 565 -595
rect 1675 2129 1995 2167
rect 1675 1893 1717 2129
rect 1954 1893 1995 2129
rect 1675 -359 1995 1893
rect 1675 -595 1717 -359
rect 1954 -595 1995 -359
rect 1675 -634 1995 -595
rect 3259 2129 3579 2167
rect 3259 1893 3301 2129
rect 3538 1893 3579 2129
rect 3259 -359 3579 1893
rect 3259 -595 3301 -359
rect 3538 -595 3579 -359
rect 3259 -634 3579 -595
rect 5352 2129 5672 2167
rect 5352 1893 5394 2129
rect 5631 1893 5672 2129
rect 5352 -359 5672 1893
rect 5352 -595 5394 -359
rect 5631 -595 5672 -359
rect 5352 -634 5672 -595
rect 10326 2129 10646 2167
rect 10326 1893 10368 2129
rect 10605 1893 10646 2129
rect 10326 -359 10646 1893
rect 10326 -595 10368 -359
rect 10605 -595 10646 -359
rect 10326 -634 10646 -595
rect 39256 2129 39576 2167
rect 39256 1893 39298 2129
rect 39534 1893 39576 2129
rect 39256 -325 39576 1893
rect 39256 -359 39578 -325
rect 39256 -595 39298 -359
rect 39534 -595 39578 -359
rect 39256 -645 39578 -595
<< labels >>
flabel metal4 -209 4434 -158 4641 0 FreeSans 480 0 0 0 t<0>
port 27 nsew
flabel poly 10608 6023 14646 6093 0 FreeSans 320 0 0 0 d<5>
port 113 nsew
flabel poly -271 5290 -201 5422 0 FreeSans 320 0 0 0 db<0>
port 117 nsew
flabel poly 657 5290 727 5422 0 FreeSans 320 0 0 0 db<1>
port 119 nsew
flabel poly 1921 5335 2375 5405 0 FreeSans 320 0 0 0 db<2>
port 121 nsew
flabel poly 3540 5335 4506 5405 0 FreeSans 320 0 0 0 db<3>
port 123 nsew
flabel metal5 245 4094 565 5026 0 FreeSans 800 0 0 0 t<1>
port 166 nsew
flabel metal5 1675 4100 1995 5026 0 FreeSans 800 0 0 0 t<2>
port 168 nsew
flabel metal5 3259 4132 3579 5026 0 FreeSans 800 0 0 0 t<3>
port 170 nsew
flabel metal5 5352 4142 5672 5026 0 FreeSans 800 0 0 0 t<4>
port 172 nsew
flabel metal5 39256 4154 39576 5026 0 FreeSans 800 0 0 0 t<6>
port 178 nsew
flabel metal4 -205 1413 -161 1543 0 FreeSans 320 0 0 0 tb<0>
port 76 nsew
flabel metal5 287 -595 524 -359 0 FreeSans 480 0 0 0 tb<1>
port 147 nsew
flabel metal5 1717 -595 1954 -359 0 FreeSans 480 0 0 0 tb<2>
port 149 nsew
flabel metal5 3301 -595 3538 -359 0 FreeSans 480 0 0 0 tb<3>
port 151 nsew
flabel metal5 5394 -595 5631 -359 0 FreeSans 480 0 0 0 tb<4>
port 153 nsew
flabel metal5 10368 -595 10605 -359 0 FreeSans 480 0 0 0 tb<5>
port 155 nsew
flabel metal5 39298 -595 39534 -359 0 FreeSans 480 0 0 0 tb<6>
port 157 nsew
flabel poly 657 5978 727 6110 0 FreeSans 320 0 0 0 d<1>
port 106 nsew
flabel poly 1409 6013 1863 6083 0 FreeSans 320 0 0 0 d<2>
port 104 nsew
flabel poly 3028 6013 3994 6083 0 FreeSans 320 0 0 0 d<3>
port 102 nsew
flabel metal5 10326 4154 10646 5026 0 FreeSans 800 0 0 0 t<5>
port 176 nsew
flabel poly 20445 6013 28579 6083 0 FreeSans 1600 0 0 0 d<6>
port 180 nsew
flabel poly 29413 5335 37547 5405 0 FreeSans 1600 0 0 0 db<6>
port 182 nsew
flabel poly 15869 5335 19907 5405 0 FreeSans 480 0 0 0 db<5>
port 184 nsew
flabel poly -271 5997 -201 6129 0 FreeSans 320 0 0 0 d<0>
port 109 nsew
flabel metal4 39154 5415 39565 6049 0 FreeSans 1600 0 0 0 VDD
port 161 nsew
flabel metal4 37909 5449 38298 6013 0 FreeSans 1600 0 0 0 VREF
port 163 nsew
flabel metal4 38589 5806 38950 6291 0 FreeSans 1600 0 0 0 VSS
port 159 nsew
flabel poly 5521 6013 7511 6083 0 FreeSans 480 0 0 0 d<4>
port 186 nsew
flabel poly 8105 5335 10095 5405 0 FreeSans 480 0 0 0 db<4>
port 188 nsew
flabel pwell 17436 439 17468 489 0 FreeSans 160 0 0 0 hgu_cdac_8bit_array_2.SUB
flabel metal4 7177 746 7228 787 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.drv<15:0>
flabel metal4 35915 746 35966 787 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.drv<63:0>
flabel metal4 12152 747 12207 786 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.drv<31:0>
flabel via4 5429 -519 5596 -436 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.tah<15:0>
flabel via4 10396 -538 10570 -438 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.tah<31:0>
flabel via4 39332 -533 39506 -433 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.tah<63:0>
flabel metal4 4022 749 4073 790 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.drv<7:0>
flabel via4 3335 -532 3509 -432 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.tah<7:0>
flabel via4 287 -595 524 -359 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.tah<1:0>
flabel metal4 966 749 1020 783 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.drv<1:0>
flabel metal4 -205 973 -156 1025 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.tah<0>
flabel metal4 -85 1097 -43 1131 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.drv<0>
flabel via4 1745 -528 1919 -428 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.tah<3:0>
flabel metal4 -75 1483 -49 1515 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.x1.CBOT
flabel metal4 -193 893 -167 925 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.x1.CTOP
flabel psubdiff -145 1149 -107 1227 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.x1.SUB
flabel psubdiff 29070 409 29112 499 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.SUB
flabel metal4 28886 485 28932 555 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.CTOP
flabel metal4 29004 1159 29050 1229 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.CTOP
flabel metal4 29126 889 29172 959 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.CBOT
flabel metal4 20532 323 20558 355 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[0].CBOT
flabel metal4 20414 -267 20440 -235 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[0].CTOP
flabel psubdiff 20462 -11 20500 67 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[0].SUB
flabel metal4 20410 1179 20436 1211 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[1].CBOT
flabel metal4 20528 1769 20554 1801 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[1].CTOP
flabel psubdiff 20468 1467 20506 1545 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[1].SUB
flabel metal4 21138 323 21164 355 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[2].CBOT
flabel metal4 21020 -267 21046 -235 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[2].CTOP
flabel psubdiff 21068 -11 21106 67 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[2].SUB
flabel metal4 21016 1179 21042 1211 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[3].CBOT
flabel metal4 21134 1769 21160 1801 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[3].CTOP
flabel psubdiff 21074 1467 21112 1545 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[3].SUB
flabel metal4 21744 323 21770 355 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[4].CBOT
flabel metal4 21626 -267 21652 -235 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[4].CTOP
flabel psubdiff 21674 -11 21712 67 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[4].SUB
flabel metal4 21622 1179 21648 1211 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[5].CBOT
flabel metal4 21740 1769 21766 1801 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[5].CTOP
flabel psubdiff 21680 1467 21718 1545 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[5].SUB
flabel metal4 22350 323 22376 355 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[6].CBOT
flabel metal4 22232 -267 22258 -235 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[6].CTOP
flabel psubdiff 22280 -11 22318 67 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[6].SUB
flabel metal4 22228 1179 22254 1211 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[7].CBOT
flabel metal4 22346 1769 22372 1801 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[7].CTOP
flabel psubdiff 22286 1467 22324 1545 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[7].SUB
flabel metal4 22956 323 22982 355 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[8].CBOT
flabel metal4 22838 -267 22864 -235 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[8].CTOP
flabel psubdiff 22886 -11 22924 67 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[8].SUB
flabel metal4 22834 1179 22860 1211 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[9].CBOT
flabel metal4 22952 1769 22978 1801 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[9].CTOP
flabel psubdiff 22892 1467 22930 1545 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[9].SUB
flabel metal4 23562 323 23588 355 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[10].CBOT
flabel metal4 23444 -267 23470 -235 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[10].CTOP
flabel psubdiff 23492 -11 23530 67 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[10].SUB
flabel metal4 23440 1179 23466 1211 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[11].CBOT
flabel metal4 23558 1769 23584 1801 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[11].CTOP
flabel psubdiff 23498 1467 23536 1545 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[11].SUB
flabel metal4 24168 323 24194 355 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[12].CBOT
flabel metal4 24050 -267 24076 -235 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[12].CTOP
flabel psubdiff 24098 -11 24136 67 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[12].SUB
flabel metal4 24046 1179 24072 1211 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[13].CBOT
flabel metal4 24164 1769 24190 1801 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[13].CTOP
flabel psubdiff 24104 1467 24142 1545 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[13].SUB
flabel metal4 24774 323 24800 355 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[14].CBOT
flabel metal4 24656 -267 24682 -235 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[14].CTOP
flabel psubdiff 24704 -11 24742 67 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[14].SUB
flabel metal4 24652 1179 24678 1211 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[15].CBOT
flabel metal4 24770 1769 24796 1801 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[15].CTOP
flabel psubdiff 24710 1467 24748 1545 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[15].SUB
flabel metal4 25380 323 25406 355 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[16].CBOT
flabel metal4 25262 -267 25288 -235 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[16].CTOP
flabel psubdiff 25310 -11 25348 67 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[16].SUB
flabel metal4 25258 1179 25284 1211 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[17].CBOT
flabel metal4 25376 1769 25402 1801 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[17].CTOP
flabel psubdiff 25316 1467 25354 1545 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[17].SUB
flabel metal4 25986 323 26012 355 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[18].CBOT
flabel metal4 25868 -267 25894 -235 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[18].CTOP
flabel psubdiff 25916 -11 25954 67 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[18].SUB
flabel metal4 25864 1179 25890 1211 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[19].CBOT
flabel metal4 25982 1769 26008 1801 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[19].CTOP
flabel psubdiff 25922 1467 25960 1545 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[19].SUB
flabel metal4 26592 323 26618 355 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[20].CBOT
flabel metal4 26474 -267 26500 -235 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[20].CTOP
flabel psubdiff 26522 -11 26560 67 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[20].SUB
flabel metal4 26470 1179 26496 1211 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[21].CBOT
flabel metal4 26588 1769 26614 1801 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[21].CTOP
flabel psubdiff 26528 1467 26566 1545 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[21].SUB
flabel metal4 27198 323 27224 355 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[22].CBOT
flabel metal4 27080 -267 27106 -235 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[22].CTOP
flabel psubdiff 27128 -11 27166 67 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[22].SUB
flabel metal4 27076 1179 27102 1211 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[23].CBOT
flabel metal4 27194 1769 27220 1801 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[23].CTOP
flabel psubdiff 27134 1467 27172 1545 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[23].SUB
flabel metal4 27804 323 27830 355 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[24].CBOT
flabel metal4 27686 -267 27712 -235 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[24].CTOP
flabel psubdiff 27734 -11 27772 67 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[24].SUB
flabel metal4 27682 1179 27708 1211 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[25].CBOT
flabel metal4 27800 1769 27826 1801 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[25].CTOP
flabel psubdiff 27740 1467 27778 1545 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[25].SUB
flabel metal4 28410 323 28436 355 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[26].CBOT
flabel metal4 28292 -267 28318 -235 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[26].CTOP
flabel psubdiff 28340 -11 28378 67 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[26].SUB
flabel metal4 28288 1179 28314 1211 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[27].CBOT
flabel metal4 28406 1769 28432 1801 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[27].CTOP
flabel psubdiff 28346 1467 28384 1545 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[27].SUB
flabel metal4 29016 323 29042 355 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[28].CBOT
flabel metal4 28898 -267 28924 -235 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[28].CTOP
flabel psubdiff 28946 -11 28984 67 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[28].SUB
flabel metal4 28894 1179 28920 1211 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[29].CBOT
flabel metal4 29012 1769 29038 1801 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[29].CTOP
flabel psubdiff 28952 1467 28990 1545 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[29].SUB
flabel metal4 29622 323 29648 355 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[30].CBOT
flabel metal4 29504 -267 29530 -235 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[30].CTOP
flabel psubdiff 29552 -11 29590 67 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[30].SUB
flabel metal4 29500 1179 29526 1211 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[31].CBOT
flabel metal4 29618 1769 29644 1801 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[31].CTOP
flabel psubdiff 29558 1467 29596 1545 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[31].SUB
flabel metal4 30228 323 30254 355 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[32].CBOT
flabel metal4 30110 -267 30136 -235 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[32].CTOP
flabel psubdiff 30158 -11 30196 67 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[32].SUB
flabel metal4 30106 1179 30132 1211 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[33].CBOT
flabel metal4 30224 1769 30250 1801 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[33].CTOP
flabel psubdiff 30164 1467 30202 1545 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[33].SUB
flabel metal4 30834 323 30860 355 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[34].CBOT
flabel metal4 30716 -267 30742 -235 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[34].CTOP
flabel psubdiff 30764 -11 30802 67 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[34].SUB
flabel metal4 30712 1179 30738 1211 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[35].CBOT
flabel metal4 30830 1769 30856 1801 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[35].CTOP
flabel psubdiff 30770 1467 30808 1545 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[35].SUB
flabel metal4 31440 323 31466 355 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[36].CBOT
flabel metal4 31322 -267 31348 -235 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[36].CTOP
flabel psubdiff 31370 -11 31408 67 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[36].SUB
flabel metal4 31318 1179 31344 1211 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[37].CBOT
flabel metal4 31436 1769 31462 1801 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[37].CTOP
flabel psubdiff 31376 1467 31414 1545 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[37].SUB
flabel metal4 32046 323 32072 355 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[38].CBOT
flabel metal4 31928 -267 31954 -235 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[38].CTOP
flabel psubdiff 31976 -11 32014 67 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[38].SUB
flabel metal4 31924 1179 31950 1211 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[39].CBOT
flabel metal4 32042 1769 32068 1801 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[39].CTOP
flabel psubdiff 31982 1467 32020 1545 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[39].SUB
flabel metal4 32652 323 32678 355 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[40].CBOT
flabel metal4 32534 -267 32560 -235 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[40].CTOP
flabel psubdiff 32582 -11 32620 67 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[40].SUB
flabel metal4 32530 1179 32556 1211 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[41].CBOT
flabel metal4 32648 1769 32674 1801 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[41].CTOP
flabel psubdiff 32588 1467 32626 1545 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[41].SUB
flabel metal4 33258 323 33284 355 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[42].CBOT
flabel metal4 33140 -267 33166 -235 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[42].CTOP
flabel psubdiff 33188 -11 33226 67 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[42].SUB
flabel metal4 33136 1179 33162 1211 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[43].CBOT
flabel metal4 33254 1769 33280 1801 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[43].CTOP
flabel psubdiff 33194 1467 33232 1545 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[43].SUB
flabel metal4 33864 323 33890 355 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[44].CBOT
flabel metal4 33746 -267 33772 -235 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[44].CTOP
flabel psubdiff 33794 -11 33832 67 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[44].SUB
flabel metal4 33742 1179 33768 1211 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[45].CBOT
flabel metal4 33860 1769 33886 1801 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[45].CTOP
flabel psubdiff 33800 1467 33838 1545 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[45].SUB
flabel metal4 34470 323 34496 355 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[46].CBOT
flabel metal4 34352 -267 34378 -235 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[46].CTOP
flabel psubdiff 34400 -11 34438 67 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[46].SUB
flabel metal4 34348 1179 34374 1211 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[47].CBOT
flabel metal4 34466 1769 34492 1801 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[47].CTOP
flabel psubdiff 34406 1467 34444 1545 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[47].SUB
flabel metal4 35076 323 35102 355 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[48].CBOT
flabel metal4 34958 -267 34984 -235 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[48].CTOP
flabel psubdiff 35006 -11 35044 67 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[48].SUB
flabel metal4 34954 1179 34980 1211 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[49].CBOT
flabel metal4 35072 1769 35098 1801 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[49].CTOP
flabel psubdiff 35012 1467 35050 1545 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[49].SUB
flabel metal4 35682 323 35708 355 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[50].CBOT
flabel metal4 35564 -267 35590 -235 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[50].CTOP
flabel psubdiff 35612 -11 35650 67 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[50].SUB
flabel metal4 35560 1179 35586 1211 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[51].CBOT
flabel metal4 35678 1769 35704 1801 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[51].CTOP
flabel psubdiff 35618 1467 35656 1545 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[51].SUB
flabel metal4 36288 323 36314 355 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[52].CBOT
flabel metal4 36170 -267 36196 -235 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[52].CTOP
flabel psubdiff 36218 -11 36256 67 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[52].SUB
flabel metal4 36166 1179 36192 1211 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[53].CBOT
flabel metal4 36284 1769 36310 1801 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[53].CTOP
flabel psubdiff 36224 1467 36262 1545 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[53].SUB
flabel metal4 36894 323 36920 355 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[54].CBOT
flabel metal4 36776 -267 36802 -235 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[54].CTOP
flabel psubdiff 36824 -11 36862 67 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[54].SUB
flabel metal4 36772 1179 36798 1211 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[55].CBOT
flabel metal4 36890 1769 36916 1801 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[55].CTOP
flabel psubdiff 36830 1467 36868 1545 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[55].SUB
flabel metal4 37500 323 37526 355 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[56].CBOT
flabel metal4 37382 -267 37408 -235 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[56].CTOP
flabel psubdiff 37430 -11 37468 67 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[56].SUB
flabel metal4 37378 1179 37404 1211 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[57].CBOT
flabel metal4 37496 1769 37522 1801 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[57].CTOP
flabel psubdiff 37436 1467 37474 1545 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[57].SUB
flabel metal4 38106 323 38132 355 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[58].CBOT
flabel metal4 37988 -267 38014 -235 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[58].CTOP
flabel psubdiff 38036 -11 38074 67 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[58].SUB
flabel metal4 37984 1179 38010 1211 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[59].CBOT
flabel metal4 38102 1769 38128 1801 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[59].CTOP
flabel psubdiff 38042 1467 38080 1545 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[59].SUB
flabel metal4 38712 323 38738 355 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[60].CBOT
flabel metal4 38594 -267 38620 -235 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[60].CTOP
flabel psubdiff 38642 -11 38680 67 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[60].SUB
flabel metal4 38590 1179 38616 1211 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[61].CBOT
flabel metal4 38708 1769 38734 1801 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[61].CTOP
flabel psubdiff 38648 1467 38686 1545 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[61].SUB
flabel metal4 39318 323 39344 355 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[62].CBOT
flabel metal4 39200 -267 39226 -235 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[62].CTOP
flabel psubdiff 39248 -11 39286 67 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[62].SUB
flabel metal4 39196 1179 39222 1211 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[63].CBOT
flabel metal4 39314 1769 39340 1801 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[63].CTOP
flabel psubdiff 39254 1467 39292 1545 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[63].SUB
flabel psubdiff 14766 621 14810 713 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.SUB
flabel metal4 14336 417 14380 509 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.CBOT
flabel metal4 14824 421 14868 513 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.CTOP
flabel metal4 14702 941 14746 1033 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.CTOP
flabel metal4 10588 1179 10614 1211 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[0].CBOT
flabel metal4 10706 1769 10732 1801 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[0].CTOP
flabel psubdiff 10646 1467 10684 1545 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[0].SUB
flabel metal4 10710 323 10736 355 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[1].CBOT
flabel metal4 10592 -267 10618 -235 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[1].CTOP
flabel psubdiff 10640 -11 10678 67 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[1].SUB
flabel metal4 11194 1179 11220 1211 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[2].CBOT
flabel metal4 11312 1769 11338 1801 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[2].CTOP
flabel psubdiff 11252 1467 11290 1545 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[2].SUB
flabel metal4 11316 323 11342 355 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[3].CBOT
flabel metal4 11198 -267 11224 -235 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[3].CTOP
flabel psubdiff 11246 -11 11284 67 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[3].SUB
flabel metal4 11800 1179 11826 1211 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[4].CBOT
flabel metal4 11918 1769 11944 1801 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[4].CTOP
flabel psubdiff 11858 1467 11896 1545 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[4].SUB
flabel metal4 11922 323 11948 355 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[5].CBOT
flabel metal4 11804 -267 11830 -235 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[5].CTOP
flabel psubdiff 11852 -11 11890 67 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[5].SUB
flabel metal4 12406 1179 12432 1211 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[6].CBOT
flabel metal4 12524 1769 12550 1801 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[6].CTOP
flabel psubdiff 12464 1467 12502 1545 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[6].SUB
flabel metal4 12528 323 12554 355 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[7].CBOT
flabel metal4 12410 -267 12436 -235 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[7].CTOP
flabel psubdiff 12458 -11 12496 67 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[7].SUB
flabel metal4 13012 1179 13038 1211 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[8].CBOT
flabel metal4 13130 1769 13156 1801 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[8].CTOP
flabel psubdiff 13070 1467 13108 1545 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[8].SUB
flabel metal4 13134 323 13160 355 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[9].CBOT
flabel metal4 13016 -267 13042 -235 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[9].CTOP
flabel psubdiff 13064 -11 13102 67 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[9].SUB
flabel metal4 13618 1179 13644 1211 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[10].CBOT
flabel metal4 13736 1769 13762 1801 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[10].CTOP
flabel psubdiff 13676 1467 13714 1545 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[10].SUB
flabel metal4 13740 323 13766 355 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[11].CBOT
flabel metal4 13622 -267 13648 -235 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[11].CTOP
flabel psubdiff 13670 -11 13708 67 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[11].SUB
flabel metal4 14224 1179 14250 1211 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[12].CBOT
flabel metal4 14342 1769 14368 1801 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[12].CTOP
flabel psubdiff 14282 1467 14320 1545 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[12].SUB
flabel metal4 14346 323 14372 355 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[13].CBOT
flabel metal4 14228 -267 14254 -235 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[13].CTOP
flabel psubdiff 14276 -11 14314 67 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[13].SUB
flabel metal4 14830 1179 14856 1211 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[14].CBOT
flabel metal4 14948 1769 14974 1801 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[14].CTOP
flabel psubdiff 14888 1467 14926 1545 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[14].SUB
flabel metal4 14952 323 14978 355 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[15].CBOT
flabel metal4 14834 -267 14860 -235 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[15].CTOP
flabel psubdiff 14882 -11 14920 67 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[15].SUB
flabel metal4 15436 1179 15462 1211 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[16].CBOT
flabel metal4 15554 1769 15580 1801 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[16].CTOP
flabel psubdiff 15494 1467 15532 1545 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[16].SUB
flabel metal4 15558 323 15584 355 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[17].CBOT
flabel metal4 15440 -267 15466 -235 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[17].CTOP
flabel psubdiff 15488 -11 15526 67 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[17].SUB
flabel metal4 16042 1179 16068 1211 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[18].CBOT
flabel metal4 16160 1769 16186 1801 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[18].CTOP
flabel psubdiff 16100 1467 16138 1545 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[18].SUB
flabel metal4 16164 323 16190 355 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[19].CBOT
flabel metal4 16046 -267 16072 -235 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[19].CTOP
flabel psubdiff 16094 -11 16132 67 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[19].SUB
flabel metal4 16648 1179 16674 1211 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[20].CBOT
flabel metal4 16766 1769 16792 1801 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[20].CTOP
flabel psubdiff 16706 1467 16744 1545 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[20].SUB
flabel metal4 16770 323 16796 355 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[21].CBOT
flabel metal4 16652 -267 16678 -235 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[21].CTOP
flabel psubdiff 16700 -11 16738 67 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[21].SUB
flabel metal4 17254 1179 17280 1211 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[22].CBOT
flabel metal4 17372 1769 17398 1801 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[22].CTOP
flabel psubdiff 17312 1467 17350 1545 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[22].SUB
flabel metal4 17376 323 17402 355 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[23].CBOT
flabel metal4 17258 -267 17284 -235 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[23].CTOP
flabel psubdiff 17306 -11 17344 67 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[23].SUB
flabel metal4 17860 1179 17886 1211 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[24].CBOT
flabel metal4 17978 1769 18004 1801 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[24].CTOP
flabel psubdiff 17918 1467 17956 1545 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[24].SUB
flabel metal4 17982 323 18008 355 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[25].CBOT
flabel metal4 17864 -267 17890 -235 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[25].CTOP
flabel psubdiff 17912 -11 17950 67 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[25].SUB
flabel metal4 18466 1179 18492 1211 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[26].CBOT
flabel metal4 18584 1769 18610 1801 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[26].CTOP
flabel psubdiff 18524 1467 18562 1545 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[26].SUB
flabel metal4 18588 323 18614 355 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[27].CBOT
flabel metal4 18470 -267 18496 -235 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[27].CTOP
flabel psubdiff 18518 -11 18556 67 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[27].SUB
flabel metal4 19072 1179 19098 1211 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[28].CBOT
flabel metal4 19190 1769 19216 1801 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[28].CTOP
flabel psubdiff 19130 1467 19168 1545 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[28].SUB
flabel metal4 19194 323 19220 355 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[29].CBOT
flabel metal4 19076 -267 19102 -235 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[29].CTOP
flabel psubdiff 19124 -11 19162 67 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[29].SUB
flabel metal4 19678 1179 19704 1211 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[30].CBOT
flabel metal4 19796 1769 19822 1801 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[30].CTOP
flabel psubdiff 19736 1467 19774 1545 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[30].SUB
flabel metal4 19800 323 19826 355 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[31].CBOT
flabel metal4 19682 -267 19708 -235 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[31].CTOP
flabel psubdiff 19730 -11 19768 67 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[31].SUB
flabel metal4 8156 583 8192 663 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.CBOT
flabel metal4 7432 553 7468 633 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.CTOP
flabel metal4 7546 925 7590 1007 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.CTOP
flabel psubdiff 7850 825 7894 907 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.SUB
flabel metal4 5614 1179 5640 1211 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[0].CBOT
flabel metal4 5732 1769 5758 1801 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[0].CTOP
flabel psubdiff 5672 1467 5710 1545 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[0].SUB
flabel metal4 5736 323 5762 355 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[1].CBOT
flabel metal4 5618 -267 5644 -235 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[1].CTOP
flabel psubdiff 5666 -11 5704 67 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[1].SUB
flabel metal4 6220 1179 6246 1211 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[2].CBOT
flabel metal4 6338 1769 6364 1801 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[2].CTOP
flabel psubdiff 6278 1467 6316 1545 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[2].SUB
flabel metal4 6342 323 6368 355 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[3].CBOT
flabel metal4 6224 -267 6250 -235 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[3].CTOP
flabel psubdiff 6272 -11 6310 67 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[3].SUB
flabel metal4 6826 1179 6852 1211 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[4].CBOT
flabel metal4 6944 1769 6970 1801 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[4].CTOP
flabel psubdiff 6884 1467 6922 1545 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[4].SUB
flabel metal4 6948 323 6974 355 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[5].CBOT
flabel metal4 6830 -267 6856 -235 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[5].CTOP
flabel psubdiff 6878 -11 6916 67 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[5].SUB
flabel metal4 7432 1179 7458 1211 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[6].CBOT
flabel metal4 7550 1769 7576 1801 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[6].CTOP
flabel psubdiff 7490 1467 7528 1545 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[6].SUB
flabel metal4 7554 323 7580 355 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[7].CBOT
flabel metal4 7436 -267 7462 -235 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[7].CTOP
flabel psubdiff 7484 -11 7522 67 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[7].SUB
flabel metal4 8038 1179 8064 1211 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[8].CBOT
flabel metal4 8156 1769 8182 1801 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[8].CTOP
flabel psubdiff 8096 1467 8134 1545 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[8].SUB
flabel metal4 8160 323 8186 355 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[9].CBOT
flabel metal4 8042 -267 8068 -235 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[9].CTOP
flabel psubdiff 8090 -11 8128 67 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[9].SUB
flabel metal4 8644 1179 8670 1211 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[10].CBOT
flabel metal4 8762 1769 8788 1801 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[10].CTOP
flabel psubdiff 8702 1467 8740 1545 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[10].SUB
flabel metal4 8766 323 8792 355 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[11].CBOT
flabel metal4 8648 -267 8674 -235 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[11].CTOP
flabel psubdiff 8696 -11 8734 67 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[11].SUB
flabel metal4 9250 1179 9276 1211 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[12].CBOT
flabel metal4 9368 1769 9394 1801 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[12].CTOP
flabel psubdiff 9308 1467 9346 1545 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[12].SUB
flabel metal4 9372 323 9398 355 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[13].CBOT
flabel metal4 9254 -267 9280 -235 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[13].CTOP
flabel psubdiff 9302 -11 9340 67 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[13].SUB
flabel metal4 9856 1179 9882 1211 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[14].CBOT
flabel metal4 9974 1769 10000 1801 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[14].CTOP
flabel psubdiff 9914 1467 9952 1545 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[14].SUB
flabel metal4 9978 323 10004 355 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[15].CBOT
flabel metal4 9860 -267 9886 -235 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[15].CTOP
flabel psubdiff 9908 -11 9946 67 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[15].SUB
flabel psubdiff 4207 621 4251 721 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_8_0.SUB
flabel metal4 4387 453 4433 545 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_8_0.CBOT
flabel metal4 3659 475 3705 567 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_8_0.CTOP
flabel metal4 3787 1313 3827 1397 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_8_0.CTOP
flabel metal4 5003 323 5029 355 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_8_0.x1[7].CBOT
flabel metal4 4885 -267 4911 -235 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_8_0.x1[7].CTOP
flabel psubdiff 4933 -11 4971 67 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_8_0.x1[7].SUB
flabel metal4 4881 1179 4907 1211 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_8_0.x1[6].CBOT
flabel metal4 4999 1769 5025 1801 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_8_0.x1[6].CTOP
flabel psubdiff 4939 1467 4977 1545 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_8_0.x1[6].SUB
flabel metal4 4397 323 4423 355 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_8_0.x1[5].CBOT
flabel metal4 4279 -267 4305 -235 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_8_0.x1[5].CTOP
flabel psubdiff 4327 -11 4365 67 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_8_0.x1[5].SUB
flabel metal4 4275 1179 4301 1211 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_8_0.x1[4].CBOT
flabel metal4 4393 1769 4419 1801 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_8_0.x1[4].CTOP
flabel psubdiff 4333 1467 4371 1545 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_8_0.x1[4].SUB
flabel metal4 3791 323 3817 355 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_8_0.x1[3].CBOT
flabel metal4 3673 -267 3699 -235 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_8_0.x1[3].CTOP
flabel psubdiff 3721 -11 3759 67 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_8_0.x1[3].SUB
flabel metal4 3669 1179 3695 1211 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_8_0.x1[2].CBOT
flabel metal4 3787 1769 3813 1801 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_8_0.x1[2].CTOP
flabel psubdiff 3727 1467 3765 1545 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_8_0.x1[2].SUB
flabel metal4 3185 323 3211 355 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_8_0.x1[1].CBOT
flabel metal4 3067 -267 3093 -235 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_8_0.x1[1].CTOP
flabel psubdiff 3115 -11 3153 67 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_8_0.x1[1].SUB
flabel metal4 3063 1179 3089 1211 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_8_0.x1[0].CBOT
flabel metal4 3181 1769 3207 1801 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_8_0.x1[0].CTOP
flabel psubdiff 3121 1467 3159 1545 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_8_0.x1[0].SUB
flabel metal4 2245 681 2297 721 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT
flabel metal4 1519 565 1571 605 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CTOP
flabel psubdiff 2069 575 2109 685 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.SUB
flabel metal4 1643 903 1681 985 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CTOP
flabel metal4 2257 323 2283 355 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.x1[3].CBOT
flabel metal4 2139 -267 2165 -235 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.x1[3].CTOP
flabel psubdiff 2187 -11 2225 67 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.x1[3].SUB
flabel metal4 2135 1179 2161 1211 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.x1[2].CBOT
flabel metal4 2253 1769 2279 1801 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.x1[2].CTOP
flabel psubdiff 2193 1467 2231 1545 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.x1[2].SUB
flabel metal4 1651 323 1677 355 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.x1[1].CBOT
flabel metal4 1533 -267 1559 -235 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.x1[1].CTOP
flabel psubdiff 1581 -11 1619 67 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.x1[1].SUB
flabel metal4 1529 1179 1555 1211 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.x1[0].CBOT
flabel metal4 1647 1769 1673 1801 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.x1[0].CTOP
flabel psubdiff 1587 1467 1625 1545 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.x1[0].SUB
flabel psubdiff 669 482 717 596 0 FreeSans 160 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_2_0.SUB
flabel metal4 733 477 769 567 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_2_0.CBOT
flabel metal4 613 35 649 137 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_2_0.CTOP
flabel metal4 731 1619 771 1697 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_2_0.CTOP
flabel metal4 739 323 765 355 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_2_0.x2.CBOT
flabel metal4 621 -267 647 -235 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_2_0.x2.CTOP
flabel psubdiff 669 -11 707 67 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_2_0.x2.SUB
flabel metal4 617 1179 643 1211 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_2_0.x1.CBOT
flabel metal4 735 1769 761 1801 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_2_0.x1.CTOP
flabel psubdiff 675 1467 713 1545 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_2_0.x1.SUB
flabel metal4 -197 19 -171 51 0 FreeSans 320 0 0 0 hgu_cdac_unit_0.CBOT
flabel metal4 -79 609 -53 641 0 FreeSans 320 0 0 0 hgu_cdac_unit_0.CTOP
flabel psubdiff -139 307 -101 385 0 FreeSans 320 0 0 0 hgu_cdac_unit_0.SUB
flabel pwell 17436 3572 17468 3622 0 FreeSans 160 0 0 0 hgu_cdac_8bit_array_3.SUB
flabel metal4 7177 3879 7228 3920 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.drv<15:0>
flabel metal4 35915 3879 35966 3920 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.drv<63:0>
flabel metal4 12152 3880 12207 3919 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.drv<31:0>
flabel via4 5429 2614 5596 2697 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.tah<15:0>
flabel via4 10396 2595 10570 2695 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.tah<31:0>
flabel via4 39332 2600 39506 2700 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.tah<63:0>
flabel metal4 4022 3882 4073 3923 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.drv<7:0>
flabel via4 3335 2601 3509 2701 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.tah<7:0>
flabel via4 287 2538 524 2774 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.tah<1:0>
flabel metal4 966 3882 1020 3916 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.drv<1:0>
flabel metal4 -205 4106 -156 4158 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.tah<0>
flabel metal4 -85 4230 -43 4264 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.drv<0>
flabel via4 1745 2605 1919 2705 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.tah<3:0>
flabel metal4 -75 4616 -49 4648 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.x1.CBOT
flabel metal4 -193 4026 -167 4058 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.x1.CTOP
flabel psubdiff -145 4282 -107 4360 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.x1.SUB
flabel psubdiff 29070 3542 29112 3632 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.SUB
flabel metal4 28886 3618 28932 3688 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.CTOP
flabel metal4 29004 4292 29050 4362 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.CTOP
flabel metal4 29126 4022 29172 4092 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.CBOT
flabel metal4 20532 3456 20558 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[0].CBOT
flabel metal4 20414 2866 20440 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[0].CTOP
flabel psubdiff 20462 3122 20500 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[0].SUB
flabel metal4 20410 4312 20436 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[1].CBOT
flabel metal4 20528 4902 20554 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[1].CTOP
flabel psubdiff 20468 4600 20506 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[1].SUB
flabel metal4 21138 3456 21164 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[2].CBOT
flabel metal4 21020 2866 21046 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[2].CTOP
flabel psubdiff 21068 3122 21106 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[2].SUB
flabel metal4 21016 4312 21042 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[3].CBOT
flabel metal4 21134 4902 21160 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[3].CTOP
flabel psubdiff 21074 4600 21112 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[3].SUB
flabel metal4 21744 3456 21770 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[4].CBOT
flabel metal4 21626 2866 21652 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[4].CTOP
flabel psubdiff 21674 3122 21712 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[4].SUB
flabel metal4 21622 4312 21648 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[5].CBOT
flabel metal4 21740 4902 21766 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[5].CTOP
flabel psubdiff 21680 4600 21718 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[5].SUB
flabel metal4 22350 3456 22376 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[6].CBOT
flabel metal4 22232 2866 22258 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[6].CTOP
flabel psubdiff 22280 3122 22318 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[6].SUB
flabel metal4 22228 4312 22254 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[7].CBOT
flabel metal4 22346 4902 22372 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[7].CTOP
flabel psubdiff 22286 4600 22324 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[7].SUB
flabel metal4 22956 3456 22982 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[8].CBOT
flabel metal4 22838 2866 22864 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[8].CTOP
flabel psubdiff 22886 3122 22924 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[8].SUB
flabel metal4 22834 4312 22860 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[9].CBOT
flabel metal4 22952 4902 22978 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[9].CTOP
flabel psubdiff 22892 4600 22930 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[9].SUB
flabel metal4 23562 3456 23588 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[10].CBOT
flabel metal4 23444 2866 23470 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[10].CTOP
flabel psubdiff 23492 3122 23530 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[10].SUB
flabel metal4 23440 4312 23466 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[11].CBOT
flabel metal4 23558 4902 23584 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[11].CTOP
flabel psubdiff 23498 4600 23536 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[11].SUB
flabel metal4 24168 3456 24194 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[12].CBOT
flabel metal4 24050 2866 24076 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[12].CTOP
flabel psubdiff 24098 3122 24136 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[12].SUB
flabel metal4 24046 4312 24072 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[13].CBOT
flabel metal4 24164 4902 24190 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[13].CTOP
flabel psubdiff 24104 4600 24142 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[13].SUB
flabel metal4 24774 3456 24800 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[14].CBOT
flabel metal4 24656 2866 24682 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[14].CTOP
flabel psubdiff 24704 3122 24742 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[14].SUB
flabel metal4 24652 4312 24678 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[15].CBOT
flabel metal4 24770 4902 24796 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[15].CTOP
flabel psubdiff 24710 4600 24748 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[15].SUB
flabel metal4 25380 3456 25406 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[16].CBOT
flabel metal4 25262 2866 25288 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[16].CTOP
flabel psubdiff 25310 3122 25348 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[16].SUB
flabel metal4 25258 4312 25284 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[17].CBOT
flabel metal4 25376 4902 25402 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[17].CTOP
flabel psubdiff 25316 4600 25354 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[17].SUB
flabel metal4 25986 3456 26012 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[18].CBOT
flabel metal4 25868 2866 25894 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[18].CTOP
flabel psubdiff 25916 3122 25954 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[18].SUB
flabel metal4 25864 4312 25890 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[19].CBOT
flabel metal4 25982 4902 26008 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[19].CTOP
flabel psubdiff 25922 4600 25960 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[19].SUB
flabel metal4 26592 3456 26618 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[20].CBOT
flabel metal4 26474 2866 26500 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[20].CTOP
flabel psubdiff 26522 3122 26560 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[20].SUB
flabel metal4 26470 4312 26496 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[21].CBOT
flabel metal4 26588 4902 26614 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[21].CTOP
flabel psubdiff 26528 4600 26566 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[21].SUB
flabel metal4 27198 3456 27224 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[22].CBOT
flabel metal4 27080 2866 27106 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[22].CTOP
flabel psubdiff 27128 3122 27166 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[22].SUB
flabel metal4 27076 4312 27102 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[23].CBOT
flabel metal4 27194 4902 27220 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[23].CTOP
flabel psubdiff 27134 4600 27172 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[23].SUB
flabel metal4 27804 3456 27830 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[24].CBOT
flabel metal4 27686 2866 27712 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[24].CTOP
flabel psubdiff 27734 3122 27772 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[24].SUB
flabel metal4 27682 4312 27708 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[25].CBOT
flabel metal4 27800 4902 27826 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[25].CTOP
flabel psubdiff 27740 4600 27778 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[25].SUB
flabel metal4 28410 3456 28436 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[26].CBOT
flabel metal4 28292 2866 28318 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[26].CTOP
flabel psubdiff 28340 3122 28378 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[26].SUB
flabel metal4 28288 4312 28314 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[27].CBOT
flabel metal4 28406 4902 28432 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[27].CTOP
flabel psubdiff 28346 4600 28384 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[27].SUB
flabel metal4 29016 3456 29042 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[28].CBOT
flabel metal4 28898 2866 28924 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[28].CTOP
flabel psubdiff 28946 3122 28984 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[28].SUB
flabel metal4 28894 4312 28920 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[29].CBOT
flabel metal4 29012 4902 29038 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[29].CTOP
flabel psubdiff 28952 4600 28990 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[29].SUB
flabel metal4 29622 3456 29648 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[30].CBOT
flabel metal4 29504 2866 29530 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[30].CTOP
flabel psubdiff 29552 3122 29590 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[30].SUB
flabel metal4 29500 4312 29526 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[31].CBOT
flabel metal4 29618 4902 29644 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[31].CTOP
flabel psubdiff 29558 4600 29596 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[31].SUB
flabel metal4 30228 3456 30254 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[32].CBOT
flabel metal4 30110 2866 30136 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[32].CTOP
flabel psubdiff 30158 3122 30196 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[32].SUB
flabel metal4 30106 4312 30132 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[33].CBOT
flabel metal4 30224 4902 30250 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[33].CTOP
flabel psubdiff 30164 4600 30202 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[33].SUB
flabel metal4 30834 3456 30860 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[34].CBOT
flabel metal4 30716 2866 30742 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[34].CTOP
flabel psubdiff 30764 3122 30802 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[34].SUB
flabel metal4 30712 4312 30738 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[35].CBOT
flabel metal4 30830 4902 30856 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[35].CTOP
flabel psubdiff 30770 4600 30808 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[35].SUB
flabel metal4 31440 3456 31466 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[36].CBOT
flabel metal4 31322 2866 31348 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[36].CTOP
flabel psubdiff 31370 3122 31408 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[36].SUB
flabel metal4 31318 4312 31344 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[37].CBOT
flabel metal4 31436 4902 31462 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[37].CTOP
flabel psubdiff 31376 4600 31414 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[37].SUB
flabel metal4 32046 3456 32072 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[38].CBOT
flabel metal4 31928 2866 31954 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[38].CTOP
flabel psubdiff 31976 3122 32014 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[38].SUB
flabel metal4 31924 4312 31950 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[39].CBOT
flabel metal4 32042 4902 32068 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[39].CTOP
flabel psubdiff 31982 4600 32020 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[39].SUB
flabel metal4 32652 3456 32678 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[40].CBOT
flabel metal4 32534 2866 32560 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[40].CTOP
flabel psubdiff 32582 3122 32620 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[40].SUB
flabel metal4 32530 4312 32556 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[41].CBOT
flabel metal4 32648 4902 32674 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[41].CTOP
flabel psubdiff 32588 4600 32626 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[41].SUB
flabel metal4 33258 3456 33284 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[42].CBOT
flabel metal4 33140 2866 33166 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[42].CTOP
flabel psubdiff 33188 3122 33226 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[42].SUB
flabel metal4 33136 4312 33162 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[43].CBOT
flabel metal4 33254 4902 33280 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[43].CTOP
flabel psubdiff 33194 4600 33232 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[43].SUB
flabel metal4 33864 3456 33890 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[44].CBOT
flabel metal4 33746 2866 33772 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[44].CTOP
flabel psubdiff 33794 3122 33832 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[44].SUB
flabel metal4 33742 4312 33768 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[45].CBOT
flabel metal4 33860 4902 33886 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[45].CTOP
flabel psubdiff 33800 4600 33838 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[45].SUB
flabel metal4 34470 3456 34496 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[46].CBOT
flabel metal4 34352 2866 34378 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[46].CTOP
flabel psubdiff 34400 3122 34438 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[46].SUB
flabel metal4 34348 4312 34374 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[47].CBOT
flabel metal4 34466 4902 34492 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[47].CTOP
flabel psubdiff 34406 4600 34444 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[47].SUB
flabel metal4 35076 3456 35102 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[48].CBOT
flabel metal4 34958 2866 34984 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[48].CTOP
flabel psubdiff 35006 3122 35044 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[48].SUB
flabel metal4 34954 4312 34980 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[49].CBOT
flabel metal4 35072 4902 35098 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[49].CTOP
flabel psubdiff 35012 4600 35050 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[49].SUB
flabel metal4 35682 3456 35708 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[50].CBOT
flabel metal4 35564 2866 35590 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[50].CTOP
flabel psubdiff 35612 3122 35650 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[50].SUB
flabel metal4 35560 4312 35586 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[51].CBOT
flabel metal4 35678 4902 35704 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[51].CTOP
flabel psubdiff 35618 4600 35656 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[51].SUB
flabel metal4 36288 3456 36314 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[52].CBOT
flabel metal4 36170 2866 36196 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[52].CTOP
flabel psubdiff 36218 3122 36256 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[52].SUB
flabel metal4 36166 4312 36192 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[53].CBOT
flabel metal4 36284 4902 36310 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[53].CTOP
flabel psubdiff 36224 4600 36262 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[53].SUB
flabel metal4 36894 3456 36920 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[54].CBOT
flabel metal4 36776 2866 36802 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[54].CTOP
flabel psubdiff 36824 3122 36862 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[54].SUB
flabel metal4 36772 4312 36798 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[55].CBOT
flabel metal4 36890 4902 36916 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[55].CTOP
flabel psubdiff 36830 4600 36868 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[55].SUB
flabel metal4 37500 3456 37526 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[56].CBOT
flabel metal4 37382 2866 37408 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[56].CTOP
flabel psubdiff 37430 3122 37468 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[56].SUB
flabel metal4 37378 4312 37404 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[57].CBOT
flabel metal4 37496 4902 37522 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[57].CTOP
flabel psubdiff 37436 4600 37474 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[57].SUB
flabel metal4 38106 3456 38132 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[58].CBOT
flabel metal4 37988 2866 38014 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[58].CTOP
flabel psubdiff 38036 3122 38074 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[58].SUB
flabel metal4 37984 4312 38010 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[59].CBOT
flabel metal4 38102 4902 38128 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[59].CTOP
flabel psubdiff 38042 4600 38080 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[59].SUB
flabel metal4 38712 3456 38738 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[60].CBOT
flabel metal4 38594 2866 38620 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[60].CTOP
flabel psubdiff 38642 3122 38680 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[60].SUB
flabel metal4 38590 4312 38616 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[61].CBOT
flabel metal4 38708 4902 38734 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[61].CTOP
flabel psubdiff 38648 4600 38686 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[61].SUB
flabel metal4 39318 3456 39344 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[62].CBOT
flabel metal4 39200 2866 39226 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[62].CTOP
flabel psubdiff 39248 3122 39286 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[62].SUB
flabel metal4 39196 4312 39222 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[63].CBOT
flabel metal4 39314 4902 39340 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[63].CTOP
flabel psubdiff 39254 4600 39292 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[63].SUB
flabel psubdiff 14766 3754 14810 3846 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.SUB
flabel metal4 14336 3550 14380 3642 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.CBOT
flabel metal4 14824 3554 14868 3646 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.CTOP
flabel metal4 14702 4074 14746 4166 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.CTOP
flabel metal4 10588 4312 10614 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[0].CBOT
flabel metal4 10706 4902 10732 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[0].CTOP
flabel psubdiff 10646 4600 10684 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[0].SUB
flabel metal4 10710 3456 10736 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[1].CBOT
flabel metal4 10592 2866 10618 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[1].CTOP
flabel psubdiff 10640 3122 10678 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[1].SUB
flabel metal4 11194 4312 11220 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[2].CBOT
flabel metal4 11312 4902 11338 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[2].CTOP
flabel psubdiff 11252 4600 11290 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[2].SUB
flabel metal4 11316 3456 11342 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[3].CBOT
flabel metal4 11198 2866 11224 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[3].CTOP
flabel psubdiff 11246 3122 11284 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[3].SUB
flabel metal4 11800 4312 11826 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[4].CBOT
flabel metal4 11918 4902 11944 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[4].CTOP
flabel psubdiff 11858 4600 11896 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[4].SUB
flabel metal4 11922 3456 11948 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[5].CBOT
flabel metal4 11804 2866 11830 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[5].CTOP
flabel psubdiff 11852 3122 11890 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[5].SUB
flabel metal4 12406 4312 12432 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[6].CBOT
flabel metal4 12524 4902 12550 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[6].CTOP
flabel psubdiff 12464 4600 12502 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[6].SUB
flabel metal4 12528 3456 12554 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[7].CBOT
flabel metal4 12410 2866 12436 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[7].CTOP
flabel psubdiff 12458 3122 12496 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[7].SUB
flabel metal4 13012 4312 13038 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[8].CBOT
flabel metal4 13130 4902 13156 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[8].CTOP
flabel psubdiff 13070 4600 13108 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[8].SUB
flabel metal4 13134 3456 13160 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[9].CBOT
flabel metal4 13016 2866 13042 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[9].CTOP
flabel psubdiff 13064 3122 13102 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[9].SUB
flabel metal4 13618 4312 13644 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[10].CBOT
flabel metal4 13736 4902 13762 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[10].CTOP
flabel psubdiff 13676 4600 13714 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[10].SUB
flabel metal4 13740 3456 13766 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[11].CBOT
flabel metal4 13622 2866 13648 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[11].CTOP
flabel psubdiff 13670 3122 13708 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[11].SUB
flabel metal4 14224 4312 14250 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[12].CBOT
flabel metal4 14342 4902 14368 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[12].CTOP
flabel psubdiff 14282 4600 14320 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[12].SUB
flabel metal4 14346 3456 14372 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[13].CBOT
flabel metal4 14228 2866 14254 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[13].CTOP
flabel psubdiff 14276 3122 14314 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[13].SUB
flabel metal4 14830 4312 14856 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[14].CBOT
flabel metal4 14948 4902 14974 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[14].CTOP
flabel psubdiff 14888 4600 14926 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[14].SUB
flabel metal4 14952 3456 14978 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[15].CBOT
flabel metal4 14834 2866 14860 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[15].CTOP
flabel psubdiff 14882 3122 14920 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[15].SUB
flabel metal4 15436 4312 15462 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[16].CBOT
flabel metal4 15554 4902 15580 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[16].CTOP
flabel psubdiff 15494 4600 15532 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[16].SUB
flabel metal4 15558 3456 15584 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[17].CBOT
flabel metal4 15440 2866 15466 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[17].CTOP
flabel psubdiff 15488 3122 15526 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[17].SUB
flabel metal4 16042 4312 16068 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[18].CBOT
flabel metal4 16160 4902 16186 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[18].CTOP
flabel psubdiff 16100 4600 16138 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[18].SUB
flabel metal4 16164 3456 16190 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[19].CBOT
flabel metal4 16046 2866 16072 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[19].CTOP
flabel psubdiff 16094 3122 16132 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[19].SUB
flabel metal4 16648 4312 16674 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[20].CBOT
flabel metal4 16766 4902 16792 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[20].CTOP
flabel psubdiff 16706 4600 16744 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[20].SUB
flabel metal4 16770 3456 16796 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[21].CBOT
flabel metal4 16652 2866 16678 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[21].CTOP
flabel psubdiff 16700 3122 16738 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[21].SUB
flabel metal4 17254 4312 17280 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[22].CBOT
flabel metal4 17372 4902 17398 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[22].CTOP
flabel psubdiff 17312 4600 17350 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[22].SUB
flabel metal4 17376 3456 17402 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[23].CBOT
flabel metal4 17258 2866 17284 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[23].CTOP
flabel psubdiff 17306 3122 17344 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[23].SUB
flabel metal4 17860 4312 17886 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[24].CBOT
flabel metal4 17978 4902 18004 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[24].CTOP
flabel psubdiff 17918 4600 17956 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[24].SUB
flabel metal4 17982 3456 18008 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[25].CBOT
flabel metal4 17864 2866 17890 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[25].CTOP
flabel psubdiff 17912 3122 17950 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[25].SUB
flabel metal4 18466 4312 18492 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[26].CBOT
flabel metal4 18584 4902 18610 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[26].CTOP
flabel psubdiff 18524 4600 18562 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[26].SUB
flabel metal4 18588 3456 18614 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[27].CBOT
flabel metal4 18470 2866 18496 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[27].CTOP
flabel psubdiff 18518 3122 18556 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[27].SUB
flabel metal4 19072 4312 19098 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[28].CBOT
flabel metal4 19190 4902 19216 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[28].CTOP
flabel psubdiff 19130 4600 19168 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[28].SUB
flabel metal4 19194 3456 19220 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[29].CBOT
flabel metal4 19076 2866 19102 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[29].CTOP
flabel psubdiff 19124 3122 19162 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[29].SUB
flabel metal4 19678 4312 19704 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[30].CBOT
flabel metal4 19796 4902 19822 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[30].CTOP
flabel psubdiff 19736 4600 19774 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[30].SUB
flabel metal4 19800 3456 19826 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[31].CBOT
flabel metal4 19682 2866 19708 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[31].CTOP
flabel psubdiff 19730 3122 19768 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[31].SUB
flabel metal4 8156 3716 8192 3796 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.CBOT
flabel metal4 7432 3686 7468 3766 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.CTOP
flabel metal4 7546 4058 7590 4140 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.CTOP
flabel psubdiff 7850 3958 7894 4040 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.SUB
flabel metal4 5614 4312 5640 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[0].CBOT
flabel metal4 5732 4902 5758 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[0].CTOP
flabel psubdiff 5672 4600 5710 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[0].SUB
flabel metal4 5736 3456 5762 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[1].CBOT
flabel metal4 5618 2866 5644 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[1].CTOP
flabel psubdiff 5666 3122 5704 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[1].SUB
flabel metal4 6220 4312 6246 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[2].CBOT
flabel metal4 6338 4902 6364 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[2].CTOP
flabel psubdiff 6278 4600 6316 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[2].SUB
flabel metal4 6342 3456 6368 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[3].CBOT
flabel metal4 6224 2866 6250 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[3].CTOP
flabel psubdiff 6272 3122 6310 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[3].SUB
flabel metal4 6826 4312 6852 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[4].CBOT
flabel metal4 6944 4902 6970 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[4].CTOP
flabel psubdiff 6884 4600 6922 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[4].SUB
flabel metal4 6948 3456 6974 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[5].CBOT
flabel metal4 6830 2866 6856 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[5].CTOP
flabel psubdiff 6878 3122 6916 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[5].SUB
flabel metal4 7432 4312 7458 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[6].CBOT
flabel metal4 7550 4902 7576 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[6].CTOP
flabel psubdiff 7490 4600 7528 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[6].SUB
flabel metal4 7554 3456 7580 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[7].CBOT
flabel metal4 7436 2866 7462 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[7].CTOP
flabel psubdiff 7484 3122 7522 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[7].SUB
flabel metal4 8038 4312 8064 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[8].CBOT
flabel metal4 8156 4902 8182 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[8].CTOP
flabel psubdiff 8096 4600 8134 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[8].SUB
flabel metal4 8160 3456 8186 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[9].CBOT
flabel metal4 8042 2866 8068 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[9].CTOP
flabel psubdiff 8090 3122 8128 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[9].SUB
flabel metal4 8644 4312 8670 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[10].CBOT
flabel metal4 8762 4902 8788 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[10].CTOP
flabel psubdiff 8702 4600 8740 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[10].SUB
flabel metal4 8766 3456 8792 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[11].CBOT
flabel metal4 8648 2866 8674 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[11].CTOP
flabel psubdiff 8696 3122 8734 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[11].SUB
flabel metal4 9250 4312 9276 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[12].CBOT
flabel metal4 9368 4902 9394 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[12].CTOP
flabel psubdiff 9308 4600 9346 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[12].SUB
flabel metal4 9372 3456 9398 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[13].CBOT
flabel metal4 9254 2866 9280 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[13].CTOP
flabel psubdiff 9302 3122 9340 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[13].SUB
flabel metal4 9856 4312 9882 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[14].CBOT
flabel metal4 9974 4902 10000 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[14].CTOP
flabel psubdiff 9914 4600 9952 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[14].SUB
flabel metal4 9978 3456 10004 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[15].CBOT
flabel metal4 9860 2866 9886 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[15].CTOP
flabel psubdiff 9908 3122 9946 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[15].SUB
flabel psubdiff 4207 3754 4251 3854 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_8_0.SUB
flabel metal4 4387 3586 4433 3678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_8_0.CBOT
flabel metal4 3659 3608 3705 3700 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_8_0.CTOP
flabel metal4 3787 4446 3827 4530 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_8_0.CTOP
flabel metal4 5003 3456 5029 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_8_0.x1[7].CBOT
flabel metal4 4885 2866 4911 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_8_0.x1[7].CTOP
flabel psubdiff 4933 3122 4971 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_8_0.x1[7].SUB
flabel metal4 4881 4312 4907 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_8_0.x1[6].CBOT
flabel metal4 4999 4902 5025 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_8_0.x1[6].CTOP
flabel psubdiff 4939 4600 4977 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_8_0.x1[6].SUB
flabel metal4 4397 3456 4423 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_8_0.x1[5].CBOT
flabel metal4 4279 2866 4305 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_8_0.x1[5].CTOP
flabel psubdiff 4327 3122 4365 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_8_0.x1[5].SUB
flabel metal4 4275 4312 4301 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_8_0.x1[4].CBOT
flabel metal4 4393 4902 4419 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_8_0.x1[4].CTOP
flabel psubdiff 4333 4600 4371 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_8_0.x1[4].SUB
flabel metal4 3791 3456 3817 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_8_0.x1[3].CBOT
flabel metal4 3673 2866 3699 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_8_0.x1[3].CTOP
flabel psubdiff 3721 3122 3759 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_8_0.x1[3].SUB
flabel metal4 3669 4312 3695 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_8_0.x1[2].CBOT
flabel metal4 3787 4902 3813 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_8_0.x1[2].CTOP
flabel psubdiff 3727 4600 3765 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_8_0.x1[2].SUB
flabel metal4 3185 3456 3211 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_8_0.x1[1].CBOT
flabel metal4 3067 2866 3093 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_8_0.x1[1].CTOP
flabel psubdiff 3115 3122 3153 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_8_0.x1[1].SUB
flabel metal4 3063 4312 3089 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_8_0.x1[0].CBOT
flabel metal4 3181 4902 3207 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_8_0.x1[0].CTOP
flabel psubdiff 3121 4600 3159 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_8_0.x1[0].SUB
flabel metal4 2245 3814 2297 3854 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT
flabel metal4 1519 3698 1571 3738 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CTOP
flabel psubdiff 2069 3708 2109 3818 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.SUB
flabel metal4 1643 4036 1681 4118 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CTOP
flabel metal4 2257 3456 2283 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.x1[3].CBOT
flabel metal4 2139 2866 2165 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.x1[3].CTOP
flabel psubdiff 2187 3122 2225 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.x1[3].SUB
flabel metal4 2135 4312 2161 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.x1[2].CBOT
flabel metal4 2253 4902 2279 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.x1[2].CTOP
flabel psubdiff 2193 4600 2231 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.x1[2].SUB
flabel metal4 1651 3456 1677 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.x1[1].CBOT
flabel metal4 1533 2866 1559 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.x1[1].CTOP
flabel psubdiff 1581 3122 1619 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.x1[1].SUB
flabel metal4 1529 4312 1555 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.x1[0].CBOT
flabel metal4 1647 4902 1673 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.x1[0].CTOP
flabel psubdiff 1587 4600 1625 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.x1[0].SUB
flabel psubdiff 669 3615 717 3729 0 FreeSans 160 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_2_0.SUB
flabel metal4 733 3610 769 3700 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_2_0.CBOT
flabel metal4 613 3168 649 3270 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_2_0.CTOP
flabel metal4 731 4752 771 4830 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_2_0.CTOP
flabel metal4 739 3456 765 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_2_0.x2.CBOT
flabel metal4 621 2866 647 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_2_0.x2.CTOP
flabel psubdiff 669 3122 707 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_2_0.x2.SUB
flabel metal4 617 4312 643 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_2_0.x1.CBOT
flabel metal4 735 4902 761 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_2_0.x1.CTOP
flabel psubdiff 675 4600 713 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_2_0.x1.SUB
flabel metal4 -197 3152 -171 3184 0 FreeSans 320 0 0 0 hgu_cdac_unit_1.CBOT
flabel metal4 -79 3742 -53 3774 0 FreeSans 320 0 0 0 hgu_cdac_unit_1.CTOP
flabel psubdiff -139 3440 -101 3518 0 FreeSans 320 0 0 0 hgu_cdac_unit_1.SUB
flabel metal1 7266 5770 7293 5785 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF
flabel metal1 7229 5696 7255 5724 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD
flabel metal1 7227 6274 7251 6304 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VSS
flabel metal1 7531 5770 7558 5785 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VREF
flabel metal1 7569 5696 7595 5724 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VDD
flabel metal1 7573 6274 7597 6304 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VSS
flabel metal1 7010 5770 7037 5785 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VREF
flabel metal1 6973 5696 6999 5724 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VDD
flabel metal1 6971 6274 6995 6304 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VSS
flabel metal1 7275 5770 7302 5785 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VREF
flabel metal1 7313 5696 7339 5724 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VDD
flabel metal1 7317 6274 7341 6304 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VSS
flabel metal1 6754 5770 6781 5785 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VREF
flabel metal1 6717 5696 6743 5724 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VDD
flabel metal1 6715 6274 6739 6304 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VSS
flabel metal1 7019 5770 7046 5785 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VREF
flabel metal1 7057 5696 7083 5724 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VDD
flabel metal1 7061 6274 7085 6304 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VSS
flabel metal1 6498 5770 6525 5785 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VREF
flabel metal1 6461 5696 6487 5724 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VDD
flabel metal1 6459 6274 6483 6304 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VSS
flabel metal1 6763 5770 6790 5785 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VREF
flabel metal1 6801 5696 6827 5724 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VDD
flabel metal1 6805 6274 6829 6304 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VSS
flabel metal1 6242 5770 6269 5785 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VREF
flabel metal1 6205 5696 6231 5724 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VDD
flabel metal1 6203 6274 6227 6304 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VSS
flabel metal1 6507 5770 6534 5785 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VREF
flabel metal1 6545 5696 6571 5724 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VDD
flabel metal1 6549 6274 6573 6304 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VSS
flabel metal1 5986 5770 6013 5785 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VREF
flabel metal1 5949 5696 5975 5724 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VDD
flabel metal1 5947 6274 5971 6304 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VSS
flabel metal1 6251 5770 6278 5785 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VREF
flabel metal1 6289 5696 6315 5724 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VDD
flabel metal1 6293 6274 6317 6304 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VSS
flabel metal1 5730 5770 5757 5785 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VREF
flabel metal1 5693 5696 5719 5724 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VDD
flabel metal1 5691 6274 5715 6304 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VSS
flabel metal1 5995 5770 6022 5785 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VREF
flabel metal1 6033 5696 6059 5724 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VDD
flabel metal1 6037 6274 6061 6304 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VSS
flabel metal1 5474 5770 5501 5785 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VREF
flabel metal1 5437 5696 5463 5724 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VDD
flabel metal1 5435 6274 5459 6304 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VSS
flabel metal1 5739 5770 5766 5785 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VREF
flabel metal1 5777 5696 5803 5724 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VDD
flabel metal1 5781 6274 5805 6304 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VSS
flabel metal1 3749 5770 3776 5785 0 FreeSans 160 0 0 0 inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF
flabel metal1 3712 5696 3738 5724 0 FreeSans 160 0 0 0 inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD
flabel metal1 3710 6274 3734 6304 0 FreeSans 160 0 0 0 inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VSS
flabel metal1 4014 5770 4041 5785 0 FreeSans 160 0 0 0 inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VREF
flabel metal1 4052 5696 4078 5724 0 FreeSans 160 0 0 0 inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VDD
flabel metal1 4056 6274 4080 6304 0 FreeSans 160 0 0 0 inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VSS
flabel metal1 3493 5770 3520 5785 0 FreeSans 160 0 0 0 inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VREF
flabel metal1 3456 5696 3482 5724 0 FreeSans 160 0 0 0 inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VDD
flabel metal1 3454 6274 3478 6304 0 FreeSans 160 0 0 0 inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VSS
flabel metal1 3758 5770 3785 5785 0 FreeSans 160 0 0 0 inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VREF
flabel metal1 3796 5696 3822 5724 0 FreeSans 160 0 0 0 inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VDD
flabel metal1 3800 6274 3824 6304 0 FreeSans 160 0 0 0 inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VSS
flabel metal1 3237 5770 3264 5785 0 FreeSans 160 0 0 0 inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VREF
flabel metal1 3200 5696 3226 5724 0 FreeSans 160 0 0 0 inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VDD
flabel metal1 3198 6274 3222 6304 0 FreeSans 160 0 0 0 inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VSS
flabel metal1 3502 5770 3529 5785 0 FreeSans 160 0 0 0 inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VREF
flabel metal1 3540 5696 3566 5724 0 FreeSans 160 0 0 0 inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VDD
flabel metal1 3544 6274 3568 6304 0 FreeSans 160 0 0 0 inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VSS
flabel metal1 2981 5770 3008 5785 0 FreeSans 160 0 0 0 inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VREF
flabel metal1 2944 5696 2970 5724 0 FreeSans 160 0 0 0 inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VDD
flabel metal1 2942 6274 2966 6304 0 FreeSans 160 0 0 0 inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VSS
flabel metal1 3246 5770 3273 5785 0 FreeSans 160 0 0 0 inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VREF
flabel metal1 3284 5696 3310 5724 0 FreeSans 160 0 0 0 inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VDD
flabel metal1 3288 6274 3312 6304 0 FreeSans 160 0 0 0 inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VSS
flabel metal1 3758 5633 3785 5648 0 FreeSans 160 0 0 0 inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VREF
flabel metal1 3796 5694 3822 5722 0 FreeSans 160 0 0 0 inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VDD
flabel metal1 3800 5114 3824 5144 0 FreeSans 160 0 0 0 inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VSS
flabel metal1 3493 5633 3520 5648 0 FreeSans 160 0 0 0 inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VREF
flabel metal1 3456 5694 3482 5722 0 FreeSans 160 0 0 0 inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VDD
flabel metal1 3454 5114 3478 5144 0 FreeSans 160 0 0 0 inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VSS
flabel metal1 4014 5633 4041 5648 0 FreeSans 160 0 0 0 inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VREF
flabel metal1 4052 5694 4078 5722 0 FreeSans 160 0 0 0 inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VDD
flabel metal1 4056 5114 4080 5144 0 FreeSans 160 0 0 0 inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VSS
flabel metal1 3749 5633 3776 5648 0 FreeSans 160 0 0 0 inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VREF
flabel metal1 3712 5694 3738 5722 0 FreeSans 160 0 0 0 inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VDD
flabel metal1 3710 5114 3734 5144 0 FreeSans 160 0 0 0 inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VSS
flabel metal1 4270 5633 4297 5648 0 FreeSans 160 0 0 0 inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VREF
flabel metal1 4308 5694 4334 5722 0 FreeSans 160 0 0 0 inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VDD
flabel metal1 4312 5114 4336 5144 0 FreeSans 160 0 0 0 inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VSS
flabel metal1 4005 5633 4032 5648 0 FreeSans 160 0 0 0 inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VREF
flabel metal1 3968 5694 3994 5722 0 FreeSans 160 0 0 0 inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VDD
flabel metal1 3966 5114 3990 5144 0 FreeSans 160 0 0 0 inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VSS
flabel metal1 4526 5633 4553 5648 0 FreeSans 160 0 0 0 inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VREF
flabel metal1 4564 5694 4590 5722 0 FreeSans 160 0 0 0 inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VDD
flabel metal1 4568 5114 4592 5144 0 FreeSans 160 0 0 0 inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VSS
flabel metal1 4261 5633 4288 5648 0 FreeSans 160 0 0 0 inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VREF
flabel metal1 4224 5694 4250 5722 0 FreeSans 160 0 0 0 inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VDD
flabel metal1 4222 5114 4246 5144 0 FreeSans 160 0 0 0 inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VSS
flabel metal1 1618 5770 1645 5785 0 FreeSans 160 0 0 0 inv_4_test_2/inv_2_test_1/x2.VREF
flabel metal1 1581 5696 1607 5724 0 FreeSans 160 0 0 0 inv_4_test_2/inv_2_test_1/x2.VDD
flabel metal1 1579 6274 1603 6304 0 FreeSans 160 0 0 0 inv_4_test_2/inv_2_test_1/x2.VSS
flabel metal1 1883 5770 1910 5785 0 FreeSans 160 0 0 0 inv_4_test_2/inv_2_test_1/x1.VREF
flabel metal1 1921 5696 1947 5724 0 FreeSans 160 0 0 0 inv_4_test_2/inv_2_test_1/x1.VDD
flabel metal1 1925 6274 1949 6304 0 FreeSans 160 0 0 0 inv_4_test_2/inv_2_test_1/x1.VSS
flabel metal1 1362 5770 1389 5785 0 FreeSans 160 0 0 0 inv_4_test_2/inv_2_test_0/x2.VREF
flabel metal1 1325 5696 1351 5724 0 FreeSans 160 0 0 0 inv_4_test_2/inv_2_test_0/x2.VDD
flabel metal1 1323 6274 1347 6304 0 FreeSans 160 0 0 0 inv_4_test_2/inv_2_test_0/x2.VSS
flabel metal1 1627 5770 1654 5785 0 FreeSans 160 0 0 0 inv_4_test_2/inv_2_test_0/x1.VREF
flabel metal1 1665 5696 1691 5724 0 FreeSans 160 0 0 0 inv_4_test_2/inv_2_test_0/x1.VDD
flabel metal1 1669 6274 1693 6304 0 FreeSans 160 0 0 0 inv_4_test_2/inv_2_test_0/x1.VSS
flabel metal1 2139 5633 2166 5648 0 FreeSans 160 0 0 0 inv_4_test_1/inv_2_test_1/x2.VREF
flabel metal1 2177 5694 2203 5722 0 FreeSans 160 0 0 0 inv_4_test_1/inv_2_test_1/x2.VDD
flabel metal1 2181 5114 2205 5144 0 FreeSans 160 0 0 0 inv_4_test_1/inv_2_test_1/x2.VSS
flabel metal1 1874 5633 1901 5648 0 FreeSans 160 0 0 0 inv_4_test_1/inv_2_test_1/x1.VREF
flabel metal1 1837 5694 1863 5722 0 FreeSans 160 0 0 0 inv_4_test_1/inv_2_test_1/x1.VDD
flabel metal1 1835 5114 1859 5144 0 FreeSans 160 0 0 0 inv_4_test_1/inv_2_test_1/x1.VSS
flabel metal1 2395 5633 2422 5648 0 FreeSans 160 0 0 0 inv_4_test_1/inv_2_test_0/x2.VREF
flabel metal1 2433 5694 2459 5722 0 FreeSans 160 0 0 0 inv_4_test_1/inv_2_test_0/x2.VDD
flabel metal1 2437 5114 2461 5144 0 FreeSans 160 0 0 0 inv_4_test_1/inv_2_test_0/x2.VSS
flabel metal1 2130 5633 2157 5648 0 FreeSans 160 0 0 0 inv_4_test_1/inv_2_test_0/x1.VREF
flabel metal1 2093 5694 2119 5722 0 FreeSans 160 0 0 0 inv_4_test_1/inv_2_test_0/x1.VDD
flabel metal1 2091 5114 2115 5144 0 FreeSans 160 0 0 0 inv_4_test_1/inv_2_test_0/x1.VSS
flabel metal1 482 5770 509 5785 0 FreeSans 160 0 0 0 inv_2_test_1/x2.VREF
flabel metal1 445 5696 471 5724 0 FreeSans 160 0 0 0 inv_2_test_1/x2.VDD
flabel metal1 443 6274 467 6304 0 FreeSans 160 0 0 0 inv_2_test_1/x2.VSS
flabel metal1 747 5770 774 5785 0 FreeSans 160 0 0 0 inv_2_test_1/x1.VREF
flabel metal1 785 5696 811 5724 0 FreeSans 160 0 0 0 inv_2_test_1/x1.VDD
flabel metal1 789 6274 813 6304 0 FreeSans 160 0 0 0 inv_2_test_1/x1.VSS
flabel metal1 875 5633 902 5648 0 FreeSans 160 0 0 0 inv_2_test_0/x2.VREF
flabel metal1 913 5694 939 5722 0 FreeSans 160 0 0 0 inv_2_test_0/x2.VDD
flabel metal1 917 5114 941 5144 0 FreeSans 160 0 0 0 inv_2_test_0/x2.VSS
flabel metal1 610 5633 637 5648 0 FreeSans 160 0 0 0 inv_2_test_0/x1.VREF
flabel metal1 573 5694 599 5722 0 FreeSans 160 0 0 0 inv_2_test_0/x1.VDD
flabel metal1 571 5114 595 5144 0 FreeSans 160 0 0 0 inv_2_test_0/x1.VSS
flabel metal1 -318 5770 -291 5785 0 FreeSans 160 0 0 0 hgu_inverter_1.VREF
flabel metal1 -355 5696 -329 5724 0 FreeSans 160 0 0 0 hgu_inverter_1.VDD
flabel metal1 -357 6274 -333 6304 0 FreeSans 160 0 0 0 hgu_inverter_1.VSS
flabel metal1 -318 5633 -291 5648 0 FreeSans 160 0 0 0 hgu_inverter_0.VREF
flabel metal1 -355 5694 -329 5722 0 FreeSans 160 0 0 0 hgu_inverter_0.VDD
flabel metal1 -357 5114 -333 5144 0 FreeSans 160 0 0 0 hgu_inverter_0.VSS
flabel metal1 16087 5633 16114 5648 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF
flabel metal1 16125 5694 16151 5722 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD
flabel metal1 16129 5114 16153 5144 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VSS
flabel metal1 15822 5633 15849 5648 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VREF
flabel metal1 15785 5694 15811 5722 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VDD
flabel metal1 15783 5114 15807 5144 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VSS
flabel metal1 16343 5633 16370 5648 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VREF
flabel metal1 16381 5694 16407 5722 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VDD
flabel metal1 16385 5114 16409 5144 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VSS
flabel metal1 16078 5633 16105 5648 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VREF
flabel metal1 16041 5694 16067 5722 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VDD
flabel metal1 16039 5114 16063 5144 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VSS
flabel metal1 16599 5633 16626 5648 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VREF
flabel metal1 16637 5694 16663 5722 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VDD
flabel metal1 16641 5114 16665 5144 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VSS
flabel metal1 16334 5633 16361 5648 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VREF
flabel metal1 16297 5694 16323 5722 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VDD
flabel metal1 16295 5114 16319 5144 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VSS
flabel metal1 16855 5633 16882 5648 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VREF
flabel metal1 16893 5694 16919 5722 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VDD
flabel metal1 16897 5114 16921 5144 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VSS
flabel metal1 16590 5633 16617 5648 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VREF
flabel metal1 16553 5694 16579 5722 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VDD
flabel metal1 16551 5114 16575 5144 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VSS
flabel metal1 17111 5633 17138 5648 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VREF
flabel metal1 17149 5694 17175 5722 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VDD
flabel metal1 17153 5114 17177 5144 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VSS
flabel metal1 16846 5633 16873 5648 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VREF
flabel metal1 16809 5694 16835 5722 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VDD
flabel metal1 16807 5114 16831 5144 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VSS
flabel metal1 17367 5633 17394 5648 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VREF
flabel metal1 17405 5694 17431 5722 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VDD
flabel metal1 17409 5114 17433 5144 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VSS
flabel metal1 17102 5633 17129 5648 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VREF
flabel metal1 17065 5694 17091 5722 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VDD
flabel metal1 17063 5114 17087 5144 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VSS
flabel metal1 17623 5633 17650 5648 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VREF
flabel metal1 17661 5694 17687 5722 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VDD
flabel metal1 17665 5114 17689 5144 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VSS
flabel metal1 17358 5633 17385 5648 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VREF
flabel metal1 17321 5694 17347 5722 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VDD
flabel metal1 17319 5114 17343 5144 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VSS
flabel metal1 17879 5633 17906 5648 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VREF
flabel metal1 17917 5694 17943 5722 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VDD
flabel metal1 17921 5114 17945 5144 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VSS
flabel metal1 17614 5633 17641 5648 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VREF
flabel metal1 17577 5694 17603 5722 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VDD
flabel metal1 17575 5114 17599 5144 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VSS
flabel metal1 18135 5633 18162 5648 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF
flabel metal1 18173 5694 18199 5722 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD
flabel metal1 18177 5114 18201 5144 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VSS
flabel metal1 17870 5633 17897 5648 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VREF
flabel metal1 17833 5694 17859 5722 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VDD
flabel metal1 17831 5114 17855 5144 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VSS
flabel metal1 18391 5633 18418 5648 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VREF
flabel metal1 18429 5694 18455 5722 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VDD
flabel metal1 18433 5114 18457 5144 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VSS
flabel metal1 18126 5633 18153 5648 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VREF
flabel metal1 18089 5694 18115 5722 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VDD
flabel metal1 18087 5114 18111 5144 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VSS
flabel metal1 18647 5633 18674 5648 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VREF
flabel metal1 18685 5694 18711 5722 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VDD
flabel metal1 18689 5114 18713 5144 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VSS
flabel metal1 18382 5633 18409 5648 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VREF
flabel metal1 18345 5694 18371 5722 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VDD
flabel metal1 18343 5114 18367 5144 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VSS
flabel metal1 18903 5633 18930 5648 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VREF
flabel metal1 18941 5694 18967 5722 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VDD
flabel metal1 18945 5114 18969 5144 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VSS
flabel metal1 18638 5633 18665 5648 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VREF
flabel metal1 18601 5694 18627 5722 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VDD
flabel metal1 18599 5114 18623 5144 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VSS
flabel metal1 19159 5633 19186 5648 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VREF
flabel metal1 19197 5694 19223 5722 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VDD
flabel metal1 19201 5114 19225 5144 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VSS
flabel metal1 18894 5633 18921 5648 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VREF
flabel metal1 18857 5694 18883 5722 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VDD
flabel metal1 18855 5114 18879 5144 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VSS
flabel metal1 19415 5633 19442 5648 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VREF
flabel metal1 19453 5694 19479 5722 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VDD
flabel metal1 19457 5114 19481 5144 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VSS
flabel metal1 19150 5633 19177 5648 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VREF
flabel metal1 19113 5694 19139 5722 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VDD
flabel metal1 19111 5114 19135 5144 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VSS
flabel metal1 19671 5633 19698 5648 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VREF
flabel metal1 19709 5694 19735 5722 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VDD
flabel metal1 19713 5114 19737 5144 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VSS
flabel metal1 19406 5633 19433 5648 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VREF
flabel metal1 19369 5694 19395 5722 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VDD
flabel metal1 19367 5114 19391 5144 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VSS
flabel metal1 19927 5633 19954 5648 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VREF
flabel metal1 19965 5694 19991 5722 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VDD
flabel metal1 19969 5114 19993 5144 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VSS
flabel metal1 19662 5633 19689 5648 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VREF
flabel metal1 19625 5694 19651 5722 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VDD
flabel metal1 19623 5114 19647 5144 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VSS
flabel metal1 14401 5770 14428 5785 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF
flabel metal1 14364 5696 14390 5724 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD
flabel metal1 14362 6274 14386 6304 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VSS
flabel metal1 14666 5770 14693 5785 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VREF
flabel metal1 14704 5696 14730 5724 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VDD
flabel metal1 14708 6274 14732 6304 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VSS
flabel metal1 14145 5770 14172 5785 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VREF
flabel metal1 14108 5696 14134 5724 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VDD
flabel metal1 14106 6274 14130 6304 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VSS
flabel metal1 14410 5770 14437 5785 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VREF
flabel metal1 14448 5696 14474 5724 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VDD
flabel metal1 14452 6274 14476 6304 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VSS
flabel metal1 13889 5770 13916 5785 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VREF
flabel metal1 13852 5696 13878 5724 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VDD
flabel metal1 13850 6274 13874 6304 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VSS
flabel metal1 14154 5770 14181 5785 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VREF
flabel metal1 14192 5696 14218 5724 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VDD
flabel metal1 14196 6274 14220 6304 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VSS
flabel metal1 13633 5770 13660 5785 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VREF
flabel metal1 13596 5696 13622 5724 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VDD
flabel metal1 13594 6274 13618 6304 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VSS
flabel metal1 13898 5770 13925 5785 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VREF
flabel metal1 13936 5696 13962 5724 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VDD
flabel metal1 13940 6274 13964 6304 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VSS
flabel metal1 13377 5770 13404 5785 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VREF
flabel metal1 13340 5696 13366 5724 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VDD
flabel metal1 13338 6274 13362 6304 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VSS
flabel metal1 13642 5770 13669 5785 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VREF
flabel metal1 13680 5696 13706 5724 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VDD
flabel metal1 13684 6274 13708 6304 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VSS
flabel metal1 13121 5770 13148 5785 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VREF
flabel metal1 13084 5696 13110 5724 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VDD
flabel metal1 13082 6274 13106 6304 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VSS
flabel metal1 13386 5770 13413 5785 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VREF
flabel metal1 13424 5696 13450 5724 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VDD
flabel metal1 13428 6274 13452 6304 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VSS
flabel metal1 12865 5770 12892 5785 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VREF
flabel metal1 12828 5696 12854 5724 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VDD
flabel metal1 12826 6274 12850 6304 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VSS
flabel metal1 13130 5770 13157 5785 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VREF
flabel metal1 13168 5696 13194 5724 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VDD
flabel metal1 13172 6274 13196 6304 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VSS
flabel metal1 12609 5770 12636 5785 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VREF
flabel metal1 12572 5696 12598 5724 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VDD
flabel metal1 12570 6274 12594 6304 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VSS
flabel metal1 12874 5770 12901 5785 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VREF
flabel metal1 12912 5696 12938 5724 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VDD
flabel metal1 12916 6274 12940 6304 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VSS
flabel metal1 12353 5770 12380 5785 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF
flabel metal1 12316 5696 12342 5724 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD
flabel metal1 12314 6274 12338 6304 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VSS
flabel metal1 12618 5770 12645 5785 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VREF
flabel metal1 12656 5696 12682 5724 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VDD
flabel metal1 12660 6274 12684 6304 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VSS
flabel metal1 12097 5770 12124 5785 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VREF
flabel metal1 12060 5696 12086 5724 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VDD
flabel metal1 12058 6274 12082 6304 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VSS
flabel metal1 12362 5770 12389 5785 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VREF
flabel metal1 12400 5696 12426 5724 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VDD
flabel metal1 12404 6274 12428 6304 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VSS
flabel metal1 11841 5770 11868 5785 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VREF
flabel metal1 11804 5696 11830 5724 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VDD
flabel metal1 11802 6274 11826 6304 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VSS
flabel metal1 12106 5770 12133 5785 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VREF
flabel metal1 12144 5696 12170 5724 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VDD
flabel metal1 12148 6274 12172 6304 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VSS
flabel metal1 11585 5770 11612 5785 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VREF
flabel metal1 11548 5696 11574 5724 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VDD
flabel metal1 11546 6274 11570 6304 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VSS
flabel metal1 11850 5770 11877 5785 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VREF
flabel metal1 11888 5696 11914 5724 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VDD
flabel metal1 11892 6274 11916 6304 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VSS
flabel metal1 11329 5770 11356 5785 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VREF
flabel metal1 11292 5696 11318 5724 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VDD
flabel metal1 11290 6274 11314 6304 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VSS
flabel metal1 11594 5770 11621 5785 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VREF
flabel metal1 11632 5696 11658 5724 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VDD
flabel metal1 11636 6274 11660 6304 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VSS
flabel metal1 11073 5770 11100 5785 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VREF
flabel metal1 11036 5696 11062 5724 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VDD
flabel metal1 11034 6274 11058 6304 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VSS
flabel metal1 11338 5770 11365 5785 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VREF
flabel metal1 11376 5696 11402 5724 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VDD
flabel metal1 11380 6274 11404 6304 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VSS
flabel metal1 10817 5770 10844 5785 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VREF
flabel metal1 10780 5696 10806 5724 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VDD
flabel metal1 10778 6274 10802 6304 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VSS
flabel metal1 11082 5770 11109 5785 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VREF
flabel metal1 11120 5696 11146 5724 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VDD
flabel metal1 11124 6274 11148 6304 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VSS
flabel metal1 10561 5770 10588 5785 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VREF
flabel metal1 10524 5696 10550 5724 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VDD
flabel metal1 10522 6274 10546 6304 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VSS
flabel metal1 10826 5770 10853 5785 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VREF
flabel metal1 10864 5696 10890 5724 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VDD
flabel metal1 10868 6274 10892 6304 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VSS
flabel metal1 8323 5633 8350 5648 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF
flabel metal1 8361 5694 8387 5722 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD
flabel metal1 8365 5114 8389 5144 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VSS
flabel metal1 8058 5633 8085 5648 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VREF
flabel metal1 8021 5694 8047 5722 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VDD
flabel metal1 8019 5114 8043 5144 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VSS
flabel metal1 8579 5633 8606 5648 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VREF
flabel metal1 8617 5694 8643 5722 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VDD
flabel metal1 8621 5114 8645 5144 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VSS
flabel metal1 8314 5633 8341 5648 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VREF
flabel metal1 8277 5694 8303 5722 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VDD
flabel metal1 8275 5114 8299 5144 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VSS
flabel metal1 8835 5633 8862 5648 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VREF
flabel metal1 8873 5694 8899 5722 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VDD
flabel metal1 8877 5114 8901 5144 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VSS
flabel metal1 8570 5633 8597 5648 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VREF
flabel metal1 8533 5694 8559 5722 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VDD
flabel metal1 8531 5114 8555 5144 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VSS
flabel metal1 9091 5633 9118 5648 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VREF
flabel metal1 9129 5694 9155 5722 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VDD
flabel metal1 9133 5114 9157 5144 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VSS
flabel metal1 8826 5633 8853 5648 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VREF
flabel metal1 8789 5694 8815 5722 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VDD
flabel metal1 8787 5114 8811 5144 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VSS
flabel metal1 9347 5633 9374 5648 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VREF
flabel metal1 9385 5694 9411 5722 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VDD
flabel metal1 9389 5114 9413 5144 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VSS
flabel metal1 9082 5633 9109 5648 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VREF
flabel metal1 9045 5694 9071 5722 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VDD
flabel metal1 9043 5114 9067 5144 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VSS
flabel metal1 9603 5633 9630 5648 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VREF
flabel metal1 9641 5694 9667 5722 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VDD
flabel metal1 9645 5114 9669 5144 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VSS
flabel metal1 9338 5633 9365 5648 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VREF
flabel metal1 9301 5694 9327 5722 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VDD
flabel metal1 9299 5114 9323 5144 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VSS
flabel metal1 9859 5633 9886 5648 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VREF
flabel metal1 9897 5694 9923 5722 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VDD
flabel metal1 9901 5114 9925 5144 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VSS
flabel metal1 9594 5633 9621 5648 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VREF
flabel metal1 9557 5694 9583 5722 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VDD
flabel metal1 9555 5114 9579 5144 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VSS
flabel metal1 10115 5633 10142 5648 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VREF
flabel metal1 10153 5694 10179 5722 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VDD
flabel metal1 10157 5114 10181 5144 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VSS
flabel metal1 9850 5633 9877 5648 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VREF
flabel metal1 9813 5694 9839 5722 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VDD
flabel metal1 9811 5114 9835 5144 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VSS
flabel metal1 24238 5770 24265 5785 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF
flabel metal1 24201 5696 24227 5724 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD
flabel metal1 24199 6274 24223 6304 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VSS
flabel metal1 24503 5770 24530 5785 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VREF
flabel metal1 24541 5696 24567 5724 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VDD
flabel metal1 24545 6274 24569 6304 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VSS
flabel metal1 23982 5770 24009 5785 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VREF
flabel metal1 23945 5696 23971 5724 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VDD
flabel metal1 23943 6274 23967 6304 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VSS
flabel metal1 24247 5770 24274 5785 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VREF
flabel metal1 24285 5696 24311 5724 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VDD
flabel metal1 24289 6274 24313 6304 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VSS
flabel metal1 23726 5770 23753 5785 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VREF
flabel metal1 23689 5696 23715 5724 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VDD
flabel metal1 23687 6274 23711 6304 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VSS
flabel metal1 23991 5770 24018 5785 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VREF
flabel metal1 24029 5696 24055 5724 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VDD
flabel metal1 24033 6274 24057 6304 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VSS
flabel metal1 23470 5770 23497 5785 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VREF
flabel metal1 23433 5696 23459 5724 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VDD
flabel metal1 23431 6274 23455 6304 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VSS
flabel metal1 23735 5770 23762 5785 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VREF
flabel metal1 23773 5696 23799 5724 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VDD
flabel metal1 23777 6274 23801 6304 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VSS
flabel metal1 23214 5770 23241 5785 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VREF
flabel metal1 23177 5696 23203 5724 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VDD
flabel metal1 23175 6274 23199 6304 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VSS
flabel metal1 23479 5770 23506 5785 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VREF
flabel metal1 23517 5696 23543 5724 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VDD
flabel metal1 23521 6274 23545 6304 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VSS
flabel metal1 22958 5770 22985 5785 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VREF
flabel metal1 22921 5696 22947 5724 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VDD
flabel metal1 22919 6274 22943 6304 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VSS
flabel metal1 23223 5770 23250 5785 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VREF
flabel metal1 23261 5696 23287 5724 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VDD
flabel metal1 23265 6274 23289 6304 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VSS
flabel metal1 22702 5770 22729 5785 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VREF
flabel metal1 22665 5696 22691 5724 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VDD
flabel metal1 22663 6274 22687 6304 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VSS
flabel metal1 22967 5770 22994 5785 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VREF
flabel metal1 23005 5696 23031 5724 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VDD
flabel metal1 23009 6274 23033 6304 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VSS
flabel metal1 22446 5770 22473 5785 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VREF
flabel metal1 22409 5696 22435 5724 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VDD
flabel metal1 22407 6274 22431 6304 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VSS
flabel metal1 22711 5770 22738 5785 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VREF
flabel metal1 22749 5696 22775 5724 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VDD
flabel metal1 22753 6274 22777 6304 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VSS
flabel metal1 22190 5770 22217 5785 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF
flabel metal1 22153 5696 22179 5724 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD
flabel metal1 22151 6274 22175 6304 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VSS
flabel metal1 22455 5770 22482 5785 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VREF
flabel metal1 22493 5696 22519 5724 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VDD
flabel metal1 22497 6274 22521 6304 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VSS
flabel metal1 21934 5770 21961 5785 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VREF
flabel metal1 21897 5696 21923 5724 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VDD
flabel metal1 21895 6274 21919 6304 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VSS
flabel metal1 22199 5770 22226 5785 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VREF
flabel metal1 22237 5696 22263 5724 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VDD
flabel metal1 22241 6274 22265 6304 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VSS
flabel metal1 21678 5770 21705 5785 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VREF
flabel metal1 21641 5696 21667 5724 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VDD
flabel metal1 21639 6274 21663 6304 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VSS
flabel metal1 21943 5770 21970 5785 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VREF
flabel metal1 21981 5696 22007 5724 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VDD
flabel metal1 21985 6274 22009 6304 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VSS
flabel metal1 21422 5770 21449 5785 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VREF
flabel metal1 21385 5696 21411 5724 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VDD
flabel metal1 21383 6274 21407 6304 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VSS
flabel metal1 21687 5770 21714 5785 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VREF
flabel metal1 21725 5696 21751 5724 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VDD
flabel metal1 21729 6274 21753 6304 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VSS
flabel metal1 21166 5770 21193 5785 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VREF
flabel metal1 21129 5696 21155 5724 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VDD
flabel metal1 21127 6274 21151 6304 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VSS
flabel metal1 21431 5770 21458 5785 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VREF
flabel metal1 21469 5696 21495 5724 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VDD
flabel metal1 21473 6274 21497 6304 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VSS
flabel metal1 20910 5770 20937 5785 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VREF
flabel metal1 20873 5696 20899 5724 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VDD
flabel metal1 20871 6274 20895 6304 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VSS
flabel metal1 21175 5770 21202 5785 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VREF
flabel metal1 21213 5696 21239 5724 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VDD
flabel metal1 21217 6274 21241 6304 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VSS
flabel metal1 20654 5770 20681 5785 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VREF
flabel metal1 20617 5696 20643 5724 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VDD
flabel metal1 20615 6274 20639 6304 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VSS
flabel metal1 20919 5770 20946 5785 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VREF
flabel metal1 20957 5696 20983 5724 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VDD
flabel metal1 20961 6274 20985 6304 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VSS
flabel metal1 20398 5770 20425 5785 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VREF
flabel metal1 20361 5696 20387 5724 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VDD
flabel metal1 20359 6274 20383 6304 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VSS
flabel metal1 20663 5770 20690 5785 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VREF
flabel metal1 20701 5696 20727 5724 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VDD
flabel metal1 20705 6274 20729 6304 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VSS
flabel metal1 28334 5770 28361 5785 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF
flabel metal1 28297 5696 28323 5724 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD
flabel metal1 28295 6274 28319 6304 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VSS
flabel metal1 28599 5770 28626 5785 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VREF
flabel metal1 28637 5696 28663 5724 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VDD
flabel metal1 28641 6274 28665 6304 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VSS
flabel metal1 28078 5770 28105 5785 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VREF
flabel metal1 28041 5696 28067 5724 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VDD
flabel metal1 28039 6274 28063 6304 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VSS
flabel metal1 28343 5770 28370 5785 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VREF
flabel metal1 28381 5696 28407 5724 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VDD
flabel metal1 28385 6274 28409 6304 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VSS
flabel metal1 27822 5770 27849 5785 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VREF
flabel metal1 27785 5696 27811 5724 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VDD
flabel metal1 27783 6274 27807 6304 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VSS
flabel metal1 28087 5770 28114 5785 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VREF
flabel metal1 28125 5696 28151 5724 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VDD
flabel metal1 28129 6274 28153 6304 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VSS
flabel metal1 27566 5770 27593 5785 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VREF
flabel metal1 27529 5696 27555 5724 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VDD
flabel metal1 27527 6274 27551 6304 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VSS
flabel metal1 27831 5770 27858 5785 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VREF
flabel metal1 27869 5696 27895 5724 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VDD
flabel metal1 27873 6274 27897 6304 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VSS
flabel metal1 27310 5770 27337 5785 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VREF
flabel metal1 27273 5696 27299 5724 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VDD
flabel metal1 27271 6274 27295 6304 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VSS
flabel metal1 27575 5770 27602 5785 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VREF
flabel metal1 27613 5696 27639 5724 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VDD
flabel metal1 27617 6274 27641 6304 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VSS
flabel metal1 27054 5770 27081 5785 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VREF
flabel metal1 27017 5696 27043 5724 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VDD
flabel metal1 27015 6274 27039 6304 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VSS
flabel metal1 27319 5770 27346 5785 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VREF
flabel metal1 27357 5696 27383 5724 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VDD
flabel metal1 27361 6274 27385 6304 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VSS
flabel metal1 26798 5770 26825 5785 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VREF
flabel metal1 26761 5696 26787 5724 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VDD
flabel metal1 26759 6274 26783 6304 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VSS
flabel metal1 27063 5770 27090 5785 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VREF
flabel metal1 27101 5696 27127 5724 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VDD
flabel metal1 27105 6274 27129 6304 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VSS
flabel metal1 26542 5770 26569 5785 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VREF
flabel metal1 26505 5696 26531 5724 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VDD
flabel metal1 26503 6274 26527 6304 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VSS
flabel metal1 26807 5770 26834 5785 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VREF
flabel metal1 26845 5696 26871 5724 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VDD
flabel metal1 26849 6274 26873 6304 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VSS
flabel metal1 26286 5770 26313 5785 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF
flabel metal1 26249 5696 26275 5724 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD
flabel metal1 26247 6274 26271 6304 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VSS
flabel metal1 26551 5770 26578 5785 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VREF
flabel metal1 26589 5696 26615 5724 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VDD
flabel metal1 26593 6274 26617 6304 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VSS
flabel metal1 26030 5770 26057 5785 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VREF
flabel metal1 25993 5696 26019 5724 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VDD
flabel metal1 25991 6274 26015 6304 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VSS
flabel metal1 26295 5770 26322 5785 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VREF
flabel metal1 26333 5696 26359 5724 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VDD
flabel metal1 26337 6274 26361 6304 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VSS
flabel metal1 25774 5770 25801 5785 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VREF
flabel metal1 25737 5696 25763 5724 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VDD
flabel metal1 25735 6274 25759 6304 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VSS
flabel metal1 26039 5770 26066 5785 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VREF
flabel metal1 26077 5696 26103 5724 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VDD
flabel metal1 26081 6274 26105 6304 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VSS
flabel metal1 25518 5770 25545 5785 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VREF
flabel metal1 25481 5696 25507 5724 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VDD
flabel metal1 25479 6274 25503 6304 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VSS
flabel metal1 25783 5770 25810 5785 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VREF
flabel metal1 25821 5696 25847 5724 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VDD
flabel metal1 25825 6274 25849 6304 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VSS
flabel metal1 25262 5770 25289 5785 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VREF
flabel metal1 25225 5696 25251 5724 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VDD
flabel metal1 25223 6274 25247 6304 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VSS
flabel metal1 25527 5770 25554 5785 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VREF
flabel metal1 25565 5696 25591 5724 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VDD
flabel metal1 25569 6274 25593 6304 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VSS
flabel metal1 25006 5770 25033 5785 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VREF
flabel metal1 24969 5696 24995 5724 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VDD
flabel metal1 24967 6274 24991 6304 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VSS
flabel metal1 25271 5770 25298 5785 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VREF
flabel metal1 25309 5696 25335 5724 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VDD
flabel metal1 25313 6274 25337 6304 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VSS
flabel metal1 24750 5770 24777 5785 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VREF
flabel metal1 24713 5696 24739 5724 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VDD
flabel metal1 24711 6274 24735 6304 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VSS
flabel metal1 25015 5770 25042 5785 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VREF
flabel metal1 25053 5696 25079 5724 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VDD
flabel metal1 25057 6274 25081 6304 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VSS
flabel metal1 24494 5770 24521 5785 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VREF
flabel metal1 24457 5696 24483 5724 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VDD
flabel metal1 24455 6274 24479 6304 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VSS
flabel metal1 24759 5770 24786 5785 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VREF
flabel metal1 24797 5696 24823 5724 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VDD
flabel metal1 24801 6274 24825 6304 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VSS
flabel metal1 33727 5633 33754 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF
flabel metal1 33765 5694 33791 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD
flabel metal1 33769 5114 33793 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VSS
flabel metal1 33462 5633 33489 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VREF
flabel metal1 33425 5694 33451 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VDD
flabel metal1 33423 5114 33447 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VSS
flabel metal1 33983 5633 34010 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VREF
flabel metal1 34021 5694 34047 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VDD
flabel metal1 34025 5114 34049 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VSS
flabel metal1 33718 5633 33745 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VREF
flabel metal1 33681 5694 33707 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VDD
flabel metal1 33679 5114 33703 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VSS
flabel metal1 34239 5633 34266 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VREF
flabel metal1 34277 5694 34303 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VDD
flabel metal1 34281 5114 34305 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VSS
flabel metal1 33974 5633 34001 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VREF
flabel metal1 33937 5694 33963 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VDD
flabel metal1 33935 5114 33959 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VSS
flabel metal1 34495 5633 34522 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VREF
flabel metal1 34533 5694 34559 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VDD
flabel metal1 34537 5114 34561 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VSS
flabel metal1 34230 5633 34257 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VREF
flabel metal1 34193 5694 34219 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VDD
flabel metal1 34191 5114 34215 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VSS
flabel metal1 34751 5633 34778 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VREF
flabel metal1 34789 5694 34815 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VDD
flabel metal1 34793 5114 34817 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VSS
flabel metal1 34486 5633 34513 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VREF
flabel metal1 34449 5694 34475 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VDD
flabel metal1 34447 5114 34471 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VSS
flabel metal1 35007 5633 35034 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VREF
flabel metal1 35045 5694 35071 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VDD
flabel metal1 35049 5114 35073 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VSS
flabel metal1 34742 5633 34769 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VREF
flabel metal1 34705 5694 34731 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VDD
flabel metal1 34703 5114 34727 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VSS
flabel metal1 35263 5633 35290 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VREF
flabel metal1 35301 5694 35327 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VDD
flabel metal1 35305 5114 35329 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VSS
flabel metal1 34998 5633 35025 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VREF
flabel metal1 34961 5694 34987 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VDD
flabel metal1 34959 5114 34983 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VSS
flabel metal1 35519 5633 35546 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VREF
flabel metal1 35557 5694 35583 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VDD
flabel metal1 35561 5114 35585 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VSS
flabel metal1 35254 5633 35281 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VREF
flabel metal1 35217 5694 35243 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VDD
flabel metal1 35215 5114 35239 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VSS
flabel metal1 35775 5633 35802 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF
flabel metal1 35813 5694 35839 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD
flabel metal1 35817 5114 35841 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VSS
flabel metal1 35510 5633 35537 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VREF
flabel metal1 35473 5694 35499 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VDD
flabel metal1 35471 5114 35495 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VSS
flabel metal1 36031 5633 36058 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VREF
flabel metal1 36069 5694 36095 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VDD
flabel metal1 36073 5114 36097 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VSS
flabel metal1 35766 5633 35793 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VREF
flabel metal1 35729 5694 35755 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VDD
flabel metal1 35727 5114 35751 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VSS
flabel metal1 36287 5633 36314 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VREF
flabel metal1 36325 5694 36351 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VDD
flabel metal1 36329 5114 36353 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VSS
flabel metal1 36022 5633 36049 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VREF
flabel metal1 35985 5694 36011 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VDD
flabel metal1 35983 5114 36007 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VSS
flabel metal1 36543 5633 36570 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VREF
flabel metal1 36581 5694 36607 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VDD
flabel metal1 36585 5114 36609 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VSS
flabel metal1 36278 5633 36305 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VREF
flabel metal1 36241 5694 36267 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VDD
flabel metal1 36239 5114 36263 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VSS
flabel metal1 36799 5633 36826 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VREF
flabel metal1 36837 5694 36863 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VDD
flabel metal1 36841 5114 36865 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VSS
flabel metal1 36534 5633 36561 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VREF
flabel metal1 36497 5694 36523 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VDD
flabel metal1 36495 5114 36519 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VSS
flabel metal1 37055 5633 37082 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VREF
flabel metal1 37093 5694 37119 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VDD
flabel metal1 37097 5114 37121 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VSS
flabel metal1 36790 5633 36817 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VREF
flabel metal1 36753 5694 36779 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VDD
flabel metal1 36751 5114 36775 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VSS
flabel metal1 37311 5633 37338 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VREF
flabel metal1 37349 5694 37375 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VDD
flabel metal1 37353 5114 37377 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VSS
flabel metal1 37046 5633 37073 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VREF
flabel metal1 37009 5694 37035 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VDD
flabel metal1 37007 5114 37031 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VSS
flabel metal1 37567 5633 37594 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VREF
flabel metal1 37605 5694 37631 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VDD
flabel metal1 37609 5114 37633 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VSS
flabel metal1 37302 5633 37329 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VREF
flabel metal1 37265 5694 37291 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VDD
flabel metal1 37263 5114 37287 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VSS
flabel metal1 29631 5633 29658 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF
flabel metal1 29669 5694 29695 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD
flabel metal1 29673 5114 29697 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VSS
flabel metal1 29366 5633 29393 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VREF
flabel metal1 29329 5694 29355 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VDD
flabel metal1 29327 5114 29351 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VSS
flabel metal1 29887 5633 29914 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VREF
flabel metal1 29925 5694 29951 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VDD
flabel metal1 29929 5114 29953 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VSS
flabel metal1 29622 5633 29649 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VREF
flabel metal1 29585 5694 29611 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VDD
flabel metal1 29583 5114 29607 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VSS
flabel metal1 30143 5633 30170 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VREF
flabel metal1 30181 5694 30207 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VDD
flabel metal1 30185 5114 30209 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VSS
flabel metal1 29878 5633 29905 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VREF
flabel metal1 29841 5694 29867 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VDD
flabel metal1 29839 5114 29863 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VSS
flabel metal1 30399 5633 30426 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VREF
flabel metal1 30437 5694 30463 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VDD
flabel metal1 30441 5114 30465 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VSS
flabel metal1 30134 5633 30161 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VREF
flabel metal1 30097 5694 30123 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VDD
flabel metal1 30095 5114 30119 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VSS
flabel metal1 30655 5633 30682 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VREF
flabel metal1 30693 5694 30719 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VDD
flabel metal1 30697 5114 30721 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VSS
flabel metal1 30390 5633 30417 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VREF
flabel metal1 30353 5694 30379 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VDD
flabel metal1 30351 5114 30375 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VSS
flabel metal1 30911 5633 30938 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VREF
flabel metal1 30949 5694 30975 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VDD
flabel metal1 30953 5114 30977 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VSS
flabel metal1 30646 5633 30673 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VREF
flabel metal1 30609 5694 30635 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VDD
flabel metal1 30607 5114 30631 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VSS
flabel metal1 31167 5633 31194 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VREF
flabel metal1 31205 5694 31231 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VDD
flabel metal1 31209 5114 31233 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VSS
flabel metal1 30902 5633 30929 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VREF
flabel metal1 30865 5694 30891 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VDD
flabel metal1 30863 5114 30887 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VSS
flabel metal1 31423 5633 31450 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VREF
flabel metal1 31461 5694 31487 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VDD
flabel metal1 31465 5114 31489 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VSS
flabel metal1 31158 5633 31185 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VREF
flabel metal1 31121 5694 31147 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VDD
flabel metal1 31119 5114 31143 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VSS
flabel metal1 31679 5633 31706 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF
flabel metal1 31717 5694 31743 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD
flabel metal1 31721 5114 31745 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VSS
flabel metal1 31414 5633 31441 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VREF
flabel metal1 31377 5694 31403 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VDD
flabel metal1 31375 5114 31399 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VSS
flabel metal1 31935 5633 31962 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VREF
flabel metal1 31973 5694 31999 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VDD
flabel metal1 31977 5114 32001 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VSS
flabel metal1 31670 5633 31697 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VREF
flabel metal1 31633 5694 31659 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VDD
flabel metal1 31631 5114 31655 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VSS
flabel metal1 32191 5633 32218 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VREF
flabel metal1 32229 5694 32255 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VDD
flabel metal1 32233 5114 32257 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VSS
flabel metal1 31926 5633 31953 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VREF
flabel metal1 31889 5694 31915 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VDD
flabel metal1 31887 5114 31911 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VSS
flabel metal1 32447 5633 32474 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VREF
flabel metal1 32485 5694 32511 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VDD
flabel metal1 32489 5114 32513 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VSS
flabel metal1 32182 5633 32209 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VREF
flabel metal1 32145 5694 32171 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VDD
flabel metal1 32143 5114 32167 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VSS
flabel metal1 32703 5633 32730 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VREF
flabel metal1 32741 5694 32767 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VDD
flabel metal1 32745 5114 32769 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VSS
flabel metal1 32438 5633 32465 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VREF
flabel metal1 32401 5694 32427 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VDD
flabel metal1 32399 5114 32423 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VSS
flabel metal1 32959 5633 32986 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VREF
flabel metal1 32997 5694 33023 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VDD
flabel metal1 33001 5114 33025 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VSS
flabel metal1 32694 5633 32721 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VREF
flabel metal1 32657 5694 32683 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VDD
flabel metal1 32655 5114 32679 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VSS
flabel metal1 33215 5633 33242 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VREF
flabel metal1 33253 5694 33279 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VDD
flabel metal1 33257 5114 33281 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VSS
flabel metal1 32950 5633 32977 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VREF
flabel metal1 32913 5694 32939 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VDD
flabel metal1 32911 5114 32935 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VSS
flabel metal1 33471 5633 33498 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VREF
flabel metal1 33509 5694 33535 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VDD
flabel metal1 33513 5114 33537 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VSS
flabel metal1 33206 5633 33233 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VREF
flabel metal1 33169 5694 33195 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VDD
flabel metal1 33167 5114 33191 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VSS
<< end >>
