magic
tech sky130A
timestamp 1697024547
<< checkpaint >>
rect -649 1202 787 1226
rect -649 1178 1082 1202
rect -649 1154 1239 1178
rect -649 1130 1396 1154
rect -649 1106 1553 1130
rect -649 1082 1848 1106
rect -649 1058 2143 1082
rect -649 1034 2438 1058
rect -649 1010 2917 1034
rect -649 986 3396 1010
rect -649 962 3875 986
rect -649 938 4354 962
rect -649 914 4511 938
rect -649 890 4990 914
rect -649 866 5469 890
rect -649 842 5626 866
rect -649 -354 5783 842
rect -630 -498 5783 -354
rect -630 -1830 730 -498
rect 864 -522 5783 -498
rect 1159 -546 5783 -522
rect 1638 -570 5783 -546
rect 2117 -594 5783 -570
rect 2596 -618 5783 -594
rect 3075 -642 5783 -618
rect 3232 -666 5783 -642
rect 3711 -690 5783 -666
rect 4190 -714 5783 -690
rect 4347 -738 5783 -714
<< metal1 >>
rect 0 0 100 100
rect 0 -200 100 -100
rect 0 -400 100 -300
rect 0 -600 100 -500
rect 0 -800 100 -700
rect 0 -1000 100 -900
rect 0 -1200 100 -1100
use sky130_fd_sc_hd__inv_1  x1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 3724 0 1 12
box -19 -24 157 296
use sky130_fd_sc_hd__buf_4  x2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 157 0 1 276
box -19 -24 295 296
use sky130_fd_sc_hd__dlymetal6s6s_1  x3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 1808 0 1 108
box -19 -24 479 296
use sky130_fd_sc_hd__buf_4  x4
timestamp 1683767628
transform 1 0 923 0 1 180
box -19 -24 295 296
use sky130_fd_sc_hd__inv_1  x5
timestamp 1683767628
transform 1 0 452 0 1 252
box -19 -24 157 296
use sky130_fd_sc_hd__dlymetal6s6s_1  x6
timestamp 1683767628
transform 1 0 2766 0 1 60
box -19 -24 479 296
use sky130_fd_sc_hd__buf_4  x7
timestamp 1683767628
transform 1 0 1218 0 1 156
box -19 -24 295 296
use sky130_fd_sc_hd__buf_4  x8
timestamp 1683767628
transform 1 0 1513 0 1 132
box -19 -24 295 296
use sky130_fd_sc_hd__dlymetal6s6s_1  x9
timestamp 1683767628
transform 1 0 3881 0 1 -12
box -19 -24 479 296
use sky130_fd_sc_hd__dlymetal6s6s_1  x10
timestamp 1683767628
transform 1 0 2287 0 1 84
box -19 -24 479 296
use sky130_fd_sc_hd__inv_1  x11
timestamp 1683767628
transform 1 0 609 0 1 228
box -19 -24 157 296
use sky130_fd_sc_hd__inv_1  x12
timestamp 1683767628
transform 1 0 766 0 1 204
box -19 -24 157 296
use sky130_fd_sc_hd__dlymetal6s6s_1  x13
timestamp 1683767628
transform 1 0 3245 0 1 36
box -19 -24 479 296
use sky130_fd_sc_hd__dlymetal6s6s_1  x14
timestamp 1683767628
transform 1 0 4360 0 1 -36
box -19 -24 479 296
use sky130_fd_sc_hd__nand2_1  x15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 4839 0 1 -60
box -19 -24 157 296
use sky130_fd_sc_hd__nand2_1  x16
timestamp 1683767628
transform 1 0 4996 0 1 -84
box -19 -24 157 296
use sky130_fd_sc_hd__inv_1  x23
timestamp 1683767628
transform 1 0 0 0 1 300
box -19 -24 157 296
<< labels >>
flabel metal1 0 0 100 100 0 FreeSans 128 0 0 0 VDD
port 0 nsew
flabel metal1 0 -200 100 -100 0 FreeSans 128 0 0 0 VSS
port 1 nsew
flabel metal1 0 -400 100 -300 0 FreeSans 128 0 0 0 phi2_n
port 2 nsew
flabel metal1 0 -600 100 -500 0 FreeSans 128 0 0 0 phi2
port 3 nsew
flabel metal1 0 -800 100 -700 0 FreeSans 128 0 0 0 phi1
port 4 nsew
flabel metal1 0 -1000 100 -900 0 FreeSans 128 0 0 0 phi1_n
port 5 nsew
flabel metal1 0 -1200 100 -1100 0 FreeSans 128 0 0 0 clk
port 6 nsew
<< end >>
