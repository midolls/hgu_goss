magic
tech sky130A
magscale 1 2
timestamp 1698609214
use inv_16_test  inv_16_test_0
timestamp 1698608947
transform 1 0 394 0 1 -2362
box 1014 2362 2652 3027
use inv_16_test  inv_16_test_1
timestamp 1698608947
transform 1 0 -1014 0 1 -2362
box 1014 2362 2652 3027
<< end >>
