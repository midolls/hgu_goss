magic
tech sky130A
magscale 1 2
timestamp 1698581447
<< nmos >>
rect -63 -42 -33 42
rect 33 -42 63 42
<< ndiff >>
rect -125 30 -63 42
rect -125 -30 -113 30
rect -79 -30 -63 30
rect -125 -42 -63 -30
rect -33 30 33 42
rect -33 -30 -17 30
rect 17 -30 33 30
rect -33 -42 33 -30
rect 63 30 125 42
rect 63 -30 79 30
rect 113 -30 125 30
rect 63 -42 125 -30
<< ndiffc >>
rect -113 -30 -79 30
rect -17 -30 17 30
rect 79 -30 113 30
<< poly >>
rect -63 42 -33 68
rect 33 42 63 68
rect -63 -57 -33 -42
rect 33 -57 63 -42
rect -63 -64 63 -57
rect -81 -87 63 -64
rect -81 -130 -15 -87
<< locali >>
rect -113 30 -79 46
rect -113 -46 -79 -30
rect -17 30 17 84
rect -17 -46 17 -30
rect 79 30 113 46
rect 79 -46 113 -30
<< viali >>
rect -113 -30 -79 30
rect 79 -30 113 30
<< metal1 >>
rect -119 30 119 42
rect -119 -30 -113 30
rect -79 -30 79 30
rect 113 -30 119 30
rect -119 -43 119 -30
<< properties >>
string FIXED_BBOX -210 -199 210 199
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.42 l 0.15 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
