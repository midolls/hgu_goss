magic
tech sky130A
magscale 1 2
timestamp 1697025759
<< error_p >>
rect -29 241 29 247
rect -29 207 -17 241
rect -29 201 29 207
rect -29 -207 29 -201
rect -29 -241 -17 -207
rect -29 -247 29 -241
<< nwell >>
rect -211 -379 211 379
<< pmos >>
rect -15 -160 15 160
<< pdiff >>
rect -73 148 -15 160
rect -73 -148 -61 148
rect -27 -148 -15 148
rect -73 -160 -15 -148
rect 15 148 73 160
rect 15 -148 27 148
rect 61 -148 73 148
rect 15 -160 73 -148
<< pdiffc >>
rect -61 -148 -27 148
rect 27 -148 61 148
<< nsubdiff >>
rect -175 309 -79 343
rect 79 309 175 343
rect -175 247 -141 309
rect 141 247 175 309
rect -175 -309 -141 -247
rect 141 -309 175 -247
rect -175 -343 -79 -309
rect 79 -343 175 -309
<< nsubdiffcont >>
rect -79 309 79 343
rect -175 -247 -141 247
rect 141 -247 175 247
rect -79 -343 79 -309
<< poly >>
rect -33 241 33 257
rect -33 207 -17 241
rect 17 207 33 241
rect -33 191 33 207
rect -15 160 15 191
rect -15 -191 15 -160
rect -33 -207 33 -191
rect -33 -241 -17 -207
rect 17 -241 33 -207
rect -33 -257 33 -241
<< polycont >>
rect -17 207 17 241
rect -17 -241 17 -207
<< locali >>
rect -175 309 -79 343
rect 79 309 175 343
rect -175 247 -141 309
rect 141 247 175 309
rect -33 207 -17 241
rect 17 207 33 241
rect -61 148 -27 164
rect -61 -164 -27 -148
rect 27 148 61 164
rect 27 -164 61 -148
rect -33 -241 -17 -207
rect 17 -241 33 -207
rect -175 -309 -141 -247
rect 141 -309 175 -247
rect -175 -343 -79 -309
rect 79 -343 175 -309
<< viali >>
rect -17 207 17 241
rect -61 -148 -27 148
rect 27 -148 61 148
rect -17 -241 17 -207
<< metal1 >>
rect -29 241 29 247
rect -29 207 -17 241
rect 17 207 29 241
rect -29 201 29 207
rect -67 148 -21 160
rect -67 -148 -61 148
rect -27 -148 -21 148
rect -67 -160 -21 -148
rect 21 148 67 160
rect 21 -148 27 148
rect 61 -148 67 148
rect 21 -160 67 -148
rect -29 -207 29 -201
rect -29 -241 -17 -207
rect 17 -241 29 -207
rect -29 -247 29 -241
<< properties >>
string FIXED_BBOX -158 -326 158 326
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.6 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
