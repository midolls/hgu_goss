magic
tech sky130A
magscale 1 2
timestamp 1698584986
<< error_p >>
rect 305 719 363 725
rect 305 685 317 719
rect 305 679 363 685
<< nwell >>
rect 49 897 341 900
rect 49 730 443 897
rect 225 729 443 730
<< pmoshvt >>
rect 144 766 174 852
rect 216 766 246 852
rect 319 766 349 850
<< pdiff >>
rect 86 839 144 852
rect 86 779 97 839
rect 131 779 144 839
rect 86 766 144 779
rect 174 766 216 852
rect 246 850 304 852
rect 246 766 319 850
rect 349 838 407 850
rect 349 778 361 838
rect 395 778 407 838
rect 349 766 407 778
<< pdiffc >>
rect 97 779 131 839
rect 361 778 395 838
<< poly >>
rect 144 852 174 883
rect 216 852 246 883
rect 319 850 349 880
rect 144 751 174 766
rect 216 751 246 766
rect 319 751 349 766
rect 144 735 349 751
rect 144 721 367 735
rect 301 719 367 721
rect 301 685 317 719
rect 351 685 367 719
rect 301 669 367 685
<< polycont >>
rect 317 685 351 719
<< locali >>
rect 97 839 131 856
rect 97 763 131 779
rect 361 838 395 854
rect 361 762 395 778
rect 301 685 317 719
rect 351 685 367 719
<< viali >>
rect 361 778 395 838
rect 317 685 351 719
<< metal1 >>
rect 355 838 401 850
rect 355 778 361 838
rect 395 778 401 838
rect 355 766 401 778
rect 305 719 363 725
rect 305 685 317 719
rect 351 685 363 719
rect 305 679 363 685
<< end >>
