magic
tech sky130A
magscale 1 2
timestamp 1700938627
<< nwell >>
rect 433 5763 438 5795
<< psubdiff >>
rect 2878 6266 2936 6312
rect 5397 6266 5429 6312
rect -109 5106 565 5152
rect 4598 5106 8013 5152
rect 10187 5106 15777 5152
rect 19999 5106 29321 5152
<< poly >>
rect -271 5997 -201 6129
rect 657 5978 727 6110
rect 1409 6013 1863 6083
rect 3028 6013 3994 6083
rect 5521 6013 7511 6083
rect 10608 6023 14646 6093
rect 20445 6013 28579 6083
rect -271 5290 -201 5422
rect 657 5290 727 5422
rect 1921 5335 2375 5405
rect 3540 5335 4506 5405
rect 8105 5335 10095 5405
rect 15869 5335 19907 5405
rect 29413 5335 37547 5405
<< locali >>
rect -109 6266 437 6312
rect 818 6266 1345 6312
rect 1955 6266 2936 6312
rect 4086 6266 5429 6312
rect 7603 6266 10516 6312
rect 14738 6266 23329 6312
rect -109 5686 565 5732
rect 947 5686 1829 5732
rect 2467 5686 3448 5732
rect 4598 5686 8013 5732
rect 10187 5686 15777 5732
rect 19393 5686 23292 5732
rect 28671 5686 29321 5732
rect -109 5106 565 5152
rect 947 5106 1829 5152
rect 2467 5106 3448 5152
rect 4598 5106 8013 5152
rect 10187 5106 15777 5152
rect 19999 5106 29321 5152
<< metal1 >>
rect 38407 6316 38471 6322
rect 38407 6314 38413 6316
rect -116 6264 440 6314
rect 818 6264 1345 6314
rect 1954 6264 2936 6314
rect 4086 6264 5429 6314
rect 7603 6264 10516 6314
rect 14738 6264 23329 6314
rect 28671 6264 38413 6314
rect 38465 6264 38471 6316
rect 38407 6258 38471 6264
rect 1268 6109 1332 6115
rect -95 6083 -31 6089
rect -95 6073 -89 6083
rect -155 6040 -89 6073
rect -95 6031 -89 6040
rect -37 6031 -31 6083
rect -95 6025 -31 6031
rect 357 6066 421 6072
rect 357 6014 363 6066
rect 415 6060 421 6066
rect 415 6024 611 6060
rect 1268 6057 1274 6109
rect 1326 6099 1332 6109
rect 2803 6112 2867 6118
rect 1326 6068 1553 6099
rect 1874 6094 1938 6100
rect 1874 6083 1880 6094
rect 1326 6057 1332 6068
rect 1268 6051 1332 6057
rect 1747 6054 1880 6083
rect 1874 6042 1880 6054
rect 1932 6042 1938 6094
rect 2803 6060 2809 6112
rect 2861 6099 2867 6112
rect 5353 6110 5417 6116
rect 2861 6070 3110 6099
rect 4015 6094 4079 6100
rect 4015 6086 4021 6094
rect 2861 6060 2867 6070
rect 2803 6054 2867 6060
rect 3912 6051 4021 6086
rect 1874 6036 1938 6042
rect 4015 6042 4021 6051
rect 4073 6042 4079 6094
rect 5353 6058 5359 6110
rect 5411 6099 5417 6110
rect 10326 6107 10390 6113
rect 5411 6061 5603 6099
rect 5960 6094 6024 6100
rect 5411 6058 5417 6061
rect 5353 6052 5417 6058
rect 4015 6036 4079 6042
rect 5960 6042 5966 6094
rect 6018 6042 6024 6094
rect 5960 6036 6024 6042
rect 6565 6094 6629 6100
rect 6565 6042 6571 6094
rect 6623 6042 6629 6094
rect 6565 6036 6629 6042
rect 7171 6093 7235 6099
rect 7171 6041 7177 6093
rect 7229 6041 7235 6093
rect 7777 6092 7841 6098
rect 7777 6091 7783 6092
rect 7429 6044 7783 6091
rect 7171 6035 7235 6041
rect 7777 6040 7783 6044
rect 7835 6040 7841 6092
rect 10326 6055 10332 6107
rect 10384 6097 10390 6107
rect 10384 6067 10690 6097
rect 10932 6094 10996 6100
rect 10384 6055 10390 6067
rect 10326 6049 10390 6055
rect 7777 6034 7841 6040
rect 10932 6042 10938 6094
rect 10990 6042 10996 6094
rect 10932 6036 10996 6042
rect 11538 6093 11602 6099
rect 11538 6041 11544 6093
rect 11596 6041 11602 6093
rect 11538 6035 11602 6041
rect 12172 6093 12236 6099
rect 12172 6041 12178 6093
rect 12230 6041 12236 6093
rect 12172 6035 12236 6041
rect 12750 6093 12814 6099
rect 14529 6093 14628 6099
rect 12750 6041 12756 6093
rect 12808 6041 12814 6093
rect 12750 6035 12814 6041
rect 13356 6087 13420 6093
rect 13356 6035 13362 6087
rect 13414 6035 13420 6087
rect 13356 6029 13420 6035
rect 13962 6087 14026 6093
rect 13962 6035 13968 6087
rect 14020 6035 14026 6087
rect 14529 6070 14570 6093
rect 14564 6041 14570 6070
rect 14622 6041 14628 6093
rect 14564 6035 14628 6041
rect 20149 6097 20213 6103
rect 20149 6045 20155 6097
rect 20207 6045 20213 6097
rect 20756 6092 20820 6098
rect 20756 6081 20762 6092
rect 20755 6052 20762 6081
rect 20149 6039 20213 6045
rect 20756 6040 20762 6052
rect 20814 6040 20820 6092
rect 21361 6092 21425 6098
rect 21361 6081 21367 6092
rect 21360 6052 21367 6081
rect 13962 6029 14026 6035
rect 20756 6034 20820 6040
rect 21361 6040 21367 6052
rect 21419 6040 21425 6092
rect 21968 6093 22032 6099
rect 21968 6082 21974 6093
rect 21967 6053 21974 6082
rect 21361 6034 21425 6040
rect 21968 6041 21974 6053
rect 22026 6041 22032 6093
rect 22574 6093 22638 6099
rect 22574 6082 22580 6093
rect 22573 6053 22580 6082
rect 21968 6035 22032 6041
rect 22574 6041 22580 6053
rect 22632 6041 22638 6093
rect 23180 6094 23244 6100
rect 23180 6083 23186 6094
rect 23179 6054 23186 6083
rect 22574 6035 22638 6041
rect 23180 6042 23186 6054
rect 23238 6042 23244 6094
rect 23792 6093 23856 6099
rect 23792 6082 23798 6093
rect 23791 6053 23798 6082
rect 23180 6036 23244 6042
rect 23792 6041 23798 6053
rect 23850 6041 23856 6093
rect 23792 6035 23856 6041
rect 24997 6093 25061 6099
rect 24997 6041 25003 6093
rect 25055 6041 25061 6093
rect 24997 6035 25061 6041
rect 25603 6093 25667 6099
rect 25603 6041 25609 6093
rect 25661 6041 25667 6093
rect 25603 6035 25667 6041
rect 26191 6092 26255 6098
rect 26191 6040 26197 6092
rect 26249 6040 26255 6092
rect 26191 6034 26255 6040
rect 26816 6093 26880 6099
rect 26816 6041 26822 6093
rect 26874 6041 26880 6093
rect 26816 6035 26880 6041
rect 27423 6093 27487 6099
rect 27423 6041 27429 6093
rect 27481 6041 27487 6093
rect 27423 6035 27487 6041
rect 28028 6094 28092 6100
rect 28028 6042 28034 6094
rect 28086 6042 28092 6094
rect 28447 6093 28696 6099
rect 28447 6070 28638 6093
rect 28028 6036 28092 6042
rect 28632 6041 28638 6070
rect 28690 6041 28696 6093
rect 28632 6035 28696 6041
rect 415 6014 421 6024
rect 357 6008 421 6014
rect 37698 5820 37762 5826
rect 37698 5795 37704 5820
rect -109 5763 438 5795
rect 819 5763 1346 5795
rect 1954 5763 2936 5795
rect 4086 5763 5429 5795
rect 7603 5763 10516 5795
rect 14738 5763 20353 5795
rect 28671 5768 37704 5795
rect 37756 5768 37762 5820
rect 28671 5763 37762 5768
rect 37698 5762 37762 5763
rect 38683 5736 38747 5742
rect 38683 5734 38689 5736
rect -109 5684 565 5734
rect 947 5684 1829 5734
rect 2467 5684 3448 5734
rect 4598 5684 8013 5734
rect 10187 5684 15777 5734
rect 19393 5732 19870 5734
rect 22898 5732 23292 5734
rect 19393 5686 23292 5732
rect 19393 5684 19870 5686
rect 22898 5684 23292 5686
rect 28670 5684 29321 5734
rect 31571 5684 31630 5734
rect 35933 5684 36046 5734
rect 36885 5684 36916 5734
rect 37076 5684 37184 5734
rect 37637 5684 38689 5734
rect 38741 5684 38747 5736
rect 38683 5678 38747 5684
rect -109 5623 565 5655
rect 947 5623 1829 5655
rect 2467 5623 3448 5655
rect 4598 5623 8013 5655
rect 10187 5623 15777 5655
rect 19393 5623 19870 5655
rect 19999 5623 29321 5655
rect 31571 5623 31630 5655
rect 35933 5623 36046 5655
rect 36885 5623 36916 5655
rect 37076 5623 37184 5655
rect 37637 5649 37762 5655
rect 37637 5623 37704 5649
rect 37698 5597 37704 5623
rect 37756 5597 37762 5649
rect 37698 5591 37762 5597
rect 962 5401 1026 5407
rect 962 5394 968 5401
rect -95 5363 -31 5369
rect -95 5356 -89 5363
rect -173 5322 -89 5356
rect -95 5311 -89 5322
rect -37 5311 -31 5363
rect 773 5358 968 5394
rect 962 5349 968 5358
rect 1020 5349 1026 5401
rect 8381 5378 8445 5384
rect 3408 5371 3472 5377
rect 2480 5364 2544 5370
rect 962 5343 1026 5349
rect 1750 5358 1814 5364
rect -95 5305 -31 5311
rect 1750 5306 1756 5358
rect 1808 5348 1814 5358
rect 2480 5354 2486 5364
rect 1808 5319 2003 5348
rect 2293 5323 2486 5354
rect 1808 5306 1814 5319
rect 2480 5312 2486 5323
rect 2538 5312 2544 5364
rect 3408 5319 3414 5371
rect 3466 5348 3472 5371
rect 4620 5359 4684 5365
rect 4620 5348 4626 5359
rect 3466 5319 3622 5348
rect 4424 5319 4626 5348
rect 3408 5313 3472 5319
rect 2480 5306 2544 5312
rect 4620 5307 4626 5319
rect 4678 5307 4684 5359
rect 1750 5300 1814 5306
rect 4620 5301 4684 5307
rect 7923 5352 7987 5358
rect 7923 5300 7929 5352
rect 7981 5347 7987 5352
rect 7981 5318 8187 5347
rect 8381 5326 8387 5378
rect 8439 5326 8445 5378
rect 8987 5377 9051 5383
rect 8446 5331 8447 5360
rect 8381 5320 8445 5326
rect 8987 5325 8993 5377
rect 9045 5325 9051 5377
rect 8987 5319 9051 5325
rect 9593 5377 9657 5383
rect 9593 5325 9599 5377
rect 9651 5325 9657 5377
rect 29846 5378 29910 5384
rect 10200 5362 10264 5368
rect 10200 5353 10206 5362
rect 9593 5319 9657 5325
rect 10013 5324 10206 5353
rect 7981 5300 7987 5318
rect 10200 5310 10206 5324
rect 10258 5310 10264 5362
rect 20023 5358 20087 5364
rect 20023 5347 20029 5358
rect 19219 5344 19271 5347
rect 19825 5318 20029 5347
rect 10200 5304 10264 5310
rect 20023 5306 20029 5318
rect 20081 5306 20087 5358
rect 20023 5300 20087 5306
rect 29239 5356 29303 5362
rect 29239 5304 29245 5356
rect 29297 5349 29303 5356
rect 29297 5320 29495 5349
rect 29846 5326 29852 5378
rect 29904 5326 29910 5378
rect 29846 5320 29910 5326
rect 30455 5377 30519 5383
rect 30455 5325 30461 5377
rect 30513 5325 30519 5377
rect 29297 5304 29303 5320
rect 30455 5319 30519 5325
rect 31057 5377 31121 5383
rect 31057 5325 31063 5377
rect 31115 5325 31121 5377
rect 31057 5319 31121 5325
rect 31663 5377 31727 5383
rect 31663 5325 31669 5377
rect 31721 5325 31727 5377
rect 31663 5319 31727 5325
rect 32269 5377 32333 5383
rect 32269 5325 32275 5377
rect 32327 5325 32333 5377
rect 32269 5319 32333 5325
rect 32885 5377 32949 5383
rect 32885 5325 32891 5377
rect 32943 5325 32949 5377
rect 32885 5319 32949 5325
rect 33481 5377 33545 5383
rect 33481 5325 33487 5377
rect 33539 5325 33545 5377
rect 33481 5319 33545 5325
rect 34087 5377 34151 5383
rect 34087 5325 34093 5377
rect 34145 5325 34151 5377
rect 34087 5319 34151 5325
rect 34694 5377 34758 5383
rect 34694 5325 34700 5377
rect 34752 5325 34758 5377
rect 34694 5319 34758 5325
rect 35291 5376 35355 5382
rect 35291 5324 35297 5376
rect 35349 5324 35355 5376
rect 35291 5318 35355 5324
rect 35906 5376 35970 5382
rect 35906 5324 35912 5376
rect 35964 5324 35970 5376
rect 35906 5318 35970 5324
rect 36512 5377 36576 5383
rect 36512 5325 36518 5377
rect 36570 5325 36576 5377
rect 36512 5319 36576 5325
rect 37118 5377 37182 5383
rect 37118 5325 37124 5377
rect 37176 5325 37182 5377
rect 37720 5359 37784 5365
rect 37720 5349 37726 5359
rect 37118 5319 37182 5325
rect 37465 5320 37726 5349
rect 7923 5294 7987 5300
rect 29239 5298 29303 5304
rect 37720 5307 37726 5320
rect 37778 5307 37784 5359
rect 37720 5301 37784 5307
rect 38407 5158 38471 5164
rect 38407 5154 38413 5158
rect -109 5104 565 5154
rect 947 5104 1829 5154
rect 2467 5104 3448 5154
rect 4598 5104 8013 5154
rect 10187 5104 15777 5154
rect 19999 5104 29321 5154
rect 31571 5104 31630 5154
rect 35933 5104 36046 5154
rect 36885 5104 36916 5154
rect 37076 5104 37184 5154
rect 37636 5106 38413 5154
rect 38465 5106 38471 5158
rect 37636 5104 38471 5106
rect 38407 5102 38471 5104
rect 150 4070 210 4078
rect 150 4018 154 4070
rect 206 4018 210 4070
rect 150 4007 210 4018
rect 162 3998 196 4007
rect 5102 3925 5169 3929
rect 5102 3873 5108 3925
rect 5160 3915 5169 3925
rect 5160 3881 5175 3915
rect 5160 3873 5169 3881
rect 5102 3869 5169 3873
rect 358 3085 418 3091
rect 358 3033 362 3085
rect 414 3033 418 3085
rect 358 3024 418 3033
rect 370 3013 404 3024
rect 358 2914 418 2920
rect 358 2862 362 2914
rect 414 2862 418 2914
rect 358 2853 418 2862
rect 1270 2914 1330 2920
rect 1270 2862 1274 2914
rect 1326 2862 1330 2914
rect 1270 2853 1330 2862
rect 1876 2913 1936 2919
rect 1876 2861 1880 2913
rect 1932 2861 1936 2913
rect 370 2842 404 2853
rect 1282 2842 1316 2853
rect 1876 2852 1936 2861
rect 2804 2912 2864 2918
rect 2804 2860 2808 2912
rect 2860 2860 2864 2912
rect 1888 2841 1922 2852
rect 2804 2849 2864 2860
rect 4016 2914 4076 2920
rect 4016 2862 4020 2914
rect 4072 2862 4076 2914
rect 4016 2853 4076 2862
rect 5352 2907 5418 2918
rect 5352 2855 5358 2907
rect 5410 2855 5418 2907
rect 2816 2840 2850 2849
rect 4028 2842 4062 2853
rect 5352 2844 5418 2855
rect 5959 2905 6023 2911
rect 5959 2853 5965 2905
rect 6017 2853 6023 2905
rect 5959 2847 6023 2853
rect 6565 2905 6629 2911
rect 6565 2853 6571 2905
rect 6623 2853 6629 2905
rect 6565 2847 6629 2853
rect 7171 2905 7235 2911
rect 7171 2853 7177 2905
rect 7229 2853 7235 2905
rect 7171 2847 7235 2853
rect 7777 2905 7841 2911
rect 7777 2853 7783 2905
rect 7835 2853 7841 2905
rect 7777 2847 7841 2853
rect 10327 2910 10391 2921
rect 10327 2858 10332 2910
rect 10384 2858 10391 2910
rect 10327 2847 10391 2858
rect 10932 2901 10998 2912
rect 10932 2849 10938 2901
rect 10990 2849 10998 2901
rect 5367 2840 5401 2844
rect 5973 2839 6007 2847
rect 6579 2839 6613 2847
rect 7185 2839 7219 2847
rect 7791 2839 7825 2847
rect 10341 2843 10375 2847
rect 10932 2838 10998 2849
rect 11538 2902 11604 2913
rect 11538 2850 11544 2902
rect 11596 2850 11604 2902
rect 11538 2839 11604 2850
rect 12144 2901 12210 2912
rect 12144 2849 12150 2901
rect 12202 2849 12210 2901
rect 12144 2838 12210 2849
rect 12750 2901 12816 2912
rect 12750 2849 12756 2901
rect 12808 2849 12816 2901
rect 12750 2838 12816 2849
rect 13356 2903 13422 2914
rect 13356 2851 13362 2903
rect 13414 2851 13422 2903
rect 13356 2840 13422 2851
rect 13962 2903 14028 2914
rect 13962 2851 13968 2903
rect 14020 2851 14028 2903
rect 13962 2840 14028 2851
rect 14568 2902 14634 2913
rect 14568 2850 14574 2902
rect 14626 2850 14634 2902
rect 14568 2839 14634 2850
rect 20149 2902 20213 2908
rect 20149 2850 20155 2902
rect 20207 2850 20213 2902
rect 20149 2844 20213 2850
rect 20755 2902 20819 2908
rect 20755 2850 20761 2902
rect 20813 2850 20819 2902
rect 20755 2844 20819 2850
rect 21361 2903 21425 2909
rect 21361 2851 21367 2903
rect 21419 2851 21425 2903
rect 21361 2845 21425 2851
rect 21967 2902 22031 2908
rect 21967 2850 21973 2902
rect 22025 2850 22031 2902
rect 20163 2839 20197 2844
rect 20769 2839 20803 2844
rect 21375 2840 21409 2845
rect 21967 2844 22031 2850
rect 22573 2902 22637 2908
rect 22573 2850 22579 2902
rect 22631 2850 22637 2902
rect 22573 2844 22637 2850
rect 23179 2902 23243 2908
rect 23179 2850 23185 2902
rect 23237 2850 23243 2902
rect 23179 2844 23243 2850
rect 23785 2902 23849 2908
rect 23785 2850 23791 2902
rect 23843 2850 23849 2902
rect 23785 2844 23849 2850
rect 24391 2902 24455 2908
rect 24391 2850 24397 2902
rect 24449 2850 24455 2902
rect 24391 2844 24455 2850
rect 24997 2902 25061 2908
rect 24997 2850 25003 2902
rect 25055 2850 25061 2902
rect 24997 2844 25061 2850
rect 25603 2902 25667 2908
rect 25603 2850 25609 2902
rect 25661 2850 25667 2902
rect 25603 2844 25667 2850
rect 26209 2902 26273 2908
rect 26209 2850 26215 2902
rect 26267 2850 26273 2902
rect 26209 2844 26273 2850
rect 26815 2902 26879 2908
rect 26815 2850 26821 2902
rect 26873 2850 26879 2902
rect 26815 2844 26879 2850
rect 27421 2902 27485 2908
rect 27421 2850 27427 2902
rect 27479 2850 27485 2902
rect 27421 2844 27485 2850
rect 28027 2902 28091 2908
rect 28027 2850 28033 2902
rect 28085 2850 28091 2902
rect 28027 2844 28091 2850
rect 28633 2902 28697 2908
rect 28633 2850 28639 2902
rect 28691 2850 28697 2902
rect 28633 2844 28697 2850
rect 21981 2839 22015 2844
rect 22587 2839 22621 2844
rect 23193 2839 23227 2844
rect 23799 2839 23833 2844
rect 24405 2839 24439 2844
rect 25011 2839 25045 2844
rect 25617 2839 25651 2844
rect 26223 2839 26257 2844
rect 26829 2839 26863 2844
rect 27435 2839 27469 2844
rect 28041 2839 28075 2844
rect 28647 2839 28681 2844
rect -93 1954 -33 1960
rect -93 1902 -89 1954
rect -37 1902 -33 1954
rect -93 1896 -33 1902
rect -81 1882 -47 1896
rect 964 1815 1024 1821
rect 964 1763 968 1815
rect 1020 1763 1024 1815
rect 964 1754 1024 1763
rect 1876 1814 1936 1820
rect 1876 1762 1880 1814
rect 1932 1762 1936 1814
rect 976 1743 1010 1754
rect 1876 1753 1936 1762
rect 2482 1815 2542 1821
rect 2482 1763 2486 1815
rect 2538 1763 2542 1815
rect 7776 1818 7842 1829
rect 2482 1754 2542 1763
rect 3408 1804 3472 1810
rect 1888 1742 1922 1753
rect 2494 1743 2528 1754
rect 3408 1752 3414 1804
rect 3466 1752 3472 1804
rect 3408 1746 3472 1752
rect 4620 1805 4684 1811
rect 4620 1753 4626 1805
rect 4678 1753 4684 1805
rect 4620 1747 4684 1753
rect 5226 1805 5290 1811
rect 5226 1753 5232 1805
rect 5284 1753 5290 1805
rect 7776 1766 7782 1818
rect 7834 1766 7842 1818
rect 7776 1755 7842 1766
rect 8382 1818 8448 1829
rect 8382 1766 8388 1818
rect 8440 1766 8448 1818
rect 8382 1755 8448 1766
rect 8988 1818 9054 1829
rect 8988 1766 8994 1818
rect 9046 1766 9054 1818
rect 8988 1755 9054 1766
rect 9594 1818 9660 1829
rect 15780 1818 15846 1829
rect 9594 1766 9600 1818
rect 9652 1766 9660 1818
rect 9594 1755 9660 1766
rect 10200 1807 10266 1818
rect 10200 1755 10206 1807
rect 10258 1755 10266 1807
rect 15780 1766 15786 1818
rect 15838 1766 15846 1818
rect 15780 1755 15846 1766
rect 16386 1817 16452 1828
rect 16386 1765 16392 1817
rect 16444 1765 16452 1817
rect 5226 1747 5290 1753
rect 3422 1738 3456 1746
rect 4634 1733 4668 1747
rect 5240 1739 5274 1747
rect 10200 1744 10266 1755
rect 16386 1754 16452 1765
rect 16992 1817 17058 1828
rect 16992 1765 16998 1817
rect 17050 1765 17058 1817
rect 16992 1754 17058 1765
rect 17598 1816 17664 1827
rect 17598 1764 17604 1816
rect 17656 1764 17664 1816
rect 17598 1753 17664 1764
rect 18204 1816 18270 1827
rect 18204 1764 18210 1816
rect 18262 1764 18270 1816
rect 18204 1753 18270 1764
rect 18810 1816 18876 1827
rect 18810 1764 18816 1816
rect 18868 1764 18876 1816
rect 18810 1753 18876 1764
rect 19416 1815 19482 1826
rect 19416 1763 19422 1815
rect 19474 1763 19482 1815
rect 19416 1752 19482 1763
rect 20023 1815 20087 1821
rect 20023 1763 20029 1815
rect 20081 1763 20087 1815
rect 20023 1757 20087 1763
rect 29239 1814 29303 1820
rect 29239 1762 29245 1814
rect 29297 1762 29303 1814
rect 20037 1752 20071 1757
rect 29239 1756 29303 1762
rect 29845 1814 29909 1820
rect 29845 1762 29851 1814
rect 29903 1762 29909 1814
rect 29845 1756 29909 1762
rect 30451 1813 30515 1819
rect 30451 1761 30457 1813
rect 30509 1761 30515 1813
rect 29253 1751 29287 1756
rect 29859 1751 29893 1756
rect 30451 1755 30515 1761
rect 31057 1814 31121 1820
rect 31057 1762 31063 1814
rect 31115 1762 31121 1814
rect 31057 1756 31121 1762
rect 31663 1814 31727 1820
rect 31663 1762 31669 1814
rect 31721 1762 31727 1814
rect 31663 1756 31727 1762
rect 32269 1814 32333 1820
rect 32269 1762 32275 1814
rect 32327 1762 32333 1814
rect 32269 1756 32333 1762
rect 32875 1814 32939 1820
rect 32875 1762 32881 1814
rect 32933 1762 32939 1814
rect 32875 1756 32939 1762
rect 33481 1814 33545 1820
rect 33481 1762 33487 1814
rect 33539 1762 33545 1814
rect 33481 1756 33545 1762
rect 34087 1814 34151 1820
rect 34087 1762 34093 1814
rect 34145 1762 34151 1814
rect 34087 1756 34151 1762
rect 34693 1814 34757 1820
rect 34693 1762 34699 1814
rect 34751 1762 34757 1814
rect 34693 1756 34757 1762
rect 35299 1814 35363 1820
rect 35299 1762 35305 1814
rect 35357 1762 35363 1814
rect 35299 1756 35363 1762
rect 35905 1813 35969 1819
rect 35905 1761 35911 1813
rect 35963 1761 35969 1813
rect 30465 1750 30499 1755
rect 31071 1751 31105 1756
rect 31677 1751 31711 1756
rect 32283 1751 32317 1756
rect 32889 1751 32923 1756
rect 33495 1751 33529 1756
rect 34101 1751 34135 1756
rect 34707 1751 34741 1756
rect 35313 1751 35347 1756
rect 35905 1755 35969 1761
rect 36511 1814 36575 1820
rect 36511 1762 36517 1814
rect 36569 1762 36575 1814
rect 36511 1756 36575 1762
rect 37117 1814 37181 1820
rect 37117 1762 37123 1814
rect 37175 1762 37181 1814
rect 37117 1756 37181 1762
rect 37723 1814 37787 1820
rect 37723 1762 37729 1814
rect 37781 1762 37787 1814
rect 37723 1756 37787 1762
rect 35919 1750 35953 1755
rect 36525 1751 36559 1756
rect 37131 1751 37165 1756
rect 37737 1751 37771 1756
rect 10215 1735 10249 1744
rect 964 1669 1024 1675
rect 964 1617 968 1669
rect 1020 1617 1024 1669
rect 964 1608 1024 1617
rect 976 1597 1010 1608
<< via1 >>
rect 38413 6264 38465 6316
rect -89 6031 -37 6083
rect 363 6014 415 6066
rect 1274 6057 1326 6109
rect 1880 6042 1932 6094
rect 2809 6060 2861 6112
rect 4021 6042 4073 6094
rect 5359 6058 5411 6110
rect 5966 6042 6018 6094
rect 6571 6042 6623 6094
rect 7177 6041 7229 6093
rect 7783 6040 7835 6092
rect 10332 6055 10384 6107
rect 10938 6042 10990 6094
rect 11544 6041 11596 6093
rect 12178 6041 12230 6093
rect 12756 6041 12808 6093
rect 13362 6035 13414 6087
rect 13968 6035 14020 6087
rect 14570 6041 14622 6093
rect 20155 6045 20207 6097
rect 20762 6040 20814 6092
rect 21367 6040 21419 6092
rect 21974 6041 22026 6093
rect 22580 6041 22632 6093
rect 23186 6042 23238 6094
rect 23798 6041 23850 6093
rect 25003 6041 25055 6093
rect 25609 6041 25661 6093
rect 26197 6040 26249 6092
rect 26822 6041 26874 6093
rect 27429 6041 27481 6093
rect 28034 6042 28086 6094
rect 28638 6041 28690 6093
rect 37704 5768 37756 5820
rect 38689 5684 38741 5736
rect 37704 5597 37756 5649
rect -89 5311 -37 5363
rect 968 5349 1020 5401
rect 1756 5306 1808 5358
rect 2486 5312 2538 5364
rect 3414 5319 3466 5371
rect 4626 5307 4678 5359
rect 7929 5300 7981 5352
rect 8387 5326 8439 5378
rect 8993 5325 9045 5377
rect 9599 5325 9651 5377
rect 10206 5310 10258 5362
rect 20029 5306 20081 5358
rect 29245 5304 29297 5356
rect 29852 5326 29904 5378
rect 30461 5325 30513 5377
rect 31063 5325 31115 5377
rect 31669 5325 31721 5377
rect 32275 5325 32327 5377
rect 32891 5325 32943 5377
rect 33487 5325 33539 5377
rect 34093 5325 34145 5377
rect 34700 5325 34752 5377
rect 35297 5324 35349 5376
rect 35912 5324 35964 5376
rect 36518 5325 36570 5377
rect 37124 5325 37176 5377
rect 37726 5307 37778 5359
rect 38413 5106 38465 5158
rect 154 4018 206 4070
rect 5108 3873 5160 3925
rect 362 3033 414 3085
rect 362 2862 414 2914
rect 1274 2862 1326 2914
rect 1880 2861 1932 2913
rect 2808 2860 2860 2912
rect 4020 2862 4072 2914
rect 5358 2855 5410 2907
rect 5965 2853 6017 2905
rect 6571 2853 6623 2905
rect 7177 2853 7229 2905
rect 7783 2853 7835 2905
rect 10332 2858 10384 2910
rect 10938 2849 10990 2901
rect 11544 2850 11596 2902
rect 12150 2849 12202 2901
rect 12756 2849 12808 2901
rect 13362 2851 13414 2903
rect 13968 2851 14020 2903
rect 14574 2850 14626 2902
rect 20155 2850 20207 2902
rect 20761 2850 20813 2902
rect 21367 2851 21419 2903
rect 21973 2850 22025 2902
rect 22579 2850 22631 2902
rect 23185 2850 23237 2902
rect 23791 2850 23843 2902
rect 24397 2850 24449 2902
rect 25003 2850 25055 2902
rect 25609 2850 25661 2902
rect 26215 2850 26267 2902
rect 26821 2850 26873 2902
rect 27427 2850 27479 2902
rect 28033 2850 28085 2902
rect 28639 2850 28691 2902
rect -89 1902 -37 1954
rect 968 1763 1020 1815
rect 1880 1762 1932 1814
rect 2486 1763 2538 1815
rect 3414 1752 3466 1804
rect 4626 1753 4678 1805
rect 5232 1753 5284 1805
rect 7782 1766 7834 1818
rect 8388 1766 8440 1818
rect 8994 1766 9046 1818
rect 9600 1766 9652 1818
rect 10206 1755 10258 1807
rect 15786 1766 15838 1818
rect 16392 1765 16444 1817
rect 16998 1765 17050 1817
rect 17604 1764 17656 1816
rect 18210 1764 18262 1816
rect 18816 1764 18868 1816
rect 19422 1763 19474 1815
rect 20029 1763 20081 1815
rect 29245 1762 29297 1814
rect 29851 1762 29903 1814
rect 30457 1761 30509 1813
rect 31063 1762 31115 1814
rect 31669 1762 31721 1814
rect 32275 1762 32327 1814
rect 32881 1762 32933 1814
rect 33487 1762 33539 1814
rect 34093 1762 34145 1814
rect 34699 1762 34751 1814
rect 35305 1762 35357 1814
rect 35911 1761 35963 1813
rect 36517 1762 36569 1814
rect 37123 1762 37175 1814
rect 37729 1762 37781 1814
rect 968 1617 1020 1669
<< metal2 >>
rect 38407 6316 38471 6322
rect 38407 6264 38413 6316
rect 38465 6264 38471 6316
rect 38407 6258 38471 6264
rect -95 6198 210 6254
rect -95 6083 -31 6198
rect -95 6031 -89 6083
rect -37 6031 -31 6083
rect -95 6025 -31 6031
rect -95 5363 -31 5369
rect -95 5311 -89 5363
rect -37 5311 -31 5363
rect -95 5305 -31 5311
rect -93 1960 -31 5305
rect 150 4072 210 6198
rect 1268 6109 1332 6115
rect 357 6066 421 6072
rect 357 6014 363 6066
rect 415 6014 421 6066
rect 1268 6057 1274 6109
rect 1326 6057 1332 6109
rect 2803 6112 2867 6118
rect 1268 6051 1332 6057
rect 1874 6094 1938 6100
rect 357 6008 421 6014
rect 150 4016 152 4072
rect 208 4016 210 4072
rect 150 4007 210 4016
rect 363 3096 414 6008
rect 962 5401 1026 5407
rect 962 5349 968 5401
rect 1020 5349 1026 5401
rect 962 5343 1026 5349
rect 358 3087 418 3096
rect 358 3031 360 3087
rect 416 3031 418 3087
rect 358 3022 418 3031
rect 363 2925 414 3022
rect 358 2916 418 2925
rect 358 2860 360 2916
rect 416 2860 418 2916
rect 358 2851 418 2860
rect -93 1956 -33 1960
rect -93 1900 -91 1956
rect -35 1900 -33 1956
rect -93 1891 -33 1900
rect 968 1826 1024 5343
rect 1274 2925 1326 6051
rect 1874 6042 1880 6094
rect 1932 6042 1938 6094
rect 2803 6060 2809 6112
rect 2861 6060 2867 6112
rect 5353 6110 5417 6116
rect 2803 6054 2867 6060
rect 4015 6094 4079 6100
rect 1874 6036 1938 6042
rect 1750 5358 1814 5364
rect 1750 5306 1756 5358
rect 1808 5306 1814 5358
rect 1750 5300 1814 5306
rect 1270 2916 1330 2925
rect 1270 2860 1272 2916
rect 1328 2860 1330 2916
rect 1270 2851 1330 2860
rect 964 1817 1024 1826
rect 964 1761 966 1817
rect 1022 1761 1024 1817
rect 1756 1814 1808 5300
rect 1880 2924 1932 6036
rect 2480 5364 2544 5370
rect 2480 5312 2486 5364
rect 2538 5312 2544 5364
rect 2480 5306 2544 5312
rect 1876 2915 1936 2924
rect 1876 2859 1878 2915
rect 1934 2859 1936 2915
rect 1876 2850 1936 2859
rect 1889 1825 1923 1829
rect 2486 1826 2538 5306
rect 2808 2923 2861 6054
rect 4015 6042 4021 6094
rect 4073 6042 5160 6094
rect 5353 6058 5359 6110
rect 5411 6058 5417 6110
rect 10326 6107 10390 6113
rect 5353 6052 5417 6058
rect 5960 6094 6024 6100
rect 4015 6036 4079 6042
rect 4867 6041 5160 6042
rect 3408 5371 3472 5377
rect 3408 5319 3414 5371
rect 3466 5319 3472 5371
rect 3408 5313 3472 5319
rect 2804 2914 2864 2923
rect 2804 2858 2806 2914
rect 2862 2858 2864 2914
rect 2804 2849 2864 2858
rect 1876 1816 1936 1825
rect 1876 1814 1878 1816
rect 1756 1762 1878 1814
rect 964 1752 1024 1761
rect 968 1680 1024 1752
rect 1876 1760 1878 1762
rect 1934 1760 1936 1816
rect 1876 1751 1936 1760
rect 2482 1817 2542 1826
rect 2482 1761 2484 1817
rect 2540 1761 2542 1817
rect 3414 1815 3466 5313
rect 4020 2925 4073 6036
rect 4620 5359 4684 5365
rect 4620 5307 4626 5359
rect 4678 5307 4684 5359
rect 4620 5301 4684 5307
rect 4016 2916 4076 2925
rect 4016 2860 4018 2916
rect 4074 2860 4076 2916
rect 4016 2851 4076 2860
rect 4626 2017 4678 5301
rect 5108 3929 5160 6041
rect 5097 3927 5171 3929
rect 5097 3926 5106 3927
rect 5094 3873 5106 3926
rect 5097 3871 5106 3873
rect 5162 3871 5171 3927
rect 5097 3869 5171 3871
rect 5358 2918 5411 6052
rect 5960 6042 5966 6094
rect 6018 6042 6024 6094
rect 5960 6036 6024 6042
rect 6565 6094 6629 6100
rect 6565 6042 6571 6094
rect 6623 6042 6629 6094
rect 6565 6036 6629 6042
rect 7171 6093 7235 6099
rect 7171 6041 7177 6093
rect 7229 6041 7235 6093
rect 5352 2909 5418 2918
rect 5965 2916 6018 6036
rect 6571 2916 6624 6036
rect 7171 6035 7235 6041
rect 7777 6092 7841 6098
rect 7777 6040 7783 6092
rect 7835 6040 7841 6092
rect 10326 6055 10332 6107
rect 10384 6055 10390 6107
rect 10326 6049 10390 6055
rect 10932 6094 10996 6100
rect 7177 2916 7230 6035
rect 7777 6034 7841 6040
rect 7783 2916 7836 6034
rect 8381 5378 8445 5384
rect 7923 5352 7987 5358
rect 7923 5300 7929 5352
rect 7981 5300 7987 5352
rect 8381 5326 8387 5378
rect 8439 5326 8445 5378
rect 8381 5320 8445 5326
rect 8987 5377 9051 5383
rect 8987 5325 8993 5377
rect 9045 5325 9051 5377
rect 7923 5294 7987 5300
rect 5352 2853 5357 2909
rect 5413 2853 5418 2909
rect 5352 2844 5418 2853
rect 5959 2907 6023 2916
rect 5959 2851 5963 2907
rect 6019 2851 6023 2907
rect 5959 2842 6023 2851
rect 6565 2907 6629 2916
rect 6565 2851 6569 2907
rect 6625 2851 6629 2907
rect 6565 2842 6629 2851
rect 7171 2907 7235 2916
rect 7171 2851 7175 2907
rect 7231 2851 7235 2907
rect 7171 2842 7235 2851
rect 7777 2907 7841 2916
rect 7777 2851 7781 2907
rect 7837 2851 7841 2907
rect 7777 2842 7841 2851
rect 4626 1965 5284 2017
rect 4626 1816 4678 1965
rect 5232 1816 5284 1965
rect 7776 1820 7842 1829
rect 2482 1752 2542 1761
rect 3408 1806 3472 1815
rect 3408 1750 3412 1806
rect 3468 1750 3472 1806
rect 3408 1741 3472 1750
rect 4620 1807 4684 1816
rect 4620 1751 4624 1807
rect 4680 1751 4684 1807
rect 4620 1742 4684 1751
rect 5226 1807 5290 1816
rect 5226 1751 5230 1807
rect 5286 1751 5290 1807
rect 7776 1764 7781 1820
rect 7837 1818 7842 1820
rect 7930 1818 7982 5294
rect 8388 1829 8440 5320
rect 8987 5319 9051 5325
rect 9593 5377 9657 5383
rect 9593 5325 9599 5377
rect 9651 5325 9657 5377
rect 9593 5319 9657 5325
rect 10200 5362 10264 5368
rect 8994 1829 9046 5319
rect 9600 1829 9652 5319
rect 10200 5310 10206 5362
rect 10258 5310 10264 5362
rect 10200 5304 10264 5310
rect 7837 1766 7982 1818
rect 8382 1820 8448 1829
rect 7837 1764 7842 1766
rect 7776 1755 7842 1764
rect 8382 1764 8387 1820
rect 8443 1764 8448 1820
rect 8382 1755 8448 1764
rect 8988 1820 9054 1829
rect 8988 1764 8993 1820
rect 9049 1764 9054 1820
rect 8988 1755 9054 1764
rect 9594 1820 9660 1829
rect 9594 1764 9599 1820
rect 9655 1764 9660 1820
rect 10206 1818 10258 5304
rect 10332 2921 10384 6049
rect 10932 6042 10938 6094
rect 10990 6042 10996 6094
rect 10932 6036 10996 6042
rect 11538 6093 11602 6099
rect 11538 6041 11544 6093
rect 11596 6041 11602 6093
rect 10327 2912 10391 2921
rect 10938 2912 10990 6036
rect 11538 6035 11602 6041
rect 12150 6093 12236 6099
rect 12150 6041 12178 6093
rect 12230 6041 12236 6093
rect 12150 6035 12236 6041
rect 12750 6093 12814 6099
rect 14564 6093 14628 6099
rect 12750 6041 12756 6093
rect 12808 6041 12814 6093
rect 12750 6035 12814 6041
rect 13356 6087 13420 6093
rect 13356 6035 13362 6087
rect 13414 6035 13420 6087
rect 11544 2913 11596 6035
rect 10327 2856 10331 2912
rect 10387 2856 10391 2912
rect 10327 2847 10391 2856
rect 10932 2903 10998 2912
rect 10932 2847 10937 2903
rect 10993 2847 10998 2903
rect 10932 2838 10998 2847
rect 11538 2904 11604 2913
rect 12150 2912 12202 6035
rect 12756 2912 12808 6035
rect 13356 6029 13420 6035
rect 13962 6087 14026 6093
rect 13962 6035 13968 6087
rect 14020 6035 14026 6087
rect 14564 6041 14570 6093
rect 14622 6041 14628 6093
rect 14564 6035 14628 6041
rect 20149 6097 20213 6103
rect 20149 6045 20155 6097
rect 20207 6045 20213 6097
rect 20149 6039 20213 6045
rect 20756 6092 20820 6098
rect 20756 6040 20762 6092
rect 20814 6040 20820 6092
rect 13962 6029 14026 6035
rect 13362 2914 13414 6029
rect 13968 2914 14020 6029
rect 11538 2848 11543 2904
rect 11599 2848 11604 2904
rect 11538 2839 11604 2848
rect 12144 2903 12210 2912
rect 12144 2847 12149 2903
rect 12205 2847 12210 2903
rect 12144 2838 12210 2847
rect 12750 2903 12816 2912
rect 12750 2847 12755 2903
rect 12811 2847 12816 2903
rect 12750 2838 12816 2847
rect 13356 2905 13422 2914
rect 13356 2849 13361 2905
rect 13417 2849 13422 2905
rect 13356 2840 13422 2849
rect 13962 2905 14028 2914
rect 14574 2913 14626 6035
rect 20023 5358 20087 5364
rect 13962 2849 13967 2905
rect 14023 2849 14028 2905
rect 13962 2840 14028 2849
rect 14568 2904 14634 2913
rect 14568 2848 14573 2904
rect 14629 2848 14634 2904
rect 14568 2839 14634 2848
rect 15786 1829 15838 5307
rect 20023 5306 20029 5358
rect 20081 5306 20087 5358
rect 15780 1820 15846 1829
rect 16392 1828 16444 5306
rect 16998 1828 17050 5306
rect 9594 1755 9660 1764
rect 10200 1809 10266 1818
rect 5226 1742 5290 1751
rect 10200 1753 10205 1809
rect 10261 1753 10266 1809
rect 15780 1764 15785 1820
rect 15841 1764 15846 1820
rect 15780 1755 15846 1764
rect 16386 1819 16452 1828
rect 16386 1763 16391 1819
rect 16447 1763 16452 1819
rect 16386 1754 16452 1763
rect 16992 1819 17058 1828
rect 17604 1827 17656 5305
rect 18210 1827 18262 5305
rect 18816 1827 18868 5305
rect 16992 1763 16997 1819
rect 17053 1763 17058 1819
rect 16992 1754 17058 1763
rect 17598 1818 17664 1827
rect 17598 1762 17603 1818
rect 17659 1762 17664 1818
rect 17598 1753 17664 1762
rect 18204 1818 18270 1827
rect 18204 1762 18209 1818
rect 18265 1762 18270 1818
rect 18204 1753 18270 1762
rect 18810 1818 18876 1827
rect 19422 1826 19474 5304
rect 20023 5300 20087 5306
rect 20029 1826 20081 5300
rect 20155 2913 20208 6039
rect 20756 6034 20820 6040
rect 21361 6092 21425 6098
rect 21361 6040 21367 6092
rect 21419 6040 21425 6092
rect 21361 6034 21425 6040
rect 21968 6093 22032 6099
rect 21968 6041 21974 6093
rect 22026 6041 22032 6093
rect 21968 6035 22032 6041
rect 22574 6093 22638 6099
rect 22574 6041 22580 6093
rect 22632 6041 22638 6093
rect 22574 6035 22638 6041
rect 23180 6094 23244 6100
rect 23180 6042 23186 6094
rect 23238 6042 23244 6094
rect 23792 6093 23856 6099
rect 23792 6062 23798 6093
rect 23180 6036 23244 6042
rect 23791 6041 23798 6062
rect 23850 6041 23856 6093
rect 20761 2913 20814 6034
rect 21367 2914 21420 6034
rect 20149 2904 20213 2913
rect 20149 2848 20153 2904
rect 20209 2848 20213 2904
rect 20149 2839 20213 2848
rect 20755 2904 20819 2913
rect 20755 2848 20759 2904
rect 20815 2848 20819 2904
rect 20755 2839 20819 2848
rect 21361 2905 21425 2914
rect 21973 2913 22026 6035
rect 22579 2913 22632 6035
rect 23185 2913 23238 6036
rect 23791 6035 23856 6041
rect 24997 6093 25061 6099
rect 24997 6041 25003 6093
rect 25055 6041 25061 6093
rect 23791 6034 23850 6035
rect 23791 2913 23844 6034
rect 24397 2913 24450 6039
rect 24997 6035 25061 6041
rect 25603 6093 25667 6099
rect 25603 6041 25609 6093
rect 25661 6041 25667 6093
rect 25603 6035 25667 6041
rect 26191 6092 26268 6098
rect 26191 6040 26197 6092
rect 26249 6040 26268 6092
rect 25003 2913 25056 6035
rect 25609 2913 25662 6035
rect 26191 6034 26268 6040
rect 26816 6093 26880 6099
rect 26816 6041 26822 6093
rect 26874 6041 26880 6093
rect 26816 6035 26880 6041
rect 27423 6093 27487 6099
rect 27423 6041 27429 6093
rect 27481 6041 27487 6093
rect 27423 6035 27487 6041
rect 28028 6094 28092 6100
rect 28028 6042 28034 6094
rect 28086 6042 28092 6094
rect 28028 6036 28092 6042
rect 28632 6093 28696 6099
rect 28632 6041 28638 6093
rect 28690 6041 28696 6093
rect 26215 2913 26268 6034
rect 26821 2913 26874 6035
rect 27427 2913 27480 6035
rect 28033 2913 28086 6036
rect 28632 6035 28696 6041
rect 38413 6078 38465 6258
rect 38520 6078 38595 6080
rect 38413 6071 38595 6078
rect 28638 2913 28691 6035
rect 38413 6015 38529 6071
rect 38585 6015 38595 6071
rect 38413 6008 38595 6015
rect 37698 5820 37762 5826
rect 37698 5768 37704 5820
rect 37756 5768 37762 5820
rect 37698 5762 37762 5768
rect 37713 5734 37747 5762
rect 37806 5744 37915 5753
rect 37806 5734 37849 5744
rect 37713 5688 37849 5734
rect 37905 5688 37915 5744
rect 37713 5683 37915 5688
rect 37713 5655 37747 5683
rect 37806 5679 37915 5683
rect 37698 5649 37762 5655
rect 37698 5597 37704 5649
rect 37756 5597 37762 5649
rect 37698 5591 37762 5597
rect 29846 5378 29910 5384
rect 29239 5356 29303 5362
rect 29239 5304 29245 5356
rect 29297 5304 29303 5356
rect 29846 5326 29852 5378
rect 29904 5326 29910 5378
rect 29846 5320 29910 5326
rect 30455 5377 30519 5383
rect 30455 5325 30461 5377
rect 30513 5325 30519 5377
rect 29239 5298 29303 5304
rect 21361 2849 21365 2905
rect 21421 2849 21425 2905
rect 21361 2840 21425 2849
rect 21967 2904 22031 2913
rect 21967 2848 21971 2904
rect 22027 2848 22031 2904
rect 21967 2839 22031 2848
rect 22573 2904 22637 2913
rect 22573 2848 22577 2904
rect 22633 2848 22637 2904
rect 22573 2839 22637 2848
rect 23179 2904 23243 2913
rect 23179 2848 23183 2904
rect 23239 2848 23243 2904
rect 23179 2839 23243 2848
rect 23785 2904 23849 2913
rect 23785 2848 23789 2904
rect 23845 2848 23849 2904
rect 23785 2839 23849 2848
rect 24391 2904 24455 2913
rect 24391 2848 24395 2904
rect 24451 2848 24455 2904
rect 24391 2839 24455 2848
rect 24997 2904 25061 2913
rect 24997 2848 25001 2904
rect 25057 2848 25061 2904
rect 24997 2839 25061 2848
rect 25603 2904 25667 2913
rect 25603 2848 25607 2904
rect 25663 2848 25667 2904
rect 25603 2839 25667 2848
rect 26209 2904 26273 2913
rect 26209 2848 26213 2904
rect 26269 2848 26273 2904
rect 26209 2839 26273 2848
rect 26815 2904 26879 2913
rect 26815 2848 26819 2904
rect 26875 2848 26879 2904
rect 26815 2839 26879 2848
rect 27421 2904 27485 2913
rect 27421 2848 27425 2904
rect 27481 2848 27485 2904
rect 27421 2839 27485 2848
rect 28027 2904 28091 2913
rect 28027 2848 28031 2904
rect 28087 2848 28091 2904
rect 28027 2839 28091 2848
rect 28633 2904 28697 2913
rect 28633 2848 28637 2904
rect 28693 2848 28697 2904
rect 28633 2839 28697 2848
rect 18810 1762 18815 1818
rect 18871 1762 18876 1818
rect 18810 1753 18876 1762
rect 19416 1817 19482 1826
rect 19416 1761 19421 1817
rect 19477 1761 19482 1817
rect 10200 1744 10266 1753
rect 19416 1752 19482 1761
rect 20023 1817 20087 1826
rect 29245 1825 29297 5298
rect 29851 1825 29903 5320
rect 30455 5319 30519 5325
rect 31057 5377 31121 5383
rect 31057 5325 31063 5377
rect 31115 5325 31121 5377
rect 31057 5319 31121 5325
rect 31663 5377 31727 5383
rect 31663 5325 31669 5377
rect 31721 5325 31727 5377
rect 31663 5319 31727 5325
rect 32269 5377 32333 5383
rect 32269 5325 32275 5377
rect 32327 5325 32333 5377
rect 32269 5319 32333 5325
rect 32885 5377 32949 5383
rect 32885 5325 32891 5377
rect 32943 5325 32949 5377
rect 32885 5320 32949 5325
rect 32881 5319 32949 5320
rect 33481 5377 33545 5383
rect 33481 5325 33487 5377
rect 33539 5325 33545 5377
rect 33481 5319 33545 5325
rect 34087 5377 34151 5383
rect 34087 5325 34093 5377
rect 34145 5325 34151 5377
rect 34087 5319 34151 5325
rect 34694 5377 34758 5383
rect 34694 5325 34700 5377
rect 34752 5325 34758 5377
rect 34694 5319 34758 5325
rect 35291 5376 35355 5382
rect 35291 5324 35297 5376
rect 35349 5324 35355 5376
rect 35291 5320 35355 5324
rect 35906 5376 35970 5382
rect 35906 5324 35912 5376
rect 35964 5324 35970 5376
rect 20023 1761 20027 1817
rect 20083 1761 20087 1817
rect 20023 1752 20087 1761
rect 29239 1816 29303 1825
rect 29239 1760 29243 1816
rect 29299 1760 29303 1816
rect 29239 1751 29303 1760
rect 29845 1816 29909 1825
rect 30457 1824 30509 5319
rect 31063 1825 31115 5319
rect 31669 1825 31721 5319
rect 32275 1825 32327 5319
rect 32881 1825 32933 5319
rect 33487 1825 33539 5319
rect 34093 1825 34145 5319
rect 34699 1825 34751 5319
rect 35291 5318 35357 5320
rect 35906 5318 35970 5324
rect 36512 5377 36576 5383
rect 36512 5325 36518 5377
rect 36570 5325 36576 5377
rect 36512 5319 36576 5325
rect 37118 5377 37182 5383
rect 37118 5325 37124 5377
rect 37176 5325 37182 5377
rect 37118 5319 37182 5325
rect 37720 5359 37784 5365
rect 35305 1825 35357 5318
rect 29845 1760 29849 1816
rect 29905 1760 29909 1816
rect 29845 1751 29909 1760
rect 30451 1815 30515 1824
rect 30451 1759 30455 1815
rect 30511 1759 30515 1815
rect 30451 1750 30515 1759
rect 31057 1816 31121 1825
rect 31057 1760 31061 1816
rect 31117 1760 31121 1816
rect 31057 1751 31121 1760
rect 31663 1816 31727 1825
rect 31663 1760 31667 1816
rect 31723 1760 31727 1816
rect 31663 1751 31727 1760
rect 32269 1816 32333 1825
rect 32269 1760 32273 1816
rect 32329 1760 32333 1816
rect 32269 1751 32333 1760
rect 32875 1816 32939 1825
rect 32875 1760 32879 1816
rect 32935 1760 32939 1816
rect 32875 1751 32939 1760
rect 33481 1816 33545 1825
rect 33481 1760 33485 1816
rect 33541 1760 33545 1816
rect 33481 1751 33545 1760
rect 34087 1816 34151 1825
rect 34087 1760 34091 1816
rect 34147 1760 34151 1816
rect 34087 1751 34151 1760
rect 34693 1816 34757 1825
rect 34693 1760 34697 1816
rect 34753 1760 34757 1816
rect 34693 1751 34757 1760
rect 35299 1816 35363 1825
rect 35911 1824 35963 5318
rect 36517 1825 36569 5319
rect 37123 1825 37175 5319
rect 37720 5307 37726 5359
rect 37778 5307 37784 5359
rect 37720 5301 37784 5307
rect 37729 1825 37781 5301
rect 38413 5164 38465 6008
rect 38520 6006 38595 6008
rect 39085 5745 39160 5747
rect 39081 5744 39160 5745
rect 38683 5738 39160 5744
rect 38683 5736 39094 5738
rect 38683 5684 38689 5736
rect 38741 5684 39094 5736
rect 38683 5682 39094 5684
rect 39150 5682 39160 5738
rect 38683 5676 39160 5682
rect 39081 5675 39160 5676
rect 39085 5673 39160 5675
rect 38407 5158 38471 5164
rect 38407 5106 38413 5158
rect 38465 5106 38471 5158
rect 38407 5102 38471 5106
rect 35299 1760 35303 1816
rect 35359 1760 35363 1816
rect 35299 1751 35363 1760
rect 35905 1815 35969 1824
rect 35905 1759 35909 1815
rect 35965 1759 35969 1815
rect 35905 1750 35969 1759
rect 36511 1816 36575 1825
rect 36511 1760 36515 1816
rect 36571 1760 36575 1816
rect 36511 1751 36575 1760
rect 37117 1816 37181 1825
rect 37117 1760 37121 1816
rect 37177 1760 37181 1816
rect 37117 1751 37181 1760
rect 37723 1816 37787 1825
rect 37723 1760 37727 1816
rect 37783 1760 37787 1816
rect 37723 1751 37787 1760
rect 964 1671 1024 1680
rect 964 1615 966 1671
rect 1022 1615 1024 1671
rect 964 1606 1024 1615
<< via2 >>
rect 152 4070 208 4072
rect 152 4018 154 4070
rect 154 4018 206 4070
rect 206 4018 208 4070
rect 152 4016 208 4018
rect 360 3085 416 3087
rect 360 3033 362 3085
rect 362 3033 414 3085
rect 414 3033 416 3085
rect 360 3031 416 3033
rect 360 2914 416 2916
rect 360 2862 362 2914
rect 362 2862 414 2914
rect 414 2862 416 2914
rect 360 2860 416 2862
rect -91 1954 -35 1956
rect -91 1902 -89 1954
rect -89 1902 -37 1954
rect -37 1902 -35 1954
rect -91 1900 -35 1902
rect 1272 2914 1328 2916
rect 1272 2862 1274 2914
rect 1274 2862 1326 2914
rect 1326 2862 1328 2914
rect 1272 2860 1328 2862
rect 966 1815 1022 1817
rect 966 1763 968 1815
rect 968 1763 1020 1815
rect 1020 1763 1022 1815
rect 966 1761 1022 1763
rect 1878 2913 1934 2915
rect 1878 2861 1880 2913
rect 1880 2861 1932 2913
rect 1932 2861 1934 2913
rect 1878 2859 1934 2861
rect 2806 2912 2862 2914
rect 2806 2860 2808 2912
rect 2808 2860 2860 2912
rect 2860 2860 2862 2912
rect 2806 2858 2862 2860
rect 1878 1814 1934 1816
rect 1878 1762 1880 1814
rect 1880 1762 1932 1814
rect 1932 1762 1934 1814
rect 1878 1760 1934 1762
rect 2484 1815 2540 1817
rect 2484 1763 2486 1815
rect 2486 1763 2538 1815
rect 2538 1763 2540 1815
rect 2484 1761 2540 1763
rect 4018 2914 4074 2916
rect 4018 2862 4020 2914
rect 4020 2862 4072 2914
rect 4072 2862 4074 2914
rect 4018 2860 4074 2862
rect 5106 3925 5162 3927
rect 5106 3873 5108 3925
rect 5108 3873 5160 3925
rect 5160 3873 5162 3925
rect 5106 3871 5162 3873
rect 5357 2907 5413 2909
rect 5357 2855 5358 2907
rect 5358 2855 5410 2907
rect 5410 2855 5413 2907
rect 5357 2853 5413 2855
rect 5963 2905 6019 2907
rect 5963 2853 5965 2905
rect 5965 2853 6017 2905
rect 6017 2853 6019 2905
rect 5963 2851 6019 2853
rect 6569 2905 6625 2907
rect 6569 2853 6571 2905
rect 6571 2853 6623 2905
rect 6623 2853 6625 2905
rect 6569 2851 6625 2853
rect 7175 2905 7231 2907
rect 7175 2853 7177 2905
rect 7177 2853 7229 2905
rect 7229 2853 7231 2905
rect 7175 2851 7231 2853
rect 7781 2905 7837 2907
rect 7781 2853 7783 2905
rect 7783 2853 7835 2905
rect 7835 2853 7837 2905
rect 7781 2851 7837 2853
rect 3412 1804 3468 1806
rect 3412 1752 3414 1804
rect 3414 1752 3466 1804
rect 3466 1752 3468 1804
rect 3412 1750 3468 1752
rect 4624 1805 4680 1807
rect 4624 1753 4626 1805
rect 4626 1753 4678 1805
rect 4678 1753 4680 1805
rect 4624 1751 4680 1753
rect 5230 1805 5286 1807
rect 5230 1753 5232 1805
rect 5232 1753 5284 1805
rect 5284 1753 5286 1805
rect 5230 1751 5286 1753
rect 7781 1818 7837 1820
rect 7781 1766 7782 1818
rect 7782 1766 7834 1818
rect 7834 1766 7837 1818
rect 7781 1764 7837 1766
rect 8387 1818 8443 1820
rect 8387 1766 8388 1818
rect 8388 1766 8440 1818
rect 8440 1766 8443 1818
rect 8387 1764 8443 1766
rect 8993 1818 9049 1820
rect 8993 1766 8994 1818
rect 8994 1766 9046 1818
rect 9046 1766 9049 1818
rect 8993 1764 9049 1766
rect 9599 1818 9655 1820
rect 9599 1766 9600 1818
rect 9600 1766 9652 1818
rect 9652 1766 9655 1818
rect 9599 1764 9655 1766
rect 10331 2910 10387 2912
rect 10331 2858 10332 2910
rect 10332 2858 10384 2910
rect 10384 2858 10387 2910
rect 10331 2856 10387 2858
rect 10937 2901 10993 2903
rect 10937 2849 10938 2901
rect 10938 2849 10990 2901
rect 10990 2849 10993 2901
rect 10937 2847 10993 2849
rect 11543 2902 11599 2904
rect 11543 2850 11544 2902
rect 11544 2850 11596 2902
rect 11596 2850 11599 2902
rect 11543 2848 11599 2850
rect 12149 2901 12205 2903
rect 12149 2849 12150 2901
rect 12150 2849 12202 2901
rect 12202 2849 12205 2901
rect 12149 2847 12205 2849
rect 12755 2901 12811 2903
rect 12755 2849 12756 2901
rect 12756 2849 12808 2901
rect 12808 2849 12811 2901
rect 12755 2847 12811 2849
rect 13361 2903 13417 2905
rect 13361 2851 13362 2903
rect 13362 2851 13414 2903
rect 13414 2851 13417 2903
rect 13361 2849 13417 2851
rect 13967 2903 14023 2905
rect 13967 2851 13968 2903
rect 13968 2851 14020 2903
rect 14020 2851 14023 2903
rect 13967 2849 14023 2851
rect 14573 2902 14629 2904
rect 14573 2850 14574 2902
rect 14574 2850 14626 2902
rect 14626 2850 14629 2902
rect 14573 2848 14629 2850
rect 10205 1807 10261 1809
rect 10205 1755 10206 1807
rect 10206 1755 10258 1807
rect 10258 1755 10261 1807
rect 10205 1753 10261 1755
rect 15785 1818 15841 1820
rect 15785 1766 15786 1818
rect 15786 1766 15838 1818
rect 15838 1766 15841 1818
rect 15785 1764 15841 1766
rect 16391 1817 16447 1819
rect 16391 1765 16392 1817
rect 16392 1765 16444 1817
rect 16444 1765 16447 1817
rect 16391 1763 16447 1765
rect 16997 1817 17053 1819
rect 16997 1765 16998 1817
rect 16998 1765 17050 1817
rect 17050 1765 17053 1817
rect 16997 1763 17053 1765
rect 17603 1816 17659 1818
rect 17603 1764 17604 1816
rect 17604 1764 17656 1816
rect 17656 1764 17659 1816
rect 17603 1762 17659 1764
rect 18209 1816 18265 1818
rect 18209 1764 18210 1816
rect 18210 1764 18262 1816
rect 18262 1764 18265 1816
rect 18209 1762 18265 1764
rect 20153 2902 20209 2904
rect 20153 2850 20155 2902
rect 20155 2850 20207 2902
rect 20207 2850 20209 2902
rect 20153 2848 20209 2850
rect 20759 2902 20815 2904
rect 20759 2850 20761 2902
rect 20761 2850 20813 2902
rect 20813 2850 20815 2902
rect 20759 2848 20815 2850
rect 38529 6015 38585 6071
rect 37849 5688 37905 5744
rect 21365 2903 21421 2905
rect 21365 2851 21367 2903
rect 21367 2851 21419 2903
rect 21419 2851 21421 2903
rect 21365 2849 21421 2851
rect 21971 2902 22027 2904
rect 21971 2850 21973 2902
rect 21973 2850 22025 2902
rect 22025 2850 22027 2902
rect 21971 2848 22027 2850
rect 22577 2902 22633 2904
rect 22577 2850 22579 2902
rect 22579 2850 22631 2902
rect 22631 2850 22633 2902
rect 22577 2848 22633 2850
rect 23183 2902 23239 2904
rect 23183 2850 23185 2902
rect 23185 2850 23237 2902
rect 23237 2850 23239 2902
rect 23183 2848 23239 2850
rect 23789 2902 23845 2904
rect 23789 2850 23791 2902
rect 23791 2850 23843 2902
rect 23843 2850 23845 2902
rect 23789 2848 23845 2850
rect 24395 2902 24451 2904
rect 24395 2850 24397 2902
rect 24397 2850 24449 2902
rect 24449 2850 24451 2902
rect 24395 2848 24451 2850
rect 25001 2902 25057 2904
rect 25001 2850 25003 2902
rect 25003 2850 25055 2902
rect 25055 2850 25057 2902
rect 25001 2848 25057 2850
rect 25607 2902 25663 2904
rect 25607 2850 25609 2902
rect 25609 2850 25661 2902
rect 25661 2850 25663 2902
rect 25607 2848 25663 2850
rect 26213 2902 26269 2904
rect 26213 2850 26215 2902
rect 26215 2850 26267 2902
rect 26267 2850 26269 2902
rect 26213 2848 26269 2850
rect 26819 2902 26875 2904
rect 26819 2850 26821 2902
rect 26821 2850 26873 2902
rect 26873 2850 26875 2902
rect 26819 2848 26875 2850
rect 27425 2902 27481 2904
rect 27425 2850 27427 2902
rect 27427 2850 27479 2902
rect 27479 2850 27481 2902
rect 27425 2848 27481 2850
rect 28031 2902 28087 2904
rect 28031 2850 28033 2902
rect 28033 2850 28085 2902
rect 28085 2850 28087 2902
rect 28031 2848 28087 2850
rect 28637 2902 28693 2904
rect 28637 2850 28639 2902
rect 28639 2850 28691 2902
rect 28691 2850 28693 2902
rect 28637 2848 28693 2850
rect 18815 1816 18871 1818
rect 18815 1764 18816 1816
rect 18816 1764 18868 1816
rect 18868 1764 18871 1816
rect 18815 1762 18871 1764
rect 19421 1815 19477 1817
rect 19421 1763 19422 1815
rect 19422 1763 19474 1815
rect 19474 1763 19477 1815
rect 19421 1761 19477 1763
rect 20027 1815 20083 1817
rect 20027 1763 20029 1815
rect 20029 1763 20081 1815
rect 20081 1763 20083 1815
rect 20027 1761 20083 1763
rect 29243 1814 29299 1816
rect 29243 1762 29245 1814
rect 29245 1762 29297 1814
rect 29297 1762 29299 1814
rect 29243 1760 29299 1762
rect 29849 1814 29905 1816
rect 29849 1762 29851 1814
rect 29851 1762 29903 1814
rect 29903 1762 29905 1814
rect 29849 1760 29905 1762
rect 30455 1813 30511 1815
rect 30455 1761 30457 1813
rect 30457 1761 30509 1813
rect 30509 1761 30511 1813
rect 30455 1759 30511 1761
rect 31061 1814 31117 1816
rect 31061 1762 31063 1814
rect 31063 1762 31115 1814
rect 31115 1762 31117 1814
rect 31061 1760 31117 1762
rect 31667 1814 31723 1816
rect 31667 1762 31669 1814
rect 31669 1762 31721 1814
rect 31721 1762 31723 1814
rect 31667 1760 31723 1762
rect 32273 1814 32329 1816
rect 32273 1762 32275 1814
rect 32275 1762 32327 1814
rect 32327 1762 32329 1814
rect 32273 1760 32329 1762
rect 32879 1814 32935 1816
rect 32879 1762 32881 1814
rect 32881 1762 32933 1814
rect 32933 1762 32935 1814
rect 32879 1760 32935 1762
rect 33485 1814 33541 1816
rect 33485 1762 33487 1814
rect 33487 1762 33539 1814
rect 33539 1762 33541 1814
rect 33485 1760 33541 1762
rect 34091 1814 34147 1816
rect 34091 1762 34093 1814
rect 34093 1762 34145 1814
rect 34145 1762 34147 1814
rect 34091 1760 34147 1762
rect 34697 1814 34753 1816
rect 34697 1762 34699 1814
rect 34699 1762 34751 1814
rect 34751 1762 34753 1814
rect 34697 1760 34753 1762
rect 39094 5682 39150 5738
rect 35303 1814 35359 1816
rect 35303 1762 35305 1814
rect 35305 1762 35357 1814
rect 35357 1762 35359 1814
rect 35303 1760 35359 1762
rect 35909 1813 35965 1815
rect 35909 1761 35911 1813
rect 35911 1761 35963 1813
rect 35963 1761 35965 1813
rect 35909 1759 35965 1761
rect 36515 1814 36571 1816
rect 36515 1762 36517 1814
rect 36517 1762 36569 1814
rect 36569 1762 36571 1814
rect 36515 1760 36571 1762
rect 37121 1814 37177 1816
rect 37121 1762 37123 1814
rect 37123 1762 37175 1814
rect 37175 1762 37177 1814
rect 37121 1760 37177 1762
rect 37727 1814 37783 1816
rect 37727 1762 37729 1814
rect 37729 1762 37781 1814
rect 37781 1762 37783 1814
rect 37727 1760 37783 1762
rect 966 1669 1022 1671
rect 966 1617 968 1669
rect 968 1617 1020 1669
rect 1020 1617 1022 1669
rect 966 1615 1022 1617
<< metal3 >>
rect 38516 6075 38613 6095
rect 38516 6011 38525 6075
rect 38589 6011 38613 6075
rect 38516 5991 38613 6011
rect 37836 5748 37933 5768
rect 37836 5684 37845 5748
rect 37909 5684 37933 5748
rect 37836 5664 37933 5684
rect 39081 5742 39178 5762
rect 39081 5678 39090 5742
rect 39154 5678 39178 5742
rect 39081 5658 39178 5678
rect 150 4072 210 4087
rect 150 4016 152 4072
rect 208 4016 210 4072
rect 150 4007 210 4016
rect 5094 3927 5175 3932
rect 5094 3871 5106 3927
rect 5162 3871 5175 3927
rect 5094 3866 5175 3871
rect 28632 3102 28633 3192
rect 31725 3183 31726 3192
rect 31663 3179 31726 3183
rect 31721 3168 31726 3179
rect 28697 3152 28698 3168
rect 31721 3123 31726 3152
rect 31663 3122 31670 3123
rect 31671 3122 31726 3123
rect 31663 3102 31726 3122
rect 355 3087 421 3097
rect 355 3031 360 3087
rect 416 3031 421 3087
rect 355 3009 421 3031
rect 358 2929 418 2931
rect 355 2916 421 2929
rect 355 2860 360 2916
rect 416 2860 421 2916
rect 355 2840 421 2860
rect 1267 2916 1333 2925
rect 1267 2860 1272 2916
rect 1328 2860 1333 2916
rect 1267 2850 1333 2860
rect 1873 2915 1939 2924
rect 1873 2859 1878 2915
rect 1934 2859 1939 2915
rect 1268 2845 1332 2850
rect 1873 2840 1939 2859
rect 2804 2914 2864 2918
rect 2804 2858 2806 2914
rect 2862 2858 2864 2914
rect 2804 2852 2864 2858
rect 4013 2916 4079 2929
rect 4013 2860 4018 2916
rect 4074 2860 4079 2916
rect 2866 2840 2867 2841
rect 4013 2839 4079 2860
rect 5352 2909 5367 2930
rect 5401 2909 5418 2930
rect 5352 2853 5357 2909
rect 5413 2853 5418 2909
rect 5352 2840 5418 2853
rect 5958 2907 6024 2916
rect 5958 2851 5963 2907
rect 6019 2851 6024 2907
rect 5958 2839 6024 2851
rect 6564 2907 6630 2916
rect 6564 2851 6569 2907
rect 6625 2851 6630 2907
rect 6564 2838 6630 2851
rect 7170 2907 7236 2916
rect 7170 2851 7175 2907
rect 7231 2851 7236 2907
rect 7170 2838 7236 2851
rect 7776 2907 7842 2916
rect 7776 2851 7781 2907
rect 7837 2851 7842 2907
rect 10932 2903 10998 2912
rect 7776 2838 7842 2851
rect 10327 2842 10391 2852
rect 10932 2847 10937 2903
rect 10993 2847 10998 2903
rect 10932 2838 10998 2847
rect 11538 2904 11604 2913
rect 11538 2848 11543 2904
rect 11599 2848 11604 2904
rect 11538 2839 11604 2848
rect 12144 2903 12210 2912
rect 12144 2847 12149 2903
rect 12205 2847 12210 2903
rect 12144 2838 12210 2847
rect 12750 2903 12816 2912
rect 12750 2847 12755 2903
rect 12811 2847 12816 2903
rect 12750 2838 12816 2847
rect 13356 2905 13422 2914
rect 13356 2849 13361 2905
rect 13417 2849 13422 2905
rect 13356 2840 13422 2849
rect 13962 2905 14028 2914
rect 13962 2849 13967 2905
rect 14023 2849 14028 2905
rect 13962 2840 14028 2849
rect 14568 2904 14634 2913
rect 14568 2848 14573 2904
rect 14629 2848 14634 2904
rect 14568 2839 14634 2848
rect 20148 2904 20214 2917
rect 20148 2848 20153 2904
rect 20209 2848 20214 2904
rect 20148 2838 20214 2848
rect 20754 2904 20820 2917
rect 20754 2848 20759 2904
rect 20815 2848 20820 2904
rect 20754 2838 20820 2848
rect 21360 2905 21426 2918
rect 21360 2849 21365 2905
rect 21421 2849 21426 2905
rect 21360 2839 21426 2849
rect 21966 2904 22032 2917
rect 21966 2848 21971 2904
rect 22027 2848 22032 2904
rect 21966 2838 22032 2848
rect 22572 2904 22638 2917
rect 22572 2848 22577 2904
rect 22633 2848 22638 2904
rect 22572 2838 22638 2848
rect 23178 2904 23244 2917
rect 23178 2848 23183 2904
rect 23239 2848 23244 2904
rect 23178 2838 23244 2848
rect 23784 2904 23850 2917
rect 23784 2848 23789 2904
rect 23845 2848 23850 2904
rect 23784 2838 23850 2848
rect 24390 2904 24456 2917
rect 24390 2848 24395 2904
rect 24451 2848 24456 2904
rect 24390 2838 24456 2848
rect 24996 2904 25062 2917
rect 24996 2848 25001 2904
rect 25057 2848 25062 2904
rect 24996 2838 25062 2848
rect 25602 2904 25668 2917
rect 25602 2848 25607 2904
rect 25663 2848 25668 2904
rect 25602 2838 25668 2848
rect 26208 2904 26274 2917
rect 26208 2848 26213 2904
rect 26269 2848 26274 2904
rect 26208 2838 26274 2848
rect 26814 2904 26880 2917
rect 26814 2848 26819 2904
rect 26875 2848 26880 2904
rect 26814 2838 26880 2848
rect 27420 2904 27486 2917
rect 27420 2848 27425 2904
rect 27481 2848 27486 2904
rect 27420 2838 27486 2848
rect 28026 2904 28092 2917
rect 28026 2848 28031 2904
rect 28087 2848 28092 2904
rect 28026 2838 28092 2848
rect 28633 2893 28635 2908
rect 28633 2882 28637 2893
rect 28633 2881 28636 2882
rect 28633 2877 28637 2881
rect 28633 2839 28635 2877
rect 28693 2883 28697 2893
rect 28694 2882 28697 2883
rect 28693 2877 28697 2882
rect 2442 1894 2545 1904
rect 964 1821 1024 1832
rect 2482 1830 2542 1832
rect 1873 1820 1939 1829
rect 964 1752 1024 1757
rect 1873 1756 1874 1820
rect 1938 1756 1939 1820
rect 1873 1739 1939 1756
rect 2479 1821 2545 1830
rect 2479 1757 2480 1821
rect 2544 1757 2545 1821
rect 2479 1740 2545 1757
rect 3407 1806 3473 1827
rect 3407 1750 3412 1806
rect 3468 1750 3473 1806
rect 3407 1738 3473 1750
rect 4620 1812 4685 1828
rect 4620 1748 4621 1812
rect 5225 1807 5291 1829
rect 5225 1751 5230 1807
rect 5286 1751 5291 1807
rect 7776 1820 7842 1829
rect 7776 1764 7781 1820
rect 7837 1764 7842 1820
rect 7776 1755 7842 1764
rect 8382 1820 8448 1829
rect 8382 1764 8387 1820
rect 8443 1764 8448 1820
rect 8382 1755 8448 1764
rect 8988 1820 9054 1829
rect 8988 1764 8993 1820
rect 9049 1764 9054 1820
rect 8988 1755 9054 1764
rect 9594 1820 9660 1829
rect 9594 1764 9599 1820
rect 9655 1764 9660 1820
rect 15780 1820 15846 1829
rect 9594 1755 9660 1764
rect 10200 1809 10266 1818
rect 4620 1733 4685 1748
rect 5225 1739 5291 1751
rect 10200 1753 10205 1809
rect 10261 1753 10266 1809
rect 15780 1764 15785 1820
rect 15841 1764 15846 1820
rect 15780 1755 15846 1764
rect 16386 1819 16452 1828
rect 16386 1763 16391 1819
rect 16447 1763 16452 1819
rect 16386 1754 16452 1763
rect 16992 1819 17058 1828
rect 16992 1763 16997 1819
rect 17053 1763 17058 1819
rect 16992 1754 17058 1763
rect 17598 1818 17664 1827
rect 17598 1762 17603 1818
rect 17659 1762 17664 1818
rect 17598 1753 17664 1762
rect 18204 1818 18270 1827
rect 18204 1762 18209 1818
rect 18265 1762 18270 1818
rect 18204 1753 18270 1762
rect 18810 1818 18876 1827
rect 18810 1762 18815 1818
rect 18871 1762 18876 1818
rect 18810 1753 18876 1762
rect 19416 1817 19482 1826
rect 19416 1761 19421 1817
rect 19477 1761 19482 1817
rect 10200 1744 10266 1753
rect 19416 1752 19482 1761
rect 20022 1821 20088 1826
rect 20022 1757 20023 1821
rect 20087 1757 20088 1821
rect 29844 1816 29910 1829
rect 29844 1760 29849 1816
rect 29905 1760 29910 1816
rect 20022 1740 20088 1757
rect 29844 1742 29910 1760
rect 30450 1815 30516 1828
rect 30450 1759 30455 1815
rect 30511 1759 30516 1815
rect 30450 1741 30516 1759
rect 31056 1816 31122 1829
rect 31056 1760 31061 1816
rect 31117 1760 31122 1816
rect 31056 1742 31122 1760
rect 31662 1816 31728 1829
rect 31662 1760 31667 1816
rect 31723 1760 31728 1816
rect 31662 1742 31728 1760
rect 32268 1816 32334 1829
rect 32268 1760 32273 1816
rect 32329 1760 32334 1816
rect 32268 1742 32334 1760
rect 32874 1816 32940 1829
rect 32874 1760 32879 1816
rect 32935 1760 32940 1816
rect 32874 1742 32940 1760
rect 33480 1816 33546 1829
rect 33480 1760 33485 1816
rect 33541 1760 33546 1816
rect 33480 1742 33546 1760
rect 34086 1816 34152 1829
rect 34086 1760 34091 1816
rect 34147 1760 34152 1816
rect 34086 1742 34152 1760
rect 34692 1816 34758 1829
rect 34692 1760 34697 1816
rect 34753 1760 34758 1816
rect 34692 1742 34758 1760
rect 35298 1816 35364 1829
rect 35298 1760 35303 1816
rect 35359 1760 35364 1816
rect 35298 1742 35364 1760
rect 35904 1815 35970 1828
rect 35904 1759 35909 1815
rect 35965 1759 35970 1815
rect 35904 1741 35970 1759
rect 36510 1816 36576 1829
rect 36510 1760 36515 1816
rect 36571 1760 36576 1816
rect 36510 1742 36576 1760
rect 37116 1816 37182 1829
rect 37116 1760 37121 1816
rect 37177 1760 37182 1816
rect 37116 1742 37182 1760
rect 37722 1816 37788 1829
rect 37722 1760 37727 1816
rect 37783 1760 37788 1816
rect 37722 1742 37788 1760
rect 961 1671 1027 1682
rect 961 1615 966 1671
rect 1022 1615 1027 1671
rect 961 1596 1027 1615
<< via3 >>
rect 38525 6071 38589 6075
rect 38525 6015 38529 6071
rect 38529 6015 38585 6071
rect 38585 6015 38589 6071
rect 38525 6011 38589 6015
rect 37845 5744 37909 5748
rect 37845 5688 37849 5744
rect 37849 5688 37905 5744
rect 37905 5688 37909 5744
rect 37845 5684 37909 5688
rect 39090 5738 39154 5742
rect 39090 5682 39094 5738
rect 39094 5682 39150 5738
rect 39150 5682 39154 5738
rect 39090 5678 39154 5682
rect 962 1817 1026 1821
rect 962 1761 966 1817
rect 966 1761 1022 1817
rect 1022 1761 1026 1817
rect 962 1757 1026 1761
rect 1874 1816 1938 1820
rect 1874 1760 1878 1816
rect 1878 1760 1934 1816
rect 1934 1760 1938 1816
rect 1874 1756 1938 1760
rect 2480 1817 2544 1821
rect 2480 1761 2484 1817
rect 2484 1761 2540 1817
rect 2540 1761 2544 1817
rect 2480 1757 2544 1761
<< metal4 >>
rect 38511 6075 38950 6291
rect 38065 6013 38298 6014
rect 37836 5748 38298 6013
rect 38511 6011 38525 6075
rect 38589 6011 38950 6075
rect 38511 5806 38950 6011
rect 37836 5684 37845 5748
rect 37909 5684 38298 5748
rect 37836 5449 38298 5684
rect 38065 5448 38298 5449
rect 39077 5742 39565 6049
rect 39077 5678 39090 5742
rect 39154 5678 39565 5742
rect 39077 5415 39565 5678
rect -209 4434 -158 4641
rect 150 3994 210 4087
rect 5094 3866 5175 3932
rect 355 3009 421 3097
rect 355 2840 421 2929
rect 1267 2842 1333 2925
rect 1873 2840 1939 2924
rect 4013 2839 4079 2929
rect 5352 2907 5367 2930
rect 5401 2907 5418 2930
rect 8383 2928 8447 2992
rect 5352 2840 5418 2907
rect 5958 2839 6024 2916
rect 6564 2838 6630 2916
rect 7170 2838 7236 2916
rect 7776 2838 7842 2916
rect 10327 2842 10391 2921
rect 10932 2838 10998 2912
rect 11538 2839 11604 2913
rect 12144 2838 12210 2912
rect 12750 2838 12816 2912
rect 13356 2840 13422 2914
rect 13962 2840 14028 2914
rect 14568 2839 14634 2913
rect 20148 2838 20214 2917
rect 20754 2838 20820 2917
rect 21360 2839 21426 2918
rect 21966 2838 22032 2917
rect 22572 2838 22638 2917
rect 23178 2838 23244 2917
rect 23784 2838 23850 2917
rect 24390 2838 24456 2917
rect 24996 2838 25062 2917
rect 25602 2838 25668 2917
rect 26208 2838 26274 2917
rect 26814 2838 26880 2917
rect 27420 2838 27486 2917
rect 28026 2838 28092 2917
rect -93 1882 -33 1897
rect 964 1821 1024 1830
rect 1873 1820 1939 1829
rect 964 1740 1024 1757
rect 1873 1756 1874 1820
rect 1938 1756 1939 1820
rect 1873 1739 1939 1756
rect 2479 1821 2545 1830
rect 2479 1757 2480 1821
rect 2544 1757 2545 1821
rect 2479 1740 2545 1757
rect 3407 1738 3473 1827
rect 4620 1812 4685 1828
rect 4620 1748 4621 1812
rect 4620 1733 4685 1748
rect 5225 1739 5291 1829
rect 7776 1755 7842 1829
rect 8382 1755 8448 1829
rect 8988 1755 9054 1829
rect 9594 1755 9660 1829
rect 10200 1744 10266 1818
rect 15780 1755 15846 1829
rect 16386 1754 16452 1828
rect 16992 1754 17058 1828
rect 17598 1753 17664 1827
rect 18204 1753 18270 1827
rect 18810 1753 18876 1827
rect 19416 1752 19482 1826
rect 20023 1821 20087 1825
rect 29238 1739 29304 1829
rect 29844 1742 29910 1829
rect 30450 1741 30516 1828
rect 31056 1742 31122 1829
rect 31662 1742 31728 1829
rect 32268 1742 32334 1829
rect 32874 1742 32940 1829
rect 33480 1742 33546 1829
rect 34086 1742 34152 1829
rect 34692 1742 34758 1829
rect 35298 1742 35364 1829
rect 35904 1741 35970 1828
rect 36510 1742 36576 1829
rect 37116 1742 37182 1829
rect 37722 1742 37788 1829
rect 961 1596 1027 1682
rect -205 1413 -161 1543
<< metal5 >>
rect 245 4094 565 5026
rect 1675 4100 1995 5026
rect 3259 4132 3579 5026
rect 5352 4142 5672 5026
rect 10326 4154 10646 5026
rect 39256 4154 39576 5026
rect 287 -595 524 -359
rect 1717 -595 1954 -359
rect 3301 -595 3538 -359
rect 5394 -595 5631 -359
rect 10368 -595 10605 -359
rect 39298 -595 39534 -359
use hgu_cdac_8bit_array  hgu_cdac_8bit_array_2
timestamp 1700813856
transform 1 0 4202 0 -1 -5445
box -4661 -7612 35404 -4800
use hgu_cdac_8bit_array  hgu_cdac_8bit_array_3
timestamp 1700813856
transform 1 0 4202 0 -1 -2312
box -4661 -7612 35404 -4800
use hgu_cdac_unit  hgu_cdac_unit_0
timestamp 1700813856
transform 1 0 -1145 0 -1 1399
box 686 598 1358 1826
use hgu_cdac_unit  hgu_cdac_unit_1
timestamp 1700813856
transform 1 0 -1145 0 -1 4532
box 686 598 1358 1826
use hgu_inverter  hgu_inverter_0
timestamp 1700938176
transform 1 0 -747 0 1 4944
box 347 160 675 824
use hgu_inverter  hgu_inverter_1
timestamp 1700938176
transform 1 0 -747 0 -1 6474
box 347 160 675 824
use inv_2_test  inv_2_test_0
timestamp 1700938176
transform 1 0 128 0 1 2744
box 400 2360 856 3024
use inv_2_test  inv_2_test_1
timestamp 1700938176
transform -1 0 1256 0 -1 8674
box 400 2360 856 3024
use inv_4_test  inv_4_test_1
timestamp 1700938176
transform 1 0 2239 0 1 3780
box -447 1324 265 1988
use inv_4_test  inv_4_test_2
timestamp 1700938176
transform -1 0 1545 0 -1 7638
box -447 1324 265 1988
use inv_8_test  inv_8_test_0
timestamp 1700938176
transform 1 0 3315 0 1 2784
box 96 2320 1320 2984
use inv_8_test  inv_8_test_1
timestamp 1700938176
transform -1 0 4219 0 -1 8634
box 96 2320 1320 2984
use inv_16_test  inv_16_test_0
timestamp 1700938176
transform 1 0 8625 0 1 5144
box -649 -40 1599 624
use inv_16_test  inv_16_test_1
timestamp 1700938176
transform -1 0 6991 0 -1 6274
box -649 -40 1599 624
use inv_32_test  inv_32_test_0
timestamp 1700938176
transform -1 0 12472 0 -1 3912
box -2303 -2402 1993 -1738
use inv_32_test  inv_32_test_1
timestamp 1700938176
transform 1 0 18043 0 1 7506
box -2303 -2402 1993 -1738
use inv_64_test  inv_64_test_0
timestamp 1700938176
transform 1 0 32867 0 1 7506
box -3583 -2402 4809 -1738
use inv_64_test  inv_64_test_1
timestamp 1700938176
transform -1 0 25125 0 -1 3912
box -3583 -2402 4809 -1738
<< labels >>
flabel metal4 -209 4434 -158 4641 0 FreeSans 480 0 0 0 t<0>
port 27 nsew
flabel poly 10608 6023 14646 6093 0 FreeSans 320 0 0 0 d<5>
port 113 nsew
flabel poly -271 5290 -201 5422 0 FreeSans 320 0 0 0 db<0>
port 117 nsew
flabel poly 657 5290 727 5422 0 FreeSans 320 0 0 0 db<1>
port 119 nsew
flabel poly 1921 5335 2375 5405 0 FreeSans 320 0 0 0 db<2>
port 121 nsew
flabel poly 3540 5335 4506 5405 0 FreeSans 320 0 0 0 db<3>
port 123 nsew
flabel metal5 245 4094 565 5026 0 FreeSans 800 0 0 0 t<1>
port 166 nsew
flabel metal5 1675 4100 1995 5026 0 FreeSans 800 0 0 0 t<2>
port 168 nsew
flabel metal5 3259 4132 3579 5026 0 FreeSans 800 0 0 0 t<3>
port 170 nsew
flabel metal5 5352 4142 5672 5026 0 FreeSans 800 0 0 0 t<4>
port 172 nsew
flabel metal5 39256 4154 39576 5026 0 FreeSans 800 0 0 0 t<6>
port 178 nsew
flabel metal4 -205 1413 -161 1543 0 FreeSans 320 0 0 0 tb<0>
port 76 nsew
flabel metal5 287 -595 524 -359 0 FreeSans 480 0 0 0 tb<1>
port 147 nsew
flabel metal5 1717 -595 1954 -359 0 FreeSans 480 0 0 0 tb<2>
port 149 nsew
flabel metal5 3301 -595 3538 -359 0 FreeSans 480 0 0 0 tb<3>
port 151 nsew
flabel metal5 5394 -595 5631 -359 0 FreeSans 480 0 0 0 tb<4>
port 153 nsew
flabel metal5 10368 -595 10605 -359 0 FreeSans 480 0 0 0 tb<5>
port 155 nsew
flabel metal5 39298 -595 39534 -359 0 FreeSans 480 0 0 0 tb<6>
port 157 nsew
flabel poly 657 5978 727 6110 0 FreeSans 320 0 0 0 d<1>
port 106 nsew
flabel poly 1409 6013 1863 6083 0 FreeSans 320 0 0 0 d<2>
port 104 nsew
flabel poly 3028 6013 3994 6083 0 FreeSans 320 0 0 0 d<3>
port 102 nsew
flabel metal5 10326 4154 10646 5026 0 FreeSans 800 0 0 0 t<5>
port 176 nsew
flabel poly 20445 6013 28579 6083 0 FreeSans 1600 0 0 0 d<6>
port 180 nsew
flabel poly 29413 5335 37547 5405 0 FreeSans 1600 0 0 0 db<6>
port 182 nsew
flabel poly 15869 5335 19907 5405 0 FreeSans 480 0 0 0 db<5>
port 184 nsew
flabel poly -271 5997 -201 6129 0 FreeSans 320 0 0 0 d<0>
port 109 nsew
flabel metal4 39154 5415 39565 6049 0 FreeSans 1600 0 0 0 VDD
port 161 nsew
flabel metal4 37909 5449 38298 6013 0 FreeSans 1600 0 0 0 VREF
port 163 nsew
flabel metal4 38589 5806 38950 6291 0 FreeSans 1600 0 0 0 VSS
port 159 nsew
flabel poly 5521 6013 7511 6083 0 FreeSans 480 0 0 0 d<4>
port 186 nsew
flabel poly 8105 5335 10095 5405 0 FreeSans 480 0 0 0 db<4>
port 188 nsew
<< end >>
