magic
tech sky130A
magscale 1 2
timestamp 1697616495
<< nmos >>
rect -369 -42 369 42
<< ndiff >>
rect -427 30 -369 42
rect -427 -30 -415 30
rect -381 -30 -369 30
rect -427 -42 -369 -30
rect 369 30 427 42
rect 369 -30 381 30
rect 415 -30 427 30
rect 369 -42 427 -30
<< ndiffc >>
rect -415 -30 -381 30
rect 381 -30 415 30
<< poly >>
rect -369 114 369 130
rect -369 80 -353 114
rect 353 80 369 114
rect -369 42 369 80
rect -369 -80 369 -42
rect -369 -114 -353 -80
rect 353 -114 369 -80
rect -369 -130 369 -114
<< polycont >>
rect -353 80 353 114
rect -353 -114 353 -80
<< locali >>
rect -369 80 -353 114
rect 353 80 369 114
rect -415 30 -381 46
rect -415 -46 -381 -30
rect 381 30 415 46
rect 381 -46 415 -30
rect -369 -114 -353 -80
rect 353 -114 369 -80
<< viali >>
rect -353 80 353 114
rect -415 -30 -381 30
rect 381 -30 415 30
rect -353 -114 353 -80
<< metal1 >>
rect -365 114 365 120
rect -365 80 -353 114
rect 353 80 365 114
rect -365 74 365 80
rect -421 30 -375 42
rect -421 -30 -415 30
rect -381 -30 -375 30
rect -421 -42 -375 -30
rect 375 30 421 42
rect 375 -30 381 30
rect 415 -30 421 30
rect 375 -42 421 -30
rect -365 -80 365 -74
rect -365 -114 -353 -80
rect 353 -114 365 -80
rect -365 -120 365 -114
<< properties >>
string FIXED_BBOX -512 -199 512 199
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.42 l 3.69 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
