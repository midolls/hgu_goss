magic
tech sky130A
magscale 1 2
timestamp 1700649561
<< nwell >>
rect -98 1976 408 2272
rect -98 1808 413 1976
rect -98 1296 408 1808
rect 47 1259 267 1296
<< pwell >>
rect -176 -206 498 1048
<< nmos >>
rect 88 992 118 1076
rect 160 992 190 1076
rect 88 854 118 938
rect 160 854 190 938
rect 88 716 118 800
rect 160 716 190 800
rect 88 578 118 662
rect 160 578 190 662
rect 88 440 118 524
rect 160 440 190 524
rect 88 302 118 386
rect 160 302 190 386
rect 88 164 118 248
rect 160 164 190 248
rect 88 26 118 110
rect 160 26 190 110
<< pmoshvt >>
rect 142 1997 172 2081
rect 142 1859 172 1943
rect 142 1721 172 1805
rect 142 1583 172 1667
rect 142 1445 172 1529
rect 142 1307 172 1391
<< ndiff >>
rect 30 1064 88 1076
rect 30 1004 42 1064
rect 76 1004 88 1064
rect 30 992 88 1004
rect 118 992 160 1076
rect 190 1064 248 1076
rect 190 1004 202 1064
rect 236 1004 248 1064
rect 190 992 248 1004
rect 30 926 88 938
rect 30 866 42 926
rect 76 866 88 926
rect 30 854 88 866
rect 118 854 160 938
rect 190 926 248 938
rect 190 866 202 926
rect 236 866 248 926
rect 190 854 248 866
rect 30 788 88 800
rect 30 728 42 788
rect 76 728 88 788
rect 30 716 88 728
rect 118 716 160 800
rect 190 788 248 800
rect 190 728 202 788
rect 236 728 248 788
rect 190 716 248 728
rect 30 650 88 662
rect 30 590 42 650
rect 76 590 88 650
rect 30 578 88 590
rect 118 578 160 662
rect 190 650 248 662
rect 190 590 202 650
rect 236 590 248 650
rect 190 578 248 590
rect 30 512 88 524
rect 30 452 42 512
rect 76 452 88 512
rect 30 440 88 452
rect 118 440 160 524
rect 190 512 248 524
rect 190 452 202 512
rect 236 452 248 512
rect 190 440 248 452
rect 30 374 88 386
rect 30 314 42 374
rect 76 314 88 374
rect 30 302 88 314
rect 118 302 160 386
rect 190 374 248 386
rect 190 314 202 374
rect 236 314 248 374
rect 190 302 248 314
rect 30 236 88 248
rect 30 176 42 236
rect 76 176 88 236
rect 30 164 88 176
rect 118 164 160 248
rect 190 236 248 248
rect 190 176 202 236
rect 236 176 248 236
rect 190 164 248 176
rect 30 98 88 110
rect 30 38 42 98
rect 76 38 88 98
rect 30 26 88 38
rect 118 26 160 110
rect 190 98 248 110
rect 190 38 202 98
rect 236 38 248 98
rect 190 26 248 38
<< pdiff >>
rect 84 2069 142 2081
rect 84 2009 96 2069
rect 130 2009 142 2069
rect 84 1997 142 2009
rect 172 2069 230 2081
rect 172 2009 184 2069
rect 218 2009 230 2069
rect 172 1997 230 2009
rect 84 1931 142 1943
rect 84 1871 96 1931
rect 130 1871 142 1931
rect 84 1859 142 1871
rect 172 1931 230 1943
rect 172 1871 184 1931
rect 218 1871 230 1931
rect 172 1859 230 1871
rect 84 1793 142 1805
rect 84 1733 96 1793
rect 130 1733 142 1793
rect 84 1721 142 1733
rect 172 1793 230 1805
rect 172 1733 184 1793
rect 218 1733 230 1793
rect 172 1721 230 1733
rect 84 1655 142 1667
rect 84 1595 96 1655
rect 130 1595 142 1655
rect 84 1583 142 1595
rect 172 1655 230 1667
rect 172 1595 184 1655
rect 218 1595 230 1655
rect 172 1583 230 1595
rect 84 1517 142 1529
rect 84 1457 96 1517
rect 130 1457 142 1517
rect 84 1445 142 1457
rect 172 1517 230 1529
rect 172 1457 184 1517
rect 218 1457 230 1517
rect 172 1445 230 1457
rect 84 1379 142 1391
rect 84 1319 96 1379
rect 130 1319 142 1379
rect 84 1307 142 1319
rect 172 1379 230 1391
rect 172 1319 184 1379
rect 218 1319 230 1379
rect 172 1307 230 1319
<< ndiffc >>
rect 42 1004 76 1064
rect 202 1004 236 1064
rect 42 866 76 926
rect 202 866 236 926
rect 42 728 76 788
rect 202 728 236 788
rect 42 590 76 650
rect 202 590 236 650
rect 42 452 76 512
rect 202 452 236 512
rect 42 314 76 374
rect 202 314 236 374
rect 42 176 76 236
rect 202 176 236 236
rect 42 38 76 98
rect 202 38 236 98
<< pdiffc >>
rect 96 2009 130 2069
rect 184 2009 218 2069
rect 96 1871 130 1931
rect 184 1871 218 1931
rect 96 1733 130 1793
rect 184 1733 218 1793
rect 96 1595 130 1655
rect 184 1595 218 1655
rect 96 1457 130 1517
rect 184 1457 218 1517
rect 96 1319 130 1379
rect 184 1319 218 1379
<< psubdiff >>
rect -135 944 -31 979
rect -135 910 -104 944
rect -70 910 -31 944
rect -135 882 -31 910
rect 329 876 433 911
rect 329 842 360 876
rect 394 842 433 876
rect 329 814 433 842
rect -151 738 -47 773
rect -151 704 -120 738
rect -86 704 -47 738
rect 321 724 425 759
rect -151 676 -47 704
rect 321 690 352 724
rect 386 690 425 724
rect 321 662 425 690
rect -147 546 -43 581
rect -147 512 -116 546
rect -82 512 -43 546
rect 329 534 433 569
rect -147 484 -43 512
rect 329 500 360 534
rect 394 500 433 534
rect 329 472 433 500
rect -129 390 -25 425
rect -129 356 -98 390
rect -64 356 -25 390
rect -129 328 -25 356
rect 345 382 449 417
rect 345 348 376 382
rect 410 348 449 382
rect 345 320 449 348
rect -131 236 -27 271
rect -131 202 -100 236
rect -66 202 -27 236
rect -131 174 -27 202
rect 319 222 423 257
rect 319 188 350 222
rect 384 188 423 222
rect 319 159 423 188
rect -133 60 -29 95
rect -133 26 -102 60
rect -68 26 -29 60
rect 333 46 437 81
rect -133 -2 -29 26
rect 333 12 364 46
rect 398 12 437 46
rect 333 -16 437 12
rect -115 -104 -11 -69
rect -115 -138 -84 -104
rect -50 -138 -11 -104
rect -115 -166 -11 -138
rect 111 -104 215 -69
rect 111 -138 142 -104
rect 176 -138 215 -104
rect 111 -166 215 -138
rect 323 -110 427 -75
rect 323 -144 354 -110
rect 388 -144 427 -110
rect 323 -172 427 -144
<< nsubdiff >>
rect 276 2203 359 2228
rect 276 2168 301 2203
rect 335 2168 359 2203
rect -60 2139 23 2164
rect 276 2144 359 2168
rect -60 2104 -35 2139
rect -1 2104 23 2139
rect -60 2080 23 2104
rect -54 1983 29 2008
rect 288 2065 371 2090
rect 288 2030 313 2065
rect 347 2030 371 2065
rect 288 2006 371 2030
rect -54 1948 -29 1983
rect 5 1948 29 1983
rect -54 1924 29 1948
rect 284 1915 367 1940
rect 284 1880 309 1915
rect 343 1880 367 1915
rect -54 1799 29 1824
rect 284 1856 367 1880
rect -54 1764 -29 1799
rect 5 1764 29 1799
rect -54 1740 29 1764
rect 284 1769 367 1794
rect 284 1734 309 1769
rect 343 1734 367 1769
rect -58 1653 25 1678
rect 284 1710 367 1734
rect -58 1618 -33 1653
rect 1 1618 25 1653
rect -58 1594 25 1618
rect 286 1623 369 1648
rect 286 1588 311 1623
rect 345 1588 369 1623
rect 286 1564 369 1588
rect -54 1471 29 1496
rect -54 1436 -29 1471
rect 5 1436 29 1471
rect 286 1471 369 1496
rect -54 1412 29 1436
rect 286 1436 311 1471
rect 345 1436 369 1471
rect 286 1412 369 1436
<< psubdiffcont >>
rect -104 910 -70 944
rect 360 842 394 876
rect -120 704 -86 738
rect 352 690 386 724
rect -116 512 -82 546
rect 360 500 394 534
rect -98 356 -64 390
rect 376 348 410 382
rect -100 202 -66 236
rect 350 188 384 222
rect -102 26 -68 60
rect 364 12 398 46
rect -84 -138 -50 -104
rect 142 -138 176 -104
rect 354 -144 388 -110
<< nsubdiffcont >>
rect 301 2168 335 2203
rect -35 2104 -1 2139
rect 313 2030 347 2065
rect -29 1948 5 1983
rect 309 1880 343 1915
rect -29 1764 5 1799
rect 309 1734 343 1769
rect -33 1618 1 1653
rect 311 1588 345 1623
rect -29 1436 5 1471
rect 311 1436 345 1471
<< poly >>
rect 142 2081 172 2111
rect 142 1943 172 1997
rect 142 1805 172 1859
rect 142 1667 172 1721
rect 142 1529 172 1583
rect 142 1391 172 1445
rect 142 1276 172 1307
rect 124 1260 190 1276
rect 124 1226 140 1260
rect 174 1226 190 1260
rect 124 1121 190 1226
rect 88 1091 190 1121
rect 88 1076 118 1091
rect 160 1076 190 1091
rect 88 938 118 992
rect 160 938 190 992
rect 88 800 118 854
rect 160 800 190 854
rect 88 662 118 716
rect 160 662 190 716
rect 88 524 118 578
rect 160 524 190 578
rect 88 386 118 440
rect 160 386 190 440
rect 88 248 118 302
rect 160 248 190 302
rect 88 110 118 164
rect 160 110 190 164
rect 88 0 118 26
rect 160 0 190 26
<< polycont >>
rect 140 1226 174 1260
<< locali >>
rect -18 2256 32 2258
rect 298 2256 348 2258
rect -18 2248 356 2256
rect -18 2228 358 2248
rect -18 2210 359 2228
rect -18 2164 32 2210
rect -60 2139 32 2164
rect 276 2203 359 2210
rect 276 2168 301 2203
rect 335 2168 359 2203
rect 276 2144 359 2168
rect -60 2104 -35 2139
rect -1 2104 32 2139
rect -60 2080 32 2104
rect 292 2090 358 2144
rect -18 2008 32 2080
rect 96 2069 130 2085
rect -54 1983 29 2008
rect -54 1948 -29 1983
rect 5 1948 29 1983
rect -54 1924 29 1948
rect 96 1931 130 2009
rect 184 2075 218 2085
rect 288 2076 371 2090
rect 253 2075 371 2076
rect 184 2069 371 2075
rect 218 2065 371 2069
rect 218 2030 313 2065
rect 347 2030 371 2065
rect 218 2009 371 2030
rect 184 2006 371 2009
rect 184 2004 354 2006
rect 184 1993 218 2004
rect -18 1824 32 1924
rect 96 1855 130 1871
rect 184 1931 218 1947
rect 297 1940 354 2004
rect -54 1799 29 1824
rect -54 1764 -29 1799
rect 5 1764 29 1799
rect -54 1740 29 1764
rect 96 1793 130 1809
rect -18 1678 32 1740
rect -58 1653 32 1678
rect -58 1618 -33 1653
rect 1 1618 32 1653
rect -58 1594 32 1618
rect -18 1496 32 1594
rect 96 1655 130 1733
rect 184 1793 218 1871
rect 284 1915 367 1940
rect 284 1880 309 1915
rect 343 1880 367 1915
rect 284 1856 367 1880
rect 298 1794 348 1856
rect 184 1717 218 1733
rect 284 1769 367 1794
rect 284 1734 309 1769
rect 343 1734 367 1769
rect 284 1710 367 1734
rect 96 1579 130 1595
rect 184 1655 218 1671
rect 298 1648 348 1710
rect -54 1471 32 1496
rect -54 1436 -29 1471
rect 5 1436 32 1471
rect -54 1412 32 1436
rect -18 1302 32 1412
rect 96 1517 130 1533
rect 96 1379 130 1457
rect 184 1517 218 1595
rect 286 1623 369 1648
rect 286 1588 311 1623
rect 345 1588 369 1623
rect 286 1564 369 1588
rect 298 1496 348 1564
rect 184 1441 218 1457
rect 286 1471 369 1496
rect 286 1436 311 1471
rect 345 1436 369 1471
rect 286 1412 369 1436
rect 96 1303 130 1319
rect 184 1379 218 1395
rect 184 1303 218 1319
rect 298 1302 348 1412
rect 124 1226 140 1260
rect 174 1226 190 1260
rect 116 1126 162 1144
rect 116 1092 122 1126
rect 156 1092 162 1126
rect 116 1080 162 1092
rect 42 1064 76 1080
rect -94 980 -44 1062
rect -114 979 -44 980
rect -136 944 -31 979
rect -136 910 -104 944
rect -70 910 -31 944
rect -136 882 -31 910
rect 42 926 76 1004
rect 202 1064 236 1080
rect 202 988 236 1004
rect -94 774 -44 882
rect 42 850 76 866
rect 202 926 236 942
rect 340 912 390 1044
rect 340 911 400 912
rect -130 773 -44 774
rect -152 738 -44 773
rect -152 704 -120 738
rect -86 704 -44 738
rect -152 676 -44 704
rect -94 582 -44 676
rect -126 581 -44 582
rect 42 788 76 804
rect 42 650 76 728
rect 202 788 236 866
rect 328 876 433 911
rect 328 842 360 876
rect 394 842 433 876
rect 328 814 433 842
rect 340 760 390 814
rect 340 759 392 760
rect 202 712 236 728
rect 320 724 425 759
rect 320 690 352 724
rect 386 690 425 724
rect -148 546 -43 581
rect 42 574 76 590
rect 202 650 236 666
rect 320 662 425 690
rect -148 512 -116 546
rect -82 512 -43 546
rect -148 484 -43 512
rect 42 512 76 528
rect -94 426 -44 484
rect -108 425 -44 426
rect -130 390 -25 425
rect -130 356 -98 390
rect -64 356 -25 390
rect -130 328 -25 356
rect 42 374 76 452
rect 202 512 236 590
rect 340 570 390 662
rect 340 569 400 570
rect 328 534 433 569
rect 328 500 360 534
rect 394 500 433 534
rect 328 472 433 500
rect 202 436 236 452
rect 340 418 390 472
rect 340 417 416 418
rect -94 272 -44 328
rect 42 298 76 314
rect 202 374 236 390
rect -110 271 -44 272
rect -132 236 -27 271
rect -132 202 -100 236
rect -66 202 -27 236
rect -132 174 -27 202
rect 42 236 76 252
rect -94 96 -44 174
rect -112 95 -44 96
rect 42 98 76 176
rect 202 236 236 314
rect 340 382 449 417
rect 340 348 376 382
rect 410 348 449 382
rect 340 320 449 348
rect 340 257 390 320
rect 202 160 236 176
rect 318 222 423 257
rect 318 188 350 222
rect 384 188 423 222
rect 318 159 423 188
rect -134 60 -29 95
rect -134 26 -102 60
rect -68 26 -29 60
rect -134 -2 -29 26
rect 42 22 76 38
rect 202 104 236 114
rect 332 104 409 159
rect 202 98 409 104
rect 236 81 409 98
rect 236 46 437 81
rect 236 38 364 46
rect 202 35 364 38
rect 202 22 236 35
rect 324 12 364 35
rect 398 12 437 46
rect -94 -69 -44 -2
rect 324 -16 437 12
rect 132 -69 182 -68
rect -116 -88 -11 -69
rect 110 -88 215 -69
rect 324 -75 410 -16
rect 322 -88 427 -75
rect -116 -104 427 -88
rect -116 -138 -84 -104
rect -50 -132 142 -104
rect -50 -138 -11 -132
rect -116 -166 -11 -138
rect 110 -138 142 -132
rect 176 -110 427 -104
rect 176 -132 354 -110
rect 176 -138 215 -132
rect 110 -166 215 -138
rect 322 -144 354 -132
rect 388 -144 427 -110
rect 322 -172 427 -144
<< viali >>
rect 96 2009 130 2069
rect 184 2009 218 2069
rect 96 1871 130 1931
rect 184 1871 218 1931
rect 96 1733 130 1793
rect 184 1733 218 1793
rect 96 1595 130 1655
rect 184 1595 218 1655
rect 96 1457 130 1517
rect 184 1457 218 1517
rect 96 1319 130 1379
rect 184 1319 218 1379
rect 140 1226 174 1260
rect 122 1092 156 1126
rect 42 1004 76 1064
rect 202 1004 236 1064
rect 42 866 76 926
rect 202 866 236 926
rect 42 728 76 788
rect 202 728 236 788
rect 42 590 76 650
rect 202 590 236 650
rect 42 452 76 512
rect 202 452 236 512
rect 42 314 76 374
rect 202 314 236 374
rect 42 176 76 236
rect 202 176 236 236
rect 42 38 76 98
rect 202 38 236 98
<< metal1 >>
rect 158 2140 252 2190
rect 90 2069 136 2081
rect 90 2009 96 2069
rect 130 2009 136 2069
rect 90 1931 136 2009
rect 178 2069 224 2140
rect 178 2009 184 2069
rect 218 2009 224 2069
rect 178 1997 224 2009
rect 90 1871 96 1931
rect 130 1871 136 1931
rect 90 1859 136 1871
rect 178 1931 224 1943
rect 178 1871 184 1931
rect 218 1871 224 1931
rect 90 1793 136 1805
rect 90 1733 96 1793
rect 130 1733 136 1793
rect 90 1655 136 1733
rect 178 1793 224 1871
rect 178 1733 184 1793
rect 218 1733 224 1793
rect 178 1721 224 1733
rect 90 1595 96 1655
rect 130 1595 136 1655
rect 90 1583 136 1595
rect 178 1655 224 1667
rect 178 1595 184 1655
rect 218 1595 224 1655
rect 90 1517 136 1529
rect 90 1457 96 1517
rect 130 1457 136 1517
rect 90 1379 136 1457
rect 178 1517 224 1595
rect 178 1457 184 1517
rect 218 1457 224 1517
rect 178 1445 224 1457
rect 90 1319 96 1379
rect 130 1319 136 1379
rect 90 1307 136 1319
rect 178 1379 224 1391
rect 178 1319 184 1379
rect 218 1336 224 1379
rect 218 1334 528 1336
rect 218 1319 548 1334
rect 178 1294 548 1319
rect 280 1292 548 1294
rect 128 1260 186 1266
rect 116 1226 140 1260
rect 174 1226 186 1260
rect 116 1220 186 1226
rect -62 1172 -6 1192
rect 116 1172 160 1220
rect 502 1208 548 1292
rect 594 1208 688 1226
rect 502 1174 688 1208
rect -62 1126 186 1172
rect -62 1104 -6 1126
rect 116 1092 122 1126
rect 156 1092 162 1126
rect 502 1096 548 1174
rect 594 1136 688 1174
rect 116 1080 162 1092
rect 36 1064 82 1076
rect 36 1004 42 1064
rect 76 1004 82 1064
rect 36 926 82 1004
rect 196 1064 548 1096
rect 196 1004 202 1064
rect 236 1054 548 1064
rect 236 1052 544 1054
rect 236 1004 242 1052
rect 196 992 242 1004
rect 36 866 42 926
rect 76 866 82 926
rect 36 854 82 866
rect 196 926 242 938
rect 196 866 202 926
rect 236 866 242 926
rect 36 788 82 800
rect 36 728 42 788
rect 76 728 82 788
rect 36 650 82 728
rect 196 788 242 866
rect 196 728 202 788
rect 236 728 242 788
rect 196 716 242 728
rect 36 590 42 650
rect 76 590 82 650
rect 36 578 82 590
rect 196 650 242 662
rect 196 590 202 650
rect 236 590 242 650
rect 36 512 82 524
rect 36 452 42 512
rect 76 452 82 512
rect 36 374 82 452
rect 196 512 242 590
rect 196 452 202 512
rect 236 452 242 512
rect 196 440 242 452
rect 36 314 42 374
rect 76 314 82 374
rect 36 302 82 314
rect 196 374 242 386
rect 196 314 202 374
rect 236 314 242 374
rect 36 236 82 248
rect 36 176 42 236
rect 76 176 82 236
rect 36 98 82 176
rect 196 236 242 314
rect 196 176 202 236
rect 236 176 242 236
rect 196 164 242 176
rect 36 38 42 98
rect 76 38 82 98
rect 36 26 82 38
rect 196 98 242 110
rect 196 38 202 98
rect 236 38 242 98
rect 196 -10 242 38
rect 182 -60 264 -10
<< labels >>
flabel metal1 182 -60 264 -10 0 FreeSans 320 0 0 0 vss
port 1 nsew
flabel metal1 -62 1104 -6 1192 0 FreeSans 320 0 0 0 input
port 2 nsew
flabel metal1 158 2140 252 2190 0 FreeSans 320 0 0 0 vdd
port 0 nsew
flabel metal1 594 1136 688 1226 0 FreeSans 320 0 0 0 output
port 4 nsew
flabel metal1 140 1226 174 1260 0 FreeSans 320 0 0 0 hgu_pfet_hvt_stack_in_delay_0.input_stack
flabel nwell 184 2009 218 2069 0 FreeSans 320 0 0 0 hgu_pfet_hvt_stack_in_delay_0.vdd
flabel metal1 178 1307 224 1319 0 FreeSans 320 0 0 0 hgu_pfet_hvt_stack_in_delay_0.output_stack
flabel poly 88 1091 190 1121 0 FreeSans 320 0 0 0 hgu_nfet_hvt_stack_in_delay_0.input_stack
flabel metal1 202 38 236 98 0 FreeSans 320 0 0 0 hgu_nfet_hvt_stack_in_delay_0.vss
flabel metal1 196 1064 242 1076 0 FreeSans 320 0 0 0 hgu_nfet_hvt_stack_in_delay_0.output_stack
<< end >>
