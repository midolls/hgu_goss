* NGSPICE file created from hgu_comp_flat.ext - technology: sky130A

.subckt hgu_comp_flat cdac_vn cdac_vp comp_outp comp_outn clk VDD VSS
X0 a_1830_n378# cdac_vn a_582_n702# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1 VSS a_476_n1721# a_564_n1266# VSS sky130_fd_pr__nfet_01v8 ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.15
X2 comp_outp a_1950_n1721# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.3 as=0.139 ps=1.17 w=0.84 l=0.15
X3 a_582_n702# cdac_vn a_1830_n378# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X4 a_1950_n1721# RS_p VDD VDD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0.244 ps=2.26 w=0.84 l=0.15
X5 a_482_n1818# a_1716_n1348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0759 pd=0.79 as=0.143 ps=1.54 w=0.46 l=0.15
X6 a_476_n1266# a_482_n1818# a_476_n1721# VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.15
X7 VDD a_1026_n1747# comp_outn VDD sky130_fd_pr__pfet_01v8 ad=0.139 pd=1.17 as=0.26 ps=2.3 w=0.84 l=0.15
X8 VSS RS_n a_1026_n1747# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X9 VDD clk a_1248_n288# VDD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X10 a_674_n702# cdac_vp a_582_n702# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.165 pd=1.33 as=0.31 ps=2.62 w=1 l=0.15
X11 VDD a_852_n296# a_476_n1721# VDD sky130_fd_pr__pfet_01v8 ad=0.139 pd=1.17 as=0.26 ps=2.3 w=0.84 l=0.15
X12 comp_outn a_1026_n1747# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.139 pd=1.17 as=0.139 ps=1.17 w=0.84 l=0.15
X13 a_476_n1721# a_852_n296# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.139 pd=1.17 as=0.139 ps=1.17 w=0.84 l=0.15
X14 a_582_n702# cdac_vn a_1830_n378# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X15 a_582_n702# cdac_vp a_674_n702# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X16 comp_outp a_1950_n1721# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.54 as=0.0759 ps=0.79 w=0.46 l=0.15
X17 VDD a_852_n296# a_476_n1721# VDD sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.3 as=0.139 ps=1.17 w=0.84 l=0.15
X18 a_674_n702# cdac_vp a_582_n702# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X19 a_1830_n378# cdac_vn a_582_n702# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X20 a_564_n1266# a_482_n1818# a_476_n1266# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.15
X21 VSS a_1026_n1747# comp_outn VSS sky130_fd_pr__nfet_01v8 ad=0.0759 pd=0.79 as=0.143 ps=1.54 w=0.46 l=0.15
X22 a_1950_n1721# RS_p VSS VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X23 a_1566_n378# clk VDD VDD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X24 VSS a_852_n296# a_476_n1721# VSS sky130_fd_pr__nfet_01v8 ad=0.0759 pd=0.79 as=0.143 ps=1.54 w=0.46 l=0.15
X25 VDD a_1248_n288# a_852_n296# VDD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0.244 ps=2.26 w=0.84 l=0.15
X26 a_482_n1818# a_1716_n1348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.54 as=0.0759 ps=0.79 w=0.46 l=0.15
X27 a_582_n702# clk VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X28 comp_outn a_1026_n1747# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0759 pd=0.79 as=0.0759 ps=0.79 w=0.46 l=0.15
X29 VSS a_1248_n288# a_852_n296# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X30 a_674_n702# cdac_vp a_582_n702# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X31 a_582_n702# cdac_vn a_1830_n378# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X32 a_1248_n288# a_1566_n378# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X33 a_1918_109# clk VDD VDD sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X34 a_582_n702# cdac_vp a_674_n702# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X35 VDD a_1026_n1747# comp_outn VDD sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.3 as=0.139 ps=1.17 w=0.84 l=0.15
X36 RS_p a_1716_n1348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.15
X37 comp_outp a_1950_n1721# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.139 pd=1.17 as=0.26 ps=2.3 w=0.84 l=0.15
X38 a_1716_n1348# a_1566_n378# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X39 VSS a_1716_n1348# a_482_n1818# VSS sky130_fd_pr__nfet_01v8 ad=0.0759 pd=0.79 as=0.0759 ps=0.79 w=0.46 l=0.15
X40 VSS clk a_582_n702# VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.31 ps=2.62 w=1 l=0.15
X41 a_582_n702# cdac_vn a_1830_n378# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.31 pd=2.62 as=0.165 ps=1.33 w=1 l=0.15
X42 VSS a_852_n296# a_476_n1721# VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.54 as=0.0759 ps=0.79 w=0.46 l=0.15
X43 a_1830_n378# a_1566_n378# a_1248_n288# VSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X44 a_852_n1721# a_476_n1266# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0.244 ps=2.26 w=0.84 l=0.15
X45 a_1830_n378# cdac_vn a_582_n702# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.165 pd=1.33 as=0.31 ps=2.62 w=1 l=0.15
X46 RS_p RS_n VDD VDD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.15
X47 VDD a_1950_n1721# comp_outp VDD sky130_fd_pr__pfet_01v8 ad=0.139 pd=1.17 as=0.139 ps=1.17 w=0.84 l=0.15
X48 a_1716_n1348# a_1566_n378# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0.244 ps=2.26 w=0.84 l=0.15
X49 a_1842_n702# clk VSS VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.165 ps=1.33 w=1 l=0.15
X50 VDD clk a_1390_109# VDD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X51 a_674_n702# cdac_vp a_582_n702# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X52 VSS a_1026_n1747# comp_outn VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.54 as=0.0759 ps=0.79 w=0.46 l=0.15
X53 comp_outp a_1950_n1721# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0759 pd=0.79 as=0.143 ps=1.54 w=0.46 l=0.15
X54 a_482_n1818# a_1716_n1348# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.139 pd=1.17 as=0.26 ps=2.3 w=0.84 l=0.15
X55 a_482_n1818# a_1716_n1348# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.3 as=0.139 ps=1.17 w=0.84 l=0.15
X56 a_582_n702# cdac_vp a_674_n702# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.31 pd=2.62 as=0.165 ps=1.33 w=1 l=0.15
X57 VSS a_852_n296# RS_n VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.15
X58 VDD a_1716_n1348# a_482_n1818# VDD sky130_fd_pr__pfet_01v8 ad=0.139 pd=1.17 as=0.139 ps=1.17 w=0.84 l=0.15
X59 a_1830_n378# cdac_vn a_582_n702# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X60 a_852_n1721# a_476_n1266# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X61 a_482_n1818# a_476_n1721# a_476_n1266# VDD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.15
X62 VSS a_1950_n1721# comp_outp VSS sky130_fd_pr__nfet_01v8 ad=0.0759 pd=0.79 as=0.0759 ps=0.79 w=0.46 l=0.15
X63 a_476_n1721# a_852_n296# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0759 pd=0.79 as=0.0759 ps=0.79 w=0.46 l=0.15
X64 VDD RS_n a_1026_n1747# VDD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0.244 ps=2.26 w=0.84 l=0.15
X65 VDD a_1248_n288# a_1566_n378# VDD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X66 a_1566_n378# a_1248_n288# a_674_n702# VSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X67 a_582_n702# cdac_vp a_674_n702# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X68 VSS clk a_582_n702# VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X69 VDD RS_p RS_n VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.15
.ends

