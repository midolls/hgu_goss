magic
tech sky130A
magscale 1 2
timestamp 1699830634
<< metal1 >>
rect 247 5371 311 5377
rect 247 5362 253 5371
rect 157 5328 253 5362
rect 247 5319 253 5328
rect 305 5319 311 5371
rect 2320 5363 2688 5392
rect 4426 5364 4669 5393
rect 1262 5360 1296 5362
rect 869 5326 1296 5360
rect 247 5313 311 5319
rect 1262 3048 1296 5326
rect 1250 3042 1314 3048
rect 1250 2990 1256 3042
rect 1308 2990 1314 3042
rect 2654 3030 2688 5363
rect 1250 2984 1314 2990
rect 2642 3024 2706 3030
rect 2642 2972 2648 3024
rect 2700 2972 2706 3024
rect 4635 2991 4669 5364
rect 8151 5354 8431 5383
rect 2642 2966 2706 2972
rect 4621 2985 4685 2991
rect 4621 2933 4627 2985
rect 4679 2933 4685 2985
rect 8397 2953 8431 5354
rect 15583 5322 15829 5351
rect 28405 5328 28681 5357
rect 4621 2927 4685 2933
rect 8383 2947 8447 2953
rect 8383 2895 8389 2947
rect 8441 2895 8447 2947
rect 15795 2940 15829 5322
rect 28647 2958 28681 5328
rect 28633 2952 28697 2958
rect 8383 2889 8447 2895
rect 15781 2934 15845 2940
rect 15781 2882 15787 2934
rect 15839 2882 15845 2934
rect 28633 2900 28639 2952
rect 28691 2900 28697 2952
rect 28633 2894 28697 2900
rect 15781 2876 15845 2882
<< via1 >>
rect 253 5319 305 5371
rect 1256 2990 1308 3042
rect 2648 2972 2700 3024
rect 4627 2933 4679 2985
rect 8389 2895 8441 2947
rect 15787 2882 15839 2934
rect 28639 2900 28691 2952
<< metal2 >>
rect 242 5373 316 5377
rect 242 5317 251 5373
rect 307 5317 316 5373
rect 242 5313 316 5317
rect 1250 3044 1314 3053
rect 1250 2988 1254 3044
rect 1310 2988 1314 3044
rect 1250 2979 1314 2988
rect 2642 3026 2706 3035
rect 2642 2970 2646 3026
rect 2702 2970 2706 3026
rect 2642 2961 2706 2970
rect 4621 2987 4685 2996
rect 4621 2931 4625 2987
rect 4681 2931 4685 2987
rect 4621 2922 4685 2931
rect 8383 2949 8447 2958
rect 8383 2893 8387 2949
rect 8443 2893 8447 2949
rect 28633 2954 28697 2963
rect 8383 2884 8447 2893
rect 15781 2936 15845 2945
rect 15781 2880 15785 2936
rect 15841 2880 15845 2936
rect 28633 2898 28637 2954
rect 28693 2898 28697 2954
rect 28633 2889 28697 2898
rect 15781 2871 15845 2880
<< via2 >>
rect 251 5371 307 5373
rect 251 5319 253 5371
rect 253 5319 305 5371
rect 305 5319 307 5371
rect 251 5317 307 5319
rect 1254 3042 1310 3044
rect 1254 2990 1256 3042
rect 1256 2990 1308 3042
rect 1308 2990 1310 3042
rect 1254 2988 1310 2990
rect 2646 3024 2702 3026
rect 2646 2972 2648 3024
rect 2648 2972 2700 3024
rect 2700 2972 2702 3024
rect 2646 2970 2702 2972
rect 4625 2985 4681 2987
rect 4625 2933 4627 2985
rect 4627 2933 4679 2985
rect 4679 2933 4681 2985
rect 4625 2931 4681 2933
rect 8387 2947 8443 2949
rect 8387 2895 8389 2947
rect 8389 2895 8441 2947
rect 8441 2895 8443 2947
rect 8387 2893 8443 2895
rect 15785 2934 15841 2936
rect 15785 2882 15787 2934
rect 15787 2882 15839 2934
rect 15839 2882 15841 2934
rect 15785 2880 15841 2882
rect 28637 2952 28693 2954
rect 28637 2900 28639 2952
rect 28639 2900 28691 2952
rect 28691 2900 28693 2952
rect 28637 2898 28693 2900
<< metal3 >>
rect 228 5373 328 5388
rect 228 5317 251 5373
rect 307 5317 328 5373
rect 228 5289 328 5317
rect 1232 3044 1331 3067
rect 1232 2988 1254 3044
rect 1310 2988 1331 3044
rect 1232 2967 1331 2988
rect 2624 3026 2723 3049
rect 2624 2970 2646 3026
rect 2702 2970 2723 3026
rect 2624 2949 2723 2970
rect 4625 2987 4681 3010
rect 4625 2910 4681 2931
rect 8387 2949 8443 2972
rect 8387 2872 8443 2893
rect 15780 2936 15846 2955
rect 15780 2880 15785 2936
rect 15841 2880 15846 2936
rect 15780 2859 15846 2880
rect 28632 2946 28633 2977
rect 28632 2932 28637 2946
rect 28632 2931 28636 2932
rect 28632 2898 28637 2931
rect 28697 2946 28698 2977
rect 28693 2933 28698 2946
rect 28694 2932 28698 2933
rect 28693 2898 28698 2932
rect 28632 2897 28642 2898
rect 28643 2897 28698 2898
rect 28632 2877 28698 2897
<< metal4 >>
rect 246 5094 312 5377
<< via4 >>
rect 1107 2839 1344 3075
rect 2505 2834 2742 3070
rect 4533 2836 4770 3072
rect 8295 2837 8532 3073
rect 15692 2837 15929 3073
rect 28546 2837 28783 3073
rect 1107 2240 1344 2476
rect 2505 2235 2742 2471
rect 4533 2237 4770 2473
rect 8295 2238 8532 2474
rect 15692 2238 15929 2474
rect 28546 2238 28783 2474
<< metal5 >>
rect 1065 3075 1388 3120
rect 1065 2839 1107 3075
rect 1344 2839 1388 3075
rect 1065 2476 1388 2839
rect 1065 2240 1107 2476
rect 1344 2240 1388 2476
rect 1065 2202 1388 2240
rect 2463 3070 2786 3115
rect 2463 2834 2505 3070
rect 2742 2834 2786 3070
rect 2463 2471 2786 2834
rect 2463 2235 2505 2471
rect 2742 2235 2786 2471
rect 2463 2197 2786 2235
rect 4491 3072 4814 3117
rect 4491 2836 4533 3072
rect 4770 2836 4814 3072
rect 4491 2473 4814 2836
rect 4491 2237 4533 2473
rect 4770 2237 4814 2473
rect 4491 2199 4814 2237
rect 8253 3073 8576 3118
rect 8253 2837 8295 3073
rect 8532 2837 8576 3073
rect 8253 2474 8576 2837
rect 8253 2238 8295 2474
rect 8532 2238 8576 2474
rect 8253 2200 8576 2238
rect 15650 3073 15973 3118
rect 15650 2837 15692 3073
rect 15929 2837 15973 3073
rect 15650 2474 15973 2837
rect 15650 2238 15692 2474
rect 15929 2238 15973 2474
rect 15650 2200 15973 2238
rect 28504 3073 28827 3118
rect 28504 2837 28546 3073
rect 28783 2837 28827 3073
rect 28504 2474 28827 2837
rect 28504 2238 28546 2474
rect 28783 2238 28827 2474
rect 28504 2200 28827 2238
use hgu_cdac_8bit_array  hgu_cdac_8bit_array_2
timestamp 1699813282
transform 1 0 4202 0 -1 -4800
box -4516 -7612 35404 -4800
use hgu_cdac_8bit_array  hgu_cdac_8bit_array_3
timestamp 1699813282
transform 1 0 4202 0 -1 -2312
box -4516 -7612 35404 -4800
use hgu_cdac_unit  hgu_cdac_unit_0
timestamp 1699173900
transform 1 0 -1000 0 -1 2044
box 686 598 1358 1826
use hgu_cdac_unit  hgu_cdac_unit_1
timestamp 1699173900
transform 1 0 -1000 0 -1 4532
box 686 598 1358 1826
use hgu_inverter  hgu_inverter_0
timestamp 1699345134
transform 1 0 -435 0 1 4948
box 347 160 675 824
use inv_2_test  inv_2_test_0
timestamp 1699782319
transform 1 0 258 0 1 2748
box 400 2360 856 3024
use inv_4_test  inv_4_test_0
timestamp 1699782319
transform 1 0 2266 0 1 3824
box -447 1324 265 1988
use inv_8_test  inv_8_test_0
timestamp 1699782319
transform 1 0 3317 0 1 2829
box 96 2320 1320 2984
use inv_16_test  inv_16_test_0
timestamp 1699782319
transform 1 0 6763 0 1 5179
box -649 -40 1599 624
use inv_32_test  inv_32_test_0
timestamp 1699782319
transform 1 0 13801 0 1 7509
box -2303 -2402 1993 -1738
use inv_64_test  inv_64_test_0
timestamp 1699782319
transform 1 0 23813 0 1 7515
box -3583 -2402 4809 -1738
<< labels >>
flabel metal1 165 5335 203 5356 0 FreeSans 160 0 0 0 d<0>
port 2 nsew
<< end >>
