magic
tech sky130A
magscale 1 2
timestamp 1697713470
<< nwell >>
rect -109 -116 110 116
<< pmos >>
rect -15 -80 15 80
<< pdiff >>
rect -73 -80 -15 80
rect 15 -80 73 80
<< poly >>
rect -15 80 15 111
rect -15 -127 15 -80
<< properties >>
string FIXED_BBOX -158 -246 158 246
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.8 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
