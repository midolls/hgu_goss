magic
tech sky130A
timestamp 1699890160
<< psubdiff >>
rect 744 2037 764 2092
<< metal4 >>
rect 469 2077 495 2097
rect 832 2019 858 2039
rect 531 1887 550 1928
use hgu_cdac_unit  x1[0]
timestamp 1699890160
transform 1 0 0 0 1 1100
box 343 299 679 913
use hgu_cdac_unit  x1[1]
timestamp 1699890160
transform -1 0 1022 0 -1 2892
box 343 299 679 913
use hgu_cdac_unit  x1[2]
timestamp 1699890160
transform 1 0 303 0 1 1100
box 343 299 679 913
use hgu_cdac_unit  x1[3]
timestamp 1699890160
transform -1 0 1325 0 -1 2892
box 343 299 679 913
<< labels >>
flabel metal4 832 2019 858 2039 0 FreeSans 160 0 0 0 CBOT
port 1 nsew
flabel metal4 469 2077 495 2097 0 FreeSans 160 0 0 0 CTOP
port 3 nsew
flabel psubdiff 744 2037 764 2092 0 FreeSans 160 0 0 0 SUB
port 5 nsew
flabel metal4 531 1887 550 1928 0 FreeSans 160 0 0 0 CTOP
port 7 nsew
<< end >>
