magic
tech sky130A
magscale 1 2
timestamp 1699172750
<< nwell >>
rect 1 80 1277 1356
rect 467 0 811 80
<< pmos >>
rect 561 49 591 133
rect 687 49 717 133
<< pdiff >>
rect 503 121 561 133
rect 503 61 515 121
rect 549 61 561 121
rect 503 49 561 61
rect 591 49 687 133
rect 717 121 775 133
rect 717 61 729 121
rect 763 61 775 121
rect 717 49 775 61
<< pdiffc >>
rect 515 61 549 121
rect 729 61 763 121
<< nsubdiff >>
rect 71 1290 609 1310
rect 71 1256 119 1290
rect 153 1256 199 1290
rect 233 1256 279 1290
rect 313 1256 359 1290
rect 393 1256 439 1290
rect 473 1256 519 1290
rect 553 1256 609 1290
rect 71 1242 609 1256
rect 669 1290 1207 1310
rect 669 1256 725 1290
rect 759 1256 805 1290
rect 839 1256 885 1290
rect 919 1256 965 1290
rect 999 1256 1045 1290
rect 1079 1256 1125 1290
rect 1159 1256 1207 1290
rect 669 1242 1207 1256
<< nsubdiffcont >>
rect 119 1256 153 1290
rect 199 1256 233 1290
rect 279 1256 313 1290
rect 359 1256 393 1290
rect 439 1256 473 1290
rect 519 1256 553 1290
rect 725 1256 759 1290
rect 805 1256 839 1290
rect 885 1256 919 1290
rect 965 1256 999 1290
rect 1045 1256 1079 1290
rect 1125 1256 1159 1290
<< poly >>
rect 543 214 609 230
rect 543 180 559 214
rect 593 180 609 214
rect 543 164 609 180
rect 669 214 735 230
rect 669 180 685 214
rect 719 180 735 214
rect 669 164 735 180
rect 561 133 591 164
rect 687 133 717 164
rect 561 21 591 49
rect 687 21 717 49
<< polycont >>
rect 559 180 593 214
rect 685 180 719 214
<< locali >>
rect 3 1290 1275 1308
rect 3 1256 119 1290
rect 155 1256 199 1290
rect 235 1256 279 1290
rect 315 1256 359 1290
rect 395 1256 439 1290
rect 475 1256 519 1290
rect 555 1256 723 1290
rect 759 1256 803 1290
rect 839 1256 883 1290
rect 919 1256 963 1290
rect 999 1256 1043 1290
rect 1079 1256 1123 1290
rect 1159 1256 1275 1290
rect 3 1242 1275 1256
rect 543 180 559 214
rect 593 180 609 214
rect 669 180 685 214
rect 719 180 735 214
rect 515 121 549 137
rect 515 45 549 61
rect 729 121 763 137
rect 729 45 763 61
<< viali >>
rect 121 1256 153 1290
rect 153 1256 155 1290
rect 201 1256 233 1290
rect 233 1256 235 1290
rect 281 1256 313 1290
rect 313 1256 315 1290
rect 361 1256 393 1290
rect 393 1256 395 1290
rect 441 1256 473 1290
rect 473 1256 475 1290
rect 521 1256 553 1290
rect 553 1256 555 1290
rect 723 1256 725 1290
rect 725 1256 757 1290
rect 803 1256 805 1290
rect 805 1256 837 1290
rect 883 1256 885 1290
rect 885 1256 917 1290
rect 963 1256 965 1290
rect 965 1256 997 1290
rect 1043 1256 1045 1290
rect 1045 1256 1077 1290
rect 1123 1256 1125 1290
rect 1125 1256 1157 1290
rect 559 180 593 214
rect 685 180 719 214
rect 515 61 549 121
rect 729 61 763 121
<< metal1 >>
rect 3 1302 1275 1308
rect 3 1250 111 1302
rect 163 1250 191 1302
rect 243 1250 271 1302
rect 323 1250 351 1302
rect 403 1250 431 1302
rect 483 1250 511 1302
rect 563 1250 715 1302
rect 767 1250 795 1302
rect 847 1250 875 1302
rect 927 1250 955 1302
rect 1007 1250 1035 1302
rect 1087 1250 1115 1302
rect 1167 1250 1275 1302
rect 3 1242 1275 1250
rect 546 214 733 220
rect 546 180 559 214
rect 593 180 685 214
rect 719 180 733 214
rect 546 173 733 180
rect 509 125 555 133
rect 723 125 769 133
rect 486 124 565 125
rect 486 60 493 124
rect 557 60 565 124
rect 713 124 792 125
rect 713 60 721 124
rect 785 60 792 124
rect 509 49 555 60
rect 723 49 769 60
<< via1 >>
rect 111 1290 163 1302
rect 111 1256 121 1290
rect 121 1256 155 1290
rect 155 1256 163 1290
rect 111 1250 163 1256
rect 191 1290 243 1302
rect 191 1256 201 1290
rect 201 1256 235 1290
rect 235 1256 243 1290
rect 191 1250 243 1256
rect 271 1290 323 1302
rect 271 1256 281 1290
rect 281 1256 315 1290
rect 315 1256 323 1290
rect 271 1250 323 1256
rect 351 1290 403 1302
rect 351 1256 361 1290
rect 361 1256 395 1290
rect 395 1256 403 1290
rect 351 1250 403 1256
rect 431 1290 483 1302
rect 431 1256 441 1290
rect 441 1256 475 1290
rect 475 1256 483 1290
rect 431 1250 483 1256
rect 511 1290 563 1302
rect 511 1256 521 1290
rect 521 1256 555 1290
rect 555 1256 563 1290
rect 511 1250 563 1256
rect 715 1290 767 1302
rect 715 1256 723 1290
rect 723 1256 757 1290
rect 757 1256 767 1290
rect 715 1250 767 1256
rect 795 1290 847 1302
rect 795 1256 803 1290
rect 803 1256 837 1290
rect 837 1256 847 1290
rect 795 1250 847 1256
rect 875 1290 927 1302
rect 875 1256 883 1290
rect 883 1256 917 1290
rect 917 1256 927 1290
rect 875 1250 927 1256
rect 955 1290 1007 1302
rect 955 1256 963 1290
rect 963 1256 997 1290
rect 997 1256 1007 1290
rect 955 1250 1007 1256
rect 1035 1290 1087 1302
rect 1035 1256 1043 1290
rect 1043 1256 1077 1290
rect 1077 1256 1087 1290
rect 1035 1250 1087 1256
rect 1115 1290 1167 1302
rect 1115 1256 1123 1290
rect 1123 1256 1157 1290
rect 1157 1256 1167 1290
rect 1115 1250 1167 1256
rect 493 121 557 124
rect 493 61 515 121
rect 515 61 549 121
rect 549 61 557 121
rect 493 60 557 61
rect 721 121 785 124
rect 721 61 729 121
rect 729 61 763 121
rect 763 61 785 121
rect 721 60 785 61
<< metal2 >>
rect 3 1304 1275 1308
rect 3 1248 107 1304
rect 163 1248 187 1304
rect 243 1248 267 1304
rect 323 1248 347 1304
rect 403 1248 427 1304
rect 483 1248 507 1304
rect 563 1248 715 1304
rect 771 1248 795 1304
rect 851 1248 875 1304
rect 931 1248 955 1304
rect 1011 1248 1035 1304
rect 1091 1248 1115 1304
rect 1171 1248 1275 1304
rect 3 1242 1275 1248
rect 486 124 565 125
rect 713 124 792 125
rect 483 60 493 124
rect 557 60 566 124
rect 712 60 721 124
rect 785 60 795 124
<< via2 >>
rect 107 1302 163 1304
rect 107 1250 111 1302
rect 111 1250 163 1302
rect 107 1248 163 1250
rect 187 1302 243 1304
rect 187 1250 191 1302
rect 191 1250 243 1302
rect 187 1248 243 1250
rect 267 1302 323 1304
rect 267 1250 271 1302
rect 271 1250 323 1302
rect 267 1248 323 1250
rect 347 1302 403 1304
rect 347 1250 351 1302
rect 351 1250 403 1302
rect 347 1248 403 1250
rect 427 1302 483 1304
rect 427 1250 431 1302
rect 431 1250 483 1302
rect 427 1248 483 1250
rect 507 1302 563 1304
rect 507 1250 511 1302
rect 511 1250 563 1302
rect 507 1248 563 1250
rect 715 1302 771 1304
rect 715 1250 767 1302
rect 767 1250 771 1302
rect 715 1248 771 1250
rect 795 1302 851 1304
rect 795 1250 847 1302
rect 847 1250 851 1302
rect 795 1248 851 1250
rect 875 1302 931 1304
rect 875 1250 927 1302
rect 927 1250 931 1302
rect 875 1248 931 1250
rect 955 1302 1011 1304
rect 955 1250 1007 1302
rect 1007 1250 1011 1302
rect 955 1248 1011 1250
rect 1035 1302 1091 1304
rect 1035 1250 1087 1302
rect 1087 1250 1091 1302
rect 1035 1248 1091 1250
rect 1115 1302 1171 1304
rect 1115 1250 1167 1302
rect 1167 1250 1171 1302
rect 1115 1248 1171 1250
rect 493 60 557 124
rect 721 60 785 124
<< metal3 >>
rect 0 1307 1278 1309
rect 0 1243 104 1307
rect 168 1243 184 1307
rect 248 1243 264 1307
rect 328 1243 344 1307
rect 408 1243 424 1307
rect 488 1243 504 1307
rect 568 1243 710 1307
rect 774 1243 790 1307
rect 854 1243 870 1307
rect 934 1243 950 1307
rect 1014 1243 1030 1307
rect 1094 1243 1110 1307
rect 1174 1243 1278 1307
rect 0 1241 1278 1243
rect 0 1087 66 1177
rect 0 1023 1 1087
rect 65 1023 66 1087
rect 0 1007 66 1023
rect 0 943 1 1007
rect 65 943 66 1007
rect 0 927 66 943
rect 0 863 1 927
rect 65 863 66 927
rect 0 847 66 863
rect 0 783 1 847
rect 65 783 66 847
rect 0 767 66 783
rect 0 703 1 767
rect 65 703 66 767
rect 0 687 66 703
rect 0 623 1 687
rect 65 623 66 687
rect 0 607 66 623
rect 0 543 1 607
rect 65 543 66 607
rect 0 527 66 543
rect 0 463 1 527
rect 65 463 66 527
rect 0 447 66 463
rect 0 383 1 447
rect 65 383 66 447
rect 0 367 66 383
rect 0 303 1 367
rect 65 303 66 367
rect 0 149 66 303
rect 126 149 186 1181
rect 246 211 306 1241
rect 366 149 426 1181
rect 486 211 546 1241
rect 606 1087 672 1177
rect 606 1023 607 1087
rect 671 1023 672 1087
rect 606 1007 672 1023
rect 606 943 607 1007
rect 671 943 672 1007
rect 606 927 672 943
rect 606 863 607 927
rect 671 863 672 927
rect 606 847 672 863
rect 606 783 607 847
rect 671 783 672 847
rect 606 767 672 783
rect 606 703 607 767
rect 671 703 672 767
rect 606 687 672 703
rect 606 623 607 687
rect 671 623 672 687
rect 606 607 672 623
rect 606 543 607 607
rect 671 543 672 607
rect 606 527 672 543
rect 606 463 607 527
rect 671 463 672 527
rect 606 447 672 463
rect 606 383 607 447
rect 671 383 672 447
rect 606 367 672 383
rect 606 303 607 367
rect 671 303 672 367
rect 606 149 672 303
rect 732 211 792 1241
rect 852 149 912 1181
rect 972 211 1032 1241
rect 1092 149 1152 1181
rect 1212 1087 1278 1177
rect 1212 1023 1213 1087
rect 1277 1023 1278 1087
rect 1212 1007 1278 1023
rect 1212 943 1213 1007
rect 1277 943 1278 1007
rect 1212 927 1278 943
rect 1212 863 1213 927
rect 1277 863 1278 927
rect 1212 847 1278 863
rect 1212 783 1213 847
rect 1277 783 1278 847
rect 1212 767 1278 783
rect 1212 703 1213 767
rect 1277 703 1278 767
rect 1212 687 1278 703
rect 1212 623 1213 687
rect 1277 623 1278 687
rect 1212 607 1278 623
rect 1212 543 1213 607
rect 1277 543 1278 607
rect 1212 527 1278 543
rect 1212 463 1213 527
rect 1277 463 1278 527
rect 1212 447 1278 463
rect 1212 383 1213 447
rect 1277 383 1278 447
rect 1212 367 1278 383
rect 1212 303 1213 367
rect 1277 303 1278 367
rect 1212 149 1278 303
rect 0 147 1278 149
rect 0 83 104 147
rect 168 83 184 147
rect 248 83 264 147
rect 328 83 344 147
rect 408 83 424 147
rect 488 124 504 147
rect 488 83 493 124
rect 568 83 710 147
rect 774 124 790 147
rect 785 83 790 124
rect 854 83 870 147
rect 934 83 950 147
rect 1014 83 1030 147
rect 1094 83 1110 147
rect 1174 83 1278 147
rect 0 81 493 83
rect 483 60 493 81
rect 557 81 721 83
rect 557 60 566 81
rect 483 55 566 60
rect 712 60 721 81
rect 785 81 1278 83
rect 785 60 795 81
rect 712 55 795 60
<< via3 >>
rect 104 1304 168 1307
rect 104 1248 107 1304
rect 107 1248 163 1304
rect 163 1248 168 1304
rect 104 1243 168 1248
rect 184 1304 248 1307
rect 184 1248 187 1304
rect 187 1248 243 1304
rect 243 1248 248 1304
rect 184 1243 248 1248
rect 264 1304 328 1307
rect 264 1248 267 1304
rect 267 1248 323 1304
rect 323 1248 328 1304
rect 264 1243 328 1248
rect 344 1304 408 1307
rect 344 1248 347 1304
rect 347 1248 403 1304
rect 403 1248 408 1304
rect 344 1243 408 1248
rect 424 1304 488 1307
rect 424 1248 427 1304
rect 427 1248 483 1304
rect 483 1248 488 1304
rect 424 1243 488 1248
rect 504 1304 568 1307
rect 504 1248 507 1304
rect 507 1248 563 1304
rect 563 1248 568 1304
rect 504 1243 568 1248
rect 710 1304 774 1307
rect 710 1248 715 1304
rect 715 1248 771 1304
rect 771 1248 774 1304
rect 710 1243 774 1248
rect 790 1304 854 1307
rect 790 1248 795 1304
rect 795 1248 851 1304
rect 851 1248 854 1304
rect 790 1243 854 1248
rect 870 1304 934 1307
rect 870 1248 875 1304
rect 875 1248 931 1304
rect 931 1248 934 1304
rect 870 1243 934 1248
rect 950 1304 1014 1307
rect 950 1248 955 1304
rect 955 1248 1011 1304
rect 1011 1248 1014 1304
rect 950 1243 1014 1248
rect 1030 1304 1094 1307
rect 1030 1248 1035 1304
rect 1035 1248 1091 1304
rect 1091 1248 1094 1304
rect 1030 1243 1094 1248
rect 1110 1304 1174 1307
rect 1110 1248 1115 1304
rect 1115 1248 1171 1304
rect 1171 1248 1174 1304
rect 1110 1243 1174 1248
rect 1 1023 65 1087
rect 1 943 65 1007
rect 1 863 65 927
rect 1 783 65 847
rect 1 703 65 767
rect 1 623 65 687
rect 1 543 65 607
rect 1 463 65 527
rect 1 383 65 447
rect 1 303 65 367
rect 607 1023 671 1087
rect 607 943 671 1007
rect 607 863 671 927
rect 607 783 671 847
rect 607 703 671 767
rect 607 623 671 687
rect 607 543 671 607
rect 607 463 671 527
rect 607 383 671 447
rect 607 303 671 367
rect 1213 1023 1277 1087
rect 1213 943 1277 1007
rect 1213 863 1277 927
rect 1213 783 1277 847
rect 1213 703 1277 767
rect 1213 623 1277 687
rect 1213 543 1277 607
rect 1213 463 1277 527
rect 1213 383 1277 447
rect 1213 303 1277 367
rect 104 83 168 147
rect 184 83 248 147
rect 264 83 328 147
rect 344 83 408 147
rect 424 83 488 147
rect 504 124 568 147
rect 504 83 557 124
rect 557 83 568 124
rect 710 124 774 147
rect 710 83 721 124
rect 721 83 774 124
rect 790 83 854 147
rect 870 83 934 147
rect 950 83 1014 147
rect 1030 83 1094 147
rect 1110 83 1174 147
<< metal4 >>
rect 3 1309 1275 1310
rect 0 1307 1278 1309
rect 0 1243 104 1307
rect 168 1243 184 1307
rect 248 1243 264 1307
rect 328 1243 344 1307
rect 408 1243 424 1307
rect 488 1243 504 1307
rect 568 1243 710 1307
rect 774 1243 790 1307
rect 854 1243 870 1307
rect 934 1243 950 1307
rect 1014 1243 1030 1307
rect 1094 1243 1110 1307
rect 1174 1243 1278 1307
rect 0 1241 1278 1243
rect 0 1087 66 1177
rect 0 1023 1 1087
rect 65 1023 66 1087
rect 0 1007 66 1023
rect 0 943 1 1007
rect 65 943 66 1007
rect 0 927 66 943
rect 0 863 1 927
rect 65 863 66 927
rect 0 847 66 863
rect 0 783 1 847
rect 65 783 66 847
rect 0 767 66 783
rect 0 703 1 767
rect 65 703 66 767
rect 0 687 66 703
rect 0 623 1 687
rect 65 623 66 687
rect 0 607 66 623
rect 0 543 1 607
rect 65 543 66 607
rect 0 527 66 543
rect 0 463 1 527
rect 65 463 66 527
rect 0 447 66 463
rect 0 383 1 447
rect 65 383 66 447
rect 0 367 66 383
rect 0 303 1 367
rect 65 303 66 367
rect 0 149 66 303
rect 126 211 186 1241
rect 246 149 306 1181
rect 366 211 426 1241
rect 486 149 546 1181
rect 606 1087 672 1177
rect 606 1023 607 1087
rect 671 1023 672 1087
rect 606 1007 672 1023
rect 606 943 607 1007
rect 671 943 672 1007
rect 606 927 672 943
rect 606 863 607 927
rect 671 863 672 927
rect 606 847 672 863
rect 606 783 607 847
rect 671 783 672 847
rect 606 767 672 783
rect 606 703 607 767
rect 671 703 672 767
rect 606 687 672 703
rect 606 623 607 687
rect 671 623 672 687
rect 606 607 672 623
rect 606 543 607 607
rect 671 543 672 607
rect 606 527 672 543
rect 606 463 607 527
rect 671 463 672 527
rect 606 447 672 463
rect 606 383 607 447
rect 671 383 672 447
rect 606 367 672 383
rect 606 303 607 367
rect 671 303 672 367
rect 606 149 672 303
rect 732 149 792 1181
rect 852 211 912 1241
rect 972 149 1032 1181
rect 1092 211 1152 1241
rect 1212 1087 1278 1177
rect 1212 1023 1213 1087
rect 1277 1023 1278 1087
rect 1212 1007 1278 1023
rect 1212 943 1213 1007
rect 1277 943 1278 1007
rect 1212 927 1278 943
rect 1212 863 1213 927
rect 1277 863 1278 927
rect 1212 847 1278 863
rect 1212 783 1213 847
rect 1277 783 1278 847
rect 1212 767 1278 783
rect 1212 703 1213 767
rect 1277 703 1278 767
rect 1212 687 1278 703
rect 1212 623 1213 687
rect 1277 623 1278 687
rect 1212 607 1278 623
rect 1212 543 1213 607
rect 1277 543 1278 607
rect 1212 527 1278 543
rect 1212 463 1213 527
rect 1277 463 1278 527
rect 1212 447 1278 463
rect 1212 383 1213 447
rect 1277 383 1278 447
rect 1212 367 1278 383
rect 1212 303 1213 367
rect 1277 303 1278 367
rect 1212 149 1278 303
rect 0 147 1278 149
rect 0 83 104 147
rect 168 83 184 147
rect 248 83 264 147
rect 328 83 344 147
rect 408 83 424 147
rect 488 83 504 147
rect 568 83 710 147
rect 774 83 790 147
rect 854 83 870 147
rect 934 83 950 147
rect 1014 83 1030 147
rect 1094 83 1110 147
rect 1174 83 1278 147
rect 0 81 1278 83
<< labels >>
flabel metal1 685 180 719 214 0 FreeSans 320 0 0 0 hgu_sw_cap_pmos_0.SW
flabel pdiff 629 49 687 133 0 FreeSans 320 0 0 0 hgu_sw_cap_pmos_0.delay_signal
flabel metal3 605 1242 1275 1310 0 FreeSans 320 0 0 0 hgu_sw_cap_pmos_0.VDD
flabel metal1 559 180 593 214 0 FreeSans 320 0 0 0 hgu_sw_cap_pmos_1.SW
flabel pdiff 591 49 649 133 0 FreeSans 320 0 0 0 hgu_sw_cap_pmos_1.delay_signal
flabel metal3 3 1242 673 1310 0 FreeSans 320 0 0 0 hgu_sw_cap_pmos_1.VDD
<< end >>
