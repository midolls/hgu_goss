magic
tech sky130A
timestamp 1698655397
<< end >>
