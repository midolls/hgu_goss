* NGSPICE file created from hgu_cdac_sw_buffer_flat.ext - technology: sky130A

.subckt hgu_cdac_sw_buffer_RC sar_val<7> sar_val<6> sar_val<5> sar_val<4> sar_val<3>
+ sw<6> sw<2> sw<3> sw<4> sw<5> VSS VDD
X0 sw<6>.t25 a_n85_n1195# VDD.t50 VDD.t49 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 VSS.t92 a_795_n2019# sw<5>.t1 VSS.t91 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 sw<6>.t24 a_n85_n1195# VDD.t48 VDD.t47 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3 VSS.t21 a_1317_n2468# x8.X VSS.t20 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X4 x11.A a_1347_n2019# VDD.t58 VDD.t57 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5 VDD.t56 a_1347_n2019# x11.A VDD.t55 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_n85_n1195# x11.A VSS.t67 VSS.t66 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 VSS.t49 a_n85_n1195# sw<6>.t2 VSS.t48 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 VDD.t46 a_n85_n1195# sw<6>.t23 VDD.t45 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_n85_n1195# x11.A VDD.t72 VDD.t71 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 VSS.t47 a_n85_n1195# sw<6>.t1 VSS.t46 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 VSS.t82 sar_val<7>.t0 a_1543_n2633# VSS.t81 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X12 VSS.t45 a_n85_n1195# sw<6>.t5 VSS.t44 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 VDD.t44 a_n85_n1195# sw<6>.t22 VDD.t43 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 x3.X a_991_n2633# VSS.t5 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X15 VDD.t42 a_n85_n1195# sw<6>.t21 VDD.t41 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 sw<2>.t0 a_n113_n2633# VSS.t69 VSS.t68 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X17 sw<6>.t0 a_n85_n1195# VSS.t43 VSS.t42 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X18 VSS.t41 a_n85_n1195# sw<6>.t28 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X19 VDD.t40 a_n85_n1195# sw<6>.t20 VDD.t39 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 VSS.t19 a_765_n2468# x12.X VSS.t18 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X21 sw<5>.t7 a_795_n2019# VDD.t88 VDD.t87 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X22 VSS.t1 sar_val<3>.t0 a_n113_n2633# VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X23 sw<6>.t19 a_n85_n1195# VDD.t38 VDD.t37 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X24 sw<3>.t0 a_163_n2633# VSS.t80 VSS.t79 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X25 VDD.t93 sar_val<6>.t0 a_991_n2633# VDD.t92 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X26 x11.A a_1347_n2019# VDD.t54 VDD.t53 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 a_n85_n1195# x11.A VSS.t65 VSS.t56 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X28 a_255_n2019# x4.X VSS.t96 VSS.t35 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X29 VSS.t64 x11.A a_n85_n1195# VSS.t63 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X30 VDD.t70 x11.A a_n85_n1195# VDD.t69 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X31 a_n85_n1195# x11.A VDD.t68 VDD.t67 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X32 VDD.t80 sar_val<4>.t0 a_163_n2633# VDD.t79 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X33 a_795_n2019# x3.X VDD.t6 VDD.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X34 sw<4>.t3 a_255_n2019# VSS.t17 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X35 a_n85_n1195# x11.A VSS.t62 VSS.t54 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X36 VSS.t61 x11.A a_n85_n1195# VSS.t52 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X37 VDD.t66 x11.A a_n85_n1195# VDD.t65 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X38 a_n85_n1195# x11.A VDD.t64 VDD.t63 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X39 x4.X a_439_n2633# VDD.t97 VDD.t96 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X40 VDD.t90 sar_val<5>.t0 a_439_n2633# VDD.t89 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X41 sw<6>.t31 a_n85_n1195# VSS.t40 VSS.t39 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X42 sw<5>.t6 a_795_n2019# VDD.t86 VDD.t85 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X43 sw<6>.t18 a_n85_n1195# VDD.t36 VDD.t35 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X44 VDD.t84 a_795_n2019# sw<5>.t5 VDD.t83 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X45 VSS.t78 VSS.t76 a_n101_n1993# VSS.t77 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X46 VDD.t82 a_795_n2019# sw<5>.t4 VDD.t81 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X47 VSS.t95 sar_val<6>.t1 a_991_n2633# VSS.t94 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X48 x7.X a_n101_n1993# VSS.t59 VSS.t58 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X49 VDD.t5 VSS.t99 a_n101_n1993# VDD.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X50 VSS.t60 x11.A a_n85_n1195# VSS.t50 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X51 sw<4>.t2 a_255_n2019# VSS.t15 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X52 VDD.t62 x11.A a_n85_n1195# VDD.t61 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X53 VSS.t84 sar_val<4>.t1 a_163_n2633# VSS.t83 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X54 x7.X a_n101_n1993# VDD.t60 VDD.t59 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X55 VSS.t13 a_255_n2019# sw<4>.t1 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X56 x4.X a_439_n2633# VSS.t98 VSS.t97 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X57 VSS.t7 sar_val<5>.t1 a_439_n2633# VSS.t6 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X58 a_255_n2019# x4.X VDD.t95 VDD.t94 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X59 sw<4>.t7 a_255_n2019# VDD.t14 VDD.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X60 a_1317_n2468# VSS.t100 VDD.t99 VDD.t98 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X61 VSS.t11 a_255_n2019# sw<4>.t0 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X62 VSS.t38 a_n85_n1195# sw<6>.t3 VSS.t37 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X63 VDD.t34 a_n85_n1195# sw<6>.t17 VDD.t33 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X64 x9.X a_1543_n2633# VDD.t1 VDD.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X65 VSS.t57 a_1347_n2019# x11.A VSS.t56 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X66 a_1347_n2019# x9.X VSS.t93 VSS.t63 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X67 a_765_n2468# VSS.t101 VDD.t101 VDD.t100 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X68 VSS.t55 a_1347_n2019# x11.A VSS.t54 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X69 x11.A a_1347_n2019# VSS.t53 VSS.t52 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X70 sw<4>.t6 a_255_n2019# VDD.t12 VDD.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X71 sw<6>.t7 a_n85_n1195# VSS.t36 VSS.t35 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X72 sw<6>.t16 a_n85_n1195# VDD.t32 VDD.t31 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X73 VDD.t10 a_255_n2019# sw<4>.t5 VDD.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X74 a_1317_n2468# VSS.t73 VSS.t75 VSS.t74 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X75 sw<6>.t29 a_n85_n1195# VSS.t34 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X76 sw<6>.t15 a_n85_n1195# VDD.t30 VDD.t29 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X77 VSS.t33 a_n85_n1195# sw<6>.t27 VSS.t32 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X78 VDD.t28 a_n85_n1195# sw<6>.t14 VDD.t27 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X79 sw<5>.t3 a_795_n2019# VSS.t90 VSS.t89 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X80 VDD.t18 a_1317_n2468# x8.X VDD.t17 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X81 x9.X a_1543_n2633# VSS.t3 VSS.t2 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X82 x11.A a_1347_n2019# VSS.t51 VSS.t50 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X83 a_765_n2468# VSS.t70 VSS.t72 VSS.t71 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X84 VDD.t103 sar_val<7>.t1 a_1543_n2633# VDD.t102 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X85 sw<6>.t9 a_n85_n1195# VSS.t31 VSS.t30 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X86 sw<6>.t13 a_n85_n1195# VDD.t26 VDD.t25 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X87 x3.X a_991_n2633# VDD.t3 VDD.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X88 sw<2>.t1 a_n113_n2633# VDD.t76 VDD.t75 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X89 VDD.t8 a_255_n2019# sw<4>.t4 VDD.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X90 a_795_n2019# x3.X VSS.t9 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X91 sw<6>.t4 a_n85_n1195# VSS.t29 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X92 VSS.t28 a_n85_n1195# sw<6>.t6 VSS.t27 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X93 sw<6>.t12 a_n85_n1195# VDD.t24 VDD.t23 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X94 VDD.t22 a_n85_n1195# sw<6>.t11 VDD.t21 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X95 VDD.t16 a_765_n2468# x12.X VDD.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X96 VDD.t74 sar_val<3>.t1 a_n113_n2633# VDD.t73 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X97 sw<3>.t1 a_163_n2633# VDD.t78 VDD.t77 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X98 sw<5>.t0 a_795_n2019# VSS.t88 VSS.t87 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X99 VDD.t52 a_1347_n2019# x11.A VDD.t51 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X100 a_1347_n2019# x9.X VDD.t91 VDD.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X101 VSS.t86 a_795_n2019# sw<5>.t2 VSS.t85 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X102 VSS.t26 a_n85_n1195# sw<6>.t26 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X103 VDD.t20 a_n85_n1195# sw<6>.t10 VDD.t19 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X104 sw<6>.t8 a_n85_n1195# VSS.t25 VSS.t24 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X105 sw<6>.t30 a_n85_n1195# VSS.t23 VSS.t22 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R0 VDD.n326 VDD.t48 201.19
R1 VDD.n316 VDD.n315 174.595
R2 VDD.n310 VDD.n309 174.595
R3 VDD.n300 VDD.n299 174.595
R4 VDD.n290 VDD.n289 174.595
R5 VDD.n280 VDD.n279 174.595
R6 VDD.n270 VDD.n269 174.595
R7 VDD.n65 VDD.n64 174.595
R8 VDD.n59 VDD.n58 174.595
R9 VDD.n36 VDD.n35 174.595
R10 VDD.n18 VDD.n17 174.595
R11 VDD.n128 VDD.n127 166.381
R12 VDD.n109 VDD.n108 166.381
R13 VDD.n175 VDD.n174 166.381
R14 VDD.n325 VDD.t47 164.006
R15 VDD.n199 VDD.n198 162.47
R16 VDD.n213 VDD.n212 162.47
R17 VDD.n231 VDD.n230 162.47
R18 VDD.n99 VDD.n95 162.47
R19 VDD.n110 VDD.n107 162.47
R20 VDD.n157 VDD.n124 162.47
R21 VDD.n132 VDD.n126 162.47
R22 VDD.n186 VDD.n185 162.47
R23 VDD.n149 VDD.n148 160.918
R24 VDD.n94 VDD.n93 160.918
R25 VDD.n181 VDD.n179 160.918
R26 VDD.n2 VDD.t70 159.46
R27 VDD.n119 VDD.t58 142.571
R28 VDD.n96 VDD.t88 142.571
R29 VDD.n183 VDD.t14 142.571
R30 VDD.n4 VDD.t69 112.367
R31 VDD.n281 VDD.t21 112.367
R32 VDD VDD.n129 111.127
R33 VDD.n4 VDD.t63 102.151
R34 VDD.n281 VDD.t37 102.151
R35 VDD.n146 VDD.n145 92.5005
R36 VDD.n147 VDD.n146 92.5005
R37 VDD.n132 VDD.n131 92.5005
R38 VDD.n131 VDD.n130 92.5005
R39 VDD.n235 VDD.n234 92.5005
R40 VDD.n236 VDD.n235 92.5005
R41 VDD.n228 VDD.n227 92.5005
R42 VDD.n227 VDD.n226 92.5005
R43 VDD.n195 VDD.n194 92.5005
R44 VDD.n194 VDD.n193 92.5005
R45 VDD.n189 VDD.n188 92.5005
R46 VDD.n188 VDD.n187 92.5005
R47 VDD.n206 VDD.n205 92.5005
R48 VDD.n207 VDD.n206 92.5005
R49 VDD.n210 VDD.n209 92.5005
R50 VDD.n209 VDD.n208 92.5005
R51 VDD.n221 VDD.n220 92.5005
R52 VDD.n220 VDD.n219 92.5005
R53 VDD.n224 VDD.n223 92.5005
R54 VDD.n225 VDD.n224 92.5005
R55 VDD.n239 VDD.n238 92.5005
R56 VDD.n238 VDD.n237 92.5005
R57 VDD.n171 VDD.n170 92.5005
R58 VDD.n170 VDD.n169 92.5005
R59 VDD.n99 VDD.n98 92.5005
R60 VDD.n98 VDD.n97 92.5005
R61 VDD.n246 VDD.n245 92.5005
R62 VDD.n247 VDD.n246 92.5005
R63 VDD.n250 VDD.n249 92.5005
R64 VDD.n249 VDD.n248 92.5005
R65 VDD.n111 VDD.n110 92.5005
R66 VDD.n112 VDD.n111 92.5005
R67 VDD.n115 VDD.n114 92.5005
R68 VDD.n114 VDD.n113 92.5005
R69 VDD.n122 VDD.n121 92.5005
R70 VDD.n121 VDD.n120 92.5005
R71 VDD.n156 VDD.n155 92.5005
R72 VDD.n155 VDD.n154 92.5005
R73 VDD.n152 VDD.n151 92.5005
R74 VDD.n153 VDD.n152 92.5005
R75 VDD.n129 VDD.n125 92.5005
R76 VDD.n323 VDD.n322 92.5005
R77 VDD.n322 VDD.n321 92.5005
R78 VDD.n319 VDD.n318 92.5005
R79 VDD.n318 VDD.n317 92.5005
R80 VDD.n313 VDD.n312 92.5005
R81 VDD.n312 VDD.n311 92.5005
R82 VDD.n307 VDD.n306 92.5005
R83 VDD.n306 VDD.n305 92.5005
R84 VDD.n303 VDD.n302 92.5005
R85 VDD.n302 VDD.n301 92.5005
R86 VDD.n297 VDD.n296 92.5005
R87 VDD.n296 VDD.n295 92.5005
R88 VDD.n293 VDD.n292 92.5005
R89 VDD.n292 VDD.n291 92.5005
R90 VDD.n287 VDD.n286 92.5005
R91 VDD.n286 VDD.n285 92.5005
R92 VDD.n283 VDD.n282 92.5005
R93 VDD.n282 VDD.n281 92.5005
R94 VDD.n277 VDD.n276 92.5005
R95 VDD.n276 VDD.n275 92.5005
R96 VDD.n273 VDD.n272 92.5005
R97 VDD.n272 VDD.n271 92.5005
R98 VDD.n75 VDD.n74 92.5005
R99 VDD.n74 VDD.n73 92.5005
R100 VDD.n68 VDD.n67 92.5005
R101 VDD.n67 VDD.n66 92.5005
R102 VDD.n6 VDD.n5 92.5005
R103 VDD.n5 VDD.n4 92.5005
R104 VDD.n21 VDD.n20 92.5005
R105 VDD.n20 VDD.n19 92.5005
R106 VDD.n25 VDD.n24 92.5005
R107 VDD.n24 VDD.n23 92.5005
R108 VDD.n40 VDD.n38 92.5005
R109 VDD.n38 VDD.n37 92.5005
R110 VDD.n47 VDD.n46 92.5005
R111 VDD.n46 VDD.n45 92.5005
R112 VDD.n61 VDD.n60 92.5005
R113 VDD.n60 VDD.t41 92.5005
R114 VDD.n327 VDD.n325 92.5005
R115 VDD.n285 VDD.t31 91.936
R116 VDD.t11 VDD.n225 87.4062
R117 VDD.t85 VDD.n247 85.9734
R118 VDD VDD.n207 85.9734
R119 VDD.n153 VDD.t53 84.5405
R120 VDD.n19 VDD.t61 81.7209
R121 VDD.n275 VDD.t43 81.7209
R122 VDD.t69 VDD 76.6134
R123 VDD.n291 VDD.t39 71.5059
R124 VDD.n187 VDD.t4 65.913
R125 VDD.n130 VDD.t0 63.0473
R126 VDD.t2 VDD.n112 63.0473
R127 VDD.n97 VDD.t100 63.0473
R128 VDD.n154 VDD.t98 61.6144
R129 VDD.n23 VDD.t67 61.2908
R130 VDD.n271 VDD.t35 61.2908
R131 VDD.n130 VDD.t55 57.3157
R132 VDD.n112 VDD.t83 57.3157
R133 VDD.n236 VDD.t7 57.3157
R134 VDD.n193 VDD.t73 54.45
R135 VDD.n226 VDD.t89 51.5842
R136 VDD.n208 VDD.t79 51.5842
R137 VDD.n295 VDD.t23 51.0758
R138 VDD.n321 VDD.t27 51.0758
R139 VDD.t96 VDD.n236 45.8527
R140 VDD.n219 VDD.t77 45.8527
R141 VDD.t0 VDD 42.9869
R142 VDD VDD.t2 42.9869
R143 VDD VDD.t94 42.9869
R144 VDD.n187 VDD.t75 42.9869
R145 VDD.n226 VDD 41.554
R146 VDD.n208 VDD 41.554
R147 VDD.n37 VDD.t65 40.8607
R148 VDD.n73 VDD.t45 40.8607
R149 VDD.t57 VDD.t17 40.1212
R150 VDD.t87 VDD.t15 40.1212
R151 VDD.n198 VDD.t76 36.1587
R152 VDD.n198 VDD.t74 36.1587
R153 VDD.n212 VDD.t78 36.1587
R154 VDD.n212 VDD.t80 36.1587
R155 VDD.n230 VDD.t97 36.1587
R156 VDD.n230 VDD.t90 36.1587
R157 VDD.n95 VDD.t101 36.1587
R158 VDD.n95 VDD.t16 36.1587
R159 VDD.n107 VDD.t3 36.1587
R160 VDD.n107 VDD.t93 36.1587
R161 VDD.n124 VDD.t99 36.1587
R162 VDD.n124 VDD.t18 36.1587
R163 VDD.n126 VDD.t1 36.1587
R164 VDD.n126 VDD.t103 36.1587
R165 VDD.n185 VDD.t60 36.1587
R166 VDD.n185 VDD.t5 36.1587
R167 VDD.t98 VDD.t51 34.3896
R168 VDD.t100 VDD.t81 34.3896
R169 VDD.n225 VDD.t9 32.9568
R170 VDD.n301 VDD.t19 30.6457
R171 VDD.n317 VDD.t49 30.6457
R172 VDD.n237 VDD 28.6581
R173 VDD.n127 VDD.t91 26.5955
R174 VDD.n127 VDD.t56 26.5955
R175 VDD.n148 VDD.t54 26.5955
R176 VDD.n148 VDD.t52 26.5955
R177 VDD.n108 VDD.t6 26.5955
R178 VDD.n108 VDD.t84 26.5955
R179 VDD.n93 VDD.t86 26.5955
R180 VDD.n93 VDD.t82 26.5955
R181 VDD.n174 VDD.t95 26.5955
R182 VDD.n174 VDD.t8 26.5955
R183 VDD.n179 VDD.t12 26.5955
R184 VDD.n179 VDD.t10 26.5955
R185 VDD.n315 VDD.t50 26.5955
R186 VDD.n315 VDD.t28 26.5955
R187 VDD.n309 VDD.t30 26.5955
R188 VDD.n309 VDD.t34 26.5955
R189 VDD.n299 VDD.t24 26.5955
R190 VDD.n299 VDD.t20 26.5955
R191 VDD.n289 VDD.t32 26.5955
R192 VDD.n289 VDD.t40 26.5955
R193 VDD.n279 VDD.t38 26.5955
R194 VDD.n279 VDD.t22 26.5955
R195 VDD.n269 VDD.t36 26.5955
R196 VDD.n269 VDD.t44 26.5955
R197 VDD.n64 VDD.t26 26.5955
R198 VDD.n64 VDD.t46 26.5955
R199 VDD.n58 VDD.t72 26.5955
R200 VDD.n58 VDD.t42 26.5955
R201 VDD.n35 VDD.t68 26.5955
R202 VDD.n35 VDD.t66 26.5955
R203 VDD.n17 VDD.t64 26.5955
R204 VDD.n17 VDD.t62 26.5955
R205 VDD VDD.n153 25.7924
R206 VDD VDD.n147 24.3595
R207 VDD.n154 VDD.t57 24.3595
R208 VDD.n113 VDD 24.3595
R209 VDD.n248 VDD 24.3595
R210 VDD.n247 VDD 24.3595
R211 VDD.n97 VDD.t87 22.9266
R212 VDD.n219 VDD.t13 22.9266
R213 VDD.t53 VDD 21.4937
R214 VDD VDD.t85 21.4937
R215 VDD.n193 VDD 21.4937
R216 VDD.n45 VDD.t71 20.4306
R217 VDD.n66 VDD.t25 20.4306
R218 VDD.t94 VDD.t96 17.1951
R219 VDD.t75 VDD.t59 17.1951
R220 VDD.n3 VDD.n2 14.6556
R221 VDD.n305 VDD.t29 10.2156
R222 VDD.n311 VDD.t33 10.2156
R223 VDD.t51 VDD 10.0307
R224 VDD.t81 VDD 10.0307
R225 VDD.n245 VDD.n99 9.05896
R226 VDD.n313 VDD.n310 8.53383
R227 VDD.n222 VDD.n221 7.87742
R228 VDD.n61 VDD.n59 7.7918
R229 VDD.n240 VDD.n239 7.6805
R230 VDD.n190 VDD.n189 7.6805
R231 VDD.n205 VDD.n184 7.58204
R232 VDD.n132 VDD 7.28665
R233 VDD.n110 VDD 7.28665
R234 VDD.n234 VDD 7.28665
R235 VDD.n68 VDD.n65 6.30775
R236 VDD.n181 VDD.n180 6.10512
R237 VDD.n2 VDD 5.78698
R238 VDD.t55 VDD.t102 5.73202
R239 VDD.t83 VDD.t92 5.73202
R240 VDD.n99 VDD.n96 5.71127
R241 VDD.n303 VDD.n300 5.56572
R242 VDD.n319 VDD.n316 5.56572
R243 VDD.n192 VDD.n191 4.6505
R244 VDD.n176 VDD.n172 4.6505
R245 VDD.n234 VDD.n233 4.6505
R246 VDD.n229 VDD.n228 4.6505
R247 VDD.n218 VDD.n217 4.6505
R248 VDD.n211 VDD.n210 4.6505
R249 VDD.n204 VDD.n203 4.6505
R250 VDD.n197 VDD.n196 4.6505
R251 VDD.n232 VDD.n231 4.6505
R252 VDD.n214 VDD.n213 4.6505
R253 VDD.n200 VDD.n199 4.6505
R254 VDD.n184 VDD.n182 4.6505
R255 VDD.n180 VDD.n178 4.6505
R256 VDD.n328 VDD.n327 4.6505
R257 VDD.n69 VDD.n68 4.6505
R258 VDD.n48 VDD.n47 4.6505
R259 VDD.n22 VDD.n21 4.6505
R260 VDD.n26 VDD.n25 4.6505
R261 VDD.n274 VDD.n273 4.6505
R262 VDD.n278 VDD.n277 4.6505
R263 VDD.n284 VDD.n283 4.6505
R264 VDD.n288 VDD.n287 4.6505
R265 VDD.n294 VDD.n293 4.6505
R266 VDD.n298 VDD.n297 4.6505
R267 VDD.n304 VDD.n303 4.6505
R268 VDD.n308 VDD.n307 4.6505
R269 VDD.n314 VDD.n313 4.6505
R270 VDD.n320 VDD.n319 4.6505
R271 VDD.n324 VDD.n323 4.6505
R272 VDD.n8 VDD.n7 4.5005
R273 VDD.n42 VDD.n41 4.5005
R274 VDD.n77 VDD.n76 4.5005
R275 VDD VDD.t11 4.29914
R276 VDD.n41 VDD.n36 3.52514
R277 VDD.n122 VDD.n119 3.34819
R278 VDD.n210 VDD.n183 3.34819
R279 VDD.n273 VDD.n270 3.33963
R280 VDD.n62 VDD.n61 3.03311
R281 VDD.n75 VDD.n72 2.96862
R282 VDD.n133 VDD.n125 2.8777
R283 VDD.n293 VDD.n290 2.5976
R284 VDD.n327 VDD.n326 2.5976
R285 VDD.n133 VDD.n132 2.3255
R286 VDD.n158 VDD.n157 2.3255
R287 VDD.n110 VDD.n92 2.3255
R288 VDD.n242 VDD.n99 2.3255
R289 VDD.n241 VDD.n240 2.3255
R290 VDD.n245 VDD.n244 2.3255
R291 VDD.n251 VDD.n250 2.3255
R292 VDD.n117 VDD.n116 2.3255
R293 VDD.n123 VDD.n122 2.3255
R294 VDD.n150 VDD.n102 2.3255
R295 VDD.n145 VDD.n144 2.3255
R296 VDD.n118 VDD.n106 1.94045
R297 VDD.n143 VDD.n142 1.94045
R298 VDD.n160 VDD.n159 1.94045
R299 VDD.n243 VDD.n168 1.94045
R300 VDD.n253 VDD.n252 1.94045
R301 VDD.n7 VDD.n6 1.85557
R302 VDD.n21 VDD.n18 1.85557
R303 VDD.n40 VDD.n39 1.85557
R304 VDD.n245 VDD.n94 1.77281
R305 VDD.n218 VDD.n181 1.77281
R306 VDD.n255 VDD.n254 1.7089
R307 VDD.n167 VDD.n164 1.7089
R308 VDD.n104 VDD.n89 1.70599
R309 VDD.n140 VDD.n139 1.70599
R310 VDD.n163 VDD.n162 1.70599
R311 VDD.n265 VDD.n263 1.70599
R312 VDD.n151 VDD.n149 1.67435
R313 VDD.n115 VDD 1.67435
R314 VDD.n15 VDD.n14 1.35607
R315 VDD.n267 VDD.n266 1.35607
R316 VDD.n34 VDD.n33 1.35607
R317 VDD.n57 VDD.n56 1.35607
R318 VDD.n6 VDD.n3 1.29905
R319 VDD.n41 VDD.n40 1.29905
R320 VDD VDD.n125 1.2805
R321 VDD.n173 VDD.n172 1.18204
R322 VDD.n204 VDD.n190 1.18204
R323 VDD.n223 VDD.n222 1.08358
R324 VDD.n14 VDD.n12 0.853
R325 VDD.n266 VDD.n265 0.853
R326 VDD.n33 VDD.n32 0.853
R327 VDD.n56 VDD.n55 0.853
R328 VDD.n168 VDD.n167 0.685162
R329 VDD.n254 VDD.n253 0.685162
R330 VDD.n161 VDD.n160 0.682811
R331 VDD.n142 VDD.n141 0.682811
R332 VDD.n106 VDD.n105 0.682811
R333 VDD VDD.n173 0.591269
R334 VDD.n132 VDD.n128 0.492808
R335 VDD.n110 VDD.n109 0.492808
R336 VDD.n234 VDD.n175 0.492808
R337 VDD.n191 VDD 0.492808
R338 VDD.n283 VDD.n280 0.371515
R339 VDD.n205 VDD.n204 0.295885
R340 VDD.n239 VDD.n172 0.197423
R341 VDD.n189 VDD.n186 0.197423
R342 VDD.n196 VDD.n195 0.197423
R343 VDD.n76 VDD.n75 0.186007
R344 VDD.n26 VDD.n22 0.120292
R345 VDD.n278 VDD.n274 0.120292
R346 VDD.n284 VDD.n278 0.120292
R347 VDD.n288 VDD.n284 0.120292
R348 VDD.n294 VDD.n288 0.120292
R349 VDD.n298 VDD.n294 0.120292
R350 VDD.n304 VDD.n298 0.120292
R351 VDD.n308 VDD.n304 0.120292
R352 VDD.n314 VDD.n308 0.120292
R353 VDD.n320 VDD.n314 0.120292
R354 VDD.n324 VDD.n320 0.120292
R355 VDD.n328 VDD.n324 0.120292
R356 VDD.n329 VDD.n328 0.120292
R357 VDD.n48 VDD.n44 0.107271
R358 VDD.n70 VDD.n69 0.0994583
R359 VDD.n151 VDD.n150 0.0989615
R360 VDD.n157 VDD.n156 0.0989615
R361 VDD.n116 VDD.n115 0.0989615
R362 VDD.n240 VDD.n171 0.0989615
R363 VDD.n223 VDD.n218 0.0989615
R364 VDD.n69 VDD.n63 0.0968542
R365 VDD VDD.n1 0.0877396
R366 VDD.n49 VDD.n48 0.0877396
R367 VDD.n274 VDD.n268 0.0851354
R368 VDD.n27 VDD.n26 0.0773229
R369 VDD.n22 VDD.n16 0.0734167
R370 VDD.n158 VDD.n123 0.0603958
R371 VDD.n117 VDD.n92 0.0603958
R372 VDD.n242 VDD.n241 0.0603958
R373 VDD VDD.n329 0.0603958
R374 VDD.n259 VDD.n258 0.0573462
R375 VDD.n144 VDD.n143 0.0564896
R376 VDD.n252 VDD.n251 0.0525833
R377 VDD.n233 VDD.n177 0.0525833
R378 VDD.n232 VDD.n229 0.0525833
R379 VDD.n216 VDD.n215 0.0525833
R380 VDD.n214 VDD.n211 0.0525833
R381 VDD.n202 VDD.n201 0.0525833
R382 VDD.n200 VDD.n197 0.0525833
R383 VDD VDD.n158 0.0493281
R384 VDD VDD.n242 0.0493281
R385 VDD.n14 VDD.n9 0.0429107
R386 VDD.n56 VDD.n50 0.0406786
R387 VDD.n52 VDD.n51 0.0406786
R388 VDD.n266 VDD.n79 0.0384464
R389 VDD.n33 VDD.n29 0.0362143
R390 VDD VDD.n102 0.0304479
R391 VDD VDD.n117 0.0304479
R392 VDD.n244 VDD 0.0304479
R393 VDD.n241 VDD 0.0304479
R394 VDD.n136 VDD 0.0302812
R395 VDD.n118 VDD 0.0265417
R396 VDD.n15 VDD.n8 0.0252396
R397 VDD.n57 VDD.n49 0.0239375
R398 VDD.n63 VDD.n62 0.0239375
R399 VDD.n33 VDD.n28 0.0228214
R400 VDD.n176 VDD 0.0226354
R401 VDD.n217 VDD 0.0226354
R402 VDD.n203 VDD 0.0226354
R403 VDD.n268 VDD.n267 0.0226354
R404 VDD.n42 VDD.n34 0.0213333
R405 VDD.n71 VDD.n70 0.0213333
R406 VDD.n266 VDD.n78 0.0205893
R407 VDD.n166 VDD.n165 0.0167692
R408 VDD.n162 VDD.n101 0.0167692
R409 VDD.n140 VDD.n134 0.0167692
R410 VDD.n104 VDD.n103 0.0167692
R411 VDD.n91 VDD.n90 0.0167692
R412 VDD.n32 VDD.n31 0.0167692
R413 VDD.n12 VDD.n10 0.0167692
R414 VDD.n12 VDD.n11 0.0167692
R415 VDD.n55 VDD.n54 0.0167692
R416 VDD.n265 VDD.n80 0.0167692
R417 VDD.n265 VDD.n264 0.0167692
R418 VDD.n14 VDD.n13 0.016125
R419 VDD.n56 VDD.n52 0.016125
R420 VDD.n8 VDD.n0 0.0135208
R421 VDD.n34 VDD.n27 0.0135208
R422 VDD.n44 VDD.n43 0.0135208
R423 VDD.n267 VDD.n77 0.0122188
R424 VDD.n144 VDD 0.0115677
R425 VDD.n251 VDD 0.0115677
R426 VDD VDD.n178 0.0115677
R427 VDD VDD.n182 0.0115677
R428 VDD.n192 VDD 0.0115677
R429 VDD.n1 VDD.n0 0.00961458
R430 VDD.n16 VDD.n15 0.00961458
R431 VDD.n43 VDD.n42 0.00961458
R432 VDD.n62 VDD.n57 0.00961458
R433 VDD.n32 VDD.n30 0.00911311
R434 VDD.n55 VDD.n53 0.00911311
R435 VDD.n244 VDD.n243 0.00896354
R436 VDD.n252 VDD.n92 0.0083125
R437 VDD.n177 VDD.n176 0.0083125
R438 VDD.n233 VDD.n232 0.0083125
R439 VDD.n229 VDD.n178 0.0083125
R440 VDD.n217 VDD.n216 0.0083125
R441 VDD.n215 VDD.n214 0.0083125
R442 VDD.n211 VDD.n182 0.0083125
R443 VDD.n203 VDD.n202 0.0083125
R444 VDD.n201 VDD.n200 0.0083125
R445 VDD.n197 VDD.n192 0.0083125
R446 VDD.n159 VDD 0.00766146
R447 VDD.n143 VDD.n133 0.00440625
R448 VDD.n159 VDD.n102 0.00440625
R449 VDD.n123 VDD.n118 0.00440625
R450 VDD.n162 VDD.n161 0.00419645
R451 VDD.n141 VDD.n140 0.00419645
R452 VDD.n105 VDD.n104 0.00419645
R453 VDD.n243 VDD 0.00310417
R454 VDD.n167 VDD.n166 0.00284309
R455 VDD.n254 VDD.n91 0.00284309
R456 VDD.n263 VDD.n262 0.00228535
R457 VDD.n139 VDD.n138 0.00228535
R458 VDD.n77 VDD.n71 0.00180208
R459 VDD.n84 VDD.n83 0.00171259
R460 VDD.n256 VDD.n255 0.00171259
R461 VDD.n87 VDD.n86 0.00107275
R462 VDD.n86 VDD.n85 0.00102425
R463 VDD.n263 VDD.n88 0.00102425
R464 VDD.n255 VDD.n89 0.00102425
R465 VDD.n164 VDD.n163 0.00102425
R466 VDD.n139 VDD.n135 0.00102425
R467 VDD.n164 VDD.n89 0.00102425
R468 VDD.n163 VDD.n100 0.00102425
R469 VDD.n257 VDD.n256 0.000645511
R470 VDD.n137 VDD.n136 0.000645511
R471 VDD.n82 VDD.n81 0.000597007
R472 VDD.n261 VDD.n260 0.000597007
R473 VDD.n135 VDD.n100 0.000597007
R474 VDD.n83 VDD.n82 0.000548504
R475 VDD.n85 VDD.n84 0.000548504
R476 VDD.n88 VDD.n87 0.000548504
R477 VDD.n262 VDD.n261 0.000548504
R478 VDD.n260 VDD.n259 0.000548504
R479 VDD.n258 VDD.n257 0.000548504
R480 VDD.n138 VDD.n137 0.000548504
R481 sw<6>.n2 sw<6>.n0 146.811
R482 sw<6>.n14 sw<6>.n13 108.412
R483 sw<6>.n2 sw<6>.n1 108.412
R484 sw<6>.n4 sw<6>.n3 108.412
R485 sw<6>.n6 sw<6>.n5 108.412
R486 sw<6>.n8 sw<6>.n7 108.412
R487 sw<6>.n10 sw<6>.n9 108.412
R488 sw<6>.n12 sw<6>.n11 108.412
R489 sw<6>.n17 sw<6>.n15 90.8321
R490 sw<6>.n17 sw<6>.n16 52.4321
R491 sw<6>.n19 sw<6>.n18 52.4321
R492 sw<6>.n21 sw<6>.n20 52.4321
R493 sw<6>.n23 sw<6>.n22 52.4321
R494 sw<6>.n25 sw<6>.n24 52.4321
R495 sw<6>.n27 sw<6>.n26 52.4321
R496 sw<6>.n29 sw<6>.n28 52.4321
R497 sw<6> sw<6>.n29 40.4711
R498 sw<6>.n4 sw<6>.n2 38.4005
R499 sw<6>.n6 sw<6>.n4 38.4005
R500 sw<6>.n8 sw<6>.n6 38.4005
R501 sw<6>.n10 sw<6>.n8 38.4005
R502 sw<6>.n12 sw<6>.n10 38.4005
R503 sw<6>.n14 sw<6>.n12 38.4005
R504 sw<6>.n19 sw<6>.n17 38.4005
R505 sw<6>.n21 sw<6>.n19 38.4005
R506 sw<6>.n23 sw<6>.n21 38.4005
R507 sw<6>.n25 sw<6>.n23 38.4005
R508 sw<6>.n27 sw<6>.n25 38.4005
R509 sw<6>.n29 sw<6>.n27 38.4005
R510 sw<6> sw<6>.n14 33.7342
R511 sw<6>.n0 sw<6>.t21 26.5955
R512 sw<6>.n0 sw<6>.t13 26.5955
R513 sw<6>.n1 sw<6>.t23 26.5955
R514 sw<6>.n1 sw<6>.t18 26.5955
R515 sw<6>.n3 sw<6>.t22 26.5955
R516 sw<6>.n3 sw<6>.t19 26.5955
R517 sw<6>.n5 sw<6>.t11 26.5955
R518 sw<6>.n5 sw<6>.t16 26.5955
R519 sw<6>.n7 sw<6>.t20 26.5955
R520 sw<6>.n7 sw<6>.t12 26.5955
R521 sw<6>.n9 sw<6>.t10 26.5955
R522 sw<6>.n9 sw<6>.t15 26.5955
R523 sw<6>.n11 sw<6>.t17 26.5955
R524 sw<6>.n11 sw<6>.t25 26.5955
R525 sw<6>.n13 sw<6>.t14 26.5955
R526 sw<6>.n13 sw<6>.t24 26.5955
R527 sw<6>.n15 sw<6>.t5 24.9236
R528 sw<6>.n15 sw<6>.t9 24.9236
R529 sw<6>.n16 sw<6>.t2 24.9236
R530 sw<6>.n16 sw<6>.t31 24.9236
R531 sw<6>.n18 sw<6>.t1 24.9236
R532 sw<6>.n18 sw<6>.t0 24.9236
R533 sw<6>.n20 sw<6>.t6 24.9236
R534 sw<6>.n20 sw<6>.t7 24.9236
R535 sw<6>.n22 sw<6>.t28 24.9236
R536 sw<6>.n22 sw<6>.t4 24.9236
R537 sw<6>.n24 sw<6>.t26 24.9236
R538 sw<6>.n24 sw<6>.t29 24.9236
R539 sw<6>.n26 sw<6>.t3 24.9236
R540 sw<6>.n26 sw<6>.t8 24.9236
R541 sw<6>.n28 sw<6>.t27 24.9236
R542 sw<6>.n28 sw<6>.t30 24.9236
R543 sw<6>.n30 sw<6> 8.08471
R544 sw<6> sw<6>.n30 3.83425
R545 sw<6>.n30 sw<6> 3.36892
R546 sw<5>.n5 sw<5>.n3 197.595
R547 sw<5> sw<5>.n4 165.219
R548 sw<5>.n2 sw<5>.n0 138.054
R549 sw<5>.n2 sw<5>.n1 107.874
R550 sw<5>.n3 sw<5>.t5 26.5955
R551 sw<5>.n3 sw<5>.t6 26.5955
R552 sw<5>.n4 sw<5>.t4 26.5955
R553 sw<5>.n4 sw<5>.t7 26.5955
R554 sw<5>.n0 sw<5>.t2 24.9236
R555 sw<5>.n0 sw<5>.t0 24.9236
R556 sw<5>.n1 sw<5>.t1 24.9236
R557 sw<5>.n1 sw<5>.t3 24.9236
R558 sw<5>.n6 sw<5> 6.98232
R559 sw<5> sw<5>.n5 6.59444
R560 sw<5> sw<5>.n6 3.83425
R561 sw<5> sw<5>.n2 2.97424
R562 sw<5>.n5 sw<5> 2.19848
R563 sw<5>.n6 sw<5> 1.8106
R564 VSS.n198 VSS 896.297
R565 VSS.n225 VSS 896.297
R566 VSS.n257 VSS 896.297
R567 VSS VSS.n265 896.297
R568 VSS.n187 VSS.t2 711.548
R569 VSS.n184 VSS.t81 512.169
R570 VSS.n199 VSS.t74 512.169
R571 VSS.n199 VSS.t20 512.169
R572 VSS.n212 VSS.t4 512.169
R573 VSS.n212 VSS.t94 512.169
R574 VSS.n226 VSS.t71 512.169
R575 VSS.n226 VSS.t18 512.169
R576 VSS.n249 VSS.t97 512.169
R577 VSS.n249 VSS.t6 512.169
R578 VSS.n274 VSS.t79 512.169
R579 VSS.n274 VSS.t83 512.169
R580 VSS.n291 VSS.t68 512.169
R581 VSS.n291 VSS.t0 512.169
R582 VSS.n43 VSS.n41 495.315
R583 VSS VSS.n41 413.536
R584 VSS.t74 VSS 337.567
R585 VSS.t71 VSS 337.567
R586 VSS.n101 VSS.t35 313.269
R587 VSS.n42 VSS.t54 306.149
R588 VSS.n188 VSS.n187 296.384
R589 VSS.n238 VSS.n237 292.5
R590 VSS.n237 VSS.n236 292.5
R591 VSS.n301 VSS.n300 292.5
R592 VSS.n302 VSS.n301 292.5
R593 VSS.n293 VSS.n292 292.5
R594 VSS.n292 VSS.n291 292.5
R595 VSS.n259 VSS.n258 292.5
R596 VSS.n258 VSS.n257 292.5
R597 VSS.n276 VSS.n275 292.5
R598 VSS.n275 VSS.n274 292.5
R599 VSS.n268 VSS.n267 292.5
R600 VSS.n267 VSS.n266 292.5
R601 VSS.n264 VSS.n263 292.5
R602 VSS.n265 VSS.n264 292.5
R603 VSS.n255 VSS.n254 292.5
R604 VSS.n256 VSS.n255 292.5
R605 VSS.n251 VSS.n250 292.5
R606 VSS.n250 VSS.n249 292.5
R607 VSS.n186 VSS.n185 292.5
R608 VSS.n185 VSS.n184 292.5
R609 VSS.n195 VSS.n194 292.5
R610 VSS.n196 VSS.n195 292.5
R611 VSS.n197 VSS.n182 292.5
R612 VSS.n198 VSS.n197 292.5
R613 VSS.n201 VSS.n200 292.5
R614 VSS.n200 VSS.n199 292.5
R615 VSS.n206 VSS.n205 292.5
R616 VSS.n205 VSS.n204 292.5
R617 VSS.n209 VSS.n208 292.5
R618 VSS.n208 VSS.n207 292.5
R619 VSS.n214 VSS.n213 292.5
R620 VSS.n213 VSS.n212 292.5
R621 VSS.n222 VSS.n221 292.5
R622 VSS.n223 VSS.n222 292.5
R623 VSS.n224 VSS.n180 292.5
R624 VSS.n225 VSS.n224 292.5
R625 VSS.n228 VSS.n227 292.5
R626 VSS.n227 VSS.n226 292.5
R627 VSS.n234 VSS.n233 292.5
R628 VSS.n233 VSS.n232 292.5
R629 VSS.n41 VSS.n40 292.5
R630 VSS.t44 VSS.n69 292.5
R631 VSS.n144 VSS.t24 292.5
R632 VSS.n145 VSS.n144 292.5
R633 VSS.n140 VSS.n139 292.5
R634 VSS.n139 VSS.n138 292.5
R635 VSS.n103 VSS.n102 292.5
R636 VSS.n102 VSS.n101 292.5
R637 VSS.n57 VSS.n56 292.5
R638 VSS.n56 VSS.n55 292.5
R639 VSS.n44 VSS.n43 292.5
R640 VSS.n43 VSS.n42 292.5
R641 VSS.n51 VSS.n50 292.5
R642 VSS.n50 VSS.n49 292.5
R643 VSS.n63 VSS.n62 292.5
R644 VSS.n62 VSS.n61 292.5
R645 VSS.n36 VSS.n35 292.5
R646 VSS.n35 VSS.n34 292.5
R647 VSS.n69 VSS.n68 292.5
R648 VSS.n72 VSS.n71 292.5
R649 VSS.n71 VSS.n70 292.5
R650 VSS.n76 VSS.n75 292.5
R651 VSS.n75 VSS.n74 292.5
R652 VSS.n85 VSS.n84 292.5
R653 VSS.n84 VSS.n83 292.5
R654 VSS.n89 VSS.n88 292.5
R655 VSS.n88 VSS.n87 292.5
R656 VSS.n95 VSS.n94 292.5
R657 VSS.n94 VSS.n93 292.5
R658 VSS.n99 VSS.n98 292.5
R659 VSS.n100 VSS.n99 292.5
R660 VSS.n14 VSS.n13 292.5
R661 VSS.n13 VSS.n12 292.5
R662 VSS.n125 VSS.n124 292.5
R663 VSS.n124 VSS.n123 292.5
R664 VSS.n131 VSS.n130 292.5
R665 VSS.n130 VSS.n129 292.5
R666 VSS.n154 VSS.n153 292.5
R667 VSS.n153 VSS.n152 292.5
R668 VSS.n305 VSS.n304 292.5
R669 VSS.n304 VSS.n303 292.5
R670 VSS.n42 VSS.t63 291.909
R671 VSS.n93 VSS.t42 291.909
R672 VSS.n70 VSS.t85 284.791
R673 VSS.n101 VSS.t10 284.791
R674 VSS.n100 VSS.t27 263.43
R675 VSS.n1 VSS.t99 260.322
R676 VSS.n189 VSS.t100 260.322
R677 VSS.n216 VSS.t101 260.322
R678 VSS.t30 VSS.t8 256.312
R679 VSS.t32 VSS.t58 256.312
R680 VSS.n74 VSS.t87 234.952
R681 VSS.n49 VSS.t50 227.833
R682 VSS.n87 VSS.t46 227.833
R683 VSS.t22 VSS.t77 227.833
R684 VSS VSS.n198 221.165
R685 VSS VSS.n225 221.165
R686 VSS.n12 VSS.t14 220.713
R687 VSS.t63 VSS 213.593
R688 VSS.t8 VSS 213.593
R689 VSS.t35 VSS 213.593
R690 VSS VSS.n302 197.885
R691 VSS.n308 VSS.t23 190.065
R692 VSS.n303 VSS 177.994
R693 VSS.n1 VSS.t76 175.169
R694 VSS.n189 VSS.t73 175.169
R695 VSS.n216 VSS.t70 175.169
R696 VSS VSS.n196 174.603
R697 VSS VSS.n223 174.603
R698 VSS VSS.n256 174.603
R699 VSS.n266 VSS 174.603
R700 VSS.n55 VSS.t56 170.875
R701 VSS.n83 VSS.t39 170.875
R702 VSS.n83 VSS.t91 170.875
R703 VSS.n123 VSS.t12 170.875
R704 VSS.n216 VSS 152.865
R705 VSS VSS.t44 128.155
R706 VSS VSS.n100 121.037
R707 VSS.n48 VSS.n47 116.219
R708 VSS.n60 VSS.n59 116.219
R709 VSS.n67 VSS.n32 116.219
R710 VSS.n31 VSS.n30 116.219
R711 VSS.n82 VSS.n81 116.219
R712 VSS.n96 VSS.n25 116.219
R713 VSS.n104 VSS.n24 116.219
R714 VSS.n122 VSS.n120 116.219
R715 VSS.n137 VSS.n136 116.219
R716 VSS.n148 VSS.n147 116.219
R717 VSS.n39 VSS.t64 114.775
R718 VSS.n61 VSS.t52 113.916
R719 VSS.n87 VSS.t89 113.916
R720 VSS.n105 VSS.n23 109.3
R721 VSS.n29 VSS.n28 109.3
R722 VSS.n38 VSS.n37 109.3
R723 VSS.n74 VSS.t48 106.796
R724 VSS.n122 VSS.n121 104.719
R725 VSS.n80 VSS.n79 104.719
R726 VSS.n54 VSS.n53 104.719
R727 VSS.n155 VSS.n151 103.942
R728 VSS.n228 VSS.n179 103.942
R729 VSS.n214 VSS.n211 103.942
R730 VSS.n201 VSS.n181 103.942
R731 VSS.n186 VSS.n183 103.942
R732 VSS.n251 VSS.n248 103.942
R733 VSS.n276 VSS.n272 103.942
R734 VSS.n293 VSS.n289 103.942
R735 VSS.n137 VSS.t17 100.21
R736 VSS.n26 VSS.t90 100.21
R737 VSS.n33 VSS.t53 100.21
R738 VSS.n129 VSS.t16 99.6769
R739 VSS.n34 VSS.t66 64.0782
R740 VSS.n70 VSS.t30 56.9584
R741 VSS.n138 VSS.t37 56.9584
R742 VSS.n152 VSS.t32 42.7189
R743 VSS.n303 VSS.t22 42.7189
R744 VSS.n151 VSS.t59 33.462
R745 VSS.n151 VSS.t78 33.462
R746 VSS.n179 VSS.t72 33.462
R747 VSS.n179 VSS.t19 33.462
R748 VSS.n211 VSS.t5 33.462
R749 VSS.n211 VSS.t95 33.462
R750 VSS.n181 VSS.t75 33.462
R751 VSS.n181 VSS.t21 33.462
R752 VSS.n183 VSS.t3 33.462
R753 VSS.n183 VSS.t82 33.462
R754 VSS.n248 VSS.t98 33.462
R755 VSS.n248 VSS.t7 33.462
R756 VSS.n272 VSS.t80 33.462
R757 VSS.n272 VSS.t84 33.462
R758 VSS.n289 VSS.t69 33.462
R759 VSS.n289 VSS.t1 33.462
R760 VSS.n308 VSS.n0 28.455
R761 VSS.n47 VSS.t62 24.9236
R762 VSS.n47 VSS.t60 24.9236
R763 VSS.n59 VSS.t65 24.9236
R764 VSS.n59 VSS.t61 24.9236
R765 VSS.n32 VSS.t67 24.9236
R766 VSS.n32 VSS.t45 24.9236
R767 VSS.n30 VSS.t31 24.9236
R768 VSS.n30 VSS.t49 24.9236
R769 VSS.n81 VSS.t40 24.9236
R770 VSS.n81 VSS.t47 24.9236
R771 VSS.n25 VSS.t43 24.9236
R772 VSS.n25 VSS.t28 24.9236
R773 VSS.n24 VSS.t36 24.9236
R774 VSS.n24 VSS.t41 24.9236
R775 VSS.n121 VSS.t15 24.9236
R776 VSS.n121 VSS.t13 24.9236
R777 VSS.n120 VSS.t29 24.9236
R778 VSS.n120 VSS.t26 24.9236
R779 VSS.n136 VSS.t34 24.9236
R780 VSS.n136 VSS.t38 24.9236
R781 VSS.n147 VSS.t25 24.9236
R782 VSS.n147 VSS.t33 24.9236
R783 VSS.n23 VSS.t96 24.9236
R784 VSS.n23 VSS.t11 24.9236
R785 VSS.n79 VSS.t88 24.9236
R786 VSS.n79 VSS.t92 24.9236
R787 VSS.n28 VSS.t9 24.9236
R788 VSS.n28 VSS.t86 24.9236
R789 VSS.n53 VSS.t51 24.9236
R790 VSS.n53 VSS.t57 24.9236
R791 VSS.n37 VSS.t93 24.9236
R792 VSS.n37 VSS.t55 24.9236
R793 VSS.n194 VSS.n182 16.8234
R794 VSS.n201 VSS.n182 16.8234
R795 VSS.n209 VSS.n206 16.8234
R796 VSS.n221 VSS.n180 16.8234
R797 VSS.n228 VSS.n180 16.8234
R798 VSS.n235 VSS.n234 16.6405
R799 VSS.n2 VSS.n1 9.28751
R800 VSS.n217 VSS.n216 8.73669
R801 VSS.n190 VSS.n189 8.16166
R802 VSS.n145 VSS.n143 7.87742
R803 VSS.n97 VSS.n96 7.6805
R804 VSS VSS.n38 6.4005
R805 VSS VSS.n29 6.4005
R806 VSS VSS.n105 6.4005
R807 VSS.n67 VSS.n66 4.92358
R808 VSS.n234 VSS.n231 4.6505
R809 VSS.n229 VSS.n228 4.6505
R810 VSS.n219 VSS.n180 4.6505
R811 VSS.n221 VSS.n220 4.6505
R812 VSS.n215 VSS.n214 4.6505
R813 VSS.n210 VSS.n209 4.6505
R814 VSS.n202 VSS.n201 4.6505
R815 VSS.n254 VSS.n253 4.6505
R816 VSS.n263 VSS.n262 4.6505
R817 VSS.n269 VSS.n268 4.6505
R818 VSS.n299 VSS.n298 4.6505
R819 VSS.n260 VSS.n259 4.6505
R820 VSS.n252 VSS.n251 4.6505
R821 VSS.n206 VSS.n203 4.6505
R822 VSS.n192 VSS.n182 4.6505
R823 VSS.n194 VSS.n193 4.6505
R824 VSS.n156 VSS.n155 4.6505
R825 VSS.n307 VSS.n306 4.6505
R826 VSS.n146 VSS.n145 4.6505
R827 VSS.n141 VSS.n140 4.6505
R828 VSS.n133 VSS.n132 4.6505
R829 VSS.n126 VSS.n125 4.6505
R830 VSS.n16 VSS.n15 4.6505
R831 VSS.n103 VSS.n22 4.6505
R832 VSS.n97 VSS.n21 4.6505
R833 VSS.n107 VSS.n106 4.6505
R834 VSS.n11 VSS.n10 4.6505
R835 VSS.n119 VSS.n118 4.6505
R836 VSS.n128 VSS.n127 4.6505
R837 VSS.n135 VSS.n134 4.6505
R838 VSS.n150 VSS.n149 4.6505
R839 VSS.n158 VSS.n157 4.6505
R840 VSS.n310 VSS.n309 4.6505
R841 VSS.n240 VSS.n239 4.5005
R842 VSS.n295 VSS.n294 4.5005
R843 VSS.n278 VSS.n277 4.5005
R844 VSS.n68 VSS.n67 4.13588
R845 VSS.n191 VSS.n190 4.07975
R846 VSS.n218 VSS.n217 3.97187
R847 VSS.n72 VSS.n31 3.34819
R848 VSS.n92 VSS.n26 3.34819
R849 VSS.n140 VSS.n137 3.34819
R850 VSS.n36 VSS.n33 3.24973
R851 VSS.n3 VSS.n2 2.95474
R852 VSS.n149 VSS.n148 2.95435
R853 VSS.n239 VSS.n238 2.92621
R854 VSS.n294 VSS.n293 2.74336
R855 VSS.n299 VSS 2.74336
R856 VSS.n188 VSS.n186 2.59307
R857 VSS.n63 VSS.n60 2.5605
R858 VSS.n40 VSS 2.43568
R859 VSS.n2 VSS 2.37344
R860 VSS.n46 VSS.n45 2.3255
R861 VSS.n52 VSS.n51 2.3255
R862 VSS.n58 VSS.n57 2.3255
R863 VSS.n64 VSS.n63 2.3255
R864 VSS.n66 VSS.n65 2.3255
R865 VSS.n68 VSS.n27 2.3255
R866 VSS.n73 VSS.n72 2.3255
R867 VSS.n78 VSS.n77 2.3255
R868 VSS.n86 VSS.n85 2.3255
R869 VSS.n90 VSS.n89 2.3255
R870 VSS.n92 VSS.n91 2.3255
R871 VSS.n217 VSS 2.04519
R872 VSS.n276 VSS.n273 2.01193
R873 VSS.n119 VSS.n117 1.94045
R874 VSS.n109 VSS.n108 1.94045
R875 VSS.n160 VSS.n159 1.94045
R876 VSS.n190 VSS 1.91099
R877 VSS.n57 VSS.n54 1.77281
R878 VSS.n68 VSS 1.77281
R879 VSS.n85 VSS.n80 1.77281
R880 VSS.n85 VSS.n82 1.77281
R881 VSS.n125 VSS.n122 1.77281
R882 VSS.n116 VSS.n113 1.7089
R883 VSS.n112 VSS.n110 1.7089
R884 VSS.n286 VSS.n284 1.70599
R885 VSS.n282 VSS.n281 1.70599
R886 VSS.n163 VSS.n162 1.70599
R887 VSS.n283 VSS.n170 1.70239
R888 VSS.n288 VSS.n287 1.35607
R889 VSS.n280 VSS.n279 1.35607
R890 VSS.n246 VSS.n245 1.35607
R891 VSS.n193 VSS.n188 1.35477
R892 VSS.n39 VSS 1.18204
R893 VSS.n277 VSS.n276 1.09764
R894 VSS VSS.n308 1.08358
R895 VSS.n51 VSS.n48 0.985115
R896 VSS.n306 VSS.n305 0.985115
R897 VSS.n72 VSS.n29 0.886654
R898 VSS.n281 VSS.n280 0.853
R899 VSS.n287 VSS.n286 0.853
R900 VSS.n245 VSS.n244 0.853
R901 VSS.n105 VSS.n104 0.689731
R902 VSS.n110 VSS.n109 0.685162
R903 VSS.n117 VSS.n116 0.685162
R904 VSS.n161 VSS.n160 0.682811
R905 VSS.n44 VSS.n38 0.591269
R906 VSS.n106 VSS 0.591269
R907 VSS.n40 VSS.n39 0.492808
R908 VSS.n293 VSS.n290 0.366214
R909 VSS.n300 VSS.n299 0.366214
R910 VSS.n45 VSS.n44 0.295885
R911 VSS.n309 VSS 0.295885
R912 VSS.n104 VSS.n103 0.197423
R913 VSS.n132 VSS.n131 0.197423
R914 VSS.n155 VSS.n154 0.197423
R915 VSS.n238 VSS.n235 0.183357
R916 VSS.n203 VSS.n202 0.120292
R917 VSS.n215 VSS.n210 0.120292
R918 VSS.n220 VSS.n215 0.120292
R919 VSS.n231 VSS.n229 0.120292
R920 VSS.n253 VSS.n252 0.120292
R921 VSS.n298 VSS.n297 0.117688
R922 VSS.n270 VSS.n269 0.105969
R923 VSS.n66 VSS.n36 0.0989615
R924 VSS.n77 VSS.n76 0.0989615
R925 VSS.n95 VSS.n92 0.0989615
R926 VSS.n96 VSS.n95 0.0989615
R927 VSS.n98 VSS.n97 0.0989615
R928 VSS.n15 VSS.n14 0.0989615
R929 VSS.n202 VSS 0.0955521
R930 VSS.n229 VSS 0.0955521
R931 VSS.n261 VSS.n260 0.078625
R932 VSS VSS.n0 0.0760208
R933 VSS.n262 VSS.n4 0.0669062
R934 VSS.n252 VSS.n247 0.0656042
R935 VSS VSS.n192 0.0603958
R936 VSS.n203 VSS 0.0603958
R937 VSS.n210 VSS 0.0603958
R938 VSS VSS.n219 0.0603958
R939 VSS.n231 VSS 0.0603958
R940 VSS.n260 VSS 0.0603958
R941 VSS.n262 VSS 0.0603958
R942 VSS.n298 VSS 0.0603958
R943 VSS.n0 VSS 0.0603958
R944 VSS.n52 VSS.n46 0.0603958
R945 VSS.n58 VSS.n52 0.0603958
R946 VSS.n64 VSS.n58 0.0603958
R947 VSS.n65 VSS.n64 0.0603958
R948 VSS.n73 VSS.n27 0.0603958
R949 VSS.n78 VSS.n73 0.0603958
R950 VSS.n86 VSS.n78 0.0603958
R951 VSS.n90 VSS.n86 0.0603958
R952 VSS.n91 VSS.n90 0.0603958
R953 VSS VSS.n230 0.0590938
R954 VSS.n167 VSS.n166 0.0567656
R955 VSS.n245 VSS.n241 0.0563036
R956 VSS.n287 VSS.n6 0.0540714
R957 VSS.n107 VSS.n22 0.0525833
R958 VSS.n16 VSS.n11 0.0525833
R959 VSS.n126 VSS.n119 0.0525833
R960 VSS.n133 VSS.n128 0.0525833
R961 VSS.n141 VSS.n135 0.0525833
R962 VSS.n156 VSS.n150 0.0525833
R963 VSS.n46 VSS 0.0486771
R964 VSS.n280 VSS.n177 0.0362143
R965 VSS.n246 VSS.n240 0.0330521
R966 VSS.n295 VSS.n288 0.03175
R967 VSS.n65 VSS 0.0304479
R968 VSS VSS.n27 0.0304479
R969 VSS.n91 VSS 0.0304479
R970 VSS.n146 VSS 0.0304479
R971 VSS.n159 VSS.n3 0.0297969
R972 VSS.n280 VSS.n176 0.0228214
R973 VSS VSS.n21 0.0226354
R974 VSS VSS.n142 0.0226354
R975 VSS VSS.n310 0.0226354
R976 VSS.n159 VSS.n158 0.0219844
R977 VSS.n191 VSS 0.0213333
R978 VSS.n218 VSS 0.0213333
R979 VSS.n240 VSS.n178 0.0213333
R980 VSS.n279 VSS.n278 0.0213333
R981 VSS.n193 VSS 0.0200312
R982 VSS.n220 VSS 0.0200312
R983 VSS.n253 VSS 0.0200312
R984 VSS.n269 VSS 0.0200312
R985 VSS.n296 VSS.n295 0.0200312
R986 VSS.n20 VSS.n19 0.0167692
R987 VSS.n115 VSS.n114 0.0167692
R988 VSS.n281 VSS.n174 0.0167692
R989 VSS.n281 VSS.n175 0.0167692
R990 VSS.n286 VSS.n7 0.0167692
R991 VSS.n286 VSS.n285 0.0167692
R992 VSS.n244 VSS.n243 0.0167692
R993 VSS.n162 VSS.n9 0.0167692
R994 VSS.n271 VSS.n270 0.0148229
R995 VSS.n279 VSS.n261 0.0135208
R996 VSS.n244 VSS.n170 0.00911311
R997 VSS.n278 VSS.n271 0.0083125
R998 VSS.n119 VSS.n16 0.0083125
R999 VSS.n128 VSS.n126 0.0083125
R1000 VSS.n135 VSS.n133 0.0083125
R1001 VSS.n142 VSS.n141 0.0083125
R1002 VSS.n150 VSS.n146 0.0083125
R1003 VSS.n158 VSS.n156 0.0083125
R1004 VSS.n310 VSS.n307 0.0083125
R1005 VSS.n108 VSS.n21 0.00701042
R1006 VSS.n287 VSS.n5 0.00496429
R1007 VSS.n192 VSS.n191 0.00440625
R1008 VSS.n219 VSS.n218 0.00440625
R1009 VSS.n162 VSS.n161 0.00419645
R1010 VSS.n288 VSS.n4 0.00310417
R1011 VSS.n297 VSS.n296 0.00310417
R1012 VSS.n110 VSS.n20 0.00284309
R1013 VSS.n116 VSS.n115 0.00284309
R1014 VSS.n245 VSS.n242 0.00273214
R1015 VSS.n164 VSS.n163 0.00232022
R1016 VSS.n230 VSS.n178 0.00180208
R1017 VSS.n247 VSS.n246 0.00180208
R1018 VSS.n108 VSS.n107 0.00180208
R1019 VSS.n307 VSS.n3 0.00180208
R1020 VSS.n113 VSS.n18 0.00174821
R1021 VSS.n173 VSS.n172 0.00174821
R1022 VSS.n169 VSS.n168 0.0017002
R1023 VSS.n171 VSS 0.00131614
R1024 VSS.n284 VSS.n283 0.00116803
R1025 VSS.n163 VSS.n8 0.001024
R1026 VSS.n284 VSS.n169 0.001024
R1027 VSS.n283 VSS.n282 0.001024
R1028 VSS.n282 VSS.n173 0.001024
R1029 VSS.n168 VSS.n167 0.000692033
R1030 VSS.n172 VSS.n171 0.000692033
R1031 VSS.n18 VSS.n17 0.000596016
R1032 VSS.n166 VSS.n165 0.000596016
R1033 VSS.n113 VSS.n112 0.000548008
R1034 VSS.n112 VSS.n111 0.000548008
R1035 VSS.n111 VSS.n8 0.000548008
R1036 VSS.n165 VSS.n164 0.000548008
R1037 sar_val<7>.n2 sar_val<7>.t1 260.322
R1038 sar_val<7>.n2 sar_val<7>.t0 175.169
R1039 sar_val<7>.n3 sar_val<7>.n2 8.30068
R1040 sar_val<7>.n7 sar_val<7>.n5 4.5005
R1041 sar_val<7>.n5 sar_val<7>.n4 2.42212
R1042 sar_val<7>.n9 sar_val<7> 1.39782
R1043 sar_val<7>.n8 sar_val<7>.n7 1.11928
R1044 sar_val<7>.n4 sar_val<7> 0.865365
R1045 sar_val<7> sar_val<7>.n9 0.752904
R1046 sar_val<7>.n5 sar_val<7>.n3 0.519419
R1047 sar_val<7>.n9 sar_val<7>.n8 0.0643193
R1048 sar_val<7>.n7 sar_val<7>.n6 0.0278438
R1049 sar_val<7>.n8 sar_val<7>.n0 0.0141422
R1050 sar_val<7>.n7 sar_val<7>.n1 0.00635938
R1051 sw<2>.t1 sw<2> 459.913
R1052 sw<2>.n4 sw<2>.t1 141.43
R1053 sw<2>.n3 sw<2>.t0 123.654
R1054 sw<2> sw<2>.n3 78.8791
R1055 sw<2>.n5 sw<2>.n1 9.31706
R1056 sw<2>.n6 sw<2>.n5 9.3005
R1057 sw<2> sw<2>.n2 7.62451
R1058 sw<2>.n4 sw<2> 6.07224
R1059 sw<2>.n3 sw<2> 5.16973
R1060 sw<2>.n6 sw<2>.n0 4.53175
R1061 sw<2>.n8 sw<2>.n7 4.5005
R1062 sw<2>.n7 sw<2>.n2 2.48005
R1063 sw<2>.n5 sw<2>.n2 1.77056
R1064 sw<2>.n1 sw<2>.n0 1.12705
R1065 sw<2>.n5 sw<2>.n4 0.0681707
R1066 sw<2>.n8 sw<2>.n0 0.0509808
R1067 sw<2> sw<2>.n8 0.0125192
R1068 sw<2>.n7 sw<2>.n6 0.0122188
R1069 sw<2>.n7 sw<2>.n1 0.00635287
R1070 sar_val<3>.n2 sar_val<3>.t1 259.736
R1071 sar_val<3>.n2 sar_val<3>.t0 175.083
R1072 sar_val<3>.n3 sar_val<3>.n2 7.36568
R1073 sar_val<3>.n7 sar_val<3>.n5 3.03311
R1074 sar_val<3>.n5 sar_val<3>.n4 2.42212
R1075 sar_val<3>.n9 sar_val<3> 1.41121
R1076 sar_val<3>.n8 sar_val<3>.n7 1.11928
R1077 sar_val<3> sar_val<3>.n9 0.760115
R1078 sar_val<3>.n4 sar_val<3> 0.692392
R1079 sar_val<3>.n5 sar_val<3>.n3 0.519419
R1080 sar_val<3>.n9 sar_val<3>.n8 0.0643193
R1081 sar_val<3>.n7 sar_val<3>.n6 0.0278438
R1082 sar_val<3>.n8 sar_val<3>.n0 0.0141422
R1083 sar_val<3>.n7 sar_val<3>.n1 0.00635938
R1084 sw<3>.t1 sw<3> 459.913
R1085 sw<3>.n4 sw<3>.t1 137.642
R1086 sw<3>.n3 sw<3>.t0 123.654
R1087 sw<3> sw<3>.n3 78.8791
R1088 sw<3>.n5 sw<3>.n1 9.31851
R1089 sw<3>.n6 sw<3>.n5 9.3005
R1090 sw<3> sw<3>.n2 7.16781
R1091 sw<3>.n4 sw<3> 6.30577
R1092 sw<3>.n3 sw<3> 5.16973
R1093 sw<3>.n6 sw<3>.n0 4.5337
R1094 sw<3>.n8 sw<3>.n7 4.5005
R1095 sw<3>.n7 sw<3>.n2 2.55168
R1096 sw<3>.n5 sw<3>.n2 2.13835
R1097 sw<3>.n1 sw<3>.n0 1.12656
R1098 sw<3>.n5 sw<3>.n4 0.0710634
R1099 sw<3>.n8 sw<3>.n0 0.0509808
R1100 sw<3> sw<3>.n8 0.0125192
R1101 sw<3>.n7 sw<3>.n6 0.0102656
R1102 sw<3>.n7 sw<3>.n1 0.00683949
R1103 sar_val<6>.n2 sar_val<6>.t0 260.322
R1104 sar_val<6>.n2 sar_val<6>.t1 175.169
R1105 sar_val<6>.n3 sar_val<6>.n2 8.30219
R1106 sar_val<6>.n7 sar_val<6>.n5 4.5005
R1107 sar_val<6>.n5 sar_val<6>.n4 2.42212
R1108 sar_val<6>.n9 sar_val<6> 1.3755
R1109 sar_val<6>.n8 sar_val<6>.n7 1.11928
R1110 sar_val<6> sar_val<6>.n9 0.740885
R1111 sar_val<6>.n4 sar_val<6> 0.692392
R1112 sar_val<6>.n5 sar_val<6>.n3 0.519419
R1113 sar_val<6>.n9 sar_val<6>.n8 0.0643193
R1114 sar_val<6>.n7 sar_val<6>.n6 0.0278438
R1115 sar_val<6>.n8 sar_val<6>.n0 0.0141422
R1116 sar_val<6>.n7 sar_val<6>.n1 0.00635938
R1117 sar_val<4>.n2 sar_val<4>.t0 259.736
R1118 sar_val<4>.n2 sar_val<4>.t1 175.083
R1119 sar_val<4>.n3 sar_val<4>.n2 7.36568
R1120 sar_val<4>.n7 sar_val<4>.n5 3.03311
R1121 sar_val<4>.n5 sar_val<4>.n4 2.42212
R1122 sar_val<4>.n9 sar_val<4> 1.41121
R1123 sar_val<4>.n8 sar_val<4>.n7 1.11928
R1124 sar_val<4> sar_val<4>.n9 0.760115
R1125 sar_val<4>.n4 sar_val<4> 0.692392
R1126 sar_val<4>.n5 sar_val<4>.n3 0.519419
R1127 sar_val<4>.n9 sar_val<4>.n8 0.0643193
R1128 sar_val<4>.n7 sar_val<4>.n6 0.0278438
R1129 sar_val<4>.n8 sar_val<4>.n0 0.0141422
R1130 sar_val<4>.n7 sar_val<4>.n1 0.00635938
R1131 sw<4>.n5 sw<4>.n3 197.595
R1132 sw<4> sw<4>.n4 165.219
R1133 sw<4>.n2 sw<4>.n0 138.054
R1134 sw<4>.n2 sw<4>.n1 107.874
R1135 sw<4>.n3 sw<4>.t4 26.5955
R1136 sw<4>.n3 sw<4>.t6 26.5955
R1137 sw<4>.n4 sw<4>.t5 26.5955
R1138 sw<4>.n4 sw<4>.t7 26.5955
R1139 sw<4>.n0 sw<4>.t0 24.9236
R1140 sw<4>.n0 sw<4>.t2 24.9236
R1141 sw<4>.n1 sw<4>.t1 24.9236
R1142 sw<4>.n1 sw<4>.t3 24.9236
R1143 sw<4> sw<4>.n6 7.1971
R1144 sw<4> sw<4>.n5 6.59444
R1145 sw<4>.n6 sw<4> 6.20656
R1146 sw<4> sw<4>.n2 2.97424
R1147 sw<4>.n6 sw<4> 2.58636
R1148 sw<4>.n5 sw<4> 2.19848
R1149 sar_val<5>.n2 sar_val<5>.t0 259.736
R1150 sar_val<5>.n2 sar_val<5>.t1 175.083
R1151 sar_val<5>.n3 sar_val<5>.n2 7.36568
R1152 sar_val<5>.n7 sar_val<5>.n5 3.03311
R1153 sar_val<5>.n5 sar_val<5>.n4 2.42212
R1154 sar_val<5>.n9 sar_val<5> 1.38889
R1155 sar_val<5>.n8 sar_val<5>.n7 1.11928
R1156 sar_val<5> sar_val<5>.n9 0.748096
R1157 sar_val<5>.n4 sar_val<5> 0.692392
R1158 sar_val<5>.n5 sar_val<5>.n3 0.519419
R1159 sar_val<5>.n9 sar_val<5>.n8 0.0643193
R1160 sar_val<5>.n7 sar_val<5>.n6 0.0278438
R1161 sar_val<5>.n8 sar_val<5>.n0 0.0141422
R1162 sar_val<5>.n7 sar_val<5>.n1 0.00635938
C0 sw<4> a_795_n2019# 3.79e-20
C1 sw<4> a_n101_n1993# 0.00188f
C2 x12.X sw<2> 2.56e-20
C3 sar_val<4> sar_val<5> 0.0642f
C4 a_n113_n2633# a_n101_n1993# 0.00305f
C5 sw<4> x11.A 1.58e-19
C6 sar_val<6> x4.X 0.00234f
C7 a_n85_n1195# sar_val<4> 0.00156f
C8 sw<4> x4.X 0.0139f
C9 a_1543_n2633# sw<2> 7.94e-21
C10 VDD sw<3> 0.389f
C11 sw<5> x3.X 0.0295f
C12 x3.X sw<2> 1.49e-20
C13 x9.X sw<2> 8.94e-22
C14 a_765_n2468# sar_val<5> 0.00206f
C15 VDD sar_val<3> 0.0917f
C16 VDD a_163_n2633# 0.201f
C17 a_1317_n2468# a_1543_n2633# 0.0873f
C18 a_n85_n1195# a_765_n2468# 5.84e-19
C19 sw<5> a_255_n2019# 0.0109f
C20 a_439_n2633# sw<2> 7.78e-20
C21 x7.X x3.X 1.65e-21
C22 a_1317_n2468# x9.X 0.0025f
C23 a_255_n2019# sw<2> 0.00224f
C24 a_1317_n2468# x3.X 0.00469f
C25 a_991_n2633# sw<2> 1.87e-20
C26 a_255_n2019# x7.X 0.0035f
C27 sw<6> sar_val<4> 2.16e-19
C28 a_1317_n2468# a_991_n2633# 0.0245f
C29 sar_val<5> sw<3> 0.0393f
C30 VDD sar_val<7> 0.138f
C31 VDD a_1347_n2019# 0.412f
C32 x12.X x3.X 0.00124f
C33 x12.X x9.X 7.31e-21
C34 a_n85_n1195# sw<3> 0.032f
C35 sw<5> a_795_n2019# 0.222f
C36 sw<5> a_n101_n1993# 1.35e-19
C37 x12.X a_439_n2633# 0.00253f
C38 a_163_n2633# sar_val<5> 0.0326f
C39 a_n101_n1993# sw<2> 0.0149f
C40 a_n85_n1195# sar_val<3> 1.1e-19
C41 a_n85_n1195# a_163_n2633# 7.15e-20
C42 sw<5> x11.A 0.0592f
C43 sw<6> a_765_n2468# 8.54e-21
C44 a_1543_n2633# x3.X 0.00126f
C45 a_1543_n2633# x9.X 0.115f
C46 x11.A sw<2> 3.52e-21
C47 VDD sar_val<6> 0.138f
C48 x7.X a_n101_n1993# 0.107f
C49 sw<5> x4.X 0.0414f
C50 sw<4> VDD 0.462f
C51 x4.X sw<2> 4.07e-20
C52 x3.X x9.X 0.0509f
C53 x11.A x7.X 3.5e-22
C54 a_1317_n2468# x11.A 5.59e-19
C55 sar_val<7> sar_val<5> 2.2e-19
C56 VDD a_n113_n2633# 0.202f
C57 x4.X x7.X 8.93e-21
C58 a_439_n2633# x3.X 1.35e-20
C59 a_n85_n1195# sar_val<7> 8.55e-20
C60 a_n85_n1195# a_1347_n2019# 4.69e-19
C61 a_1317_n2468# x4.X 2.9e-20
C62 a_255_n2019# x3.X 2.69e-19
C63 a_991_n2633# x3.X 0.115f
C64 a_991_n2633# x9.X 2.38e-20
C65 sw<6> sw<3> 0.0492f
C66 a_255_n2019# a_439_n2633# 4.95e-19
C67 sar_val<3> sw<6> 8.15e-20
C68 sar_val<6> sar_val<5> 0.028f
C69 x4.X x12.X 0.186f
C70 x8.X sar_val<7> 0.0023f
C71 a_n85_n1195# sar_val<6> 2.78e-19
C72 sw<4> sar_val<5> 0.00144f
C73 a_n85_n1195# sw<4> 0.0152f
C74 a_795_n2019# x3.X 0.211f
C75 a_n101_n1993# x3.X 2.99e-21
C76 a_795_n2019# x9.X 1.45e-19
C77 x11.A a_1543_n2633# 3.2e-19
C78 a_n85_n1195# a_n113_n2633# 2.13e-19
C79 x4.X a_1543_n2633# 1.86e-20
C80 x11.A x3.X 0.0356f
C81 x11.A x9.X 0.0328f
C82 sar_val<6> x8.X 0.00243f
C83 a_795_n2019# a_255_n2019# 6.6e-19
C84 a_255_n2019# a_n101_n1993# 0.0151f
C85 a_795_n2019# a_991_n2633# 2.72e-19
C86 x4.X x9.X 1.74e-19
C87 x4.X x3.X 0.0501f
C88 x11.A a_255_n2019# 2.45e-20
C89 sw<5> VDD 0.618f
C90 x4.X a_439_n2633# 0.112f
C91 x4.X a_255_n2019# 0.211f
C92 VDD sw<2> 0.376f
C93 x4.X a_991_n2633# 0.00178f
C94 sar_val<6> sw<6> 2.85e-19
C95 VDD x7.X 0.159f
C96 sw<4> sw<6> 0.0317f
C97 a_795_n2019# a_n101_n1993# 6.3e-20
C98 a_1317_n2468# VDD 0.223f
C99 sar_val<4> sw<3> 0.00504f
C100 x11.A a_795_n2019# 0.0107f
C101 x11.A a_n101_n1993# 4.97e-20
C102 sar_val<3> sar_val<4> 0.0647f
C103 a_163_n2633# sar_val<4> 0.205f
C104 a_795_n2019# x4.X 0.0254f
C105 x4.X a_n101_n1993# 1.4e-20
C106 VDD x12.X 0.101f
C107 sar_val<5> sw<2> 3.04e-20
C108 sw<5> a_n85_n1195# 0.0497f
C109 x11.A x4.X 1.31e-19
C110 a_n85_n1195# sw<2> 0.0222f
C111 a_n85_n1195# x7.X 0.0011f
C112 VDD a_1543_n2633# 0.219f
C113 a_1317_n2468# a_n85_n1195# 4.16e-20
C114 VDD x3.X 0.546f
C115 VDD x9.X 0.436f
C116 x8.X sw<2> 7.97e-21
C117 x12.X sar_val<5> 0.00246f
C118 VDD a_439_n2633# 0.2f
C119 VDD a_255_n2019# 0.437f
C120 a_n85_n1195# x12.X 1.25e-19
C121 sar_val<6> sar_val<4> 1.47e-20
C122 VDD a_991_n2633# 0.222f
C123 a_1317_n2468# x8.X 0.107f
C124 sar_val<3> sw<3> 1.27e-20
C125 a_163_n2633# sw<3> 0.11f
C126 sw<5> sw<6> 0.0587f
C127 sw<4> sar_val<4> 0.0018f
C128 sw<6> sw<2> 0.122f
C129 a_n113_n2633# sar_val<4> 0.0326f
C130 sar_val<3> a_163_n2633# 1.71e-19
C131 a_n85_n1195# a_1543_n2633# 1.92e-20
C132 sar_val<5> x3.X 5.16e-21
C133 sar_val<6> a_765_n2468# 0.00483f
C134 a_n85_n1195# x3.X 0.00507f
C135 VDD a_795_n2019# 0.463f
C136 VDD a_n101_n1993# 0.207f
C137 sar_val<5> a_439_n2633# 0.205f
C138 a_255_n2019# sar_val<5> 0.00467f
C139 a_n85_n1195# a_439_n2633# 5.15e-19
C140 VDD x11.A 0.839f
C141 a_n85_n1195# a_255_n2019# 0.0196f
C142 a_n85_n1195# a_991_n2633# 3.66e-19
C143 VDD x4.X 0.402f
C144 x8.X x9.X 0.00126f
C145 x8.X x3.X 0.186f
C146 sar_val<6> sw<3> 9.58e-21
C147 sw<4> sw<3> 0.365f
C148 x8.X a_991_n2633# 0.00253f
C149 sar_val<6> sar_val<3> 8.41e-21
C150 sar_val<6> a_163_n2633# 1.49e-20
C151 sar_val<7> a_1347_n2019# 0.00496f
C152 a_n113_n2633# sw<3> 3.5e-20
C153 a_n85_n1195# a_795_n2019# 0.0136f
C154 a_n85_n1195# a_n101_n1993# 0.00329f
C155 sw<6> x3.X 0.00185f
C156 sw<4> a_163_n2633# 0.00127f
C157 sar_val<3> a_n113_n2633# 0.205f
C158 sw<6> a_439_n2633# 8.67e-21
C159 a_n113_n2633# a_163_n2633# 5.3e-19
C160 sar_val<4> sw<2> 0.0393f
C161 a_n85_n1195# x11.A 0.652f
C162 x4.X sar_val<5> 0.00504f
C163 sw<6> a_255_n2019# 7.21e-19
C164 sw<6> a_991_n2633# 5.23e-21
C165 a_n85_n1195# x4.X 0.00512f
C166 sar_val<6> sar_val<7> 0.0325f
C167 sw<4> a_1347_n2019# 3.61e-21
C168 x11.A x8.X 1.41e-19
C169 sw<5> a_765_n2468# 2.62e-20
C170 a_765_n2468# sw<2> 2.92e-20
C171 x4.X x8.X 2.54e-20
C172 sw<6> a_795_n2019# 0.00155f
C173 sw<6> a_n101_n1993# 1.06e-19
C174 x11.A sw<6> 0.00792f
C175 sar_val<6> a_n113_n2633# 8.03e-21
C176 sw<5> sw<3> 0.0876f
C177 sw<6> x4.X 3.1e-19
C178 sw<3> sw<2> 0.106f
C179 x12.X a_765_n2468# 0.107f
C180 sar_val<4> x3.X 2.73e-21
C181 x7.X sw<3> 0.00116f
C182 sar_val<3> sw<2> 0.00505f
C183 a_163_n2633# sw<2> 0.111f
C184 sar_val<4> a_439_n2633# 1.5e-19
C185 VDD sar_val<5> 0.0973f
C186 a_n85_n1195# VDD 1.47f
C187 a_765_n2468# x9.X 1.47e-20
C188 a_765_n2468# x3.X 0.00246f
C189 sw<5> a_1347_n2019# 6.21e-19
C190 sar_val<7> sw<2> 3.34e-21
C191 a_765_n2468# a_439_n2633# 0.0245f
C192 a_991_n2633# a_765_n2468# 0.0873f
C193 VDD x8.X 0.114f
C194 a_1317_n2468# sar_val<7> 0.00464f
C195 a_1317_n2468# a_1347_n2019# 0.00179f
C196 sw<5> sar_val<6> 0.00165f
C197 sar_val<6> sw<2> 1.27e-20
C198 x3.X sw<3> 9.76e-21
C199 sw<5> sw<4> 0.00156f
C200 sw<4> sw<2> 0.352f
C201 a_439_n2633# sw<3> 0.111f
C202 VDD sw<6> 1.71f
C203 sar_val<3> x3.X 1.67e-21
C204 a_163_n2633# x3.X 6.99e-21
C205 a_1317_n2468# sar_val<6> 0.00205f
C206 a_255_n2019# sw<3> 0.0227f
C207 a_795_n2019# a_765_n2468# 0.00179f
C208 a_n113_n2633# sw<2> 0.11f
C209 sw<4> x7.X 0.0205f
C210 a_163_n2633# a_439_n2633# 5.3e-19
C211 a_255_n2019# a_163_n2633# 0.00206f
C212 sar_val<7> a_1543_n2633# 0.205f
C213 a_1543_n2633# a_1347_n2019# 2.72e-19
C214 sar_val<6> x12.X 0.00236f
C215 x4.X a_765_n2468# 0.00552f
C216 sar_val<7> x3.X 0.00213f
C217 sar_val<7> x9.X 0.00539f
C218 x3.X a_1347_n2019# 0.0242f
C219 a_1347_n2019# x9.X 0.211f
C220 a_795_n2019# sw<3> 6.25e-19
C221 a_n101_n1993# sw<3> 3.7e-20
C222 a_991_n2633# sar_val<7> 0.00178f
C223 sar_val<6> a_1543_n2633# 8.56e-20
C224 a_n85_n1195# sw<6> 1.71f
C225 x11.A sw<3> 7.33e-21
C226 sar_val<3> a_n101_n1993# 0.001f
C227 x4.X sw<3> 0.12f
C228 sar_val<6> x9.X 9.3e-21
C229 sar_val<6> x3.X 0.0053f
C230 sw<4> x3.X 1.96e-20
C231 sar_val<6> a_439_n2633# 0.00172f
C232 sar_val<6> a_991_n2633# 0.205f
C233 a_n113_n2633# x3.X 4.23e-21
C234 sw<5> sw<2> 1.58e-21
C235 a_795_n2019# a_1347_n2019# 6.05e-19
C236 VDD sar_val<4> 0.0978f
C237 sw<4> a_255_n2019# 0.223f
C238 a_n101_n1993# a_1347_n2019# 7.93e-21
C239 sw<5> x7.X 2.1e-21
C240 x11.A sar_val<7> 0.00181f
C241 x11.A a_1347_n2019# 0.24f
C242 x7.X sw<2> 0.0208f
C243 a_1317_n2468# sw<2> 1.06e-20
C244 x4.X sar_val<7> 7.79e-21
C245 x4.X a_1347_n2019# 5.03e-21
C246 sar_val<6> a_795_n2019# 0.00499f
C247 VDD a_765_n2468# 0.216f
C248 x8.X VSS 0.0754f
C249 x12.X VSS 0.0809f
C250 sw<3> VSS 0.429f
C251 sw<2> VSS 0.583f
C252 a_1543_n2633# VSS 0.258f
C253 sar_val<7> VSS 0.436f
C254 a_1317_n2468# VSS 0.435f
C255 a_991_n2633# VSS 0.237f
C256 sar_val<6> VSS 0.405f
C257 a_765_n2468# VSS 0.437f
C258 a_439_n2633# VSS 0.245f
C259 sar_val<5> VSS 0.342f
C260 a_163_n2633# VSS 0.238f
C261 sar_val<4> VSS 0.33f
C262 a_n113_n2633# VSS 0.301f
C263 sar_val<3> VSS 0.404f
C264 sw<5> VSS 0.553f
C265 sw<4> VSS 0.543f
C266 x7.X VSS 0.119f
C267 x9.X VSS 0.479f
C268 a_1347_n2019# VSS 0.571f
C269 x3.X VSS 0.257f
C270 a_795_n2019# VSS 0.544f
C271 x4.X VSS 0.324f
C272 a_255_n2019# VSS 0.574f
C273 a_n101_n1993# VSS 0.518f
C274 sw<6> VSS 1.47f
C275 x11.A VSS 1.24f
C276 a_n85_n1195# VSS 2.15f
C277 VDD VSS 10.2f
.ends

