magic
tech sky130A
timestamp 1699450567
<< end >>
