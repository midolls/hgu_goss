* NGSPICE file created from hgu_cdac_cap_2.ext - technology: sky130A


* Top level circuit hgu_cdac_cap_2

C0 hgu_cdac_unit_1.C0 hgu_cdac_unit_1.C1 4.31f
C1 hgu_cdac_unit_0.C1 hgu_cdac_unit_1.C1 4.47f
C2 hgu_cdac_unit_1.C1 VSUBS 1.26f $ **FLOATING
C3 hgu_cdac_unit_0.C1 VSUBS 1.24f $ **FLOATING
.end

