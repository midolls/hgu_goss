magic
tech sky130A
magscale 1 2
timestamp 1697026607
<< checkpaint >>
rect 866 -1074 3808 2480
<< error_p >>
rect 4962 7292 4997 7301
rect 4926 7267 4997 7292
rect 4323 7251 4358 7256
rect 4287 7222 4358 7251
rect 4287 6783 4357 7222
rect 4287 6747 4340 6783
rect 4926 6730 4996 7267
rect 5658 7056 5692 7110
rect 6080 7092 6115 7097
rect 6044 7063 6115 7092
rect 4926 6694 4979 6730
rect 5677 6677 5692 7056
rect 5711 7022 5746 7056
rect 5711 6677 5745 7022
rect 5857 6954 5915 6960
rect 5857 6920 5869 6954
rect 5857 6914 5915 6920
rect 5857 6760 5915 6766
rect 5857 6726 5869 6760
rect 5857 6720 5915 6726
rect 5711 6643 5726 6677
rect 6044 6624 6114 7063
rect 6226 6995 6284 7001
rect 6226 6961 6238 6995
rect 6396 6986 6430 7001
rect 6818 6986 6853 6991
rect 6226 6955 6284 6961
rect 6396 6950 6466 6986
rect 6782 6957 6853 6986
rect 7133 6964 7168 6982
rect 7556 6964 7590 6982
rect 7133 6957 7204 6964
rect 6413 6916 6484 6950
rect 6226 6707 6284 6713
rect 6226 6673 6238 6707
rect 6226 6667 6284 6673
rect 6044 6588 6097 6624
rect 6413 6571 6483 6916
rect 6595 6848 6653 6854
rect 6595 6814 6607 6848
rect 6595 6808 6653 6814
rect 6595 6654 6653 6660
rect 6595 6620 6607 6654
rect 6595 6614 6653 6620
rect 6413 6535 6466 6571
rect 6782 6518 6852 6957
rect 7134 6928 7204 6957
rect 6964 6889 7022 6895
rect 7151 6894 7222 6928
rect 6964 6855 6976 6889
rect 6964 6849 7022 6855
rect 6964 6601 7022 6607
rect 6964 6567 6976 6601
rect 6964 6561 7022 6567
rect 6782 6482 6835 6518
rect 7151 6465 7221 6894
rect 7333 6826 7391 6832
rect 7333 6792 7345 6826
rect 7333 6786 7391 6792
rect 7333 6548 7391 6554
rect 7333 6514 7345 6548
rect 7333 6508 7391 6514
rect 7151 6429 7204 6465
rect 7520 6412 7590 6964
rect 7702 6943 7760 6949
rect 7702 6909 7714 6943
rect 7702 6903 7760 6909
rect 7702 6495 7760 6501
rect 7702 6461 7714 6495
rect 7702 6455 7760 6461
rect 7520 6376 7573 6412
<< error_s >>
rect 2544 2901 2585 2933
rect 640 1422 682 1478
rect 676 1339 684 1391
rect 827 1340 885 1346
rect 196 1305 226 1315
rect 190 1289 226 1305
rect 190 1285 224 1289
rect 190 1271 226 1285
rect 234 1271 264 1289
rect 274 1271 304 1305
rect 642 1271 666 1305
rect 156 1243 186 1271
rect 196 1237 226 1247
rect 158 1209 188 1219
rect 152 1184 188 1209
rect 190 1203 226 1237
rect 234 1243 270 1271
rect 510 1257 540 1267
rect 234 1209 264 1243
rect 504 1241 540 1257
rect 504 1237 538 1241
rect 196 1184 226 1193
rect 234 1184 266 1209
rect 274 1203 304 1237
rect 152 1175 266 1184
rect 118 1147 275 1175
rect 318 1147 324 1237
rect 504 1223 540 1237
rect 548 1223 578 1241
rect 588 1223 618 1257
rect 676 1237 700 1339
rect 827 1306 839 1340
rect 827 1300 885 1306
rect 352 1175 358 1209
rect 470 1195 500 1223
rect 510 1189 540 1199
rect 472 1161 502 1171
rect 147 1137 275 1147
rect 152 1133 275 1137
rect 466 1136 502 1161
rect 504 1155 540 1189
rect 548 1195 584 1223
rect 548 1161 578 1195
rect 510 1136 540 1145
rect 548 1136 580 1161
rect 588 1155 618 1189
rect 676 1137 684 1237
rect 1570 1232 1628 1238
rect 1570 1198 1582 1232
rect 1570 1192 1628 1198
rect 152 1107 384 1133
rect 466 1127 580 1136
rect 144 1091 182 1103
rect 188 1091 384 1107
rect 432 1099 589 1127
rect 106 1088 121 1090
rect 144 1088 384 1091
rect 461 1089 589 1099
rect 72 993 73 1079
rect 106 1071 384 1088
rect 466 1071 592 1089
rect 676 1071 710 1089
rect 106 1049 710 1071
rect 104 1045 710 1049
rect 106 995 107 1045
rect 109 1041 710 1045
rect 114 1011 710 1041
rect 123 1003 710 1011
rect 140 995 710 1003
rect 68 992 73 993
rect 118 992 710 995
rect 68 945 710 992
rect 1002 1005 1036 1023
rect 1424 1005 1458 1023
rect 1002 969 1072 1005
rect 68 851 73 945
rect 102 911 107 945
rect 113 909 710 945
rect 113 899 331 909
rect 382 899 390 905
rect 80 839 331 899
rect 377 840 390 899
rect 416 897 424 909
rect 448 903 540 909
rect 448 897 510 903
rect 407 888 510 897
rect 407 865 534 888
rect 407 863 504 865
rect 407 861 502 863
rect 548 861 578 909
rect 588 903 618 909
rect 623 903 710 909
rect 623 891 630 903
rect 401 857 479 861
rect 401 852 491 857
rect 497 852 502 861
rect 401 847 502 852
rect 510 849 540 859
rect 589 857 600 891
rect 623 887 634 891
rect 640 887 710 903
rect 401 846 454 847
rect 80 817 320 839
rect 68 813 320 817
rect 68 809 86 813
rect 102 809 120 813
rect 106 783 113 809
rect 166 801 240 813
rect 248 809 255 813
rect 297 809 320 813
rect 405 829 454 846
rect 405 813 445 829
rect 457 813 502 847
rect 405 812 502 813
rect 188 783 240 801
rect 411 807 502 812
rect 509 813 543 849
rect 549 823 581 857
rect 106 775 158 783
rect 68 763 86 775
rect 102 743 158 775
rect 167 763 240 783
rect 167 747 248 763
rect 167 743 240 747
rect 102 729 167 743
rect 68 713 79 729
rect 102 713 113 729
rect 143 714 259 729
rect 148 713 259 714
rect 297 603 303 783
rect 411 779 497 807
rect 411 761 445 779
rect 411 745 453 761
rect 472 756 497 779
rect 457 745 497 756
rect 411 727 497 745
rect 411 711 462 727
rect 263 535 276 569
rect 297 501 310 603
rect 318 597 331 699
rect 411 673 445 711
rect 472 695 497 727
rect 509 779 546 813
rect 550 807 580 823
rect 589 795 600 823
rect 623 791 710 887
rect 509 761 543 779
rect 623 761 634 791
rect 509 745 545 761
rect 509 711 546 745
rect 497 669 502 695
rect 509 673 543 711
rect 352 631 365 665
rect 381 657 415 665
rect 473 657 507 665
rect 381 635 544 657
rect 565 635 581 665
rect 410 631 544 635
rect 444 597 510 623
rect 460 593 494 597
rect 640 487 710 791
rect 1019 935 1090 969
rect 827 570 885 576
rect 827 536 839 570
rect 827 530 885 536
rect 640 451 693 487
rect 1019 434 1089 935
rect 1201 867 1259 873
rect 1201 833 1213 867
rect 1201 827 1259 833
rect 1201 517 1259 523
rect 1201 483 1213 517
rect 1201 477 1259 483
rect 1019 398 1072 434
rect 1388 381 1458 1005
rect 1740 859 1774 877
rect 1740 823 1810 859
rect 1757 789 1828 823
rect 1570 464 1628 470
rect 1570 430 1582 464
rect 1570 424 1628 430
rect 1388 345 1441 381
rect 1757 328 1827 789
rect 1939 721 1997 727
rect 1939 687 1951 721
rect 1939 681 1997 687
rect 1939 411 1997 417
rect 1939 377 1951 411
rect 1939 371 1997 377
rect 1757 292 1810 328
use hgu_clk_div  x1
timestamp 1697026605
transform 1 0 152 0 1 2088
box -152 -1488 3058 1192
use hgu_delay  x2
timestamp 1697026606
transform 1 0 3263 0 1 6200
box -53 -5600 4679 1137
use sky130_fd_sc_hd__nand2_1  x3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 0 0 1 552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x7 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 7942 0 1 600
box -38 -48 314 592
use sky130_fd_pr__nfet_01v8_723X3M  XM1
timestamp 0
transform 1 0 477 0 1 761
box -216 -310 216 310
use sky130_fd_pr__pfet_01v8_BMSA97  XM2
timestamp 0
transform 1 0 856 0 1 938
box -216 -540 216 540
use sky130_fd_pr__nfet_01v8_8X7SK7  XM3
timestamp 0
transform 1 0 1230 0 1 675
box -211 -330 211 330
use sky130_fd_pr__pfet_01v8_U4MAJH  XM4
timestamp 0
transform 1 0 1599 0 1 831
box -211 -539 211 539
use sky130_fd_pr__nfet_01v8_648S5X  XM5
timestamp 0
transform 1 0 1968 0 1 549
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_MYDY2X  XM6
timestamp 0
transform 1 0 2337 0 1 703
box -211 -517 211 517
<< end >>
