magic
tech sky130A
magscale 1 2
timestamp 1698501754
<< ndiff >>
rect 791 827 825 843
rect 791 757 825 771
<< ndiffc >>
rect 94 771 128 827
rect 791 771 825 827
<< poly >>
rect 135 888 179 903
rect 135 858 780 888
<< locali >>
rect 94 827 128 843
rect 94 693 128 771
rect 791 827 825 905
rect 791 755 825 771
use sky130_fd_pr__nfet_01v8_56T3VD  XM1
timestamp 1698498532
transform -1 0 693 0 1 800
box -73 -69 73 69
use sky130_fd_pr__nfet_01v8_56T3VD  XM2
timestamp 1698498532
transform -1 0 621 0 1 800
box -73 -69 73 69
use sky130_fd_pr__nfet_01v8_56T3VD  XM3
timestamp 1698498532
transform -1 0 549 0 1 800
box -73 -69 73 69
use sky130_fd_pr__nfet_01v8_56T3VD  XM4
timestamp 1698498532
transform -1 0 477 0 1 800
box -73 -69 73 69
use sky130_fd_pr__nfet_01v8_56T3VD  XM5
timestamp 1698498532
transform -1 0 405 0 1 800
box -73 -69 73 69
use sky130_fd_pr__nfet_01v8_56T3VD  XM6
timestamp 1698498532
transform -1 0 765 0 1 800
box -73 -69 73 69
use sky130_fd_pr__nfet_01v8_L7T3GD  XM7
timestamp 1698498532
transform -1 0 302 0 1 799
box -73 -68 73 68
use sky130_fd_pr__nfet_01v8_L7T3GD  XM8
timestamp 1698498532
transform -1 0 230 0 1 799
box -73 -68 73 68
use sky130_fd_pr__nfet_01v8_L7T3GD  XM9
timestamp 1698498532
transform -1 0 158 0 1 799
box -73 -68 73 68
<< end >>
