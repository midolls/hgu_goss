magic
tech sky130A
magscale 1 2
timestamp 1699322317
<< checkpaint >>
rect -1313 2258 1629 2311
rect -1313 2205 1998 2258
rect -1313 2152 2367 2205
rect -1313 2099 2736 2152
rect -1313 2046 3105 2099
rect -1313 1993 3474 2046
rect -1313 1940 3843 1993
rect -1313 1887 4212 1940
rect -1313 1834 4581 1887
rect -1313 1781 4950 1834
rect -1313 1728 5319 1781
rect -1313 1675 5688 1728
rect -1313 1622 6057 1675
rect -1313 1569 6426 1622
rect -1313 1516 6795 1569
rect -1313 -713 7164 1516
rect -944 -766 7164 -713
rect -575 -819 7164 -766
rect -206 -872 7164 -819
rect 163 -925 7164 -872
rect 532 -978 7164 -925
rect 901 -1031 7164 -978
rect 1270 -1084 7164 -1031
rect 1639 -1137 7164 -1084
rect 2008 -1190 7164 -1137
rect 2377 -1243 7164 -1190
rect 2746 -1296 7164 -1243
rect 3115 -1349 7164 -1296
rect 3484 -1402 7164 -1349
rect 3853 -1455 7164 -1402
rect 4222 -1508 7164 -1455
<< error_s >>
rect 298 981 333 1015
rect 299 962 333 981
rect 129 913 187 919
rect 129 879 141 913
rect 318 879 333 962
rect 129 873 187 879
rect 215 769 219 840
rect 223 769 225 841
rect 215 719 233 769
rect 251 729 253 841
rect 265 753 291 845
rect 93 703 169 719
rect 173 703 233 719
rect 110 691 213 703
rect 103 685 213 691
rect 103 671 143 685
rect 85 619 143 671
rect 173 671 191 685
rect 265 671 291 707
rect 299 671 333 879
rect 173 619 215 671
rect 245 619 333 671
rect 265 617 291 619
rect 299 617 333 619
rect 31 583 333 617
rect 352 928 387 962
rect 667 928 702 962
rect 352 583 386 928
rect 668 909 702 928
rect 498 860 556 866
rect 498 826 510 860
rect 498 820 556 826
rect 498 666 556 672
rect 498 632 510 666
rect 498 626 556 632
rect 97 565 131 569
rect 257 565 291 569
rect 85 558 143 565
rect 173 558 215 565
rect 245 558 303 565
rect 97 549 131 558
rect 257 549 291 558
rect 352 549 367 583
rect 352 530 357 549
rect 687 530 702 909
rect 721 875 756 909
rect 1036 875 1071 909
rect 721 530 755 875
rect 1037 856 1071 875
rect 867 807 925 813
rect 867 773 879 807
rect 867 767 925 773
rect 867 613 925 619
rect 867 579 879 613
rect 867 573 925 579
rect 721 496 736 530
rect 1056 477 1071 856
rect 1090 822 1125 856
rect 1405 822 1440 856
rect 1090 477 1124 822
rect 1406 803 1440 822
rect 1236 754 1294 760
rect 1236 720 1248 754
rect 1236 714 1294 720
rect 1236 560 1294 566
rect 1236 526 1248 560
rect 1236 520 1294 526
rect 1090 443 1105 477
rect 1425 424 1440 803
rect 1459 769 1494 803
rect 1774 769 1809 803
rect 1459 424 1493 769
rect 1775 750 1809 769
rect 1605 701 1663 707
rect 1605 667 1617 701
rect 1605 661 1663 667
rect 1605 507 1663 513
rect 1605 473 1617 507
rect 1605 467 1663 473
rect 1459 390 1474 424
rect 1794 371 1809 750
rect 1828 716 1863 750
rect 2143 716 2178 750
rect 1828 371 1862 716
rect 2144 697 2178 716
rect 1974 648 2032 654
rect 1974 614 1986 648
rect 1974 608 2032 614
rect 1974 454 2032 460
rect 1974 420 1986 454
rect 1974 414 2032 420
rect 1828 337 1843 371
rect 2163 318 2178 697
rect 2197 663 2232 697
rect 2512 663 2547 697
rect 2197 318 2231 663
rect 2513 644 2547 663
rect 2343 595 2401 601
rect 2343 561 2355 595
rect 2343 555 2401 561
rect 2343 401 2401 407
rect 2343 367 2355 401
rect 2343 361 2401 367
rect 2197 284 2212 318
rect 2532 265 2547 644
rect 2566 610 2601 644
rect 2881 610 2916 644
rect 2566 265 2600 610
rect 2882 591 2916 610
rect 2712 542 2770 548
rect 2712 508 2724 542
rect 2712 502 2770 508
rect 2712 348 2770 354
rect 2712 314 2724 348
rect 2712 308 2770 314
rect 2566 231 2581 265
rect 91 205 137 228
rect 2901 212 2916 591
rect 2935 557 2970 591
rect 3250 557 3285 591
rect 2935 212 2969 557
rect 3251 538 3285 557
rect 3081 489 3139 495
rect 3081 455 3093 489
rect 3081 449 3139 455
rect 3081 295 3139 301
rect 3081 261 3093 295
rect 3081 255 3139 261
rect 63 177 165 200
rect 2935 178 2950 212
rect 3270 159 3285 538
rect 3304 504 3339 538
rect 3619 504 3654 538
rect 3304 159 3338 504
rect 3620 485 3654 504
rect 3450 436 3508 442
rect 3450 402 3462 436
rect 3450 396 3508 402
rect 3450 242 3508 248
rect 3450 208 3462 242
rect 3450 202 3508 208
rect 3304 125 3319 159
rect 3639 106 3654 485
rect 3673 451 3708 485
rect 3988 451 4023 485
rect 3673 106 3707 451
rect 3989 432 4023 451
rect 3819 383 3877 389
rect 3819 349 3831 383
rect 3819 343 3877 349
rect 3819 189 3877 195
rect 3819 155 3831 189
rect 3819 149 3877 155
rect 3673 72 3688 106
rect 4008 53 4023 432
rect 4042 398 4077 432
rect 4357 398 4392 432
rect 4042 53 4076 398
rect 4358 379 4392 398
rect 4188 330 4246 336
rect 4188 296 4200 330
rect 4188 290 4246 296
rect 4188 136 4246 142
rect 4188 102 4200 136
rect 4188 96 4246 102
rect 4042 19 4057 53
rect 4377 0 4392 379
rect 4411 345 4446 379
rect 4726 345 4761 379
rect 4411 0 4445 345
rect 4727 326 4761 345
rect 4557 277 4615 283
rect 4557 243 4569 277
rect 4557 237 4615 243
rect 4557 83 4615 89
rect 4557 49 4569 83
rect 4557 43 4615 49
rect 4411 -34 4426 0
rect 4746 -53 4761 326
rect 4780 292 4815 326
rect 5095 292 5130 326
rect 4780 -53 4814 292
rect 5096 273 5130 292
rect 4926 224 4984 230
rect 4926 190 4938 224
rect 4926 184 4984 190
rect 4926 30 4984 36
rect 4926 -4 4938 30
rect 4926 -10 4984 -4
rect 4780 -87 4795 -53
rect 5115 -106 5130 273
rect 5149 239 5184 273
rect 5149 -106 5183 239
rect 5295 171 5353 177
rect 5295 137 5307 171
rect 5295 131 5353 137
rect 5295 -23 5353 -17
rect 5295 -57 5307 -23
rect 5295 -63 5353 -57
rect 5149 -140 5164 -106
<< nmos >>
rect 143 757 173 841
rect 215 757 245 841
rect 143 619 173 703
rect 215 619 245 703
rect 143 481 173 565
rect 215 481 245 565
rect 143 343 173 427
rect 215 343 245 427
rect 143 205 173 289
rect 215 205 245 289
rect 143 67 173 151
rect 215 67 245 151
rect 143 -71 173 13
rect 215 -71 245 13
rect 143 -209 173 -125
rect 215 -209 245 -125
<< ndiff >>
rect 85 829 143 841
rect 85 769 97 829
rect 131 769 143 829
rect 85 757 143 769
rect 173 757 215 841
rect 245 829 303 841
rect 245 769 257 829
rect 291 769 303 829
rect 245 757 303 769
rect 85 691 143 703
rect 85 631 97 691
rect 131 631 143 691
rect 85 619 143 631
rect 173 619 215 703
rect 245 691 303 703
rect 245 631 257 691
rect 291 631 303 691
rect 245 619 303 631
rect 85 553 143 565
rect 85 493 97 553
rect 131 493 143 553
rect 85 481 143 493
rect 173 481 215 565
rect 245 553 303 565
rect 245 493 257 553
rect 291 493 303 553
rect 245 481 303 493
rect 85 415 143 427
rect 85 355 97 415
rect 131 355 143 415
rect 85 343 143 355
rect 173 343 215 427
rect 245 415 303 427
rect 245 355 257 415
rect 291 355 303 415
rect 245 343 303 355
rect 85 277 143 289
rect 85 217 97 277
rect 131 217 143 277
rect 85 205 143 217
rect 173 205 215 289
rect 245 277 303 289
rect 245 217 257 277
rect 291 217 303 277
rect 245 205 303 217
rect 85 139 143 151
rect 85 79 97 139
rect 131 79 143 139
rect 85 67 143 79
rect 173 67 215 151
rect 245 139 303 151
rect 245 79 257 139
rect 291 79 303 139
rect 245 67 303 79
rect 85 1 143 13
rect 85 -59 97 1
rect 131 -59 143 1
rect 85 -71 143 -59
rect 173 -71 215 13
rect 245 1 303 13
rect 245 -59 257 1
rect 291 -59 303 1
rect 245 -71 303 -59
rect 85 -137 143 -125
rect 85 -197 97 -137
rect 131 -197 143 -137
rect 85 -209 143 -197
rect 173 -209 215 -125
rect 245 -137 303 -125
rect 245 -197 257 -137
rect 291 -197 303 -137
rect 245 -209 303 -197
<< ndiffc >>
rect 97 769 131 829
rect 257 769 291 829
rect 97 631 131 691
rect 257 631 291 691
rect 97 493 131 553
rect 257 493 291 553
rect 97 355 131 415
rect 257 355 291 415
rect 97 217 131 277
rect 257 217 291 277
rect 97 79 131 139
rect 257 79 291 139
rect 97 -59 131 1
rect 257 -59 291 1
rect 97 -197 131 -137
rect 257 -197 291 -137
<< psubdiff >>
rect -90 -13 14 22
rect -90 -47 -51 -13
rect -17 -47 14 -13
rect -90 -76 14 -47
<< psubdiffcont >>
rect -51 -47 -17 -13
<< poly >>
rect 143 856 245 886
rect 143 841 173 856
rect 215 841 245 856
rect 143 703 173 757
rect 215 703 245 757
rect 143 565 173 619
rect 215 565 245 619
rect 143 427 173 481
rect 215 427 245 481
rect 143 289 173 343
rect 215 289 245 343
rect 143 151 173 205
rect 215 151 245 205
rect 143 13 173 67
rect 215 13 245 67
rect 143 -125 173 -71
rect 215 -125 245 -71
rect 143 -235 173 -209
rect 215 -235 245 -209
<< locali >>
rect 97 829 131 845
rect 97 753 131 769
rect 257 829 291 845
rect 257 753 291 769
rect 97 691 131 707
rect 97 615 131 631
rect 257 691 291 707
rect 257 615 291 631
rect 97 553 131 569
rect 97 477 131 493
rect 257 553 291 569
rect 257 477 291 493
rect 97 415 131 431
rect 97 339 131 355
rect 257 415 291 431
rect 257 339 291 355
rect 97 277 131 293
rect 97 201 131 217
rect 257 277 291 293
rect 257 201 291 217
rect 97 139 131 155
rect 97 63 131 79
rect 257 139 291 155
rect 257 63 291 79
rect -90 -13 15 22
rect -90 -47 -51 -13
rect -17 -47 15 -13
rect -90 -76 15 -47
rect 97 1 131 17
rect 97 -75 131 -59
rect 257 1 291 17
rect 257 -75 291 -59
rect -76 -131 1 -76
rect 97 -131 131 -121
rect -76 -137 131 -131
rect -76 -197 97 -137
rect -76 -200 131 -197
rect 97 -213 131 -200
rect 257 -137 291 -121
rect 257 -213 291 -197
<< viali >>
rect 97 769 131 829
rect 257 769 291 829
rect 97 631 131 691
rect 257 631 291 691
rect 97 493 131 553
rect 257 493 291 553
rect 97 355 131 415
rect 257 355 291 415
rect 97 217 131 277
rect 257 217 291 277
rect 97 79 131 139
rect 257 79 291 139
rect 97 -59 131 1
rect 257 -59 291 1
rect 97 -197 131 -137
rect 257 -197 291 -137
<< metal1 >>
rect 91 829 137 841
rect 91 769 97 829
rect 131 769 137 829
rect 91 757 137 769
rect 251 829 297 841
rect 251 769 257 829
rect 291 769 297 829
rect 91 691 137 703
rect 91 631 97 691
rect 131 631 137 691
rect 91 553 137 631
rect 251 691 297 769
rect 251 631 257 691
rect 291 631 297 691
rect 251 619 297 631
rect 91 493 97 553
rect 131 493 137 553
rect 91 481 137 493
rect 251 553 297 565
rect 251 493 257 553
rect 291 493 297 553
rect 91 415 137 427
rect 91 355 97 415
rect 131 355 137 415
rect 91 277 137 355
rect 251 415 297 493
rect 251 355 257 415
rect 291 355 297 415
rect 251 343 297 355
rect 91 217 97 277
rect 131 217 137 277
rect 91 205 137 217
rect 251 277 297 289
rect 251 217 257 277
rect 291 217 297 277
rect 0 139 200 200
rect 0 79 97 139
rect 131 79 200 139
rect 0 1 200 79
rect 251 139 297 217
rect 251 79 257 139
rect 291 79 297 139
rect 251 67 297 79
rect 0 0 97 1
rect 91 -59 97 0
rect 131 0 200 1
rect 251 1 297 13
rect 131 -59 137 0
rect 91 -71 137 -59
rect 251 -59 257 1
rect 291 -59 297 1
rect 91 -137 137 -125
rect 91 -197 97 -137
rect 131 -197 137 -137
rect 91 -200 137 -197
rect 251 -137 297 -59
rect 251 -197 257 -137
rect 291 -197 297 -137
rect 0 -400 200 -200
rect 251 -209 297 -197
rect 0 -800 200 -600
use sky130_fd_pr__nfet_01v8_L7T3GD  XM1
timestamp 1698825334
transform 1 0 158 0 1 799
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_L7T3GD  XM2
timestamp 1698825334
transform 1 0 527 0 1 746
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_L7T3GD  XM3
timestamp 1698825334
transform 1 0 896 0 1 693
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_L7T3GD  XM4
timestamp 1698825334
transform 1 0 1265 0 1 640
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_L7T3GD  XM5
timestamp 1698825334
transform 1 0 1634 0 1 587
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_L7T3GD  XM6
timestamp 1698825334
transform 1 0 2003 0 1 534
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_L7T3GD  XM7
timestamp 1698825334
transform 1 0 2372 0 1 481
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_L7T3GD  XM8
timestamp 1698825334
transform 1 0 2741 0 1 428
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_L7T3GD  XM9
timestamp 1698825334
transform 1 0 3110 0 1 375
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_L7T3GD  XM10
timestamp 1698825334
transform 1 0 3479 0 1 322
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_L7T3GD  XM11
timestamp 1698825334
transform 1 0 3848 0 1 269
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_L7T3GD  XM12
timestamp 1698825334
transform 1 0 4217 0 1 216
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_L7T3GD  XM13
timestamp 1698825334
transform 1 0 4586 0 1 163
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_L7T3GD  XM14
timestamp 1698825334
transform 1 0 4955 0 1 110
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_L7T3GD  XM15
timestamp 1698825334
transform 1 0 5324 0 1 57
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_L7T3GD  XM16
timestamp 1698825334
transform 1 0 5693 0 1 4
box -211 -252 211 252
<< labels >>
flabel poly 143 856 245 886 0 FreeSans 320 0 0 0 input_stack
port 0 nsew
flabel metal1 97 -197 131 -137 0 FreeSans 320 0 0 0 vss
port 3 nsew
flabel metal1 91 829 137 841 0 FreeSans 320 0 0 0 output_stack
port 5 nsew
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 input_stack
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 output_stack
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 VSS
port 2 nsew
<< end >>
