* NGSPICE file created from hgu_sarlogic_sw_ctrl_flat.ext - technology: sky130A

.subckt hgu_sarlogic_sw_ctrl_flat VSS_SW[1] VSS_SW[2] VSS_SW[3] VSS_SW[4] VSS_SW[5]
+ VSS_SW[6] VSS_SW[7] VDD_SW[2] VDD_SW[3] VDD_SW[4] VDD_SW[5] VDD_SW[6] VDD_SW[7]
+ D[2] D[3] D[4] D[5] D[6] D[7] check[0] check[1] check[2] check[3] check[4] check[5]
+ check[6] VDD_SW_b[1] VDD_SW_b[2] VDD_SW_b[3] VDD_SW_b[4] VDD_SW_b[5] VDD_SW_b[6]
+ VDD_SW_b[7] VSS_SW_b[1] VSS_SW_b[2] VSS_SW_b[3] VSS_SW_b[4] VSS_SW_b[5] VSS_SW_b[6]
+ VSS_SW_b[7] D[1] VDD_SW[1] ready reset VSS VDD
X0 a_3420_212# x9.X VSS.t258 VSS.t257 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 VSS.t85 VDD.t753 a_10509_601# VSS.t84 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X2 a_11539_1642# VSS.t718 a_11325_1642# VDD.t566 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.193 ps=1.34 w=0.42 l=0.15
X3 VSS.t87 VDD.t754 a_7769_n62# VSS.t86 sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.109 ps=1.03 w=0.42 l=0.15
X4 VDD.t503 a_15293_601# a_16024_909# VDD.t502 sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X5 VSS.t166 a_5812_212# a_5813_n88# VSS.t165 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6 a_5927_n62# a_5812_212# a_5504_106# VSS.t164 sky130_fd_pr__nfet_01v8 ad=0.116 pd=1.09 as=0.0486 ps=0.63 w=0.36 l=0.15
X7 a_5323_2457# x30.A VSS.t632 VSS.t631 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 VDD.t688 x3.X a_939_2457# VDD.t687 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_5271_n62# x2.X.t32 VSS.t112 VSS.t111 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X10 a_13300_993# a_11987_627# a_13216_993# VDD.t585 sky130_fd_pr__pfet_01v8_hvt ad=0.0787 pd=0.795 as=0.0567 ps=0.69 w=0.42 l=0.15
X11 VDD.t149 VDD.t147 a_10509_601# VDD.t148 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.17 ps=1.81 w=0.64 l=0.15
X12 VDD.t617 x16.X a_11987_627# VDD.t616 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X13 a_14887_1642# x9.A1.t32 a_14428_1467# VDD.t34 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X14 a_7896_106# a_8205_n88# a_8140_n62# VSS.t110 sky130_fd_pr__nfet_01v8 ad=0.0486 pd=0.63 as=0.066 ps=0.745 w=0.36 l=0.15
X15 VSS.t441 a_9742_n88# VSS_SW_b[3].t1 VSS.t440 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X16 VSS.t347 a_14857_1289# a_14791_1315# VSS.t346 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X17 VDD.t280 a_1415_895# a_2136_627# VDD.t279 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X18 VDD.t238 a_8591_895# a_8516_993# VDD.t237 sky130_fd_pr__pfet_01v8_hvt ad=0.0956 pd=0.875 as=0.0787 ps=0.795 w=0.42 l=0.15
X19 x7.X a_1757_1642# VSS.t662 VSS.t661 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.113 ps=1.04 w=0.65 l=0.15
X20 a_1501_122# a_1029_n88# a_1745_304# VDD.t474 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X21 a_8933_1642# x9.A1.t33 a_8861_1642# VDD.t35 sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X22 a_8933_1315# a_8679_1642# VSS.t306 VSS.t305 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.145 ps=1.11 w=0.42 l=0.15
X23 a_9154_1315# x9.A1.t34 a_8933_1642# VSS.t195 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X24 VSS.t364 D[6].t0 a_4338_n62# VSS.t363 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X25 VDD.t218 check[1].t0 a_13461_1642# VDD.t217 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.118 ps=1.4 w=0.42 l=0.15
X26 a_10983_895# a_10824_993# a_11123_627# VSS.t19 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.109 ps=1.03 w=0.64 l=0.15
X27 VSS.t160 check[1].t1 a_13461_1642# VSS.t159 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.109 ps=1.36 w=0.42 l=0.15
X28 VDD.t216 D[2].t0 a_13906_n62# VDD.t215 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X29 a_16298_n62# a_15381_n88# a_15853_122# VSS.t656 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0675 ps=0.735 w=0.36 l=0.15
X30 a_15518_304# a_15381_n88# a_15072_106# VDD.t691 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X31 VDD_SW_b[6].t0 a_3807_895# VDD.t354 VDD.t353 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X32 a_8731_627# a_8117_601# a_8591_895# VSS.t664 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X33 a_10041_993# a_9595_627# a_9949_627# VDD.t266 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0651 ps=0.73 w=0.42 l=0.15
X34 a_5462_220# a_5271_n62# VDD.t494 VDD.t493 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X35 VSS.t582 x16.X a_11987_627# VSS.t581 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X36 x9.A1.t31 a_5323_2457# VSS.t506 VSS.t505 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X37 a_15608_993# a_14545_627# a_15464_909# VDD.t638 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X38 a_9949_627# D[3].t0 VDD.t75 VDD.t74 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X39 VDD.t245 a_76_1467# x6.X VDD.t244 sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X40 VDD.t501 a_15293_601# a_15243_909# VDD.t500 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X41 a_8545_n62# a_8677_122# a_8409_n88# VSS.t637 sky130_fd_pr__nfet_01v8 ad=0.0974 pd=0.97 as=0.0864 ps=0.91 w=0.64 l=0.15
X42 a_11325_1642# x9.A1.t35 a_11253_1642# VDD.t255 sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X43 VDD.t719 a_12134_n88# VSS_SW_b[2].t0 VDD.t718 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X44 a_15585_n88# a_15853_122# a_15799_220# VDD.t600 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X45 a_11325_1315# a_11071_1642# VSS.t567 VSS.t566 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.145 ps=1.11 w=0.42 l=0.15
X46 VDD.t206 a_13193_n88# a_13126_304# VDD.t205 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X47 VDD.t663 x30.A a_5323_2457# VDD.t662 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X48 a_10532_n62# a_9742_n88# VSS.t439 VSS.t438 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0703 ps=0.755 w=0.42 l=0.15
X49 a_1028_212# x7.X VSS.t284 VSS.t283 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X50 a_5319_1642# x9.A1.t36 a_4860_1467# VDD.t256 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X51 a_10801_n88# a_10055_n62# a_10937_n62# VSS.t49 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X52 a_8921_304# a_8409_n88# VDD.t303 VDD.t302 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X53 VSS.t92 a_3420_212# a_3421_n88# VSS.t91 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X54 VSS.t427 a_5289_1289# a_5223_1315# VSS.t426 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X55 a_3807_895# x2.X.t33 VDD.t169 VDD.t168 sky130_fd_pr__pfet_01v8_hvt ad=0.132 pd=1.22 as=0.0956 ps=0.875 w=0.42 l=0.15
X56 a_15380_212# x20.X VSS.t609 VSS.t608 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X57 VSS.t141 a_7823_601# a_7757_627# VSS.t140 sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0671 ps=0.75 w=0.42 l=0.15
X58 a_2773_627# D[6].t1 VSS.t366 VSS.t365 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X59 a_12433_993# a_12153_627# a_12341_627# VSS.t83 sky130_fd_pr__nfet_01v8 ad=0.0675 pd=0.735 as=0.066 ps=0.745 w=0.36 l=0.15
X60 VDD.t298 check[4].t0 a_6753_1642# VDD.t297 sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.0767 ps=0.785 w=0.42 l=0.15
X61 VSS.t658 VDD.t755 a_8545_n62# VSS.t657 sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0974 ps=0.97 w=0.42 l=0.15
X62 a_12134_n88# a_12680_106# a_12638_220# VDD.t310 sky130_fd_pr__pfet_01v8_hvt ad=0.132 pd=1.22 as=0.0882 ps=1.05 w=0.84 l=0.15
X63 VSS.t230 check[4].t1 a_6760_1315# VSS.t229 sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.0693 ps=0.75 w=0.42 l=0.15
X64 VSS.t451 a_305_2457# x3.X VSS.t450 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X65 VDD.t372 a_12607_601# a_12517_993# VDD.t371 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X66 a_6753_1642# VSS.t719 a_6539_1642# VDD.t565 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.193 ps=1.34 w=0.42 l=0.15
X67 a_7757_627# a_7203_627# a_7649_993# VSS.t674 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0675 ps=0.735 w=0.36 l=0.15
X68 VDD_SW[4].t1 a_9312_627# VSS.t5 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X69 VSS.t660 VDD.t756 a_8117_601# VSS.t659 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X70 VSS.t653 x3.X a_939_2457# VSS.t652 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X71 a_2927_1642# x9.A1.t37 a_2468_1467# VDD.t453 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X72 a_4862_90# a_4958_n88# VDD.t65 VDD.t64 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X73 VDD.t464 a_13375_895# a_14096_627# VDD.t463 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X74 VSS.t69 D[7].t0 a_1946_n62# VSS.t68 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X75 a_487_n62# x2.X.t34 VSS.t465 VSS.t464 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X76 x30.A a_4689_2457# VDD.t159 VDD.t158 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X77 VDD.t546 a_5323_2457# x9.A1.t15 VDD.t545 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X78 x9.A1.t30 a_5323_2457# VSS.t504 VSS.t503 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X79 VSS.t557 a_2897_1289# a_2831_1315# VSS.t556 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X80 VDD.t79 check[3].t0 a_8679_1642# VDD.t78 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.118 ps=1.4 w=0.42 l=0.15
X81 VDD.t146 VDD.t144 a_1233_n88# VDD.t145 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X82 VDD.t247 a_7681_1289# a_7711_1642# VDD.t246 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X83 VSS.t77 check[3].t1 a_8679_1642# VSS.t76 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.109 ps=1.36 w=0.42 l=0.15
X84 VDD.t602 check[0].t0 a_16323_1642# VDD.t601 sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.0767 ps=0.785 w=0.42 l=0.15
X85 VSS.t706 VDD.t757 a_941_601# VSS.t705 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X86 VSS.t570 check[0].t1 a_16330_1315# VSS.t569 sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.0693 ps=0.75 w=0.42 l=0.15
X87 a_6730_n62# a_5813_n88# a_6285_122# VSS.t412 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0675 ps=0.735 w=0.36 l=0.15
X88 a_10596_212# x15.X VDD.t191 VDD.t190 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X89 a_5950_304# a_5813_n88# a_5504_106# VDD.t452 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X90 a_15143_627# a_15293_601# a_14999_601# VSS.t463 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X91 a_3732_993# a_2419_627# a_3648_993# VDD.t183 sky130_fd_pr__pfet_01v8_hvt ad=0.0787 pd=0.795 as=0.0567 ps=0.69 w=0.42 l=0.15
X92 a_13126_304# a_12989_n88# a_12680_106# VDD.t395 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X93 VSS.t400 a_939_2457# x2.X.t31 VSS.t399 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X94 a_16323_1642# VSS.t720 a_16109_1642# VDD.t564 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.193 ps=1.34 w=0.42 l=0.15
X95 VDD.t143 VDD.t141 a_941_601# VDD.t142 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.17 ps=1.81 w=0.64 l=0.15
X96 a_3070_220# a_2879_n62# VDD.t622 VDD.t621 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X97 VDD.t574 reset.t0 a_29_2457# VDD.t573 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X98 a_13216_993# a_12153_627# a_13072_909# VDD.t81 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X99 a_7557_627# D[4].t0 VDD.t338 VDD.t337 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X100 VSS.t641 a_14428_1467# x18.X VSS.t640 sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X101 a_14945_n62# a_15072_106# a_14526_n88# VSS.t617 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.03 as=0.0864 ps=0.91 w=0.64 l=0.15
X102 x9.A1.t29 a_5323_2457# VSS.t502 VSS.t501 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X103 VSS.t178 a_8591_895# a_8539_627# VSS.t177 sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.066 ps=0.745 w=0.42 l=0.15
X104 VDD.t189 a_6199_895# a_6124_993# VDD.t188 sky130_fd_pr__pfet_01v8_hvt ad=0.0956 pd=0.875 as=0.0787 ps=0.795 w=0.42 l=0.15
X105 VSS.t601 a_7350_n88# VSS_SW_b[4].t1 VSS.t600 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X106 VDD_SW_b[1].t0 a_15767_895# VDD.t316 VDD.t315 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X107 VSS.t235 a_8409_n88# a_8319_n62# VSS.t234 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.116 ps=1.09 w=0.64 l=0.15
X108 a_13193_n88# a_13461_122# a_13407_220# VDD.t744 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X109 VDD.t661 x30.A a_5323_2457# VDD.t660 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X110 VSS.t398 a_939_2457# x2.X.t30 VSS.t397 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X111 a_678_220# a_487_n62# VDD.t729 VDD.t728 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X112 a_1415_895# x2.X.t35 VDD.t505 VDD.t504 sky130_fd_pr__pfet_01v8_hvt ad=0.132 pd=1.22 as=0.0956 ps=0.875 w=0.42 l=0.15
X113 VDD.t140 VDD.t138 a_8117_601# VDD.t139 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.17 ps=1.81 w=0.64 l=0.15
X114 a_9644_1467# VSS.t721 a_9786_1642# VDD.t563 sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X115 a_12937_304# a_12134_n88# VDD.t717 VDD.t716 sky130_fd_pr__pfet_01v8_hvt ad=0.0787 pd=0.795 as=0.0956 ps=0.875 w=0.42 l=0.15
X116 a_4862_90# a_4958_n88# VSS.t63 VSS.t62 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X117 a_12988_212# x17.X VSS.t304 VSS.t303 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X118 VSS.t433 a_10983_895# a_11704_627# VSS.t432 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X119 VSS.t555 a_5431_601# a_5365_627# VSS.t554 sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0671 ps=0.75 w=0.42 l=0.15
X120 a_15495_n62# a_15380_212# a_15072_106# VSS.t182 sky130_fd_pr__nfet_01v8 ad=0.116 pd=1.09 as=0.0486 ps=0.63 w=0.36 l=0.15
X121 VSS.t181 a_15380_212# a_15381_n88# VSS.t180 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X122 VDD.t77 D[3].t1 a_11514_n62# VDD.t76 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X123 a_10041_993# a_9761_627# a_9949_627# VSS.t443 sky130_fd_pr__nfet_01v8 ad=0.0675 pd=0.735 as=0.066 ps=0.745 w=0.36 l=0.15
X124 VSS.t708 VDD.t758 a_6153_n62# VSS.t707 sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0974 ps=0.97 w=0.42 l=0.15
X125 VDD.t624 a_9644_1467# x14.X VDD.t623 sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X126 a_9786_1642# check[2].t0 VDD.t444 VDD.t443 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X127 VDD.t393 a_14857_1289# a_14887_1642# VDD.t392 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X128 x2.X.t15 a_939_2457# VDD.t440 VDD.t439 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X129 a_9786_1315# check[2].t1 VSS.t404 VSS.t403 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X130 x17.X a_13715_1642# VDD.t268 VDD.t267 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.158 ps=1.39 w=1 l=0.15
X131 VDD.t364 a_10215_601# a_10125_993# VDD.t363 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X132 a_7769_n62# a_7896_106# a_7350_n88# VSS.t654 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.03 as=0.0864 ps=0.91 w=0.64 l=0.15
X133 a_939_2457# x3.X VDD.t686 VDD.t685 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X134 VDD.t290 a_5725_601# a_5675_909# VDD.t289 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X135 a_5365_627# a_4811_627# a_5257_993# VSS.t270 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0675 ps=0.735 w=0.36 l=0.15
X136 VDD_SW[5].t1 a_6920_627# VSS.t199 VSS.t198 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X137 a_8140_n62# a_7350_n88# VSS.t599 VSS.t598 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0703 ps=0.755 w=0.42 l=0.15
X138 a_14733_627# D[1].t0 VSS.t57 VSS.t56 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X139 VDD.t544 a_5323_2457# x9.A1.t14 VDD.t543 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X140 a_6153_n62# a_6285_122# a_6017_n88# VSS.t419 sky130_fd_pr__nfet_01v8 ad=0.0974 pd=0.97 as=0.0864 ps=0.91 w=0.64 l=0.15
X141 VSS.t282 x3.A a_305_2457# VSS.t281 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X142 a_2470_90# a_2566_n88# VDD.t214 VDD.t213 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X143 a_8409_n88# a_7663_n62# a_8545_n62# VSS.t360 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X144 VSS.t158 D[2].t1 a_13906_n62# VSS.t157 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X145 a_11069_122# a_10597_n88# a_11313_304# VDD.t73 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X146 a_76_1467# x9.A1.t38 a_218_1315# VSS.t413 sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X147 a_15799_220# a_14839_n62# VDD.t7 VDD.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X148 x9.A1.t28 a_5323_2457# VSS.t500 VSS.t499 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X149 VDD.t230 a_3333_601# a_4064_909# VDD.t229 sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X150 a_10931_627# a_9761_627# a_10824_993# VSS.t442 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0486 ps=0.63 w=0.36 l=0.15
X151 a_6529_304# a_6017_n88# VDD.t752 VDD.t751 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X152 VSS.t694 a_1028_212# a_1029_n88# VSS.t693 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X153 a_7615_1315# VSS.t539 a_7252_1467# VSS.t540 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X154 a_1340_993# a_27_627# a_1256_993# VDD.t552 sky130_fd_pr__pfet_01v8_hvt ad=0.0787 pd=0.795 as=0.0567 ps=0.69 w=0.42 l=0.15
X155 VDD.t542 a_5323_2457# x9.A1.t13 VDD.t541 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X156 a_1978_1315# x9.A1.t39 a_1757_1642# VSS.t414 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X157 a_12036_1467# VSS.t722 a_12178_1642# VDD.t562 sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X158 a_5165_627# D[5].t0 VDD.t570 VDD.t569 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X159 x2.X.t14 a_939_2457# VDD.t438 VDD.t437 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X160 VSS.t396 a_939_2457# x2.X.t29 VSS.t395 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X161 VDD_SW[6].t0 a_4528_627# VDD.t37 VDD.t36 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X162 VSS.t133 a_6199_895# a_6147_627# VSS.t132 sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.066 ps=0.745 w=0.42 l=0.15
X163 a_9742_n88# a_10288_106# a_10246_220# VDD.t325 sky130_fd_pr__pfet_01v8_hvt ad=0.132 pd=1.22 as=0.0882 ps=1.05 w=0.84 l=0.15
X164 a_15030_220# a_14839_n62# VDD.t5 VDD.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X165 VSS.t61 a_4958_n88# VSS_SW_b[5].t1 VSS.t60 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X166 VSS.t114 reset.t1 a_29_2457# VSS.t113 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X167 VDD.t137 VDD.t135 a_14526_n88# VDD.t136 sky130_fd_pr__pfet_01v8_hvt ad=0.0956 pd=0.875 as=0.132 ps=1.22 w=0.42 l=0.15
X168 VSS.t717 a_6017_n88# a_5927_n62# VSS.t716 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.116 ps=1.09 w=0.64 l=0.15
X169 a_8335_627# a_7823_601# VSS.t139 VSS.t138 sky130_fd_pr__nfet_01v8 ad=0.116 pd=1.09 as=0.166 ps=1.8 w=0.64 l=0.15
X170 a_8921_n62# a_8409_n88# VSS.t233 VSS.t232 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0882 ps=0.84 w=0.42 l=0.15
X171 x9.A1.t27 a_5323_2457# VSS.t498 VSS.t497 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X172 a_13715_1642# x9.A1.t40 a_13643_1642# VDD.t618 sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X173 VSS.t211 a_2468_1467# x8.X VSS.t210 sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X174 a_13715_1315# a_13461_1642# VSS.t474 VSS.t473 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.145 ps=1.11 w=0.42 l=0.15
X175 a_8848_909# a_8432_993# a_8591_895# VDD.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.132 ps=1.22 w=0.84 l=0.15
X176 a_10545_304# a_9742_n88# VDD.t480 VDD.t479 sky130_fd_pr__pfet_01v8_hvt ad=0.0787 pd=0.795 as=0.0956 ps=0.875 w=0.42 l=0.15
X177 a_2470_90# a_2566_n88# VSS.t156 VSS.t155 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X178 VDD.t659 x30.A a_5323_2457# VDD.t658 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X179 VSS.t394 a_939_2457# x2.X.t28 VSS.t393 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X180 VDD.t701 a_941_601# a_891_909# VDD.t700 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X181 a_581_627# a_27_627# a_473_993# VSS.t512 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0675 ps=0.735 w=0.36 l=0.15
X182 a_4338_n62# a_3421_n88# a_3893_122# VSS.t194 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0675 ps=0.735 w=0.36 l=0.15
X183 x9.A1.t26 a_5323_2457# VSS.t496 VSS.t495 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X184 a_5575_627# a_5725_601# a_5431_601# VSS.t222 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X185 a_13103_n62# a_12988_212# a_12680_106# VSS.t192 sky130_fd_pr__nfet_01v8 ad=0.116 pd=1.09 as=0.0486 ps=0.63 w=0.36 l=0.15
X186 a_3558_304# a_3421_n88# a_3112_106# VDD.t254 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X187 VDD.t296 a_10596_212# a_10597_n88# VDD.t295 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X188 a_15072_106# a_15381_n88# a_15316_n62# VSS.t655 sky130_fd_pr__nfet_01v8 ad=0.0486 pd=0.63 as=0.066 ps=0.745 w=0.36 l=0.15
X189 x3.X a_305_2457# VDD.t490 VDD.t489 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X190 a_3648_993# a_2585_627# a_3504_909# VDD.t193 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X191 a_8677_122# a_8204_212# a_8921_n62# VSS.t565 sky130_fd_pr__nfet_01v8 ad=0.0675 pd=0.735 as=0.0671 ps=0.75 w=0.36 l=0.15
X192 a_5504_106# a_5812_212# a_5761_304# VDD.t224 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0787 ps=0.795 w=0.42 l=0.15
X193 VSS.t150 a_12036_1467# x16.X VSS.t149 sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X194 a_5377_n62# a_5504_106# a_4958_n88# VSS.t319 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.03 as=0.0864 ps=0.91 w=0.64 l=0.15
X195 a_12341_627# D[2].t2 VSS.t65 VSS.t64 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X196 a_939_2457# x3.X VDD.t684 VDD.t683 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X197 VDD.t228 a_3333_601# a_3283_909# VDD.t227 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X198 a_7350_n88# a_7663_n62# a_7769_n62# VSS.t359 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X199 a_5675_909# a_5257_993# a_5431_601# VDD.t735 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X200 a_7967_627# x2.X.t36 VSS.t467 VSS.t466 sky130_fd_pr__nfet_01v8 ad=0.0974 pd=0.97 as=0.0882 ps=0.84 w=0.42 l=0.15
X201 VDD.t540 a_5323_2457# x9.A1.t12 VDD.t539 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X202 VDD.t591 a_2897_1289# a_2927_1642# VDD.t590 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X203 a_10801_n88# a_11069_122# a_11015_220# VDD.t248 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X204 VDD.t538 a_5323_2457# x9.A1.t11 VDD.t537 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X205 a_9761_627# a_9595_627# VDD.t265 VDD.t264 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X206 a_13407_220# a_12447_n62# VDD.t348 VDD.t347 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X207 a_381_627# D[7].t1 VDD.t71 VDD.t70 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X208 VSS.t580 a_647_601# a_581_627# VSS.t579 sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0671 ps=0.75 w=0.42 l=0.15
X209 VSS.t176 a_8591_895# a_9312_627# VSS.t175 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X210 VDD.t406 check[2].t2 a_11539_1642# VDD.t405 sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.0767 ps=0.785 w=0.42 l=0.15
X211 a_14430_90# a_14526_n88# VDD.t47 VDD.t46 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X212 a_8204_212# x13.X VDD.t258 VDD.t257 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X213 VDD.t340 D[4].t1 a_9122_n62# VDD.t339 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X214 VSS.t362 check[2].t3 a_11546_1315# VSS.t361 sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.0693 ps=0.75 w=0.42 l=0.15
X215 VSS.t27 VDD.t759 a_14945_n62# VSS.t26 sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.109 ps=1.03 w=0.42 l=0.15
X216 VSS.t245 a_174_n88# VSS_SW_b[7].t1 VSS.t244 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X217 VSS.t576 a_3039_601# a_2973_627# VSS.t575 sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0671 ps=0.75 w=0.42 l=0.15
X218 x13.X a_8933_1642# VSS.t14 VSS.t13 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.113 ps=1.04 w=0.65 l=0.15
X219 VSS.t191 a_12988_212# a_12989_n88# VSS.t190 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X220 VDD.t536 a_5323_2457# x9.A1.t10 VDD.t535 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X221 VSS.t449 a_305_2457# x3.X VSS.t448 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X222 VDD_SW[7].t0 a_2136_627# VDD.t446 VDD.t445 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X223 VDD_SW_b[5].t1 a_6199_895# VSS.t131 VSS.t130 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X224 VDD.t134 VDD.t132 a_4958_n88# VDD.t133 sky130_fd_pr__pfet_01v8_hvt ad=0.0956 pd=0.875 as=0.132 ps=1.22 w=0.42 l=0.15
X225 a_8677_122# a_8205_n88# a_8921_304# VDD.t167 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X226 VSS.t392 a_939_2457# x2.X.t27 VSS.t391 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X227 a_16037_1642# a_15855_1642# VDD.t324 VDD.t323 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X228 a_14857_1289# check[0].t2 VDD.t640 VDD.t639 sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X229 VDD_SW[1].t0 a_16488_627# VDD.t15 VDD.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X230 x30.A a_4689_2457# VDD.t157 VDD.t156 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X231 a_791_627# a_941_601# a_647_601# VSS.t666 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X232 x2.X.t13 a_939_2457# VDD.t436 VDD.t435 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X233 a_14857_1289# check[0].t3 VSS.t607 VSS.t606 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X234 a_4149_1642# VSS.t537 a_4149_1315# VSS.t538 sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X235 x20.X a_16109_1642# VDD.t232 VDD.t231 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.158 ps=1.39 w=1 l=0.15
X236 a_7823_601# x2.X.t37 VDD.t379 VDD.t378 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X237 a_9761_627# a_9595_627# VSS.t205 VSS.t204 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X238 a_6456_909# a_6040_993# a_6199_895# VDD.t651 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.132 ps=1.22 w=0.84 l=0.15
X239 VSS.t349 D[3].t2 a_11514_n62# VSS.t348 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X240 x9.A1.t25 a_5323_2457# VSS.t494 VSS.t493 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X241 a_8731_627# x2.X.t38 VSS.t329 VSS.t328 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.03 as=0.0703 ps=0.755 w=0.42 l=0.15
X242 a_891_909# a_473_993# a_647_601# VDD.t82 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X243 a_3183_627# a_3333_601# a_3039_601# VSS.t170 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X244 a_10824_993# a_9595_627# a_10727_627# VSS.t203 sky130_fd_pr__nfet_01v8 ad=0.0486 pd=0.63 as=0.116 ps=1.09 w=0.36 l=0.15
X245 VSS.t390 a_939_2457# x2.X.t26 VSS.t389 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X246 a_1166_304# a_1029_n88# a_720_106# VDD.t473 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X247 a_10983_895# x2.X.t39 VDD.t381 VDD.t380 sky130_fd_pr__pfet_01v8_hvt ad=0.132 pd=1.22 as=0.0956 ps=0.875 w=0.42 l=0.15
X248 a_5431_601# a_5257_993# a_5575_627# VSS.t696 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.0974 ps=0.97 w=0.64 l=0.15
X249 a_14430_90# a_14526_n88# VSS.t47 VSS.t46 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X250 VDD.t334 a_9646_90# VSS_SW[3].t0 VDD.t333 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X251 a_1256_993# a_193_627# a_1112_909# VDD.t725 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X252 a_6285_122# a_5812_212# a_6529_n62# VSS.t163 sky130_fd_pr__nfet_01v8 ad=0.0675 pd=0.735 as=0.0671 ps=0.75 w=0.36 l=0.15
X253 VSS.t51 a_4862_90# VSS_SW[5].t1 VSS.t50 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X254 a_3112_106# a_3420_212# a_3369_304# VDD.t86 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0787 ps=0.795 w=0.42 l=0.15
X255 VSS.t201 x27.A a_4689_2457# VSS.t200 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X256 a_12465_1289# check[1].t2 VDD.t383 VDD.t382 sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X257 a_2985_n62# a_3112_106# a_2566_n88# VSS.t695 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.03 as=0.0864 ps=0.91 w=0.64 l=0.15
X258 VDD.t646 check[6].t0 a_1971_1642# VDD.t645 sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.0767 ps=0.785 w=0.42 l=0.15
X259 a_7252_1467# x9.A1.t41 a_7394_1315# VSS.t583 sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X260 a_12465_1289# check[1].t3 VSS.t337 VSS.t336 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X261 a_5896_909# a_5431_601# VDD.t589 VDD.t588 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X262 a_15907_627# a_15293_601# a_15767_895# VSS.t462 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X263 a_1757_1642# VSS.t535 a_1757_1315# VSS.t536 sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X264 VSS.t615 check[6].t1 a_1978_1315# VSS.t614 sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.0693 ps=0.75 w=0.42 l=0.15
X265 a_3283_909# a_2865_993# a_3039_601# VDD.t512 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X266 a_5575_627# x2.X.t40 VSS.t469 VSS.t468 sky130_fd_pr__nfet_01v8 ad=0.0974 pd=0.97 as=0.0882 ps=0.84 w=0.42 l=0.15
X267 a_1233_n88# a_1501_122# a_1447_220# VDD.t400 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X268 a_939_2457# x3.X VDD.t682 VDD.t681 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X269 a_6529_n62# a_6017_n88# VSS.t715 VSS.t714 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0882 ps=0.84 w=0.42 l=0.15
X270 a_8153_304# a_7350_n88# VDD.t634 VDD.t633 sky130_fd_pr__pfet_01v8_hvt ad=0.0787 pd=0.795 as=0.0956 ps=0.875 w=0.42 l=0.15
X271 VSS.t388 a_939_2457# x2.X.t25 VSS.t387 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X272 a_8539_627# a_7369_627# a_8432_993# VSS.t168 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0486 ps=0.63 w=0.36 l=0.15
X273 a_12038_90# a_12134_n88# VDD.t715 VDD.t714 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X274 a_7733_993# a_7369_627# a_7649_993# VDD.t226 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X275 a_5812_212# x11.X VDD.t548 VDD.t547 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X276 VSS.t29 VDD.t760 a_5377_n62# VSS.t28 sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.109 ps=1.03 w=0.42 l=0.15
X277 VDD.t202 a_12901_601# a_13632_909# VDD.t201 sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X278 VDD.t597 a_8204_212# a_8205_n88# VDD.t596 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X279 a_593_n62# a_720_106# a_174_n88# VSS.t142 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.03 as=0.0864 ps=0.91 w=0.64 l=0.15
X280 a_2831_1315# VSS.t533 a_2468_1467# VSS.t534 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X281 VDD.t327 ready.t0 a_4413_2457# VDD.t326 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X282 a_3535_n62# a_3420_212# a_3112_106# VSS.t90 sky130_fd_pr__nfet_01v8 ad=0.116 pd=1.09 as=0.0486 ps=0.63 w=0.36 l=0.15
X283 x2.X.t12 a_939_2457# VDD.t434 VDD.t433 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X284 a_16097_304# a_15585_n88# VDD.t667 VDD.t666 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X285 VSS.t713 a_14999_601# a_14933_627# VSS.t712 sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0671 ps=0.75 w=0.42 l=0.15
X286 a_5504_106# a_5813_n88# a_5748_n62# VSS.t411 sky130_fd_pr__nfet_01v8 ad=0.0486 pd=0.63 as=0.066 ps=0.745 w=0.36 l=0.15
X287 VDD_SW_b[6].t1 a_3807_895# VSS.t292 VSS.t291 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X288 a_16330_1315# x9.A1.t42 a_16109_1642# VSS.t584 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X289 a_7663_n62# x2.X.t41 VDD.t507 VDD.t506 sky130_fd_pr__pfet_01v8_hvt ad=0.17 pd=1.81 as=0.154 ps=1.34 w=0.64 l=0.15
X290 VSS.t252 a_15767_895# a_15715_627# VSS.t251 sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.066 ps=0.745 w=0.42 l=0.15
X291 VDD.t534 a_5323_2457# x9.A1.t9 VDD.t533 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X292 a_5323_2457# x30.A VSS.t630 VSS.t629 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X293 VDD.t131 VDD.t129 a_8409_n88# VDD.t130 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X294 VSS.t636 a_15585_n88# a_15495_n62# VSS.t635 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.116 ps=1.09 w=0.64 l=0.15
X295 VSS.t185 a_76_1467# x6.X VSS.t184 sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X296 a_4958_n88# a_5271_n62# a_5377_n62# VSS.t453 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X297 VDD_SW[2].t0 a_14096_627# VDD.t713 VDD.t712 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X298 a_5431_601# x2.X.t42 VDD.t509 VDD.t508 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X299 a_4064_909# a_3648_993# a_3807_895# VDD.t299 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.132 ps=1.22 w=0.84 l=0.15
X300 a_3839_220# a_2879_n62# VDD.t620 VDD.t619 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X301 x2.X.t11 a_939_2457# VDD.t432 VDD.t431 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X302 a_4077_1642# a_3895_1642# VDD.t220 VDD.t219 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X303 a_7369_627# a_7203_627# VDD.t709 VDD.t708 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X304 a_14428_1467# x9.A1.t43 a_14570_1315# VSS.t458 sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X305 a_2897_1289# check[5].t0 VDD.t397 VDD.t396 sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X306 VDD.t450 x14.X a_9595_627# VDD.t449 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X307 VDD.t128 VDD.t126 a_174_n88# VDD.t127 sky130_fd_pr__pfet_01v8_hvt ad=0.0956 pd=0.875 as=0.132 ps=1.22 w=0.42 l=0.15
X308 VDD.t532 a_5323_2457# x9.A1.t8 VDD.t531 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X309 x9.A1.t24 a_5323_2457# VSS.t492 VSS.t491 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X310 a_2897_1289# check[5].t1 VSS.t355 VSS.t354 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X311 a_791_627# x2.X.t43 VSS.t331 VSS.t330 sky130_fd_pr__nfet_01v8 ad=0.0974 pd=0.97 as=0.0882 ps=0.84 w=0.42 l=0.15
X312 a_13906_n62# a_12989_n88# a_13461_122# VSS.t353 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0675 ps=0.735 w=0.36 l=0.15
X313 x9.X a_4149_1642# VDD.t408 VDD.t407 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.158 ps=1.39 w=1 l=0.15
X314 a_10908_993# a_9595_627# a_10824_993# VDD.t263 sky130_fd_pr__pfet_01v8_hvt ad=0.0787 pd=0.795 as=0.0567 ps=0.69 w=0.42 l=0.15
X315 a_12038_90# a_12134_n88# VSS.t684 VSS.t683 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X316 VDD.t650 a_7254_90# VSS_SW[4].t0 VDD.t649 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X317 a_2879_n62# x2.X.t44 VSS.t333 VSS.t332 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X318 a_720_106# a_1028_212# a_977_304# VDD.t733 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0787 ps=0.795 w=0.42 l=0.15
X319 VSS.t298 a_2470_90# VSS_SW[6].t1 VSS.t297 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X320 VDD_SW_b[7].t0 a_1415_895# VDD.t278 VDD.t277 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X321 a_6339_627# a_5725_601# a_6199_895# VSS.t221 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X322 a_3504_909# a_3039_601# VDD.t611 VDD.t610 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X323 VDD.t125 VDD.t123 a_2566_n88# VDD.t124 sky130_fd_pr__pfet_01v8_hvt ad=0.0956 pd=0.875 as=0.132 ps=1.22 w=0.42 l=0.15
X324 a_3183_627# x2.X.t45 VSS.t335 VSS.t334 sky130_fd_pr__nfet_01v8 ad=0.0974 pd=0.97 as=0.0882 ps=0.84 w=0.42 l=0.15
X325 a_15072_106# a_15380_212# a_15329_304# VDD.t242 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0787 ps=0.795 w=0.42 l=0.15
X326 VSS.t325 D[4].t2 a_9122_n62# VSS.t324 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X327 VSS.t386 a_939_2457# x2.X.t24 VSS.t385 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X328 a_12495_1642# x9.A1.t44 a_12036_1467# VDD.t497 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X329 a_1685_1642# a_1503_1642# VDD.t11 VDD.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X330 VSS.t471 a_12465_1289# a_12399_1315# VSS.t470 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X331 a_6147_627# a_4977_627# a_6040_993# VSS.t294 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0486 ps=0.63 w=0.36 l=0.15
X332 a_15243_909# a_14825_993# a_14999_601# VDD.t581 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X333 a_218_1642# check[6].t2 VDD.t743 VDD.t742 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X334 a_647_601# a_473_993# a_791_627# VSS.t88 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.0974 ps=0.97 w=0.64 l=0.15
X335 a_5341_993# a_4977_627# a_5257_993# VDD.t356 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X336 a_7369_627# a_7203_627# VSS.t673 VSS.t672 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X337 a_8432_993# a_7203_627# a_8335_627# VSS.t671 sky130_fd_pr__nfet_01v8 ad=0.0486 pd=0.63 as=0.116 ps=1.09 w=0.36 l=0.15
X338 VDD.t286 a_10509_601# a_11240_909# VDD.t285 sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X339 a_218_1315# check[6].t3 VSS.t704 VSS.t703 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X340 VSS.t410 x14.X a_9595_627# VSS.t409 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X341 a_13929_1642# VSS.t723 a_13715_1642# VDD.t561 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.193 ps=1.34 w=0.42 l=0.15
X342 a_1143_n62# a_1028_212# a_720_106# VSS.t692 sky130_fd_pr__nfet_01v8 ad=0.116 pd=1.09 as=0.0486 ps=0.63 w=0.36 l=0.15
X343 a_174_n88# a_487_n62# a_593_n62# VSS.t690 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X344 a_6339_627# x2.X.t46 VSS.t23 VSS.t22 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.03 as=0.0703 ps=0.755 w=0.42 l=0.15
X345 a_3112_106# a_3421_n88# a_3356_n62# VSS.t193 sky130_fd_pr__nfet_01v8 ad=0.0486 pd=0.63 as=0.066 ps=0.745 w=0.36 l=0.15
X346 a_647_601# x2.X.t47 VDD.t29 VDD.t28 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X347 a_3039_601# a_2865_993# a_3183_627# VSS.t472 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.0974 ps=0.97 w=0.64 l=0.15
X348 VDD.t478 a_9742_n88# VSS_SW_b[3].t0 VDD.t477 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X349 VSS.t611 ready.t1 a_4413_2457# VSS.t610 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X350 a_16298_n62# a_15380_212# a_15853_122# VDD.t241 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.0567 ps=0.69 w=0.42 l=0.15
X351 a_5271_n62# x2.X.t48 VDD.t31 VDD.t30 sky130_fd_pr__pfet_01v8_hvt ad=0.17 pd=1.81 as=0.154 ps=1.34 w=0.64 l=0.15
X352 VSS.t148 a_13193_n88# a_13103_n62# VSS.t147 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.116 ps=1.09 w=0.64 l=0.15
X353 VDD.t122 VDD.t120 a_6017_n88# VDD.t121 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X354 VDD.t175 check[0].t4 a_15855_1642# VDD.t174 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.118 ps=1.4 w=0.42 l=0.15
X355 a_4860_1467# x9.A1.t45 a_5002_1315# VSS.t459 sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X356 VSS.t120 check[0].t5 a_15855_1642# VSS.t119 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.109 ps=1.36 w=0.42 l=0.15
X357 a_15511_627# a_14999_601# VSS.t711 VSS.t710 sky130_fd_pr__nfet_01v8 ad=0.116 pd=1.09 as=0.166 ps=1.8 w=0.64 l=0.15
X358 a_5323_2457# x30.A VSS.t628 VSS.t627 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X359 a_15316_n62# a_14526_n88# VSS.t45 VSS.t44 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0703 ps=0.755 w=0.42 l=0.15
X360 a_2566_n88# a_2879_n62# a_2985_n62# VSS.t586 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X361 VSS.t71 VDD.t761 a_593_n62# VSS.t70 sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.109 ps=1.03 w=0.42 l=0.15
X362 VDD_SW_b[1].t1 a_15767_895# VSS.t250 VSS.t249 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X363 VDD.t472 a_10983_895# a_11704_627# VDD.t471 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X364 a_4370_1315# x9.A1.t46 a_4149_1642# VSS.t589 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X365 a_8591_895# a_8432_993# a_8731_627# VSS.t12 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.109 ps=1.03 w=0.64 l=0.15
X366 a_3039_601# x2.X.t49 VDD.t496 VDD.t495 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X367 x3.X a_305_2457# VSS.t447 VSS.t446 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X368 VDD.t22 a_10801_n88# a_10734_304# VDD.t21 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X369 a_1447_220# a_487_n62# VDD.t727 VDD.t726 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X370 a_16024_909# a_15608_993# a_15767_895# VDD.t647 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.132 ps=1.22 w=0.84 l=0.15
X371 a_6539_1642# VSS.t531 a_6539_1315# VSS.t532 sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X372 VDD.t292 x12.X a_7203_627# VDD.t291 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X373 VSS.t73 VDD.t762 a_2985_n62# VSS.t72 sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.109 ps=1.03 w=0.42 l=0.15
X374 x2.X.t10 a_939_2457# VDD.t430 VDD.t429 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X375 VDD.t155 a_4689_2457# x30.A VDD.t154 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X376 VSS.t651 x3.X a_939_2457# VSS.t650 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X377 a_11514_n62# a_10597_n88# a_11069_122# VSS.t75 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0675 ps=0.735 w=0.36 l=0.15
X378 a_7649_993# a_7203_627# a_7557_627# VDD.t707 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0651 ps=0.73 w=0.42 l=0.15
X379 a_2468_1467# x9.A1.t47 a_2610_1315# VSS.t590 sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X380 a_10824_993# a_9761_627# a_10680_909# VDD.t482 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X381 VSS.t588 a_9644_1467# x14.X VSS.t587 sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X382 a_1112_909# a_647_601# VDD.t615 VDD.t614 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X383 a_14839_n62# x2.X.t50 VSS.t455 VSS.t454 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X384 VSS.t425 a_13375_895# a_13323_627# VSS.t424 sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.066 ps=0.745 w=0.42 l=0.15
X385 VDD_SW_b[2].t0 a_13375_895# VDD.t462 VDD.t461 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X386 x2.X.t23 a_939_2457# VSS.t384 VSS.t383 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X387 x17.X a_13715_1642# VSS.t207 VSS.t206 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.113 ps=1.04 w=0.65 l=0.15
X388 a_16109_1642# VSS.t529 a_16109_1315# VSS.t530 sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X389 a_12680_106# a_12988_212# a_12937_304# VDD.t252 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0787 ps=0.795 w=0.42 l=0.15
X390 VSS.t461 a_14430_90# VSS_SW[1].t1 VSS.t460 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X391 a_15853_122# a_15380_212# a_16097_n62# VSS.t179 sky130_fd_pr__nfet_01v8 ad=0.0675 pd=0.735 as=0.0671 ps=0.75 w=0.36 l=0.15
X392 VSS.t37 VDD.t763 a_5725_601# VSS.t36 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X393 a_15464_909# a_14999_601# VDD.t748 VDD.t747 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X394 a_15143_627# x2.X.t51 VSS.t457 VSS.t456 sky130_fd_pr__nfet_01v8 ad=0.0974 pd=0.97 as=0.0882 ps=0.84 w=0.42 l=0.15
X395 a_6040_993# a_4811_627# a_5943_627# VSS.t269 sky130_fd_pr__nfet_01v8 ad=0.0486 pd=0.63 as=0.116 ps=1.09 w=0.36 l=0.15
X396 a_16097_n62# a_15585_n88# VSS.t634 VSS.t633 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0882 ps=0.84 w=0.42 l=0.15
X397 VSS.t224 x12.X a_7203_627# VSS.t223 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X398 a_8516_993# a_7203_627# a_8432_993# VDD.t706 sky130_fd_pr__pfet_01v8_hvt ad=0.0787 pd=0.795 as=0.0567 ps=0.69 w=0.42 l=0.15
X399 VDD.t119 VDD.t117 a_5725_601# VDD.t118 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.17 ps=1.81 w=0.64 l=0.15
X400 a_10596_212# x15.X VSS.t135 VSS.t134 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X401 a_11546_1315# x9.A1.t48 a_11325_1642# VSS.t591 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X402 VDD.t466 a_5289_1289# a_5319_1642# VDD.t465 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X403 a_5323_2457# x30.A VDD.t657 VDD.t656 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X404 VSS.t39 VDD.t764 a_3761_n62# VSS.t38 sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0974 ps=0.97 w=0.42 l=0.15
X405 VSS.t102 a_4689_2457# x30.A VSS.t101 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X406 a_193_627# a_27_627# VDD.t551 VDD.t550 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X407 a_2973_627# a_2419_627# a_2865_993# VSS.t127 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0675 ps=0.735 w=0.36 l=0.15
X408 VDD_SW[6].t1 a_4528_627# VSS.t31 VSS.t30 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X409 a_12553_n62# a_12680_106# a_12134_n88# VSS.t246 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.03 as=0.0864 ps=0.91 w=0.64 l=0.15
X410 a_557_993# a_193_627# a_473_993# VDD.t724 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X411 a_3947_627# a_3333_601# a_3807_895# VSS.t169 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X412 a_14999_601# a_14825_993# a_15143_627# VSS.t547 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.0974 ps=0.97 w=0.64 l=0.15
X413 a_14526_n88# a_14839_n62# a_14945_n62# VSS.t3 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X414 a_3761_n62# a_3893_122# a_3625_n88# VSS.t183 sky130_fd_pr__nfet_01v8 ad=0.0974 pd=0.97 as=0.0864 ps=0.91 w=0.64 l=0.15
X415 a_6199_895# a_6040_993# a_6339_627# VSS.t620 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.109 ps=1.03 w=0.64 l=0.15
X416 VDD.t173 check[5].t2 a_3895_1642# VDD.t172 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.118 ps=1.4 w=0.42 l=0.15
X417 a_14791_1315# VSS.t527 a_14428_1467# VSS.t528 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X418 a_4149_1642# x9.A1.t49 a_4077_1642# VDD.t604 sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X419 VSS.t118 check[5].t3 a_3895_1642# VSS.t117 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.109 ps=1.36 w=0.42 l=0.15
X420 a_6467_1642# a_6285_1642# VDD.t385 VDD.t384 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X421 VDD.t699 a_941_601# a_1672_909# VDD.t698 sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X422 a_7649_993# a_7369_627# a_7557_627# VSS.t167 sky130_fd_pr__nfet_01v8 ad=0.0675 pd=0.735 as=0.066 ps=0.745 w=0.36 l=0.15
X423 a_6017_n88# a_5271_n62# a_6153_n62# VSS.t452 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X424 a_4149_1315# a_3895_1642# VSS.t162 VSS.t161 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.145 ps=1.11 w=0.42 l=0.15
X425 a_14999_601# x2.X.t52 VDD.t1 VDD.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X426 a_5257_993# a_4811_627# a_5165_627# VDD.t332 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0651 ps=0.73 w=0.42 l=0.15
X427 VSS.t296 a_78_90# VSS_SW[7].t1 VSS.t295 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X428 a_487_n62# x2.X.t53 VDD.t3 VDD.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.17 pd=1.81 as=0.154 ps=1.34 w=0.64 l=0.15
X429 VDD.t197 a_7823_601# a_7733_993# VDD.t196 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X430 x11.X a_6539_1642# VDD.t336 VDD.t335 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.158 ps=1.39 w=1 l=0.15
X431 a_7252_1467# VSS.t724 a_7394_1642# VDD.t560 sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X432 a_2773_627# D[6].t2 VDD.t672 VDD.t671 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X433 a_4137_304# a_3625_n88# VDD.t389 VDD.t388 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X434 a_193_627# a_27_627# VSS.t511 VSS.t510 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X435 VDD.t236 a_8591_895# a_9312_627# VDD.t235 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X436 a_6730_n62# a_5812_212# a_6285_122# VDD.t223 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.0567 ps=0.69 w=0.42 l=0.15
X437 a_720_106# a_1029_n88# a_964_n62# VSS.t435 sky130_fd_pr__nfet_01v8 ad=0.0486 pd=0.63 as=0.066 ps=0.745 w=0.36 l=0.15
X438 VSS.t290 a_3807_895# a_3755_627# VSS.t289 sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.066 ps=0.745 w=0.42 l=0.15
X439 a_12447_n62# x2.X.t54 VSS.t1 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X440 VDD.t632 a_7350_n88# VSS_SW_b[4].t0 VDD.t631 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X441 VSS.t154 a_2566_n88# VSS_SW_b[6].t1 VSS.t153 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X442 x9.A1.t7 a_5323_2457# VDD.t530 VDD.t529 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X443 VDD.t116 VDD.t114 a_12134_n88# VDD.t115 sky130_fd_pr__pfet_01v8_hvt ad=0.0956 pd=0.875 as=0.132 ps=1.22 w=0.42 l=0.15
X444 VSS.t343 a_3625_n88# a_3535_n62# VSS.t342 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.116 ps=1.09 w=0.64 l=0.15
X445 a_15853_122# a_15381_n88# a_16097_304# VDD.t690 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X446 VDD.t301 a_8409_n88# a_8342_304# VDD.t300 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X447 VDD.t55 a_7252_1467# x12.X VDD.t54 sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X448 a_7394_1642# check[3].t2 VDD.t576 VDD.t575 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X449 VDD.t511 a_12465_1289# a_12495_1642# VDD.t510 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X450 a_5943_627# a_5431_601# VSS.t553 VSS.t552 sky130_fd_pr__nfet_01v8 ad=0.116 pd=1.09 as=0.166 ps=1.8 w=0.64 l=0.15
X451 a_13119_627# a_12607_601# VSS.t310 VSS.t309 sky130_fd_pr__nfet_01v8 ad=0.116 pd=1.09 as=0.166 ps=1.8 w=0.64 l=0.15
X452 a_1757_1642# x9.A1.t50 a_1685_1642# VDD.t605 sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X453 a_7394_1315# check[3].t3 VSS.t544 VSS.t543 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X454 a_5748_n62# a_4958_n88# VSS.t59 VSS.t58 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0703 ps=0.755 w=0.42 l=0.15
X455 x2.X.t22 a_939_2457# VSS.t382 VSS.t381 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X456 VSS.t237 VDD.t765 a_3333_601# VSS.t236 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X457 VDD.t314 a_15767_895# a_15692_993# VDD.t313 sky130_fd_pr__pfet_01v8_hvt ad=0.0956 pd=0.875 as=0.0787 ps=0.795 w=0.42 l=0.15
X458 a_13072_909# a_12607_601# VDD.t370 VDD.t369 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X459 a_1757_1315# a_1503_1642# VSS.t7 VSS.t6 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.145 ps=1.11 w=0.42 l=0.15
X460 a_15715_627# a_14545_627# a_15608_993# VSS.t605 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0486 ps=0.63 w=0.36 l=0.15
X461 a_9122_n62# a_8205_n88# a_8677_122# VSS.t109 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0675 ps=0.735 w=0.36 l=0.15
X462 a_6124_993# a_4811_627# a_6040_993# VDD.t331 sky130_fd_pr__pfet_01v8_hvt ad=0.0787 pd=0.795 as=0.0567 ps=0.69 w=0.42 l=0.15
X463 VSS.t649 x3.X a_939_2457# VSS.t648 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X464 VDD.t113 VDD.t111 a_3333_601# VDD.t112 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.17 ps=1.81 w=0.64 l=0.15
X465 a_10711_n62# a_10596_212# a_10288_106# VSS.t228 sky130_fd_pr__nfet_01v8 ad=0.116 pd=1.09 as=0.0486 ps=0.63 w=0.36 l=0.15
X466 a_7350_n88# a_7896_106# a_7854_220# VDD.t689 sky130_fd_pr__pfet_01v8_hvt ad=0.132 pd=1.22 as=0.0882 ps=1.05 w=0.84 l=0.15
X467 a_1946_n62# a_1029_n88# a_1501_122# VSS.t434 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0675 ps=0.735 w=0.36 l=0.15
X468 a_15907_627# x2.X.t55 VSS.t274 VSS.t273 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.03 as=0.0703 ps=0.755 w=0.42 l=0.15
X469 VDD.t41 a_4860_1467# x10.X VDD.t40 sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X470 a_5002_1642# check[4].t2 VDD.t703 VDD.t702 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X471 a_5002_1315# check[4].t3 VSS.t668 VSS.t667 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X472 a_5223_1315# VSS.t525 a_4860_1467# VSS.t526 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X473 a_9147_1642# VSS.t725 a_8933_1642# VDD.t559 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.193 ps=1.34 w=0.42 l=0.15
X474 VDD_SW[7].t1 a_2136_627# VSS.t406 VSS.t405 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X475 VSS.t239 VDD.t766 a_15721_n62# VSS.t238 sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0974 ps=0.97 w=0.42 l=0.15
X476 a_10161_n62# a_10288_106# a_9742_n88# VSS.t261 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.03 as=0.0864 ps=0.91 w=0.64 l=0.15
X477 VDD_SW_b[3].t0 a_10983_895# VDD.t470 VDD.t469 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X478 a_12638_220# a_12447_n62# VDD.t346 VDD.t345 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X479 VSS.t94 a_12038_90# VSS_SW[2].t1 VSS.t93 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X480 VDD.t488 a_305_2457# x3.X VDD.t487 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X481 a_473_993# a_27_627# a_381_627# VDD.t549 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0651 ps=0.73 w=0.42 l=0.15
X482 a_3807_895# a_3648_993# a_3947_627# VSS.t231 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.109 ps=1.03 w=0.64 l=0.15
X483 a_14933_627# a_14379_627# a_14825_993# VSS.t595 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0675 ps=0.735 w=0.36 l=0.15
X484 VDD.t680 x3.X a_939_2457# VDD.t679 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X485 a_6760_1315# x9.A1.t51 a_6539_1642# VSS.t572 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X486 VSS.t129 a_6199_895# a_6920_627# VSS.t128 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X487 a_15329_304# a_14526_n88# VDD.t45 VDD.t44 sky130_fd_pr__pfet_01v8_hvt ad=0.0787 pd=0.795 as=0.0956 ps=0.875 w=0.42 l=0.15
X488 a_11015_220# a_10055_n62# VDD.t51 VDD.t50 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X489 VDD_SW[1].t1 a_16488_627# VSS.t11 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X490 a_15721_n62# a_15853_122# a_15585_n88# VSS.t568 sky130_fd_pr__nfet_01v8 ad=0.0974 pd=0.97 as=0.0864 ps=0.91 w=0.64 l=0.15
X491 a_5257_993# a_4977_627# a_5165_627# VSS.t293 sky130_fd_pr__nfet_01v8 ad=0.0675 pd=0.735 as=0.066 ps=0.745 w=0.36 l=0.15
X492 VDD.t572 D[5].t1 a_6730_n62# VDD.t571 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X493 x9.A1.t6 a_5323_2457# VDD.t528 VDD.t527 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X494 x20.X a_16109_1642# VSS.t172 VSS.t171 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.113 ps=1.04 w=0.65 l=0.15
X495 VSS.t316 VDD.t767 a_12553_n62# VSS.t315 sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.109 ps=1.03 w=0.42 l=0.15
X496 a_14909_993# a_14545_627# a_14825_993# VDD.t637 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X497 a_535_1642# x9.A1.t52 a_76_1467# VDD.t178 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X498 VDD.t587 a_5431_601# a_5341_993# VDD.t586 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X499 a_964_n62# a_174_n88# VSS.t243 VSS.t242 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0703 ps=0.755 w=0.42 l=0.15
X500 VSS.t408 a_505_1289# a_439_1315# VSS.t407 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X501 VSS.t227 a_10596_212# a_10597_n88# VSS.t226 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X502 a_12680_106# a_12989_n88# a_12924_n62# VSS.t352 sky130_fd_pr__nfet_01v8 ad=0.0486 pd=0.63 as=0.066 ps=0.745 w=0.36 l=0.15
X503 a_4338_n62# a_3420_212# a_3893_122# VDD.t85 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.0567 ps=0.69 w=0.42 l=0.15
X504 VDD.t428 a_939_2457# x2.X.t9 VDD.t427 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X505 a_10055_n62# x2.X.t56 VSS.t276 VSS.t275 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X506 VDD.t63 a_4958_n88# VSS_SW_b[5].t0 VDD.t62 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X507 VDD.t110 VDD.t108 a_9742_n88# VDD.t109 sky130_fd_pr__pfet_01v8_hvt ad=0.0956 pd=0.875 as=0.132 ps=1.22 w=0.42 l=0.15
X508 a_8409_n88# a_8677_122# a_8623_220# VDD.t668 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X509 VDD.t750 a_6017_n88# a_5950_304# VDD.t749 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X510 VSS.t418 a_1233_n88# a_1143_n62# VSS.t417 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.116 ps=1.09 w=0.64 l=0.15
X511 a_3551_627# a_3039_601# VSS.t574 VSS.t573 sky130_fd_pr__nfet_01v8 ad=0.116 pd=1.09 as=0.166 ps=1.8 w=0.64 l=0.15
X512 a_14733_627# D[1].t1 VDD.t59 VDD.t58 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X513 x9.A1.t5 a_5323_2457# VDD.t526 VDD.t525 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X514 VSS.t626 x30.A a_5323_2457# VSS.t625 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X515 a_3356_n62# a_2566_n88# VSS.t152 VSS.t151 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0703 ps=0.755 w=0.42 l=0.15
X516 VSS.t43 a_14526_n88# VSS_SW_b[1].t1 VSS.t42 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X517 VDD.t460 a_13375_895# a_13300_993# VDD.t459 sky130_fd_pr__pfet_01v8_hvt ad=0.0956 pd=0.875 as=0.0787 ps=0.795 w=0.42 l=0.15
X518 a_13323_627# a_12153_627# a_13216_993# VSS.t82 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0486 ps=0.63 w=0.36 l=0.15
X519 VDD.t33 check[6].t4 a_1503_1642# VDD.t32 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.118 ps=1.4 w=0.42 l=0.15
X520 a_12399_1315# VSS.t523 a_12036_1467# VSS.t524 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X521 VSS.t25 check[6].t5 a_1503_1642# VSS.t24 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.109 ps=1.36 w=0.42 l=0.15
X522 a_8204_212# x13.X VSS.t197 VSS.t196 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X523 VSS.t318 VDD.t768 a_15293_601# VSS.t317 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X524 VDD.t426 a_939_2457# x2.X.t8 VDD.t425 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X525 a_13515_627# x2.X.t57 VSS.t278 VSS.t277 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.03 as=0.0703 ps=0.755 w=0.42 l=0.15
X526 a_13936_1315# x9.A1.t53 a_13715_1642# VSS.t123 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X527 VDD.t107 VDD.t105 a_15293_601# VDD.t106 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.17 ps=1.81 w=0.64 l=0.15
X528 a_9949_627# D[3].t3 VSS.t351 VSS.t350 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X529 VSS.t79 VDD.t769 a_13329_n62# VSS.t78 sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0974 ps=0.97 w=0.42 l=0.15
X530 a_7681_1289# check[3].t4 VDD.t670 VDD.t669 sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X531 VSS.t217 a_1415_895# a_1363_627# VSS.t216 sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.066 ps=0.745 w=0.42 l=0.15
X532 a_10246_220# a_10055_n62# VDD.t49 VDD.t48 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X533 a_3893_122# a_3420_212# a_4137_n62# VSS.t89 sky130_fd_pr__nfet_01v8 ad=0.0675 pd=0.735 as=0.0671 ps=0.75 w=0.36 l=0.15
X534 a_13515_627# a_12901_601# a_13375_895# VSS.t144 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X535 a_7681_1289# check[3].t5 VSS.t639 VSS.t638 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X536 a_6285_122# a_5813_n88# a_6529_304# VDD.t451 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X537 a_15767_895# a_15608_993# a_15907_627# VSS.t616 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.109 ps=1.03 w=0.64 l=0.15
X538 x30.A a_4689_2457# VSS.t100 VSS.t99 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X539 VSS.t490 a_5323_2457# x9.A1.t23 VSS.t489 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X540 a_5761_304# a_4958_n88# VDD.t61 VDD.t60 sky130_fd_pr__pfet_01v8_hvt ad=0.0787 pd=0.795 as=0.0956 ps=0.875 w=0.42 l=0.15
X541 VDD_SW[2].t1 a_14096_627# VSS.t678 VSS.t677 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X542 a_12541_627# a_11987_627# a_12433_993# VSS.t551 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0675 ps=0.735 w=0.36 l=0.15
X543 VSS.t288 a_3807_895# a_4528_627# VSS.t287 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X544 VDD.t200 a_12901_601# a_12851_909# VDD.t199 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X545 VDD.t342 x3.A a_305_2457# VDD.t341 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X546 a_76_1467# VSS.t726 a_218_1642# VDD.t558 sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X547 a_13329_n62# a_13461_122# a_13193_n88# VSS.t709 sky130_fd_pr__nfet_01v8 ad=0.0974 pd=0.97 as=0.0864 ps=0.91 w=0.64 l=0.15
X548 a_15585_n88# a_14839_n62# a_15721_n62# VSS.t2 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X549 a_4137_n62# a_3625_n88# VSS.t341 VSS.t340 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0882 ps=0.84 w=0.42 l=0.15
X550 a_3420_212# x9.X VDD.t322 VDD.t321 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X551 VDD.t309 a_174_n88# VSS_SW_b[7].t0 VDD.t308 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X552 a_12517_993# a_12153_627# a_12433_993# VDD.t80 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X553 a_6539_1642# x9.A1.t54 a_6467_1642# VDD.t179 sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X554 a_8591_895# x2.X.t58 VDD.t25 VDD.t24 sky130_fd_pr__pfet_01v8_hvt ad=0.132 pd=1.22 as=0.0956 ps=0.875 w=0.42 l=0.15
X555 a_6539_1315# a_6285_1642# VSS.t339 VSS.t338 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.145 ps=1.11 w=0.42 l=0.15
X556 VDD.t222 a_5812_212# a_5813_n88# VDD.t221 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X557 a_14825_993# a_14379_627# a_14733_627# VDD.t628 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0651 ps=0.73 w=0.42 l=0.15
X558 x9.A1.t4 a_5323_2457# VDD.t524 VDD.t523 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X559 a_13705_304# a_13193_n88# VDD.t204 VDD.t203 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X560 VDD_SW_b[4].t0 a_8591_895# VDD.t234 VDD.t233 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X561 x9.X a_4149_1642# VSS.t368 VSS.t367 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.113 ps=1.04 w=0.65 l=0.15
X562 a_10288_106# a_10597_n88# a_10532_n62# VSS.t74 sky130_fd_pr__nfet_01v8 ad=0.0486 pd=0.63 as=0.066 ps=0.745 w=0.36 l=0.15
X563 a_6017_n88# a_6285_122# a_6231_220# VDD.t458 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X564 a_8623_220# a_7663_n62# VDD.t404 VDD.t403 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X565 VSS.t308 a_12607_601# a_12541_627# VSS.t307 sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0671 ps=0.75 w=0.42 l=0.15
X566 a_12341_627# D[2].t3 VDD.t67 VDD.t66 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X567 VDD.t424 a_939_2457# x2.X.t7 VDD.t423 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X568 a_11253_1642# a_11071_1642# VDD.t599 VDD.t598 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X569 a_16109_1642# x9.A1.t55 a_16037_1642# VDD.t281 sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X570 a_473_993# a_193_627# a_381_627# VSS.t688 sky130_fd_pr__nfet_01v8 ad=0.0675 pd=0.735 as=0.066 ps=0.745 w=0.36 l=0.15
X571 VDD_SW_b[7].t1 a_1415_895# VSS.t215 VSS.t214 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X572 a_9646_90# a_9742_n88# VDD.t476 VDD.t475 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X573 VDD_SW[3].t0 a_11704_627# VDD.t644 VDD.t643 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X574 VSS.t682 a_12134_n88# VSS_SW_b[2].t1 VSS.t681 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X575 a_10073_1289# check[2].t4 VDD.t442 VDD.t441 sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X576 a_16109_1315# a_15855_1642# VSS.t260 VSS.t259 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.145 ps=1.11 w=0.42 l=0.15
X577 x9.A1.t3 a_5323_2457# VDD.t522 VDD.t521 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X578 VSS.t624 x30.A a_5323_2457# VSS.t623 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X579 a_10073_1289# check[2].t5 VSS.t402 VSS.t401 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X580 x15.X a_11325_1642# VDD.t320 VDD.t319 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.158 ps=1.39 w=1 l=0.15
X581 VDD.t613 a_647_601# a_557_993# VDD.t612 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X582 a_1672_909# a_1256_993# a_1415_895# VDD.t705 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.132 ps=1.22 w=0.84 l=0.15
X583 a_4977_627# a_4811_627# VDD.t330 VDD.t329 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X584 a_5812_212# x11.X VSS.t508 VSS.t507 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X585 VSS.t564 a_8204_212# a_8205_n88# VSS.t563 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X586 a_8319_n62# a_8204_212# a_7896_106# VSS.t562 sky130_fd_pr__nfet_01v8 ad=0.116 pd=1.09 as=0.0486 ps=0.63 w=0.36 l=0.15
X587 a_11123_627# x2.X.t59 VSS.t21 VSS.t20 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.03 as=0.0703 ps=0.755 w=0.42 l=0.15
X588 VDD.t422 a_939_2457# x2.X.t6 VDD.t421 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X589 x2.X.t21 a_939_2457# VSS.t380 VSS.t379 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X590 VDD.t609 a_3039_601# a_2949_993# VDD.t608 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X591 VDD.t53 a_4862_90# VSS_SW[5].t0 VDD.t52 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X592 a_7557_627# D[4].t3 VSS.t327 VSS.t326 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X593 x9.A1.t2 a_5323_2457# VDD.t520 VDD.t519 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X594 a_12751_627# a_12901_601# a_12607_601# VSS.t143 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X595 a_939_2457# x3.X VSS.t647 VSS.t646 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X596 VSS.t488 a_5323_2457# x9.A1.t22 VSS.t487 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X597 a_10734_304# a_10597_n88# a_10288_106# VDD.t72 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X598 a_11123_627# a_10509_601# a_10983_895# VSS.t220 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X599 VSS.t321 D[5].t2 a_6730_n62# VSS.t320 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X600 a_3893_122# a_3421_n88# a_4137_304# VDD.t253 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X601 a_13375_895# a_13216_993# a_13515_627# VSS.t262 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.109 ps=1.03 w=0.64 l=0.15
X602 a_1159_627# a_647_601# VSS.t578 VSS.t577 sky130_fd_pr__nfet_01v8 ad=0.116 pd=1.09 as=0.166 ps=1.8 w=0.64 l=0.15
X603 VDD.t352 a_3807_895# a_3732_993# VDD.t351 sky130_fd_pr__pfet_01v8_hvt ad=0.0956 pd=0.875 as=0.0787 ps=0.795 w=0.42 l=0.15
X604 VDD.t284 a_10509_601# a_10459_909# VDD.t283 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X605 a_10937_n62# a_11069_122# a_10801_n88# VSS.t188 sky130_fd_pr__nfet_01v8 ad=0.0974 pd=0.97 as=0.0864 ps=0.91 w=0.64 l=0.15
X606 a_3755_627# a_2585_627# a_3648_993# VSS.t137 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0486 ps=0.63 w=0.36 l=0.15
X607 a_12851_909# a_12433_993# a_12607_601# VDD.t317 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X608 a_13193_n88# a_12447_n62# a_13329_n62# VSS.t286 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X609 a_4977_627# a_4811_627# VSS.t268 VSS.t267 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X610 a_6199_895# x2.X.t60 VDD.t27 VDD.t26 sky130_fd_pr__pfet_01v8_hvt ad=0.132 pd=1.22 as=0.0956 ps=0.875 w=0.42 l=0.15
X611 a_10125_993# a_9761_627# a_10041_993# VDD.t481 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X612 a_1028_212# x7.X VDD.t344 VDD.t343 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X613 VDD.t84 a_3420_212# a_3421_n88# VDD.t83 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X614 VSS.t486 a_5323_2457# x9.A1.t21 VSS.t485 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X615 a_9646_90# a_9742_n88# VSS.t437 VSS.t436 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X616 VSS.t248 a_15767_895# a_16488_627# VSS.t247 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X617 VDD.t165 D[1].t2 a_16298_n62# VDD.t164 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X618 a_3947_627# x2.X.t61 VSS.t559 VSS.t558 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.03 as=0.0703 ps=0.755 w=0.42 l=0.15
X619 a_15380_212# x20.X VDD.t642 VDD.t641 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X620 a_11313_304# a_10801_n88# VDD.t20 VDD.t19 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X621 x2.X.t20 a_939_2457# VSS.t378 VSS.t377 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X622 a_12036_1467# x9.A1.t56 a_12178_1315# VSS.t218 sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X623 a_2879_n62# x2.X.t62 VDD.t593 VDD.t592 sky130_fd_pr__pfet_01v8_hvt ad=0.17 pd=1.81 as=0.154 ps=1.34 w=0.64 l=0.15
X624 a_977_304# a_174_n88# VDD.t307 VDD.t306 sky130_fd_pr__pfet_01v8_hvt ad=0.0787 pd=0.795 as=0.0956 ps=0.875 w=0.42 l=0.15
X625 x7.X a_1757_1642# VDD.t693 VDD.t692 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.158 ps=1.39 w=1 l=0.15
X626 VDD.t163 check[1].t4 a_13929_1642# VDD.t162 sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.0767 ps=0.785 w=0.42 l=0.15
X627 VSS.t302 a_10215_601# a_10149_627# VSS.t301 sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0671 ps=0.75 w=0.42 l=0.15
X628 VSS.t81 VDD.t770 a_10937_n62# VSS.t80 sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0974 ps=0.97 w=0.42 l=0.15
X629 VDD.t486 a_305_2457# x3.X VDD.t485 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X630 VSS.t106 check[1].t5 a_13936_1315# VSS.t105 sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.0693 ps=0.75 w=0.42 l=0.15
X631 a_7254_90# a_7350_n88# VDD.t630 VDD.t629 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X632 a_12924_n62# a_12134_n88# VSS.t680 VSS.t679 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0703 ps=0.755 w=0.42 l=0.15
X633 VDD_SW_b[2].t1 a_13375_895# VSS.t423 VSS.t422 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X634 VDD.t697 a_8117_601# a_8848_909# VDD.t696 sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X635 VDD.t104 VDD.t102 a_3625_n88# VDD.t103 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X636 VDD.t420 a_939_2457# x2.X.t5 VDD.t419 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X637 a_3369_304# a_2566_n88# VDD.t212 VDD.t211 sky130_fd_pr__pfet_01v8_hvt ad=0.0787 pd=0.795 as=0.0956 ps=0.875 w=0.42 l=0.15
X638 a_10149_627# a_9595_627# a_10041_993# VSS.t202 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0675 ps=0.735 w=0.36 l=0.15
X639 a_10103_1642# x9.A1.t57 a_9644_1467# VDD.t282 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X640 a_2585_627# a_2419_627# VDD.t182 VDD.t181 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X641 VSS.t213 a_1415_895# a_2136_627# VSS.t212 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X642 VSS.t622 x30.A a_5323_2457# VSS.t621 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X643 VSS.t67 a_10073_1289# a_10007_1315# VSS.t66 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X644 VDD.t739 x10.X a_4811_627# VDD.t738 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X645 a_2949_993# a_2585_627# a_2865_993# VDD.t192 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X646 a_14825_993# a_14545_627# a_14733_627# VSS.t604 sky130_fd_pr__nfet_01v8 ad=0.0675 pd=0.735 as=0.066 ps=0.745 w=0.36 l=0.15
X647 a_505_1289# check[6].t6 VDD.t376 VDD.t375 sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X648 a_505_1289# check[6].t7 VSS.t314 VSS.t313 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X649 a_13632_909# a_13216_993# a_13375_895# VDD.t328 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.132 ps=1.22 w=0.84 l=0.15
X650 x9.A1.t1 a_5323_2457# VDD.t518 VDD.t517 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X651 x3.X a_305_2457# VSS.t445 VSS.t444 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X652 VDD.t360 a_2470_90# VSS_SW[6].t0 VDD.t359 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X653 a_5165_627# D[5].t3 VSS.t323 VSS.t322 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X654 VDD.t746 a_14999_601# a_14909_993# VDD.t745 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X655 a_14526_n88# a_15072_106# a_15030_220# VDD.t648 sky130_fd_pr__pfet_01v8_hvt ad=0.132 pd=1.22 as=0.0882 ps=1.05 w=0.84 l=0.15
X656 x3.A a_29_2457# VDD.t13 VDD.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X657 VDD.t418 a_939_2457# x2.X.t4 VDD.t417 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X658 a_939_2457# x3.X VSS.t645 VSS.t644 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X659 a_13906_n62# a_12988_212# a_13461_122# VDD.t251 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.0567 ps=0.69 w=0.42 l=0.15
X660 VDD.t262 x27.A a_4689_2457# VDD.t261 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X661 VSS.t484 a_5323_2457# x9.A1.t20 VSS.t483 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X662 a_10288_106# a_10596_212# a_10545_304# VDD.t294 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0787 ps=0.795 w=0.42 l=0.15
X663 VSS.t431 a_10983_895# a_10931_627# VSS.t430 sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.066 ps=0.745 w=0.42 l=0.15
X664 a_13461_122# a_12988_212# a_13705_n62# VSS.t189 sky130_fd_pr__nfet_01v8 ad=0.0675 pd=0.735 as=0.0671 ps=0.75 w=0.36 l=0.15
X665 VSS.t482 a_5323_2457# x9.A1.t19 VSS.t481 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X666 VDD.t276 a_1415_895# a_1340_993# VDD.t275 sky130_fd_pr__pfet_01v8_hvt ad=0.0956 pd=0.875 as=0.0787 ps=0.795 w=0.42 l=0.15
X667 a_1363_627# a_193_627# a_1256_993# VSS.t687 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0486 ps=0.63 w=0.36 l=0.15
X668 a_2585_627# a_2419_627# VSS.t126 VSS.t125 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X669 a_12751_627# x2.X.t63 VSS.t561 VSS.t560 sky130_fd_pr__nfet_01v8 ad=0.0974 pd=0.97 as=0.0882 ps=0.84 w=0.42 l=0.15
X670 a_3648_993# a_2419_627# a_3551_627# VSS.t124 sky130_fd_pr__nfet_01v8 ad=0.0486 pd=0.63 as=0.116 ps=1.09 w=0.36 l=0.15
X671 a_13705_n62# a_13193_n88# VSS.t146 VSS.t145 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0882 ps=0.84 w=0.42 l=0.15
X672 VDD.t416 a_939_2457# x2.X.t3 VDD.t415 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X673 VSS.t700 x10.X a_4811_627# VSS.t699 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X674 a_7254_90# a_7350_n88# VSS.t597 VSS.t596 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X675 VSS.t480 a_5323_2457# x9.A1.t18 VSS.t479 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X676 a_1555_627# x2.X.t64 VSS.t209 VSS.t208 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.03 as=0.0703 ps=0.755 w=0.42 l=0.15
X677 a_12988_212# x17.X VDD.t366 VDD.t365 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X678 a_8342_304# a_8205_n88# a_7896_106# VDD.t166 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X679 a_8432_993# a_7369_627# a_8288_909# VDD.t225 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X680 VDD.t240 a_15380_212# a_15381_n88# VDD.t239 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X681 x11.X a_6539_1642# VSS.t280 VSS.t279 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.113 ps=1.04 w=0.65 l=0.15
X682 a_8933_1642# VSS.t521 a_8933_1315# VSS.t522 sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X683 a_439_1315# VSS.t519 a_76_1467# VSS.t520 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X684 VDD.t695 a_8117_601# a_8067_909# VDD.t694 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X685 VDD.t399 check[3].t6 a_9147_1642# VDD.t398 sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.0767 ps=0.785 w=0.42 l=0.15
X686 VDD_SW[4].t0 a_9312_627# VDD.t9 VDD.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X687 VSS.t264 VDD.t771 a_1369_n62# VSS.t263 sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0974 ps=0.97 w=0.42 l=0.15
X688 a_10359_627# a_10509_601# a_10215_601# VSS.t219 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X689 x30.A a_4689_2457# VSS.t98 VSS.t97 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X690 VSS.t357 check[3].t7 a_9154_1315# VSS.t356 sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.0693 ps=0.75 w=0.42 l=0.15
X691 a_1555_627# a_941_601# a_1415_895# VSS.t665 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X692 a_12607_601# a_12433_993# a_12751_627# VSS.t253 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.0974 ps=0.97 w=0.64 l=0.15
X693 a_5323_2457# x30.A VDD.t655 VDD.t654 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X694 x2.X.t19 a_939_2457# VSS.t376 VSS.t375 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X695 a_13643_1642# a_13461_1642# VDD.t514 VDD.t513 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X696 a_14839_n62# x2.X.t65 VDD.t270 VDD.t269 sky130_fd_pr__pfet_01v8_hvt ad=0.17 pd=1.81 as=0.154 ps=1.34 w=0.64 l=0.15
X697 VSS.t53 a_7252_1467# x12.X VSS.t52 sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X698 VDD.t101 VDD.t99 a_15585_n88# VDD.t100 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X699 a_381_627# D[7].t2 VSS.t122 VSS.t121 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X700 a_1369_n62# a_1501_122# a_1233_n88# VSS.t358 sky130_fd_pr__nfet_01v8 ad=0.0974 pd=0.97 as=0.0864 ps=0.91 w=0.64 l=0.15
X701 a_12134_n88# a_12447_n62# a_12553_n62# VSS.t285 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X702 a_10007_1315# VSS.t517 a_9644_1467# VSS.t518 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X703 VDD.t161 x8.X a_2419_627# VDD.t160 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X704 a_10459_909# a_10041_993# a_10215_601# VDD.t318 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X705 a_3625_n88# a_2879_n62# a_3761_n62# VSS.t585 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X706 a_14428_1467# VSS.t727 a_14570_1642# VDD.t557 sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X707 a_12607_601# x2.X.t66 VDD.t272 VDD.t271 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X708 a_2865_993# a_2419_627# a_2773_627# VDD.t180 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0651 ps=0.73 w=0.42 l=0.15
X709 VDD.t732 a_1028_212# a_1029_n88# VDD.t731 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X710 VSS.t421 a_13375_895# a_14096_627# VSS.t420 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X711 a_14545_627# a_14379_627# VDD.t627 VDD.t626 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X712 a_11240_909# a_10824_993# a_10983_895# VDD.t23 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.132 ps=1.22 w=0.84 l=0.15
X713 VDD.t676 a_14428_1467# x18.X VDD.t675 sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X714 a_14570_1642# check[0].t6 VDD.t711 VDD.t710 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X715 a_1745_304# a_1233_n88# VDD.t457 VDD.t456 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X716 x9.A1.t0 a_5323_2457# VDD.t516 VDD.t515 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X717 a_14570_1315# check[0].t7 VSS.t676 VSS.t675 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X718 VDD.t187 a_6199_895# a_6920_627# VDD.t186 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X719 a_11514_n62# a_10596_212# a_11069_122# VDD.t293 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.0567 ps=0.69 w=0.42 l=0.15
X720 VSS.t41 a_4860_1467# x10.X VSS.t40 sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X721 VDD.t499 a_14430_90# VSS_SW[1].t0 VDD.t498 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X722 a_939_2457# x3.X VSS.t643 VSS.t642 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X723 a_13461_122# a_12989_n88# a_13705_304# VDD.t394 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X724 x3.A a_29_2457# VSS.t9 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X725 a_11325_1642# VSS.t515 a_11325_1315# VSS.t516 sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X726 a_10727_627# a_10215_601# VSS.t300 VSS.t299 sky130_fd_pr__nfet_01v8 ad=0.116 pd=1.09 as=0.166 ps=1.8 w=0.64 l=0.15
X727 a_10680_909# a_10215_601# VDD.t362 VDD.t361 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X728 VDD_SW_b[3].t1 a_10983_895# VSS.t429 VSS.t428 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X729 VDD.t414 a_939_2457# x2.X.t2 VDD.t413 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X730 VDD.t288 a_5725_601# a_6456_909# VDD.t287 sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X731 VSS.t108 D[1].t3 a_16298_n62# VSS.t107 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X732 a_11313_n62# a_10801_n88# VSS.t18 VSS.t17 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0882 ps=0.84 w=0.42 l=0.15
X733 VSS.t104 x8.X a_2419_627# VSS.t103 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X734 x2.X.t18 a_939_2457# VSS.t374 VSS.t373 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X735 a_15608_993# a_14379_627# a_15511_627# VSS.t594 sky130_fd_pr__nfet_01v8 ad=0.0486 pd=0.63 as=0.116 ps=1.09 w=0.36 l=0.15
X736 a_14545_627# a_14379_627# VSS.t593 VSS.t592 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X737 a_6040_993# a_4977_627# a_5896_909# VDD.t355 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X738 VSS.t478 a_5323_2457# x9.A1.t17 VSS.t477 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X739 a_4958_n88# a_5504_106# a_5462_220# VDD.t377 sky130_fd_pr__pfet_01v8_hvt ad=0.132 pd=1.22 as=0.0882 ps=1.05 w=0.84 l=0.15
X740 VDD_SW[5].t0 a_6920_627# VDD.t260 VDD.t259 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X741 a_10215_601# a_10041_993# a_10359_627# VSS.t254 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.0974 ps=0.97 w=0.64 l=0.15
X742 a_4860_1467# VSS.t728 a_5002_1642# VDD.t556 sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X743 a_1415_895# a_1256_993# a_1555_627# VSS.t670 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.109 ps=1.03 w=0.64 l=0.15
X744 a_11069_122# a_10596_212# a_11313_n62# VSS.t225 sky130_fd_pr__nfet_01v8 ad=0.0675 pd=0.735 as=0.0671 ps=0.75 w=0.36 l=0.15
X745 a_8861_1642# a_8679_1642# VDD.t368 VDD.t367 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X746 VDD.t171 check[2].t6 a_11071_1642# VDD.t170 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.118 ps=1.4 w=0.42 l=0.15
X747 a_5323_2457# x30.A VDD.t653 VDD.t652 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X748 x2.X.t17 a_939_2457# VSS.t372 VSS.t371 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X749 a_9742_n88# a_10055_n62# a_10161_n62# VSS.t48 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X750 VDD.t69 a_10073_1289# a_10103_1642# VDD.t68 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X751 VSS.t116 check[2].t7 a_11071_1642# VSS.t115 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.109 ps=1.36 w=0.42 l=0.15
X752 a_1233_n88# a_487_n62# a_1369_n62# VSS.t689 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X753 a_10359_627# x2.X.t67 VSS.t546 VSS.t545 sky130_fd_pr__nfet_01v8 ad=0.0974 pd=0.97 as=0.0882 ps=0.84 w=0.42 l=0.15
X754 x3.X a_305_2457# VDD.t484 VDD.t483 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X755 a_1256_993# a_27_627# a_1159_627# VSS.t509 sky130_fd_pr__nfet_01v8 ad=0.0486 pd=0.63 as=0.116 ps=1.09 w=0.36 l=0.15
X756 a_10215_601# x2.X.t68 VDD.t578 VDD.t577 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X757 VSS.t476 a_5323_2457# x9.A1.t16 VSS.t475 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X758 VDD.t358 a_78_90# VSS_SW[7].t0 VDD.t357 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X759 x27.A a_4413_2457# VDD.t39 VDD.t38 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X760 a_15767_895# x2.X.t69 VDD.t580 VDD.t579 sky130_fd_pr__pfet_01v8_hvt ad=0.132 pd=1.22 as=0.0956 ps=0.875 w=0.42 l=0.15
X761 a_12153_627# a_11987_627# VDD.t584 VDD.t583 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X762 a_7967_627# a_8117_601# a_7823_601# VSS.t663 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X763 VDD.t674 D[6].t3 a_4338_n62# VDD.t673 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X764 VDD.t568 x18.X a_14379_627# VDD.t567 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X765 VDD.t678 x3.X a_939_2457# VDD.t677 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X766 VSS.t266 VDD.t772 a_10161_n62# VSS.t265 sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.109 ps=1.03 w=0.42 l=0.15
X767 a_78_90# a_174_n88# VDD.t305 VDD.t304 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X768 a_2468_1467# VSS.t729 a_2610_1642# VDD.t555 sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X769 VDD.t250 a_12988_212# a_12989_n88# VDD.t249 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X770 VSS.t272 a_9646_90# VSS_SW[3].t1 VSS.t271 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X771 a_7896_106# a_8204_212# a_8153_304# VDD.t595 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0787 ps=0.795 w=0.42 l=0.15
X772 VDD.t350 a_3807_895# a_4528_627# VDD.t349 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X773 VDD.t210 a_2566_n88# VSS_SW_b[6].t0 VDD.t209 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X774 VDD.t387 a_3625_n88# a_3558_304# VDD.t386 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X775 VDD.t274 a_2468_1467# x8.X VDD.t273 sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X776 a_2610_1642# check[5].t4 VDD.t374 VDD.t373 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X777 a_8067_909# a_7649_993# a_7823_601# VDD.t704 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X778 x2.X.t1 a_939_2457# VDD.t412 VDD.t411 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X779 a_2610_1315# check[5].t5 VSS.t312 VSS.t311 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X780 VDD.t468 a_10983_895# a_10908_993# VDD.t467 sky130_fd_pr__pfet_01v8_hvt ad=0.0956 pd=0.875 as=0.0787 ps=0.795 w=0.42 l=0.15
X781 a_12447_n62# x2.X.t70 VDD.t721 VDD.t720 sky130_fd_pr__pfet_01v8_hvt ad=0.17 pd=1.81 as=0.154 ps=1.34 w=0.64 l=0.15
X782 VDD.t98 VDD.t96 a_13193_n88# VDD.t97 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X783 a_174_n88# a_720_106# a_678_220# VDD.t198 sky130_fd_pr__pfet_01v8_hvt ad=0.132 pd=1.22 as=0.0882 ps=1.05 w=0.84 l=0.15
X784 VSS.t35 VDD.t773 a_12901_601# VSS.t34 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X785 a_2865_993# a_2585_627# a_2773_627# VSS.t136 sky130_fd_pr__nfet_01v8 ad=0.0675 pd=0.735 as=0.066 ps=0.745 w=0.36 l=0.15
X786 a_12153_627# a_11987_627# VSS.t550 VSS.t549 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X787 a_7663_n62# x2.X.t71 VSS.t686 VSS.t685 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X788 a_9122_n62# a_8204_212# a_8677_122# VDD.t594 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.0567 ps=0.69 w=0.42 l=0.15
X789 a_15692_993# a_14379_627# a_15608_993# VDD.t625 sky130_fd_pr__pfet_01v8_hvt ad=0.0787 pd=0.795 as=0.0567 ps=0.69 w=0.42 l=0.15
X790 VSS.t542 x18.X a_14379_627# VSS.t541 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X791 VDD.t741 check[5].t6 a_4363_1642# VDD.t740 sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.0767 ps=0.785 w=0.42 l=0.15
X792 VDD.t95 VDD.t93 a_12901_601# VDD.t94 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.17 ps=1.81 w=0.64 l=0.15
X793 VDD.t208 a_12036_1467# x16.X VDD.t207 sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X794 a_12178_1642# check[1].t6 VDD.t636 VDD.t635 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X795 a_9644_1467# x9.A1.t58 a_9786_1315# VSS.t571 sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X796 VSS.t702 check[5].t7 a_4370_1315# VSS.t701 sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.0693 ps=0.75 w=0.42 l=0.15
X797 a_12178_1315# check[1].t7 VSS.t603 VSS.t602 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X798 a_2566_n88# a_3112_106# a_3070_220# VDD.t734 sky130_fd_pr__pfet_01v8_hvt ad=0.132 pd=1.22 as=0.0882 ps=1.05 w=0.84 l=0.15
X799 VDD_SW_b[4].t1 a_8591_895# VSS.t174 VSS.t173 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X800 VDD.t153 a_4689_2457# x30.A VDD.t152 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X801 VDD.t92 VDD.t90 a_7350_n88# VDD.t91 sky130_fd_pr__pfet_01v8_hvt ad=0.0956 pd=0.875 as=0.132 ps=1.22 w=0.42 l=0.15
X802 a_1946_n62# a_1028_212# a_1501_122# VDD.t730 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.0567 ps=0.69 w=0.42 l=0.15
X803 a_4363_1642# VSS.t730 a_4149_1642# VDD.t554 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.193 ps=1.34 w=0.42 l=0.15
X804 VDD.t151 a_12038_90# VSS_SW[2].t0 VDD.t150 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X805 a_1501_122# a_1028_212# a_1745_n62# VSS.t691 sky130_fd_pr__nfet_01v8 ad=0.0675 pd=0.735 as=0.0671 ps=0.75 w=0.36 l=0.15
X806 a_78_90# a_174_n88# VSS.t241 VSS.t240 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X807 VDD.t737 x6.X a_27_627# VDD.t736 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X808 VDD_SW[3].t1 a_11704_627# VSS.t613 VSS.t612 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X809 x2.X.t16 a_939_2457# VSS.t370 VSS.t369 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X810 a_7711_1642# x9.A1.t59 a_7252_1467# VDD.t603 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X811 a_1745_n62# a_1233_n88# VSS.t416 VSS.t415 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0882 ps=0.84 w=0.42 l=0.15
X812 VSS.t96 a_4689_2457# x30.A VSS.t95 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X813 x15.X a_11325_1642# VSS.t256 VSS.t255 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.113 ps=1.04 w=0.65 l=0.15
X814 VSS.t187 a_7681_1289# a_7615_1315# VSS.t186 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X815 a_13375_895# x2.X.t72 VDD.t723 VDD.t722 sky130_fd_pr__pfet_01v8_hvt ad=0.132 pd=1.22 as=0.0956 ps=0.875 w=0.42 l=0.15
X816 VDD.t177 D[7].t3 a_1946_n62# VDD.t176 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X817 VDD.t448 a_505_1289# a_535_1642# VDD.t447 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X818 x13.X a_8933_1642# VDD.t18 VDD.t17 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.158 ps=1.39 w=1 l=0.15
X819 a_13216_993# a_11987_627# a_13119_627# VSS.t548 sky130_fd_pr__nfet_01v8 ad=0.0486 pd=0.63 as=0.116 ps=1.09 w=0.36 l=0.15
X820 a_7823_601# a_7649_993# a_7967_627# VSS.t669 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.0974 ps=0.97 w=0.64 l=0.15
X821 x27.A a_4413_2457# VSS.t33 VSS.t32 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X822 a_1971_1642# VSS.t731 a_1757_1642# VDD.t553 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.193 ps=1.34 w=0.42 l=0.15
X823 VDD_SW_b[5].t0 a_6199_895# VDD.t185 VDD.t184 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X824 VSS.t619 a_7254_90# VSS_SW[4].t1 VSS.t618 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X825 a_12433_993# a_11987_627# a_12341_627# VDD.t582 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0651 ps=0.73 w=0.42 l=0.15
X826 a_7854_220# a_7663_n62# VDD.t402 VDD.t401 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X827 VDD.t57 check[4].t4 a_6285_1642# VDD.t56 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.118 ps=1.4 w=0.42 l=0.15
X828 a_3625_n88# a_3893_122# a_3839_220# VDD.t243 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X829 VSS.t55 check[4].t5 a_6285_1642# VSS.t54 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.109 ps=1.36 w=0.42 l=0.15
X830 VDD.t455 a_1233_n88# a_1166_304# VDD.t454 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X831 a_8288_909# a_7823_601# VDD.t195 VDD.t194 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X832 a_13715_1642# VSS.t513 a_13715_1315# VSS.t514 sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X833 VDD.t43 a_14526_n88# VSS_SW_b[1].t0 VDD.t42 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X834 VDD.t312 a_15767_895# a_16488_627# VDD.t311 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X835 a_10055_n62# x2.X.t73 VDD.t607 VDD.t606 sky130_fd_pr__pfet_01v8_hvt ad=0.17 pd=1.81 as=0.154 ps=1.34 w=0.64 l=0.15
X836 VSS.t698 x6.X a_27_627# VSS.t697 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X837 VSS.t16 a_10801_n88# a_10711_n62# VSS.t15 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.116 ps=1.09 w=0.64 l=0.15
X838 VDD.t665 a_15585_n88# a_15518_304# VDD.t664 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X839 VDD.t89 VDD.t87 a_10801_n88# VDD.t88 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X840 a_6231_220# a_5271_n62# VDD.t492 VDD.t491 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X841 a_5289_1289# check[4].t6 VDD.t391 VDD.t390 sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X842 x2.X.t0 a_939_2457# VDD.t410 VDD.t409 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X843 a_5289_1289# check[4].t7 VSS.t345 VSS.t344 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
R0 VSS VSS.n983 18062.3
R1 VSS.n4255 VSS.n4254 16202.7
R2 VSS.n3669 VSS.n3668 15745.9
R3 VSS.n3499 VSS.n3498 4543.55
R4 VSS.n1063 VSS.n1055 2992
R5 VSS.n3670 VSS.n3669 1854.77
R6 VSS.n990 VSS.n983 1757.32
R7 VSS VSS.n4255 1609.76
R8 VSS.n2561 VSS 1056
R9 VSS VSS.n4746 1056
R10 VSS VSS.n1347 1006.1
R11 VSS.n2421 VSS 1006.1
R12 VSS.n669 VSS 1006.1
R13 VSS VSS.n4817 1006.1
R14 VSS VSS.n4621 1006.1
R15 VSS.n4091 VSS 1006.1
R16 VSS VSS.n4657 1001.85
R17 VSS VSS.n3869 1001.85
R18 VSS VSS.n1477 817.779
R19 VSS VSS.n104 817.779
R20 VSS VSS.n321 817.779
R21 VSS.n4914 VSS 817.779
R22 VSS VSS.n3137 817.779
R23 VSS VSS.n4406 817.779
R24 VSS.t640 VSS.n1759 744.615
R25 VSS.t149 VSS.n2249 744.615
R26 VSS.n3668 VSS 692.958
R27 VSS.n4738 VSS.t279 649.846
R28 VSS.t541 VSS 643.903
R29 VSS VSS.t581 643.903
R30 VSS VSS.t409 643.903
R31 VSS.t223 VSS 643.903
R32 VSS.t699 VSS 643.903
R33 VSS VSS.t103 643.903
R34 VSS VSS.t697 643.903
R35 VSS.n1363 VSS.t604 603.659
R36 VSS.n2395 VSS.t83 603.659
R37 VSS.n654 VSS.t443 603.659
R38 VSS.n4788 VSS.t167 603.659
R39 VSS.n2872 VSS.t293 603.659
R40 VSS.n4065 VSS.t136 603.659
R41 VSS.n4269 VSS.t688 603.659
R42 VSS.n4670 VSS.t40 595.692
R43 VSS.n3776 VSS.t538 595.692
R44 VSS.t210 VSS.n3856 595.692
R45 VSS.n3722 VSS.t536 595.692
R46 VSS.t184 VSS.n3301 595.692
R47 VSS.n994 VSS.t10 590.245
R48 VSS.n1305 VSS.t56 590.245
R49 VSS.n1348 VSS.t541 590.245
R50 VSS.n1338 VSS.t677 590.245
R51 VSS.n2403 VSS.t64 590.245
R52 VSS.n2412 VSS.t581 590.245
R53 VSS.n2425 VSS.t612 590.245
R54 VSS.n774 VSS.t350 590.245
R55 VSS.t409 VSS.n668 590.245
R56 VSS.n671 VSS.t4 590.245
R57 VSS.n483 VSS.t326 590.245
R58 VSS.n4818 VSS.t223 590.245
R59 VSS.n471 VSS.t198 590.245
R60 VSS.n4591 VSS.t322 590.245
R61 VSS.n4622 VSS.t699 590.245
R62 VSS.n4603 VSS.t30 590.245
R63 VSS.n4073 VSS.t365 590.245
R64 VSS.n4082 VSS.t103 590.245
R65 VSS.n3984 VSS.t405 590.245
R66 VSS.n4131 VSS.t121 590.245
R67 VSS.t697 VSS.n4139 590.245
R68 VSS.n1083 VSS.t569 582.154
R69 VSS.n935 VSS.t105 568.615
R70 VSS.n2527 VSS.t518 568.615
R71 VSS.n2748 VSS.t540 568.615
R72 VSS.n999 VSS.t247 550
R73 VSS.n1333 VSS.t420 550
R74 VSS.n2431 VSS.t432 550
R75 VSS.n760 VSS.t175 550
R76 VSS.n467 VSS.t128 550
R77 VSS.n4565 VSS.t287 550
R78 VSS.n3980 VSS.t212 550
R79 VSS.n3784 VSS.t161 541.538
R80 VSS.n3734 VSS.t6 541.538
R81 VSS.n1348 VSS.t592 536.586
R82 VSS.n2412 VSS.t549 536.586
R83 VSS.n668 VSS.t204 536.586
R84 VSS.n4818 VSS.t672 536.586
R85 VSS.n4622 VSS.t267 536.586
R86 VSS.n4082 VSS.t125 536.586
R87 VSS.n4139 VSS.t510 536.586
R88 VSS.n3655 VSS.n3652 533.059
R89 VSS.n1138 VSS.t584 528
R90 VSS.n1745 VSS.t675 514.462
R91 VSS.n1822 VSS.t123 514.462
R92 VSS.n2272 VSS.t602 514.462
R93 VSS.n592 VSS.t401 514.462
R94 VSS.n594 VSS.t66 514.462
R95 VSS.n2729 VSS.t638 514.462
R96 VSS.n2731 VSS.t186 514.462
R97 VSS VSS.n4669 514.462
R98 VSS.n3857 VSS 514.462
R99 VSS.n3670 VSS 514.462
R100 VSS.n1249 VSS.t616 509.757
R101 VSS.n1922 VSS.t262 509.757
R102 VSS.n2461 VSS.t19 509.757
R103 VSS.n739 VSS.t12 509.757
R104 VSS.n446 VSS.t620 509.757
R105 VSS.n4012 VSS.t231 509.757
R106 VSS.n4110 VSS.t670 509.757
R107 VSS.n1103 VSS.t249 496.341
R108 VSS.n1312 VSS.t422 496.341
R109 VSS.n2439 VSS.t428 496.341
R110 VSS.n676 VSS.t173 496.341
R111 VSS.n431 VSS.t130 496.341
R112 VSS.n4571 VSS.t291 496.341
R113 VSS.n3950 VSS.t214 496.341
R114 VSS.n1068 VSS 487.385
R115 VSS.n3782 VSS.t117 487.385
R116 VSS.n3732 VSS.t24 487.385
R117 VSS.n1787 VSS 473.846
R118 VSS.n501 VSS.n500 473.24
R119 VSS.n3500 VSS.n3499 473.24
R120 VSS.n1709 VSS.t727 471.289
R121 VSS.n2294 VSS.t722 471.289
R122 VSS.n3683 VSS.t726 471.289
R123 VSS.n3898 VSS.t731 471.289
R124 VSS.n3836 VSS.t729 471.289
R125 VSS.n3763 VSS.t730 471.289
R126 VSS.n1145 VSS.t720 471.289
R127 VSS.n1845 VSS.t723 471.289
R128 VSS.n2179 VSS.t718 471.289
R129 VSS.n2533 VSS.t721 471.289
R130 VSS.n2615 VSS.t725 471.289
R131 VSS.n2738 VSS.t724 471.289
R132 VSS.n4719 VSS.t719 471.289
R133 VSS.n2791 VSS.t728 471.289
R134 VSS.n1731 VSS.t458 460.308
R135 VSS.n2286 VSS.t218 460.308
R136 VSS.n1115 VSS.t317 456.099
R137 VSS.n1873 VSS.t34 456.099
R138 VSS.n2445 VSS.t84 456.099
R139 VSS.n751 VSS.t659 456.099
R140 VSS.n458 VSS.t36 456.099
R141 VSS.n3991 VSS.t236 456.099
R142 VSS.n3958 VSS.t705 456.099
R143 VSS.n1367 VSS.t595 429.269
R144 VSS.n2391 VSS.t551 429.269
R145 VSS.n828 VSS.t202 429.269
R146 VSS.n4783 VSS.t674 429.269
R147 VSS.n2866 VSS.t270 429.269
R148 VSS.n4061 VSS.t127 429.269
R149 VSS.n4273 VSS.t512 429.269
R150 VSS.n3428 VSS 428.17
R151 VSS VSS.n3456 428.17
R152 VSS.n3629 VSS 428.17
R153 VSS.n3654 VSS 428.17
R154 VSS.n2229 VSS.t255 406.154
R155 VSS.t13 VSS.n2575 406.154
R156 VSS.n1245 VSS.t462 402.44
R157 VSS.n1878 VSS.t144 402.44
R158 VSS.n2453 VSS.t220 402.44
R159 VSS.n743 VSS.t664 402.44
R160 VSS.n450 VSS.t221 402.44
R161 VSS.n4008 VSS.t169 402.44
R162 VSS.n4104 VSS.t665 402.44
R163 VSS.n1179 VSS.t656 400
R164 VSS.n1533 VSS.t353 400
R165 VSS.n5054 VSS.t75 400
R166 VSS.n343 VSS.t109 400
R167 VSS.n2906 VSS.t412 400
R168 VSS.n3174 VSS.t194 400
R169 VSS.n4434 VSS.t434 400
R170 VSS.n1022 VSS.t608 391.111
R171 VSS.n1029 VSS.t107 391.111
R172 VSS.n1505 VSS.t460 391.111
R173 VSS.n1523 VSS.t303 391.111
R174 VSS.n1542 VSS.t157 391.111
R175 VSS.n94 VSS.t93 391.111
R176 VSS.t134 VSS.n110 391.111
R177 VSS.n126 VSS.t348 391.111
R178 VSS.n312 VSS.t271 391.111
R179 VSS.n322 VSS.t196 391.111
R180 VSS.n5002 VSS.t324 391.111
R181 VSS.n4918 VSS.t618 391.111
R182 VSS.t507 VSS.n4913 391.111
R183 VSS.n4885 VSS.t320 391.111
R184 VSS.n3096 VSS.t50 391.111
R185 VSS.t257 VSS.n3138 391.111
R186 VSS.n3146 VSS.t363 391.111
R187 VSS.n4393 VSS.t297 391.111
R188 VSS.t283 VSS.n4407 391.111
R189 VSS.n4424 VSS.t68 391.111
R190 VSS.n4245 VSS.t295 391.111
R191 VSS.n3498 VSS 388.733
R192 VSS.n2216 VSS.t361 379.077
R193 VSS.n2593 VSS.t356 379.077
R194 VSS.n1373 VSS.t712 375.611
R195 VSS.n2387 VSS.t307 375.611
R196 VSS.n822 VSS.t301 375.611
R197 VSS.n683 VSS.t140 375.611
R198 VSS.n2862 VSS.t554 375.611
R199 VSS.n4057 VSS.t575 375.611
R200 VSS.n4279 VSS.t579 375.611
R201 VSS.n4730 VSS.t229 365.538
R202 VSS.n4676 VSS.t667 365.538
R203 VSS.n3847 VSS.t311 365.538
R204 VSS.n3675 VSS.t703 365.538
R205 VSS.n1500 VSS.t46 364.445
R206 VSS.n80 VSS.t683 364.445
R207 VSS.n301 VSS.t436 364.445
R208 VSS.n4925 VSS.t596 364.445
R209 VSS.n3103 VSS.t62 364.445
R210 VSS.n4382 VSS.t155 364.445
R211 VSS.n4241 VSS.t240 364.445
R212 VSS.n1022 VSS.t180 355.557
R213 VSS.n1523 VSS.t190 355.557
R214 VSS.n110 VSS.t226 355.557
R215 VSS.n322 VSS.t563 355.557
R216 VSS.n4913 VSS.t165 355.557
R217 VSS.n3138 VSS.t91 355.557
R218 VSS.n4407 VSS.t693 355.557
R219 VSS.n1446 VSS.t617 337.779
R220 VSS.n12 VSS.t246 337.779
R221 VSS.n205 VSS.t261 337.779
R222 VSS.n4967 VSS.t654 337.779
R223 VSS.n3027 VSS.t319 337.779
R224 VSS.n3219 VSS.t695 337.779
R225 VSS.n4205 VSS.t142 337.779
R226 VSS.n1489 VSS.t42 328.889
R227 VSS.n69 VSS.t681 328.889
R228 VSS.n289 VSS.t440 328.889
R229 VSS.n4937 VSS.t600 328.889
R230 VSS.n3053 VSS.t60 328.889
R231 VSS.n3248 VSS.t153 328.889
R232 VSS.n4230 VSS.t244 328.889
R233 VSS VSS.t171 324.923
R234 VSS VSS.t206 324.923
R235 VSS.t255 VSS 324.923
R236 VSS.n2202 VSS.t591 324.923
R237 VSS VSS.t13 324.923
R238 VSS.n2607 VSS.t195 324.923
R239 VSS.t279 VSS 324.923
R240 VSS.n4726 VSS.t572 311.385
R241 VSS.n2813 VSS.t459 311.385
R242 VSS.n3843 VSS.t590 311.385
R243 VSS.n3679 VSS.t413 311.385
R244 VSS.n1478 VSS.t454 302.223
R245 VSS.n61 VSS.t0 302.223
R246 VSS.n284 VSS.t275 302.223
R247 VSS.n4873 VSS.t685 302.223
R248 VSS.n3060 VSS.t111 302.223
R249 VSS.n3242 VSS.t332 302.223
R250 VSS.n4149 VSS.t464 302.223
R251 VSS.n1298 VSS.t273 295.123
R252 VSS.n1398 VSS.t594 295.123
R253 VSS.n1930 VSS.t277 295.123
R254 VSS.n842 VSS.t548 295.123
R255 VSS.n2467 VSS.t20 295.123
R256 VSS.n2492 VSS.t203 295.123
R257 VSS.n733 VSS.t328 295.123
R258 VSS.n721 VSS.t671 295.123
R259 VSS.n440 VSS.t22 295.123
R260 VSS.n2835 VSS.t269 295.123
R261 VSS.n4016 VSS.t558 295.123
R262 VSS.n4030 VSS.t124 295.123
R263 VSS.n3922 VSS.t208 295.123
R264 VSS.n4125 VSS.t509 295.123
R265 VSS.n3737 VSS.n3733 294.007
R266 VSS.n3787 VSS.n3783 294.007
R267 VSS.n597 VSS.n593 294.007
R268 VSS.n2734 VSS.n2730 294.007
R269 VSS.n3707 VSS.n3706 292.5
R270 VSS.n3706 VSS.n3705 292.5
R271 VSS.n3704 VSS.n3703 292.5
R272 VSS.n3703 VSS.n3702 292.5
R273 VSS.n3701 VSS.n3700 292.5
R274 VSS.n3700 VSS.n3699 292.5
R275 VSS.n3279 VSS.n3278 292.5
R276 VSS.n3278 VSS.n3277 292.5
R277 VSS.n3282 VSS.n3281 292.5
R278 VSS.n3281 VSS.n3280 292.5
R279 VSS.n3285 VSS.n3284 292.5
R280 VSS.n3284 VSS.n3283 292.5
R281 VSS.n3288 VSS.n3287 292.5
R282 VSS.n3287 VSS.n3286 292.5
R283 VSS.n3274 VSS.n3273 292.5
R284 VSS.n3273 VSS.n3272 292.5
R285 VSS.n3733 VSS.n3732 292.5
R286 VSS.n3736 VSS.n3735 292.5
R287 VSS.n3735 VSS.n3734 292.5
R288 VSS.n3724 VSS.n3723 292.5
R289 VSS.n3723 VSS.n3722 292.5
R290 VSS.n3897 VSS.n3896 292.5
R291 VSS.n3896 VSS.n3895 292.5
R292 VSS.n3889 VSS.n3888 292.5
R293 VSS.n3888 VSS.n3887 292.5
R294 VSS.n3868 VSS.n3867 292.5
R295 VSS.n3869 VSS.n3868 292.5
R296 VSS.n3872 VSS.n3871 292.5
R297 VSS.n3871 VSS.n3870 292.5
R298 VSS.n3865 VSS.n3864 292.5
R299 VSS.n3864 VSS.n3863 292.5
R300 VSS.n3862 VSS.n3861 292.5
R301 VSS.n3861 VSS.n3860 292.5
R302 VSS.n3817 VSS.n3816 292.5
R303 VSS.n3816 VSS.n3815 292.5
R304 VSS.n3814 VSS.n3813 292.5
R305 VSS.n3813 VSS.n3812 292.5
R306 VSS.n3797 VSS.n3796 292.5
R307 VSS.n3796 VSS.n3795 292.5
R308 VSS.n3800 VSS.n3799 292.5
R309 VSS.n3799 VSS.n3798 292.5
R310 VSS.n3803 VSS.n3802 292.5
R311 VSS.n3802 VSS.n3801 292.5
R312 VSS.n3806 VSS.n3805 292.5
R313 VSS.n3805 VSS.n3804 292.5
R314 VSS.n3809 VSS.n3808 292.5
R315 VSS.n3808 VSS.n3807 292.5
R316 VSS.n3794 VSS.n3793 292.5
R317 VSS.n3793 VSS.n3792 292.5
R318 VSS.n3783 VSS.n3782 292.5
R319 VSS.n3786 VSS.n3785 292.5
R320 VSS.n3785 VSS.n3784 292.5
R321 VSS.n3778 VSS.n3777 292.5
R322 VSS.n3777 VSS.n3776 292.5
R323 VSS.n3753 VSS.n3752 292.5
R324 VSS.n3752 VSS.n3751 292.5
R325 VSS.n3760 VSS.n3759 292.5
R326 VSS.n3759 VSS.n3758 292.5
R327 VSS.n4656 VSS.n4655 292.5
R328 VSS.n4657 VSS.n4656 292.5
R329 VSS.n4660 VSS.n4659 292.5
R330 VSS.n4659 VSS.n4658 292.5
R331 VSS.n2821 VSS.n2820 292.5
R332 VSS.n2820 VSS.n2819 292.5
R333 VSS.n4666 VSS.n4665 292.5
R334 VSS.n4665 VSS.n4664 292.5
R335 VSS.n4701 VSS.n4700 292.5
R336 VSS.n4700 VSS.n4699 292.5
R337 VSS.n4743 VSS.n4742 292.5
R338 VSS.n4742 VSS.n4741 292.5
R339 VSS.n4745 VSS.n4744 292.5
R340 VSS.n4746 VSS.n4745 292.5
R341 VSS.n4749 VSS.n4748 292.5
R342 VSS.n4748 VSS.n4747 292.5
R343 VSS.n2776 VSS.n2775 292.5
R344 VSS.n2775 VSS.n2774 292.5
R345 VSS.n2769 VSS.n2768 292.5
R346 VSS.n2768 VSS.n2767 292.5
R347 VSS.n2743 VSS.n2742 292.5
R348 VSS.n2742 VSS.n2741 292.5
R349 VSS.n2750 VSS.n2749 292.5
R350 VSS.n2749 VSS.n2748 292.5
R351 VSS.n2733 VSS.n2732 292.5
R352 VSS.n2732 VSS.n2731 292.5
R353 VSS.n2730 VSS.n2729 292.5
R354 VSS.n2709 VSS.n2708 292.5
R355 VSS.n2708 VSS.n2707 292.5
R356 VSS.n2706 VSS.n2705 292.5
R357 VSS.n2705 VSS.n2704 292.5
R358 VSS.n2703 VSS.n2702 292.5
R359 VSS.n2702 VSS.n2701 292.5
R360 VSS.n2700 VSS.n2699 292.5
R361 VSS.n2699 VSS.n2698 292.5
R362 VSS.n2697 VSS.n2696 292.5
R363 VSS.n2696 VSS.n2695 292.5
R364 VSS.n2694 VSS.n2693 292.5
R365 VSS.n2693 VSS.n2692 292.5
R366 VSS.n2675 VSS.n2674 292.5
R367 VSS.n2674 VSS.n2673 292.5
R368 VSS.n2678 VSS.n2677 292.5
R369 VSS.n2677 VSS.n2676 292.5
R370 VSS.n2563 VSS.n2562 292.5
R371 VSS.n2562 VSS.n2561 292.5
R372 VSS.n2551 VSS.n2550 292.5
R373 VSS.n2550 VSS.n2549 292.5
R374 VSS.n2559 VSS.n2558 292.5
R375 VSS.n2560 VSS.n2559 292.5
R376 VSS.n2554 VSS.n2553 292.5
R377 VSS.n2553 VSS.n2552 292.5
R378 VSS.n2543 VSS.n2542 292.5
R379 VSS.n2542 VSS.n2541 292.5
R380 VSS.n2538 VSS.n2537 292.5
R381 VSS.n2537 VSS.n2536 292.5
R382 VSS.n2529 VSS.n2528 292.5
R383 VSS.n2528 VSS.n2527 292.5
R384 VSS.n593 VSS.n592 292.5
R385 VSS.n596 VSS.n595 292.5
R386 VSS.n595 VSS.n594 292.5
R387 VSS.n626 VSS.n625 292.5
R388 VSS.n625 VSS.n624 292.5
R389 VSS.n2113 VSS.n2112 292.5
R390 VSS.n2112 VSS.n2111 292.5
R391 VSS.n2110 VSS.n2109 292.5
R392 VSS.n2109 VSS.n2108 292.5
R393 VSS.n2107 VSS.n2106 292.5
R394 VSS.n2106 VSS.n2105 292.5
R395 VSS.n612 VSS.n611 292.5
R396 VSS.n611 VSS.n610 292.5
R397 VSS.n615 VSS.n614 292.5
R398 VSS.n614 VSS.n613 292.5
R399 VSS.n618 VSS.n617 292.5
R400 VSS.n617 VSS.n616 292.5
R401 VSS.n621 VSS.n620 292.5
R402 VSS.n620 VSS.n619 292.5
R403 VSS.n1639 VSS.n1638 292.5
R404 VSS.n1638 VSS.n1637 292.5
R405 VSS.n1636 VSS.n1635 292.5
R406 VSS.n1635 VSS.n1634 292.5
R407 VSS.n1633 VSS.n1632 292.5
R408 VSS.n1632 VSS.n1631 292.5
R409 VSS.n1630 VSS.n1629 292.5
R410 VSS.n1629 VSS.n1628 292.5
R411 VSS.n1627 VSS.n1626 292.5
R412 VSS.n1626 VSS.n1625 292.5
R413 VSS.n1653 VSS.n1652 292.5
R414 VSS.n1652 VSS.n1651 292.5
R415 VSS.n1770 VSS.n1769 292.5
R416 VSS.n1769 VSS.n1768 292.5
R417 VSS.n1767 VSS.n1766 292.5
R418 VSS.n1766 VSS.n1765 292.5
R419 VSS.n1989 VSS.n1988 292.5
R420 VSS.n1988 VSS.n1987 292.5
R421 VSS.n1986 VSS.n1985 292.5
R422 VSS.n1985 VSS.n1984 292.5
R423 VSS.n1983 VSS.n1982 292.5
R424 VSS.n1982 VSS.n1981 292.5
R425 VSS.n2343 VSS.n2342 292.5
R426 VSS.n2342 VSS.n2341 292.5
R427 VSS.n2346 VSS.n2345 292.5
R428 VSS.n2345 VSS.n2344 292.5
R429 VSS.n2349 VSS.n2348 292.5
R430 VSS.n2348 VSS.n2347 292.5
R431 VSS.n2257 VSS.n2256 292.5
R432 VSS.n2256 VSS.n2255 292.5
R433 VSS.n1185 VSS.t179 284.445
R434 VSS.n1896 VSS.t189 284.445
R435 VSS.n5049 VSS.t225 284.445
R436 VSS.n347 VSS.t565 284.445
R437 VSS.n2901 VSS.t163 284.445
R438 VSS.n4520 VSS.t89 284.445
R439 VSS.n4355 VSS.t691 284.445
R440 VSS VSS.n2228 284.308
R441 VSS.n2578 VSS 284.308
R442 VSS.t608 VSS 275.557
R443 VSS.t303 VSS 275.557
R444 VSS VSS.t134 275.557
R445 VSS.t196 VSS 275.557
R446 VSS VSS.t507 275.557
R447 VSS VSS.t257 275.557
R448 VSS VSS.t283 275.557
R449 VSS VSS.n4737 270.769
R450 VSS.n3654 VSS.t8 270.423
R451 VSS.n1451 VSS.t3 266.668
R452 VSS.n46 VSS.t285 266.668
R453 VSS.n147 VSS.t48 266.668
R454 VSS.n4851 VSS.t359 266.668
R455 VSS.n3043 VSS.t453 266.668
R456 VSS.n4471 VSS.t586 266.668
R457 VSS.n4140 VSS.t690 266.668
R458 VSS.n1264 VSS.t633 248.889
R459 VSS.n1902 VSS.t145 248.889
R460 VSS.n5040 VSS.t17 248.889
R461 VSS.n361 VSS.t232 248.889
R462 VSS.n2922 VSS.t714 248.889
R463 VSS.n4528 VSS.t340 248.889
R464 VSS.n4363 VSS.t415 248.889
R465 VSS.n517 VSS.t493 247.887
R466 VSS.n3411 VSS.t627 247.887
R467 VSS.n3463 VSS.t200 247.887
R468 VSS.n3446 VSS.t32 247.887
R469 VSS.n3446 VSS.t610 247.887
R470 VSS.n3333 VSS.t383 247.887
R471 VSS.n3617 VSS.t646 247.887
R472 VSS.n3646 VSS.t281 247.887
R473 VSS.n3659 VSS.t113 247.887
R474 VSS.n969 VSS.t119 243.692
R475 VSS.n4658 VSS 243.692
R476 VSS.n3870 VSS 243.692
R477 VSS.n913 VSS.t159 230.155
R478 VSS.n2541 VSS.t571 230.155
R479 VSS.n2767 VSS.t583 230.155
R480 VSS.n1406 VSS.t251 228.049
R481 VSS.n873 VSS.t424 228.049
R482 VSS.n2474 VSS.t430 228.049
R483 VSS.n729 VSS.t177 228.049
R484 VSS.n436 VSS.t132 228.049
R485 VSS.n4022 VSS.t289 228.049
R486 VSS.n3932 VSS.t216 228.049
R487 VSS.n517 VSS.t487 225.352
R488 VSS.n3411 VSS.t621 225.352
R489 VSS.n3463 VSS.t99 225.352
R490 VSS.n3333 VSS.t399 225.352
R491 VSS.n3617 VSS.t648 225.352
R492 VSS.n3646 VSS.t444 225.352
R493 VSS.n1064 VSS.n1063 216.615
R494 VSS.n1068 VSS.n1067 216.615
R495 VSS.n1083 VSS.n1082 216.615
R496 VSS.n1138 VSS.n1137 216.615
R497 VSS.n1154 VSS.n1153 216.615
R498 VSS.n1208 VSS.n1207 216.615
R499 VSS.n1228 VSS.n1227 216.615
R500 VSS.n969 VSS.n968 216.615
R501 VSS.n1646 VSS.n1645 216.615
R502 VSS.t206 VSS.n1784 216.615
R503 VSS.n2230 VSS.n2229 216.615
R504 VSS.n2082 VSS.n2081 216.615
R505 VSS.n2215 VSS.n2214 216.615
R506 VSS.n2201 VSS.n2200 216.615
R507 VSS.n2150 VSS.n2149 216.615
R508 VSS.n2133 VSS.n2132 216.615
R509 VSS.n2119 VSS.n2118 216.615
R510 VSS.n2575 VSS.n2574 216.615
R511 VSS.n2577 VSS.n2576 216.615
R512 VSS.n2592 VSS.n2591 216.615
R513 VSS.n2606 VSS.n2605 216.615
R514 VSS.n2646 VSS.n2645 216.615
R515 VSS.n2664 VSS.n2663 216.615
R516 VSS.n2684 VSS.n2683 216.615
R517 VSS.t171 VSS.n1065 203.077
R518 VSS.n1783 VSS.n1782 203.077
R519 VSS.n1787 VSS.n1786 203.077
R520 VSS.n935 VSS.n934 203.077
R521 VSS.n1822 VSS.n1821 203.077
R522 VSS.n1853 VSS.n1852 203.077
R523 VSS.n1836 VSS.n1835 203.077
R524 VSS.n898 VSS.n897 203.077
R525 VSS.n913 VSS.n912 203.077
R526 VSS.n1996 VSS.n1995 203.077
R527 VSS.n3751 VSS.t589 203.077
R528 VSS.n3887 VSS.t414 203.077
R529 VSS.n521 VSS.t477 202.817
R530 VSS.n3324 VSS.t385 202.817
R531 VSS.n1592 VSS.t182 195.556
R532 VSS.n1431 VSS.t26 195.556
R533 VSS.n2023 VSS.t192 195.556
R534 VSS.n18 VSS.t315 195.556
R535 VSS.n222 VSS.t228 195.556
R536 VSS.n199 VSS.t265 195.556
R537 VSS.n410 VSS.t562 195.556
R538 VSS.n4961 VSS.t86 195.556
R539 VSS.n2991 VSS.t164 195.556
R540 VSS.n3023 VSS.t28 195.556
R541 VSS.n3195 VSS.t90 195.556
R542 VSS.n3225 VSS.t72 195.556
R543 VSS.n4171 VSS.t692 195.556
R544 VSS.n4199 VSS.t70 195.556
R545 VSS.n3504 VSS.t388 190.065
R546 VSS.n505 VSS.t476 190.065
R547 VSS.n4715 VSS.t338 189.538
R548 VSS.n2800 VSS.t426 189.538
R549 VSS.n3832 VSS.t556 189.538
R550 VSS.n3690 VSS.t407 189.538
R551 VSS.n4295 VSS.t578 189.362
R552 VSS.n4038 VSS.t574 189.362
R553 VSS.n2843 VSS.t553 189.362
R554 VSS.n712 VSS.t139 189.362
R555 VSS.n2477 VSS.t300 189.362
R556 VSS.n856 VSS.t310 189.362
R557 VSS.n1389 VSS.t711 189.362
R558 VSS.n4163 VSS.t418 189.362
R559 VSS.n396 VSS.t235 189.362
R560 VSS.n245 VSS.t16 189.362
R561 VSS.n1579 VSS.t636 189.362
R562 VSS.n1402 VSS.t605 187.805
R563 VSS.n879 VSS.t82 187.805
R564 VSS.n2496 VSS.t442 187.805
R565 VSS.n725 VSS.t168 187.805
R566 VSS.n2831 VSS.t294 187.805
R567 VSS.n4026 VSS.t137 187.805
R568 VSS.n3927 VSS.t687 187.805
R569 VSS.n4503 VSS.t343 187.167
R570 VSS.n2975 VSS.t717 187.167
R571 VSS.n2020 VSS.t148 187.167
R572 VSS.n511 VSS.t491 180.282
R573 VSS.n3405 VSS.t629 180.282
R574 VSS.n3468 VSS.t95 180.282
R575 VSS.n3568 VSS.t381 180.282
R576 VSS.n3613 VSS.t642 180.282
R577 VSS.n3640 VSS.t450 180.282
R578 VSS.n1674 VSS.t606 176
R579 VSS.n2333 VSS.t336 176
R580 VSS.n2552 VSS.t403 176
R581 VSS.n2774 VSS.t543 176
R582 VSS.n2170 VSS.t566 162.463
R583 VSS.n2637 VSS.t305 162.463
R584 VSS.n506 VSS.t475 157.746
R585 VSS.n527 VSS.t497 157.746
R586 VSS.n3505 VSS.t387 157.746
R587 VSS.n3538 VSS.t369 157.746
R588 VSS.n1424 VSS.t44 151.112
R589 VSS.n7 VSS.t679 151.112
R590 VSS.n231 VSS.t438 151.112
R591 VSS.n400 VSS.t598 151.112
R592 VSS.n2996 VSS.t58 151.112
R593 VSS.n3214 VSS.t151 151.112
R594 VSS.n4176 VSS.t242 151.112
R595 VSS.n1660 VSS.n1659 148.923
R596 VSS.n1674 VSS.n1673 148.923
R597 VSS.n1688 VSS.n1687 148.923
R598 VSS.n1717 VSS.n1716 148.923
R599 VSS.n1731 VSS.n1730 148.923
R600 VSS.n1745 VSS.n1744 148.923
R601 VSS.n1759 VSS.n957 148.923
R602 VSS.n1762 VSS.n1761 148.923
R603 VSS.n2356 VSS.n2355 148.923
R604 VSS.n2333 VSS.n2332 148.923
R605 VSS.n2070 VSS.n2069 148.923
R606 VSS.n2302 VSS.n2301 148.923
R607 VSS.n2286 VSS.n2285 148.923
R608 VSS.n2272 VSS.n2271 148.923
R609 VSS.n2249 VSS.n2243 148.923
R610 VSS.n2252 VSS.n2251 148.923
R611 VSS.n4657 VSS.t701 148.923
R612 VSS.n3869 VSS.t614 148.923
R613 VSS.n1709 VSS.t527 148.35
R614 VSS.n2294 VSS.t523 148.35
R615 VSS.n3683 VSS.t519 148.35
R616 VSS.n3898 VSS.t535 148.35
R617 VSS.n3836 VSS.t533 148.35
R618 VSS.n3763 VSS.t537 148.35
R619 VSS.n1145 VSS.t529 148.35
R620 VSS.n1845 VSS.t513 148.35
R621 VSS.n2179 VSS.t515 148.35
R622 VSS.n2533 VSS.t517 148.35
R623 VSS.n2615 VSS.t521 148.35
R624 VSS.n2738 VSS.t539 148.35
R625 VSS.n4719 VSS.t531 148.35
R626 VSS.n2791 VSS.t525 148.35
R627 VSS.n4134 VSS.t122 145.006
R628 VSS.n4076 VSS.t366 145.006
R629 VSS.n777 VSS.t351 145.006
R630 VSS.n2406 VSS.t65 145.006
R631 VSS.n1308 VSS.t57 145.006
R632 VSS.n4427 VSS.t69 145.006
R633 VSS.n3149 VSS.t364 145.006
R634 VSS.n4888 VSS.t321 145.006
R635 VSS.n5005 VSS.t325 145.006
R636 VSS.n129 VSS.t349 145.006
R637 VSS.n1545 VSS.t158 145.006
R638 VSS.n1032 VSS.t108 145.006
R639 VSS.n4596 VSS.t323 143.871
R640 VSS.n482 VSS.t327 143.871
R641 VSS VSS.t640 135.386
R642 VSS.n1760 VSS 135.386
R643 VSS VSS.t149 135.386
R644 VSS.n2250 VSS 135.386
R645 VSS VSS.t587 135.386
R646 VSS.t52 VSS 135.386
R647 VSS.n4722 VSS.t532 135.386
R648 VSS.n2794 VSS.t526 135.386
R649 VSS.t40 VSS 135.386
R650 VSS.n3839 VSS.t534 135.386
R651 VSS VSS.t210 135.386
R652 VSS.n3686 VSS.t520 135.386
R653 VSS VSS.t184 135.386
R654 VSS.n3370 VSS.t481 135.212
R655 VSS.n3399 VSS.t623 135.212
R656 VSS.n3472 VSS.t97 135.212
R657 VSS.n3575 VSS.t395 135.212
R658 VSS.n3607 VSS.t650 135.212
R659 VSS.n3634 VSS.t446 135.212
R660 VSS.n1385 VSS.t463 134.147
R661 VSS.n862 VSS.t143 134.147
R662 VSS.n793 VSS.t219 134.147
R663 VSS.n708 VSS.t663 134.147
R664 VSS.n2848 VSS.t222 134.147
R665 VSS.n4043 VSS.t170 134.147
R666 VSS.n4291 VSS.t666 134.147
R667 VSS.n1587 VSS.t655 124.445
R668 VSS.n3 VSS.t352 124.445
R669 VSS.n227 VSS.t74 124.445
R670 VSS.n406 VSS.t110 124.445
R671 VSS.n3002 VSS.t411 124.445
R672 VSS.n3201 VSS.t193 124.445
R673 VSS.n4181 VSS.t435 124.445
R674 VSS.n3514 VSS.n3513 116.219
R675 VSS.n3524 VSS.n3523 116.219
R676 VSS.n3530 VSS.n3529 116.219
R677 VSS.n3537 VSS.n3536 116.219
R678 VSS.n3331 VSS.n3330 116.219
R679 VSS.n3574 VSS.n3573 116.219
R680 VSS.n3304 VSS.n3303 116.219
R681 VSS.n3315 VSS.n3314 116.219
R682 VSS.n3601 VSS.n3600 116.219
R683 VSS.n3612 VSS.n3611 116.219
R684 VSS.n552 VSS.n551 116.219
R685 VSS.n546 VSS.n545 116.219
R686 VSS.n536 VSS.n535 116.219
R687 VSS.n526 VSS.n525 116.219
R688 VSS.n516 VSS.n515 116.219
R689 VSS.n3369 VSS.n3368 116.219
R690 VSS.n3379 VSS.n3378 116.219
R691 VSS.n3385 VSS.n3384 116.219
R692 VSS.n3394 VSS.n3393 116.219
R693 VSS.n3404 VSS.n3403 116.219
R694 VSS.n3302 VSS.t647 114.775
R695 VSS.n3367 VSS.t628 114.775
R696 VSS.n4278 VSS.n4277 113.207
R697 VSS.n4056 VSS.n4055 113.207
R698 VSS.n2861 VSS.n2860 113.207
R699 VSS.n688 VSS.n687 113.207
R700 VSS.n817 VSS.n816 113.207
R701 VSS.n2386 VSS.n2385 113.207
R702 VSS.n1372 VSS.n1371 113.207
R703 VSS.n4362 VSS.n4361 113.207
R704 VSS.n4527 VSS.n4526 113.207
R705 VSS.n2927 VSS.n2926 113.207
R706 VSS.n366 VSS.n365 113.207
R707 VSS.n5034 VSS.n5033 113.207
R708 VSS.n1944 VSS.n1943 113.207
R709 VSS.n1270 VSS.n1269 113.207
R710 VSS.n559 VSS.t495 112.677
R711 VSS.n531 VSS.t479 112.677
R712 VSS.n3509 VSS.t377 112.677
R713 VSS.n3544 VSS.t389 112.677
R714 VSS.n3462 VSS.n3461 109.3
R715 VSS.n3645 VSS.n3644 109.3
R716 VSS.n4249 VSS.n4248 109.231
R717 VSS.n3988 VSS.n3987 109.231
R718 VSS.n4607 VSS.n4606 109.231
R719 VSS.n475 VSS.n474 109.231
R720 VSS.n675 VSS.n674 109.231
R721 VSS.n2429 VSS.n2428 109.231
R722 VSS.n1342 VSS.n1341 109.231
R723 VSS.n998 VSS.n997 109.231
R724 VSS.n4397 VSS.n4396 109.231
R725 VSS.n3100 VSS.n3099 109.231
R726 VSS.n4922 VSS.n4921 109.231
R727 VSS.n316 VSS.n315 109.231
R728 VSS.n1509 VSS.n1508 109.231
R729 VSS.n3921 VSS.n3920 109.043
R730 VSS.n4019 VSS.n4018 109.043
R731 VSS.n443 VSS.n442 109.043
R732 VSS.n736 VSS.n735 109.043
R733 VSS.n2470 VSS.n2469 109.043
R734 VSS.n1929 VSS.n1928 109.043
R735 VSS.n1303 VSS.n1302 109.043
R736 VSS.n3022 VSS.n3021 109.043
R737 VSS.n23 VSS.n22 109.043
R738 VSS.n3954 VSS.n3953 108.689
R739 VSS.n4575 VSS.n4574 108.689
R740 VSS.n435 VSS.n434 108.689
R741 VSS.n680 VSS.n679 108.689
R742 VSS.n2443 VSS.n2442 108.689
R743 VSS.n1316 VSS.n1315 108.689
R744 VSS.n1107 VSS.n1106 108.689
R745 VSS.n3252 VSS.n3251 108.689
R746 VSS.n293 VSS.n292 108.689
R747 VSS.n73 VSS.n72 108.591
R748 VSS.t346 VSS.n1700 108.308
R749 VSS.t470 VSS.n2315 108.308
R750 VSS.n2187 VSS.t516 108.308
R751 VSS.t516 VSS.n2186 108.308
R752 VSS.n2623 VSS.t522 108.308
R753 VSS.t522 VSS.n2622 108.308
R754 VSS.n3476 VSS.n3475 108.254
R755 VSS.n3638 VSS.n3637 108.254
R756 VSS.n93 VSS.n92 107.903
R757 VSS.n3662 VSS.n3658 107.478
R758 VSS.n4136 VSS.n4135 107.478
R759 VSS.n4086 VSS.n4085 107.478
R760 VSS.n4626 VSS.n4625 107.478
R761 VSS.n4822 VSS.n4821 107.478
R762 VSS.n664 VSS.n663 107.478
R763 VSS.n2416 VSS.n2415 107.478
R764 VSS.n1352 VSS.n1351 107.478
R765 VSS.n3298 VSS.n3297 107.478
R766 VSS.n3853 VSS.n3852 107.478
R767 VSS.n4674 VSS.n4673 107.478
R768 VSS.n2780 VSS.n2779 107.478
R769 VSS.n4412 VSS.n4411 107.478
R770 VSS.n3143 VSS.n3142 107.478
R771 VSS.n4880 VSS.n4879 107.478
R772 VSS.n283 VSS.n282 107.478
R773 VSS.n107 VSS.n106 107.478
R774 VSS.n1527 VSS.n1526 107.478
R775 VSS.n1026 VSS.n1025 107.478
R776 VSS.n3052 VSS.n3051 107.398
R777 VSS.n4936 VSS.n4935 107.398
R778 VSS.n1488 VSS.n1487 107.398
R779 VSS.n4229 VSS.n4228 107.398
R780 VSS.n3749 VSS.n3748 107.24
R781 VSS.n4653 VSS.n2822 107.24
R782 VSS.n2556 VSS.n2555 107.24
R783 VSS.n4751 VSS.n2773 107.24
R784 VSS.n1755 VSS.n960 106.731
R785 VSS.n2075 VSS.n2074 106.731
R786 VSS.n2225 VSS.n2224 106.731
R787 VSS.n2583 VSS.n2582 106.731
R788 VSS.n4197 VSS.n4196 106.678
R789 VSS.n3231 VSS.n3230 106.678
R790 VSS.n4959 VSS.n4958 106.678
R791 VSS.n197 VSS.n196 106.678
R792 VSS.n1437 VSS.n1436 106.678
R793 VSS.n3445 VSS.n3444 106.27
R794 VSS.n1051 VSS.n1050 106.27
R795 VSS.n946 VSS.n945 106.27
R796 VSS.n3626 VSS.t449 105.835
R797 VSS.n3366 VSS.t102 105.835
R798 VSS.n3731 VSS.t7 93.2783
R799 VSS.n3781 VSS.t162 93.2783
R800 VSS.n1219 VSS.t260 93.2783
R801 VSS.n891 VSS.t474 93.2783
R802 VSS.n2147 VSS.t567 93.2783
R803 VSS.n2653 VSS.t306 93.2783
R804 VSS.n2784 VSS.t339 93.2783
R805 VSS.n3295 VSS.t408 93.2779
R806 VSS.n3829 VSS.t557 93.2779
R807 VSS.n1682 VSS.t347 93.2779
R808 VSS.n2064 VSS.t471 93.2779
R809 VSS.n591 VSS.t67 93.2779
R810 VSS.n2728 VSS.t187 93.2779
R811 VSS.n2789 VSS.t427 93.2779
R812 VSS.n1062 VSS.n1057 92.7064
R813 VSS.n1069 VSS.n1054 92.7064
R814 VSS.n1084 VSS.n1080 92.7064
R815 VSS.n1139 VSS.n1135 92.7064
R816 VSS.n1155 VSS.n1151 92.7064
R817 VSS.n1209 VSS.n1205 92.7064
R818 VSS.n1229 VSS.n1225 92.7064
R819 VSS.n970 VSS.n966 92.7064
R820 VSS.n1647 VSS.n1643 92.7064
R821 VSS.n2080 VSS.n2079 92.7064
R822 VSS.n2213 VSS.n2212 92.7064
R823 VSS.n2199 VSS.n2198 92.7064
R824 VSS.n2185 VSS.n2184 92.7064
R825 VSS.n2168 VSS.n2167 92.7064
R826 VSS.n2154 VSS.n2153 92.7064
R827 VSS.n2131 VSS.n2130 92.7064
R828 VSS.n2117 VSS.n2116 92.7064
R829 VSS.n589 VSS.n588 92.7064
R830 VSS.n2590 VSS.n2589 92.7064
R831 VSS.n2604 VSS.n2603 92.7064
R832 VSS.n2621 VSS.n2620 92.7064
R833 VSS.n2635 VSS.n2634 92.7064
R834 VSS.n2650 VSS.n2649 92.7064
R835 VSS.n2662 VSS.n2661 92.7064
R836 VSS.n2682 VSS.n2681 92.7064
R837 VSS.n3374 VSS.t503 90.1413
R838 VSS.n3395 VSS.t631 90.1413
R839 VSS VSS.n3427 90.1413
R840 VSS.n3434 VSS.t101 90.1413
R841 VSS.n3457 VSS 90.1413
R842 VSS.n3579 VSS.t373 90.1413
R843 VSS.n3602 VSS.t644 90.1413
R844 VSS VSS.n3628 90.1413
R845 VSS.n3623 VSS.t448 90.1413
R846 VSS VSS.n3653 90.1413
R847 VSS.n1275 VSS.t2 88.8894
R848 VSS.n1950 VSS.t286 88.8894
R849 VSS.n173 VSS.t49 88.8894
R850 VSS.n390 VSS.t360 88.8894
R851 VSS.n2952 VSS.t452 88.8894
R852 VSS.n4545 VSS.t585 88.8894
R853 VSS.n4323 VSS.t689 88.8894
R854 VSS.n1781 VSS.n949 86.9123
R855 VSS.n936 VSS.n932 86.9123
R856 VSS.n1823 VSS.n1819 86.9123
R857 VSS.n1854 VSS.n1850 86.9123
R858 VSS.n1837 VSS.n1833 86.9123
R859 VSS.n899 VSS.n895 86.9123
R860 VSS.n914 VSS.n910 86.9123
R861 VSS.n1997 VSS.n1993 86.9123
R862 VSS VSS.n3497 84.5075
R863 VSS VSS.n3667 84.5075
R864 VSS.n4277 VSS.t580 81.4291
R865 VSS.n4055 VSS.t576 81.4291
R866 VSS.n2860 VSS.t555 81.4291
R867 VSS.n687 VSS.t141 81.4291
R868 VSS.n816 VSS.t302 81.4291
R869 VSS.n2385 VSS.t308 81.4291
R870 VSS.n1371 VSS.t713 81.4291
R871 VSS.n4361 VSS.t416 81.4291
R872 VSS.n4526 VSS.t341 81.4291
R873 VSS.n2926 VSS.t715 81.4291
R874 VSS.n365 VSS.t233 81.4291
R875 VSS.n5033 VSS.t18 81.4291
R876 VSS.n1943 VSS.t146 81.4291
R877 VSS.n1269 VSS.t634 81.4291
R878 VSS.n1154 VSS.t530 81.2313
R879 VSS.n1659 VSS.n1658 81.2313
R880 VSS.n1673 VSS.n1672 81.2313
R881 VSS.n1687 VSS.n1686 81.2313
R882 VSS.n1700 VSS.n1699 81.2313
R883 VSS.n1716 VSS.n1715 81.2313
R884 VSS.n1730 VSS.n1729 81.2313
R885 VSS.n1744 VSS.n1743 81.2313
R886 VSS.n957 VSS.n956 81.2313
R887 VSS.n1761 VSS.n1760 81.2313
R888 VSS.n2355 VSS.n2354 81.2313
R889 VSS.n2332 VSS.n2331 81.2313
R890 VSS.n2069 VSS.n2068 81.2313
R891 VSS.n2315 VSS.n2314 81.2313
R892 VSS.n2301 VSS.n2300 81.2313
R893 VSS.n2285 VSS.n2284 81.2313
R894 VSS.n2271 VSS.n2270 81.2313
R895 VSS.n2243 VSS.n2242 81.2313
R896 VSS.n2251 VSS.n2250 81.2313
R897 VSS.n4658 VSS.t367 81.2313
R898 VSS.n3870 VSS.t661 81.2313
R899 VSS.n1394 VSS.t710 80.4883
R900 VSS.n1377 VSS.t456 80.4883
R901 VSS.n850 VSS.t309 80.4883
R902 VSS.n2381 VSS.t560 80.4883
R903 VSS.n2484 VSS.t299 80.4883
R904 VSS.n814 VSS.t545 80.4883
R905 VSS.n717 VSS.t138 80.4883
R906 VSS.n699 VSS.t466 80.4883
R907 VSS.n2839 VSS.t552 80.4883
R908 VSS.n2856 VSS.t468 80.4883
R909 VSS.n4034 VSS.t573 80.4883
R910 VSS.n4051 VSS.t334 80.4883
R911 VSS.n4300 VSS.t577 80.4883
R912 VSS.n4283 VSS.t330 80.4883
R913 VSS.n1710 VSS.n1709 76.0005
R914 VSS.n2295 VSS.n2294 76.0005
R915 VSS.n3684 VSS.n3683 76.0005
R916 VSS.n3899 VSS.n3898 76.0005
R917 VSS.n3837 VSS.n3836 76.0005
R918 VSS.n3764 VSS.n3763 76.0005
R919 VSS.n1146 VSS.n1145 76.0005
R920 VSS.n1846 VSS.n1845 76.0005
R921 VSS.n2180 VSS.n2179 76.0005
R922 VSS.n2534 VSS.n2533 76.0005
R923 VSS.n2616 VSS.n2615 76.0005
R924 VSS.n2739 VSS.n2738 76.0005
R925 VSS.n4720 VSS.n4719 76.0005
R926 VSS.n2792 VSS.n2791 76.0005
R927 VSS.n3297 VSS.t704 74.2862
R928 VSS.n3748 VSS.t615 74.2862
R929 VSS.n3852 VSS.t312 74.2862
R930 VSS.n2822 VSS.t702 74.2862
R931 VSS.n4673 VSS.t668 74.2862
R932 VSS.n1050 VSS.t570 74.2862
R933 VSS.n960 VSS.t676 74.2862
R934 VSS.n945 VSS.t106 74.2862
R935 VSS.n2074 VSS.t603 74.2862
R936 VSS.n2224 VSS.t362 74.2862
R937 VSS.n2555 VSS.t404 74.2862
R938 VSS.n2582 VSS.t357 74.2862
R939 VSS.n2773 VSS.t544 74.2862
R940 VSS.n2779 VSS.t230 74.2862
R941 VSS.n3295 VSS.t314 70.4212
R942 VSS.n3829 VSS.t355 70.4212
R943 VSS.n1682 VSS.t607 70.4212
R944 VSS.n2064 VSS.t337 70.4212
R945 VSS.n591 VSS.t402 70.4212
R946 VSS.n2728 VSS.t639 70.4212
R947 VSS.n2789 VSS.t345 70.4212
R948 VSS.n3731 VSS.t25 70.4207
R949 VSS.n3781 VSS.t118 70.4207
R950 VSS.n1219 VSS.t120 70.4207
R951 VSS.n891 VSS.t160 70.4207
R952 VSS.n2147 VSS.t116 70.4207
R953 VSS.n2653 VSS.t77 70.4207
R954 VSS.n2784 VSS.t55 70.4207
R955 VSS.n1853 VSS.t514 67.6928
R956 VSS.n553 VSS.t489 67.6061
R957 VSS.n537 VSS.t501 67.6061
R958 VSS.n3515 VSS.t397 67.6061
R959 VSS.n3531 VSS.t371 67.6061
R960 VSS.n1791 VSS.n1790 65.5422
R961 VSS.n1661 VSS.n1657 63.7358
R962 VSS.n1675 VSS.n1671 63.7358
R963 VSS.n1689 VSS.n1685 63.7358
R964 VSS.n1702 VSS.n1698 63.7358
R965 VSS.n1718 VSS.n1714 63.7358
R966 VSS.n1732 VSS.n1728 63.7358
R967 VSS.n1746 VSS.n1742 63.7358
R968 VSS.n1763 VSS.n955 63.7358
R969 VSS.n2357 VSS.n2353 63.7358
R970 VSS.n2334 VSS.n2330 63.7358
R971 VSS.n2071 VSS.n2067 63.7358
R972 VSS.n2317 VSS.n2313 63.7358
R973 VSS.n2303 VSS.n2299 63.7358
R974 VSS.n2287 VSS.n2283 63.7358
R975 VSS.n2273 VSS.n2269 63.7358
R976 VSS.n2253 VSS.n2241 63.7358
R977 VSS.n3920 VSS.t217 57.1434
R978 VSS.n4018 VSS.t290 57.1434
R979 VSS.n442 VSS.t133 57.1434
R980 VSS.n735 VSS.t178 57.1434
R981 VSS.n2469 VSS.t431 57.1434
R982 VSS.n1928 VSS.t425 57.1434
R983 VSS.n1302 VSS.t252 57.1434
R984 VSS.n4196 VSS.t243 57.1434
R985 VSS.n3230 VSS.t152 57.1434
R986 VSS.n3021 VSS.t59 57.1434
R987 VSS.n4958 VSS.t599 57.1434
R988 VSS.n196 VSS.t439 57.1434
R989 VSS.n22 VSS.t680 57.1434
R990 VSS.n1436 VSS.t45 57.1434
R991 VSS.n2084 VSS.n2083 55.7517
R992 VSS.n586 VSS.n585 55.7517
R993 VSS.n4248 VSS.t241 54.2862
R994 VSS.n3953 VSS.t706 54.2862
R995 VSS.n3987 VSS.t213 54.2862
R996 VSS.n4574 VSS.t237 54.2862
R997 VSS.n4606 VSS.t288 54.2862
R998 VSS.n434 VSS.t37 54.2862
R999 VSS.n474 VSS.t129 54.2862
R1000 VSS.n679 VSS.t660 54.2862
R1001 VSS.n674 VSS.t176 54.2862
R1002 VSS.n2442 VSS.t85 54.2862
R1003 VSS.n2428 VSS.t433 54.2862
R1004 VSS.n1315 VSS.t35 54.2862
R1005 VSS.n1341 VSS.t421 54.2862
R1006 VSS.n1106 VSS.t318 54.2862
R1007 VSS.n997 VSS.t248 54.2862
R1008 VSS.n4396 VSS.t156 54.2862
R1009 VSS.n3251 VSS.t333 54.2862
R1010 VSS.n3099 VSS.t63 54.2862
R1011 VSS.n3051 VSS.t112 54.2862
R1012 VSS.n4921 VSS.t597 54.2862
R1013 VSS.n4935 VSS.t686 54.2862
R1014 VSS.n315 VSS.t437 54.2862
R1015 VSS.n292 VSS.t276 54.2862
R1016 VSS.n92 VSS.t684 54.2862
R1017 VSS.n72 VSS.t1 54.2862
R1018 VSS.n1508 VSS.t47 54.2862
R1019 VSS.n1487 VSS.t455 54.2862
R1020 VSS.n4228 VSS.t465 54.2862
R1021 VSS.t566 VSS.n2169 54.1543
R1022 VSS.t587 VSS.n2560 54.1543
R1023 VSS.t305 VSS.n2636 54.1543
R1024 VSS.n4747 VSS.t52 54.1543
R1025 VSS.n1271 VSS.t238 53.3338
R1026 VSS.n1582 VSS.t635 53.3338
R1027 VSS.n1945 VSS.t78 53.3338
R1028 VSS.n2027 VSS.t147 53.3338
R1029 VSS.n5035 VSS.t80 53.3338
R1030 VSS.n253 VSS.t15 53.3338
R1031 VSS.n374 VSS.t657 53.3338
R1032 VSS.n415 VSS.t234 53.3338
R1033 VSS.n2930 VSS.t707 53.3338
R1034 VSS.n2977 VSS.t716 53.3338
R1035 VSS.n4533 VSS.t38 53.3338
R1036 VSS.n4505 VSS.t342 53.3338
R1037 VSS.n4318 VSS.t263 53.3338
R1038 VSS.n4167 VSS.t417 53.3338
R1039 VSS.n1757 VSS.n959 51.0906
R1040 VSS.n2247 VSS.n2245 51.0906
R1041 VSS.n3380 VSS.t483 45.0709
R1042 VSS.n3389 VSS.t625 45.0709
R1043 VSS.n3305 VSS.t391 45.0709
R1044 VSS.n3596 VSS.t652 45.0709
R1045 VSS.n3296 VSS.n3295 41.945
R1046 VSS.n3830 VSS.n3829 41.945
R1047 VSS.n2785 VSS.n2784 41.945
R1048 VSS.n2790 VSS.n2789 41.945
R1049 VSS.n3738 VSS.n3731 41.7468
R1050 VSS.n3788 VSS.n3781 41.7468
R1051 VSS.n598 VSS.n591 41.7468
R1052 VSS.n2735 VSS.n2728 41.7468
R1053 VSS.n1719 VSS.n1710 41.6587
R1054 VSS.n2304 VSS.n2295 41.6587
R1055 VSS.n3685 VSS.n3684 41.6587
R1056 VSS.n3900 VSS.n3899 41.6587
R1057 VSS.n3838 VSS.n3837 41.6587
R1058 VSS.n3765 VSS.n3764 41.6587
R1059 VSS.n1147 VSS.n1146 41.6587
R1060 VSS.n1856 VSS.n1846 41.6587
R1061 VSS.n2182 VSS.n2180 41.6587
R1062 VSS.n2535 VSS.n2534 41.6587
R1063 VSS.n2618 VSS.n2616 41.6587
R1064 VSS.n2740 VSS.n2739 41.6587
R1065 VSS.n4721 VSS.n4720 41.6587
R1066 VSS.n2793 VSS.n2792 41.6587
R1067 VSS.n1691 VSS.n1682 41.4233
R1068 VSS.n901 VSS.n891 41.4233
R1069 VSS.n2073 VSS.n2064 41.4233
R1070 VSS.n2654 VSS.n2653 41.4233
R1071 VSS.n1220 VSS.n1219 41.1193
R1072 VSS.n2148 VSS.n2147 41.1193
R1073 VSS.n1701 VSS.t346 40.6159
R1074 VSS.n2316 VSS.t470 40.6159
R1075 VSS.n2134 VSS.t115 40.6159
R1076 VSS.n2665 VSS.t76 40.6159
R1077 VSS.n4135 VSS.t511 38.5719
R1078 VSS.n4135 VSS.t698 38.5719
R1079 VSS.n4277 VSS.t331 38.5719
R1080 VSS.n3920 VSS.t209 38.5719
R1081 VSS.n4085 VSS.t126 38.5719
R1082 VSS.n4085 VSS.t104 38.5719
R1083 VSS.n4055 VSS.t335 38.5719
R1084 VSS.n4018 VSS.t559 38.5719
R1085 VSS.n4625 VSS.t268 38.5719
R1086 VSS.n4625 VSS.t700 38.5719
R1087 VSS.n2860 VSS.t469 38.5719
R1088 VSS.n442 VSS.t23 38.5719
R1089 VSS.n4821 VSS.t673 38.5719
R1090 VSS.n4821 VSS.t224 38.5719
R1091 VSS.n687 VSS.t467 38.5719
R1092 VSS.n735 VSS.t329 38.5719
R1093 VSS.n663 VSS.t205 38.5719
R1094 VSS.n663 VSS.t410 38.5719
R1095 VSS.n816 VSS.t546 38.5719
R1096 VSS.n2469 VSS.t21 38.5719
R1097 VSS.n2415 VSS.t550 38.5719
R1098 VSS.n2415 VSS.t582 38.5719
R1099 VSS.n2385 VSS.t561 38.5719
R1100 VSS.n1928 VSS.t278 38.5719
R1101 VSS.n1351 VSS.t593 38.5719
R1102 VSS.n1351 VSS.t542 38.5719
R1103 VSS.n1371 VSS.t457 38.5719
R1104 VSS.n1302 VSS.t274 38.5719
R1105 VSS.n4196 VSS.t71 38.5719
R1106 VSS.n4361 VSS.t264 38.5719
R1107 VSS.n4411 VSS.t284 38.5719
R1108 VSS.n4411 VSS.t694 38.5719
R1109 VSS.n3230 VSS.t73 38.5719
R1110 VSS.n4526 VSS.t39 38.5719
R1111 VSS.n3142 VSS.t258 38.5719
R1112 VSS.n3142 VSS.t92 38.5719
R1113 VSS.n3021 VSS.t29 38.5719
R1114 VSS.n2926 VSS.t708 38.5719
R1115 VSS.n4879 VSS.t508 38.5719
R1116 VSS.n4879 VSS.t166 38.5719
R1117 VSS.n4958 VSS.t87 38.5719
R1118 VSS.n365 VSS.t658 38.5719
R1119 VSS.n282 VSS.t197 38.5719
R1120 VSS.n282 VSS.t564 38.5719
R1121 VSS.n196 VSS.t266 38.5719
R1122 VSS.n5033 VSS.t81 38.5719
R1123 VSS.n106 VSS.t135 38.5719
R1124 VSS.n106 VSS.t227 38.5719
R1125 VSS.n22 VSS.t316 38.5719
R1126 VSS.n1943 VSS.t79 38.5719
R1127 VSS.n1526 VSS.t304 38.5719
R1128 VSS.n1526 VSS.t191 38.5719
R1129 VSS.n1436 VSS.t27 38.5719
R1130 VSS.n1269 VSS.t239 38.5719
R1131 VSS.n1025 VSS.t609 38.5719
R1132 VSS.n1025 VSS.t181 38.5719
R1133 VSS.n1657 VSS.n1656 34.7652
R1134 VSS.n1671 VSS.n1670 34.7652
R1135 VSS.n1698 VSS.n1697 34.7652
R1136 VSS.n1714 VSS.n1713 34.7652
R1137 VSS.n1728 VSS.n1727 34.7652
R1138 VSS.n1742 VSS.n1741 34.7652
R1139 VSS.n959 VSS.n958 34.7652
R1140 VSS.n955 VSS.n954 34.7652
R1141 VSS.n2353 VSS.n2352 34.7652
R1142 VSS.n2330 VSS.n2329 34.7652
R1143 VSS.n2313 VSS.n2312 34.7652
R1144 VSS.n2299 VSS.n2298 34.7652
R1145 VSS.n2283 VSS.n2282 34.7652
R1146 VSS.n2269 VSS.n2268 34.7652
R1147 VSS.n2245 VSS.n2244 34.7652
R1148 VSS.n2241 VSS.n2240 34.7652
R1149 VSS.n3444 VSS.t33 33.462
R1150 VSS.n3444 VSS.t611 33.462
R1151 VSS.n3658 VSS.t9 33.462
R1152 VSS.n3658 VSS.t114 33.462
R1153 VSS.n2258 VSS.n2257 31.2934
R1154 VSS.n2085 VSS.n2084 28.1212
R1155 VSS.n587 VSS.n586 28.1212
R1156 VSS.n1208 VSS.t259 27.0774
R1157 VSS.n1784 VSS.n1783 27.0774
R1158 VSS.n1786 VSS.n1785 27.0774
R1159 VSS.n934 VSS.n933 27.0774
R1160 VSS.n1821 VSS.n1820 27.0774
R1161 VSS.n1852 VSS.n1851 27.0774
R1162 VSS.n1835 VSS.n1834 27.0774
R1163 VSS.n897 VSS.n896 27.0774
R1164 VSS.n912 VSS.n911 27.0774
R1165 VSS.n1995 VSS.n1994 27.0774
R1166 VSS.n4710 VSS.t54 27.0774
R1167 VSS.n4695 VSS.t344 27.0774
R1168 VSS.n3822 VSS.t354 27.0774
R1169 VSS.n3695 VSS.t313 27.0774
R1170 VSS.n1381 VSS.t547 26.8298
R1171 VSS.n2377 VSS.t253 26.8298
R1172 VSS.n799 VSS.t254 26.8298
R1173 VSS.n703 VSS.t669 26.8298
R1174 VSS.n2852 VSS.t696 26.8298
R1175 VSS.n4047 VSS.t472 26.8298
R1176 VSS.n4287 VSS.t88 26.8298
R1177 VSS.n4248 VSS.t296 25.9346
R1178 VSS.n3953 VSS.t215 25.9346
R1179 VSS.n3987 VSS.t406 25.9346
R1180 VSS.n4574 VSS.t292 25.9346
R1181 VSS.n4606 VSS.t31 25.9346
R1182 VSS.n434 VSS.t131 25.9346
R1183 VSS.n474 VSS.t199 25.9346
R1184 VSS.n679 VSS.t174 25.9346
R1185 VSS.n674 VSS.t5 25.9346
R1186 VSS.n2442 VSS.t429 25.9346
R1187 VSS.n2428 VSS.t613 25.9346
R1188 VSS.n1315 VSS.t423 25.9346
R1189 VSS.n1341 VSS.t678 25.9346
R1190 VSS.n1106 VSS.t250 25.9346
R1191 VSS.n997 VSS.t11 25.9346
R1192 VSS.n4396 VSS.t298 25.9346
R1193 VSS.n3251 VSS.t154 25.9346
R1194 VSS.n3099 VSS.t51 25.9346
R1195 VSS.n3051 VSS.t61 25.9346
R1196 VSS.n4921 VSS.t619 25.9346
R1197 VSS.n4935 VSS.t601 25.9346
R1198 VSS.n315 VSS.t272 25.9346
R1199 VSS.n292 VSS.t441 25.9346
R1200 VSS.n92 VSS.t94 25.9346
R1201 VSS.n72 VSS.t682 25.9346
R1202 VSS.n1508 VSS.t461 25.9346
R1203 VSS.n1487 VSS.t43 25.9346
R1204 VSS.n4228 VSS.t245 25.9346
R1205 VSS.n3297 VSS.t185 25.4291
R1206 VSS.n3748 VSS.t662 25.4291
R1207 VSS.n3852 VSS.t211 25.4291
R1208 VSS.n2822 VSS.t368 25.4291
R1209 VSS.n4673 VSS.t41 25.4291
R1210 VSS.n1050 VSS.t172 25.4291
R1211 VSS.n960 VSS.t641 25.4291
R1212 VSS.n945 VSS.t207 25.4291
R1213 VSS.n2074 VSS.t150 25.4291
R1214 VSS.n2224 VSS.t256 25.4291
R1215 VSS.n2555 VSS.t588 25.4291
R1216 VSS.n2582 VSS.t14 25.4291
R1217 VSS.n2773 VSS.t53 25.4291
R1218 VSS.n2779 VSS.t280 25.4291
R1219 VSS.n3475 VSS.t98 24.9236
R1220 VSS.n3475 VSS.t96 24.9236
R1221 VSS.n3461 VSS.t100 24.9236
R1222 VSS.n3461 VSS.t201 24.9236
R1223 VSS.n3513 VSS.t378 24.9236
R1224 VSS.n3513 VSS.t398 24.9236
R1225 VSS.n3523 VSS.t376 24.9236
R1226 VSS.n3523 VSS.t394 24.9236
R1227 VSS.n3529 VSS.t372 24.9236
R1228 VSS.n3529 VSS.t390 24.9236
R1229 VSS.n3536 VSS.t370 24.9236
R1230 VSS.n3536 VSS.t386 24.9236
R1231 VSS.n3330 VSS.t384 24.9236
R1232 VSS.n3330 VSS.t400 24.9236
R1233 VSS.n3573 VSS.t382 24.9236
R1234 VSS.n3573 VSS.t396 24.9236
R1235 VSS.n3303 VSS.t374 24.9236
R1236 VSS.n3303 VSS.t392 24.9236
R1237 VSS.n3314 VSS.t380 24.9236
R1238 VSS.n3314 VSS.t653 24.9236
R1239 VSS.n3600 VSS.t645 24.9236
R1240 VSS.n3600 VSS.t651 24.9236
R1241 VSS.n3611 VSS.t643 24.9236
R1242 VSS.n3611 VSS.t649 24.9236
R1243 VSS.n3637 VSS.t447 24.9236
R1244 VSS.n3637 VSS.t451 24.9236
R1245 VSS.n3644 VSS.t445 24.9236
R1246 VSS.n3644 VSS.t282 24.9236
R1247 VSS.n551 VSS.t496 24.9236
R1248 VSS.n551 VSS.t490 24.9236
R1249 VSS.n545 VSS.t506 24.9236
R1250 VSS.n545 VSS.t486 24.9236
R1251 VSS.n535 VSS.t502 24.9236
R1252 VSS.n535 VSS.t480 24.9236
R1253 VSS.n525 VSS.t498 24.9236
R1254 VSS.n525 VSS.t478 24.9236
R1255 VSS.n515 VSS.t494 24.9236
R1256 VSS.n515 VSS.t488 24.9236
R1257 VSS.n3368 VSS.t492 24.9236
R1258 VSS.n3368 VSS.t482 24.9236
R1259 VSS.n3378 VSS.t504 24.9236
R1260 VSS.n3378 VSS.t484 24.9236
R1261 VSS.n3384 VSS.t500 24.9236
R1262 VSS.n3384 VSS.t626 24.9236
R1263 VSS.n3393 VSS.t632 24.9236
R1264 VSS.n3393 VSS.t624 24.9236
R1265 VSS.n3403 VSS.t630 24.9236
R1266 VSS.n3403 VSS.t622 24.9236
R1267 VSS.n3288 VSS.n3285 24.0332
R1268 VSS.n3285 VSS.n3282 24.0332
R1269 VSS.n3282 VSS.n3279 24.0332
R1270 VSS.n3704 VSS.n3701 24.0332
R1271 VSS.n3707 VSS.n3704 24.0332
R1272 VSS.n3809 VSS.n3806 24.0332
R1273 VSS.n3806 VSS.n3803 24.0332
R1274 VSS.n3803 VSS.n3800 24.0332
R1275 VSS.n3800 VSS.n3797 24.0332
R1276 VSS.n3817 VSS.n3814 24.0332
R1277 VSS.n1639 VSS.n1636 24.0332
R1278 VSS.n1636 VSS.n1633 24.0332
R1279 VSS.n1633 VSS.n1630 24.0332
R1280 VSS.n1630 VSS.n1627 24.0332
R1281 VSS.n1770 VSS.n1767 24.0332
R1282 VSS.n1989 VSS.n1986 24.0332
R1283 VSS.n1986 VSS.n1983 24.0332
R1284 VSS.n2346 VSS.n2343 24.0332
R1285 VSS.n2349 VSS.n2346 24.0332
R1286 VSS.n2113 VSS.n2110 24.0332
R1287 VSS.n2110 VSS.n2107 24.0332
R1288 VSS.n615 VSS.n612 24.0332
R1289 VSS.n618 VSS.n615 24.0332
R1290 VSS.n621 VSS.n618 24.0332
R1291 VSS.n2678 VSS.n2675 24.0332
R1292 VSS.n2697 VSS.n2694 24.0332
R1293 VSS.n2700 VSS.n2697 24.0332
R1294 VSS.n2703 VSS.n2700 24.0332
R1295 VSS.n2706 VSS.n2703 24.0332
R1296 VSS.n2563 VSS.n2551 23.7899
R1297 VSS.n4744 VSS.n4743 23.7899
R1298 VSS.n3865 VSS.n3862 23.7089
R1299 VSS.n1640 VSS.n1639 23.245
R1300 VSS.n1990 VSS.n1989 22.9432
R1301 VSS.n547 VSS.t505 22.5357
R1302 VSS.n541 VSS.t485 22.5357
R1303 VSS.n3519 VSS.t375 22.5357
R1304 VSS.n3525 VSS.t393 22.5357
R1305 VSS.n2066 VSS.n2065 22.2537
R1306 VSS.n1684 VSS.n1683 22.2537
R1307 VSS.n3710 VSS.n3707 22.1686
R1308 VSS.n3862 VSS.n3859 22.1686
R1309 VSS.n3820 VSS.n3817 22.1686
R1310 VSS.n4667 VSS.n4666 22.1686
R1311 VSS.n4743 VSS.n4740 22.1686
R1312 VSS.n4704 VSS.n4701 22.1686
R1313 VSS.n1654 VSS.n1653 21.7362
R1314 VSS.n2350 VSS.n2349 21.7362
R1315 VSS.n3631 VSS.n3622 20.3039
R1316 VSS.n2114 VSS.n2113 18.7186
R1317 VSS.n2679 VSS.n2678 18.7186
R1318 VSS.n2551 VSS.n590 18.1151
R1319 VSS.n1279 VSS.t568 17.7783
R1320 VSS.n1955 VSS.t709 17.7783
R1321 VSS.n167 VSS.t188 17.7783
R1322 VSS.n370 VSS.t637 17.7783
R1323 VSS.n2946 VSS.t419 17.7783
R1324 VSS.n4539 VSS.t183 17.7783
R1325 VSS.n4328 VSS.t358 17.7783
R1326 VSS.n3454 VSS 16.7729
R1327 VSS.n3656 VSS 16.7729
R1328 VSS.n4093 VSS 16.5522
R1329 VSS.n4619 VSS 16.5522
R1330 VSS VSS.n766 16.5522
R1331 VSS.n2423 VSS 16.5522
R1332 VSS.n1771 VSS.n1770 15.0975
R1333 VSS.n1767 VSS.n950 13.8904
R1334 VSS.n1065 VSS.n1064 13.539
R1335 VSS.n1067 VSS.n1066 13.539
R1336 VSS.n1082 VSS.n1081 13.539
R1337 VSS.n1137 VSS.n1136 13.539
R1338 VSS.n1153 VSS.n1152 13.539
R1339 VSS.n1207 VSS.n1206 13.539
R1340 VSS.n1227 VSS.n1226 13.539
R1341 VSS.n968 VSS.n967 13.539
R1342 VSS.n1645 VSS.n1644 13.539
R1343 VSS.n1717 VSS.t528 13.539
R1344 VSS.n1836 VSS.t473 13.539
R1345 VSS.n2302 VSS.t524 13.539
R1346 VSS.n2231 VSS.n2230 13.539
R1347 VSS.n2228 VSS.n2082 13.539
R1348 VSS.n2216 VSS.n2215 13.539
R1349 VSS.n2202 VSS.n2201 13.539
R1350 VSS.n2188 VSS.n2187 13.539
R1351 VSS.n2171 VSS.n2170 13.539
R1352 VSS.n2151 VSS.n2150 13.539
R1353 VSS.n2134 VSS.n2133 13.539
R1354 VSS.n2120 VSS.n2119 13.539
R1355 VSS.n2574 VSS.n2573 13.539
R1356 VSS.n2578 VSS.n2577 13.539
R1357 VSS.n2593 VSS.n2592 13.539
R1358 VSS.n2607 VSS.n2606 13.539
R1359 VSS.n2624 VSS.n2623 13.539
R1360 VSS.n2638 VSS.n2637 13.539
R1361 VSS.n2647 VSS.n2646 13.539
R1362 VSS.n2665 VSS.n2664 13.539
R1363 VSS.n2685 VSS.n2684 13.539
R1364 VSS.n4826 VSS 13.4626
R1365 VSS.n4740 VSS.n2778 12.5798
R1366 VSS.n3810 VSS.n3809 12.242
R1367 VSS.n3873 VSS.n3872 11.9177
R1368 VSS.n4661 VSS.n4660 11.9177
R1369 VSS.n2710 VSS.n2706 11.7196
R1370 VSS.n949 VSS.n948 11.5887
R1371 VSS.n1790 VSS.n1789 11.5887
R1372 VSS.n932 VSS.n931 11.5887
R1373 VSS.n1819 VSS.n1818 11.5887
R1374 VSS.n1850 VSS.n1849 11.5887
R1375 VSS.n1833 VSS.n1832 11.5887
R1376 VSS.n910 VSS.n909 11.5887
R1377 VSS.n1993 VSS.n1992 11.5887
R1378 VSS.n622 VSS.n621 11.4989
R1379 VSS.n1685 VSS.n1684 11.1906
R1380 VSS.n2067 VSS.n2066 11.1906
R1381 VSS.n818 VSS.n817 10.5936
R1382 VSS.n5037 VSS.n5034 10.5936
R1383 VSS.n1947 VSS.n1944 10.5936
R1384 VSS.n1273 VSS.n1270 10.5936
R1385 VSS.n3289 VSS.n3288 10.2558
R1386 VSS.n3527 VSS.n3524 10.1522
R1387 VSS.n549 VSS.n546 10.1522
R1388 VSS.n2581 VSS.n2580 9.93153
R1389 VSS.n4281 VSS.n4278 9.71084
R1390 VSS.n4059 VSS.n4056 9.71084
R1391 VSS.n2864 VSS.n2861 9.71084
R1392 VSS.n2389 VSS.n2386 9.71084
R1393 VSS.n1375 VSS.n1372 9.71084
R1394 VSS.n4365 VSS.n4362 9.71084
R1395 VSS.n4530 VSS.n4527 9.71084
R1396 VSS.n2136 VSS.n2135 9.3005
R1397 VSS.n2135 VSS.n2134 9.3005
R1398 VSS.n2152 VSS.n2151 9.3005
R1399 VSS.n2173 VSS.n2172 9.3005
R1400 VSS.n2172 VSS.n2171 9.3005
R1401 VSS.n2190 VSS.n2189 9.3005
R1402 VSS.n2189 VSS.n2188 9.3005
R1403 VSS.n2204 VSS.n2203 9.3005
R1404 VSS.n2203 VSS.n2202 9.3005
R1405 VSS.n2218 VSS.n2217 9.3005
R1406 VSS.n2217 VSS.n2216 9.3005
R1407 VSS.n2227 VSS.n2226 9.3005
R1408 VSS.n2228 VSS.n2227 9.3005
R1409 VSS.n2233 VSS.n2232 9.3005
R1410 VSS.n2232 VSS.n2231 9.3005
R1411 VSS.n2254 VSS.n2253 9.3005
R1412 VSS.n2253 VSS.n2252 9.3005
R1413 VSS.n2249 VSS.n2248 9.3005
R1414 VSS.n2274 VSS.n2273 9.3005
R1415 VSS.n2273 VSS.n2272 9.3005
R1416 VSS.n2288 VSS.n2287 9.3005
R1417 VSS.n2287 VSS.n2286 9.3005
R1418 VSS.n2304 VSS.n2303 9.3005
R1419 VSS.n2303 VSS.n2302 9.3005
R1420 VSS.n2318 VSS.n2317 9.3005
R1421 VSS.n2317 VSS.n2316 9.3005
R1422 VSS.n2072 VSS.n2071 9.3005
R1423 VSS.n2071 VSS.n2070 9.3005
R1424 VSS.n2335 VSS.n2334 9.3005
R1425 VSS.n2334 VSS.n2333 9.3005
R1426 VSS.n2358 VSS.n2357 9.3005
R1427 VSS.n2357 VSS.n2356 9.3005
R1428 VSS.n1998 VSS.n1997 9.3005
R1429 VSS.n1997 VSS.n1996 9.3005
R1430 VSS.n915 VSS.n914 9.3005
R1431 VSS.n914 VSS.n913 9.3005
R1432 VSS.n900 VSS.n899 9.3005
R1433 VSS.n899 VSS.n898 9.3005
R1434 VSS.n1838 VSS.n1837 9.3005
R1435 VSS.n1837 VSS.n1836 9.3005
R1436 VSS.n1855 VSS.n1854 9.3005
R1437 VSS.n1854 VSS.n1853 9.3005
R1438 VSS.n1824 VSS.n1823 9.3005
R1439 VSS.n1823 VSS.n1822 9.3005
R1440 VSS.n937 VSS.n936 9.3005
R1441 VSS.n936 VSS.n935 9.3005
R1442 VSS.n1788 VSS.n1787 9.3005
R1443 VSS.n1781 VSS.n1780 9.3005
R1444 VSS.n1782 VSS.n1781 9.3005
R1445 VSS.n1764 VSS.n1763 9.3005
R1446 VSS.n1763 VSS.n1762 9.3005
R1447 VSS.n1759 VSS.n1758 9.3005
R1448 VSS.n1747 VSS.n1746 9.3005
R1449 VSS.n1746 VSS.n1745 9.3005
R1450 VSS.n1733 VSS.n1732 9.3005
R1451 VSS.n1732 VSS.n1731 9.3005
R1452 VSS.n1719 VSS.n1718 9.3005
R1453 VSS.n1718 VSS.n1717 9.3005
R1454 VSS.n1703 VSS.n1702 9.3005
R1455 VSS.n1702 VSS.n1701 9.3005
R1456 VSS.n1690 VSS.n1689 9.3005
R1457 VSS.n1689 VSS.n1688 9.3005
R1458 VSS.n1676 VSS.n1675 9.3005
R1459 VSS.n1675 VSS.n1674 9.3005
R1460 VSS.n1662 VSS.n1661 9.3005
R1461 VSS.n1661 VSS.n1660 9.3005
R1462 VSS.n1649 VSS.n1648 9.3005
R1463 VSS.n1648 VSS.n1647 9.3005
R1464 VSS.n1647 VSS.n1646 9.3005
R1465 VSS.n971 VSS.n970 9.3005
R1466 VSS.n970 VSS.n969 9.3005
R1467 VSS.n1230 VSS.n1229 9.3005
R1468 VSS.n1229 VSS.n1228 9.3005
R1469 VSS.n1210 VSS.n1209 9.3005
R1470 VSS.n1209 VSS.n1208 9.3005
R1471 VSS.n1157 VSS.n1156 9.3005
R1472 VSS.n1156 VSS.n1155 9.3005
R1473 VSS.n1155 VSS.n1154 9.3005
R1474 VSS.n1140 VSS.n1139 9.3005
R1475 VSS.n1139 VSS.n1138 9.3005
R1476 VSS.n1085 VSS.n1084 9.3005
R1477 VSS.n1084 VSS.n1083 9.3005
R1478 VSS.n1072 VSS.n1069 9.3005
R1479 VSS.n1069 VSS.n1068 9.3005
R1480 VSS.n1062 VSS.n1061 9.3005
R1481 VSS.n1063 VSS.n1062 9.3005
R1482 VSS.n2581 VSS.n2579 9.3005
R1483 VSS.n2579 VSS.n2578 9.3005
R1484 VSS.n2609 VSS.n2608 9.3005
R1485 VSS.n2608 VSS.n2607 9.3005
R1486 VSS.n2640 VSS.n2639 9.3005
R1487 VSS.n2639 VSS.n2638 9.3005
R1488 VSS.n2667 VSS.n2666 9.3005
R1489 VSS.n2666 VSS.n2665 9.3005
R1490 VSS.n2687 VSS.n2686 9.3005
R1491 VSS.n2686 VSS.n2685 9.3005
R1492 VSS.n2648 VSS.n2647 9.3005
R1493 VSS.n2626 VSS.n2625 9.3005
R1494 VSS.n2625 VSS.n2624 9.3005
R1495 VSS.n2595 VSS.n2594 9.3005
R1496 VSS.n2594 VSS.n2593 9.3005
R1497 VSS.n2572 VSS.n2571 9.3005
R1498 VSS.n2573 VSS.n2572 9.3005
R1499 VSS.n2122 VSS.n2121 9.3005
R1500 VSS.n2121 VSS.n2120 9.3005
R1501 VSS.n3387 VSS.n3385 9.26947
R1502 VSS.n2928 VSS.n2927 9.26947
R1503 VSS.n473 VSS.n472 9.01861
R1504 VSS.n2427 VSS.n2426 9.01861
R1505 VSS.n3250 VSS.n3249 9.01852
R1506 VSS.n4939 VSS.n4938 9.01852
R1507 VSS.n3636 VSS.n3635 9.01832
R1508 VSS.n4820 VSS.n4819 9.01832
R1509 VSS.n4410 VSS.n4375 9.01832
R1510 VSS.n485 VSS.n484 9.01815
R1511 VSS.n4426 VSS.n4425 9.01815
R1512 VSS.n1544 VSS.n1543 9.01815
R1513 VSS.n4247 VSS.n4246 9.01761
R1514 VSS.n3986 VSS.n3985 9.01761
R1515 VSS.n4605 VSS.n4604 9.01761
R1516 VSS.n673 VSS.n672 9.01761
R1517 VSS.n1340 VSS.n1339 9.01761
R1518 VSS.n4395 VSS.n4394 9.01761
R1519 VSS.n3098 VSS.n3097 9.01761
R1520 VSS.n4920 VSS.n4919 9.01761
R1521 VSS.n314 VSS.n313 9.01761
R1522 VSS.n96 VSS.n95 9.01761
R1523 VSS.n1507 VSS.n1506 9.01761
R1524 VSS.n4232 VSS.n4231 9.01754
R1525 VSS.n3952 VSS.n3951 9.01752
R1526 VSS.n4573 VSS.n4572 9.01752
R1527 VSS.n433 VSS.n432 9.01752
R1528 VSS.n678 VSS.n677 9.01752
R1529 VSS.n2441 VSS.n2440 9.01752
R1530 VSS.n1314 VSS.n1313 9.01752
R1531 VSS.n3055 VSS.n3054 9.01752
R1532 VSS.n291 VSS.n290 9.01752
R1533 VSS.n71 VSS.n70 9.01752
R1534 VSS.n1491 VSS.n1490 9.01752
R1535 VSS.n3661 VSS.n3660 9.01734
R1536 VSS.n3448 VSS.n3447 9.01732
R1537 VSS.n4138 VSS.n4137 9.01732
R1538 VSS.n4084 VSS.n4083 9.01732
R1539 VSS.n4624 VSS.n4623 9.01732
R1540 VSS.n667 VSS.n666 9.01732
R1541 VSS.n2414 VSS.n2413 9.01732
R1542 VSS.n1350 VSS.n1349 9.01732
R1543 VSS.n3141 VSS.n3116 9.01732
R1544 VSS.n4912 VSS.n4911 9.01732
R1545 VSS.n324 VSS.n323 9.01732
R1546 VSS.n109 VSS.n108 9.01732
R1547 VSS.n1525 VSS.n1524 9.01732
R1548 VSS.n1024 VSS.n1023 9.01732
R1549 VSS.n4133 VSS.n4132 9.01716
R1550 VSS.n4075 VSS.n4074 9.01716
R1551 VSS.n4593 VSS.n4592 9.01716
R1552 VSS.n776 VSS.n775 9.01716
R1553 VSS.n2405 VSS.n2404 9.01716
R1554 VSS.n1307 VSS.n1306 9.01716
R1555 VSS.n3148 VSS.n3147 9.01716
R1556 VSS.n4887 VSS.n4886 9.01716
R1557 VSS.n5004 VSS.n5003 9.01716
R1558 VSS.n128 VSS.n127 9.01716
R1559 VSS.n1031 VSS.n1030 9.01716
R1560 VSS.n996 VSS.n995 9.01662
R1561 VSS.n1105 VSS.n1104 9.01654
R1562 VSS.n3474 VSS.n3473 9.01634
R1563 VSS.n3300 VSS.n3299 9.01634
R1564 VSS.n3855 VSS.n3854 9.01634
R1565 VSS.n4672 VSS.n4671 9.01634
R1566 VSS.n4736 VSS.n2778 9.01634
R1567 VSS.n3294 VSS.n3293 9.01549
R1568 VSS.n3828 VSS.n3827 9.01549
R1569 VSS.n2783 VSS.n2782 9.01549
R1570 VSS.n2788 VSS.n2787 9.01549
R1571 VSS.n3436 VSS.n3435 9.01392
R1572 VSS.n3435 VSS.n3434 9.01392
R1573 VSS.n3465 VSS.n3464 9.01392
R1574 VSS.n3459 VSS.n3458 9.01392
R1575 VSS.n3455 VSS.n3454 9.01392
R1576 VSS.n3470 VSS.n3469 9.01392
R1577 VSS.n503 VSS.n502 9.01392
R1578 VSS.n508 VSS.n507 9.01392
R1579 VSS.n561 VSS.n560 9.01392
R1580 VSS.n555 VSS.n554 9.01392
R1581 VSS.n549 VSS.n548 9.01392
R1582 VSS.n543 VSS.n542 9.01392
R1583 VSS.n539 VSS.n538 9.01392
R1584 VSS.n533 VSS.n532 9.01392
R1585 VSS.n529 VSS.n528 9.01392
R1586 VSS.n523 VSS.n522 9.01392
R1587 VSS.n519 VSS.n518 9.01392
R1588 VSS.n513 VSS.n512 9.01392
R1589 VSS.n3372 VSS.n3371 9.01392
R1590 VSS.n3376 VSS.n3375 9.01392
R1591 VSS.n3382 VSS.n3381 9.01392
R1592 VSS.n3387 VSS.n3386 9.01392
R1593 VSS.n3386 VSS.t499 9.01392
R1594 VSS.n3391 VSS.n3390 9.01392
R1595 VSS.n3397 VSS.n3396 9.01392
R1596 VSS.n3401 VSS.n3400 9.01392
R1597 VSS.n3407 VSS.n3406 9.01392
R1598 VSS.n3413 VSS.n3412 9.01392
R1599 VSS.n3426 VSS.n3425 9.01392
R1600 VSS.n3430 VSS.n3429 9.01392
R1601 VSS.n3660 VSS.n3659 9.01392
R1602 VSS.n3502 VSS.n3501 9.01392
R1603 VSS.n3507 VSS.n3506 9.01392
R1604 VSS.n3511 VSS.n3510 9.01392
R1605 VSS.n3517 VSS.n3516 9.01392
R1606 VSS.n3521 VSS.n3520 9.01392
R1607 VSS.n3527 VSS.n3526 9.01392
R1608 VSS.n3533 VSS.n3532 9.01392
R1609 VSS.n3546 VSS.n3545 9.01392
R1610 VSS.n3540 VSS.n3539 9.01392
R1611 VSS.n3326 VSS.n3325 9.01392
R1612 VSS.n3335 VSS.n3334 9.01392
R1613 VSS.n3570 VSS.n3569 9.01392
R1614 VSS.n3577 VSS.n3576 9.01392
R1615 VSS.n3581 VSS.n3580 9.01392
R1616 VSS.n3307 VSS.n3306 9.01392
R1617 VSS.n3312 VSS.n3311 9.01392
R1618 VSS.n3311 VSS.t379 9.01392
R1619 VSS.n3598 VSS.n3597 9.01392
R1620 VSS.n3604 VSS.n3603 9.01392
R1621 VSS.n3609 VSS.n3608 9.01392
R1622 VSS.n3615 VSS.n3614 9.01392
R1623 VSS.n3619 VSS.n3618 9.01392
R1624 VSS.n3627 VSS.n3622 9.01392
R1625 VSS.n3631 VSS.n3630 9.01392
R1626 VSS.n3625 VSS.n3624 9.01392
R1627 VSS.n3642 VSS.n3641 9.01392
R1628 VSS.n3648 VSS.n3647 9.01392
R1629 VSS.n3652 VSS.n3651 9.01392
R1630 VSS.n3656 VSS.n3655 9.01392
R1631 VSS.n3697 VSS.n3696 9.01392
R1632 VSS.n3692 VSS.n3691 9.01392
R1633 VSS.n3688 VSS.n3687 9.01392
R1634 VSS.n3681 VSS.n3680 9.01392
R1635 VSS.n3677 VSS.n3676 9.01392
R1636 VSS.n3710 VSS.n3709 9.01392
R1637 VSS.n3859 VSS.n3858 9.01392
R1638 VSS.n3849 VSS.n3848 9.01392
R1639 VSS.n3845 VSS.n3844 9.01392
R1640 VSS.n3834 VSS.n3833 9.01392
R1641 VSS.n4668 VSS.n4667 9.01392
R1642 VSS.n4697 VSS.n4696 9.01392
R1643 VSS.n2802 VSS.n2801 9.01392
R1644 VSS.n2796 VSS.n2795 9.01392
R1645 VSS.n2815 VSS.n2814 9.01392
R1646 VSS.n4678 VSS.n4677 9.01392
R1647 VSS.n4704 VSS.n4703 9.01392
R1648 VSS.n4732 VSS.n4731 9.01392
R1649 VSS.n4728 VSS.n4727 9.01392
R1650 VSS.n4724 VSS.n4723 9.01392
R1651 VSS.n4717 VSS.n4716 9.01392
R1652 VSS.n4712 VSS.n4711 9.01392
R1653 VSS.n4708 VSS.n4707 9.01392
R1654 VSS.n4740 VSS.n4739 9.01392
R1655 VSS.n992 VSS.n991 9.01392
R1656 VSS.n991 VSS.n990 9.01392
R1657 VSS.n1408 VSS.n1407 9.01392
R1658 VSS.n1036 VSS.n1035 9.01392
R1659 VSS.n1035 VSS.n1034 9.01392
R1660 VSS.n4239 VSS.n4238 9.01392
R1661 VSS.n4231 VSS.n4230 9.01392
R1662 VSS.n3429 VSS.n3428 9.01392
R1663 VSS.n3427 VSS.n3426 9.01392
R1664 VSS.n3412 VSS.n3411 9.01392
R1665 VSS.n3406 VSS.n3405 9.01392
R1666 VSS.n3400 VSS.n3399 9.01392
R1667 VSS.n3396 VSS.n3395 9.01392
R1668 VSS.n3390 VSS.n3389 9.01392
R1669 VSS.n3381 VSS.n3380 9.01392
R1670 VSS.n3375 VSS.n3374 9.01392
R1671 VSS.n3371 VSS.n3370 9.01392
R1672 VSS.n512 VSS.n511 9.01392
R1673 VSS.n518 VSS.n517 9.01392
R1674 VSS.n522 VSS.n521 9.01392
R1675 VSS.n528 VSS.n527 9.01392
R1676 VSS.n532 VSS.n531 9.01392
R1677 VSS.n538 VSS.n537 9.01392
R1678 VSS.n542 VSS.n541 9.01392
R1679 VSS.n548 VSS.n547 9.01392
R1680 VSS.n554 VSS.n553 9.01392
R1681 VSS.n560 VSS.n559 9.01392
R1682 VSS.n507 VSS.n506 9.01392
R1683 VSS.n502 VSS.n501 9.01392
R1684 VSS.n3469 VSS.n3468 9.01392
R1685 VSS.n3464 VSS.n3463 9.01392
R1686 VSS.n3458 VSS.n3457 9.01392
R1687 VSS.n3456 VSS.n3455 9.01392
R1688 VSS.n3447 VSS.n3446 9.01392
R1689 VSS.n3496 VSS.n3495 9.01392
R1690 VSS.n3497 VSS.n3496 9.01392
R1691 VSS.n3473 VSS.n3472 9.01392
R1692 VSS.n3655 VSS.n3654 9.01392
R1693 VSS.n3653 VSS.n3652 9.01392
R1694 VSS.n3647 VSS.n3646 9.01392
R1695 VSS.n3641 VSS.n3640 9.01392
R1696 VSS.n3635 VSS.n3634 9.01392
R1697 VSS.n3624 VSS.n3623 9.01392
R1698 VSS.n3630 VSS.n3629 9.01392
R1699 VSS.n3628 VSS.n3627 9.01392
R1700 VSS.n3618 VSS.n3617 9.01392
R1701 VSS.n3614 VSS.n3613 9.01392
R1702 VSS.n3608 VSS.n3607 9.01392
R1703 VSS.n3603 VSS.n3602 9.01392
R1704 VSS.n3597 VSS.n3596 9.01392
R1705 VSS.n3306 VSS.n3305 9.01392
R1706 VSS.n3580 VSS.n3579 9.01392
R1707 VSS.n3576 VSS.n3575 9.01392
R1708 VSS.n3569 VSS.n3568 9.01392
R1709 VSS.n3334 VSS.n3333 9.01392
R1710 VSS.n3325 VSS.n3324 9.01392
R1711 VSS.n3539 VSS.n3538 9.01392
R1712 VSS.n3545 VSS.n3544 9.01392
R1713 VSS.n3532 VSS.n3531 9.01392
R1714 VSS.n3526 VSS.n3525 9.01392
R1715 VSS.n3520 VSS.n3519 9.01392
R1716 VSS.n3516 VSS.n3515 9.01392
R1717 VSS.n3510 VSS.n3509 9.01392
R1718 VSS.n3506 VSS.n3505 9.01392
R1719 VSS.n3666 VSS.n3665 9.01392
R1720 VSS.n3667 VSS.n3666 9.01392
R1721 VSS.n3501 VSS.n3500 9.01392
R1722 VSS.n4739 VSS.n4738 9.01392
R1723 VSS.n4737 VSS.n4736 9.01392
R1724 VSS.n4731 VSS.n4730 9.01392
R1725 VSS.n4727 VSS.n4726 9.01392
R1726 VSS.n4723 VSS.n4722 9.01392
R1727 VSS.n4716 VSS.n4715 9.01392
R1728 VSS.n2782 VSS.n2781 9.01392
R1729 VSS.n4711 VSS.n4710 9.01392
R1730 VSS.n4707 VSS.n4706 9.01392
R1731 VSS.n4703 VSS.n4702 9.01392
R1732 VSS.n4696 VSS.n4695 9.01392
R1733 VSS.n2787 VSS.n2786 9.01392
R1734 VSS.n2801 VSS.n2800 9.01392
R1735 VSS.n2795 VSS.n2794 9.01392
R1736 VSS.n2814 VSS.n2813 9.01392
R1737 VSS.n4677 VSS.n4676 9.01392
R1738 VSS.n4669 VSS.n4668 9.01392
R1739 VSS.n3827 VSS.n3826 9.01392
R1740 VSS.n3833 VSS.n3832 9.01392
R1741 VSS.n3844 VSS.n3843 9.01392
R1742 VSS.n3848 VSS.n3847 9.01392
R1743 VSS.n3858 VSS.n3857 9.01392
R1744 VSS.n3709 VSS.n3708 9.01392
R1745 VSS.n3696 VSS.n3695 9.01392
R1746 VSS.n3293 VSS.n3292 9.01392
R1747 VSS.n3691 VSS.n3690 9.01392
R1748 VSS.n3687 VSS.n3686 9.01392
R1749 VSS.n3680 VSS.n3679 9.01392
R1750 VSS.n3676 VSS.n3675 9.01392
R1751 VSS.n3301 VSS.n3300 9.01392
R1752 VSS.n3672 VSS.n3671 9.01392
R1753 VSS.n3671 VSS.n3670 9.01392
R1754 VSS.n3856 VSS.n3855 9.01392
R1755 VSS.n3841 VSS.n3840 9.01392
R1756 VSS.n3840 VSS.n3839 9.01392
R1757 VSS.n3824 VSS.n3823 9.01392
R1758 VSS.n3823 VSS.n3822 9.01392
R1759 VSS.n3820 VSS.n3819 9.01392
R1760 VSS.n3819 VSS.n3818 9.01392
R1761 VSS.n4671 VSS.n4670 9.01392
R1762 VSS.n1030 VSS.n1029 9.01392
R1763 VSS.n1177 VSS.n1176 9.01392
R1764 VSS.n1176 VSS.n1175 9.01392
R1765 VSS.n1188 VSS.n1186 9.01392
R1766 VSS.n1186 VSS.n1185 9.01392
R1767 VSS.n1266 VSS.n1265 9.01392
R1768 VSS.n1265 VSS.n1264 9.01392
R1769 VSS.n1273 VSS.n1272 9.01392
R1770 VSS.n1272 VSS.n1271 9.01392
R1771 VSS.n1281 VSS.n1280 9.01392
R1772 VSS.n1280 VSS.n1279 9.01392
R1773 VSS.n1580 VSS.n1578 9.01392
R1774 VSS.n1578 VSS.n1577 9.01392
R1775 VSS.n1584 VSS.n1583 9.01392
R1776 VSS.n1583 VSS.n1582 9.01392
R1777 VSS.n1595 VSS.n1593 9.01392
R1778 VSS.n1593 VSS.n1592 9.01392
R1779 VSS.n1426 VSS.n1425 9.01392
R1780 VSS.n1425 VSS.n1424 9.01392
R1781 VSS.n1434 VSS.n1432 9.01392
R1782 VSS.n1432 VSS.n1431 9.01392
R1783 VSS.n1453 VSS.n1452 9.01392
R1784 VSS.n1452 VSS.n1451 9.01392
R1785 VSS.n1457 VSS.n1456 9.01392
R1786 VSS.n1456 VSS.n1455 9.01392
R1787 VSS.n1490 VSS.n1489 9.01392
R1788 VSS.n1498 VSS.n1497 9.01392
R1789 VSS.n1497 VSS.n1496 9.01392
R1790 VSS.n1506 VSS.n1505 9.01392
R1791 VSS.n1512 VSS.n1511 9.01392
R1792 VSS.n1511 VSS.n1477 9.01392
R1793 VSS.n1524 VSS.n1523 9.01392
R1794 VSS.n1532 VSS.n1531 9.01392
R1795 VSS.n1531 VSS.n1530 9.01392
R1796 VSS.n1898 VSS.n1897 9.01392
R1797 VSS.n1897 VSS.n1896 9.01392
R1798 VSS.n1905 VSS.n1903 9.01392
R1799 VSS.n1903 VSS.n1902 9.01392
R1800 VSS.n1947 VSS.n1946 9.01392
R1801 VSS.n1946 VSS.n1945 9.01392
R1802 VSS.n1957 VSS.n1956 9.01392
R1803 VSS.n1956 VSS.n1955 9.01392
R1804 VSS.n1952 VSS.n1951 9.01392
R1805 VSS.n1951 VSS.n1950 9.01392
R1806 VSS.n2018 VSS.n2016 9.01392
R1807 VSS.n2016 VSS.n2015 9.01392
R1808 VSS.n2029 VSS.n2028 9.01392
R1809 VSS.n2028 VSS.n2027 9.01392
R1810 VSS.n5 VSS.n4 9.01392
R1811 VSS.n4 VSS.n3 9.01392
R1812 VSS.n9 VSS.n8 9.01392
R1813 VSS.n8 VSS.n7 9.01392
R1814 VSS.n14 VSS.n13 9.01392
R1815 VSS.n13 VSS.n12 9.01392
R1816 VSS.n48 VSS.n47 9.01392
R1817 VSS.n47 VSS.n46 9.01392
R1818 VSS.n82 VSS.n81 9.01392
R1819 VSS.n81 VSS.n80 9.01392
R1820 VSS.n95 VSS.n94 9.01392
R1821 VSS.n112 VSS.n111 9.01392
R1822 VSS.n111 VSS 9.01392
R1823 VSS.n110 VSS.n109 9.01392
R1824 VSS.n248 VSS.n247 9.01392
R1825 VSS.n247 VSS.n246 9.01392
R1826 VSS.n175 VSS.n174 9.01392
R1827 VSS.n174 VSS.n173 9.01392
R1828 VSS.n169 VSS.n168 9.01392
R1829 VSS.n168 VSS.n167 9.01392
R1830 VSS.n5037 VSS.n5036 9.01392
R1831 VSS.n5036 VSS.n5035 9.01392
R1832 VSS.n5043 VSS.n5041 9.01392
R1833 VSS.n5041 VSS.n5040 9.01392
R1834 VSS.n5051 VSS.n5050 9.01392
R1835 VSS.n5050 VSS.n5049 9.01392
R1836 VSS.n5057 VSS.n5055 9.01392
R1837 VSS.n5055 VSS.n5054 9.01392
R1838 VSS.n5030 VSS.n5029 9.01392
R1839 VSS.n5029 VSS.n5028 9.01392
R1840 VSS.n127 VSS.n126 9.01392
R1841 VSS.n201 VSS.n200 9.01392
R1842 VSS.n200 VSS.n199 9.01392
R1843 VSS.n207 VSS.n206 9.01392
R1844 VSS.n206 VSS.n205 9.01392
R1845 VSS.n155 VSS.n154 9.01392
R1846 VSS.n154 VSS.n153 9.01392
R1847 VSS.n286 VSS.n285 9.01392
R1848 VSS.n285 VSS.n284 9.01392
R1849 VSS.n320 VSS.n319 9.01392
R1850 VSS.n321 VSS.n320 9.01392
R1851 VSS.n326 VSS.n280 9.01392
R1852 VSS VSS.n280 9.01392
R1853 VSS.n363 VSS.n362 9.01392
R1854 VSS.n362 VSS.n361 9.01392
R1855 VSS.n376 VSS.n375 9.01392
R1856 VSS.n375 VSS.n374 9.01392
R1857 VSS.n372 VSS.n371 9.01392
R1858 VSS.n371 VSS.n370 9.01392
R1859 VSS.n392 VSS.n391 9.01392
R1860 VSS.n391 VSS.n390 9.01392
R1861 VSS.n397 VSS.n395 9.01392
R1862 VSS.n395 VSS.n394 9.01392
R1863 VSS.n418 VSS.n416 9.01392
R1864 VSS.n416 VSS.n415 9.01392
R1865 VSS.n412 VSS.n411 9.01392
R1866 VSS.n411 VSS.n410 9.01392
R1867 VSS.n408 VSS.n407 9.01392
R1868 VSS.n407 VSS.n406 9.01392
R1869 VSS.n402 VSS.n401 9.01392
R1870 VSS.n401 VSS.n400 9.01392
R1871 VSS.n4963 VSS.n4962 9.01392
R1872 VSS.n4962 VSS.n4961 9.01392
R1873 VSS.n4969 VSS.n4968 9.01392
R1874 VSS.n4968 VSS.n4967 9.01392
R1875 VSS.n4859 VSS.n4858 9.01392
R1876 VSS.n4858 VSS.n4857 9.01392
R1877 VSS.n4875 VSS.n4874 9.01392
R1878 VSS.n4874 VSS.n4873 9.01392
R1879 VSS.n4919 VSS.n4918 9.01392
R1880 VSS.n4916 VSS.n4915 9.01392
R1881 VSS.n4915 VSS.n4914 9.01392
R1882 VSS.n4894 VSS.n4892 9.01392
R1883 VSS.n4892 VSS.n4891 9.01392
R1884 VSS.n4886 VSS.n4885 9.01392
R1885 VSS.n2908 VSS.n2907 9.01392
R1886 VSS.n2907 VSS.n2906 9.01392
R1887 VSS.n2903 VSS.n2902 9.01392
R1888 VSS.n2902 VSS.n2901 9.01392
R1889 VSS.n2932 VSS.n2931 9.01392
R1890 VSS.n2931 VSS.n2930 9.01392
R1891 VSS.n2948 VSS.n2947 9.01392
R1892 VSS.n2947 VSS.n2946 9.01392
R1893 VSS.n2979 VSS.n2978 9.01392
R1894 VSS.n2978 VSS.n2977 9.01392
R1895 VSS.n2993 VSS.n2992 9.01392
R1896 VSS.n2992 VSS.n2991 9.01392
R1897 VSS.n2998 VSS.n2997 9.01392
R1898 VSS.n2997 VSS.n2996 9.01392
R1899 VSS.n3025 VSS.n3024 9.01392
R1900 VSS.n3024 VSS.n3023 9.01392
R1901 VSS.n3029 VSS.n3028 9.01392
R1902 VSS.n3028 VSS.n3027 9.01392
R1903 VSS.n3045 VSS.n3044 9.01392
R1904 VSS.n3044 VSS.n3043 9.01392
R1905 VSS.n3066 VSS.n3065 9.01392
R1906 VSS.n3065 VSS.n3064 9.01392
R1907 VSS.n3062 VSS.n3061 9.01392
R1908 VSS.n3061 VSS.n3060 9.01392
R1909 VSS.n3054 VSS.n3053 9.01392
R1910 VSS.n3093 VSS.n3092 9.01392
R1911 VSS.n3092 VSS.n3091 9.01392
R1912 VSS.n3105 VSS.n3104 9.01392
R1913 VSS.n3104 VSS.n3103 9.01392
R1914 VSS.n3097 VSS.n3096 9.01392
R1915 VSS.n3136 VSS.n3135 9.01392
R1916 VSS.n3137 VSS.n3136 9.01392
R1917 VSS.n3140 VSS.n3139 9.01392
R1918 VSS.n3139 VSS 9.01392
R1919 VSS.n3138 VSS.n3116 9.01392
R1920 VSS.n3155 VSS.n3153 9.01392
R1921 VSS.n3153 VSS.n3152 9.01392
R1922 VSS.n3147 VSS.n3146 9.01392
R1923 VSS.n3170 VSS.n3169 9.01392
R1924 VSS.n3169 VSS.n3168 9.01392
R1925 VSS.n3177 VSS.n3175 9.01392
R1926 VSS.n3175 VSS.n3174 9.01392
R1927 VSS.n4530 VSS.n4529 9.01392
R1928 VSS.n4529 VSS.n4528 9.01392
R1929 VSS.n4535 VSS.n4534 9.01392
R1930 VSS.n4534 VSS.n4533 9.01392
R1931 VSS.n4357 VSS.n4356 9.01392
R1932 VSS.n4356 VSS.n4355 9.01392
R1933 VSS.n4365 VSS.n4364 9.01392
R1934 VSS.n4364 VSS.n4363 9.01392
R1935 VSS.n4331 VSS.n4329 9.01392
R1936 VSS.n4329 VSS.n4328 9.01392
R1937 VSS.n4325 VSS.n4324 9.01392
R1938 VSS.n4324 VSS.n4323 9.01392
R1939 VSS.n4164 VSS.n4162 9.01392
R1940 VSS.n4162 VSS.n4161 9.01392
R1941 VSS.n4169 VSS.n4168 9.01392
R1942 VSS.n4168 VSS.n4167 9.01392
R1943 VSS.n4173 VSS.n4172 9.01392
R1944 VSS.n4172 VSS.n4171 9.01392
R1945 VSS.n4183 VSS.n4182 9.01392
R1946 VSS.n4182 VSS.n4181 9.01392
R1947 VSS.n4178 VSS.n4177 9.01392
R1948 VSS.n4177 VSS.n4176 9.01392
R1949 VSS.n4201 VSS.n4200 9.01392
R1950 VSS.n4200 VSS.n4199 9.01392
R1951 VSS.n4207 VSS.n4206 9.01392
R1952 VSS.n4206 VSS.n4205 9.01392
R1953 VSS.n4142 VSS.n4141 9.01392
R1954 VSS.n4141 VSS.n4140 9.01392
R1955 VSS.n4147 VSS.n4146 9.01392
R1956 VSS.n4146 VSS.n4145 9.01392
R1957 VSS.n4151 VSS.n4150 9.01392
R1958 VSS.n4150 VSS.n4149 9.01392
R1959 VSS.n4243 VSS.n4242 9.01392
R1960 VSS.n4242 VSS.n4241 9.01392
R1961 VSS.n4246 VSS.n4245 9.01392
R1962 VSS.n4253 VSS.n4252 9.01392
R1963 VSS.n4254 VSS.n4253 9.01392
R1964 VSS.n4238 VSS.n4237 9.01392
R1965 VSS.n4320 VSS.n4319 9.01392
R1966 VSS.n4319 VSS.n4318 9.01392
R1967 VSS.n4432 VSS.n4431 9.01392
R1968 VSS.n4431 VSS.n4430 9.01392
R1969 VSS.n4425 VSS.n4424 9.01392
R1970 VSS.n4421 VSS.n4419 9.01392
R1971 VSS.n4419 VSS.n4418 9.01392
R1972 VSS.n4407 VSS.n4375 9.01392
R1973 VSS.n4409 VSS.n4408 9.01392
R1974 VSS.n4408 VSS 9.01392
R1975 VSS.n4405 VSS.n4404 9.01392
R1976 VSS.n4406 VSS.n4405 9.01392
R1977 VSS.n4394 VSS.n4393 9.01392
R1978 VSS.n4384 VSS.n4383 9.01392
R1979 VSS.n4383 VSS.n4382 9.01392
R1980 VSS.n4378 VSS.n4377 9.01392
R1981 VSS.n4377 VSS.n4376 9.01392
R1982 VSS.n3249 VSS.n3248 9.01392
R1983 VSS.n3244 VSS.n3243 9.01392
R1984 VSS.n3243 VSS.n3242 9.01392
R1985 VSS.n4479 VSS.n4478 9.01392
R1986 VSS.n4478 VSS.n4477 9.01392
R1987 VSS.n4473 VSS.n4472 9.01392
R1988 VSS.n4472 VSS.n4471 9.01392
R1989 VSS.n3221 VSS.n3220 9.01392
R1990 VSS.n3220 VSS.n3219 9.01392
R1991 VSS.n3228 VSS.n3226 9.01392
R1992 VSS.n3226 VSS.n3225 9.01392
R1993 VSS.n3216 VSS.n3215 9.01392
R1994 VSS.n3215 VSS.n3214 9.01392
R1995 VSS.n3204 VSS.n3202 9.01392
R1996 VSS.n3202 VSS.n3201 9.01392
R1997 VSS.n3197 VSS.n3196 9.01392
R1998 VSS.n3196 VSS.n3195 9.01392
R1999 VSS.n4507 VSS.n4506 9.01392
R2000 VSS.n4506 VSS.n4505 9.01392
R2001 VSS.n4501 VSS.n4499 9.01392
R2002 VSS.n4499 VSS.n4498 9.01392
R2003 VSS.n4547 VSS.n4546 9.01392
R2004 VSS.n4546 VSS.n4545 9.01392
R2005 VSS.n4541 VSS.n4540 9.01392
R2006 VSS.n4540 VSS.n4539 9.01392
R2007 VSS.n4436 VSS.n4435 9.01392
R2008 VSS.n4435 VSS.n4434 9.01392
R2009 VSS.n4522 VSS.n4521 9.01392
R2010 VSS.n4521 VSS.n4520 9.01392
R2011 VSS.n3004 VSS.n3003 9.01392
R2012 VSS.n3003 VSS.n3002 9.01392
R2013 VSS.n2954 VSS.n2953 9.01392
R2014 VSS.n2953 VSS.n2952 9.01392
R2015 VSS.n2973 VSS.n2972 9.01392
R2016 VSS.n2972 VSS.n2971 9.01392
R2017 VSS.n2924 VSS.n2923 9.01392
R2018 VSS.n2923 VSS.n2922 9.01392
R2019 VSS.n2898 VSS.n2897 9.01392
R2020 VSS.n2897 VSS.n2896 9.01392
R2021 VSS.n4909 VSS.n4878 9.01392
R2022 VSS VSS.n4878 9.01392
R2023 VSS.n4913 VSS.n4912 9.01392
R2024 VSS.n4931 VSS.n4930 9.01392
R2025 VSS.n4930 VSS.n4929 9.01392
R2026 VSS.n4938 VSS.n4937 9.01392
R2027 VSS.n4927 VSS.n4926 9.01392
R2028 VSS.n4926 VSS.n4925 9.01392
R2029 VSS.n4853 VSS.n4852 9.01392
R2030 VSS.n4852 VSS.n4851 9.01392
R2031 VSS.n345 VSS.n344 9.01392
R2032 VSS.n344 VSS.n343 9.01392
R2033 VSS.n340 VSS.n339 9.01392
R2034 VSS.n339 VSS.n338 9.01392
R2035 VSS.n5003 VSS.n5002 9.01392
R2036 VSS.n5010 VSS.n5009 9.01392
R2037 VSS.n5009 VSS.n5008 9.01392
R2038 VSS.n323 VSS.n322 9.01392
R2039 VSS.n349 VSS.n348 9.01392
R2040 VSS.n348 VSS.n347 9.01392
R2041 VSS.n303 VSS.n302 9.01392
R2042 VSS.n302 VSS.n301 9.01392
R2043 VSS.n297 VSS.n296 9.01392
R2044 VSS.n296 VSS.n295 9.01392
R2045 VSS.n290 VSS.n289 9.01392
R2046 VSS.n313 VSS.n312 9.01392
R2047 VSS.n149 VSS.n148 9.01392
R2048 VSS.n148 VSS.n147 9.01392
R2049 VSS.n229 VSS.n228 9.01392
R2050 VSS.n228 VSS.n227 9.01392
R2051 VSS.n224 VSS.n223 9.01392
R2052 VSS.n223 VSS.n222 9.01392
R2053 VSS.n233 VSS.n232 9.01392
R2054 VSS.n232 VSS.n231 9.01392
R2055 VSS.n124 VSS.n123 9.01392
R2056 VSS.n123 VSS.n122 9.01392
R2057 VSS.n255 VSS.n254 9.01392
R2058 VSS.n254 VSS.n253 9.01392
R2059 VSS.n103 VSS.n102 9.01392
R2060 VSS.n104 VSS.n103 9.01392
R2061 VSS.n70 VSS.n69 9.01392
R2062 VSS.n63 VSS.n62 9.01392
R2063 VSS.n62 VSS.n61 9.01392
R2064 VSS.n59 VSS.n58 9.01392
R2065 VSS.n58 VSS.n57 9.01392
R2066 VSS.n78 VSS.n77 9.01392
R2067 VSS.n77 VSS.n76 9.01392
R2068 VSS.n20 VSS.n19 9.01392
R2069 VSS.n19 VSS.n18 9.01392
R2070 VSS.n2025 VSS.n2024 9.01392
R2071 VSS.n2024 VSS.n2023 9.01392
R2072 VSS.n1540 VSS.n1539 9.01392
R2073 VSS.n1539 VSS.n1538 9.01392
R2074 VSS.n1543 VSS.n1542 9.01392
R2075 VSS.n1535 VSS.n1534 9.01392
R2076 VSS.n1534 VSS.n1533 9.01392
R2077 VSS.n1522 VSS.n1521 9.01392
R2078 VSS VSS.n1522 9.01392
R2079 VSS.n1502 VSS.n1501 9.01392
R2080 VSS.n1501 VSS.n1500 9.01392
R2081 VSS.n1480 VSS.n1479 9.01392
R2082 VSS.n1479 VSS.n1478 9.01392
R2083 VSS.n1448 VSS.n1447 9.01392
R2084 VSS.n1447 VSS.n1446 9.01392
R2085 VSS.n1589 VSS.n1588 9.01392
R2086 VSS.n1588 VSS.n1587 9.01392
R2087 VSS.n1277 VSS.n1276 9.01392
R2088 VSS.n1276 VSS.n1275 9.01392
R2089 VSS.n1181 VSS.n1180 9.01392
R2090 VSS.n1180 VSS.n1179 9.01392
R2091 VSS.n1023 VSS.n1022 9.01392
R2092 VSS.n1021 VSS.n1020 9.01392
R2093 VSS VSS.n1021 9.01392
R2094 VSS.n995 VSS.n994 9.01392
R2095 VSS.n1001 VSS.n1000 9.01392
R2096 VSS.n1000 VSS.n999 9.01392
R2097 VSS.n1101 VSS.n1100 9.01392
R2098 VSS.n1100 VSS.n1099 9.01392
R2099 VSS.n1104 VSS.n1103 9.01392
R2100 VSS.n1117 VSS.n1116 9.01392
R2101 VSS.n1116 VSS.n1115 9.01392
R2102 VSS.n1112 VSS.n1111 9.01392
R2103 VSS.n1111 VSS.n1110 9.01392
R2104 VSS.n1300 VSS.n1299 9.01392
R2105 VSS.n1299 VSS.n1298 9.01392
R2106 VSS.n1407 VSS.n1406 9.01392
R2107 VSS.n1400 VSS.n1399 9.01392
R2108 VSS.n1399 VSS.n1398 9.01392
R2109 VSS.n1396 VSS.n1395 9.01392
R2110 VSS.n1395 VSS.n1394 9.01392
R2111 VSS.n1387 VSS.n1386 9.01392
R2112 VSS.n1386 VSS.n1385 9.01392
R2113 VSS.n1383 VSS.n1382 9.01392
R2114 VSS.n1382 VSS.n1381 9.01392
R2115 VSS.n1375 VSS.n1374 9.01392
R2116 VSS.n1374 VSS.n1373 9.01392
R2117 VSS.n1369 VSS.n1368 9.01392
R2118 VSS.n1368 VSS.n1367 9.01392
R2119 VSS.n1361 VSS.n1360 9.01392
R2120 VSS.n1360 VSS.n1359 9.01392
R2121 VSS.n1306 VSS.n1305 9.01392
R2122 VSS.n1349 VSS.n1348 9.01392
R2123 VSS.n1311 VSS.n1310 9.01392
R2124 VSS VSS.n1311 9.01392
R2125 VSS.n1339 VSS.n1338 9.01392
R2126 VSS.n1335 VSS.n1334 9.01392
R2127 VSS.n1334 VSS.n1333 9.01392
R2128 VSS.n1320 VSS.n1319 9.01392
R2129 VSS.n1319 VSS.n1318 9.01392
R2130 VSS.n1875 VSS.n1874 9.01392
R2131 VSS.n1874 VSS.n1873 9.01392
R2132 VSS.n1885 VSS.n1884 9.01392
R2133 VSS.n1884 VSS.n1883 9.01392
R2134 VSS.n859 VSS.n858 9.01392
R2135 VSS.n858 VSS.n857 9.01392
R2136 VSS.n852 VSS.n851 9.01392
R2137 VSS.n851 VSS.n850 9.01392
R2138 VSS.n844 VSS.n843 9.01392
R2139 VSS.n843 VSS.n842 9.01392
R2140 VSS.n881 VSS.n880 9.01392
R2141 VSS.n880 VSS.n879 9.01392
R2142 VSS.n875 VSS.n874 9.01392
R2143 VSS.n874 VSS.n873 9.01392
R2144 VSS.n824 VSS.n823 9.01392
R2145 VSS.n823 VSS.n822 9.01392
R2146 VSS.n818 VSS.n815 9.01392
R2147 VSS.n815 VSS.n814 9.01392
R2148 VSS.n802 VSS.n800 9.01392
R2149 VSS.n800 VSS.n799 9.01392
R2150 VSS.n795 VSS.n794 9.01392
R2151 VSS.n794 VSS.n793 9.01392
R2152 VSS.n2480 VSS.n2479 9.01392
R2153 VSS.n2479 VSS.n2478 9.01392
R2154 VSS.n2486 VSS.n2485 9.01392
R2155 VSS.n2485 VSS.n2484 9.01392
R2156 VSS.n2494 VSS.n2493 9.01392
R2157 VSS.n2493 VSS.n2492 9.01392
R2158 VSS.n2498 VSS.n2497 9.01392
R2159 VSS.n2497 VSS.n2496 9.01392
R2160 VSS.n2476 VSS.n2475 9.01392
R2161 VSS.n2475 VSS.n2474 9.01392
R2162 VSS.n2471 VSS.n2468 9.01392
R2163 VSS.n2468 VSS.n2467 9.01392
R2164 VSS.n2464 VSS.n2462 9.01392
R2165 VSS.n2462 VSS.n2461 9.01392
R2166 VSS.n772 VSS.n771 9.01392
R2167 VSS.n771 VSS.n770 9.01392
R2168 VSS.n668 VSS.n667 9.01392
R2169 VSS.n767 VSS.n665 9.01392
R2170 VSS VSS.n665 9.01392
R2171 VSS.n766 VSS.n670 9.01392
R2172 VSS.n670 VSS.n669 9.01392
R2173 VSS.n672 VSS.n671 9.01392
R2174 VSS.n762 VSS.n761 9.01392
R2175 VSS.n761 VSS.n760 9.01392
R2176 VSS.n758 VSS.n757 9.01392
R2177 VSS.n757 VSS.n756 9.01392
R2178 VSS.n677 VSS.n676 9.01392
R2179 VSS.n753 VSS.n752 9.01392
R2180 VSS.n752 VSS.n751 9.01392
R2181 VSS.n749 VSS.n748 9.01392
R2182 VSS.n748 VSS.n747 9.01392
R2183 VSS.n745 VSS.n744 9.01392
R2184 VSS.n744 VSS.n743 9.01392
R2185 VSS.n741 VSS.n740 9.01392
R2186 VSS.n740 VSS.n739 9.01392
R2187 VSS.n737 VSS.n734 9.01392
R2188 VSS.n734 VSS.n733 9.01392
R2189 VSS.n731 VSS.n730 9.01392
R2190 VSS.n730 VSS.n729 9.01392
R2191 VSS.n727 VSS.n726 9.01392
R2192 VSS.n726 VSS.n725 9.01392
R2193 VSS.n723 VSS.n722 9.01392
R2194 VSS.n722 VSS.n721 9.01392
R2195 VSS.n719 VSS.n718 9.01392
R2196 VSS.n718 VSS.n717 9.01392
R2197 VSS.n715 VSS.n714 9.01392
R2198 VSS.n714 VSS.n713 9.01392
R2199 VSS.n710 VSS.n709 9.01392
R2200 VSS.n709 VSS.n708 9.01392
R2201 VSS.n705 VSS.n704 9.01392
R2202 VSS.n704 VSS.n703 9.01392
R2203 VSS.n4825 VSS.n479 9.01392
R2204 VSS VSS.n479 9.01392
R2205 VSS.n4819 VSS.n4818 9.01392
R2206 VSS.n4812 VSS.n4811 9.01392
R2207 VSS.n4811 VSS.n4810 9.01392
R2208 VSS.n484 VSS.n483 9.01392
R2209 VSS.n4794 VSS.n4793 9.01392
R2210 VSS.n4793 VSS.n4792 9.01392
R2211 VSS.n4623 VSS.n4622 9.01392
R2212 VSS.n4601 VSS.n4600 9.01392
R2213 VSS VSS.n4600 9.01392
R2214 VSS.n4620 VSS.n4619 9.01392
R2215 VSS.n4621 VSS.n4620 9.01392
R2216 VSS.n4604 VSS.n4603 9.01392
R2217 VSS.n4579 VSS.n4578 9.01392
R2218 VSS.n4578 VSS.n4577 9.01392
R2219 VSS.n4572 VSS.n4571 9.01392
R2220 VSS.n3997 VSS.n3996 9.01392
R2221 VSS.n3996 VSS.n3995 9.01392
R2222 VSS.n4010 VSS.n4009 9.01392
R2223 VSS.n4009 VSS.n4008 9.01392
R2224 VSS.n4014 VSS.n4013 9.01392
R2225 VSS.n4013 VSS.n4012 9.01392
R2226 VSS.n4020 VSS.n4017 9.01392
R2227 VSS.n4017 VSS.n4016 9.01392
R2228 VSS.n4024 VSS.n4023 9.01392
R2229 VSS.n4023 VSS.n4022 9.01392
R2230 VSS.n4028 VSS.n4027 9.01392
R2231 VSS.n4027 VSS.n4026 9.01392
R2232 VSS.n4032 VSS.n4031 9.01392
R2233 VSS.n4031 VSS.n4030 9.01392
R2234 VSS.n4036 VSS.n4035 9.01392
R2235 VSS.n4035 VSS.n4034 9.01392
R2236 VSS.n4041 VSS.n4040 9.01392
R2237 VSS.n4040 VSS.n4039 9.01392
R2238 VSS.n4045 VSS.n4044 9.01392
R2239 VSS.n4044 VSS.n4043 9.01392
R2240 VSS.n4049 VSS.n4048 9.01392
R2241 VSS.n4048 VSS.n4047 9.01392
R2242 VSS.n4053 VSS.n4052 9.01392
R2243 VSS.n4052 VSS.n4051 9.01392
R2244 VSS.n4059 VSS.n4058 9.01392
R2245 VSS.n4058 VSS.n4057 9.01392
R2246 VSS.n4063 VSS.n4062 9.01392
R2247 VSS.n4062 VSS.n4061 9.01392
R2248 VSS.n4067 VSS.n4066 9.01392
R2249 VSS.n4066 VSS.n4065 9.01392
R2250 VSS.n4071 VSS.n4070 9.01392
R2251 VSS.n4070 VSS.n4069 9.01392
R2252 VSS.n4074 VSS.n4073 9.01392
R2253 VSS.n4080 VSS.n4079 9.01392
R2254 VSS.n4079 VSS.n4078 9.01392
R2255 VSS.n4083 VSS.n4082 9.01392
R2256 VSS.n4090 VSS.n4089 9.01392
R2257 VSS VSS.n4090 9.01392
R2258 VSS.n4093 VSS.n4092 9.01392
R2259 VSS.n4092 VSS.n4091 9.01392
R2260 VSS.n3985 VSS.n3984 9.01392
R2261 VSS.n3948 VSS.n3947 9.01392
R2262 VSS.n3947 VSS.n3946 9.01392
R2263 VSS.n3951 VSS.n3950 9.01392
R2264 VSS.n3966 VSS.n3965 9.01392
R2265 VSS.n3965 VSS.n3964 9.01392
R2266 VSS.n4106 VSS.n4105 9.01392
R2267 VSS.n4105 VSS.n4104 9.01392
R2268 VSS.n4139 VSS.n4138 9.01392
R2269 VSS.n4262 VSS.n4261 9.01392
R2270 VSS.n4261 VSS.n4260 9.01392
R2271 VSS.n4132 VSS.n4131 9.01392
R2272 VSS.n4267 VSS.n4266 9.01392
R2273 VSS.n4266 VSS.n4265 9.01392
R2274 VSS.n4271 VSS.n4270 9.01392
R2275 VSS.n4270 VSS.n4269 9.01392
R2276 VSS.n4275 VSS.n4274 9.01392
R2277 VSS.n4274 VSS.n4273 9.01392
R2278 VSS.n4281 VSS.n4280 9.01392
R2279 VSS.n4280 VSS.n4279 9.01392
R2280 VSS.n4285 VSS.n4284 9.01392
R2281 VSS.n4284 VSS.n4283 9.01392
R2282 VSS.n4289 VSS.n4288 9.01392
R2283 VSS.n4288 VSS.n4287 9.01392
R2284 VSS.n4293 VSS.n4292 9.01392
R2285 VSS.n4292 VSS.n4291 9.01392
R2286 VSS.n4298 VSS.n4297 9.01392
R2287 VSS.n4297 VSS.n4296 9.01392
R2288 VSS.n4302 VSS.n4301 9.01392
R2289 VSS.n4301 VSS.n4300 9.01392
R2290 VSS.n4127 VSS.n4126 9.01392
R2291 VSS.n4126 VSS.n4125 9.01392
R2292 VSS.n3929 VSS.n3928 9.01392
R2293 VSS.n3928 VSS.n3927 9.01392
R2294 VSS.n3935 VSS.n3933 9.01392
R2295 VSS.n3933 VSS.n3932 9.01392
R2296 VSS.n3924 VSS.n3923 9.01392
R2297 VSS.n3923 VSS.n3922 9.01392
R2298 VSS.n4112 VSS.n4111 9.01392
R2299 VSS.n4111 VSS.n4110 9.01392
R2300 VSS.n4257 VSS.n4256 9.01392
R2301 VSS.n4256 VSS 9.01392
R2302 VSS.n3960 VSS.n3959 9.01392
R2303 VSS.n3959 VSS.n3958 9.01392
R2304 VSS.n3982 VSS.n3981 9.01392
R2305 VSS.n3981 VSS.n3980 9.01392
R2306 VSS.n3993 VSS.n3992 9.01392
R2307 VSS.n3992 VSS.n3991 9.01392
R2308 VSS.n4567 VSS.n4566 9.01392
R2309 VSS.n4566 VSS.n4565 9.01392
R2310 VSS.n4592 VSS.n4591 9.01392
R2311 VSS.n2880 VSS.n2879 9.01392
R2312 VSS.n2879 VSS.n2878 9.01392
R2313 VSS.n2874 VSS.n2873 9.01392
R2314 VSS.n2873 VSS.n2872 9.01392
R2315 VSS.n2868 VSS.n2867 9.01392
R2316 VSS.n2867 VSS.n2866 9.01392
R2317 VSS.n2864 VSS.n2863 9.01392
R2318 VSS.n2863 VSS.n2862 9.01392
R2319 VSS.n2858 VSS.n2857 9.01392
R2320 VSS.n2857 VSS.n2856 9.01392
R2321 VSS.n2854 VSS.n2853 9.01392
R2322 VSS.n2853 VSS.n2852 9.01392
R2323 VSS.n2850 VSS.n2849 9.01392
R2324 VSS.n2849 VSS.n2848 9.01392
R2325 VSS.n2846 VSS.n2845 9.01392
R2326 VSS.n2845 VSS.n2844 9.01392
R2327 VSS.n2841 VSS.n2840 9.01392
R2328 VSS.n2840 VSS.n2839 9.01392
R2329 VSS.n2837 VSS.n2836 9.01392
R2330 VSS.n2836 VSS.n2835 9.01392
R2331 VSS.n2833 VSS.n2832 9.01392
R2332 VSS.n2832 VSS.n2831 9.01392
R2333 VSS.n438 VSS.n437 9.01392
R2334 VSS.n437 VSS.n436 9.01392
R2335 VSS.n444 VSS.n441 9.01392
R2336 VSS.n441 VSS.n440 9.01392
R2337 VSS.n448 VSS.n447 9.01392
R2338 VSS.n447 VSS.n446 9.01392
R2339 VSS.n452 VSS.n451 9.01392
R2340 VSS.n451 VSS.n450 9.01392
R2341 VSS.n456 VSS.n455 9.01392
R2342 VSS.n455 VSS.n454 9.01392
R2343 VSS.n460 VSS.n459 9.01392
R2344 VSS.n459 VSS.n458 9.01392
R2345 VSS.n432 VSS.n431 9.01392
R2346 VSS.n465 VSS.n464 9.01392
R2347 VSS.n464 VSS.n463 9.01392
R2348 VSS.n469 VSS.n468 9.01392
R2349 VSS.n468 VSS.n467 9.01392
R2350 VSS.n472 VSS.n471 9.01392
R2351 VSS.n4630 VSS.n4629 9.01392
R2352 VSS.n4629 VSS.n4628 9.01392
R2353 VSS.n4790 VSS.n4789 9.01392
R2354 VSS.n4789 VSS.n4788 9.01392
R2355 VSS.n4785 VSS.n4784 9.01392
R2356 VSS.n4784 VSS.n4783 9.01392
R2357 VSS.n685 VSS.n684 9.01392
R2358 VSS.n684 VSS.n683 9.01392
R2359 VSS.n701 VSS.n700 9.01392
R2360 VSS.n700 VSS.n699 9.01392
R2361 VSS.n4816 VSS.n4815 9.01392
R2362 VSS.n4817 VSS.n4816 9.01392
R2363 VSS.n661 VSS.n660 9.01392
R2364 VSS.n660 VSS.n659 9.01392
R2365 VSS.n656 VSS.n655 9.01392
R2366 VSS.n655 VSS.n654 9.01392
R2367 VSS.n775 VSS.n774 9.01392
R2368 VSS.n2455 VSS.n2454 9.01392
R2369 VSS.n2454 VSS.n2453 9.01392
R2370 VSS.n2451 VSS.n2450 9.01392
R2371 VSS.n2450 VSS.n2449 9.01392
R2372 VSS.n2447 VSS.n2446 9.01392
R2373 VSS.n2446 VSS.n2445 9.01392
R2374 VSS.n2440 VSS.n2439 9.01392
R2375 VSS.n2437 VSS.n2436 9.01392
R2376 VSS.n2436 VSS.n2435 9.01392
R2377 VSS.n2433 VSS.n2432 9.01392
R2378 VSS.n2432 VSS.n2431 9.01392
R2379 VSS.n2426 VSS.n2425 9.01392
R2380 VSS.n2423 VSS.n2422 9.01392
R2381 VSS.n2422 VSS.n2421 9.01392
R2382 VSS.n2420 VSS.n2419 9.01392
R2383 VSS VSS.n2420 9.01392
R2384 VSS.n2413 VSS.n2412 9.01392
R2385 VSS.n2410 VSS.n2409 9.01392
R2386 VSS.n2409 VSS.n2408 9.01392
R2387 VSS.n2404 VSS.n2403 9.01392
R2388 VSS.n2401 VSS.n2400 9.01392
R2389 VSS.n2400 VSS.n2399 9.01392
R2390 VSS.n2397 VSS.n2396 9.01392
R2391 VSS.n2396 VSS.n2395 9.01392
R2392 VSS.n2393 VSS.n2392 9.01392
R2393 VSS.n2392 VSS.n2391 9.01392
R2394 VSS.n2389 VSS.n2388 9.01392
R2395 VSS.n2388 VSS.n2387 9.01392
R2396 VSS.n2383 VSS.n2382 9.01392
R2397 VSS.n2382 VSS.n2381 9.01392
R2398 VSS.n2379 VSS.n2378 9.01392
R2399 VSS.n2378 VSS.n2377 9.01392
R2400 VSS.n830 VSS.n829 9.01392
R2401 VSS.n829 VSS.n828 9.01392
R2402 VSS.n1932 VSS.n1931 9.01392
R2403 VSS.n1931 VSS.n1930 9.01392
R2404 VSS.n1924 VSS.n1923 9.01392
R2405 VSS.n1923 VSS.n1922 9.01392
R2406 VSS.n1880 VSS.n1879 9.01392
R2407 VSS.n1879 VSS.n1878 9.01392
R2408 VSS.n864 VSS.n863 9.01392
R2409 VSS.n863 VSS.n862 9.01392
R2410 VSS.n1313 VSS.n1312 9.01392
R2411 VSS.n1346 VSS.n1345 9.01392
R2412 VSS.n1347 VSS.n1346 9.01392
R2413 VSS.n1356 VSS.n1355 9.01392
R2414 VSS.n1355 VSS.n1354 9.01392
R2415 VSS.n1365 VSS.n1364 9.01392
R2416 VSS.n1364 VSS.n1363 9.01392
R2417 VSS.n1379 VSS.n1378 9.01392
R2418 VSS.n1378 VSS.n1377 9.01392
R2419 VSS.n1392 VSS.n1391 9.01392
R2420 VSS.n1391 VSS.n1390 9.01392
R2421 VSS.n1404 VSS.n1403 9.01392
R2422 VSS.n1403 VSS.n1402 9.01392
R2423 VSS.n1247 VSS.n1246 9.01392
R2424 VSS.n1246 VSS.n1245 9.01392
R2425 VSS.n1251 VSS.n1250 9.01392
R2426 VSS.n1250 VSS.n1249 9.01392
R2427 VSS.n2156 VSS.n2155 8.84709
R2428 VSS.n2652 VSS.n2651 8.84709
R2429 VSS.n689 VSS.n688 8.82809
R2430 VSS.n2530 VSS.n2529 8.82809
R2431 VSS.n2539 VSS.n2538 8.82809
R2432 VSS.n2544 VSS.n2543 8.82809
R2433 VSS.n2564 VSS.n2563 8.82809
R2434 VSS.n2710 VSS.n2709 8.82809
R2435 VSS.n2744 VSS.n2743 8.82809
R2436 VSS.n4744 VSS.n2777 8.82809
R2437 VSS.n3316 VSS.n3315 8.82809
R2438 VSS.n4410 VSS 8.82809
R2439 VSS.n3141 VSS 8.82809
R2440 VSS.n4911 VSS 8.82809
R2441 VSS VSS.n324 8.82809
R2442 VSS.n108 VSS 8.82809
R2443 VSS.n2226 VSS.n2086 8.6074
R2444 VSS.n2581 VSS.n584 8.6074
R2445 VSS.n3890 VSS.n3889 8.38671
R2446 VSS.n3725 VSS.n3724 8.38671
R2447 VSS.n3873 VSS.n3865 8.38671
R2448 VSS.n3810 VSS.n3794 8.38671
R2449 VSS.n3754 VSS.n3753 8.38671
R2450 VSS.n3779 VSS.n3778 8.38671
R2451 VSS.n4661 VSS.n2821 8.38671
R2452 VSS.n367 VSS.n366 7.72464
R2453 VSS.n894 VSS.n893 7.61156
R2454 VSS.n3307 VSS.n3304 7.50395
R2455 VSS.n3382 VSS.n3379 7.50395
R2456 VSS.n2247 VSS.n2246 7.4558
R2457 VSS.n1757 VSS.n1756 7.4558
R2458 VSS.n1793 VSS.n1791 7.01424
R2459 VSS.n3275 VSS.n3274 6.62119
R2460 VSS.n3517 VSS.n3514 6.62119
R2461 VSS.n3533 VSS.n3530 6.62119
R2462 VSS.n555 VSS.n552 6.62119
R2463 VSS.n539 VSS.n536 6.62119
R2464 VSS.n2770 VSS.n2769 6.4005
R2465 VSS.n3761 VSS.n3760 5.95912
R2466 VSS.n1710 VSS 5.81868
R2467 VSS.n2295 VSS 5.81868
R2468 VSS.n3684 VSS 5.81868
R2469 VSS.n3899 VSS 5.81868
R2470 VSS.n3837 VSS 5.81868
R2471 VSS.n3764 VSS 5.81868
R2472 VSS.n1146 VSS 5.81868
R2473 VSS.n1846 VSS 5.81868
R2474 VSS.n2180 VSS 5.81868
R2475 VSS.n2534 VSS 5.81868
R2476 VSS.n2616 VSS 5.81868
R2477 VSS.n2739 VSS 5.81868
R2478 VSS.n4720 VSS 5.81868
R2479 VSS.n2792 VSS 5.81868
R2480 VSS.n1057 VSS.n1056 5.79462
R2481 VSS.n1054 VSS.n1053 5.79462
R2482 VSS.n1080 VSS.n1079 5.79462
R2483 VSS.n1135 VSS.n1134 5.79462
R2484 VSS.n1151 VSS.n1150 5.79462
R2485 VSS.n1205 VSS.n1204 5.79462
R2486 VSS.n966 VSS.n965 5.79462
R2487 VSS.n1643 VSS.n1642 5.79462
R2488 VSS.n2232 VSS.n2080 5.79462
R2489 VSS.n2227 VSS.n2085 5.79462
R2490 VSS.n2217 VSS.n2213 5.79462
R2491 VSS.n2203 VSS.n2199 5.79462
R2492 VSS.n2189 VSS.n2185 5.79462
R2493 VSS.n2172 VSS.n2168 5.79462
R2494 VSS.n2135 VSS.n2131 5.79462
R2495 VSS.n2121 VSS.n2117 5.79462
R2496 VSS.n2572 VSS.n589 5.79462
R2497 VSS.n2579 VSS.n587 5.79462
R2498 VSS.n2594 VSS.n2590 5.79462
R2499 VSS.n2608 VSS.n2604 5.79462
R2500 VSS.n2625 VSS.n2621 5.79462
R2501 VSS.n2639 VSS.n2635 5.79462
R2502 VSS.n2666 VSS.n2662 5.79462
R2503 VSS.n2686 VSS.n2682 5.79462
R2504 VSS.n3604 VSS.n3601 5.73843
R2505 VSS.n3397 VSS.n3394 5.73843
R2506 VSS.n1793 VSS.n947 5.51774
R2507 VSS.n3626 VSS.n3625 5.51774
R2508 VSS.n2155 VSS.n2154 5.51232
R2509 VSS.n2651 VSS.n2650 5.51232
R2510 VSS.n3903 VSS.n3897 5.29705
R2511 VSS.n1072 VSS.n1052 5.29705
R2512 VSS.n627 VSS.n626 5.29705
R2513 VSS.n2751 VSS.n2750 5.29705
R2514 VSS.n3867 VSS.n3866 5.07636
R2515 VSS.n4655 VSS.n4654 5.07636
R2516 VSS.n900 VSS.n892 5.07636
R2517 VSS.n1230 VSS.n1222 4.85567
R2518 VSS.n2138 VSS.n2137 4.6505
R2519 VSS.n1840 VSS.n1839 4.6505
R2520 VSS.n1826 VSS.n1825 4.6505
R2521 VSS.n939 VSS.n938 4.6505
R2522 VSS.n1778 VSS.n1777 4.6505
R2523 VSS.n1773 VSS.n1772 4.6505
R2524 VSS.n1750 VSS.n1749 4.6505
R2525 VSS.n1736 VSS.n1735 4.6505
R2526 VSS.n1722 VSS.n1721 4.6505
R2527 VSS.n1706 VSS.n1705 4.6505
R2528 VSS.n1679 VSS.n1678 4.6505
R2529 VSS.n1665 VSS.n1664 4.6505
R2530 VSS.n2175 VSS.n2174 4.6505
R2531 VSS.n2192 VSS.n2191 4.6505
R2532 VSS.n2206 VSS.n2205 4.6505
R2533 VSS.n2220 VSS.n2219 4.6505
R2534 VSS.n2235 VSS.n2234 4.6505
R2535 VSS.n2260 VSS.n2259 4.6505
R2536 VSS.n2277 VSS.n2276 4.6505
R2537 VSS.n2291 VSS.n2290 4.6505
R2538 VSS.n2307 VSS.n2306 4.6505
R2539 VSS.n2321 VSS.n2320 4.6505
R2540 VSS.n2338 VSS.n2337 4.6505
R2541 VSS.n2361 VSS.n2360 4.6505
R2542 VSS.n973 VSS.n972 4.6505
R2543 VSS.n1212 VSS.n1211 4.6505
R2544 VSS.n1142 VSS.n1141 4.6505
R2545 VSS.n1087 VSS.n1086 4.6505
R2546 VSS.n2000 VSS.n1999 4.6505
R2547 VSS.n4752 VSS.n4751 4.6505
R2548 VSS.n3729 VSS.n3728 4.6505
R2549 VSS.n3726 VSS.n3725 4.6505
R2550 VSS.n3891 VSS.n3890 4.6505
R2551 VSS.n3878 VSS.n3877 4.6505
R2552 VSS.n3874 VSS.n3873 4.6505
R2553 VSS.n3811 VSS.n3810 4.6505
R2554 VSS.n3791 VSS.n3790 4.6505
R2555 VSS.n3789 VSS.n3788 4.6505
R2556 VSS.n3780 VSS.n3779 4.6505
R2557 VSS.n3755 VSS.n3754 4.6505
R2558 VSS.n2824 VSS.n2823 4.6505
R2559 VSS.n4662 VSS.n4661 4.6505
R2560 VSS.n2777 VSS.n2772 4.6505
R2561 VSS.n4754 VSS.n4753 4.6505
R2562 VSS.n2745 VSS.n2744 4.6505
R2563 VSS.n2736 VSS.n2735 4.6505
R2564 VSS.n2711 VSS.n2710 4.6505
R2565 VSS.n2689 VSS.n2688 4.6505
R2566 VSS.n2669 VSS.n2668 4.6505
R2567 VSS.n2642 VSS.n2641 4.6505
R2568 VSS.n2628 VSS.n2627 4.6505
R2569 VSS.n2611 VSS.n2610 4.6505
R2570 VSS.n2597 VSS.n2596 4.6505
R2571 VSS.n2569 VSS.n2568 4.6505
R2572 VSS.n2565 VSS.n2564 4.6505
R2573 VSS.n2556 VSS.n2548 4.6505
R2574 VSS.n2547 VSS.n2546 4.6505
R2575 VSS.n2545 VSS.n2544 4.6505
R2576 VSS.n2540 VSS.n2539 4.6505
R2577 VSS.n599 VSS.n598 4.6505
R2578 VSS.n630 VSS.n629 4.6505
R2579 VSS.n2124 VSS.n2123 4.6505
R2580 VSS.n3479 VSS.n3436 4.6505
R2581 VSS.n3414 VSS.n3413 4.6505
R2582 VSS.n562 VSS.n561 4.6505
R2583 VSS.n3313 VSS.n3312 4.6505
R2584 VSS.n3336 VSS.n3335 4.6505
R2585 VSS.n3547 VSS.n3546 4.6505
R2586 VSS.n2803 VSS.n2802 4.6505
R2587 VSS.n2816 VSS.n2815 4.6505
R2588 VSS.n1435 VSS.n1434 4.6505
R2589 VSS.n170 VSS.n169 4.6505
R2590 VSS.n5044 VSS.n5043 4.6505
R2591 VSS.n5058 VSS.n5057 4.6505
R2592 VSS.n2949 VSS.n2948 4.6505
R2593 VSS.n4202 VSS.n4201 4.6505
R2594 VSS.n4332 VSS.n4331 4.6505
R2595 VSS.n4358 VSS.n4357 4.6505
R2596 VSS.n4422 VSS.n4421 4.6505
R2597 VSS.n4385 VSS.n4384 4.6505
R2598 VSS.n3245 VSS.n3244 4.6505
R2599 VSS.n4474 VSS.n4473 4.6505
R2600 VSS.n3229 VSS.n3228 4.6505
R2601 VSS.n3205 VSS.n3204 4.6505
R2602 VSS.n4542 VSS.n4541 4.6505
R2603 VSS.n3178 VSS.n3177 4.6505
R2604 VSS.n3156 VSS.n3155 4.6505
R2605 VSS.n3135 VSS.n3134 4.6505
R2606 VSS.n3046 VSS.n3045 4.6505
R2607 VSS.n3005 VSS.n3004 4.6505
R2608 VSS.n2974 VSS.n2973 4.6505
R2609 VSS.n2925 VSS.n2924 4.6505
R2610 VSS.n4895 VSS.n4894 4.6505
R2611 VSS.n4909 VSS.n4908 4.6505
R2612 VSS.n4964 VSS.n4963 4.6505
R2613 VSS.n419 VSS.n418 4.6505
R2614 VSS.n364 VSS.n363 4.6505
R2615 VSS.n327 VSS.n326 4.6505
R2616 VSS.n304 VSS.n303 4.6505
R2617 VSS.n150 VSS.n149 4.6505
R2618 VSS.n202 VSS.n201 4.6505
R2619 VSS.n256 VSS.n255 4.6505
R2620 VSS.n49 VSS.n48 4.6505
R2621 VSS.n21 VSS.n20 4.6505
R2622 VSS.n2019 VSS.n2018 4.6505
R2623 VSS.n1906 VSS.n1905 4.6505
R2624 VSS.n1596 VSS.n1595 4.6505
R2625 VSS.n1189 VSS.n1188 4.6505
R2626 VSS.n853 VSS.n852 4.6505
R2627 VSS.n876 VSS.n875 4.6505
R2628 VSS.n825 VSS.n824 4.6505
R2629 VSS.n803 VSS.n802 4.6505
R2630 VSS.n2487 VSS.n2486 4.6505
R2631 VSS.n4107 VSS.n4106 4.6505
R2632 VSS.n4128 VSS.n4127 4.6505
R2633 VSS.n3936 VSS.n3935 4.6505
R2634 VSS.n3961 VSS.n3960 4.6505
R2635 VSS.n4568 VSS.n4567 4.6505
R2636 VSS.n2875 VSS.n2874 4.6505
R2637 VSS.n686 VSS.n685 4.6505
R2638 VSS.n4815 VSS.n478 4.6505
R2639 VSS.n2465 VSS.n2464 4.6505
R2640 VSS.n1925 VSS.n1924 4.6505
R2641 VSS.n1336 VSS.n1335 4.6505
R2642 VSS.n1301 VSS.n1300 4.6505
R2643 VSS.n2557 VSS.n2554 4.63498
R2644 VSS.n4750 VSS.n2776 4.63498
R2645 VSS.n2818 VSS.n2817 4.5005
R2646 VSS.n2805 VSS.n2804 4.5005
R2647 VSS.n2771 VSS.n2770 4.5005
R2648 VSS.n2754 VSS.n2753 4.5005
R2649 VSS.n2158 VSS.n2157 4.5005
R2650 VSS.n1795 VSS.n1794 4.5005
R2651 VSS.n1621 VSS.n1620 4.5005
R2652 VSS.n1232 VSS.n1231 4.5005
R2653 VSS.n1165 VSS.n1164 4.5005
R2654 VSS.n1074 VSS.n1073 4.5005
R2655 VSS.n2718 VSS.n2717 4.5005
R2656 VSS.n628 VSS.n627 4.5005
R2657 VSS.n3290 VSS.n3289 4.5005
R2658 VSS.n3904 VSS.n3903 4.5005
R2659 VSS.n3767 VSS.n3766 4.5005
R2660 VSS.n3317 VSS.n3316 4.5005
R2661 VSS.n3338 VSS.n3337 4.5005
R2662 VSS.n3450 VSS.n3449 4.5005
R2663 VSS.n3549 VSS.n3548 4.5005
R2664 VSS.n564 VSS.n563 4.5005
R2665 VSS.n3416 VSS.n3415 4.5005
R2666 VSS.n3481 VSS.n3480 4.5005
R2667 VSS.n4234 VSS.n4233 4.5005
R2668 VSS.n4204 VSS.n4203 4.5005
R2669 VSS.n4334 VSS.n4333 4.5005
R2670 VSS.n3247 VSS.n3246 4.5005
R2671 VSS.n3232 VSS.n3231 4.5005
R2672 VSS.n3133 VSS.n3132 4.5005
R2673 VSS.n3048 VSS.n3047 4.5005
R2674 VSS.n204 VSS.n203 4.5005
R2675 VSS.n25 VSS.n24 4.5005
R2676 VSS.n1908 VSS.n1907 4.5005
R2677 VSS.n2021 VSS.n2020 4.5005
R2678 VSS.n1598 VSS.n1597 4.5005
R2679 VSS.n1191 VSS.n1190 4.5005
R2680 VSS.n98 VSS.n97 4.5005
R2681 VSS.n5060 VSS.n5059 4.5005
R2682 VSS.n5046 VSS.n5045 4.5005
R2683 VSS.n172 VSS.n171 4.5005
R2684 VSS.n152 VSS.n151 4.5005
R2685 VSS.n4856 VSS.n4855 4.5005
R2686 VSS.n4966 VSS.n4965 4.5005
R2687 VSS.n421 VSS.n420 4.5005
R2688 VSS.n368 VSS.n367 4.5005
R2689 VSS.n306 VSS.n305 4.5005
R2690 VSS.n4941 VSS.n4940 4.5005
R2691 VSS.n4884 VSS.n4883 4.5005
R2692 VSS.n4897 VSS.n4896 4.5005
R2693 VSS.n2929 VSS.n2928 4.5005
R2694 VSS.n2951 VSS.n2950 4.5005
R2695 VSS.n2976 VSS.n2975 4.5005
R2696 VSS.n3007 VSS.n3006 4.5005
R2697 VSS.n3180 VSS.n3179 4.5005
R2698 VSS.n3158 VSS.n3157 4.5005
R2699 VSS.n3057 VSS.n3056 4.5005
R2700 VSS.n4417 VSS.n4416 4.5005
R2701 VSS.n4360 VSS.n4359 4.5005
R2702 VSS.n4387 VSS.n4386 4.5005
R2703 VSS.n4476 VSS.n4475 4.5005
R2704 VSS.n3207 VSS.n3206 4.5005
R2705 VSS.n4504 VSS.n4503 4.5005
R2706 VSS.n4544 VSS.n4543 4.5005
R2707 VSS.n329 VSS.n328 4.5005
R2708 VSS.n258 VSS.n257 4.5005
R2709 VSS.n51 VSS.n50 4.5005
R2710 VSS.n1493 VSS.n1492 4.5005
R2711 VSS.n1438 VSS.n1437 4.5005
R2712 VSS.n3938 VSS.n3937 4.5005
R2713 VSS.n4109 VSS.n4108 4.5005
R2714 VSS.n4000 VSS.n3999 4.5005
R2715 VSS.n4570 VSS.n4569 4.5005
R2716 VSS.n805 VSS.n804 4.5005
R2717 VSS.n878 VSS.n877 4.5005
R2718 VSS.n1331 VSS.n1330 4.5005
R2719 VSS.n1927 VSS.n1926 4.5005
R2720 VSS.n849 VSS.n848 4.5005
R2721 VSS.n2460 VSS.n2459 4.5005
R2722 VSS.n2489 VSS.n2488 4.5005
R2723 VSS.n827 VSS.n826 4.5005
R2724 VSS.n690 VSS.n689 4.5005
R2725 VSS.n487 VSS.n486 4.5005
R2726 VSS.n2877 VSS.n2876 4.5005
R2727 VSS.n4598 VSS.n4597 4.5005
R2728 VSS.n3963 VSS.n3962 4.5005
R2729 VSS.n4130 VSS.n4129 4.5005
R2730 VSS.n4827 VSS.n4826 4.5005
R2731 VSS.n1304 VSS.n1303 4.5005
R2732 VSS.n902 VSS.n901 4.49926
R2733 VSS.n1692 VSS.n1691 4.49926
R2734 VSS.n2324 VSS.n2073 4.49926
R2735 VSS.n2655 VSS.n2654 4.49926
R2736 VSS.n2225 VSS.n2223 4.42059
R2737 VSS.n1755 VSS.n1754 4.42059
R2738 VSS.n2263 VSS.n2075 4.42059
R2739 VSS.n2584 VSS.n2583 4.42059
R2740 VSS.n4595 VSS.n4594 4.16651
R2741 VSS.n3577 VSS.n3574 3.97291
R2742 VSS.n3372 VSS.n3369 3.97291
R2743 VSS.n1061 VSS 3.88975
R2744 VSS.n1224 VSS.n1223 3.8312
R2745 VSS.n895 VSS.n894 3.82791
R2746 VSS.n4257 VSS 3.75222
R2747 VSS.n4089 VSS 3.75222
R2748 VSS VSS.n4601 3.75222
R2749 VSS VSS.n4825 3.75222
R2750 VSS.n767 VSS 3.75222
R2751 VSS.n2419 VSS 3.75222
R2752 VSS VSS.n4409 3.75222
R2753 VSS VSS.n3140 3.75222
R2754 VSS.n112 VSS 3.75222
R2755 VSS.n3459 VSS 3.53153
R2756 VSS.n1061 VSS.n1058 3.53153
R2757 VSS.n1086 VSS.n1085 3.53153
R2758 VSS.n1085 VSS.n1078 3.53153
R2759 VSS.n1141 VSS.n1140 3.53153
R2760 VSS.n1140 VSS.n1133 3.53153
R2761 VSS.n1156 VSS.n1149 3.53153
R2762 VSS.n1211 VSS.n1210 3.53153
R2763 VSS.n972 VSS.n971 3.53153
R2764 VSS.n971 VSS.n964 3.53153
R2765 VSS.n1648 VSS.n1641 3.53153
R2766 VSS.n2234 VSS.n2077 3.53153
R2767 VSS.n2086 VSS.n2078 3.53153
R2768 VSS.n2219 VSS.n2209 3.53153
R2769 VSS.n2211 VSS.n2210 3.53153
R2770 VSS.n2205 VSS.n2195 3.53153
R2771 VSS.n2197 VSS.n2196 3.53153
R2772 VSS.n2191 VSS.n2178 3.53153
R2773 VSS.n2174 VSS.n2164 3.53153
R2774 VSS.n2166 VSS.n2165 3.53153
R2775 VSS.n2137 VSS.n2127 3.53153
R2776 VSS.n2129 VSS.n2128 3.53153
R2777 VSS.n2123 VSS.n2104 3.53153
R2778 VSS.n2115 VSS.n2114 3.53153
R2779 VSS.n627 VSS.n623 3.53153
R2780 VSS.n2569 VSS.n590 3.53153
R2781 VSS.n2570 VSS.n584 3.53153
R2782 VSS.n2588 VSS.n2587 3.53153
R2783 VSS.n2610 VSS.n2600 3.53153
R2784 VSS.n2602 VSS.n2601 3.53153
R2785 VSS.n2627 VSS.n2614 3.53153
R2786 VSS.n2641 VSS.n2631 3.53153
R2787 VSS.n2633 VSS.n2632 3.53153
R2788 VSS.n2668 VSS.n2658 3.53153
R2789 VSS.n2660 VSS.n2659 3.53153
R2790 VSS.n2688 VSS.n2672 3.53153
R2791 VSS.n2680 VSS.n2679 3.53153
R2792 VSS.n2752 VSS.n2751 3.53153
R2793 VSS.n3651 VSS 3.53153
R2794 VSS.n4473 VSS.n4470 3.53153
R2795 VSS.n20 VSS.n17 3.53153
R2796 VSS.n3495 VSS 3.31084
R2797 VSS.n3665 VSS 3.31084
R2798 VSS.n1780 VSS.n1778 3.31084
R2799 VSS.n1780 VSS.n1779 3.31084
R2800 VSS.n938 VSS.n937 3.31084
R2801 VSS.n937 VSS.n930 3.31084
R2802 VSS.n1825 VSS.n1824 3.31084
R2803 VSS.n1824 VSS.n1817 3.31084
R2804 VSS.n1855 VSS.n1848 3.31084
R2805 VSS.n1839 VSS.n1838 3.31084
R2806 VSS.n1838 VSS.n1831 3.31084
R2807 VSS.n916 VSS.n915 3.31084
R2808 VSS.n915 VSS.n908 3.31084
R2809 VSS.n1999 VSS.n1998 3.31084
R2810 VSS.n1998 VSS.n1991 3.31084
R2811 VSS.n3312 VSS.n3310 3.31084
R2812 VSS.n2924 VSS.n2921 3.31084
R2813 VSS.n4894 VSS.n4893 3.31084
R2814 VSS.n326 VSS.n325 3.31084
R2815 VSS.n3657 VSS.n3656 3.1005
R2816 VSS.n3665 VSS.n3664 3.1005
R2817 VSS.n3454 VSS.n3453 3.1005
R2818 VSS.n3495 VSS.n3494 3.1005
R2819 VSS.n3431 VSS.n3430 3.1005
R2820 VSS.n3425 VSS.n3424 3.1005
R2821 VSS.n3408 VSS.n3407 3.1005
R2822 VSS.n3402 VSS.n3401 3.1005
R2823 VSS.n3398 VSS.n3397 3.1005
R2824 VSS.n3392 VSS.n3391 3.1005
R2825 VSS.n3388 VSS.n3387 3.1005
R2826 VSS.n3383 VSS.n3382 3.1005
R2827 VSS.n3377 VSS.n3376 3.1005
R2828 VSS.n3373 VSS.n3372 3.1005
R2829 VSS.n514 VSS.n513 3.1005
R2830 VSS.n520 VSS.n519 3.1005
R2831 VSS.n524 VSS.n523 3.1005
R2832 VSS.n530 VSS.n529 3.1005
R2833 VSS.n534 VSS.n533 3.1005
R2834 VSS.n540 VSS.n539 3.1005
R2835 VSS.n544 VSS.n543 3.1005
R2836 VSS.n550 VSS.n549 3.1005
R2837 VSS.n556 VSS.n555 3.1005
R2838 VSS.n509 VSS.n508 3.1005
R2839 VSS.n504 VSS.n503 3.1005
R2840 VSS.n3471 VSS.n3470 3.1005
R2841 VSS.n3466 VSS.n3465 3.1005
R2842 VSS.n3460 VSS.n3459 3.1005
R2843 VSS.n3651 VSS.n3650 3.1005
R2844 VSS.n3649 VSS.n3648 3.1005
R2845 VSS.n3643 VSS.n3642 3.1005
R2846 VSS.n3632 VSS.n3631 3.1005
R2847 VSS.n3622 VSS.n3621 3.1005
R2848 VSS.n3620 VSS.n3619 3.1005
R2849 VSS.n3616 VSS.n3615 3.1005
R2850 VSS.n3610 VSS.n3609 3.1005
R2851 VSS.n3605 VSS.n3604 3.1005
R2852 VSS.n3599 VSS.n3598 3.1005
R2853 VSS.n3308 VSS.n3307 3.1005
R2854 VSS.n3582 VSS.n3581 3.1005
R2855 VSS.n3571 VSS.n3570 3.1005
R2856 VSS.n3327 VSS.n3326 3.1005
R2857 VSS.n3541 VSS.n3540 3.1005
R2858 VSS.n3534 VSS.n3533 3.1005
R2859 VSS.n3528 VSS.n3527 3.1005
R2860 VSS.n3522 VSS.n3521 3.1005
R2861 VSS.n3518 VSS.n3517 3.1005
R2862 VSS.n3512 VSS.n3511 3.1005
R2863 VSS.n3508 VSS.n3507 3.1005
R2864 VSS.n3503 VSS.n3502 3.1005
R2865 VSS.n4740 VSS.n4735 3.1005
R2866 VSS.n4733 VSS.n4732 3.1005
R2867 VSS.n4729 VSS.n4728 3.1005
R2868 VSS.n4725 VSS.n4724 3.1005
R2869 VSS.n4718 VSS.n4717 3.1005
R2870 VSS.n4713 VSS.n4712 3.1005
R2871 VSS.n4709 VSS.n4708 3.1005
R2872 VSS.n4705 VSS.n4704 3.1005
R2873 VSS.n4698 VSS.n4697 3.1005
R2874 VSS.n2797 VSS.n2796 3.1005
R2875 VSS.n4679 VSS.n4678 3.1005
R2876 VSS.n4667 VSS.n4663 3.1005
R2877 VSS.n3835 VSS.n3834 3.1005
R2878 VSS.n3846 VSS.n3845 3.1005
R2879 VSS.n3850 VSS.n3849 3.1005
R2880 VSS.n3859 VSS.n3750 3.1005
R2881 VSS.n3711 VSS.n3710 3.1005
R2882 VSS.n3698 VSS.n3697 3.1005
R2883 VSS.n3693 VSS.n3692 3.1005
R2884 VSS.n3689 VSS.n3688 3.1005
R2885 VSS.n3682 VSS.n3681 3.1005
R2886 VSS.n3678 VSS.n3677 3.1005
R2887 VSS.n3673 VSS.n3672 3.1005
R2888 VSS.n3842 VSS.n3841 3.1005
R2889 VSS.n3825 VSS.n3824 3.1005
R2890 VSS.n3821 VSS.n3820 3.1005
R2891 VSS.n1499 VSS.n1498 3.1005
R2892 VSS.n5038 VSS.n5037 3.1005
R2893 VSS.n5052 VSS.n5051 3.1005
R2894 VSS.n4240 VSS.n4239 3.1005
R2895 VSS.n4252 VSS.n4251 3.1005
R2896 VSS.n4244 VSS.n4243 3.1005
R2897 VSS.n4152 VSS.n4151 3.1005
R2898 VSS.n4148 VSS.n4147 3.1005
R2899 VSS.n4143 VSS.n4142 3.1005
R2900 VSS.n4208 VSS.n4207 3.1005
R2901 VSS.n4179 VSS.n4178 3.1005
R2902 VSS.n4174 VSS.n4173 3.1005
R2903 VSS.n4170 VSS.n4169 3.1005
R2904 VSS.n4165 VSS.n4164 3.1005
R2905 VSS.n4326 VSS.n4325 3.1005
R2906 VSS.n4321 VSS.n4320 3.1005
R2907 VSS.n4366 VSS.n4365 3.1005
R2908 VSS.n4409 VSS.n4374 3.1005
R2909 VSS.n4508 VSS.n4507 3.1005
R2910 VSS.n3198 VSS.n3197 3.1005
R2911 VSS.n4404 VSS.n4403 3.1005
R2912 VSS.n4379 VSS.n4378 3.1005
R2913 VSS.n4480 VSS.n4479 3.1005
R2914 VSS.n3222 VSS.n3221 3.1005
R2915 VSS.n3217 VSS.n3216 3.1005
R2916 VSS.n4502 VSS.n4501 3.1005
R2917 VSS.n4548 VSS.n4547 3.1005
R2918 VSS.n4536 VSS.n4535 3.1005
R2919 VSS.n4437 VSS.n4436 3.1005
R2920 VSS.n4523 VSS.n4522 3.1005
R2921 VSS.n3171 VSS.n3170 3.1005
R2922 VSS.n3140 VSS.n3115 3.1005
R2923 VSS.n3094 VSS.n3093 3.1005
R2924 VSS.n3063 VSS.n3062 3.1005
R2925 VSS.n3067 VSS.n3066 3.1005
R2926 VSS.n3030 VSS.n3029 3.1005
R2927 VSS.n2999 VSS.n2998 3.1005
R2928 VSS.n2994 VSS.n2993 3.1005
R2929 VSS.n2980 VSS.n2979 3.1005
R2930 VSS.n2955 VSS.n2954 3.1005
R2931 VSS.n2933 VSS.n2932 3.1005
R2932 VSS.n2904 VSS.n2903 3.1005
R2933 VSS.n2899 VSS.n2898 3.1005
R2934 VSS.n4917 VSS.n4916 3.1005
R2935 VSS.n4932 VSS.n4931 3.1005
R2936 VSS.n4928 VSS.n4927 3.1005
R2937 VSS.n4876 VSS.n4875 3.1005
R2938 VSS.n4860 VSS.n4859 3.1005
R2939 VSS.n4854 VSS.n4853 3.1005
R2940 VSS.n4970 VSS.n4969 3.1005
R2941 VSS.n403 VSS.n402 3.1005
R2942 VSS.n413 VSS.n412 3.1005
R2943 VSS.n398 VSS.n397 3.1005
R2944 VSS.n393 VSS.n392 3.1005
R2945 VSS.n373 VSS.n372 3.1005
R2946 VSS.n377 VSS.n376 3.1005
R2947 VSS.n341 VSS.n340 3.1005
R2948 VSS.n350 VSS.n349 3.1005
R2949 VSS.n319 VSS.n318 3.1005
R2950 VSS.n298 VSS.n297 3.1005
R2951 VSS.n287 VSS.n286 3.1005
R2952 VSS.n156 VSS.n155 3.1005
R2953 VSS.n208 VSS.n207 3.1005
R2954 VSS.n225 VSS.n224 3.1005
R2955 VSS.n234 VSS.n233 3.1005
R2956 VSS.n249 VSS.n248 3.1005
R2957 VSS.n176 VSS.n175 3.1005
R2958 VSS.n5031 VSS.n5030 3.1005
R2959 VSS.n102 VSS.n101 3.1005
R2960 VSS.n83 VSS.n82 3.1005
R2961 VSS.n64 VSS.n63 3.1005
R2962 VSS.n60 VSS.n59 3.1005
R2963 VSS.n79 VSS.n78 3.1005
R2964 VSS.n15 VSS.n14 3.1005
R2965 VSS.n10 VSS.n9 3.1005
R2966 VSS.n6 VSS.n5 3.1005
R2967 VSS.n2026 VSS.n2025 3.1005
R2968 VSS.n2030 VSS.n2029 3.1005
R2969 VSS.n1953 VSS.n1952 3.1005
R2970 VSS.n1948 VSS.n1947 3.1005
R2971 VSS.n1899 VSS.n1898 3.1005
R2972 VSS.n1541 VSS.n1540 3.1005
R2973 VSS.n1536 VSS.n1535 3.1005
R2974 VSS.n1513 VSS.n1512 3.1005
R2975 VSS.n1503 VSS.n1502 3.1005
R2976 VSS.n1481 VSS.n1480 3.1005
R2977 VSS.n1458 VSS.n1457 3.1005
R2978 VSS.n1449 VSS.n1448 3.1005
R2979 VSS.n1427 VSS.n1426 3.1005
R2980 VSS.n1590 VSS.n1589 3.1005
R2981 VSS.n1585 VSS.n1584 3.1005
R2982 VSS.n1581 VSS.n1580 3.1005
R2983 VSS.n1278 VSS.n1277 3.1005
R2984 VSS.n1282 VSS.n1281 3.1005
R2985 VSS.n1267 VSS.n1266 3.1005
R2986 VSS.n1182 VSS.n1181 3.1005
R2987 VSS.n1178 VSS.n1177 3.1005
R2988 VSS.n1409 VSS.n1408 3.1005
R2989 VSS.n860 VSS.n859 3.1005
R2990 VSS.n2495 VSS.n2494 3.1005
R2991 VSS.n2499 VSS.n2498 3.1005
R2992 VSS.n4825 VSS.n4824 3.1005
R2993 VSS.n4813 VSS.n4812 3.1005
R2994 VSS.n4263 VSS.n4262 3.1005
R2995 VSS.n4268 VSS.n4267 3.1005
R2996 VSS.n4272 VSS.n4271 3.1005
R2997 VSS.n4276 VSS.n4275 3.1005
R2998 VSS.n4282 VSS.n4281 3.1005
R2999 VSS.n4286 VSS.n4285 3.1005
R3000 VSS.n4290 VSS.n4289 3.1005
R3001 VSS.n4294 VSS.n4293 3.1005
R3002 VSS.n4299 VSS.n4298 3.1005
R3003 VSS.n4303 VSS.n4302 3.1005
R3004 VSS.n3930 VSS.n3929 3.1005
R3005 VSS.n3925 VSS.n3924 3.1005
R3006 VSS.n4113 VSS.n4112 3.1005
R3007 VSS.n4258 VSS.n4257 3.1005
R3008 VSS.n3967 VSS.n3966 3.1005
R3009 VSS.n3949 VSS.n3948 3.1005
R3010 VSS.n3983 VSS.n3982 3.1005
R3011 VSS.n4089 VSS.n4088 3.1005
R3012 VSS.n4081 VSS.n4080 3.1005
R3013 VSS.n4072 VSS.n4071 3.1005
R3014 VSS.n4068 VSS.n4067 3.1005
R3015 VSS.n4064 VSS.n4063 3.1005
R3016 VSS.n4060 VSS.n4059 3.1005
R3017 VSS.n4054 VSS.n4053 3.1005
R3018 VSS.n4050 VSS.n4049 3.1005
R3019 VSS.n4046 VSS.n4045 3.1005
R3020 VSS.n4042 VSS.n4041 3.1005
R3021 VSS.n4037 VSS.n4036 3.1005
R3022 VSS.n4033 VSS.n4032 3.1005
R3023 VSS.n4029 VSS.n4028 3.1005
R3024 VSS.n4025 VSS.n4024 3.1005
R3025 VSS.n4021 VSS.n4020 3.1005
R3026 VSS.n4015 VSS.n4014 3.1005
R3027 VSS.n4011 VSS.n4010 3.1005
R3028 VSS.n3998 VSS.n3997 3.1005
R3029 VSS.n3994 VSS.n3993 3.1005
R3030 VSS.n4580 VSS.n4579 3.1005
R3031 VSS.n4601 VSS.n4599 3.1005
R3032 VSS.n2881 VSS.n2880 3.1005
R3033 VSS.n2869 VSS.n2868 3.1005
R3034 VSS.n2865 VSS.n2864 3.1005
R3035 VSS.n2859 VSS.n2858 3.1005
R3036 VSS.n2855 VSS.n2854 3.1005
R3037 VSS.n2851 VSS.n2850 3.1005
R3038 VSS.n2847 VSS.n2846 3.1005
R3039 VSS.n2842 VSS.n2841 3.1005
R3040 VSS.n2838 VSS.n2837 3.1005
R3041 VSS.n2834 VSS.n2833 3.1005
R3042 VSS.n439 VSS.n438 3.1005
R3043 VSS.n445 VSS.n444 3.1005
R3044 VSS.n449 VSS.n448 3.1005
R3045 VSS.n453 VSS.n452 3.1005
R3046 VSS.n457 VSS.n456 3.1005
R3047 VSS.n461 VSS.n460 3.1005
R3048 VSS.n466 VSS.n465 3.1005
R3049 VSS.n470 VSS.n469 3.1005
R3050 VSS.n4631 VSS.n4630 3.1005
R3051 VSS.n4795 VSS.n4794 3.1005
R3052 VSS.n4786 VSS.n4785 3.1005
R3053 VSS.n702 VSS.n701 3.1005
R3054 VSS.n706 VSS.n705 3.1005
R3055 VSS.n711 VSS.n710 3.1005
R3056 VSS.n716 VSS.n715 3.1005
R3057 VSS.n720 VSS.n719 3.1005
R3058 VSS.n724 VSS.n723 3.1005
R3059 VSS.n728 VSS.n727 3.1005
R3060 VSS.n732 VSS.n731 3.1005
R3061 VSS.n738 VSS.n737 3.1005
R3062 VSS.n742 VSS.n741 3.1005
R3063 VSS.n746 VSS.n745 3.1005
R3064 VSS.n750 VSS.n749 3.1005
R3065 VSS.n754 VSS.n753 3.1005
R3066 VSS.n759 VSS.n758 3.1005
R3067 VSS.n763 VSS.n762 3.1005
R3068 VSS.n766 VSS.n765 3.1005
R3069 VSS.n768 VSS.n767 3.1005
R3070 VSS.n773 VSS.n772 3.1005
R3071 VSS.n657 VSS.n656 3.1005
R3072 VSS.n796 VSS.n795 3.1005
R3073 VSS.n2481 VSS.n2480 3.1005
R3074 VSS.n819 VSS.n818 3.1005
R3075 VSS.n2472 VSS.n2471 3.1005
R3076 VSS.n2456 VSS.n2455 3.1005
R3077 VSS.n2452 VSS.n2451 3.1005
R3078 VSS.n2448 VSS.n2447 3.1005
R3079 VSS.n2438 VSS.n2437 3.1005
R3080 VSS.n2434 VSS.n2433 3.1005
R3081 VSS.n2424 VSS.n2423 3.1005
R3082 VSS.n2419 VSS.n2418 3.1005
R3083 VSS.n2411 VSS.n2410 3.1005
R3084 VSS.n2402 VSS.n2401 3.1005
R3085 VSS.n2398 VSS.n2397 3.1005
R3086 VSS.n2394 VSS.n2393 3.1005
R3087 VSS.n2390 VSS.n2389 3.1005
R3088 VSS.n2384 VSS.n2383 3.1005
R3089 VSS.n2380 VSS.n2379 3.1005
R3090 VSS.n831 VSS.n830 3.1005
R3091 VSS.n845 VSS.n844 3.1005
R3092 VSS.n882 VSS.n881 3.1005
R3093 VSS.n1933 VSS.n1932 3.1005
R3094 VSS.n1881 VSS.n1880 3.1005
R3095 VSS.n1876 VSS.n1875 3.1005
R3096 VSS.n1321 VSS.n1320 3.1005
R3097 VSS.n1345 VSS.n1344 3.1005
R3098 VSS.n1310 VSS.n1309 3.1005
R3099 VSS.n1357 VSS.n1356 3.1005
R3100 VSS.n1362 VSS.n1361 3.1005
R3101 VSS.n1366 VSS.n1365 3.1005
R3102 VSS.n1370 VSS.n1369 3.1005
R3103 VSS.n1376 VSS.n1375 3.1005
R3104 VSS.n1380 VSS.n1379 3.1005
R3105 VSS.n1384 VSS.n1383 3.1005
R3106 VSS.n1388 VSS.n1387 3.1005
R3107 VSS.n1393 VSS.n1392 3.1005
R3108 VSS.n1397 VSS.n1396 3.1005
R3109 VSS.n1401 VSS.n1400 3.1005
R3110 VSS.n1405 VSS.n1404 3.1005
R3111 VSS.n1252 VSS.n1251 3.1005
R3112 VSS.n1113 VSS.n1112 3.1005
R3113 VSS.n1102 VSS.n1101 3.1005
R3114 VSS.n1002 VSS.n1001 3.1005
R3115 VSS.n1300 VSS.n1297 3.09016
R3116 VSS.n3903 VSS.n3902 3.09016
R3117 VSS.n3507 VSS.n3504 3.09016
R3118 VSS.n3546 VSS.n3543 3.09016
R3119 VSS.n3540 VSS.n3537 3.09016
R3120 VSS.n508 VSS.n505 3.09016
R3121 VSS.n529 VSS.n526 3.09016
R3122 VSS.n3228 VSS.n3227 3.09016
R3123 VSS.n5043 VSS.n5042 3.09016
R3124 VSS.n917 VSS.n916 3.03311
R3125 VSS.n1858 VSS.n1857 3.03311
R3126 VSS.n3739 VSS.n3738 3.03311
R3127 VSS.n2531 VSS.n2530 3.03311
R3128 VSS.n4567 VSS.n4564 2.86947
R3129 VSS.n685 VSS.n682 2.86947
R3130 VSS.n1164 VSS.n1163 2.86947
R3131 VSS.n2716 VSS.n2715 2.86947
R3132 VSS.n4331 VSS.n4330 2.86947
R3133 VSS.n4541 VSS.n4538 2.86947
R3134 VSS.n1756 VSS.n1755 2.7891
R3135 VSS.n2246 VSS.n2075 2.7891
R3136 VSS.n2226 VSS.n2225 2.7891
R3137 VSS.n2583 VSS.n2581 2.7891
R3138 VSS.n3694 VSS.n3296 2.68147
R3139 VSS.n3831 VSS.n3830 2.68147
R3140 VSS.n4694 VSS.n2790 2.68147
R3141 VSS.n4714 VSS.n2785 2.68147
R3142 VSS.n1924 VSS.n1921 2.64878
R3143 VSS.n1335 VSS.n1332 2.64878
R3144 VSS.n1857 VSS.n1856 2.64878
R3145 VSS.n4724 VSS.n4721 2.64878
R3146 VSS.n2802 VSS.n2799 2.64878
R3147 VSS.n3335 VSS.n3332 2.64878
R3148 VSS.n3135 VSS.n3117 2.64878
R3149 VSS.n1020 VSS.n1019 2.62699
R3150 VSS.n97 VSS.n96 2.60389
R3151 VSS.n4889 VSS.n4888 2.52719
R3152 VSS.n4428 VSS.n4427 2.52719
R3153 VSS.n1546 VSS.n1545 2.52719
R3154 VSS.n1358 VSS.n1308 2.52719
R3155 VSS.n778 VSS.n777 2.52719
R3156 VSS.n1033 VSS.n1032 2.52719
R3157 VSS.n130 VSS.n129 2.52719
R3158 VSS.n3150 VSS.n3149 2.52719
R3159 VSS.n5006 VSS.n5005 2.52719
R3160 VSS.n4077 VSS.n4076 2.52719
R3161 VSS.n4264 VSS.n4134 2.52719
R3162 VSS.n2407 VSS.n2406 2.52719
R3163 VSS.n3056 VSS.n3055 2.51853
R3164 VSS.n4940 VSS.n4939 2.51853
R3165 VSS.n1492 VSS.n1491 2.51853
R3166 VSS.n4233 VSS.n4232 2.51853
R3167 VSS.n4675 VSS.n4674 2.49102
R3168 VSS.n3853 VSS.n3851 2.49102
R3169 VSS.n3674 VSS.n3298 2.49102
R3170 VSS.n4734 VSS.n2780 2.49102
R3171 VSS.n3639 VSS.n3638 2.49102
R3172 VSS.n3477 VSS.n3476 2.49102
R3173 VSS.n1528 VSS.n1527 2.49102
R3174 VSS.n107 VSS.n105 2.49102
R3175 VSS.n4906 VSS.n4880 2.49102
R3176 VSS.n3144 VSS.n3143 2.49102
R3177 VSS.n4413 VSS.n4412 2.49102
R3178 VSS.n283 VSS.n281 2.49102
R3179 VSS.n1027 VSS.n1026 2.49102
R3180 VSS.n1353 VSS.n1352 2.49102
R3181 VSS.n769 VSS.n664 2.49102
R3182 VSS.n4823 VSS.n4822 2.49102
R3183 VSS.n4627 VSS.n4626 2.49102
R3184 VSS.n4087 VSS.n4086 2.49102
R3185 VSS.n4259 VSS.n4136 2.49102
R3186 VSS.n2417 VSS.n2416 2.49102
R3187 VSS.n3663 VSS.n3662 2.49101
R3188 VSS.n3253 VSS.n3252 2.45
R3189 VSS.n294 VSS.n293 2.45
R3190 VSS.n1108 VSS.n1107 2.45
R3191 VSS.n1317 VSS.n1316 2.45
R3192 VSS.n755 VSS.n680 2.45
R3193 VSS.n4576 VSS.n4575 2.45
R3194 VSS.n3955 VSS.n3954 2.45
R3195 VSS.n462 VSS.n435 2.45
R3196 VSS.n2444 VSS.n2443 2.45
R3197 VSS.n1510 VSS.n1509 2.43201
R3198 VSS.n317 VSS.n316 2.43201
R3199 VSS.n4923 VSS.n4922 2.43201
R3200 VSS.n3101 VSS.n3100 2.43201
R3201 VSS.n4250 VSS.n4249 2.43201
R3202 VSS.n4398 VSS.n4397 2.43201
R3203 VSS.n1003 VSS.n998 2.43201
R3204 VSS.n1343 VSS.n1342 2.43201
R3205 VSS.n764 VSS.n675 2.43201
R3206 VSS.n4608 VSS.n4607 2.43201
R3207 VSS.n3989 VSS.n3988 2.43201
R3208 VSS.n476 VSS.n475 2.43201
R3209 VSS.n2430 VSS.n2429 2.43201
R3210 VSS.n3935 VSS.n3934 2.42809
R3211 VSS.n3688 VSS.n3685 2.42809
R3212 VSS.n3841 VSS.n3838 2.42809
R3213 VSS.n3762 VSS.n3761 2.42809
R3214 VSS.n1618 VSS.n1617 2.42809
R3215 VSS.n1662 VSS.n1655 2.42809
R3216 VSS.n1664 VSS.n1662 2.42809
R3217 VSS.n1676 VSS.n1669 2.42809
R3218 VSS.n1678 VSS.n1676 2.42809
R3219 VSS.n1703 VSS.n1696 2.42809
R3220 VSS.n1705 VSS.n1703 2.42809
R3221 VSS.n1719 VSS.n1712 2.42809
R3222 VSS.n1721 VSS.n1719 2.42809
R3223 VSS.n1733 VSS.n1726 2.42809
R3224 VSS.n1735 VSS.n1733 2.42809
R3225 VSS.n1747 VSS.n1740 2.42809
R3226 VSS.n1749 VSS.n1747 2.42809
R3227 VSS.n1764 VSS.n953 2.42809
R3228 VSS.n1772 VSS.n1764 2.42809
R3229 VSS.n2358 VSS.n2351 2.42809
R3230 VSS.n2360 VSS.n2358 2.42809
R3231 VSS.n2335 VSS.n2328 2.42809
R3232 VSS.n2337 VSS.n2335 2.42809
R3233 VSS.n2318 VSS.n2311 2.42809
R3234 VSS.n2320 VSS.n2318 2.42809
R3235 VSS.n2304 VSS.n2297 2.42809
R3236 VSS.n2306 VSS.n2304 2.42809
R3237 VSS.n2288 VSS.n2281 2.42809
R3238 VSS.n2290 VSS.n2288 2.42809
R3239 VSS.n2274 VSS.n2267 2.42809
R3240 VSS.n2276 VSS.n2274 2.42809
R3241 VSS.n2254 VSS.n2239 2.42809
R3242 VSS.n2259 VSS.n2254 2.42809
R3243 VSS.n2539 VSS.n2535 2.42809
R3244 VSS.n2744 VSS.n2740 2.42809
R3245 VSS.n2770 VSS.n2766 2.42809
R3246 VSS.n2796 VSS.n2793 2.42809
R3247 VSS.n1905 VSS.n1904 2.42809
R3248 VSS.n1595 VSS.n1594 2.42809
R3249 VSS.n4198 VSS.n4197 2.36358
R3250 VSS.n4960 VSS.n4959 2.36358
R3251 VSS.n198 VSS.n197 2.36358
R3252 VSS.n3449 VSS.n3448 2.32777
R3253 VSS.n3866 VSS.n3749 2.32777
R3254 VSS.n4654 VSS.n4653 2.32777
R3255 VSS.n1073 VSS.n1072 2.32777
R3256 VSS.n1794 VSS.n1793 2.32777
R3257 VSS.n2557 VSS.n2556 2.32777
R3258 VSS.n4751 VSS.n4750 2.32777
R3259 VSS.n3578 VSS.n3577 2.28739
R3260 VSS.n1037 VSS.n1036 2.28739
R3261 VSS.n1548 VSS.n1532 2.28739
R3262 VSS.n4433 VSS.n4432 2.28739
R3263 VSS.n4531 VSS.n4530 2.28739
R3264 VSS.n3106 VSS.n3105 2.28739
R3265 VSS.n3026 VSS.n3025 2.28739
R3266 VSS.n2909 VSS.n2908 2.28739
R3267 VSS.n409 VSS.n408 2.28739
R3268 VSS.n346 VSS.n345 2.28739
R3269 VSS.n5011 VSS.n5010 2.28739
R3270 VSS.n230 VSS.n229 2.28739
R3271 VSS.n125 VSS.n124 2.28739
R3272 VSS.n113 VSS.n112 2.28739
R3273 VSS.n1958 VSS.n1957 2.28739
R3274 VSS.n1521 VSS.n1520 2.28739
R3275 VSS.n1454 VSS.n1453 2.28739
R3276 VSS.n1274 VSS.n1273 2.28739
R3277 VSS.n4184 VSS.n4183 2.28739
R3278 VSS.n993 VSS.n992 2.28739
R3279 VSS.n1886 VSS.n1885 2.28739
R3280 VSS.n2501 VSS.n2476 2.28739
R3281 VSS.n4094 VSS.n4093 2.28739
R3282 VSS.n4619 VSS.n4618 2.28739
R3283 VSS.n4791 VSS.n4790 2.28739
R3284 VSS.n662 VSS.n661 2.28739
R3285 VSS.n2375 VSS.n864 2.28739
R3286 VSS.n1248 VSS.n1247 2.28739
R3287 VSS.n1118 VSS.n1117 2.28739
R3288 VSS.n4653 VSS.n4652 2.28336
R3289 VSS.n3875 VSS.n3749 2.28314
R3290 VSS.n2183 VSS.n2182 2.2074
R3291 VSS.n2619 VSS.n2618 2.2074
R3292 VSS.n3615 VSS.n3612 2.2074
R3293 VSS.n3407 VSS.n3404 2.2074
R3294 VSS.n3413 VSS.n3410 2.2074
R3295 VSS.n4384 VSS.n4381 2.2074
R3296 VSS.n418 VSS.n417 2.2074
R3297 VSS.n1020 VSS.n984 2.2074
R3298 VSS.n486 VSS.n485 2.16388
R3299 VSS.n1791 VSS.n1788 2.06672
R3300 VSS.n4127 VSS.n4124 1.98671
R3301 VSS.n3465 VSS.n3462 1.98671
R3302 VSS.n3289 VSS.n3276 1.98671
R3303 VSS.n3901 VSS.n3900 1.98671
R3304 VSS.n3648 VSS.n3645 1.98671
R3305 VSS.n3436 VSS.n3433 1.98671
R3306 VSS.n2948 VSS.n2945 1.98671
R3307 VSS VSS.n4910 1.98671
R3308 VSS.n2364 VSS.n2363 1.94045
R3309 VSS.n2042 VSS.n2041 1.94045
R3310 VSS.n2003 VSS.n2002 1.94045
R3311 VSS.n3712 VSS.n3291 1.94045
R3312 VSS.n2518 VSS.n2517 1.94045
R3313 VSS.n2102 VSS.n2101 1.94045
R3314 VSS.n3493 VSS.n3492 1.94045
R3315 VSS VSS.n4402 1.94045
R3316 VSS.n1225 VSS.n1224 1.92698
R3317 VSS.n1691 VSS.n1690 1.81037
R3318 VSS.n901 VSS.n900 1.81037
R3319 VSS.n2073 VSS.n2072 1.81037
R3320 VSS.n2654 VSS.n2652 1.81037
R3321 VSS.n824 VSS.n821 1.76602
R3322 VSS.n3276 VSS.n3275 1.76602
R3323 VSS.n4421 VSS.n4420 1.76602
R3324 VSS.n3004 VSS.n3001 1.76602
R3325 VSS.n4910 VSS.n4909 1.76602
R3326 VSS.n363 VSS.n360 1.76602
R3327 VSS.n73 VSS.n71 1.76531
R3328 VSS.n74 VSS.n73 1.75392
R3329 VSS.n3988 VSS.n3986 1.72554
R3330 VSS.n4607 VSS.n4605 1.72554
R3331 VSS.n675 VSS.n673 1.72554
R3332 VSS.n1342 VSS.n1340 1.72554
R3333 VSS.n998 VSS.n996 1.72554
R3334 VSS.n3100 VSS.n3098 1.72554
R3335 VSS.n4922 VSS.n4920 1.72554
R3336 VSS.n1509 VSS.n1507 1.72554
R3337 VSS.n4249 VSS.n4247 1.72554
R3338 VSS.n4397 VSS.n4395 1.72554
R3339 VSS.n316 VSS.n314 1.72554
R3340 VSS.n475 VSS.n473 1.72554
R3341 VSS.n2429 VSS.n2427 1.72554
R3342 VSS.n680 VSS.n678 1.67882
R3343 VSS.n2443 VSS.n2441 1.67882
R3344 VSS.n1107 VSS.n1105 1.67882
R3345 VSS.n293 VSS.n291 1.67882
R3346 VSS.n3252 VSS.n3250 1.67882
R3347 VSS.n4575 VSS.n4573 1.67882
R3348 VSS.n3954 VSS.n3952 1.67882
R3349 VSS.n435 VSS.n433 1.67882
R3350 VSS.n1316 VSS.n1314 1.67882
R3351 VSS.n1758 VSS.n1757 1.61124
R3352 VSS.n2248 VSS.n2247 1.61124
R3353 VSS.n4137 VSS.n4136 1.57241
R3354 VSS.n4086 VSS.n4084 1.57241
R3355 VSS.n4626 VSS.n4624 1.57241
R3356 VSS.n666 VSS.n664 1.57241
R3357 VSS.n2416 VSS.n2414 1.57241
R3358 VSS.n1352 VSS.n1350 1.57241
R3359 VSS.n3476 VSS.n3474 1.57241
R3360 VSS.n3638 VSS.n3636 1.57241
R3361 VSS.n2780 VSS.n2778 1.57241
R3362 VSS.n3299 VSS.n3298 1.57241
R3363 VSS.n3854 VSS.n3853 1.57241
R3364 VSS.n4674 VSS.n4672 1.57241
R3365 VSS.n3143 VSS.n3141 1.57241
R3366 VSS.n1527 VSS.n1525 1.57241
R3367 VSS.n1026 VSS.n1024 1.57241
R3368 VSS.n108 VSS.n107 1.57241
R3369 VSS.n4412 VSS.n4410 1.57241
R3370 VSS.n4911 VSS.n4880 1.57241
R3371 VSS.n324 VSS.n283 1.57241
R3372 VSS.n4822 VSS.n4820 1.57241
R3373 VSS.n3662 VSS.n3661 1.57193
R3374 VSS.n4298 VSS.n4295 1.54533
R3375 VSS.n3960 VSS.n3957 1.54533
R3376 VSS.n4041 VSS.n4038 1.54533
R3377 VSS.n2846 VSS.n2843 1.54533
R3378 VSS.n715 VSS.n712 1.54533
R3379 VSS.n2480 VSS.n2477 1.54533
R3380 VSS.n859 VSS.n856 1.54533
R3381 VSS.n1392 VSS.n1389 1.54533
R3382 VSS.n4357 VSS.n4354 1.54533
R3383 VSS.n4164 VSS.n4163 1.54533
R3384 VSS.n4501 VSS.n4500 1.54533
R3385 VSS.n2973 VSS.n2970 1.54533
R3386 VSS.n397 VSS.n396 1.54533
R3387 VSS.n169 VSS.n166 1.54533
R3388 VSS.n248 VSS.n245 1.54533
R3389 VSS.n2018 VSS.n2017 1.54533
R3390 VSS.n1580 VSS.n1579 1.54533
R3391 VSS.n3738 VSS.n3737 1.50638
R3392 VSS.n3788 VSS.n3787 1.50638
R3393 VSS.n1231 VSS.n1230 1.50638
R3394 VSS.n2157 VSS.n2156 1.50638
R3395 VSS.n598 VSS.n597 1.50638
R3396 VSS.n2735 VSS.n2734 1.50638
R3397 VSS.n4134 VSS.n4133 1.47868
R3398 VSS.n4076 VSS.n4075 1.47868
R3399 VSS.n2406 VSS.n2405 1.47868
R3400 VSS.n3149 VSS.n3148 1.47868
R3401 VSS.n5005 VSS.n5004 1.47868
R3402 VSS.n129 VSS.n128 1.47868
R3403 VSS.n1032 VSS.n1031 1.47868
R3404 VSS.n4888 VSS.n4887 1.47868
R3405 VSS.n4427 VSS.n4426 1.47868
R3406 VSS.n1545 VSS.n1544 1.47868
R3407 VSS.n1308 VSS.n1307 1.47868
R3408 VSS.n777 VSS.n776 1.47868
R3409 VSS.n2721 VSS.n2719 1.35607
R3410 VSS.n2526 VSS.n2525 1.35607
R3411 VSS.n1091 VSS.n1090 1.35607
R3412 VSS.n1167 VSS.n1166 1.35607
R3413 VSS.n1616 VSS.n1615 1.35607
R3414 VSS.n1797 VSS.n1796 1.35607
R3415 VSS.n2146 VSS.n2145 1.35607
R3416 VSS.n1863 VSS.n1860 1.35607
R3417 VSS.n1976 VSS.n1975 1.35607
R3418 VSS.n3774 VSS.n3773 1.35607
R3419 VSS.n3881 VSS.n3880 1.35607
R3420 VSS.n3906 VSS.n3905 1.35607
R3421 VSS.n3741 VSS.n3740 1.35607
R3422 VSS.n3715 VSS.n3714 1.35607
R3423 VSS.n634 VSS.n632 1.35607
R3424 VSS.n4757 VSS.n4756 1.35607
R3425 VSS.n4692 VSS.n4691 1.35607
R3426 VSS.n4650 VSS.n4649 1.35607
R3427 VSS.n3422 VSS.n3421 1.35607
R3428 VSS.n3484 VSS.n3482 1.35607
R3429 VSS.n567 VSS.n565 1.35607
R3430 VSS.n3443 VSS.n3442 1.35607
R3431 VSS.n3552 VSS.n3550 1.35607
R3432 VSS.n3586 VSS.n3584 1.35607
R3433 VSS.n4483 VSS.n4482 1.35607
R3434 VSS.n4551 VSS.n4550 1.35607
R3435 VSS.n4511 VSS.n4510 1.35607
R3436 VSS.n3010 VSS.n3008 1.35607
R3437 VSS.n55 VSS.n54 1.35607
R3438 VSS.n1519 VSS.n1518 1.35607
R3439 VSS.n1440 VSS.n1439 1.35607
R3440 VSS.n115 VSS.n114 1.35607
R3441 VSS.n261 VSS.n259 1.35607
R3442 VSS.n4391 VSS.n4390 1.35607
R3443 VSS.n3209 VSS.n3208 1.35607
R3444 VSS.n354 VSS.n352 1.35607
R3445 VSS.n160 VSS.n158 1.35607
R3446 VSS.n212 VSS.n210 1.35607
R3447 VSS.n4944 VSS.n4942 1.35607
R3448 VSS.n4904 VSS.n4903 1.35607
R3449 VSS.n332 VSS.n330 1.35607
R3450 VSS.n381 VSS.n379 1.35607
R3451 VSS.n2959 VSS.n2957 1.35607
R3452 VSS.n4369 VSS.n4368 1.35607
R3453 VSS.n3071 VSS.n3069 1.35607
R3454 VSS.n3131 VSS.n3130 1.35607
R3455 VSS.n4864 VSS.n4862 1.35607
R3456 VSS.n424 VSS.n422 1.35607
R3457 VSS.n310 VSS.n309 1.35607
R3458 VSS.n180 VSS.n178 1.35607
R3459 VSS.n134 VSS.n132 1.35607
R3460 VSS.n1486 VSS.n1485 1.35607
R3461 VSS.n1040 VSS.n1038 1.35607
R3462 VSS.n1194 VSS.n1192 1.35607
R3463 VSS.n1462 VSS.n1460 1.35607
R3464 VSS.n2034 VSS.n2032 1.35607
R3465 VSS.n1962 VSS.n1959 1.35607
R3466 VSS.n1911 VSS.n1909 1.35607
R3467 VSS.n28 VSS.n26 1.35607
R3468 VSS.n3235 VSS.n3233 1.35607
R3469 VSS.n3257 VSS.n3255 1.35607
R3470 VSS.n4337 VSS.n4335 1.35607
R3471 VSS.n4212 VSS.n4210 1.35607
R3472 VSS.n4186 VSS.n4185 1.35607
R3473 VSS.n4830 VSS.n4828 1.35607
R3474 VSS.n1006 VSS.n1005 1.35607
R3475 VSS.n1255 VSS.n1254 1.35607
R3476 VSS.n1888 VSS.n1887 1.35607
R3477 VSS.n2885 VSS.n2883 1.35607
R3478 VSS.n4635 VSS.n4633 1.35607
R3479 VSS.n4307 VSS.n4305 1.35607
R3480 VSS.n4117 VSS.n4115 1.35607
R3481 VSS.n4006 VSS.n4005 1.35607
R3482 VSS.n3971 VSS.n3969 1.35607
R3483 VSS.n697 VSS.n696 1.35607
R3484 VSS.n4799 VSS.n4797 1.35607
R3485 VSS.n782 VSS.n780 1.35607
R3486 VSS.n1937 VSS.n1935 1.35607
R3487 VSS.n886 VSS.n884 1.35607
R3488 VSS.n1412 VSS.n1411 1.35607
R3489 VSS.n1235 VSS.n1233 1.35607
R3490 VSS.n2756 VSS.n2755 1.35607
R3491 VSS.n4683 VSS.n4681 1.35607
R3492 VSS.n3341 VSS.n3339 1.35607
R3493 VSS.n3594 VSS.n3593 1.35607
R3494 VSS.n4441 VSS.n4439 1.35607
R3495 VSS.n3182 VSS.n3181 1.35607
R3496 VSS.n3160 VSS.n3159 1.35607
R3497 VSS.n3108 VSS.n3107 1.35607
R3498 VSS.n3033 VSS.n3032 1.35607
R3499 VSS.n2983 VSS.n2982 1.35607
R3500 VSS.n5013 VSS.n5012 1.35607
R3501 VSS.n4973 VSS.n4972 1.35607
R3502 VSS.n2911 VSS.n2910 1.35607
R3503 VSS.n2936 VSS.n2935 1.35607
R3504 VSS.n237 VSS.n236 1.35607
R3505 VSS.n5063 VSS.n5061 1.35607
R3506 VSS.n91 VSS.n90 1.35607
R3507 VSS.n1286 VSS.n1284 1.35607
R3508 VSS.n1601 VSS.n1599 1.35607
R3509 VSS.n4227 VSS.n4226 1.35607
R3510 VSS.n4617 VSS.n4616 1.35607
R3511 VSS.n4808 VSS.n4807 1.35607
R3512 VSS.n834 VSS.n833 1.35607
R3513 VSS.n1122 VSS.n1119 1.35607
R3514 VSS.n1329 VSS.n1328 1.35607
R3515 VSS.n807 VSS.n806 1.35607
R3516 VSS.n4583 VSS.n4582 1.35607
R3517 VSS.n4096 VSS.n4095 1.35607
R3518 VSS.n3940 VSS.n3939 1.35607
R3519 VSS.n2874 VSS.n2871 1.32464
R3520 VSS.n3766 VSS.n3762 1.32464
R3521 VSS.n3766 VSS.n3765 1.32464
R3522 VSS.n1655 VSS.n1654 1.32464
R3523 VSS.n1664 VSS.n1663 1.32464
R3524 VSS.n1669 VSS.n1668 1.32464
R3525 VSS.n1678 VSS.n1677 1.32464
R3526 VSS.n1696 VSS.n1695 1.32464
R3527 VSS.n1705 VSS.n1704 1.32464
R3528 VSS.n1712 VSS.n1711 1.32464
R3529 VSS.n1721 VSS.n1720 1.32464
R3530 VSS.n1726 VSS.n1725 1.32464
R3531 VSS.n1735 VSS.n1734 1.32464
R3532 VSS.n1740 VSS.n1739 1.32464
R3533 VSS.n1749 VSS.n1748 1.32464
R3534 VSS.n953 VSS.n952 1.32464
R3535 VSS.n1772 VSS.n1771 1.32464
R3536 VSS.n2351 VSS.n2350 1.32464
R3537 VSS.n2360 VSS.n2359 1.32464
R3538 VSS.n2328 VSS.n2327 1.32464
R3539 VSS.n2337 VSS.n2336 1.32464
R3540 VSS.n2311 VSS.n2310 1.32464
R3541 VSS.n2320 VSS.n2319 1.32464
R3542 VSS.n2297 VSS.n2296 1.32464
R3543 VSS.n2306 VSS.n2305 1.32464
R3544 VSS.n2281 VSS.n2280 1.32464
R3545 VSS.n2290 VSS.n2289 1.32464
R3546 VSS.n2267 VSS.n2266 1.32464
R3547 VSS.n2276 VSS.n2275 1.32464
R3548 VSS.n2239 VSS.n2238 1.32464
R3549 VSS.n2259 VSS.n2258 1.32464
R3550 VSS.n2182 VSS.n2181 1.32464
R3551 VSS.n2618 VSS.n2617 1.32464
R3552 VSS.n2766 VSS.n2765 1.32464
R3553 VSS.n3622 VSS.n3302 1.32464
R3554 VSS.n3425 VSS.n3367 1.32464
R3555 VSS.n3204 VSS.n3203 1.32464
R3556 VSS.n3045 VSS.n3042 1.32464
R3557 VSS.n1188 VSS.n1187 1.32464
R3558 VSS.n3744 VSS.n3266 1.13857
R3559 VSS.n4401 VSS.n4349 1.13857
R3560 VSS.n216 VSS.n186 1.13845
R3561 VSS.n4765 VSS.n4764 1.13845
R3562 VSS.n4779 VSS.n4778 1.13845
R3563 VSS.n4977 VSS.n4842 1.13845
R3564 VSS.n3491 VSS.n3488 1.13845
R3565 VSS.n3563 VSS.n3558 1.13845
R3566 VSS.n4348 VSS.n4347 1.13845
R3567 VSS.n495 VSS.n494 1.13746
R3568 VSS.n2096 VSS.n2095 1.13469
R3569 VSS.n2522 VSS.n2521 1.13469
R3570 VSS.n2098 VSS.n2097 1.13469
R3571 VSS.n837 VSS.n836 1.13469
R3572 VSS.n2505 VSS.n2504 1.13469
R3573 VSS.n810 VSS.n809 1.13469
R3574 VSS.n240 VSS.n239 1.13469
R3575 VSS.n2759 VSS.n2758 1.13469
R3576 VSS.n4804 VSS.n4803 1.13469
R3577 VSS.n4976 VSS.n4953 1.13469
R3578 VSS.n4976 VSS.n4975 1.13469
R3579 VSS.n574 VSS.n573 1.13469
R3580 VSS.n4687 VSS.n4686 1.13469
R3581 VSS.n4613 VSS.n4588 1.13469
R3582 VSS.n4586 VSS.n4585 1.13469
R3583 VSS.n3185 VSS.n3184 1.13469
R3584 VSS.n3163 VSS.n3162 1.13469
R3585 VSS.n3111 VSS.n3110 1.13469
R3586 VSS.n3363 VSS.n3362 1.13469
R3587 VSS.n3589 VSS.n3344 1.13469
R3588 VSS.n3590 VSS.n3589 1.13469
R3589 VSS.n3744 VSS.n3717 1.13469
R3590 VSS.n3744 VSS.n3743 1.13469
R3591 VSS.n3909 VSS.n3908 1.13469
R3592 VSS.n4099 VSS.n4098 1.13469
R3593 VSS.n4445 VSS.n4444 1.13469
R3594 VSS.n3974 VSS.n3973 1.13458
R3595 VSS.n4120 VSS.n4119 1.13458
R3596 VSS.n4310 VSS.n4309 1.13458
R3597 VSS.n4445 VSS.n4371 1.13458
R3598 VSS.n4452 VSS.n4451 1.13458
R3599 VSS.n4348 VSS.n4339 1.13458
R3600 VSS.n3564 VSS.n3554 1.13458
R3601 VSS.n3589 VSS.n3588 1.13458
R3602 VSS.n3487 VSS.n3486 1.13458
R3603 VSS.n3164 VSS.n3086 1.13458
R3604 VSS.n3185 VSS.n3079 1.13458
R3605 VSS.n3128 VSS.n3127 1.13458
R3606 VSS.n4638 VSS.n4637 1.13458
R3607 VSS.n3909 VSS.n3883 1.13458
R3608 VSS.n3771 VSS.n2809 1.13458
R3609 VSS.n4947 VSS.n4946 1.13458
R3610 VSS.n4976 VSS.n4848 1.13458
R3611 VSS.n4870 VSS.n4866 1.13458
R3612 VSS.n4802 VSS.n4801 1.13458
R3613 VSS.n4833 VSS.n4832 1.13458
R3614 VSS.n694 VSS.n427 1.13458
R3615 VSS.n2724 VSS.n2723 1.13458
R3616 VSS.n574 VSS.n569 1.13458
R3617 VSS.n241 VSS.n162 1.13458
R3618 VSS.n217 VSS.n182 1.13458
R3619 VSS.n215 VSS.n214 1.13458
R3620 VSS.n242 VSS.n142 1.13458
R3621 VSS.n264 VSS.n263 1.13458
R3622 VSS.n2523 VSS.n2522 1.13458
R3623 VSS.n637 VSS.n636 1.13458
R3624 VSS.n2516 VSS.n638 1.13458
R3625 VSS.n838 VSS.n644 1.13458
R3626 VSS.n837 VSS.n650 1.13458
R3627 VSS.n789 VSS.n784 1.13458
R3628 VSS.n4760 VSS.n4759 1.13458
R3629 VSS.n4688 VSS.n4687 1.13458
R3630 VSS.n4647 VSS.n4646 1.13458
R3631 VSS.n4638 VSS.n2887 1.13458
R3632 VSS.n4587 VSS.n2888 1.13458
R3633 VSS.n3440 VSS.n3351 1.13458
R3634 VSS.n3487 VSS.n3352 1.13458
R3635 VSS.n3943 VSS.n3942 1.13458
R3636 VSS.n1620 VSS.n1619 1.10395
R3637 VSS.n2558 VSS.n2557 1.10395
R3638 VSS.n4750 VSS.n4749 1.10395
R3639 VSS.n3177 VSS.n3176 1.10395
R3640 VSS.n255 VSS.n252 1.10395
R3641 VSS.n97 VSS.n93 1.08525
R3642 VSS.n2785 VSS.n2783 1.0798
R3643 VSS.n2790 VSS.n2788 1.0798
R3644 VSS.n3830 VSS.n3828 1.0798
R3645 VSS.n3296 VSS.n3294 1.0798
R3646 VSS.n1017 VSS.n1016 1.06282
R3647 VSS.n3056 VSS.n3052 1.04968
R3648 VSS.n4940 VSS.n4936 1.04968
R3649 VSS.n1492 VSS.n1488 1.04968
R3650 VSS.n4233 VSS.n4229 1.04968
R3651 VSS.n74 VSS.n68 1.04225
R3652 VSS.n2375 VSS.n2374 1.04225
R3653 VSS.n1550 VSS.n1548 1.04225
R3654 VSS.n2502 VSS.n2501 1.04225
R3655 VSS.n3449 VSS.n3445 0.970197
R3656 VSS.n1073 VSS.n1051 0.970197
R3657 VSS.n1794 VSS.n946 0.970197
R3658 VSS.n4594 VSS.n4593 0.969987
R3659 VSS.n4597 VSS.n4596 0.901908
R3660 VSS.n486 VSS.n482 0.901908
R3661 VSS.n2486 VSS.n2483 0.883259
R3662 VSS.n1156 VSS.n1147 0.883259
R3663 VSS.n2717 VSS.n2716 0.883259
R3664 VSS.n3244 VSS.n3241 0.883259
R3665 VSS.n2973 VSS.n2969 0.883259
R3666 VSS.n5057 VSS.n5056 0.883259
R3667 VSS.n1938 VSS.n1937 0.853
R3668 VSS.n1889 VSS.n1888 0.853
R3669 VSS.n1256 VSS.n1255 0.853
R3670 VSS.n1007 VSS.n1006 0.853
R3671 VSS.n887 VSS.n886 0.853
R3672 VSS.n2374 VSS.n2373 0.853
R3673 VSS.n3972 VSS.n3971 0.853
R3674 VSS.n4118 VSS.n4117 0.853
R3675 VSS.n4308 VSS.n4307 0.853
R3676 VSS.n1485 VSS.n1466 0.853
R3677 VSS.n4370 VSS.n4369 0.853
R3678 VSS.n3210 VSS.n3209 0.853
R3679 VSS.n4390 VSS.n3261 0.853
R3680 VSS.n4450 VSS.n4449 0.853
R3681 VSS.n135 VSS.n134 0.853
R3682 VSS.n116 VSS.n115 0.853
R3683 VSS.n68 VSS.n36 0.853
R3684 VSS.n1441 VSS.n1440 0.853
R3685 VSS.n1041 VSS.n1040 0.853
R3686 VSS.n1015 VSS.n1013 0.853
R3687 VSS.n1195 VSS.n1194 0.853
R3688 VSS.n1463 VSS.n1462 0.853
R3689 VSS.n1518 VSS.n1473 0.853
R3690 VSS.n2035 VSS.n2034 0.853
R3691 VSS.n1963 VSS.n1962 0.853
R3692 VSS.n1912 VSS.n1911 0.853
R3693 VSS.n29 VSS.n28 0.853
R3694 VSS.n54 VSS.n33 0.853
R3695 VSS.n4512 VSS.n4511 0.853
R3696 VSS.n4552 VSS.n4551 0.853
R3697 VSS.n3236 VSS.n3235 0.853
R3698 VSS.n4484 VSS.n4483 0.853
R3699 VSS.n3258 VSS.n3257 0.853
R3700 VSS.n4338 VSS.n4337 0.853
R3701 VSS.n4213 VSS.n4212 0.853
R3702 VSS.n3553 VSS.n3552 0.853
R3703 VSS.n3587 VSS.n3586 0.853
R3704 VSS.n3485 VSS.n3484 0.853
R3705 VSS.n3085 VSS.n3084 0.853
R3706 VSS.n3078 VSS.n3077 0.853
R3707 VSS.n3130 VSS.n3129 0.853
R3708 VSS.n4636 VSS.n4635 0.853
R3709 VSS.n3716 VSS.n3715 0.853
R3710 VSS.n3742 VSS.n3741 0.853
R3711 VSS.n3907 VSS.n3906 0.853
R3712 VSS.n3882 VSS.n3881 0.853
R3713 VSS.n3773 VSS.n3772 0.853
R3714 VSS.n1864 VSS.n1863 0.853
R3715 VSS.n1975 VSS.n1973 0.853
R3716 VSS.n1798 VSS.n1797 0.853
R3717 VSS.n1615 VSS.n1614 0.853
R3718 VSS.n1168 VSS.n1167 0.853
R3719 VSS.n1092 VSS.n1091 0.853
R3720 VSS.n4945 VSS.n4944 0.853
R3721 VSS.n4847 VSS.n4846 0.853
R3722 VSS.n4865 VSS.n4864 0.853
R3723 VSS.n4800 VSS.n4799 0.853
R3724 VSS.n4831 VSS.n4830 0.853
R3725 VSS.n696 VSS.n695 0.853
R3726 VSS.n2722 VSS.n2721 0.853
R3727 VSS.n568 VSS.n567 0.853
R3728 VSS.n355 VSS.n354 0.853
R3729 VSS.n333 VSS.n332 0.853
R3730 VSS.n425 VSS.n424 0.853
R3731 VSS.n382 VSS.n381 0.853
R3732 VSS.n309 VSS.n274 0.853
R3733 VSS.n161 VSS.n160 0.853
R3734 VSS.n181 VSS.n180 0.853
R3735 VSS.n213 VSS.n212 0.853
R3736 VSS.n141 VSS.n140 0.853
R3737 VSS.n262 VSS.n261 0.853
R3738 VSS.n2525 VSS.n2524 0.853
R3739 VSS.n635 VSS.n634 0.853
R3740 VSS.n2145 VSS.n2144 0.853
R3741 VSS.n643 VSS.n642 0.853
R3742 VSS.n649 VSS.n648 0.853
R3743 VSS.n783 VSS.n782 0.853
R3744 VSS.n4903 VSS.n4902 0.853
R3745 VSS.n3011 VSS.n3010 0.853
R3746 VSS.n2960 VSS.n2959 0.853
R3747 VSS.n3072 VSS.n3071 0.853
R3748 VSS.n3073 VSS.n3072 0.853
R3749 VSS.n2961 VSS.n2960 0.853
R3750 VSS.n3012 VSS.n3011 0.853
R3751 VSS.n3035 VSS.n3034 0.853
R3752 VSS.n2985 VSS.n2984 0.853
R3753 VSS.n4902 VSS.n426 0.853
R3754 VSS.n2913 VSS.n2912 0.853
R3755 VSS.n2938 VSS.n2937 0.853
R3756 VSS.n5021 VSS.n274 0.853
R3757 VSS.n4990 VSS.n382 0.853
R3758 VSS.n4987 VSS.n386 0.853
R3759 VSS.n4984 VSS.n425 0.853
R3760 VSS.n5018 VSS.n333 0.853
R3761 VSS.n4993 VSS.n355 0.853
R3762 VSS.n5015 VSS.n5014 0.853
R3763 VSS.n4758 VSS.n4757 0.853
R3764 VSS.n4691 VSS.n4689 0.853
R3765 VSS.n2757 VSS.n2756 0.853
R3766 VSS.n4649 VSS.n4648 0.853
R3767 VSS.n2886 VSS.n2885 0.853
R3768 VSS.n4005 VSS.n4004 0.853
R3769 VSS.n3442 VSS.n3441 0.853
R3770 VSS.n4685 VSS.n4683 0.853
R3771 VSS.n3421 VSS.n3420 0.853
R3772 VSS.n3183 VSS.n3182 0.853
R3773 VSS.n3161 VSS.n3160 0.853
R3774 VSS.n3109 VSS.n3108 0.853
R3775 VSS.n3034 VSS.n3033 0.853
R3776 VSS.n2984 VSS.n2983 0.853
R3777 VSS.n4952 VSS.n4951 0.853
R3778 VSS.n5014 VSS.n5013 0.853
R3779 VSS.n4974 VSS.n4973 0.853
R3780 VSS.n2912 VSS.n2911 0.853
R3781 VSS.n2937 VSS.n2936 0.853
R3782 VSS.n238 VSS.n237 0.853
R3783 VSS.n4188 VSS.n4186 0.853
R3784 VSS.n4189 VSS.n4188 0.853
R3785 VSS.n4214 VSS.n4213 0.853
R3786 VSS.n4221 VSS.n4220 0.853
R3787 VSS.n4226 VSS.n4225 0.853
R3788 VSS.n4459 VSS.n3261 0.853
R3789 VSS.n4491 VSS.n3210 0.853
R3790 VSS.n4488 VSS.n3236 0.853
R3791 VSS.n4462 VSS.n3258 0.853
R3792 VSS.n4485 VSS.n4484 0.853
R3793 VSS.n4513 VSS.n4512 0.853
R3794 VSS.n4553 VSS.n4552 0.853
R3795 VSS.n3343 VSS.n3341 0.853
R3796 VSS.n3593 VSS.n3592 0.853
R3797 VSS.n4443 VSS.n4441 0.853
R3798 VSS.n4616 VSS.n4615 0.853
R3799 VSS.n4807 VSS.n4806 0.853
R3800 VSS.n835 VSS.n834 0.853
R3801 VSS.n2503 VSS.n2502 0.853
R3802 VSS.n808 VSS.n807 0.853
R3803 VSS.n4584 VSS.n4583 0.853
R3804 VSS.n4097 VSS.n4096 0.853
R3805 VSS.n3941 VSS.n3940 0.853
R3806 VSS.n1414 VSS.n1412 0.853
R3807 VSS.n1415 VSS.n1414 0.853
R3808 VSS.n1257 VSS.n1256 0.853
R3809 VSS.n1614 VSS.n1612 0.853
R3810 VSS.n1237 VSS.n1235 0.853
R3811 VSS.n1238 VSS.n1237 0.853
R3812 VSS.n1093 VSS.n1092 0.853
R3813 VSS.n1169 VSS.n1168 0.853
R3814 VSS.n1124 VSS.n1122 0.853
R3815 VSS.n1125 VSS.n1124 0.853
R3816 VSS.n1008 VSS.n1007 0.853
R3817 VSS.n1042 VSS.n1041 0.853
R3818 VSS.n1196 VSS.n1195 0.853
R3819 VSS.n1288 VSS.n1286 0.853
R3820 VSS.n1289 VSS.n1288 0.853
R3821 VSS.n1562 VSS.n1470 0.853
R3822 VSS.n1565 VSS.n1466 0.853
R3823 VSS.n1571 VSS.n1441 0.853
R3824 VSS.n1568 VSS.n1463 0.853
R3825 VSS.n1607 VSS.n1419 0.853
R3826 VSS.n1559 VSS.n1473 0.853
R3827 VSS.n1603 VSS.n1601 0.853
R3828 VSS.n1604 VSS.n1603 0.853
R3829 VSS.n888 VSS.n887 0.853
R3830 VSS.n1890 VSS.n1889 0.853
R3831 VSS.n1939 VSS.n1938 0.853
R3832 VSS.n1799 VSS.n1798 0.853
R3833 VSS.n1973 VSS.n1971 0.853
R3834 VSS.n1865 VSS.n1864 0.853
R3835 VSS.n2045 VSS.n2044 0.853
R3836 VSS.n2367 VSS.n2366 0.853
R3837 VSS.n2006 VSS.n2005 0.853
R3838 VSS.n2373 VSS.n2371 0.853
R3839 VSS.n2051 VSS.n2049 0.853
R3840 VSS.n2052 VSS.n2051 0.853
R3841 VSS.n1328 VSS.n1327 0.853
R3842 VSS.n1327 VSS.n921 0.853
R3843 VSS.n1967 VSS.n1963 0.853
R3844 VSS.n1808 VSS.n1807 0.853
R3845 VSS.n1913 VSS.n1912 0.853
R3846 VSS.n30 VSS.n29 0.853
R3847 VSS.n2036 VSS.n2035 0.853
R3848 VSS.n2059 VSS.n2058 0.853
R3849 VSS.n1552 VSS.n1550 0.853
R3850 VSS.n1553 VSS.n1552 0.853
R3851 VSS.n5072 VSS.n116 0.853
R3852 VSS.n5078 VSS.n36 0.853
R3853 VSS.n5081 VSS.n33 0.853
R3854 VSS.n5069 VSS.n135 0.853
R3855 VSS.n5065 VSS.n5063 0.853
R3856 VSS.n5066 VSS.n5065 0.853
R3857 VSS.n90 VSS.n89 0.853
R3858 VSS.n3821 VSS 0.849458
R3859 VSS VSS.n4705 0.846854
R3860 VSS.n1650 VSS 0.835135
R3861 VSS.n3291 VSS.n3266 0.685913
R3862 VSS.n4402 VSS.n4401 0.685913
R3863 VSS.n4224 VSS.n4223 0.685559
R3864 VSS.n4347 VSS.n4346 0.685246
R3865 VSS.n3558 VSS.n3557 0.685246
R3866 VSS.n4842 VSS.n4841 0.685246
R3867 VSS.n4778 VSS.n4777 0.685246
R3868 VSS.n4764 VSS.n4763 0.685246
R3869 VSS.n186 VSS.n185 0.685246
R3870 VSS.n3492 VSS.n3491 0.685246
R3871 VSS.n571 VSS.n570 0.682731
R3872 VSS.n2519 VSS.n2518 0.682731
R3873 VSS.n2093 VSS.n2092 0.682731
R3874 VSS.n2101 VSS.n2100 0.682731
R3875 VSS.n3360 VSS.n3359 0.682731
R3876 VSS.n4219 VSS.n4218 0.682471
R3877 VSS.n1418 VSS.n1417 0.682471
R3878 VSS.n1469 VSS.n1468 0.682471
R3879 VSS.n2057 VSS.n2056 0.682471
R3880 VSS.n1806 VSS.n1805 0.682471
R3881 VSS.n2004 VSS.n2003 0.682471
R3882 VSS.n2043 VSS.n2042 0.682471
R3883 VSS.n2365 VSS.n2364 0.682471
R3884 VSS.n493 VSS.n492 0.682471
R3885 VSS.n385 VSS.n384 0.682471
R3886 VSS.n1011 VSS.n1010 0.680783
R3887 VSS.n2691 VSS 0.664562
R3888 VSS.n4106 VSS.n4103 0.662569
R3889 VSS.n3924 VSS.n3921 0.662569
R3890 VSS.n4020 VSS.n4019 0.662569
R3891 VSS.n444 VSS.n443 0.662569
R3892 VSS.n4815 VSS.n4814 0.662569
R3893 VSS.n737 VSS.n736 0.662569
R3894 VSS.n2471 VSS.n2470 0.662569
R3895 VSS.n1932 VSS.n1929 0.662569
R3896 VSS.n3902 VSS.n3901 0.662569
R3897 VSS.n3872 VSS.n3866 0.662569
R3898 VSS.n4660 VSS.n4654 0.662569
R3899 VSS.n1162 VSS.n1161 0.662569
R3900 VSS.n1856 VSS.n1855 0.662569
R3901 VSS.n597 VSS.n596 0.662569
R3902 VSS.n2734 VSS.n2733 0.662569
R3903 VSS.n2815 VSS.n2812 0.662569
R3904 VSS.n4201 VSS.n4198 0.662569
R3905 VSS.n3228 VSS.n3224 0.662569
R3906 VSS.n3155 VSS.n3154 0.662569
R3907 VSS.n3025 VSS.n3022 0.662569
R3908 VSS.n4963 VSS.n4960 0.662569
R3909 VSS.n303 VSS.n300 0.662569
R3910 VSS.n201 VSS.n198 0.662569
R3911 VSS.n149 VSS.n146 0.662569
R3912 VSS.n48 VSS.n45 0.662569
R3913 VSS.n2018 VSS.n2014 0.662569
R3914 VSS.n1434 VSS.n1430 0.662569
R3915 VSS.n1231 VSS.n1220 0.627951
R3916 VSS.n2157 VSS.n2148 0.627951
R3917 VSS.n3712 VSS.n3711 0.591646
R3918 VSS.n802 VSS.n801 0.441879
R3919 VSS.n856 VSS.n855 0.441879
R3920 VSS.n1778 VSS.n950 0.441879
R3921 VSS.n1779 VSS.n947 0.441879
R3922 VSS.n938 VSS.n928 0.441879
R3923 VSS.n930 VSS.n929 0.441879
R3924 VSS.n1825 VSS.n1815 0.441879
R3925 VSS.n1817 VSS.n1816 0.441879
R3926 VSS.n1857 VSS.n1844 0.441879
R3927 VSS.n1848 VSS.n1847 0.441879
R3928 VSS.n1839 VSS.n1830 0.441879
R3929 VSS.n916 VSS.n906 0.441879
R3930 VSS.n908 VSS.n907 0.441879
R3931 VSS.n1999 VSS.n1980 0.441879
R3932 VSS.n1991 VSS.n1990 0.441879
R3933 VSS.n3335 VSS.n3331 0.441879
R3934 VSS.n561 VSS.n558 0.441879
R3935 VSS.n519 VSS.n516 0.441879
R3936 VSS.n325 VSS 0.441879
R3937 VSS.n24 VSS.n23 0.441879
R3938 VSS.n1434 VSS.n1433 0.441879
R3939 VSS.n1557 VSS 0.267519
R3940 VSS VSS.n3712 0.258312
R3941 VSS.n608 VSS.n607 0.241385
R3942 VSS.n4735 VSS 0.232271
R3943 VSS.n1775 VSS 0.229667
R3944 VSS VSS.n4662 0.229667
R3945 VSS.n3874 VSS 0.229667
R3946 VSS.n2363 VSS.n2362 0.227062
R3947 VSS.n2464 VSS.n2463 0.22119
R3948 VSS.n875 VSS.n872 0.22119
R3949 VSS.n3737 VSS.n3736 0.22119
R3950 VSS.n3787 VSS.n3786 0.22119
R3951 VSS.n1058 VSS.n1052 0.22119
R3952 VSS.n1072 VSS.n1071 0.22119
R3953 VSS.n1071 VSS.n1070 0.22119
R3954 VSS.n1086 VSS.n1076 0.22119
R3955 VSS.n1078 VSS.n1077 0.22119
R3956 VSS.n1141 VSS.n1131 0.22119
R3957 VSS.n1133 VSS.n1132 0.22119
R3958 VSS.n1163 VSS.n1162 0.22119
R3959 VSS.n1149 VSS.n1148 0.22119
R3960 VSS.n1211 VSS.n1203 0.22119
R3961 VSS.n1222 VSS.n1221 0.22119
R3962 VSS.n972 VSS.n962 0.22119
R3963 VSS.n964 VSS.n963 0.22119
R3964 VSS.n1619 VSS.n1618 0.22119
R3965 VSS.n1641 VSS.n1640 0.22119
R3966 VSS.n1793 VSS.n1792 0.22119
R3967 VSS.n2234 VSS.n2233 0.22119
R3968 VSS.n2233 VSS.n2078 0.22119
R3969 VSS.n2219 VSS.n2218 0.22119
R3970 VSS.n2218 VSS.n2211 0.22119
R3971 VSS.n2205 VSS.n2204 0.22119
R3972 VSS.n2204 VSS.n2197 0.22119
R3973 VSS.n2191 VSS.n2190 0.22119
R3974 VSS.n2190 VSS.n2183 0.22119
R3975 VSS.n2174 VSS.n2173 0.22119
R3976 VSS.n2173 VSS.n2166 0.22119
R3977 VSS.n2137 VSS.n2136 0.22119
R3978 VSS.n2136 VSS.n2129 0.22119
R3979 VSS.n2123 VSS.n2122 0.22119
R3980 VSS.n2122 VSS.n2115 0.22119
R3981 VSS.n623 VSS.n622 0.22119
R3982 VSS.n2571 VSS.n2569 0.22119
R3983 VSS.n2571 VSS.n2570 0.22119
R3984 VSS.n2596 VSS.n2595 0.22119
R3985 VSS.n2595 VSS.n2588 0.22119
R3986 VSS.n2610 VSS.n2609 0.22119
R3987 VSS.n2609 VSS.n2602 0.22119
R3988 VSS.n2627 VSS.n2626 0.22119
R3989 VSS.n2626 VSS.n2619 0.22119
R3990 VSS.n2641 VSS.n2640 0.22119
R3991 VSS.n2640 VSS.n2633 0.22119
R3992 VSS.n2668 VSS.n2667 0.22119
R3993 VSS.n2667 VSS.n2660 0.22119
R3994 VSS.n2688 VSS.n2687 0.22119
R3995 VSS.n2687 VSS.n2680 0.22119
R3996 VSS.n2753 VSS.n2752 0.22119
R3997 VSS.n3631 VSS.n3626 0.22119
R3998 VSS.n3430 VSS.n3366 0.22119
R3999 VSS VSS.n2236 0.208833
R4000 VSS.n2566 VSS 0.208833
R4001 VSS.n2711 VSS.n2691 0.185396
R4002 VSS.n2651 VSS.n2648 0.175241
R4003 VSS.n2155 VSS.n2152 0.175241
R4004 VSS VSS.n3493 0.172375
R4005 VSS.n2545 VSS.n2540 0.120292
R4006 VSS.n2547 VSS.n2545 0.120292
R4007 VSS.n2548 VSS.n2547 0.120292
R4008 VSS.n2565 VSS.n2548 0.120292
R4009 VSS.n4754 VSS.n4752 0.120292
R4010 VSS.n4752 VSS.n2772 0.120292
R4011 VSS.n4734 VSS.n4733 0.120292
R4012 VSS.n4733 VSS.n4729 0.120292
R4013 VSS.n4729 VSS.n4725 0.120292
R4014 VSS.n4725 VSS.n4718 0.120292
R4015 VSS.n4718 VSS.n4714 0.120292
R4016 VSS.n4714 VSS.n4713 0.120292
R4017 VSS.n4713 VSS.n4709 0.120292
R4018 VSS.n4705 VSS.n4698 0.120292
R4019 VSS.n4698 VSS.n4694 0.120292
R4020 VSS.n4679 VSS.n4675 0.120292
R4021 VSS.n4675 VSS.n4663 0.120292
R4022 VSS.n3789 VSS.n3780 0.120292
R4023 VSS.n3791 VSS.n3789 0.120292
R4024 VSS.n3811 VSS.n3791 0.120292
R4025 VSS.n3825 VSS.n3821 0.120292
R4026 VSS.n3831 VSS.n3825 0.120292
R4027 VSS.n3835 VSS.n3831 0.120292
R4028 VSS.n3842 VSS.n3835 0.120292
R4029 VSS.n3846 VSS.n3842 0.120292
R4030 VSS.n3850 VSS.n3846 0.120292
R4031 VSS.n3851 VSS.n3850 0.120292
R4032 VSS.n3851 VSS.n3750 0.120292
R4033 VSS.n3711 VSS.n3698 0.120292
R4034 VSS.n3698 VSS.n3694 0.120292
R4035 VSS.n3694 VSS.n3693 0.120292
R4036 VSS.n3693 VSS.n3689 0.120292
R4037 VSS.n3689 VSS.n3682 0.120292
R4038 VSS.n3682 VSS.n3678 0.120292
R4039 VSS.n3678 VSS.n3674 0.120292
R4040 VSS.n3674 VSS.n3673 0.120292
R4041 VSS.n509 VSS.n504 0.120292
R4042 VSS.n556 VSS.n550 0.120292
R4043 VSS.n550 VSS.n544 0.120292
R4044 VSS.n544 VSS.n540 0.120292
R4045 VSS.n540 VSS.n534 0.120292
R4046 VSS.n534 VSS.n530 0.120292
R4047 VSS.n530 VSS.n524 0.120292
R4048 VSS.n524 VSS.n520 0.120292
R4049 VSS.n520 VSS.n514 0.120292
R4050 VSS.n3377 VSS.n3373 0.120292
R4051 VSS.n3383 VSS.n3377 0.120292
R4052 VSS.n3388 VSS.n3383 0.120292
R4053 VSS.n3392 VSS.n3388 0.120292
R4054 VSS.n3398 VSS.n3392 0.120292
R4055 VSS.n3402 VSS.n3398 0.120292
R4056 VSS.n3408 VSS.n3402 0.120292
R4057 VSS.n3477 VSS.n3471 0.120292
R4058 VSS.n3466 VSS.n3460 0.120292
R4059 VSS.n3508 VSS.n3503 0.120292
R4060 VSS.n3512 VSS.n3508 0.120292
R4061 VSS.n3518 VSS.n3512 0.120292
R4062 VSS.n3522 VSS.n3518 0.120292
R4063 VSS.n3528 VSS.n3522 0.120292
R4064 VSS.n3534 VSS.n3528 0.120292
R4065 VSS.n3605 VSS.n3599 0.120292
R4066 VSS.n3616 VSS.n3610 0.120292
R4067 VSS.n3620 VSS.n3616 0.120292
R4068 VSS.n3621 VSS.n3620 0.120292
R4069 VSS.n3633 VSS.n3632 0.120292
R4070 VSS.n3639 VSS.n3633 0.120292
R4071 VSS.n3643 VSS.n3639 0.120292
R4072 VSS.n3649 VSS.n3643 0.120292
R4073 VSS.n3650 VSS.n3649 0.120292
R4074 VSS.n3663 VSS.n3657 0.120292
R4075 VSS.n3664 VSS.n3663 0.120292
R4076 VSS.n1037 VSS.n1033 0.120292
R4077 VSS.n1182 VSS.n1178 0.120292
R4078 VSS.n1282 VSS.n1278 0.120292
R4079 VSS.n1585 VSS.n1581 0.120292
R4080 VSS.n1503 VSS.n1499 0.120292
R4081 VSS.n1513 VSS.n1510 0.120292
R4082 VSS.n1546 VSS.n1541 0.120292
R4083 VSS.n2030 VSS.n2026 0.120292
R4084 VSS.n10 VSS.n6 0.120292
R4085 VSS.n64 VSS.n60 0.120292
R4086 VSS.n83 VSS.n79 0.120292
R4087 VSS.n298 VSS.n294 0.120292
R4088 VSS.n318 VSS.n317 0.120292
R4089 VSS.n377 VSS.n373 0.120292
R4090 VSS.n398 VSS.n393 0.120292
R4091 VSS.n413 VSS.n409 0.120292
R4092 VSS.n4932 VSS.n4928 0.120292
R4093 VSS.n4923 VSS.n4917 0.120292
R4094 VSS.n3067 VSS.n3063 0.120292
R4095 VSS.n3144 VSS.n3115 0.120292
R4096 VSS.n4403 VSS.n4398 0.120292
R4097 VSS.n4413 VSS.n4374 0.120292
R4098 VSS.n4174 VSS.n4170 0.120292
R4099 VSS.n4152 VSS.n4148 0.120292
R4100 VSS.n4244 VSS.n4240 0.120292
R4101 VSS.n4250 VSS.n4244 0.120292
R4102 VSS.n4251 VSS.n4250 0.120292
R4103 VSS.n1003 VSS.n1002 0.120292
R4104 VSS.n1108 VSS.n1102 0.120292
R4105 VSS.n1409 VSS.n1405 0.120292
R4106 VSS.n1405 VSS.n1401 0.120292
R4107 VSS.n1401 VSS.n1397 0.120292
R4108 VSS.n1397 VSS.n1393 0.120292
R4109 VSS.n1393 VSS.n1388 0.120292
R4110 VSS.n1388 VSS.n1384 0.120292
R4111 VSS.n1384 VSS.n1380 0.120292
R4112 VSS.n1380 VSS.n1376 0.120292
R4113 VSS.n1376 VSS.n1370 0.120292
R4114 VSS.n1370 VSS.n1366 0.120292
R4115 VSS.n1366 VSS.n1362 0.120292
R4116 VSS.n1362 VSS.n1358 0.120292
R4117 VSS.n1358 VSS.n1357 0.120292
R4118 VSS.n1357 VSS.n1353 0.120292
R4119 VSS.n1353 VSS.n1309 0.120292
R4120 VSS.n1344 VSS.n1343 0.120292
R4121 VSS.n1321 VSS.n1317 0.120292
R4122 VSS.n2384 VSS.n2380 0.120292
R4123 VSS.n2390 VSS.n2384 0.120292
R4124 VSS.n2394 VSS.n2390 0.120292
R4125 VSS.n2398 VSS.n2394 0.120292
R4126 VSS.n2402 VSS.n2398 0.120292
R4127 VSS.n2407 VSS.n2402 0.120292
R4128 VSS.n2411 VSS.n2407 0.120292
R4129 VSS.n2417 VSS.n2411 0.120292
R4130 VSS.n2418 VSS.n2417 0.120292
R4131 VSS.n2430 VSS.n2424 0.120292
R4132 VSS.n2434 VSS.n2430 0.120292
R4133 VSS.n2438 VSS.n2434 0.120292
R4134 VSS.n2444 VSS.n2438 0.120292
R4135 VSS.n2448 VSS.n2444 0.120292
R4136 VSS.n2452 VSS.n2448 0.120292
R4137 VSS.n2456 VSS.n2452 0.120292
R4138 VSS.n2499 VSS.n2495 0.120292
R4139 VSS.n778 VSS.n773 0.120292
R4140 VSS.n773 VSS.n769 0.120292
R4141 VSS.n769 VSS.n768 0.120292
R4142 VSS.n765 VSS.n764 0.120292
R4143 VSS.n764 VSS.n763 0.120292
R4144 VSS.n763 VSS.n759 0.120292
R4145 VSS.n759 VSS.n755 0.120292
R4146 VSS.n755 VSS.n754 0.120292
R4147 VSS.n754 VSS.n750 0.120292
R4148 VSS.n750 VSS.n746 0.120292
R4149 VSS.n746 VSS.n742 0.120292
R4150 VSS.n742 VSS.n738 0.120292
R4151 VSS.n738 VSS.n732 0.120292
R4152 VSS.n732 VSS.n728 0.120292
R4153 VSS.n728 VSS.n724 0.120292
R4154 VSS.n724 VSS.n720 0.120292
R4155 VSS.n720 VSS.n716 0.120292
R4156 VSS.n716 VSS.n711 0.120292
R4157 VSS.n706 VSS.n702 0.120292
R4158 VSS.n4823 VSS.n4813 0.120292
R4159 VSS.n4824 VSS.n4823 0.120292
R4160 VSS.n476 VSS.n470 0.120292
R4161 VSS.n470 VSS.n466 0.120292
R4162 VSS.n466 VSS.n462 0.120292
R4163 VSS.n462 VSS.n461 0.120292
R4164 VSS.n461 VSS.n457 0.120292
R4165 VSS.n457 VSS.n453 0.120292
R4166 VSS.n453 VSS.n449 0.120292
R4167 VSS.n449 VSS.n445 0.120292
R4168 VSS.n445 VSS.n439 0.120292
R4169 VSS.n2838 VSS.n2834 0.120292
R4170 VSS.n2842 VSS.n2838 0.120292
R4171 VSS.n2847 VSS.n2842 0.120292
R4172 VSS.n2851 VSS.n2847 0.120292
R4173 VSS.n2855 VSS.n2851 0.120292
R4174 VSS.n2859 VSS.n2855 0.120292
R4175 VSS.n2865 VSS.n2859 0.120292
R4176 VSS.n2869 VSS.n2865 0.120292
R4177 VSS.n4631 VSS.n4627 0.120292
R4178 VSS.n4627 VSS.n4599 0.120292
R4179 VSS.n4580 VSS.n4576 0.120292
R4180 VSS.n3998 VSS.n3994 0.120292
R4181 VSS.n4015 VSS.n4011 0.120292
R4182 VSS.n4021 VSS.n4015 0.120292
R4183 VSS.n4025 VSS.n4021 0.120292
R4184 VSS.n4029 VSS.n4025 0.120292
R4185 VSS.n4033 VSS.n4029 0.120292
R4186 VSS.n4037 VSS.n4033 0.120292
R4187 VSS.n4042 VSS.n4037 0.120292
R4188 VSS.n4046 VSS.n4042 0.120292
R4189 VSS.n4050 VSS.n4046 0.120292
R4190 VSS.n4054 VSS.n4050 0.120292
R4191 VSS.n4060 VSS.n4054 0.120292
R4192 VSS.n4064 VSS.n4060 0.120292
R4193 VSS.n4068 VSS.n4064 0.120292
R4194 VSS.n4072 VSS.n4068 0.120292
R4195 VSS.n4077 VSS.n4072 0.120292
R4196 VSS.n4081 VSS.n4077 0.120292
R4197 VSS.n4087 VSS.n4081 0.120292
R4198 VSS.n4088 VSS.n4087 0.120292
R4199 VSS.n3989 VSS.n3983 0.120292
R4200 VSS.n3955 VSS.n3949 0.120292
R4201 VSS.n4303 VSS.n4299 0.120292
R4202 VSS.n4299 VSS.n4294 0.120292
R4203 VSS.n4294 VSS.n4290 0.120292
R4204 VSS.n4290 VSS.n4286 0.120292
R4205 VSS.n4286 VSS.n4282 0.120292
R4206 VSS.n4282 VSS.n4276 0.120292
R4207 VSS.n4276 VSS.n4272 0.120292
R4208 VSS.n4272 VSS.n4268 0.120292
R4209 VSS.n4268 VSS.n4264 0.120292
R4210 VSS.n4264 VSS.n4263 0.120292
R4211 VSS.n4263 VSS.n4259 0.120292
R4212 VSS.n4259 VSS.n4258 0.120292
R4213 VSS.n2472 VSS.n2466 0.11899
R4214 VSS.n557 VSS.n556 0.117688
R4215 VSS.n299 VSS.n298 0.116385
R4216 VSS.n3151 VSS.n3150 0.116385
R4217 VSS.n477 VSS.n476 0.116385
R4218 VSS.n5053 VSS.n5052 0.115083
R4219 VSS.n4933 VSS.n4932 0.115083
R4220 VSS.n2482 VSS.n2481 0.115083
R4221 VSS.n4240 VSS.n4236 0.113781
R4222 VSS.n2870 VSS.n2869 0.112479
R4223 VSS.n3956 VSS.n3955 0.111177
R4224 VSS.n4907 VSS.n4906 0.109875
R4225 VSS.n3000 VSS.n2999 0.109875
R4226 VSS.n4428 VSS.n4423 0.109875
R4227 VSS.n820 VSS.n819 0.109875
R4228 VSS.n3478 VSS.n3477 0.108573
R4229 VSS.n1499 VSS.n1495 0.108573
R4230 VSS.n3409 VSS.n3408 0.107271
R4231 VSS.n414 VSS.n413 0.107271
R4232 VSS.n4380 VSS.n4379 0.107271
R4233 VSS.n3756 VSS.n3755 0.105969
R4234 VSS.n3453 VSS.n3452 0.105969
R4235 VSS.n1591 VSS.n1590 0.105969
R4236 VSS.n3931 VSS.n3930 0.105969
R4237 VSS.n2798 VSS.n2797 0.104667
R4238 VSS.n101 VSS.n100 0.104667
R4239 VSS.n1343 VSS.n1337 0.104667
R4240 VSS.n4537 VSS.n4536 0.103365
R4241 VSS.n4327 VSS.n4326 0.103365
R4242 VSS.n860 VSS.n854 0.103365
R4243 VSS.n3875 VSS 0.102083
R4244 VSS.n3542 VSS.n3541 0.102062
R4245 VSS.n5039 VSS.n5038 0.102062
R4246 VSS.n3223 VSS.n3222 0.102062
R4247 VSS.n3309 VSS.n3308 0.10076
R4248 VSS.n281 VSS.n279 0.10076
R4249 VSS.n4890 VSS.n4889 0.10076
R4250 VSS.n2746 VSS.n2745 0.0994583
R4251 VSS.n16 VSS.n15 0.0994583
R4252 VSS.n1667 VSS.n1666 0.0981562
R4253 VSS.n1681 VSS.n1680 0.0981562
R4254 VSS.n1694 VSS.n1693 0.0981562
R4255 VSS.n1708 VSS.n1707 0.0981562
R4256 VSS.n1724 VSS.n1723 0.0981562
R4257 VSS.n1738 VSS.n1737 0.0981562
R4258 VSS.n1752 VSS.n1751 0.0981562
R4259 VSS.n1753 VSS.n951 0.0981562
R4260 VSS.n941 VSS.n940 0.0981562
R4261 VSS.n2340 VSS.n2339 0.0981562
R4262 VSS.n2326 VSS.n2325 0.0981562
R4263 VSS.n2323 VSS.n2322 0.0981562
R4264 VSS.n2309 VSS.n2308 0.0981562
R4265 VSS.n2293 VSS.n2292 0.0981562
R4266 VSS.n2279 VSS.n2278 0.0981562
R4267 VSS.n2265 VSS.n2264 0.0981562
R4268 VSS.n2262 VSS.n2261 0.0981562
R4269 VSS.n2222 VSS.n2221 0.0981562
R4270 VSS.n2208 VSS.n2207 0.0981562
R4271 VSS.n2194 VSS.n2193 0.0981562
R4272 VSS.n2177 VSS.n2176 0.0981562
R4273 VSS.n2163 VSS.n2162 0.0981562
R4274 VSS.n2126 VSS.n2125 0.0981562
R4275 VSS.n2586 VSS.n2585 0.0981562
R4276 VSS.n2599 VSS.n2598 0.0981562
R4277 VSS.n2613 VSS.n2612 0.0981562
R4278 VSS.n2630 VSS.n2629 0.0981562
R4279 VSS.n2644 VSS.n2643 0.0981562
R4280 VSS.n2657 VSS.n2656 0.0981562
R4281 VSS.n2671 VSS.n2670 0.0981562
R4282 VSS.n1027 VSS 0.0981562
R4283 VSS.n4787 VSS.n4786 0.0981562
R4284 VSS.n4652 VSS 0.0975498
R4285 VSS.n2540 VSS.n2532 0.0968542
R4286 VSS VSS.n4734 0.0968542
R4287 VSS.n3730 VSS.n3729 0.0968542
R4288 VSS.n1450 VSS.n1449 0.0968542
R4289 VSS.n1954 VSS.n1953 0.0968542
R4290 VSS.n105 VSS.n43 0.0968542
R4291 VSS.n4429 VSS.n4428 0.0968542
R4292 VSS.n658 VSS.n657 0.0968542
R4293 VSS.n3572 VSS.n3571 0.0955521
R4294 VSS.n1268 VSS.n1267 0.0955521
R4295 VSS.n1528 VSS.n1476 0.0955521
R4296 VSS.n5007 VSS.n5006 0.0955521
R4297 VSS.n2905 VSS.n2904 0.0955521
R4298 VSS.n4180 VSS.n4179 0.0955521
R4299 VSS.n3990 VSS.n3989 0.0955521
R4300 VSS.n1842 VSS.n1841 0.09425
R4301 VSS.n226 VSS.n225 0.09425
R4302 VSS.n342 VSS.n341 0.09425
R4303 VSS.n3102 VSS.n3101 0.09425
R4304 VSS.n1114 VSS.n1113 0.09425
R4305 VSS.n1882 VSS.n1881 0.09425
R4306 VSS.n1529 VSS.n1528 0.0929479
R4307 VSS.n65 VSS.n64 0.0929479
R4308 VSS.n4536 VSS.n4532 0.0929479
R4309 VSS.n861 VSS.n860 0.0929479
R4310 VSS.n2473 VSS.n2472 0.0929479
R4311 VSS.n2002 VSS 0.0916458
R4312 VSS.n1547 VSS.n1546 0.0916458
R4313 VSS.n79 VSS.n75 0.0916458
R4314 VSS.n4524 VSS.n4523 0.0916458
R4315 VSS.n2380 VSS.n2376 0.0916458
R4316 VSS.n2500 VSS.n2499 0.0916458
R4317 VSS.n131 VSS.n130 0.0903438
R4318 VSS.n235 VSS.n234 0.0903438
R4319 VSS.n351 VSS.n350 0.0903438
R4320 VSS.n3095 VSS.n3094 0.0903438
R4321 VSS.n1109 VSS.n1108 0.0903438
R4322 VSS.n1877 VSS.n1876 0.0903438
R4323 VSS.n3583 VSS.n3582 0.0890417
R4324 VSS.n1283 VSS.n1282 0.0890417
R4325 VSS.n2900 VSS.n2899 0.0890417
R4326 VSS.n4175 VSS.n4174 0.0890417
R4327 VSS.n4609 VSS.n4608 0.0890417
R4328 VSS.n600 VSS.n599 0.0877396
R4329 VSS.n3727 VSS.n3726 0.0877396
R4330 VSS.n1459 VSS.n1458 0.0877396
R4331 VSS.n1949 VSS.n1948 0.0877396
R4332 VSS.n3031 VSS.n3030 0.0877396
R4333 VSS.n4438 VSS.n4437 0.0877396
R4334 VSS.n1253 VSS.n1252 0.0877396
R4335 VSS.n779 VSS.n778 0.0877396
R4336 VSS.n1028 VSS.n1027 0.0864375
R4337 VSS.n404 VSS.n403 0.0864375
R4338 VSS.n1004 VSS.n1003 0.0864375
R4339 VSS.n4796 VSS.n4795 0.0864375
R4340 VSS.n1979 VSS.n1978 0.0851354
R4341 VSS.n2737 VSS.n2736 0.0851354
R4342 VSS.n11 VSS.n10 0.0851354
R4343 VSS.n4481 VSS.n4480 0.0851354
R4344 VSS.n3599 VSS.n3595 0.0838333
R4345 VSS.n4906 VSS.n4905 0.0838333
R4346 VSS.n2934 VSS.n2933 0.0838333
R4347 VSS.n3535 VSS.n3534 0.0825312
R4348 VSS.n5052 VSS.n5048 0.0825312
R4349 VSS.n3218 VSS.n3217 0.0825312
R4350 VSS.n1410 VSS.n1409 0.0825312
R4351 VSS.n2712 VSS.n2711 0.0812292
R4352 VSS.n4549 VSS.n4548 0.0812292
R4353 VSS.n4322 VSS.n4321 0.0812292
R4354 VSS.n4209 VSS.n4208 0.0812292
R4355 VSS.n846 VSS.n845 0.0812292
R4356 VSS.n702 VSS.n698 0.0812292
R4357 VSS.n4581 VSS.n4580 0.0812292
R4358 VSS VSS.n1060 0.0799271
R4359 VSS.n1089 VSS.n1088 0.0799271
R4360 VSS.n4694 VSS.n4693 0.0799271
R4361 VSS.n2825 VSS.n2824 0.0799271
R4362 VSS.n3328 VSS.n3327 0.0799271
R4363 VSS.n84 VSS.n83 0.0799271
R4364 VSS.n1322 VSS.n1321 0.0799271
R4365 VSS.n1934 VSS.n1933 0.0799271
R4366 VSS.n3780 VSS.n3775 0.078625
R4367 VSS.n504 VSS.n499 0.078625
R4368 VSS.n3494 VSS.n3347 0.078625
R4369 VSS.n1586 VSS.n1585 0.078625
R4370 VSS.n1900 VSS.n1899 0.078625
R4371 VSS.n3926 VSS.n3925 0.078625
R4372 VSS.n904 VSS.n903 0.0773229
R4373 VSS.n3424 VSS.n3423 0.0773229
R4374 VSS.n209 VSS.n208 0.0773229
R4375 VSS.n399 VSS.n398 0.0773229
R4376 VSS.n4398 VSS.n4392 0.0773229
R4377 VSS.n2087 VSS 0.0760208
R4378 VSS VSS.n583 0.0760208
R4379 VSS.n3432 VSS.n3431 0.0760208
R4380 VSS.n1482 VSS.n1481 0.0760208
R4381 VSS.n2956 VSS.n2955 0.0760208
R4382 VSS.n4304 VSS.n4303 0.0760208
R4383 VSS.n378 VSS.n377 0.0747188
R4384 VSS.n2995 VSS.n2994 0.0747188
R4385 VSS.n4414 VSS.n4413 0.0747188
R4386 VSS.n832 VSS.n831 0.0747188
R4387 VSS.n3879 VSS.n3878 0.0734167
R4388 VSS.n177 VSS.n176 0.0734167
R4389 VSS.n4367 VSS.n4366 0.0734167
R4390 VSS.n3968 VSS.n3967 0.0734167
R4391 VSS.n4755 VSS.n4754 0.0721146
R4392 VSS.n1183 VSS.n1182 0.0721146
R4393 VSS.n3068 VSS.n3067 0.0721146
R4394 VSS.n3199 VSS.n3198 0.0721146
R4395 VSS.n4813 VSS.n4809 0.0721146
R4396 VSS.n2882 VSS.n2881 0.0721146
R4397 VSS.n250 VSS.n249 0.0708125
R4398 VSS.n3172 VSS.n3171 0.0708125
R4399 VSS.n4153 VSS.n4152 0.0708125
R4400 VSS.n5032 VSS.n5031 0.0695104
R4401 VSS.n4877 VSS.n4876 0.0695104
R4402 VSS.n2981 VSS.n2980 0.0695104
R4403 VSS.n3254 VSS.n3253 0.0695104
R4404 VSS.n2495 VSS.n2491 0.0695104
R4405 VSS.n1828 VSS.n1827 0.0682083
R4406 VSS.n4680 VSS.n4679 0.0682083
R4407 VSS.n3892 VSS.n3891 0.0682083
R4408 VSS.n2031 VSS.n2030 0.0682083
R4409 VSS.n60 VSS.n56 0.0682083
R4410 VSS.n157 VSS.n156 0.0682083
R4411 VSS.n317 VSS.n311 0.0682083
R4412 VSS.n4971 VSS.n4970 0.0682083
R4413 VSS.n3145 VSS.n3144 0.0682083
R4414 VSS.n4114 VSS.n4113 0.0682083
R4415 VSS.n510 VSS.n509 0.0669062
R4416 VSS.n1428 VSS.n1427 0.0669062
R4417 VSS.n3063 VSS.n3059 0.0669062
R4418 VSS.n797 VSS.n796 0.0669062
R4419 VSS.n631 VSS.n630 0.0656042
R4420 VSS.n883 VSS.n882 0.0656042
R4421 VSS.n2457 VSS.n2456 0.0656042
R4422 VSS.n1537 VSS.n1536 0.0643021
R4423 VSS.n4861 VSS.n4860 0.0643021
R4424 VSS.n4509 VSS.n4508 0.0643021
R4425 VSS.n4170 VSS.n4166 0.0643021
R4426 VSS.n4632 VSS.n4631 0.0643021
R4427 VSS.n4011 VSS.n4007 0.0643021
R4428 VSS.n4148 VSS.n4144 0.063
R4429 VSS.n3467 VSS.n3466 0.0616979
R4430 VSS.n3606 VSS.n3605 0.0616979
R4431 VSS.n1581 VSS.n1576 0.0616979
R4432 VSS.n1510 VSS.n1504 0.0616979
R4433 VSS.n288 VSS.n287 0.0616979
R4434 VSS.n373 VSS.n369 0.0616979
R4435 VSS.n4924 VSS.n4923 0.0616979
R4436 VSS.n711 VSS.n707 0.0616979
R4437 VSS.n4709 VSS 0.0603958
R4438 VSS VSS.n3811 0.0603958
R4439 VSS.n3431 VSS 0.0603958
R4440 VSS.n3460 VSS 0.0603958
R4441 VSS.n3453 VSS 0.0603958
R4442 VSS.n3494 VSS 0.0603958
R4443 VSS.n3632 VSS 0.0603958
R4444 VSS.n3650 VSS 0.0603958
R4445 VSS.n3657 VSS 0.0603958
R4446 VSS.n3664 VSS 0.0603958
R4447 VSS VSS.n1513 0.0603958
R4448 VSS.n101 VSS 0.0603958
R4449 VSS.n318 VSS 0.0603958
R4450 VSS.n4917 VSS 0.0603958
R4451 VSS VSS.n3115 0.0603958
R4452 VSS.n4403 VSS 0.0603958
R4453 VSS VSS.n4374 0.0603958
R4454 VSS.n4251 VSS 0.0603958
R4455 VSS.n1344 VSS 0.0603958
R4456 VSS.n2418 VSS 0.0603958
R4457 VSS.n2424 VSS 0.0603958
R4458 VSS.n768 VSS 0.0603958
R4459 VSS.n765 VSS 0.0603958
R4460 VSS.n4824 VSS 0.0603958
R4461 VSS VSS.n4599 0.0603958
R4462 VSS.n4088 VSS 0.0603958
R4463 VSS.n4258 VSS 0.0603958
R4464 VSS.n2103 VSS 0.0590938
R4465 VSS VSS.n2690 0.0590938
R4466 VSS.n3471 VSS.n3467 0.0590938
R4467 VSS.n3610 VSS.n3606 0.0590938
R4468 VSS.n1504 VSS.n1503 0.0590938
R4469 VSS.n294 VSS.n288 0.0590938
R4470 VSS.n4928 VSS.n4924 0.0590938
R4471 VSS.n707 VSS.n706 0.0590938
R4472 VSS.n975 VSS.n974 0.0577917
R4473 VSS VSS.n926 0.0577917
R4474 VSS.n4144 VSS.n4143 0.0577917
R4475 VSS.n1541 VSS.n1537 0.0564896
R4476 VSS.n2026 VSS.n2022 0.0564896
R4477 VSS.n4166 VSS.n4165 0.0564896
R4478 VSS.n1609 VSS 0.0560545
R4479 VSS.n1214 VSS.n1213 0.0512812
R4480 VSS.n1144 VSS.n1143 0.047375
R4481 VSS.n2140 VSS.n2139 0.0447708
R4482 VSS.n886 VSS.n870 0.0427297
R4483 VSS.n4511 VSS.n4496 0.0427297
R4484 VSS.n3077 VSS.n3076 0.0427297
R4485 VSS.n4635 VSS.n4590 0.0427297
R4486 VSS.n4864 VSS.n4850 0.0427297
R4487 VSS.n567 VSS.n566 0.0427297
R4488 VSS.n648 VSS.n647 0.0427297
R4489 VSS.n807 VSS.n792 0.0427297
R4490 VSS.n4005 VSS.n4001 0.0427297
R4491 VSS.n1440 VSS.n1423 0.0410405
R4492 VSS.n3160 VSS.n3114 0.0410405
R4493 VSS.n634 VSS.n606 0.0410405
R4494 VSS.n2145 VSS.n2141 0.0410405
R4495 VSS VSS.n2001 0.0408646
R4496 VSS VSS.n1649 0.0395625
R4497 VSS.n5063 VSS.n5062 0.0393514
R4498 VSS.n54 VSS.n52 0.0393514
R4499 VSS.n3906 VSS.n3886 0.0393514
R4500 VSS.n1167 VSS.n1129 0.0393514
R4501 VSS.n4944 VSS.n4943 0.0393514
R4502 VSS.n4973 VSS.n4955 0.0393514
R4503 VSS.n4830 VSS.n4829 0.0393514
R4504 VSS.n160 VSS.n144 0.0393514
R4505 VSS.n2374 VSS.n866 0.0376622
R4506 VSS.n4117 VSS.n4101 0.0376622
R4507 VSS.n68 VSS.n67 0.0376622
R4508 VSS.n1550 VSS.n1549 0.0376622
R4509 VSS.n2034 VSS.n2012 0.0376622
R4510 VSS.n3257 VSS.n3239 0.0376622
R4511 VSS.n309 VSS.n307 0.0376622
R4512 VSS.n642 VSS.n641 0.0376622
R4513 VSS.n2502 VSS.n841 0.0376622
R4514 VSS.n2983 VSS.n2966 0.0376622
R4515 VSS.n4683 VSS.n2810 0.0376622
R4516 VSS.n3560 VSS.n3559 0.0372251
R4517 VSS.n577 VSS.n576 0.0370556
R4518 VSS.n3355 VSS.n3354 0.0368521
R4519 VSS.n2374 VSS.n865 0.035973
R4520 VSS.n134 VSS.n133 0.035973
R4521 VSS.n68 VSS.n66 0.035973
R4522 VSS.n1550 VSS.n1475 0.035973
R4523 VSS.n3084 VSS.n3081 0.035973
R4524 VSS.n3083 VSS.n3082 0.035973
R4525 VSS.n3182 VSS.n3167 0.035973
R4526 VSS.n1235 VSS.n1234 0.035973
R4527 VSS.n354 VSS.n353 0.035973
R4528 VSS.n261 VSS.n260 0.035973
R4529 VSS.n2502 VSS.n840 0.035973
R4530 VSS.n4226 VSS.n4155 0.035973
R4531 VSS.n4602 VSS 0.0356562
R4532 VSS.n1888 VSS.n1870 0.0342838
R4533 VSS.n1872 VSS.n1871 0.0342838
R4534 VSS.n1121 VSS.n1120 0.0342838
R4535 VSS.n3209 VSS.n3194 0.0342838
R4536 VSS.n120 VSS.n119 0.0342838
R4537 VSS.n1194 VSS.n1193 0.0342838
R4538 VSS.n1286 VSS.n1285 0.0342838
R4539 VSS.n3108 VSS.n3088 0.0342838
R4540 VSS.n3090 VSS.n3089 0.0342838
R4541 VSS.n4616 VSS.n4612 0.0342838
R4542 VSS.n337 VSS.n336 0.0342838
R4543 VSS.n220 VSS.n219 0.0342838
R4544 VSS.n237 VSS.n221 0.0342838
R4545 VSS.n3071 VSS.n3040 0.0342838
R4546 VSS.n4757 VSS.n2761 0.0342838
R4547 VSS.n2890 VSS.n2889 0.0334
R4548 VSS.n4995 VSS.n4994 0.0332531
R4549 VSS.n565 VSS.n564 0.0330521
R4550 VSS.n4862 VSS.n4856 0.0330521
R4551 VSS.n3058 VSS.n3057 0.0330521
R4552 VSS.n4510 VSS.n4504 0.0330521
R4553 VSS.n884 VSS.n878 0.0330521
R4554 VSS.n2460 VSS.n2458 0.0330521
R4555 VSS.n806 VSS.n805 0.0330521
R4556 VSS.n4633 VSS.n4598 0.0330521
R4557 VSS.n4006 VSS.n4000 0.0330521
R4558 VSS.n1122 VSS.n1098 0.0325946
R4559 VSS.n3978 VSS.n3977 0.0325946
R4560 VSS.n4369 VSS.n4351 0.0325946
R4561 VSS.n1263 VSS.n1262 0.0325946
R4562 VSS.n1518 VSS.n1515 0.0325946
R4563 VSS.n1517 VSS.n1516 0.0325946
R4564 VSS.n3567 VSS.n3566 0.0325946
R4565 VSS.n3586 VSS.n3585 0.0325946
R4566 VSS.n4611 VSS.n4610 0.0325946
R4567 VSS.n1975 VSS.n1974 0.0325946
R4568 VSS.n4951 VSS.n4950 0.0325946
R4569 VSS.n4807 VSS.n488 0.0325946
R4570 VSS.n5013 VSS.n4998 0.0325946
R4571 VSS.n5000 VSS.n4999 0.0325946
R4572 VSS.n3033 VSS.n3019 0.0325946
R4573 VSS.n2911 VSS.n2893 0.0325946
R4574 VSS.n2895 VSS.n2894 0.0325946
R4575 VSS.n2885 VSS.n2830 0.0325946
R4576 VSS.n4186 VSS.n4158 0.0325946
R4577 VSS.n4160 VSS.n4159 0.0325946
R4578 VSS.n2158 VSS.n2146 0.03175
R4579 VSS.n632 VSS.n628 0.03175
R4580 VSS.n1439 VSS.n1438 0.03175
R4581 VSS.n3159 VSS.n3158 0.03175
R4582 VSS.n1242 VSS.n1241 0.0309054
R4583 VSS.n1255 VSS.n1243 0.0309054
R4584 VSS.n3971 VSS.n3945 0.0309054
R4585 VSS.n4096 VSS.n3976 0.0309054
R4586 VSS.n4373 VSS.n4372 0.0309054
R4587 VSS.n4441 VSS.n4440 0.0309054
R4588 VSS.n4449 VSS.n4448 0.0309054
R4589 VSS.n115 VSS.n39 0.0309054
R4590 VSS.n41 VSS.n40 0.0309054
R4591 VSS.n1445 VSS.n1444 0.0309054
R4592 VSS.n1462 VSS.n1461 0.0309054
R4593 VSS.n1961 VSS.n1960 0.0309054
R4594 VSS.n3715 VSS.n3268 0.0309054
R4595 VSS.n3721 VSS.n3720 0.0309054
R4596 VSS.n3881 VSS.n3746 0.0309054
R4597 VSS.n1862 VSS.n1861 0.0309054
R4598 VSS.n919 VSS.n918 0.0309054
R4599 VSS.n4799 VSS.n4798 0.0309054
R4600 VSS.n180 VSS.n164 0.0309054
R4601 VSS.n2525 VSS.n601 0.0309054
R4602 VSS.n603 VSS.n602 0.0309054
R4603 VSS.n653 VSS.n652 0.0309054
R4604 VSS.n782 VSS.n781 0.0309054
R4605 VSS.n3018 VSS.n3017 0.0309054
R4606 VSS.n3010 VSS.n3009 0.0309054
R4607 VSS.n1166 VSS.n1165 0.0304479
R4608 VSS.n3905 VSS.n3904 0.0304479
R4609 VSS.n55 VSS.n51 0.0304479
R4610 VSS.n5061 VSS.n5060 0.0304479
R4611 VSS.n158 VSS.n152 0.0304479
R4612 VSS.n4972 VSS.n4966 0.0304479
R4613 VSS.n4942 VSS.n4941 0.0304479
R4614 VSS.n4828 VSS.n4827 0.0304479
R4615 VSS.n4461 VSS.n4460 0.0303156
R4616 VSS.n1573 VSS.n1572 0.0295812
R4617 VSS.n5077 VSS.n5076 0.0292875
R4618 VSS.n1006 VSS.n989 0.0292162
R4619 VSS.n1485 VSS.n1484 0.0292162
R4620 VSS.n1040 VSS.n982 0.0292162
R4621 VSS.n1015 VSS.n1014 0.0292162
R4622 VSS.n1962 VSS.n1942 0.0292162
R4623 VSS.n3484 VSS.n3483 0.0292162
R4624 VSS.n3741 VSS.n3719 0.0292162
R4625 VSS.n1863 VSS.n1813 0.0292162
R4626 VSS.n4846 VSS.n4845 0.0292162
R4627 VSS.n4782 VSS.n4781 0.0292162
R4628 VSS.n424 VSS.n423 0.0292162
R4629 VSS.n381 VSS.n358 0.0292162
R4630 VSS.n834 VSS.n812 0.0292162
R4631 VSS.n4681 VSS.n2818 0.0291458
R4632 VSS.n1514 VSS 0.0291458
R4633 VSS.n1548 VSS.n1547 0.0291458
R4634 VSS.n2032 VSS.n2021 0.0291458
R4635 VSS.n75 VSS.n74 0.0291458
R4636 VSS.n310 VSS.n306 0.0291458
R4637 VSS.n2982 VSS.n2976 0.0291458
R4638 VSS.n3255 VSS.n3247 0.0291458
R4639 VSS.n2376 VSS.n2375 0.0291458
R4640 VSS.n2501 VSS.n2500 0.0291458
R4641 VSS.n2490 VSS.n2489 0.0291458
R4642 VSS VSS.n3979 0.0291458
R4643 VSS.n4115 VSS.n4109 0.0291458
R4644 VSS.n1564 VSS.n1563 0.0289937
R4645 VSS.n1233 VSS.n1232 0.0278438
R4646 VSS.n1548 VSS.n1529 0.0278438
R4647 VSS.n74 VSS.n65 0.0278438
R4648 VSS VSS.n42 0.0278438
R4649 VSS.n132 VSS.n131 0.0278438
R4650 VSS.n259 VSS.n258 0.0278438
R4651 VSS.n352 VSS.n351 0.0278438
R4652 VSS.n3181 VSS.n3180 0.0278438
R4653 VSS.n4525 VSS.n4524 0.0278438
R4654 VSS.n4532 VSS.n4531 0.0278438
R4655 VSS.n4234 VSS.n4227 0.0278438
R4656 VSS.n2375 VSS.n861 0.0278438
R4657 VSS.n2501 VSS.n2473 0.0278438
R4658 VSS.n4307 VSS.n4122 0.027527
R4659 VSS.n4483 VSS.n4468 0.027527
R4660 VSS.n3593 VSS.n3319 0.027527
R4661 VSS.n1615 VSS.n977 0.027527
R4662 VSS.n212 VSS.n194 0.027527
R4663 VSS.n2959 VSS.n2943 0.027527
R4664 VSS.n1567 VSS.n1566 0.027525
R4665 VSS.n5068 VSS.n5067 0.0266437
R4666 VSS.n4756 VSS.n2771 0.0265417
R4667 VSS.n1192 VSS.n1191 0.0265417
R4668 VSS.n1284 VSS.n1283 0.0265417
R4669 VSS.n125 VSS.n121 0.0265417
R4670 VSS.n230 VSS.n226 0.0265417
R4671 VSS.n236 VSS.n235 0.0265417
R4672 VSS.n346 VSS.n342 0.0265417
R4673 VSS.n3069 VSS.n3048 0.0265417
R4674 VSS.n3107 VSS.n3095 0.0265417
R4675 VSS.n3106 VSS.n3102 0.0265417
R4676 VSS.n3208 VSS.n3207 0.0265417
R4677 VSS.n1118 VSS.n1114 0.0265417
R4678 VSS.n1887 VSS.n1877 0.0265417
R4679 VSS.n1886 VSS.n1882 0.0265417
R4680 VSS.n4617 VSS.n4609 0.0265417
R4681 VSS.n5080 VSS 0.0264969
R4682 VSS.n5083 VSS.n5082 0.0259094
R4683 VSS.n4390 VSS.n4388 0.0258378
R4684 VSS.n90 VSS.n86 0.0258378
R4685 VSS.n1601 VSS.n1600 0.0258378
R4686 VSS.n1911 VSS.n1910 0.0258378
R4687 VSS.n28 VSS.n2 0.0258378
R4688 VSS.n3341 VSS.n3340 0.0258378
R4689 VSS.n2756 VSS.n2726 0.0258378
R4690 VSS.n2936 VSS.n2919 0.0258378
R4691 VSS.n4903 VSS.n4898 0.0258378
R4692 VSS.n3442 VSS.n3437 0.0258378
R4693 VSS.n3421 VSS.n3417 0.0258378
R4694 VSS.n3940 VSS.n3919 0.0258378
R4695 VSS.n1412 VSS.n1295 0.0258378
R4696 VSS.n1570 VSS.n1569 0.0254688
R4697 VSS.n3578 VSS.n3572 0.0252396
R4698 VSS.n3584 VSS.n3583 0.0252396
R4699 VSS.n1274 VSS.n1268 0.0252396
R4700 VSS.n1519 VSS.n1514 0.0252396
R4701 VSS.n5012 VSS.n5001 0.0252396
R4702 VSS.n5011 VSS.n5007 0.0252396
R4703 VSS.n4884 VSS.n4882 0.0252396
R4704 VSS.n2910 VSS.n2900 0.0252396
R4705 VSS.n2909 VSS.n2905 0.0252396
R4706 VSS.n3032 VSS.n3031 0.0252396
R4707 VSS.n4368 VSS.n4360 0.0252396
R4708 VSS.n4185 VSS.n4175 0.0252396
R4709 VSS.n4184 VSS.n4180 0.0252396
R4710 VSS.n1119 VSS.n1109 0.0252396
R4711 VSS.n4808 VSS.n487 0.0252396
R4712 VSS.n2883 VSS.n2877 0.0252396
R4713 VSS.n4618 VSS.n4602 0.0252396
R4714 VSS.n4094 VSS.n3990 0.0252396
R4715 VSS.n5020 VSS.n5019 0.0248813
R4716 VSS.n1561 VSS.n1560 0.0248813
R4717 VSS.n4551 VSS.n4519 0.0241486
R4718 VSS.n3235 VSS.n3213 0.0241486
R4719 VSS.n3552 VSS.n3346 0.0241486
R4720 VSS.n3773 VSS.n3768 0.0241486
R4721 VSS.n1091 VSS.n1048 0.0241486
R4722 VSS.n696 VSS.n692 0.0241486
R4723 VSS.n2721 VSS.n2720 0.0241486
R4724 VSS.n332 VSS.n277 0.0241486
R4725 VSS.n4691 VSS.n4690 0.0241486
R4726 VSS.n2526 VSS.n600 0.0239375
R4727 VSS.n2532 VSS.n2531 0.0239375
R4728 VSS.n4735 VSS 0.0239375
R4729 VSS.n4662 VSS 0.0239375
R4730 VSS VSS.n3874 0.0239375
R4731 VSS.n3880 VSS.n3876 0.0239375
R4732 VSS.n3739 VSS.n3730 0.0239375
R4733 VSS.n3714 VSS.n3290 0.0239375
R4734 VSS.n1454 VSS.n1450 0.0239375
R4735 VSS.n1460 VSS.n1459 0.0239375
R4736 VSS.n1958 VSS.n1954 0.0239375
R4737 VSS.n114 VSS.n42 0.0239375
R4738 VSS.n113 VSS.n43 0.0239375
R4739 VSS.n178 VSS.n172 0.0239375
R4740 VSS VSS.n278 0.0239375
R4741 VSS.n3008 VSS.n3007 0.0239375
R4742 VSS.n3026 VSS.n3020 0.0239375
R4743 VSS.n4417 VSS.n4415 0.0239375
R4744 VSS.n4433 VSS.n4429 0.0239375
R4745 VSS.n4439 VSS.n4438 0.0239375
R4746 VSS.n1248 VSS.n1244 0.0239375
R4747 VSS.n1254 VSS.n1253 0.0239375
R4748 VSS.n662 VSS.n658 0.0239375
R4749 VSS.n780 VSS.n779 0.0239375
R4750 VSS.n4797 VSS.n4796 0.0239375
R4751 VSS.n4095 VSS.n3979 0.0239375
R4752 VSS.n3969 VSS.n3963 0.0239375
R4753 VSS.n3014 VSS.n3013 0.0235594
R4754 VSS.n2987 VSS.n2986 0.0231188
R4755 VSS.n4216 VSS.n4215 0.0226781
R4756 VSS.n1860 VSS.n1828 0.0226354
R4757 VSS VSS.n2076 0.0226354
R4758 VSS.n2567 VSS 0.0226354
R4759 VSS.n3740 VSS.n3727 0.0226354
R4760 VSS.n3482 VSS.n3481 0.0226354
R4761 VSS.n1038 VSS.n1028 0.0226354
R4762 VSS.n1493 VSS.n1486 0.0226354
R4763 VSS.n1520 VSS 0.0226354
R4764 VSS.n1959 VSS.n1949 0.0226354
R4765 VSS.n379 VSS.n368 0.0226354
R4766 VSS.n422 VSS.n421 0.0226354
R4767 VSS.n405 VSS.n404 0.0226354
R4768 VSS.n4856 VSS.n4854 0.0226354
R4769 VSS.n4504 VSS.n4502 0.0226354
R4770 VSS.n1005 VSS.n1004 0.0226354
R4771 VSS VSS.n1309 0.0226354
R4772 VSS.n833 VSS.n827 0.0226354
R4773 VSS.n4791 VSS.n4787 0.0226354
R4774 VSS.n4598 VSS.n4595 0.0226354
R4775 VSS.n4000 VSS.n3998 0.0226354
R4776 VSS.n4515 VSS.n4514 0.0225312
R4777 VSS.n4487 VSS.n4486 0.0225312
R4778 VSS.n1606 VSS.n1605 0.0225312
R4779 VSS.n2049 VSS.n2047 0.0224595
R4780 VSS.n2049 VSS.n2048 0.0224595
R4781 VSS.n1937 VSS.n1919 0.0224595
R4782 VSS.n1937 VSS.n1936 0.0224595
R4783 VSS.n1328 VSS.n1323 0.0224595
R4784 VSS.n1328 VSS.n1324 0.0224595
R4785 VSS.n4337 VSS.n4317 0.0224595
R4786 VSS.n4337 VSS.n4336 0.0224595
R4787 VSS.n4212 VSS.n4194 0.0224595
R4788 VSS.n4212 VSS.n4211 0.0224595
R4789 VSS.n3130 VSS.n3120 0.0224595
R4790 VSS.n3130 VSS.n3121 0.0224595
R4791 VSS.n1797 VSS.n924 0.0224595
R4792 VSS.n1797 VSS.n925 0.0224595
R4793 VSS.n140 VSS.n138 0.0224595
R4794 VSS.n140 VSS.n139 0.0224595
R4795 VSS.n4649 VSS.n2826 0.0224595
R4796 VSS.n4649 VSS.n2827 0.0224595
R4797 VSS.n4583 VSS.n4561 0.0224595
R4798 VSS.n4583 VSS.n4562 0.0224595
R4799 VSS.n3037 VSS.n3036 0.0223844
R4800 VSS.n4992 VSS.n4991 0.0222375
R4801 VSS.n4464 VSS.n4463 0.0222375
R4802 VSS.n4191 VSS.n4190 0.0219438
R4803 VSS.n4989 VSS.n4988 0.0217969
R4804 VSS.n4986 VSS.n4985 0.0217969
R4805 VSS.n5025 VSS.n5024 0.02165
R4806 VSS.n4493 VSS.n4492 0.0215031
R4807 VSS.n2511 VSS.n2510 0.0214906
R4808 VSS.n4770 VSS.n4769 0.0214906
R4809 VSS.n4643 VSS.n4642 0.0214567
R4810 VSS.n3912 VSS.n3911 0.0214567
R4811 VSS.n2915 VSS.n2914 0.0213563
R4812 VSS.n1087 VSS.n1075 0.0213333
R4813 VSS.n1143 VSS.n1142 0.0213333
R4814 VSS.n1213 VSS.n1212 0.0213333
R4815 VSS.n974 VSS.n973 0.0213333
R4816 VSS.n1621 VSS.n1616 0.0213333
R4817 VSS.n905 VSS.n904 0.0213333
R4818 VSS.n2236 VSS.n2235 0.0213333
R4819 VSS.n2223 VSS.n2087 0.0213333
R4820 VSS.n2221 VSS.n2220 0.0213333
R4821 VSS.n2207 VSS.n2206 0.0213333
R4822 VSS.n2193 VSS.n2192 0.0213333
R4823 VSS.n2176 VSS.n2175 0.0213333
R4824 VSS.n2139 VSS.n2138 0.0213333
R4825 VSS.n2125 VSS.n2124 0.0213333
R4826 VSS.n628 VSS.n609 0.0213333
R4827 VSS VSS.n2565 0.0213333
R4828 VSS.n2568 VSS.n2566 0.0213333
R4829 VSS.n2584 VSS.n583 0.0213333
R4830 VSS.n2597 VSS.n2586 0.0213333
R4831 VSS.n2611 VSS.n2599 0.0213333
R4832 VSS.n2628 VSS.n2613 0.0213333
R4833 VSS.n2642 VSS.n2630 0.0213333
R4834 VSS.n2655 VSS.n2644 0.0213333
R4835 VSS.n2669 VSS.n2657 0.0213333
R4836 VSS.n2689 VSS.n2671 0.0213333
R4837 VSS.n2747 VSS.n2746 0.0213333
R4838 VSS VSS.n2772 0.0213333
R4839 VSS.n4663 VSS 0.0213333
R4840 VSS.n3750 VSS 0.0213333
R4841 VSS.n3673 VSS 0.0213333
R4842 VSS.n3424 VSS 0.0213333
R4843 VSS.n3595 VSS.n3594 0.0213333
R4844 VSS.n3621 VSS 0.0213333
R4845 VSS.n21 VSS.n16 0.0213333
R4846 VSS.n210 VSS.n204 0.0213333
R4847 VSS.n2957 VSS.n2951 0.0213333
R4848 VSS.n4474 VSS.n4469 0.0213333
R4849 VSS.n4482 VSS.n4481 0.0213333
R4850 VSS.n878 VSS.n876 0.0213333
R4851 VSS.n2465 VSS.n2460 0.0213333
R4852 VSS.n4305 VSS.n4130 0.0213333
R4853 VSS.n4490 VSS.n4489 0.0210625
R4854 VSS.n4223 VSS.n4222 0.0209156
R4855 VSS.n4551 VSS.n4518 0.0207703
R4856 VSS.n3235 VSS.n3234 0.0207703
R4857 VSS.n3552 VSS.n3551 0.0207703
R4858 VSS.n3773 VSS.n3769 0.0207703
R4859 VSS.n1091 VSS.n1047 0.0207703
R4860 VSS.n696 VSS.n691 0.0207703
R4861 VSS.n2721 VSS.n582 0.0207703
R4862 VSS.n332 VSS.n331 0.0207703
R4863 VSS.n4691 VSS.n2806 0.0207703
R4864 VSS.n4982 VSS.n4838 0.0206429
R4865 VSS.n5074 VSS.n5073 0.0206219
R4866 VSS.n4556 VSS.n4555 0.0205411
R4867 VSS.n5023 VSS.n136 0.0205072
R4868 VSS.n4457 VSS.n4315 0.0205072
R4869 VSS.n2940 VSS.n2939 0.0203281
R4870 VSS.n2963 VSS.n2962 0.0203281
R4871 VSS.n5017 VSS.n5016 0.0200344
R4872 VSS.n5071 VSS.n5070 0.0200344
R4873 VSS.n1777 VSS.n1776 0.0200312
R4874 VSS.n939 VSS.n927 0.0200312
R4875 VSS.n1827 VSS.n1826 0.0200312
R4876 VSS.n1858 VSS.n1843 0.0200312
R4877 VSS.n1840 VSS.n1829 0.0200312
R4878 VSS.n903 VSS.n902 0.0200312
R4879 VSS.n2001 VSS.n2000 0.0200312
R4880 VSS.n2162 VSS.n2161 0.0200312
R4881 VSS.n2159 VSS.n2158 0.0200312
R4882 VSS.n2755 VSS.n2737 0.0200312
R4883 VSS.n564 VSS.n562 0.0200312
R4884 VSS.n3422 VSS.n3416 0.0200312
R4885 VSS.n3450 VSS.n3443 0.0200312
R4886 VSS.n3339 VSS.n3338 0.0200312
R4887 VSS.n3313 VSS.n3309 0.0200312
R4888 VSS.n1599 VSS.n1598 0.0200312
R4889 VSS.n1438 VSS.n1435 0.0200312
R4890 VSS.n1909 VSS.n1908 0.0200312
R4891 VSS.n26 VSS.n11 0.0200312
R4892 VSS.n98 VSS.n91 0.0200312
R4893 VSS.n327 VSS.n279 0.0200312
R4894 VSS.n4905 VSS.n4904 0.0200312
R4895 VSS.n4895 VSS.n4890 0.0200312
R4896 VSS.n2925 VSS.n2920 0.0200312
R4897 VSS.n2935 VSS.n2934 0.0200312
R4898 VSS.n3057 VSS.n3050 0.0200312
R4899 VSS.n3119 VSS 0.0200312
R4900 VSS.n4391 VSS.n4387 0.0200312
R4901 VSS.n1411 VSS.n1410 0.0200312
R4902 VSS.n805 VSS.n803 0.0200312
R4903 VSS.n3939 VSS.n3938 0.0200312
R4904 VSS.n4390 VSS.n4389 0.0190811
R4905 VSS.n90 VSS.n85 0.0190811
R4906 VSS.n1601 VSS.n1575 0.0190811
R4907 VSS.n1911 VSS.n1895 0.0190811
R4908 VSS.n28 VSS.n27 0.0190811
R4909 VSS.n3341 VSS.n3323 0.0190811
R4910 VSS.n2756 VSS.n2727 0.0190811
R4911 VSS.n2936 VSS.n2918 0.0190811
R4912 VSS.n4903 VSS.n4899 0.0190811
R4913 VSS.n3442 VSS.n3438 0.0190811
R4914 VSS.n3421 VSS.n3418 0.0190811
R4915 VSS.n3940 VSS.n3918 0.0190811
R4916 VSS.n1412 VSS.n1294 0.0190811
R4917 VSS.n1090 VSS.n1089 0.0187292
R4918 VSS.n2719 VSS.n2718 0.0187292
R4919 VSS.n4692 VSS.n2805 0.0187292
R4920 VSS.n2818 VSS.n2816 0.0187292
R4921 VSS.n3774 VSS.n3767 0.0187292
R4922 VSS.n3904 VSS.n3894 0.0187292
R4923 VSS.n3550 VSS.n3535 0.0187292
R4924 VSS.n3547 VSS.n3542 0.0187292
R4925 VSS.n2021 VSS.n2019 0.0187292
R4926 VSS.n51 VSS.n49 0.0187292
R4927 VSS.n5044 VSS.n5039 0.0187292
R4928 VSS.n152 VSS.n150 0.0187292
R4929 VSS.n306 VSS.n304 0.0187292
R4930 VSS.n330 VSS.n278 0.0187292
R4931 VSS.n4966 VSS.n4964 0.0187292
R4932 VSS.n3158 VSS.n3156 0.0187292
R4933 VSS.n4550 VSS.n4549 0.0187292
R4934 VSS.n3233 VSS.n3218 0.0187292
R4935 VSS.n3229 VSS.n3223 0.0187292
R4936 VSS.n1301 VSS.n1296 0.0187292
R4937 VSS.n697 VSS.n690 0.0187292
R4938 VSS.n4827 VSS.n478 0.0187292
R4939 VSS.n4109 VSS.n4107 0.0187292
R4940 VSS.n1019 VSS.n1018 0.0179804
R4941 VSS.n4555 VSS.n4554 0.0178313
R4942 VSS.n1165 VSS.n1160 0.0174271
R4943 VSS.n1796 VSS.n926 0.0174271
R4944 VSS.n1796 VSS.n1795 0.0174271
R4945 VSS.n943 VSS.n942 0.0174271
R4946 VSS.n2714 VSS.n2713 0.0174271
R4947 VSS.n4651 VSS.n4650 0.0174271
R4948 VSS.n4650 VSS.n2825 0.0174271
R4949 VSS.n5060 VSS.n5058 0.0174271
R4950 VSS.n5048 VSS.n5047 0.0174271
R4951 VSS.n5047 VSS.n5046 0.0174271
R4952 VSS.n4941 VSS.n4934 0.0174271
R4953 VSS.n2976 VSS.n2974 0.0174271
R4954 VSS.n3133 VSS.n3131 0.0174271
R4955 VSS.n3131 VSS.n3119 0.0174271
R4956 VSS.n4542 VSS.n4537 0.0174271
R4957 VSS.n3247 VSS.n3245 0.0174271
R4958 VSS.n4335 VSS.n4322 0.0174271
R4959 VSS.n4335 VSS.n4334 0.0174271
R4960 VSS.n4332 VSS.n4327 0.0174271
R4961 VSS.n4202 VSS.n4195 0.0174271
R4962 VSS.n4210 VSS.n4204 0.0174271
R4963 VSS.n4210 VSS.n4209 0.0174271
R4964 VSS.n1331 VSS.n1329 0.0174271
R4965 VSS.n1329 VSS.n1322 0.0174271
R4966 VSS.n1935 VSS.n1927 0.0174271
R4967 VSS.n1935 VSS.n1934 0.0174271
R4968 VSS.n847 VSS.n846 0.0174271
R4969 VSS.n849 VSS.n847 0.0174271
R4970 VSS.n854 VSS.n853 0.0174271
R4971 VSS.n2489 VSS.n2487 0.0174271
R4972 VSS.n686 VSS.n681 0.0174271
R4973 VSS.n4568 VSS.n4563 0.0174271
R4974 VSS.n4582 VSS.n4570 0.0174271
R4975 VSS.n4582 VSS.n4581 0.0174271
R4976 VSS.n1158 VSS.n1157 0.0174271
R4977 VSS.n4307 VSS.n4306 0.0173919
R4978 VSS.n4483 VSS.n4467 0.0173919
R4979 VSS.n3593 VSS.n3318 0.0173919
R4980 VSS.n1615 VSS.n976 0.0173919
R4981 VSS.n212 VSS.n211 0.0173919
R4982 VSS.n2959 VSS.n2958 0.0173919
R4983 VSS.n5023 VSS.n5022 0.0172437
R4984 VSS.n1060 VSS.n1059 0.016125
R4985 VSS.n1090 VSS.n1074 0.016125
R4986 VSS.n2719 VSS.n2712 0.016125
R4987 VSS.n4693 VSS.n4692 0.016125
R4988 VSS.n2803 VSS.n2798 0.016125
R4989 VSS.n3775 VSS.n3774 0.016125
R4990 VSS.n3550 VSS.n3549 0.016125
R4991 VSS.n3336 VSS.n3329 0.016125
R4992 VSS.n100 VSS.n99 0.016125
R4993 VSS.n258 VSS.n256 0.016125
R4994 VSS.n330 VSS.n329 0.016125
R4995 VSS.n3134 VSS.n3118 0.016125
R4996 VSS.n3180 VSS.n3178 0.016125
R4997 VSS.n4550 VSS.n4544 0.016125
R4998 VSS.n3233 VSS.n3232 0.016125
R4999 VSS.n4235 VSS.n4234 0.016125
R5000 VSS.n1337 VSS.n1336 0.016125
R5001 VSS.n1925 VSS.n1920 0.016125
R5002 VSS.n698 VSS.n697 0.016125
R5003 VSS.n1006 VSS.n988 0.0157027
R5004 VSS.n1485 VSS.n1483 0.0157027
R5005 VSS.n1040 VSS.n1039 0.0157027
R5006 VSS.n3484 VSS.n3365 0.0157027
R5007 VSS.n4846 VSS.n4844 0.0157027
R5008 VSS.n424 VSS.n389 0.0157027
R5009 VSS.n381 VSS.n380 0.0157027
R5010 VSS.n834 VSS.n813 0.0157027
R5011 VSS.n2051 VSS.n2046 0.0152558
R5012 VSS.n2051 VSS.n2050 0.0152558
R5013 VSS.n1938 VSS.n1917 0.0152558
R5014 VSS.n1938 VSS.n1918 0.0152558
R5015 VSS.n1889 VSS.n1868 0.0152558
R5016 VSS.n1889 VSS.n1869 0.0152558
R5017 VSS.n1256 VSS.n1239 0.0152558
R5018 VSS.n1256 VSS.n1240 0.0152558
R5019 VSS.n1124 VSS.n1097 0.0152558
R5020 VSS.n1124 VSS.n1123 0.0152558
R5021 VSS.n1007 VSS.n986 0.0152558
R5022 VSS.n1007 VSS.n987 0.0152558
R5023 VSS.n1327 VSS.n1325 0.0152558
R5024 VSS.n1327 VSS.n1326 0.0152558
R5025 VSS.n887 VSS.n868 0.0152558
R5026 VSS.n887 VSS.n869 0.0152558
R5027 VSS.n2373 VSS.n867 0.0152558
R5028 VSS.n2373 VSS.n2372 0.0152558
R5029 VSS.n3972 VSS.n3944 0.0152558
R5030 VSS.n4097 VSS.n3975 0.0152558
R5031 VSS.n4118 VSS.n4100 0.0152558
R5032 VSS.n4308 VSS.n4121 0.0152558
R5033 VSS.n4220 VSS.n4217 0.0152558
R5034 VSS.n4345 VSS.n4344 0.0152558
R5035 VSS.n1419 VSS.n1416 0.0152558
R5036 VSS.n1466 VSS.n1464 0.0152558
R5037 VSS.n1466 VSS.n1465 0.0152558
R5038 VSS.n1470 VSS.n1467 0.0152558
R5039 VSS.n4370 VSS.n4350 0.0152558
R5040 VSS.n4443 VSS.n4442 0.0152558
R5041 VSS.n3210 VSS.n3191 0.0152558
R5042 VSS.n3210 VSS.n3192 0.0152558
R5043 VSS.n3261 VSS.n3259 0.0152558
R5044 VSS.n3261 VSS.n3260 0.0152558
R5045 VSS.n4450 VSS.n4446 0.0152558
R5046 VSS.n5065 VSS.n5026 0.0152558
R5047 VSS.n5065 VSS.n5064 0.0152558
R5048 VSS.n135 VSS.n117 0.0152558
R5049 VSS.n135 VSS.n118 0.0152558
R5050 VSS.n116 VSS.n37 0.0152558
R5051 VSS.n116 VSS.n38 0.0152558
R5052 VSS.n89 VSS.n87 0.0152558
R5053 VSS.n89 VSS.n88 0.0152558
R5054 VSS.n2058 VSS.n2055 0.0152558
R5055 VSS.n36 VSS.n34 0.0152558
R5056 VSS.n36 VSS.n35 0.0152558
R5057 VSS.n1441 VSS.n1420 0.0152558
R5058 VSS.n1441 VSS.n1421 0.0152558
R5059 VSS.n1041 VSS.n980 0.0152558
R5060 VSS.n1041 VSS.n981 0.0152558
R5061 VSS.n1013 VSS.n1012 0.0152558
R5062 VSS.n1195 VSS.n1172 0.0152558
R5063 VSS.n1195 VSS.n1173 0.0152558
R5064 VSS.n1288 VSS.n1261 0.0152558
R5065 VSS.n1288 VSS.n1287 0.0152558
R5066 VSS.n1603 VSS.n1574 0.0152558
R5067 VSS.n1603 VSS.n1602 0.0152558
R5068 VSS.n1463 VSS.n1442 0.0152558
R5069 VSS.n1463 VSS.n1443 0.0152558
R5070 VSS.n1473 VSS.n1471 0.0152558
R5071 VSS.n1473 VSS.n1472 0.0152558
R5072 VSS.n1552 VSS.n1474 0.0152558
R5073 VSS.n1552 VSS.n1551 0.0152558
R5074 VSS.n2035 VSS.n2010 0.0152558
R5075 VSS.n2035 VSS.n2011 0.0152558
R5076 VSS.n1963 VSS.n1940 0.0152558
R5077 VSS.n1963 VSS.n1941 0.0152558
R5078 VSS.n1912 VSS.n1893 0.0152558
R5079 VSS.n1912 VSS.n1894 0.0152558
R5080 VSS.n1807 VSS.n1804 0.0152558
R5081 VSS.n29 VSS.n0 0.0152558
R5082 VSS.n29 VSS.n1 0.0152558
R5083 VSS.n33 VSS.n31 0.0152558
R5084 VSS.n33 VSS.n32 0.0152558
R5085 VSS.n4512 VSS.n4494 0.0152558
R5086 VSS.n4512 VSS.n4495 0.0152558
R5087 VSS.n4552 VSS.n4516 0.0152558
R5088 VSS.n4552 VSS.n4517 0.0152558
R5089 VSS.n3236 VSS.n3211 0.0152558
R5090 VSS.n3236 VSS.n3212 0.0152558
R5091 VSS.n4484 VSS.n4465 0.0152558
R5092 VSS.n4484 VSS.n4466 0.0152558
R5093 VSS.n3258 VSS.n3237 0.0152558
R5094 VSS.n3258 VSS.n3238 0.0152558
R5095 VSS.n4400 VSS.n4399 0.0152558
R5096 VSS.n4338 VSS.n4316 0.0152558
R5097 VSS.n4213 VSS.n4192 0.0152558
R5098 VSS.n4213 VSS.n4193 0.0152558
R5099 VSS.n3556 VSS.n3555 0.0152558
R5100 VSS.n3553 VSS.n3345 0.0152558
R5101 VSS.n3343 VSS.n3342 0.0152558
R5102 VSS.n3587 VSS.n3565 0.0152558
R5103 VSS.n3592 VSS.n3591 0.0152558
R5104 VSS.n3485 VSS.n3364 0.0152558
R5105 VSS.n3109 VSS.n3087 0.0152558
R5106 VSS.n3161 VSS.n3112 0.0152558
R5107 VSS.n3085 VSS.n3080 0.0152558
R5108 VSS.n3183 VSS.n3165 0.0152558
R5109 VSS.n3078 VSS.n3074 0.0152558
R5110 VSS.n3129 VSS.n3122 0.0152558
R5111 VSS.n4615 VSS.n4614 0.0152558
R5112 VSS.n4636 VSS.n4589 0.0152558
R5113 VSS.n3265 VSS.n3264 0.0152558
R5114 VSS.n3716 VSS.n3267 0.0152558
R5115 VSS.n3742 VSS.n3718 0.0152558
R5116 VSS.n3907 VSS.n3884 0.0152558
R5117 VSS.n3882 VSS.n3745 0.0152558
R5118 VSS.n3772 VSS.n3770 0.0152558
R5119 VSS.n2005 VSS.n889 0.0152558
R5120 VSS.n1237 VSS.n1200 0.0152558
R5121 VSS.n1237 VSS.n1236 0.0152558
R5122 VSS.n2044 VSS.n2040 0.0152558
R5123 VSS.n2366 VSS.n2063 0.0152558
R5124 VSS.n1864 VSS.n1811 0.0152558
R5125 VSS.n1864 VSS.n1812 0.0152558
R5126 VSS.n1973 VSS.n920 0.0152558
R5127 VSS.n1973 VSS.n1972 0.0152558
R5128 VSS.n1798 VSS.n922 0.0152558
R5129 VSS.n1798 VSS.n923 0.0152558
R5130 VSS.n1614 VSS.n978 0.0152558
R5131 VSS.n1614 VSS.n1613 0.0152558
R5132 VSS.n1168 VSS.n1126 0.0152558
R5133 VSS.n1168 VSS.n1127 0.0152558
R5134 VSS.n1092 VSS.n1045 0.0152558
R5135 VSS.n1092 VSS.n1046 0.0152558
R5136 VSS.n4952 VSS.n4948 0.0152558
R5137 VSS.n4945 VSS.n4871 0.0152558
R5138 VSS.n4974 VSS.n4954 0.0152558
R5139 VSS.n4847 VSS.n4843 0.0152558
R5140 VSS.n4865 VSS.n4849 0.0152558
R5141 VSS.n4840 VSS.n4839 0.0152558
R5142 VSS.n2757 VSS.n2725 0.0152558
R5143 VSS.n4806 VSS.n4805 0.0152558
R5144 VSS.n4800 VSS.n4780 0.0152558
R5145 VSS.n4831 VSS.n428 0.0152558
R5146 VSS.n695 VSS.n693 0.0152558
R5147 VSS.n4776 VSS.n4775 0.0152558
R5148 VSS.n4762 VSS.n4761 0.0152558
R5149 VSS.n2722 VSS.n581 0.0152558
R5150 VSS.n568 VSS.n497 0.0152558
R5151 VSS.n494 VSS.n491 0.0152558
R5152 VSS.n355 VSS.n334 0.0152558
R5153 VSS.n355 VSS.n335 0.0152558
R5154 VSS.n5014 VSS.n4996 0.0152558
R5155 VSS.n5014 VSS.n4997 0.0152558
R5156 VSS.n333 VSS.n275 0.0152558
R5157 VSS.n333 VSS.n276 0.0152558
R5158 VSS.n425 VSS.n387 0.0152558
R5159 VSS.n425 VSS.n388 0.0152558
R5160 VSS.n386 VSS.n383 0.0152558
R5161 VSS.n382 VSS.n356 0.0152558
R5162 VSS.n382 VSS.n357 0.0152558
R5163 VSS.n274 VSS.n272 0.0152558
R5164 VSS.n274 VSS.n273 0.0152558
R5165 VSS.n184 VSS.n183 0.0152558
R5166 VSS.n161 VSS.n143 0.0152558
R5167 VSS.n238 VSS.n218 0.0152558
R5168 VSS.n181 VSS.n163 0.0152558
R5169 VSS.n213 VSS.n193 0.0152558
R5170 VSS.n141 VSS.n137 0.0152558
R5171 VSS.n262 VSS.n243 0.0152558
R5172 VSS.n2524 VSS.n604 0.0152558
R5173 VSS.n635 VSS.n605 0.0152558
R5174 VSS.n2144 VSS.n2143 0.0152558
R5175 VSS.n835 VSS.n811 0.0152558
R5176 VSS.n643 VSS.n639 0.0152558
R5177 VSS.n2503 VSS.n839 0.0152558
R5178 VSS.n649 VSS.n645 0.0152558
R5179 VSS.n808 VSS.n790 0.0152558
R5180 VSS.n783 VSS.n651 0.0152558
R5181 VSS.n2937 VSS.n2916 0.0152558
R5182 VSS.n2937 VSS.n2917 0.0152558
R5183 VSS.n4902 VSS.n4900 0.0152558
R5184 VSS.n4902 VSS.n4901 0.0152558
R5185 VSS.n3034 VSS.n3015 0.0152558
R5186 VSS.n3034 VSS.n3016 0.0152558
R5187 VSS.n3011 VSS.n2988 0.0152558
R5188 VSS.n3011 VSS.n2989 0.0152558
R5189 VSS.n2984 VSS.n2964 0.0152558
R5190 VSS.n2984 VSS.n2965 0.0152558
R5191 VSS.n2960 VSS.n2941 0.0152558
R5192 VSS.n2960 VSS.n2942 0.0152558
R5193 VSS.n2912 VSS.n2891 0.0152558
R5194 VSS.n2912 VSS.n2892 0.0152558
R5195 VSS.n3072 VSS.n3038 0.0152558
R5196 VSS.n3072 VSS.n3039 0.0152558
R5197 VSS.n4758 VSS.n2760 0.0152558
R5198 VSS.n4689 VSS.n2807 0.0152558
R5199 VSS.n4685 VSS.n4684 0.0152558
R5200 VSS.n4648 VSS.n2828 0.0152558
R5201 VSS.n2886 VSS.n2829 0.0152558
R5202 VSS.n4584 VSS.n4560 0.0152558
R5203 VSS.n4004 VSS.n4003 0.0152558
R5204 VSS.n3441 VSS.n3439 0.0152558
R5205 VSS.n3490 VSS.n3489 0.0152558
R5206 VSS.n3420 VSS.n3419 0.0152558
R5207 VSS.n4225 VSS.n4156 0.0152558
R5208 VSS.n4188 VSS.n4157 0.0152558
R5209 VSS.n4188 VSS.n4187 0.0152558
R5210 VSS.n3941 VSS.n3917 0.0152558
R5211 VSS.n1414 VSS.n1293 0.0152558
R5212 VSS.n1414 VSS.n1413 0.0152558
R5213 VSS.n1624 VSS.n1623 0.0148229
R5214 VSS.n1665 VSS.n1650 0.0148229
R5215 VSS.n1679 VSS.n1667 0.0148229
R5216 VSS.n1692 VSS.n1681 0.0148229
R5217 VSS.n1706 VSS.n1694 0.0148229
R5218 VSS.n1722 VSS.n1708 0.0148229
R5219 VSS.n1736 VSS.n1724 0.0148229
R5220 VSS.n1750 VSS.n1738 0.0148229
R5221 VSS.n1754 VSS.n1752 0.0148229
R5222 VSS.n1773 VSS.n951 0.0148229
R5223 VSS.n2362 VSS.n2361 0.0148229
R5224 VSS.n2339 VSS.n2338 0.0148229
R5225 VSS.n2325 VSS.n2324 0.0148229
R5226 VSS.n2322 VSS.n2321 0.0148229
R5227 VSS.n2308 VSS.n2307 0.0148229
R5228 VSS.n2292 VSS.n2291 0.0148229
R5229 VSS.n2278 VSS.n2277 0.0148229
R5230 VSS.n2264 VSS.n2263 0.0148229
R5231 VSS.n2261 VSS.n2260 0.0148229
R5232 VSS.n2755 VSS.n2754 0.0148229
R5233 VSS.n2771 VSS.n2764 0.0148229
R5234 VSS.n3757 VSS.n3756 0.0148229
R5235 VSS.n3713 VSS 0.0148229
R5236 VSS.n3423 VSS.n3422 0.0148229
R5237 VSS.n3452 VSS.n3451 0.0148229
R5238 VSS.n3443 VSS.n3347 0.0148229
R5239 VSS.n3339 VSS.n3328 0.0148229
R5240 VSS.n1191 VSS.n1189 0.0148229
R5241 VSS.n1599 VSS.n1586 0.0148229
R5242 VSS.n1596 VSS.n1591 0.0148229
R5243 VSS.n1909 VSS.n1900 0.0148229
R5244 VSS.n1906 VSS.n1901 0.0148229
R5245 VSS.n26 VSS.n25 0.0148229
R5246 VSS.n91 VSS.n84 0.0148229
R5247 VSS.n4881 VSS 0.0148229
R5248 VSS.n4904 VSS.n4897 0.0148229
R5249 VSS.n2935 VSS.n2929 0.0148229
R5250 VSS.n3048 VSS.n3046 0.0148229
R5251 VSS.n3207 VSS.n3205 0.0148229
R5252 VSS.n4392 VSS.n4391 0.0148229
R5253 VSS.n1411 VSS.n1304 0.0148229
R5254 VSS.n487 VSS.n481 0.0148229
R5255 VSS.n2877 VSS.n2875 0.0148229
R5256 VSS.n3939 VSS.n3926 0.0148229
R5257 VSS.n3936 VSS.n3931 0.0148229
R5258 VSS.n3971 VSS.n3970 0.0140135
R5259 VSS.n4449 VSS.n4447 0.0140135
R5260 VSS.n1962 VSS.n1961 0.0140135
R5261 VSS.n3715 VSS.n3269 0.0140135
R5262 VSS.n3741 VSS.n3721 0.0140135
R5263 VSS.n3881 VSS.n3747 0.0140135
R5264 VSS.n1863 VSS.n1862 0.0140135
R5265 VSS.n4799 VSS.n4782 0.0140135
R5266 VSS.n180 VSS.n179 0.0140135
R5267 VSS.n3010 VSS.n2990 0.0140135
R5268 VSS.n1232 VSS.n1218 0.0135208
R5269 VSS.n1216 VSS.n1215 0.0135208
R5270 VSS.n1616 VSS.n975 0.0135208
R5271 VSS VSS.n1774 0.0135208
R5272 VSS.n1978 VSS.n1977 0.0135208
R5273 VSS.n2237 VSS 0.0135208
R5274 VSS.n3414 VSS.n3409 0.0135208
R5275 VSS.n3594 VSS.n3317 0.0135208
R5276 VSS.n172 VSS.n170 0.0135208
R5277 VSS.n202 VSS.n195 0.0135208
R5278 VSS.n210 VSS.n209 0.0135208
R5279 VSS.n419 VSS.n414 0.0135208
R5280 VSS.n2957 VSS.n2956 0.0135208
R5281 VSS.n4482 VSS.n4476 0.0135208
R5282 VSS.n4385 VSS.n4380 0.0135208
R5283 VSS.n4360 VSS.n4358 0.0135208
R5284 VSS.n3963 VSS.n3961 0.0135208
R5285 VSS.n4305 VSS.n4304 0.0135208
R5286 VSS.n1255 VSS.n1242 0.0123243
R5287 VSS.n4369 VSS.n4352 0.0123243
R5288 VSS.n4441 VSS.n4373 0.0123243
R5289 VSS.n115 VSS.n41 0.0123243
R5290 VSS.n1462 VSS.n1445 0.0123243
R5291 VSS.n4951 VSS.n4949 0.0123243
R5292 VSS.n4807 VSS.n489 0.0123243
R5293 VSS.n2525 VSS.n603 0.0123243
R5294 VSS.n782 VSS.n653 0.0123243
R5295 VSS.n2885 VSS.n2884 0.0123243
R5296 VSS.n1977 VSS.n1976 0.0122188
R5297 VSS.n3290 VSS.n3271 0.0122188
R5298 VSS.n3482 VSS.n3432 0.0122188
R5299 VSS.n3479 VSS.n3478 0.0122188
R5300 VSS.n1038 VSS.n1037 0.0122188
R5301 VSS.n1486 VSS.n1482 0.0122188
R5302 VSS.n1495 VSS.n1494 0.0122188
R5303 VSS.n368 VSS.n364 0.0122188
R5304 VSS.n379 VSS.n378 0.0122188
R5305 VSS.n422 VSS.n399 0.0122188
R5306 VSS.n409 VSS.n405 0.0122188
R5307 VSS.n4908 VSS.n4884 0.0122188
R5308 VSS.n2949 VSS.n2944 0.0122188
R5309 VSS.n3007 VSS.n3005 0.0122188
R5310 VSS.n4422 VSS.n4417 0.0122188
R5311 VSS.n1005 VSS.n993 0.0122188
R5312 VSS.n827 VSS.n825 0.0122188
R5313 VSS.n833 VSS.n832 0.0122188
R5314 VSS.n4128 VSS.n4123 0.0122188
R5315 VSS.n4458 VSS.n4457 0.0113687
R5316 VSS.n3880 VSS.n3879 0.0109167
R5317 VSS.n3740 VSS.n3739 0.0109167
R5318 VSS.n3271 VSS.n3270 0.0109167
R5319 VSS.n3714 VSS.n3713 0.0109167
R5320 VSS.n3481 VSS.n3479 0.0109167
R5321 VSS.n1494 VSS.n1493 0.0109167
R5322 VSS.n1959 VSS.n1958 0.0109167
R5323 VSS.n178 VSS.n177 0.0109167
R5324 VSS.n364 VSS.n359 0.0109167
R5325 VSS.n4908 VSS.n4907 0.0109167
R5326 VSS.n2951 VSS.n2949 0.0109167
R5327 VSS.n3008 VSS.n2995 0.0109167
R5328 VSS.n3005 VSS.n3000 0.0109167
R5329 VSS.n4415 VSS.n4414 0.0109167
R5330 VSS.n4423 VSS.n4422 0.0109167
R5331 VSS.n825 VSS.n820 0.0109167
R5332 VSS.n4797 VSS.n4791 0.0109167
R5333 VSS.n3969 VSS.n3968 0.0109167
R5334 VSS.n4130 VSS.n4128 0.0109167
R5335 VSS.n4096 VSS.n3978 0.0106351
R5336 VSS.n3209 VSS.n3193 0.0106351
R5337 VSS.n1194 VSS.n1174 0.0106351
R5338 VSS.n1975 VSS.n919 0.0106351
R5339 VSS.n3033 VSS.n3018 0.0106351
R5340 VSS.n3071 VSS.n3070 0.0106351
R5341 VSS.n4757 VSS.n2762 0.0106351
R5342 VSS.n3876 VSS.n3875 0.0102525
R5343 VSS.n2531 VSS.n2526 0.00961458
R5344 VSS.n3416 VSS.n3414 0.00961458
R5345 VSS.n1018 VSS 0.00961458
R5346 VSS.n1460 VSS.n1454 0.00961458
R5347 VSS.n114 VSS.n113 0.00961458
R5348 VSS.n170 VSS.n165 0.00961458
R5349 VSS.n204 VSS.n202 0.00961458
R5350 VSS.n421 VSS.n419 0.00961458
R5351 VSS.n4882 VSS.n4881 0.00961458
R5352 VSS.n4387 VSS.n4385 0.00961458
R5353 VSS.n4439 VSS.n4433 0.00961458
R5354 VSS.n4358 VSS.n4353 0.00961458
R5355 VSS.n4368 VSS.n4367 0.00961458
R5356 VSS.n1254 VSS.n1248 0.00961458
R5357 VSS.n780 VSS.n662 0.00961458
R5358 VSS.n4809 VSS.n4808 0.00961458
R5359 VSS.n2883 VSS.n2882 0.00961458
R5360 VSS.n3961 VSS.n3956 0.00961458
R5361 VSS.n1518 VSS.n1517 0.00894595
R5362 VSS.n3586 VSS.n3567 0.00894595
R5363 VSS.n3182 VSS.n3166 0.00894595
R5364 VSS.n1235 VSS.n1201 0.00894595
R5365 VSS.n5013 VSS.n5000 0.00894595
R5366 VSS.n261 VSS.n244 0.00894595
R5367 VSS.n2911 VSS.n2895 0.00894595
R5368 VSS.n4226 VSS.n4154 0.00894595
R5369 VSS.n4186 VSS.n4160 0.00894595
R5370 VSS.n1558 VSS.n1557 0.00887187
R5371 VSS.n1217 VSS.n1216 0.0083125
R5372 VSS.n1666 VSS.n1665 0.0083125
R5373 VSS.n1680 VSS.n1679 0.0083125
R5374 VSS.n1693 VSS.n1692 0.0083125
R5375 VSS.n1707 VSS.n1706 0.0083125
R5376 VSS.n1723 VSS.n1722 0.0083125
R5377 VSS.n1737 VSS.n1736 0.0083125
R5378 VSS.n1751 VSS.n1750 0.0083125
R5379 VSS.n1754 VSS.n1753 0.0083125
R5380 VSS.n1774 VSS.n1773 0.0083125
R5381 VSS.n1860 VSS.n1859 0.0083125
R5382 VSS.n1976 VSS.n917 0.0083125
R5383 VSS.n2361 VSS.n2340 0.0083125
R5384 VSS.n2338 VSS.n2326 0.0083125
R5385 VSS.n2324 VSS.n2323 0.0083125
R5386 VSS.n2321 VSS.n2309 0.0083125
R5387 VSS.n2307 VSS.n2293 0.0083125
R5388 VSS.n2291 VSS.n2279 0.0083125
R5389 VSS.n2277 VSS.n2265 0.0083125
R5390 VSS.n2263 VSS.n2262 0.0083125
R5391 VSS.n2260 VSS.n2237 0.0083125
R5392 VSS.n2764 VSS.n2763 0.0083125
R5393 VSS.n4756 VSS.n4755 0.0083125
R5394 VSS.n3767 VSS.n3757 0.0083125
R5395 VSS.n3451 VSS.n3450 0.0083125
R5396 VSS.n1192 VSS.n1183 0.0083125
R5397 VSS.n1189 VSS.n1184 0.0083125
R5398 VSS.n1598 VSS.n1596 0.0083125
R5399 VSS.n1908 VSS.n1906 0.0083125
R5400 VSS.n3032 VSS.n3026 0.0083125
R5401 VSS.n3046 VSS.n3041 0.0083125
R5402 VSS.n3069 VSS.n3068 0.0083125
R5403 VSS.n3208 VSS.n3199 0.0083125
R5404 VSS.n3205 VSS.n3200 0.0083125
R5405 VSS.n481 VSS.n480 0.0083125
R5406 VSS VSS.n430 0.0083125
R5407 VSS.n2875 VSS.n2870 0.0083125
R5408 VSS.n4095 VSS.n4094 0.0083125
R5409 VSS.n3938 VSS.n3936 0.0083125
R5410 VSS.n4652 VSS.n4651 0.00827766
R5411 VSS.n4983 VSS.n4982 0.0081375
R5412 VSS VSS.n5084 0.00763422
R5413 VSS.n1122 VSS.n1121 0.00725676
R5414 VSS.n4117 VSS.n4116 0.00725676
R5415 VSS.n1286 VSS.n1263 0.00725676
R5416 VSS.n2034 VSS.n2033 0.00725676
R5417 VSS.n3257 VSS.n3256 0.00725676
R5418 VSS.n4616 VSS.n4611 0.00725676
R5419 VSS.n309 VSS.n308 0.00725676
R5420 VSS.n642 VSS.n640 0.00725676
R5421 VSS.n2983 VSS.n2967 0.00725676
R5422 VSS.n4683 VSS.n4682 0.00725676
R5423 VSS.n1233 VSS.n1214 0.00701042
R5424 VSS.n1622 VSS.n1621 0.00701042
R5425 VSS.n1649 VSS.n1624 0.00701042
R5426 VSS.n2805 VSS.n2803 0.00701042
R5427 VSS.n3338 VSS.n3336 0.00701042
R5428 VSS.n3584 VSS.n3578 0.00701042
R5429 VSS.n1520 VSS.n1519 0.00701042
R5430 VSS.n99 VSS.n98 0.00701042
R5431 VSS.n259 VSS.n250 0.00701042
R5432 VSS.n256 VSS.n251 0.00701042
R5433 VSS.n5012 VSS.n5011 0.00701042
R5434 VSS.n2910 VSS.n2909 0.00701042
R5435 VSS.n3134 VSS.n3133 0.00701042
R5436 VSS.n3181 VSS.n3172 0.00701042
R5437 VSS.n3178 VSS.n3173 0.00701042
R5438 VSS.n4185 VSS.n4184 0.00701042
R5439 VSS.n4227 VSS.n4153 0.00701042
R5440 VSS.n4236 VSS.n4235 0.00701042
R5441 VSS.n1336 VSS.n1331 0.00701042
R5442 VSS.n1927 VSS.n1925 0.00701042
R5443 VSS.n4098 VSS.n4097 0.00623493
R5444 VSS.n4444 VSS.n4443 0.00623493
R5445 VSS.n3344 VSS.n3343 0.00623493
R5446 VSS.n3592 VSS.n3590 0.00623493
R5447 VSS.n3110 VSS.n3109 0.00623493
R5448 VSS.n3162 VSS.n3161 0.00623493
R5449 VSS.n3184 VSS.n3183 0.00623493
R5450 VSS.n4615 VSS.n4613 0.00623493
R5451 VSS.n3717 VSS.n3716 0.00623493
R5452 VSS.n3743 VSS.n3742 0.00623493
R5453 VSS.n3908 VSS.n3907 0.00623493
R5454 VSS.n573 VSS.n572 0.00623493
R5455 VSS.n4953 VSS.n4952 0.00623493
R5456 VSS.n4975 VSS.n4974 0.00623493
R5457 VSS.n2758 VSS.n2757 0.00623493
R5458 VSS.n4806 VSS.n4804 0.00623493
R5459 VSS.n239 VSS.n238 0.00623493
R5460 VSS.n2521 VSS.n2520 0.00623493
R5461 VSS.n2095 VSS.n2094 0.00623493
R5462 VSS.n2099 VSS.n2098 0.00623493
R5463 VSS.n836 VSS.n835 0.00623493
R5464 VSS.n2504 VSS.n2503 0.00623493
R5465 VSS.n809 VSS.n808 0.00623493
R5466 VSS.n4686 VSS.n4685 0.00623493
R5467 VSS.n4585 VSS.n4584 0.00623493
R5468 VSS.n3362 VSS.n3361 0.00623493
R5469 VSS.n1019 VSS.n1017 0.00614727
R5470 VSS.n2524 VSS.n2523 0.00590289
R5471 VSS.n636 VSS.n635 0.00590289
R5472 VSS.n2144 VSS.n638 0.00590289
R5473 VSS.n644 VSS.n643 0.00590289
R5474 VSS.n650 VSS.n649 0.00590289
R5475 VSS.n784 VSS.n783 0.00590289
R5476 VSS.n263 VSS.n262 0.00590289
R5477 VSS.n142 VSS.n141 0.00590289
R5478 VSS.n214 VSS.n213 0.00590289
R5479 VSS.n162 VSS.n161 0.00590289
R5480 VSS.n182 VSS.n181 0.00590289
R5481 VSS.n569 VSS.n568 0.00590289
R5482 VSS.n2723 VSS.n2722 0.00590289
R5483 VSS.n695 VSS.n694 0.00590289
R5484 VSS.n4832 VSS.n4831 0.00590289
R5485 VSS.n4801 VSS.n4800 0.00590289
R5486 VSS.n4848 VSS.n4847 0.00590289
R5487 VSS.n4946 VSS.n4945 0.00590289
R5488 VSS.n4866 VSS.n4865 0.00590289
R5489 VSS.n4759 VSS.n4758 0.00590289
R5490 VSS.n3441 VSS.n3440 0.00590289
R5491 VSS.n4648 VSS.n4647 0.00590289
R5492 VSS.n3772 VSS.n3771 0.00590289
R5493 VSS.n4689 VSS.n4688 0.00590289
R5494 VSS.n4637 VSS.n4636 0.00590289
R5495 VSS.n2887 VSS.n2886 0.00590289
R5496 VSS.n4004 VSS.n2888 0.00590289
R5497 VSS.n3129 VSS.n3128 0.00590289
R5498 VSS.n3079 VSS.n3078 0.00590289
R5499 VSS.n3086 VSS.n3085 0.00590289
R5500 VSS.n3486 VSS.n3485 0.00590289
R5501 VSS.n3420 VSS.n3352 0.00590289
R5502 VSS.n4309 VSS.n4308 0.00590289
R5503 VSS.n3554 VSS.n3553 0.00590289
R5504 VSS.n3588 VSS.n3587 0.00590289
R5505 VSS.n3883 VSS.n3882 0.00590289
R5506 VSS.n3973 VSS.n3972 0.00590289
R5507 VSS.n4119 VSS.n4118 0.00590289
R5508 VSS.n4451 VSS.n4450 0.00590289
R5509 VSS.n4339 VSS.n4338 0.00590289
R5510 VSS.n4371 VSS.n4370 0.00590289
R5511 VSS.n3942 VSS.n3941 0.00590289
R5512 VSS.n1074 VSS.n1049 0.00570833
R5513 VSS.n2718 VSS.n2714 0.00570833
R5514 VSS.n4681 VSS.n4680 0.00570833
R5515 VSS.n1284 VSS.n1274 0.00570833
R5516 VSS.n2032 VSS.n2031 0.00570833
R5517 VSS.n5058 VSS.n5053 0.00570833
R5518 VSS.n311 VSS.n310 0.00570833
R5519 VSS.n4934 VSS.n4933 0.00570833
R5520 VSS.n2974 VSS.n2968 0.00570833
R5521 VSS.n2982 VSS.n2981 0.00570833
R5522 VSS.n4544 VSS.n4542 0.00570833
R5523 VSS.n3245 VSS.n3240 0.00570833
R5524 VSS.n3255 VSS.n3254 0.00570833
R5525 VSS.n4334 VSS.n4332 0.00570833
R5526 VSS.n4204 VSS.n4202 0.00570833
R5527 VSS.n1119 VSS.n1118 0.00570833
R5528 VSS.n853 VSS.n849 0.00570833
R5529 VSS.n2491 VSS.n2490 0.00570833
R5530 VSS.n2487 VSS.n2482 0.00570833
R5531 VSS.n690 VSS.n686 0.00570833
R5532 VSS.n4618 VSS.n4617 0.00570833
R5533 VSS.n4570 VSS.n4568 0.00570833
R5534 VSS.n4115 VSS.n4114 0.00570833
R5535 VSS.n1888 VSS.n1872 0.00556757
R5536 VSS.n5063 VSS.n5027 0.00556757
R5537 VSS.n54 VSS.n53 0.00556757
R5538 VSS.n3108 VSS.n3090 0.00556757
R5539 VSS.n3906 VSS.n3885 0.00556757
R5540 VSS.n1167 VSS.n1128 0.00556757
R5541 VSS.n4944 VSS.n4872 0.00556757
R5542 VSS.n4973 VSS.n4956 0.00556757
R5543 VSS.n4830 VSS.n429 0.00556757
R5544 VSS.n160 VSS.n159 0.00556757
R5545 VSS.n237 VSS.n220 0.00556757
R5546 VSS.n2889 VSS.n426 0.00490625
R5547 VSS.n2913 VSS.n2890 0.00490625
R5548 VSS.n2914 VSS.n2913 0.00490625
R5549 VSS.n2938 VSS.n2915 0.00490625
R5550 VSS.n2939 VSS.n2938 0.00490625
R5551 VSS.n2961 VSS.n2940 0.00490625
R5552 VSS.n2962 VSS.n2961 0.00490625
R5553 VSS.n2985 VSS.n2963 0.00490625
R5554 VSS.n2986 VSS.n2985 0.00490625
R5555 VSS.n3012 VSS.n2987 0.00490625
R5556 VSS.n3013 VSS.n3012 0.00490625
R5557 VSS.n3035 VSS.n3014 0.00490625
R5558 VSS.n3036 VSS.n3035 0.00490625
R5559 VSS.n3073 VSS.n3037 0.00490625
R5560 VSS.n5022 VSS.n5021 0.00490625
R5561 VSS.n5021 VSS.n5020 0.00490625
R5562 VSS.n5019 VSS.n5018 0.00490625
R5563 VSS.n5018 VSS.n5017 0.00490625
R5564 VSS.n5016 VSS.n5015 0.00490625
R5565 VSS.n5015 VSS.n4995 0.00490625
R5566 VSS.n4994 VSS.n4993 0.00490625
R5567 VSS.n4993 VSS.n4992 0.00490625
R5568 VSS.n4991 VSS.n4990 0.00490625
R5569 VSS.n4990 VSS.n4989 0.00490625
R5570 VSS.n4988 VSS.n4987 0.00490625
R5571 VSS.n4987 VSS.n4986 0.00490625
R5572 VSS.n4985 VSS.n4984 0.00490625
R5573 VSS.n4984 VSS.n4983 0.00490625
R5574 VSS.n4189 VSS.n3262 0.00490625
R5575 VSS.n4190 VSS.n4189 0.00490625
R5576 VSS.n4214 VSS.n4191 0.00490625
R5577 VSS.n4215 VSS.n4214 0.00490625
R5578 VSS.n4221 VSS.n4216 0.00490625
R5579 VSS.n4222 VSS.n4221 0.00490625
R5580 VSS.n4554 VSS.n4553 0.00490625
R5581 VSS.n4553 VSS.n4515 0.00490625
R5582 VSS.n4514 VSS.n4513 0.00490625
R5583 VSS.n4513 VSS.n4493 0.00490625
R5584 VSS.n4492 VSS.n4491 0.00490625
R5585 VSS.n4491 VSS.n4490 0.00490625
R5586 VSS.n4489 VSS.n4488 0.00490625
R5587 VSS.n4488 VSS.n4487 0.00490625
R5588 VSS.n4486 VSS.n4485 0.00490625
R5589 VSS.n4485 VSS.n4464 0.00490625
R5590 VSS.n4463 VSS.n4462 0.00490625
R5591 VSS.n4462 VSS.n4461 0.00490625
R5592 VSS.n4460 VSS.n4459 0.00490625
R5593 VSS.n4459 VSS.n4458 0.00490625
R5594 VSS.n1608 VSS.n1607 0.00490625
R5595 VSS.n1607 VSS.n1606 0.00490625
R5596 VSS.n1605 VSS.n1604 0.00490625
R5597 VSS.n1604 VSS.n1573 0.00490625
R5598 VSS.n1572 VSS.n1571 0.00490625
R5599 VSS.n1571 VSS.n1570 0.00490625
R5600 VSS.n1569 VSS.n1568 0.00490625
R5601 VSS.n1568 VSS.n1567 0.00490625
R5602 VSS.n1566 VSS.n1565 0.00490625
R5603 VSS.n1565 VSS.n1564 0.00490625
R5604 VSS.n1563 VSS.n1562 0.00490625
R5605 VSS.n1562 VSS.n1561 0.00490625
R5606 VSS.n1560 VSS.n1559 0.00490625
R5607 VSS.n1559 VSS.n1558 0.00490625
R5608 VSS.n5082 VSS.n5081 0.00490625
R5609 VSS.n5081 VSS.n5080 0.00490625
R5610 VSS.n5079 VSS.n5078 0.00490625
R5611 VSS.n5078 VSS.n5077 0.00490625
R5612 VSS.n5076 VSS.n5075 0.00490625
R5613 VSS.n5075 VSS.n5074 0.00490625
R5614 VSS.n5073 VSS.n5072 0.00490625
R5615 VSS.n5072 VSS.n5071 0.00490625
R5616 VSS.n5070 VSS.n5069 0.00490625
R5617 VSS.n5069 VSS.n5068 0.00490625
R5618 VSS.n5067 VSS.n5066 0.00490625
R5619 VSS.n5066 VSS.n5025 0.00490625
R5620 VSS.n4225 VSS.n4224 0.00483277
R5621 VSS.n2094 VSS.n2093 0.00480456
R5622 VSS.n2520 VSS.n2519 0.00480456
R5623 VSS.n2100 VSS.n2099 0.00480456
R5624 VSS.n572 VSS.n571 0.00480456
R5625 VSS.n3361 VSS.n3360 0.00480456
R5626 VSS.n1016 VSS.n1015 0.00450332
R5627 VSS.n1166 VSS.n1144 0.00440625
R5628 VSS.n1159 VSS.n1158 0.00440625
R5629 VSS.n1776 VSS 0.00440625
R5630 VSS.n1843 VSS.n1842 0.00440625
R5631 VSS.n2816 VSS.n2811 0.00440625
R5632 VSS.n3905 VSS.n3892 0.00440625
R5633 VSS.n3894 VSS.n3893 0.00440625
R5634 VSS.n3549 VSS.n3547 0.00440625
R5635 VSS.n2019 VSS.n2013 0.00440625
R5636 VSS.n49 VSS.n44 0.00440625
R5637 VSS.n56 VSS.n55 0.00440625
R5638 VSS.n5061 VSS.n5032 0.00440625
R5639 VSS.n5046 VSS.n5044 0.00440625
R5640 VSS.n236 VSS.n230 0.00440625
R5641 VSS.n150 VSS.n145 0.00440625
R5642 VSS.n158 VSS.n157 0.00440625
R5643 VSS.n304 VSS.n299 0.00440625
R5644 VSS.n4964 VSS.n4957 0.00440625
R5645 VSS.n4972 VSS.n4971 0.00440625
R5646 VSS.n4942 VSS.n4877 0.00440625
R5647 VSS.n3107 VSS.n3106 0.00440625
R5648 VSS.n3156 VSS.n3151 0.00440625
R5649 VSS.n3232 VSS.n3229 0.00440625
R5650 VSS.n1304 VSS.n1301 0.00440625
R5651 VSS.n1887 VSS.n1886 0.00440625
R5652 VSS.n4828 VSS.n430 0.00440625
R5653 VSS.n478 VSS.n477 0.00440625
R5654 VSS.n4107 VSS.n4102 0.00440625
R5655 VSS.n5024 VSS.n5023 0.004025
R5656 VSS.n1013 VSS.n1011 0.00393951
R5657 VSS.n4220 VSS.n4219 0.00390995
R5658 VSS.n1419 VSS.n1418 0.00390995
R5659 VSS.n1470 VSS.n1469 0.00390995
R5660 VSS.n2058 VSS.n2057 0.00390995
R5661 VSS.n1807 VSS.n1806 0.00390995
R5662 VSS.n2005 VSS.n2004 0.00390995
R5663 VSS.n2044 VSS.n2043 0.00390995
R5664 VSS.n2366 VSS.n2365 0.00390995
R5665 VSS.n494 VSS.n493 0.00390995
R5666 VSS.n386 VSS.n385 0.00390995
R5667 VSS.n134 VSS.n120 0.00387838
R5668 VSS.n1440 VSS.n1422 0.00387838
R5669 VSS.n3160 VSS.n3113 0.00387838
R5670 VSS.n354 VSS.n337 0.00387838
R5671 VSS.n634 VSS.n633 0.00387838
R5672 VSS.n2145 VSS.n2142 0.00387838
R5673 VSS.n5084 VSS.n5083 0.00373125
R5674 VSS.n1095 VSS.n1094 0.00310928
R5675 VSS.n1777 VSS.n1775 0.00310417
R5676 VSS.n1795 VSS.n944 0.00310417
R5677 VSS.n944 VSS.n943 0.00310417
R5678 VSS.n942 VSS.n941 0.00310417
R5679 VSS.n940 VSS.n939 0.00310417
R5680 VSS.n1826 VSS.n1814 0.00310417
R5681 VSS.n1859 VSS.n1858 0.00310417
R5682 VSS.n1841 VSS.n1840 0.00310417
R5683 VSS.n902 VSS.n890 0.00310417
R5684 VSS.n917 VSS.n905 0.00310417
R5685 VSS.n2000 VSS.n1979 0.00310417
R5686 VSS.n2146 VSS.n2140 0.00310417
R5687 VSS VSS.n2102 0.00310417
R5688 VSS.n632 VSS.n631 0.00310417
R5689 VSS.n562 VSS.n557 0.00310417
R5690 VSS.n3317 VSS.n3313 0.00310417
R5691 VSS.n1439 VSS.n1428 0.00310417
R5692 VSS.n1435 VSS.n1429 0.00310417
R5693 VSS VSS.n1476 0.00310417
R5694 VSS.n132 VSS.n125 0.00310417
R5695 VSS.n329 VSS.n327 0.00310417
R5696 VSS.n352 VSS.n346 0.00310417
R5697 VSS.n4897 VSS.n4895 0.00310417
R5698 VSS.n2929 VSS.n2925 0.00310417
R5699 VSS.n3050 VSS.n3049 0.00310417
R5700 VSS.n3159 VSS.n3145 0.00310417
R5701 VSS.n803 VSS.n798 0.00310417
R5702 VSS.n4457 VSS.n3262 0.00299688
R5703 VSS.n1803 VSS.n1802 0.00287807
R5704 VSS.n4982 VSS.n426 0.00270313
R5705 VSS.n4555 VSS.n3073 0.00270313
R5706 VSS.n4401 VSS.n4400 0.00246557
R5707 VSS.n3266 VSS.n3265 0.00246557
R5708 VSS.n985 VSS.n979 0.00225053
R5709 VSS.n886 VSS.n885 0.00218919
R5710 VSS.n4511 VSS.n4497 0.00218919
R5711 VSS.n3084 VSS.n3083 0.00218919
R5712 VSS.n3077 VSS.n3075 0.00218919
R5713 VSS.n4635 VSS.n4634 0.00218919
R5714 VSS.n4864 VSS.n4863 0.00218919
R5715 VSS.n567 VSS.n498 0.00218919
R5716 VSS.n648 VSS.n646 0.00218919
R5717 VSS.n807 VSS.n791 0.00218919
R5718 VSS.n4005 VSS.n4002 0.00218919
R5719 VSS.n4347 VSS.n4345 0.00213281
R5720 VSS.n3558 VSS.n3556 0.00213281
R5721 VSS.n4842 VSS.n4840 0.00213281
R5722 VSS.n4778 VSS.n4776 0.00213281
R5723 VSS.n4764 VSS.n4762 0.00213281
R5724 VSS.n186 VSS.n184 0.00213281
R5725 VSS.n3491 VSS.n3490 0.00213281
R5726 VSS.n1966 VSS.n1965 0.00183767
R5727 VSS.n2061 VSS.n2060 0.00182115
R5728 VSS.n1059 VSS.n1049 0.00180208
R5729 VSS.n1088 VSS.n1087 0.00180208
R5730 VSS.n1142 VSS.n1130 0.00180208
R5731 VSS.n1160 VSS.n1159 0.00180208
R5732 VSS.n1212 VSS.n1202 0.00180208
R5733 VSS.n1218 VSS.n1217 0.00180208
R5734 VSS.n973 VSS.n961 0.00180208
R5735 VSS.n1623 VSS.n1622 0.00180208
R5736 VSS.n2235 VSS.n2076 0.00180208
R5737 VSS.n2223 VSS.n2222 0.00180208
R5738 VSS.n2220 VSS.n2208 0.00180208
R5739 VSS.n2206 VSS.n2194 0.00180208
R5740 VSS.n2192 VSS.n2177 0.00180208
R5741 VSS.n2175 VSS.n2163 0.00180208
R5742 VSS.n2161 VSS.n2160 0.00180208
R5743 VSS.n2160 VSS.n2159 0.00180208
R5744 VSS.n2138 VSS.n2126 0.00180208
R5745 VSS.n2124 VSS.n2103 0.00180208
R5746 VSS.n609 VSS.n608 0.00180208
R5747 VSS.n2568 VSS.n2567 0.00180208
R5748 VSS.n2585 VSS.n2584 0.00180208
R5749 VSS.n2598 VSS.n2597 0.00180208
R5750 VSS.n2612 VSS.n2611 0.00180208
R5751 VSS.n2629 VSS.n2628 0.00180208
R5752 VSS.n2643 VSS.n2642 0.00180208
R5753 VSS.n2656 VSS.n2655 0.00180208
R5754 VSS.n2670 VSS.n2669 0.00180208
R5755 VSS.n2690 VSS.n2689 0.00180208
R5756 VSS.n2754 VSS.n2747 0.00180208
R5757 VSS.n565 VSS.n510 0.00180208
R5758 VSS.n25 VSS.n21 0.00180208
R5759 VSS.n4862 VSS.n4861 0.00180208
R5760 VSS.n3059 VSS.n3058 0.00180208
R5761 VSS.n4531 VSS.n4525 0.00180208
R5762 VSS.n4510 VSS.n4509 0.00180208
R5763 VSS.n4476 VSS.n4474 0.00180208
R5764 VSS.n876 VSS.n871 0.00180208
R5765 VSS.n884 VSS.n883 0.00180208
R5766 VSS.n2458 VSS.n2457 0.00180208
R5767 VSS.n2466 VSS.n2465 0.00180208
R5768 VSS.n806 VSS.n797 0.00180208
R5769 VSS.n4633 VSS.n4632 0.00180208
R5770 VSS.n4007 VSS.n4006 0.00180208
R5771 VSS.n1557 VSS.n1556 0.00168904
R5772 VSS.n1915 VSS.n1914 0.00167252
R5773 VSS.n1198 VSS.n1197 0.00163949
R5774 VSS.n495 VSS.n490 0.00163288
R5775 VSS.n2038 VSS.n2037 0.00160647
R5776 VSS.n1609 VSS.n1608 0.00152813
R5777 VSS.n575 VSS.n574 0.00144949
R5778 VSS.n4555 VSS.n3190 0.00144949
R5779 VSS.n5023 VSS.n271 0.00141558
R5780 VSS.n4982 VSS.n4981 0.00141558
R5781 VSS.n1610 VSS.n1609 0.00139178
R5782 VSS.n4978 VSS.n4977 0.00138167
R5783 VSS.n4870 VSS.n4869 0.00138167
R5784 VSS.n3589 VSS.n3322 0.00138167
R5785 VSS.n3563 VSS.n3562 0.00138167
R5786 VSS.n3744 VSS.n3263 0.00138167
R5787 VSS.n3910 VSS.n3909 0.00138167
R5788 VSS.n4687 VSS.n2808 0.00134776
R5789 VSS.n4646 VSS.n4645 0.00134776
R5790 VSS.n496 VSS.n495 0.00131643
R5791 VSS.n4457 VSS.n4456 0.00131385
R5792 VSS.n4779 VSS.n4774 0.00127994
R5793 VSS.n4834 VSS.n4833 0.00127994
R5794 VSS.n3186 VSS.n3185 0.00127994
R5795 VSS.n3127 VSS.n3126 0.00127994
R5796 VSS.n4453 VSS.n4452 0.00127994
R5797 VSS.n4348 VSS.n4343 0.00127994
R5798 VSS.n2724 VSS.n580 0.00121212
R5799 VSS.n4766 VSS.n4765 0.00121212
R5800 VSS.n1291 VSS.n1290 0.0011936
R5801 VSS.n4639 VSS.n4638 0.00117821
R5802 VSS.n4586 VSS.n4559 0.00117821
R5803 VSS.n2096 VSS.n2091 0.0011443
R5804 VSS.n2516 VSS.n2515 0.0011443
R5805 VSS.n2506 VSS.n2505 0.0011443
R5806 VSS.n789 VSS.n788 0.0011443
R5807 VSS.n265 VSS.n264 0.0011443
R5808 VSS.n215 VSS.n192 0.0011443
R5809 VSS.n3943 VSS.n3916 0.00111039
R5810 VSS.n4311 VSS.n4310 0.00111039
R5811 VSS.n3351 VSS.n3350 0.00104257
R5812 VSS.n3363 VSS.n3358 0.00104257
R5813 VSS.n1008 VSS.n985 0.000995432
R5814 VSS.n1042 VSS.n979 0.000995432
R5815 VSS.n1043 VSS.n1042 0.000995432
R5816 VSS.n1093 VSS.n1044 0.000995432
R5817 VSS.n1094 VSS.n1093 0.000995432
R5818 VSS.n1196 VSS.n1171 0.000995432
R5819 VSS.n1197 VSS.n1196 0.000995432
R5820 VSS.n1289 VSS.n1260 0.000995432
R5821 VSS.n1290 VSS.n1289 0.000995432
R5822 VSS.n1808 VSS.n1803 0.000995432
R5823 VSS.n1809 VSS.n1808 0.000995432
R5824 VSS.n1865 VSS.n1810 0.000995432
R5825 VSS.n1891 VSS.n1890 0.000995432
R5826 VSS.n1913 VSS.n1892 0.000995432
R5827 VSS.n1914 VSS.n1913 0.000995432
R5828 VSS.n1967 VSS.n1966 0.000995432
R5829 VSS.n2036 VSS.n2009 0.000995432
R5830 VSS.n2037 VSS.n2036 0.000995432
R5831 VSS.n2059 VSS.n2054 0.000995432
R5832 VSS.n2060 VSS.n2059 0.000995432
R5833 VSS.n2368 VSS.n30 0.000995432
R5834 VSS.n1238 VSS.n1199 0.000978918
R5835 VSS.n1258 VSS.n1257 0.000978918
R5836 VSS.n1260 VSS.n1259 0.000978918
R5837 VSS.n2367 VSS.n2062 0.000978918
R5838 VSS.n2371 VSS.n2370 0.000978918
R5839 VSS.n1415 VSS.n1292 0.000962403
R5840 VSS.n1612 VSS.n1611 0.000962403
R5841 VSS.n1916 VSS.n1915 0.000962403
R5842 VSS.n1971 VSS.n1939 0.000962403
R5843 VSS.n1010 VSS.n1009 0.000945889
R5844 VSS.n1866 VSS.n1865 0.000945889
R5845 VSS.n1890 VSS.n1867 0.000945889
R5846 VSS.n2045 VSS.n2039 0.000929375
R5847 VSS.n2053 VSS.n2052 0.000929375
R5848 VSS.n1125 VSS.n1096 0.00091286
R5849 VSS.n1170 VSS.n1169 0.00091286
R5850 VSS.n1965 VSS.n1964 0.000879831
R5851 VSS.n2006 VSS.n888 0.000879831
R5852 VSS.n2008 VSS.n2007 0.000879831
R5853 VSS.n1969 VSS.n1968 0.000863317
R5854 VSS.n1810 VSS.n1809 0.000846803
R5855 VSS.n2369 VSS.n2368 0.000830288
R5856 VSS.n1556 VSS.n1555 0.000797259
R5857 VSS.n1553 VSS.n921 0.000797259
R5858 VSS.n1801 VSS.n1800 0.000797259
R5859 VSS VSS.n5079 0.00079375
R5860 VSS.n1892 VSS.n1891 0.000731202
R5861 VSS.n3350 VSS.n3349 0.000703463
R5862 VSS.n3487 VSS.n3363 0.000703463
R5863 VSS.n3356 VSS.n3355 0.000703463
R5864 VSS.n4641 VSS.n4640 0.000703463
R5865 VSS.n4588 VSS.n4587 0.000703463
R5866 VSS.n4558 VSS.n4557 0.000703463
R5867 VSS.n3913 VSS.n3912 0.000703463
R5868 VSS.n3974 VSS.n3943 0.000703463
R5869 VSS.n4312 VSS.n4311 0.000703463
R5870 VSS.n266 VSS.n265 0.000669553
R5871 VSS.n216 VSS.n215 0.000669553
R5872 VSS.n579 VSS.n578 0.000669553
R5873 VSS.n4760 VSS.n2759 0.000669553
R5874 VSS.n4768 VSS.n4767 0.000669553
R5875 VSS.n3349 VSS.n3348 0.000669553
R5876 VSS.n3488 VSS.n3487 0.000669553
R5877 VSS.n3357 VSS.n3356 0.000669553
R5878 VSS.n4456 VSS.n4455 0.000669553
R5879 VSS.n4452 VSS.n4445 0.000669553
R5880 VSS.n4343 VSS.n4342 0.000669553
R5881 VSS.n2508 VSS.n2507 0.000635642
R5882 VSS.n837 VSS.n810 0.000635642
R5883 VSS.n786 VSS.n785 0.000635642
R5884 VSS.n3354 VSS.n3353 0.000635642
R5885 VSS.n4687 VSS.n2809 0.000635642
R5886 VSS.n4645 VSS.n4644 0.000635642
R5887 VSS.n3188 VSS.n3187 0.000635642
R5888 VSS.n3163 VSS.n3111 0.000635642
R5889 VSS.n3124 VSS.n3123 0.000635642
R5890 VSS.n3559 VSS.n3263 0.000635642
R5891 VSS.n3909 VSS.n3744 0.000635642
R5892 VSS.n3911 VSS.n3910 0.000635642
R5893 VSS.n1968 VSS.n1967 0.000632115
R5894 VSS.n5084 VSS.n30 0.000632115
R5895 VSS.n1554 VSS.n1553 0.000615601
R5896 VSS.n1800 VSS.n1799 0.000615601
R5897 VSS.n1964 VSS.n888 0.000615601
R5898 VSS.n2007 VSS.n2006 0.000615601
R5899 VSS.n2089 VSS.n2088 0.000601732
R5900 VSS.n2090 VSS.n2089 0.000601732
R5901 VSS.n2091 VSS.n2090 0.000601732
R5902 VSS.n2097 VSS.n637 0.000601732
R5903 VSS.n2522 VSS.n637 0.000601732
R5904 VSS.n2522 VSS.n2516 0.000601732
R5905 VSS.n2514 VSS.n2513 0.000601732
R5906 VSS.n2513 VSS.n2512 0.000601732
R5907 VSS.n2512 VSS.n2511 0.000601732
R5908 VSS.n2510 VSS.n2509 0.000601732
R5909 VSS.n2507 VSS.n2506 0.000601732
R5910 VSS.n2505 VSS.n838 0.000601732
R5911 VSS.n810 VSS.n789 0.000601732
R5912 VSS.n788 VSS.n787 0.000601732
R5913 VSS.n785 VSS.n136 0.000601732
R5914 VSS.n4773 VSS.n4772 0.000601732
R5915 VSS.n4803 VSS.n427 0.000601732
R5916 VSS.n4837 VSS.n4836 0.000601732
R5917 VSS.n3488 VSS.n3351 0.000601732
R5918 VSS.n3358 VSS.n3357 0.000601732
R5919 VSS.n1970 VSS.n1969 0.000599086
R5920 VSS.n1096 VSS.n1095 0.000582572
R5921 VSS.n1169 VSS.n1125 0.000582572
R5922 VSS.n1171 VSS.n1170 0.000582572
R5923 VSS.n1555 VSS.n1554 0.000582572
R5924 VSS.n1799 VSS.n921 0.000582572
R5925 VSS.n1802 VSS.n1801 0.000582572
R5926 VSS.n2097 VSS.n2096 0.000567821
R5927 VSS.n2515 VSS.n2514 0.000567821
R5928 VSS.n267 VSS.n266 0.000567821
R5929 VSS.n217 VSS.n216 0.000567821
R5930 VSS.n188 VSS.n187 0.000567821
R5931 VSS.n574 VSS.n496 0.000567821
R5932 VSS.n576 VSS.n575 0.000567821
R5933 VSS.n578 VSS.n577 0.000567821
R5934 VSS.n580 VSS.n579 0.000567821
R5935 VSS.n2759 VSS.n2724 0.000567821
R5936 VSS.n4765 VSS.n4760 0.000567821
R5937 VSS.n4767 VSS.n4766 0.000567821
R5938 VSS.n4769 VSS.n4768 0.000567821
R5939 VSS.n4771 VSS.n4770 0.000567821
R5940 VSS.n4802 VSS.n4779 0.000567821
R5941 VSS.n4835 VSS.n4834 0.000567821
R5942 VSS.n4981 VSS.n4980 0.000567821
R5943 VSS.n4977 VSS.n4976 0.000567821
R5944 VSS.n4869 VSS.n4868 0.000567821
R5945 VSS.n4642 VSS.n4641 0.000567821
R5946 VSS.n4640 VSS.n4639 0.000567821
R5947 VSS.n4638 VSS.n4588 0.000567821
R5948 VSS.n4587 VSS.n4586 0.000567821
R5949 VSS.n4559 VSS.n4558 0.000567821
R5950 VSS.n4557 VSS.n4556 0.000567821
R5951 VSS.n3321 VSS.n3320 0.000567821
R5952 VSS.n3322 VSS.n3321 0.000567821
R5953 VSS.n3589 VSS.n3564 0.000567821
R5954 VSS.n3564 VSS.n3563 0.000567821
R5955 VSS.n3562 VSS.n3561 0.000567821
R5956 VSS.n3561 VSS.n3560 0.000567821
R5957 VSS.n3914 VSS.n3913 0.000567821
R5958 VSS.n3915 VSS.n3914 0.000567821
R5959 VSS.n3916 VSS.n3915 0.000567821
R5960 VSS.n4099 VSS.n3974 0.000567821
R5961 VSS.n4120 VSS.n4099 0.000567821
R5962 VSS.n4310 VSS.n4120 0.000567821
R5963 VSS.n4313 VSS.n4312 0.000567821
R5964 VSS.n4314 VSS.n4313 0.000567821
R5965 VSS.n4315 VSS.n4314 0.000567821
R5966 VSS.n2009 VSS.n2008 0.000566058
R5967 VSS.n2039 VSS.n2038 0.000566058
R5968 VSS.n2052 VSS.n2045 0.000566058
R5969 VSS.n2054 VSS.n2053 0.000566058
R5970 VSS.n1009 VSS.n1008 0.000549543
R5971 VSS.n1044 VSS.n1043 0.000549543
R5972 VSS.n1867 VSS.n1866 0.000549543
R5973 VSS.n2509 VSS.n2508 0.000533911
R5974 VSS.n838 VSS.n837 0.000533911
R5975 VSS.n787 VSS.n786 0.000533911
R5976 VSS.n271 VSS.n270 0.000533911
R5977 VSS.n270 VSS.n269 0.000533911
R5978 VSS.n269 VSS.n268 0.000533911
R5979 VSS.n268 VSS.n267 0.000533911
R5980 VSS.n264 VSS.n242 0.000533911
R5981 VSS.n242 VSS.n241 0.000533911
R5982 VSS.n241 VSS.n240 0.000533911
R5983 VSS.n240 VSS.n217 0.000533911
R5984 VSS.n192 VSS.n191 0.000533911
R5985 VSS.n191 VSS.n190 0.000533911
R5986 VSS.n190 VSS.n189 0.000533911
R5987 VSS.n189 VSS.n188 0.000533911
R5988 VSS.n4772 VSS.n4771 0.000533911
R5989 VSS.n4774 VSS.n4773 0.000533911
R5990 VSS.n4803 VSS.n4802 0.000533911
R5991 VSS.n4833 VSS.n427 0.000533911
R5992 VSS.n4836 VSS.n4835 0.000533911
R5993 VSS.n4838 VSS.n4837 0.000533911
R5994 VSS.n4980 VSS.n4979 0.000533911
R5995 VSS.n4979 VSS.n4978 0.000533911
R5996 VSS.n4976 VSS.n4947 0.000533911
R5997 VSS.n4947 VSS.n4870 0.000533911
R5998 VSS.n4868 VSS.n4867 0.000533911
R5999 VSS.n3353 VSS.n2808 0.000533911
R6000 VSS.n4646 VSS.n2809 0.000533911
R6001 VSS.n4644 VSS.n4643 0.000533911
R6002 VSS.n3190 VSS.n3189 0.000533911
R6003 VSS.n3189 VSS.n3188 0.000533911
R6004 VSS.n3187 VSS.n3186 0.000533911
R6005 VSS.n3185 VSS.n3164 0.000533911
R6006 VSS.n3164 VSS.n3163 0.000533911
R6007 VSS.n3127 VSS.n3111 0.000533911
R6008 VSS.n3126 VSS.n3125 0.000533911
R6009 VSS.n3125 VSS.n3124 0.000533911
R6010 VSS.n4455 VSS.n4454 0.000533911
R6011 VSS.n4454 VSS.n4453 0.000533911
R6012 VSS.n4445 VSS.n4349 0.000533911
R6013 VSS.n4349 VSS.n4348 0.000533911
R6014 VSS.n4342 VSS.n4341 0.000533911
R6015 VSS.n4341 VSS.n4340 0.000533911
R6016 VSS.n1292 VSS.n1291 0.000533029
R6017 VSS.n1612 VSS.n1415 0.000533029
R6018 VSS.n1611 VSS.n1610 0.000533029
R6019 VSS.n1939 VSS.n1916 0.000533029
R6020 VSS.n1971 VSS.n1970 0.000533029
R6021 VSS.n1199 VSS.n1198 0.000516514
R6022 VSS.n1257 VSS.n1238 0.000516514
R6023 VSS.n1259 VSS.n1258 0.000516514
R6024 VSS.n2062 VSS.n2061 0.000516514
R6025 VSS.n2371 VSS.n2367 0.000516514
R6026 VSS.n2370 VSS.n2369 0.000516514
R6027 VDD.n4125 VDD.t729 507.748
R6028 VDD.n1832 VDD.t697 500.865
R6029 VDD.n1975 VDD.t286 500.865
R6030 VDD.n983 VDD.t202 500.865
R6031 VDD.n449 VDD.t503 500.865
R6032 VDD.n3745 VDD.t288 500.865
R6033 VDD.n3940 VDD.t230 500.865
R6034 VDD.n4026 VDD.t699 500.865
R6035 VDD.n697 VDD.t5 500.865
R6036 VDD.n1075 VDD.t346 500.865
R6037 VDD.n2055 VDD.t49 500.865
R6038 VDD.n4655 VDD.t402 500.865
R6039 VDD.n4513 VDD.t494 500.865
R6040 VDD.n4402 VDD.t622 500.865
R6041 VDD.n1801 VDD.n1800 440.25
R6042 VDD.n1776 VDD.n1775 440.25
R6043 VDD.n972 VDD.n971 440.25
R6044 VDD.n438 VDD.n437 440.25
R6045 VDD.n3728 VDD.n3727 440.25
R6046 VDD.n3927 VDD.n3926 440.25
R6047 VDD.n4015 VDD.n4014 440.25
R6048 VDD.n720 VDD.n719 440.25
R6049 VDD.n1559 VDD.n1558 440.25
R6050 VDD.n2030 VDD.n2029 440.25
R6051 VDD.n4640 VDD.n4639 440.25
R6052 VDD.n4496 VDD.n4495 440.25
R6053 VDD.n4368 VDD.n4367 440.25
R6054 VDD.n4144 VDD.n4143 440.25
R6055 VDD.t99 VDD.n539 396.851
R6056 VDD.t96 VDD.n1146 396.851
R6057 VDD.t87 VDD.n2109 396.851
R6058 VDD.t129 VDD.n2497 396.851
R6059 VDD.t120 VDD.n2559 396.851
R6060 VDD.t102 VDD.n4443 396.851
R6061 VDD.t144 VDD.n4265 396.851
R6062 VDD.n531 VDD.t135 391.606
R6063 VDD.n1138 VDD.t114 391.606
R6064 VDD.n2101 VDD.t108 391.606
R6065 VDD.n2489 VDD.t90 391.606
R6066 VDD.n2551 VDD.t132 391.606
R6067 VDD.n4435 VDD.t123 391.606
R6068 VDD.n4257 VDD.t126 391.606
R6069 VDD.n1794 VDD.t75 374.084
R6070 VDD.n1722 VDD.t67 374.084
R6071 VDD.n3893 VDD.t570 374.084
R6072 VDD.n3695 VDD.t338 374.084
R6073 VDD.n2632 VDD.t177 374.084
R6074 VDD.n2597 VDD.t674 374.084
R6075 VDD.n4610 VDD.t572 374.084
R6076 VDD.n2354 VDD.t340 374.084
R6077 VDD.n1609 VDD.t77 374.084
R6078 VDD.n1172 VDD.t216 374.084
R6079 VDD.n511 VDD.t165 374.084
R6080 VDD.n294 VDD.t59 372.949
R6081 VDD.n3244 VDD.t71 372.949
R6082 VDD.n2676 VDD.t672 372.949
R6083 VDD.n3284 VDD.n3283 337.3
R6084 VDD.n3340 VDD.n3339 337.3
R6085 VDD.n3414 VDD.n3413 337.3
R6086 VDD.n3486 VDD.n3485 337.3
R6087 VDD.n2704 VDD.n2703 337.3
R6088 VDD.n402 VDD.n401 337.3
R6089 VDD.n840 VDD.n839 337.3
R6090 VDD.n1304 VDD.n1303 337.3
R6091 VDD.n1394 VDD.n1393 337.3
R6092 VDD.n2186 VDD.n2185 337.3
R6093 VDD.n2259 VDD.n2258 337.3
R6094 VDD.n2439 VDD.n2438 337.3
R6095 VDD.n4729 VDD.n4728 337.3
R6096 VDD.n4816 VDD.n4815 337.3
R6097 VDD.n450 VDD.t106 327.223
R6098 VDD.n984 VDD.t94 327.223
R6099 VDD.n1976 VDD.t148 327.223
R6100 VDD.n1833 VDD.t139 327.223
R6101 VDD.n3741 VDD.t118 327.223
R6102 VDD.n3938 VDD.t112 327.223
R6103 VDD.n4027 VDD.t142 327.223
R6104 VDD.n3248 VDD.n3247 312.132
R6105 VDD.n3991 VDD.n3987 312.132
R6106 VDD.n3903 VDD.n3899 312.132
R6107 VDD.n3704 VDD.n3703 312.132
R6108 VDD.n948 VDD.n944 312.132
R6109 VDD.n1733 VDD.n1729 312.132
R6110 VDD.n1796 VDD.n1795 312.132
R6111 VDD.n2628 VDD.n2627 312.132
R6112 VDD.n2593 VDD.n2592 312.132
R6113 VDD.n4617 VDD.n4616 312.132
R6114 VDD.n2345 VDD.n180 312.132
R6115 VDD.n1596 VDD.n1533 312.132
R6116 VDD.n1074 VDD.n1073 312.132
R6117 VDD.n502 VDD.n496 312.132
R6118 VDD.n1790 VDD.n1786 307.212
R6119 VDD.n3876 VDD.n3872 307.212
R6120 VDD.n3678 VDD.n3674 307.212
R6121 VDD.n4097 VDD.n4093 307.13
R6122 VDD.n4274 VDD.n4273 306.985
R6123 VDD.n4452 VDD.n4451 306.985
R6124 VDD.n2546 VDD.n2545 306.985
R6125 VDD.n2485 VDD.n2484 306.985
R6126 VDD.n2118 VDD.n2117 306.985
R6127 VDD.n1155 VDD.n1154 306.985
R6128 VDD.n527 VDD.n526 306.985
R6129 VDD.n1043 VDD.n1042 306.142
R6130 VDD.n630 VDD.n629 306.142
R6131 VDD.n3600 VDD.n3599 306.142
R6132 VDD.n2471 VDD.n2467 305.529
R6133 VDD.n1785 VDD.n1781 305.529
R6134 VDD.n1000 VDD.n996 305.529
R6135 VDD.n4043 VDD.n4039 305.529
R6136 VDD.n3955 VDD.n3951 305.529
R6137 VDD.n3802 VDD.n3798 305.529
R6138 VDD.n466 VDD.n462 305.529
R6139 VDD.n2642 VDD.n2638 305.529
R6140 VDD.n4672 VDD.n4668 305.529
R6141 VDD.n2009 VDD.n2005 305.529
R6142 VDD.n1104 VDD.n1100 305.529
R6143 VDD.n684 VDD.n680 305.529
R6144 VDD.n4340 VDD.n4339 304.459
R6145 VDD.n4532 VDD.n4531 304.459
R6146 VDD.n4020 VDD.t141 287.159
R6147 VDD.n1820 VDD.t138 287.159
R6148 VDD.n1984 VDD.t147 287.159
R6149 VDD.n443 VDD.t105 286.277
R6150 VDD.n977 VDD.t93 286.277
R6151 VDD.n3932 VDD.t111 286.277
R6152 VDD.n3733 VDD.t117 286.277
R6153 VDD.n546 VDD.t100 278.947
R6154 VDD.n1132 VDD.t97 278.947
R6155 VDD.n2095 VDD.t88 278.947
R6156 VDD.n2510 VDD.t130 278.947
R6157 VDD.n4553 VDD.t121 278.947
R6158 VDD.n4429 VDD.t103 278.947
R6159 VDD.n4251 VDD.t145 278.947
R6160 VDD.n1182 VDD 242.106
R6161 VDD VDD.n1534 242.106
R6162 VDD VDD.n181 242.106
R6163 VDD VDD.n2532 242.106
R6164 VDD.n4475 VDD 242.106
R6165 VDD.n4297 VDD 242.106
R6166 VDD.n3460 VDD 219.232
R6167 VDD.n3364 VDD 219.232
R6168 VDD.n1819 VDD.t756 202.559
R6169 VDD.n1983 VDD.t753 202.559
R6170 VDD.n976 VDD.t773 202.559
R6171 VDD.n442 VDD.t768 202.559
R6172 VDD.n3732 VDD.t763 202.559
R6173 VDD.n3931 VDD.t765 202.559
R6174 VDD.n4019 VDD.t757 202.559
R6175 VDD.n2 VDD.t532 201.19
R6176 VDD.n2911 VDD.t416 201.19
R6177 VDD.n2843 VDD 200.556
R6178 VDD.n2888 VDD 200.556
R6179 VDD.n3128 VDD 200.556
R6180 VDD VDD.n3185 200.556
R6181 VDD.n953 VDD 197.917
R6182 VDD.n1738 VDD 197.917
R6183 VDD VDD.n1909 197.917
R6184 VDD.n3709 VDD 197.917
R6185 VDD.n3908 VDD 197.917
R6186 VDD.n3996 VDD 197.917
R6187 VDD VDD.n1207 185
R6188 VDD VDD.n1508 185
R6189 VDD.n2292 VDD 177.474
R6190 VDD.n4770 VDD 177.474
R6191 VDD.n2817 VDD.n2816 174.595
R6192 VDD.n48 VDD.n47 174.595
R6193 VDD.n42 VDD.n41 174.595
R6194 VDD.n32 VDD.n31 174.595
R6195 VDD.n84 VDD.n83 174.595
R6196 VDD.n67 VDD.n66 174.595
R6197 VDD.n125 VDD.n124 174.595
R6198 VDD.n111 VDD.n110 174.595
R6199 VDD.n102 VDD.n101 174.595
R6200 VDD.n4858 VDD.n4857 174.595
R6201 VDD.n3109 VDD.n3108 174.595
R6202 VDD.n2780 VDD.n2779 174.595
R6203 VDD.n3081 VDD.n3080 174.595
R6204 VDD.n3067 VDD.n3066 174.595
R6205 VDD.n3042 VDD.n3041 174.595
R6206 VDD.n3027 VDD.n3026 174.595
R6207 VDD.n2987 VDD.n2986 174.595
R6208 VDD.n2980 VDD.n2979 174.595
R6209 VDD.n2956 VDD.n2955 174.595
R6210 VDD.n2949 VDD.n2948 174.595
R6211 VDD.t138 VDD.n1819 173.638
R6212 VDD.t147 VDD.n1983 173.638
R6213 VDD.t93 VDD.n976 173.638
R6214 VDD.t105 VDD.n442 173.638
R6215 VDD.t117 VDD.n3732 173.638
R6216 VDD.t111 VDD.n3931 173.638
R6217 VDD.t141 VDD.n4019 173.638
R6218 VDD.n521 VDD.t666 168.422
R6219 VDD.n1157 VDD.t203 168.422
R6220 VDD.n2120 VDD.t19 168.422
R6221 VDD.n2366 VDD.t302 168.422
R6222 VDD.n2536 VDD.t751 168.422
R6223 VDD.n4454 VDD.t388 168.422
R6224 VDD.n4276 VDD.t456 168.422
R6225 VDD.n1941 VDD.n1940 166.542
R6226 VDD.n1023 VDD.n1022 166.542
R6227 VDD.n595 VDD.n594 166.542
R6228 VDD.n4066 VDD.n4065 166.542
R6229 VDD.n3531 VDD.n3530 166.542
R6230 VDD.n3849 VDD.n3848 166.542
R6231 VDD.n3661 VDD.n3660 166.542
R6232 VDD.n551 VDD.n550 166.542
R6233 VDD.n4246 VDD.n4245 166.542
R6234 VDD.n4423 VDD.n4422 166.542
R6235 VDD.n4576 VDD.n4575 166.542
R6236 VDD.n2507 VDD.n2506 166.542
R6237 VDD.n2090 VDD.n2089 166.542
R6238 VDD.n1127 VDD.n1126 166.542
R6239 VDD.n2879 VDD.n2878 166.381
R6240 VDD.n3191 VDD.n3190 166.381
R6241 VDD.n3180 VDD.n3176 166.006
R6242 VDD.n4001 VDD.n4000 165.578
R6243 VDD.n3913 VDD.n3912 165.578
R6244 VDD.n3714 VDD.n3713 165.578
R6245 VDD.n424 VDD.n423 165.578
R6246 VDD.n958 VDD.n957 165.578
R6247 VDD.n1743 VDD.n1742 165.578
R6248 VDD.n1901 VDD.n1900 165.578
R6249 VDD.n4184 VDD.n4183 165.578
R6250 VDD.n4302 VDD.n4301 165.578
R6251 VDD.n4480 VDD.n4479 165.578
R6252 VDD.n4626 VDD.n4625 165.578
R6253 VDD.n2014 VDD.n2013 165.578
R6254 VDD.n1574 VDD.n1573 165.578
R6255 VDD.n1062 VDD.n1061 165.578
R6256 VDD.n2931 VDD.n2930 164.797
R6257 VDD.n2860 VDD.n2856 164.453
R6258 VDD.n3143 VDD.n3139 164.453
R6259 VDD.n2835 VDD.t653 159.46
R6260 VDD.n3120 VDD.t686 159.46
R6261 VDD.n2846 VDD.t153 148.195
R6262 VDD.n2775 VDD.t486 148.195
R6263 VDD.n1147 VDD.t96 146.554
R6264 VDD.n2560 VDD.t120 146.553
R6265 VDD.n4266 VDD.t144 146.553
R6266 VDD.n4444 VDD.t102 146.553
R6267 VDD.n2498 VDD.t129 146.553
R6268 VDD.n2110 VDD.t87 146.553
R6269 VDD.n433 VDD.t315 145.139
R6270 VDD.n967 VDD.t461 145.139
R6271 VDD.n1754 VDD.t469 145.139
R6272 VDD.n1806 VDD.t233 145.139
R6273 VDD.n3723 VDD.t184 145.139
R6274 VDD.n3922 VDD.t353 145.139
R6275 VDD.n4010 VDD.t277 145.139
R6276 VDD.t675 VDD.n1206 143.544
R6277 VDD.t207 VDD.n1507 143.544
R6278 VDD.n540 VDD.t99 142.458
R6279 VDD.n531 VDD.t759 137.93
R6280 VDD.n1138 VDD.t767 137.93
R6281 VDD.n2101 VDD.t772 137.93
R6282 VDD.n2489 VDD.t754 137.93
R6283 VDD.n2551 VDD.t760 137.93
R6284 VDD.n4435 VDD.t762 137.93
R6285 VDD.n4257 VDD.t761 137.93
R6286 VDD.n261 VDD.n260 137.606
R6287 VDD.n3215 VDD.n3214 137.606
R6288 VDD.n3361 VDD.n3360 137.606
R6289 VDD.n3444 VDD.n3443 137.606
R6290 VDD.n3456 VDD.n3454 137.606
R6291 VDD.n2736 VDD.n2735 137.606
R6292 VDD.n314 VDD.n313 137.606
R6293 VDD.n281 VDD.n279 137.606
R6294 VDD.n1500 VDD.n1498 137.606
R6295 VDD.n1444 VDD.n1440 137.606
R6296 VDD.n2288 VDD.n221 137.606
R6297 VDD.n2318 VDD.n209 137.606
R6298 VDD.n4766 VDD.n4764 137.606
R6299 VDD.n173 VDD.n172 137.606
R6300 VDD.n539 VDD.t766 134.047
R6301 VDD.n1146 VDD.t769 134.047
R6302 VDD.n2109 VDD.t770 134.047
R6303 VDD.n2497 VDD.t755 134.047
R6304 VDD.n2559 VDD.t758 134.047
R6305 VDD.n4443 VDD.t764 134.047
R6306 VDD.n4265 VDD.t771 134.047
R6307 VDD VDD.t567 126.668
R6308 VDD VDD.t616 126.668
R6309 VDD VDD.t449 126.668
R6310 VDD VDD.t291 126.668
R6311 VDD VDD.t738 126.668
R6312 VDD VDD.t160 126.668
R6313 VDD VDD.t736 126.668
R6314 VDD.t335 VDD.n4778 125.275
R6315 VDD.n260 VDD.t163 123.496
R6316 VDD.n3214 VDD.t743 123.496
R6317 VDD.n3360 VDD.t646 123.496
R6318 VDD.n3443 VDD.t703 123.496
R6319 VDD.n3454 VDD.t741 123.496
R6320 VDD.n2735 VDD.t374 123.496
R6321 VDD.n313 VDD.t602 123.496
R6322 VDD.n279 VDD.t711 123.496
R6323 VDD.n1498 VDD.t636 123.496
R6324 VDD.n1440 VDD.t406 123.496
R6325 VDD.n221 VDD.t444 123.496
R6326 VDD.n209 VDD.t399 123.496
R6327 VDD.n4764 VDD.t576 123.496
R6328 VDD.n172 VDD.t298 123.496
R6329 VDD.n1781 VDD.t468 121.953
R6330 VDD.n996 VDD.t460 121.953
R6331 VDD.n4039 VDD.t276 121.953
R6332 VDD.n3951 VDD.t352 121.953
R6333 VDD.n3798 VDD.t189 121.953
R6334 VDD.n2467 VDD.t238 121.953
R6335 VDD.n462 VDD.t314 121.953
R6336 VDD.n680 VDD.t45 121.953
R6337 VDD.n2638 VDD.t307 121.953
R6338 VDD.n4339 VDD.t212 121.953
R6339 VDD.n4531 VDD.t61 121.953
R6340 VDD.n4668 VDD.t634 121.953
R6341 VDD.n2005 VDD.t480 121.953
R6342 VDD.n1100 VDD.t717 121.953
R6343 VDD.n324 VDD 120.055
R6344 VDD.n454 VDD.t647 118.751
R6345 VDD.n988 VDD.t328 118.751
R6346 VDD.n1971 VDD.t23 118.751
R6347 VDD.n1827 VDD.t16 118.751
R6348 VDD.n3778 VDD.t651 118.751
R6349 VDD.n3943 VDD.t299 118.751
R6350 VDD.n4031 VDD.t705 118.751
R6351 VDD.n692 VDD.t648 118.421
R6352 VDD.n1091 VDD.t310 118.421
R6353 VDD.n2060 VDD.t325 118.421
R6354 VDD.n4660 VDD.t689 118.421
R6355 VDD.n4518 VDD.t377 118.421
R6356 VDD.n4398 VDD.t734 118.421
R6357 VDD.n4121 VDD.t198 118.421
R6358 VDD.n1239 VDD 117.445
R6359 VDD.n425 VDD.t14 116.112
R6360 VDD.n657 VDD.t628 116.112
R6361 VDD.n291 VDD.t58 116.112
R6362 VDD.n945 VDD.t567 116.112
R6363 VDD.n959 VDD.t712 116.112
R6364 VDD.n1715 VDD.t582 116.112
R6365 VDD.n1719 VDD.t66 116.112
R6366 VDD.n1730 VDD.t616 116.112
R6367 VDD.n1744 VDD.t643 116.112
R6368 VDD.n1919 VDD.t266 116.112
R6369 VDD.n1791 VDD.t74 116.112
R6370 VDD.t449 VDD.n1799 116.112
R6371 VDD.n1902 VDD.t8 116.112
R6372 VDD.n3688 VDD.t707 116.112
R6373 VDD.n3692 VDD.t337 116.112
R6374 VDD.t291 VDD.n3707 116.112
R6375 VDD.n3715 VDD.t259 116.112
R6376 VDD.n3886 VDD.t332 116.112
R6377 VDD.n3890 VDD.t569 116.112
R6378 VDD.n3900 VDD.t738 116.112
R6379 VDD.n3914 VDD.t36 116.112
R6380 VDD.n3619 VDD.t180 116.112
R6381 VDD.n2673 VDD.t671 116.112
R6382 VDD.n3988 VDD.t160 116.112
R6383 VDD.n4002 VDD.t445 116.112
R6384 VDD.n2657 VDD.t549 116.112
R6385 VDD.n3241 VDD.t70 116.112
R6386 VDD.t736 VDD.n3251 116.112
R6387 VDD.n68 VDD.t517 116.112
R6388 VDD.n2820 VDD.t652 116.112
R6389 VDD.n2880 VDD.t261 116.112
R6390 VDD.n2927 VDD.t38 116.112
R6391 VDD.n2927 VDD.t326 116.112
R6392 VDD.n3022 VDD.t411 116.112
R6393 VDD.n3114 VDD.t685 116.112
R6394 VDD.n3192 VDD.t341 116.112
R6395 VDD.n3177 VDD.t12 116.112
R6396 VDD.n3177 VDD.t573 116.112
R6397 VDD.n499 VDD.t641 115.79
R6398 VDD.n508 VDD.t164 115.79
R6399 VDD.n513 VDD.t241 115.79
R6400 VDD.n1063 VDD.t498 115.79
R6401 VDD.n1070 VDD.t365 115.79
R6402 VDD.n1169 VDD.t215 115.79
R6403 VDD.n1165 VDD.t251 115.79
R6404 VDD.n1575 VDD.t150 115.79
R6405 VDD.n1593 VDD.t190 115.79
R6406 VDD.n1606 VDD.t76 115.79
R6407 VDD.n2000 VDD.t293 115.79
R6408 VDD.n2015 VDD.t333 115.79
R6409 VDD.n2342 VDD.t257 115.79
R6410 VDD.n2351 VDD.t339 115.79
R6411 VDD.n2356 VDD.t594 115.79
R6412 VDD.n4623 VDD.t649 115.79
R6413 VDD.n2533 VDD.t547 115.79
R6414 VDD.n4607 VDD.t571 115.79
R6415 VDD.n4603 VDD.t223 115.79
R6416 VDD.n4481 VDD.t52 115.79
R6417 VDD.n2589 VDD.t321 115.79
R6418 VDD.n2594 VDD.t673 115.79
R6419 VDD.n4462 VDD.t85 115.79
R6420 VDD.n4303 VDD.t359 115.79
R6421 VDD.n2624 VDD.t343 115.79
R6422 VDD.n2629 VDD.t176 115.79
R6423 VDD.n4284 VDD.t730 115.79
R6424 VDD.n4185 VDD.t357 115.79
R6425 VDD.t40 VDD.n3447 114.835
R6426 VDD.n3380 VDD.t273 114.835
R6427 VDD.t244 VDD.n3219 114.835
R6428 VDD.n338 VDD.t601 112.225
R6429 VDD.n1253 VDD.t162 109.615
R6430 VDD.n429 VDD.t311 108.195
R6431 VDD.n963 VDD.t463 108.195
R6432 VDD.n1748 VDD.t471 108.195
R6433 VDD.n1896 VDD.t235 108.195
R6434 VDD.n3719 VDD.t186 108.195
R6435 VDD.n3918 VDD.t349 108.195
R6436 VDD.n4006 VDD.t279 108.195
R6437 VDD.n703 VDD.t46 107.895
R6438 VDD.n1569 VDD.t714 107.895
R6439 VDD.n2019 VDD.t475 107.895
R6440 VDD.n4629 VDD.t629 107.895
R6441 VDD.n4485 VDD.t64 107.895
R6442 VDD.n4307 VDD.t213 107.895
R6443 VDD.n4179 VDD.t304 107.895
R6444 VDD.n945 VDD.t626 105.556
R6445 VDD.n1730 VDD.t583 105.556
R6446 VDD.n1799 VDD.t264 105.556
R6447 VDD.n3707 VDD.t708 105.556
R6448 VDD.n3900 VDD.t329 105.556
R6449 VDD.n3988 VDD.t181 105.556
R6450 VDD.n3251 VDD.t550 105.556
R6451 VDD.n68 VDD.t543 105.556
R6452 VDD.n2820 VDD.t658 105.556
R6453 VDD.n2880 VDD.t158 105.556
R6454 VDD.n3022 VDD.t427 105.556
R6455 VDD.n3114 VDD.t687 105.556
R6456 VDD.n3192 VDD.t489 105.556
R6457 VDD.n499 VDD.t239 105.263
R6458 VDD.n1070 VDD.t249 105.263
R6459 VDD.n1593 VDD.t295 105.263
R6460 VDD.n2342 VDD.t596 105.263
R6461 VDD.n2533 VDD.t221 105.263
R6462 VDD.n2589 VDD.t83 105.263
R6463 VDD.n2624 VDD.t731 105.263
R6464 VDD.n3480 VDD.t604 104.397
R6465 VDD.n3336 VDD.t605 104.397
R6466 VDD.n589 VDD.t747 102.918
R6467 VDD.n1018 VDD.t369 102.918
R6468 VDD.n1946 VDD.t361 102.918
R6469 VDD.n3656 VDD.t194 102.918
R6470 VDD.n3844 VDD.t588 102.918
R6471 VDD.n3563 VDD.t610 102.918
R6472 VDD.n4061 VDD.t614 102.918
R6473 VDD.n556 VDD.t664 102.632
R6474 VDD.n1122 VDD.t205 102.632
R6475 VDD.n2085 VDD.t21 102.632
R6476 VDD.n4691 VDD.t300 102.632
R6477 VDD.n4568 VDD.t749 102.632
R6478 VDD.n2603 VDD.t386 102.632
R6479 VDD.n4241 VDD.t454 102.632
R6480 VDD.n4374 VDD.t209 100.001
R6481 VDD.n890 VDD.t710 99.1763
R6482 VDD.n1671 VDD.t635 99.1763
R6483 VDD.n2253 VDD.t441 99.1763
R6484 VDD.n2260 VDD.t282 99.1763
R6485 VDD.n4730 VDD.t669 99.1763
R6486 VDD.n4735 VDD.t603 99.1763
R6487 VDD.n1560 VDD.t718 97.3689
R6488 VDD.n4646 VDD.t631 97.3689
R6489 VDD.n662 VDD.t637 95.0005
R6490 VDD.n1711 VDD.t80 95.0005
R6491 VDD.n1923 VDD.t481 95.0005
R6492 VDD.n3684 VDD.t226 95.0005
R6493 VDD.n3882 VDD.t356 95.0005
R6494 VDD.n3615 VDD.t192 95.0005
R6495 VDD.n2651 VDD.t724 95.0005
R6496 VDD.n119 VDD.t533 95.0005
R6497 VDD.n3011 VDD.t413 95.0005
R6498 VDD.n517 VDD.t690 94.7373
R6499 VDD.n1161 VDD.t394 94.7373
R6500 VDD.n2125 VDD.t73 94.7373
R6501 VDD.n2360 VDD.t167 94.7373
R6502 VDD.n4598 VDD.t451 94.7373
R6503 VDD.n4458 VDD.t253 94.7373
R6504 VDD.n4280 VDD.t474 94.7373
R6505 VDD.n3487 VDD.t172 93.9565
R6506 VDD.n3331 VDD.t32 93.9565
R6507 VDD.n2752 VDD.n2751 92.5005
R6508 VDD.n2751 VDD.n2750 92.5005
R6509 VDD.n2749 VDD.n2748 92.5005
R6510 VDD.n2748 VDD.n2747 92.5005
R6511 VDD.n2746 VDD.n2745 92.5005
R6512 VDD.n2745 VDD.n2744 92.5005
R6513 VDD.n2743 VDD.n2742 92.5005
R6514 VDD.n2742 VDD.n2741 92.5005
R6515 VDD.n2740 VDD.n2739 92.5005
R6516 VDD.n2739 VDD.n2738 92.5005
R6517 VDD.n3325 VDD.n3324 92.5005
R6518 VDD.n3324 VDD.n3323 92.5005
R6519 VDD.n3328 VDD.n3327 92.5005
R6520 VDD.n3327 VDD.n3326 92.5005
R6521 VDD.n3322 VDD.n3321 92.5005
R6522 VDD.n3321 VDD.n3320 92.5005
R6523 VDD.n3333 VDD.n3332 92.5005
R6524 VDD.n3332 VDD.n3331 92.5005
R6525 VDD.n3338 VDD.n3337 92.5005
R6526 VDD.n3337 VDD.n3336 92.5005
R6527 VDD.n3345 VDD.n3344 92.5005
R6528 VDD.n3344 VDD.n3343 92.5005
R6529 VDD.n3350 VDD.n3349 92.5005
R6530 VDD.n3349 VDD.n3348 92.5005
R6531 VDD.n3355 VDD.n3354 92.5005
R6532 VDD.n3354 VDD.n3353 92.5005
R6533 VDD.n3366 VDD.n3365 92.5005
R6534 VDD.n3365 VDD.n3364 92.5005
R6535 VDD.n3362 VDD.n2737 92.5005
R6536 VDD.n3363 VDD.n3362 92.5005
R6537 VDD.n3373 VDD.n3372 92.5005
R6538 VDD.n3372 VDD.n3371 92.5005
R6539 VDD.n3376 VDD.n3375 92.5005
R6540 VDD.n3375 VDD.n3374 92.5005
R6541 VDD.n2692 VDD.n2691 92.5005
R6542 VDD.n2691 VDD.n2690 92.5005
R6543 VDD.n2689 VDD.n2688 92.5005
R6544 VDD.n2688 VDD.n2687 92.5005
R6545 VDD.n2686 VDD.n2685 92.5005
R6546 VDD.n2685 VDD.n2684 92.5005
R6547 VDD.n3497 VDD.n3496 92.5005
R6548 VDD.n3496 VDD.n3495 92.5005
R6549 VDD.n3500 VDD.n3499 92.5005
R6550 VDD.n3499 VDD.n3498 92.5005
R6551 VDD.n3503 VDD.n3502 92.5005
R6552 VDD.n3502 VDD.n3501 92.5005
R6553 VDD.n3506 VDD.n3505 92.5005
R6554 VDD.n3505 VDD.n3504 92.5005
R6555 VDD.n3494 VDD.n3493 92.5005
R6556 VDD.n3493 VDD.n3492 92.5005
R6557 VDD.n3489 VDD.n3488 92.5005
R6558 VDD.n3488 VDD.n3487 92.5005
R6559 VDD.n3482 VDD.n3481 92.5005
R6560 VDD.n3481 VDD.n3480 92.5005
R6561 VDD.n3477 VDD.n3476 92.5005
R6562 VDD.n3476 VDD.n3475 92.5005
R6563 VDD.n3472 VDD.n3471 92.5005
R6564 VDD.n3471 VDD.n3470 92.5005
R6565 VDD.n3467 VDD.n3466 92.5005
R6566 VDD.n3466 VDD.n3465 92.5005
R6567 VDD.n3462 VDD.n3461 92.5005
R6568 VDD.n3461 VDD.n3460 92.5005
R6569 VDD.n3458 VDD.n3457 92.5005
R6570 VDD.n3459 VDD.n3458 92.5005
R6571 VDD.n3403 VDD.n3402 92.5005
R6572 VDD.n3402 VDD.n3401 92.5005
R6573 VDD.n3442 VDD.n3441 92.5005
R6574 VDD.n3441 VDD.n3440 92.5005
R6575 VDD.n3408 VDD.n3407 92.5005
R6576 VDD.n3407 VDD.n3406 92.5005
R6577 VDD.n809 VDD.n808 92.5005
R6578 VDD.n808 VDD.n807 92.5005
R6579 VDD.n806 VDD.n805 92.5005
R6580 VDD.n805 VDD.n804 92.5005
R6581 VDD.n803 VDD.n802 92.5005
R6582 VDD.n802 VDD.n801 92.5005
R6583 VDD.n800 VDD.n799 92.5005
R6584 VDD.n799 VDD.n798 92.5005
R6585 VDD.n797 VDD.n796 92.5005
R6586 VDD.n796 VDD.n795 92.5005
R6587 VDD.n794 VDD.n793 92.5005
R6588 VDD.n793 VDD.n792 92.5005
R6589 VDD.n1217 VDD.n1216 92.5005
R6590 VDD.n1216 VDD.n1215 92.5005
R6591 VDD.n1214 VDD.n1213 92.5005
R6592 VDD.n1213 VDD.n1212 92.5005
R6593 VDD.n1335 VDD.n1334 92.5005
R6594 VDD.n1334 VDD.n1333 92.5005
R6595 VDD.n1351 VDD.n1350 92.5005
R6596 VDD.n1350 VDD.n1349 92.5005
R6597 VDD.n1354 VDD.n1353 92.5005
R6598 VDD.n1353 VDD.n1352 92.5005
R6599 VDD.n1357 VDD.n1356 92.5005
R6600 VDD.n1356 VDD.n1355 92.5005
R6601 VDD.n1360 VDD.n1359 92.5005
R6602 VDD.n1359 VDD.n1358 92.5005
R6603 VDD.n1363 VDD.n1362 92.5005
R6604 VDD.n1362 VDD.n1361 92.5005
R6605 VDD.n1515 VDD.n1514 92.5005
R6606 VDD.n1514 VDD.n1513 92.5005
R6607 VDD.n2247 VDD.n2246 92.5005
R6608 VDD.n2246 VDD.n2245 92.5005
R6609 VDD.n2244 VDD.n2243 92.5005
R6610 VDD.n2243 VDD.n2242 92.5005
R6611 VDD.n2241 VDD.n2240 92.5005
R6612 VDD.n2240 VDD.n2239 92.5005
R6613 VDD.n2238 VDD.n2237 92.5005
R6614 VDD.n2237 VDD.n2236 92.5005
R6615 VDD.n2217 VDD.n2216 92.5005
R6616 VDD.n2216 VDD.n2215 92.5005
R6617 VDD.n2220 VDD.n2219 92.5005
R6618 VDD.n2219 VDD.n2218 92.5005
R6619 VDD.n2223 VDD.n2222 92.5005
R6620 VDD.n2222 VDD.n2221 92.5005
R6621 VDD.n2294 VDD.n2293 92.5005
R6622 VDD.n2293 VDD.n2292 92.5005
R6623 VDD.n2290 VDD.n2289 92.5005
R6624 VDD.n2291 VDD.n2290 92.5005
R6625 VDD.n2282 VDD.n2281 92.5005
R6626 VDD.n2281 VDD.n2280 92.5005
R6627 VDD.n2277 VDD.n2276 92.5005
R6628 VDD.n2276 VDD.n2275 92.5005
R6629 VDD.n2272 VDD.n2271 92.5005
R6630 VDD.n2271 VDD.n2270 92.5005
R6631 VDD.n2267 VDD.n2266 92.5005
R6632 VDD.n2266 VDD.n2265 92.5005
R6633 VDD.n2262 VDD.n2261 92.5005
R6634 VDD.n2261 VDD.n2260 92.5005
R6635 VDD.n2255 VDD.n2254 92.5005
R6636 VDD.n2254 VDD.n2253 92.5005
R6637 VDD.n2250 VDD.n2249 92.5005
R6638 VDD.n2249 VDD.n2248 92.5005
R6639 VDD.n220 VDD.n219 92.5005
R6640 VDD.n219 VDD.n218 92.5005
R6641 VDD.n2408 VDD.n2407 92.5005
R6642 VDD.n2407 VDD.n2406 92.5005
R6643 VDD.n2405 VDD.n2404 92.5005
R6644 VDD.n2404 VDD.n2403 92.5005
R6645 VDD.n2402 VDD.n2401 92.5005
R6646 VDD.n2401 VDD.n2400 92.5005
R6647 VDD.n4713 VDD.n4712 92.5005
R6648 VDD.n4712 VDD.n4711 92.5005
R6649 VDD.n4716 VDD.n4715 92.5005
R6650 VDD.n4715 VDD.n4714 92.5005
R6651 VDD.n4719 VDD.n4718 92.5005
R6652 VDD.n4718 VDD.n4717 92.5005
R6653 VDD.n4722 VDD.n4721 92.5005
R6654 VDD.n4721 VDD.n4720 92.5005
R6655 VDD.n4772 VDD.n4771 92.5005
R6656 VDD.n4771 VDD.n4770 92.5005
R6657 VDD.n4768 VDD.n4767 92.5005
R6658 VDD.n4769 VDD.n4768 92.5005
R6659 VDD.n4757 VDD.n4756 92.5005
R6660 VDD.n4756 VDD.n4755 92.5005
R6661 VDD.n4752 VDD.n4751 92.5005
R6662 VDD.n4751 VDD.n4750 92.5005
R6663 VDD.n4747 VDD.n4746 92.5005
R6664 VDD.n4746 VDD.n4745 92.5005
R6665 VDD.n4737 VDD.n4736 92.5005
R6666 VDD.n4736 VDD.n4735 92.5005
R6667 VDD.n4742 VDD.n4741 92.5005
R6668 VDD.n4741 VDD.n4740 92.5005
R6669 VDD.n4732 VDD.n4731 92.5005
R6670 VDD.n4731 VDD.n4730 92.5005
R6671 VDD.n4725 VDD.n4724 92.5005
R6672 VDD.n4724 VDD.n4723 92.5005
R6673 VDD.n4763 VDD.n4762 92.5005
R6674 VDD.n4762 VDD.n4761 92.5005
R6675 VDD.n4167 VDD.t2 92.1058
R6676 VDD.n1786 VDD.t578 91.4648
R6677 VDD.n1781 VDD.t381 91.4648
R6678 VDD.n1042 VDD.t272 91.4648
R6679 VDD.n996 VDD.t723 91.4648
R6680 VDD.n629 VDD.t1 91.4648
R6681 VDD.n4093 VDD.t29 91.4648
R6682 VDD.n4039 VDD.t505 91.4648
R6683 VDD.n3599 VDD.t496 91.4648
R6684 VDD.n3951 VDD.t169 91.4648
R6685 VDD.n3872 VDD.t509 91.4648
R6686 VDD.n3798 VDD.t27 91.4648
R6687 VDD.n3674 VDD.t379 91.4648
R6688 VDD.n2467 VDD.t25 91.4648
R6689 VDD.n462 VDD.t580 91.4648
R6690 VDD.n680 VDD.t137 91.4648
R6691 VDD.n2638 VDD.t128 91.4648
R6692 VDD.n4273 VDD.t146 91.4648
R6693 VDD.n4339 VDD.t125 91.4648
R6694 VDD.n4451 VDD.t104 91.4648
R6695 VDD.n4531 VDD.t134 91.4648
R6696 VDD.n2545 VDD.t122 91.4648
R6697 VDD.n4668 VDD.t92 91.4648
R6698 VDD.n2484 VDD.t131 91.4648
R6699 VDD.n2005 VDD.t110 91.4648
R6700 VDD.n2117 VDD.t89 91.4648
R6701 VDD.n1100 VDD.t116 91.4648
R6702 VDD.n1154 VDD.t98 91.4648
R6703 VDD.n526 VDD.t101 91.4648
R6704 VDD.n2260 VDD.t68 88.7368
R6705 VDD.n4735 VDD.t246 88.7368
R6706 VDD.n463 VDD.t579 87.0838
R6707 VDD.n997 VDD.t722 87.0838
R6708 VDD.n1782 VDD.t380 87.0838
R6709 VDD.n2468 VDD.t24 87.0838
R6710 VDD.n3799 VDD.t26 87.0838
R6711 VDD.n3952 VDD.t168 87.0838
R6712 VDD.n4040 VDD.t504 87.0838
R6713 VDD.n681 VDD.t136 86.8426
R6714 VDD.n1101 VDD.t115 86.8426
R6715 VDD.n2006 VDD.t109 86.8426
R6716 VDD.n4669 VDD.t91 86.8426
R6717 VDD.n4528 VDD.t133 86.8426
R6718 VDD.n4336 VDD.t124 86.8426
R6719 VDD.n2639 VDD.t127 86.8426
R6720 VDD.n3283 VDD.t448 86.7743
R6721 VDD.n3339 VDD.t11 86.7743
R6722 VDD.n3413 VDD.t466 86.7743
R6723 VDD.n3485 VDD.t220 86.7743
R6724 VDD.n2703 VDD.t591 86.7743
R6725 VDD.n401 VDD.t324 86.7743
R6726 VDD.n839 VDD.t393 86.7743
R6727 VDD.n1303 VDD.t514 86.7743
R6728 VDD.n1393 VDD.t511 86.7743
R6729 VDD.n2185 VDD.t599 86.7743
R6730 VDD.n2258 VDD.t69 86.7743
R6731 VDD.n2438 VDD.t368 86.7743
R6732 VDD.n4728 VDD.t247 86.7743
R6733 VDD.n4815 VDD.t385 86.7743
R6734 VDD.n1786 VDD.t364 86.7743
R6735 VDD.n1940 VDD.t362 86.7743
R6736 VDD.n1042 VDD.t372 86.7743
R6737 VDD.n1022 VDD.t370 86.7743
R6738 VDD.n629 VDD.t746 86.7743
R6739 VDD.n594 VDD.t748 86.7743
R6740 VDD.n4093 VDD.t613 86.7743
R6741 VDD.n4065 VDD.t615 86.7743
R6742 VDD.n3599 VDD.t609 86.7743
R6743 VDD.n3530 VDD.t611 86.7743
R6744 VDD.n3872 VDD.t587 86.7743
R6745 VDD.n3848 VDD.t589 86.7743
R6746 VDD.n3674 VDD.t197 86.7743
R6747 VDD.n3660 VDD.t195 86.7743
R6748 VDD.n550 VDD.t665 86.7743
R6749 VDD.n4245 VDD.t455 86.7743
R6750 VDD.n4273 VDD.t457 86.7743
R6751 VDD.n4422 VDD.t387 86.7743
R6752 VDD.n4451 VDD.t389 86.7743
R6753 VDD.n4575 VDD.t750 86.7743
R6754 VDD.n2545 VDD.t752 86.7743
R6755 VDD.n2506 VDD.t301 86.7743
R6756 VDD.n2484 VDD.t303 86.7743
R6757 VDD.n2089 VDD.t22 86.7743
R6758 VDD.n2117 VDD.t20 86.7743
R6759 VDD.n1126 VDD.t206 86.7743
R6760 VDD.n1154 VDD.t204 86.7743
R6761 VDD.n526 VDD.t667 86.7743
R6762 VDD.n72 VDD.t515 84.4449
R6763 VDD.n2814 VDD.t654 84.4449
R6764 VDD.n2801 VDD.t154 84.4449
R6765 VDD.n3016 VDD.t409 84.4449
R6766 VDD.n3106 VDD.t681 84.4449
R6767 VDD.n3154 VDD.t487 84.4449
R6768 VDD.n739 VDD.t269 84.211
R6769 VDD.n2051 VDD.t606 84.211
R6770 VDD.n4651 VDD.t506 84.211
R6771 VDD.n4509 VDD.t30 84.211
R6772 VDD.n4357 VDD.t592 84.211
R6773 VDD.n352 VDD.t564 83.517
R6774 VDD.n3480 VDD.t219 83.517
R6775 VDD.n3336 VDD.t10 83.517
R6776 VDD.t641 VDD 81.5794
R6777 VDD.t365 VDD 81.5794
R6778 VDD.t190 VDD 81.5794
R6779 VDD.t257 VDD 81.5794
R6780 VDD.t547 VDD 81.5794
R6781 VDD.t321 VDD 81.5794
R6782 VDD.t343 VDD 81.5794
R6783 VDD.n3220 VDD 81.5278
R6784 VDD.n1267 VDD.t561 80.9071
R6785 VDD VDD.n1477 80.9071
R6786 VDD.n2314 VDD 80.9071
R6787 VDD.n1478 VDD.t319 78.2972
R6788 VDD.t17 VDD.n2311 78.2972
R6789 VDD.n4779 VDD 78.2972
R6790 VDD.n1819 VDD 78.1104
R6791 VDD.n1983 VDD 78.1104
R6792 VDD.n976 VDD 78.1104
R6793 VDD.n442 VDD 78.1104
R6794 VDD.n3732 VDD 78.1104
R6795 VDD.n3931 VDD 78.1104
R6796 VDD.n4019 VDD 78.1104
R6797 VDD.n3 VDD.t531 77.5227
R6798 VDD.n2913 VDD.t415 77.5227
R6799 VDD.n626 VDD.t745 73.8894
R6800 VDD.n1039 VDD.t371 73.8894
R6801 VDD.n1787 VDD.t363 73.8894
R6802 VDD.n3675 VDD.t196 73.8894
R6803 VDD.n3873 VDD.t586 73.8894
R6804 VDD.n3605 VDD.t608 73.8894
R6805 VDD.n4094 VDD.t612 73.8894
R6806 VDD.n127 VDD.t521 73.8894
R6807 VDD.n2988 VDD.t429 73.8894
R6808 VDD.n1459 VDD.t405 73.0774
R6809 VDD.n199 VDD.t398 73.0774
R6810 VDD.n3448 VDD 73.0774
R6811 VDD VDD.n3379 73.0774
R6812 VDD.n454 VDD.t502 71.2505
R6813 VDD.n988 VDD.t201 71.2505
R6814 VDD.n1971 VDD.t285 71.2505
R6815 VDD.n1827 VDD.t696 71.2505
R6816 VDD.n3778 VDD.t287 71.2505
R6817 VDD.n3943 VDD.t229 71.2505
R6818 VDD.n4031 VDD.t698 71.2505
R6819 VDD.n692 VDD.t4 71.0531
R6820 VDD.n1091 VDD.t345 71.0531
R6821 VDD.n2060 VDD.t48 71.0531
R6822 VDD.n4660 VDD.t401 71.0531
R6823 VDD.n4518 VDD.t493 71.0531
R6824 VDD.n4398 VDD.t621 71.0531
R6825 VDD.n4121 VDD.t728 71.0531
R6826 VDD.n910 VDD.t557 70.4675
R6827 VDD.n1687 VDD.t562 70.4675
R6828 VDD.n4783 VDD.t297 70.4675
R6829 VDD.n3435 VDD.t702 70.4675
R6830 VDD.n3384 VDD.t373 70.4675
R6831 VDD.n3305 VDD.t742 70.4675
R6832 VDD.n3283 VDD.t376 68.0124
R6833 VDD.n3339 VDD.t33 68.0124
R6834 VDD.n3413 VDD.t391 68.0124
R6835 VDD.n3485 VDD.t173 68.0124
R6836 VDD.n2703 VDD.t397 68.0124
R6837 VDD.n401 VDD.t175 68.0124
R6838 VDD.n839 VDD.t640 68.0124
R6839 VDD.n1303 VDD.t218 68.0124
R6840 VDD.n1393 VDD.t383 68.0124
R6841 VDD.n2185 VDD.t171 68.0124
R6842 VDD.n2258 VDD.t442 68.0124
R6843 VDD.n2438 VDD.t79 68.0124
R6844 VDD.n4728 VDD.t670 68.0124
R6845 VDD.n4815 VDD.t57 68.0124
R6846 VDD.n79 VDD.t537 63.3338
R6847 VDD.n141 VDD.t660 63.3338
R6848 VDD.n2857 VDD.t156 63.3338
R6849 VDD.n3044 VDD.t423 63.3338
R6850 VDD.n2783 VDD.t677 63.3338
R6851 VDD.n3140 VDD.t483 63.3338
R6852 VDD.n1800 VDD.t140 63.1021
R6853 VDD.n1775 VDD.t149 63.1021
R6854 VDD.n971 VDD.t95 63.1021
R6855 VDD.n437 VDD.t107 63.1021
R6856 VDD.n3727 VDD.t119 63.1021
R6857 VDD.n3926 VDD.t113 63.1021
R6858 VDD.n4014 VDD.t143 63.1021
R6859 VDD.n719 VDD.t270 63.1021
R6860 VDD.n1558 VDD.t721 63.1021
R6861 VDD.n2029 VDD.t607 63.1021
R6862 VDD.n4639 VDD.t507 63.1021
R6863 VDD.n4495 VDD.t31 63.1021
R6864 VDD.n4367 VDD.t593 63.1021
R6865 VDD.n4143 VDD.t3 63.1021
R6866 VDD.n2275 VDD.t563 62.6379
R6867 VDD.n4750 VDD.t560 62.6379
R6868 VDD.n1547 VDD.n1544 60.0005
R6869 VDD.n725 VDD.n722 60.0005
R6870 VDD.n4000 VDD.t280 58.4849
R6871 VDD.n3912 VDD.t350 58.4849
R6872 VDD.n3713 VDD.t187 58.4849
R6873 VDD.n423 VDD.t312 58.4849
R6874 VDD.n957 VDD.t464 58.4849
R6875 VDD.n1742 VDD.t472 58.4849
R6876 VDD.n1900 VDD.t236 58.4849
R6877 VDD.n4183 VDD.t305 58.4849
R6878 VDD.n4301 VDD.t214 58.4849
R6879 VDD.n4479 VDD.t65 58.4849
R6880 VDD.n4625 VDD.t630 58.4849
R6881 VDD.n2013 VDD.t476 58.4849
R6882 VDD.n1573 VDD.t715 58.4849
R6883 VDD.n1061 VDD.t47 58.4849
R6884 VDD.n394 VDD.t323 57.4181
R6885 VDD.n3465 VDD.t554 57.4181
R6886 VDD.n3353 VDD.t553 57.4181
R6887 VDD.n1435 VDD.n1434 56.4711
R6888 VDD.n1439 VDD.n1438 56.4711
R6889 VDD.n1456 VDD.n1455 56.4711
R6890 VDD.n230 VDD.n229 56.4711
R6891 VDD.n2160 VDD.n2159 56.4711
R6892 VDD.n2174 VDD.n2173 56.4711
R6893 VDD.n2190 VDD.n2189 56.4711
R6894 VDD.n2204 VDD.n2203 56.4711
R6895 VDD.n2227 VDD.n2226 56.4711
R6896 VDD.n215 VDD.n214 56.4711
R6897 VDD.n213 VDD.n212 56.4711
R6898 VDD.n196 VDD.n195 56.4711
R6899 VDD.n1853 VDD.n1852 56.4711
R6900 VDD.n1871 VDD.n1870 56.4711
R6901 VDD.n2387 VDD.n2386 56.4711
R6902 VDD.n2444 VDD.n2443 56.4711
R6903 VDD.n2426 VDD.n2425 56.4711
R6904 VDD.n2412 VDD.n2411 56.4711
R6905 VDD.n325 VDD.n312 56.4711
R6906 VDD.n339 VDD.n335 56.4711
R6907 VDD.n353 VDD.n349 56.4711
R6908 VDD.n367 VDD.n363 56.4711
R6909 VDD.n381 VDD.n377 56.4711
R6910 VDD.n395 VDD.n391 56.4711
R6911 VDD.n409 VDD.n405 56.4711
R6912 VDD.n788 VDD.n784 56.4711
R6913 VDD.n2048 VDD.n2047 56.4711
R6914 VDD.n2034 VDD.n2033 56.4711
R6915 VDD.n4643 VDD.n4642 56.4711
R6916 VDD.n4500 VDD.n4499 56.4711
R6917 VDD.n4354 VDD.n4353 56.4711
R6918 VDD.n4371 VDD.n4370 56.4711
R6919 VDD.n736 VDD.n735 56.4711
R6920 VDD.n4148 VDD.n4147 54.8576
R6921 VDD.n1311 VDD.t513 54.8082
R6922 VDD.n1233 VDD.n267 52.9417
R6923 VDD.n1240 VDD.n265 52.9417
R6924 VDD.n1254 VDD.n1250 52.9417
R6925 VDD.n1268 VDD.n1264 52.9417
R6926 VDD.n1282 VDD.n1278 52.9417
R6927 VDD.n1296 VDD.n1292 52.9417
R6928 VDD.n1312 VDD.n1308 52.9417
R6929 VDD.n1326 VDD.n1322 52.9417
R6930 VDD.n1343 VDD.n1339 52.9417
R6931 VDD.n4851 VDD.t519 52.7783
R6932 VDD.n114 VDD.t535 52.7783
R6933 VDD.n2944 VDD.t437 52.7783
R6934 VDD.n2994 VDD.t417 52.7783
R6935 VDD VDD.t675 52.1983
R6936 VDD VDD.t207 52.1983
R6937 VDD VDD.t623 52.1983
R6938 VDD VDD.t54 52.1983
R6939 VDD VDD.t40 52.1983
R6940 VDD.t273 VDD 52.1983
R6941 VDD VDD.t244 52.1983
R6942 VDD.n723 VDD.t42 50.0005
R6943 VDD.n2035 VDD.t477 50.0005
R6944 VDD.n4501 VDD.t62 50.0005
R6945 VDD.n4149 VDD.t308 47.3689
R6946 VDD.n408 VDD.t174 46.9785
R6947 VDD.n2921 VDD 44.8616
R6948 VDD.n3162 VDD 44.8616
R6949 VDD.n724 VDD.n723 44.7373
R6950 VDD.n1546 VDD.n1545 44.7373
R6951 VDD.n4164 VDD.n4163 44.5719
R6952 VDD.n847 VDD.t392 44.3686
R6953 VDD.n1325 VDD.t217 44.3686
R6954 VDD.n1405 VDD.t510 44.3686
R6955 VDD.n233 VDD.t566 44.3686
R6956 VDD.n1856 VDD.t559 44.3686
R6957 VDD.n20 VDD.t527 42.2227
R6958 VDD.n49 VDD.t656 42.2227
R6959 VDD VDD.n2842 42.2227
R6960 VDD.n2850 VDD.t152 42.2227
R6961 VDD VDD.n2887 42.2227
R6962 VDD.n3050 VDD.t433 42.2227
R6963 VDD.n2777 VDD.t683 42.2227
R6964 VDD VDD.n3127 42.2227
R6965 VDD.n3133 VDD.t485 42.2227
R6966 VDD.n3186 VDD 42.2227
R6967 VDD.n738 VDD.n737 42.1058
R6968 VDD.n2050 VDD.n2049 42.1058
R6969 VDD.n2036 VDD.n2035 42.1058
R6970 VDD.n4645 VDD.n4644 42.1058
R6971 VDD.n4502 VDD.n4501 42.1058
R6972 VDD.n4356 VDD.n4355 42.1058
R6973 VDD.n4373 VDD.n4372 42.1058
R6974 VDD.n4150 VDD.n4149 42.1058
R6975 VDD.n324 VDD.n323 41.7587
R6976 VDD.n338 VDD.n337 41.7587
R6977 VDD.n352 VDD.n351 41.7587
R6978 VDD.n366 VDD.n365 41.7587
R6979 VDD.n380 VDD.n379 41.7587
R6980 VDD.n394 VDD.n393 41.7587
R6981 VDD.n408 VDD.n407 41.7587
R6982 VDD.n787 VDD.n786 41.7587
R6983 VDD.t267 VDD.n1236 41.7587
R6984 VDD.n1479 VDD.n1478 41.7587
R6985 VDD.n1437 VDD.n1436 41.7587
R6986 VDD.n1458 VDD.n1457 41.7587
R6987 VDD.n232 VDD.n231 41.7587
R6988 VDD.n2162 VDD.n2161 41.7587
R6989 VDD.n2192 VDD.n2191 41.7587
R6990 VDD.n2206 VDD.n2205 41.7587
R6991 VDD.n2229 VDD.n2228 41.7587
R6992 VDD.n2311 VDD.n2310 41.7587
R6993 VDD.n2313 VDD.n2312 41.7587
R6994 VDD.n198 VDD.n197 41.7587
R6995 VDD.n1855 VDD.n1854 41.7587
R6996 VDD.n1873 VDD.n1872 41.7587
R6997 VDD.n2446 VDD.n2445 41.7587
R6998 VDD.n2428 VDD.n2427 41.7587
R6999 VDD.n2414 VDD.n2413 41.7587
R7000 VDD.n4787 VDD.t565 41.7587
R7001 VDD.n3431 VDD.t556 41.7587
R7002 VDD.n3389 VDD.t555 41.7587
R7003 VDD.n3299 VDD.t558 41.7587
R7004 VDD.n1795 VDD.t265 41.5552
R7005 VDD.n1795 VDD.t450 41.5552
R7006 VDD.n944 VDD.t627 41.5552
R7007 VDD.n944 VDD.t568 41.5552
R7008 VDD.n3247 VDD.t551 41.5552
R7009 VDD.n3247 VDD.t737 41.5552
R7010 VDD.n3987 VDD.t182 41.5552
R7011 VDD.n3987 VDD.t161 41.5552
R7012 VDD.n3899 VDD.t330 41.5552
R7013 VDD.n3899 VDD.t739 41.5552
R7014 VDD.n3703 VDD.t709 41.5552
R7015 VDD.n3703 VDD.t292 41.5552
R7016 VDD.n1729 VDD.t584 41.5552
R7017 VDD.n1729 VDD.t617 41.5552
R7018 VDD.n2627 VDD.t344 41.5552
R7019 VDD.n2627 VDD.t732 41.5552
R7020 VDD.n2592 VDD.t322 41.5552
R7021 VDD.n2592 VDD.t84 41.5552
R7022 VDD.n4616 VDD.t548 41.5552
R7023 VDD.n4616 VDD.t222 41.5552
R7024 VDD.n180 VDD.t258 41.5552
R7025 VDD.n180 VDD.t597 41.5552
R7026 VDD.n1533 VDD.t191 41.5552
R7027 VDD.n1533 VDD.t296 41.5552
R7028 VDD.n1073 VDD.t366 41.5552
R7029 VDD.n1073 VDD.t250 41.5552
R7030 VDD.n496 VDD.t642 41.5552
R7031 VDD.n496 VDD.t240 41.5552
R7032 VDD.t231 VDD.n321 39.1488
R7033 VDD.n1235 VDD.n1234 39.1488
R7034 VDD.n1239 VDD.n1238 39.1488
R7035 VDD.n1253 VDD.n1252 39.1488
R7036 VDD.n1267 VDD.n1266 39.1488
R7037 VDD.n1281 VDD.n1280 39.1488
R7038 VDD.n1295 VDD.n1294 39.1488
R7039 VDD.n1311 VDD.n1310 39.1488
R7040 VDD.n1325 VDD.n1324 39.1488
R7041 VDD.n1342 VDD.n1341 39.1488
R7042 VDD.n817 VDD.n813 38.824
R7043 VDD.n831 VDD.n827 38.824
R7044 VDD.n848 VDD.n844 38.824
R7045 VDD.n862 VDD.n858 38.824
R7046 VDD.n876 VDD.n872 38.824
R7047 VDD.n911 VDD.n907 38.824
R7048 VDD.n891 VDD.n887 38.824
R7049 VDD.n1205 VDD.n276 38.824
R7050 VDD.n1210 VDD.n272 38.824
R7051 VDD.n1371 VDD.n1367 38.824
R7052 VDD.n1388 VDD.n1384 38.824
R7053 VDD.n1406 VDD.n1402 38.824
R7054 VDD.n1643 VDD.n1639 38.824
R7055 VDD.n1657 VDD.n1653 38.824
R7056 VDD.n1688 VDD.n1684 38.824
R7057 VDD.n1672 VDD.n1668 38.824
R7058 VDD.n1506 VDD.n1495 38.824
R7059 VDD.n1511 VDD.n1491 38.824
R7060 VDD.n1940 VDD.t284 38.6969
R7061 VDD.n1022 VDD.t200 38.6969
R7062 VDD.n594 VDD.t501 38.6969
R7063 VDD.n4065 VDD.t701 38.6969
R7064 VDD.n3530 VDD.t228 38.6969
R7065 VDD.n3848 VDD.t290 38.6969
R7066 VDD.n3660 VDD.t695 38.6969
R7067 VDD.n550 VDD.t7 38.6969
R7068 VDD.n4245 VDD.t727 38.6969
R7069 VDD.n4422 VDD.t620 38.6969
R7070 VDD.n4575 VDD.t492 38.6969
R7071 VDD.n2506 VDD.t404 38.6969
R7072 VDD.n2089 VDD.t51 38.6969
R7073 VDD.n1126 VDD.t348 38.6969
R7074 VDD.n619 VDD.t0 36.9449
R7075 VDD.n1032 VDD.t271 36.9449
R7076 VDD.n1932 VDD.t577 36.9449
R7077 VDD.n3670 VDD.t378 36.9449
R7078 VDD.n3866 VDD.t508 36.9449
R7079 VDD.n3539 VDD.t495 36.9449
R7080 VDD.n4088 VDD.t28 36.9449
R7081 VDD.n1545 VDD.t720 36.8426
R7082 VDD VDD.t231 36.539
R7083 VDD VDD.t267 36.539
R7084 VDD.t319 VDD 36.539
R7085 VDD VDD.t17 36.539
R7086 VDD VDD.t335 36.539
R7087 VDD.n4796 VDD.t179 36.539
R7088 VDD.n3423 VDD.t256 36.539
R7089 VDD.n2707 VDD.t453 36.539
R7090 VDD.n3289 VDD.t178 36.539
R7091 VDD.n2930 VDD.t39 36.1587
R7092 VDD.n2930 VDD.t327 36.1587
R7093 VDD.n3176 VDD.t13 36.1587
R7094 VDD.n3176 VDD.t574 36.1587
R7095 VDD.n4166 VDD.n4165 34.211
R7096 VDD.n830 VDD.t639 33.9291
R7097 VDD.n1387 VDD.t382 33.9291
R7098 VDD.n2280 VDD.t443 33.9291
R7099 VDD.n4755 VDD.t575 33.9291
R7100 VDD.n4000 VDD.t446 31.831
R7101 VDD.n3912 VDD.t37 31.831
R7102 VDD.n3713 VDD.t260 31.831
R7103 VDD.n423 VDD.t15 31.831
R7104 VDD.n957 VDD.t713 31.831
R7105 VDD.n1742 VDD.t644 31.831
R7106 VDD.n1900 VDD.t9 31.831
R7107 VDD.n4183 VDD.t358 31.831
R7108 VDD.n4301 VDD.t360 31.831
R7109 VDD.n4479 VDD.t53 31.831
R7110 VDD.n4625 VDD.t650 31.831
R7111 VDD.n2013 VDD.t334 31.831
R7112 VDD.n1573 VDD.t151 31.831
R7113 VDD.n1061 VDD.t499 31.831
R7114 VDD.n4859 VDD.t545 31.6672
R7115 VDD.n108 VDD.t525 31.6672
R7116 VDD.n2950 VDD.t425 31.6672
R7117 VDD.n2981 VDD.t431 31.6672
R7118 VDD.n2176 VDD.t255 31.3192
R7119 VDD.n2389 VDD.t35 31.3192
R7120 VDD.n1516 VDD.n1515 30.4106
R7121 VDD.n260 VDD.t268 28.7575
R7122 VDD.n3214 VDD.t245 28.7575
R7123 VDD.n3360 VDD.t693 28.7575
R7124 VDD.n3443 VDD.t41 28.7575
R7125 VDD.n3454 VDD.t408 28.7575
R7126 VDD.n2735 VDD.t274 28.7575
R7127 VDD.n313 VDD.t232 28.7575
R7128 VDD.n279 VDD.t676 28.7575
R7129 VDD.n1498 VDD.t208 28.7575
R7130 VDD.n1440 VDD.t320 28.7575
R7131 VDD.n221 VDD.t624 28.7575
R7132 VDD.n209 VDD.t18 28.7575
R7133 VDD.n4764 VDD.t55 28.7575
R7134 VDD.n172 VDD.t336 28.7575
R7135 VDD.n816 VDD.n815 28.7093
R7136 VDD.n830 VDD.n829 28.7093
R7137 VDD.n847 VDD.n846 28.7093
R7138 VDD.n875 VDD.n874 28.7093
R7139 VDD.n910 VDD.n909 28.7093
R7140 VDD.n890 VDD.n889 28.7093
R7141 VDD.n1206 VDD.n274 28.7093
R7142 VDD.n1209 VDD.n1208 28.7093
R7143 VDD.n1370 VDD.n1369 28.7093
R7144 VDD.n1387 VDD.n1386 28.7093
R7145 VDD.n1405 VDD.n1404 28.7093
R7146 VDD.n1656 VDD.n1655 28.7093
R7147 VDD.n1687 VDD.n1686 28.7093
R7148 VDD.n1671 VDD.n1670 28.7093
R7149 VDD.n1507 VDD.n1493 28.7093
R7150 VDD.n1510 VDD.n1509 28.7093
R7151 VDD.n3460 VDD.t740 28.7093
R7152 VDD.n3364 VDD.t645 28.7093
R7153 VDD.n1800 VDD.t234 28.0332
R7154 VDD.n1775 VDD.t470 28.0332
R7155 VDD.n971 VDD.t462 28.0332
R7156 VDD.n437 VDD.t316 28.0332
R7157 VDD.n3727 VDD.t185 28.0332
R7158 VDD.n3926 VDD.t354 28.0332
R7159 VDD.n4014 VDD.t278 28.0332
R7160 VDD.n719 VDD.t43 28.0332
R7161 VDD.n1558 VDD.t719 28.0332
R7162 VDD.n2029 VDD.t478 28.0332
R7163 VDD.n4639 VDD.t632 28.0332
R7164 VDD.n4495 VDD.t63 28.0332
R7165 VDD.n4367 VDD.t210 28.0332
R7166 VDD.n4143 VDD.t309 28.0332
R7167 VDD.n2878 VDD.t159 26.5955
R7168 VDD.n2878 VDD.t262 26.5955
R7169 VDD.n2856 VDD.t157 26.5955
R7170 VDD.n2856 VDD.t155 26.5955
R7171 VDD.n2816 VDD.t655 26.5955
R7172 VDD.n2816 VDD.t659 26.5955
R7173 VDD.n47 VDD.t657 26.5955
R7174 VDD.n47 VDD.t661 26.5955
R7175 VDD.n41 VDD.t524 26.5955
R7176 VDD.n41 VDD.t663 26.5955
R7177 VDD.n31 VDD.t528 26.5955
R7178 VDD.n31 VDD.t540 26.5955
R7179 VDD.n83 VDD.t516 26.5955
R7180 VDD.n83 VDD.t538 26.5955
R7181 VDD.n66 VDD.t518 26.5955
R7182 VDD.n66 VDD.t544 26.5955
R7183 VDD.n124 VDD.t522 26.5955
R7184 VDD.n124 VDD.t534 26.5955
R7185 VDD.n110 VDD.t526 26.5955
R7186 VDD.n110 VDD.t536 26.5955
R7187 VDD.n101 VDD.t530 26.5955
R7188 VDD.n101 VDD.t542 26.5955
R7189 VDD.n4857 VDD.t520 26.5955
R7190 VDD.n4857 VDD.t546 26.5955
R7191 VDD.n3190 VDD.t490 26.5955
R7192 VDD.n3190 VDD.t342 26.5955
R7193 VDD.n3139 VDD.t484 26.5955
R7194 VDD.n3139 VDD.t488 26.5955
R7195 VDD.n3108 VDD.t682 26.5955
R7196 VDD.n3108 VDD.t688 26.5955
R7197 VDD.n2779 VDD.t684 26.5955
R7198 VDD.n2779 VDD.t678 26.5955
R7199 VDD.n3080 VDD.t440 26.5955
R7200 VDD.n3080 VDD.t680 26.5955
R7201 VDD.n3066 VDD.t434 26.5955
R7202 VDD.n3066 VDD.t420 26.5955
R7203 VDD.n3041 VDD.t410 26.5955
R7204 VDD.n3041 VDD.t424 26.5955
R7205 VDD.n3026 VDD.t412 26.5955
R7206 VDD.n3026 VDD.t428 26.5955
R7207 VDD.n2986 VDD.t430 26.5955
R7208 VDD.n2986 VDD.t414 26.5955
R7209 VDD.n2979 VDD.t432 26.5955
R7210 VDD.n2979 VDD.t418 26.5955
R7211 VDD.n2955 VDD.t436 26.5955
R7212 VDD.n2955 VDD.t422 26.5955
R7213 VDD.n2948 VDD.t438 26.5955
R7214 VDD.n2948 VDD.t426 26.5955
R7215 VDD.n321 VDD.n320 26.2219
R7216 VDD.n320 VDD.n319 26.1149
R7217 VDD.n3328 VDD.n3325 24.0332
R7218 VDD.n2743 VDD.n2740 24.0332
R7219 VDD.n2746 VDD.n2743 24.0332
R7220 VDD.n2749 VDD.n2746 24.0332
R7221 VDD.n2752 VDD.n2749 24.0332
R7222 VDD.n3506 VDD.n3503 24.0332
R7223 VDD.n3503 VDD.n3500 24.0332
R7224 VDD.n3500 VDD.n3497 24.0332
R7225 VDD.n2689 VDD.n2686 24.0332
R7226 VDD.n2692 VDD.n2689 24.0332
R7227 VDD.n797 VDD.n794 24.0332
R7228 VDD.n800 VDD.n797 24.0332
R7229 VDD.n803 VDD.n800 24.0332
R7230 VDD.n806 VDD.n803 24.0332
R7231 VDD.n809 VDD.n806 24.0332
R7232 VDD.n1217 VDD.n1214 24.0332
R7233 VDD.n1354 VDD.n1351 24.0332
R7234 VDD.n1357 VDD.n1354 24.0332
R7235 VDD.n1360 VDD.n1357 24.0332
R7236 VDD.n1363 VDD.n1360 24.0332
R7237 VDD.n2223 VDD.n2220 24.0332
R7238 VDD.n2220 VDD.n2217 24.0332
R7239 VDD.n2241 VDD.n2238 24.0332
R7240 VDD.n2244 VDD.n2241 24.0332
R7241 VDD.n2247 VDD.n2244 24.0332
R7242 VDD.n2408 VDD.n2405 24.0332
R7243 VDD.n2405 VDD.n2402 24.0332
R7244 VDD.n4716 VDD.n4713 24.0332
R7245 VDD.n4719 VDD.n4716 24.0332
R7246 VDD.n4722 VDD.n4719 24.0332
R7247 VDD.n2294 VDD.n220 23.7899
R7248 VDD.n4772 VDD.n4763 23.7899
R7249 VDD.n472 VDD.t625 23.7505
R7250 VDD.n1006 VDD.t585 23.7505
R7251 VDD.n1958 VDD.t263 23.7505
R7252 VDD.n3644 VDD.t706 23.7505
R7253 VDD.n3819 VDD.t331 23.7505
R7254 VDD.n3965 VDD.t183 23.7505
R7255 VDD.n4049 VDD.t552 23.7505
R7256 VDD.n320 VDD.n317 23.7154
R7257 VDD.n3376 VDD.n3373 23.7089
R7258 VDD.n568 VDD.t242 23.6847
R7259 VDD.n1110 VDD.t252 23.6847
R7260 VDD.n2073 VDD.t294 23.6847
R7261 VDD.n4678 VDD.t595 23.6847
R7262 VDD.n2580 VDD.t224 23.6847
R7263 VDD.n4325 VDD.t86 23.6847
R7264 VDD.n4229 VDD.t733 23.6847
R7265 VDD.n794 VDD.n791 23.245
R7266 VDD.n1336 VDD.n1335 22.9432
R7267 VDD.n2755 VDD.n2752 22.1686
R7268 VDD.n3377 VDD.n3376 22.1686
R7269 VDD.n3411 VDD.n3408 22.1686
R7270 VDD.n3450 VDD.n3442 22.1686
R7271 VDD.n2695 VDD.n2692 22.1686
R7272 VDD.n810 VDD.n809 21.7362
R7273 VDD.n1364 VDD.n1363 21.7362
R7274 VDD.n813 VDD.n812 21.177
R7275 VDD.n827 VDD.n826 21.177
R7276 VDD.n844 VDD.n843 21.177
R7277 VDD.n858 VDD.n857 21.177
R7278 VDD.n872 VDD.n871 21.177
R7279 VDD.n907 VDD.n906 21.177
R7280 VDD.n887 VDD.n886 21.177
R7281 VDD.n276 VDD.n275 21.177
R7282 VDD.n1207 VDD.n272 21.177
R7283 VDD.n1367 VDD.n1366 21.177
R7284 VDD.n1384 VDD.n1383 21.177
R7285 VDD.n1402 VDD.n1401 21.177
R7286 VDD.n1639 VDD.n1638 21.177
R7287 VDD.n1653 VDD.n1652 21.177
R7288 VDD.n1684 VDD.n1683 21.177
R7289 VDD.n1668 VDD.n1667 21.177
R7290 VDD.n1495 VDD.n1494 21.177
R7291 VDD.n1508 VDD.n1491 21.177
R7292 VDD.n27 VDD.t539 21.1116
R7293 VDD.n54 VDD.t662 21.1116
R7294 VDD.n3069 VDD.t419 21.1116
R7295 VDD.n3076 VDD.t679 21.1116
R7296 VDD.t34 VDD.n860 20.8796
R7297 VDD.t497 VDD.n1641 20.8796
R7298 VDD VDD.n3459 20.8796
R7299 VDD VDD.n3363 20.8796
R7300 VDD.n3711 VDD.n3630 20.3039
R7301 VDD.n4621 VDD.n4620 20.3039
R7302 VDD.n4776 VDD.n173 19.8626
R7303 VDD.n2224 VDD.n2223 18.7186
R7304 VDD.n2409 VDD.n2408 18.7186
R7305 VDD.n2193 VDD.t598 18.2697
R7306 VDD.n2447 VDD.t367 18.2697
R7307 VDD.n3183 VDD 16.7729
R7308 VDD.n597 VDD.t500 15.8338
R7309 VDD.n1024 VDD.t199 15.8338
R7310 VDD.n1942 VDD.t283 15.8338
R7311 VDD.n3662 VDD.t694 15.8338
R7312 VDD.n3850 VDD.t289 15.8338
R7313 VDD.n3532 VDD.t227 15.8338
R7314 VDD.n4067 VDD.t700 15.8338
R7315 VDD.n552 VDD.t6 15.79
R7316 VDD.n1128 VDD.t347 15.79
R7317 VDD.n2091 VDD.t50 15.79
R7318 VDD.n2504 VDD.t403 15.79
R7319 VDD.n4573 VDD.t491 15.79
R7320 VDD.n4424 VDD.t619 15.79
R7321 VDD.n4247 VDD.t726 15.79
R7322 VDD.n815 VDD.n814 15.6598
R7323 VDD.n829 VDD.n828 15.6598
R7324 VDD.n846 VDD.n845 15.6598
R7325 VDD.n860 VDD.n859 15.6598
R7326 VDD.n874 VDD.n873 15.6598
R7327 VDD.n909 VDD.n908 15.6598
R7328 VDD.n889 VDD.n888 15.6598
R7329 VDD.n274 VDD.n273 15.6598
R7330 VDD.n1208 VDD 15.6598
R7331 VDD.n1369 VDD.n1368 15.6598
R7332 VDD.n1386 VDD.n1385 15.6598
R7333 VDD.n1404 VDD.n1403 15.6598
R7334 VDD.n1641 VDD.n1640 15.6598
R7335 VDD.n1655 VDD.n1654 15.6598
R7336 VDD.n1686 VDD.n1685 15.6598
R7337 VDD.n1670 VDD.n1669 15.6598
R7338 VDD.n1493 VDD.n1492 15.6598
R7339 VDD.n1509 VDD 15.6598
R7340 VDD.n4792 VDD.t384 15.6598
R7341 VDD.n3419 VDD.t465 15.6598
R7342 VDD.n3459 VDD.t407 15.6598
R7343 VDD.n2711 VDD.t590 15.6598
R7344 VDD.n3363 VDD.t692 15.6598
R7345 VDD.n3285 VDD.t447 15.6598
R7346 VDD.n1214 VDD.n268 13.8904
R7347 VDD.n1218 VDD.n1217 13.7733
R7348 VDD.n4168 VDD.n4164 13.7148
R7349 VDD.n537 VDD 13.6005
R7350 VDD.n1144 VDD 13.6005
R7351 VDD.n2107 VDD 13.6005
R7352 VDD.n2495 VDD 13.6005
R7353 VDD.n2557 VDD 13.6005
R7354 VDD.n4441 VDD 13.6005
R7355 VDD.n4263 VDD 13.6005
R7356 VDD.n306 VDD.n305 12.8005
R7357 VDD.n1230 VDD.n261 12.8005
R7358 VDD.n1442 VDD.n1441 12.8005
R7359 VDD.n2305 VDD.n208 12.8005
R7360 VDD.n315 VDD.n314 12.5798
R7361 VDD.n501 VDD.n497 12.5798
R7362 VDD.n4295 VDD.n2626 12.5798
R7363 VDD.n4473 VDD.n2591 12.5798
R7364 VDD.n4620 VDD.n2535 12.5798
R7365 VDD.n1180 VDD.n1072 12.5798
R7366 VDD.n3329 VDD.n3328 12.242
R7367 VDD.n3507 VDD.n3506 12.242
R7368 VDD.n3370 VDD.n2737 11.9177
R7369 VDD.n3367 VDD.n3366 11.9177
R7370 VDD.n3457 VDD.n3453 11.9177
R7371 VDD.n2251 VDD.n2247 11.7196
R7372 VDD.n4726 VDD.n4722 11.7196
R7373 VDD.n468 VDD.t313 10.5561
R7374 VDD.n1002 VDD.t459 10.5561
R7375 VDD.n1962 VDD.t467 10.5561
R7376 VDD.n3633 VDD.t237 10.5561
R7377 VDD.n3804 VDD.t188 10.5561
R7378 VDD.n3959 VDD.t351 10.5561
R7379 VDD.n4045 VDD.t275 10.5561
R7380 VDD.n97 VDD.t529 10.5561
R7381 VDD.n103 VDD.t541 10.5561
R7382 VDD.n2963 VDD.t435 10.5561
R7383 VDD.n2957 VDD.t421 10.5561
R7384 VDD.n675 VDD.t44 10.5268
R7385 VDD.n1106 VDD.t716 10.5268
R7386 VDD.n2069 VDD.t479 10.5268
R7387 VDD.n4674 VDD.t633 10.5268
R7388 VDD.n2584 VDD.t60 10.5268
R7389 VDD.n4329 VDD.t211 10.5268
R7390 VDD.n4224 VDD.t306 10.5268
R7391 VDD.n4167 VDD.n4166 10.5268
R7392 VDD.t255 VDD.n2175 10.4401
R7393 VDD.t623 VDD.n2291 10.4401
R7394 VDD.t35 VDD.n2388 10.4401
R7395 VDD.t54 VDD.n4769 10.4401
R7396 VDD.n3287 VDD.n3284 10.1522
R7397 VDD.n3341 VDD.n3340 10.1522
R7398 VDD.n3417 VDD.n3414 10.1522
R7399 VDD.n2263 VDD.n2259 10.1522
R7400 VDD.n4819 VDD.n4816 10.1522
R7401 VDD.n105 VDD.n102 10.1522
R7402 VDD.n2959 VDD.n2956 10.1522
R7403 VDD.n403 VDD.n402 9.93153
R7404 VDD.n535 VDD.n534 9.3005
R7405 VDD.n534 VDD.n532 9.3005
R7406 VDD.n1142 VDD.n1141 9.3005
R7407 VDD.n1141 VDD.n1139 9.3005
R7408 VDD.n2105 VDD.n2104 9.3005
R7409 VDD.n2104 VDD.n2102 9.3005
R7410 VDD.n2493 VDD.n2492 9.3005
R7411 VDD.n2492 VDD.n2490 9.3005
R7412 VDD.n2555 VDD.n2554 9.3005
R7413 VDD.n2554 VDD.n2552 9.3005
R7414 VDD.n4439 VDD.n4438 9.3005
R7415 VDD.n4438 VDD.n4436 9.3005
R7416 VDD.n4261 VDD.n4260 9.3005
R7417 VDD.n4260 VDD.n4258 9.3005
R7418 VDD.n741 VDD.n740 9.3005
R7419 VDD.n740 VDD.n739 9.3005
R7420 VDD.n4153 VDD.n4152 9.3005
R7421 VDD.n4152 VDD.n4151 9.3005
R7422 VDD.n4169 VDD.n4168 9.3005
R7423 VDD.n4168 VDD.n4167 9.3005
R7424 VDD.n4376 VDD.n4375 9.3005
R7425 VDD.n4375 VDD.n4374 9.3005
R7426 VDD.n4359 VDD.n4358 9.3005
R7427 VDD.n4358 VDD.n4357 9.3005
R7428 VDD.n4505 VDD.n4504 9.3005
R7429 VDD.n4504 VDD.n4503 9.3005
R7430 VDD.n4649 VDD.n4647 9.3005
R7431 VDD.n4647 VDD.n4646 9.3005
R7432 VDD.n2039 VDD.n2038 9.3005
R7433 VDD.n2038 VDD.n2037 9.3005
R7434 VDD.n2053 VDD.n2052 9.3005
R7435 VDD.n2052 VDD.n2051 9.3005
R7436 VDD.n789 VDD.n788 9.3005
R7437 VDD.n788 VDD.n787 9.3005
R7438 VDD.n410 VDD.n409 9.3005
R7439 VDD.n409 VDD.n408 9.3005
R7440 VDD.n396 VDD.n395 9.3005
R7441 VDD.n395 VDD.n394 9.3005
R7442 VDD.n382 VDD.n381 9.3005
R7443 VDD.n381 VDD.n380 9.3005
R7444 VDD.n368 VDD.n367 9.3005
R7445 VDD.n367 VDD.n366 9.3005
R7446 VDD.n354 VDD.n353 9.3005
R7447 VDD.n353 VDD.n352 9.3005
R7448 VDD.n340 VDD.n339 9.3005
R7449 VDD.n339 VDD.n338 9.3005
R7450 VDD.n326 VDD.n325 9.3005
R7451 VDD.n325 VDD.n324 9.3005
R7452 VDD.n818 VDD.n817 9.3005
R7453 VDD.n817 VDD.n816 9.3005
R7454 VDD.n849 VDD.n848 9.3005
R7455 VDD.n848 VDD.n847 9.3005
R7456 VDD.n863 VDD.n862 9.3005
R7457 VDD.n862 VDD.n861 9.3005
R7458 VDD.n877 VDD.n876 9.3005
R7459 VDD.n876 VDD.n875 9.3005
R7460 VDD.n912 VDD.n911 9.3005
R7461 VDD.n911 VDD.n910 9.3005
R7462 VDD.n892 VDD.n891 9.3005
R7463 VDD.n891 VDD.n890 9.3005
R7464 VDD.n1205 VDD.n1204 9.3005
R7465 VDD.n1206 VDD.n1205 9.3005
R7466 VDD.n1211 VDD.n1210 9.3005
R7467 VDD.n1210 VDD.n1209 9.3005
R7468 VDD.n1233 VDD.n1232 9.3005
R7469 VDD.n1234 VDD.n1233 9.3005
R7470 VDD.n1241 VDD.n1240 9.3005
R7471 VDD.n1240 VDD.n1239 9.3005
R7472 VDD.n1255 VDD.n1254 9.3005
R7473 VDD.n1254 VDD.n1253 9.3005
R7474 VDD.n1269 VDD.n1268 9.3005
R7475 VDD.n1268 VDD.n1267 9.3005
R7476 VDD.n1283 VDD.n1282 9.3005
R7477 VDD.n1282 VDD.n1281 9.3005
R7478 VDD.n1297 VDD.n1296 9.3005
R7479 VDD.n1296 VDD.n1295 9.3005
R7480 VDD.n1313 VDD.n1312 9.3005
R7481 VDD.n1312 VDD.n1311 9.3005
R7482 VDD.n1327 VDD.n1326 9.3005
R7483 VDD.n1326 VDD.n1325 9.3005
R7484 VDD.n1344 VDD.n1343 9.3005
R7485 VDD.n1343 VDD.n1342 9.3005
R7486 VDD.n1372 VDD.n1371 9.3005
R7487 VDD.n1371 VDD.n1370 9.3005
R7488 VDD.n1389 VDD.n1388 9.3005
R7489 VDD.n1388 VDD.n1387 9.3005
R7490 VDD.n1407 VDD.n1406 9.3005
R7491 VDD.n1406 VDD.n1405 9.3005
R7492 VDD.n1876 VDD.n1875 9.3005
R7493 VDD.n1875 VDD.n1874 9.3005
R7494 VDD.n1858 VDD.n1857 9.3005
R7495 VDD.n1857 VDD.n1856 9.3005
R7496 VDD.n201 VDD.n200 9.3005
R7497 VDD.n200 VDD.n199 9.3005
R7498 VDD.n2316 VDD.n2315 9.3005
R7499 VDD.n2315 VDD.n2314 9.3005
R7500 VDD.n2308 VDD.n2307 9.3005
R7501 VDD.n2309 VDD.n2308 9.3005
R7502 VDD.n2232 VDD.n2231 9.3005
R7503 VDD.n2231 VDD.n2230 9.3005
R7504 VDD.n2209 VDD.n2208 9.3005
R7505 VDD.n2208 VDD.n2207 9.3005
R7506 VDD.n2195 VDD.n2194 9.3005
R7507 VDD.n2194 VDD.n2193 9.3005
R7508 VDD.n2179 VDD.n2178 9.3005
R7509 VDD.n2178 VDD.n2177 9.3005
R7510 VDD.n2165 VDD.n2164 9.3005
R7511 VDD.n2164 VDD.n2163 9.3005
R7512 VDD.n223 VDD.n222 9.3005
R7513 VDD.n235 VDD.n234 9.3005
R7514 VDD.n234 VDD.n233 9.3005
R7515 VDD.n1461 VDD.n1460 9.3005
R7516 VDD.n1460 VDD.n1459 9.3005
R7517 VDD.n1476 VDD.n1475 9.3005
R7518 VDD.n1477 VDD.n1476 9.3005
R7519 VDD.n1482 VDD.n1481 9.3005
R7520 VDD.n1481 VDD.n1480 9.3005
R7521 VDD.n1512 VDD.n1511 9.3005
R7522 VDD.n1511 VDD.n1510 9.3005
R7523 VDD.n1506 VDD.n1505 9.3005
R7524 VDD.n1507 VDD.n1506 9.3005
R7525 VDD.n1673 VDD.n1672 9.3005
R7526 VDD.n1672 VDD.n1671 9.3005
R7527 VDD.n1689 VDD.n1688 9.3005
R7528 VDD.n1688 VDD.n1687 9.3005
R7529 VDD.n1658 VDD.n1657 9.3005
R7530 VDD.n1657 VDD.n1656 9.3005
R7531 VDD.n1644 VDD.n1643 9.3005
R7532 VDD.n1643 VDD.n1642 9.3005
R7533 VDD.n2392 VDD.n2391 9.3005
R7534 VDD.n2391 VDD.n2390 9.3005
R7535 VDD.n2449 VDD.n2448 9.3005
R7536 VDD.n2448 VDD.n2447 9.3005
R7537 VDD.n2431 VDD.n2430 9.3005
R7538 VDD.n2430 VDD.n2429 9.3005
R7539 VDD.n2417 VDD.n2416 9.3005
R7540 VDD.n2416 VDD.n2415 9.3005
R7541 VDD.n832 VDD.n831 9.3005
R7542 VDD.n831 VDD.n830 9.3005
R7543 VDD.n44 VDD.n42 9.26947
R7544 VDD.n3083 VDD.n3081 9.26947
R7545 VDD.n539 VDD.n538 8.94661
R7546 VDD.n1146 VDD.n1145 8.94661
R7547 VDD.n2109 VDD.n2108 8.94661
R7548 VDD.n2497 VDD.n2496 8.94661
R7549 VDD.n2559 VDD.n2558 8.94661
R7550 VDD.n4443 VDD.n4442 8.94661
R7551 VDD.n4265 VDD.n4264 8.94661
R7552 VDD.n2251 VDD.n2250 8.82809
R7553 VDD.n2256 VDD.n2255 8.82809
R7554 VDD.n2263 VDD.n2262 8.82809
R7555 VDD.n2268 VDD.n2267 8.82809
R7556 VDD.n2273 VDD.n2272 8.82809
R7557 VDD.n2278 VDD.n2277 8.82809
R7558 VDD.n2283 VDD.n2282 8.82809
R7559 VDD.n4726 VDD.n4725 8.82809
R7560 VDD.n4733 VDD.n4732 8.82809
R7561 VDD.n4738 VDD.n4737 8.82809
R7562 VDD.n4743 VDD.n4742 8.82809
R7563 VDD.n4748 VDD.n4747 8.82809
R7564 VDD.n4753 VDD.n4752 8.82809
R7565 VDD.n4758 VDD.n4757 8.82809
R7566 VDD.n4773 VDD.n4772 8.82809
R7567 VDD.n1395 VDD.n1394 8.6074
R7568 VDD.n947 VDD.n946 8.47281
R7569 VDD.n1732 VDD.n1731 8.47281
R7570 VDD.n1798 VDD.n1797 8.47281
R7571 VDD.n2929 VDD.n2928 8.47281
R7572 VDD.n3179 VDD.n3178 8.47281
R7573 VDD.n3706 VDD.n3705 8.47276
R7574 VDD.n2859 VDD.n2858 8.47276
R7575 VDD.n3142 VDD.n3141 8.47276
R7576 VDD.n1072 VDD.n1071 8.47276
R7577 VDD.n3990 VDD.n3989 8.47181
R7578 VDD.n3250 VDD.n3249 8.47181
R7579 VDD.n3902 VDD.n3901 8.47181
R7580 VDD.n501 VDD.n500 8.47181
R7581 VDD.n2626 VDD.n2625 8.47181
R7582 VDD.n2591 VDD.n2590 8.47181
R7583 VDD.n2535 VDD.n2534 8.47181
R7584 VDD.n2344 VDD.n2343 8.47181
R7585 VDD.n1595 VDD.n1594 8.47181
R7586 VDD.n510 VDD.n509 8.47137
R7587 VDD.n293 VDD.n292 8.47133
R7588 VDD.n1793 VDD.n1792 8.47133
R7589 VDD.n3694 VDD.n3693 8.47133
R7590 VDD.n1721 VDD.n1720 8.47133
R7591 VDD.n1171 VDD.n1170 8.47133
R7592 VDD.n2675 VDD.n2674 8.47037
R7593 VDD.n3243 VDD.n3242 8.47037
R7594 VDD.n3892 VDD.n3891 8.47037
R7595 VDD.n2631 VDD.n2630 8.47037
R7596 VDD.n2596 VDD.n2595 8.47037
R7597 VDD.n4609 VDD.n4608 8.47037
R7598 VDD.n2353 VDD.n2352 8.47037
R7599 VDD.n1608 VDD.n1607 8.47037
R7600 VDD.n4096 VDD.n4095 8.47012
R7601 VDD.n2470 VDD.n2469 8.47011
R7602 VDD.n683 VDD.n682 8.47011
R7603 VDD.n465 VDD.n464 8.47007
R7604 VDD.n628 VDD.n627 8.47007
R7605 VDD.n1784 VDD.n1783 8.47007
R7606 VDD.n1789 VDD.n1788 8.47007
R7607 VDD.n3677 VDD.n3676 8.47007
R7608 VDD.n1041 VDD.n1040 8.47007
R7609 VDD.n999 VDD.n998 8.47007
R7610 VDD.n3954 VDD.n3953 8.46911
R7611 VDD.n4042 VDD.n4041 8.46911
R7612 VDD.n3875 VDD.n3874 8.46911
R7613 VDD.n3801 VDD.n3800 8.46911
R7614 VDD.n1103 VDD.n1102 8.46911
R7615 VDD.n2641 VDD.n2640 8.46911
R7616 VDD.n4338 VDD.n4337 8.46911
R7617 VDD.n4530 VDD.n4529 8.46911
R7618 VDD.n4671 VDD.n4670 8.46911
R7619 VDD.n2008 VDD.n2007 8.46911
R7620 VDD.n4128 VDD.n4127 8.46584
R7621 VDD.n2701 VDD.n2700 8.45089
R7622 VDD.n2700 VDD.n2699 8.45089
R7623 VDD.n3379 VDD.n3378 8.45089
R7624 VDD.n3381 VDD.n3380 8.45089
R7625 VDD.n3385 VDD.n3384 8.45089
R7626 VDD.n3390 VDD.n3389 8.45089
R7627 VDD.n2730 VDD.n2729 8.45089
R7628 VDD.n2708 VDD.n2707 8.45089
R7629 VDD.n2712 VDD.n2711 8.45089
R7630 VDD.n3278 VDD.n3277 8.45089
R7631 VDD.n3290 VDD.n3289 8.45089
R7632 VDD.n3300 VDD.n3299 8.45089
R7633 VDD.n3219 VDD.n3218 8.45089
R7634 VDD.n3306 VDD.n3305 8.45089
R7635 VDD.n3294 VDD.n3293 8.45089
R7636 VDD.n3286 VDD.n3285 8.45089
R7637 VDD.n2754 VDD.n2753 8.45089
R7638 VDD.n2694 VDD.n2693 8.45089
R7639 VDD.n3410 VDD.n3409 8.45089
R7640 VDD.n3449 VDD.n3448 8.45089
R7641 VDD.n3447 VDD.n3446 8.45089
R7642 VDD.n3436 VDD.n3435 8.45089
R7643 VDD.n3432 VDD.n3431 8.45089
R7644 VDD.n3428 VDD.n3427 8.45089
R7645 VDD.n3424 VDD.n3423 8.45089
R7646 VDD.n3420 VDD.n3419 8.45089
R7647 VDD.n3416 VDD.n3415 8.45089
R7648 VDD.n4780 VDD.n4779 8.45089
R7649 VDD.n4784 VDD.n4783 8.45089
R7650 VDD.n4803 VDD.n4802 8.45089
R7651 VDD.n4797 VDD.n4796 8.45089
R7652 VDD.n4818 VDD.n4817 8.45089
R7653 VDD.n4824 VDD.n4823 8.45089
R7654 VDD.n4793 VDD.n4792 8.45089
R7655 VDD.n4788 VDD.n4787 8.45089
R7656 VDD.n4778 VDD.n4777 8.45089
R7657 VDD.n2469 VDD.n2468 8.45089
R7658 VDD.n3646 VDD.n3645 8.45089
R7659 VDD.n3645 VDD.n3644 8.45089
R7660 VDD.n3649 VDD.n3648 8.45089
R7661 VDD.n3534 VDD.n3533 8.45089
R7662 VDD.n3533 VDD.n3532 8.45089
R7663 VDD.n3564 VDD.n3563 8.45089
R7664 VDD.n3569 VDD.n3568 8.45089
R7665 VDD.n3559 VDD.n3558 8.45089
R7666 VDD.n3966 VDD.n3965 8.45089
R7667 VDD.n3960 VDD.n3959 8.45089
R7668 VDD.n3953 VDD.n3952 8.45089
R7669 VDD.n3948 VDD.n3947 8.45089
R7670 VDD.n3944 VDD.n3943 8.45089
R7671 VDD.n3939 VDD.n3938 8.45089
R7672 VDD.n3546 VDD.n3545 8.45089
R7673 VDD.n3606 VDD.n3605 8.45089
R7674 VDD.n3611 VDD.n3610 8.45089
R7675 VDD.n2674 VDD.n2673 8.45089
R7676 VDD.n3620 VDD.n3619 8.45089
R7677 VDD.n3616 VDD.n3615 8.45089
R7678 VDD.n3984 VDD.n3983 8.45089
R7679 VDD.n3989 VDD.n3988 8.45089
R7680 VDD.n3997 VDD.n3996 8.45089
R7681 VDD.n4003 VDD.n4002 8.45089
R7682 VDD.n4011 VDD.n4010 8.45089
R7683 VDD.n4033 VDD.n4032 8.45089
R7684 VDD.n4032 VDD.n4031 8.45089
R7685 VDD.n4041 VDD.n4040 8.45089
R7686 VDD.n4050 VDD.n4049 8.45089
R7687 VDD.n4058 VDD.n4057 8.45089
R7688 VDD.n4068 VDD.n4067 8.45089
R7689 VDD.n4089 VDD.n4088 8.45089
R7690 VDD.n4100 VDD.n4099 8.45089
R7691 VDD.n2658 VDD.n2657 8.45089
R7692 VDD.n3242 VDD.n3241 8.45089
R7693 VDD.n3251 VDD.n3250 8.45089
R7694 VDD.n3257 VDD.n3256 8.45089
R7695 VDD.n2652 VDD.n2651 8.45089
R7696 VDD.n4095 VDD.n4094 8.45089
R7697 VDD.n4075 VDD.n4074 8.45089
R7698 VDD.n4062 VDD.n4061 8.45089
R7699 VDD.n4054 VDD.n4053 8.45089
R7700 VDD.n4046 VDD.n4045 8.45089
R7701 VDD.n4036 VDD.n4035 8.45089
R7702 VDD.n4028 VDD.n4027 8.45089
R7703 VDD.n4007 VDD.n4006 8.45089
R7704 VDD.n3540 VDD.n3539 8.45089
R7705 VDD.n3924 VDD.n3923 8.45089
R7706 VDD.n3923 VDD.n3922 8.45089
R7707 VDD.n3919 VDD.n3918 8.45089
R7708 VDD.n3915 VDD.n3914 8.45089
R7709 VDD.n3909 VDD.n3908 8.45089
R7710 VDD.n3901 VDD.n3900 8.45089
R7711 VDD.n3896 VDD.n3895 8.45089
R7712 VDD.n3891 VDD.n3890 8.45089
R7713 VDD.n3887 VDD.n3886 8.45089
R7714 VDD.n3883 VDD.n3882 8.45089
R7715 VDD.n3879 VDD.n3878 8.45089
R7716 VDD.n3874 VDD.n3873 8.45089
R7717 VDD.n3867 VDD.n3866 8.45089
R7718 VDD.n3855 VDD.n3854 8.45089
R7719 VDD.n3851 VDD.n3850 8.45089
R7720 VDD.n3845 VDD.n3844 8.45089
R7721 VDD.n3839 VDD.n3838 8.45089
R7722 VDD.n3825 VDD.n3824 8.45089
R7723 VDD.n3820 VDD.n3819 8.45089
R7724 VDD.n3805 VDD.n3804 8.45089
R7725 VDD.n3800 VDD.n3799 8.45089
R7726 VDD.n3785 VDD.n3784 8.45089
R7727 VDD.n3779 VDD.n3778 8.45089
R7728 VDD.n3742 VDD.n3741 8.45089
R7729 VDD.n3724 VDD.n3723 8.45089
R7730 VDD.n3720 VDD.n3719 8.45089
R7731 VDD.n3716 VDD.n3715 8.45089
R7732 VDD.n3710 VDD.n3709 8.45089
R7733 VDD.n3707 VDD.n3706 8.45089
R7734 VDD.n3698 VDD.n3697 8.45089
R7735 VDD.n3693 VDD.n3692 8.45089
R7736 VDD.n3689 VDD.n3688 8.45089
R7737 VDD.n3685 VDD.n3684 8.45089
R7738 VDD.n3681 VDD.n3680 8.45089
R7739 VDD.n3676 VDD.n3675 8.45089
R7740 VDD.n3671 VDD.n3670 8.45089
R7741 VDD.n3667 VDD.n3666 8.45089
R7742 VDD.n3663 VDD.n3662 8.45089
R7743 VDD.n3657 VDD.n3656 8.45089
R7744 VDD.n3653 VDD.n3652 8.45089
R7745 VDD.n3634 VDD.n3633 8.45089
R7746 VDD.n435 VDD.n434 8.45089
R7747 VDD.n434 VDD.n433 8.45089
R7748 VDD.n430 VDD.n429 8.45089
R7749 VDD.n426 VDD.n425 8.45089
R7750 VDD.n486 VDD.n485 8.45089
R7751 VDD.n485 VDD.n484 8.45089
R7752 VDD.n479 VDD.n478 8.45089
R7753 VDD.n473 VDD.n472 8.45089
R7754 VDD.n469 VDD.n468 8.45089
R7755 VDD.n464 VDD.n463 8.45089
R7756 VDD.n459 VDD.n458 8.45089
R7757 VDD.n455 VDD.n454 8.45089
R7758 VDD.n590 VDD.n589 8.45089
R7759 VDD.n604 VDD.n603 8.45089
R7760 VDD.n620 VDD.n619 8.45089
R7761 VDD.n653 VDD.n652 8.45089
R7762 VDD.n941 VDD.n940 8.45089
R7763 VDD.n292 VDD.n291 8.45089
R7764 VDD.n658 VDD.n657 8.45089
R7765 VDD.n663 VDD.n662 8.45089
R7766 VDD.n627 VDD.n626 8.45089
R7767 VDD.n598 VDD.n597 8.45089
R7768 VDD.n451 VDD.n450 8.45089
R7769 VDD.n946 VDD.n945 8.45089
R7770 VDD.n954 VDD.n953 8.45089
R7771 VDD.n960 VDD.n959 8.45089
R7772 VDD.n968 VDD.n967 8.45089
R7773 VDD.n964 VDD.n963 8.45089
R7774 VDD.n986 VDD.n985 8.45089
R7775 VDD.n985 VDD.n984 8.45089
R7776 VDD.n993 VDD.n992 8.45089
R7777 VDD.n998 VDD.n997 8.45089
R7778 VDD.n1007 VDD.n1006 8.45089
R7779 VDD.n1011 VDD.n1010 8.45089
R7780 VDD.n1019 VDD.n1018 8.45089
R7781 VDD.n1025 VDD.n1024 8.45089
R7782 VDD.n1033 VDD.n1032 8.45089
R7783 VDD.n1040 VDD.n1039 8.45089
R7784 VDD.n1712 VDD.n1711 8.45089
R7785 VDD.n1720 VDD.n1719 8.45089
R7786 VDD.n1726 VDD.n1725 8.45089
R7787 VDD.n1716 VDD.n1715 8.45089
R7788 VDD.n246 VDD.n245 8.45089
R7789 VDD.n1029 VDD.n1028 8.45089
R7790 VDD.n1015 VDD.n1014 8.45089
R7791 VDD.n1003 VDD.n1002 8.45089
R7792 VDD.n989 VDD.n988 8.45089
R7793 VDD.n1731 VDD.n1730 8.45089
R7794 VDD.n1755 VDD.n1754 8.45089
R7795 VDD.n1749 VDD.n1748 8.45089
R7796 VDD.n1745 VDD.n1744 8.45089
R7797 VDD.n1739 VDD.n1738 8.45089
R7798 VDD.n1978 VDD.n1977 8.45089
R7799 VDD.n1977 VDD.n1976 8.45089
R7800 VDD.n1972 VDD.n1971 8.45089
R7801 VDD.n1968 VDD.n1967 8.45089
R7802 VDD.n1783 VDD.n1782 8.45089
R7803 VDD.n1959 VDD.n1958 8.45089
R7804 VDD.n1951 VDD.n1950 8.45089
R7805 VDD.n1943 VDD.n1942 8.45089
R7806 VDD.n1933 VDD.n1932 8.45089
R7807 VDD.n1928 VDD.n1927 8.45089
R7808 VDD.n1920 VDD.n1919 8.45089
R7809 VDD.n1792 VDD.n1791 8.45089
R7810 VDD.n1915 VDD.n1914 8.45089
R7811 VDD.n1924 VDD.n1923 8.45089
R7812 VDD.n1788 VDD.n1787 8.45089
R7813 VDD.n1937 VDD.n1936 8.45089
R7814 VDD.n1947 VDD.n1946 8.45089
R7815 VDD.n1955 VDD.n1954 8.45089
R7816 VDD.n1963 VDD.n1962 8.45089
R7817 VDD.n1799 VDD.n1798 8.45089
R7818 VDD.n1909 VDD.n1908 8.45089
R7819 VDD.n1903 VDD.n1902 8.45089
R7820 VDD.n1807 VDD.n1806 8.45089
R7821 VDD.n1897 VDD.n1896 8.45089
R7822 VDD.n1834 VDD.n1833 8.45089
R7823 VDD.n1828 VDD.n1827 8.45089
R7824 VDD.n2465 VDD.n2464 8.45089
R7825 VDD.n2464 VDD.n2463 8.45089
R7826 VDD.n116 VDD.n115 8.45089
R7827 VDD.n115 VDD.n114 8.45089
R7828 VDD.n109 VDD.n108 8.45089
R7829 VDD.n104 VDD.n103 8.45089
R7830 VDD.n98 VDD.n97 8.45089
R7831 VDD.n4860 VDD.n4859 8.45089
R7832 VDD.n4852 VDD.n4851 8.45089
R7833 VDD.n128 VDD.n127 8.45089
R7834 VDD.n69 VDD.n68 8.45089
R7835 VDD.n80 VDD.n79 8.45089
R7836 VDD.n28 VDD.n27 8.45089
R7837 VDD.n43 VDD.t523 8.45089
R7838 VDD.n50 VDD.n49 8.45089
R7839 VDD.n55 VDD.n54 8.45089
R7840 VDD.n142 VDD.n141 8.45089
R7841 VDD.n2821 VDD.n2820 8.45089
R7842 VDD.n2881 VDD.n2880 8.45089
R7843 VDD.n2802 VDD.n2801 8.45089
R7844 VDD.n2858 VDD.n2857 8.45089
R7845 VDD.n2851 VDD.n2850 8.45089
R7846 VDD.n2844 VDD.n2843 8.45089
R7847 VDD.n2842 VDD.n2841 8.45089
R7848 VDD.n2887 VDD.n2886 8.45089
R7849 VDD.n2923 VDD.n2922 8.45089
R7850 VDD.n2922 VDD.n2921 8.45089
R7851 VDD.n2889 VDD.n2888 8.45089
R7852 VDD.n2815 VDD.n2814 8.45089
R7853 VDD.n21 VDD.n20 8.45089
R7854 VDD.n73 VDD.n72 8.45089
R7855 VDD.n120 VDD.n119 8.45089
R7856 VDD.n2928 VDD.n2927 8.45089
R7857 VDD.n3083 VDD.n3082 8.45089
R7858 VDD.n3082 VDD.t439 8.45089
R7859 VDD.n3070 VDD.n3069 8.45089
R7860 VDD.n3051 VDD.n3050 8.45089
R7861 VDD.n2945 VDD.n2944 8.45089
R7862 VDD.n2951 VDD.n2950 8.45089
R7863 VDD.n2958 VDD.n2957 8.45089
R7864 VDD.n2995 VDD.n2994 8.45089
R7865 VDD.n3012 VDD.n3011 8.45089
R7866 VDD.n3017 VDD.n3016 8.45089
R7867 VDD.n3077 VDD.n3076 8.45089
R7868 VDD.n2784 VDD.n2783 8.45089
R7869 VDD.n3115 VDD.n3114 8.45089
R7870 VDD.n3127 VDD.n3126 8.45089
R7871 VDD.n3134 VDD.n3133 8.45089
R7872 VDD.n3141 VDD.n3140 8.45089
R7873 VDD.n3193 VDD.n3192 8.45089
R7874 VDD.n3185 VDD.n3184 8.45089
R7875 VDD.n3187 VDD.n3186 8.45089
R7876 VDD.n3155 VDD.n3154 8.45089
R7877 VDD.n3129 VDD.n3128 8.45089
R7878 VDD.n3107 VDD.n3106 8.45089
R7879 VDD.n2778 VDD.n2777 8.45089
R7880 VDD.n3045 VDD.n3044 8.45089
R7881 VDD.n3023 VDD.n3022 8.45089
R7882 VDD.n2989 VDD.n2988 8.45089
R7883 VDD.n2982 VDD.n2981 8.45089
R7884 VDD.n2964 VDD.n2963 8.45089
R7885 VDD.n3178 VDD.n3177 8.45089
R7886 VDD.n3164 VDD.n3163 8.45089
R7887 VDD.n3163 VDD.n3162 8.45089
R7888 VDD.n1130 VDD.n1129 8.45089
R7889 VDD.n1129 VDD.n1128 8.45089
R7890 VDD.n1119 VDD.n1118 8.45089
R7891 VDD.n1115 VDD.n1114 8.45089
R7892 VDD.n1107 VDD.n1106 8.45089
R7893 VDD.n1102 VDD.n1101 8.45089
R7894 VDD.n1092 VDD.n1091 8.45089
R7895 VDD.n1077 VDD.n1076 8.45089
R7896 VDD.n4127 VDD.n4126 8.45089
R7897 VDD.n4122 VDD.n4121 8.45089
R7898 VDD.n2635 VDD.n2634 8.45089
R7899 VDD.n2640 VDD.n2639 8.45089
R7900 VDD.n4225 VDD.n4224 8.45089
R7901 VDD.n4230 VDD.n4229 8.45089
R7902 VDD.n4234 VDD.n4233 8.45089
R7903 VDD.n4238 VDD.n4237 8.45089
R7904 VDD.n4242 VDD.n4241 8.45089
R7905 VDD.n4248 VDD.n4247 8.45089
R7906 VDD.n4180 VDD.n4179 8.45089
R7907 VDD.n4137 VDD.n4136 8.45089
R7908 VDD.n4186 VDD.n4185 8.45089
R7909 VDD.n4252 VDD.n4251 8.45089
R7910 VDD.n4278 VDD.n4277 8.45089
R7911 VDD.n4277 VDD.n4276 8.45089
R7912 VDD.n4281 VDD.n4280 8.45089
R7913 VDD.n4285 VDD.n4284 8.45089
R7914 VDD.n2630 VDD.n2629 8.45089
R7915 VDD.n4290 VDD.n4289 8.45089
R7916 VDD.n2625 VDD.n2624 8.45089
R7917 VDD.n4298 VDD.n4297 8.45089
R7918 VDD.n4304 VDD.n4303 8.45089
R7919 VDD.n4308 VDD.n4307 8.45089
R7920 VDD.n2619 VDD.n2618 8.45089
R7921 VDD.n4337 VDD.n4336 8.45089
R7922 VDD.n4330 VDD.n4329 8.45089
R7923 VDD.n4326 VDD.n4325 8.45089
R7924 VDD.n4322 VDD.n4321 8.45089
R7925 VDD.n2600 VDD.n2599 8.45089
R7926 VDD.n2604 VDD.n2603 8.45089
R7927 VDD.n4425 VDD.n4424 8.45089
R7928 VDD.n4394 VDD.n4393 8.45089
R7929 VDD.n4404 VDD.n4403 8.45089
R7930 VDD.n4399 VDD.n4398 8.45089
R7931 VDD.n4430 VDD.n4429 8.45089
R7932 VDD.n4456 VDD.n4455 8.45089
R7933 VDD.n4455 VDD.n4454 8.45089
R7934 VDD.n4459 VDD.n4458 8.45089
R7935 VDD.n4463 VDD.n4462 8.45089
R7936 VDD.n2595 VDD.n2594 8.45089
R7937 VDD.n4468 VDD.n4467 8.45089
R7938 VDD.n2590 VDD.n2589 8.45089
R7939 VDD.n4476 VDD.n4475 8.45089
R7940 VDD.n4482 VDD.n4481 8.45089
R7941 VDD.n4486 VDD.n4485 8.45089
R7942 VDD.n4490 VDD.n4489 8.45089
R7943 VDD.n4510 VDD.n4509 8.45089
R7944 VDD.n4515 VDD.n4514 8.45089
R7945 VDD.n4519 VDD.n4518 8.45089
R7946 VDD.n4523 VDD.n4522 8.45089
R7947 VDD.n4529 VDD.n4528 8.45089
R7948 VDD.n2585 VDD.n2584 8.45089
R7949 VDD.n2581 VDD.n2580 8.45089
R7950 VDD.n2577 VDD.n2576 8.45089
R7951 VDD.n4564 VDD.n4563 8.45089
R7952 VDD.n4569 VDD.n4568 8.45089
R7953 VDD.n4574 VDD.n4573 8.45089
R7954 VDD.n4600 VDD.n4599 8.45089
R7955 VDD.n4599 VDD.n4598 8.45089
R7956 VDD.n4604 VDD.n4603 8.45089
R7957 VDD.n4608 VDD.n4607 8.45089
R7958 VDD.n4613 VDD.n4612 8.45089
R7959 VDD.n2534 VDD.n2533 8.45089
R7960 VDD.n2532 VDD.n2530 8.45089
R7961 VDD.n4624 VDD.n4623 8.45089
R7962 VDD.n4630 VDD.n4629 8.45089
R7963 VDD.n4634 VDD.n4633 8.45089
R7964 VDD.n4652 VDD.n4651 8.45089
R7965 VDD.n4657 VDD.n4656 8.45089
R7966 VDD.n4661 VDD.n4660 8.45089
R7967 VDD.n4665 VDD.n4664 8.45089
R7968 VDD.n4670 VDD.n4669 8.45089
R7969 VDD.n4675 VDD.n4674 8.45089
R7970 VDD.n4679 VDD.n4678 8.45089
R7971 VDD.n4683 VDD.n4682 8.45089
R7972 VDD.n4687 VDD.n4686 8.45089
R7973 VDD.n4692 VDD.n4691 8.45089
R7974 VDD.n2505 VDD.n2504 8.45089
R7975 VDD.n2511 VDD.n2510 8.45089
R7976 VDD.n2368 VDD.n2367 8.45089
R7977 VDD.n2367 VDD.n2366 8.45089
R7978 VDD.n2361 VDD.n2360 8.45089
R7979 VDD.n2357 VDD.n2356 8.45089
R7980 VDD.n2352 VDD.n2351 8.45089
R7981 VDD.n2348 VDD.n2347 8.45089
R7982 VDD.n2343 VDD.n2342 8.45089
R7983 VDD.n2010 VDD.n181 8.45089
R7984 VDD.n2016 VDD.n2015 8.45089
R7985 VDD.n2020 VDD.n2019 8.45089
R7986 VDD.n2024 VDD.n2023 8.45089
R7987 VDD.n2057 VDD.n2056 8.45089
R7988 VDD.n2061 VDD.n2060 8.45089
R7989 VDD.n2065 VDD.n2064 8.45089
R7990 VDD.n2007 VDD.n2006 8.45089
R7991 VDD.n2070 VDD.n2069 8.45089
R7992 VDD.n2074 VDD.n2073 8.45089
R7993 VDD.n2078 VDD.n2077 8.45089
R7994 VDD.n2082 VDD.n2081 8.45089
R7995 VDD.n2086 VDD.n2085 8.45089
R7996 VDD.n2092 VDD.n2091 8.45089
R7997 VDD.n2096 VDD.n2095 8.45089
R7998 VDD.n2121 VDD.n2120 8.45089
R7999 VDD.n2126 VDD.n2125 8.45089
R8000 VDD.n2001 VDD.n2000 8.45089
R8001 VDD.n1607 VDD.n1606 8.45089
R8002 VDD.n1601 VDD.n1600 8.45089
R8003 VDD.n1594 VDD.n1593 8.45089
R8004 VDD.n1579 VDD.n1534 8.45089
R8005 VDD.n1576 VDD.n1575 8.45089
R8006 VDD.n1570 VDD.n1569 8.45089
R8007 VDD.n1565 VDD.n1564 8.45089
R8008 VDD.n1561 VDD.n1560 8.45089
R8009 VDD.n1547 VDD.n1546 8.45089
R8010 VDD.n2537 VDD.n2536 8.45089
R8011 VDD.n4554 VDD.n4553 8.45089
R8012 VDD.n1097 VDD.n1096 8.45089
R8013 VDD.n1111 VDD.n1110 8.45089
R8014 VDD.n1123 VDD.n1122 8.45089
R8015 VDD.n1133 VDD.n1132 8.45089
R8016 VDD.n500 VDD.n499 8.45089
R8017 VDD.n506 VDD.n505 8.45089
R8018 VDD.n505 VDD.n504 8.45089
R8019 VDD.n498 VDD.n497 8.45089
R8020 VDD.n509 VDD.n508 8.45089
R8021 VDD.n518 VDD.n517 8.45089
R8022 VDD.n522 VDD.n521 8.45089
R8023 VDD.n514 VDD.n513 8.45089
R8024 VDD.n548 VDD.n547 8.45089
R8025 VDD.n547 VDD.n546 8.45089
R8026 VDD.n553 VDD.n552 8.45089
R8027 VDD.n563 VDD.n562 8.45089
R8028 VDD.n569 VDD.n568 8.45089
R8029 VDD.n1175 VDD.n1174 8.45089
R8030 VDD.n1170 VDD.n1169 8.45089
R8031 VDD.n1162 VDD.n1161 8.45089
R8032 VDD.n1158 VDD.n1157 8.45089
R8033 VDD.n1166 VDD.n1165 8.45089
R8034 VDD.n1071 VDD.n1070 8.45089
R8035 VDD.n676 VDD.n675 8.45089
R8036 VDD.n573 VDD.n572 8.45089
R8037 VDD.n557 VDD.n556 8.45089
R8038 VDD.n682 VDD.n681 8.45089
R8039 VDD.n693 VDD.n692 8.45089
R8040 VDD.n687 VDD.n686 8.45089
R8041 VDD.n725 VDD.n724 8.45089
R8042 VDD.n699 VDD.n698 8.45089
R8043 VDD.n704 VDD.n703 8.45089
R8044 VDD.n1064 VDD.n1063 8.45089
R8045 VDD.n1183 VDD.n1182 8.45089
R8046 VDD.n713 VDD.n712 8.45089
R8047 VDD.n480 VDD.n479 8.45089
R8048 VDD.n474 VDD.n473 8.45089
R8049 VDD.n470 VDD.n469 8.45089
R8050 VDD.n460 VDD.n459 8.45089
R8051 VDD.n456 VDD.n455 8.45089
R8052 VDD.n452 VDD.n451 8.45089
R8053 VDD.n599 VDD.n598 8.45089
R8054 VDD.n605 VDD.n604 8.45089
R8055 VDD.n942 VDD.n941 8.45089
R8056 VDD.n659 VDD.n658 8.45089
R8057 VDD.n952 VDD.n951 8.45089
R8058 VDD VDD.n952 8.45089
R8059 VDD.n955 VDD.n954 8.45089
R8060 VDD.n965 VDD.n964 8.45089
R8061 VDD.n969 VDD.n968 8.45089
R8062 VDD.n990 VDD.n989 8.45089
R8063 VDD.n994 VDD.n993 8.45089
R8064 VDD.n1004 VDD.n1003 8.45089
R8065 VDD.n1008 VDD.n1007 8.45089
R8066 VDD.n1016 VDD.n1015 8.45089
R8067 VDD.n1020 VDD.n1019 8.45089
R8068 VDD.n1030 VDD.n1029 8.45089
R8069 VDD.n1034 VDD.n1033 8.45089
R8070 VDD.n247 VDD.n246 8.45089
R8071 VDD.n1717 VDD.n1716 8.45089
R8072 VDD.n1757 VDD.n1755 8.45089
R8073 VDD.n1973 VDD.n1972 8.45089
R8074 VDD.n1964 VDD.n1963 8.45089
R8075 VDD.n1956 VDD.n1955 8.45089
R8076 VDD.n1948 VDD.n1947 8.45089
R8077 VDD.n1938 VDD.n1937 8.45089
R8078 VDD.n1925 VDD.n1924 8.45089
R8079 VDD.n1916 VDD.n1915 8.45089
R8080 VDD.n1911 VDD.n1910 8.45089
R8081 VDD.n1910 VDD 8.45089
R8082 VDD.n1904 VDD.n1903 8.45089
R8083 VDD.n1898 VDD.n1897 8.45089
R8084 VDD.n1835 VDD.n1834 8.45089
R8085 VDD.n3635 VDD.n3634 8.45089
R8086 VDD.n3565 VDD.n3564 8.45089
R8087 VDD.n3571 VDD.n3569 8.45089
R8088 VDD.n3560 VDD.n3559 8.45089
R8089 VDD.n3967 VDD.n3966 8.45089
R8090 VDD.n3961 VDD.n3960 8.45089
R8091 VDD.n3949 VDD.n3948 8.45089
R8092 VDD.n3945 VDD.n3944 8.45089
R8093 VDD.n3541 VDD.n3540 8.45089
R8094 VDD.n3621 VDD.n3620 8.45089
R8095 VDD.n3995 VDD.n3994 8.45089
R8096 VDD VDD.n3995 8.45089
R8097 VDD.n4004 VDD.n4003 8.45089
R8098 VDD.n4008 VDD.n4007 8.45089
R8099 VDD.n4029 VDD.n4028 8.45089
R8100 VDD.n4037 VDD.n4036 8.45089
R8101 VDD.n4047 VDD.n4046 8.45089
R8102 VDD.n4055 VDD.n4054 8.45089
R8103 VDD.n4063 VDD.n4062 8.45089
R8104 VDD.n4076 VDD.n4075 8.45089
R8105 VDD.n2653 VDD.n2652 8.45089
R8106 VDD.n3258 VDD.n3257 8.45089
R8107 VDD.n3253 VDD.n3252 8.45089
R8108 VDD.n3252 VDD 8.45089
R8109 VDD.n2659 VDD.n2658 8.45089
R8110 VDD.n4101 VDD.n4100 8.45089
R8111 VDD.n4090 VDD.n4089 8.45089
R8112 VDD.n4069 VDD.n4068 8.45089
R8113 VDD.n4059 VDD.n4058 8.45089
R8114 VDD.n4051 VDD.n4050 8.45089
R8115 VDD.n4012 VDD.n4011 8.45089
R8116 VDD.n3998 VDD.n3997 8.45089
R8117 VDD.n3985 VDD.n3984 8.45089
R8118 VDD.n3617 VDD.n3616 8.45089
R8119 VDD.n3612 VDD.n3611 8.45089
R8120 VDD.n3547 VDD.n3546 8.45089
R8121 VDD.n3941 VDD.n3939 8.45089
R8122 VDD.n3920 VDD.n3919 8.45089
R8123 VDD.n3916 VDD.n3915 8.45089
R8124 VDD.n3910 VDD.n3909 8.45089
R8125 VDD.n3907 VDD.n3906 8.45089
R8126 VDD VDD.n3907 8.45089
R8127 VDD.n3897 VDD.n3896 8.45089
R8128 VDD.n3888 VDD.n3887 8.45089
R8129 VDD.n3884 VDD.n3883 8.45089
R8130 VDD.n3880 VDD.n3879 8.45089
R8131 VDD.n3869 VDD.n3867 8.45089
R8132 VDD.n3856 VDD.n3855 8.45089
R8133 VDD.n3852 VDD.n3851 8.45089
R8134 VDD.n3846 VDD.n3845 8.45089
R8135 VDD.n3841 VDD.n3839 8.45089
R8136 VDD.n3826 VDD.n3825 8.45089
R8137 VDD.n3821 VDD.n3820 8.45089
R8138 VDD.n3806 VDD.n3805 8.45089
R8139 VDD.n3786 VDD.n3785 8.45089
R8140 VDD.n3780 VDD.n3779 8.45089
R8141 VDD.n3743 VDD.n3742 8.45089
R8142 VDD.n3725 VDD.n3724 8.45089
R8143 VDD.n3721 VDD.n3720 8.45089
R8144 VDD.n3717 VDD.n3716 8.45089
R8145 VDD.n3711 VDD.n3710 8.45089
R8146 VDD.n3708 VDD.n3630 8.45089
R8147 VDD VDD.n3708 8.45089
R8148 VDD.n3699 VDD.n3698 8.45089
R8149 VDD.n3690 VDD.n3689 8.45089
R8150 VDD.n3686 VDD.n3685 8.45089
R8151 VDD.n3682 VDD.n3681 8.45089
R8152 VDD.n3672 VDD.n3671 8.45089
R8153 VDD.n3668 VDD.n3667 8.45089
R8154 VDD.n3664 VDD.n3663 8.45089
R8155 VDD.n3658 VDD.n3657 8.45089
R8156 VDD.n3654 VDD.n3653 8.45089
R8157 VDD.n3650 VDD.n3649 8.45089
R8158 VDD.n1829 VDD.n1828 8.45089
R8159 VDD.n1808 VDD.n1807 8.45089
R8160 VDD.n1908 VDD.n1907 8.45089
R8161 VDD.n1921 VDD.n1920 8.45089
R8162 VDD.n1929 VDD.n1928 8.45089
R8163 VDD.n1934 VDD.n1933 8.45089
R8164 VDD.n1944 VDD.n1943 8.45089
R8165 VDD.n1952 VDD.n1951 8.45089
R8166 VDD.n1960 VDD.n1959 8.45089
R8167 VDD.n1969 VDD.n1968 8.45089
R8168 VDD.n1750 VDD.n1749 8.45089
R8169 VDD.n1746 VDD.n1745 8.45089
R8170 VDD.n1740 VDD.n1739 8.45089
R8171 VDD.n1737 VDD.n1736 8.45089
R8172 VDD VDD.n1737 8.45089
R8173 VDD.n1727 VDD.n1726 8.45089
R8174 VDD.n1713 VDD.n1712 8.45089
R8175 VDD.n1026 VDD.n1025 8.45089
R8176 VDD.n1012 VDD.n1011 8.45089
R8177 VDD.n961 VDD.n960 8.45089
R8178 VDD.n665 VDD.n663 8.45089
R8179 VDD.n654 VDD.n653 8.45089
R8180 VDD.n621 VDD.n620 8.45089
R8181 VDD.n591 VDD.n590 8.45089
R8182 VDD.n431 VDD.n430 8.45089
R8183 VDD.n427 VDD.n426 8.45089
R8184 VDD.n422 VDD.n421 8.45089
R8185 VDD.n112 VDD.n109 8.45089
R8186 VDD.n105 VDD.n104 8.45089
R8187 VDD.n99 VDD.n98 8.45089
R8188 VDD.n4861 VDD.n4860 8.45089
R8189 VDD.n4853 VDD.n4852 8.45089
R8190 VDD.n5 VDD.n4 8.45089
R8191 VDD.n121 VDD.n120 8.45089
R8192 VDD.n74 VDD.n73 8.45089
R8193 VDD.n22 VDD.n21 8.45089
R8194 VDD.n29 VDD.n28 8.45089
R8195 VDD.n51 VDD.n50 8.45089
R8196 VDD.n2818 VDD.n2815 8.45089
R8197 VDD.n2882 VDD.n2881 8.45089
R8198 VDD.n2803 VDD.n2802 8.45089
R8199 VDD.n2852 VDD.n2851 8.45089
R8200 VDD.n2847 VDD.n2844 8.45089
R8201 VDD.n2890 VDD.n2889 8.45089
R8202 VDD.n3071 VDD.n3070 8.45089
R8203 VDD.n3052 VDD.n3051 8.45089
R8204 VDD.n2946 VDD.n2945 8.45089
R8205 VDD.n2915 VDD.n2914 8.45089
R8206 VDD.n2965 VDD.n2964 8.45089
R8207 VDD.n2983 VDD.n2982 8.45089
R8208 VDD.n2990 VDD.n2989 8.45089
R8209 VDD.n3024 VDD.n3023 8.45089
R8210 VDD.n3046 VDD.n3045 8.45089
R8211 VDD.n2781 VDD.n2778 8.45089
R8212 VDD.n3111 VDD.n3107 8.45089
R8213 VDD.n3116 VDD.n3115 8.45089
R8214 VDD.n3130 VDD.n3129 8.45089
R8215 VDD.n3135 VDD.n3134 8.45089
R8216 VDD.n3156 VDD.n3155 8.45089
R8217 VDD.n3188 VDD.n3187 8.45089
R8218 VDD.n3184 VDD.n3183 8.45089
R8219 VDD.n3194 VDD.n3193 8.45089
R8220 VDD.n3126 VDD.n3125 8.45089
R8221 VDD.n2785 VDD.n2784 8.45089
R8222 VDD.n3078 VDD.n3077 8.45089
R8223 VDD.n3018 VDD.n3017 8.45089
R8224 VDD.n3013 VDD.n3012 8.45089
R8225 VDD.n2996 VDD.n2995 8.45089
R8226 VDD.n2959 VDD.n2958 8.45089
R8227 VDD.n2952 VDD.n2951 8.45089
R8228 VDD.n2886 VDD.n2885 8.45089
R8229 VDD.n2841 VDD.n2840 8.45089
R8230 VDD.n2822 VDD.n2821 8.45089
R8231 VDD.n143 VDD.n142 8.45089
R8232 VDD.n56 VDD.n55 8.45089
R8233 VDD.n44 VDD.n43 8.45089
R8234 VDD.n81 VDD.n80 8.45089
R8235 VDD.n70 VDD.n69 8.45089
R8236 VDD.n129 VDD.n128 8.45089
R8237 VDD VDD.n498 8.45089
R8238 VDD.n515 VDD.n514 8.45089
R8239 VDD.n523 VDD.n522 8.45089
R8240 VDD.n558 VDD.n557 8.45089
R8241 VDD.n574 VDD.n573 8.45089
R8242 VDD.n677 VDD.n676 8.45089
R8243 VDD.n688 VDD.n687 8.45089
R8244 VDD.n700 VDD.n699 8.45089
R8245 VDD.n714 VDD.n713 8.45089
R8246 VDD.n705 VDD.n704 8.45089
R8247 VDD.n1184 VDD.n1183 8.45089
R8248 VDD.n1176 VDD.n1175 8.45089
R8249 VDD.n1167 VDD.n1166 8.45089
R8250 VDD.n1163 VDD.n1162 8.45089
R8251 VDD.n1134 VDD.n1133 8.45089
R8252 VDD.n1124 VDD.n1123 8.45089
R8253 VDD.n1120 VDD.n1119 8.45089
R8254 VDD.n1112 VDD.n1111 8.45089
R8255 VDD.n1108 VDD.n1107 8.45089
R8256 VDD.n1098 VDD.n1097 8.45089
R8257 VDD.n1093 VDD.n1092 8.45089
R8258 VDD.n1078 VDD.n1077 8.45089
R8259 VDD.n1116 VDD.n1115 8.45089
R8260 VDD.n1159 VDD.n1158 8.45089
R8261 VDD.n1181 VDD.n1180 8.45089
R8262 VDD VDD.n1181 8.45089
R8263 VDD.n1065 VDD.n1064 8.45089
R8264 VDD.n726 VDD.n725 8.45089
R8265 VDD.n694 VDD.n693 8.45089
R8266 VDD.n570 VDD.n569 8.45089
R8267 VDD.n564 VDD.n563 8.45089
R8268 VDD.n554 VDD.n553 8.45089
R8269 VDD.n519 VDD.n518 8.45089
R8270 VDD.n1548 VDD.n1547 8.45089
R8271 VDD.n2538 VDD.n2537 8.45089
R8272 VDD.n4138 VDD.n4137 8.45089
R8273 VDD.n4123 VDD.n4122 8.45089
R8274 VDD.n2636 VDD.n2635 8.45089
R8275 VDD.n4226 VDD.n4225 8.45089
R8276 VDD.n4231 VDD.n4230 8.45089
R8277 VDD.n4235 VDD.n4234 8.45089
R8278 VDD.n4239 VDD.n4238 8.45089
R8279 VDD.n4243 VDD.n4242 8.45089
R8280 VDD.n4249 VDD.n4248 8.45089
R8281 VDD.n4253 VDD.n4252 8.45089
R8282 VDD.n4187 VDD.n4186 8.45089
R8283 VDD.n4191 VDD.n4190 8.45089
R8284 VDD.n4181 VDD.n4180 8.45089
R8285 VDD.n4282 VDD.n4281 8.45089
R8286 VDD.n4286 VDD.n4285 8.45089
R8287 VDD.n4291 VDD.n4290 8.45089
R8288 VDD.n4296 VDD.n4295 8.45089
R8289 VDD VDD.n4296 8.45089
R8290 VDD.n4299 VDD.n4298 8.45089
R8291 VDD.n4305 VDD.n4304 8.45089
R8292 VDD.n4309 VDD.n4308 8.45089
R8293 VDD.n2620 VDD.n2619 8.45089
R8294 VDD.n4331 VDD.n4330 8.45089
R8295 VDD.n4327 VDD.n4326 8.45089
R8296 VDD.n4323 VDD.n4322 8.45089
R8297 VDD.n2601 VDD.n2600 8.45089
R8298 VDD.n2605 VDD.n2604 8.45089
R8299 VDD.n4426 VDD.n4425 8.45089
R8300 VDD.n4431 VDD.n4430 8.45089
R8301 VDD.n4400 VDD.n4399 8.45089
R8302 VDD.n4405 VDD.n4404 8.45089
R8303 VDD.n4395 VDD.n4394 8.45089
R8304 VDD.n4460 VDD.n4459 8.45089
R8305 VDD.n4464 VDD.n4463 8.45089
R8306 VDD.n4469 VDD.n4468 8.45089
R8307 VDD.n4474 VDD.n4473 8.45089
R8308 VDD VDD.n4474 8.45089
R8309 VDD.n4477 VDD.n4476 8.45089
R8310 VDD.n4483 VDD.n4482 8.45089
R8311 VDD.n4487 VDD.n4486 8.45089
R8312 VDD.n4491 VDD.n4490 8.45089
R8313 VDD.n4511 VDD.n4510 8.45089
R8314 VDD.n4516 VDD.n4515 8.45089
R8315 VDD.n4520 VDD.n4519 8.45089
R8316 VDD.n4524 VDD.n4523 8.45089
R8317 VDD.n2586 VDD.n2585 8.45089
R8318 VDD.n2582 VDD.n2581 8.45089
R8319 VDD.n2578 VDD.n2577 8.45089
R8320 VDD.n4565 VDD.n4564 8.45089
R8321 VDD.n4570 VDD.n4569 8.45089
R8322 VDD.n4578 VDD.n4574 8.45089
R8323 VDD.n4605 VDD.n4604 8.45089
R8324 VDD.n4614 VDD.n4613 8.45089
R8325 VDD.n4620 VDD.n2531 8.45089
R8326 VDD VDD.n2531 8.45089
R8327 VDD.n4621 VDD.n2530 8.45089
R8328 VDD.n4627 VDD.n4624 8.45089
R8329 VDD.n4631 VDD.n4630 8.45089
R8330 VDD.n4635 VDD.n4634 8.45089
R8331 VDD.n4653 VDD.n4652 8.45089
R8332 VDD.n4658 VDD.n4657 8.45089
R8333 VDD.n4662 VDD.n4661 8.45089
R8334 VDD.n4666 VDD.n4665 8.45089
R8335 VDD.n4676 VDD.n4675 8.45089
R8336 VDD.n4680 VDD.n4679 8.45089
R8337 VDD.n4684 VDD.n4683 8.45089
R8338 VDD.n4688 VDD.n4687 8.45089
R8339 VDD.n4694 VDD.n4692 8.45089
R8340 VDD.n2508 VDD.n2505 8.45089
R8341 VDD.n2512 VDD.n2511 8.45089
R8342 VDD.n2362 VDD.n2361 8.45089
R8343 VDD.n2358 VDD.n2357 8.45089
R8344 VDD.n2349 VDD.n2348 8.45089
R8345 VDD.n2341 VDD.n2340 8.45089
R8346 VDD VDD.n2341 8.45089
R8347 VDD.n2011 VDD.n2010 8.45089
R8348 VDD.n2017 VDD.n2016 8.45089
R8349 VDD.n2021 VDD.n2020 8.45089
R8350 VDD.n2025 VDD.n2024 8.45089
R8351 VDD.n2058 VDD.n2057 8.45089
R8352 VDD.n2062 VDD.n2061 8.45089
R8353 VDD.n2066 VDD.n2065 8.45089
R8354 VDD.n2071 VDD.n2070 8.45089
R8355 VDD.n2075 VDD.n2074 8.45089
R8356 VDD.n2079 VDD.n2078 8.45089
R8357 VDD.n2083 VDD.n2082 8.45089
R8358 VDD.n2087 VDD.n2086 8.45089
R8359 VDD.n2093 VDD.n2092 8.45089
R8360 VDD.n2097 VDD.n2096 8.45089
R8361 VDD.n2122 VDD.n2121 8.45089
R8362 VDD.n2127 VDD.n2126 8.45089
R8363 VDD.n2002 VDD.n2001 8.45089
R8364 VDD.n1602 VDD.n1601 8.45089
R8365 VDD.n1592 VDD.n1591 8.45089
R8366 VDD VDD.n1592 8.45089
R8367 VDD.n1580 VDD.n1579 8.45089
R8368 VDD.n1577 VDD.n1576 8.45089
R8369 VDD.n1571 VDD.n1570 8.45089
R8370 VDD.n1566 VDD.n1565 8.45089
R8371 VDD.n1562 VDD.n1561 8.45089
R8372 VDD.n4555 VDD.n4554 8.45089
R8373 VDD.n4777 VDD.n4776 8.45089
R8374 VDD.n4781 VDD.n4780 8.45089
R8375 VDD.n4789 VDD.n4788 8.45089
R8376 VDD.n4804 VDD.n4803 8.45089
R8377 VDD.n4794 VDD.n4793 8.45089
R8378 VDD.n4825 VDD.n4824 8.45089
R8379 VDD.n3411 VDD.n3410 8.45089
R8380 VDD.n3450 VDD.n3449 8.45089
R8381 VDD.n3446 VDD.n3445 8.45089
R8382 VDD.n3437 VDD.n3436 8.45089
R8383 VDD.n3433 VDD.n3432 8.45089
R8384 VDD.n3429 VDD.n3428 8.45089
R8385 VDD.n3425 VDD.n3424 8.45089
R8386 VDD.n3421 VDD.n3420 8.45089
R8387 VDD.n2695 VDD.n2694 8.45089
R8388 VDD.n3378 VDD.n3377 8.45089
R8389 VDD.n3382 VDD.n3381 8.45089
R8390 VDD.n3386 VDD.n3385 8.45089
R8391 VDD.n3392 VDD.n3390 8.45089
R8392 VDD.n2731 VDD.n2730 8.45089
R8393 VDD.n2709 VDD.n2708 8.45089
R8394 VDD.n2755 VDD.n2754 8.45089
R8395 VDD.n3287 VDD.n3286 8.45089
R8396 VDD.n3295 VDD.n3294 8.45089
R8397 VDD.n3307 VDD.n3306 8.45089
R8398 VDD.n3221 VDD.n3220 8.45089
R8399 VDD.n3218 VDD.n3217 8.45089
R8400 VDD.n3301 VDD.n3300 8.45089
R8401 VDD.n3291 VDD.n3290 8.45089
R8402 VDD.n3279 VDD.n3278 8.45089
R8403 VDD.n2713 VDD.n2712 8.45089
R8404 VDD.n3417 VDD.n3416 8.45089
R8405 VDD.n4819 VDD.n4818 8.45089
R8406 VDD.n4798 VDD.n4797 8.45089
R8407 VDD.n4785 VDD.n4784 8.45089
R8408 VDD.n3607 VDD.n3606 8.44032
R8409 VDD.n3373 VDD.n3370 8.38671
R8410 VDD.n3356 VDD.n3355 8.38671
R8411 VDD.n3351 VDD.n3350 8.38671
R8412 VDD.n3346 VDD.n3345 8.38671
R8413 VDD.n3341 VDD.n3338 8.38671
R8414 VDD.n3334 VDD.n3333 8.38671
R8415 VDD.n3329 VDD.n3322 8.38671
R8416 VDD.n3453 VDD.n3403 8.38671
R8417 VDD.n3463 VDD.n3462 8.38671
R8418 VDD.n3468 VDD.n3467 8.38671
R8419 VDD.n3473 VDD.n3472 8.38671
R8420 VDD.n3478 VDD.n3477 8.38671
R8421 VDD.n3483 VDD.n3482 8.38671
R8422 VDD.n3490 VDD.n3489 8.38671
R8423 VDD.n3507 VDD.n3494 8.38671
R8424 VDD.n2289 VDD.n2288 8.38671
R8425 VDD.n4767 VDD.n4766 8.38671
R8426 VDD.n3361 VDD.n2737 7.94533
R8427 VDD.n3457 VDD.n3456 7.94533
R8428 VDD.n2705 VDD.n2704 7.94533
R8429 VDD.n861 VDD.t34 7.83017
R8430 VDD.n1642 VDD.t497 7.83017
R8431 VDD.n2207 VDD.t170 7.83017
R8432 VDD.n2429 VDD.t78 7.83017
R8433 VDD.n267 VDD.n266 7.05932
R8434 VDD.n265 VDD.n264 7.05932
R8435 VDD.n1250 VDD.n1249 7.05932
R8436 VDD.n1264 VDD.n1263 7.05932
R8437 VDD.n1278 VDD.n1277 7.05932
R8438 VDD.n1292 VDD.n1291 7.05932
R8439 VDD.n1308 VDD.n1307 7.05932
R8440 VDD.n1322 VDD.n1321 7.05932
R8441 VDD.n1339 VDD.n1338 7.05932
R8442 VDD.n534 VDD.n531 6.80365
R8443 VDD.n1141 VDD.n1138 6.80365
R8444 VDD.n2104 VDD.n2101 6.80365
R8445 VDD.n2492 VDD.n2489 6.80365
R8446 VDD.n2554 VDD.n2551 6.80365
R8447 VDD.n4438 VDD.n4435 6.80365
R8448 VDD.n4260 VDD.n4257 6.80365
R8449 VDD.n2295 VDD.n2294 6.62119
R8450 VDD.n4861 VDD.n4858 6.62119
R8451 VDD.n112 VDD.n111 6.62119
R8452 VDD.n2952 VDD.n2949 6.62119
R8453 VDD.n2983 VDD.n2980 6.62119
R8454 VDD.n3068 VDD.n3067 6.62119
R8455 VDD.n2187 VDD.n2186 6.17981
R8456 VDD.n2440 VDD.n2439 6.17981
R8457 VDD.n33 VDD.n32 5.73843
R8458 VDD.n51 VDD.n48 5.73843
R8459 VDD.n2781 VDD.n2780 5.73843
R8460 VDD.n603 VDD.t581 5.27828
R8461 VDD.n1028 VDD.t317 5.27828
R8462 VDD.n1936 VDD.t318 5.27828
R8463 VDD.n3666 VDD.t704 5.27828
R8464 VDD.n3854 VDD.t735 5.27828
R8465 VDD.n3545 VDD.t512 5.27828
R8466 VDD.n4074 VDD.t82 5.27828
R8467 VDD.n546 VDD.t600 5.26366
R8468 VDD.n1132 VDD.t744 5.26366
R8469 VDD.n2095 VDD.t248 5.26366
R8470 VDD.n2510 VDD.t668 5.26366
R8471 VDD.n4553 VDD.t458 5.26366
R8472 VDD.n4429 VDD.t243 5.26366
R8473 VDD.n4251 VDD.t400 5.26366
R8474 VDD.n380 VDD.t281 5.22028
R8475 VDD.n1236 VDD.n1235 5.22028
R8476 VDD.n1238 VDD.n1237 5.22028
R8477 VDD.n1252 VDD.n1251 5.22028
R8478 VDD.n1266 VDD.n1265 5.22028
R8479 VDD.n1280 VDD.n1279 5.22028
R8480 VDD.n1294 VDD.n1293 5.22028
R8481 VDD.n1310 VDD.n1309 5.22028
R8482 VDD.n1324 VDD.n1323 5.22028
R8483 VDD.n1341 VDD.n1340 5.22028
R8484 VDD.n4817 VDD.t56 5.22028
R8485 VDD.n3415 VDD.t390 5.22028
R8486 VDD.n2699 VDD.t396 5.22028
R8487 VDD.n3277 VDD.t375 5.22028
R8488 VDD.n3608 VDD.n3607 4.7844
R8489 VDD.n4 VDD.n3 4.69636
R8490 VDD.n2914 VDD.n2913 4.69636
R8491 VDD.n1803 VDD.n1802 4.6505
R8492 VDD.n1824 VDD.n1823 4.6505
R8493 VDD.n4017 VDD.n4016 4.6505
R8494 VDD.n4024 VDD.n4023 4.6505
R8495 VDD.n4077 VDD.n4076 4.6505
R8496 VDD.n2654 VDD.n2653 4.6505
R8497 VDD.n3548 VDD.n3547 4.6505
R8498 VDD.n3730 VDD.n3729 4.6505
R8499 VDD.n3737 VDD.n3736 4.6505
R8500 VDD.n3744 VDD.n3743 4.6505
R8501 VDD.n3787 VDD.n3786 4.6505
R8502 VDD.n3870 VDD.n3869 4.6505
R8503 VDD.n3929 VDD.n3928 4.6505
R8504 VDD.n3936 VDD.n3935 4.6505
R8505 VDD.n3962 VDD.n3961 4.6505
R8506 VDD.n3572 VDD.n3571 4.6505
R8507 VDD.n3636 VDD.n3635 4.6505
R8508 VDD.n1809 VDD.n1808 4.6505
R8509 VDD.n1778 VDD.n1777 4.6505
R8510 VDD.n1758 VDD.n1757 4.6505
R8511 VDD.n981 VDD.n980 4.6505
R8512 VDD.n974 VDD.n973 4.6505
R8513 VDD.n666 VDD.n665 4.6505
R8514 VDD.n600 VDD.n599 4.6505
R8515 VDD.n440 VDD.n439 4.6505
R8516 VDD.n447 VDD.n446 4.6505
R8517 VDD.n481 VDD.n480 4.6505
R8518 VDD.n3166 VDD.n3164 4.6505
R8519 VDD.n30 VDD.n29 4.6505
R8520 VDD.n2966 VDD.n2965 4.6505
R8521 VDD.n3025 VDD.n3024 4.6505
R8522 VDD.n3047 VDD.n3046 4.6505
R8523 VDD.n3136 VDD.n3135 4.6505
R8524 VDD.n3157 VDD.n3156 4.6505
R8525 VDD.n3125 VDD.n3124 4.6505
R8526 VDD.n3112 VDD.n3111 4.6505
R8527 VDD.n2997 VDD.n2996 4.6505
R8528 VDD.n2916 VDD.n2915 4.6505
R8529 VDD.n3072 VDD.n3071 4.6505
R8530 VDD.n2840 VDD.n2839 4.6505
R8531 VDD.n2853 VDD.n2852 4.6505
R8532 VDD.n2804 VDD.n2803 4.6505
R8533 VDD.n144 VDD.n143 4.6505
R8534 VDD.n82 VDD.n81 4.6505
R8535 VDD.n130 VDD.n129 4.6505
R8536 VDD.n4854 VDD.n4853 4.6505
R8537 VDD.n728 VDD.n727 4.6505
R8538 VDD.n1185 VDD.n1184 4.6505
R8539 VDD.n1094 VDD.n1093 4.6505
R8540 VDD.n1151 VDD.n1150 4.6505
R8541 VDD.n1156 VDD.n1155 4.6505
R8542 VDD.n715 VDD.n714 4.6505
R8543 VDD.n565 VDD.n564 4.6505
R8544 VDD.n544 VDD.n543 4.6505
R8545 VDD.n528 VDD.n527 4.6505
R8546 VDD.n4360 VDD.n4359 4.6505
R8547 VDD.n1591 VDD.n1590 4.6505
R8548 VDD.n1603 VDD.n1602 4.6505
R8549 VDD.n2119 VDD.n2118 4.6505
R8550 VDD.n2114 VDD.n2113 4.6505
R8551 VDD.n2041 VDD.n2040 4.6505
R8552 VDD.n2340 VDD.n2339 4.6505
R8553 VDD.n2486 VDD.n2485 4.6505
R8554 VDD.n2502 VDD.n2501 4.6505
R8555 VDD.n4601 VDD.n4600 4.6505
R8556 VDD.n4579 VDD.n4578 4.6505
R8557 VDD.n4566 VDD.n4565 4.6505
R8558 VDD.n4507 VDD.n4506 4.6505
R8559 VDD.n4453 VDD.n4452 4.6505
R8560 VDD.n4448 VDD.n4447 4.6505
R8561 VDD.n4379 VDD.n4378 4.6505
R8562 VDD.n2621 VDD.n2620 4.6505
R8563 VDD.n4275 VDD.n4274 4.6505
R8564 VDD.n4270 VDD.n4269 4.6505
R8565 VDD.n4227 VDD.n4226 4.6505
R8566 VDD.n4155 VDD.n4154 4.6505
R8567 VDD.n4139 VDD.n4138 4.6505
R8568 VDD.n2564 VDD.n2563 4.6505
R8569 VDD.n4805 VDD.n4804 4.6505
R8570 VDD.n4826 VDD.n4825 4.6505
R8571 VDD.n2702 VDD.n2701 4.6505
R8572 VDD.n3302 VDD.n3301 4.6505
R8573 VDD.n3393 VDD.n3392 4.6505
R8574 VDD.n3370 VDD.n3369 4.6505
R8575 VDD.n3368 VDD.n3367 4.6505
R8576 VDD.n3359 VDD.n3358 4.6505
R8577 VDD.n3357 VDD.n3356 4.6505
R8578 VDD.n3352 VDD.n3351 4.6505
R8579 VDD.n3347 VDD.n3346 4.6505
R8580 VDD.n3342 VDD.n3341 4.6505
R8581 VDD.n3335 VDD.n3334 4.6505
R8582 VDD.n3330 VDD.n3329 4.6505
R8583 VDD.n3453 VDD.n3452 4.6505
R8584 VDD.n3455 VDD.n3400 4.6505
R8585 VDD.n3464 VDD.n3463 4.6505
R8586 VDD.n3469 VDD.n3468 4.6505
R8587 VDD.n3474 VDD.n3473 4.6505
R8588 VDD.n3479 VDD.n3478 4.6505
R8589 VDD.n3484 VDD.n3483 4.6505
R8590 VDD.n3491 VDD.n3490 4.6505
R8591 VDD.n3508 VDD.n3507 4.6505
R8592 VDD.n4774 VDD.n4773 4.6505
R8593 VDD.n4765 VDD.n4760 4.6505
R8594 VDD.n4759 VDD.n4758 4.6505
R8595 VDD.n4754 VDD.n4753 4.6505
R8596 VDD.n4749 VDD.n4748 4.6505
R8597 VDD.n4744 VDD.n4743 4.6505
R8598 VDD.n4739 VDD.n4738 4.6505
R8599 VDD.n4734 VDD.n4733 4.6505
R8600 VDD.n4727 VDD.n4726 4.6505
R8601 VDD.n2419 VDD.n2418 4.6505
R8602 VDD.n2433 VDD.n2432 4.6505
R8603 VDD.n2394 VDD.n2393 4.6505
R8604 VDD.n1647 VDD.n1646 4.6505
R8605 VDD.n1661 VDD.n1660 4.6505
R8606 VDD.n1676 VDD.n1675 4.6505
R8607 VDD.n1504 VDD.n1503 4.6505
R8608 VDD.n1484 VDD.n1483 4.6505
R8609 VDD.n1463 VDD.n1462 4.6505
R8610 VDD.n2167 VDD.n2166 4.6505
R8611 VDD.n2181 VDD.n2180 4.6505
R8612 VDD.n2197 VDD.n2196 4.6505
R8613 VDD.n2211 VDD.n2210 4.6505
R8614 VDD.n2234 VDD.n2233 4.6505
R8615 VDD.n2252 VDD.n2251 4.6505
R8616 VDD.n2257 VDD.n2256 4.6505
R8617 VDD.n2264 VDD.n2263 4.6505
R8618 VDD.n2269 VDD.n2268 4.6505
R8619 VDD.n2274 VDD.n2273 4.6505
R8620 VDD.n2279 VDD.n2278 4.6505
R8621 VDD.n2284 VDD.n2283 4.6505
R8622 VDD.n2287 VDD.n2286 4.6505
R8623 VDD.n2304 VDD.n2303 4.6505
R8624 VDD.n203 VDD.n202 4.6505
R8625 VDD.n1860 VDD.n1859 4.6505
R8626 VDD.n1410 VDD.n1409 4.6505
R8627 VDD.n1375 VDD.n1374 4.6505
R8628 VDD.n1346 VDD.n1345 4.6505
R8629 VDD.n1329 VDD.n1328 4.6505
R8630 VDD.n1315 VDD.n1314 4.6505
R8631 VDD.n1299 VDD.n1298 4.6505
R8632 VDD.n1285 VDD.n1284 4.6505
R8633 VDD.n1271 VDD.n1270 4.6505
R8634 VDD.n1257 VDD.n1256 4.6505
R8635 VDD.n1243 VDD.n1242 4.6505
R8636 VDD.n1229 VDD.n1228 4.6505
R8637 VDD.n1203 VDD.n1202 4.6505
R8638 VDD.n895 VDD.n894 4.6505
R8639 VDD.n880 VDD.n879 4.6505
R8640 VDD.n866 VDD.n865 4.6505
R8641 VDD.n852 VDD.n851 4.6505
R8642 VDD.n835 VDD.n834 4.6505
R8643 VDD.n821 VDD.n820 4.6505
R8644 VDD.n328 VDD.n327 4.6505
R8645 VDD.n342 VDD.n341 4.6505
R8646 VDD.n356 VDD.n355 4.6505
R8647 VDD.n370 VDD.n369 4.6505
R8648 VDD.n384 VDD.n383 4.6505
R8649 VDD.n398 VDD.n397 4.6505
R8650 VDD.n412 VDD.n411 4.6505
R8651 VDD.n782 VDD.n781 4.6505
R8652 VDD.n533 VDD.n530 4.53646
R8653 VDD.n1140 VDD.n1137 4.53646
R8654 VDD.n2103 VDD.n2100 4.53646
R8655 VDD.n2491 VDD.n2488 4.53646
R8656 VDD.n2553 VDD.n2550 4.53646
R8657 VDD.n4437 VDD.n4434 4.53646
R8658 VDD.n4259 VDD.n4256 4.53646
R8659 VDD.n1811 VDD.n1810 4.5005
R8660 VDD.n1990 VDD.n1989 4.5005
R8661 VDD.n1760 VDD.n1759 4.5005
R8662 VDD.n1045 VDD.n1044 4.5005
R8663 VDD.n632 VDD.n631 4.5005
R8664 VDD.n602 VDD.n601 4.5005
R8665 VDD.n483 VDD.n482 4.5005
R8666 VDD.n668 VDD.n667 4.5005
R8667 VDD.n296 VDD.n295 4.5005
R8668 VDD.n3638 VDD.n3637 4.5005
R8669 VDD.n3574 VDD.n3573 4.5005
R8670 VDD.n3964 VDD.n3963 4.5005
R8671 VDD.n3865 VDD.n3864 4.5005
R8672 VDD.n3837 VDD.n3836 4.5005
R8673 VDD.n3817 VDD.n3816 4.5005
R8674 VDD.n3789 VDD.n3788 4.5005
R8675 VDD.n3747 VDD.n3746 4.5005
R8676 VDD.n3550 VDD.n3549 4.5005
R8677 VDD.n2656 VDD.n2655 4.5005
R8678 VDD.n4079 VDD.n4078 4.5005
R8679 VDD.n2678 VDD.n2677 4.5005
R8680 VDD.n3602 VDD.n3601 4.5005
R8681 VDD.n3246 VDD.n3245 4.5005
R8682 VDD.n3159 VDD.n3158 4.5005
R8683 VDD.n3138 VDD.n3137 4.5005
R8684 VDD.n2968 VDD.n2967 4.5005
R8685 VDD.n2933 VDD.n2932 4.5005
R8686 VDD.n146 VDD.n145 4.5005
R8687 VDD.n4856 VDD.n4855 4.5005
R8688 VDD.n86 VDD.n85 4.5005
R8689 VDD.n132 VDD.n131 4.5005
R8690 VDD.n2837 VDD.n2836 4.5005
R8691 VDD.n2855 VDD.n2854 4.5005
R8692 VDD.n2806 VDD.n2805 4.5005
R8693 VDD.n2910 VDD.n2909 4.5005
R8694 VDD.n2999 VDD.n2998 4.5005
R8695 VDD.n3049 VDD.n3048 4.5005
R8696 VDD.n3105 VDD.n3104 4.5005
R8697 VDD.n3074 VDD.n3073 4.5005
R8698 VDD.n3122 VDD.n3121 4.5005
R8699 VDD.n34 VDD.n33 4.5005
R8700 VDD.n3168 VDD.n3167 4.5005
R8701 VDD.n3029 VDD.n3028 4.5005
R8702 VDD.n1187 VDD.n1186 4.5005
R8703 VDD.n710 VDD.n709 4.5005
R8704 VDD.n567 VDD.n566 4.5005
R8705 VDD.n1089 VDD.n1088 4.5005
R8706 VDD.n1551 VDD.n1550 4.5005
R8707 VDD.n4194 VDD.n4193 4.5005
R8708 VDD.n4363 VDD.n4362 4.5005
R8709 VDD.n4342 VDD.n4341 4.5005
R8710 VDD.n4534 VDD.n4533 4.5005
R8711 VDD.n4581 VDD.n4580 4.5005
R8712 VDD.n4596 VDD.n4595 4.5005
R8713 VDD.n2337 VDD.n2336 4.5005
R8714 VDD.n4134 VDD.n4133 4.5005
R8715 VDD.n1588 VDD.n1587 4.5005
R8716 VDD.n1605 VDD.n1604 4.5005
R8717 VDD.n2371 VDD.n2370 4.5005
R8718 VDD.n4697 VDD.n4696 4.5005
R8719 VDD.n4561 VDD.n4560 4.5005
R8720 VDD.n4222 VDD.n4221 4.5005
R8721 VDD.n2623 VDD.n2622 4.5005
R8722 VDD.n4828 VDD.n4827 4.5005
R8723 VDD.n4807 VDD.n4806 4.5005
R8724 VDD.n2320 VDD.n2319 4.5005
R8725 VDD.n1222 VDD.n1221 4.5005
R8726 VDD.n914 VDD.n913 4.5005
R8727 VDD.n1396 VDD.n1395 4.5005
R8728 VDD.n1694 VDD.n1693 4.5005
R8729 VDD.n1520 VDD.n1519 4.5005
R8730 VDD.n1474 VDD.n1473 4.5005
R8731 VDD.n239 VDD.n238 4.5005
R8732 VDD.n2298 VDD.n2297 4.5005
R8733 VDD.n3395 VDD.n3394 4.5005
R8734 VDD.n3225 VDD.n3224 4.5005
R8735 VDD.n3304 VDD.n3303 4.5005
R8736 VDD.n2706 VDD.n2705 4.5005
R8737 VDD.n1879 VDD.n1878 4.5005
R8738 VDD.n841 VDD.n840 3.97291
R8739 VDD.n317 VDD 3.89041
R8740 VDD.n4129 VDD.n4125 3.78744
R8741 VDD.n317 VDD.n316 3.53153
R8742 VDD.n327 VDD.n326 3.53153
R8743 VDD.n326 VDD.n310 3.53153
R8744 VDD.n341 VDD.n340 3.53153
R8745 VDD.n340 VDD.n333 3.53153
R8746 VDD.n355 VDD.n354 3.53153
R8747 VDD.n354 VDD.n347 3.53153
R8748 VDD.n369 VDD.n368 3.53153
R8749 VDD.n368 VDD.n361 3.53153
R8750 VDD.n383 VDD.n382 3.53153
R8751 VDD.n382 VDD.n375 3.53153
R8752 VDD.n397 VDD.n396 3.53153
R8753 VDD.n396 VDD.n389 3.53153
R8754 VDD.n411 VDD.n410 3.53153
R8755 VDD.n789 VDD.n782 3.53153
R8756 VDD.n790 VDD.n789 3.53153
R8757 VDD.n1483 VDD.n1432 3.53153
R8758 VDD.n1441 VDD.n1433 3.53153
R8759 VDD.n1474 VDD.n1446 3.53153
R8760 VDD.n1462 VDD.n1452 3.53153
R8761 VDD.n1454 VDD.n1453 3.53153
R8762 VDD.n2166 VDD.n2156 3.53153
R8763 VDD.n2158 VDD.n2157 3.53153
R8764 VDD.n2180 VDD.n2170 3.53153
R8765 VDD.n2172 VDD.n2171 3.53153
R8766 VDD.n2196 VDD.n2184 3.53153
R8767 VDD.n2188 VDD.n2187 3.53153
R8768 VDD.n2210 VDD.n2200 3.53153
R8769 VDD.n2202 VDD.n2201 3.53153
R8770 VDD.n2233 VDD.n2214 3.53153
R8771 VDD.n2225 VDD.n2224 3.53153
R8772 VDD.n2304 VDD.n216 3.53153
R8773 VDD.n2306 VDD.n2305 3.53153
R8774 VDD.n211 VDD.n210 3.53153
R8775 VDD.n202 VDD.n192 3.53153
R8776 VDD.n194 VDD.n193 3.53153
R8777 VDD.n1859 VDD.n1849 3.53153
R8778 VDD.n1851 VDD.n1850 3.53153
R8779 VDD.n2393 VDD.n2383 3.53153
R8780 VDD.n2385 VDD.n2384 3.53153
R8781 VDD.n2450 VDD.n2437 3.53153
R8782 VDD.n2432 VDD.n2422 3.53153
R8783 VDD.n2424 VDD.n2423 3.53153
R8784 VDD.n2418 VDD.n2399 3.53153
R8785 VDD.n2410 VDD.n2409 3.53153
R8786 VDD.n3188 VDD 3.53153
R8787 VDD.n4226 VDD.n4223 3.53153
R8788 VDD.n4600 VDD.n4597 3.53153
R8789 VDD.n1481 VDD.n1435 3.52991
R8790 VDD.n1476 VDD.n1439 3.52991
R8791 VDD.n1460 VDD.n1456 3.52991
R8792 VDD.n234 VDD.n230 3.52991
R8793 VDD.n2164 VDD.n2160 3.52991
R8794 VDD.n2178 VDD.n2174 3.52991
R8795 VDD.n2194 VDD.n2190 3.52991
R8796 VDD.n2208 VDD.n2204 3.52991
R8797 VDD.n2231 VDD.n2227 3.52991
R8798 VDD.n2308 VDD.n215 3.52991
R8799 VDD.n2315 VDD.n213 3.52991
R8800 VDD.n200 VDD.n196 3.52991
R8801 VDD.n1857 VDD.n1853 3.52991
R8802 VDD.n1875 VDD.n1871 3.52991
R8803 VDD.n2391 VDD.n2387 3.52991
R8804 VDD.n2448 VDD.n2444 3.52991
R8805 VDD.n2430 VDD.n2426 3.52991
R8806 VDD.n2416 VDD.n2412 3.52991
R8807 VDD.n319 VDD.n318 3.52991
R8808 VDD.n312 VDD.n311 3.52991
R8809 VDD.n335 VDD.n334 3.52991
R8810 VDD.n349 VDD.n348 3.52991
R8811 VDD.n363 VDD.n362 3.52991
R8812 VDD.n377 VDD.n376 3.52991
R8813 VDD.n391 VDD.n390 3.52991
R8814 VDD.n405 VDD.n404 3.52991
R8815 VDD.n784 VDD.n783 3.52991
R8816 VDD.n2052 VDD.n2048 3.52991
R8817 VDD.n2038 VDD.n2034 3.52991
R8818 VDD.n4647 VDD.n4643 3.52991
R8819 VDD.n4504 VDD.n4500 3.52991
R8820 VDD.n4358 VDD.n4354 3.52991
R8821 VDD.n4375 VDD.n4371 3.52991
R8822 VDD.n740 VDD.n736 3.52991
R8823 VDD.n4152 VDD.n4148 3.42907
R8824 VDD.n1232 VDD.n1229 3.31084
R8825 VDD.n1232 VDD.n1231 3.31084
R8826 VDD.n1242 VDD.n1241 3.31084
R8827 VDD.n1241 VDD.n263 3.31084
R8828 VDD.n1256 VDD.n1255 3.31084
R8829 VDD.n1255 VDD.n1248 3.31084
R8830 VDD.n1270 VDD.n1269 3.31084
R8831 VDD.n1269 VDD.n1262 3.31084
R8832 VDD.n1284 VDD.n1283 3.31084
R8833 VDD.n1283 VDD.n1276 3.31084
R8834 VDD.n1298 VDD.n1297 3.31084
R8835 VDD.n1297 VDD.n1290 3.31084
R8836 VDD.n1314 VDD.n1313 3.31084
R8837 VDD.n1313 VDD.n1306 3.31084
R8838 VDD.n1328 VDD.n1327 3.31084
R8839 VDD.n1327 VDD.n1320 3.31084
R8840 VDD.n1345 VDD.n1344 3.31084
R8841 VDD.n1344 VDD.n1337 3.31084
R8842 VDD.n2442 VDD.n2441 3.31084
R8843 VDD.n665 VDD.n664 3.31084
R8844 VDD.n2653 VDD.n2650 3.31084
R8845 VDD.n3635 VDD.n3632 3.31084
R8846 VDD.n2846 VDD.n2845 3.31084
R8847 VDD.n2840 VDD.n2813 3.31084
R8848 VDD.n2996 VDD.n2993 3.31084
R8849 VDD.n3125 VDD.n2776 3.31084
R8850 VDD.n4192 VDD.n4191 3.27033
R8851 VDD.n428 VDD.n422 3.22029
R8852 VDD.n497 VDD 3.12264
R8853 VDD.n537 VDD 3.10353
R8854 VDD.n1144 VDD 3.10353
R8855 VDD.n2107 VDD 3.10353
R8856 VDD.n2495 VDD 3.10353
R8857 VDD.n2557 VDD 3.10353
R8858 VDD.n4441 VDD 3.10353
R8859 VDD.n4263 VDD 3.10353
R8860 VDD.n1979 VDD.n1978 3.1005
R8861 VDD.n487 VDD.n486 3.1005
R8862 VDD.n606 VDD.n605 3.1005
R8863 VDD.n987 VDD.n986 3.1005
R8864 VDD.n1035 VDD.n1034 3.1005
R8865 VDD.n248 VDD.n247 3.1005
R8866 VDD.n1974 VDD.n1973 3.1005
R8867 VDD.n1965 VDD.n1964 3.1005
R8868 VDD.n1957 VDD.n1956 3.1005
R8869 VDD.n1949 VDD.n1948 3.1005
R8870 VDD.n1939 VDD.n1938 3.1005
R8871 VDD.n1926 VDD.n1925 3.1005
R8872 VDD.n1917 VDD.n1916 3.1005
R8873 VDD.n1912 VDD.n1911 3.1005
R8874 VDD.n1905 VDD.n1904 3.1005
R8875 VDD.n1899 VDD.n1898 3.1005
R8876 VDD.n3647 VDD.n3646 3.1005
R8877 VDD.n3994 VDD.n3993 3.1005
R8878 VDD.n4005 VDD.n4004 3.1005
R8879 VDD.n4009 VDD.n4008 3.1005
R8880 VDD.n4030 VDD.n4029 3.1005
R8881 VDD.n4038 VDD.n4037 3.1005
R8882 VDD.n4048 VDD.n4047 3.1005
R8883 VDD.n4056 VDD.n4055 3.1005
R8884 VDD.n4064 VDD.n4063 3.1005
R8885 VDD.n3259 VDD.n3258 3.1005
R8886 VDD.n3254 VDD.n3253 3.1005
R8887 VDD.n2660 VDD.n2659 3.1005
R8888 VDD.n4102 VDD.n4101 3.1005
R8889 VDD.n4091 VDD.n4090 3.1005
R8890 VDD.n4070 VDD.n4069 3.1005
R8891 VDD.n4060 VDD.n4059 3.1005
R8892 VDD.n4052 VDD.n4051 3.1005
R8893 VDD.n4034 VDD.n4033 3.1005
R8894 VDD.n4013 VDD.n4012 3.1005
R8895 VDD.n3999 VDD.n3998 3.1005
R8896 VDD.n3986 VDD.n3985 3.1005
R8897 VDD.n3622 VDD.n3621 3.1005
R8898 VDD.n3613 VDD.n3612 3.1005
R8899 VDD.n3542 VDD.n3541 3.1005
R8900 VDD.n3655 VDD.n3654 3.1005
R8901 VDD.n3659 VDD.n3658 3.1005
R8902 VDD.n3665 VDD.n3664 3.1005
R8903 VDD.n3669 VDD.n3668 3.1005
R8904 VDD.n3673 VDD.n3672 3.1005
R8905 VDD.n3683 VDD.n3682 3.1005
R8906 VDD.n3687 VDD.n3686 3.1005
R8907 VDD.n3691 VDD.n3690 3.1005
R8908 VDD.n3700 VDD.n3699 3.1005
R8909 VDD.n3701 VDD.n3630 3.1005
R8910 VDD.n3712 VDD.n3711 3.1005
R8911 VDD.n3718 VDD.n3717 3.1005
R8912 VDD.n3722 VDD.n3721 3.1005
R8913 VDD.n3726 VDD.n3725 3.1005
R8914 VDD.n3781 VDD.n3780 3.1005
R8915 VDD.n3807 VDD.n3806 3.1005
R8916 VDD.n3822 VDD.n3821 3.1005
R8917 VDD.n3827 VDD.n3826 3.1005
R8918 VDD.n3842 VDD.n3841 3.1005
R8919 VDD.n3847 VDD.n3846 3.1005
R8920 VDD.n3853 VDD.n3852 3.1005
R8921 VDD.n3857 VDD.n3856 3.1005
R8922 VDD.n3881 VDD.n3880 3.1005
R8923 VDD.n3885 VDD.n3884 3.1005
R8924 VDD.n3889 VDD.n3888 3.1005
R8925 VDD.n3898 VDD.n3897 3.1005
R8926 VDD.n3906 VDD.n3905 3.1005
R8927 VDD.n3911 VDD.n3910 3.1005
R8928 VDD.n3917 VDD.n3916 3.1005
R8929 VDD.n3921 VDD.n3920 3.1005
R8930 VDD.n3925 VDD.n3924 3.1005
R8931 VDD.n3942 VDD.n3941 3.1005
R8932 VDD.n3946 VDD.n3945 3.1005
R8933 VDD.n3950 VDD.n3949 3.1005
R8934 VDD.n3968 VDD.n3967 3.1005
R8935 VDD.n3561 VDD.n3560 3.1005
R8936 VDD.n3566 VDD.n3565 3.1005
R8937 VDD.n3535 VDD.n3534 3.1005
R8938 VDD.n3651 VDD.n3650 3.1005
R8939 VDD.n1830 VDD.n1829 3.1005
R8940 VDD.n1907 VDD.n1906 3.1005
R8941 VDD.n1922 VDD.n1921 3.1005
R8942 VDD.n1930 VDD.n1929 3.1005
R8943 VDD.n1935 VDD.n1934 3.1005
R8944 VDD.n1945 VDD.n1944 3.1005
R8945 VDD.n1953 VDD.n1952 3.1005
R8946 VDD.n1961 VDD.n1960 3.1005
R8947 VDD.n1970 VDD.n1969 3.1005
R8948 VDD.n1728 VDD.n1727 3.1005
R8949 VDD.n1736 VDD.n1735 3.1005
R8950 VDD.n1741 VDD.n1740 3.1005
R8951 VDD.n1747 VDD.n1746 3.1005
R8952 VDD.n1751 VDD.n1750 3.1005
R8953 VDD.n1718 VDD.n1717 3.1005
R8954 VDD.n1031 VDD.n1030 3.1005
R8955 VDD.n1021 VDD.n1020 3.1005
R8956 VDD.n1027 VDD.n1026 3.1005
R8957 VDD.n1017 VDD.n1016 3.1005
R8958 VDD.n1009 VDD.n1008 3.1005
R8959 VDD.n1013 VDD.n1012 3.1005
R8960 VDD.n1005 VDD.n1004 3.1005
R8961 VDD.n995 VDD.n994 3.1005
R8962 VDD.n991 VDD.n990 3.1005
R8963 VDD.n970 VDD.n969 3.1005
R8964 VDD.n966 VDD.n965 3.1005
R8965 VDD.n956 VDD.n955 3.1005
R8966 VDD.n962 VDD.n961 3.1005
R8967 VDD.n951 VDD.n950 3.1005
R8968 VDD.n660 VDD.n659 3.1005
R8969 VDD.n943 VDD.n942 3.1005
R8970 VDD.n655 VDD.n654 3.1005
R8971 VDD.n622 VDD.n621 3.1005
R8972 VDD.n592 VDD.n591 3.1005
R8973 VDD.n428 VDD.n427 3.1005
R8974 VDD.n432 VDD.n431 3.1005
R8975 VDD.n436 VDD.n435 3.1005
R8976 VDD.n453 VDD.n452 3.1005
R8977 VDD.n457 VDD.n456 3.1005
R8978 VDD.n461 VDD.n460 3.1005
R8979 VDD.n471 VDD.n470 3.1005
R8980 VDD.n475 VDD.n474 3.1005
R8981 VDD.n117 VDD.n116 3.1005
R8982 VDD.n122 VDD.n121 3.1005
R8983 VDD.n75 VDD.n74 3.1005
R8984 VDD.n2924 VDD.n2923 3.1005
R8985 VDD.n3084 VDD.n3083 3.1005
R8986 VDD.n2984 VDD.n2983 3.1005
R8987 VDD.n2991 VDD.n2990 3.1005
R8988 VDD.n3117 VDD.n3116 3.1005
R8989 VDD.n3183 VDD.n3182 3.1005
R8990 VDD.n3189 VDD.n3188 3.1005
R8991 VDD.n3195 VDD.n3194 3.1005
R8992 VDD.n3131 VDD.n3130 3.1005
R8993 VDD.n2782 VDD.n2781 3.1005
R8994 VDD.n2786 VDD.n2785 3.1005
R8995 VDD.n3079 VDD.n3078 3.1005
R8996 VDD.n3019 VDD.n3018 3.1005
R8997 VDD.n3014 VDD.n3013 3.1005
R8998 VDD.n2960 VDD.n2959 3.1005
R8999 VDD.n2953 VDD.n2952 3.1005
R9000 VDD.n2919 VDD.n2918 3.1005
R9001 VDD.n2947 VDD.n2946 3.1005
R9002 VDD.n3053 VDD.n3052 3.1005
R9003 VDD.n2891 VDD.n2890 3.1005
R9004 VDD.n2885 VDD.n2884 3.1005
R9005 VDD.n2848 VDD.n2847 3.1005
R9006 VDD.n2883 VDD.n2882 3.1005
R9007 VDD.n2819 VDD.n2818 3.1005
R9008 VDD.n2823 VDD.n2822 3.1005
R9009 VDD.n52 VDD.n51 3.1005
R9010 VDD.n45 VDD.n44 3.1005
R9011 VDD.n23 VDD.n22 3.1005
R9012 VDD.n71 VDD.n70 3.1005
R9013 VDD.n8 VDD.n7 3.1005
R9014 VDD.n6 VDD.n5 3.1005
R9015 VDD.n4862 VDD.n4861 3.1005
R9016 VDD.n100 VDD.n99 3.1005
R9017 VDD.n106 VDD.n105 3.1005
R9018 VDD.n113 VDD.n112 3.1005
R9019 VDD.n549 VDD.n548 3.1005
R9020 VDD.n507 VDD.n506 3.1005
R9021 VDD.n516 VDD.n515 3.1005
R9022 VDD.n524 VDD.n523 3.1005
R9023 VDD.n559 VDD.n558 3.1005
R9024 VDD.n575 VDD.n574 3.1005
R9025 VDD.n678 VDD.n677 3.1005
R9026 VDD.n706 VDD.n705 3.1005
R9027 VDD.n1131 VDD.n1130 3.1005
R9028 VDD.n1079 VDD.n1078 3.1005
R9029 VDD.n1099 VDD.n1098 3.1005
R9030 VDD.n1109 VDD.n1108 3.1005
R9031 VDD.n1113 VDD.n1112 3.1005
R9032 VDD.n1121 VDD.n1120 3.1005
R9033 VDD.n1117 VDD.n1116 3.1005
R9034 VDD.n1125 VDD.n1124 3.1005
R9035 VDD.n1135 VDD.n1134 3.1005
R9036 VDD.n1164 VDD.n1163 3.1005
R9037 VDD.n1160 VDD.n1159 3.1005
R9038 VDD.n1168 VDD.n1167 3.1005
R9039 VDD.n1177 VDD.n1176 3.1005
R9040 VDD.n1180 VDD.n1179 3.1005
R9041 VDD.n1066 VDD.n1065 3.1005
R9042 VDD.n701 VDD.n700 3.1005
R9043 VDD.n689 VDD.n688 3.1005
R9044 VDD.n571 VDD.n570 3.1005
R9045 VDD.n555 VDD.n554 3.1005
R9046 VDD.n520 VDD.n519 3.1005
R9047 VDD.n4188 VDD.n4187 3.1005
R9048 VDD.n4182 VDD.n4181 3.1005
R9049 VDD.n4406 VDD.n4405 3.1005
R9050 VDD.n4396 VDD.n4395 3.1005
R9051 VDD.n1563 VDD.n1562 3.1005
R9052 VDD.n1567 VDD.n1566 3.1005
R9053 VDD.n1572 VDD.n1571 3.1005
R9054 VDD.n1578 VDD.n1577 3.1005
R9055 VDD.n1581 VDD.n1580 3.1005
R9056 VDD.n2003 VDD.n2002 3.1005
R9057 VDD.n2123 VDD.n2122 3.1005
R9058 VDD.n2098 VDD.n2097 3.1005
R9059 VDD.n2094 VDD.n2093 3.1005
R9060 VDD.n2088 VDD.n2087 3.1005
R9061 VDD.n2084 VDD.n2083 3.1005
R9062 VDD.n2080 VDD.n2079 3.1005
R9063 VDD.n2076 VDD.n2075 3.1005
R9064 VDD.n2072 VDD.n2071 3.1005
R9065 VDD.n2067 VDD.n2066 3.1005
R9066 VDD.n2063 VDD.n2062 3.1005
R9067 VDD.n2059 VDD.n2058 3.1005
R9068 VDD.n2054 VDD.n2053 3.1005
R9069 VDD.n2026 VDD.n2025 3.1005
R9070 VDD.n2022 VDD.n2021 3.1005
R9071 VDD.n2018 VDD.n2017 3.1005
R9072 VDD.n2012 VDD.n2011 3.1005
R9073 VDD.n2350 VDD.n2349 3.1005
R9074 VDD.n2359 VDD.n2358 3.1005
R9075 VDD.n2363 VDD.n2362 3.1005
R9076 VDD.n2369 VDD.n2368 3.1005
R9077 VDD.n2513 VDD.n2512 3.1005
R9078 VDD.n2509 VDD.n2508 3.1005
R9079 VDD.n4695 VDD.n4694 3.1005
R9080 VDD.n4689 VDD.n4688 3.1005
R9081 VDD.n4685 VDD.n4684 3.1005
R9082 VDD.n4681 VDD.n4680 3.1005
R9083 VDD.n4677 VDD.n4676 3.1005
R9084 VDD.n4667 VDD.n4666 3.1005
R9085 VDD.n4663 VDD.n4662 3.1005
R9086 VDD.n4659 VDD.n4658 3.1005
R9087 VDD.n4654 VDD.n4653 3.1005
R9088 VDD.n4650 VDD.n4649 3.1005
R9089 VDD.n4636 VDD.n4635 3.1005
R9090 VDD.n4632 VDD.n4631 3.1005
R9091 VDD.n4628 VDD.n4627 3.1005
R9092 VDD.n4622 VDD.n4621 3.1005
R9093 VDD.n4620 VDD.n4619 3.1005
R9094 VDD.n4615 VDD.n4614 3.1005
R9095 VDD.n4606 VDD.n4605 3.1005
R9096 VDD.n4556 VDD.n4555 3.1005
R9097 VDD.n4571 VDD.n4570 3.1005
R9098 VDD.n2579 VDD.n2578 3.1005
R9099 VDD.n2583 VDD.n2582 3.1005
R9100 VDD.n2587 VDD.n2586 3.1005
R9101 VDD.n4525 VDD.n4524 3.1005
R9102 VDD.n4521 VDD.n4520 3.1005
R9103 VDD.n4517 VDD.n4516 3.1005
R9104 VDD.n4512 VDD.n4511 3.1005
R9105 VDD.n4492 VDD.n4491 3.1005
R9106 VDD.n4488 VDD.n4487 3.1005
R9107 VDD.n4484 VDD.n4483 3.1005
R9108 VDD.n4478 VDD.n4477 3.1005
R9109 VDD.n4473 VDD.n4472 3.1005
R9110 VDD.n4470 VDD.n4469 3.1005
R9111 VDD.n4465 VDD.n4464 3.1005
R9112 VDD.n4461 VDD.n4460 3.1005
R9113 VDD.n4457 VDD.n4456 3.1005
R9114 VDD.n4432 VDD.n4431 3.1005
R9115 VDD.n2606 VDD.n2605 3.1005
R9116 VDD.n2602 VDD.n2601 3.1005
R9117 VDD.n4324 VDD.n4323 3.1005
R9118 VDD.n4328 VDD.n4327 3.1005
R9119 VDD.n4332 VDD.n4331 3.1005
R9120 VDD.n4310 VDD.n4309 3.1005
R9121 VDD.n4306 VDD.n4305 3.1005
R9122 VDD.n4300 VDD.n4299 3.1005
R9123 VDD.n4295 VDD.n4294 3.1005
R9124 VDD.n4292 VDD.n4291 3.1005
R9125 VDD.n4287 VDD.n4286 3.1005
R9126 VDD.n4283 VDD.n4282 3.1005
R9127 VDD.n4279 VDD.n4278 3.1005
R9128 VDD.n4254 VDD.n4253 3.1005
R9129 VDD.n4250 VDD.n4249 3.1005
R9130 VDD.n4244 VDD.n4243 3.1005
R9131 VDD.n4240 VDD.n4239 3.1005
R9132 VDD.n4236 VDD.n4235 3.1005
R9133 VDD.n4232 VDD.n4231 3.1005
R9134 VDD.n2637 VDD.n2636 3.1005
R9135 VDD.n4124 VDD.n4123 3.1005
R9136 VDD.n2539 VDD.n2538 3.1005
R9137 VDD.n4795 VDD.n4794 3.1005
R9138 VDD.n2696 VDD.n2695 3.1005
R9139 VDD.n2756 VDD.n2755 3.1005
R9140 VDD.n3296 VDD.n3295 3.1005
R9141 VDD.n3308 VDD.n3307 3.1005
R9142 VDD.n3217 VDD.n3216 3.1005
R9143 VDD.n3292 VDD.n3291 3.1005
R9144 VDD.n3280 VDD.n3279 3.1005
R9145 VDD.n2714 VDD.n2713 3.1005
R9146 VDD.n2710 VDD.n2709 3.1005
R9147 VDD.n2732 VDD.n2731 3.1005
R9148 VDD.n3387 VDD.n3386 3.1005
R9149 VDD.n3383 VDD.n3382 3.1005
R9150 VDD.n3377 VDD.n2734 3.1005
R9151 VDD.n3418 VDD.n3417 3.1005
R9152 VDD.n3422 VDD.n3421 3.1005
R9153 VDD.n3426 VDD.n3425 3.1005
R9154 VDD.n3430 VDD.n3429 3.1005
R9155 VDD.n3434 VDD.n3433 3.1005
R9156 VDD.n3438 VDD.n3437 3.1005
R9157 VDD.n3445 VDD.n3439 3.1005
R9158 VDD.n3451 VDD.n3450 3.1005
R9159 VDD.n3412 VDD.n3411 3.1005
R9160 VDD.n4820 VDD.n4819 3.1005
R9161 VDD.n4799 VDD.n4798 3.1005
R9162 VDD.n4790 VDD.n4789 3.1005
R9163 VDD.n4782 VDD.n4781 3.1005
R9164 VDD.n4786 VDD.n4785 3.1005
R9165 VDD.n4776 VDD.n4775 3.1005
R9166 VDD.n3392 VDD.n3391 3.09016
R9167 VDD.n1305 VDD.n1304 3.09016
R9168 VDD.n5 VDD.n2 3.09016
R9169 VDD.n2965 VDD.n2962 3.09016
R9170 VDD.n2990 VDD.n2987 3.09016
R9171 VDD.n3024 VDD.n3021 3.09016
R9172 VDD VDD.n536 3.08979
R9173 VDD VDD.n1143 3.08979
R9174 VDD VDD.n2106 3.08979
R9175 VDD VDD.n2494 3.08979
R9176 VDD VDD.n2556 3.08979
R9177 VDD VDD.n4440 3.08979
R9178 VDD VDD.n4262 3.08979
R9179 VDD.n4170 VDD.n4169 3.03311
R9180 VDD.n2451 VDD.n2450 3.03311
R9181 VDD.n1444 VDD.n1443 2.86947
R9182 VDD.n238 VDD.n236 2.86947
R9183 VDD.n2319 VDD.n2318 2.86947
R9184 VDD.n143 VDD.n140 2.86947
R9185 VDD.n3156 VDD.n3153 2.86947
R9186 VDD.n3046 VDD.n3043 2.86947
R9187 VDD.n714 VDD.n711 2.86947
R9188 VDD.n1184 VDD.n1069 2.86947
R9189 VDD.n4138 VDD.n4135 2.82084
R9190 VDD.n1868 VDD.n1867 2.64878
R9191 VDD.n2912 VDD.n2911 2.64878
R9192 VDD.n1602 VDD.n1599 2.64878
R9193 VDD.n4130 VDD.n4129 2.64594
R9194 VDD.n478 VDD.t638 2.63939
R9195 VDD.n1010 VDD.t81 2.63939
R9196 VDD.n1954 VDD.t482 2.63939
R9197 VDD.n3648 VDD.t225 2.63939
R9198 VDD.n3824 VDD.t355 2.63939
R9199 VDD.n3558 VDD.t193 2.63939
R9200 VDD.n4053 VDD.t725 2.63939
R9201 VDD.n572 VDD.t691 2.63208
R9202 VDD.n739 VDD.n738 2.63208
R9203 VDD.n1114 VDD.t395 2.63208
R9204 VDD.n2077 VDD.t72 2.63208
R9205 VDD.n2051 VDD.n2050 2.63208
R9206 VDD.n2037 VDD.n2036 2.63208
R9207 VDD.n4682 VDD.t166 2.63208
R9208 VDD.n4646 VDD.n4645 2.63208
R9209 VDD.n2576 VDD.t452 2.63208
R9210 VDD.n4503 VDD.n4502 2.63208
R9211 VDD.n4321 VDD.t254 2.63208
R9212 VDD.n4357 VDD.n4356 2.63208
R9213 VDD.n4374 VDD.n4373 2.63208
R9214 VDD.n4233 VDD.t473 2.63208
R9215 VDD.n4151 VDD.n4150 2.63208
R9216 VDD.n323 VDD.n322 2.61039
R9217 VDD.n337 VDD.n336 2.61039
R9218 VDD.n351 VDD.n350 2.61039
R9219 VDD.n365 VDD.n364 2.61039
R9220 VDD.n379 VDD.n378 2.61039
R9221 VDD.n393 VDD.n392 2.61039
R9222 VDD.n407 VDD.n406 2.61039
R9223 VDD.n786 VDD.n785 2.61039
R9224 VDD.n1295 VDD.t618 2.61039
R9225 VDD.n1480 VDD.n1479 2.61039
R9226 VDD.n1477 VDD.n1437 2.61039
R9227 VDD.n1459 VDD.n1458 2.61039
R9228 VDD.n233 VDD.n232 2.61039
R9229 VDD.n2163 VDD.n2162 2.61039
R9230 VDD.n2177 VDD.n2176 2.61039
R9231 VDD.n2193 VDD.n2192 2.61039
R9232 VDD.n2207 VDD.n2206 2.61039
R9233 VDD.n2230 VDD.n2229 2.61039
R9234 VDD.n2310 VDD.n2309 2.61039
R9235 VDD.n2314 VDD.n2313 2.61039
R9236 VDD.n199 VDD.n198 2.61039
R9237 VDD.n1856 VDD.n1855 2.61039
R9238 VDD.n1874 VDD.n1873 2.61039
R9239 VDD.n2390 VDD.n2389 2.61039
R9240 VDD.n2447 VDD.n2446 2.61039
R9241 VDD.n2429 VDD.n2428 2.61039
R9242 VDD.n2415 VDD.n2414 2.61039
R9243 VDD.n1001 VDD.n1000 2.55931
R9244 VDD.n1966 VDD.n1785 2.55931
R9245 VDD.n1931 VDD.n1790 2.55931
R9246 VDD.n4044 VDD.n4043 2.55931
R9247 VDD.n3679 VDD.n3678 2.55931
R9248 VDD.n3803 VDD.n3802 2.55931
R9249 VDD.n3877 VDD.n3876 2.55931
R9250 VDD.n3956 VDD.n3955 2.55931
R9251 VDD.n467 VDD.n466 2.55931
R9252 VDD.n1105 VDD.n1104 2.55931
R9253 VDD.n685 VDD.n684 2.55931
R9254 VDD.n2068 VDD.n2009 2.55931
R9255 VDD.n4673 VDD.n4672 2.55931
R9256 VDD.n2643 VDD.n2642 2.55931
R9257 VDD.n2472 VDD.n2471 2.5593
R9258 VDD.n1723 VDD.n1722 2.52719
R9259 VDD.n1918 VDD.n1794 2.52719
R9260 VDD.n3696 VDD.n3695 2.52719
R9261 VDD.n3894 VDD.n3893 2.52719
R9262 VDD.n1173 VDD.n1172 2.52719
R9263 VDD.n512 VDD.n511 2.52719
R9264 VDD.n1610 VDD.n1609 2.52719
R9265 VDD.n2355 VDD.n2354 2.52719
R9266 VDD.n4611 VDD.n4610 2.52719
R9267 VDD.n4466 VDD.n2597 2.52719
R9268 VDD.n4288 VDD.n2632 2.52719
R9269 VDD.n949 VDD.n948 2.49102
R9270 VDD.n3992 VDD.n3991 2.49102
R9271 VDD.n3255 VDD.n3248 2.49102
R9272 VDD.n3704 VDD.n3702 2.49102
R9273 VDD.n3904 VDD.n3903 2.49102
R9274 VDD.n1913 VDD.n1796 2.49102
R9275 VDD.n1734 VDD.n1733 2.49102
R9276 VDD.n3181 VDD.n3180 2.49102
R9277 VDD.n3144 VDD.n3143 2.49102
R9278 VDD.n2861 VDD.n2860 2.49102
R9279 VDD.n1178 VDD.n1074 2.49102
R9280 VDD.n503 VDD.n502 2.49102
R9281 VDD.n1597 VDD.n1596 2.49102
R9282 VDD.n2346 VDD.n2345 2.49102
R9283 VDD.n4618 VDD.n4617 2.49102
R9284 VDD.n4471 VDD.n2593 2.49102
R9285 VDD.n4293 VDD.n2628 2.49102
R9286 VDD.n533 VDD 2.46127
R9287 VDD.n1140 VDD 2.46127
R9288 VDD.n2103 VDD 2.46127
R9289 VDD.n2491 VDD 2.46127
R9290 VDD.n2553 VDD 2.46127
R9291 VDD.n4437 VDD 2.46127
R9292 VDD.n4259 VDD 2.46127
R9293 VDD.n818 VDD.n811 2.42809
R9294 VDD.n820 VDD.n818 2.42809
R9295 VDD.n832 VDD.n825 2.42809
R9296 VDD.n834 VDD.n832 2.42809
R9297 VDD.n849 VDD.n842 2.42809
R9298 VDD.n851 VDD.n849 2.42809
R9299 VDD.n863 VDD.n856 2.42809
R9300 VDD.n865 VDD.n863 2.42809
R9301 VDD.n877 VDD.n870 2.42809
R9302 VDD.n879 VDD.n877 2.42809
R9303 VDD.n912 VDD.n905 2.42809
R9304 VDD.n892 VDD.n885 2.42809
R9305 VDD.n894 VDD.n892 2.42809
R9306 VDD.n1204 VDD.n278 2.42809
R9307 VDD.n1204 VDD.n1203 2.42809
R9308 VDD.n1211 VDD.n271 2.42809
R9309 VDD.n1372 VDD.n1365 2.42809
R9310 VDD.n1374 VDD.n1372 2.42809
R9311 VDD.n1389 VDD.n1382 2.42809
R9312 VDD.n1407 VDD.n1400 2.42809
R9313 VDD.n1409 VDD.n1407 2.42809
R9314 VDD.n1644 VDD.n1637 2.42809
R9315 VDD.n1646 VDD.n1644 2.42809
R9316 VDD.n1658 VDD.n1651 2.42809
R9317 VDD.n1660 VDD.n1658 2.42809
R9318 VDD.n1689 VDD.n1682 2.42809
R9319 VDD.n1673 VDD.n1666 2.42809
R9320 VDD.n1675 VDD.n1673 2.42809
R9321 VDD.n1505 VDD.n1497 2.42809
R9322 VDD.n1505 VDD.n1504 2.42809
R9323 VDD.n1512 VDD.n1490 2.42809
R9324 VDD.n1878 VDD.n1877 2.42809
R9325 VDD.n3547 VDD.n3544 2.42809
R9326 VDD.n126 VDD.n125 2.42809
R9327 VDD.n3161 VDD 2.42809
R9328 VDD.n1093 VDD.n1090 2.42809
R9329 VDD.n2932 VDD.n2929 2.32777
R9330 VDD.n2466 VDD.n2465 2.28739
R9331 VDD.n1836 VDD.n1835 2.28739
R9332 VDD.n3618 VDD.n3617 2.28739
R9333 VDD.n1714 VDD.n1713 2.28739
R9334 VDD.n57 VDD.n56 2.28739
R9335 VDD.n742 VDD.n741 2.28739
R9336 VDD.n695 VDD.n694 2.28739
R9337 VDD.n4401 VDD.n4400 2.28739
R9338 VDD.n2128 VDD.n2127 2.28739
R9339 VDD.n4427 VDD.n4426 2.28739
R9340 VDD.n3288 VDD.n3287 2.28739
R9341 VDD.n3222 VDD.n3221 2.28739
R9342 VDD.n2547 VDD.n2546 2.28323
R9343 VDD.n1391 VDD.n1390 2.2074
R9344 VDD.n2296 VDD.n2295 2.2074
R9345 VDD.n2818 VDD.n2817 2.2074
R9346 VDD.n4269 VDD.n4268 2.2074
R9347 VDD.n4447 VDD.n4446 2.2074
R9348 VDD.n2563 VDD.n2562 2.2074
R9349 VDD.n2501 VDD.n2500 2.2074
R9350 VDD.n2113 VDD.n2112 2.2074
R9351 VDD.n1150 VDD.n1149 2.2074
R9352 VDD.n543 VDD.n542 2.2074
R9353 VDD.n4029 VDD.n4026 2.19751
R9354 VDD.n3941 VDD.n3940 2.19751
R9355 VDD.n452 VDD.n449 2.19751
R9356 VDD.n986 VDD.n983 2.19751
R9357 VDD.n1978 VDD.n1975 2.19751
R9358 VDD.n1835 VDD.n1832 2.19751
R9359 VDD.n4405 VDD.n4402 2.19751
R9360 VDD.n4516 VDD.n4513 2.19751
R9361 VDD.n4658 VDD.n4655 2.19751
R9362 VDD.n2058 VDD.n2055 2.19751
R9363 VDD.n1078 VDD.n1075 2.19751
R9364 VDD.n700 VDD.n697 2.19751
R9365 VDD.n295 VDD.n293 2.16388
R9366 VDD.n3245 VDD.n3243 2.16388
R9367 VDD.n2677 VDD.n2675 2.16388
R9368 VDD.n1044 VDD.n1041 2.02155
R9369 VDD.n631 VDD.n628 2.02155
R9370 VDD.n4274 VDD.n4272 2.02155
R9371 VDD.n4341 VDD.n4338 2.02155
R9372 VDD.n4452 VDD.n4450 2.02155
R9373 VDD.n4533 VDD.n4530 2.02155
R9374 VDD.n2546 VDD.n2544 2.02155
R9375 VDD.n2485 VDD.n2483 2.02155
R9376 VDD.n2118 VDD.n2116 2.02155
R9377 VDD.n1155 VDD.n1153 2.02155
R9378 VDD.n527 VDD.n525 2.02155
R9379 VDD.n9 VDD.n8 2.01076
R9380 VDD.n1693 VDD.n1692 1.98671
R9381 VDD.n4804 VDD.n4801 1.98671
R9382 VDD.n1944 VDD.n1941 1.98671
R9383 VDD.n1026 VDD.n1023 1.98671
R9384 VDD.n4069 VDD.n4066 1.98671
R9385 VDD.n3534 VDD.n3531 1.98671
R9386 VDD.n3571 VDD.n3570 1.98671
R9387 VDD.n3852 VDD.n3849 1.98671
R9388 VDD.n3841 VDD.n3840 1.98671
R9389 VDD.n3664 VDD.n3661 1.98671
R9390 VDD.n29 VDD.n26 1.98671
R9391 VDD.n2775 VDD.n2774 1.98671
R9392 VDD.n4249 VDD.n4246 1.98671
R9393 VDD.n4426 VDD.n4423 1.98671
R9394 VDD.n2508 VDD.n2507 1.98671
R9395 VDD.n2093 VDD.n2090 1.98671
R9396 VDD.n1130 VDD.n1127 1.98671
R9397 VDD.n554 VDD.n551 1.98671
R9398 VDD.n3815 VDD.n3814 1.94045
R9399 VDD.n3835 VDD.n3834 1.94045
R9400 VDD.n4866 VDD.n4864 1.94045
R9401 VDD.n2374 VDD.n2373 1.94045
R9402 VDD.n2515 VDD.n2514 1.94045
R9403 VDD.n4699 VDD.n4698 1.94045
R9404 VDD.n4710 VDD.n4709 1.94045
R9405 VDD.n3319 VDD.n3318 1.94045
R9406 VDD.n3515 VDD.n3514 1.94045
R9407 VDD.n3513 VDD.n3512 1.94045
R9408 VDD.n3405 VDD.n3404 1.94045
R9409 VDD.n583 VDD.n582 1.94045
R9410 VDD.n4837 VDD.n4836 1.94045
R9411 VDD.n779 VDD.n778 1.94045
R9412 VDD VDD.n2920 1.92238
R9413 VDD.n538 VDD 1.91393
R9414 VDD.n1145 VDD 1.91393
R9415 VDD.n2108 VDD 1.91393
R9416 VDD.n2496 VDD 1.91393
R9417 VDD.n2558 VDD 1.91393
R9418 VDD.n4442 VDD 1.91393
R9419 VDD.n4264 VDD 1.91393
R9420 VDD.n4098 VDD.n4097 1.84226
R9421 VDD.n3489 VDD.n3486 1.76602
R9422 VDD.n913 VDD.n902 1.76602
R9423 VDD.n480 VDD.n477 1.76602
R9424 VDD.n534 VDD.n533 1.75668
R9425 VDD.n1141 VDD.n1140 1.75668
R9426 VDD.n2104 VDD.n2103 1.75668
R9427 VDD.n2492 VDD.n2491 1.75668
R9428 VDD.n2554 VDD.n2553 1.75668
R9429 VDD.n4438 VDD.n4437 1.75668
R9430 VDD.n4260 VDD.n4259 1.75668
R9431 VDD.n4649 VDD.n4648 1.62438
R9432 VDD.n2053 VDD.n2046 1.62438
R9433 VDD.n741 VDD.n734 1.62438
R9434 VDD.n726 VDD.n721 1.62438
R9435 VDD.n1797 VDD.n1796 1.57241
R9436 VDD.n1733 VDD.n1732 1.57241
R9437 VDD.n3903 VDD.n3902 1.57241
R9438 VDD.n3249 VDD.n3248 1.57241
R9439 VDD.n3991 VDD.n3990 1.57241
R9440 VDD.n3705 VDD.n3704 1.57241
R9441 VDD.n948 VDD.n947 1.57241
R9442 VDD.n3143 VDD.n3142 1.57241
R9443 VDD.n2860 VDD.n2859 1.57241
R9444 VDD.n3180 VDD.n3179 1.57241
R9445 VDD.n1074 VDD.n1072 1.57241
R9446 VDD.n502 VDD.n501 1.57241
R9447 VDD.n2345 VDD.n2344 1.57241
R9448 VDD.n1596 VDD.n1595 1.57241
R9449 VDD.n2593 VDD.n2591 1.57241
R9450 VDD.n2628 VDD.n2626 1.57241
R9451 VDD.n2701 VDD.n2698 1.54533
R9452 VDD.n1519 VDD.n1518 1.54533
R9453 VDD.n2297 VDD.n2296 1.54533
R9454 VDD.n3604 VDD.n3603 1.54533
R9455 VDD.n3821 VDD.n3818 1.54533
R9456 VDD.n564 VDD.n561 1.54533
R9457 VDD.n4269 VDD.n4267 1.54533
R9458 VDD.n4447 VDD.n4445 1.54533
R9459 VDD.n2563 VDD.n2561 1.54533
R9460 VDD.n2501 VDD.n2499 1.54533
R9461 VDD.n2113 VDD.n2111 1.54533
R9462 VDD.n1150 VDD.n1148 1.54533
R9463 VDD.n543 VDD.n541 1.54533
R9464 VDD.n4023 VDD.n4021 1.52886
R9465 VDD.n3935 VDD.n3933 1.52886
R9466 VDD.n3736 VDD.n3734 1.52886
R9467 VDD.n446 VDD.n444 1.52886
R9468 VDD.n980 VDD.n978 1.52886
R9469 VDD.n1823 VDD.n1821 1.52886
R9470 VDD.n4378 VDD.n4377 1.52886
R9471 VDD.n4498 VDD.n4497 1.52886
R9472 VDD.n2045 VDD.n2044 1.52886
R9473 VDD.n2032 VDD.n2031 1.52886
R9474 VDD.n733 VDD.n732 1.52886
R9475 VDD.n4146 VDD.n4145 1.51754
R9476 VDD.n1794 VDD.n1793 1.47868
R9477 VDD.n3893 VDD.n3892 1.47868
R9478 VDD.n3695 VDD.n3694 1.47868
R9479 VDD.n1722 VDD.n1721 1.47868
R9480 VDD.n511 VDD.n510 1.47868
R9481 VDD.n1172 VDD.n1171 1.47868
R9482 VDD.n4610 VDD.n4609 1.47868
R9483 VDD.n2354 VDD.n2353 1.47868
R9484 VDD.n1609 VDD.n1608 1.47868
R9485 VDD.n2597 VDD.n2596 1.47868
R9486 VDD.n2632 VDD.n2631 1.47868
R9487 VDD.n4097 VDD.n4096 1.47016
R9488 VDD.n1542 VDD.n1541 1.43334
R9489 VDD.n1550 VDD.n1548 1.43334
R9490 VDD.n1785 VDD.n1784 1.39551
R9491 VDD.n1790 VDD.n1789 1.39551
R9492 VDD.n3876 VDD.n3875 1.39551
R9493 VDD.n3955 VDD.n3954 1.39551
R9494 VDD.n4043 VDD.n4042 1.39551
R9495 VDD.n3678 VDD.n3677 1.39551
R9496 VDD.n3802 VDD.n3801 1.39551
R9497 VDD.n1000 VDD.n999 1.39551
R9498 VDD.n466 VDD.n465 1.39551
R9499 VDD.n684 VDD.n683 1.39551
R9500 VDD.n1104 VDD.n1103 1.39551
R9501 VDD.n4672 VDD.n4671 1.39551
R9502 VDD.n2009 VDD.n2008 1.39551
R9503 VDD.n2642 VDD.n2641 1.39551
R9504 VDD.n2471 VDD.n2470 1.39505
R9505 VDD.n670 VDD.n669 1.35607
R9506 VDD.n3552 VDD.n3551 1.35607
R9507 VDD.n3625 VDD.n3624 1.35607
R9508 VDD.n4081 VDD.n4080 1.35607
R9509 VDD.n3981 VDD.n3980 1.35607
R9510 VDD.n2664 VDD.n2662 1.35607
R9511 VDD.n4106 VDD.n4104 1.35607
R9512 VDD.n3776 VDD.n3775 1.35607
R9513 VDD.n3577 VDD.n3575 1.35607
R9514 VDD.n938 VDD.n937 1.35607
R9515 VDD.n491 VDD.n489 1.35607
R9516 VDD.n610 VDD.n608 1.35607
R9517 VDD.n635 VDD.n633 1.35607
R9518 VDD.n1048 VDD.n1046 1.35607
R9519 VDD.n1993 VDD.n1991 1.35607
R9520 VDD.n1894 VDD.n1893 1.35607
R9521 VDD.n1840 VDD.n1837 1.35607
R9522 VDD.n3262 VDD.n3261 1.35607
R9523 VDD.n3174 VDD.n3173 1.35607
R9524 VDD.n134 VDD.n133 1.35607
R9525 VDD.n36 VDD.n35 1.35607
R9526 VDD.n2834 VDD.n2833 1.35607
R9527 VDD.n2908 VDD.n2907 1.35607
R9528 VDD.n3088 VDD.n3086 1.35607
R9529 VDD.n3057 VDD.n3055 1.35607
R9530 VDD.n2876 VDD.n2875 1.35607
R9531 VDD.n2865 VDD.n2863 1.35607
R9532 VDD.n2936 VDD.n2934 1.35607
R9533 VDD.n3148 VDD.n3146 1.35607
R9534 VDD.n3031 VDD.n3030 1.35607
R9535 VDD.n1087 VDD.n1086 1.35607
R9536 VDD.n579 VDD.n577 1.35607
R9537 VDD.n1555 VDD.n1554 1.35607
R9538 VDD.n1586 VDD.n1585 1.35607
R9539 VDD.n1613 VDD.n1612 1.35607
R9540 VDD.n2130 VDD.n2129 1.35607
R9541 VDD.n4197 VDD.n4195 1.35607
R9542 VDD.n4409 VDD.n4408 1.35607
R9543 VDD.n4421 VDD.n4420 1.35607
R9544 VDD.n2335 VDD.n2334 1.35607
R9545 VDD.n4594 VDD.n4593 1.35607
R9546 VDD.n4537 VDD.n4535 1.35607
R9547 VDD.n4345 VDD.n4343 1.35607
R9548 VDD.n4313 VDD.n4312 1.35607
R9549 VDD.n4834 VDD.n4833 1.35607
R9550 VDD.n1414 VDD.n1413 1.35607
R9551 VDD.n2136 VDD.n217 1.35607
R9552 VDD.n4810 VDD.n4808 1.35607
R9553 VDD.n2718 VDD.n2716 1.35607
R9554 VDD.n3226 VDD.n3223 1.35607
R9555 VDD.n2153 VDD.n2152 1.35607
R9556 VDD.n1524 VDD.n1522 1.35607
R9557 VDD.n917 VDD.n915 1.35607
R9558 VDD.n1199 VDD.n1198 1.35607
R9559 VDD.n2454 VDD.n2452 1.35607
R9560 VDD.n3796 VDD.n3795 1.35607
R9561 VDD.n3972 VDD.n3970 1.35607
R9562 VDD.n3642 VDD.n3641 1.35607
R9563 VDD.n1710 VDD.n1709 1.35607
R9564 VDD.n1763 VDD.n1761 1.35607
R9565 VDD.n2476 VDD.n2474 1.35607
R9566 VDD.n3103 VDD.n3102 1.35607
R9567 VDD.n3002 VDD.n3000 1.35607
R9568 VDD.n61 VDD.n58 1.35607
R9569 VDD.n89 VDD.n87 1.35607
R9570 VDD.n150 VDD.n148 1.35607
R9571 VDD.n2971 VDD.n2969 1.35607
R9572 VDD.n3199 VDD.n3197 1.35607
R9573 VDD.n1190 VDD.n1188 1.35607
R9574 VDD.n4172 VDD.n4171 1.35607
R9575 VDD.n4220 VDD.n4219 1.35607
R9576 VDD.n2569 VDD.n2567 1.35607
R9577 VDD.n4584 VDD.n4582 1.35607
R9578 VDD.n4384 VDD.n4382 1.35607
R9579 VDD.n3311 VDD.n3310 1.35607
R9580 VDD.n3397 VDD.n3396 1.35607
R9581 VDD.n1883 VDD.n1881 1.35607
R9582 VDD.n1472 VDD.n1471 1.35607
R9583 VDD.n1698 VDD.n1696 1.35607
R9584 VDD.n2324 VDD.n2322 1.35607
R9585 VDD.n1989 VDD.n1985 1.33781
R9586 VDD.n1987 VDD.n1986 1.33781
R9587 VDD.n4162 VDD.n4161 1.32791
R9588 VDD.n811 VDD.n810 1.32464
R9589 VDD.n820 VDD.n819 1.32464
R9590 VDD.n825 VDD.n824 1.32464
R9591 VDD.n834 VDD.n833 1.32464
R9592 VDD.n842 VDD.n841 1.32464
R9593 VDD.n851 VDD.n850 1.32464
R9594 VDD.n856 VDD.n855 1.32464
R9595 VDD.n865 VDD.n864 1.32464
R9596 VDD.n870 VDD.n869 1.32464
R9597 VDD.n879 VDD.n878 1.32464
R9598 VDD.n902 VDD.n901 1.32464
R9599 VDD.n885 VDD.n884 1.32464
R9600 VDD.n894 VDD.n893 1.32464
R9601 VDD.n278 VDD.n277 1.32464
R9602 VDD.n271 VDD.n270 1.32464
R9603 VDD.n1221 VDD.n1211 1.32464
R9604 VDD.n1220 VDD.n1219 1.32464
R9605 VDD.n1219 VDD.n1218 1.32464
R9606 VDD.n1365 VDD.n1364 1.32464
R9607 VDD.n1374 VDD.n1373 1.32464
R9608 VDD.n1382 VDD.n1381 1.32464
R9609 VDD.n1392 VDD.n1391 1.32464
R9610 VDD.n1400 VDD.n1399 1.32464
R9611 VDD.n1409 VDD.n1408 1.32464
R9612 VDD.n1637 VDD.n1636 1.32464
R9613 VDD.n1646 VDD.n1645 1.32464
R9614 VDD.n1651 VDD.n1650 1.32464
R9615 VDD.n1660 VDD.n1659 1.32464
R9616 VDD.n1682 VDD.n1681 1.32464
R9617 VDD.n1692 VDD.n1691 1.32464
R9618 VDD.n1666 VDD.n1665 1.32464
R9619 VDD.n1675 VDD.n1674 1.32464
R9620 VDD.n1497 VDD.n1496 1.32464
R9621 VDD.n1490 VDD.n1489 1.32464
R9622 VDD.n1518 VDD.n1517 1.32464
R9623 VDD.n4732 VDD.n4729 1.32464
R9624 VDD.n4825 VDD.n4822 1.32464
R9625 VDD.n599 VDD.n596 1.32464
R9626 VDD.n4004 VDD.n4001 1.32464
R9627 VDD.n3961 VDD.n3958 1.32464
R9628 VDD.n3916 VDD.n3913 1.32464
R9629 VDD.n3717 VDD.n3714 1.32464
R9630 VDD.n427 VDD.n424 1.32464
R9631 VDD.n961 VDD.n958 1.32464
R9632 VDD.n1746 VDD.n1743 1.32464
R9633 VDD.n1904 VDD.n1901 1.32464
R9634 VDD.n85 VDD.n84 1.32464
R9635 VDD.n3111 VDD.n3110 1.32464
R9636 VDD.n3164 VDD.n3161 1.32464
R9637 VDD.n4305 VDD.n4302 1.32464
R9638 VDD.n4483 VDD.n4480 1.32464
R9639 VDD.n4578 VDD.n4577 1.32464
R9640 VDD.n4627 VDD.n4626 1.32464
R9641 VDD.n2017 VDD.n2014 1.32464
R9642 VDD.n1577 VDD.n1574 1.32464
R9643 VDD.n1065 VDD.n1062 1.32464
R9644 VDD.n4187 VDD.n4184 1.30219
R9645 VDD.n4368 VDD.n4366 1.24229
R9646 VDD.n4160 VDD.n4159 1.23309
R9647 VDD.n4129 VDD.n4128 1.17153
R9648 VDD.n4351 VDD.n4350 1.14677
R9649 VDD.n4640 VDD.n4638 1.14677
R9650 VDD.n4416 VDD.n4415 1.13857
R9651 VDD.n2902 VDD.n2901 1.13857
R9652 VDD.n2770 VDD.n2769 1.13845
R9653 VDD.n3511 VDD.n2725 1.13845
R9654 VDD.n4814 VDD.n168 1.13845
R9655 VDD.n159 VDD.n158 1.13845
R9656 VDD.n2906 VDD.n2904 1.13745
R9657 VDD.n4175 VDD.n4174 1.13469
R9658 VDD.n4216 VDD.n4215 1.13469
R9659 VDD.n3315 VDD.n3314 1.13469
R9660 VDD.n3314 VDD.n3313 1.13469
R9661 VDD.n4214 VDD.n4213 1.13469
R9662 VDD.n3203 VDD.n3202 1.13469
R9663 VDD.n3555 VDD.n3554 1.13469
R9664 VDD.n3519 VDD.n3399 1.13469
R9665 VDD.n2725 VDD.n2724 1.13469
R9666 VDD.n3519 VDD.n3518 1.13469
R9667 VDD.n3976 VDD.n3975 1.13469
R9668 VDD.n4388 VDD.n4387 1.13469
R9669 VDD.n4841 VDD.n4840 1.13469
R9670 VDD.n2573 VDD.n2572 1.13469
R9671 VDD.n4588 VDD.n4587 1.13469
R9672 VDD.n4550 VDD.n4549 1.13469
R9673 VDD.n93 VDD.n64 1.13469
R9674 VDD.n93 VDD.n92 1.13469
R9675 VDD.n137 VDD.n136 1.13469
R9676 VDD.n154 VDD.n153 1.13469
R9677 VDD.n4813 VDD.n4812 1.13458
R9678 VDD.n2725 VDD.n2720 1.13458
R9679 VDD.n4590 VDD.n4589 1.13458
R9680 VDD.n4551 VDD.n4539 1.13458
R9681 VDD.n4418 VDD.n4417 1.13458
R9682 VDD.n4388 VDD.n4347 1.13458
R9683 VDD.n4416 VDD.n4411 1.13458
R9684 VDD.n3594 VDD.n3593 1.13458
R9685 VDD.n3977 VDD.n3976 1.13458
R9686 VDD.n2667 VDD.n2666 1.13458
R9687 VDD.n4109 VDD.n4108 1.13458
R9688 VDD.n4084 VDD.n4083 1.13458
R9689 VDD.n3628 VDD.n3627 1.13458
R9690 VDD.n3772 VDD.n3771 1.13458
R9691 VDD.n3580 VDD.n3579 1.13458
R9692 VDD.n3265 VDD.n3264 1.13458
R9693 VDD.n3273 VDD.n3235 1.13458
R9694 VDD.n3229 VDD.n3228 1.13458
R9695 VDD.n4214 VDD.n4199 1.13458
R9696 VDD.n2770 VDD.n2765 1.13458
R9697 VDD.n39 VDD.n38 1.13458
R9698 VDD.n3203 VDD.n3150 1.13458
R9699 VDD.n3203 VDD.n2771 1.13458
R9700 VDD.n4209 VDD.n4205 1.13458
R9701 VDD.n4388 VDD.n4315 1.13458
R9702 VDD.n4841 VDD.n165 1.13458
R9703 VDD.n1221 VDD.n1220 1.10395
R9704 VDD.n1878 VDD.n1866 1.10395
R9705 VDD.n1757 VDD.n1756 1.10395
R9706 VDD.n2882 VDD.n2879 1.10395
R9707 VDD.n81 VDD.n78 1.10395
R9708 VDD.n3194 VDD.n3191 1.10395
R9709 VDD.n3043 VDD.n3042 1.10395
R9710 VDD.n2368 VDD.n2365 1.10395
R9711 VDD.n2340 VDD.n182 1.10395
R9712 VDD.n1591 VDD.n1535 1.10395
R9713 VDD.n4496 VDD.n4494 1.05125
R9714 VDD.n2030 VDD.n2028 1.05125
R9715 VDD.n720 VDD.n718 1.05125
R9716 VDD.n3863 VDD.n3862 1.04225
R9717 VDD.n744 VDD.n742 1.04225
R9718 VDD.n2932 VDD.n2931 0.970197
R9719 VDD.n3746 VDD.n3745 0.955724
R9720 VDD.n4144 VDD.n4142 0.948648
R9721 VDD.n295 VDD.n294 0.901908
R9722 VDD.n3245 VDD.n3244 0.901908
R9723 VDD.n2677 VDD.n2676 0.901908
R9724 VDD.n281 VDD.n280 0.883259
R9725 VDD.n1500 VDD.n1499 0.883259
R9726 VDD.n1519 VDD.n1512 0.883259
R9727 VDD.n1517 VDD.n1516 0.883259
R9728 VDD.n1869 VDD.n1868 0.883259
R9729 VDD.n4853 VDD.n4850 0.883259
R9730 VDD.n2836 VDD.n2835 0.883259
R9731 VDD.n3071 VDD.n3068 0.883259
R9732 VDD.n3110 VDD.n3109 0.883259
R9733 VDD.n3121 VDD.n3120 0.883259
R9734 VDD.n4694 VDD.n4693 0.883259
R9735 VDD.n1055 VDD 0.867705
R9736 VDD.n2152 VDD.n2150 0.853
R9737 VDD.n1525 VDD.n1524 0.853
R9738 VDD.n918 VDD.n917 0.853
R9739 VDD.n1198 VDD.n1196 0.853
R9740 VDD.n2137 VDD.n2136 0.853
R9741 VDD.n1415 VDD.n1414 0.853
R9742 VDD.n2455 VDD.n2454 0.853
R9743 VDD.n4811 VDD.n4810 0.853
R9744 VDD.n2719 VDD.n2718 0.853
R9745 VDD.n2334 VDD.n2332 0.853
R9746 VDD.n4593 VDD.n4591 0.853
R9747 VDD.n4538 VDD.n4537 0.853
R9748 VDD.n4420 VDD.n4419 0.853
R9749 VDD.n4346 VDD.n4345 0.853
R9750 VDD.n4410 VDD.n4409 0.853
R9751 VDD.n3592 VDD.n3591 0.853
R9752 VDD.n3980 VDD.n3978 0.853
R9753 VDD.n2665 VDD.n2664 0.853
R9754 VDD.n4107 VDD.n4106 0.853
R9755 VDD.n4082 VDD.n4081 0.853
R9756 VDD.n3626 VDD.n3625 0.853
R9757 VDD.n3775 VDD.n3773 0.853
R9758 VDD.n3814 VDD.n3813 0.853
R9759 VDD.n3578 VDD.n3577 0.853
R9760 VDD.n3553 VDD.n3552 0.853
R9761 VDD.n3641 VDD.n2524 0.853
R9762 VDD.n937 VDD.n935 0.853
R9763 VDD.n671 VDD.n670 0.853
R9764 VDD.n492 VDD.n491 0.853
R9765 VDD.n611 VDD.n610 0.853
R9766 VDD.n636 VDD.n635 0.853
R9767 VDD.n1049 VDD.n1048 0.853
R9768 VDD.n1994 VDD.n1993 0.853
R9769 VDD.n1893 VDD.n1891 0.853
R9770 VDD.n1841 VDD.n1840 0.853
R9771 VDD.n3263 VDD.n3262 0.853
R9772 VDD.n3234 VDD.n3233 0.853
R9773 VDD.n3227 VDD.n3226 0.853
R9774 VDD.n4198 VDD.n4197 0.853
R9775 VDD.n2764 VDD.n2763 0.853
R9776 VDD.n3089 VDD.n3088 0.853
R9777 VDD.n3058 VDD.n3057 0.853
R9778 VDD.n2907 VDD.n2906 0.853
R9779 VDD.n2875 VDD.n2873 0.853
R9780 VDD.n2866 VDD.n2865 0.853
R9781 VDD.n2833 VDD.n2832 0.853
R9782 VDD.n37 VDD.n36 0.853
R9783 VDD.n135 VDD.n134 0.853
R9784 VDD.n2937 VDD.n2936 0.853
R9785 VDD.n3149 VDD.n3148 0.853
R9786 VDD.n3173 VDD.n3172 0.853
R9787 VDD.n3033 VDD.n3031 0.853
R9788 VDD.n3034 VDD.n3033 0.853
R9789 VDD.n3090 VDD.n3089 0.853
R9790 VDD.n3059 VDD.n3058 0.853
R9791 VDD.n3097 VDD.n3096 0.853
R9792 VDD.n3102 VDD.n3101 0.853
R9793 VDD.n3101 VDD.n3100 0.853
R9794 VDD.n3004 VDD.n3002 0.853
R9795 VDD.n3005 VDD.n3004 0.853
R9796 VDD.n2973 VDD.n2971 0.853
R9797 VDD.n2974 VDD.n2973 0.853
R9798 VDD.n3201 VDD.n3199 0.853
R9799 VDD.n4204 VDD.n4203 0.853
R9800 VDD.n4548 VDD.n4547 0.853
R9801 VDD.n4700 VDD.n4699 0.853
R9802 VDD.n2375 VDD.n2374 0.853
R9803 VDD.n2131 VDD.n2130 0.853
R9804 VDD.n1614 VDD.n1613 0.853
R9805 VDD.n1585 VDD.n1528 0.853
R9806 VDD.n1554 VDD.n1422 0.853
R9807 VDD.n1086 VDD.n1085 0.853
R9808 VDD.n643 VDD.n642 0.853
R9809 VDD.n580 VDD.n579 0.853
R9810 VDD.n745 VDD.n744 0.853
R9811 VDD.n928 VDD.n927 0.853
R9812 VDD.n4173 VDD.n4172 0.853
R9813 VDD.n4219 VDD.n4218 0.853
R9814 VDD.n4314 VDD.n4313 0.853
R9815 VDD.n3974 VDD.n3972 0.853
R9816 VDD.n4386 VDD.n4384 0.853
R9817 VDD.n2938 VDD.n2937 0.853
R9818 VDD.n2832 VDD.n2830 0.853
R9819 VDD.n2873 VDD.n2871 0.853
R9820 VDD.n2867 VDD.n2866 0.853
R9821 VDD.n4872 VDD.n11 0.853
R9822 VDD.n4868 VDD.n4866 0.853
R9823 VDD.n4869 VDD.n4868 0.853
R9824 VDD.n3795 VDD.n3794 0.853
R9825 VDD.n3834 VDD.n3833 0.853
R9826 VDD.n2571 VDD.n2569 0.853
R9827 VDD.n4586 VDD.n4584 0.853
R9828 VDD.n63 VDD.n61 0.853
R9829 VDD.n91 VDD.n89 0.853
R9830 VDD.n152 VDD.n150 0.853
R9831 VDD.n4833 VDD.n4831 0.853
R9832 VDD.n3312 VDD.n3311 0.853
R9833 VDD.n3398 VDD.n3397 0.853
R9834 VDD.n776 VDD.n775 0.853
R9835 VDD.n766 VDD.n585 0.853
R9836 VDD.n753 VDD.n647 0.853
R9837 VDD.n919 VDD.n918 0.853
R9838 VDD.n1196 VDD.n1194 0.853
R9839 VDD.n935 VDD.n933 0.853
R9840 VDD.n774 VDD.n492 0.853
R9841 VDD.n765 VDD.n611 0.853
R9842 VDD.n759 VDD.n636 0.853
R9843 VDD.n756 VDD.n643 0.853
R9844 VDD.n764 VDD.n615 0.853
R9845 VDD.n773 VDD.n580 0.853
R9846 VDD.n748 VDD.n745 0.853
R9847 VDD.n929 VDD.n928 0.853
R9848 VDD.n749 VDD.n671 0.853
R9849 VDD.n1192 VDD.n1190 0.853
R9850 VDD.n1193 VDD.n1192 0.853
R9851 VDD.n1085 VDD.n254 0.853
R9852 VDD.n1704 VDD.n1422 0.853
R9853 VDD.n1621 VDD.n1528 0.853
R9854 VDD.n1618 VDD.n1614 0.853
R9855 VDD.n2146 VDD.n2131 0.853
R9856 VDD.n2147 VDD.n1994 0.853
R9857 VDD.n1631 VDD.n1426 0.853
R9858 VDD.n1053 VDD.n1049 0.853
R9859 VDD.n1416 VDD.n1415 0.853
R9860 VDD.n1624 VDD.n1525 0.853
R9861 VDD.n2150 VDD.n2148 0.853
R9862 VDD.n1471 VDD.n1470 0.853
R9863 VDD.n1470 VDD.n242 0.853
R9864 VDD.n1700 VDD.n1698 0.853
R9865 VDD.n1701 VDD.n1700 0.853
R9866 VDD.n1709 VDD.n1708 0.853
R9867 VDD.n1708 VDD.n1707 0.853
R9868 VDD.n1765 VDD.n1763 0.853
R9869 VDD.n1766 VDD.n1765 0.853
R9870 VDD.n1631 VDD.n1630 0.853
R9871 VDD.n2332 VDD.n2330 0.853
R9872 VDD.n1891 VDD.n1889 0.853
R9873 VDD.n1843 VDD.n1841 0.853
R9874 VDD.n4705 VDD.n2524 0.853
R9875 VDD.n2456 VDD.n2455 0.853
R9876 VDD.n2139 VDD.n2137 0.853
R9877 VDD.n4707 VDD.n4706 0.853
R9878 VDD.n1885 VDD.n1883 0.853
R9879 VDD.n1886 VDD.n1885 0.853
R9880 VDD.n2326 VDD.n2324 0.853
R9881 VDD.n2327 VDD.n2326 0.853
R9882 VDD.n2478 VDD.n2476 0.853
R9883 VDD.n2479 VDD.n2478 0.853
R9884 VDD.n2376 VDD.n2375 0.853
R9885 VDD.n2518 VDD.n2517 0.853
R9886 VDD.n4701 VDD.n4700 0.853
R9887 VDD.n2252 VDD 0.849458
R9888 VDD.n1044 VDD.n1043 0.842605
R9889 VDD.n631 VDD.n630 0.842605
R9890 VDD.n4341 VDD.n4340 0.842605
R9891 VDD.n4533 VDD.n4532 0.842605
R9892 VDD.n4727 VDD.n4710 0.833833
R9893 VDD.n1348 VDD 0.832531
R9894 VDD VDD.n3319 0.793469
R9895 VDD.n538 VDD.n537 0.750619
R9896 VDD.n1145 VDD.n1144 0.750619
R9897 VDD.n2108 VDD.n2107 0.750619
R9898 VDD.n2496 VDD.n2495 0.750619
R9899 VDD.n2558 VDD.n2557 0.750619
R9900 VDD.n4442 VDD.n4441 0.750619
R9901 VDD.n4264 VDD.n4263 0.750619
R9902 VDD.n4415 VDD.n4414 0.685913
R9903 VDD.n2901 VDD.n2900 0.685913
R9904 VDD.n3404 VDD.n168 0.685246
R9905 VDD.n3512 VDD.n3511 0.685246
R9906 VDD.n158 VDD.n157 0.685246
R9907 VDD.n2769 VDD.n2768 0.685246
R9908 VDD.n4838 VDD.n4837 0.682731
R9909 VDD.n2722 VDD.n2721 0.682731
R9910 VDD.n3516 VDD.n3515 0.682731
R9911 VDD.n3318 VDD.n3317 0.682731
R9912 VDD.n4211 VDD.n4210 0.682731
R9913 VDD.n646 VDD.n645 0.682471
R9914 VDD.n584 VDD.n583 0.682471
R9915 VDD.n4709 VDD.n4708 0.682471
R9916 VDD.n1629 VDD.n1628 0.682471
R9917 VDD.n1425 VDD.n1424 0.682471
R9918 VDD.n3862 VDD.n3860 0.682471
R9919 VDD.n10 VDD.n9 0.682471
R9920 VDD.n3095 VDD.n3094 0.682471
R9921 VDD.n2516 VDD.n2515 0.682471
R9922 VDD.n614 VDD.n613 0.682471
R9923 VDD.n778 VDD.n777 0.682471
R9924 VDD.n1537 VDD 0.678885
R9925 VDD.n3601 VDD.n3600 0.674184
R9926 VDD.n3301 VDD.n3298 0.662569
R9927 VDD.n913 VDD.n912 0.662569
R9928 VDD.n905 VDD.n904 0.662569
R9929 VDD.n904 VDD.n903 0.662569
R9930 VDD.n238 VDD.n237 0.662569
R9931 VDD.n596 VDD.n595 0.662569
R9932 VDD.n4076 VDD.n4073 0.662569
R9933 VDD.n1808 VDD.n1805 0.662569
R9934 VDD.n129 VDD.n126 0.662569
R9935 VDD.n4565 VDD.n4562 0.662569
R9936 VDD.n4577 VDD.n4576 0.662569
R9937 VDD.n1557 VDD 0.546892
R9938 VDD.n4016 VDD.n4015 0.478112
R9939 VDD.n3928 VDD.n3927 0.478112
R9940 VDD.n3729 VDD.n3728 0.478112
R9941 VDD.n439 VDD.n438 0.478112
R9942 VDD.n973 VDD.n972 0.478112
R9943 VDD.n1777 VDD.n1776 0.478112
R9944 VDD.n1802 VDD.n1801 0.478112
R9945 VDD.n4362 VDD.n4361 0.478112
R9946 VDD.n4506 VDD.n4496 0.478112
R9947 VDD.n2040 VDD.n2030 0.478112
R9948 VDD.n1562 VDD.n1559 0.478112
R9949 VDD.n727 VDD.n720 0.478112
R9950 VDD.n4154 VDD.n4144 0.474574
R9951 VDD.n3217 VDD.n3215 0.441879
R9952 VDD.n3367 VDD.n3361 0.441879
R9953 VDD.n3445 VDD.n3444 0.441879
R9954 VDD.n3456 VDD.n3455 0.441879
R9955 VDD.n3382 VDD.n2736 0.441879
R9956 VDD.n1203 VDD.n281 0.441879
R9957 VDD.n1229 VDD.n268 0.441879
R9958 VDD.n1231 VDD.n1230 0.441879
R9959 VDD.n1242 VDD.n261 0.441879
R9960 VDD.n263 VDD.n262 0.441879
R9961 VDD.n1256 VDD.n1246 0.441879
R9962 VDD.n1248 VDD.n1247 0.441879
R9963 VDD.n1270 VDD.n1260 0.441879
R9964 VDD.n1262 VDD.n1261 0.441879
R9965 VDD.n1284 VDD.n1274 0.441879
R9966 VDD.n1276 VDD.n1275 0.441879
R9967 VDD.n1298 VDD.n1288 0.441879
R9968 VDD.n1290 VDD.n1289 0.441879
R9969 VDD.n1314 VDD.n1302 0.441879
R9970 VDD.n1306 VDD.n1305 0.441879
R9971 VDD.n1328 VDD.n1318 0.441879
R9972 VDD.n1320 VDD.n1319 0.441879
R9973 VDD.n1345 VDD.n1332 0.441879
R9974 VDD.n1337 VDD.n1336 0.441879
R9975 VDD.n1693 VDD.n1689 0.441879
R9976 VDD.n1691 VDD.n1690 0.441879
R9977 VDD.n1504 VDD.n1500 0.441879
R9978 VDD.n1445 VDD.n1444 0.441879
R9979 VDD.n228 VDD.n227 0.441879
R9980 VDD.n2288 VDD.n2287 0.441879
R9981 VDD.n2318 VDD.n2317 0.441879
R9982 VDD.n4766 VDD.n4765 0.441879
R9983 VDD.n4781 VDD.n173 0.441879
R9984 VDD.n2803 VDD.n2800 0.441879
R9985 VDD.n70 VDD.n67 0.441879
R9986 VDD.n2915 VDD.n2912 0.441879
R9987 VDD.n2620 VDD.n2617 0.441879
R9988 VDD.n2141 VDD 0.403719
R9989 VDD.n3743 VDD.n3740 0.38259
R9990 VDD.n4352 VDD.n4351 0.38259
R9991 VDD.n4641 VDD.n4640 0.38259
R9992 VDD.n4169 VDD.n4160 0.379759
R9993 VDD.n541 VDD.n540 0.332294
R9994 VDD.n1148 VDD.n1147 0.332063
R9995 VDD.n4267 VDD.n4266 0.331593
R9996 VDD.n4445 VDD.n4444 0.331593
R9997 VDD.n2561 VDD.n2560 0.331593
R9998 VDD.n2499 VDD.n2498 0.331593
R9999 VDD.n2111 VDD.n2110 0.331593
R10000 VDD VDD.n3513 0.310396
R10001 VDD.n4836 VDD 0.297375
R10002 VDD.n4369 VDD.n4368 0.287067
R10003 VDD.n4169 VDD.n4162 0.284944
R10004 VDD VDD.n779 0.277844
R10005 VDD.n536 VDD 0.259429
R10006 VDD.n1143 VDD 0.259429
R10007 VDD.n2106 VDD 0.259429
R10008 VDD.n2494 VDD 0.259429
R10009 VDD.n2556 VDD 0.259429
R10010 VDD.n4440 VDD 0.259429
R10011 VDD.n4262 VDD 0.259429
R10012 VDD.n1056 VDD.n1055 0.245153
R10013 VDD.n2142 VDD.n2141 0.245153
R10014 VDD.n4775 VDD 0.232271
R10015 VDD.n1226 VDD 0.229667
R10016 VDD.n3452 VDD 0.229667
R10017 VDD.n3369 VDD 0.229667
R10018 VDD.n3933 VDD.n3932 0.225571
R10019 VDD.n3734 VDD.n3733 0.225571
R10020 VDD.n444 VDD.n443 0.225571
R10021 VDD.n978 VDD.n977 0.225571
R10022 VDD.n4021 VDD.n4020 0.225256
R10023 VDD.n1821 VDD.n1820 0.225256
R10024 VDD.n1985 VDD.n1984 0.224793
R10025 VDD.n316 VDD.n315 0.22119
R10026 VDD.n314 VDD.n308 0.22119
R10027 VDD.n327 VDD.n308 0.22119
R10028 VDD.n310 VDD.n309 0.22119
R10029 VDD.n341 VDD.n331 0.22119
R10030 VDD.n333 VDD.n332 0.22119
R10031 VDD.n355 VDD.n345 0.22119
R10032 VDD.n347 VDD.n346 0.22119
R10033 VDD.n369 VDD.n359 0.22119
R10034 VDD.n361 VDD.n360 0.22119
R10035 VDD.n383 VDD.n373 0.22119
R10036 VDD.n375 VDD.n374 0.22119
R10037 VDD.n397 VDD.n387 0.22119
R10038 VDD.n389 VDD.n388 0.22119
R10039 VDD.n411 VDD.n403 0.22119
R10040 VDD.n305 VDD.n304 0.22119
R10041 VDD.n782 VDD.n306 0.22119
R10042 VDD.n791 VDD.n790 0.22119
R10043 VDD.n1390 VDD.n1389 0.22119
R10044 VDD.n1395 VDD.n1392 0.22119
R10045 VDD.n1483 VDD.n1482 0.22119
R10046 VDD.n1482 VDD.n1433 0.22119
R10047 VDD.n1443 VDD.n1442 0.22119
R10048 VDD.n1475 VDD.n1445 0.22119
R10049 VDD.n1475 VDD.n1474 0.22119
R10050 VDD.n1462 VDD.n1461 0.22119
R10051 VDD.n1461 VDD.n1454 0.22119
R10052 VDD.n235 VDD.n228 0.22119
R10053 VDD.n236 VDD.n235 0.22119
R10054 VDD.n2166 VDD.n2165 0.22119
R10055 VDD.n2165 VDD.n2158 0.22119
R10056 VDD.n2180 VDD.n2179 0.22119
R10057 VDD.n2179 VDD.n2172 0.22119
R10058 VDD.n2196 VDD.n2195 0.22119
R10059 VDD.n2195 VDD.n2188 0.22119
R10060 VDD.n2210 VDD.n2209 0.22119
R10061 VDD.n2209 VDD.n2202 0.22119
R10062 VDD.n2233 VDD.n2232 0.22119
R10063 VDD.n2232 VDD.n2225 0.22119
R10064 VDD.n2307 VDD.n2304 0.22119
R10065 VDD.n2307 VDD.n2306 0.22119
R10066 VDD.n2319 VDD.n208 0.22119
R10067 VDD.n2317 VDD.n2316 0.22119
R10068 VDD.n2316 VDD.n211 0.22119
R10069 VDD.n202 VDD.n201 0.22119
R10070 VDD.n201 VDD.n194 0.22119
R10071 VDD.n1859 VDD.n1858 0.22119
R10072 VDD.n1858 VDD.n1851 0.22119
R10073 VDD.n1877 VDD.n1876 0.22119
R10074 VDD.n1876 VDD.n1869 0.22119
R10075 VDD.n2393 VDD.n2392 0.22119
R10076 VDD.n2392 VDD.n2385 0.22119
R10077 VDD.n2450 VDD.n2449 0.22119
R10078 VDD.n2449 VDD.n2442 0.22119
R10079 VDD.n2441 VDD.n2440 0.22119
R10080 VDD.n2432 VDD.n2431 0.22119
R10081 VDD.n2431 VDD.n2424 0.22119
R10082 VDD.n2418 VDD.n2417 0.22119
R10083 VDD.n2417 VDD.n2410 0.22119
R10084 VDD.n3869 VDD.n3868 0.22119
R10085 VDD.n3786 VDD.n3783 0.22119
R10086 VDD.n2847 VDD.n2846 0.22119
R10087 VDD.n3028 VDD.n3027 0.22119
R10088 VDD.n3130 VDD.n2775 0.22119
R10089 VDD VDD.n1485 0.208833
R10090 VDD.n2301 VDD 0.208833
R10091 VDD.n2696 VDD.n2683 0.193208
R10092 VDD.n1989 VDD.n1988 0.191545
R10093 VDD.n1550 VDD.n1549 0.191545
R10094 VDD.n4154 VDD.n4153 0.19013
R10095 VDD.n4874 VDD 0.184386
R10096 VDD.n2920 VDD.n2919 0.133312
R10097 VDD.n432 VDD.n428 0.120292
R10098 VDD.n436 VDD.n432 0.120292
R10099 VDD.n440 VDD.n436 0.120292
R10100 VDD.n457 VDD.n453 0.120292
R10101 VDD.n461 VDD.n457 0.120292
R10102 VDD.n467 VDD.n461 0.120292
R10103 VDD.n471 VDD.n467 0.120292
R10104 VDD.n475 VDD.n471 0.120292
R10105 VDD.n949 VDD.n943 0.120292
R10106 VDD.n950 VDD.n949 0.120292
R10107 VDD.n962 VDD.n956 0.120292
R10108 VDD.n966 VDD.n962 0.120292
R10109 VDD.n970 VDD.n966 0.120292
R10110 VDD.n974 VDD.n970 0.120292
R10111 VDD.n991 VDD.n987 0.120292
R10112 VDD.n995 VDD.n991 0.120292
R10113 VDD.n1001 VDD.n995 0.120292
R10114 VDD.n1005 VDD.n1001 0.120292
R10115 VDD.n1009 VDD.n1005 0.120292
R10116 VDD.n1013 VDD.n1009 0.120292
R10117 VDD.n1017 VDD.n1013 0.120292
R10118 VDD.n1021 VDD.n1017 0.120292
R10119 VDD.n1027 VDD.n1021 0.120292
R10120 VDD.n1031 VDD.n1027 0.120292
R10121 VDD.n1035 VDD.n1031 0.120292
R10122 VDD.n1718 VDD.n1714 0.120292
R10123 VDD.n1723 VDD.n1718 0.120292
R10124 VDD.n1734 VDD.n1728 0.120292
R10125 VDD.n1735 VDD.n1734 0.120292
R10126 VDD.n1747 VDD.n1741 0.120292
R10127 VDD.n1751 VDD.n1747 0.120292
R10128 VDD.n1979 VDD.n1974 0.120292
R10129 VDD.n1974 VDD.n1970 0.120292
R10130 VDD.n1970 VDD.n1966 0.120292
R10131 VDD.n1966 VDD.n1965 0.120292
R10132 VDD.n1965 VDD.n1961 0.120292
R10133 VDD.n1961 VDD.n1957 0.120292
R10134 VDD.n1957 VDD.n1953 0.120292
R10135 VDD.n1953 VDD.n1949 0.120292
R10136 VDD.n1949 VDD.n1945 0.120292
R10137 VDD.n1945 VDD.n1939 0.120292
R10138 VDD.n1939 VDD.n1935 0.120292
R10139 VDD.n1935 VDD.n1931 0.120292
R10140 VDD.n1931 VDD.n1930 0.120292
R10141 VDD.n1930 VDD.n1926 0.120292
R10142 VDD.n1926 VDD.n1922 0.120292
R10143 VDD.n1922 VDD.n1918 0.120292
R10144 VDD.n1918 VDD.n1917 0.120292
R10145 VDD.n1917 VDD.n1913 0.120292
R10146 VDD.n1913 VDD.n1912 0.120292
R10147 VDD.n1906 VDD.n1905 0.120292
R10148 VDD.n1905 VDD.n1899 0.120292
R10149 VDD.n3651 VDD.n3647 0.120292
R10150 VDD.n3655 VDD.n3651 0.120292
R10151 VDD.n3659 VDD.n3655 0.120292
R10152 VDD.n3665 VDD.n3659 0.120292
R10153 VDD.n3669 VDD.n3665 0.120292
R10154 VDD.n3673 VDD.n3669 0.120292
R10155 VDD.n3679 VDD.n3673 0.120292
R10156 VDD.n3683 VDD.n3679 0.120292
R10157 VDD.n3687 VDD.n3683 0.120292
R10158 VDD.n3691 VDD.n3687 0.120292
R10159 VDD.n3696 VDD.n3691 0.120292
R10160 VDD.n3700 VDD.n3696 0.120292
R10161 VDD.n3702 VDD.n3700 0.120292
R10162 VDD.n3702 VDD.n3701 0.120292
R10163 VDD.n3718 VDD.n3712 0.120292
R10164 VDD.n3722 VDD.n3718 0.120292
R10165 VDD.n3726 VDD.n3722 0.120292
R10166 VDD.n3730 VDD.n3726 0.120292
R10167 VDD.n3807 VDD.n3803 0.120292
R10168 VDD.n3853 VDD.n3847 0.120292
R10169 VDD.n3857 VDD.n3853 0.120292
R10170 VDD.n3881 VDD.n3877 0.120292
R10171 VDD.n3885 VDD.n3881 0.120292
R10172 VDD.n3889 VDD.n3885 0.120292
R10173 VDD.n3894 VDD.n3889 0.120292
R10174 VDD.n3898 VDD.n3894 0.120292
R10175 VDD.n3904 VDD.n3898 0.120292
R10176 VDD.n3905 VDD.n3904 0.120292
R10177 VDD.n3917 VDD.n3911 0.120292
R10178 VDD.n3921 VDD.n3917 0.120292
R10179 VDD.n3925 VDD.n3921 0.120292
R10180 VDD.n3929 VDD.n3925 0.120292
R10181 VDD.n3946 VDD.n3942 0.120292
R10182 VDD.n3950 VDD.n3946 0.120292
R10183 VDD.n3956 VDD.n3950 0.120292
R10184 VDD.n3992 VDD.n3986 0.120292
R10185 VDD.n3993 VDD.n3992 0.120292
R10186 VDD.n4005 VDD.n3999 0.120292
R10187 VDD.n4009 VDD.n4005 0.120292
R10188 VDD.n4013 VDD.n4009 0.120292
R10189 VDD.n4017 VDD.n4013 0.120292
R10190 VDD.n4034 VDD.n4030 0.120292
R10191 VDD.n4038 VDD.n4034 0.120292
R10192 VDD.n4044 VDD.n4038 0.120292
R10193 VDD.n4048 VDD.n4044 0.120292
R10194 VDD.n4052 VDD.n4048 0.120292
R10195 VDD.n4056 VDD.n4052 0.120292
R10196 VDD.n4060 VDD.n4056 0.120292
R10197 VDD.n4064 VDD.n4060 0.120292
R10198 VDD.n4070 VDD.n4064 0.120292
R10199 VDD.n3259 VDD.n3255 0.120292
R10200 VDD.n3255 VDD.n3254 0.120292
R10201 VDD.n8 VDD.n6 0.120292
R10202 VDD.n106 VDD.n100 0.120292
R10203 VDD.n117 VDD.n113 0.120292
R10204 VDD.n75 VDD.n71 0.120292
R10205 VDD.n2823 VDD.n2819 0.120292
R10206 VDD.n2884 VDD.n2883 0.120292
R10207 VDD.n2953 VDD.n2947 0.120292
R10208 VDD.n3084 VDD.n3079 0.120292
R10209 VDD.n2786 VDD.n2782 0.120292
R10210 VDD.n3195 VDD.n3189 0.120292
R10211 VDD.n3182 VDD.n3181 0.120292
R10212 VDD.n507 VDD.n503 0.120292
R10213 VDD.n512 VDD.n507 0.120292
R10214 VDD.n516 VDD.n512 0.120292
R10215 VDD.n520 VDD.n516 0.120292
R10216 VDD.n524 VDD.n520 0.120292
R10217 VDD.n528 VDD.n524 0.120292
R10218 VDD.n555 VDD.n549 0.120292
R10219 VDD.n559 VDD.n555 0.120292
R10220 VDD.n575 VDD.n571 0.120292
R10221 VDD.n689 VDD.n685 0.120292
R10222 VDD.n1178 VDD.n1177 0.120292
R10223 VDD.n1177 VDD.n1173 0.120292
R10224 VDD.n1173 VDD.n1168 0.120292
R10225 VDD.n1168 VDD.n1164 0.120292
R10226 VDD.n1164 VDD.n1160 0.120292
R10227 VDD.n1160 VDD.n1156 0.120292
R10228 VDD.n1135 VDD.n1131 0.120292
R10229 VDD.n1131 VDD.n1125 0.120292
R10230 VDD.n1125 VDD.n1121 0.120292
R10231 VDD.n1121 VDD.n1117 0.120292
R10232 VDD.n1117 VDD.n1113 0.120292
R10233 VDD.n1113 VDD.n1109 0.120292
R10234 VDD.n1109 VDD.n1105 0.120292
R10235 VDD.n1105 VDD.n1099 0.120292
R10236 VDD.n1567 VDD.n1563 0.120292
R10237 VDD.n1578 VDD.n1572 0.120292
R10238 VDD.n1581 VDD.n1578 0.120292
R10239 VDD.n2123 VDD.n2119 0.120292
R10240 VDD.n2098 VDD.n2094 0.120292
R10241 VDD.n2094 VDD.n2088 0.120292
R10242 VDD.n2088 VDD.n2084 0.120292
R10243 VDD.n2084 VDD.n2080 0.120292
R10244 VDD.n2080 VDD.n2076 0.120292
R10245 VDD.n2076 VDD.n2072 0.120292
R10246 VDD.n2072 VDD.n2068 0.120292
R10247 VDD.n2068 VDD.n2067 0.120292
R10248 VDD.n2067 VDD.n2063 0.120292
R10249 VDD.n2063 VDD.n2059 0.120292
R10250 VDD.n2059 VDD.n2054 0.120292
R10251 VDD.n2026 VDD.n2022 0.120292
R10252 VDD.n2022 VDD.n2018 0.120292
R10253 VDD.n2018 VDD.n2012 0.120292
R10254 VDD.n2350 VDD.n2346 0.120292
R10255 VDD.n2355 VDD.n2350 0.120292
R10256 VDD.n2359 VDD.n2355 0.120292
R10257 VDD.n2363 VDD.n2359 0.120292
R10258 VDD.n2513 VDD.n2509 0.120292
R10259 VDD.n4689 VDD.n4685 0.120292
R10260 VDD.n4685 VDD.n4681 0.120292
R10261 VDD.n4681 VDD.n4677 0.120292
R10262 VDD.n4677 VDD.n4673 0.120292
R10263 VDD.n4673 VDD.n4667 0.120292
R10264 VDD.n4667 VDD.n4663 0.120292
R10265 VDD.n4663 VDD.n4659 0.120292
R10266 VDD.n4659 VDD.n4654 0.120292
R10267 VDD.n4654 VDD.n4650 0.120292
R10268 VDD.n4636 VDD.n4632 0.120292
R10269 VDD.n4632 VDD.n4628 0.120292
R10270 VDD.n4628 VDD.n4622 0.120292
R10271 VDD.n4618 VDD.n4615 0.120292
R10272 VDD.n4615 VDD.n4611 0.120292
R10273 VDD.n4611 VDD.n4606 0.120292
R10274 VDD.n2583 VDD.n2579 0.120292
R10275 VDD.n2587 VDD.n2583 0.120292
R10276 VDD.n4525 VDD.n4521 0.120292
R10277 VDD.n4521 VDD.n4517 0.120292
R10278 VDD.n4517 VDD.n4512 0.120292
R10279 VDD.n4492 VDD.n4488 0.120292
R10280 VDD.n4488 VDD.n4484 0.120292
R10281 VDD.n4484 VDD.n4478 0.120292
R10282 VDD.n4471 VDD.n4470 0.120292
R10283 VDD.n4470 VDD.n4466 0.120292
R10284 VDD.n4466 VDD.n4465 0.120292
R10285 VDD.n4465 VDD.n4461 0.120292
R10286 VDD.n4461 VDD.n4457 0.120292
R10287 VDD.n4457 VDD.n4453 0.120292
R10288 VDD.n2606 VDD.n2602 0.120292
R10289 VDD.n4328 VDD.n4324 0.120292
R10290 VDD.n4332 VDD.n4328 0.120292
R10291 VDD.n4310 VDD.n4306 0.120292
R10292 VDD.n4306 VDD.n4300 0.120292
R10293 VDD.n4293 VDD.n4292 0.120292
R10294 VDD.n4292 VDD.n4288 0.120292
R10295 VDD.n4288 VDD.n4287 0.120292
R10296 VDD.n4287 VDD.n4283 0.120292
R10297 VDD.n4283 VDD.n4279 0.120292
R10298 VDD.n4279 VDD.n4275 0.120292
R10299 VDD.n4254 VDD.n4250 0.120292
R10300 VDD.n4250 VDD.n4244 0.120292
R10301 VDD.n4244 VDD.n4240 0.120292
R10302 VDD.n4240 VDD.n4236 0.120292
R10303 VDD.n4236 VDD.n4232 0.120292
R10304 VDD.n2643 VDD.n2637 0.120292
R10305 VDD.n4130 VDD.n4124 0.120292
R10306 VDD.n4188 VDD.n4182 0.120292
R10307 VDD.n2257 VDD.n2252 0.120292
R10308 VDD.n2264 VDD.n2257 0.120292
R10309 VDD.n2269 VDD.n2264 0.120292
R10310 VDD.n2274 VDD.n2269 0.120292
R10311 VDD.n2279 VDD.n2274 0.120292
R10312 VDD.n2284 VDD.n2279 0.120292
R10313 VDD.n2286 VDD.n2284 0.120292
R10314 VDD.n4734 VDD.n4727 0.120292
R10315 VDD.n4739 VDD.n4734 0.120292
R10316 VDD.n4744 VDD.n4739 0.120292
R10317 VDD.n4749 VDD.n4744 0.120292
R10318 VDD.n4754 VDD.n4749 0.120292
R10319 VDD.n4759 VDD.n4754 0.120292
R10320 VDD.n4760 VDD.n4759 0.120292
R10321 VDD.n4774 VDD.n4760 0.120292
R10322 VDD.n4786 VDD.n4782 0.120292
R10323 VDD.n4790 VDD.n4786 0.120292
R10324 VDD.n4799 VDD.n4795 0.120292
R10325 VDD.n3418 VDD.n3412 0.120292
R10326 VDD.n3422 VDD.n3418 0.120292
R10327 VDD.n3426 VDD.n3422 0.120292
R10328 VDD.n3430 VDD.n3426 0.120292
R10329 VDD.n3434 VDD.n3430 0.120292
R10330 VDD.n3438 VDD.n3434 0.120292
R10331 VDD.n3439 VDD.n3438 0.120292
R10332 VDD.n3451 VDD.n3439 0.120292
R10333 VDD.n3464 VDD.n3400 0.120292
R10334 VDD.n3469 VDD.n3464 0.120292
R10335 VDD.n3474 VDD.n3469 0.120292
R10336 VDD.n3479 VDD.n3474 0.120292
R10337 VDD.n3484 VDD.n3479 0.120292
R10338 VDD.n3491 VDD.n3484 0.120292
R10339 VDD.n3508 VDD.n3491 0.120292
R10340 VDD.n2714 VDD.n2710 0.120292
R10341 VDD.n3387 VDD.n3383 0.120292
R10342 VDD.n3383 VDD.n2734 0.120292
R10343 VDD.n3368 VDD.n3359 0.120292
R10344 VDD.n3359 VDD.n3357 0.120292
R10345 VDD.n3357 VDD.n3352 0.120292
R10346 VDD.n3352 VDD.n3347 0.120292
R10347 VDD.n3347 VDD.n3342 0.120292
R10348 VDD.n3342 VDD.n3335 0.120292
R10349 VDD.n3335 VDD.n3330 0.120292
R10350 VDD.n3292 VDD.n3288 0.120292
R10351 VDD.n3296 VDD.n3292 0.120292
R10352 VDD.n453 VDD.n448 0.11899
R10353 VDD.n987 VDD.n982 0.11899
R10354 VDD.n3782 VDD.n3781 0.11899
R10355 VDD.n3877 VDD.n3871 0.11899
R10356 VDD.n3942 VDD.n3937 0.11899
R10357 VDD.n4030 VDD.n4025 0.11899
R10358 VDD.n2027 VDD.n2026 0.11899
R10359 VDD.n4493 VDD.n4492 0.11899
R10360 VDD.n2919 VDD.n2917 0.117688
R10361 VDD.n1056 VDD 0.117476
R10362 VDD.n1804 VDD.n1803 0.116385
R10363 VDD.n123 VDD.n122 0.116385
R10364 VDD.n4571 VDD.n4567 0.116385
R10365 VDD.n3297 VDD.n3296 0.116385
R10366 VDD.n4690 VDD.n4689 0.115083
R10367 VDD.n3739 VDD.n3738 0.113781
R10368 VDD.n2364 VDD.n2363 0.113781
R10369 VDD.n593 VDD.n592 0.112479
R10370 VDD.n3957 VDD.n3956 0.112479
R10371 VDD.n3117 VDD.n3113 0.112479
R10372 VDD.n4572 VDD.n4571 0.112479
R10373 VDD.n4526 VDD.n4525 0.112479
R10374 VDD.n4821 VDD.n4820 0.112479
R10375 VDD.n3827 VDD.n3823 0.111177
R10376 VDD.n529 VDD.n528 0.111177
R10377 VDD.n560 VDD.n559 0.111177
R10378 VDD.n1156 VDD.n1152 0.111177
R10379 VDD.n2119 VDD.n2115 0.111177
R10380 VDD.n2487 VDD.n2486 0.111177
R10381 VDD.n4453 VDD.n4449 0.111177
R10382 VDD.n4275 VDD.n4271 0.111177
R10383 VDD.n2697 VDD.n2696 0.111177
R10384 VDD.n476 VDD.n475 0.109875
R10385 VDD.n3847 VDD.n3843 0.108573
R10386 VDD.n3567 VDD.n3566 0.108573
R10387 VDD.n4800 VDD.n4799 0.108573
R10388 VDD.n2849 VDD.n2848 0.107271
R10389 VDD.n549 VDD.n545 0.107271
R10390 VDD.n1136 VDD.n1135 0.107271
R10391 VDD.n2099 VDD.n2098 0.107271
R10392 VDD.n4433 VDD.n4432 0.107271
R10393 VDD.n4255 VDD.n4254 0.107271
R10394 VDD.n3543 VDD.n3542 0.105969
R10395 VDD.n2925 VDD.n2924 0.105969
R10396 VDD.n1099 VDD.n1095 0.105969
R10397 VDD.n1598 VDD.n1597 0.104667
R10398 VDD.n2961 VDD.n2960 0.102062
R10399 VDD.n3020 VDD.n3019 0.102062
R10400 VDD.n717 VDD.n716 0.102062
R10401 VDD.n3388 VDD.n3387 0.102062
R10402 VDD.n661 VDD.n660 0.10076
R10403 VDD.n1980 VDD.n1979 0.10076
R10404 VDD.n2992 VDD.n2991 0.10076
R10405 VDD.n4141 VDD.n4140 0.10076
R10406 VDD.n441 VDD.n440 0.0994583
R10407 VDD.n975 VDD.n974 0.0994583
R10408 VDD.n3731 VDD.n3730 0.0994583
R10409 VDD.n3930 VDD.n3929 0.0994583
R10410 VDD.n3613 VDD.n3609 0.0994583
R10411 VDD.n4018 VDD.n4017 0.0994583
R10412 VDD.n3132 VDD.n3131 0.0994583
R10413 VDD.n4606 VDD.n4602 0.0994583
R10414 VDD.n4512 VDD.n4508 0.0994583
R10415 VDD.n4232 VDD.n4228 0.0994583
R10416 VDD.n4092 VDD.n4091 0.0981562
R10417 VDD.n503 VDD 0.0981562
R10418 VDD VDD.n1178 0.0981562
R10419 VDD.n1597 VDD 0.0981562
R10420 VDD.n2346 VDD 0.0981562
R10421 VDD.n4637 VDD.n4636 0.0981562
R10422 VDD VDD.n4618 0.0981562
R10423 VDD VDD.n4471 0.0981562
R10424 VDD VDD.n4293 0.0981562
R10425 VDD.n330 VDD.n329 0.0981562
R10426 VDD.n344 VDD.n343 0.0981562
R10427 VDD.n358 VDD.n357 0.0981562
R10428 VDD.n372 VDD.n371 0.0981562
R10429 VDD.n386 VDD.n385 0.0981562
R10430 VDD.n400 VDD.n399 0.0981562
R10431 VDD.n414 VDD.n413 0.0981562
R10432 VDD.n823 VDD.n822 0.0981562
R10433 VDD.n854 VDD.n853 0.0981562
R10434 VDD.n868 VDD.n867 0.0981562
R10435 VDD.n897 VDD.n896 0.0981562
R10436 VDD.n1245 VDD.n1244 0.0981562
R10437 VDD.n1259 VDD.n1258 0.0981562
R10438 VDD.n1273 VDD.n1272 0.0981562
R10439 VDD.n1287 VDD.n1286 0.0981562
R10440 VDD.n1301 VDD.n1300 0.0981562
R10441 VDD.n1317 VDD.n1316 0.0981562
R10442 VDD.n1331 VDD.n1330 0.0981562
R10443 VDD.n1377 VDD.n1376 0.0981562
R10444 VDD.n1398 VDD.n1397 0.0981562
R10445 VDD.n1649 VDD.n1648 0.0981562
R10446 VDD.n2169 VDD.n2168 0.0981562
R10447 VDD.n2183 VDD.n2182 0.0981562
R10448 VDD.n2199 VDD.n2198 0.0981562
R10449 VDD.n2213 VDD.n2212 0.0981562
R10450 VDD.n2421 VDD.n2420 0.0981562
R10451 VDD.n53 VDD.n52 0.0968542
R10452 VDD.n4432 VDD.n4428 0.0968542
R10453 VDD.n4397 VDD.n4396 0.0968542
R10454 VDD.n205 VDD.n204 0.0968542
R10455 VDD.n4782 VDD 0.0968542
R10456 VDD VDD.n3400 0.0968542
R10457 VDD VDD.n3368 0.0968542
R10458 VDD.n4023 VDD.n4022 0.0960224
R10459 VDD.n3935 VDD.n3934 0.0960224
R10460 VDD.n3736 VDD.n3735 0.0960224
R10461 VDD.n446 VDD.n445 0.0960224
R10462 VDD.n980 VDD.n979 0.0960224
R10463 VDD.n1988 VDD.n1987 0.0960224
R10464 VDD.n1823 VDD.n1822 0.0960224
R10465 VDD.n4359 VDD.n4352 0.0960224
R10466 VDD.n4376 VDD.n4369 0.0960224
R10467 VDD.n4378 VDD.n4376 0.0960224
R10468 VDD.n4506 VDD.n4505 0.0960224
R10469 VDD.n4505 VDD.n4498 0.0960224
R10470 VDD.n4649 VDD.n4641 0.0960224
R10471 VDD.n2053 VDD.n2045 0.0960224
R10472 VDD.n2040 VDD.n2039 0.0960224
R10473 VDD.n2039 VDD.n2032 0.0960224
R10474 VDD.n1543 VDD.n1542 0.0960224
R10475 VDD.n1548 VDD.n1543 0.0960224
R10476 VDD.n741 VDD.n733 0.0960224
R10477 VDD.n727 VDD.n726 0.0960224
R10478 VDD.n701 VDD.n696 0.0955521
R10479 VDD VDD.n307 0.0955521
R10480 VDD.n1678 VDD.n1677 0.0955521
R10481 VDD.n4153 VDD.n4146 0.0953148
R10482 VDD.n1831 VDD.n1830 0.09425
R10483 VDD.n3614 VDD.n3613 0.09425
R10484 VDD VDD.n259 0.09425
R10485 VDD.n702 VDD.n701 0.0929479
R10486 VDD.n2124 VDD.n2123 0.0929479
R10487 VDD.n3216 VDD.n3213 0.0929479
R10488 VDD.n2004 VDD.n2003 0.0916458
R10489 VDD.n3623 VDD.n3622 0.0903438
R10490 VDD.n1826 VDD.n1825 0.0890417
R10491 VDD.n690 VDD.n689 0.0890417
R10492 VDD.n2473 VDD.n2472 0.0877396
R10493 VDD.n46 VDD.n45 0.0877396
R10494 VDD.n2607 VDD.n2606 0.0877396
R10495 VDD.n4407 VDD.n4406 0.0877396
R10496 VDD.n249 VDD.n248 0.0864375
R10497 VDD.n4103 VDD.n4102 0.0864375
R10498 VDD.n3281 VDD.n3280 0.0864375
R10499 VDD.n3542 VDD.n3538 0.0851354
R10500 VDD.n3145 VDD.n3144 0.0851354
R10501 VDD.n2540 VDD.n2539 0.0851354
R10502 VDD.n2644 VDD.n2643 0.0851354
R10503 VDD.n2396 VDD.n2395 0.0851354
R10504 VDD.n656 VDD.n655 0.0838333
R10505 VDD.n1779 VDD.n1778 0.0838333
R10506 VDD.n3647 VDD.n3643 0.0838333
R10507 VDD.n2661 VDD.n2660 0.0838333
R10508 VDD.n2824 VDD.n2823 0.0838333
R10509 VDD.n2985 VDD.n2984 0.0838333
R10510 VDD.n3118 VDD.n3117 0.0838333
R10511 VDD.n2954 VDD.n2953 0.0825312
R10512 VDD.n3015 VDD.n3014 0.0825312
R10513 VDD.n4131 VDD.n4130 0.0825312
R10514 VDD.n4157 VDD.n4156 0.0825312
R10515 VDD.n2733 VDD.n2732 0.0825312
R10516 VDD.n2940 VDD.n2939 0.0818688
R10517 VDD.n3054 VDD.n3053 0.0812292
R10518 VDD.n3196 VDD.n3195 0.0812292
R10519 VDD.n707 VDD.n706 0.0812292
R10520 VDD.n1067 VDD.n1066 0.0812292
R10521 VDD.n4182 VDD.n4178 0.0812292
R10522 VDD.n1611 VDD.n1610 0.0799271
R10523 VDD.n3536 VDD.n3535 0.078625
R10524 VDD.n2892 VDD.n2891 0.078625
R10525 VDD.n1080 VDD.n1079 0.078625
R10526 VDD.n2862 VDD.n2861 0.0773229
R10527 VDD.n2043 VDD.n2042 0.0773229
R10528 VDD.n2286 VDD.n2285 0.0773229
R10529 VDD.n2435 VDD.n2434 0.0773229
R10530 VDD.n3828 VDD.n3827 0.0760208
R10531 VDD.n3562 VDD.n3561 0.0760208
R10532 VDD.n24 VDD.n23 0.0760208
R10533 VDD.n1447 VDD 0.0760208
R10534 VDD.n4791 VDD.n4790 0.0760208
R10535 VDD.n488 VDD.n487 0.0747188
R10536 VDD.n4333 VDD.n4332 0.0747188
R10537 VDD.n4189 VDD.n4188 0.0747188
R10538 VDD.n536 VDD.n535 0.0738696
R10539 VDD.n1143 VDD.n1142 0.0738696
R10540 VDD.n2106 VDD.n2105 0.0738696
R10541 VDD.n2494 VDD.n2493 0.0738696
R10542 VDD.n2556 VDD.n2555 0.0738696
R10543 VDD.n4440 VDD.n4439 0.0738696
R10544 VDD.n4262 VDD.n4261 0.0738696
R10545 VDD.n1036 VDD.n1035 0.0734167
R10546 VDD.n3808 VDD.n3807 0.0734167
R10547 VDD.n576 VDD.n575 0.0734167
R10548 VDD.n3412 VDD.n3405 0.0734167
R10549 VDD.n2715 VDD.n2714 0.0734167
R10550 VDD.n607 VDD.n606 0.0721146
R10551 VDD.n3969 VDD.n3968 0.0721146
R10552 VDD.n3260 VDD.n3259 0.0721146
R10553 VDD.n2787 VDD.n2786 0.0721146
R10554 VDD.n3181 VDD.n3175 0.0721146
R10555 VDD.n4557 VDD.n4556 0.0721146
R10556 VDD.n2588 VDD.n2587 0.0721146
R10557 VDD.n1201 VDD.n1200 0.0721146
R10558 VDD.n1752 VDD.n1751 0.0708125
R10559 VDD.n76 VDD.n75 0.0708125
R10560 VDD.n730 VDD.n729 0.0708125
R10561 VDD.n1862 VDD.n1861 0.0708125
R10562 VDD.n943 VDD.n939 0.0695104
R10563 VDD.n3781 VDD.n3777 0.0695104
R10564 VDD.n3986 VDD.n3982 0.0695104
R10565 VDD.n4863 VDD.n4862 0.0695104
R10566 VDD.n3085 VDD.n3084 0.0695104
R10567 VDD.n4381 VDD.n4380 0.0695104
R10568 VDD.n1502 VDD.n1430 0.0695104
R10569 VDD.n2142 VDD 0.0686608
R10570 VDD.n623 VDD.n622 0.0682083
R10571 VDD.n1899 VDD.n1895 0.0682083
R10572 VDD.n4071 VDD.n4070 0.0682083
R10573 VDD.n118 VDD.n117 0.0682083
R10574 VDD.n3309 VDD.n3308 0.0682083
R10575 VDD.n2883 VDD.n2877 0.0669062
R10576 VDD.n4311 VDD.n4310 0.0669062
R10577 VDD.n1663 VDD.n1662 0.0669062
R10578 VDD.n3803 VDD.n3797 0.0656042
R10579 VDD.n3863 VDD.n3857 0.0656042
R10580 VDD.n2566 VDD.n2565 0.0656042
R10581 VDD.n107 VDD.n106 0.0643021
R10582 VDD.n679 VDD.n678 0.0643021
R10583 VDD.n1412 VDD.n1411 0.063
R10584 VDD.n1465 VDD.n1464 0.063
R10585 VDD.n956 VDD 0.0603958
R10586 VDD.n1724 VDD.n1723 0.0603958
R10587 VDD.n1728 VDD.n1724 0.0603958
R10588 VDD.n1741 VDD 0.0603958
R10589 VDD.n1906 VDD 0.0603958
R10590 VDD.n3712 VDD 0.0603958
R10591 VDD.n3911 VDD 0.0603958
R10592 VDD.n3999 VDD 0.0603958
R10593 VDD.n2848 VDD 0.0603958
R10594 VDD.n2891 VDD 0.0603958
R10595 VDD.n3131 VDD 0.0603958
R10596 VDD.n3182 VDD 0.0603958
R10597 VDD.n1179 VDD 0.0603958
R10598 VDD.n1568 VDD.n1567 0.0603958
R10599 VDD.n1572 VDD.n1568 0.0603958
R10600 VDD VDD.n1581 0.0603958
R10601 VDD.n2012 VDD 0.0603958
R10602 VDD.n4622 VDD 0.0603958
R10603 VDD.n4619 VDD 0.0603958
R10604 VDD.n4478 VDD 0.0603958
R10605 VDD.n4472 VDD 0.0603958
R10606 VDD.n2602 VDD.n2598 0.0603958
R10607 VDD.n4300 VDD 0.0603958
R10608 VDD.n4294 VDD 0.0603958
R10609 VDD.n882 VDD.n881 0.0603958
R10610 VDD.n3330 VDD 0.0603958
R10611 VDD.n3079 VDD.n3075 0.0590938
R10612 VDD VDD.n2235 0.0590938
R10613 VDD.n2398 VDD 0.0590938
R10614 VDD.n4192 VDD 0.0578029
R10615 VDD.n3514 VDD.n3508 0.0577917
R10616 VDD.n113 VDD.n107 0.0564896
R10617 VDD.n3189 VDD.n3160 0.0564896
R10618 VDD.n685 VDD.n679 0.0564896
R10619 VDD.n2514 VDD.n2513 0.0564896
R10620 VDD.n2637 VDD.n2633 0.0564896
R10621 VDD.n3319 VDD.n2756 0.0564896
R10622 VDD.n3165 VDD 0.0525833
R10623 VDD.n1557 VDD.n1556 0.0520464
R10624 VDD.n2514 VDD.n2503 0.0512812
R10625 VDD.n838 VDD.n837 0.0499792
R10626 VDD.n837 VDD.n836 0.0486771
R10627 VDD.n2155 VDD.n2154 0.0460729
R10628 VDD.n3862 VDD.n3861 0.0444189
R10629 VDD VDD.n1068 0.0434688
R10630 VDD VDD.n190 0.0434688
R10631 VDD.n3795 VDD.n3790 0.0427297
R10632 VDD.n3207 VDD.n3206 0.0423356
R10633 VDD.n532 VDD.n530 0.0412609
R10634 VDD.n1139 VDD.n1137 0.0412609
R10635 VDD.n2102 VDD.n2100 0.0412609
R10636 VDD.n2490 VDD.n2488 0.0412609
R10637 VDD.n2552 VDD.n2550 0.0412609
R10638 VDD.n4436 VDD.n4434 0.0412609
R10639 VDD.n4258 VDD.n4256 0.0412609
R10640 VDD.n2152 VDD.n240 0.0410405
R10641 VDD.n917 VDD.n916 0.0410405
R10642 VDD.n2324 VDD.n2323 0.0410405
R10643 VDD.n1893 VDD.n1892 0.0410405
R10644 VDD.n134 VDD.n96 0.0410405
R10645 VDD.n1554 VDD.n1552 0.0410405
R10646 VDD VDD.n1347 0.0408646
R10647 VDD.n780 VDD 0.0395625
R10648 VDD.n4081 VDD.n2670 0.0393514
R10649 VDD.n635 VDD.n634 0.0393514
R10650 VDD.n3311 VDD.n3275 0.0393514
R10651 VDD.n2907 VDD.n2894 0.0393514
R10652 VDD.n2875 VDD.n2807 0.0393514
R10653 VDD.n4313 VDD.n2614 0.0393514
R10654 VDD.n532 VDD 0.0385435
R10655 VDD.n1139 VDD 0.0385435
R10656 VDD.n2102 VDD 0.0385435
R10657 VDD.n2490 VDD 0.0385435
R10658 VDD.n2552 VDD 0.0385435
R10659 VDD.n4436 VDD 0.0385435
R10660 VDD.n4258 VDD 0.0385435
R10661 VDD.n937 VDD.n297 0.0376622
R10662 VDD.n89 VDD.n88 0.0376622
R10663 VDD.n4866 VDD.n4848 0.0376622
R10664 VDD.n4547 VDD.n4545 0.0376622
R10665 VDD.n4699 VDD.n2528 0.0376622
R10666 VDD.n744 VDD.n743 0.0376622
R10667 VDD.n2870 VDD.n2795 0.036925
R10668 VDD.n1883 VDD.n1882 0.035973
R10669 VDD.n2334 VDD.n2333 0.035973
R10670 VDD.n4584 VDD.n4583 0.035973
R10671 VDD.n4537 VDD.n4536 0.035973
R10672 VDD.n3980 VDD.n2679 0.035973
R10673 VDD.n3775 VDD.n3748 0.035973
R10674 VDD.n1763 VDD.n1762 0.035973
R10675 VDD.n3212 VDD.n3211 0.035973
R10676 VDD.n3226 VDD.n3225 0.035973
R10677 VDD.n3088 VDD.n3064 0.035973
R10678 VDD.n3102 VDD.n2789 0.035973
R10679 VDD.n2374 VDD.n178 0.035973
R10680 VDD.n1999 VDD.n1998 0.035973
R10681 VDD.n1585 VDD.n1584 0.035973
R10682 VDD.n744 VDD.n674 0.035973
R10683 VDD.n2940 VDD.n2794 0.0358009
R10684 VDD.n4845 VDD.n4844 0.0356652
R10685 VDD.n3865 VDD.n3863 0.0343542
R10686 VDD.n4384 VDD.n4348 0.0342838
R10687 VDD.n3597 VDD.n3596 0.0342838
R10688 VDD.n3625 VDD.n3598 0.0342838
R10689 VDD.n3814 VDD.n3810 0.0342838
R10690 VDD.n3972 VDD.n3629 0.0342838
R10691 VDD.n1840 VDD.n1817 0.0342838
R10692 VDD.n1839 VDD.n1838 0.0342838
R10693 VDD.n3262 VDD.n3237 0.0342838
R10694 VDD.n3173 VDD.n3170 0.0342838
R10695 VDD.n2130 VDD.n1997 0.0342838
R10696 VDD.n3796 VDD.n3789 0.0330521
R10697 VDD.n1698 VDD.n1697 0.0325946
R10698 VDD.n4420 VDD.n2610 0.0325946
R10699 VDD.n4409 VDD.n4392 0.0325946
R10700 VDD.n610 VDD.n588 0.0325946
R10701 VDD.n1048 VDD.n1047 0.0325946
R10702 VDD.n641 VDD.n640 0.0325946
R10703 VDD.n579 VDD.n495 0.0325946
R10704 VDD.n4833 VDD.n4829 0.0325946
R10705 VDD.n2976 VDD.n2975 0.0323719
R10706 VDD.n3007 VDD.n3006 0.0319313
R10707 VDD.n4871 VDD.n4870 0.0317844
R10708 VDD.n1894 VDD.n1811 0.03175
R10709 VDD.n133 VDD.n132 0.03175
R10710 VDD.n915 VDD.n914 0.03175
R10711 VDD.n2153 VDD.n239 0.03175
R10712 VDD.n3224 VDD 0.03175
R10713 VDD.n1555 VDD.n1551 0.0314278
R10714 VDD.n2718 VDD.n2682 0.0309054
R10715 VDD.n2569 VDD.n2543 0.0309054
R10716 VDD.n2609 VDD.n2608 0.0309054
R10717 VDD.n4345 VDD.n4344 0.0309054
R10718 VDD.n4391 VDD.n4390 0.0309054
R10719 VDD.n4106 VDD.n4105 0.0309054
R10720 VDD.n3577 VDD.n3576 0.0309054
R10721 VDD.n2461 VDD.n2460 0.0309054
R10722 VDD.n2476 VDD.n2475 0.0309054
R10723 VDD.n4197 VDD.n4196 0.0309054
R10724 VDD.n61 VDD.n40 0.0309054
R10725 VDD.n60 VDD.n59 0.0309054
R10726 VDD.n642 VDD.n639 0.0309054
R10727 VDD.n633 VDD.n632 0.0304479
R10728 VDD.n4080 VDD.n4079 0.0304479
R10729 VDD.n2876 VDD.n2806 0.0304479
R10730 VDD.n2910 VDD.n2908 0.0304479
R10731 VDD.n4312 VDD.n2623 0.0304479
R10732 VDD.n2322 VDD.n2321 0.0304479
R10733 VDD.n3310 VDD.n3304 0.0304479
R10734 VDD.n3607 VDD.n3604 0.0301109
R10735 VDD.n1524 VDD.n1523 0.0292162
R10736 VDD.n4810 VDD.n4809 0.0292162
R10737 VDD.n4593 VDD.n4592 0.0292162
R10738 VDD.n4087 VDD.n4086 0.0292162
R10739 VDD.n3834 VDD.n3830 0.0292162
R10740 VDD.n491 VDD.n420 0.0292162
R10741 VDD.n1709 VDD.n250 0.0292162
R10742 VDD.n3233 VDD.n3231 0.0292162
R10743 VDD.n36 VDD.n19 0.0292162
R10744 VDD.n3148 VDD.n3147 0.0292162
R10745 VDD.n938 VDD.n296 0.0291458
R10746 VDD.n4864 VDD.n4856 0.0291458
R10747 VDD.n87 VDD.n86 0.0291458
R10748 VDD.n4698 VDD.n4697 0.0291458
R10749 VDD.n4561 VDD.n4559 0.0291458
R10750 VDD.n1761 VDD.n1760 0.0278438
R10751 VDD.n3776 VDD.n3747 0.0278438
R10752 VDD.n3981 VDD.n2678 0.0278438
R10753 VDD.n3086 VDD.n3074 0.0278438
R10754 VDD.n3105 VDD.n3103 0.0278438
R10755 VDD.n742 VDD.n702 0.0278438
R10756 VDD.n1588 VDD.n1586 0.0278438
R10757 VDD.n2128 VDD.n2124 0.0278438
R10758 VDD.n2337 VDD.n2335 0.0278438
R10759 VDD.n2373 VDD.n2371 0.0278438
R10760 VDD.n4582 VDD.n4581 0.0278438
R10761 VDD.n4535 VDD.n4534 0.0278438
R10762 VDD.n3222 VDD.n3213 0.0278438
R10763 VDD.n2828 VDD.n12 0.0278187
R10764 VDD.n2136 VDD.n2135 0.027527
R10765 VDD.n1414 VDD.n257 0.027527
R10766 VDD.n2454 VDD.n2381 0.027527
R10767 VDD.n4219 VDD.n2646 0.027527
R10768 VDD.n3591 VDD.n3589 0.027527
R10769 VDD.n3552 VDD.n3529 0.027527
R10770 VDD.n2936 VDD.n2935 0.027527
R10771 VDD.n1837 VDD.n1826 0.0265417
R10772 VDD.n1836 VDD.n1831 0.0265417
R10773 VDD.n3817 VDD.n3815 0.0265417
R10774 VDD.n3970 VDD.n3964 0.0265417
R10775 VDD.n3618 VDD.n3614 0.0265417
R10776 VDD.n3624 VDD.n3623 0.0265417
R10777 VDD.n3261 VDD.n3246 0.0265417
R10778 VDD.n3174 VDD.n3168 0.0265417
R10779 VDD.n2129 VDD.n2004 0.0265417
R10780 VDD.n1471 VDD.n1467 0.0258378
R10781 VDD.n2664 VDD.n2663 0.0258378
R10782 VDD.n3641 VDD.n3640 0.0258378
R10783 VDD.n1993 VDD.n1774 0.0258378
R10784 VDD.n2865 VDD.n2812 0.0258378
R10785 VDD.n2833 VDD.n2825 0.0258378
R10786 VDD.n4114 VDD.n4113 0.0254412
R10787 VDD.n3270 VDD.n3269 0.0253211
R10788 VDD.n608 VDD.n602 0.0252396
R10789 VDD.n1046 VDD.n1045 0.0252396
R10790 VDD.n577 VDD.n567 0.0252396
R10791 VDD.n696 VDD.n695 0.0252396
R10792 VDD.n4421 VDD.n2607 0.0252396
R10793 VDD.n4408 VDD.n4407 0.0252396
R10794 VDD.n4834 VDD.n4828 0.0252396
R10795 VDD.n1198 VDD.n1197 0.0241486
R10796 VDD.n3397 VDD.n2727 0.0241486
R10797 VDD.n4172 VDD.n4119 0.0241486
R10798 VDD.n670 VDD.n650 0.0241486
R10799 VDD.n2763 VDD.n2761 0.0241486
R10800 VDD.n3002 VDD.n2978 0.0241486
R10801 VDD.n2971 VDD.n2943 0.0241486
R10802 VDD.n3199 VDD.n3198 0.0241486
R10803 VDD.n4203 VDD.n4202 0.0241486
R10804 VDD.n1086 VDD.n1081 0.0241486
R10805 VDD.n927 VDD.n926 0.0241486
R10806 VDD.n1190 VDD.n1189 0.0241486
R10807 VDD.n2466 VDD.n2462 0.0239375
R10808 VDD.n2474 VDD.n2473 0.0239375
R10809 VDD.n3575 VDD.n3574 0.0239375
R10810 VDD.n4104 VDD.n4103 0.0239375
R10811 VDD.n58 VDD.n46 0.0239375
R10812 VDD.n57 VDD.n53 0.0239375
R10813 VDD.n691 VDD.n690 0.0239375
R10814 VDD.n2567 VDD.n2548 0.0239375
R10815 VDD.n4428 VDD.n4427 0.0239375
R10816 VDD.n4343 VDD.n4342 0.0239375
R10817 VDD.n4401 VDD.n4397 0.0239375
R10818 VDD.n4195 VDD.n4194 0.0239375
R10819 VDD.n4775 VDD 0.0239375
R10820 VDD.n3452 VDD 0.0239375
R10821 VDD.n2716 VDD.n2706 0.0239375
R10822 VDD.n3369 VDD 0.0239375
R10823 VDD.n2829 VDD.n2809 0.0238531
R10824 VDD.n3036 VDD.n3035 0.0235594
R10825 VDD.n489 VDD.n483 0.0226354
R10826 VDD.n950 VDD 0.0226354
R10827 VDD.n1710 VDD.n249 0.0226354
R10828 VDD.n1735 VDD 0.0226354
R10829 VDD.n1912 VDD 0.0226354
R10830 VDD.n3701 VDD 0.0226354
R10831 VDD.n3837 VDD.n3835 0.0226354
R10832 VDD.n3905 VDD 0.0226354
R10833 VDD.n3993 VDD 0.0226354
R10834 VDD.n4098 VDD.n4092 0.0226354
R10835 VDD.n3254 VDD 0.0226354
R10836 VDD.n35 VDD.n34 0.0226354
R10837 VDD.n2924 VDD 0.0226354
R10838 VDD.n3146 VDD.n3145 0.0226354
R10839 VDD.n742 VDD.n731 0.0226354
R10840 VDD.n1179 VDD 0.0226354
R10841 VDD.n2054 VDD.n2043 0.0226354
R10842 VDD.n4650 VDD.n4637 0.0226354
R10843 VDD.n4619 VDD 0.0226354
R10844 VDD.n4594 VDD.n2540 0.0226354
R10845 VDD.n4472 VDD 0.0226354
R10846 VDD.n4294 VDD 0.0226354
R10847 VDD.n1696 VDD.n1695 0.0226354
R10848 VDD VDD.n1431 0.0226354
R10849 VDD.n2302 VDD 0.0226354
R10850 VDD.n4808 VDD.n4807 0.0226354
R10851 VDD.n3282 VDD.n3281 0.0226354
R10852 VDD.n3057 VDD.n3039 0.0224595
R10853 VDD.n3057 VDD.n3056 0.0224595
R10854 VDD.n150 VDD.n138 0.0224595
R10855 VDD.n150 VDD.n149 0.0224595
R10856 VDD.n3031 VDD.n3009 0.0224595
R10857 VDD.n3031 VDD.n3010 0.0224595
R10858 VDD.n1613 VDD.n1531 0.0224595
R10859 VDD.n1613 VDD.n1532 0.0224595
R10860 VDD.n3522 VDD.n3521 0.0216602
R10861 VDD.n3752 VDD.n3751 0.0216602
R10862 VDD.n3583 VDD.n3582 0.0214906
R10863 VDD.n3762 VDD.n3761 0.0214228
R10864 VDD.n447 VDD.n441 0.0213333
R10865 VDD.n981 VDD.n975 0.0213333
R10866 VDD.n1824 VDD.n1818 0.0213333
R10867 VDD.n3737 VDD.n3731 0.0213333
R10868 VDD.n3789 VDD.n3787 0.0213333
R10869 VDD.n3870 VDD.n3865 0.0213333
R10870 VDD.n3936 VDD.n3930 0.0213333
R10871 VDD.n3551 VDD.n3550 0.0213333
R10872 VDD.n3538 VDD.n3537 0.0213333
R10873 VDD.n3609 VDD.n3608 0.0213333
R10874 VDD.n4024 VDD.n4018 0.0213333
R10875 VDD.n2884 VDD 0.0213333
R10876 VDD.n2934 VDD.n2933 0.0213333
R10877 VDD.n3136 VDD.n3132 0.0213333
R10878 VDD.n729 VDD.n728 0.0213333
R10879 VDD.n2042 VDD.n2041 0.0213333
R10880 VDD.n4602 VDD.n4601 0.0213333
R10881 VDD.n4508 VDD.n4507 0.0213333
R10882 VDD.n4379 VDD.n4365 0.0213333
R10883 VDD.n4228 VDD.n4227 0.0213333
R10884 VDD.n4220 VDD.n2644 0.0213333
R10885 VDD.n329 VDD.n328 0.0213333
R10886 VDD.n343 VDD.n342 0.0213333
R10887 VDD.n357 VDD.n356 0.0213333
R10888 VDD.n371 VDD.n370 0.0213333
R10889 VDD.n385 VDD.n384 0.0213333
R10890 VDD.n399 VDD.n398 0.0213333
R10891 VDD.n413 VDD.n412 0.0213333
R10892 VDD.n781 VDD.n780 0.0213333
R10893 VDD.n1413 VDD.n1396 0.0213333
R10894 VDD.n1485 VDD.n1484 0.0213333
R10895 VDD.n1464 VDD.n1463 0.0213333
R10896 VDD.n2167 VDD.n2155 0.0213333
R10897 VDD.n2181 VDD.n2169 0.0213333
R10898 VDD.n2197 VDD.n2183 0.0213333
R10899 VDD.n2211 VDD.n2199 0.0213333
R10900 VDD.n2234 VDD.n2213 0.0213333
R10901 VDD.n2298 VDD.n217 0.0213333
R10902 VDD.n2303 VDD.n2301 0.0213333
R10903 VDD.n204 VDD.n203 0.0213333
R10904 VDD.n1860 VDD.n1848 0.0213333
R10905 VDD.n1881 VDD.n1880 0.0213333
R10906 VDD.n2394 VDD.n2382 0.0213333
R10907 VDD.n2436 VDD.n2435 0.0213333
R10908 VDD.n2434 VDD.n2433 0.0213333
R10909 VDD.n2420 VDD.n2419 0.0213333
R10910 VDD VDD.n4774 0.0213333
R10911 VDD VDD.n3451 0.0213333
R10912 VDD VDD.n2734 0.0213333
R10913 VDD.n3061 VDD.n3060 0.0212094
R10914 VDD.n2869 VDD.n2868 0.0210625
R10915 VDD.n3099 VDD.n3098 0.0209156
R10916 VDD.n1198 VDD.n283 0.0207703
R10917 VDD.n3397 VDD.n2728 0.0207703
R10918 VDD.n4172 VDD.n4120 0.0207703
R10919 VDD.n670 VDD.n651 0.0207703
R10920 VDD.n2763 VDD.n2762 0.0207703
R10921 VDD.n3002 VDD.n3001 0.0207703
R10922 VDD.n2971 VDD.n2970 0.0207703
R10923 VDD.n3199 VDD.n3151 0.0207703
R10924 VDD.n4203 VDD.n4201 0.0207703
R10925 VDD.n1086 VDD.n1082 0.0207703
R10926 VDD.n927 VDD.n925 0.0207703
R10927 VDD.n1190 VDD.n1060 0.0207703
R10928 VDD.n3092 VDD.n3091 0.0203281
R10929 VDD.n666 VDD.n661 0.0200312
R10930 VDD.n3636 VDD.n3631 0.0200312
R10931 VDD.n3643 VDD.n3642 0.0200312
R10932 VDD.n2654 VDD.n2649 0.0200312
R10933 VDD.n2662 VDD.n2661 0.0200312
R10934 VDD.n2834 VDD.n2824 0.0200312
R10935 VDD.n2839 VDD.n2838 0.0200312
R10936 VDD.n2863 VDD.n2855 0.0200312
R10937 VDD.n2806 VDD.n2804 0.0200312
R10938 VDD.n2916 VDD.n2910 0.0200312
R10939 VDD.n2997 VDD.n2992 0.0200312
R10940 VDD.n3124 VDD.n3123 0.0200312
R10941 VDD.n4382 VDD.n4364 0.0200312
R10942 VDD.n2623 VDD.n2621 0.0200312
R10943 VDD.n4156 VDD.n4155 0.0200312
R10944 VDD.n1228 VDD.n1227 0.0200312
R10945 VDD.n1244 VDD.n1243 0.0200312
R10946 VDD.n1258 VDD.n1257 0.0200312
R10947 VDD.n1272 VDD.n1271 0.0200312
R10948 VDD.n1286 VDD.n1285 0.0200312
R10949 VDD.n1300 VDD.n1299 0.0200312
R10950 VDD.n1316 VDD.n1315 0.0200312
R10951 VDD.n1330 VDD.n1329 0.0200312
R10952 VDD.n1347 VDD.n1346 0.0200312
R10953 VDD.n1449 VDD.n1448 0.0200312
R10954 VDD.n1472 VDD.n1465 0.0200312
R10955 VDD.n2320 VDD.n207 0.0200312
R10956 VDD VDD.n3223 0.0200312
R10957 VDD VDD.n4874 0.0198461
R10958 VDD.n1551 VDD.n1540 0.0198299
R10959 VDD.n1471 VDD.n1466 0.0190811
R10960 VDD.n2664 VDD.n2648 0.0190811
R10961 VDD.n3641 VDD.n3639 0.0190811
R10962 VDD.n1993 VDD.n1992 0.0190811
R10963 VDD.n2865 VDD.n2864 0.0190811
R10964 VDD.n2833 VDD.n2826 0.0190811
R10965 VDD.n632 VDD.n625 0.0187292
R10966 VDD.n669 VDD.n656 0.0187292
R10967 VDD.n1981 VDD.n1980 0.0187292
R10968 VDD.n1811 VDD.n1809 0.0187292
R10969 VDD.n4079 VDD.n4077 0.0187292
R10970 VDD.n132 VDD.n130 0.0187292
R10971 VDD.n2969 VDD.n2954 0.0187292
R10972 VDD.n2966 VDD.n2961 0.0187292
R10973 VDD.n3000 VDD.n2985 0.0187292
R10974 VDD.n3025 VDD.n3020 0.0187292
R10975 VDD.n3119 VDD.n3118 0.0187292
R10976 VDD.n3197 VDD.n3196 0.0187292
R10977 VDD.n708 VDD.n707 0.0187292
R10978 VDD.n1188 VDD.n1187 0.0187292
R10979 VDD.n1089 VDD.n1087 0.0187292
R10980 VDD.n4566 VDD.n4561 0.0187292
R10981 VDD.n4171 VDD.n4131 0.0187292
R10982 VDD.n4158 VDD.n4157 0.0187292
R10983 VDD.n224 VDD.n223 0.0187292
R10984 VDD.n239 VDD.n226 0.0187292
R10985 VDD.n3396 VDD.n2733 0.0187292
R10986 VDD.n3393 VDD.n3388 0.0187292
R10987 VDD.n3304 VDD.n3302 0.0187292
R10988 VDD.n1538 VDD.n1537 0.0185412
R10989 VDD.n296 VDD.n290 0.0174271
R10990 VDD.n3747 VDD.n3744 0.0174271
R10991 VDD.n2678 VDD.n2672 0.0174271
R10992 VDD.n4856 VDD.n4854 0.0174271
R10993 VDD.n144 VDD.n139 0.0174271
R10994 VDD.n148 VDD.n146 0.0174271
R10995 VDD.n148 VDD.n147 0.0174271
R10996 VDD.n3030 VDD.n3015 0.0174271
R10997 VDD.n3030 VDD.n3029 0.0174271
R10998 VDD.n3047 VDD.n3040 0.0174271
R10999 VDD.n3055 VDD.n3049 0.0174271
R11000 VDD.n3055 VDD.n3054 0.0174271
R11001 VDD.n3074 VDD.n3072 0.0174271
R11002 VDD.n3157 VDD.n3152 0.0174271
R11003 VDD.n716 VDD.n715 0.0174271
R11004 VDD.n1185 VDD.n1068 0.0174271
R11005 VDD.n1612 VDD.n1605 0.0174271
R11006 VDD.n1612 VDD.n1611 0.0174271
R11007 VDD.n4697 VDD.n4695 0.0174271
R11008 VDD.n4140 VDD.n4139 0.0174271
R11009 VDD.n1522 VDD.n1521 0.0174271
R11010 VDD.n2136 VDD.n2134 0.0173919
R11011 VDD.n1414 VDD.n258 0.0173919
R11012 VDD.n2454 VDD.n2453 0.0173919
R11013 VDD.n4219 VDD.n2645 0.0173919
R11014 VDD.n3591 VDD.n3590 0.0173919
R11015 VDD.n3552 VDD.n3528 0.0173919
R11016 VDD.n2936 VDD.n2798 0.0173919
R11017 VDD.n669 VDD.n668 0.016125
R11018 VDD.n1760 VDD.n1758 0.016125
R11019 VDD.n1780 VDD.n1779 0.016125
R11020 VDD.n86 VDD.n82 0.016125
R11021 VDD.n2969 VDD.n2968 0.016125
R11022 VDD.n3000 VDD.n2999 0.016125
R11023 VDD.n3122 VDD.n3119 0.016125
R11024 VDD.n3197 VDD.n3159 0.016125
R11025 VDD.n710 VDD.n708 0.016125
R11026 VDD.n1188 VDD.n1067 0.016125
R11027 VDD.n1087 VDD.n1080 0.016125
R11028 VDD.n1590 VDD.n1588 0.016125
R11029 VDD.n1589 VDD 0.016125
R11030 VDD.n1603 VDD.n1598 0.016125
R11031 VDD.n2339 VDD.n2337 0.016125
R11032 VDD.n2338 VDD 0.016125
R11033 VDD.n2371 VDD.n2369 0.016125
R11034 VDD.n4363 VDD.n4360 0.016125
R11035 VDD.n4171 VDD.n4170 0.016125
R11036 VDD.n4134 VDD.n4132 0.016125
R11037 VDD.n1200 VDD.n1199 0.016125
R11038 VDD.n4710 VDD 0.016125
R11039 VDD.n3396 VDD.n3395 0.016125
R11040 VDD.n4194 VDD.n4192 0.0158047
R11041 VDD.n1524 VDD.n1429 0.0157027
R11042 VDD.n4810 VDD.n171 0.0157027
R11043 VDD.n4593 VDD.n2541 0.0157027
R11044 VDD.n3834 VDD.n3829 0.0157027
R11045 VDD.n491 VDD.n490 0.0157027
R11046 VDD.n1709 VDD.n251 0.0157027
R11047 VDD.n3233 VDD.n3232 0.0157027
R11048 VDD.n36 VDD.n18 0.0157027
R11049 VDD.n3148 VDD.n2773 0.0157027
R11050 VDD.n647 VDD.n644 0.0152558
R11051 VDD.n585 VDD.n581 0.0152558
R11052 VDD.n1885 VDD.n1846 0.0152558
R11053 VDD.n1885 VDD.n1884 0.0152558
R11054 VDD.n2150 VDD.n241 0.0152558
R11055 VDD.n2150 VDD.n2149 0.0152558
R11056 VDD.n1470 VDD.n1468 0.0152558
R11057 VDD.n1470 VDD.n1469 0.0152558
R11058 VDD.n1525 VDD.n1427 0.0152558
R11059 VDD.n1525 VDD.n1428 0.0152558
R11060 VDD.n1700 VDD.n1634 0.0152558
R11061 VDD.n1700 VDD.n1699 0.0152558
R11062 VDD.n918 VDD.n300 0.0152558
R11063 VDD.n918 VDD.n301 0.0152558
R11064 VDD.n1196 VDD.n284 0.0152558
R11065 VDD.n1196 VDD.n1195 0.0152558
R11066 VDD.n2137 VDD.n2132 0.0152558
R11067 VDD.n2137 VDD.n2133 0.0152558
R11068 VDD.n1415 VDD.n255 0.0152558
R11069 VDD.n1415 VDD.n256 0.0152558
R11070 VDD.n2326 VDD.n188 0.0152558
R11071 VDD.n2326 VDD.n2325 0.0152558
R11072 VDD.n2455 VDD.n2379 0.0152558
R11073 VDD.n2455 VDD.n2380 0.0152558
R11074 VDD.n4707 VDD.n174 0.0152558
R11075 VDD.n167 VDD.n166 0.0152558
R11076 VDD.n4811 VDD.n170 0.0152558
R11077 VDD.n3398 VDD.n2726 0.0152558
R11078 VDD.n2719 VDD.n2681 0.0152558
R11079 VDD.n3510 VDD.n3509 0.0152558
R11080 VDD.n1630 VDD.n1627 0.0152558
R11081 VDD.n4413 VDD.n4412 0.0152558
R11082 VDD.n2332 VDD.n185 0.0152558
R11083 VDD.n2332 VDD.n2331 0.0152558
R11084 VDD.n2571 VDD.n2570 0.0152558
R11085 VDD.n4591 VDD.n2542 0.0152558
R11086 VDD.n4586 VDD.n4585 0.0152558
R11087 VDD.n4538 VDD.n2574 0.0152558
R11088 VDD.n4419 VDD.n2611 0.0152558
R11089 VDD.n4346 VDD.n4319 0.0152558
R11090 VDD.n4410 VDD.n4389 0.0152558
R11091 VDD.n4386 VDD.n4385 0.0152558
R11092 VDD.n4218 VDD.n4217 0.0152558
R11093 VDD.n4173 VDD.n4118 0.0152558
R11094 VDD.n1426 VDD.n1423 0.0152558
R11095 VDD.n3592 VDD.n3588 0.0152558
R11096 VDD.n3978 VDD.n2680 0.0152558
R11097 VDD.n2665 VDD.n2647 0.0152558
R11098 VDD.n4107 VDD.n4085 0.0152558
R11099 VDD.n4082 VDD.n2668 0.0152558
R11100 VDD.n3626 VDD.n3595 0.0152558
R11101 VDD.n3773 VDD.n3749 0.0152558
R11102 VDD.n3794 VDD.n3793 0.0152558
R11103 VDD.n3813 VDD.n3811 0.0152558
R11104 VDD.n3833 VDD.n3832 0.0152558
R11105 VDD.n3974 VDD.n3973 0.0152558
R11106 VDD.n3578 VDD.n3556 0.0152558
R11107 VDD.n3553 VDD.n3527 0.0152558
R11108 VDD.n2524 VDD.n2522 0.0152558
R11109 VDD.n2524 VDD.n2523 0.0152558
R11110 VDD.n935 VDD.n298 0.0152558
R11111 VDD.n935 VDD.n934 0.0152558
R11112 VDD.n671 VDD.n648 0.0152558
R11113 VDD.n671 VDD.n649 0.0152558
R11114 VDD.n492 VDD.n418 0.0152558
R11115 VDD.n492 VDD.n419 0.0152558
R11116 VDD.n611 VDD.n586 0.0152558
R11117 VDD.n611 VDD.n587 0.0152558
R11118 VDD.n636 VDD.n616 0.0152558
R11119 VDD.n636 VDD.n617 0.0152558
R11120 VDD.n1049 VDD.n286 0.0152558
R11121 VDD.n1049 VDD.n287 0.0152558
R11122 VDD.n1708 VDD.n252 0.0152558
R11123 VDD.n1708 VDD.n253 0.0152558
R11124 VDD.n1765 VDD.n243 0.0152558
R11125 VDD.n1765 VDD.n1764 0.0152558
R11126 VDD.n1994 VDD.n1772 0.0152558
R11127 VDD.n1994 VDD.n1773 0.0152558
R11128 VDD.n1891 VDD.n1813 0.0152558
R11129 VDD.n1891 VDD.n1890 0.0152558
R11130 VDD.n1841 VDD.n1815 0.0152558
R11131 VDD.n1841 VDD.n1816 0.0152558
R11132 VDD.n2478 VDD.n2459 0.0152558
R11133 VDD.n2478 VDD.n2477 0.0152558
R11134 VDD.n3263 VDD.n3236 0.0152558
R11135 VDD.n3234 VDD.n3230 0.0152558
R11136 VDD.n3312 VDD.n3274 0.0152558
R11137 VDD.n3227 VDD.n3210 0.0152558
R11138 VDD.n4198 VDD.n4176 0.0152558
R11139 VDD.n156 VDD.n155 0.0152558
R11140 VDD.n11 VDD.n1 0.0152558
R11141 VDD.n2767 VDD.n2766 0.0152558
R11142 VDD.n2764 VDD.n2760 0.0152558
R11143 VDD.n3089 VDD.n3062 0.0152558
R11144 VDD.n3089 VDD.n3063 0.0152558
R11145 VDD.n3096 VDD.n3093 0.0152558
R11146 VDD.n3101 VDD.n2790 0.0152558
R11147 VDD.n3101 VDD.n2791 0.0152558
R11148 VDD.n3058 VDD.n3037 0.0152558
R11149 VDD.n3058 VDD.n3038 0.0152558
R11150 VDD.n3004 VDD.n2977 0.0152558
R11151 VDD.n3004 VDD.n3003 0.0152558
R11152 VDD.n2906 VDD.n2896 0.0152558
R11153 VDD.n2906 VDD.n2905 0.0152558
R11154 VDD.n2873 VDD.n2808 0.0152558
R11155 VDD.n2873 VDD.n2872 0.0152558
R11156 VDD.n2866 VDD.n2810 0.0152558
R11157 VDD.n2866 VDD.n2811 0.0152558
R11158 VDD.n2832 VDD.n2827 0.0152558
R11159 VDD.n2832 VDD.n2831 0.0152558
R11160 VDD.n63 VDD.n62 0.0152558
R11161 VDD.n37 VDD.n17 0.0152558
R11162 VDD.n91 VDD.n90 0.0152558
R11163 VDD.n4868 VDD.n4847 0.0152558
R11164 VDD.n4868 VDD.n4867 0.0152558
R11165 VDD.n135 VDD.n94 0.0152558
R11166 VDD.n152 VDD.n151 0.0152558
R11167 VDD.n2937 VDD.n2796 0.0152558
R11168 VDD.n2937 VDD.n2797 0.0152558
R11169 VDD.n2899 VDD.n2898 0.0152558
R11170 VDD.n2973 VDD.n2942 0.0152558
R11171 VDD.n2973 VDD.n2972 0.0152558
R11172 VDD.n3149 VDD.n2772 0.0152558
R11173 VDD.n3201 VDD.n3200 0.0152558
R11174 VDD.n3172 VDD.n3171 0.0152558
R11175 VDD.n3033 VDD.n3008 0.0152558
R11176 VDD.n3033 VDD.n3032 0.0152558
R11177 VDD.n4204 VDD.n4200 0.0152558
R11178 VDD.n4548 VDD.n4544 0.0152558
R11179 VDD.n4700 VDD.n2525 0.0152558
R11180 VDD.n4700 VDD.n2526 0.0152558
R11181 VDD.n2517 VDD.n2482 0.0152558
R11182 VDD.n2375 VDD.n176 0.0152558
R11183 VDD.n2375 VDD.n177 0.0152558
R11184 VDD.n2131 VDD.n1995 0.0152558
R11185 VDD.n2131 VDD.n1996 0.0152558
R11186 VDD.n1614 VDD.n1529 0.0152558
R11187 VDD.n1614 VDD.n1530 0.0152558
R11188 VDD.n1528 VDD.n1526 0.0152558
R11189 VDD.n1528 VDD.n1527 0.0152558
R11190 VDD.n1422 VDD.n1420 0.0152558
R11191 VDD.n1422 VDD.n1421 0.0152558
R11192 VDD.n615 VDD.n612 0.0152558
R11193 VDD.n1085 VDD.n1083 0.0152558
R11194 VDD.n1085 VDD.n1084 0.0152558
R11195 VDD.n643 VDD.n637 0.0152558
R11196 VDD.n643 VDD.n638 0.0152558
R11197 VDD.n580 VDD.n493 0.0152558
R11198 VDD.n580 VDD.n494 0.0152558
R11199 VDD.n745 VDD.n672 0.0152558
R11200 VDD.n745 VDD.n673 0.0152558
R11201 VDD.n928 VDD.n923 0.0152558
R11202 VDD.n928 VDD.n924 0.0152558
R11203 VDD.n1192 VDD.n1059 0.0152558
R11204 VDD.n1192 VDD.n1191 0.0152558
R11205 VDD.n4314 VDD.n2613 0.0152558
R11206 VDD.n4831 VDD.n4830 0.0152558
R11207 VDD.n776 VDD.n415 0.0152558
R11208 VDD.n602 VDD.n600 0.0148229
R11209 VDD.n1991 VDD.n1990 0.0148229
R11210 VDD.n3642 VDD.n3638 0.0148229
R11211 VDD.n3964 VDD.n3962 0.0148229
R11212 VDD.n3548 VDD.n3543 0.0148229
R11213 VDD.n2662 VDD.n2656 0.0148229
R11214 VDD.n3246 VDD.n3240 0.0148229
R11215 VDD.n2837 VDD.n2834 0.0148229
R11216 VDD.n2863 VDD.n2862 0.0148229
R11217 VDD.n2926 VDD.n2925 0.0148229
R11218 VDD.n3112 VDD.n3105 0.0148229
R11219 VDD.n3168 VDD.n3166 0.0148229
R11220 VDD.n1095 VDD.n1094 0.0148229
R11221 VDD.n4581 VDD.n4579 0.0148229
R11222 VDD.n4534 VDD.n4527 0.0148229
R11223 VDD.n821 VDD.n303 0.0148229
R11224 VDD.n835 VDD.n823 0.0148229
R11225 VDD.n852 VDD.n838 0.0148229
R11226 VDD.n866 VDD.n854 0.0148229
R11227 VDD.n880 VDD.n868 0.0148229
R11228 VDD.n900 VDD.n899 0.0148229
R11229 VDD.n896 VDD.n895 0.0148229
R11230 VDD.n1202 VDD.n282 0.0148229
R11231 VDD.n1375 VDD.n1348 0.0148229
R11232 VDD.n1411 VDD.n1410 0.0148229
R11233 VDD.n1661 VDD.n1649 0.0148229
R11234 VDD.n1677 VDD.n1676 0.0148229
R11235 VDD.n1503 VDD.n1501 0.0148229
R11236 VDD.n1473 VDD.n1472 0.0148229
R11237 VDD.n1879 VDD.n1865 0.0148229
R11238 VDD.n4828 VDD.n4826 0.0148229
R11239 VDD.n2718 VDD.n2717 0.0140135
R11240 VDD.n2569 VDD.n2568 0.0140135
R11241 VDD.n4345 VDD.n4320 0.0140135
R11242 VDD.n4106 VDD.n4087 0.0140135
R11243 VDD.n3577 VDD.n3557 0.0140135
R11244 VDD.n4197 VDD.n4177 0.0140135
R11245 VDD.n2941 VDD.n2940 0.0138656
R11246 VDD.n1045 VDD.n1038 0.0135208
R11247 VDD.n3822 VDD.n3817 0.0135208
R11248 VDD.n3551 VDD.n3536 0.0135208
R11249 VDD.n2853 VDD.n2849 0.0135208
R11250 VDD.n2934 VDD.n2892 0.0135208
R11251 VDD.n545 VDD.n544 0.0135208
R11252 VDD.n567 VDD.n565 0.0135208
R11253 VDD.n1151 VDD.n1136 0.0135208
R11254 VDD.n1563 VDD.n1557 0.0135208
R11255 VDD.n2114 VDD.n2099 0.0135208
R11256 VDD.n2503 VDD.n2502 0.0135208
R11257 VDD.n2564 VDD.n2549 0.0135208
R11258 VDD.n4448 VDD.n4433 0.0135208
R11259 VDD.n4270 VDD.n4255 0.0135208
R11260 VDD.n4222 VDD.n4220 0.0135208
R11261 VDD.n1379 VDD.n1378 0.0135208
R11262 VDD.n1413 VDD.n1412 0.0135208
R11263 VDD.n2285 VDD.n217 0.0135208
R11264 VDD.n2300 VDD.n2299 0.0135208
R11265 VDD.n2397 VDD.n2396 0.0135208
R11266 VDD.n2452 VDD.n2451 0.0135208
R11267 VDD.n2706 VDD.n2702 0.0135208
R11268 VDD.n1698 VDD.n1635 0.0123243
R11269 VDD.n610 VDD.n609 0.0123243
R11270 VDD.n1048 VDD.n288 0.0123243
R11271 VDD.n2476 VDD.n2461 0.0123243
R11272 VDD.n61 VDD.n60 0.0123243
R11273 VDD.n579 VDD.n578 0.0123243
R11274 VDD.n4833 VDD.n4832 0.0123243
R11275 VDD.n483 VDD.n481 0.0122188
R11276 VDD.n489 VDD.n488 0.0122188
R11277 VDD.n1714 VDD.n1710 0.0122188
R11278 VDD.n3835 VDD.n3828 0.0122188
R11279 VDD.n3843 VDD.n3842 0.0122188
R11280 VDD.n3572 VDD.n3567 0.0122188
R11281 VDD.n35 VDD.n24 0.0122188
R11282 VDD.n30 VDD.n25 0.0122188
R11283 VDD.n3146 VDD.n3138 0.0122188
R11284 VDD.n4596 VDD.n4594 0.0122188
R11285 VDD.n4342 VDD.n4335 0.0122188
R11286 VDD.n1694 VDD.n1680 0.0122188
R11287 VDD.n1522 VDD.n1430 0.0122188
R11288 VDD.n4808 VDD.n4791 0.0122188
R11289 VDD.n4805 VDD.n4800 0.0122188
R11290 VDD VDD.n4835 0.0122188
R11291 VDD.n3288 VDD.n3282 0.0122188
R11292 VDD.n481 VDD.n476 0.0109167
R11293 VDD.n3842 VDD.n3837 0.0109167
R11294 VDD.n3575 VDD.n3562 0.0109167
R11295 VDD.n3574 VDD.n3572 0.0109167
R11296 VDD.n4104 VDD.n4098 0.0109167
R11297 VDD.n34 VDD.n30 0.0109167
R11298 VDD.n1582 VDD 0.0109167
R11299 VDD VDD.n183 0.0109167
R11300 VDD.n2567 VDD.n2566 0.0109167
R11301 VDD.n4343 VDD.n4333 0.0109167
R11302 VDD.n4335 VDD.n4334 0.0109167
R11303 VDD.n4195 VDD.n4189 0.0109167
R11304 VDD.n1199 VDD.n269 0.0109167
R11305 VDD.n4807 VDD.n4805 0.0109167
R11306 VDD.n2716 VDD.n2715 0.0109167
R11307 VDD.n4420 VDD.n2609 0.0106351
R11308 VDD.n4409 VDD.n4391 0.0106351
R11309 VDD.n4384 VDD.n4383 0.0106351
R11310 VDD.n3814 VDD.n3809 0.0106351
R11311 VDD.n3972 VDD.n3971 0.0106351
R11312 VDD.n3262 VDD.n3238 0.0106351
R11313 VDD.n3173 VDD.n3169 0.0106351
R11314 VDD.n642 VDD.n641 0.0106351
R11315 VDD.n2548 VDD.n2547 0.00993343
R11316 VDD.n608 VDD.n607 0.00961458
R11317 VDD.n1046 VDD.n1036 0.00961458
R11318 VDD.n1038 VDD.n1037 0.00961458
R11319 VDD.n2474 VDD.n2466 0.00961458
R11320 VDD.n3823 VDD.n3822 0.00961458
R11321 VDD.n58 VDD.n57 0.00961458
R11322 VDD.n2855 VDD.n2853 0.00961458
R11323 VDD.n544 VDD.n529 0.00961458
R11324 VDD.n565 VDD.n560 0.00961458
R11325 VDD.n577 VDD.n576 0.00961458
R11326 VDD.n1152 VDD.n1151 0.00961458
R11327 VDD.n2115 VDD.n2114 0.00961458
R11328 VDD.n2502 VDD.n2487 0.00961458
R11329 VDD.n2565 VDD.n2564 0.00961458
R11330 VDD.n4449 VDD.n4448 0.00961458
R11331 VDD.n4271 VDD.n4270 0.00961458
R11332 VDD.n1696 VDD.n1663 0.00961458
R11333 VDD.n1520 VDD.n1488 0.00961458
R11334 VDD.n2299 VDD.n2298 0.00961458
R11335 VDD.n4835 VDD.n4834 0.00961458
R11336 VDD.n2702 VDD.n2697 0.00961458
R11337 VDD.n1883 VDD.n1847 0.00894595
R11338 VDD.n2334 VDD.n184 0.00894595
R11339 VDD.n4584 VDD.n4552 0.00894595
R11340 VDD.n4537 VDD.n2575 0.00894595
R11341 VDD.n3980 VDD.n3979 0.00894595
R11342 VDD.n3775 VDD.n3774 0.00894595
R11343 VDD.n1763 VDD.n244 0.00894595
R11344 VDD.n3088 VDD.n3087 0.00894595
R11345 VDD.n3102 VDD.n2788 0.00894595
R11346 VDD.n2374 VDD.n179 0.00894595
R11347 VDD.n1585 VDD.n1583 0.00894595
R11348 VDD.n600 VDD.n593 0.0083125
R11349 VDD.n3815 VDD.n3808 0.0083125
R11350 VDD.n3962 VDD.n3957 0.0083125
R11351 VDD.n3970 VDD.n3969 0.0083125
R11352 VDD.n3550 VDD.n3548 0.0083125
R11353 VDD.n3240 VDD.n3239 0.0083125
R11354 VDD.n3261 VDD.n3260 0.0083125
R11355 VDD.n2933 VDD.n2926 0.0083125
R11356 VDD.n3113 VDD.n3112 0.0083125
R11357 VDD.n3175 VDD.n3174 0.0083125
R11358 VDD.n3166 VDD.n3165 0.0083125
R11359 VDD.n695 VDD.n691 0.0083125
R11360 VDD.n1094 VDD.n1089 0.0083125
R11361 VDD.n4579 VDD.n4572 0.0083125
R11362 VDD.n4527 VDD.n4526 0.0083125
R11363 VDD.n4427 VDD.n4421 0.0083125
R11364 VDD.n4408 VDD.n4401 0.0083125
R11365 VDD.n4382 VDD.n4381 0.0083125
R11366 VDD.n822 VDD.n821 0.0083125
R11367 VDD.n836 VDD.n835 0.0083125
R11368 VDD.n853 VDD.n852 0.0083125
R11369 VDD.n867 VDD.n866 0.0083125
R11370 VDD.n881 VDD.n880 0.0083125
R11371 VDD.n895 VDD.n883 0.0083125
R11372 VDD.n1202 VDD.n1201 0.0083125
R11373 VDD.n1222 VDD.n269 0.0083125
R11374 VDD.n1224 VDD.n1223 0.0083125
R11375 VDD.n1225 VDD.n1224 0.0083125
R11376 VDD.n1376 VDD.n1375 0.0083125
R11377 VDD.n1380 VDD.n1379 0.0083125
R11378 VDD.n1410 VDD.n1398 0.0083125
R11379 VDD.n1648 VDD.n1647 0.0083125
R11380 VDD.n1662 VDD.n1661 0.0083125
R11381 VDD.n1680 VDD.n1679 0.0083125
R11382 VDD.n1676 VDD.n1664 0.0083125
R11383 VDD.n1503 VDD.n1502 0.0083125
R11384 VDD.n1488 VDD.n1487 0.0083125
R11385 VDD.n1486 VDD 0.0083125
R11386 VDD VDD.n2300 0.0083125
R11387 VDD.n2452 VDD.n2397 0.0083125
R11388 VDD.n4826 VDD.n4821 0.0083125
R11389 VDD.n3224 VDD 0.0083125
R11390 VDD.n4846 VDD.n4845 0.00769688
R11391 VDD.n937 VDD.n936 0.00725676
R11392 VDD.n89 VDD.n65 0.00725676
R11393 VDD.n4866 VDD.n4865 0.00725676
R11394 VDD.n4547 VDD.n4546 0.00725676
R11395 VDD.n4699 VDD.n2527 0.00725676
R11396 VDD.n1761 VDD.n1752 0.00701042
R11397 VDD.n1758 VDD.n1753 0.00701042
R11398 VDD.n3777 VDD.n3776 0.00701042
R11399 VDD.n3982 VDD.n3981 0.00701042
R11400 VDD.n82 VDD.n77 0.00701042
R11401 VDD.n3086 VDD.n3085 0.00701042
R11402 VDD.n3103 VDD.n2787 0.00701042
R11403 VDD.n731 VDD.n730 0.00701042
R11404 VDD.n1586 VDD.n1582 0.00701042
R11405 VDD.n1590 VDD.n1589 0.00701042
R11406 VDD.n1605 VDD.n1603 0.00701042
R11407 VDD.n2335 VDD.n183 0.00701042
R11408 VDD.n2339 VDD.n2338 0.00701042
R11409 VDD.n2369 VDD.n2364 0.00701042
R11410 VDD.n2373 VDD.n2372 0.00701042
R11411 VDD.n4582 VDD.n4557 0.00701042
R11412 VDD.n4535 VDD.n2588 0.00701042
R11413 VDD.n4360 VDD.n4349 0.00701042
R11414 VDD.n4364 VDD.n4363 0.00701042
R11415 VDD.n1223 VDD.n1222 0.00701042
R11416 VDD.n1881 VDD.n1862 0.00701042
R11417 VDD.n1880 VDD.n1879 0.00701042
R11418 VDD.n1864 VDD.n1863 0.00701042
R11419 VDD.n4840 VDD.n4839 0.00623493
R11420 VDD.n2724 VDD.n2723 0.00623493
R11421 VDD.n3399 VDD.n3398 0.00623493
R11422 VDD.n3518 VDD.n3517 0.00623493
R11423 VDD.n2572 VDD.n2571 0.00623493
R11424 VDD.n4587 VDD.n4586 0.00623493
R11425 VDD.n4387 VDD.n4386 0.00623493
R11426 VDD.n3316 VDD.n3315 0.00623493
R11427 VDD.n4218 VDD.n4216 0.00623493
R11428 VDD.n4174 VDD.n4173 0.00623493
R11429 VDD.n3794 VDD.n3792 0.00623493
R11430 VDD.n3833 VDD.n3831 0.00623493
R11431 VDD.n3975 VDD.n3974 0.00623493
R11432 VDD.n3554 VDD.n3553 0.00623493
R11433 VDD.n3313 VDD.n3312 0.00623493
R11434 VDD.n4213 VDD.n4212 0.00623493
R11435 VDD.n64 VDD.n63 0.00623493
R11436 VDD.n92 VDD.n91 0.00623493
R11437 VDD.n136 VDD.n135 0.00623493
R11438 VDD.n153 VDD.n152 0.00623493
R11439 VDD.n3202 VDD.n3201 0.00623493
R11440 VDD.n4549 VDD.n4548 0.00623493
R11441 VDD.n535 VDD.n530 0.00593478
R11442 VDD.n1142 VDD.n1137 0.00593478
R11443 VDD.n2105 VDD.n2100 0.00593478
R11444 VDD.n2493 VDD.n2488 0.00593478
R11445 VDD.n2555 VDD.n2550 0.00593478
R11446 VDD.n4439 VDD.n4434 0.00593478
R11447 VDD.n4261 VDD.n4256 0.00593478
R11448 VDD.n3264 VDD.n3263 0.00590289
R11449 VDD.n2666 VDD.n2665 0.00590289
R11450 VDD.n4083 VDD.n4082 0.00590289
R11451 VDD.n4108 VDD.n4107 0.00590289
R11452 VDD.n3235 VDD.n3234 0.00590289
R11453 VDD.n3228 VDD.n3227 0.00590289
R11454 VDD.n4199 VDD.n4198 0.00590289
R11455 VDD.n2765 VDD.n2764 0.00590289
R11456 VDD.n3150 VDD.n3149 0.00590289
R11457 VDD.n3172 VDD.n2771 0.00590289
R11458 VDD.n4205 VDD.n4204 0.00590289
R11459 VDD.n3593 VDD.n3592 0.00590289
R11460 VDD.n3627 VDD.n3626 0.00590289
R11461 VDD.n3978 VDD.n3977 0.00590289
R11462 VDD.n4419 VDD.n4418 0.00590289
R11463 VDD.n4411 VDD.n4410 0.00590289
R11464 VDD.n2720 VDD.n2719 0.00590289
R11465 VDD.n3579 VDD.n3578 0.00590289
R11466 VDD.n4347 VDD.n4346 0.00590289
R11467 VDD.n4315 VDD.n4314 0.00590289
R11468 VDD.n4812 VDD.n4811 0.00590289
R11469 VDD.n3773 VDD.n3772 0.00590289
R11470 VDD.n3813 VDD.n3812 0.00590289
R11471 VDD.n3859 VDD.n3858 0.00590289
R11472 VDD.n4591 VDD.n4590 0.00590289
R11473 VDD.n4539 VDD.n4538 0.00590289
R11474 VDD.n38 VDD.n37 0.00590289
R11475 VDD.n4831 VDD.n165 0.00590289
R11476 VDD.n290 VDD.n289 0.00570833
R11477 VDD.n939 VDD.n938 0.00570833
R11478 VDD.n3744 VDD.n3739 0.00570833
R11479 VDD.n2672 VDD.n2671 0.00570833
R11480 VDD.n4854 VDD.n4849 0.00570833
R11481 VDD.n4864 VDD.n4863 0.00570833
R11482 VDD.n87 VDD.n76 0.00570833
R11483 VDD.n146 VDD.n144 0.00570833
R11484 VDD.n3049 VDD.n3047 0.00570833
R11485 VDD.n3072 VDD.n3065 0.00570833
R11486 VDD.n3159 VDD.n3157 0.00570833
R11487 VDD.n715 VDD.n710 0.00570833
R11488 VDD.n1187 VDD.n1185 0.00570833
R11489 VDD.n4698 VDD.n2529 0.00570833
R11490 VDD.n4695 VDD.n4690 0.00570833
R11491 VDD.n4559 VDD.n4558 0.00570833
R11492 VDD.n4139 VDD.n4134 0.00570833
R11493 VDD VDD.n1225 0.00570833
R11494 VDD.n1521 VDD.n1520 0.00570833
R11495 VDD.n1487 VDD.n1486 0.00570833
R11496 VDD.n4081 VDD.n2669 0.00556757
R11497 VDD.n3625 VDD.n3597 0.00556757
R11498 VDD.n635 VDD.n618 0.00556757
R11499 VDD.n1840 VDD.n1839 0.00556757
R11500 VDD.n3311 VDD.n3276 0.00556757
R11501 VDD.n2907 VDD.n2895 0.00556757
R11502 VDD.n2875 VDD.n2874 0.00556757
R11503 VDD.n4313 VDD.n2615 0.00556757
R11504 VDD.n3206 VDD.n2757 0.0052
R11505 VDD.n2974 VDD.n2941 0.00490625
R11506 VDD.n2975 VDD.n2974 0.00490625
R11507 VDD.n3005 VDD.n2976 0.00490625
R11508 VDD.n3006 VDD.n3005 0.00490625
R11509 VDD.n3034 VDD.n3007 0.00490625
R11510 VDD.n3035 VDD.n3034 0.00490625
R11511 VDD.n3059 VDD.n3036 0.00490625
R11512 VDD.n3060 VDD.n3059 0.00490625
R11513 VDD.n3090 VDD.n3061 0.00490625
R11514 VDD.n3091 VDD.n3090 0.00490625
R11515 VDD.n3097 VDD.n3092 0.00490625
R11516 VDD.n3098 VDD.n3097 0.00490625
R11517 VDD.n3100 VDD.n3099 0.00490625
R11518 VDD.n3100 VDD.n2757 0.00490625
R11519 VDD.n2830 VDD.n2828 0.00490625
R11520 VDD.n2830 VDD.n2829 0.00490625
R11521 VDD.n2867 VDD.n2809 0.00490625
R11522 VDD.n2868 VDD.n2867 0.00490625
R11523 VDD.n2871 VDD.n2869 0.00490625
R11524 VDD.n2871 VDD.n2870 0.00490625
R11525 VDD.n2938 VDD.n2795 0.00490625
R11526 VDD.n2939 VDD.n2938 0.00490625
R11527 VDD.n4873 VDD.n4872 0.00490625
R11528 VDD.n4872 VDD.n4871 0.00490625
R11529 VDD.n4870 VDD.n4869 0.00490625
R11530 VDD.n4869 VDD.n4846 0.00490625
R11531 VDD.n4212 VDD.n4211 0.00480456
R11532 VDD.n3317 VDD.n3316 0.00480456
R11533 VDD.n2723 VDD.n2722 0.00480456
R11534 VDD.n3517 VDD.n3516 0.00480456
R11535 VDD.n4839 VDD.n4838 0.00480456
R11536 VDD.n633 VDD.n623 0.00440625
R11537 VDD.n625 VDD.n624 0.00440625
R11538 VDD.n1991 VDD.n1780 0.00440625
R11539 VDD.n1809 VDD.n1804 0.00440625
R11540 VDD.n1837 VDD.n1836 0.00440625
R11541 VDD.n3624 VDD.n3618 0.00440625
R11542 VDD.n4080 VDD.n4071 0.00440625
R11543 VDD.n4077 VDD.n4072 0.00440625
R11544 VDD.n130 VDD.n123 0.00440625
R11545 VDD.n2877 VDD.n2876 0.00440625
R11546 VDD.n2908 VDD.n2893 0.00440625
R11547 VDD.n2968 VDD.n2966 0.00440625
R11548 VDD.n3029 VDD.n3025 0.00440625
R11549 VDD VDD.n3160 0.00440625
R11550 VDD.n4567 VDD.n4566 0.00440625
R11551 VDD.n4312 VDD.n4311 0.00440625
R11552 VDD.n4170 VDD.n4158 0.00440625
R11553 VDD.n914 VDD.n900 0.00440625
R11554 VDD.n899 VDD.n898 0.00440625
R11555 VDD.n898 VDD.n897 0.00440625
R11556 VDD.n1227 VDD 0.00440625
R11557 VDD.n3395 VDD.n3393 0.00440625
R11558 VDD.n3302 VDD.n3297 0.00440625
R11559 VDD.n3310 VDD.n3309 0.00440625
R11560 VDD.n770 VDD.n769 0.00409617
R11561 VDD.n647 VDD.n646 0.00390995
R11562 VDD.n585 VDD.n584 0.00390995
R11563 VDD.n4708 VDD.n4707 0.00390995
R11564 VDD.n1630 VDD.n1629 0.00390995
R11565 VDD.n1426 VDD.n1425 0.00390995
R11566 VDD.n3860 VDD.n3859 0.00390995
R11567 VDD.n11 VDD.n10 0.00390995
R11568 VDD.n3096 VDD.n3095 0.00390995
R11569 VDD.n2517 VDD.n2516 0.00390995
R11570 VDD.n615 VDD.n614 0.00390995
R11571 VDD.n777 VDD.n776 0.00390995
R11572 VDD.n2152 VDD.n2151 0.00387838
R11573 VDD.n917 VDD.n302 0.00387838
R11574 VDD.n2324 VDD.n189 0.00387838
R11575 VDD.n1893 VDD.n1812 0.00387838
R11576 VDD.n134 VDD.n95 0.00387838
R11577 VDD.n2130 VDD.n1999 0.00387838
R11578 VDD.n1554 VDD.n1553 0.00387838
R11579 VDD.n1620 VDD.n1619 0.00341357
R11580 VDD.n1888 VDD.n1887 0.00329702
R11581 VDD.n4845 VDD.n12 0.00329063
R11582 VDD.n931 VDD.n930 0.00319713
R11583 VDD.n2141 VDD.n2140 0.00314718
R11584 VDD.n668 VDD.n666 0.00310417
R11585 VDD.n1990 VDD.n1982 0.00310417
R11586 VDD.n1895 VDD.n1894 0.00310417
R11587 VDD.n3638 VDD.n3636 0.00310417
R11588 VDD.n2656 VDD.n2654 0.00310417
R11589 VDD.n133 VDD.n118 0.00310417
R11590 VDD.n2839 VDD.n2837 0.00310417
R11591 VDD.n2804 VDD.n2799 0.00310417
R11592 VDD.n2917 VDD.n2916 0.00310417
R11593 VDD.n2999 VDD.n2997 0.00310417
R11594 VDD.n3124 VDD.n3122 0.00310417
R11595 VDD.n2129 VDD.n2128 0.00310417
R11596 VDD.n2621 VDD.n2616 0.00310417
R11597 VDD.n4155 VDD.n4141 0.00310417
R11598 VDD.n915 VDD.n882 0.00310417
R11599 VDD.n1228 VDD.n1226 0.00310417
R11600 VDD.n1243 VDD.n259 0.00310417
R11601 VDD.n1257 VDD.n1245 0.00310417
R11602 VDD.n1271 VDD.n1259 0.00310417
R11603 VDD.n1285 VDD.n1273 0.00310417
R11604 VDD.n1299 VDD.n1287 0.00310417
R11605 VDD.n1315 VDD.n1301 0.00310417
R11606 VDD.n1329 VDD.n1317 0.00310417
R11607 VDD.n1346 VDD.n1331 0.00310417
R11608 VDD.n1695 VDD.n1694 0.00310417
R11609 VDD.n1679 VDD.n1678 0.00310417
R11610 VDD.n225 VDD.n224 0.00310417
R11611 VDD.n2154 VDD.n2153 0.00310417
R11612 VDD.n2322 VDD.n190 0.00310417
R11613 VDD.n3514 VDD 0.00310417
R11614 VDD.n2329 VDD.n2328 0.00309724
R11615 VDD.n1556 VDD.n1555 0.00307732
R11616 VDD.n1626 VDD.n1625 0.00293075
R11617 VDD.n1769 VDD.n1768 0.00286415
R11618 VDD.n761 VDD.n760 0.00266436
R11619 VDD.n4415 VDD.n4413 0.00246557
R11620 VDD.n2901 VDD.n2899 0.00246557
R11621 VDD.n3795 VDD.n3791 0.00218919
R11622 VDD.n3226 VDD.n3212 0.00218919
R11623 VDD.n168 VDD.n167 0.00213281
R11624 VDD.n3511 VDD.n3510 0.00213281
R11625 VDD.n158 VDD.n156 0.00213281
R11626 VDD.n2769 VDD.n2767 0.00213281
R11627 VDD.n3206 VDD.n3205 0.00206133
R11628 VDD.n1419 VDD.n1418 0.0020317
R11629 VDD.n746 VDD.n299 0.00193181
R11630 VDD.n1057 VDD.n1056 0.00186521
R11631 VDD.n2520 VDD.n2519 0.00181527
R11632 VDD.n448 VDD.n447 0.00180208
R11633 VDD.n982 VDD.n981 0.00180208
R11634 VDD.n1982 VDD.n1981 0.00180208
R11635 VDD.n1825 VDD.n1824 0.00180208
R11636 VDD.n3738 VDD.n3737 0.00180208
R11637 VDD.n3787 VDD.n3782 0.00180208
R11638 VDD.n3797 VDD.n3796 0.00180208
R11639 VDD.n3871 VDD.n3870 0.00180208
R11640 VDD.n3937 VDD.n3936 0.00180208
R11641 VDD.n3608 VDD.n3602 0.00180208
R11642 VDD.n4025 VDD.n4024 0.00180208
R11643 VDD.n2838 VDD 0.00180208
R11644 VDD.n3123 VDD 0.00180208
R11645 VDD.n3138 VDD.n3136 0.00180208
R11646 VDD.n728 VDD.n717 0.00180208
R11647 VDD.n1537 VDD.n1536 0.00180208
R11648 VDD.n2041 VDD.n2027 0.00180208
R11649 VDD.n4601 VDD.n4596 0.00180208
R11650 VDD.n4507 VDD.n4493 0.00180208
R11651 VDD.n4380 VDD.n4379 0.00180208
R11652 VDD.n4227 VDD.n4222 0.00180208
R11653 VDD.n328 VDD.n307 0.00180208
R11654 VDD.n342 VDD.n330 0.00180208
R11655 VDD.n356 VDD.n344 0.00180208
R11656 VDD.n370 VDD.n358 0.00180208
R11657 VDD.n384 VDD.n372 0.00180208
R11658 VDD.n398 VDD.n386 0.00180208
R11659 VDD.n412 VDD.n400 0.00180208
R11660 VDD.n781 VDD.n414 0.00180208
R11661 VDD.n1378 VDD.n1377 0.00180208
R11662 VDD.n1396 VDD.n1380 0.00180208
R11663 VDD.n1484 VDD.n1431 0.00180208
R11664 VDD.n1448 VDD.n1447 0.00180208
R11665 VDD.n1450 VDD.n1449 0.00180208
R11666 VDD.n1473 VDD.n1450 0.00180208
R11667 VDD.n1463 VDD.n1451 0.00180208
R11668 VDD.n226 VDD.n225 0.00180208
R11669 VDD.n2168 VDD.n2167 0.00180208
R11670 VDD.n2182 VDD.n2181 0.00180208
R11671 VDD.n2198 VDD.n2197 0.00180208
R11672 VDD.n2212 VDD.n2211 0.00180208
R11673 VDD.n2235 VDD.n2234 0.00180208
R11674 VDD.n2303 VDD.n2302 0.00180208
R11675 VDD.n2321 VDD.n2320 0.00180208
R11676 VDD.n207 VDD.n206 0.00180208
R11677 VDD.n206 VDD.n205 0.00180208
R11678 VDD.n203 VDD.n191 0.00180208
R11679 VDD.n1861 VDD.n1860 0.00180208
R11680 VDD.n1865 VDD.n1864 0.00180208
R11681 VDD.n2395 VDD.n2394 0.00180208
R11682 VDD.n2451 VDD.n2436 0.00180208
R11683 VDD.n2433 VDD.n2421 0.00180208
R11684 VDD.n2419 VDD.n2398 0.00180208
R11685 VDD.n3223 VDD.n3222 0.00180208
R11686 VDD.n1539 VDD.n1538 0.00178866
R11687 VDD.n1540 VDD.n1539 0.00178866
R11688 VDD.n2940 VDD.n2792 0.0017886
R11689 VDD.n4874 VDD.n0 0.00174867
R11690 VDD.n4845 VDD.n164 0.00165296
R11691 VDD.n2770 VDD.n2759 0.00162095
R11692 VDD.n3204 VDD.n3203 0.00162095
R11693 VDD.n752 VDD.n751 0.00161548
R11694 VDD.n3229 VDD.n3209 0.00158092
R11695 VDD.n3273 VDD.n3272 0.00158092
R11696 VDD.n2902 VDD.n2897 0.00148341
R11697 VDD.n2793 VDD.n2725 0.00144949
R11698 VDD.n3520 VDD.n3519 0.00144949
R11699 VDD.n1703 VDD.n1702 0.00143234
R11700 VDD.n3266 VDD.n3265 0.00142078
R11701 VDD.n4110 VDD.n4109 0.00142078
R11702 VDD.n4175 VDD.n4117 0.00142078
R11703 VDD.n4209 VDD.n4208 0.00142078
R11704 VDD.n2143 VDD.n2142 0.00139904
R11705 VDD.n39 VDD.n16 0.00138167
R11706 VDD.n160 VDD.n159 0.00138167
R11707 VDD.n2904 VDD.n2903 0.00132774
R11708 VDD.n1055 VDD.n1054 0.0013158
R11709 VDD.n4417 VDD.n2612 0.00124603
R11710 VDD.n4388 VDD.n4318 0.00124603
R11711 VDD.n4842 VDD.n4841 0.00121212
R11712 VDD.n4813 VDD.n169 0.00121212
R11713 VDD.n3771 VDD.n3756 0.00121212
R11714 VDD.n3767 VDD.n3766 0.00121212
R11715 VDD.n3757 VDD.n2573 0.00121212
R11716 VDD.n4550 VDD.n4543 0.00121212
R11717 VDD.n3555 VDD.n3526 0.00117821
R11718 VDD.n3594 VDD.n3587 0.00117821
R11719 VDD.n760 VDD.n759 0.000999469
R11720 VDD.n753 VDD.n752 0.000999469
R11721 VDD.n919 VDD.n299 0.000999469
R11722 VDD.n1054 VDD.n1053 0.000999469
R11723 VDD.n1707 VDD.n1419 0.000999469
R11724 VDD.n1704 VDD.n1703 0.000999469
R11725 VDD.n1702 VDD.n1701 0.000999469
R11726 VDD.n1701 VDD.n1633 0.000999469
R11727 VDD.n1632 VDD.n1631 0.000999469
R11728 VDD.n1631 VDD.n1626 0.000999469
R11729 VDD.n1625 VDD.n1624 0.000999469
R11730 VDD.n1624 VDD.n1623 0.000999469
R11731 VDD.n1622 VDD.n1621 0.000999469
R11732 VDD.n1621 VDD.n1620 0.000999469
R11733 VDD.n1619 VDD.n1618 0.000999469
R11734 VDD.n2140 VDD.n2139 0.000999469
R11735 VDD.n2139 VDD.n2138 0.000999469
R11736 VDD.n2330 VDD.n186 0.000999469
R11737 VDD.n2330 VDD.n2329 0.000999469
R11738 VDD.n2328 VDD.n2327 0.000999469
R11739 VDD.n1889 VDD.n1888 0.000999469
R11740 VDD.n1887 VDD.n1886 0.000999469
R11741 VDD.n1886 VDD.n1845 0.000999469
R11742 VDD.n1844 VDD.n1843 0.000999469
R11743 VDD.n2377 VDD.n2376 0.000999469
R11744 VDD.n2456 VDD.n2378 0.000999469
R11745 VDD.n2457 VDD.n2456 0.000999469
R11746 VDD.n2479 VDD.n2458 0.000999469
R11747 VDD.n2519 VDD.n2518 0.000999469
R11748 VDD.n4701 VDD.n0 0.000999469
R11749 VDD.n758 VDD.n757 0.00098282
R11750 VDD.n1194 VDD.n285 0.00098282
R11751 VDD.n1193 VDD.n1058 0.00098282
R11752 VDD.n1417 VDD.n1416 0.000949522
R11753 VDD.n2378 VDD.n2377 0.000949522
R11754 VDD.n2327 VDD.n187 0.000916224
R11755 VDD.n1889 VDD.n1814 0.000916224
R11756 VDD.n920 VDD.n919 0.000899575
R11757 VDD.n1842 VDD.n175 0.000899575
R11758 VDD.n1623 VDD.n1622 0.000882926
R11759 VDD.n1845 VDD.n1844 0.000882926
R11760 VDD.n775 VDD.n417 0.000866277
R11761 VDD.n773 VDD.n772 0.000866277
R11762 VDD.n1767 VDD.n1766 0.000866277
R11763 VDD.n2138 VDD.n186 0.000866277
R11764 VDD.n4706 VDD.n2521 0.000849628
R11765 VDD.n768 VDD.n767 0.00081633
R11766 VDD.n765 VDD.n764 0.00081633
R11767 VDD.n762 VDD.n761 0.00081633
R11768 VDD.n756 VDD.n755 0.00081633
R11769 VDD.n754 VDD.n753 0.00081633
R11770 VDD.n933 VDD.n929 0.00081633
R11771 VDD.n932 VDD.n931 0.00081633
R11772 VDD.n1053 VDD.n1052 0.00081633
R11773 VDD.n1050 VDD.n254 0.00081633
R11774 VDD.n1707 VDD.n1706 0.00081633
R11775 VDD.n1705 VDD.n1704 0.00081633
R11776 VDD.n1616 VDD.n1615 0.00081633
R11777 VDD.n2481 VDD.n2480 0.000799681
R11778 VDD VDD.n4873 0.00079375
R11779 VDD.n2148 VDD.n1771 0.000783032
R11780 VDD.n2146 VDD.n2145 0.000783032
R11781 VDD.n750 VDD.n749 0.000766383
R11782 VDD.n748 VDD.n747 0.000766383
R11783 VDD.n751 VDD.n750 0.000733085
R11784 VDD.n749 VDD.n748 0.000733085
R11785 VDD.n747 VDD.n746 0.000733085
R11786 VDD.n1633 VDD.n1632 0.000733085
R11787 VDD.n4705 VDD.n4704 0.000733085
R11788 VDD.n4702 VDD.n4701 0.000733085
R11789 VDD.n922 VDD.n921 0.000716436
R11790 VDD.n4843 VDD.n4842 0.000703463
R11791 VDD.n4814 VDD.n4813 0.000703463
R11792 VDD.n3751 VDD.n3750 0.000703463
R11793 VDD.n2480 VDD.n2479 0.000699787
R11794 VDD.n2518 VDD.n2481 0.000699787
R11795 VDD.n755 VDD.n754 0.000683139
R11796 VDD.n929 VDD.n922 0.000683139
R11797 VDD.n933 VDD.n932 0.000683139
R11798 VDD.n1706 VDD.n1705 0.000683139
R11799 VDD.n1771 VDD.n1770 0.000683139
R11800 VDD.n2147 VDD.n2146 0.000683139
R11801 VDD.n2144 VDD.n2143 0.000683139
R11802 VDD.n2458 VDD.n2457 0.000683139
R11803 VDD.n3582 VDD.n3581 0.000669553
R11804 VDD.n4417 VDD.n4416 0.000669553
R11805 VDD.n4318 VDD.n4317 0.000669553
R11806 VDD.n767 VDD.n766 0.00066649
R11807 VDD.n764 VDD.n763 0.00066649
R11808 VDD.n3269 VDD.n3268 0.000660136
R11809 VDD.n3265 VDD.n2667 0.000660136
R11810 VDD.n4111 VDD.n4110 0.000660136
R11811 VDD.n4117 VDD.n4116 0.000660136
R11812 VDD.n4214 VDD.n4209 0.000660136
R11813 VDD.n2521 VDD.n2520 0.000649841
R11814 VDD.n4706 VDD.n4705 0.000649841
R11815 VDD.n4703 VDD.n4702 0.000649841
R11816 VDD.n1051 VDD.n1050 0.000633192
R11817 VDD.n1617 VDD.n1616 0.000633192
R11818 VDD.n1766 VDD.n242 0.000633192
R11819 VDD.n1768 VDD.n1767 0.000633192
R11820 VDD.n4704 VDD.n4703 0.000616543
R11821 VDD.n3525 VDD.n3524 0.000601732
R11822 VDD.n3526 VDD.n3525 0.000601732
R11823 VDD.n3976 VDD.n3628 0.000601732
R11824 VDD.n3628 VDD.n3594 0.000601732
R11825 VDD.n3585 VDD.n3584 0.000601732
R11826 VDD.n3584 VDD.n3583 0.000601732
R11827 VDD.n3581 VDD.n2612 0.000601732
R11828 VDD.n4416 VDD.n4388 0.000601732
R11829 VDD.n4317 VDD.n4316 0.000601732
R11830 VDD.n4844 VDD.n4843 0.000601732
R11831 VDD.n4841 VDD.n4814 0.000601732
R11832 VDD.n3750 VDD.n169 0.000601732
R11833 VDD.n3755 VDD.n3754 0.000601732
R11834 VDD.n3769 VDD.n3768 0.000601732
R11835 VDD.n3764 VDD.n3763 0.000601732
R11836 VDD.n3761 VDD.n3760 0.000601732
R11837 VDD.n4589 VDD.n2573 0.000601732
R11838 VDD.n4543 VDD.n4542 0.000601732
R11839 VDD.n921 VDD.n920 0.000599894
R11840 VDD.n1843 VDD.n1842 0.000599894
R11841 VDD.n2376 VDD.n175 0.000599894
R11842 VDD.n775 VDD.n774 0.000583245
R11843 VDD.n772 VDD.n771 0.000583245
R11844 VDD.n1814 VDD.n187 0.000583245
R11845 VDD.n2759 VDD.n2758 0.000580068
R11846 VDD.n3203 VDD.n2770 0.000580068
R11847 VDD.n3205 VDD.n3204 0.000580068
R11848 VDD.n3208 VDD.n3207 0.000580068
R11849 VDD.n3314 VDD.n3229 0.000580068
R11850 VDD.n3272 VDD.n3271 0.000580068
R11851 VDD.n3268 VDD.n3267 0.000580068
R11852 VDD.n4084 VDD.n2667 0.000580068
R11853 VDD.n4112 VDD.n4111 0.000580068
R11854 VDD.n4115 VDD.n4114 0.000580068
R11855 VDD.n4215 VDD.n4175 0.000580068
R11856 VDD.n4208 VDD.n4207 0.000580068
R11857 VDD.n2794 VDD.n2793 0.000567821
R11858 VDD.n3519 VDD.n2725 0.000567821
R11859 VDD.n3521 VDD.n3520 0.000567821
R11860 VDD.n3523 VDD.n3522 0.000567821
R11861 VDD.n3524 VDD.n3523 0.000567821
R11862 VDD.n3580 VDD.n3555 0.000567821
R11863 VDD.n3976 VDD.n3580 0.000567821
R11864 VDD.n3587 VDD.n3586 0.000567821
R11865 VDD.n3586 VDD.n3585 0.000567821
R11866 VDD.n3753 VDD.n3752 0.000567821
R11867 VDD.n3754 VDD.n3753 0.000567821
R11868 VDD.n3756 VDD.n3755 0.000567821
R11869 VDD.n3771 VDD.n3770 0.000567821
R11870 VDD.n3770 VDD.n3769 0.000567821
R11871 VDD.n3768 VDD.n3767 0.000567821
R11872 VDD.n3766 VDD.n3765 0.000567821
R11873 VDD.n3765 VDD.n3764 0.000567821
R11874 VDD.n3763 VDD.n3762 0.000567821
R11875 VDD.n3760 VDD.n3759 0.000567821
R11876 VDD.n3759 VDD.n3758 0.000567821
R11877 VDD.n3758 VDD.n3757 0.000567821
R11878 VDD.n4589 VDD.n4588 0.000567821
R11879 VDD.n4588 VDD.n4551 0.000567821
R11880 VDD.n4551 VDD.n4550 0.000567821
R11881 VDD.n4542 VDD.n4541 0.000567821
R11882 VDD.n4541 VDD.n4540 0.000567821
R11883 VDD.n417 VDD.n416 0.000549947
R11884 VDD.n774 VDD.n773 0.000549947
R11885 VDD.n771 VDD.n770 0.000549947
R11886 VDD.n1052 VDD.n1051 0.000549947
R11887 VDD.n1416 VDD.n254 0.000549947
R11888 VDD.n1418 VDD.n1417 0.000549947
R11889 VDD.n1618 VDD.n1617 0.000549947
R11890 VDD.n1615 VDD.n242 0.000549947
R11891 VDD.n3209 VDD.n3208 0.000540034
R11892 VDD.n3314 VDD.n3273 0.000540034
R11893 VDD.n3271 VDD.n3270 0.000540034
R11894 VDD.n3267 VDD.n3266 0.000540034
R11895 VDD.n4109 VDD.n4084 0.000540034
R11896 VDD.n4113 VDD.n4112 0.000540034
R11897 VDD.n4116 VDD.n4115 0.000540034
R11898 VDD.n4215 VDD.n4214 0.000540034
R11899 VDD.n4207 VDD.n4206 0.000540034
R11900 VDD.n2903 VDD.n2902 0.000533911
R11901 VDD.n2897 VDD.n2792 0.000533911
R11902 VDD.n14 VDD.n13 0.000533911
R11903 VDD.n15 VDD.n14 0.000533911
R11904 VDD.n16 VDD.n15 0.000533911
R11905 VDD.n93 VDD.n39 0.000533911
R11906 VDD.n137 VDD.n93 0.000533911
R11907 VDD.n154 VDD.n137 0.000533911
R11908 VDD.n159 VDD.n154 0.000533911
R11909 VDD.n161 VDD.n160 0.000533911
R11910 VDD.n162 VDD.n161 0.000533911
R11911 VDD.n163 VDD.n162 0.000533911
R11912 VDD.n164 VDD.n163 0.000533911
R11913 VDD.n1770 VDD.n1769 0.000533298
R11914 VDD.n2148 VDD.n2147 0.000533298
R11915 VDD.n2145 VDD.n2144 0.000533298
R11916 VDD.n769 VDD.n768 0.000516649
R11917 VDD.n766 VDD.n765 0.000516649
R11918 VDD.n763 VDD.n762 0.000516649
R11919 VDD.n759 VDD.n758 0.000516649
R11920 VDD.n757 VDD.n756 0.000516649
R11921 VDD.n930 VDD.n285 0.000516649
R11922 VDD.n1194 VDD.n1193 0.000516649
R11923 VDD.n1058 VDD.n1057 0.000516649
R11924 x2.X.n138 x2.X.t47 396.834
R11925 x2.X.n117 x2.X.t49 396.834
R11926 x2.X.n96 x2.X.t42 396.834
R11927 x2.X.n75 x2.X.t37 396.834
R11928 x2.X.n54 x2.X.t68 396.834
R11929 x2.X.n33 x2.X.t66 396.834
R11930 x2.X.n13 x2.X.t52 396.834
R11931 x2.X.n133 x2.X.t35 381.228
R11932 x2.X.n112 x2.X.t33 381.228
R11933 x2.X.n91 x2.X.t60 381.228
R11934 x2.X.n70 x2.X.t58 381.228
R11935 x2.X.n49 x2.X.t39 381.228
R11936 x2.X.n28 x2.X.t72 381.228
R11937 x2.X.n8 x2.X.t69 381.228
R11938 x2.X.n127 x2.X.t44 198.335
R11939 x2.X.n106 x2.X.t32 198.335
R11940 x2.X.n85 x2.X.t71 198.335
R11941 x2.X.n64 x2.X.t56 198.335
R11942 x2.X.n43 x2.X.t54 198.335
R11943 x2.X.n23 x2.X.t50 198.335
R11944 x2.X.n148 x2.X.t34 198.025
R11945 x2.X.n149 x2.X.t53 172.463
R11946 x2.X.n128 x2.X.t62 171.875
R11947 x2.X.n107 x2.X.t48 171.875
R11948 x2.X.n86 x2.X.t41 171.875
R11949 x2.X.n65 x2.X.t73 171.875
R11950 x2.X.n44 x2.X.t70 171.875
R11951 x2.X.n24 x2.X.t65 171.875
R11952 x2.X.n135 x2.X.n134 152
R11953 x2.X.n114 x2.X.n113 152
R11954 x2.X.n93 x2.X.n92 152
R11955 x2.X.n72 x2.X.n71 152
R11956 x2.X.n51 x2.X.n50 152
R11957 x2.X.n30 x2.X.n29 152
R11958 x2.X.n10 x2.X.n9 152
R11959 x2.X.n161 x2.X.n160 146.812
R11960 x2.X.n135 x2.X.t64 136.745
R11961 x2.X.n114 x2.X.t61 136.745
R11962 x2.X.n93 x2.X.t46 136.745
R11963 x2.X.n72 x2.X.t38 136.745
R11964 x2.X.n51 x2.X.t59 136.745
R11965 x2.X.n30 x2.X.t57 136.745
R11966 x2.X.n10 x2.X.t55 136.745
R11967 x2.X.n138 x2.X.t43 134.065
R11968 x2.X.n117 x2.X.t45 134.065
R11969 x2.X.n96 x2.X.t40 134.065
R11970 x2.X.n75 x2.X.t36 134.065
R11971 x2.X.n54 x2.X.t67 134.065
R11972 x2.X.n33 x2.X.t63 134.065
R11973 x2.X.n13 x2.X.t51 134.065
R11974 x2.X.n167 x2.X.n153 108.412
R11975 x2.X.n166 x2.X.n154 108.412
R11976 x2.X.n165 x2.X.n155 108.412
R11977 x2.X.n164 x2.X.n156 108.412
R11978 x2.X.n163 x2.X.n157 108.412
R11979 x2.X.n162 x2.X.n158 108.412
R11980 x2.X.n161 x2.X.n159 108.412
R11981 x2.X.n171 x2.X.n169 90.8321
R11982 x2.X.n133 x2.X.n132 75.1188
R11983 x2.X.n112 x2.X.n111 75.1188
R11984 x2.X.n91 x2.X.n90 75.1188
R11985 x2.X.n70 x2.X.n69 75.1188
R11986 x2.X.n49 x2.X.n48 75.1188
R11987 x2.X.n28 x2.X.n27 75.1188
R11988 x2.X.n8 x2.X.n7 75.1188
R11989 x2.X.n171 x2.X.n170 52.4321
R11990 x2.X.n173 x2.X.n172 52.4321
R11991 x2.X.n175 x2.X.n174 52.4321
R11992 x2.X.n177 x2.X.n176 52.4321
R11993 x2.X.n179 x2.X.n178 52.4321
R11994 x2.X.n181 x2.X.n180 52.4321
R11995 x2.X.n183 x2.X.n182 52.4321
R11996 x2.X x2.X.n183 40.4711
R11997 x2.X.n173 x2.X.n171 38.4005
R11998 x2.X.n175 x2.X.n173 38.4005
R11999 x2.X.n177 x2.X.n175 38.4005
R12000 x2.X.n179 x2.X.n177 38.4005
R12001 x2.X.n181 x2.X.n179 38.4005
R12002 x2.X.n183 x2.X.n181 38.4005
R12003 x2.X.n167 x2.X.n166 38.4005
R12004 x2.X.n166 x2.X.n165 38.4005
R12005 x2.X.n165 x2.X.n164 38.4005
R12006 x2.X.n164 x2.X.n163 38.4005
R12007 x2.X.n163 x2.X.n162 38.4005
R12008 x2.X.n162 x2.X.n161 38.4005
R12009 x2.X x2.X.n167 33.7342
R12010 x2.X.n168 x2.X.n152 26.8074
R12011 x2.X.n153 x2.X.t3 26.5955
R12012 x2.X.n153 x2.X.t14 26.5955
R12013 x2.X.n154 x2.X.t8 26.5955
R12014 x2.X.n154 x2.X.t13 26.5955
R12015 x2.X.n155 x2.X.t6 26.5955
R12016 x2.X.n155 x2.X.t11 26.5955
R12017 x2.X.n156 x2.X.t4 26.5955
R12018 x2.X.n156 x2.X.t10 26.5955
R12019 x2.X.n157 x2.X.t2 26.5955
R12020 x2.X.n157 x2.X.t1 26.5955
R12021 x2.X.n158 x2.X.t9 26.5955
R12022 x2.X.n158 x2.X.t0 26.5955
R12023 x2.X.n159 x2.X.t7 26.5955
R12024 x2.X.n159 x2.X.t12 26.5955
R12025 x2.X.n160 x2.X.t5 26.5955
R12026 x2.X.n160 x2.X.t15 26.5955
R12027 x2.X.n169 x2.X.t27 24.9236
R12028 x2.X.n169 x2.X.t21 24.9236
R12029 x2.X.n170 x2.X.t29 24.9236
R12030 x2.X.n170 x2.X.t18 24.9236
R12031 x2.X.n172 x2.X.t31 24.9236
R12032 x2.X.n172 x2.X.t22 24.9236
R12033 x2.X.n174 x2.X.t24 24.9236
R12034 x2.X.n174 x2.X.t23 24.9236
R12035 x2.X.n176 x2.X.t26 24.9236
R12036 x2.X.n176 x2.X.t16 24.9236
R12037 x2.X.n178 x2.X.t28 24.9236
R12038 x2.X.n178 x2.X.t17 24.9236
R12039 x2.X.n180 x2.X.t30 24.9236
R12040 x2.X.n180 x2.X.t19 24.9236
R12041 x2.X.n182 x2.X.t25 24.9236
R12042 x2.X.n182 x2.X.t20 24.9236
R12043 x2.X.n140 x2.X 13.6005
R12044 x2.X.n119 x2.X 13.6005
R12045 x2.X.n98 x2.X 13.6005
R12046 x2.X.n77 x2.X 13.6005
R12047 x2.X.n56 x2.X 13.6005
R12048 x2.X.n35 x2.X 13.6005
R12049 x2.X.n15 x2.X 13.6005
R12050 x2.X.n135 x2.X.n133 13.3692
R12051 x2.X.n114 x2.X.n112 13.3692
R12052 x2.X.n93 x2.X.n91 13.3692
R12053 x2.X.n72 x2.X.n70 13.3692
R12054 x2.X.n51 x2.X.n49 13.3692
R12055 x2.X.n30 x2.X.n28 13.3692
R12056 x2.X.n10 x2.X.n8 13.3692
R12057 x2.X.n47 x2.X.n26 13.2412
R12058 x2.X.n152 x2.X.n151 11.2004
R12059 x2.X.n134 x2.X 11.055
R12060 x2.X.n113 x2.X 11.055
R12061 x2.X.n92 x2.X 11.055
R12062 x2.X.n71 x2.X 11.055
R12063 x2.X.n50 x2.X 11.055
R12064 x2.X.n29 x2.X 11.055
R12065 x2.X.n9 x2.X 11.055
R12066 x2.X.n136 x2.X.n135 9.3005
R12067 x2.X.n150 x2.X.n149 9.3005
R12068 x2.X.n115 x2.X.n114 9.3005
R12069 x2.X.n129 x2.X.n128 9.3005
R12070 x2.X.n94 x2.X.n93 9.3005
R12071 x2.X.n108 x2.X.n107 9.3005
R12072 x2.X.n73 x2.X.n72 9.3005
R12073 x2.X.n87 x2.X.n86 9.3005
R12074 x2.X.n52 x2.X.n51 9.3005
R12075 x2.X.n66 x2.X.n65 9.3005
R12076 x2.X.n31 x2.X.n30 9.3005
R12077 x2.X.n45 x2.X.n44 9.3005
R12078 x2.X.n11 x2.X.n10 9.3005
R12079 x2.X.n25 x2.X.n24 9.3005
R12080 x2.X.n151 x2.X.n150 9.23046
R12081 x2.X.n46 x2.X.n45 9.10496
R12082 x2.X.n26 x2.X.n25 9.10496
R12083 x2.X.n109 x2.X.n108 9.10363
R12084 x2.X.n88 x2.X.n87 9.10363
R12085 x2.X.n67 x2.X.n66 9.1023
R12086 x2.X.n130 x2.X.n129 8.98032
R12087 x2.X.n168 x2.X 8.75839
R12088 x2.X.n89 x2.X.n68 8.70611
R12089 x2.X.n68 x2.X.n47 8.70243
R12090 x2.X.n131 x2.X.n110 8.70243
R12091 x2.X.n110 x2.X.n89 8.69014
R12092 x2.X.n139 x2.X.n138 6.98562
R12093 x2.X.n118 x2.X.n117 6.98562
R12094 x2.X.n97 x2.X.n96 6.98562
R12095 x2.X.n76 x2.X.n75 6.98562
R12096 x2.X.n55 x2.X.n54 6.98562
R12097 x2.X.n34 x2.X.n33 6.98562
R12098 x2.X.n14 x2.X.n13 6.98562
R12099 x2.X.n128 x2.X.n127 5.7706
R12100 x2.X.n107 x2.X.n106 5.7706
R12101 x2.X.n86 x2.X.n85 5.7706
R12102 x2.X.n65 x2.X.n64 5.7706
R12103 x2.X.n44 x2.X.n43 5.7706
R12104 x2.X.n24 x2.X.n23 5.7706
R12105 x2.X.n149 x2.X.n148 5.46089
R12106 x2.X.n131 x2.X.n130 4.53188
R12107 x2.X.n110 x2.X.n109 4.53188
R12108 x2.X.n89 x2.X.n88 4.53188
R12109 x2.X.n68 x2.X.n67 4.53188
R12110 x2.X.n47 x2.X.n46 4.53188
R12111 x2.X.n0 x2.X.n141 4.46483
R12112 x2.X.n1 x2.X.n120 4.46483
R12113 x2.X.n2 x2.X.n99 4.46483
R12114 x2.X.n3 x2.X.n78 4.46483
R12115 x2.X.n4 x2.X.n57 4.46483
R12116 x2.X.n5 x2.X.n36 4.46483
R12117 x2.X.n6 x2.X.n16 4.46483
R12118 x2.X.n126 x2.X.n125 4.17441
R12119 x2.X.n105 x2.X.n104 4.17441
R12120 x2.X.n63 x2.X.n62 4.17441
R12121 x2.X.n22 x2.X.n21 4.17441
R12122 x2.X.n147 x2.X.n146 3.89615
R12123 x2.X.n84 x2.X.n83 3.89615
R12124 x2.X.n42 x2.X.n41 3.89615
R12125 x2.X.n134 x2.X.n132 2.90959
R12126 x2.X.n113 x2.X.n111 2.90959
R12127 x2.X.n92 x2.X.n90 2.90959
R12128 x2.X.n71 x2.X.n69 2.90959
R12129 x2.X.n50 x2.X.n48 2.90959
R12130 x2.X.n29 x2.X.n27 2.90959
R12131 x2.X.n9 x2.X.n7 2.90959
R12132 x2.X.n141 x2.X 2.89456
R12133 x2.X.n120 x2.X 2.89456
R12134 x2.X.n99 x2.X 2.89456
R12135 x2.X.n78 x2.X 2.89456
R12136 x2.X.n57 x2.X 2.89456
R12137 x2.X.n36 x2.X 2.89456
R12138 x2.X.n16 x2.X 2.89456
R12139 x2.X x2.X.n136 2.75432
R12140 x2.X x2.X.n115 2.75432
R12141 x2.X x2.X.n94 2.75432
R12142 x2.X x2.X.n73 2.75432
R12143 x2.X x2.X.n52 2.75432
R12144 x2.X x2.X.n31 2.75432
R12145 x2.X x2.X.n11 2.75432
R12146 x2.X x2.X.n168 2.69524
R12147 x2.X.n140 x2.X.n139 2.52171
R12148 x2.X.n119 x2.X.n118 2.52171
R12149 x2.X.n98 x2.X.n97 2.52171
R12150 x2.X.n77 x2.X.n76 2.52171
R12151 x2.X.n56 x2.X.n55 2.52171
R12152 x2.X.n35 x2.X.n34 2.52171
R12153 x2.X.n15 x2.X.n14 2.52171
R12154 x2.X.n146 x2.X 2.50485
R12155 x2.X.n83 x2.X 2.50485
R12156 x2.X.n41 x2.X 2.50485
R12157 x2.X.n151 x2.X.n145 2.2505
R12158 x2.X.n130 x2.X.n124 2.2505
R12159 x2.X.n109 x2.X.n103 2.2505
R12160 x2.X.n88 x2.X.n82 2.2505
R12161 x2.X.n67 x2.X.n61 2.2505
R12162 x2.X.n46 x2.X.n40 2.2505
R12163 x2.X.n26 x2.X.n20 2.2505
R12164 x2.X.n125 x2.X 2.22659
R12165 x2.X.n104 x2.X 2.22659
R12166 x2.X.n62 x2.X 2.22659
R12167 x2.X.n21 x2.X 2.22659
R12168 x2.X.n152 x2.X.n131 1.94561
R12169 x2.X.n137 x2.X 1.89782
R12170 x2.X.n53 x2.X 1.89782
R12171 x2.X.n32 x2.X 1.89782
R12172 x2.X.n12 x2.X 1.89782
R12173 x2.X.n116 x2.X 1.89336
R12174 x2.X.n95 x2.X 1.89336
R12175 x2.X.n74 x2.X 1.89336
R12176 x2.X.n116 x2.X 1.45586
R12177 x2.X.n95 x2.X 1.45586
R12178 x2.X.n74 x2.X 1.45586
R12179 x2.X.n137 x2.X 1.45139
R12180 x2.X.n53 x2.X 1.45139
R12181 x2.X.n32 x2.X 1.45139
R12182 x2.X.n12 x2.X 1.45139
R12183 x2.X.n123 x2.X.n122 0.955857
R12184 x2.X.n102 x2.X.n101 0.955857
R12185 x2.X.n81 x2.X.n80 0.955857
R12186 x2.X.n144 x2.X.n143 0.951393
R12187 x2.X.n60 x2.X.n59 0.951393
R12188 x2.X.n39 x2.X.n38 0.951393
R12189 x2.X.n19 x2.X.n18 0.951393
R12190 x2.X.n150 x2.X.n147 0.835283
R12191 x2.X.n87 x2.X.n84 0.835283
R12192 x2.X.n45 x2.X.n42 0.835283
R12193 x2.X.n129 x2.X.n126 0.557022
R12194 x2.X.n108 x2.X.n105 0.557022
R12195 x2.X.n66 x2.X.n63 0.557022
R12196 x2.X.n25 x2.X.n22 0.557022
R12197 x2.X.n123 x2.X 0.53175
R12198 x2.X.n102 x2.X 0.53175
R12199 x2.X.n81 x2.X 0.53175
R12200 x2.X.n144 x2.X 0.529797
R12201 x2.X.n39 x2.X 0.529797
R12202 x2.X.n19 x2.X 0.529797
R12203 x2.X.n60 x2.X 0.513758
R12204 x2.X.n136 x2.X.n132 0.388379
R12205 x2.X.n115 x2.X.n111 0.388379
R12206 x2.X.n94 x2.X.n90 0.388379
R12207 x2.X.n73 x2.X.n69 0.388379
R12208 x2.X.n52 x2.X.n48 0.388379
R12209 x2.X.n31 x2.X.n27 0.388379
R12210 x2.X.n11 x2.X.n7 0.388379
R12211 x2.X.n141 x2.X.n140 0.373349
R12212 x2.X.n120 x2.X.n119 0.373349
R12213 x2.X.n99 x2.X.n98 0.373349
R12214 x2.X.n78 x2.X.n77 0.373349
R12215 x2.X.n57 x2.X.n56 0.373349
R12216 x2.X.n36 x2.X.n35 0.373349
R12217 x2.X.n16 x2.X.n15 0.373349
R12218 x2.X.n143 x2.X 0.259429
R12219 x2.X.n122 x2.X 0.259429
R12220 x2.X.n101 x2.X 0.259429
R12221 x2.X.n80 x2.X 0.259429
R12222 x2.X.n59 x2.X 0.259429
R12223 x2.X.n38 x2.X 0.259429
R12224 x2.X.n18 x2.X 0.259429
R12225 x2.X.n143 x2.X.n0 0.076587
R12226 x2.X.n122 x2.X.n1 0.076587
R12227 x2.X.n101 x2.X.n2 0.076587
R12228 x2.X.n80 x2.X.n3 0.076587
R12229 x2.X.n59 x2.X.n4 0.076587
R12230 x2.X.n38 x2.X.n5 0.076587
R12231 x2.X.n18 x2.X.n6 0.076587
R12232 x2.X.n145 x2.X.n137 0.0532344
R12233 x2.X.n145 x2.X.n144 0.0532344
R12234 x2.X.n124 x2.X.n116 0.0532344
R12235 x2.X.n124 x2.X.n123 0.0532344
R12236 x2.X.n103 x2.X.n95 0.0532344
R12237 x2.X.n103 x2.X.n102 0.0532344
R12238 x2.X.n82 x2.X.n74 0.0532344
R12239 x2.X.n82 x2.X.n81 0.0532344
R12240 x2.X.n40 x2.X.n32 0.0532344
R12241 x2.X.n40 x2.X.n39 0.0532344
R12242 x2.X.n20 x2.X.n12 0.0532344
R12243 x2.X.n20 x2.X.n19 0.0532344
R12244 x2.X.n61 x2.X.n53 0.0516364
R12245 x2.X.n61 x2.X.n60 0.0516364
R12246 x2.X.n6 x2.X.n17 0.0466957
R12247 x2.X.n5 x2.X.n37 0.0466957
R12248 x2.X.n4 x2.X.n58 0.0466957
R12249 x2.X.n3 x2.X.n79 0.0466957
R12250 x2.X.n2 x2.X.n100 0.0466957
R12251 x2.X.n1 x2.X.n121 0.0466957
R12252 x2.X.n0 x2.X.n142 0.0466957
R12253 x2.X.n142 x2.X 0.0358261
R12254 x2.X.n121 x2.X 0.0358261
R12255 x2.X.n100 x2.X 0.0358261
R12256 x2.X.n79 x2.X 0.0358261
R12257 x2.X.n58 x2.X 0.0358261
R12258 x2.X.n37 x2.X 0.0358261
R12259 x2.X.n17 x2.X 0.0358261
R12260 x9.A1.n88 x9.A1.t41 327.974
R12261 x9.A1.n105 x9.A1.t45 327.961
R12262 x9.A1.n121 x9.A1.t47 327.961
R12263 x9.A1.n137 x9.A1.t38 327.599
R12264 x9.A1.n70 x9.A1.t58 327.584
R12265 x9.A1.n34 x9.A1.t43 327.584
R12266 x9.A1.n52 x9.A1.t56 327.57
R12267 x9.A1.n76 x9.A1.t34 327.361
R12268 x9.A1.n40 x9.A1.t53 327.361
R12269 x9.A1.n110 x9.A1.t46 327.337
R12270 x9.A1.n126 x9.A1.t39 327.337
R12271 x9.A1.n94 x9.A1.t51 326.986
R12272 x9.A1.n58 x9.A1.t48 326.986
R12273 x9.A1.n23 x9.A1.t42 326.986
R12274 x9.A1.n50 x9.A1.t44 151.681
R12275 x9.A1.n103 x9.A1.t36 150.825
R12276 x9.A1.n119 x9.A1.t37 150.825
R12277 x9.A1.n86 x9.A1.t59 150.81
R12278 x9.A1.n68 x9.A1.t57 150.794
R12279 x9.A1.n32 x9.A1.t32 150.794
R12280 x9.A1.n111 x9.A1.t49 150.78
R12281 x9.A1.n127 x9.A1.t50 150.78
R12282 x9.A1.n135 x9.A1.t52 150.78
R12283 x9.A1.n77 x9.A1.t33 149.893
R12284 x9.A1.n41 x9.A1.t40 149.893
R12285 x9.A1.n95 x9.A1.t54 149.862
R12286 x9.A1.n59 x9.A1.t35 149.862
R12287 x9.A1.n24 x9.A1.t55 149.862
R12288 x9.A1.n10 x9.A1.n8 146.811
R12289 x9.A1.n20 x9.A1.n19 108.412
R12290 x9.A1.n21 x9.A1.n7 108.412
R12291 x9.A1.n10 x9.A1.n9 108.412
R12292 x9.A1.n12 x9.A1.n11 108.412
R12293 x9.A1.n14 x9.A1.n13 108.412
R12294 x9.A1.n16 x9.A1.n15 108.412
R12295 x9.A1.n18 x9.A1.n17 108.412
R12296 x9.A1.n150 x9.A1.n148 90.8321
R12297 x9.A1.n150 x9.A1.n149 52.4321
R12298 x9.A1.n152 x9.A1.n151 52.4321
R12299 x9.A1.n154 x9.A1.n153 52.4321
R12300 x9.A1.n156 x9.A1.n155 52.4321
R12301 x9.A1.n158 x9.A1.n157 52.4321
R12302 x9.A1.n160 x9.A1.n159 52.4321
R12303 x9.A1.n162 x9.A1.n161 52.4321
R12304 x9.A1 x9.A1.n162 40.4711
R12305 x9.A1.n152 x9.A1.n150 38.4005
R12306 x9.A1.n154 x9.A1.n152 38.4005
R12307 x9.A1.n156 x9.A1.n154 38.4005
R12308 x9.A1.n158 x9.A1.n156 38.4005
R12309 x9.A1.n160 x9.A1.n158 38.4005
R12310 x9.A1.n162 x9.A1.n160 38.4005
R12311 x9.A1.n12 x9.A1.n10 38.4005
R12312 x9.A1.n14 x9.A1.n12 38.4005
R12313 x9.A1.n16 x9.A1.n14 38.4005
R12314 x9.A1.n18 x9.A1.n16 38.4005
R12315 x9.A1.n20 x9.A1.n18 38.4005
R12316 x9.A1.n21 x9.A1.n20 38.4005
R12317 x9.A1 x9.A1.n21 33.7342
R12318 x9.A1.n95 x9.A1 29.1167
R12319 x9.A1.n59 x9.A1 29.1167
R12320 x9.A1.n24 x9.A1 29.1167
R12321 x9.A1.n77 x9.A1 28.9113
R12322 x9.A1.n41 x9.A1 28.9113
R12323 x9.A1.n111 x9.A1 28.5657
R12324 x9.A1.n127 x9.A1 28.5657
R12325 x9.A1.n135 x9.A1 28.5657
R12326 x9.A1.n86 x9.A1 28.3628
R12327 x9.A1.n68 x9.A1 28.246
R12328 x9.A1.n32 x9.A1 28.246
R12329 x9.A1.n103 x9.A1 28.0462
R12330 x9.A1.n119 x9.A1 28.0462
R12331 x9.A1.n50 x9.A1 27.901
R12332 x9.A1.n7 x9.A1.t8 26.5955
R12333 x9.A1.n7 x9.A1.t2 26.5955
R12334 x9.A1.n8 x9.A1.t12 26.5955
R12335 x9.A1.n8 x9.A1.t4 26.5955
R12336 x9.A1.n9 x9.A1.t11 26.5955
R12337 x9.A1.n9 x9.A1.t6 26.5955
R12338 x9.A1.n11 x9.A1.t14 26.5955
R12339 x9.A1.n11 x9.A1.t0 26.5955
R12340 x9.A1.n13 x9.A1.t9 26.5955
R12341 x9.A1.n13 x9.A1.t1 26.5955
R12342 x9.A1.n15 x9.A1.t10 26.5955
R12343 x9.A1.n15 x9.A1.t3 26.5955
R12344 x9.A1.n17 x9.A1.t13 26.5955
R12345 x9.A1.n17 x9.A1.t5 26.5955
R12346 x9.A1.n19 x9.A1.t15 26.5955
R12347 x9.A1.n19 x9.A1.t7 26.5955
R12348 x9.A1.n148 x9.A1.t20 24.9236
R12349 x9.A1.n148 x9.A1.t28 24.9236
R12350 x9.A1.n149 x9.A1.t19 24.9236
R12351 x9.A1.n149 x9.A1.t30 24.9236
R12352 x9.A1.n151 x9.A1.t22 24.9236
R12353 x9.A1.n151 x9.A1.t24 24.9236
R12354 x9.A1.n153 x9.A1.t17 24.9236
R12355 x9.A1.n153 x9.A1.t25 24.9236
R12356 x9.A1.n155 x9.A1.t18 24.9236
R12357 x9.A1.n155 x9.A1.t27 24.9236
R12358 x9.A1.n157 x9.A1.t21 24.9236
R12359 x9.A1.n157 x9.A1.t29 24.9236
R12360 x9.A1.n159 x9.A1.t23 24.9236
R12361 x9.A1.n159 x9.A1.t31 24.9236
R12362 x9.A1.n161 x9.A1.t16 24.9236
R12363 x9.A1.n161 x9.A1.t26 24.9236
R12364 x9.A1.n147 x9.A1.n146 11.2712
R12365 x9.A1.n147 x9.A1 8.42155
R12366 x9.A1.n38 x9.A1.n30 8.31458
R12367 x9.A1.n141 x9.A1.n140 8.3109
R12368 x9.A1.n74 x9.A1.n66 4.55989
R12369 x9.A1.n143 x9.A1.n142 4.55254
R12370 x9.A1.n92 x9.A1.n84 4.55254
R12371 x9.A1.n145 x9.A1.n144 4.54886
R12372 x9.A1.n56 x9.A1.n48 4.54886
R12373 x9.A1.n48 x9.A1.n38 4.07827
R12374 x9.A1.n142 x9.A1.n141 4.07459
R12375 x9.A1.n144 x9.A1.n143 4.07459
R12376 x9.A1.n84 x9.A1.n74 4.07092
R12377 x9.A1.n66 x9.A1.n56 4.06724
R12378 x9.A1.n145 x9.A1.n101 3.75519
R12379 x9.A1.n144 x9.A1.n108 3.75519
R12380 x9.A1.n143 x9.A1.n117 3.75519
R12381 x9.A1.n142 x9.A1.n124 3.75519
R12382 x9.A1.n141 x9.A1.n133 3.75519
R12383 x9.A1.n92 x9.A1.n91 3.75519
R12384 x9.A1.n84 x9.A1.n83 3.75519
R12385 x9.A1.n74 x9.A1.n73 3.75519
R12386 x9.A1.n66 x9.A1.n65 3.75519
R12387 x9.A1.n56 x9.A1.n55 3.75519
R12388 x9.A1.n48 x9.A1.n47 3.75519
R12389 x9.A1.n38 x9.A1.n37 3.75519
R12390 x9.A1.n138 x9.A1.n137 3.44665
R12391 x9.A1.n89 x9.A1.n88 3.44665
R12392 x9.A1.n106 x9.A1.n105 3.38163
R12393 x9.A1.n122 x9.A1.n121 3.38163
R12394 x9.A1.n71 x9.A1.n70 3.38163
R12395 x9.A1.n35 x9.A1.n34 3.38163
R12396 x9.A1.n53 x9.A1.n52 3.31902
R12397 x9.A1.n146 x9.A1.n145 3.25601
R12398 x9.A1.n98 x9.A1.n97 3.03311
R12399 x9.A1.n0 x9.A1.n106 3.03311
R12400 x9.A1.n114 x9.A1.n113 3.03311
R12401 x9.A1.n1 x9.A1.n122 3.03311
R12402 x9.A1.n130 x9.A1.n129 3.03311
R12403 x9.A1.n2 x9.A1.n138 3.03311
R12404 x9.A1.n3 x9.A1.n89 3.03311
R12405 x9.A1.n80 x9.A1.n79 3.03311
R12406 x9.A1.n4 x9.A1.n71 3.03311
R12407 x9.A1.n62 x9.A1.n61 3.03311
R12408 x9.A1.n5 x9.A1.n53 3.03311
R12409 x9.A1.n44 x9.A1.n43 3.03311
R12410 x9.A1.n6 x9.A1.n35 3.03311
R12411 x9.A1.n27 x9.A1.n26 3.03311
R12412 x9.A1 x9.A1.n147 3.03208
R12413 x9.A1.n97 x9.A1.n94 3.01226
R12414 x9.A1.n79 x9.A1.n76 3.01226
R12415 x9.A1.n61 x9.A1.n58 3.01226
R12416 x9.A1.n43 x9.A1.n40 3.01226
R12417 x9.A1.n26 x9.A1.n23 3.01226
R12418 x9.A1.n113 x9.A1.n110 2.95435
R12419 x9.A1.n129 x9.A1.n126 2.95435
R12420 x9.A1.n107 x9.A1.n0 1.50871
R12421 x9.A1.n123 x9.A1.n1 1.50871
R12422 x9.A1.n139 x9.A1.n2 1.50871
R12423 x9.A1.n90 x9.A1.n3 1.50871
R12424 x9.A1.n72 x9.A1.n4 1.50871
R12425 x9.A1.n54 x9.A1.n5 1.50871
R12426 x9.A1.n36 x9.A1.n6 1.50871
R12427 x9.A1.n100 x9.A1.n99 1.50153
R12428 x9.A1.n116 x9.A1.n115 1.50153
R12429 x9.A1.n132 x9.A1.n131 1.50153
R12430 x9.A1.n82 x9.A1.n81 1.50153
R12431 x9.A1.n64 x9.A1.n63 1.50153
R12432 x9.A1.n46 x9.A1.n45 1.50153
R12433 x9.A1.n29 x9.A1.n28 1.50153
R12434 x9.A1.n97 x9.A1.n96 1.2554
R12435 x9.A1.n79 x9.A1.n78 1.2554
R12436 x9.A1.n61 x9.A1.n60 1.2554
R12437 x9.A1.n43 x9.A1.n42 1.2554
R12438 x9.A1.n26 x9.A1.n25 1.2554
R12439 x9.A1.n113 x9.A1.n112 1.23127
R12440 x9.A1.n129 x9.A1.n128 1.23127
R12441 x9.A1.n146 x9.A1.n92 0.741309
R12442 x9.A1.n138 x9.A1.n136 0.738962
R12443 x9.A1.n89 x9.A1.n87 0.738962
R12444 x9.A1.n106 x9.A1.n104 0.725028
R12445 x9.A1.n122 x9.A1.n120 0.725028
R12446 x9.A1.n71 x9.A1.n69 0.725028
R12447 x9.A1.n35 x9.A1.n33 0.725028
R12448 x9.A1.n53 x9.A1.n51 0.711611
R12449 x9.A1.n96 x9.A1.n95 0.213762
R12450 x9.A1.n60 x9.A1.n59 0.213762
R12451 x9.A1.n25 x9.A1.n24 0.213762
R12452 x9.A1.n78 x9.A1.n77 0.178608
R12453 x9.A1.n42 x9.A1.n41 0.178608
R12454 x9.A1.n112 x9.A1.n111 0.178047
R12455 x9.A1.n128 x9.A1.n127 0.178047
R12456 x9.A1.n136 x9.A1.n135 0.178047
R12457 x9.A1.n69 x9.A1.n68 0.161787
R12458 x9.A1.n33 x9.A1.n32 0.161787
R12459 x9.A1.n51 x9.A1.n50 0.161251
R12460 x9.A1.n87 x9.A1.n86 0.143169
R12461 x9.A1.n104 x9.A1.n103 0.127479
R12462 x9.A1.n120 x9.A1.n119 0.127479
R12463 x9.A1.n6 x9.A1.n31 0.0373802
R12464 x9.A1.n5 x9.A1.n49 0.0373802
R12465 x9.A1.n4 x9.A1.n67 0.0373802
R12466 x9.A1.n3 x9.A1.n85 0.0373802
R12467 x9.A1.n2 x9.A1.n134 0.0373802
R12468 x9.A1.n1 x9.A1.n118 0.0373802
R12469 x9.A1.n0 x9.A1.n102 0.0373802
R12470 x9.A1.n101 x9.A1.n100 0.0226928
R12471 x9.A1.n108 x9.A1.n107 0.0226928
R12472 x9.A1.n117 x9.A1.n116 0.0226928
R12473 x9.A1.n124 x9.A1.n123 0.0226928
R12474 x9.A1.n133 x9.A1.n132 0.0226928
R12475 x9.A1.n140 x9.A1.n139 0.0226928
R12476 x9.A1.n91 x9.A1.n90 0.0226928
R12477 x9.A1.n83 x9.A1.n82 0.0226928
R12478 x9.A1.n73 x9.A1.n72 0.0226928
R12479 x9.A1.n65 x9.A1.n64 0.0226928
R12480 x9.A1.n55 x9.A1.n54 0.0226928
R12481 x9.A1.n47 x9.A1.n46 0.0226928
R12482 x9.A1.n37 x9.A1.n36 0.0226928
R12483 x9.A1.n30 x9.A1.n29 0.0226928
R12484 x9.A1.n98 x9.A1.n93 0.0125192
R12485 x9.A1.n114 x9.A1.n109 0.0125192
R12486 x9.A1.n130 x9.A1.n125 0.0125192
R12487 x9.A1.n80 x9.A1.n75 0.0125192
R12488 x9.A1.n62 x9.A1.n57 0.0125192
R12489 x9.A1.n44 x9.A1.n39 0.0125192
R12490 x9.A1.n27 x9.A1.n22 0.0125192
R12491 x9.A1.n99 x9.A1.n98 0.0109043
R12492 x9.A1.n115 x9.A1.n114 0.0109043
R12493 x9.A1.n131 x9.A1.n130 0.0109043
R12494 x9.A1.n81 x9.A1.n80 0.0109043
R12495 x9.A1.n63 x9.A1.n62 0.0109043
R12496 x9.A1.n45 x9.A1.n44 0.0109043
R12497 x9.A1.n28 x9.A1.n27 0.0109043
R12498 VSS_SW_b[3].n4 VSS_SW_b[3].n3 641.827
R12499 VSS_SW_b[3] VSS_SW_b[3].t0 422.656
R12500 VSS_SW_b[3].t0 VSS_SW_b[3].n5 121.231
R12501 VSS_SW_b[3].n2 VSS_SW_b[3].t1 117.424
R12502 VSS_SW_b[3].n3 VSS_SW_b[3].n2 77.418
R12503 VSS_SW_b[3].n6 VSS_SW_b[3] 11.3827
R12504 VSS_SW_b[3].n5 VSS_SW_b[3].n0 9.15497
R12505 VSS_SW_b[3].n5 VSS_SW_b[3].n4 7.57742
R12506 VSS_SW_b[3].n2 VSS_SW_b[3] 5.61454
R12507 VSS_SW_b[3].n8 VSS_SW_b[3].n6 2.47092
R12508 VSS_SW_b[3].n3 VSS_SW_b[3] 2.02155
R12509 VSS_SW_b[3].n12 VSS_SW_b[3] 1.6999
R12510 VSS_SW_b[3].n6 VSS_SW_b[3].n0 1.50964
R12511 VSS_SW_b[3].n10 VSS_SW_b[3].n9 1.5083
R12512 VSS_SW_b[3] VSS_SW_b[3].n12 1.3731
R12513 VSS_SW_b[3] VSS_SW_b[3].n1 1.34787
R12514 VSS_SW_b[3].n1 VSS_SW_b[3].n0 0.449623
R12515 VSS_SW_b[3].n12 VSS_SW_b[3].n11 0.0501381
R12516 VSS_SW_b[3].n11 VSS_SW_b[3].n10 0.0260996
R12517 VSS_SW_b[3].n8 VSS_SW_b[3].n7 0.0219844
R12518 VSS_SW_b[3].n9 VSS_SW_b[3].n8 0.00489987
R12519 D[6].n0 D[6].t2 331.51
R12520 D[6].n5 D[6].t3 331.51
R12521 D[6].n0 D[6].t1 209.403
R12522 D[6].n5 D[6].t0 209.403
R12523 D[6].n1 D[6].n0 76.0005
R12524 D[6].n6 D[6].n5 76.0005
R12525 D[6].n3 D[6].n2 14.0187
R12526 D[6].n2 D[6].n1 8.11757
R12527 D[6].n4 D[6] 7.49318
R12528 D[6].n4 D[6].n3 6.97656
R12529 D[6].n1 D[6] 2.02977
R12530 D[6] D[6].n6 2.02977
R12531 D[6].n6 D[6].n4 1.09318
R12532 D[6].n2 D[6] 0.468793
R12533 D[6].n3 D[6] 0.0519212
R12534 check[1] check[1].n3 363.457
R12535 check[1] check[1].n1 352.005
R12536 check[1].n0 check[1].t3 329.762
R12537 check[1].n7 check[1].t1 328.118
R12538 check[1].n3 check[1].t4 272.062
R12539 check[1].n1 check[1].t6 272.062
R12540 check[1].n3 check[1].t5 206.19
R12541 check[1].n1 check[1].t7 206.19
R12542 check[1].n0 check[1].t2 147.188
R12543 check[1].n6 check[1].t0 141.374
R12544 check[1].n16 check[1] 28.0657
R12545 check[1].n4 check[1] 15.1584
R12546 check[1].n8 check[1].n7 9.3005
R12547 check[1].n7 check[1].n6 8.19823
R12548 check[1] check[1].n0 7.17927
R12549 check[1].n5 check[1].n4 5.05313
R12550 check[1].n10 check[1].n9 5.05313
R12551 check[1].n16 check[1].n15 4.77557
R12552 check[1].n9 check[1] 4.37945
R12553 check[1].n13 check[1].n10 3.03311
R12554 check[1] check[1].n16 1.31653
R12555 check[1].n8 check[1].n5 0.674184
R12556 check[1].n10 check[1].n8 0.674184
R12557 check[1].n13 check[1].n12 0.166613
R12558 check[1].n12 check[1] 0.0531797
R12559 check[1].n14 check[1].n13 0.0352222
R12560 check[1].n15 check[1].n14 0.0167037
R12561 check[1].n12 check[1].n11 0.00485575
R12562 check[1].n13 check[1].n2 0.00331272
R12563 D[2].n0 D[2].t3 331.51
R12564 D[2].n5 D[2].t0 331.51
R12565 D[2].n0 D[2].t2 209.403
R12566 D[2].n5 D[2].t1 209.403
R12567 D[2].n1 D[2].n0 76.0005
R12568 D[2].n6 D[2].n5 76.0005
R12569 D[2].n3 D[2].n2 14.0187
R12570 D[2].n2 D[2].n1 8.27367
R12571 D[2].n4 D[2] 7.49318
R12572 D[2].n4 D[2].n3 6.97953
R12573 D[2].n1 D[2] 2.02977
R12574 D[2] D[2].n6 2.02977
R12575 D[2].n6 D[2].n4 1.09318
R12576 D[2].n2 D[2] 0.312695
R12577 D[2].n3 D[2] 0.051922
R12578 VDD_SW_b[6].n3 VDD_SW_b[6].t1 117.424
R12579 VDD_SW_b[6].n0 VDD_SW_b[6].t0 100.715
R12580 VDD_SW_b[6].n4 VDD_SW_b[6].n3 76.5198
R12581 VDD_SW_b[6].n0 VDD_SW_b[6] 10.2646
R12582 VDD_SW_b[6].n6 VDD_SW_b[6].n4 9.3005
R12583 VDD_SW_b[6].n3 VDD_SW_b[6] 5.61454
R12584 VDD_SW_b[6].n6 VDD_SW_b[6].n2 4.5005
R12585 VDD_SW_b[6].n1 VDD_SW_b[6].n0 3.75113
R12586 VDD_SW_b[6].n10 VDD_SW_b[6] 3.66121
R12587 VDD_SW_b[6] VDD_SW_b[6].n10 2.95723
R12588 VDD_SW_b[6].n4 VDD_SW_b[6] 2.9198
R12589 VDD_SW_b[6].n8 VDD_SW_b[6].n7 1.50505
R12590 VDD_SW_b[6].n2 VDD_SW_b[6].n1 0.449623
R12591 VDD_SW_b[6] VDD_SW_b[6].n2 0.449623
R12592 VDD_SW_b[6].n10 VDD_SW_b[6].n9 0.0501381
R12593 VDD_SW_b[6].n9 VDD_SW_b[6].n8 0.0260996
R12594 VDD_SW_b[6].n6 VDD_SW_b[6].n5 0.0122188
R12595 VDD_SW_b[6].n7 VDD_SW_b[6].n6 0.00814977
R12596 D[3].n0 D[3].t0 331.51
R12597 D[3].n5 D[3].t1 331.51
R12598 D[3].n0 D[3].t3 209.403
R12599 D[3].n5 D[3].t2 209.403
R12600 D[3].n1 D[3].n0 76.0005
R12601 D[3].n6 D[3].n5 76.0005
R12602 D[3].n3 D[3].n2 14.0217
R12603 D[3].n2 D[3].n1 8.11757
R12604 D[3].n4 D[3] 7.49318
R12605 D[3].n4 D[3].n3 6.97953
R12606 D[3].n1 D[3] 2.02977
R12607 D[3] D[3].n6 2.02977
R12608 D[3].n6 D[3].n4 1.09318
R12609 D[3].n2 D[3] 0.468793
R12610 D[3].n3 D[3] 0.051922
R12611 VSS_SW_b[2].n4 VSS_SW_b[2].n3 638.038
R12612 VSS_SW_b[2] VSS_SW_b[2].t0 422.656
R12613 VSS_SW_b[2].t0 VSS_SW_b[2].n5 117.442
R12614 VSS_SW_b[2].n2 VSS_SW_b[2].t1 117.424
R12615 VSS_SW_b[2].n3 VSS_SW_b[2].n2 77.6426
R12616 VSS_SW_b[2].n5 VSS_SW_b[2].n4 11.3659
R12617 VSS_SW_b[2].n6 VSS_SW_b[2] 11.1582
R12618 VSS_SW_b[2].n5 VSS_SW_b[2].n0 9.15497
R12619 VSS_SW_b[2].n2 VSS_SW_b[2] 5.61454
R12620 VSS_SW_b[2].n8 VSS_SW_b[2].n6 2.47092
R12621 VSS_SW_b[2].n3 VSS_SW_b[2] 1.79699
R12622 VSS_SW_b[2].n12 VSS_SW_b[2] 1.70288
R12623 VSS_SW_b[2].n6 VSS_SW_b[2].n0 1.50964
R12624 VSS_SW_b[2].n10 VSS_SW_b[2].n9 1.5083
R12625 VSS_SW_b[2] VSS_SW_b[2].n12 1.3755
R12626 VSS_SW_b[2] VSS_SW_b[2].n1 1.34787
R12627 VSS_SW_b[2].n1 VSS_SW_b[2].n0 0.674184
R12628 VSS_SW_b[2].n12 VSS_SW_b[2].n11 0.0501381
R12629 VSS_SW_b[2].n11 VSS_SW_b[2].n10 0.0260996
R12630 VSS_SW_b[2].n8 VSS_SW_b[2].n7 0.0219844
R12631 VSS_SW_b[2].n9 VSS_SW_b[2].n8 0.00489987
R12632 check[4] check[4].n3 363.457
R12633 check[4] check[4].n1 352.005
R12634 check[4].n0 check[4].t7 328.911
R12635 check[4].n7 check[4].t5 328.118
R12636 check[4].n3 check[4].t0 272.062
R12637 check[4].n1 check[4].t2 272.062
R12638 check[4].n3 check[4].t1 206.19
R12639 check[4].n1 check[4].t3 206.19
R12640 check[4].n0 check[4].t6 148.035
R12641 check[4].n6 check[4].t4 141.374
R12642 check[4].n16 check[4] 28.0656
R12643 check[4].n4 check[4] 15.1584
R12644 check[4].n8 check[4].n7 9.3005
R12645 check[4].n7 check[4].n6 8.19823
R12646 check[4] check[4].n0 7.14463
R12647 check[4].n10 check[4].n9 5.38997
R12648 check[4].n16 check[4].n15 5.06786
R12649 check[4].n5 check[4].n4 5.05313
R12650 check[4].n9 check[4] 4.37945
R12651 check[4].n13 check[4].n10 3.03311
R12652 check[4] check[4].n16 1.31656
R12653 check[4].n8 check[4].n5 0.674184
R12654 check[4].n10 check[4].n8 0.337342
R12655 check[4].n13 check[4].n12 0.166613
R12656 check[4].n12 check[4] 0.0531797
R12657 check[4].n14 check[4].n13 0.037537
R12658 check[4].n15 check[4].n14 0.0143889
R12659 check[4].n12 check[4].n11 0.00485575
R12660 check[4].n13 check[4].n2 0.00215636
R12661 VDD_SW[4].n8 VDD_SW[4].t1 117.424
R12662 VDD_SW[4].n6 VDD_SW[4].t0 75.7697
R12663 VDD_SW[4].n7 VDD_SW[4].n6 73.0808
R12664 VDD_SW[4] VDD_SW[4].n8 67.6928
R12665 VDD_SW[4].n10 VDD_SW[4].n9 13.0467
R12666 VDD_SW[4].n8 VDD_SW[4] 6.64665
R12667 VDD_SW[4].n5 VDD_SW[4].n4 2.82795
R12668 VDD_SW[4] VDD_SW[4].n7 2.2023
R12669 VDD_SW[4] VDD_SW[4].n10 1.96973
R12670 VDD_SW[4].n9 VDD_SW[4] 1.72358
R12671 VDD_SW[4].n3 VDD_SW[4].n1 1.49691
R12672 VDD_SW[4].n1 VDD_SW[4] 0.0595299
R12673 VDD_SW[4].n1 VDD_SW[4].n0 0.0177811
R12674 VDD_SW[4].n7 VDD_SW[4].n5 0.0146776
R12675 VDD_SW[4].n3 VDD_SW[4].n2 0.0102656
R12676 VDD_SW[4].n4 VDD_SW[4].n3 0.00635152
R12677 D[7].n0 D[7].t1 331.51
R12678 D[7].n5 D[7].t3 331.51
R12679 D[7].n0 D[7].t2 209.403
R12680 D[7].n5 D[7].t0 209.403
R12681 D[7].n1 D[7].n0 76.0005
R12682 D[7].n6 D[7].n5 76.0005
R12683 D[7].n3 D[7].n2 14.0187
R12684 D[7].n2 D[7].n1 8.11757
R12685 D[7].n4 D[7] 7.49318
R12686 D[7].n4 D[7].n3 6.97656
R12687 D[7].n1 D[7] 2.02977
R12688 D[7] D[7].n6 2.02977
R12689 D[7].n6 D[7].n4 1.09318
R12690 D[7].n2 D[7] 0.468793
R12691 D[7].n3 D[7] 0.0519212
R12692 check[3] check[3].n3 363.457
R12693 check[3] check[3].n1 352.005
R12694 check[3].n7 check[3].t1 329.01
R12695 check[3].n0 check[3].t5 328.911
R12696 check[3].n3 check[3].t6 272.062
R12697 check[3].n1 check[3].t2 272.062
R12698 check[3].n3 check[3].t7 206.19
R12699 check[3].n1 check[3].t3 206.19
R12700 check[3].n0 check[3].t4 148.035
R12701 check[3].n6 check[3].t0 140.888
R12702 check[3].n16 check[3] 28.1395
R12703 check[3].n4 check[3] 15.1584
R12704 check[3].n8 check[3].n7 9.3005
R12705 check[3].n7 check[3].n6 7.71392
R12706 check[3] check[3].n0 7.14463
R12707 check[3].n10 check[3].n9 5.38997
R12708 check[3].n5 check[3].n4 5.05313
R12709 check[3].n16 check[3].n15 4.87033
R12710 check[3].n9 check[3] 4.37945
R12711 check[3].n13 check[3].n10 3.03311
R12712 check[3] check[3].n16 1.15253
R12713 check[3].n8 check[3].n5 0.674184
R12714 check[3].n10 check[3].n8 0.337342
R12715 check[3].n13 check[3].n12 0.166613
R12716 check[3].n12 check[3] 0.0531806
R12717 check[3].n14 check[3].n13 0.037537
R12718 check[3].n15 check[3].n14 0.0143889
R12719 check[3].n12 check[3].n11 0.00485575
R12720 check[3].n13 check[3].n2 0.00215636
R12721 check[0] check[0].n3 363.457
R12722 check[0] check[0].n1 352.005
R12723 check[0].n0 check[0].t3 329.762
R12724 check[0].n7 check[0].t5 329.01
R12725 check[0].n3 check[0].t0 272.062
R12726 check[0].n1 check[0].t6 272.062
R12727 check[0].n3 check[0].t1 206.19
R12728 check[0].n1 check[0].t7 206.19
R12729 check[0].n0 check[0].t2 147.188
R12730 check[0].n6 check[0].t4 140.888
R12731 check[0].n16 check[0] 28.1411
R12732 check[0].n4 check[0] 15.1584
R12733 check[0].n8 check[0].n7 9.3005
R12734 check[0].n7 check[0].n6 7.71392
R12735 check[0] check[0].n0 7.17927
R12736 check[0].n10 check[0].n9 5.38997
R12737 check[0].n5 check[0].n4 5.05313
R12738 check[0].n16 check[0].n15 4.81189
R12739 check[0].n9 check[0] 4.37945
R12740 check[0].n13 check[0].n10 3.03311
R12741 check[0] check[0].n16 1.15191
R12742 check[0].n8 check[0].n5 0.674184
R12743 check[0].n10 check[0].n8 0.337342
R12744 check[0].n13 check[0].n12 0.166613
R12745 check[0].n12 check[0] 0.0531806
R12746 check[0].n14 check[0].n13 0.037537
R12747 check[0].n15 check[0].n14 0.0143889
R12748 check[0].n12 check[0].n11 0.00485575
R12749 check[0].n13 check[0].n2 0.00215636
R12750 reset.n2 reset.t0 255.25
R12751 reset.n0 reset.t1 169.462
R12752 reset.n3 reset.n2 9.3005
R12753 reset.n1 reset.n0 5.70839
R12754 reset.n3 reset 5.61776
R12755 reset.n2 reset.n1 5.07418
R12756 reset.n5 reset.n4 1.69462
R12757 reset.n4 reset.n3 1.50638
R12758 reset reset.n5 0.376971
R12759 D[4].n0 D[4].t0 331.51
R12760 D[4].n5 D[4].t1 331.51
R12761 D[4].n0 D[4].t3 209.403
R12762 D[4].n5 D[4].t2 209.403
R12763 D[4].n1 D[4].n0 76.0005
R12764 D[4].n6 D[4].n5 76.0005
R12765 D[4].n3 D[4].n2 14.0157
R12766 D[4].n2 D[4].n1 8.27367
R12767 D[4].n4 D[4] 7.49318
R12768 D[4].n4 D[4].n3 6.97656
R12769 D[4].n1 D[4] 2.02977
R12770 D[4] D[4].n6 2.02977
R12771 D[4].n6 D[4].n4 1.09318
R12772 D[4].n2 D[4] 0.312695
R12773 D[4].n3 D[4] 0.0519212
R12774 VSS_SW_b[4].n4 VSS_SW_b[4].n3 641.827
R12775 VSS_SW_b[4] VSS_SW_b[4].t0 422.656
R12776 VSS_SW_b[4].t0 VSS_SW_b[4].n5 121.231
R12777 VSS_SW_b[4].n2 VSS_SW_b[4].t1 117.424
R12778 VSS_SW_b[4].n3 VSS_SW_b[4].n2 77.418
R12779 VSS_SW_b[4].n6 VSS_SW_b[4] 11.3827
R12780 VSS_SW_b[4].n5 VSS_SW_b[4].n0 9.15497
R12781 VSS_SW_b[4].n5 VSS_SW_b[4].n4 7.57742
R12782 VSS_SW_b[4].n2 VSS_SW_b[4] 5.61454
R12783 VSS_SW_b[4].n8 VSS_SW_b[4].n6 2.47092
R12784 VSS_SW_b[4].n3 VSS_SW_b[4] 2.02155
R12785 VSS_SW_b[4].n12 VSS_SW_b[4] 1.6999
R12786 VSS_SW_b[4].n6 VSS_SW_b[4].n0 1.50964
R12787 VSS_SW_b[4].n10 VSS_SW_b[4].n9 1.5083
R12788 VSS_SW_b[4] VSS_SW_b[4].n12 1.3731
R12789 VSS_SW_b[4] VSS_SW_b[4].n1 1.34787
R12790 VSS_SW_b[4].n1 VSS_SW_b[4].n0 0.449623
R12791 VSS_SW_b[4].n12 VSS_SW_b[4].n11 0.0501381
R12792 VSS_SW_b[4].n11 VSS_SW_b[4].n10 0.0260996
R12793 VSS_SW_b[4].n8 VSS_SW_b[4].n7 0.0219844
R12794 VSS_SW_b[4].n9 VSS_SW_b[4].n8 0.00489987
R12795 VDD_SW_b[1].n3 VDD_SW_b[1].t1 117.424
R12796 VDD_SW_b[1].n0 VDD_SW_b[1].t0 100.715
R12797 VDD_SW_b[1].n4 VDD_SW_b[1].n3 76.5198
R12798 VDD_SW_b[1].n0 VDD_SW_b[1] 10.2646
R12799 VDD_SW_b[1].n6 VDD_SW_b[1].n4 9.3005
R12800 VDD_SW_b[1].n3 VDD_SW_b[1] 5.61454
R12801 VDD_SW_b[1].n6 VDD_SW_b[1].n2 4.5005
R12802 VDD_SW_b[1].n1 VDD_SW_b[1].n0 3.75113
R12803 VDD_SW_b[1].n10 VDD_SW_b[1] 3.66419
R12804 VDD_SW_b[1] VDD_SW_b[1].n10 2.95963
R12805 VDD_SW_b[1].n4 VDD_SW_b[1] 2.9198
R12806 VDD_SW_b[1].n8 VDD_SW_b[1].n7 1.50505
R12807 VDD_SW_b[1] VDD_SW_b[1].n2 0.674184
R12808 VDD_SW_b[1].n2 VDD_SW_b[1].n1 0.225061
R12809 VDD_SW_b[1].n10 VDD_SW_b[1].n9 0.0501381
R12810 VDD_SW_b[1].n9 VDD_SW_b[1].n8 0.0260996
R12811 VDD_SW_b[1].n6 VDD_SW_b[1].n5 0.0122188
R12812 VDD_SW_b[1].n7 VDD_SW_b[1].n6 0.00814977
R12813 check[2] check[2].n3 363.457
R12814 check[2] check[2].n1 352.005
R12815 check[2].n0 check[2].t5 329.762
R12816 check[2].n7 check[2].t7 328.118
R12817 check[2].n3 check[2].t2 272.062
R12818 check[2].n1 check[2].t0 272.062
R12819 check[2].n3 check[2].t3 206.19
R12820 check[2].n1 check[2].t1 206.19
R12821 check[2].n0 check[2].t4 147.188
R12822 check[2].n6 check[2].t6 141.374
R12823 check[2].n16 check[2] 28.0653
R12824 check[2].n4 check[2] 15.1584
R12825 check[2].n8 check[2].n7 9.3005
R12826 check[2].n7 check[2].n6 8.19823
R12827 check[2] check[2].n0 7.17927
R12828 check[2].n10 check[2].n9 5.38997
R12829 check[2].n5 check[2].n4 5.05313
R12830 check[2].n16 check[2].n15 4.97041
R12831 check[2].n9 check[2] 4.37945
R12832 check[2].n13 check[2].n10 3.03311
R12833 check[2] check[2].n16 1.31669
R12834 check[2].n8 check[2].n5 0.674184
R12835 check[2].n10 check[2].n8 0.337342
R12836 check[2].n13 check[2].n12 0.166613
R12837 check[2].n12 check[2] 0.0531797
R12838 check[2].n14 check[2].n13 0.037537
R12839 check[2].n15 check[2].n14 0.0143889
R12840 check[2].n12 check[2].n11 0.00485575
R12841 check[2].n13 check[2].n2 0.00215636
R12842 VDD_SW[5].n8 VDD_SW[5].t1 117.424
R12843 VDD_SW[5].n6 VDD_SW[5].t0 75.7697
R12844 VDD_SW[5].n7 VDD_SW[5].n6 73.0808
R12845 VDD_SW[5] VDD_SW[5].n8 67.6928
R12846 VDD_SW[5].n10 VDD_SW[5].n9 13.0467
R12847 VDD_SW[5].n8 VDD_SW[5] 6.64665
R12848 VDD_SW[5].n5 VDD_SW[5].n4 2.82795
R12849 VDD_SW[5] VDD_SW[5].n7 2.2023
R12850 VDD_SW[5] VDD_SW[5].n10 1.96973
R12851 VDD_SW[5].n9 VDD_SW[5] 1.72358
R12852 VDD_SW[5].n3 VDD_SW[5].n1 1.49691
R12853 VDD_SW[5].n1 VDD_SW[5] 0.0595299
R12854 VDD_SW[5].n1 VDD_SW[5].n0 0.0177811
R12855 VDD_SW[5].n7 VDD_SW[5].n5 0.0146776
R12856 VDD_SW[5].n3 VDD_SW[5].n2 0.0102656
R12857 VDD_SW[5].n4 VDD_SW[5].n3 0.00635152
R12858 D[1].n0 D[1].t1 331.51
R12859 D[1].n5 D[1].t2 331.51
R12860 D[1].n0 D[1].t0 209.403
R12861 D[1].n5 D[1].t3 209.403
R12862 D[1].n1 D[1].n0 76.0005
R12863 D[1].n6 D[1].n5 76.0005
R12864 D[1].n3 D[1].n2 14.0217
R12865 D[1].n2 D[1].n1 8.11757
R12866 D[1].n4 D[1] 7.49318
R12867 D[1].n4 D[1].n3 6.97953
R12868 D[1].n1 D[1] 2.02977
R12869 D[1] D[1].n6 2.02977
R12870 D[1].n6 D[1].n4 1.09318
R12871 D[1].n2 D[1] 0.468793
R12872 D[1].n3 D[1] 0.051922
R12873 D[5].n0 D[5].t0 331.51
R12874 D[5].n5 D[5].t1 331.51
R12875 D[5].n0 D[5].t3 209.403
R12876 D[5].n5 D[5].t2 209.403
R12877 D[5].n1 D[5].n0 76.0005
R12878 D[5].n6 D[5].n5 76.0005
R12879 D[5].n3 D[5].n2 14.0187
R12880 D[5].n2 D[5].n1 8.27367
R12881 D[5].n4 D[5].n3 7.5711
R12882 D[5].n4 D[5] 7.33709
R12883 D[5].n1 D[5] 2.02977
R12884 D[5] D[5].n6 2.02977
R12885 D[5].n6 D[5].n4 1.24928
R12886 D[5].n2 D[5] 0.312695
R12887 D[5].n3 D[5] 0.051922
R12888 VDD_SW[6].n8 VDD_SW[6].t1 117.424
R12889 VDD_SW[6].n6 VDD_SW[6].t0 75.7697
R12890 VDD_SW[6].n7 VDD_SW[6].n6 73.0808
R12891 VDD_SW[6] VDD_SW[6].n8 67.6928
R12892 VDD_SW[6].n10 VDD_SW[6].n9 13.0467
R12893 VDD_SW[6].n8 VDD_SW[6] 6.64665
R12894 VDD_SW[6].n5 VDD_SW[6].n4 2.82795
R12895 VDD_SW[6] VDD_SW[6].n7 2.2023
R12896 VDD_SW[6] VDD_SW[6].n10 1.96973
R12897 VDD_SW[6].n9 VDD_SW[6] 1.72358
R12898 VDD_SW[6].n3 VDD_SW[6].n1 1.49691
R12899 VDD_SW[6].n1 VDD_SW[6] 0.0595299
R12900 VDD_SW[6].n1 VDD_SW[6].n0 0.0177811
R12901 VDD_SW[6].n7 VDD_SW[6].n5 0.0146776
R12902 VDD_SW[6].n3 VDD_SW[6].n2 0.0102656
R12903 VDD_SW[6].n4 VDD_SW[6].n3 0.00635152
R12904 VSS_SW_b[5].n4 VSS_SW_b[5].n3 641.827
R12905 VSS_SW_b[5] VSS_SW_b[5].t0 422.656
R12906 VSS_SW_b[5].t0 VSS_SW_b[5].n5 121.231
R12907 VSS_SW_b[5].n2 VSS_SW_b[5].t1 117.424
R12908 VSS_SW_b[5].n3 VSS_SW_b[5].n2 77.418
R12909 VSS_SW_b[5].n6 VSS_SW_b[5] 11.3827
R12910 VSS_SW_b[5].n5 VSS_SW_b[5].n0 9.15497
R12911 VSS_SW_b[5].n5 VSS_SW_b[5].n4 7.57742
R12912 VSS_SW_b[5].n2 VSS_SW_b[5] 5.61454
R12913 VSS_SW_b[5].n8 VSS_SW_b[5].n6 2.47092
R12914 VSS_SW_b[5].n3 VSS_SW_b[5] 2.02155
R12915 VSS_SW_b[5].n12 VSS_SW_b[5] 1.6999
R12916 VSS_SW_b[5].n6 VSS_SW_b[5].n0 1.50964
R12917 VSS_SW_b[5].n10 VSS_SW_b[5].n9 1.5083
R12918 VSS_SW_b[5] VSS_SW_b[5].n12 1.3731
R12919 VSS_SW_b[5] VSS_SW_b[5].n1 1.34787
R12920 VSS_SW_b[5].n1 VSS_SW_b[5].n0 0.449623
R12921 VSS_SW_b[5].n12 VSS_SW_b[5].n11 0.0501381
R12922 VSS_SW_b[5].n11 VSS_SW_b[5].n10 0.0260996
R12923 VSS_SW_b[5].n8 VSS_SW_b[5].n7 0.0219844
R12924 VSS_SW_b[5].n9 VSS_SW_b[5].n8 0.00489987
R12925 VSS_SW_b[7].n4 VSS_SW_b[7].n3 641.827
R12926 VSS_SW_b[7] VSS_SW_b[7].t0 422.656
R12927 VSS_SW_b[7].t0 VSS_SW_b[7].n5 121.231
R12928 VSS_SW_b[7].n2 VSS_SW_b[7].t1 117.424
R12929 VSS_SW_b[7].n3 VSS_SW_b[7].n2 77.418
R12930 VSS_SW_b[7].n6 VSS_SW_b[7] 11.3827
R12931 VSS_SW_b[7].n5 VSS_SW_b[7].n0 9.15497
R12932 VSS_SW_b[7].n5 VSS_SW_b[7].n4 7.57742
R12933 VSS_SW_b[7].n2 VSS_SW_b[7] 5.61454
R12934 VSS_SW_b[7].n8 VSS_SW_b[7].n6 2.47092
R12935 VSS_SW_b[7].n3 VSS_SW_b[7] 2.02155
R12936 VSS_SW_b[7].n12 VSS_SW_b[7] 1.6999
R12937 VSS_SW_b[7].n6 VSS_SW_b[7].n0 1.50964
R12938 VSS_SW_b[7].n10 VSS_SW_b[7].n9 1.5083
R12939 VSS_SW_b[7] VSS_SW_b[7].n12 1.3731
R12940 VSS_SW_b[7] VSS_SW_b[7].n1 1.34787
R12941 VSS_SW_b[7].n1 VSS_SW_b[7].n0 0.449623
R12942 VSS_SW_b[7].n12 VSS_SW_b[7].n11 0.0501381
R12943 VSS_SW_b[7].n11 VSS_SW_b[7].n10 0.0260996
R12944 VSS_SW_b[7].n8 VSS_SW_b[7].n7 0.0219844
R12945 VSS_SW_b[7].n9 VSS_SW_b[7].n8 0.00489987
R12946 VDD_SW[7].n8 VDD_SW[7].t1 117.424
R12947 VDD_SW[7].n6 VDD_SW[7].t0 75.7697
R12948 VDD_SW[7].n7 VDD_SW[7].n6 73.0808
R12949 VDD_SW[7] VDD_SW[7].n8 67.6928
R12950 VDD_SW[7].n10 VDD_SW[7].n9 13.0467
R12951 VDD_SW[7].n8 VDD_SW[7] 6.64665
R12952 VDD_SW[7].n5 VDD_SW[7].n4 2.82795
R12953 VDD_SW[7] VDD_SW[7].n7 2.2023
R12954 VDD_SW[7] VDD_SW[7].n10 1.96973
R12955 VDD_SW[7].n9 VDD_SW[7] 1.72358
R12956 VDD_SW[7].n3 VDD_SW[7].n1 1.49691
R12957 VDD_SW[7].n1 VDD_SW[7] 0.0595299
R12958 VDD_SW[7].n1 VDD_SW[7].n0 0.0177811
R12959 VDD_SW[7].n7 VDD_SW[7].n5 0.0146776
R12960 VDD_SW[7].n3 VDD_SW[7].n2 0.0102656
R12961 VDD_SW[7].n4 VDD_SW[7].n3 0.00635152
R12962 VDD_SW_b[5].n3 VDD_SW_b[5].t1 117.424
R12963 VDD_SW_b[5].n0 VDD_SW_b[5].t0 100.715
R12964 VDD_SW_b[5].n4 VDD_SW_b[5].n3 76.5198
R12965 VDD_SW_b[5].n0 VDD_SW_b[5] 10.2646
R12966 VDD_SW_b[5].n6 VDD_SW_b[5].n4 9.3005
R12967 VDD_SW_b[5].n3 VDD_SW_b[5] 5.61454
R12968 VDD_SW_b[5].n6 VDD_SW_b[5].n2 4.5005
R12969 VDD_SW_b[5].n1 VDD_SW_b[5].n0 3.75113
R12970 VDD_SW_b[5].n10 VDD_SW_b[5] 3.66121
R12971 VDD_SW_b[5] VDD_SW_b[5].n10 2.95723
R12972 VDD_SW_b[5].n4 VDD_SW_b[5] 2.9198
R12973 VDD_SW_b[5].n8 VDD_SW_b[5].n7 1.5044
R12974 VDD_SW_b[5].n2 VDD_SW_b[5].n1 0.449623
R12975 VDD_SW_b[5] VDD_SW_b[5].n2 0.449623
R12976 VDD_SW_b[5].n10 VDD_SW_b[5].n9 0.0501381
R12977 VDD_SW_b[5].n9 VDD_SW_b[5].n8 0.0260996
R12978 VDD_SW_b[5].n6 VDD_SW_b[5].n5 0.0102656
R12979 VDD_SW_b[5].n7 VDD_SW_b[5].n6 0.00879975
R12980 VDD_SW[1].n8 VDD_SW[1].t1 117.424
R12981 VDD_SW[1].n6 VDD_SW[1].t0 75.7697
R12982 VDD_SW[1].n7 VDD_SW[1].n6 73.0808
R12983 VDD_SW[1] VDD_SW[1].n8 67.6928
R12984 VDD_SW[1].n10 VDD_SW[1].n9 13.0467
R12985 VDD_SW[1].n8 VDD_SW[1] 6.64665
R12986 VDD_SW[1].n5 VDD_SW[1].n4 2.82795
R12987 VDD_SW[1] VDD_SW[1].n7 2.2023
R12988 VDD_SW[1] VDD_SW[1].n10 1.96973
R12989 VDD_SW[1].n9 VDD_SW[1] 1.72358
R12990 VDD_SW[1].n3 VDD_SW[1].n1 1.49691
R12991 VDD_SW[1].n1 VDD_SW[1] 0.0595299
R12992 VDD_SW[1].n1 VDD_SW[1].n0 0.0177811
R12993 VDD_SW[1].n7 VDD_SW[1].n5 0.0146776
R12994 VDD_SW[1].n3 VDD_SW[1].n2 0.0102656
R12995 VDD_SW[1].n4 VDD_SW[1].n3 0.00635152
R12996 VSS_SW[3].n3 VSS_SW[3].n2 585
R12997 VSS_SW[3].n1 VSS_SW[3].t0 417.519
R12998 VSS_SW[3].n0 VSS_SW[3].t1 117.424
R12999 VSS_SW[3].n4 VSS_SW[3].n3 73.4178
R13000 VSS_SW[3].n3 VSS_SW[3].t0 68.1928
R13001 VSS_SW[3] VSS_SW[3].n0 67.6928
R13002 VSS_SW[3].n2 VSS_SW[3].n1 12.5543
R13003 VSS_SW[3].n0 VSS_SW[3] 6.64665
R13004 VSS_SW[3] VSS_SW[3].n4 3.039
R13005 VSS_SW[3].n2 VSS_SW[3] 2.46204
R13006 VSS_SW[3].n4 VSS_SW[3] 1.72358
R13007 VSS_SW[3].n1 VSS_SW[3] 1.72358
R13008 VSS_SW[5].n3 VSS_SW[5].n0 585
R13009 VSS_SW[5].n2 VSS_SW[5].t0 417.519
R13010 VSS_SW[5].n1 VSS_SW[5].t1 117.424
R13011 VSS_SW[5].n4 VSS_SW[5].n0 73.2739
R13012 VSS_SW[5].t0 VSS_SW[5].n0 71.9813
R13013 VSS_SW[5] VSS_SW[5].n1 67.6928
R13014 VSS_SW[5].n3 VSS_SW[5].n2 12.8005
R13015 VSS_SW[5].n1 VSS_SW[5] 6.64665
R13016 VSS_SW[5] VSS_SW[5].n4 3.04482
R13017 VSS_SW[5] VSS_SW[5].n3 2.21588
R13018 VSS_SW[5].n4 VSS_SW[5] 1.9648
R13019 VSS_SW[5].n2 VSS_SW[5] 1.72358
R13020 check[6] check[6].n3 363.457
R13021 check[6] check[6].n1 352.005
R13022 check[6].n7 check[6].t5 329.01
R13023 check[6].n0 check[6].t7 328.911
R13024 check[6].n3 check[6].t0 272.062
R13025 check[6].n1 check[6].t2 272.062
R13026 check[6].n3 check[6].t1 206.19
R13027 check[6].n1 check[6].t3 206.19
R13028 check[6].n0 check[6].t6 148.035
R13029 check[6].n6 check[6].t4 140.888
R13030 check[6].n16 check[6] 28.1391
R13031 check[6].n4 check[6] 15.1584
R13032 check[6].n8 check[6].n7 9.3005
R13033 check[6].n7 check[6].n6 7.71392
R13034 check[6] check[6].n0 7.14463
R13035 check[6].n10 check[6].n9 5.38997
R13036 check[6].n5 check[6].n4 5.05313
R13037 check[6].n16 check[6].n15 4.76728
R13038 check[6].n9 check[6] 4.37945
R13039 check[6].n13 check[6].n10 3.03311
R13040 check[6] check[6].n16 1.15267
R13041 check[6].n8 check[6].n5 0.674184
R13042 check[6].n10 check[6].n8 0.337342
R13043 check[6].n13 check[6].n12 0.166672
R13044 check[6].n12 check[6] 0.0532291
R13045 check[6].n14 check[6].n13 0.037537
R13046 check[6].n15 check[6].n14 0.0143889
R13047 check[6].n12 check[6].n11 0.00481511
R13048 check[6].n13 check[6].n2 0.00215119
R13049 ready.n0 ready.t0 259.723
R13050 ready.n0 ready.t1 175.108
R13051 ready.n1 ready 19.9175
R13052 ready.n1 ready.n0 8.27037
R13053 ready ready.n1 1.16637
R13054 VDD_SW[2].n8 VDD_SW[2].t1 117.424
R13055 VDD_SW[2].n6 VDD_SW[2].t0 75.7697
R13056 VDD_SW[2].n7 VDD_SW[2].n6 73.0808
R13057 VDD_SW[2] VDD_SW[2].n8 67.6928
R13058 VDD_SW[2].n10 VDD_SW[2].n9 13.0467
R13059 VDD_SW[2].n8 VDD_SW[2] 6.64665
R13060 VDD_SW[2].n5 VDD_SW[2].n4 2.82795
R13061 VDD_SW[2] VDD_SW[2].n7 2.2023
R13062 VDD_SW[2] VDD_SW[2].n10 1.96973
R13063 VDD_SW[2].n9 VDD_SW[2] 1.72358
R13064 VDD_SW[2].n3 VDD_SW[2].n1 1.49691
R13065 VDD_SW[2].n1 VDD_SW[2] 0.0595299
R13066 VDD_SW[2].n1 VDD_SW[2].n0 0.0177811
R13067 VDD_SW[2].n7 VDD_SW[2].n5 0.0146776
R13068 VDD_SW[2].n3 VDD_SW[2].n2 0.0102656
R13069 VDD_SW[2].n4 VDD_SW[2].n3 0.00635152
R13070 check[5] check[5].n3 363.457
R13071 check[5] check[5].n1 352.005
R13072 check[5].n0 check[5].t1 328.911
R13073 check[5].n7 check[5].t3 328.118
R13074 check[5].n3 check[5].t6 272.062
R13075 check[5].n1 check[5].t4 272.062
R13076 check[5].n3 check[5].t7 206.19
R13077 check[5].n1 check[5].t5 206.19
R13078 check[5].n0 check[5].t0 148.035
R13079 check[5].n6 check[5].t2 141.374
R13080 check[5].n16 check[5] 28.1388
R13081 check[5].n4 check[5] 15.1584
R13082 check[5].n8 check[5].n7 9.3005
R13083 check[5].n7 check[5].n6 8.19823
R13084 check[5] check[5].n0 7.14463
R13085 check[5].n10 check[5].n9 5.38997
R13086 check[5].n5 check[5].n4 5.05313
R13087 check[5].n16 check[5].n15 4.76129
R13088 check[5].n9 check[5] 4.37945
R13089 check[5].n13 check[5].n10 3.03311
R13090 check[5] check[5].n16 1.15277
R13091 check[5].n8 check[5].n5 0.674184
R13092 check[5].n10 check[5].n8 0.337342
R13093 check[5].n13 check[5].n12 0.166672
R13094 check[5].n12 check[5] 0.0532282
R13095 check[5].n14 check[5].n13 0.037537
R13096 check[5].n15 check[5].n14 0.0143889
R13097 check[5].n12 check[5].n11 0.00481511
R13098 check[5].n13 check[5].n2 0.00215119
R13099 VSS_SW[4].n3 VSS_SW[4].n0 585
R13100 VSS_SW[4].n2 VSS_SW[4].t0 417.519
R13101 VSS_SW[4].n1 VSS_SW[4].t1 117.424
R13102 VSS_SW[4].n4 VSS_SW[4].n0 73.2739
R13103 VSS_SW[4].t0 VSS_SW[4].n0 71.9813
R13104 VSS_SW[4] VSS_SW[4].n1 67.6928
R13105 VSS_SW[4].n3 VSS_SW[4].n2 12.8005
R13106 VSS_SW[4].n1 VSS_SW[4] 6.64665
R13107 VSS_SW[4] VSS_SW[4].n4 3.04482
R13108 VSS_SW[4] VSS_SW[4].n3 2.21588
R13109 VSS_SW[4].n4 VSS_SW[4] 1.9648
R13110 VSS_SW[4].n2 VSS_SW[4] 1.72358
R13111 VSS_SW[6].n3 VSS_SW[6].n0 585
R13112 VSS_SW[6].n2 VSS_SW[6].t0 417.519
R13113 VSS_SW[6].n1 VSS_SW[6].t1 117.424
R13114 VSS_SW[6].n4 VSS_SW[6].n0 73.2739
R13115 VSS_SW[6].t0 VSS_SW[6].n0 71.9813
R13116 VSS_SW[6] VSS_SW[6].n1 67.6928
R13117 VSS_SW[6].n3 VSS_SW[6].n2 12.8005
R13118 VSS_SW[6].n1 VSS_SW[6] 6.64665
R13119 VSS_SW[6] VSS_SW[6].n4 3.04482
R13120 VSS_SW[6] VSS_SW[6].n3 2.21588
R13121 VSS_SW[6].n4 VSS_SW[6] 1.9648
R13122 VSS_SW[6].n2 VSS_SW[6] 1.72358
R13123 VDD_SW_b[7].n3 VDD_SW_b[7].t1 117.424
R13124 VDD_SW_b[7].n0 VDD_SW_b[7].t0 102.686
R13125 VDD_SW_b[7].n4 VDD_SW_b[7].n3 76.2952
R13126 VDD_SW_b[7].n0 VDD_SW_b[7] 10.3552
R13127 VDD_SW_b[7].n6 VDD_SW_b[7].n4 9.3005
R13128 VDD_SW_b[7].n3 VDD_SW_b[7] 5.61454
R13129 VDD_SW_b[7].n6 VDD_SW_b[7].n2 4.5005
R13130 VDD_SW_b[7].n1 VDD_SW_b[7].n0 3.87653
R13131 VDD_SW_b[7].n10 VDD_SW_b[7] 3.65824
R13132 VDD_SW_b[7].n4 VDD_SW_b[7] 3.14436
R13133 VDD_SW_b[7] VDD_SW_b[7].n10 2.95483
R13134 VDD_SW_b[7].n8 VDD_SW_b[7].n7 1.50505
R13135 VDD_SW_b[7].n2 VDD_SW_b[7].n1 0.449623
R13136 VDD_SW_b[7] VDD_SW_b[7].n2 0.225061
R13137 VDD_SW_b[7].n10 VDD_SW_b[7].n9 0.0501381
R13138 VDD_SW_b[7].n9 VDD_SW_b[7].n8 0.0260996
R13139 VDD_SW_b[7].n6 VDD_SW_b[7].n5 0.0122188
R13140 VDD_SW_b[7].n7 VDD_SW_b[7].n6 0.00814977
R13141 VDD_SW_b[2].n3 VDD_SW_b[2].t1 117.424
R13142 VDD_SW_b[2].n0 VDD_SW_b[2].t0 102.686
R13143 VDD_SW_b[2].n4 VDD_SW_b[2].n3 76.2952
R13144 VDD_SW_b[2].n0 VDD_SW_b[2] 10.3552
R13145 VDD_SW_b[2].n6 VDD_SW_b[2].n4 9.3005
R13146 VDD_SW_b[2].n3 VDD_SW_b[2] 5.61454
R13147 VDD_SW_b[2].n6 VDD_SW_b[2].n2 4.5005
R13148 VDD_SW_b[2].n1 VDD_SW_b[2].n0 3.87653
R13149 VDD_SW_b[2].n10 VDD_SW_b[2] 3.65824
R13150 VDD_SW_b[2].n4 VDD_SW_b[2] 3.14436
R13151 VDD_SW_b[2] VDD_SW_b[2].n10 2.95483
R13152 VDD_SW_b[2].n8 VDD_SW_b[2].n7 1.50505
R13153 VDD_SW_b[2].n2 VDD_SW_b[2].n1 0.449623
R13154 VDD_SW_b[2] VDD_SW_b[2].n2 0.225061
R13155 VDD_SW_b[2].n10 VDD_SW_b[2].n9 0.0501381
R13156 VDD_SW_b[2].n9 VDD_SW_b[2].n8 0.0260996
R13157 VDD_SW_b[2].n6 VDD_SW_b[2].n5 0.0122188
R13158 VDD_SW_b[2].n7 VDD_SW_b[2].n6 0.00814977
R13159 VSS_SW[1].n3 VSS_SW[1].n0 585
R13160 VSS_SW[1].n2 VSS_SW[1].t0 417.519
R13161 VSS_SW[1].n1 VSS_SW[1].t1 117.424
R13162 VSS_SW[1].n4 VSS_SW[1].n0 73.2739
R13163 VSS_SW[1].t0 VSS_SW[1].n0 71.9813
R13164 VSS_SW[1] VSS_SW[1].n1 67.6928
R13165 VSS_SW[1].n3 VSS_SW[1].n2 12.8005
R13166 VSS_SW[1].n1 VSS_SW[1] 6.64665
R13167 VSS_SW[1] VSS_SW[1].n4 3.11587
R13168 VSS_SW[1] VSS_SW[1].n3 2.21588
R13169 VSS_SW[1].n4 VSS_SW[1] 1.9648
R13170 VSS_SW[1].n2 VSS_SW[1] 1.72358
R13171 VSS_SW[7].n3 VSS_SW[7].n0 585
R13172 VSS_SW[7].n2 VSS_SW[7].t0 417.519
R13173 VSS_SW[7].n1 VSS_SW[7].t1 117.424
R13174 VSS_SW[7].n4 VSS_SW[7].n0 73.2739
R13175 VSS_SW[7].t0 VSS_SW[7].n0 71.9813
R13176 VSS_SW[7] VSS_SW[7].n1 67.6928
R13177 VSS_SW[7].n3 VSS_SW[7].n2 12.8005
R13178 VSS_SW[7].n1 VSS_SW[7] 6.64665
R13179 VSS_SW[7] VSS_SW[7].n4 3.04482
R13180 VSS_SW[7] VSS_SW[7].n3 2.21588
R13181 VSS_SW[7].n4 VSS_SW[7] 1.9648
R13182 VSS_SW[7].n2 VSS_SW[7] 1.72358
R13183 VSS_SW_b[6].n4 VSS_SW_b[6].n3 641.827
R13184 VSS_SW_b[6] VSS_SW_b[6].t0 422.656
R13185 VSS_SW_b[6].t0 VSS_SW_b[6].n5 121.231
R13186 VSS_SW_b[6].n2 VSS_SW_b[6].t1 117.424
R13187 VSS_SW_b[6].n3 VSS_SW_b[6].n2 77.418
R13188 VSS_SW_b[6].n6 VSS_SW_b[6] 11.3827
R13189 VSS_SW_b[6].n5 VSS_SW_b[6].n0 9.15497
R13190 VSS_SW_b[6].n5 VSS_SW_b[6].n4 7.57742
R13191 VSS_SW_b[6].n2 VSS_SW_b[6] 5.61454
R13192 VSS_SW_b[6].n8 VSS_SW_b[6].n6 2.47092
R13193 VSS_SW_b[6].n3 VSS_SW_b[6] 2.02155
R13194 VSS_SW_b[6].n12 VSS_SW_b[6] 1.6999
R13195 VSS_SW_b[6].n6 VSS_SW_b[6].n0 1.50964
R13196 VSS_SW_b[6].n10 VSS_SW_b[6].n9 1.5083
R13197 VSS_SW_b[6] VSS_SW_b[6].n12 1.3731
R13198 VSS_SW_b[6] VSS_SW_b[6].n1 1.34787
R13199 VSS_SW_b[6].n1 VSS_SW_b[6].n0 0.449623
R13200 VSS_SW_b[6].n12 VSS_SW_b[6].n11 0.0501381
R13201 VSS_SW_b[6].n11 VSS_SW_b[6].n10 0.0260996
R13202 VSS_SW_b[6].n8 VSS_SW_b[6].n7 0.0219844
R13203 VSS_SW_b[6].n9 VSS_SW_b[6].n8 0.00489987
R13204 VDD_SW_b[3].n3 VDD_SW_b[3].t1 117.424
R13205 VDD_SW_b[3].n0 VDD_SW_b[3].t0 100.715
R13206 VDD_SW_b[3].n4 VDD_SW_b[3].n3 76.5198
R13207 VDD_SW_b[3].n0 VDD_SW_b[3] 10.2646
R13208 VDD_SW_b[3].n6 VDD_SW_b[3].n4 9.3005
R13209 VDD_SW_b[3].n3 VDD_SW_b[3] 5.61454
R13210 VDD_SW_b[3].n6 VDD_SW_b[3].n2 4.5005
R13211 VDD_SW_b[3].n1 VDD_SW_b[3].n0 3.75113
R13212 VDD_SW_b[3].n10 VDD_SW_b[3] 3.66121
R13213 VDD_SW_b[3] VDD_SW_b[3].n10 2.95723
R13214 VDD_SW_b[3].n4 VDD_SW_b[3] 2.9198
R13215 VDD_SW_b[3].n8 VDD_SW_b[3].n7 1.5044
R13216 VDD_SW_b[3].n2 VDD_SW_b[3].n1 0.449623
R13217 VDD_SW_b[3] VDD_SW_b[3].n2 0.449623
R13218 VDD_SW_b[3].n10 VDD_SW_b[3].n9 0.0501381
R13219 VDD_SW_b[3].n9 VDD_SW_b[3].n8 0.0260996
R13220 VDD_SW_b[3].n6 VDD_SW_b[3].n5 0.0102656
R13221 VDD_SW_b[3].n7 VDD_SW_b[3].n6 0.00879975
R13222 VSS_SW[2].n3 VSS_SW[2].n0 585
R13223 VSS_SW[2].n2 VSS_SW[2].t0 417.519
R13224 VSS_SW[2].n1 VSS_SW[2].t1 117.424
R13225 VSS_SW[2].n4 VSS_SW[2].n0 73.2739
R13226 VSS_SW[2].t0 VSS_SW[2].n0 71.9813
R13227 VSS_SW[2] VSS_SW[2].n1 67.6928
R13228 VSS_SW[2].n3 VSS_SW[2].n2 12.8005
R13229 VSS_SW[2].n1 VSS_SW[2] 6.64665
R13230 VSS_SW[2] VSS_SW[2].n4 3.11587
R13231 VSS_SW[2] VSS_SW[2].n3 2.21588
R13232 VSS_SW[2].n4 VSS_SW[2] 1.9648
R13233 VSS_SW[2].n2 VSS_SW[2] 1.72358
R13234 VSS_SW_b[1].n4 VSS_SW_b[1].n3 641.827
R13235 VSS_SW_b[1] VSS_SW_b[1].t0 422.656
R13236 VSS_SW_b[1].t0 VSS_SW_b[1].n5 121.231
R13237 VSS_SW_b[1].n2 VSS_SW_b[1].t1 117.424
R13238 VSS_SW_b[1].n3 VSS_SW_b[1].n2 77.418
R13239 VSS_SW_b[1].n6 VSS_SW_b[1] 11.3827
R13240 VSS_SW_b[1].n5 VSS_SW_b[1].n0 9.15497
R13241 VSS_SW_b[1].n5 VSS_SW_b[1].n4 7.57742
R13242 VSS_SW_b[1].n2 VSS_SW_b[1] 5.61454
R13243 VSS_SW_b[1].n8 VSS_SW_b[1].n6 2.47092
R13244 VSS_SW_b[1].n3 VSS_SW_b[1] 2.02155
R13245 VSS_SW_b[1].n12 VSS_SW_b[1] 1.6999
R13246 VSS_SW_b[1].n6 VSS_SW_b[1].n0 1.50964
R13247 VSS_SW_b[1].n10 VSS_SW_b[1].n9 1.5083
R13248 VSS_SW_b[1] VSS_SW_b[1].n12 1.3731
R13249 VSS_SW_b[1] VSS_SW_b[1].n1 1.34787
R13250 VSS_SW_b[1].n1 VSS_SW_b[1].n0 0.449623
R13251 VSS_SW_b[1].n12 VSS_SW_b[1].n11 0.0501381
R13252 VSS_SW_b[1].n11 VSS_SW_b[1].n10 0.0260996
R13253 VSS_SW_b[1].n8 VSS_SW_b[1].n7 0.0219844
R13254 VSS_SW_b[1].n9 VSS_SW_b[1].n8 0.00489987
R13255 VDD_SW_b[4].n3 VDD_SW_b[4].t1 117.424
R13256 VDD_SW_b[4].n0 VDD_SW_b[4].t0 100.715
R13257 VDD_SW_b[4].n4 VDD_SW_b[4].n3 76.5198
R13258 VDD_SW_b[4].n0 VDD_SW_b[4] 10.2646
R13259 VDD_SW_b[4].n6 VDD_SW_b[4].n4 9.3005
R13260 VDD_SW_b[4].n3 VDD_SW_b[4] 5.61454
R13261 VDD_SW_b[4].n6 VDD_SW_b[4].n2 4.5005
R13262 VDD_SW_b[4].n1 VDD_SW_b[4].n0 3.75113
R13263 VDD_SW_b[4].n10 VDD_SW_b[4] 3.66419
R13264 VDD_SW_b[4] VDD_SW_b[4].n10 2.95963
R13265 VDD_SW_b[4].n4 VDD_SW_b[4] 2.9198
R13266 VDD_SW_b[4].n8 VDD_SW_b[4].n7 1.50505
R13267 VDD_SW_b[4] VDD_SW_b[4].n2 0.674184
R13268 VDD_SW_b[4].n2 VDD_SW_b[4].n1 0.225061
R13269 VDD_SW_b[4].n10 VDD_SW_b[4].n9 0.0501381
R13270 VDD_SW_b[4].n9 VDD_SW_b[4].n8 0.0260996
R13271 VDD_SW_b[4].n6 VDD_SW_b[4].n5 0.0122188
R13272 VDD_SW_b[4].n7 VDD_SW_b[4].n6 0.00814977
R13273 VDD_SW[3].n8 VDD_SW[3].t1 117.424
R13274 VDD_SW[3].n6 VDD_SW[3].t0 75.7697
R13275 VDD_SW[3].n7 VDD_SW[3].n6 73.0808
R13276 VDD_SW[3] VDD_SW[3].n8 67.6928
R13277 VDD_SW[3].n10 VDD_SW[3].n9 13.0467
R13278 VDD_SW[3].n8 VDD_SW[3] 6.64665
R13279 VDD_SW[3].n5 VDD_SW[3].n4 2.82795
R13280 VDD_SW[3] VDD_SW[3].n7 2.2023
R13281 VDD_SW[3] VDD_SW[3].n10 1.96973
R13282 VDD_SW[3].n9 VDD_SW[3] 1.72358
R13283 VDD_SW[3].n3 VDD_SW[3].n1 1.49691
R13284 VDD_SW[3].n1 VDD_SW[3] 0.0595299
R13285 VDD_SW[3].n1 VDD_SW[3].n0 0.0177811
R13286 VDD_SW[3].n7 VDD_SW[3].n5 0.0146776
R13287 VDD_SW[3].n3 VDD_SW[3].n2 0.0102656
R13288 VDD_SW[3].n4 VDD_SW[3].n3 0.00635152
C0 x9.A1 a_14545_627# 2.37e-19
C1 check[2] m1_95_2154# 0.0352f
C2 a_27_627# VDD_SW[7] 3.29e-20
C3 D[7] a_1363_627# 2e-19
C4 check[5] a_3421_n88# 2.51e-20
C5 a_12901_601# a_14545_627# 5.92e-20
C6 a_720_106# a_977_304# 0.00857f
C7 a_487_n62# a_1166_304# 0.00652f
C8 D[7] a_557_993# 8.11e-19
C9 a_27_627# a_891_909# 2.46e-19
C10 VDD a_8731_627# 0.0174f
C11 a_11546_1315# VDD_SW_b[3] 3.97e-20
C12 D[4] a_10509_601# 3.09e-21
C13 a_8140_n62# a_8545_n62# 2.46e-21
C14 x8.X a_941_601# 0.00123f
C15 x13.X a_8933_1315# 2.09e-19
C16 x2.X a_12638_220# 0.0028f
C17 a_12134_n88# a_12553_n62# 0.0383f
C18 x2.X a_2419_627# 0.355f
C19 VDD a_5365_627# 1.44e-20
C20 check[4] a_5725_601# 1.55e-19
C21 a_11514_n62# VSS_SW_b[2] 2.8e-19
C22 a_14857_1289# a_14825_993# 4.54e-19
C23 a_14545_627# a_14909_993# 0.0018f
C24 a_14999_601# a_14733_627# 8.07e-20
C25 a_15293_601# a_15767_895# 0.265f
C26 x9.A1 a_9122_n62# 1.9e-20
C27 VDD_SW_b[3] a_10597_n88# 0.0406f
C28 a_5813_n88# a_8204_212# 4.92e-22
C29 a_7615_1315# D[4] 0.00202f
C30 a_5812_212# a_8205_n88# 5.48e-21
C31 x2.X m1_95_2154# 6.31f
C32 x2.X a_535_1642# 2.63e-19
C33 a_1233_n88# a_1143_n62# 9.75e-19
C34 VSS_SW_b[7] a_593_n62# 0.00335f
C35 a_1028_212# VSS_SW[6] 0.0872f
C36 a_1029_n88# a_1369_n62# 6.04e-20
C37 x10.X a_4149_1315# 1.78e-20
C38 a_193_627# a_2136_627# 2.2e-20
C39 VSS_SW[1] VSS_SW_b[1] 0.00717f
C40 a_4413_2457# m1_95_2154# 1.41e-19
C41 VDD a_10824_993# 0.189f
C42 a_9595_627# a_10801_n88# 0.00204f
C43 x9.A1 a_4860_1467# 0.197f
C44 a_4811_627# a_5813_n88# 1.06e-19
C45 D[5] a_5812_212# 0.157f
C46 a_473_993# a_941_601# 0.0633f
C47 a_193_627# a_1256_993# 0.0334f
C48 a_8432_993# VDD_SW[4] 3.28e-20
C49 VDD_SW_b[2] a_12988_212# 0.0416f
C50 a_4860_1467# a_5002_1315# 0.00783f
C51 a_13461_1642# a_12988_212# 1.39e-21
C52 VDD a_2610_1642# 0.00363f
C53 x2.X a_3558_304# 0.00338f
C54 a_2419_627# a_4977_627# 1.09e-20
C55 a_2585_627# a_4811_627# 1.36e-20
C56 VDD a_15721_n62# 0.0301f
C57 a_2419_627# VSS_SW[5] 4.66e-21
C58 a_7203_627# D[4] 0.138f
C59 a_7203_627# VSS_SW[4] 0.0576f
C60 x9.A1 a_1415_895# 2.64e-19
C61 a_14428_1467# m1_95_2154# 8.35e-20
C62 x2.X a_1112_909# 0.00309f
C63 VDD a_9154_1315# 0.00109f
C64 a_4977_627# m1_95_2154# 2.61e-20
C65 a_891_909# VDD_SW[7] 1.01e-20
C66 a_4811_627# a_6920_627# 1.75e-19
C67 VSS_SW[5] m1_95_2154# 0.0337f
C68 a_76_1467# check[6] 0.318f
C69 a_647_601# VDD_SW_b[7] 1.36e-20
C70 a_941_601# a_1159_627# 3.73e-19
C71 a_1256_993# a_791_627# 0.00316f
C72 x7.X a_3333_601# 4.31e-21
C73 x16.X a_12465_1289# 1.54e-19
C74 a_10055_n62# a_10596_212# 0.138f
C75 x12.X a_7369_627# 0.00315f
C76 x2.X a_4149_1642# 5.23e-19
C77 x2.X a_5257_993# 0.15f
C78 a_9122_n62# a_9742_n88# 8.26e-21
C79 a_4413_2457# a_4149_1642# 9.92e-19
C80 a_12988_212# a_15072_106# 5.86e-20
C81 a_12989_n88# a_14839_n62# 4.56e-21
C82 a_4689_2457# x9.A1 5.5e-19
C83 a_3420_212# VSS_SW_b[5] 0.00377f
C84 a_9312_627# m1_95_2154# 1.66e-20
C85 a_3558_304# VSS_SW[5] 2.76e-20
C86 a_1503_1642# a_941_601# 0.00263f
C87 check[6] a_174_n88# 5.27e-19
C88 x9.A1 a_11514_n62# 1.9e-20
C89 x9.A1 VDD_SW_b[7] 1.17e-20
C90 a_3333_601# a_3420_212# 6.03e-19
C91 a_2773_627# a_2566_n88# 3.32e-19
C92 a_3648_993# a_2879_n62# 3.59e-19
C93 check[4] a_5271_n62# 1.31e-20
C94 x9.A1 a_6285_1642# 0.101f
C95 VDD a_1757_1642# 0.115f
C96 x2.X a_8539_627# 0.00111f
C97 check[3] a_7681_1289# 0.249f
C98 a_2468_1467# x8.X 0.0876f
C99 x9.A1 check[5] 0.412f
C100 VDD a_2773_627# 0.126f
C101 a_8933_1642# a_9644_1467# 0.00963f
C102 a_12433_993# m1_95_1942# 2.74e-20
C103 a_3895_1642# a_3893_122# 1.57e-21
C104 a_487_n62# a_2566_n88# 5.13e-21
C105 a_11987_627# m1_95_2154# 3.53e-20
C106 a_4977_627# a_5257_993# 0.15f
C107 x2.X a_5943_627# 0.00702f
C108 VDD_SW_b[3] m1_95_2154# 1.28e-20
C109 a_5257_993# VSS_SW[5] 0.003f
C110 a_12901_601# a_12751_627# 0.00926f
C111 a_12153_627# a_13632_909# 7.17e-20
C112 a_13216_993# a_13072_909# 0.00412f
C113 a_12433_993# a_12541_627# 0.00807f
C114 a_12465_1289# a_12153_627# 0.00323f
C115 a_12607_601# a_13119_627# 9.75e-19
C116 a_8117_601# a_9595_627# 3.84e-19
C117 VDD a_487_n62# 0.348f
C118 a_193_627# VSS_SW[7] 0.023f
C119 x15.X D[2] 2.14e-19
C120 a_7663_n62# VSS_SW_b[3] 1.03e-20
C121 a_11325_1315# D[3] 0.00195f
C122 a_4689_2457# a_5323_2457# 8.37e-20
C123 VDD_SW_b[6] a_3112_106# 5.23e-19
C124 a_6285_1642# a_6040_993# 0.00181f
C125 a_15855_1642# m1_95_1942# 2.26e-19
C126 x2.X a_11313_304# 3.34e-19
C127 check[6] a_2897_1289# 3.63e-21
C128 check[0] a_15721_n62# 9.72e-20
C129 VSS_SW[2] a_12134_n88# 0.00676f
C130 a_76_1467# D[7] 0.0183f
C131 x2.X a_5289_1289# 0.0112f
C132 a_5323_2457# a_6285_1642# 0.00184f
C133 a_6730_n62# a_8204_212# 2.79e-22
C134 a_14379_627# a_15293_601# 0.14f
C135 D[1] a_14825_993# 0.00887f
C136 x9.A1 VDD_SW_b[1] 1.67e-20
C137 x9.A1 x20.X 5.49e-19
C138 a_1233_n88# VSS_SW_b[6] 4.54e-20
C139 a_10801_n88# VSS_SW[2] 8.39e-20
C140 VSS_SW_b[3] a_10711_n62# 5.24e-19
C141 VDD_SW_b[2] a_15293_601# 8.35e-20
C142 a_1946_n62# VSS_SW[6] 6.09e-20
C143 a_11069_122# a_10937_n62# 0.025f
C144 a_27_627# a_2773_627# 4.46e-21
C145 a_5257_993# a_5575_627# 0.025f
C146 a_4977_627# a_5943_627# 2.14e-20
C147 a_5725_601# a_6124_993# 9.41e-19
C148 a_5165_627# a_5341_993# 8.99e-19
C149 D[5] a_6529_304# 8.39e-19
C150 a_10983_895# a_10596_212# 0.00165f
C151 a_10509_601# a_10597_n88# 3.89e-19
C152 a_2897_1289# a_2879_n62# 3.44e-19
C153 x8.X a_3039_601# 2.4e-20
C154 D[3] a_10596_212# 0.158f
C155 VDD a_10734_304# 0.0164f
C156 a_791_627# VSS_SW[7] 0.0012f
C157 a_14430_90# a_14526_n88# 0.0967f
C158 x9.X x10.X 0.111f
C159 VSS_SW_b[2] a_13705_n62# 6.93e-20
C160 x2.X a_13300_993# 4.66e-19
C161 a_27_627# a_487_n62# 7.27e-19
C162 D[7] a_174_n88# 0.00506f
C163 x2.X a_4958_n88# 0.178f
C164 a_12036_1467# a_12038_90# 1e-19
C165 x9.A1 a_11123_627# 5.3e-20
C166 a_6539_1642# check[3] 1.64e-19
C167 VDD_SW[3] a_12607_601# 7.64e-20
C168 a_4149_1642# a_4370_1315# 0.00783f
C169 x9.A1 x12.X 0.00117f
C170 a_5289_1289# a_4977_627# 0.00323f
C171 D[6] a_3807_895# 0.0294f
C172 a_2419_627# a_3648_993# 0.14f
C173 VDD a_5462_220# 0.00458f
C174 x15.X a_10055_n62# 0.002f
C175 x9.X D[5] 2.11e-19
C176 a_5289_1289# VSS_SW[5] 0.00187f
C177 a_12036_1467# m1_95_1942# 1.97e-19
C178 VDD a_12851_909# 0.00988f
C179 VSS_SW_b[1] a_16097_n62# 6.94e-20
C180 a_5896_909# VDD_SW_b[5] 7.05e-21
C181 a_5575_627# a_5943_627# 3.34e-19
C182 a_9147_1642# VDD_SW[4] 5.38e-19
C183 a_76_1467# m1_95_2154# 4.76e-20
C184 a_14857_1289# a_14526_n88# 5.67e-21
C185 a_76_1467# a_535_1642# 6.64e-19
C186 a_15767_895# a_14839_n62# 0.00219f
C187 a_14999_601# a_15381_n88# 0.00322f
C188 a_14545_627# a_15585_n88# 8.75e-19
C189 a_15293_601# a_15072_106# 3.46e-19
C190 a_941_601# a_2585_627# 6.03e-20
C191 x2.X a_16024_909# 4.02e-19
C192 VDD a_29_2457# 0.222f
C193 a_3807_895# m1_95_1942# 8.62e-20
C194 x13.X a_8204_212# 0.245f
C195 a_3648_993# m1_95_2154# 4.11e-21
C196 a_13216_993# VDD_SW[2] 3.28e-20
C197 reset m1_95_1942# 2.37e-20
C198 x9.A1 a_6285_122# 3.53e-20
C199 a_4977_627# a_4958_n88# 4.91e-19
C200 a_29_2457# x6.X 6.01e-21
C201 VSS_SW[5] a_4958_n88# 0.00686f
C202 a_2897_1289# D[7] 5.1e-21
C203 x12.X a_6040_993# 2.81e-19
C204 VDD a_12399_1315# 0.00136f
C205 VDD a_14933_627# 9.37e-19
C206 x9.A1 a_2865_993# 1.16e-19
C207 VDD D[4] 1.22f
C208 x2.X a_2949_993# 5.29e-19
C209 a_1757_1642# VDD_SW[7] 0.00511f
C210 x11.X a_6017_n88# 1.87e-19
C211 x2.X a_11704_627# 3.88e-19
C212 D[6] VDD_SW_b[6] 0.453f
C213 a_16488_627# m1_95_1942# 2.45e-20
C214 VDD VSS_SW[4] 0.608f
C215 a_12988_212# a_13461_122# 0.159f
C216 VSS_SW[2] a_12937_304# 8.24e-20
C217 a_12989_n88# a_13193_n88# 0.117f
C218 a_12680_106# VSS_SW_b[2] 0.00322f
C219 a_6285_1642# a_5812_212# 1.39e-21
C220 VDD_SW[7] a_2773_627# 6.11e-20
C221 VDD_SW[2] a_15464_909# 2.77e-20
C222 x18.X a_15293_601# 4.9e-20
C223 VDD a_4528_627# 0.194f
C224 x2.X a_720_106# 0.0385f
C225 a_2831_1315# D[6] 0.00202f
C226 a_1028_212# a_1745_n62# 0.00206f
C227 VDD_SW_b[6] m1_95_1942# 1.99e-20
C228 a_9595_627# a_10125_993# 4.45e-20
C229 D[3] a_9949_627# 0.161f
C230 check[3] VSS_SW[3] 1.4e-19
C231 a_29_2457# a_27_627# 1.01e-19
C232 a_1555_627# a_1028_212# 7.07e-21
C233 a_6040_993# a_6285_122# 1.51e-20
C234 a_5575_627# a_4958_n88# 1.08e-19
C235 a_2897_1289# a_2419_627# 0.00104f
C236 a_1415_895# a_1233_n88# 4.26e-19
C237 a_941_601# a_1501_122# 2.7e-19
C238 VDD a_1447_220# 0.00986f
C239 x7.X VSS_SW[6] 0.138f
C240 check[3] m1_95_1942# 0.034f
C241 a_11325_1642# VDD_SW[3] 0.00506f
C242 a_8117_601# a_10041_993# 1.29e-20
C243 a_8342_304# VSS_SW_b[3] 8.9e-21
C244 a_10509_601# m1_95_2154# 2.82e-20
C245 a_3807_895# a_5725_601# 1.38e-20
C246 D[2] a_13072_909# 8.51e-19
C247 a_11987_627# a_13300_993# 2.13e-19
C248 ready VDD_SW[6] 0.00397f
C249 D[4] a_7733_993# 8.11e-19
C250 a_7203_627# a_8067_909# 2.46e-19
C251 a_2897_1289# m1_95_2154# 1.04e-19
C252 x15.X a_10983_895# 0.0066f
C253 x15.X D[3] 0.0855f
C254 a_7350_n88# a_8677_122# 4.59e-22
C255 a_7896_106# a_8205_n88# 0.0327f
C256 a_7663_n62# a_8409_n88# 0.199f
C257 VSS_SW[6] a_3420_212# 1.18e-21
C258 a_6199_895# VDD_SW[5] 0.00356f
C259 check[1] m1_95_2154# 0.0352f
C260 a_6040_993# a_6147_627# 0.00707f
C261 a_15143_627# VSS_SW[1] 0.0012f
C262 a_13715_1315# D[2] 0.00195f
C263 VDD_SW_b[7] a_1233_n88# 0.00132f
C264 a_12465_1289# a_13461_1642# 0.0146f
C265 a_10596_212# a_10545_304# 2.13e-19
C266 a_10597_n88# a_10246_220# 4.48e-20
C267 a_13632_909# VDD_SW_b[2] 3.14e-20
C268 a_10288_106# a_10734_304# 0.00412f
C269 a_10055_n62# a_11015_220# 1.21e-20
C270 D[7] a_1166_304# 9.67e-19
C271 x2.X a_5761_304# 0.00166f
C272 VDD_SW_b[6] a_5725_601# 5.2e-20
C273 VSS_SW_b[2] a_13407_220# 1.2e-20
C274 a_13461_122# a_13705_304# 0.00972f
C275 a_13193_n88# a_13906_n62# 8.07e-20
C276 a_12989_n88# a_14430_90# 5.39e-19
C277 a_13375_895# a_12447_n62# 0.00219f
C278 a_12153_627# a_13193_n88# 8.75e-19
C279 a_12901_601# a_12680_106# 3.46e-19
C280 a_12607_601# a_12989_n88# 0.00322f
C281 x3.A x2.X 2.91e-19
C282 a_11704_627# a_11987_627# 0.0011f
C283 a_7203_627# m1_95_2154# 3.53e-20
C284 a_305_2457# ready 0.0596f
C285 VDD_SW_b[3] a_11704_627# 0.185f
C286 x3.X a_939_2457# 0.619f
C287 x9.A1 VSS_SW_b[3] 2.86e-19
C288 a_4860_1467# x9.X 4.97e-19
C289 VDD_SW_b[5] VDD_SW[5] 3.63e-19
C290 check[2] a_11069_122# 5.3e-20
C291 a_15381_n88# m1_95_1942# 1.16e-21
C292 x13.X a_10596_212# 8.4e-22
C293 check[3] VDD_SW[4] 0.00393f
C294 a_14379_627# a_14839_n62# 7.27e-19
C295 D[1] a_14526_n88# 0.00508f
C296 a_5504_106# VSS_SW_b[5] 0.00321f
C297 a_5812_212# a_6285_122# 0.159f
C298 VSS_SW[5] a_5761_304# 8.37e-20
C299 a_5813_n88# a_6017_n88# 0.117f
C300 a_9644_1467# a_9786_1642# 0.00557f
C301 D[2] VDD_SW[2] 0.246f
C302 VSS_SW[7] a_1029_n88# 9.29e-21
C303 x16.X a_12607_601# 2.69e-20
C304 x2.X a_3947_627# 0.0151f
C305 D[4] a_10288_106# 1.39e-21
C306 a_6539_1315# D[5] 0.00195f
C307 x11.X a_7254_90# 0.0273f
C308 x2.X a_12447_n62# 0.371f
C309 VDD check[6] 1.85f
C310 a_8591_895# a_7663_n62# 0.00219f
C311 a_7369_627# a_8409_n88# 8.75e-19
C312 VDD a_11546_1315# 0.00115f
C313 a_8117_601# a_7896_106# 3.46e-19
C314 a_7823_601# a_8205_n88# 0.00322f
C315 a_2585_627# a_3039_601# 0.117f
C316 x2.X a_1745_304# 3.34e-19
C317 VDD_SW_b[1] a_15585_n88# 0.00131f
C318 x2.X a_11069_122# 0.0043f
C319 x20.X a_15585_n88# 1.87e-19
C320 a_1946_n62# a_1745_n62# 3.81e-19
C321 a_2566_n88# a_2879_n62# 0.245f
C322 a_11514_n62# VSS_SW[2] 6.06e-20
C323 x6.X check[6] 0.00903f
C324 a_10215_601# a_10459_909# 0.0104f
C325 a_10041_993# a_10125_993# 0.00972f
C326 D[3] a_11015_220# 7.13e-19
C327 VDD a_2879_n62# 0.367f
C328 x14.X a_7369_627# 6.29e-20
C329 a_193_627# VSS_SW[6] 5.36e-21
C330 a_10215_601# VSS_SW[3] 6.23e-19
C331 a_14839_n62# a_15072_106# 0.124f
C332 a_14526_n88# a_15380_212# 0.0319f
C333 check[4] a_6467_1642# 0.00577f
C334 a_9742_n88# VSS_SW_b[3] 0.135f
C335 VDD a_10597_n88# 0.699f
C336 a_10215_601# m1_95_1942# 3.42e-20
C337 D[4] a_8731_627# 0.00431f
C338 check[5] x9.X 0.00967f
C339 a_8204_212# a_10596_212# 9.5e-22
C340 a_12153_627# a_12607_601# 0.117f
C341 a_12751_627# VSS_SW[2] 0.0012f
C342 VDD_SW_b[4] a_7663_n62# 5.22e-19
C343 a_8205_n88# a_8623_220# 0.00276f
C344 a_7350_n88# a_7769_n62# 0.0383f
C345 a_8204_212# a_8921_304# 4.45e-20
C346 x9.A1 a_8679_1642# 0.101f
C347 VSS_SW_b[4] a_7854_220# 5.34e-20
C348 a_8409_n88# a_8342_304# 9.46e-19
C349 a_7663_n62# a_9646_90# 6.12e-21
C350 a_3333_601# a_3504_909# 0.00652f
C351 check[6] a_27_627# 0.00121f
C352 a_3039_601# a_3183_627# 0.0697f
C353 a_3625_n88# VSS_SW_b[6] 9.21e-19
C354 check[3] a_10073_1289# 3.63e-21
C355 VDD_SW_b[5] a_5748_n62# 8.12e-20
C356 VDD_SW_b[7] a_593_n62# 4.77e-19
C357 D[7] a_2566_n88# 4.33e-19
C358 a_11325_1642# x16.X 7.78e-19
C359 x9.A1 a_14825_993# 8.95e-20
C360 VDD_SW[6] a_5896_909# 2.77e-20
C361 a_13216_993# a_14545_627# 4.03e-21
C362 a_12901_601# a_14825_993# 1.11e-20
C363 x17.X D[2] 0.0854f
C364 a_174_n88# a_720_106# 0.207f
C365 VDD D[7] 1.06f
C366 VDD a_8067_909# 0.00984f
C367 x2.X a_13126_304# 0.00338f
C368 a_3283_909# VDD_SW_b[6] 3.01e-21
C369 VDD a_6529_n62# 2.27e-19
C370 a_12680_106# a_12553_n62# 0.0256f
C371 a_12447_n62# a_12924_n62# 1.96e-20
C372 a_7369_627# a_8591_895# 0.0494f
C373 a_7823_601# a_8117_601# 0.199f
C374 a_11987_627# a_12447_n62# 7.27e-19
C375 D[2] a_12134_n88# 0.00506f
C376 x6.X D[7] 0.00886f
C377 x2.X a_7681_1289# 0.0113f
C378 VDD_SW_b[1] a_14945_n62# 4.77e-19
C379 a_15293_601# a_14733_627# 1.24e-20
C380 a_15767_895# a_15608_993# 0.207f
C381 a_14999_601# a_15243_909# 0.0104f
C382 a_14825_993# a_14909_993# 0.00972f
C383 check[6] a_218_1642# 0.00688f
C384 a_14545_627# a_15464_909# 0.00907f
C385 a_15855_1642# a_15293_601# 0.00263f
C386 a_10509_601# a_11704_627# 5.73e-19
C387 a_2419_627# a_2566_n88# 0.00176f
C388 x10.X a_4862_90# 0.00259f
C389 VDD_SW_b[3] a_11069_122# 0.00446f
C390 VDD a_12638_220# 0.00643f
C391 a_9154_1315# D[4] 0.0012f
C392 x9.A1 a_8409_n88# 1.66e-20
C393 a_15072_106# a_15518_304# 0.00412f
C394 a_15381_n88# a_15030_220# 4.71e-20
C395 a_14839_n62# a_15799_220# 1.21e-20
C396 a_15380_212# a_15329_304# 2.13e-19
C397 a_5504_106# a_5748_n62# 0.00707f
C398 a_6017_n88# a_6730_n62# 8.07e-20
C399 a_5813_n88# a_7254_90# 5.39e-19
C400 a_6285_122# a_6529_304# 0.00972f
C401 a_5271_n62# a_5927_n62# 3.73e-19
C402 VSS_SW_b[5] a_6231_220# 1.12e-20
C403 VDD_SW[4] a_10215_601# 7.64e-20
C404 a_9595_627# VSS_SW_b[3] 1.08e-19
C405 VDD a_2419_627# 0.463f
C406 a_939_2457# x8.X 8.68e-19
C407 a_1501_122# VSS_SW_b[7] 7.15e-19
C408 x2.X a_14999_601# 0.2f
C409 x9.A1 a_7252_1467# 0.197f
C410 a_13461_1642# a_13193_n88# 4.63e-19
C411 check[6] VDD_SW[7] 0.00393f
C412 VDD_SW_b[2] a_13193_n88# 0.00132f
C413 VDD a_8545_n62# 0.0342f
C414 a_8933_1642# a_9147_1642# 0.00557f
C415 a_27_627# D[7] 0.138f
C416 VDD a_4077_1642# 8.63e-19
C417 x9.A1 x14.X 8.85e-19
C418 a_8432_993# a_8516_993# 0.00857f
C419 a_7369_627# VDD_SW_b[4] 0.00231f
C420 x3.A a_76_1467# 2.66e-20
C421 VDD m1_95_2154# 0.264f
C422 VDD a_535_1642# 0.0019f
C423 x11.X D[5] 0.1f
C424 x2.X a_3112_106# 0.0385f
C425 x12.X a_7394_1315# 8.34e-19
C426 x10.X a_5165_627# 6.12e-19
C427 a_10161_n62# a_10532_n62# 4.19e-20
C428 a_14096_627# m1_95_2154# 1.66e-20
C429 x17.X VSS_SW_b[1] 0.0172f
C430 a_10055_n62# a_12134_n88# 3.08e-21
C431 ready a_647_601# 3.47e-22
C432 VDD a_3558_304# 0.0224f
C433 a_305_2457# VSS_SW[7] 0.0177f
C434 a_27_627# a_2419_627# 1.63e-20
C435 D[5] a_5165_627# 0.161f
C436 a_4811_627# a_5341_993# 4.45e-20
C437 a_10055_n62# a_10801_n88# 0.199f
C438 a_10288_106# a_10597_n88# 0.0327f
C439 VDD a_1112_909# 0.0164f
C440 x2.X a_6539_1642# 5.27e-19
C441 a_12989_n88# a_15380_212# 8.02e-22
C442 a_12988_212# a_15381_n88# 5.48e-21
C443 a_8205_n88# a_10055_n62# 4.56e-21
C444 a_3333_601# VDD_SW[6] 1.79e-19
C445 a_3648_993# a_3947_627# 0.0256f
C446 ready x9.A1 3.55e-19
C447 a_27_627# m1_95_2154# 3.53e-20
C448 a_3420_212# a_3761_n62# 0.00134f
C449 a_3112_106# VSS_SW[5] 9.05e-21
C450 a_3421_n88# a_3535_n62# 2.14e-20
C451 a_14545_627# VDD_SW[1] 1.85e-20
C452 a_15293_601# a_16488_627# 5.84e-19
C453 x9.A1 a_5319_1642# 5.26e-19
C454 VDD a_5257_993# 0.195f
C455 VDD a_4149_1642# 0.115f
C456 a_10073_1289# a_10215_601# 8.76e-20
C457 check[3] a_7394_1642# 0.00688f
C458 check[2] VSS_SW[3] 0.0493f
C459 x9.A1 a_8591_895# 2.41e-19
C460 x2.X a_8288_909# 0.00309f
C461 a_13375_895# m1_95_1942# 8.63e-20
C462 x2.X a_7854_220# 0.00279f
C463 check[2] m1_95_1942# 0.034f
C464 D[7] VDD_SW[7] 0.227f
C465 a_14379_627# a_14430_90# 6.13e-19
C466 check[5] a_3625_n88# 2.51e-19
C467 a_720_106# a_1166_304# 0.00412f
C468 a_1028_212# a_977_304# 2.13e-19
C469 a_1029_n88# a_678_220# 4.48e-20
C470 a_487_n62# a_1447_220# 1.21e-20
C471 D[2] a_14545_627# 7.7e-21
C472 ready a_505_1289# 2.39e-20
C473 a_939_2457# a_1503_1642# 0.00188f
C474 VDD_SW_b[2] a_14430_90# 0.00345f
C475 D[7] a_891_909# 6.77e-19
C476 a_27_627# a_1112_909# 1.09e-19
C477 x11.X a_8117_601# 4.02e-21
C478 a_13216_993# a_12751_627# 0.00316f
C479 a_12465_1289# a_12433_993# 4.54e-19
C480 VDD a_8539_627# 0.00132f
C481 a_12901_601# a_13119_627# 3.73e-19
C482 a_12607_601# VDD_SW_b[2] 1.36e-20
C483 a_8319_n62# a_8545_n62# 3.34e-19
C484 a_4064_909# VDD_SW[6] 2.12e-20
C485 x8.X a_1415_895# 0.00864f
C486 x30.A x2.X 0.002f
C487 a_4413_2457# x30.A 6.66e-19
C488 x27.A a_4689_2457# 0.3f
C489 ready a_5323_2457# 4.34e-19
C490 x2.X D[6] 0.177f
C491 VDD a_5943_627# 0.00711f
C492 x2.X a_10459_909# 0.00138f
C493 x2.X a_12038_90# 0.00366f
C494 check[4] a_6199_895# 0.00218f
C495 VSS_SW[2] a_12680_106# 4.62e-19
C496 a_4413_2457# D[6] 0.0191f
C497 D[6] a_3070_220# 2.03e-20
C498 check[0] m1_95_2154# 0.0352f
C499 a_5725_601# a_7557_627# 2.42e-20
C500 a_6199_895# a_8432_993# 1.86e-21
C501 x9.A1 VDD_SW_b[4] 1.72e-20
C502 VDD_SW[7] a_2419_627# 0.0865f
C503 a_10596_212# a_11313_n62# 0.00206f
C504 x2.X VSS_SW[3] 0.0816f
C505 a_14857_1289# a_14379_627# 0.00104f
C506 D[1] a_15767_895# 0.0295f
C507 a_14379_627# a_15608_993# 0.14f
C508 D[3] a_12134_n88# 4.32e-19
C509 a_5813_n88# a_8205_n88# 1.33e-19
C510 a_5271_n62# VSS_SW_b[4] 8.69e-21
C511 x10.X a_2585_627# 6.35e-20
C512 VSS_SW_b[7] a_964_n62# 1.68e-19
C513 a_10983_895# a_10801_n88# 4.26e-19
C514 x2.X m1_95_1942# 0.251f
C515 a_1029_n88# VSS_SW[6] 9.23e-19
C516 a_1233_n88# a_1369_n62# 0.0697f
C517 a_10509_601# a_11069_122# 2.7e-19
C518 x15.X a_11325_1315# 1.98e-19
C519 D[3] a_10801_n88# 0.00547f
C520 a_4413_2457# m1_95_1942# 6.42e-20
C521 VDD a_11313_304# 0.00494f
C522 D[5] a_5813_n88# 0.159f
C523 a_13906_n62# a_15380_212# 5.58e-22
C524 a_4811_627# a_6017_n88# 0.00204f
C525 a_647_601# a_1256_993# 0.00189f
C526 a_193_627# a_381_627# 0.189f
C527 VDD_SW[7] m1_95_2154# 0.0327f
C528 x9.A1 a_14526_n88# 7.4e-19
C529 VDD a_5289_1289# 0.212f
C530 a_4860_1467# a_4862_90# 1e-19
C531 x8.X VDD_SW_b[7] 7.23e-19
C532 x2.X a_12541_627# 3.94e-19
C533 x30.A a_4977_627# 1.19e-21
C534 a_3895_1642# x10.X 1.14e-20
C535 check[1] a_12447_n62# 1.39e-20
C536 x30.A VSS_SW[5] 0.0445f
C537 x9.A1 VDD_SW[3] 0.0329f
C538 a_8933_1642# check[3] 0.318f
C539 VDD_SW[3] a_12901_601# 2.46e-20
C540 x2.X a_3839_220# 9.61e-19
C541 D[6] a_4977_627# 6.42e-21
C542 check[4] VDD_SW_b[5] 0.00213f
C543 D[6] VSS_SW[5] 4.85e-19
C544 a_15143_627# a_15511_627# 3.34e-19
C545 a_15464_909# VDD_SW_b[1] 9.36e-21
C546 x8.X check[5] 0.00903f
C547 x9.A1 a_2136_627# 2e-20
C548 x15.X a_10596_212# 0.245f
C549 D[4] VSS_SW[4] 0.118f
C550 a_5002_1642# VSS_SW[5] 0.00105f
C551 x2.X a_1340_993# 4.67e-19
C552 a_14428_1467# m1_95_1942# 1.97e-19
C553 x12.X a_6539_1315# 2.36e-20
C554 x9.A1 a_1256_993# 4.84e-21
C555 a_76_1467# a_218_1315# 0.00783f
C556 VDD a_13300_993# 0.00284f
C557 check[2] VDD_SW[4] 4.35e-19
C558 x14.X a_9595_627# 0.236f
C559 VDD a_4958_n88# 0.703f
C560 a_4977_627# m1_95_1942# 3.82e-20
C561 a_5431_601# m1_95_2154# 2.34e-20
C562 a_14545_627# VSS_SW_b[1] 1.51e-20
C563 a_14857_1289# a_15072_106# 5.3e-21
C564 a_15767_895# a_15380_212# 0.00165f
C565 a_15293_601# a_15381_n88# 3.89e-19
C566 VSS_SW[5] m1_95_1942# 0.033f
C567 a_1112_909# VDD_SW[7] 2.82e-20
C568 a_1757_1642# check[6] 0.318f
C569 D[5] a_6920_627# 0.00234f
C570 x18.X a_14430_90# 0.00259f
C571 a_473_993# VDD_SW_b[7] 3.93e-21
C572 a_941_601# a_1672_909# 0.0016f
C573 x18.X a_12607_601# 1.98e-20
C574 a_9312_627# VSS_SW[3] 0.00166f
C575 VDD_SW_b[4] a_9742_n88# 5.91e-19
C576 x12.X a_7823_601# 2.7e-20
C577 x2.X a_5725_601# 0.119f
C578 a_9646_90# a_9742_n88# 0.0967f
C579 check[3] a_7350_n88# 5.26e-19
C580 a_3839_220# VSS_SW[5] 1.57e-20
C581 a_3421_n88# VSS_SW_b[5] 0.00486f
C582 a_9312_627# m1_95_1942# 2.45e-20
C583 VDD a_13936_1315# 3.62e-19
C584 VDD a_16024_909# 0.00438f
C585 a_1503_1642# a_1415_895# 5.45e-19
C586 x2.X a_10931_627# 0.00111f
C587 VSS_SW[2] a_13407_220# 6.42e-21
C588 check[6] a_487_n62# 1.41e-20
C589 a_12989_n88# VSS_SW_b[2] 7.6e-19
C590 a_13193_n88# a_13461_122# 0.206f
C591 a_16109_1642# VDD_SW_b[1] 1.85e-19
C592 a_3333_601# a_3421_n88# 3.89e-19
C593 a_3807_895# a_3420_212# 0.00165f
C594 a_16109_1642# x20.X 0.0846f
C595 a_2585_627# VSS_SW_b[6] 3.72e-20
C596 a_11987_627# a_12038_90# 6.13e-19
C597 a_939_2457# a_2585_627# 4.92e-21
C598 check[4] a_5504_106# 7.9e-22
C599 VDD_SW_b[3] a_12038_90# 0.00346f
C600 a_10459_909# VDD_SW_b[3] 3.01e-21
C601 x18.X a_14857_1289# 1.51e-19
C602 x2.X VDD_SW[4] 0.0327f
C603 a_4370_1315# D[6] 0.0012f
C604 a_2610_1315# VSS_SW[6] 7.95e-19
C605 VDD a_2949_993# 0.00571f
C606 a_9595_627# a_10680_909# 1.09e-19
C607 VDD a_11704_627# 0.222f
C608 a_720_106# a_2566_n88# 1.86e-21
C609 a_6285_1642# x11.X 1.3e-19
C610 a_11987_627# m1_95_1942# 5.19e-20
C611 x2.X a_6456_909# 3.99e-19
C612 a_5431_601# a_5257_993# 0.206f
C613 VDD_SW_b[3] m1_95_1942# 1.88e-20
C614 a_4977_627# a_5725_601# 0.126f
C615 a_5725_601# VSS_SW[5] 2.18e-19
C616 a_10824_993# m1_95_2154# 4.11e-21
C617 VDD a_720_106# 0.373f
C618 a_8117_601# D[3] 8.74e-19
C619 a_647_601# VSS_SW[7] 6.23e-19
C620 a_8591_895# a_9595_627# 6.9e-19
C621 a_11987_627# a_12541_627# 0.00206f
C622 x9.A1 a_11071_1642# 0.101f
C623 VDD_SW_b[1] VDD_SW[1] 3.65e-19
C624 a_16330_1315# VDD_SW_b[1] 1.33e-20
C625 x20.X a_16330_1315# 0.00143f
C626 x20.X VDD_SW[1] 0.175f
C627 check[2] a_10073_1289# 0.248f
C628 VDD_SW_b[6] a_3420_212# 0.0418f
C629 VDD_SW[5] a_7369_627# 9.25e-19
C630 a_6920_627# a_8117_601# 1.71e-20
C631 a_1503_1642# check[5] 1.16e-20
C632 a_1757_1642# D[7] 0.0607f
C633 a_7254_90# a_8204_212# 1.66e-20
C634 a_14825_993# a_14945_n62# 6.88e-22
C635 a_6730_n62# a_8205_n88# 3.67e-21
C636 a_5950_304# VSS_SW_b[4] 9.89e-21
C637 x9.A1 VSS_SW[7] 0.0981f
C638 a_1501_122# VSS_SW_b[6] 1.09e-20
C639 a_2470_90# VSS_SW[6] 0.082f
C640 a_14379_627# D[1] 0.138f
C641 VDD_SW_b[2] D[1] 1.5e-19
C642 a_5257_993# a_5365_627# 0.00807f
C643 a_6040_993# a_5896_909# 0.00412f
C644 a_5725_601# a_5575_627# 0.00926f
C645 a_5431_601# a_5943_627# 9.75e-19
C646 a_4977_627# a_6456_909# 7.17e-20
C647 a_10596_212# a_11015_220# 2.46e-19
C648 a_10055_n62# a_11514_n62# 3.79e-20
C649 a_10597_n88# a_10734_304# 0.00907f
C650 D[5] a_6730_n62# 0.158f
C651 x8.X a_2865_993# 9.17e-20
C652 a_2897_1289# a_3112_106# 5.3e-21
C653 a_581_627# VSS_SW[7] 3.79e-19
C654 a_9312_627# VDD_SW[4] 0.0729f
C655 x2.X a_15030_220# 0.0028f
C656 a_8731_627# a_8539_627# 4.19e-20
C657 VDD_SW_b[4] a_9595_627# 5.97e-19
C658 a_7681_1289# a_7203_627# 0.00104f
C659 a_9595_627# a_9646_90# 6.13e-19
C660 a_29_2457# check[6] 7.65e-19
C661 a_27_627# a_720_106# 3.88e-21
C662 D[7] a_487_n62# 0.00257f
C663 x2.X a_5271_n62# 0.373f
C664 x9.A1 a_12989_n88# 6.75e-21
C665 x2.X a_10073_1289# 0.0112f
C666 a_13375_895# a_12988_212# 0.00165f
C667 a_12153_627# VSS_SW_b[2] 4.44e-20
C668 a_12901_601# a_12989_n88# 3.89e-19
C669 a_505_1289# VSS_SW[7] 0.00189f
C670 a_11240_909# VDD_SW[3] 2.12e-20
C671 a_5289_1289# a_5431_601# 8.76e-20
C672 VDD a_5761_304# 0.00302f
C673 D[6] a_3648_993# 0.00608f
C674 a_2419_627# a_2773_627# 0.0455f
C675 x14.X a_10041_993# 9.14e-20
C676 a_2468_1467# a_2927_1642# 6.64e-19
C677 a_9595_627# VDD_SW[3] 3.29e-20
C678 x11.X x12.X 0.11f
C679 a_76_1467# m1_95_1942# 1.09e-19
C680 a_1757_1642# m1_95_2154# 8.35e-20
C681 a_941_601# a_3039_601# 1.52e-20
C682 a_1415_895# a_2585_627# 2.96e-19
C683 a_14379_627# a_15380_212# 6.99e-20
C684 D[1] a_15072_106# 8.75e-19
C685 VDD x3.A 0.186f
C686 VDD_SW[2] VSS_SW[1] 0.412f
C687 VDD_SW_b[2] a_15380_212# 4.59e-22
C688 x13.X a_8205_n88# 0.019f
C689 a_3648_993# m1_95_1942# 5.78e-21
C690 a_7252_1467# a_7394_1315# 0.00783f
C691 x9.A1 VSS_SW_b[5] 2.15e-19
C692 a_4977_627# a_5271_n62# 2.38e-19
C693 a_5431_601# a_4958_n88# 4.37e-19
C694 x9.A1 x16.X 8.83e-19
C695 x16.X a_12901_601# 4.99e-20
C696 VSS_SW[5] a_5271_n62# 3.44e-19
C697 a_4338_n62# VSS_SW_b[5] 2.64e-19
C698 D[4] a_10597_n88# 4.83e-22
C699 x9.A1 a_3333_601# 0.00103f
C700 x2.X a_3283_909# 0.00137f
C701 x11.X a_6285_122# 2.61e-19
C702 x2.X a_12988_212# 0.0126f
C703 a_3039_601# a_2985_n62# 1.07e-20
C704 VDD_SW[7] a_2949_993# 6.61e-21
C705 x2.X a_1028_212# 0.0128f
C706 VDD a_3947_627# 0.00233f
C707 VDD_SW_b[7] a_2585_627# 0.00329f
C708 x18.X D[1] 0.00892f
C709 a_10509_601# a_10459_909# 1.21e-20
C710 a_10983_895# a_11514_n62# 4.06e-19
C711 D[3] a_11514_n62# 0.158f
C712 D[3] a_10125_993# 8.11e-19
C713 x9.A1 VDD_SW[5] 0.0926f
C714 VDD a_12447_n62# 0.344f
C715 a_14839_n62# a_15381_n88# 0.125f
C716 a_15072_106# a_15380_212# 0.14f
C717 a_10509_601# VSS_SW[3] 2.13e-19
C718 a_2897_1289# D[6] 0.0661f
C719 check[5] a_2585_627# 5.42e-19
C720 a_1415_895# a_1501_122# 4.53e-22
C721 VDD a_1745_304# 0.00424f
C722 a_1256_993# a_1233_n88# 1.86e-19
C723 VDD a_11069_122# 0.321f
C724 a_8591_895# a_10041_993# 8e-21
C725 a_8623_220# VSS_SW_b[3] 3.75e-21
C726 a_10509_601# m1_95_1942# 4.09e-20
C727 x9.A1 a_13906_n62# 1.56e-20
C728 x9.A1 a_12153_627# 2.37e-19
C729 a_12153_627# a_12901_601# 0.126f
C730 a_12607_601# a_12433_993# 0.206f
C731 x7.X a_1978_1315# 0.00146f
C732 check[1] a_12038_90# 2.5e-20
C733 x9.A1 a_7711_1642# 5.26e-19
C734 check[5] a_3895_1642# 0.257f
C735 a_7203_627# a_8288_909# 1.09e-19
C736 D[4] a_8067_909# 6.77e-19
C737 a_2897_1289# m1_95_1942# 2.26e-19
C738 a_8204_212# a_8205_n88# 0.784f
C739 a_7663_n62# a_8677_122# 0.0633f
C740 a_7896_106# a_8409_n88# 0.00189f
C741 a_7350_n88# VSS_SW_b[4] 0.135f
C742 x10.X a_4811_627# 0.236f
C743 check[4] VDD_SW[6] 4.33e-19
C744 VSS_SW[6] a_3421_n88# 9.29e-21
C745 D[1] a_15799_220# 7.1e-19
C746 check[1] m1_95_1942# 0.034f
C747 a_6040_993# VDD_SW[5] 3.28e-20
C748 D[5] a_8204_212# 7.45e-22
C749 x17.X VSS_SW[1] 0.138f
C750 x13.X a_8117_601# 1.31e-19
C751 VDD_SW_b[7] a_1501_122# 0.00445f
C752 x9.A1 a_15767_895# 2.64e-19
C753 a_5323_2457# VDD_SW[5] 0.0154f
C754 a_13375_895# a_15293_601# 1.42e-20
C755 VDD_SW_b[4] a_10041_993# 8.2e-21
C756 D[7] a_1447_220# 7.11e-19
C757 a_29_2457# m1_95_2154# 1.41e-19
C758 a_4811_627# D[5] 0.137f
C759 x2.X a_5950_304# 0.00334f
C760 a_7369_627# a_9761_627# 2.62e-19
C761 x2.X a_13705_304# 3.38e-19
C762 a_12134_n88# VSS_SW[1] 4.28e-21
C763 a_12680_106# a_13103_n62# 0.00386f
C764 a_12447_n62# a_13329_n62# 0.00926f
C765 a_7203_627# VSS_SW[3] 4.95e-21
C766 D[2] a_12680_106# 8.76e-19
C767 a_11987_627# a_12988_212# 6.99e-20
C768 a_2419_627# a_4528_627# 1.75e-19
C769 x3.X ready 0.127f
C770 VDD_SW_b[1] a_15495_n62# 5.19e-19
C771 D[4] m1_95_2154# 0.0344f
C772 VDD_SW_b[3] a_12988_212# 4.59e-22
C773 a_7203_627# m1_95_1942# 5.19e-20
C774 VDD_SW[3] VSS_SW[2] 0.411f
C775 VSS_SW[4] m1_95_2154# 0.0283f
C776 a_14545_627# a_15143_627# 6.04e-20
C777 a_14857_1289# a_15855_1642# 0.0146f
C778 a_15855_1642# a_15608_993# 0.00176f
C779 a_15293_601# a_15243_909# 1.21e-20
C780 a_10983_895# a_11123_627# 0.0383f
C781 a_10509_601# a_10931_627# 1.96e-20
C782 a_10041_993# VDD_SW[3] 4.17e-21
C783 D[3] a_11123_627# 0.00433f
C784 VDD a_13126_304# 0.0164f
C785 a_15380_212# a_15799_220# 2.46e-19
C786 a_14839_n62# a_16298_n62# 3.79e-20
C787 a_14526_n88# a_14945_n62# 0.0383f
C788 a_15381_n88# a_15518_304# 0.00907f
C789 a_4528_627# m1_95_2154# 1.66e-20
C790 x13.X a_9122_n62# 0.0016f
C791 VDD_SW[4] a_10509_601# 2.55e-20
C792 VDD a_7681_1289# 0.193f
C793 x2.X a_15293_601# 0.119f
C794 a_5812_212# VSS_SW_b[5] 0.00119f
C795 a_5813_n88# a_6285_122# 0.15f
C796 VSS_SW[5] a_5950_304# 1.97e-20
C797 x9.A1 a_9644_1467# 0.197f
C798 a_8933_1642# check[2] 1.62e-19
C799 VSS_SW[7] a_1233_n88# 9.92e-21
C800 VDD a_218_1315# 0.00205f
C801 a_6539_1642# a_6760_1315# 0.00783f
C802 x12.X a_6920_627# 0.0285f
C803 x2.X a_3755_627# 0.00111f
C804 a_8117_601# a_8204_212# 6.03e-19
C805 a_7557_627# a_7350_n88# 3.32e-19
C806 a_8432_993# a_7663_n62# 3.59e-19
C807 VDD a_14999_601# 0.349f
C808 x6.X a_218_1315# 8.34e-19
C809 x16.X a_9595_627# 0.00117f
C810 a_2585_627# a_2865_993# 0.15f
C811 x2.X a_1946_n62# 1.87e-19
C812 a_2566_n88# a_3112_106# 0.207f
C813 a_5725_601# a_7203_627# 3.81e-19
C814 a_10215_601# a_10161_n62# 1.07e-20
C815 a_10596_212# a_12134_n88# 6.15e-19
C816 VDD_SW[5] a_5812_212# 3.18e-19
C817 a_6339_627# a_6017_n88# 7.32e-20
C818 x14.X a_7823_601# 1.98e-20
C819 VDD a_3112_106# 0.369f
C820 a_10596_212# a_10801_n88# 0.15f
C821 VSS_SW[3] a_10246_220# 4.25e-19
C822 a_10055_n62# VSS_SW_b[3] 0.0142f
C823 x2.X a_8933_1642# 5.21e-19
C824 a_4149_1642# a_4528_627# 5.9e-19
C825 a_8205_n88# a_10596_212# 4.01e-22
C826 a_7203_627# VDD_SW[4] 3.29e-20
C827 D[4] a_8539_627# 2e-19
C828 D[2] a_13407_220# 7.11e-19
C829 VDD_SW_b[4] a_7896_106# 5.23e-19
C830 a_8204_212# a_9122_n62# 0.0453f
C831 a_8205_n88# a_8921_304# 0.0018f
C832 a_7663_n62# a_7769_n62# 0.0526f
C833 a_8409_n88# a_8623_220# 0.0104f
C834 x9.A1 VSS_SW[6] 0.102f
C835 a_2865_993# a_3183_627# 0.025f
C836 a_3333_601# a_3732_993# 9.41e-19
C837 a_2585_627# a_3551_627# 2.14e-20
C838 check[6] D[7] 0.445f
C839 a_2773_627# a_2949_993# 8.99e-19
C840 a_14825_993# VDD_SW[1] 4.17e-21
C841 a_15293_601# a_15715_627# 1.96e-20
C842 a_9644_1467# a_9742_n88# 6.87e-20
C843 a_15767_895# a_15907_627# 0.0383f
C844 a_3893_122# VSS_SW_b[6] 7.15e-19
C845 x9.A1 a_9761_627# 2.37e-19
C846 VDD a_6539_1642# 0.137f
C847 a_9595_627# a_12153_627# 1.09e-20
C848 check[3] a_8861_1642# 0.00577f
C849 VDD_SW_b[5] a_5927_n62# 5.21e-19
C850 VDD_SW_b[7] a_964_n62# 8.1e-20
C851 x3.X a_1256_993# 9.79e-21
C852 a_11325_1642# a_12036_1467# 0.00963f
C853 a_14545_627# VSS_SW[1] 0.023f
C854 D[7] a_2879_n62# 3.12e-21
C855 x2.X a_7350_n88# 0.178f
C856 x9.A1 a_14379_627# 7.95e-19
C857 a_4958_n88# a_5462_220# 0.00869f
C858 a_12901_601# a_14379_627# 3.77e-19
C859 a_4860_1467# a_4811_627# 5.32e-19
C860 x9.A1 VDD_SW_b[2] 2.34e-20
C861 x9.A1 a_13461_1642# 0.101f
C862 a_13375_895# a_13632_909# 0.00869f
C863 a_13216_993# a_13119_627# 0.00386f
C864 a_12341_627# a_12541_627# 3.81e-19
C865 a_12901_601# VDD_SW_b[2] 0.00647f
C866 a_13461_1642# a_12901_601# 0.00263f
C867 a_174_n88# a_1028_212# 0.0319f
C868 a_487_n62# a_720_106# 0.124f
C869 check[2] a_12465_1289# 4.15e-21
C870 VDD a_8288_909# 0.0168f
C871 a_3183_627# a_3551_627# 3.34e-19
C872 VDD a_7854_220# 0.00413f
C873 a_3504_909# VDD_SW_b[6] 7.04e-21
C874 ready x27.A 0.00414f
C875 a_7649_993# a_8117_601# 0.0633f
C876 a_7369_627# a_8432_993# 0.0334f
C877 a_8933_1642# a_9312_627# 5.9e-19
C878 x2.X a_10908_993# 4.67e-19
C879 VSS_SW[2] a_12989_n88# 9.3e-21
C880 check[6] m1_95_2154# 0.0352f
C881 check[6] a_535_1642# 0.00526f
C882 a_2419_627# a_2879_n62# 7.27e-19
C883 D[6] a_2566_n88# 0.00507f
C884 a_14379_627# a_14909_993# 4.45e-20
C885 a_15855_1642# D[1] 0.0681f
C886 D[1] a_14733_627# 0.161f
C887 check[0] a_14999_601# 0.00262f
C888 D[3] a_12680_106# 2.77e-21
C889 x2.X a_439_1315# 3.2e-19
C890 VDD x30.A 0.783f
C891 x9.A1 a_8677_122# 8.99e-21
C892 x2.X x7.X 0.00459f
C893 a_10359_627# a_9742_n88# 1.08e-19
C894 a_10824_993# a_11069_122# 1.51e-20
C895 a_5504_106# a_5927_n62# 0.00386f
C896 a_6285_122# a_6730_n62# 0.0369f
C897 a_5271_n62# a_6153_n62# 0.00926f
C898 a_4958_n88# VSS_SW[4] 4.28e-21
C899 D[3] VSS_SW_b[3] 5.32e-19
C900 VDD D[6] 1.09f
C901 ready x8.X 2.31e-20
C902 VDD a_12038_90# 0.203f
C903 VDD a_10459_909# 0.00984f
C904 a_9761_627# a_9742_n88# 4.91e-19
C905 a_14430_90# a_15381_n88# 9.87e-21
C906 a_13407_220# VSS_SW_b[1] 3.96e-21
C907 VDD a_5002_1642# 0.00198f
C908 x2.X a_12465_1289# 0.0112f
C909 x2.X a_13632_909# 4.01e-19
C910 VDD VSS_SW[3] 0.782f
C911 a_4689_2457# a_4811_627# 3.76e-19
C912 check[1] a_12988_212# 1.79e-20
C913 a_8117_601# a_8335_627# 3.73e-19
C914 a_7823_601# VDD_SW_b[4] 2.14e-20
C915 a_8432_993# a_7967_627# 0.00316f
C916 VDD_SW[3] a_13216_993# 1.08e-20
C917 x15.X a_12134_n88# 0.00865f
C918 a_7252_1467# x11.X 4.9e-19
C919 x16.X VSS_SW[2] 0.249f
C920 VDD m1_95_1942# 6.23f
C921 VDD a_1685_1642# 8.63e-19
C922 a_9644_1467# a_9595_627# 5.32e-19
C923 x16.X a_10041_993# 1.56e-20
C924 x2.X a_3420_212# 0.0127f
C925 a_3112_106# a_3369_304# 0.00857f
C926 x15.X a_10801_n88# 1.87e-19
C927 a_2879_n62# a_3558_304# 0.00652f
C928 x9.X VSS_SW_b[5] 0.0173f
C929 VDD a_12541_627# 0.00108f
C930 a_14096_627# m1_95_1942# 2.45e-20
C931 ready a_473_993# 7.59e-22
C932 a_15293_601# a_15853_122# 2.7e-19
C933 a_939_2457# a_941_601# 2.13e-20
C934 a_15855_1642# a_15380_212# 1.39e-21
C935 a_15767_895# a_15585_n88# 4.26e-19
C936 VDD a_3839_220# 0.012f
C937 a_12036_1467# a_12178_1642# 0.00557f
C938 x9.X a_3333_601# 1.27e-19
C939 x3.X VSS_SW[7] 0.0128f
C940 a_13715_1642# VDD_SW_b[2] 2.58e-19
C941 x9.A1 x18.X 8.79e-19
C942 D[7] a_2419_627# 9.98e-20
C943 a_27_627# D[6] 1.19e-20
C944 D[5] a_5341_993# 8.11e-19
C945 x18.X a_12901_601# 0.00129f
C946 a_4811_627# a_5675_909# 2.46e-19
C947 a_13072_909# VDD_SW[2] 2.82e-20
C948 VDD a_1340_993# 0.00284f
C949 x14.X a_9786_1315# 8.2e-19
C950 x2.X a_14839_n62# 0.371f
C951 a_9122_n62# a_10596_212# 2.79e-22
C952 a_8677_122# a_9742_n88# 8e-21
C953 a_8921_304# a_9122_n62# 8.99e-19
C954 a_3807_895# VDD_SW[6] 0.00356f
C955 a_3648_993# a_3755_627# 0.00707f
C956 a_27_627# m1_95_1942# 5.19e-20
C957 D[7] m1_95_2154# 0.0344f
C958 a_3421_n88# a_3761_n62# 6.04e-20
C959 a_3625_n88# a_3535_n62# 9.75e-19
C960 a_13461_122# VSS_SW_b[2] 7.16e-19
C961 a_535_1642# D[7] 5.72e-19
C962 VSS_SW_b[6] a_2985_n62# 0.00335f
C963 a_3420_212# VSS_SW[5] 0.0872f
C964 a_12153_627# VSS_SW[2] 0.0232f
C965 a_14570_1315# D[1] 7.54e-19
C966 D[1] a_16488_627# 0.00233f
C967 VDD a_5725_601# 0.536f
C968 VDD_SW_b[5] VSS_SW_b[4] 0.0325f
C969 x9.A1 check[4] 0.473f
C970 a_9761_627# a_11240_909# 7.17e-20
C971 x9.A1 a_8432_993# 4.84e-21
C972 x2.X a_8516_993# 4.67e-19
C973 a_9595_627# a_10359_627# 0.00134f
C974 x2.X a_8153_304# 0.00166f
C975 a_9595_627# a_9761_627# 0.786f
C976 check[5] a_3893_122# 6.44e-20
C977 ready a_1503_1642# 9.79e-21
C978 a_1028_212# a_1166_304# 1.09e-19
C979 VDD_SW_b[2] a_12553_n62# 4.77e-19
C980 a_2419_627# m1_95_2154# 3.53e-20
C981 a_8117_601# a_9949_627# 2.42e-20
C982 a_27_627# a_1340_993# 2.13e-19
C983 D[7] a_1112_909# 8.51e-19
C984 VDD VDD_SW[4] 0.605f
C985 x8.X a_2136_627# 0.0285f
C986 D[2] a_13119_627# 6.12e-19
C987 x9.A1 a_10103_1642# 5.26e-19
C988 VDD_SW_b[6] VDD_SW[6] 3.64e-19
C989 a_12465_1289# a_11987_627# 0.00104f
C990 x8.X a_1256_993# 2.81e-19
C991 check[2] a_9786_1642# 0.00688f
C992 x12.X a_4811_627# 0.00117f
C993 VDD a_6456_909# 0.00652f
C994 check[4] a_6040_993# 1.76e-19
C995 x2.X a_10161_n62# 5.57e-20
C996 reset a_305_2457# 0.0023f
C997 a_29_2457# x3.A 0.129f
C998 check[0] m1_95_1942# 0.034f
C999 a_6199_895# a_7557_627# 8.26e-21
C1000 a_16488_627# a_15380_212# 6.63e-19
C1001 VDD_SW[7] D[6] 4.48e-19
C1002 a_5323_2457# check[4] 0.0505f
C1003 a_13715_1642# x18.X 7.95e-19
C1004 x2.X a_193_627# 0.0537f
C1005 x10.X a_3039_601# 1.98e-20
C1006 a_1233_n88# VSS_SW[6] 8.81e-20
C1007 a_10596_212# a_11514_n62# 0.0453f
C1008 VSS_SW_b[7] a_1143_n62# 5.24e-19
C1009 a_1501_122# a_1369_n62# 0.025f
C1010 a_10597_n88# a_11313_304# 0.0018f
C1011 a_10801_n88# a_11015_220# 0.0104f
C1012 x2.X a_15518_304# 0.00338f
C1013 D[5] a_6017_n88# 0.00547f
C1014 a_941_601# a_1415_895# 0.265f
C1015 a_193_627# a_557_993# 0.0018f
C1016 a_647_601# a_381_627# 8.07e-20
C1017 VDD_SW[7] m1_95_1942# 0.0331f
C1018 VSS_SW[3] a_10288_106# 4.65e-19
C1019 x30.A a_5431_601# 7.99e-20
C1020 D[2] a_14526_n88# 4.33e-19
C1021 a_939_2457# a_2468_1467# 0.0011f
C1022 a_10288_106# m1_95_1942# 4.96e-22
C1023 a_2468_1467# VSS_SW_b[6] 1.54e-19
C1024 x9.A1 a_13461_122# 2.1e-20
C1025 a_12901_601# a_13461_122# 2.7e-19
C1026 x9.A1 a_1745_n62# 5.7e-21
C1027 a_13375_895# a_13193_n88# 4.26e-19
C1028 x2.X a_4137_304# 3.38e-19
C1029 a_2879_n62# a_4958_n88# 5.13e-21
C1030 VDD_SW[3] D[2] 4.58e-19
C1031 x9.A1 a_1555_627# 5.22e-20
C1032 x18.X a_14791_1315# 2.35e-19
C1033 VDD a_15030_220# 0.00684f
C1034 VDD_SW_b[5] a_7557_627# 9.3e-21
C1035 x17.X a_13715_1315# 2.08e-19
C1036 x9.A1 a_381_627# 4.11e-19
C1037 x2.X a_791_627# 0.0388f
C1038 a_4149_1642# a_4077_1642# 6.64e-19
C1039 x13.X VSS_SW_b[3] 0.0171f
C1040 x14.X D[3] 0.00895f
C1041 VDD a_5271_n62# 0.351f
C1042 a_5431_601# m1_95_1942# 3.42e-20
C1043 a_5257_993# m1_95_2154# 1.86e-20
C1044 a_4149_1642# m1_95_2154# 8.35e-20
C1045 VDD a_10073_1289# 0.191f
C1046 a_791_627# a_1363_627# 2.46e-21
C1047 D[5] a_6339_627# 0.00433f
C1048 D[1] a_15381_n88# 0.158f
C1049 a_14379_627# a_15585_n88# 0.00204f
C1050 a_381_627# a_581_627# 3.81e-19
C1051 a_1415_895# a_1672_909# 0.00869f
C1052 a_1256_993# a_1159_627# 0.00386f
C1053 a_941_601# VDD_SW_b[7] 0.00647f
C1054 a_11325_1642# a_11539_1642# 0.00557f
C1055 x12.X a_7649_993# 1.03e-19
C1056 x2.X a_6199_895# 0.148f
C1057 a_9646_90# a_10055_n62# 4.24e-20
C1058 check[3] a_7663_n62# 1.36e-20
C1059 x14.X a_8933_1315# 1.48e-20
C1060 a_3625_n88# VSS_SW_b[5] 4.55e-20
C1061 a_2985_n62# a_3356_n62# 4.19e-20
C1062 a_4137_304# VSS_SW[5] 6.58e-21
C1063 a_1503_1642# a_1256_993# 0.00176f
C1064 x7.X a_174_n88# 1.64e-21
C1065 x2.X a_13193_n88# 0.00372f
C1066 check[6] a_720_106# 8.67e-22
C1067 ready a_2585_627# 9.49e-21
C1068 a_11514_n62# a_11313_n62# 3.81e-19
C1069 a_3333_601# a_3625_n88# 0.00251f
C1070 a_3648_993# a_3420_212# 8.94e-21
C1071 a_3807_895# a_3421_n88# 6.35e-19
C1072 check[4] a_5812_212# 2.05e-20
C1073 VDD_SW_b[3] a_10161_n62# 4.78e-19
C1074 a_10041_993# a_10359_627# 0.025f
C1075 a_11123_627# a_10596_212# 7.07e-21
C1076 a_9949_627# a_10125_993# 8.99e-19
C1077 a_10509_601# a_10908_993# 9.41e-19
C1078 a_9761_627# VSS_SW[2] 5.1e-21
C1079 x17.X VDD_SW[2] 0.177f
C1080 VDD a_3283_909# 0.0143f
C1081 D[3] a_10680_909# 8.53e-19
C1082 a_1672_909# VDD_SW_b[7] 3.14e-20
C1083 VDD a_12988_212# 0.689f
C1084 a_9761_627# a_10041_993# 0.15f
C1085 ready a_3895_1642# 4.05e-20
C1086 a_1028_212# a_2566_n88# 6.15e-19
C1087 a_14526_n88# VSS_SW_b[1] 0.135f
C1088 a_14839_n62# a_15853_122# 0.0633f
C1089 a_15072_106# a_15585_n88# 0.00189f
C1090 a_15380_212# a_15381_n88# 0.785f
C1091 x2.X VDD_SW_b[5] 7.37e-19
C1092 a_5431_601# a_5725_601# 0.199f
C1093 a_4977_627# a_6199_895# 0.0494f
C1094 a_12036_1467# VSS_SW_b[2] 1.87e-19
C1095 a_10824_993# m1_95_1942# 5.78e-21
C1096 VDD a_1028_212# 0.688f
C1097 a_473_993# VSS_SW[7] 0.00296f
C1098 a_8591_895# D[3] 2.1e-19
C1099 a_8432_993# a_9595_627# 7.56e-20
C1100 x9.A1 a_12433_993# 8.96e-20
C1101 a_14096_627# a_12988_212# 6.63e-19
C1102 a_8204_212# VSS_SW_b[3] 0.00374f
C1103 a_5289_1289# m1_95_2154# 1.04e-19
C1104 a_12153_627# a_13216_993# 0.0334f
C1105 a_12433_993# a_12901_601# 0.0633f
C1106 check[5] a_2927_1642# 0.00526f
C1107 VDD_SW_b[6] a_3421_n88# 0.0406f
C1108 x15.X a_11514_n62# 0.00162f
C1109 VDD_SW[5] a_7823_601# 7.64e-20
C1110 a_8679_1642# x13.X 1.35e-19
C1111 a_7203_627# a_7350_n88# 0.00176f
C1112 a_5812_212# a_7769_n62# 1.09e-19
C1113 a_7254_90# a_8205_n88# 9.87e-21
C1114 a_6231_220# VSS_SW_b[4] 3.96e-21
C1115 D[1] a_16298_n62# 0.158f
C1116 a_964_n62# a_1369_n62# 2.46e-21
C1117 a_4977_627# VDD_SW_b[5] 0.00226f
C1118 x9.A1 a_15855_1642# 0.101f
C1119 a_6040_993# a_6124_993# 0.00857f
C1120 x9.A1 a_14733_627# 4.11e-19
C1121 D[5] a_7254_90# 8.71e-19
C1122 a_13375_895# a_15608_993# 1.86e-21
C1123 a_12901_601# a_14733_627# 2.27e-20
C1124 x8.X a_3333_601# 4.9e-20
C1125 check[1] a_12465_1289# 0.248f
C1126 VDD_SW_b[4] D[3] 1.51e-19
C1127 a_7681_1289# D[4] 0.0662f
C1128 check[3] a_7369_627# 5.38e-19
C1129 x3.A check[6] 9.84e-19
C1130 a_7681_1289# VSS_SW[4] 0.0019f
C1131 a_27_627# a_1028_212# 6.99e-20
C1132 D[7] a_720_106# 8.74e-19
C1133 x2.X a_5504_106# 0.0385f
C1134 x2.X a_14430_90# 0.00368f
C1135 a_3420_212# a_4137_n62# 0.00206f
C1136 x2.X a_12607_601# 0.2f
C1137 a_12988_212# a_13329_n62# 0.00134f
C1138 a_12989_n88# a_13103_n62# 2.14e-20
C1139 a_12680_106# VSS_SW[1] 9.06e-21
C1140 a_1757_1642# D[6] 1.69e-19
C1141 D[2] a_12989_n88# 0.158f
C1142 a_11987_627# a_13193_n88# 0.00204f
C1143 VDD_SW_b[1] a_16097_n62# 5.21e-19
C1144 a_5289_1289# a_5257_993# 4.54e-19
C1145 VDD a_5950_304# 0.0227f
C1146 D[6] a_2773_627# 0.161f
C1147 a_2419_627# a_2949_993# 4.45e-20
C1148 a_14825_993# a_15143_627# 0.025f
C1149 a_14545_627# a_15511_627# 2.14e-20
C1150 a_14733_627# a_14909_993# 8.99e-19
C1151 a_15293_601# a_15692_993# 9.41e-19
C1152 a_10983_895# VDD_SW[3] 0.00356f
C1153 a_10824_993# a_10931_627# 0.00707f
C1154 a_2136_627# a_2585_627# 5.39e-19
C1155 a_2468_1467# check[5] 0.318f
C1156 a_10073_1289# a_10288_106# 5.3e-21
C1157 D[3] VDD_SW[3] 0.235f
C1158 VDD a_13705_304# 0.00422f
C1159 a_1757_1642# a_1685_1642# 6.64e-19
C1160 a_1757_1642# m1_95_1942# 1.97e-19
C1161 a_14839_n62# a_15316_n62# 1.96e-20
C1162 a_15072_106# a_14945_n62# 0.0256f
C1163 a_15585_n88# a_15799_220# 0.0104f
C1164 a_15380_212# a_16298_n62# 0.0453f
C1165 a_941_601# a_2865_993# 1.11e-20
C1166 a_1256_993# a_2585_627# 4.03e-21
C1167 a_15381_n88# a_16097_304# 0.0018f
C1168 VDD_SW[4] a_10824_993# 1.08e-20
C1169 VDD a_7394_1642# 0.00177f
C1170 x2.X a_15608_993# 0.187f
C1171 x2.X a_14857_1289# 0.0112f
C1172 x9.A1 a_12036_1467# 0.197f
C1173 x13.X a_8409_n88# 1.81e-19
C1174 a_14428_1467# a_14430_90# 1e-19
C1175 a_11704_627# m1_95_2154# 1.66e-20
C1176 a_5257_993# a_4958_n88# 8.71e-20
C1177 a_5431_601# a_5271_n62# 0.0026f
C1178 a_11325_1642# check[2] 0.318f
C1179 a_8679_1642# a_8204_212# 1.39e-21
C1180 x17.X a_12134_n88# 1.64e-21
C1181 a_4862_90# VSS_SW_b[5] 0.191f
C1182 VSS_SW[5] a_5504_106# 4.64e-19
C1183 a_193_627# a_174_n88# 4.91e-19
C1184 x16.X D[2] 0.00861f
C1185 x9.A1 a_3807_895# 2.64e-19
C1186 x2.X a_3504_909# 0.0031f
C1187 x13.X x14.X 0.11f
C1188 reset x9.A1 3.51e-20
C1189 VDD a_15293_601# 0.485f
C1190 a_3807_895# a_4338_n62# 4.06e-19
C1191 a_2865_993# a_2985_n62# 6.88e-22
C1192 a_6285_1642# a_6017_n88# 4.63e-19
C1193 VDD_SW[7] a_3283_909# 2.16e-20
C1194 a_10711_n62# a_10937_n62# 3.34e-19
C1195 VDD_SW_b[7] a_3039_601# 1.99e-20
C1196 VDD a_3755_627# 0.00146f
C1197 x2.X a_1029_n88# 0.0213f
C1198 a_16109_1642# a_15767_895# 0.00232f
C1199 a_6539_1642# D[4] 1.68e-19
C1200 x9.A1 a_16488_627# 2e-20
C1201 a_10596_212# a_12680_106# 5.86e-20
C1202 a_1946_n62# a_2566_n88# 8.26e-21
C1203 a_10597_n88# a_12447_n62# 4.56e-21
C1204 VDD_SW[2] a_14545_627# 9.25e-19
C1205 a_14096_627# a_15293_601# 1.84e-20
C1206 x3.A D[7] 1.17e-20
C1207 a_1555_627# a_1233_n88# 7.32e-20
C1208 a_5165_627# VSS_SW_b[5] 3.23e-19
C1209 a_10597_n88# a_11069_122# 0.15f
C1210 a_10596_212# VSS_SW_b[3] 0.00119f
C1211 VSS_SW[3] a_10734_304# 1.97e-20
C1212 check[5] a_3039_601# 0.00264f
C1213 VDD a_1946_n62# 0.109f
C1214 x2.X a_11325_1642# 5.18e-19
C1215 a_791_627# a_174_n88# 1.08e-19
C1216 a_1256_993# a_1501_122# 1.51e-20
C1217 x9.X check[4] 5.57e-19
C1218 x11.X VDD_SW[5] 0.176f
C1219 a_13407_220# VSS_SW[1] 1.77e-20
C1220 a_12989_n88# VSS_SW_b[1] 0.00485f
C1221 a_3807_895# a_6040_993# 1.86e-21
C1222 a_3333_601# a_5165_627# 2.42e-20
C1223 x9.A1 VDD_SW_b[6] 1.63e-20
C1224 a_12433_993# a_12553_n62# 6.88e-22
C1225 a_6285_1642# a_6339_627# 1.92e-20
C1226 VDD_SW_b[6] a_4338_n62# 0.0144f
C1227 D[2] a_13906_n62# 0.158f
C1228 a_11987_627# a_12607_601# 0.149f
C1229 D[2] a_12153_627# 0.168f
C1230 a_7203_627# a_8516_993# 2.13e-19
C1231 D[4] a_8288_909# 8.51e-19
C1232 VDD_SW_b[3] a_12607_601# 2.22e-20
C1233 x9.A1 check[3] 0.402f
C1234 a_15855_1642# a_15907_627# 1.92e-20
C1235 a_15767_895# VDD_SW[1] 0.00356f
C1236 D[4] a_7854_220# 1.98e-20
C1237 a_15608_993# a_15715_627# 0.00707f
C1238 x9.A1 a_2831_1315# 0.00507f
C1239 a_11071_1642# a_10983_895# 5.45e-19
C1240 a_7663_n62# VSS_SW_b[4] 0.0142f
C1241 VDD a_8933_1642# 0.151f
C1242 a_8204_212# a_8409_n88# 0.15f
C1243 VSS_SW[4] a_7854_220# 4.25e-19
C1244 x10.X D[5] 0.00864f
C1245 a_11071_1642# D[3] 0.0682f
C1246 a_5289_1289# a_4958_n88# 5.67e-21
C1247 VSS_SW[6] a_3625_n88# 9.92e-21
C1248 a_16097_304# a_16298_n62# 8.99e-19
C1249 x13.X a_8591_895# 0.00658f
C1250 a_14825_993# VSS_SW[1] 0.00296f
C1251 a_13375_895# D[1] 2.1e-19
C1252 x9.A1 a_12495_1642# 5.26e-19
C1253 a_13216_993# a_14379_627# 7.56e-20
C1254 D[7] a_1745_304# 8.38e-19
C1255 x3.A m1_95_2154# 1.87e-19
C1256 a_29_2457# m1_95_1942# 6.42e-20
C1257 a_13461_1642# a_13216_993# 0.00181f
C1258 x2.X a_6231_220# 9.51e-19
C1259 a_13216_993# VDD_SW_b[2] 4.35e-20
C1260 D[4] VSS_SW[3] 4.86e-19
C1261 VDD a_7350_n88# 0.691f
C1262 D[6] a_4528_627# 0.00235f
C1263 x2.X a_10149_627# 3.99e-19
C1264 a_12447_n62# a_12638_220# 3.3e-19
C1265 VSS_SW[2] a_13461_122# 2.79e-21
C1266 D[4] m1_95_1942# 0.0335f
C1267 VSS_SW[4] m1_95_1942# 0.033f
C1268 VSS_SW_b[3] a_11313_n62# 6.94e-20
C1269 check[0] a_15293_601# 2.14e-19
C1270 a_14887_1642# D[1] 5.74e-19
C1271 a_14379_627# a_15464_909# 1.09e-19
C1272 D[1] a_15243_909# 6.78e-19
C1273 D[3] a_12989_n88# 9.65e-22
C1274 x17.X a_14545_627# 1.68e-19
C1275 x13.X VDD_SW_b[4] 0.242f
C1276 VDD_SW_b[2] a_15464_909# 1.97e-21
C1277 a_9949_627# VSS_SW_b[3] 5.82e-19
C1278 x13.X a_9646_90# 0.0273f
C1279 a_4528_627# m1_95_1942# 2.45e-20
C1280 VDD a_10908_993# 0.00283f
C1281 a_6017_n88# a_6285_122# 0.206f
C1282 a_5813_n88# VSS_SW_b[5] 7.55e-19
C1283 a_13906_n62# VSS_SW_b[1] 2.63e-19
C1284 VSS_SW[5] a_6231_220# 6.42e-21
C1285 x2.X D[1] 0.175f
C1286 x9.A1 a_15381_n88# 8.52e-21
C1287 x8.X VSS_SW[6] 0.253f
C1288 VDD a_6467_1642# 0.00176f
C1289 x7.X a_2566_n88# 0.00862f
C1290 a_78_90# VSS_SW_b[7] 0.19f
C1291 VSS_SW[7] a_1501_122# 2.79e-21
C1292 a_11325_1642# VDD_SW_b[3] 1.69e-19
C1293 VDD a_439_1315# 0.0017f
C1294 x2.X VDD_SW[6] 0.0327f
C1295 check[1] a_13193_n88# 1.52e-20
C1296 a_4413_2457# VDD_SW[6] 0.0115f
C1297 VDD_SW[3] a_12517_993# 6.61e-21
C1298 VDD x7.X 0.461f
C1299 x16.X a_10983_895# 0.00865f
C1300 x6.X a_439_1315# 2.41e-19
C1301 a_8591_895# a_8204_212# 0.00165f
C1302 a_8117_601# a_8205_n88# 3.89e-19
C1303 x16.X D[3] 7.79e-19
C1304 a_7369_627# VSS_SW_b[4] 2.92e-20
C1305 a_3039_601# a_2865_993# 0.206f
C1306 x2.X a_2470_90# 0.00368f
C1307 a_2585_627# a_3333_601# 0.126f
C1308 VDD a_12465_1289# 0.216f
C1309 VDD a_13632_909# 0.00439f
C1310 a_2879_n62# a_3112_106# 0.124f
C1311 a_2566_n88# a_3420_212# 0.0319f
C1312 D[5] a_8117_601# 2.67e-21
C1313 a_5725_601# D[4] 9.63e-19
C1314 a_6199_895# a_7203_627# 6.86e-19
C1315 a_15855_1642# a_15585_n88# 4.63e-19
C1316 a_15143_627# a_14526_n88# 1.08e-19
C1317 a_15608_993# a_15853_122# 1.51e-20
C1318 a_14428_1467# D[1] 0.0177f
C1319 a_9644_1467# a_9786_1315# 0.00783f
C1320 a_6199_895# a_6153_n62# 1.65e-20
C1321 a_5725_601# VSS_SW[4] 2.9e-20
C1322 a_6339_627# a_6285_122# 2.54e-20
C1323 VDD a_3420_212# 0.698f
C1324 x14.X a_7649_993# 1.56e-20
C1325 x18.X a_13216_993# 2.78e-19
C1326 a_3895_1642# a_3333_601# 0.00263f
C1327 VDD_SW[6] a_4977_627# 9.25e-19
C1328 a_4528_627# a_5725_601# 1.71e-20
C1329 x2.X a_15380_212# 0.0122f
C1330 VDD_SW[6] VSS_SW[5] 0.394f
C1331 VDD_SW_b[6] a_5812_212# 2.3e-22
C1332 a_218_1315# D[7] 7.54e-19
C1333 D[4] VDD_SW[4] 0.236f
C1334 VDD_SW_b[4] a_8204_212# 0.0416f
C1335 x7.X a_27_627# 2.67e-20
C1336 a_8409_n88# a_8921_304# 6.69e-20
C1337 a_8205_n88# a_9122_n62# 0.189f
C1338 VSS_SW_b[4] a_8342_304# 3.58e-20
C1339 a_8204_212# a_9646_90# 0.00101f
C1340 a_2865_993# a_2973_627# 0.00807f
C1341 a_3333_601# a_3183_627# 0.00926f
C1342 a_7663_n62# a_8140_n62# 1.96e-20
C1343 a_2585_627# a_4064_909# 7.17e-20
C1344 a_3039_601# a_3551_627# 9.75e-19
C1345 a_7896_106# a_7769_n62# 0.0256f
C1346 a_3648_993# a_3504_909# 0.00412f
C1347 a_305_2457# x2.X 0.00106f
C1348 a_12433_993# VSS_SW[2] 0.003f
C1349 a_16109_1315# D[1] 0.00195f
C1350 a_4860_1467# x10.X 0.0876f
C1351 x9.A1 a_10215_601# 2.81e-20
C1352 a_14379_627# VDD_SW[1] 3.29e-20
C1353 a_1757_1642# a_1028_212# 1.17e-22
C1354 D[1] a_15715_627# 2e-19
C1355 VDD_SW_b[5] a_7203_627# 5.95e-19
C1356 a_6339_627# a_6147_627# 4.19e-20
C1357 a_10983_895# a_12153_627# 2.8e-19
C1358 a_6920_627# VDD_SW[5] 0.0729f
C1359 a_10509_601# a_12607_601# 1.55e-20
C1360 VDD a_14839_n62# 0.357f
C1361 D[3] a_12153_627# 6.4e-21
C1362 VDD_SW_b[5] a_6153_n62# 0.00179f
C1363 a_9595_627# a_10727_627# 0.00272f
C1364 VDD_SW_b[7] a_1143_n62# 5.2e-19
C1365 x9.A1 a_16298_n62# 1.9e-20
C1366 D[7] a_3112_106# 2.77e-21
C1367 x2.X a_7663_n62# 0.373f
C1368 a_4860_1467# D[5] 0.0184f
C1369 VDD_SW_b[2] a_13103_n62# 5.2e-19
C1370 a_5271_n62# a_5462_220# 3.24e-19
C1371 a_7681_1289# m1_95_2154# 1.04e-19
C1372 D[2] a_14379_627# 1e-19
C1373 a_11987_627# D[1] 1.27e-20
C1374 a_13461_1642# D[2] 0.0681f
C1375 check[1] a_12607_601# 0.00262f
C1376 a_487_n62# a_1028_212# 0.138f
C1377 check[6] D[6] 3.68e-20
C1378 a_174_n88# a_1029_n88# 0.0477f
C1379 D[2] VDD_SW_b[2] 0.453f
C1380 VDD a_8516_993# 0.00437f
C1381 x12.X a_7254_90# 0.00259f
C1382 VDD a_8153_304# 0.00272f
C1383 check[2] a_11253_1642# 0.00577f
C1384 a_7369_627# a_7557_627# 0.189f
C1385 a_7823_601# a_8432_993# 0.00189f
C1386 check[6] m1_95_1942# 0.034f
C1387 check[6] a_1685_1642# 0.00577f
C1388 D[6] a_2879_n62# 0.00257f
C1389 a_2419_627# a_3112_106# 3.88e-21
C1390 a_14999_601# m1_95_2154# 2.34e-20
C1391 a_11514_n62# a_12134_n88# 8.26e-21
C1392 x2.X a_1757_1315# 2.32e-19
C1393 a_4689_2457# x10.X 5.56e-19
C1394 check[1] a_14857_1289# 5.99e-21
C1395 x9.A1 VSS_SW_b[4] 2.06e-19
C1396 a_10801_n88# a_11514_n62# 8.07e-20
C1397 a_10597_n88# a_12038_90# 5.39e-19
C1398 VSS_SW_b[3] a_11015_220# 1.12e-20
C1399 a_11069_122# a_11313_304# 0.00972f
C1400 a_5271_n62# VSS_SW[4] 1.46e-20
C1401 a_5812_212# a_5927_n62# 0.00272f
C1402 a_5504_106# a_6153_n62# 0.00316f
C1403 VDD a_10161_n62# 0.0133f
C1404 x2.X a_16097_304# 3.38e-19
C1405 a_10215_601# a_9742_n88# 4.37e-19
C1406 a_9761_627# a_10055_n62# 2.38e-19
C1407 VSS_SW[1] a_14526_n88# 0.00667f
C1408 x10.X a_6285_1642# 2.02e-20
C1409 VSS_SW[3] a_10597_n88# 9.29e-21
C1410 x7.X VDD_SW[7] 0.174f
C1411 a_12036_1467# VSS_SW[2] 0.0274f
C1412 D[2] a_15072_106# 2.77e-21
C1413 VDD a_193_627# 0.728f
C1414 a_8117_601# a_8848_909# 0.0016f
C1415 a_10597_n88# m1_95_1942# 1.16e-21
C1416 check[5] x10.X 5.87e-19
C1417 a_7649_993# VDD_SW_b[4] 5.9e-21
C1418 a_12751_627# a_12134_n88# 1.08e-19
C1419 a_13216_993# a_13461_122# 1.51e-20
C1420 a_11325_1642# a_10509_601# 7.12e-21
C1421 a_7823_601# a_7769_n62# 1.07e-20
C1422 a_9644_1467# D[3] 0.0182f
C1423 x6.X a_193_627# 0.00315f
C1424 x2.X a_3421_n88# 0.0207f
C1425 VDD a_15518_304# 0.023f
C1426 a_2879_n62# a_3839_220# 1.21e-20
C1427 a_3112_106# a_3558_304# 0.00412f
C1428 a_3421_n88# a_3070_220# 4.71e-20
C1429 a_6285_1642# D[5] 0.0682f
C1430 a_3420_212# a_3369_304# 2.13e-19
C1431 x14.X a_9949_627# 6.07e-19
C1432 a_6539_1642# m1_95_2154# 8.35e-20
C1433 VDD a_9786_1642# 0.00265f
C1434 check[5] D[5] 3.88e-20
C1435 VDD a_4137_304# 0.00423f
C1436 a_939_2457# a_1415_895# 0.00134f
C1437 x9.X a_3807_895# 0.00641f
C1438 D[1] a_15853_122# 0.00923f
C1439 a_14379_627# VSS_SW_b[1] 3.11e-20
C1440 check[0] a_14839_n62# 1.32e-20
C1441 x2.X a_7369_627# 0.0537f
C1442 a_11325_1642# check[1] 1.57e-19
C1443 VDD_SW_b[2] VSS_SW_b[1] 0.0325f
C1444 D[7] D[6] 0.00183f
C1445 D[5] a_5675_909# 6.77e-19
C1446 a_4811_627# a_5896_909# 1.09e-19
C1447 a_8933_1642# a_9154_1315# 0.00783f
C1448 x18.X D[2] 0.00106f
C1449 a_6760_1315# VDD_SW_b[5] 1.32e-20
C1450 VDD a_791_627# 0.0105f
C1451 VDD_SW_b[4] a_10596_212# 2.3e-22
C1452 a_9646_90# a_10596_212# 1.66e-20
C1453 a_27_627# a_193_627# 0.786f
C1454 a_3648_993# VDD_SW[6] 3.28e-20
C1455 x2.X VSS_SW_b[2] 0.0278f
C1456 D[7] m1_95_1942# 0.0335f
C1457 a_1685_1642# D[7] 5.72e-19
C1458 a_3625_n88# a_3761_n62# 0.0697f
C1459 VSS_SW_b[6] a_3356_n62# 1.68e-19
C1460 a_3421_n88# VSS_SW[5] 9.22e-19
C1461 VDD a_6199_895# 0.721f
C1462 VDD_SW_b[3] a_10711_n62# 5.21e-19
C1463 a_2419_627# D[6] 0.138f
C1464 a_939_2457# VDD_SW_b[7] 6.41e-21
C1465 a_2585_627# VSS_SW[6] 0.023f
C1466 VDD_SW_b[7] VSS_SW_b[6] 0.0322f
C1467 x9.X VDD_SW_b[6] 0.218f
C1468 check[4] a_4862_90# 2.5e-20
C1469 a_10824_993# a_10908_993# 0.00857f
C1470 x16.X a_12178_1315# 8.32e-19
C1471 x9.A1 a_7557_627# 4.11e-19
C1472 x2.X a_7967_627# 0.0388f
C1473 a_4977_627# a_7369_627# 2.94e-19
C1474 VDD_SW[3] a_10596_212# 2.77e-19
C1475 a_11123_627# a_10801_n88# 7.32e-20
C1476 x2.X a_8342_304# 0.00334f
C1477 VDD a_13193_n88# 0.48f
C1478 a_9761_627# a_10983_895# 0.0494f
C1479 a_15380_212# a_15853_122# 0.159f
C1480 VSS_SW[1] a_15329_304# 8.23e-20
C1481 a_15381_n88# a_15585_n88# 0.117f
C1482 D[3] a_9761_627# 0.168f
C1483 a_15072_106# VSS_SW_b[1] 0.00322f
C1484 a_9595_627# a_10215_601# 0.149f
C1485 x30.A m1_95_2154# 0.00106f
C1486 check[4] x11.X 0.00964f
C1487 a_939_2457# check[5] 0.00134f
C1488 check[5] VSS_SW_b[6] 2.02e-20
C1489 a_4077_1642# D[6] 5.72e-19
C1490 a_487_n62# a_1946_n62# 3.79e-20
C1491 a_1028_212# a_1447_220# 2.46e-19
C1492 a_1029_n88# a_1166_304# 0.00907f
C1493 a_27_627# a_791_627# 0.00134f
C1494 D[7] a_1340_993# 2.53e-19
C1495 a_8591_895# a_9949_627# 8.26e-21
C1496 a_2419_627# m1_95_1942# 5.19e-20
C1497 D[6] m1_95_2154# 0.0343f
C1498 x9.A1 a_13375_895# 2.41e-19
C1499 a_12901_601# a_13375_895# 0.265f
C1500 a_12153_627# a_12517_993# 0.0018f
C1501 a_12607_601# a_12341_627# 8.07e-20
C1502 x9.A1 check[2] 0.41f
C1503 a_7369_627# a_9312_627# 1.79e-20
C1504 a_305_2457# a_76_1467# 1.82e-20
C1505 VSS_SW[3] m1_95_2154# 0.0337f
C1506 x9.A1 a_5223_1315# 0.00507f
C1507 check[5] a_4363_1642# 0.00688f
C1508 x12.X D[5] 7.76e-19
C1509 VDD VDD_SW_b[5] 0.195f
C1510 a_3183_627# VSS_SW[6] 0.0012f
C1511 D[6] a_3558_304# 9.67e-19
C1512 m1_95_2154# m1_95_1942# 0.00289f
C1513 reset x3.X 0.00166f
C1514 x2.X a_647_601# 0.2f
C1515 a_5812_212# VSS_SW_b[4] 0.00378f
C1516 a_5950_304# VSS_SW[4] 2.77e-20
C1517 x10.X a_2865_993# 1.55e-20
C1518 x9.A1 a_14887_1642# 5.26e-19
C1519 a_10288_106# a_10161_n62# 0.0256f
C1520 a_10055_n62# a_10532_n62# 1.96e-20
C1521 a_1501_122# VSS_SW[6] 6.66e-20
C1522 VSS_SW_b[7] a_1369_n62# 5.35e-19
C1523 check[1] D[1] 3.82e-20
C1524 a_193_627# VDD_SW[7] 2.07e-20
C1525 a_941_601# a_2136_627# 5.61e-19
C1526 VDD_SW_b[4] a_9949_627# 9.33e-21
C1527 check[1] a_12178_1642# 0.00688f
C1528 D[5] a_6285_122# 0.00938f
C1529 a_4811_627# VSS_SW_b[5] 8.3e-20
C1530 a_941_601# a_1256_993# 0.13f
C1531 a_473_993# a_381_627# 0.0369f
C1532 a_647_601# a_557_993# 6.69e-20
C1533 a_193_627# a_891_909# 0.00276f
C1534 a_8067_909# VDD_SW[4] 1.01e-20
C1535 a_7394_1642# VSS_SW[4] 0.00105f
C1536 a_4689_2457# a_4860_1467# 0.00106f
C1537 x30.A a_5257_993# 5.04e-19
C1538 x2.X x9.A1 0.626f
C1539 x2.X a_12901_601# 0.119f
C1540 a_12989_n88# VSS_SW[1] 9.23e-19
C1541 a_13193_n88# a_13329_n62# 0.0697f
C1542 VSS_SW_b[2] a_12924_n62# 1.68e-19
C1543 a_4413_2457# x9.A1 1.84e-19
C1544 x2.X a_4338_n62# 1.9e-19
C1545 a_3333_601# a_4811_627# 3.81e-19
C1546 a_4149_1642# D[6] 0.0607f
C1547 D[2] a_13461_122# 0.00928f
C1548 a_11987_627# VSS_SW_b[2] 9.17e-20
C1549 a_3112_106# a_4958_n88# 1.86e-21
C1550 VDD_SW_b[3] VSS_SW_b[2] 0.0324f
C1551 a_15608_993# a_15692_993# 0.00857f
C1552 x20.X a_14545_627# 1.02e-20
C1553 a_14545_627# VDD_SW_b[1] 0.00231f
C1554 x2.X a_581_627# 3.94e-19
C1555 VDD a_5504_106# 0.366f
C1556 a_11071_1642# a_10596_212# 1.39e-21
C1557 VDD a_14430_90# 0.202f
C1558 a_4860_1467# check[5] 1.56e-19
C1559 check[2] a_9742_n88# 5.26e-19
C1560 a_4149_1642# m1_95_1942# 1.97e-19
C1561 a_1757_1642# x7.X 0.0843f
C1562 a_5725_601# m1_95_2154# 2.84e-20
C1563 VDD a_12607_601# 0.326f
C1564 a_5257_993# m1_95_1942# 2.74e-20
C1565 a_15072_106# a_15495_n62# 0.00386f
C1566 a_15853_122# a_16097_304# 0.00972f
C1567 VSS_SW_b[1] a_15799_220# 1.12e-20
C1568 a_14839_n62# a_15721_n62# 0.00926f
C1569 a_15585_n88# a_16298_n62# 8.07e-20
C1570 a_4811_627# VDD_SW[5] 3.29e-20
C1571 D[5] a_6147_627# 2e-19
C1572 VDD a_8861_1642# 0.00181f
C1573 a_1415_895# VDD_SW_b[7] 0.128f
C1574 x2.X a_14909_993# 5.31e-19
C1575 x2.X a_505_1289# 0.0112f
C1576 x9.A1 a_14428_1467# 0.197f
C1577 a_13715_1642# a_13375_895# 0.00226f
C1578 x12.X a_8117_601# 5e-20
C1579 x9.A1 a_4977_627# 2.59e-19
C1580 x17.X a_12680_106# 2.38e-20
C1581 x2.X a_6040_993# 0.187f
C1582 a_9644_1467# x13.X 4.97e-19
C1583 check[3] a_7896_106# 8.41e-22
C1584 a_1503_1642# a_1555_627# 1.92e-20
C1585 x9.A1 VSS_SW[5] 0.116f
C1586 x15.X VDD_SW[3] 0.176f
C1587 VDD_SW[4] m1_95_2154# 0.0327f
C1588 a_3893_122# VSS_SW_b[5] 1.09e-20
C1589 a_4338_n62# VSS_SW[5] 6.06e-20
C1590 a_5323_2457# x2.X 0.00627f
C1591 x7.X a_487_n62# 0.00192f
C1592 a_5002_1315# VSS_SW[5] 7.96e-19
C1593 a_4413_2457# a_5323_2457# 2.64e-19
C1594 check[6] a_1028_212# 3.24e-20
C1595 VDD a_14857_1289# 0.222f
C1596 VDD a_15608_993# 0.197f
C1597 a_3333_601# a_3893_122# 2.7e-19
C1598 a_3807_895# a_3625_n88# 4.26e-19
C1599 ready a_3039_601# 7.34e-21
C1600 check[4] a_5813_n88# 1.15e-20
C1601 a_12134_n88# a_12680_106# 0.207f
C1602 x9.A1 a_9312_627# 2e-20
C1603 a_14428_1467# a_14570_1642# 0.00557f
C1604 x2.X a_9742_n88# 0.178f
C1605 a_8933_1642# D[4] 0.0607f
C1606 x30.A a_5289_1289# 0.00187f
C1607 x9.A1 a_16109_1315# 0.00496f
C1608 a_10596_212# a_12989_n88# 5.48e-21
C1609 a_10597_n88# a_12988_212# 8.02e-22
C1610 VDD_SW[2] a_14825_993# 7.03e-20
C1611 VDD a_3504_909# 0.0248f
C1612 a_1028_212# a_2879_n62# 2.62e-19
C1613 a_10215_601# a_10041_993# 0.206f
C1614 a_1029_n88# a_2566_n88# 1.98e-19
C1615 x16.X a_11325_1315# 2.37e-20
C1616 a_5257_993# a_5725_601# 0.0633f
C1617 a_4977_627# a_6040_993# 0.0334f
C1618 a_10801_n88# VSS_SW_b[3] 9.21e-19
C1619 x2.X a_13715_1642# 5.28e-19
C1620 a_13906_n62# VSS_SW[1] 6.09e-20
C1621 a_13461_122# VSS_SW_b[1] 1.09e-20
C1622 a_941_601# VSS_SW[7] 2.13e-19
C1623 VDD a_1029_n88# 0.661f
C1624 a_5323_2457# a_4977_627# 7.32e-19
C1625 a_12153_627# VSS_SW[1] 5.36e-21
C1626 a_3895_1642# check[4] 6.17e-21
C1627 a_5323_2457# VSS_SW[5] 0.0134f
C1628 a_8205_n88# VSS_SW_b[3] 0.00484f
C1629 a_5289_1289# m1_95_1942# 2.26e-19
C1630 x9.A1 a_11987_627# 7.96e-19
C1631 a_11987_627# a_12901_601# 0.14f
C1632 D[2] a_12433_993# 0.00874f
C1633 x9.A1 VDD_SW_b[3] 1.54e-20
C1634 D[6] a_4958_n88# 4.32e-19
C1635 VDD_SW_b[6] a_3625_n88# 0.00132f
C1636 VDD_SW_b[3] a_12901_601# 5.19e-20
C1637 x27.A a_3807_895# 7.61e-21
C1638 VDD_SW[5] a_7649_993# 7.03e-20
C1639 VDD a_11325_1642# 0.152f
C1640 a_7203_627# a_7663_n62# 7.27e-19
C1641 D[4] a_7350_n88# 0.00506f
C1642 a_10103_1642# D[3] 5.74e-19
C1643 check[2] a_9595_627# 0.0012f
C1644 x13.X a_9761_627# 1.68e-19
C1645 VSS_SW[4] a_7350_n88# 0.00677f
C1646 a_1143_n62# a_1369_n62# 3.34e-19
C1647 a_13715_1642# a_14428_1467# 0.00957f
C1648 x2.X a_14791_1315# 3.2e-19
C1649 x2.X a_15907_627# 0.0151f
C1650 a_6040_993# a_5575_627# 0.00316f
C1651 a_7252_1467# a_7254_90# 1e-19
C1652 a_5431_601# VDD_SW_b[5] 1.75e-20
C1653 a_5725_601# a_5943_627# 3.73e-19
C1654 a_10073_1289# m1_95_2154# 1.04e-19
C1655 check[0] a_14430_90# 2.5e-20
C1656 check[3] a_7823_601# 0.00263f
C1657 D[7] a_1028_212# 0.158f
C1658 a_27_627# a_1029_n88# 1.06e-19
C1659 a_11071_1642# x15.X 1.31e-19
C1660 x2.X a_5812_212# 0.0129f
C1661 x2.X a_12553_n62# 5.25e-20
C1662 a_12447_n62# a_13126_304# 0.00652f
C1663 x2.X a_11240_909# 4.02e-19
C1664 a_12680_106# a_12937_304# 0.00857f
C1665 VDD a_6231_220# 0.0132f
C1666 D[6] a_2949_993# 8.11e-19
C1667 a_16109_1642# a_16488_627# 5.9e-19
C1668 a_2419_627# a_3283_909# 2.46e-19
C1669 x2.X a_4149_1315# 2.33e-19
C1670 a_14379_627# a_15143_627# 0.00134f
C1671 check[0] a_15608_993# 3.41e-19
C1672 a_16323_1642# D[1] 0.00164f
C1673 D[1] a_15692_993# 2.52e-19
C1674 x2.X a_9595_627# 0.355f
C1675 check[0] a_14857_1289# 0.245f
C1676 VDD_SW_b[3] a_9742_n88# 3.21e-19
C1677 a_1415_895# a_2865_993# 8e-21
C1678 a_193_627# a_2773_627# 3.67e-21
C1679 a_941_601# a_3333_601# 9.37e-21
C1680 a_6285_1642# x12.X 1.51e-20
C1681 x13.X a_8677_122# 2.79e-19
C1682 a_11704_627# m1_95_1942# 2.45e-20
C1683 x9.A1 a_15853_122# 3.99e-20
C1684 a_5257_993# a_5271_n62# 2.63e-19
C1685 a_5431_601# a_5504_106# 1.01e-19
C1686 VDD a_2610_1315# 0.0018f
C1687 a_5725_601# a_4958_n88# 0.00259f
C1688 a_4977_627# a_5812_212# 1.02e-19
C1689 a_12036_1467# D[2] 0.0182f
C1690 x9.A1 a_76_1467# 0.197f
C1691 VSS_SW[5] a_5812_212# 5.9e-22
C1692 a_647_601# a_174_n88# 4.37e-19
C1693 a_193_627# a_487_n62# 2.38e-19
C1694 x8.X a_2831_1315# 2.41e-19
C1695 check[1] VSS_SW_b[2] 2.7e-20
C1696 VDD_SW[3] a_13072_909# 2.77e-20
C1697 a_16488_627# VDD_SW[1] 0.0729f
C1698 a_15907_627# a_15715_627# 4.19e-20
C1699 x9.A1 a_3648_993# 4.84e-21
C1700 x2.X a_3732_993# 4.68e-19
C1701 a_720_106# m1_95_1942# 4.96e-22
C1702 x20.X VDD_SW_b[1] 0.243f
C1703 a_4528_627# a_3420_212# 6.63e-19
C1704 a_6285_1642# a_6285_122# 1.57e-21
C1705 VDD D[1] 0.9f
C1706 a_7203_627# a_7369_627# 0.786f
C1707 VDD_SW[7] a_3504_909# 2.77e-20
C1708 VDD a_12178_1642# 0.00346f
C1709 VDD VDD_SW[6] 0.471f
C1710 x9.A1 a_174_n88# 7.34e-19
C1711 VDD_SW_b[7] a_2865_993# 8.2e-21
C1712 x2.X a_1233_n88# 0.00369f
C1713 a_14733_627# VSS_SW_b[1] 7.36e-20
C1714 a_1501_122# a_1745_n62# 0.00807f
C1715 a_2470_90# a_2566_n88# 0.0967f
C1716 a_13715_1642# a_13929_1642# 0.00557f
C1717 a_13515_627# a_14379_627# 1.09e-19
C1718 a_14096_627# D[1] 4.27e-19
C1719 a_1555_627# a_1501_122# 2.54e-20
C1720 a_13461_1642# a_13515_627# 1.92e-20
C1721 check[5] a_2865_993# 7.19e-20
C1722 a_9312_627# a_9595_627# 0.00111f
C1723 VDD a_2470_90# 0.199f
C1724 x15.X x16.X 0.11f
C1725 x2.X a_15585_n88# 0.00368f
C1726 a_9122_n62# VSS_SW_b[3] 2.62e-19
C1727 a_12553_n62# a_12924_n62# 4.19e-20
C1728 a_3807_895# a_5165_627# 8.26e-21
C1729 VDD_SW_b[6] a_4862_90# 0.00345f
C1730 a_7203_627# a_7967_627# 0.00134f
C1731 D[4] a_8516_993# 2.53e-19
C1732 a_505_1289# a_174_n88# 5.67e-21
C1733 check[2] VSS_SW[2] 1.44e-19
C1734 x9.A1 a_10509_601# 0.00103f
C1735 a_7896_106# VSS_SW_b[4] 0.00322f
C1736 a_8205_n88# a_8409_n88# 0.117f
C1737 VSS_SW[4] a_8153_304# 8.35e-20
C1738 a_8204_212# a_8677_122# 0.159f
C1739 a_11240_909# VDD_SW_b[3] 3.4e-20
C1740 a_10509_601# a_12901_601# 9.37e-21
C1741 a_10983_895# a_12433_993# 8e-21
C1742 a_5289_1289# a_5271_n62# 3.44e-19
C1743 VDD a_15380_212# 0.692f
C1744 VSS_SW[6] a_3893_122# 2.79e-21
C1745 check[2] a_10041_993# 6.72e-20
C1746 a_9595_627# a_11987_627# 1.63e-20
C1747 a_9595_627# VDD_SW_b[3] 1.12e-19
C1748 x11.X check[3] 5.57e-19
C1749 x9.A1 a_2897_1289# 0.104f
C1750 VDD a_305_2457# 0.405f
C1751 a_14379_627# VSS_SW[1] 0.0564f
C1752 a_7252_1467# D[5] 2.96e-19
C1753 VDD_SW_b[2] VSS_SW[1] 0.00248f
C1754 a_8679_1642# a_8117_601# 0.00263f
C1755 D[7] a_1946_n62# 0.158f
C1756 x3.A m1_95_1942# 8.75e-20
C1757 x2.X a_6529_304# 3.34e-19
C1758 VDD_SW_b[6] a_5165_627# 9.33e-21
C1759 x9.A1 a_4137_n62# 5.7e-21
C1760 x9.A1 check[1] 0.409f
C1761 check[1] a_12901_601# 1.67e-19
C1762 a_12495_1642# D[2] 5.74e-19
C1763 a_4958_n88# a_5271_n62# 0.245f
C1764 a_4338_n62# a_4137_n62# 3.81e-19
C1765 x9.A1 a_7615_1315# 0.00507f
C1766 x15.X a_12153_627# 1.68e-19
C1767 D[6] a_3947_627# 0.00431f
C1768 VDD a_7663_n62# 0.338f
C1769 x2.X VSS_SW[2] 0.0778f
C1770 a_15907_627# a_15853_122# 2.54e-20
C1771 a_15293_601# m1_95_2154# 2.82e-20
C1772 check[6] x7.X 0.00967f
C1773 x2.X a_10041_993# 0.15f
C1774 a_12038_90# a_12447_n62# 4.24e-20
C1775 x2.X x9.X 0.00459f
C1776 check[0] D[1] 0.461f
C1777 a_14545_627# a_14825_993# 0.15f
C1778 a_4413_2457# x9.X 4.53e-20
C1779 x9.A1 a_7203_627# 7.89e-19
C1780 a_305_2457# a_27_627# 1.18e-19
C1781 VDD a_10711_n62# 0.00521f
C1782 a_9761_627# a_10596_212# 1.02e-19
C1783 x2.X a_14945_n62# 5.25e-20
C1784 a_10509_601# a_9742_n88# 0.00259f
C1785 a_6017_n88# VSS_SW_b[5] 9.2e-19
C1786 VSS_SW[3] a_11069_122# 2.79e-21
C1787 VSS_SW[1] a_15072_106# 4.61e-19
C1788 x7.X a_2879_n62# 4.41e-20
C1789 VSS_SW[7] VSS_SW_b[7] 0.0072f
C1790 D[2] a_15381_n88# 9.66e-22
C1791 a_12341_627# VSS_SW_b[2] 4.17e-19
C1792 x8.X a_1978_1315# 3.75e-20
C1793 a_12036_1467# D[3] 2.97e-19
C1794 VDD a_16097_304# 0.0042f
C1795 a_8591_895# a_8205_n88# 6.35e-19
C1796 a_8117_601# a_8409_n88# 0.00251f
C1797 a_8432_993# a_8204_212# 8.94e-21
C1798 a_5319_1642# D[5] 5.74e-19
C1799 a_2585_627# a_3807_895# 0.0494f
C1800 a_3039_601# a_3333_601# 0.199f
C1801 x2.X a_593_n62# 5.57e-20
C1802 check[4] a_4811_627# 0.0012f
C1803 x9.X a_4977_627# 1.69e-19
C1804 a_2566_n88# a_3421_n88# 0.0477f
C1805 a_2879_n62# a_3420_212# 0.138f
C1806 x9.X VSS_SW[5] 0.138f
C1807 a_8933_1642# m1_95_2154# 8.35e-20
C1808 a_6199_895# D[4] 2.17e-19
C1809 a_6040_993# a_7203_627# 7.46e-20
C1810 VDD a_11253_1642# 9.05e-19
C1811 check[0] a_15380_212# 3.24e-20
C1812 a_6199_895# VSS_SW[4] 7.03e-21
C1813 x17.X a_14526_n88# 0.00864f
C1814 x18.X VSS_SW[1] 0.248f
C1815 a_13715_1642# check[1] 0.318f
C1816 VDD a_3421_n88# 0.684f
C1817 a_1415_895# a_1369_n62# 1.65e-20
C1818 a_941_601# VSS_SW[6] 2.81e-20
C1819 x14.X a_8117_601# 0.0013f
C1820 a_3895_1642# a_3807_895# 5.45e-19
C1821 VDD_SW[6] a_5431_601# 7.64e-20
C1822 VDD_SW_b[6] a_5813_n88# 2.44e-21
C1823 a_439_1315# D[7] 0.00202f
C1824 VDD_SW_b[4] a_8205_n88# 0.0406f
C1825 VDD a_7369_627# 0.667f
C1826 x7.X D[7] 0.0855f
C1827 a_8409_n88# a_9122_n62# 8.07e-20
C1828 a_8205_n88# a_9646_90# 5.39e-19
C1829 a_8677_122# a_8921_304# 0.00972f
C1830 a_7896_106# a_8140_n62# 0.00707f
C1831 a_7663_n62# a_8319_n62# 3.73e-19
C1832 VSS_SW_b[4] a_8623_220# 1.12e-20
C1833 a_3648_993# a_3732_993# 0.00857f
C1834 x3.X x2.X 0.00477f
C1835 a_2585_627# VDD_SW_b[6] 0.00226f
C1836 a_939_2457# ready 0.262f
C1837 a_11987_627# VSS_SW[2] 0.0579f
C1838 VDD_SW_b[3] VSS_SW[2] 0.00249f
C1839 VDD_SW_b[5] D[4] 1.57e-19
C1840 VDD_SW_b[5] VSS_SW[4] 0.00249f
C1841 a_10041_993# VDD_SW_b[3] 4.92e-21
C1842 a_10509_601# a_11240_909# 0.0016f
C1843 D[3] a_10727_627# 6.13e-19
C1844 VDD_SW_b[7] a_1369_n62# 0.00179f
C1845 VDD VSS_SW_b[2] 0.126f
C1846 a_9761_627# a_9949_627# 0.189f
C1847 check[3] D[3] 3.87e-20
C1848 a_15585_n88# a_15853_122# 0.206f
C1849 VSS_SW[1] a_15799_220# 6.42e-21
C1850 a_15381_n88# VSS_SW_b[1] 7.59e-19
C1851 D[7] a_3420_212# 5.78e-20
C1852 a_9595_627# a_10509_601# 0.14f
C1853 x2.X a_7896_106# 0.0385f
C1854 x9.X a_4370_1315# 0.00145f
C1855 x7.X a_2419_627# 0.00295f
C1856 a_7681_1289# m1_95_1942# 2.26e-19
C1857 a_487_n62# a_1029_n88# 0.125f
C1858 a_720_106# a_1028_212# 0.14f
C1859 a_13515_627# a_13461_122# 2.54e-20
C1860 x9.A1 a_12341_627# 4.11e-19
C1861 a_13375_895# a_13216_993# 0.207f
C1862 a_12153_627# a_13072_909# 0.00907f
C1863 a_12607_601# a_12851_909# 0.0104f
C1864 a_12901_601# a_12341_627# 1.15e-20
C1865 VDD a_7967_627# 2.35e-19
C1866 a_12433_993# a_12517_993# 0.00972f
C1867 VDD a_8342_304# 0.018f
C1868 a_8117_601# a_8591_895# 0.265f
C1869 a_7823_601# a_7557_627# 8.07e-20
C1870 a_7369_627# a_7733_993# 0.0018f
C1871 check[6] a_193_627# 5.41e-19
C1872 x15.X a_9761_627# 1.08e-20
C1873 x7.X m1_95_2154# 1.31e-20
C1874 a_14999_601# m1_95_1942# 3.42e-20
C1875 a_2419_627# a_3420_212# 6.99e-20
C1876 D[6] a_3112_106# 8.76e-19
C1877 a_12465_1289# m1_95_2154# 1.04e-19
C1878 a_10055_n62# a_10937_n62# 0.00926f
C1879 a_10288_106# a_10711_n62# 0.00386f
C1880 a_5812_212# a_6153_n62# 0.00134f
C1881 a_5504_106# VSS_SW[4] 9.06e-21
C1882 a_5813_n88# a_5927_n62# 2.14e-20
C1883 check[1] a_13643_1642# 0.00577f
C1884 a_10215_601# a_10055_n62# 0.0026f
C1885 a_9742_n88# a_10246_220# 0.00869f
C1886 a_8861_1642# D[4] 5.72e-19
C1887 a_3112_106# m1_95_1942# 4.96e-22
C1888 x11.X VSS_SW_b[4] 0.017f
C1889 VDD a_647_601# 0.345f
C1890 a_13461_122# VSS_SW[1] 6.77e-20
C1891 VSS_SW_b[2] a_13329_n62# 5.34e-19
C1892 a_7203_627# a_9595_627# 1.74e-20
C1893 x2.X a_13216_993# 0.187f
C1894 a_8591_895# a_8848_909# 0.00869f
C1895 a_7557_627# a_7757_627# 3.81e-19
C1896 a_8117_601# VDD_SW_b[4] 0.00623f
C1897 a_8432_993# a_8335_627# 0.00386f
C1898 a_7649_993# a_7769_n62# 6.88e-22
C1899 a_8591_895# a_9122_n62# 4.06e-19
C1900 a_2468_1467# VSS_SW[6] 0.0274f
C1901 x2.X a_6539_1315# 2.34e-19
C1902 x6.X a_647_601# 2.4e-20
C1903 x9.A1 a_2566_n88# 7.35e-19
C1904 x2.X a_3625_n88# 0.00371f
C1905 a_4860_1467# a_5319_1642# 6.64e-19
C1906 a_3420_212# a_3558_304# 1.09e-19
C1907 a_15293_601# a_16024_909# 0.0016f
C1908 a_14825_993# VDD_SW_b[1] 5.89e-21
C1909 a_939_2457# a_2136_627# 6.01e-19
C1910 a_11071_1642# a_10801_n88# 4.63e-19
C1911 a_6539_1642# m1_95_1942# 1.97e-19
C1912 VDD x9.A1 5.78f
C1913 x12.X a_8679_1642# 1.98e-20
C1914 a_15381_n88# a_15495_n62# 2.14e-20
C1915 VDD a_12901_601# 0.462f
C1916 a_15380_212# a_15721_n62# 0.00134f
C1917 a_939_2457# a_1256_993# 4.83e-21
C1918 ready a_1415_895# 3.23e-21
C1919 VDD a_4338_n62# 0.109f
C1920 VDD a_5002_1315# 6.18e-19
C1921 a_14545_627# a_14526_n88# 4.91e-19
C1922 x2.X a_7823_601# 0.2f
C1923 x2.X a_15464_909# 0.00309f
C1924 x9.A1 x6.X 6.9e-19
C1925 a_4811_627# a_6124_993# 2.13e-19
C1926 D[5] a_5896_909# 8.45e-19
C1927 VDD a_581_627# 9.97e-19
C1928 x9.A1 a_14096_627# 2e-20
C1929 a_12153_627# VDD_SW[2] 2.07e-20
C1930 a_12901_601# a_14096_627# 5.61e-19
C1931 x17.X a_12989_n88# 0.019f
C1932 a_8848_909# VDD_SW_b[4] 3.66e-20
C1933 D[7] a_193_627# 0.168f
C1934 a_27_627# a_647_601# 0.149f
C1935 VDD_SW_b[4] a_9122_n62# 0.0144f
C1936 a_4149_1642# a_3420_212# 1.17e-22
C1937 VSS_SW_b[6] a_3535_n62# 5.24e-19
C1938 a_3893_122# a_3761_n62# 0.025f
C1939 a_3625_n88# VSS_SW[5] 8.78e-20
C1940 x27.A x2.X 2.91e-19
C1941 VDD a_14909_993# 0.00586f
C1942 VDD a_14570_1642# 0.00332f
C1943 a_4413_2457# x27.A 0.129f
C1944 ready a_4689_2457# 0.00228f
C1945 VDD a_505_1289# 0.222f
C1946 a_12134_n88# a_12989_n88# 0.0477f
C1947 a_12447_n62# a_12988_212# 0.138f
C1948 VDD a_6040_993# 0.225f
C1949 a_3039_601# VSS_SW[6] 6.25e-19
C1950 ready VDD_SW_b[7] 5.69e-21
C1951 a_12036_1467# a_12178_1315# 0.00783f
C1952 x6.X a_505_1289# 1.51e-19
C1953 a_10983_895# a_10937_n62# 1.65e-20
C1954 x9.A1 a_27_627# 7.67e-19
C1955 a_10509_601# VSS_SW[2] 2.89e-20
C1956 x2.X a_7757_627# 3.94e-19
C1957 VDD_SW[2] a_15767_895# 1.27e-20
C1958 VDD a_5323_2457# 1.55f
C1959 x2.X a_8623_220# 9.43e-19
C1960 a_10041_993# a_10509_601# 0.0633f
C1961 x2.X x8.X 5.54e-19
C1962 D[3] a_10215_601# 0.00583f
C1963 x30.A m1_95_1942# 4.93e-19
C1964 a_193_627# a_2419_627# 1.58e-20
C1965 ready check[5] 0.0417f
C1966 a_6539_1642# a_5725_601# 7.56e-21
C1967 a_174_n88# a_593_n62# 0.0383f
C1968 a_487_n62# a_2470_90# 6.12e-21
C1969 a_1029_n88# a_1447_220# 0.00276f
C1970 a_1233_n88# a_1166_304# 9.46e-19
C1971 VSS_SW_b[7] a_678_220# 5.34e-20
C1972 a_1028_212# a_1745_304# 4.45e-20
C1973 x2.X a_16109_1642# 5.24e-19
C1974 D[6] m1_95_1942# 0.0335f
C1975 a_27_627# a_581_627# 0.00206f
C1976 VDD a_9742_n88# 0.692f
C1977 a_2897_1289# x9.X 1.75e-20
C1978 a_11987_627# a_13216_993# 0.14f
C1979 D[2] a_13375_895# 0.0294f
C1980 check[1] VSS_SW[2] 0.0496f
C1981 VSS_SW[3] m1_95_1942# 0.0329f
C1982 x27.A VSS_SW[5] 6.7e-19
C1983 a_193_627# m1_95_2154# 2.61e-20
C1984 a_7252_1467# x12.X 0.0876f
C1985 check[2] D[2] 3.87e-20
C1986 a_15243_909# VDD_SW[1] 1.01e-20
C1987 a_505_1289# a_27_627# 0.00104f
C1988 a_2973_627# VSS_SW[6] 3.79e-19
C1989 D[6] a_3839_220# 7.11e-19
C1990 VDD a_13715_1642# 0.115f
C1991 a_9595_627# a_12341_627# 4.46e-21
C1992 check[3] x13.X 0.00968f
C1993 a_11539_1642# D[3] 0.00162f
C1994 a_14945_n62# a_15316_n62# 4.19e-20
C1995 x2.X a_473_993# 0.15f
C1996 a_6231_220# VSS_SW[4] 1.57e-20
C1997 a_5813_n88# VSS_SW_b[4] 0.00486f
C1998 x2.X VDD_SW[1] 0.0322f
C1999 x10.X a_3333_601# 0.00124f
C2000 a_14733_627# VSS_SW[1] 0.00595f
C2001 a_939_2457# VSS_SW[7] 0.00403f
C2002 a_13715_1642# a_14096_627# 5.84e-19
C2003 x9.A1 a_218_1642# 8.64e-19
C2004 a_941_601# a_1555_627# 0.0526f
C2005 a_1415_895# a_2136_627# 0.0967f
C2006 x9.A1 check[0] 0.407f
C2007 a_647_601# VDD_SW[7] 2.07e-20
C2008 x17.X a_13906_n62# 0.0016f
C2009 x9.A1 a_10007_1315# 0.00504f
C2010 x17.X a_12153_627# 1.13e-20
C2011 a_12751_627# a_13119_627# 3.34e-19
C2012 a_13072_909# VDD_SW_b[2] 4.69e-21
C2013 D[5] VSS_SW_b[5] 5.31e-19
C2014 a_1415_895# a_1256_993# 0.207f
C2015 a_473_993# a_557_993# 0.00972f
C2016 a_647_601# a_891_909# 0.0104f
C2017 a_193_627# a_1112_909# 0.00907f
C2018 a_941_601# a_381_627# 1.24e-20
C2019 a_8288_909# VDD_SW[4] 2.82e-20
C2020 x30.A a_5725_601# 2.1e-19
C2021 VDD a_15907_627# 6.88e-19
C2022 VDD a_14791_1315# 0.00121f
C2023 a_3333_601# D[5] 9.63e-19
C2024 D[6] a_5725_601# 2.67e-21
C2025 a_3807_895# a_4811_627# 6.86e-19
C2026 x2.X a_4862_90# 0.00369f
C2027 x2.X D[2] 0.18f
C2028 a_3420_212# a_4958_n88# 6.15e-19
C2029 a_12988_212# a_13126_304# 1.09e-19
C2030 a_12153_627# a_12134_n88# 4.91e-19
C2031 x9.A1 VDD_SW[7] 0.0329f
C2032 VDD_SW_b[5] a_8067_909# 2.62e-21
C2033 VDD_SW_b[5] a_6529_n62# 5.22e-19
C2034 x2.X x11.X 0.00457f
C2035 x2.X a_1159_627# 0.00702f
C2036 a_14379_627# a_15511_627# 0.00272f
C2037 check[0] a_14570_1642# 0.00688f
C2038 VDD a_5812_212# 0.709f
C2039 VDD a_12553_n62# 0.0152f
C2040 a_5725_601# m1_95_1942# 4.12e-20
C2041 a_6199_895# m1_95_2154# 5.86e-20
C2042 check[2] a_10055_n62# 1.35e-20
C2043 VDD_SW_b[7] a_2136_627# 0.185f
C2044 D[5] VDD_SW[5] 0.226f
C2045 VDD_SW[4] a_10459_909# 2.16e-20
C2046 VDD a_11240_909# 0.0044f
C2047 a_1256_993# VDD_SW_b[7] 4.35e-20
C2048 x2.X a_1503_1642# 0.00652f
C2049 VDD_SW[4] VSS_SW[3] 0.412f
C2050 a_14428_1467# D[2] 2.85e-19
C2051 x2.X a_5165_627# 0.0014f
C2052 VDD a_9595_627# 0.411f
C2053 x9.A1 a_5431_601# 3.62e-20
C2054 check[3] a_8204_212# 1.76e-20
C2055 VDD_SW_b[6] a_4811_627# 5.96e-19
C2056 a_4528_627# VDD_SW[6] 0.0729f
C2057 a_3947_627# a_3755_627# 4.19e-20
C2058 VDD_SW[4] m1_95_1942# 0.0331f
C2059 a_4862_90# VSS_SW[5] 0.082f
C2060 x7.X a_720_106# 2.38e-20
C2061 check[6] a_1029_n88# 2.51e-20
C2062 x11.X a_4977_627# 1.08e-20
C2063 a_3648_993# a_3625_n88# 1.86e-19
C2064 a_3807_895# a_3893_122# 4.53e-22
C2065 ready a_2865_993# 5.7e-21
C2066 VDD a_13643_1642# 8.63e-19
C2067 check[4] a_6017_n88# 6e-20
C2068 VDD_SW_b[5] m1_95_2154# 1.95e-20
C2069 a_29_2457# a_305_2457# 0.00202f
C2070 x9.A1 a_8731_627# 1.09e-20
C2071 x2.X a_10055_n62# 0.373f
C2072 VDD_SW_b[1] a_14526_n88# 3.21e-19
C2073 x20.X a_14526_n88# 1.53e-21
C2074 a_14570_1315# VSS_SW[1] 7.95e-19
C2075 a_13715_1642# check[0] 1.46e-19
C2076 VDD a_3732_993# 0.0044f
C2077 a_11325_1642# a_11546_1315# 0.00783f
C2078 VDD_SW[2] a_14379_627# 0.0865f
C2079 a_1029_n88# a_2879_n62# 4.56e-21
C2080 a_1745_304# a_1946_n62# 8.99e-19
C2081 a_1028_212# a_3112_106# 5.86e-20
C2082 VDD_SW_b[2] VDD_SW[2] 3.64e-19
C2083 a_5431_601# a_6040_993# 0.00189f
C2084 a_4977_627# a_5165_627# 0.189f
C2085 a_5165_627# VSS_SW[5] 0.00596f
C2086 a_9742_n88# a_10288_106# 0.207f
C2087 x2.X VSS_SW_b[1] 0.0278f
C2088 VDD a_1233_n88# 0.48f
C2089 a_5323_2457# a_5431_601# 4.92e-19
C2090 a_8409_n88# VSS_SW_b[3] 4.04e-20
C2091 check[4] a_6339_627# 1.61e-19
C2092 VDD_SW_b[6] a_3893_122# 0.00445f
C2093 D[6] a_5271_n62# 1.56e-21
C2094 a_11987_627# D[2] 0.137f
C2095 a_12341_627# VSS_SW[2] 0.00596f
C2096 VDD_SW_b[3] D[2] 1.57e-19
C2097 x9.A1 a_10824_993# 4.84e-21
C2098 check[0] a_15907_627# 4.05e-19
C2099 VDD_SW[5] a_8117_601# 2.46e-20
C2100 D[4] a_7663_n62# 0.00257f
C2101 VDD a_15585_n88# 0.483f
C2102 a_7203_627# a_7896_106# 3.88e-21
C2103 x18.X a_13715_1315# 1.47e-20
C2104 check[2] a_10983_895# 0.00235f
C2105 a_6730_n62# VSS_SW_b[4] 2.78e-19
C2106 VSS_SW[4] a_7663_n62# 3.44e-19
C2107 check[2] D[3] 0.463f
C2108 a_10073_1289# VSS_SW[3] 0.00187f
C2109 x9.A1 a_2610_1642# 8.62e-19
C2110 a_14428_1467# VSS_SW_b[1] 7.31e-20
C2111 a_5257_993# VDD_SW_b[5] 4.92e-21
C2112 a_5725_601# a_6456_909# 0.0016f
C2113 a_10073_1289# m1_95_1942# 2.26e-19
C2114 a_12607_601# m1_95_2154# 2.34e-20
C2115 a_4860_1467# VSS_SW_b[5] 1.56e-19
C2116 a_12153_627# a_14545_627# 3.26e-19
C2117 check[3] a_7649_993# 6.94e-20
C2118 a_13929_1642# D[2] 0.00166f
C2119 check[1] a_13216_993# 1.83e-19
C2120 D[7] a_1029_n88# 0.158f
C2121 a_27_627# a_1233_n88# 0.00204f
C2122 x2.X a_5813_n88# 0.0213f
C2123 x2.X a_2585_627# 0.0537f
C2124 a_2419_627# a_3504_909# 1.09e-19
C2125 D[6] a_3283_909# 6.77e-19
C2126 VDD a_6529_304# 0.00566f
C2127 x2.X a_10983_895# 0.148f
C2128 a_15608_993# m1_95_2154# 4.11e-21
C2129 a_14857_1289# m1_95_2154# 1.04e-19
C2130 a_10734_304# VSS_SW_b[2] 1.09e-20
C2131 a_12038_90# a_12988_212# 2.02e-20
C2132 a_11514_n62# a_12989_n88# 3.67e-21
C2133 x2.X D[3] 0.177f
C2134 a_14545_627# a_15767_895# 0.0494f
C2135 a_14999_601# a_15293_601# 0.199f
C2136 x17.X a_14379_627# 0.00295f
C2137 x18.X VDD_SW[2] 0.305f
C2138 a_1415_895# a_3333_601# 1.42e-20
C2139 VDD_SW_b[3] a_10055_n62# 5.23e-19
C2140 x17.X VDD_SW_b[2] 0.22f
C2141 x2.X a_3895_1642# 0.00651f
C2142 a_13461_1642# x17.X 1.37e-19
C2143 x9.X a_2566_n88# 1.49e-21
C2144 VDD VSS_SW[2] 0.944f
C2145 a_9761_627# a_10801_n88# 8.75e-19
C2146 VSS_SW[1] a_15381_n88# 9.29e-21
C2147 a_12988_212# m1_95_1942# 6.77e-21
C2148 x2.X a_6920_627# 3.85e-19
C2149 a_9595_627# a_10288_106# 3.88e-21
C2150 VDD a_10041_993# 0.18f
C2151 a_4977_627# a_5813_n88# 1.27e-19
C2152 a_5431_601# a_5812_212# 4.51e-19
C2153 a_5257_993# a_5504_106# 4.96e-20
C2154 a_5725_601# a_5271_n62# 3.74e-20
C2155 a_8679_1642# a_8409_n88# 4.63e-19
C2156 x9.A1 a_1757_1642# 0.195f
C2157 VSS_SW[5] a_5813_n88# 9.3e-21
C2158 a_473_993# a_174_n88# 8.71e-20
C2159 a_647_601# a_487_n62# 0.0026f
C2160 VDD x9.X 0.46f
C2161 x2.X a_8933_1315# 2.32e-19
C2162 a_8204_212# a_8921_n62# 0.00206f
C2163 a_78_90# VSS_SW[7] 0.082f
C2164 VDD_SW_b[2] a_12134_n88# 3.21e-19
C2165 a_12465_1289# a_12447_n62# 3.44e-19
C2166 a_1028_212# m1_95_1942# 6.77e-21
C2167 a_2585_627# a_4977_627# 2.94e-19
C2168 x2.X a_3183_627# 0.0388f
C2169 x9.A1 a_2773_627# 4.11e-19
C2170 a_2585_627# VSS_SW[5] 5.1e-21
C2171 a_11071_1642# a_11123_627# 1.92e-20
C2172 a_3947_627# a_3420_212# 7.07e-21
C2173 x8.X a_2897_1289# 1.51e-19
C2174 VDD a_14945_n62# 0.0149f
C2175 a_6753_1642# D[5] 0.00164f
C2176 a_7203_627# a_7823_601# 0.149f
C2177 D[4] a_7369_627# 0.168f
C2178 a_8679_1642# x14.X 9.51e-21
C2179 a_7369_627# VSS_SW[4] 0.023f
C2180 VDD a_7394_1315# 4.95e-19
C2181 x2.X a_1501_122# 0.0043f
C2182 VDD_SW_b[7] a_3333_601# 8.35e-20
C2183 a_11325_1642# m1_95_2154# 8.35e-20
C2184 a_2470_90# a_2879_n62# 4.24e-20
C2185 VSS_SW_b[7] a_1745_n62# 6.94e-20
C2186 check[0] a_15585_n88# 2.51e-19
C2187 a_4977_627# a_6920_627# 2e-20
C2188 VDD_SW_b[5] a_4958_n88# 3.23e-19
C2189 a_12036_1467# x15.X 4.97e-19
C2190 check[5] a_3333_601# 2.14e-19
C2191 a_8731_627# a_9595_627# 1.09e-19
C2192 a_9312_627# D[3] 4.28e-19
C2193 VDD_SW_b[4] VSS_SW_b[3] 0.0323f
C2194 VDD a_593_n62# 0.0155f
C2195 a_381_627# VSS_SW_b[7] 7.36e-20
C2196 a_305_2457# check[6] 0.00376f
C2197 a_9646_90# VSS_SW_b[3] 0.19f
C2198 a_7681_1289# a_7350_n88# 5.67e-21
C2199 a_12680_106# a_14526_n88# 1.86e-21
C2200 VDD_SW_b[6] a_2985_n62# 4.77e-19
C2201 a_7203_627# a_7757_627# 0.00206f
C2202 a_505_1289# a_487_n62# 3.44e-19
C2203 D[4] a_8342_304# 9.58e-19
C2204 a_7967_627# VSS_SW[4] 0.0012f
C2205 a_8204_212# VSS_SW_b[4] 0.00119f
C2206 a_8205_n88# a_8677_122# 0.15f
C2207 VSS_SW[4] a_8342_304# 1.97e-20
C2208 a_5289_1289# a_5504_106# 5.3e-21
C2209 a_10509_601# D[2] 9.63e-19
C2210 a_939_2457# VSS_SW[6] 0.0213f
C2211 a_10983_895# a_11987_627# 6.86e-19
C2212 VSS_SW[6] VSS_SW_b[6] 0.0072f
C2213 a_10983_895# VDD_SW_b[3] 0.129f
C2214 D[3] a_11987_627# 9.94e-20
C2215 x17.X x18.X 0.109f
C2216 a_5675_909# VDD_SW[5] 1.01e-20
C2217 D[3] VDD_SW_b[3] 0.453f
C2218 VDD x3.X 0.787f
C2219 a_15853_122# VSS_SW_b[1] 7.15e-19
C2220 a_9595_627# a_10824_993# 0.14f
C2221 a_8679_1642# a_8591_895# 5.45e-19
C2222 D[7] a_2470_90# 8.78e-19
C2223 x2.X a_6730_n62# 1.83e-19
C2224 a_4958_n88# a_5504_106# 0.207f
C2225 a_8117_601# a_9761_627# 6.5e-20
C2226 a_12901_601# a_12851_909# 1.21e-20
C2227 a_12153_627# a_12751_627# 6.04e-20
C2228 check[1] D[2] 0.46f
C2229 a_29_2457# x9.A1 9.28e-20
C2230 x13.X check[2] 5.59e-19
C2231 a_2419_627# VDD_SW[6] 3.29e-20
C2232 VDD a_7896_106# 0.356f
C2233 D[6] a_3755_627# 2e-19
C2234 x2.X a_10545_304# 0.00167f
C2235 a_15293_601# m1_95_1942# 4.09e-20
C2236 D[1] m1_95_2154# 0.0343f
C2237 a_2419_627# a_2470_90# 6.13e-19
C2238 a_14379_627# a_14545_627# 0.786f
C2239 x9.A1 a_12399_1315# 0.00504f
C2240 a_10288_106# VSS_SW[2] 9.05e-21
C2241 a_10597_n88# a_10711_n62# 2.14e-20
C2242 VDD_SW[6] m1_95_2154# 0.0327f
C2243 a_10596_212# a_10937_n62# 0.00134f
C2244 VDD_SW_b[2] a_14545_627# 0.00329f
C2245 x9.A1 D[4] 0.253f
C2246 a_305_2457# D[7] 1.02e-19
C2247 x3.X a_27_627# 5.4e-19
C2248 x9.A1 VSS_SW[4] 0.403f
C2249 a_10215_601# a_10596_212# 4.51e-19
C2250 a_10041_993# a_10288_106# 4.96e-20
C2251 a_10509_601# a_10055_n62# 3.74e-20
C2252 a_6285_122# VSS_SW_b[5] 7.14e-19
C2253 x10.X check[4] 0.00903f
C2254 x12.X VDD_SW[5] 0.305f
C2255 x11.X a_7203_627# 0.00295f
C2256 x9.A1 a_4528_627# 2e-20
C2257 x2.X a_12517_993# 5.32e-19
C2258 x2.X x13.X 0.00458f
C2259 a_6539_1642# a_6467_1642# 6.64e-19
C2260 a_8591_895# a_8409_n88# 4.26e-19
C2261 a_8117_601# a_8677_122# 2.7e-19
C2262 a_15767_895# VDD_SW_b[1] 0.128f
C2263 x20.X a_15767_895# 0.00655f
C2264 a_7350_n88# a_7854_220# 0.00869f
C2265 a_2585_627# a_3648_993# 0.0334f
C2266 a_2865_993# a_3333_601# 0.0633f
C2267 x2.X a_964_n62# 3.68e-20
C2268 check[4] D[5] 0.452f
C2269 a_3112_106# a_3420_212# 0.14f
C2270 a_2879_n62# a_3421_n88# 0.125f
C2271 a_8933_1642# m1_95_1942# 1.97e-19
C2272 a_15585_n88# a_15721_n62# 0.0697f
C2273 VDD a_13216_993# 0.189f
C2274 VSS_SW_b[1] a_15316_n62# 1.68e-19
C2275 a_4811_627# a_7557_627# 4.46e-21
C2276 VDD a_6539_1315# 0.00149f
C2277 a_14825_993# a_14526_n88# 8.71e-20
C2278 a_14999_601# a_14839_n62# 0.0026f
C2279 a_1415_895# VSS_SW[6] 7.03e-21
C2280 VDD a_3625_n88# 0.491f
C2281 x2.X a_15143_627# 0.0388f
C2282 x14.X a_8591_895# 0.00863f
C2283 a_3895_1642# a_3648_993# 0.00176f
C2284 a_5323_2457# VSS_SW[4] 2.07e-19
C2285 a_305_2457# m1_95_2154# 6.79e-19
C2286 a_12901_601# a_13323_627# 1.96e-20
C2287 a_12433_993# VDD_SW[2] 4.17e-21
C2288 x17.X a_13461_122# 2.79e-19
C2289 a_4149_1642# VDD_SW[6] 0.00511f
C2290 VDD_SW[6] a_5257_993# 7.03e-20
C2291 a_13375_895# a_13515_627# 0.0383f
C2292 a_1757_1315# D[7] 0.00195f
C2293 VDD_SW_b[4] a_8409_n88# 0.00132f
C2294 D[4] a_9742_n88# 4.32e-19
C2295 VDD a_7823_601# 0.313f
C2296 VDD a_16037_1642# 8.63e-19
C2297 a_8677_122# a_9122_n62# 0.0369f
C2298 VDD a_15464_909# 0.0225f
C2299 a_7350_n88# VSS_SW[3] 4.28e-21
C2300 a_7663_n62# a_8545_n62# 0.00926f
C2301 a_7896_106# a_8319_n62# 0.00386f
C2302 a_3648_993# a_3183_627# 0.00316f
C2303 a_3333_601# a_3551_627# 3.73e-19
C2304 a_3039_601# VDD_SW_b[6] 1.75e-20
C2305 a_12134_n88# a_13461_122# 4.59e-22
C2306 a_12447_n62# a_13193_n88# 0.199f
C2307 a_12680_106# a_12989_n88# 0.0327f
C2308 a_16109_1642# a_16323_1642# 0.00557f
C2309 a_10597_n88# VSS_SW_b[2] 0.00487f
C2310 x18.X a_14545_627# 0.00314f
C2311 VDD_SW[2] a_14733_627# 6.11e-20
C2312 x13.X a_9312_627# 0.0338f
C2313 x14.X VDD_SW_b[4] 7.27e-19
C2314 VDD_SW_b[7] VSS_SW[6] 0.00248f
C2315 VDD x27.A 0.174f
C2316 a_9761_627# a_10125_993# 0.0018f
C2317 a_10215_601# a_9949_627# 8.07e-20
C2318 a_10509_601# a_10983_895# 0.265f
C2319 x14.X a_9646_90# 0.00259f
C2320 D[7] a_3421_n88# 9.66e-22
C2321 D[3] a_10509_601# 0.0191f
C2322 x2.X a_8204_212# 0.0128f
C2323 a_13906_n62# a_13705_n62# 3.81e-19
C2324 a_5271_n62# a_5950_304# 0.00652f
C2325 a_2897_1289# a_2585_627# 0.00323f
C2326 a_5504_106# a_5761_304# 0.00857f
C2327 x7.X D[6] 2.1e-19
C2328 check[5] VSS_SW[6] 0.034f
C2329 a_487_n62# a_1233_n88# 0.199f
C2330 x2.X a_13515_627# 0.0151f
C2331 a_174_n88# a_1501_122# 4.59e-22
C2332 a_720_106# a_1029_n88# 0.0327f
C2333 a_13375_895# VSS_SW[1] 7.03e-21
C2334 a_11325_1642# a_11704_627# 5.9e-19
C2335 x2.X a_4811_627# 0.354f
C2336 D[2] a_12341_627# 0.161f
C2337 a_11987_627# a_12517_993# 4.45e-20
C2338 VDD a_8623_220# 0.0117f
C2339 VDD x8.X 0.346f
C2340 a_2897_1289# a_3895_1642# 0.0146f
C2341 a_15143_627# a_15715_627# 2.46e-21
C2342 check[6] a_647_601# 0.00263f
C2343 a_7649_993# a_7557_627# 0.0369f
C2344 a_8117_601# a_8432_993# 0.13f
C2345 a_7823_601# a_7733_993# 6.69e-20
C2346 a_7369_627# a_8067_909# 0.00276f
C2347 a_16323_1642# VDD_SW[1] 5.32e-19
C2348 VDD a_16109_1642# 0.111f
C2349 a_8933_1642# VDD_SW[4] 0.00511f
C2350 x7.X m1_95_1942# 2.51e-20
C2351 check[1] D[3] 6.16e-20
C2352 a_16298_n62# a_16097_n62# 3.81e-19
C2353 x11.X a_6760_1315# 0.00143f
C2354 D[6] a_3420_212# 0.158f
C2355 a_2419_627# a_3421_n88# 1.06e-19
C2356 a_12465_1289# m1_95_1942# 2.26e-19
C2357 VSS_SW_b[5] a_5377_n62# 0.00334f
C2358 a_5813_n88# a_6153_n62# 6.04e-20
C2359 a_6017_n88# a_5927_n62# 9.75e-19
C2360 a_5812_212# VSS_SW[4] 0.0872f
C2361 VDD_SW_b[4] a_10680_909# 3.95e-21
C2362 x9.A1 check[6] 0.411f
C2363 a_10055_n62# a_10246_220# 3.24e-19
C2364 a_3420_212# m1_95_1942# 6.77e-21
C2365 a_4811_627# a_4977_627# 0.786f
C2366 VDD a_473_993# 0.218f
C2367 a_4811_627# VSS_SW[5] 0.0578f
C2368 x2.X VSS_SW[1] 0.0814f
C2369 VDD a_16330_1315# 3.48e-19
C2370 a_7203_627# D[3] 1.27e-20
C2371 VDD VDD_SW[1] 0.278f
C2372 a_8591_895# VDD_SW_b[4] 0.129f
C2373 D[4] a_9595_627# 1e-19
C2374 a_9312_627# a_8204_212# 6.63e-19
C2375 x8.X a_27_627# 0.00117f
C2376 VSS_SW_b[2] a_12638_220# 5.56e-20
C2377 a_12989_n88# a_13407_220# 0.00276f
C2378 a_12447_n62# a_14430_90# 6.12e-21
C2379 a_13193_n88# a_13126_304# 9.46e-19
C2380 a_12988_212# a_13705_304# 4.45e-20
C2381 x6.X a_473_993# 9.17e-20
C2382 a_12433_993# a_12134_n88# 8.71e-20
C2383 a_12607_601# a_12447_n62# 0.0026f
C2384 x2.X a_3893_122# 0.0043f
C2385 x9.A1 a_2879_n62# 8.79e-21
C2386 a_3421_n88# a_3558_304# 0.00907f
C2387 a_3420_212# a_3839_220# 2.46e-19
C2388 a_2879_n62# a_4338_n62# 3.79e-20
C2389 a_7369_627# m1_95_2154# 2.61e-20
C2390 a_4860_1467# check[4] 0.318f
C2391 a_10680_909# VDD_SW[3] 2.82e-20
C2392 check[0] a_16037_1642# 0.00577f
C2393 a_6920_627# a_7203_627# 0.0011f
C2394 x20.X a_14379_627# 2.67e-20
C2395 x9.A1 a_10597_n88# 8.52e-21
C2396 a_14379_627# VDD_SW_b[1] 1.15e-19
C2397 D[1] a_16024_909# 8.04e-19
C2398 check[6] a_505_1289# 0.25f
C2399 VDD a_13103_n62# 0.00521f
C2400 check[2] a_10596_212# 2.72e-20
C2401 VDD a_4862_90# 0.189f
C2402 VDD D[2] 0.968f
C2403 x2.X a_7649_993# 0.15f
C2404 a_14428_1467# VSS_SW[1] 0.0273f
C2405 a_4811_627# a_5575_627# 0.00134f
C2406 D[5] a_6124_993# 2.48e-19
C2407 VDD x11.X 0.474f
C2408 x2.X a_11325_1315# 2.32e-19
C2409 VDD a_1159_627# 6.2e-19
C2410 D[2] a_14096_627# 0.00238f
C2411 D[7] a_647_601# 0.00584f
C2412 a_27_627# a_473_993# 0.159f
C2413 VDD_SW_b[4] a_9646_90# 0.00345f
C2414 check[3] a_7254_90# 2.5e-20
C2415 x14.X a_11071_1642# 1.97e-20
C2416 VSS_SW_b[6] a_3761_n62# 5.35e-19
C2417 a_3893_122# VSS_SW[5] 6.63e-20
C2418 VDD a_1503_1642# 0.194f
C2419 VDD a_9786_1315# 0.00121f
C2420 VDD a_5165_627# 0.109f
C2421 a_2865_993# VSS_SW[6] 0.00296f
C2422 x6.X a_1503_1642# 1.98e-20
C2423 a_16109_1642# check[0] 0.318f
C2424 x20.X a_15072_106# 1.89e-20
C2425 x9.A1 D[7] 0.268f
C2426 x2.X a_10596_212# 0.0128f
C2427 VDD_SW_b[1] a_15072_106# 5.22e-19
C2428 a_4689_2457# check[4] 0.00137f
C2429 x2.X a_8335_627# 0.00702f
C2430 a_10734_304# VSS_SW[2] 2.76e-20
C2431 x9.A1 a_6529_n62# 5.7e-21
C2432 x2.X a_8921_304# 3.27e-19
C2433 a_5271_n62# a_7350_n88# 3.08e-21
C2434 a_6539_1642# a_6199_895# 0.00226f
C2435 D[3] a_10246_220# 1.98e-20
C2436 a_1028_212# a_1946_n62# 0.0453f
C2437 a_1233_n88# a_1447_220# 0.0104f
C2438 a_487_n62# a_593_n62# 0.0526f
C2439 a_1029_n88# a_1745_304# 0.0018f
C2440 check[4] a_6285_1642# 0.256f
C2441 a_27_627# a_1159_627# 0.00272f
C2442 a_9742_n88# a_10597_n88# 0.0477f
C2443 x8.X VDD_SW[7] 0.305f
C2444 a_13103_n62# a_13329_n62# 3.34e-19
C2445 VDD a_10055_n62# 0.326f
C2446 a_12036_1467# a_12134_n88# 6.87e-20
C2447 a_11987_627# VSS_SW[1] 4.95e-21
C2448 check[5] check[4] 0.00523f
C2449 a_193_627# m1_95_1942# 3.82e-20
C2450 a_647_601# m1_95_2154# 2.34e-20
C2451 a_9644_1467# VSS_SW_b[3] 2.13e-19
C2452 x9.A1 a_2419_627# 7.97e-19
C2453 a_505_1289# D[7] 0.0661f
C2454 check[0] VDD_SW[1] 0.00392f
C2455 D[6] a_4137_304# 8.38e-19
C2456 a_10983_895# a_12341_627# 8.26e-21
C2457 VDD VSS_SW_b[1] 0.133f
C2458 x13.X a_10509_601# 4.31e-21
C2459 x2.X a_941_601# 0.119f
C2460 a_9786_1642# VSS_SW[3] 0.00105f
C2461 x9.A1 a_4077_1642# 5.26e-19
C2462 a_6017_n88# VSS_SW_b[4] 4.54e-20
C2463 a_5377_n62# a_5748_n62# 4.19e-20
C2464 a_6529_304# VSS_SW[4] 6.59e-21
C2465 x10.X a_3807_895# 0.00864f
C2466 a_6539_1642# VDD_SW_b[5] 2.59e-19
C2467 ready VSS_SW[7] 0.0387f
C2468 x9.A1 a_535_1642# 5.26e-19
C2469 x9.A1 m1_95_2154# 6.12f
C2470 a_941_601# a_1363_627# 1.96e-20
C2471 a_473_993# VDD_SW[7] 4.17e-21
C2472 a_1415_895# a_1555_627# 0.0383f
C2473 VDD_SW_b[2] a_13705_n62# 5.22e-19
C2474 a_12901_601# m1_95_2154# 2.84e-20
C2475 check[0] D[2] 5.94e-20
C2476 a_647_601# a_1112_909# 9.46e-19
C2477 a_7967_627# a_8539_627# 2.46e-21
C2478 check[2] x15.X 0.00965f
C2479 x2.X a_2985_n62# 5.25e-20
C2480 a_3648_993# a_4811_627# 7.46e-20
C2481 a_3807_895# D[5] 2.17e-19
C2482 a_3421_n88# a_4958_n88# 1.98e-19
C2483 a_3420_212# a_5271_n62# 2.62e-19
C2484 VDD_SW_b[5] a_8288_909# 2.96e-21
C2485 x2.X a_9949_627# 0.00141f
C2486 x2.X a_1672_909# 4.02e-19
C2487 a_505_1289# m1_95_2154# 1.04e-19
C2488 VDD a_5813_n88# 0.714f
C2489 x9.X a_4528_627# 0.0337f
C2490 VDD_SW_b[7] a_1745_n62# 5.22e-19
C2491 a_2585_627# a_2566_n88# 4.91e-19
C2492 x10.X VDD_SW_b[6] 7.23e-19
C2493 a_14857_1289# a_14999_601# 8.76e-20
C2494 a_14999_601# a_15608_993# 0.00189f
C2495 a_14545_627# a_14733_627# 0.189f
C2496 a_6199_895# m1_95_1942# 8.63e-20
C2497 a_6040_993# m1_95_2154# 4.11e-21
C2498 a_7252_1467# VDD_SW[5] 0.00487f
C2499 x2.X a_2927_1642# 2.62e-19
C2500 VDD_SW_b[3] a_10596_212# 0.0417f
C2501 a_7394_1315# D[4] 7.54e-19
C2502 check[4] x12.X 5.98e-19
C2503 a_14839_n62# a_15030_220# 3.3e-19
C2504 VDD a_2585_627# 0.749f
C2505 a_7394_1315# VSS_SW[4] 7.95e-19
C2506 a_9761_627# VSS_SW_b[3] 5.23e-20
C2507 a_5323_2457# m1_95_2154# 0.00298f
C2508 x13.X a_7203_627# 2.67e-20
C2509 VSS_SW[1] a_15853_122# 2.79e-21
C2510 a_9595_627# a_10597_n88# 1.06e-19
C2511 VDD a_10983_895# 0.687f
C2512 x2.X a_5341_993# 5.3e-19
C2513 VDD D[3] 1.17f
C2514 x9.A1 a_4149_1642# 0.195f
C2515 x9.A1 a_5257_993# 9.52e-20
C2516 check[3] a_8205_n88# 7.34e-21
C2517 x2.X x15.X 0.00458f
C2518 VDD_SW_b[6] D[5] 1.57e-19
C2519 a_3356_n62# a_3761_n62# 2.46e-21
C2520 a_7252_1467# a_7711_1642# 6.64e-19
C2521 VDD_SW_b[2] a_12680_106# 5.23e-19
C2522 VDD a_3895_1642# 0.212f
C2523 x7.X a_1028_212# 0.245f
C2524 check[6] a_1233_n88# 2.51e-19
C2525 check[3] D[5] 6.36e-20
C2526 VDD a_6920_627# 0.198f
C2527 VDD a_15495_n62# 0.00713f
C2528 ready a_3333_601# 5.7e-21
C2529 a_3183_627# a_2566_n88# 1.08e-19
C2530 a_3648_993# a_3893_122# 1.51e-20
C2531 reset a_939_2457# 4.31e-19
C2532 a_29_2457# x3.X 6.66e-19
C2533 x3.A a_305_2457# 0.3f
C2534 check[4] a_6285_122# 2.99e-20
C2535 VDD_SW_b[5] m1_95_1942# 2.88e-20
C2536 VDD a_8933_1315# 0.00183f
C2537 a_13715_1642# m1_95_2154# 8.35e-20
C2538 check[0] VSS_SW_b[1] 9.18e-21
C2539 VDD a_3183_627# 0.00932f
C2540 a_5812_212# a_6529_n62# 0.00206f
C2541 check[5] a_3761_n62# 9.81e-20
C2542 a_1028_212# a_3420_212# 1.9e-21
C2543 a_1029_n88# a_3112_106# 1.67e-21
C2544 a_1501_122# a_2566_n88# 8e-21
C2545 a_27_627# a_2585_627# 1.15e-20
C2546 a_5725_601# a_6199_895# 0.265f
C2547 check[1] a_13515_627# 1.9e-19
C2548 a_5431_601# a_5165_627# 8.07e-20
C2549 a_4977_627# a_5341_993# 0.0018f
C2550 a_10055_n62# a_10288_106# 0.124f
C2551 VDD a_1501_122# 0.313f
C2552 x2.X a_2468_1467# 3.56e-19
C2553 a_5323_2457# a_5257_993# 8.63e-21
C2554 a_8677_122# VSS_SW_b[3] 1.02e-20
C2555 a_12988_212# a_14839_n62# 2.62e-19
C2556 a_12989_n88# a_14526_n88# 1.98e-19
C2557 D[6] a_5504_106# 1.39e-21
C2558 VDD_SW_b[3] a_11313_n62# 5.22e-19
C2559 x9.A1 a_11313_304# 8.15e-21
C2560 VDD_SW[5] a_8591_895# 1.27e-20
C2561 a_7203_627# a_8204_212# 6.99e-20
C2562 D[4] a_7896_106# 8.71e-19
C2563 a_14545_627# a_16488_627# 1.79e-20
C2564 x9.A1 a_5289_1289# 0.105f
C2565 a_7254_90# VSS_SW_b[4] 0.19f
C2566 VSS_SW[4] a_7896_106# 4.63e-19
C2567 a_1757_1642# x8.X 7.97e-19
C2568 a_5504_106# m1_95_1942# 4.96e-22
C2569 a_5725_601# VDD_SW_b[5] 0.00636f
C2570 a_4811_627# a_7203_627# 1.63e-20
C2571 a_6040_993# a_5943_627# 0.00386f
C2572 a_6199_895# a_6456_909# 0.00869f
C2573 a_5165_627# a_5365_627# 3.81e-19
C2574 a_12607_601# m1_95_1942# 3.42e-20
C2575 x8.X a_2773_627# 6.12e-19
C2576 check[3] a_8117_601# 1.7e-19
C2577 check[1] VSS_SW[1] 1.4e-19
C2578 a_9644_1467# x14.X 0.0877f
C2579 D[7] a_1233_n88# 0.00546f
C2580 x9.A1 a_4958_n88# 7.34e-19
C2581 x2.X a_6017_n88# 0.00369f
C2582 a_12433_993# a_12751_627# 0.025f
C2583 a_12153_627# a_13119_627# 2.14e-20
C2584 a_12901_601# a_13300_993# 9.41e-19
C2585 a_12341_627# a_12517_993# 8.99e-19
C2586 x16.X VDD_SW[3] 0.307f
C2587 x15.X a_11987_627# 0.00297f
C2588 a_3893_122# a_4137_n62# 0.00807f
C2589 a_9595_627# m1_95_2154# 3.53e-20
C2590 a_4338_n62# a_4958_n88# 8.26e-21
C2591 x15.X VDD_SW_b[3] 0.219f
C2592 a_10007_1315# D[3] 0.00202f
C2593 x2.X a_3039_601# 0.2f
C2594 VDD a_6730_n62# 0.111f
C2595 D[6] a_3504_909# 8.51e-19
C2596 a_2419_627# a_3732_993# 2.13e-19
C2597 x2.X a_11015_220# 9.52e-19
C2598 a_14857_1289# m1_95_1942# 2.26e-19
C2599 a_15608_993# m1_95_1942# 5.78e-21
C2600 VDD_SW[7] a_2585_627# 9.25e-19
C2601 a_2136_627# a_3333_601# 1.84e-20
C2602 a_6456_909# VDD_SW_b[5] 3.4e-20
C2603 a_5323_2457# a_5289_1289# 6.83e-20
C2604 D[1] a_14999_601# 0.00585f
C2605 a_14379_627# a_14825_993# 0.159f
C2606 a_10597_n88# VSS_SW[2] 9.22e-19
C2607 a_10801_n88# a_10937_n62# 0.0697f
C2608 VSS_SW_b[3] a_10532_n62# 1.68e-19
C2609 VDD_SW_b[2] a_14825_993# 8.2e-21
C2610 x9.X a_2879_n62# 0.00192f
C2611 a_10509_601# a_10596_212# 6.03e-19
C2612 a_10824_993# a_10055_n62# 3.59e-19
C2613 x2.X a_6339_627# 0.0151f
C2614 D[3] a_10288_106# 8.76e-19
C2615 VDD a_10545_304# 0.00269f
C2616 a_5725_601# a_5504_106# 3.46e-19
C2617 a_6199_895# a_5271_n62# 0.00219f
C2618 a_5431_601# a_5813_n88# 0.00322f
C2619 a_4977_627# a_6017_n88# 8.75e-19
C2620 a_8679_1642# a_8677_122# 1.57e-21
C2621 VSS_SW[5] a_6017_n88# 9.93e-21
C2622 a_193_627# a_1028_212# 1.02e-19
C2623 a_647_601# a_720_106# 1.01e-19
C2624 a_13461_122# a_13705_n62# 0.00807f
C2625 a_13906_n62# a_14526_n88# 8.26e-21
C2626 a_473_993# a_487_n62# 2.63e-19
C2627 a_941_601# a_174_n88# 0.00259f
C2628 x7.X a_1946_n62# 0.0016f
C2629 x2.X a_13072_909# 0.00309f
C2630 a_1029_n88# m1_95_1942# 1.16e-21
C2631 x2.X a_2973_627# 3.94e-19
C2632 x9.A1 a_11704_627# 2e-20
C2633 a_11704_627# a_12901_601# 1.71e-20
C2634 VDD_SW[3] a_12153_627# 9.25e-19
C2635 D[4] a_7823_601# 0.00584f
C2636 a_7203_627# a_7649_993# 0.159f
C2637 a_15855_1642# x20.X 1.31e-19
C2638 a_7823_601# VSS_SW[4] 6.25e-19
C2639 x14.X a_9761_627# 0.00312f
C2640 x2.X VSS_SW_b[7] 0.0279f
C2641 a_11325_1642# m1_95_1942# 1.97e-19
C2642 VDD a_12517_993# 0.00579f
C2643 VSS_SW_b[1] a_15721_n62# 5.35e-19
C2644 a_15853_122# a_16097_n62# 0.00807f
C2645 a_1946_n62# a_3420_212# 5.58e-22
C2646 VDD x13.X 0.632f
C2647 a_15293_601# a_14839_n62# 3.74e-20
C2648 a_14825_993# a_15072_106# 4.96e-20
C2649 x2.X a_13715_1315# 2.33e-19
C2650 a_14545_627# a_15381_n88# 1.27e-19
C2651 x2.X a_15511_627# 0.00702f
C2652 a_14999_601# a_15380_212# 4.51e-19
C2653 VDD_SW_b[5] a_5271_n62# 5.28e-19
C2654 check[5] a_3807_895# 0.00272f
C2655 VDD a_964_n62# 0.00116f
C2656 a_13375_895# VDD_SW[2] 0.00356f
C2657 a_13216_993# a_13323_627# 0.00707f
C2658 x3.X check[6] 0.0144f
C2659 a_7681_1289# a_7663_n62# 3.44e-19
C2660 a_11071_1642# x16.X 1.52e-20
C2661 VDD_SW_b[6] a_3356_n62# 8.1e-20
C2662 x27.A a_4528_627# 1.61e-19
C2663 VDD a_15143_627# 0.00929f
C2664 a_7203_627# a_8335_627# 0.00272f
C2665 VDD a_12178_1315# 0.00189f
C2666 a_505_1289# a_720_106# 5.3e-21
C2667 D[4] a_8623_220# 7.05e-19
C2668 a_7757_627# VSS_SW[4] 3.79e-19
C2669 a_12988_212# a_13193_n88# 0.15f
C2670 VSS_SW[2] a_12638_220# 4.26e-19
C2671 a_12447_n62# VSS_SW_b[2] 0.0142f
C2672 VSS_SW[4] a_8623_220# 6.42e-21
C2673 a_8205_n88# VSS_SW_b[4] 7.59e-19
C2674 a_8409_n88# a_8677_122# 0.206f
C2675 a_9644_1467# a_9646_90# 1e-19
C2676 a_13715_1642# a_13936_1315# 0.00783f
C2677 ready VSS_SW[6] 0.0361f
C2678 x18.X a_14825_993# 9.17e-20
C2679 a_5896_909# VDD_SW[5] 2.82e-20
C2680 a_11069_122# VSS_SW_b[2] 1.16e-20
C2681 VDD_SW[2] a_15243_909# 2.16e-20
C2682 a_2610_1315# D[6] 7.54e-19
C2683 a_10509_601# a_9949_627# 1.24e-20
C2684 a_10983_895# a_10824_993# 0.207f
C2685 a_9761_627# a_10680_909# 0.00907f
C2686 D[5] VSS_SW_b[4] 2.02e-19
C2687 check[5] VDD_SW_b[6] 0.00208f
C2688 a_6285_1642# check[3] 9.11e-21
C2689 D[3] a_10824_993# 0.00609f
C2690 a_10149_627# VSS_SW[3] 3.79e-19
C2691 x9.X a_2419_627# 2.64e-20
C2692 a_8679_1642# a_8432_993# 0.00176f
C2693 x2.X a_7254_90# 0.00368f
C2694 VDD_SW_b[6] a_5675_909# 2.62e-21
C2695 VSS_SW[2] m1_95_2154# 0.0337f
C2696 x2.X VDD_SW[2] 0.0327f
C2697 a_8117_601# a_10215_601# 1.75e-20
C2698 a_4958_n88# a_5812_212# 0.0319f
C2699 a_5271_n62# a_5504_106# 0.124f
C2700 a_8591_895# a_9761_627# 2.64e-19
C2701 a_10041_993# m1_95_2154# 1.86e-20
C2702 x30.A VDD_SW[6] 0.0077f
C2703 a_11987_627# a_13072_909# 1.09e-19
C2704 D[2] a_12851_909# 6.77e-19
C2705 x9.X m1_95_2154# 1.31e-20
C2706 VDD_SW_b[3] a_13072_909# 2.96e-21
C2707 x20.X a_16488_627# 0.0338f
C2708 D[6] VDD_SW[6] 0.227f
C2709 VDD a_8204_212# 0.712f
C2710 x3.A x9.A1 1.27e-19
C2711 VDD_SW_b[1] a_16488_627# 0.186f
C2712 x15.X a_10509_601# 1.29e-19
C2713 VDD a_13515_627# 6.99e-19
C2714 a_15495_n62# a_15721_n62# 3.34e-19
C2715 D[1] m1_95_1942# 0.0335f
C2716 VDD a_4811_627# 0.426f
C2717 a_14428_1467# VDD_SW[2] 0.00484f
C2718 VDD_SW[6] m1_95_1942# 0.0331f
C2719 x3.X D[7] 1.77e-19
C2720 a_12399_1315# D[2] 0.00202f
C2721 x17.X a_13375_895# 0.00662f
C2722 a_10288_106# a_10545_304# 0.00857f
C2723 a_10055_n62# a_10734_304# 0.00652f
C2724 VDD_SW_b[4] a_9761_627# 0.00344f
C2725 x15.X check[1] 5.58e-19
C2726 x7.X a_3420_212# 1.68e-21
C2727 a_7681_1289# a_7369_627# 0.00323f
C2728 a_9122_n62# a_8921_n62# 3.81e-19
C2729 a_7203_627# a_9949_627# 4.74e-21
C2730 x11.X D[4] 2.11e-19
C2731 x9.A1 a_3947_627# 5.22e-20
C2732 x11.X VSS_SW[4] 0.138f
C2733 a_12989_n88# a_13906_n62# 0.189f
C2734 a_13193_n88# a_13705_304# 6.69e-20
C2735 a_12988_212# a_14430_90# 0.00101f
C2736 VSS_SW_b[2] a_13126_304# 3.87e-20
C2737 a_12607_601# a_12988_212# 4.51e-19
C2738 a_12153_627# a_12989_n88# 1.27e-19
C2739 a_12901_601# a_12447_n62# 3.74e-20
C2740 a_12433_993# a_12680_106# 4.96e-20
C2741 a_8432_993# a_8409_n88# 1.86e-19
C2742 a_8591_895# a_8677_122# 4.53e-22
C2743 a_7252_1467# check[4] 1.57e-19
C2744 a_2585_627# a_2773_627# 0.189f
C2745 a_7663_n62# a_7854_220# 3.24e-19
C2746 x9.A1 a_1745_304# 6.9e-21
C2747 a_3039_601# a_3648_993# 0.00189f
C2748 a_4149_1642# x9.X 0.0841f
C2749 x9.A1 a_11069_122# 3.99e-20
C2750 a_3112_106# a_3421_n88# 0.0327f
C2751 a_2566_n88# a_3893_122# 4.59e-22
C2752 VDD VSS_SW[1] 0.98f
C2753 a_2879_n62# a_3625_n88# 0.199f
C2754 a_9761_627# VDD_SW[3] 1.96e-20
C2755 check[2] a_10801_n88# 2.02e-19
C2756 a_15380_212# m1_95_1942# 6.77e-21
C2757 a_9595_627# a_11704_627# 1.75e-19
C2758 x12.X check[3] 0.00903f
C2759 a_2136_627# VSS_SW[6] 0.00164f
C2760 x10.X a_5223_1315# 2.41e-19
C2761 VDD a_3893_122# 0.314f
C2762 x14.X a_8432_993# 2.78e-19
C2763 a_14379_627# a_14526_n88# 0.00176f
C2764 VDD_SW_b[2] a_14526_n88# 5.91e-19
C2765 x2.X x17.X 0.00464f
C2766 a_14096_627# VSS_SW[1] 0.00166f
C2767 x3.X m1_95_2154# 0.00106f
C2768 a_305_2457# m1_95_1942# 3.15e-19
C2769 VDD_SW[6] a_5725_601# 2.46e-20
C2770 a_11987_627# VDD_SW[2] 3.29e-20
C2771 D[2] a_13323_627# 2e-19
C2772 x16.X a_12153_627# 0.00313f
C2773 a_5223_1315# D[5] 0.00202f
C2774 D[4] a_10055_n62# 1.56e-21
C2775 VDD_SW_b[4] a_8677_122# 0.00445f
C2776 VDD a_7649_993# 0.18f
C2777 a_8204_212# a_8319_n62# 0.00272f
C2778 a_3333_601# a_4064_909# 0.0016f
C2779 a_7663_n62# VSS_SW[3] 1.64e-20
C2780 a_7896_106# a_8545_n62# 0.00316f
C2781 a_2865_993# VDD_SW_b[6] 4.91e-21
C2782 x2.X a_12134_n88# 0.178f
C2783 VDD a_11325_1315# 4.79e-19
C2784 a_76_1467# VSS_SW_b[7] 7.31e-20
C2785 check[6] x8.X 5.86e-19
C2786 x2.X a_10801_n88# 0.00369f
C2787 x20.X a_15381_n88# 0.0189f
C2788 VDD_SW_b[1] a_15381_n88# 0.0406f
C2789 x2.X x10.X 3.64e-19
C2790 a_11313_304# VSS_SW[2] 6.58e-21
C2791 a_14428_1467# x17.X 4.9e-19
C2792 a_10215_601# a_10125_993# 6.69e-20
C2793 a_13929_1642# VDD_SW[2] 5.15e-19
C2794 D[3] a_10734_304# 9.69e-19
C2795 x2.X a_8205_n88# 0.0213f
C2796 a_2897_1289# a_3039_601# 8.76e-20
C2797 a_1978_1315# VDD_SW_b[7] 2.64e-20
C2798 a_5271_n62# a_6231_220# 1.21e-20
C2799 a_5812_212# a_5761_304# 2.13e-19
C2800 check[4] a_5319_1642# 0.00526f
C2801 a_14526_n88# a_15072_106# 0.207f
C2802 a_5813_n88# a_5462_220# 4.48e-20
C2803 a_5504_106# a_5950_304# 0.00412f
C2804 a_9742_n88# a_11069_122# 4.59e-22
C2805 a_1028_212# a_1029_n88# 0.784f
C2806 VDD a_10596_212# 0.704f
C2807 VSS_SW[7] a_678_220# 4.25e-19
C2808 a_487_n62# a_1501_122# 0.0633f
C2809 a_720_106# a_1233_n88# 0.00189f
C2810 a_174_n88# VSS_SW_b[7] 0.135f
C2811 VDD a_8335_627# 0.00124f
C2812 x2.X D[5] 0.18f
C2813 VDD a_8921_304# 0.0062f
C2814 x7.X a_193_627# 1.13e-20
C2815 a_8204_212# a_10288_106# 5.86e-20
C2816 a_7369_627# a_8288_909# 0.00907f
C2817 a_7823_601# a_8067_909# 0.0104f
C2818 a_7649_993# a_7733_993# 0.00972f
C2819 a_8591_895# a_8432_993# 0.207f
C2820 a_8117_601# a_7557_627# 1.15e-20
C2821 check[6] a_473_993# 7.17e-20
C2822 x9.A1 a_7681_1289# 0.105f
C2823 x10.X a_4977_627# 0.00315f
C2824 a_2419_627# a_3625_n88# 0.00204f
C2825 D[6] a_3421_n88# 0.158f
C2826 x10.X VSS_SW[5] 0.251f
C2827 x9.X a_4958_n88# 0.00863f
C2828 D[1] a_15030_220# 2.03e-20
C2829 check[0] VSS_SW[1] 0.0493f
C2830 a_6017_n88# a_6153_n62# 0.0697f
C2831 a_5813_n88# VSS_SW[4] 9.23e-19
C2832 VSS_SW_b[5] a_5748_n62# 1.68e-19
C2833 a_13216_993# m1_95_2154# 4.11e-21
C2834 x9.A1 a_14999_601# 2.81e-20
C2835 a_12901_601# a_14999_601# 1.52e-20
C2836 a_13375_895# a_14545_627# 2.96e-19
C2837 D[5] a_4977_627# 0.168f
C2838 x17.X a_11987_627# 2.67e-20
C2839 a_3421_n88# m1_95_1942# 1.16e-21
C2840 a_4811_627# a_5431_601# 0.149f
C2841 D[5] VSS_SW[5] 0.119f
C2842 VDD a_941_601# 0.474f
C2843 D[4] D[3] 0.00183f
C2844 a_8432_993# VDD_SW_b[4] 5.63e-20
C2845 x13.X a_9154_1315# 0.00146f
C2846 x2.X a_12937_304# 0.00168f
C2847 a_8731_627# a_8204_212# 7.07e-21
C2848 a_7369_627# VSS_SW[3] 4.78e-21
C2849 x8.X D[7] 9.68e-19
C2850 a_12447_n62# a_12553_n62# 0.0526f
C2851 x2.X VSS_SW_b[6] 0.0278f
C2852 x6.X a_941_601# 4.9e-20
C2853 a_939_2457# x2.X 1.72f
C2854 a_2585_627# a_4528_627# 2e-20
C2855 x20.X a_16298_n62# 0.00153f
C2856 a_7369_627# m1_95_1942# 3.82e-20
C2857 a_2566_n88# a_2985_n62# 0.0383f
C2858 a_11987_627# a_12134_n88# 0.00176f
C2859 a_3421_n88# a_3839_220# 0.00276f
C2860 VSS_SW_b[6] a_3070_220# 5.34e-20
C2861 a_3625_n88# a_3558_304# 9.46e-19
C2862 a_3420_212# a_4137_304# 4.45e-20
C2863 a_2879_n62# a_4862_90# 6.12e-21
C2864 a_7823_601# m1_95_2154# 2.34e-20
C2865 VDD_SW_b[1] a_16298_n62# 0.0143f
C2866 a_12038_90# VSS_SW_b[2] 0.191f
C2867 a_6339_627# a_7203_627# 1.09e-19
C2868 a_6920_627# D[4] 4.42e-19
C2869 a_11704_627# VSS_SW[2] 0.00163f
C2870 VDD_SW_b[3] a_12134_n88# 5.9e-19
C2871 a_14545_627# a_15243_909# 0.00276f
C2872 a_15293_601# a_15608_993# 0.13f
C2873 a_6920_627# VSS_SW[4] 0.00164f
C2874 a_14999_601# a_14909_993# 6.69e-20
C2875 check[6] a_1503_1642# 0.257f
C2876 VDD_SW_b[5] a_7350_n88# 5.9e-19
C2877 a_14825_993# a_14733_627# 0.0369f
C2878 VDD_SW_b[3] a_10801_n88# 0.00132f
C2879 VDD a_2985_n62# 0.0149f
C2880 a_8933_1315# D[4] 0.00195f
C2881 x2.X a_8117_601# 0.119f
C2882 a_14839_n62# a_15518_304# 0.00652f
C2883 a_15072_106# a_15329_304# 0.00857f
C2884 a_4811_627# a_5365_627# 0.00206f
C2885 x27.A m1_95_2154# 1.87e-19
C2886 x10.X a_4370_1315# 3.75e-20
C2887 VDD a_9949_627# 0.11f
C2888 x2.X a_14545_627# 0.0537f
C2889 VDD a_1672_909# 0.0044f
C2890 x8.X a_2419_627# 0.236f
C2891 x9.A1 a_6539_1642# 0.195f
C2892 VDD_SW_b[4] a_7769_n62# 4.77e-19
C2893 a_27_627# a_941_601# 0.14f
C2894 D[7] a_473_993# 0.00884f
C2895 a_8933_1642# a_8861_1642# 6.64e-19
C2896 VDD_SW_b[2] a_12989_n88# 0.0406f
C2897 a_8342_304# VSS_SW[3] 2.77e-20
C2898 a_3283_909# VDD_SW[6] 1.01e-20
C2899 VDD a_2927_1642# 0.00171f
C2900 x16.X a_9761_627# 6.37e-20
C2901 x8.X m1_95_2154# 6.47e-20
C2902 VDD a_5341_993# 0.00431f
C2903 a_16109_1642# m1_95_2154# 8.35e-20
C2904 a_3333_601# VSS_SW[6] 2.13e-19
C2905 VDD x15.X 0.671f
C2906 a_5725_601# a_7369_627# 6.25e-20
C2907 x2.X a_8848_909# 4.02e-19
C2908 x2.X a_9122_n62# 1.87e-19
C2909 a_5504_106# a_7350_n88# 1.86e-21
C2910 check[1] VDD_SW[2] 0.00389f
C2911 a_720_106# a_593_n62# 0.0256f
C2912 a_487_n62# a_964_n62# 1.96e-20
C2913 VSS_SW_b[7] a_1166_304# 3.58e-20
C2914 a_1028_212# a_2470_90# 0.00101f
C2915 a_1233_n88# a_1745_304# 6.69e-20
C2916 a_1029_n88# a_1946_n62# 0.189f
C2917 x16.X a_13461_1642# 2.02e-20
C2918 D[7] a_1159_627# 6.12e-19
C2919 a_10288_106# a_10596_212# 0.14f
C2920 a_10055_n62# a_10597_n88# 0.125f
C2921 a_5323_2457# a_6539_1642# 0.00112f
C2922 x2.X a_4860_1467# 2.87e-19
C2923 a_13461_122# a_14526_n88# 8e-21
C2924 a_8117_601# a_9312_627# 5.84e-19
C2925 a_12989_n88# a_15072_106# 1.67e-21
C2926 a_6753_1642# VDD_SW[5] 5.3e-19
C2927 a_12988_212# a_15380_212# 1.9e-21
C2928 a_7369_627# VDD_SW[4] 1.85e-20
C2929 x30.A x9.A1 0.00323f
C2930 a_473_993# m1_95_2154# 1.86e-20
C2931 a_647_601# m1_95_1942# 3.42e-20
C2932 a_2468_1467# a_2566_n88# 6.87e-20
C2933 D[2] a_12638_220# 2.03e-20
C2934 x9.A1 D[6] 0.268f
C2935 VDD_SW[1] m1_95_2154# 0.0325f
C2936 a_1503_1642# D[7] 0.0682f
C2937 D[6] a_4338_n62# 0.158f
C2938 x9.A1 a_5002_1642# 8.62e-19
C2939 a_9761_627# a_12153_627# 2.94e-19
C2940 VDD a_2468_1467# 0.145f
C2941 x9.A1 VSS_SW[3] 0.113f
C2942 a_7203_627# a_7254_90# 6.13e-19
C2943 check[3] a_8679_1642# 0.257f
C2944 x2.X a_1415_895# 0.148f
C2945 a_6285_122# VSS_SW_b[4] 1.09e-20
C2946 a_6730_n62# VSS_SW[4] 6.09e-20
C2947 x10.X a_3648_993# 2.81e-19
C2948 x9.A1 m1_95_1942# 6.52f
C2949 x9.A1 a_1685_1642# 5.26e-19
C2950 a_12901_601# m1_95_1942# 4.12e-20
C2951 a_941_601# VDD_SW[7] 1.75e-19
C2952 a_1256_993# a_1555_627# 0.0256f
C2953 D[2] m1_95_2154# 0.0344f
C2954 a_193_627# a_791_627# 6.04e-20
C2955 a_941_601# a_891_909# 1.21e-20
C2956 VDD_SW_b[2] a_13906_n62# 0.0144f
C2957 a_4860_1467# VSS_SW[5] 0.0274f
C2958 a_11987_627# a_14545_627# 1.2e-20
C2959 a_12153_627# a_14379_627# 1.58e-20
C2960 a_12465_1289# a_12607_601# 8.76e-20
C2961 a_12153_627# VDD_SW_b[2] 0.0022f
C2962 x11.X m1_95_2154# 1.32e-20
C2963 a_13216_993# a_13300_993# 0.00857f
C2964 x2.X a_3356_n62# 3.67e-20
C2965 a_2419_627# a_5165_627# 4.46e-21
C2966 x30.A a_5323_2457# 0.619f
C2967 a_11546_1315# D[3] 0.0012f
C2968 a_3421_n88# a_5271_n62# 4.56e-21
C2969 a_4689_2457# x2.X 0.00106f
C2970 a_3420_212# a_5504_106# 5.86e-20
C2971 a_4413_2457# a_4689_2457# 0.00202f
C2972 x2.X a_11514_n62# 1.83e-19
C2973 x2.X a_10125_993# 5.31e-19
C2974 x2.X VDD_SW_b[7] 7.26e-19
C2975 a_505_1289# m1_95_1942# 2.26e-19
C2976 a_1503_1642# m1_95_2154# 1.04e-19
C2977 VSS_SW[2] a_12447_n62# 3.44e-19
C2978 a_2585_627# a_2879_n62# 2.38e-19
C2979 a_3039_601# a_2566_n88# 4.37e-19
C2980 VDD a_6017_n88# 0.504f
C2981 x2.X a_6285_1642# 0.00651f
C2982 a_6040_993# m1_95_1942# 5.78e-21
C2983 a_14379_627# a_15767_895# 0.0321f
C2984 D[1] a_15293_601# 0.0189f
C2985 a_1672_909# VDD_SW[7] 2.12e-20
C2986 a_11069_122# VSS_SW[2] 6.75e-20
C2987 VSS_SW_b[3] a_10937_n62# 5.35e-19
C2988 check[1] x17.X 0.00967f
C2989 x2.X check[5] 0.16f
C2990 a_5323_2457# m1_95_1942# 0.00139f
C2991 VDD a_3039_601# 0.353f
C2992 a_10983_895# a_10597_n88# 6.35e-19
C2993 a_10824_993# a_10596_212# 8.94e-21
C2994 a_10509_601# a_10801_n88# 0.00251f
C2995 a_4413_2457# check[5] 8.52e-19
C2996 D[3] a_10597_n88# 0.159f
C2997 x13.X D[4] 0.0851f
C2998 VDD a_11015_220# 0.00986f
C2999 x12.X a_7557_627# 6.12e-19
C3000 x2.X a_5675_909# 0.00137f
C3001 x9.A1 a_5725_601# 9.33e-19
C3002 check[3] a_8409_n88# 1.55e-20
C3003 a_14430_90# a_14839_n62# 4.24e-20
C3004 VSS_SW[3] a_9742_n88# 0.00683f
C3005 x2.X a_12751_627# 0.0388f
C3006 a_4689_2457# a_4977_627# 1.38e-20
C3007 a_3535_n62# a_3761_n62# 3.34e-19
C3008 x7.X a_1029_n88# 0.019f
C3009 check[1] a_12134_n88# 5.26e-19
C3010 a_4689_2457# VSS_SW[5] 0.0227f
C3011 a_7252_1467# check[3] 0.318f
C3012 VDD_SW[3] a_12433_993# 7.03e-20
C3013 check[6] a_1501_122# 6.43e-20
C3014 VDD a_6339_627# 0.0135f
C3015 check[2] a_11123_627# 2.62e-19
C3016 a_15243_909# VDD_SW_b[1] 3.6e-21
C3017 ready a_3807_895# 2.44e-19
C3018 check[4] VSS_SW_b[5] 2.08e-20
C3019 reset ready 0.0713f
C3020 x3.A x3.X 4.66e-19
C3021 x15.X a_10288_106# 1.89e-20
C3022 check[3] x14.X 5.82e-19
C3023 x9.A1 VDD_SW[4] 0.0329f
C3024 a_13715_1642# m1_95_1942# 1.97e-19
C3025 VDD a_13072_909# 0.0164f
C3026 x2.X a_78_90# 0.00367f
C3027 VDD a_2973_627# 9.86e-19
C3028 a_14733_627# a_14526_n88# 3.32e-19
C3029 check[5] VSS_SW[5] 1.43e-19
C3030 a_15293_601# a_15380_212# 6.03e-19
C3031 a_14857_1289# a_14839_n62# 3.44e-19
C3032 a_15608_993# a_14839_n62# 3.59e-19
C3033 x2.X VDD_SW_b[1] 6.63e-19
C3034 a_1029_n88# a_3420_212# 8.02e-22
C3035 a_1028_212# a_3421_n88# 5.48e-21
C3036 x2.X x20.X 1.55e-19
C3037 D[7] a_2585_627# 7.7e-21
C3038 a_5257_993# a_5165_627# 0.0369f
C3039 a_5725_601# a_6040_993# 0.13f
C3040 a_4977_627# a_5675_909# 0.00276f
C3041 a_5431_601# a_5341_993# 6.69e-20
C3042 x18.X a_12153_627# 6.35e-20
C3043 VDD VSS_SW_b[7] 0.133f
C3044 a_381_627# VSS_SW[7] 0.00595f
C3045 a_5323_2457# a_5725_601# 4.01e-19
C3046 VDD a_15511_627# 0.007f
C3047 check[4] VDD_SW[5] 0.0039f
C3048 ready VDD_SW_b[6] 1.5e-20
C3049 a_2468_1467# VDD_SW[7] 0.00487f
C3050 D[6] a_5812_212# 2.89e-20
C3051 x2.X a_11123_627# 0.0151f
C3052 a_12988_212# VSS_SW_b[2] 0.00119f
C3053 a_12989_n88# a_13461_122# 0.15f
C3054 VSS_SW[2] a_13126_304# 1.97e-20
C3055 VDD_SW[5] a_8432_993# 1.08e-20
C3056 x2.X x12.X 3.64e-19
C3057 a_7203_627# a_8205_n88# 1.06e-19
C3058 D[4] a_8204_212# 0.158f
C3059 VSS_SW[4] a_8204_212# 5.9e-22
C3060 VDD_SW_b[3] a_11514_n62# 0.0145f
C3061 a_2419_627# a_2585_627# 0.786f
C3062 a_4149_1315# D[6] 0.00195f
C3063 a_5812_212# m1_95_1942# 6.77e-21
C3064 a_9761_627# a_10359_627# 6.04e-20
C3065 a_4811_627# D[4] 1.19e-20
C3066 D[5] a_7203_627# 9.94e-20
C3067 a_6199_895# VDD_SW_b[5] 0.129f
C3068 a_9595_627# a_10459_909# 2.46e-19
C3069 a_4811_627# VSS_SW[4] 4.66e-21
C3070 a_5289_1289# x11.X 1.7e-20
C3071 check[3] a_8591_895# 0.00206f
C3072 a_9595_627# VSS_SW[3] 0.0577f
C3073 a_2585_627# m1_95_2154# 2.61e-20
C3074 a_12036_1467# VDD_SW[3] 0.00487f
C3075 D[7] a_1501_122# 0.00928f
C3076 a_8117_601# a_10509_601# 1.08e-20
C3077 a_27_627# VSS_SW_b[7] 3.11e-20
C3078 a_4528_627# a_4811_627# 0.0011f
C3079 x2.X a_6285_122# 0.0043f
C3080 a_10983_895# m1_95_2154# 5.86e-20
C3081 D[2] a_13300_993# 2.53e-19
C3082 a_11987_627# a_12751_627# 0.00134f
C3083 a_4862_90# a_4958_n88# 0.0967f
C3084 a_9595_627# m1_95_1942# 5.19e-20
C3085 D[3] m1_95_2154# 0.0344f
C3086 VSS_SW_b[6] a_4137_n62# 6.94e-20
C3087 x9.A1 a_10073_1289# 0.104f
C3088 a_16024_909# VDD_SW[1] 2.12e-20
C3089 x20.X a_16109_1315# 1.98e-19
C3090 x12.X a_4977_627# 6.35e-20
C3091 a_3895_1642# m1_95_2154# 1.04e-19
C3092 x2.X a_2865_993# 0.15f
C3093 x11.X a_4958_n88# 1.53e-21
C3094 a_2419_627# a_3183_627# 0.00134f
C3095 VDD a_7254_90# 0.189f
C3096 D[6] a_3732_993# 2.53e-19
C3097 VDD VDD_SW[2] 0.511f
C3098 a_1757_1642# a_941_601# 7.12e-21
C3099 a_6920_627# m1_95_2154# 1.66e-20
C3100 VDD_SW[7] a_3039_601# 7.64e-20
C3101 a_14999_601# a_14945_n62# 1.07e-20
C3102 a_14933_627# VSS_SW[1] 3.79e-19
C3103 a_941_601# a_2773_627# 2.34e-20
C3104 a_1415_895# a_3648_993# 1.86e-21
C3105 x9.X a_3112_106# 2.38e-20
C3106 a_13515_627# a_13323_627# 4.19e-20
C3107 VDD_SW_b[2] a_14379_627# 5.97e-19
C3108 a_13936_1315# D[2] 0.0012f
C3109 a_14096_627# VDD_SW[2] 0.0729f
C3110 a_10596_212# a_10734_304# 1.09e-19
C3111 check[3] VDD_SW_b[4] 0.0021f
C3112 x2.X a_6147_627# 0.00111f
C3113 a_6040_993# a_5271_n62# 3.59e-19
C3114 a_5725_601# a_5812_212# 6.03e-19
C3115 a_5165_627# a_4958_n88# 3.32e-19
C3116 VSS_SW[5] a_6285_122# 2.79e-21
C3117 a_473_993# a_720_106# 4.96e-20
C3118 a_193_627# a_1029_n88# 1.27e-19
C3119 a_647_601# a_1028_212# 4.51e-19
C3120 a_941_601# a_487_n62# 3.74e-20
C3121 x7.X a_2470_90# 0.0273f
C3122 a_13461_122# a_13906_n62# 0.0369f
C3123 x2.X a_3551_627# 0.00702f
C3124 x9.A1 a_12988_212# 6.23e-21
C3125 a_13216_993# a_12447_n62# 3.59e-19
C3126 a_12341_627# a_12134_n88# 3.32e-19
C3127 a_12901_601# a_12988_212# 6.03e-19
C3128 a_3947_627# a_3625_n88# 7.32e-20
C3129 a_11123_627# a_11987_627# 1.09e-19
C3130 a_11704_627# D[2] 4.42e-19
C3131 a_7203_627# a_8117_601# 0.14f
C3132 D[4] a_7649_993# 0.00874f
C3133 a_7649_993# VSS_SW[4] 0.00299f
C3134 a_7350_n88# a_7663_n62# 0.245f
C3135 a_6730_n62# a_6529_n62# 3.81e-19
C3136 x9.A1 a_1028_212# 1.41e-20
C3137 x14.X a_10215_601# 2.39e-20
C3138 check[2] VSS_SW_b[3] 3.18e-20
C3139 a_2468_1467# a_2610_1642# 0.00557f
C3140 a_2470_90# a_3420_212# 2.02e-20
C3141 a_1166_304# VSS_SW_b[6] 9.89e-21
C3142 a_1946_n62# a_3421_n88# 3.67e-21
C3143 a_10073_1289# a_9742_n88# 5.67e-21
C3144 a_14379_627# a_15072_106# 3.88e-21
C3145 D[1] a_14839_n62# 0.00257f
C3146 VDD_SW_b[5] a_5504_106# 5.26e-19
C3147 check[5] a_3648_993# 3.41e-19
C3148 VDD_SW[4] a_9595_627# 0.0865f
C3149 VDD a_1143_n62# 0.00521f
C3150 VDD_SW_b[7] a_174_n88# 3.21e-19
C3151 a_9644_1467# a_10103_1642# 6.64e-19
C3152 a_7681_1289# a_7896_106# 5.3e-21
C3153 x16.X a_12433_993# 1.03e-19
C3154 VDD_SW_b[6] a_3535_n62# 5.2e-19
C3155 a_6760_1315# D[5] 0.00121f
C3156 D[4] a_10596_212# 2.89e-20
C3157 D[4] a_8335_627# 6.12e-19
C3158 x2.X a_12680_106# 0.0385f
C3159 D[4] a_8921_304# 8.28e-19
C3160 a_8409_n88# VSS_SW_b[4] 9.21e-19
C3161 VDD x17.X 0.495f
C3162 x2.X VSS_SW_b[3] 0.0279f
C3163 VDD_SW_b[1] a_15853_122# 0.00443f
C3164 x20.X a_15853_122# 2.61e-19
C3165 a_12038_90# VSS_SW[2] 0.082f
C3166 a_76_1467# a_78_90# 1e-19
C3167 a_5575_627# a_6147_627# 2.46e-21
C3168 a_7252_1467# VSS_SW_b[4] 1.4e-19
C3169 x18.X a_14379_627# 0.236f
C3170 check[0] VDD_SW[2] 4.27e-19
C3171 a_10215_601# a_10680_909# 9.46e-19
C3172 a_13461_1642# x18.X 9.44e-21
C3173 x18.X VDD_SW_b[2] 7.23e-19
C3174 x17.X a_14096_627# 0.0338f
C3175 D[3] a_11313_304# 8.39e-19
C3176 VDD a_12134_n88# 0.712f
C3177 x9.X D[6] 0.0847f
C3178 reset VSS_SW[7] 0.0145f
C3179 a_14839_n62# a_15380_212# 0.138f
C3180 a_14526_n88# a_15381_n88# 0.0477f
C3181 check[4] a_6753_1642# 0.00688f
C3182 a_10041_993# VSS_SW[3] 0.00296f
C3183 a_1757_1642# a_2468_1467# 0.00963f
C3184 VDD_SW_b[6] a_5896_909# 2.96e-21
C3185 x2.X a_5377_n62# 5.57e-20
C3186 VSS_SW[2] m1_95_1942# 0.033f
C3187 VDD a_10801_n88# 0.48f
C3188 a_4958_n88# a_5813_n88# 0.0477f
C3189 a_5271_n62# a_5812_212# 0.138f
C3190 a_8432_993# a_9761_627# 3.24e-21
C3191 a_10041_993# m1_95_1942# 2.74e-20
C3192 VDD x10.X 0.34f
C3193 a_78_90# a_174_n88# 0.0967f
C3194 a_8204_212# a_10597_n88# 5.48e-21
C3195 a_12153_627# a_12433_993# 0.15f
C3196 x9.X m1_95_1942# 2.51e-20
C3197 a_12541_627# VSS_SW[2] 3.8e-19
C3198 x7.X a_1757_1315# 2.09e-19
C3199 VDD a_8205_n88# 0.703f
C3200 x9.A1 a_7394_1642# 9.48e-19
C3201 check[5] a_2897_1289# 0.251f
C3202 a_8679_1642# check[2] 8.62e-21
C3203 a_7369_627# a_7350_n88# 4.91e-19
C3204 VDD D[5] 1.27f
C3205 a_10073_1289# a_9595_627# 0.00104f
C3206 D[1] a_15518_304# 9.65e-19
C3207 a_12036_1467# x16.X 0.0876f
C3208 x9.A1 a_15293_601# 0.00103f
C3209 a_12901_601# a_15293_601# 9.37e-21
C3210 x13.X m1_95_2154# 1.03e-20
C3211 a_12153_627# a_14733_627# 3.67e-21
C3212 a_13375_895# a_14825_993# 8e-21
C3213 VDD_SW_b[4] a_8921_n62# 5.22e-19
C3214 VDD_SW_b[4] a_10215_601# 2.46e-20
C3215 a_7681_1289# a_7823_601# 8.76e-20
C3216 x2.X a_13407_220# 9.61e-19
C3217 a_12680_106# a_12924_n62# 0.00707f
C3218 a_12447_n62# a_13103_n62# 3.73e-19
C3219 a_7967_627# a_7350_n88# 1.08e-19
C3220 a_8432_993# a_8677_122# 1.51e-20
C3221 D[2] a_12447_n62# 0.00257f
C3222 a_11987_627# a_12680_106# 3.88e-21
C3223 VDD_SW_b[1] a_15316_n62# 8.09e-20
C3224 x2.X a_8679_1642# 0.00649f
C3225 a_3333_601# a_3807_895# 0.265f
C3226 a_2585_627# a_2949_993# 0.0018f
C3227 x9.A1 a_1946_n62# 1.9e-20
C3228 a_3039_601# a_2773_627# 8.07e-20
C3229 x9.X a_5725_601# 4.04e-21
C3230 a_2566_n88# VSS_SW_b[6] 0.135f
C3231 a_3112_106# a_3625_n88# 0.00189f
C3232 a_2879_n62# a_3893_122# 0.0633f
C3233 a_3420_212# a_3421_n88# 0.785f
C3234 a_14999_601# a_15464_909# 9.46e-19
C3235 a_15855_1642# a_15767_895# 5.45e-19
C3236 a_10983_895# a_11704_627# 0.0967f
C3237 a_10509_601# a_11123_627# 0.0526f
C3238 a_10215_601# VDD_SW[3] 2.07e-20
C3239 x17.X check[0] 5.47e-19
C3240 D[3] a_11704_627# 0.00234f
C3241 VDD a_12937_304# 0.00268f
C3242 a_15380_212# a_15518_304# 1.09e-19
C3243 VDD a_939_2457# 1.49f
C3244 VDD VSS_SW_b[6] 0.129f
C3245 a_305_2457# a_193_627# 8.93e-22
C3246 VDD_SW[4] a_10041_993# 7.03e-20
C3247 x2.X a_14825_993# 0.15f
C3248 x3.X m1_95_1942# 4.93e-19
C3249 VDD_SW[6] a_6199_895# 1.27e-20
C3250 x9.A1 a_8933_1642# 0.195f
C3251 VDD_SW_b[6] VSS_SW_b[5] 0.0323f
C3252 VDD_SW_b[2] a_13461_122# 0.00445f
C3253 a_13461_1642# a_13461_122# 1.57e-21
C3254 VDD a_4363_1642# 0.00177f
C3255 VDD a_8117_601# 0.519f
C3256 a_11539_1642# VDD_SW[3] 5.44e-19
C3257 a_8205_n88# a_8319_n62# 2.14e-20
C3258 a_8204_212# a_8545_n62# 0.00134f
C3259 a_7896_106# VSS_SW[3] 9.06e-21
C3260 a_3648_993# a_3551_627# 0.00386f
C3261 a_3807_895# a_4064_909# 0.00869f
C3262 x14.X check[2] 0.00901f
C3263 a_2419_627# a_4811_627# 1.63e-20
C3264 a_3333_601# VDD_SW_b[6] 0.00635f
C3265 a_2773_627# a_2973_627# 3.81e-19
C3266 x12.X a_7615_1315# 2.41e-19
C3267 VDD a_14545_627# 0.746f
C3268 a_7896_106# m1_95_1942# 4.96e-22
C3269 a_4811_627# m1_95_2154# 3.53e-20
C3270 a_10288_106# a_12134_n88# 1.86e-21
C3271 a_14096_627# a_14545_627# 5.39e-19
C3272 a_939_2457# a_27_627# 1.42e-20
C3273 x2.X a_8409_n88# 0.00368f
C3274 x9.A1 a_7350_n88# 7.35e-19
C3275 a_5812_212# a_5950_304# 1.09e-19
C3276 a_2897_1289# a_2865_993# 4.54e-19
C3277 a_10288_106# a_10801_n88# 0.00189f
C3278 a_10055_n62# a_11069_122# 0.0633f
C3279 a_10596_212# a_10597_n88# 0.784f
C3280 VSS_SW[7] a_977_304# 8.35e-20
C3281 a_1028_212# a_1233_n88# 0.15f
C3282 a_487_n62# VSS_SW_b[7] 0.0142f
C3283 x2.X a_7252_1467# 2.92e-19
C3284 x12.X a_7203_627# 0.236f
C3285 check[3] VDD_SW[5] 4.37e-19
C3286 a_12989_n88# a_15381_n88# 1.33e-19
C3287 VDD a_8848_909# 0.00609f
C3288 a_12447_n62# VSS_SW_b[1] 1.09e-20
C3289 VDD a_9122_n62# 0.112f
C3290 a_4064_909# VDD_SW_b[6] 3.4e-20
C3291 a_8205_n88# a_10288_106# 1.67e-21
C3292 D[2] a_13126_304# 9.67e-19
C3293 a_7823_601# a_8288_909# 9.46e-19
C3294 x2.X x14.X 3.4e-19
C3295 check[6] a_941_601# 2.14e-19
C3296 a_15767_895# a_16488_627# 0.0967f
C3297 a_14999_601# VDD_SW[1] 2.07e-20
C3298 a_15293_601# a_15907_627# 0.0526f
C3299 x9.A1 a_6467_1642# 5.26e-19
C3300 x10.X a_5431_601# 2.7e-20
C3301 D[6] a_3625_n88# 0.00546f
C3302 a_10073_1289# a_10041_993# 4.54e-19
C3303 VDD a_4860_1467# 0.115f
C3304 x9.X a_5271_n62# 4.43e-20
C3305 check[3] a_7711_1642# 0.00526f
C3306 x9.A1 a_439_1315# 0.00504f
C3307 VSS_SW[1] m1_95_2154# 0.0337f
C3308 a_13216_993# m1_95_1942# 5.78e-21
C3309 a_6285_122# a_6153_n62# 0.025f
C3310 x9.A1 x7.X 6.79e-19
C3311 VSS_SW_b[5] a_5927_n62# 5.23e-19
C3312 a_6017_n88# VSS_SW[4] 8.81e-20
C3313 a_4811_627# a_5257_993# 0.159f
C3314 D[5] a_5431_601# 0.00583f
C3315 x9.A1 a_12465_1289# 0.104f
C3316 a_12901_601# a_13632_909# 0.0016f
C3317 a_12433_993# VDD_SW_b[2] 3.93e-21
C3318 VDD a_1415_895# 0.672f
C3319 ready x2.X 0.437f
C3320 x27.A x30.A 4.66e-19
C3321 x9.A1 a_3420_212# 1.26e-20
C3322 a_2879_n62# a_2985_n62# 0.0526f
C3323 a_3625_n88# a_3839_220# 0.0104f
C3324 ready a_4413_2457# 0.202f
C3325 a_7823_601# m1_95_1942# 3.42e-20
C3326 a_3420_212# a_4338_n62# 0.0453f
C3327 a_7649_993# m1_95_2154# 1.86e-20
C3328 a_3421_n88# a_4137_304# 0.0018f
C3329 x2.X a_10680_909# 0.00309f
C3330 x27.A D[6] 0.00836f
C3331 VSS_SW[2] a_12988_212# 1.18e-21
C3332 a_505_1289# x7.X 1.75e-20
C3333 a_939_2457# VDD_SW[7] 0.0315f
C3334 x2.X a_5319_1642# 2.62e-19
C3335 a_14857_1289# D[1] 0.0662f
C3336 D[1] a_15608_993# 0.00606f
C3337 a_14379_627# a_14733_627# 0.0455f
C3338 check[0] a_14545_627# 5.41e-19
C3339 VDD_SW_b[7] a_2566_n88# 5.91e-19
C3340 D[3] a_12447_n62# 3.12e-21
C3341 VDD a_3356_n62# 8.23e-19
C3342 x14.X a_9312_627# 0.0285f
C3343 a_3895_1642# a_3947_627# 1.92e-20
C3344 VDD_SW_b[2] a_14733_627# 9.33e-21
C3345 check[2] a_9646_90# 2.5e-20
C3346 VDD a_4689_2457# 0.387f
C3347 x2.X a_8591_895# 0.148f
C3348 a_10983_895# a_11069_122# 4.53e-22
C3349 a_10824_993# a_10801_n88# 1.86e-19
C3350 a_4811_627# a_5943_627# 0.00272f
C3351 x15.X a_11546_1315# 0.00143f
C3352 x27.A m1_95_1942# 8.75e-20
C3353 D[3] a_11069_122# 0.00933f
C3354 VDD a_10125_993# 0.00421f
C3355 VDD a_11514_n62# 0.113f
C3356 VDD VDD_SW_b[7] 0.156f
C3357 x8.X D[6] 0.00886f
C3358 a_14430_90# a_15380_212# 2.02e-20
C3359 a_13906_n62# a_15381_n88# 3.67e-21
C3360 check[5] a_2566_n88# 5.27e-19
C3361 a_12988_212# a_14945_n62# 1.09e-19
C3362 a_13126_304# VSS_SW_b[1] 9.89e-21
C3363 VDD a_6285_1642# 0.225f
C3364 x2.X a_13119_627# 0.00702f
C3365 a_27_627# a_1415_895# 0.0321f
C3366 D[7] a_941_601# 0.019f
C3367 VDD_SW_b[4] a_8140_n62# 8.1e-20
C3368 a_8623_220# VSS_SW[3] 1.57e-20
C3369 a_3504_909# VDD_SW[6] 2.82e-20
C3370 check[1] a_12680_106# 8.64e-22
C3371 a_9644_1467# check[3] 1.56e-19
C3372 VDD_SW[3] a_13375_895# 1.27e-20
C3373 VDD check[5] 1.91f
C3374 ready VSS_SW[5] 2e-19
C3375 a_6539_1642# x11.X 0.0845f
C3376 check[2] VDD_SW[3] 0.00394f
C3377 x8.X m1_95_1942# 1.18e-19
C3378 x16.X a_10215_601# 1.98e-20
C3379 x15.X a_10597_n88# 0.0189f
C3380 VDD a_5675_909# 0.0125f
C3381 a_5289_1289# a_4811_627# 0.00104f
C3382 a_16109_1642# m1_95_1942# 1.97e-19
C3383 x12.X a_6760_1315# 4.97e-20
C3384 VDD a_12751_627# 0.00141f
C3385 a_6199_895# a_7369_627# 2.8e-19
C3386 a_5725_601# a_7823_601# 1.55e-20
C3387 x2.X VDD_SW_b[4] 7.37e-19
C3388 a_15608_993# a_15380_212# 8.94e-21
C3389 x2.X a_9646_90# 0.00368f
C3390 a_15767_895# a_15381_n88# 6.35e-19
C3391 a_15293_601# a_15585_n88# 0.00251f
C3392 a_5812_212# a_7350_n88# 6.19e-19
C3393 a_2468_1467# check[6] 1.54e-19
C3394 a_941_601# a_2419_627# 3.79e-19
C3395 a_1029_n88# a_2470_90# 5.39e-19
C3396 a_487_n62# a_1143_n62# 3.73e-19
C3397 a_720_106# a_964_n62# 0.00707f
C3398 a_1233_n88# a_1946_n62# 8.07e-20
C3399 VSS_SW_b[7] a_1447_220# 1.12e-20
C3400 a_1501_122# a_1745_304# 0.00972f
C3401 x18.X a_12433_993# 1.55e-20
C3402 a_12851_909# VDD_SW[2] 1.01e-20
C3403 D[7] a_1672_909# 8.06e-19
C3404 a_27_627# VDD_SW_b[7] 1.09e-19
C3405 a_4811_627# a_4958_n88# 0.00176f
C3406 x2.X a_14526_n88# 0.178f
C3407 a_193_627# a_647_601# 0.117f
C3408 a_7823_601# VDD_SW[4] 2.07e-20
C3409 a_8591_895# a_9312_627# 0.0967f
C3410 a_8117_601# a_8731_627# 0.0526f
C3411 VDD a_78_90# 0.203f
C3412 VDD x20.X 0.438f
C3413 VDD VDD_SW_b[1] 0.156f
C3414 a_473_993# m1_95_1942# 2.74e-20
C3415 a_941_601# m1_95_2154# 2.82e-20
C3416 VDD_SW[1] m1_95_1942# 0.0329f
C3417 x2.X VDD_SW[3] 0.0327f
C3418 a_13193_n88# VSS_SW_b[2] 9.26e-19
C3419 D[6] a_4862_90# 8.78e-19
C3420 x6.X a_78_90# 0.00259f
C3421 x2.X a_2136_627# 4.01e-19
C3422 a_14379_627# a_16488_627# 1.75e-19
C3423 VDD_SW_b[5] a_7369_627# 0.00336f
C3424 a_10359_627# a_10727_627# 3.34e-19
C3425 a_10680_909# VDD_SW_b[3] 7.05e-21
C3426 x18.X a_14733_627# 6.12e-19
C3427 x18.X a_15855_1642# 1.97e-20
C3428 x9.A1 a_193_627# 1.78e-19
C3429 x2.X a_1256_993# 0.187f
C3430 a_7254_90# VSS_SW[4] 0.082f
C3431 a_9761_627# a_10727_627# 2.14e-20
C3432 a_9595_627# a_10908_993# 2.13e-19
C3433 VDD a_11123_627# 0.00162f
C3434 a_1256_993# a_1363_627# 0.00707f
C3435 a_14428_1467# a_14526_n88# 6.87e-20
C3436 a_1415_895# VDD_SW[7] 0.00356f
C3437 D[2] m1_95_1942# 0.0335f
C3438 VDD x12.X 0.341f
C3439 a_647_601# a_791_627# 0.0697f
C3440 a_941_601# a_1112_909# 0.00652f
C3441 VDD_SW_b[4] a_9312_627# 0.186f
C3442 x11.X m1_95_1942# 2.53e-20
C3443 a_11987_627# a_13119_627# 0.00272f
C3444 x9.A1 a_9786_1642# 8.64e-19
C3445 a_27_627# a_78_90# 6.13e-19
C3446 x9.A1 a_4137_304# 6.9e-21
C3447 check[2] a_11071_1642# 0.257f
C3448 a_3420_212# a_5812_212# 9.5e-22
C3449 a_3893_122# a_4958_n88# 8e-21
C3450 a_4137_304# a_4338_n62# 8.99e-19
C3451 a_3421_n88# a_5504_106# 1.67e-21
C3452 a_505_1289# a_193_627# 0.00323f
C3453 a_9786_1315# VSS_SW[3] 7.95e-19
C3454 a_1503_1642# m1_95_1942# 2.26e-19
C3455 a_2865_993# a_2566_n88# 8.71e-20
C3456 VDD a_6285_122# 0.332f
C3457 a_2468_1467# D[7] 2.91e-19
C3458 a_3039_601# a_2879_n62# 0.0026f
C3459 a_15767_895# a_16298_n62# 4.06e-19
C3460 VDD_SW_b[7] VDD_SW[7] 3.64e-19
C3461 x15.X m1_95_2154# 1.32e-20
C3462 a_891_909# VDD_SW_b[7] 2.4e-21
C3463 a_10055_n62# a_12038_90# 3.67e-21
C3464 VSS_SW_b[3] a_10246_220# 5.34e-20
C3465 a_10596_212# a_11313_304# 4.45e-20
C3466 a_9742_n88# a_10161_n62# 0.0383f
C3467 VDD a_2865_993# 0.222f
C3468 a_10597_n88# a_11015_220# 0.00276f
C3469 a_10801_n88# a_10734_304# 9.46e-19
C3470 x2.X a_15329_304# 0.00168f
C3471 x9.A1 a_6199_895# 2.41e-19
C3472 check[5] VDD_SW[7] 4.38e-19
C3473 x2.X a_5896_909# 0.00309f
C3474 VSS_SW[3] a_10055_n62# 3.44e-19
C3475 check[3] a_8677_122# 2.04e-20
C3476 ready a_76_1467# 3.18e-21
C3477 a_939_2457# a_1757_1642# 0.0012f
C3478 x7.X a_1233_n88# 1.81e-19
C3479 x9.A1 a_13193_n88# 3.88e-20
C3480 x2.X a_11071_1642# 0.00647f
C3481 a_13216_993# a_12988_212# 8.94e-21
C3482 a_2468_1467# a_2419_627# 5.32e-19
C3483 a_13375_895# a_12989_n88# 6.35e-19
C3484 a_12901_601# a_13193_n88# 0.00251f
C3485 check[6] VSS_SW_b[7] 9.18e-21
C3486 x11.X a_5725_601# 1.29e-19
C3487 VDD a_6147_627# 0.00101f
C3488 VDD_SW[3] a_11987_627# 0.0865f
C3489 a_2773_627# VSS_SW_b[6] 2.36e-19
C3490 a_939_2457# a_2773_627# 1.54e-21
C3491 VDD_SW_b[3] VDD_SW[3] 3.63e-19
C3492 x18.X a_14570_1315# 8.21e-19
C3493 check[0] x20.X 0.00965f
C3494 check[0] VDD_SW_b[1] 0.00207f
C3495 x14.X a_10509_601# 4.89e-20
C3496 a_2468_1467# m1_95_2154# 8.35e-20
C3497 x2.X VSS_SW[7] 0.0768f
C3498 VDD a_3551_627# 0.00717f
C3499 a_6539_1642# a_6920_627# 5.84e-19
C3500 a_1029_n88# a_3421_n88# 1.33e-19
C3501 a_487_n62# VSS_SW_b[6] 1.09e-20
C3502 a_14379_627# a_15381_n88# 1.06e-19
C3503 D[1] a_15380_212# 0.157f
C3504 VDD_SW_b[2] a_15381_n88# 2.44e-21
C3505 a_5257_993# a_5341_993# 0.00972f
C3506 a_6199_895# a_6040_993# 0.207f
C3507 a_4977_627# a_5896_909# 0.00907f
C3508 a_5725_601# a_5165_627# 1.15e-20
C3509 a_5431_601# a_5675_909# 0.0104f
C3510 x9.A1 VDD_SW_b[5] 1.13e-19
C3511 D[5] a_5462_220# 1.98e-20
C3512 a_11325_1642# a_11253_1642# 6.64e-19
C3513 a_5323_2457# a_6199_895# 0.00152f
C3514 check[2] x16.X 6.04e-19
C3515 D[6] a_5813_n88# 4.83e-22
C3516 x2.X a_12989_n88# 0.0207f
C3517 VDD_SW[5] a_7557_627# 6.11e-20
C3518 D[4] a_8205_n88# 0.158f
C3519 a_7203_627# a_8409_n88# 0.00204f
C3520 VSS_SW[4] a_8205_n88# 9.29e-21
C3521 a_2419_627# a_3039_601# 0.149f
C3522 D[6] a_2585_627# 0.168f
C3523 x10.X a_4528_627# 0.0285f
C3524 a_7252_1467# a_7203_627# 5.32e-19
C3525 a_10509_601# a_10680_909# 0.00652f
C3526 a_5813_n88# m1_95_1942# 1.16e-21
C3527 a_11704_627# a_10596_212# 6.63e-19
C3528 a_10215_601# a_10359_627# 0.0697f
C3529 D[5] D[4] 0.00183f
C3530 a_6040_993# VDD_SW_b[5] 5e-20
C3531 D[3] a_10459_909# 6.77e-19
C3532 D[3] a_12038_90# 8.76e-19
C3533 D[5] VSS_SW[4] 4.85e-19
C3534 VDD a_12680_106# 0.36f
C3535 check[4] check[3] 0.00525f
C3536 a_9761_627# a_10215_601# 0.117f
C3537 ready a_2897_1289# 4.05e-20
C3538 a_14526_n88# a_15853_122# 4.59e-22
C3539 a_14839_n62# a_15585_n88# 0.199f
C3540 a_15072_106# a_15381_n88# 0.0327f
C3541 x14.X a_7203_627# 0.00113f
C3542 a_3895_1642# D[6] 0.0681f
C3543 a_5323_2457# VDD_SW_b[5] 1.07e-20
C3544 a_2585_627# m1_95_1942# 3.82e-20
C3545 a_3039_601# m1_95_2154# 2.34e-20
C3546 check[3] a_8432_993# 2.28e-19
C3547 D[3] VSS_SW[3] 0.134f
C3548 VDD VSS_SW_b[3] 0.101f
C3549 D[7] VSS_SW_b[7] 5.32e-19
C3550 a_8591_895# a_10509_601# 1.54e-20
C3551 x2.X x16.X 3.45e-19
C3552 x2.X VSS_SW_b[5] 0.0278f
C3553 a_4528_627# D[5] 4.42e-19
C3554 a_3947_627# a_4811_627# 1.09e-19
C3555 a_10983_895# m1_95_1942# 8.62e-20
C3556 a_13375_895# a_13906_n62# 4.06e-19
C3557 D[3] m1_95_1942# 0.0335f
C3558 a_4862_90# a_5271_n62# 4.24e-20
C3559 x9.A1 a_12607_601# 2.81e-20
C3560 a_12465_1289# VSS_SW[2] 0.00187f
C3561 a_12153_627# a_13375_895# 0.0494f
C3562 a_12607_601# a_12901_601# 0.199f
C3563 x9.A1 a_8861_1642# 5.26e-19
C3564 check[5] a_2610_1642# 0.00688f
C3565 x12.X a_5431_601# 1.98e-20
C3566 x2.X a_3333_601# 0.119f
C3567 a_3895_1642# m1_95_1942# 2.26e-19
C3568 x11.X a_5271_n62# 0.002f
C3569 VDD a_5377_n62# 0.0139f
C3570 a_2419_627# a_2973_627# 0.00206f
C3571 a_29_2457# a_939_2457# 2.64e-19
C3572 a_7681_1289# x13.X 1.75e-20
C3573 a_6920_627# m1_95_1942# 2.45e-20
C3574 a_1757_1642# a_1415_895# 0.00232f
C3575 VDD_SW[7] a_2865_993# 7.03e-20
C3576 D[1] a_16097_304# 8.37e-19
C3577 a_1415_895# a_2773_627# 8.26e-21
C3578 x9.A1 a_14857_1289# 0.105f
C3579 x9.X a_3420_212# 0.244f
C3580 x9.A1 a_15608_993# 4.84e-21
C3581 x2.X VDD_SW[5] 0.0327f
C3582 VDD_SW_b[4] a_10509_601# 2.26e-20
C3583 a_6199_895# a_5812_212# 0.00165f
C3584 a_4977_627# VSS_SW_b[5] 4.03e-20
C3585 a_5725_601# a_5813_n88# 3.89e-19
C3586 VSS_SW[5] VSS_SW_b[5] 0.00723f
C3587 a_1415_895# a_487_n62# 0.00219f
C3588 a_193_627# a_1233_n88# 8.75e-19
C3589 a_941_601# a_720_106# 3.46e-19
C3590 a_647_601# a_1029_n88# 0.00322f
C3591 a_8677_122# a_8921_n62# 0.00807f
C3592 x2.X a_13906_n62# 1.9e-19
C3593 a_12988_212# a_13103_n62# 0.00272f
C3594 a_12447_n62# VSS_SW[1] 1.64e-20
C3595 a_3333_601# a_4977_627# 6.25e-20
C3596 x2.X a_4064_909# 4.04e-19
C3597 a_12680_106# a_13329_n62# 0.00316f
C3598 x2.X a_12153_627# 0.0537f
C3599 a_3333_601# VSS_SW[5] 2.89e-20
C3600 a_3807_895# a_3761_n62# 1.65e-20
C3601 a_3947_627# a_3893_122# 2.54e-20
C3602 a_11987_627# a_12989_n88# 1.06e-19
C3603 a_1757_1642# VDD_SW_b[7] 1.29e-19
C3604 D[2] a_12988_212# 0.158f
C3605 x2.X a_7711_1642# 2.63e-19
C3606 VDD_SW_b[1] a_15721_n62# 0.00178f
C3607 a_7203_627# a_8591_895# 0.0321f
C3608 D[4] a_8117_601# 0.0191f
C3609 VDD_SW_b[3] a_12989_n88# 2.44e-21
C3610 a_8117_601# VSS_SW[4] 2.17e-19
C3611 a_7350_n88# a_7896_106# 0.207f
C3612 a_15293_601# a_15464_909# 0.00652f
C3613 a_14999_601# a_15143_627# 0.0697f
C3614 VDD_SW_b[7] a_2773_627# 9.33e-21
C3615 a_10509_601# VDD_SW[3] 1.79e-19
C3616 a_10824_993# a_11123_627# 0.0256f
C3617 x9.A1 a_1029_n88# 8.52e-21
C3618 a_2470_90# a_3421_n88# 9.87e-21
C3619 a_10073_1289# a_10055_n62# 3.44e-19
C3620 D[3] a_10931_627# 2e-19
C3621 a_1757_1642# check[5] 1.67e-19
C3622 a_1447_220# VSS_SW_b[6] 3.96e-21
C3623 VDD a_13407_220# 0.00985f
C3624 a_15381_n88# a_15799_220# 0.00276f
C3625 a_14839_n62# a_14945_n62# 0.0526f
C3626 a_4977_627# VDD_SW[5] 1.96e-20
C3627 a_15585_n88# a_15518_304# 9.46e-19
C3628 a_15380_212# a_16097_304# 4.45e-20
C3629 a_5725_601# a_6920_627# 5.73e-19
C3630 VSS_SW_b[1] a_15030_220# 5.34e-20
C3631 VDD_SW_b[5] a_5812_212# 0.0417f
C3632 VDD_SW[4] a_10983_895# 1.27e-20
C3633 VDD a_8679_1642# 0.219f
C3634 x9.A1 a_11325_1642# 0.195f
C3635 x2.X a_15767_895# 0.148f
C3636 VDD_SW[4] D[3] 4.43e-19
C3637 VDD_SW_b[7] a_487_n62# 5.22e-19
C3638 VDD a_1369_n62# 0.0301f
C3639 a_9644_1467# check[2] 0.318f
C3640 x16.X a_11987_627# 0.236f
C3641 check[1] VDD_SW[3] 4.32e-19
C3642 VDD_SW_b[6] a_3761_n62# 0.00179f
C3643 x15.X a_11704_627# 0.0338f
C3644 x16.X VDD_SW_b[3] 7.25e-19
C3645 a_7203_627# VDD_SW_b[4] 1.15e-19
C3646 D[4] a_8848_909# 8.06e-19
C3647 a_1503_1642# a_1028_212# 1.39e-21
C3648 D[4] a_9122_n62# 0.158f
C3649 a_8677_122# VSS_SW_b[4] 7.15e-19
C3650 VDD a_14825_993# 0.218f
C3651 a_10532_n62# a_10937_n62# 2.46e-21
C3652 a_76_1467# VSS_SW[7] 0.0271f
C3653 VDD_SW[2] m1_95_2154# 0.0327f
C3654 a_16109_1642# a_15293_601# 7.12e-21
C3655 a_10596_212# a_12447_n62# 2.62e-19
C3656 a_10597_n88# a_12134_n88# 1.98e-19
C3657 a_10041_993# a_10161_n62# 6.88e-22
C3658 a_10596_212# a_11069_122# 0.159f
C3659 a_10597_n88# a_10801_n88# 0.117f
C3660 VSS_SW[3] a_10545_304# 8.35e-20
C3661 a_10288_106# VSS_SW_b[3] 0.00322f
C3662 x2.X a_5748_n62# 3.68e-20
C3663 x2.X a_9644_1467# 2.88e-19
C3664 a_5504_106# a_5812_212# 0.14f
C3665 a_5271_n62# a_5813_n88# 0.125f
C3666 a_13126_304# VSS_SW[1] 2.77e-20
C3667 a_12988_212# VSS_SW_b[1] 0.00377f
C3668 VSS_SW[7] a_174_n88# 0.00677f
C3669 a_78_90# a_487_n62# 4.24e-20
C3670 a_12607_601# a_12553_n62# 1.07e-20
C3671 a_8205_n88# a_10597_n88# 1.33e-19
C3672 D[2] a_13705_304# 8.38e-19
C3673 a_11987_627# a_12153_627# 0.786f
C3674 VDD a_8409_n88# 0.501f
C3675 VDD_SW_b[3] a_12153_627# 0.00336f
C3676 a_15608_993# a_15907_627# 0.0256f
C3677 a_15293_601# VDD_SW[1] 1.83e-19
C3678 a_7823_601# a_7350_n88# 4.37e-19
C3679 VDD a_7252_1467# 0.114f
C3680 a_7369_627# a_7663_n62# 2.38e-19
C3681 a_11071_1642# a_10509_601# 0.00263f
C3682 check[3] a_9147_1642# 0.00688f
C3683 x2.X a_678_220# 0.00279f
C3684 check[2] a_9761_627# 5.35e-19
C3685 a_10073_1289# D[3] 0.0662f
C3686 VDD x14.X 0.415f
C3687 x13.X VSS_SW[3] 0.138f
C3688 a_14999_601# VSS_SW[1] 6.23e-19
C3689 a_5431_601# a_5377_n62# 1.07e-20
C3690 x13.X m1_95_1942# 1.97e-20
C3691 x9.A1 D[1] 0.268f
C3692 a_12901_601# D[1] 8.7e-19
C3693 x9.A1 a_12178_1642# 8.64e-19
C3694 a_13375_895# a_14379_627# 6.9e-19
C3695 D[2] a_15293_601# 2.67e-21
C3696 a_939_2457# check[6] 0.0505f
C3697 a_7681_1289# a_7649_993# 4.54e-19
C3698 a_13375_895# VDD_SW_b[2] 0.128f
C3699 a_13461_1642# a_13375_895# 5.55e-19
C3700 x9.A1 VDD_SW[6] 0.0329f
C3701 a_11071_1642# check[1] 6.17e-21
C3702 a_4689_2457# a_4528_627# 4.35e-21
C3703 x2.X a_10359_627# 0.0391f
C3704 a_12134_n88# a_12638_220# 0.00869f
C3705 a_7896_106# a_8153_304# 0.00857f
C3706 a_7663_n62# a_8342_304# 0.00652f
C3707 x2.X VSS_SW[6] 0.18f
C3708 a_2865_993# a_2773_627# 0.0369f
C3709 a_3333_601# a_3648_993# 0.13f
C3710 VSS_SW[2] a_13193_n88# 9.93e-21
C3711 a_3039_601# a_2949_993# 6.69e-20
C3712 a_2585_627# a_3283_909# 0.00276f
C3713 a_2879_n62# VSS_SW_b[6] 0.0142f
C3714 x2.X a_9761_627# 0.0537f
C3715 VSS_SW[6] a_3070_220# 4.25e-19
C3716 a_3420_212# a_3625_n88# 0.15f
C3717 x17.X m1_95_2154# 1.31e-20
C3718 a_11069_122# a_11313_n62# 0.00807f
C3719 a_14379_627# a_15243_909# 2.46e-19
C3720 check[0] a_14825_993# 7.14e-20
C3721 D[1] a_14909_993# 8.12e-19
C3722 D[3] a_12988_212# 5.78e-20
C3723 VDD_SW_b[2] a_15243_909# 2.1e-21
C3724 VDD ready 0.792f
C3725 x3.X a_193_627# 5.4e-19
C3726 a_305_2457# a_647_601# 1.12e-19
C3727 x10.X a_2419_627# 0.00117f
C3728 VDD a_10680_909# 0.0164f
C3729 VDD_SW[6] a_6040_993# 1.08e-20
C3730 ready x6.X 4.55e-23
C3731 x2.X a_14379_627# 0.354f
C3732 VDD a_5319_1642# 8.63e-19
C3733 x9.A1 a_15380_212# 1.41e-20
C3734 x2.X a_13461_1642# 0.00643f
C3735 x2.X VDD_SW_b[2] 7.31e-19
C3736 x30.A a_4811_627# 2.63e-21
C3737 check[1] a_12989_n88# 7.54e-21
C3738 VDD a_8591_895# 0.721f
C3739 VDD_SW[3] a_12341_627# 6.11e-20
C3740 x15.X a_12447_n62# 4.73e-20
C3741 x10.X m1_95_2154# 6.47e-20
C3742 VDD a_1971_1642# 0.00177f
C3743 a_8204_212# VSS_SW[3] 0.0872f
C3744 a_8409_n88# a_8319_n62# 9.75e-19
C3745 a_8205_n88# a_8545_n62# 6.04e-20
C3746 a_305_2457# x9.A1 0.00214f
C3747 VSS_SW_b[4] a_7769_n62# 0.00335f
C3748 a_3807_895# VDD_SW_b[6] 0.129f
C3749 D[6] a_4811_627# 9.98e-20
C3750 a_2419_627# D[5] 1.19e-20
C3751 x7.X x8.X 0.11f
C3752 x16.X a_10509_601# 0.00124f
C3753 x15.X a_11069_122# 2.61e-19
C3754 a_8204_212# m1_95_1942# 6.77e-21
C3755 VDD a_13119_627# 6.2e-19
C3756 x13.X VDD_SW[4] 0.176f
C3757 a_15767_895# a_15853_122# 4.53e-22
C3758 a_15608_993# a_15585_n88# 1.86e-19
C3759 a_13715_1642# D[1] 1.62e-19
C3760 D[5] m1_95_2154# 0.0344f
C3761 a_14428_1467# a_14379_627# 5.32e-19
C3762 a_4811_627# m1_95_1942# 5.19e-20
C3763 a_12036_1467# a_12495_1642# 6.64e-19
C3764 ready a_27_627# 1.42e-21
C3765 a_8679_1642# a_8731_627# 1.92e-20
C3766 a_939_2457# D[7] 0.0344f
C3767 D[7] VSS_SW_b[6] 2.02e-19
C3768 x2.X a_8677_122# 0.00429f
C3769 a_5812_212# a_6231_220# 2.46e-19
C3770 x18.X a_13375_895# 0.00863f
C3771 a_5813_n88# a_5950_304# 0.00907f
C3772 a_5271_n62# a_6730_n62# 3.79e-20
C3773 a_12751_627# a_13323_627# 2.46e-21
C3774 x16.X check[1] 0.00902f
C3775 a_9312_627# a_9761_627# 5.39e-19
C3776 VSS_SW[7] a_1166_304# 1.97e-20
C3777 a_1029_n88# a_1233_n88# 0.117f
C3778 a_305_2457# a_505_1289# 0.00165f
C3779 a_720_106# VSS_SW_b[7] 0.00322f
C3780 a_1028_212# a_1501_122# 0.159f
C3781 x14.X a_10007_1315# 2.35e-19
C3782 x12.X D[4] 0.00875f
C3783 VDD VDD_SW_b[4] 0.218f
C3784 a_9122_n62# a_10597_n88# 3.67e-21
C3785 x2.X a_15072_106# 0.0385f
C3786 x11.X a_7350_n88# 0.00864f
C3787 x12.X VSS_SW[4] 0.253f
C3788 VDD a_9646_90# 0.196f
C3789 check[6] a_1415_895# 0.00271f
C3790 a_7369_627# a_7967_627# 6.04e-20
C3791 a_8117_601# a_8067_909# 1.21e-20
C3792 a_12607_601# VSS_SW[2] 6.25e-19
C3793 x10.X a_5257_993# 1.03e-19
C3794 a_4149_1642# x10.X 7.97e-19
C3795 a_14791_1315# D[1] 0.00202f
C3796 D[1] a_15907_627# 0.0043f
C3797 a_939_2457# a_2419_627# 2.48e-19
C3798 D[6] a_3893_122# 0.00928f
C3799 a_10509_601# a_12153_627# 6.25e-20
C3800 a_2419_627# VSS_SW_b[6] 7.68e-20
C3801 VDD a_14526_n88# 0.723f
C3802 a_9761_627# a_11987_627# 1.36e-20
C3803 x9.A1 a_1757_1315# 0.00499f
C3804 a_9761_627# VDD_SW_b[3] 0.00226f
C3805 VSS_SW[1] m1_95_1942# 0.0329f
C3806 a_9595_627# a_10149_627# 0.00206f
C3807 VDD VDD_SW[3] 0.603f
C3808 VSS_SW_b[5] a_6153_n62# 5.34e-19
C3809 a_6285_122# VSS_SW[4] 6.66e-20
C3810 x9.A1 a_16097_304# 8.15e-21
C3811 VDD a_2136_627# 0.194f
C3812 x2.X x18.X 3.35e-19
C3813 a_939_2457# m1_95_2154# 0.00298f
C3814 a_4149_1642# D[5] 1.74e-19
C3815 D[5] a_5257_993# 0.00874f
C3816 a_4811_627# a_5725_601# 0.14f
C3817 VDD_SW_b[2] a_12924_n62# 8.1e-20
C3818 a_11987_627# a_14379_627# 1.74e-20
C3819 VDD a_1256_993# 0.189f
C3820 x9.A1 a_11253_1642# 5.26e-19
C3821 check[1] a_12153_627# 5.41e-19
C3822 a_11987_627# VDD_SW_b[2] 1.09e-19
C3823 a_12465_1289# D[2] 0.0662f
C3824 D[2] a_13632_909# 8.06e-19
C3825 check[6] VDD_SW_b[7] 0.00177f
C3826 VDD_SW[4] a_8204_212# 2.77e-19
C3827 check[2] a_10103_1642# 0.00526f
C3828 a_8731_627# a_8409_n88# 7.32e-20
C3829 x9.A1 a_3421_n88# 6.68e-21
C3830 a_7663_n62# a_9742_n88# 5.13e-21
C3831 a_7649_993# m1_95_1942# 2.74e-20
C3832 a_8117_601# m1_95_2154# 2.82e-20
C3833 a_2879_n62# a_3356_n62# 1.96e-20
C3834 a_3421_n88# a_4338_n62# 0.189f
C3835 VSS_SW_b[6] a_3558_304# 3.58e-20
C3836 a_3420_212# a_4862_90# 0.00101f
C3837 a_3625_n88# a_4137_304# 6.69e-20
C3838 a_3112_106# a_2985_n62# 0.0256f
C3839 x2.X a_10532_n62# 3.68e-20
C3840 check[6] check[5] 0.00521f
C3841 a_1503_1642# x7.X 1.35e-19
C3842 VDD_SW[5] a_7203_627# 0.0865f
C3843 ready VDD_SW[7] 0.0363f
C3844 a_15907_627# a_15380_212# 7.07e-21
C3845 a_14545_627# m1_95_2154# 2.61e-20
C3846 x2.X check[4] 0.141f
C3847 VDD a_3535_n62# 0.00731f
C3848 a_14428_1467# x18.X 0.0878f
C3849 x9.A1 a_7369_627# 2.6e-19
C3850 x2.X a_8432_993# 0.187f
C3851 a_10597_n88# a_11514_n62# 0.189f
C3852 VSS_SW_b[3] a_10734_304# 3.58e-20
C3853 a_10596_212# a_12038_90# 0.00101f
C3854 a_10801_n88# a_11313_304# 6.69e-20
C3855 D[5] a_5943_627# 6.13e-19
C3856 a_27_627# a_2136_627# 1.75e-19
C3857 x2.X a_15799_220# 9.58e-19
C3858 x10.X a_5289_1289# 1.54e-19
C3859 check[5] a_2879_n62# 1.43e-20
C3860 VSS_SW[3] a_10596_212# 5.9e-22
C3861 a_174_n88# a_678_220# 0.00869f
C3862 a_1971_1642# VDD_SW[7] 5.38e-19
C3863 D[7] a_1415_895# 0.0294f
C3864 a_27_627# a_1256_993# 0.14f
C3865 VDD_SW_b[4] a_8319_n62# 5.2e-19
C3866 D[2] a_14839_n62# 3.12e-21
C3867 a_8921_304# VSS_SW[3] 6.59e-21
C3868 a_3183_627# a_3755_627# 2.46e-21
C3869 a_7769_n62# a_8140_n62# 4.19e-20
C3870 x2.X a_10103_1642# 2.63e-19
C3871 a_10596_212# m1_95_1942# 6.77e-21
C3872 x8.X a_193_627# 6.39e-20
C3873 x9.A1 VSS_SW_b[2] 2.54e-19
C3874 a_13375_895# a_13461_122# 4.53e-22
C3875 a_13216_993# a_13193_n88# 1.86e-19
C3876 a_8933_1642# D[3] 1.65e-19
C3877 check[6] a_78_90# 2.5e-20
C3878 VDD a_15329_304# 0.00298f
C3879 VDD a_5896_909# 0.0245f
C3880 check[4] a_4977_627# 5.33e-19
C3881 x17.X a_13936_1315# 0.00145f
C3882 a_5289_1289# D[5] 0.0662f
C3883 a_4149_1642# a_4363_1642# 0.00557f
C3884 check[4] VSS_SW[5] 0.0443f
C3885 a_5725_601# a_7649_993# 1.11e-20
C3886 a_6040_993# a_7369_627# 3.63e-21
C3887 VDD a_11071_1642# 0.191f
C3888 a_4860_1467# m1_95_2154# 8.35e-20
C3889 x2.X a_7769_n62# 5.57e-20
C3890 a_1415_895# a_2419_627# 6.86e-19
C3891 D[1] a_15585_n88# 0.00544f
C3892 check[0] a_14526_n88# 5.26e-19
C3893 a_941_601# D[6] 9.16e-19
C3894 a_5813_n88# a_7350_n88# 1.98e-19
C3895 a_5812_212# a_7663_n62# 2.63e-19
C3896 a_720_106# a_1143_n62# 0.00386f
C3897 a_1501_122# a_1946_n62# 0.0369f
C3898 a_487_n62# a_1369_n62# 0.00926f
C3899 a_174_n88# VSS_SW[6] 4.28e-21
C3900 D[7] VDD_SW_b[7] 0.453f
C3901 x18.X a_11987_627# 0.00113f
C3902 x16.X a_12341_627# 6.07e-19
C3903 a_4811_627# a_5271_n62# 7.27e-19
C3904 D[5] a_4958_n88# 0.00506f
C3905 a_193_627# a_473_993# 0.15f
C3906 VDD VSS_SW[7] 1.11f
C3907 a_8591_895# a_8731_627# 0.0383f
C3908 D[4] VSS_SW_b[3] 1.99e-19
C3909 x14.X a_9154_1315# 3.14e-20
C3910 a_8117_601# a_8539_627# 1.96e-20
C3911 a_7649_993# VDD_SW[4] 4.17e-21
C3912 check[5] D[7] 6.16e-20
C3913 a_1415_895# m1_95_2154# 5.86e-20
C3914 a_941_601# m1_95_1942# 4.09e-20
C3915 x2.X a_13461_122# 0.0043f
C3916 x6.X VSS_SW[7] 0.249f
C3917 x2.X a_1555_627# 0.0151f
C3918 VDD_SW_b[5] a_7823_601# 2.22e-20
C3919 VDD_SW_b[3] a_10532_n62# 8.12e-20
C3920 x2.X a_381_627# 0.00139f
C3921 x9.A1 a_647_601# 2.81e-20
C3922 a_5748_n62# a_6153_n62# 2.46e-21
C3923 VDD_SW_b[7] a_2419_627# 5.96e-19
C3924 a_2136_627# VDD_SW[7] 0.0729f
C3925 a_1555_627# a_1363_627# 4.19e-20
C3926 a_10041_993# a_10149_627# 0.00807f
C3927 a_10824_993# a_10680_909# 0.00412f
C3928 a_10215_601# a_10727_627# 9.75e-19
C3929 a_10509_601# a_10359_627# 0.00926f
C3930 D[3] a_10908_993# 2.53e-19
C3931 VDD a_12989_n88# 0.661f
C3932 a_1256_993# VDD_SW[7] 3.28e-20
C3933 a_9761_627# a_10509_601# 0.126f
C3934 VSS_SW[1] a_15030_220# 4.25e-19
C3935 a_14839_n62# VSS_SW_b[1] 0.0142f
C3936 a_15380_212# a_15585_n88# 0.15f
C3937 a_4689_2457# m1_95_2154# 6.79e-19
C3938 a_2927_1642# D[6] 5.72e-19
C3939 a_9949_627# VSS_SW[3] 0.00595f
C3940 a_4149_1642# a_4860_1467# 0.00963f
C3941 a_193_627# a_1159_627# 2.14e-20
C3942 a_381_627# a_557_993# 8.99e-19
C3943 a_473_993# a_791_627# 0.025f
C3944 a_941_601# a_1340_993# 9.41e-19
C3945 x7.X a_2585_627# 1.68e-19
C3946 a_2897_1289# VSS_SW[6] 0.00189f
C3947 check[5] a_2419_627# 0.00121f
C3948 a_8591_895# a_10824_993# 1.86e-21
C3949 VDD_SW_b[7] m1_95_2154# 9.75e-21
C3950 x9.A1 a_12901_601# 0.00103f
C3951 a_13515_627# a_12988_212# 7.07e-21
C3952 a_27_627# VSS_SW[7] 0.0565f
C3953 x9.A1 a_4338_n62# 1.9e-20
C3954 a_6285_1642# m1_95_2154# 1.04e-19
C3955 a_12153_627# a_12341_627# 0.189f
C3956 a_12607_601# a_13216_993# 0.00189f
C3957 a_12178_1642# VSS_SW[2] 0.00105f
C3958 check[5] a_4077_1642# 0.00577f
C3959 a_3421_n88# a_5812_212# 4.01e-22
C3960 a_3420_212# a_5813_n88# 5.48e-21
C3961 a_505_1289# a_647_601# 8.76e-20
C3962 x15.X a_12038_90# 0.0273f
C3963 a_12465_1289# D[3] 5.1e-21
C3964 check[5] m1_95_2154# 0.0352f
C3965 VDD VSS_SW_b[5] 0.0985f
C3966 a_2585_627# a_3420_212# 1.02e-19
C3967 a_2865_993# a_2879_n62# 2.63e-19
C3968 a_3039_601# a_3112_106# 1.01e-19
C3969 VDD x16.X 0.418f
C3970 x9.X VDD_SW[6] 0.176f
C3971 a_3333_601# a_2566_n88# 0.00259f
C3972 x15.X m1_95_1942# 2.53e-20
C3973 a_791_627# a_1159_627# 3.34e-19
C3974 a_1112_909# VDD_SW_b[7] 4.69e-21
C3975 VDD a_3333_601# 0.494f
C3976 x9.A1 a_14570_1642# 8.64e-19
C3977 x9.A1 a_505_1289# 0.104f
C3978 a_10055_n62# a_10161_n62# 0.0526f
C3979 a_13375_895# a_14733_627# 8.26e-21
C3980 check[1] VDD_SW_b[2] 0.0021f
C3981 check[1] a_13461_1642# 0.257f
C3982 a_3895_1642# a_3420_212# 1.39e-21
C3983 x2.X a_6124_993# 4.54e-19
C3984 x9.A1 a_6040_993# 4.84e-21
C3985 a_8679_1642# D[4] 0.0682f
C3986 check[3] VSS_SW_b[4] 1.77e-20
C3987 a_7203_627# a_9761_627# 1.08e-20
C3988 a_7369_627# a_9595_627# 1.14e-20
C3989 a_5323_2457# x9.A1 1.72f
C3990 x7.X a_1501_122# 2.79e-19
C3991 x2.X a_12433_993# 0.15f
C3992 a_12988_212# VSS_SW[1] 0.0872f
C3993 VSS_SW_b[2] a_12553_n62# 0.00334f
C3994 a_13193_n88# a_13103_n62# 9.75e-19
C3995 a_12989_n88# a_13329_n62# 6.04e-20
C3996 a_2468_1467# D[6] 0.0183f
C3997 x11.X a_6199_895# 0.00663f
C3998 VDD VDD_SW[5] 0.495f
C3999 a_218_1642# VSS_SW[7] 0.00105f
C4000 D[2] a_13193_n88# 0.00546f
C4001 x20.X m1_95_2154# 1.32e-20
C4002 VDD_SW_b[1] m1_95_2154# 1.39e-20
C4003 a_14545_627# a_16024_909# 7.17e-20
C4004 a_9154_1315# VDD_SW_b[4] 2.65e-20
C4005 a_15293_601# a_15143_627# 0.00926f
C4006 a_15608_993# a_15464_909# 0.00412f
C4007 a_14999_601# a_15511_627# 9.75e-19
C4008 a_14825_993# a_14933_627# 0.00807f
C4009 a_10824_993# VDD_SW[3] 3.28e-20
C4010 x9.A1 a_9742_n88# 7.4e-19
C4011 VDD a_13906_n62# 0.109f
C4012 a_4149_1642# check[5] 0.318f
C4013 VDD a_4064_909# 0.0044f
C4014 a_2468_1467# m1_95_1942# 1.97e-19
C4015 a_6285_122# a_6529_n62# 0.00807f
C4016 a_6730_n62# a_7350_n88# 8.26e-21
C4017 VDD a_12153_627# 0.722f
C4018 a_1757_1642# a_1971_1642# 0.00557f
C4019 a_14839_n62# a_15495_n62# 3.73e-19
C4020 a_15585_n88# a_16097_304# 6.69e-20
C4021 VSS_SW_b[1] a_15518_304# 3.58e-20
C4022 a_15072_106# a_15316_n62# 0.00707f
C4023 a_15381_n88# a_16298_n62# 0.189f
C4024 a_1166_304# VSS_SW[6] 2.77e-20
C4025 VDD_SW[4] a_9949_627# 6.11e-20
C4026 a_5431_601# a_5896_909# 9.46e-19
C4027 VDD a_7711_1642# 8.63e-19
C4028 x2.X a_14733_627# 0.00139f
C4029 x2.X a_15855_1642# 0.00645f
C4030 x9.A1 a_13715_1642# 0.195f
C4031 a_13715_1642# a_12901_601# 7.56e-21
C4032 a_4860_1467# a_4958_n88# 6.87e-20
C4033 a_12036_1467# check[2] 1.58e-19
C4034 a_5323_2457# a_6040_993# 2.04e-19
C4035 x17.X a_12447_n62# 0.00192f
C4036 a_8933_1642# x13.X 0.0843f
C4037 x12.X m1_95_2154# 6.47e-20
C4038 a_12153_627# a_14096_627# 2.2e-20
C4039 x11.X VDD_SW_b[5] 0.24f
C4040 VDD a_15767_895# 0.671f
C4041 VDD_SW[5] a_7733_993# 6.61e-21
C4042 D[4] a_8409_n88# 0.00544f
C4043 a_12134_n88# a_12447_n62# 0.245f
C4044 a_2419_627# a_2865_993# 0.159f
C4045 D[6] a_3039_601# 0.00583f
C4046 VSS_SW[4] a_8409_n88# 9.92e-21
C4047 a_7252_1467# D[4] 0.0183f
C4048 x9.A1 a_14791_1315# 0.00504f
C4049 x9.A1 a_15907_627# 5.3e-20
C4050 a_7252_1467# VSS_SW[4] 0.0274f
C4051 a_10597_n88# a_12680_106# 1.67e-21
C4052 a_11313_304# a_11514_n62# 8.99e-19
C4053 a_11069_122# a_12134_n88# 8e-21
C4054 a_10596_212# a_12988_212# 1.9e-21
C4055 VDD_SW[2] a_14999_601# 7.64e-20
C4056 check[1] x18.X 5.77e-19
C4057 a_193_627# a_2585_627# 3.26e-19
C4058 x14.X D[4] 0.00106f
C4059 a_10801_n88# a_11069_122# 0.206f
C4060 VSS_SW[3] a_11015_220# 6.42e-21
C4061 a_10597_n88# VSS_SW_b[3] 7.59e-19
C4062 a_5289_1289# a_6285_1642# 0.0146f
C4063 x13.X a_7350_n88# 1.64e-21
C4064 x2.X a_12036_1467# 2.86e-19
C4065 a_3039_601# m1_95_1942# 3.42e-20
C4066 a_2865_993# m1_95_2154# 1.86e-20
C4067 x9.A1 a_5812_212# 1.28e-20
C4068 a_13193_n88# VSS_SW_b[1] 4.54e-20
C4069 a_13705_304# VSS_SW[1] 6.59e-21
C4070 check[5] a_5289_1289# 4.15e-21
C4071 a_4338_n62# a_5812_212# 2.79e-22
C4072 D[2] a_14430_90# 8.78e-19
C4073 D[2] a_12607_601# 0.00583f
C4074 a_11987_627# a_12433_993# 0.159f
C4075 x12.X a_5257_993# 1.55e-20
C4076 VDD_SW_b[3] a_12433_993# 8.18e-21
C4077 a_1757_1642# a_2136_627# 5.9e-19
C4078 x2.X a_3807_895# 0.148f
C4079 x11.X a_5504_106# 1.89e-20
C4080 a_15608_993# VDD_SW[1] 3.28e-20
C4081 a_2419_627# a_3551_627# 0.00272f
C4082 a_4413_2457# a_3807_895# 7.82e-20
C4083 reset x2.X 1.3e-19
C4084 VDD a_5748_n62# 8.82e-19
C4085 x9.A1 a_4149_1315# 0.00499f
C4086 VDD a_9644_1467# 0.132f
C4087 check[3] check[2] 0.00521f
C4088 a_9761_627# a_12341_627# 3.67e-21
C4089 a_305_2457# x3.X 0.236f
C4090 a_11071_1642# a_10824_993# 0.00176f
C4091 a_29_2457# ready 0.0408f
C4092 x9.A1 a_9595_627# 7.95e-19
C4093 VDD_SW[7] a_3333_601# 2.55e-20
C4094 a_8933_1642# a_8204_212# 1.17e-22
C4095 x2.X a_16488_627# 3.63e-19
C4096 x9.X a_3421_n88# 0.0186f
C4097 a_15293_601# VSS_SW[1] 2.13e-19
C4098 a_6040_993# a_5812_212# 8.94e-21
C4099 a_14857_1289# D[2] 5.1e-21
C4100 a_11987_627# a_14733_627# 4.74e-21
C4101 a_5725_601# a_6017_n88# 0.00251f
C4102 a_6199_895# a_5813_n88# 6.35e-19
C4103 x9.A1 a_13643_1642# 5.26e-19
C4104 a_941_601# a_1028_212# 6.03e-19
C4105 a_1256_993# a_487_n62# 3.59e-19
C4106 a_381_627# a_174_n88# 3.32e-19
C4107 VDD a_678_220# 0.00634f
C4108 VSS_SW_b[4] a_8921_n62# 6.94e-20
C4109 a_10073_1289# x15.X 1.7e-20
C4110 check[6] a_1369_n62# 9.72e-20
C4111 a_3333_601# a_5431_601# 1.55e-20
C4112 x2.X VDD_SW_b[6] 7.3e-19
C4113 a_3807_895# a_4977_627# 2.8e-19
C4114 a_3807_895# VSS_SW[5] 7.52e-21
C4115 a_4413_2457# VDD_SW_b[6] 6.5e-20
C4116 check[4] a_6153_n62# 1.5e-20
C4117 x2.X a_10727_627# 0.00706f
C4118 a_7203_627# a_8432_993# 0.14f
C4119 D[4] a_8591_895# 0.0294f
C4120 VSS_SW[2] VSS_SW_b[2] 0.00722f
C4121 x2.X check[3] 0.142f
C4122 a_14428_1467# a_14570_1315# 0.00783f
C4123 x2.X a_2831_1315# 3.19e-19
C4124 x9.A1 a_1233_n88# 3.89e-20
C4125 a_7663_n62# a_7896_106# 0.124f
C4126 a_7350_n88# a_8204_212# 0.0319f
C4127 D[1] a_15464_909# 8.49e-19
C4128 check[0] a_15767_895# 0.00271f
C4129 a_14379_627# a_15692_993# 2.13e-19
C4130 a_16037_1642# D[1] 5.74e-19
C4131 VSS_SW[6] a_2566_n88# 0.00677f
C4132 a_1028_212# a_2985_n62# 1.09e-19
C4133 a_5431_601# VDD_SW[5] 2.07e-20
C4134 a_6199_895# a_6920_627# 0.0967f
C4135 a_5725_601# a_6339_627# 0.0526f
C4136 VDD_SW_b[5] a_5813_n88# 0.0406f
C4137 VDD a_10359_627# 1.8e-19
C4138 VDD_SW_b[7] a_720_106# 5.23e-19
C4139 VDD VSS_SW[6] 0.865f
C4140 x9.A1 a_15585_n88# 3.88e-20
C4141 a_14430_90# VSS_SW_b[1] 0.19f
C4142 a_9595_627# a_9742_n88# 0.00176f
C4143 VDD a_9761_627# 0.669f
C4144 VDD a_6753_1642# 0.00244f
C4145 a_11325_1642# D[2] 1.73e-19
C4146 a_12036_1467# a_11987_627# 5.32e-19
C4147 x2.X a_12495_1642# 2.63e-19
C4148 VDD_SW_b[6] a_4977_627# 0.00337f
C4149 x8.X a_2610_1315# 8.34e-19
C4150 check[1] a_13461_122# 2.02e-20
C4151 VDD_SW_b[6] VSS_SW[5] 0.00248f
C4152 x15.X a_12988_212# 1.68e-21
C4153 VDD_SW[3] a_12851_909# 2.16e-20
C4154 x27.A VDD_SW[6] 0.0227f
C4155 D[4] VDD_SW_b[4] 0.454f
C4156 a_16024_909# VDD_SW_b[1] 3.65e-20
C4157 D[4] a_9646_90# 8.78e-19
C4158 a_7681_1289# D[5] 1.02e-20
C4159 x16.X a_10824_993# 2.81e-19
C4160 VDD a_14379_627# 0.475f
C4161 VDD VDD_SW_b[2] 0.157f
C4162 VDD a_13461_1642# 0.191f
C4163 VDD_SW_b[5] a_6920_627# 0.185f
C4164 VDD_SW[2] m1_95_1942# 0.0331f
C4165 a_15855_1642# a_15853_122# 1.57e-21
C4166 a_16109_1642# D[1] 0.061f
C4167 a_13715_1642# a_13643_1642# 6.64e-19
C4168 a_14096_627# a_14379_627# 0.00111f
C4169 VDD_SW_b[2] a_14096_627# 0.185f
C4170 a_27_627# VSS_SW[6] 4.66e-21
C4171 x9.A1 a_6529_304# 5.63e-21
C4172 a_4958_n88# a_6285_122# 4.59e-22
C4173 a_5504_106# a_5813_n88# 0.0327f
C4174 a_5271_n62# a_6017_n88# 0.199f
C4175 x2.X a_15381_n88# 0.0206f
C4176 x8.X a_2470_90# 0.00259f
C4177 VSS_SW[7] a_487_n62# 3.44e-19
C4178 VDD a_8677_122# 0.334f
C4179 x9.A1 VSS_SW[2] 0.103f
C4180 a_12901_601# VSS_SW[2] 2.17e-19
C4181 check[2] a_10937_n62# 8.72e-20
C4182 a_7649_993# a_7350_n88# 8.71e-20
C4183 a_4370_1315# VDD_SW_b[6] 2.65e-20
C4184 a_7823_601# a_7663_n62# 0.0026f
C4185 a_16330_1315# D[1] 0.0012f
C4186 D[1] VDD_SW[1] 0.246f
C4187 x9.A1 a_10041_993# 8.95e-20
C4188 a_10824_993# a_12153_627# 3.63e-21
C4189 a_10509_601# a_12433_993# 1.11e-20
C4190 VDD a_15072_106# 0.37f
C4191 check[2] a_10215_601# 0.00262f
C4192 x2.X a_977_304# 0.00167f
C4193 x9.A1 x9.X 6.77e-19
C4194 x9.X a_4338_n62# 0.00158f
C4195 a_16109_1642# a_15380_212# 1.17e-22
C4196 a_6199_895# a_6730_n62# 4.06e-19
C4197 a_5257_993# a_5377_n62# 6.88e-22
C4198 a_647_601# a_593_n62# 1.07e-20
C4199 a_6539_1642# D[5] 0.0605f
C4200 VDD_SW_b[2] a_13329_n62# 0.00179f
C4201 a_8679_1642# m1_95_2154# 1.04e-19
C4202 ready check[6] 0.0393f
C4203 D[2] D[1] 0.00183f
C4204 check[1] a_12433_993# 7.12e-20
C4205 x9.A1 a_7394_1315# 4.35e-20
C4206 check[2] a_11539_1642# 0.00688f
C4207 reset a_76_1467# 8.22e-19
C4208 a_7557_627# VSS_SW_b[4] 1.42e-19
C4209 VDD x18.X 0.421f
C4210 a_2585_627# a_3504_909# 0.00907f
C4211 a_2865_993# a_2949_993# 0.00972f
C4212 a_3333_601# a_2773_627# 1.24e-20
C4213 a_3807_895# a_3648_993# 0.207f
C4214 a_8205_n88# a_7854_220# 4.48e-20
C4215 a_3039_601# a_3283_909# 0.0104f
C4216 a_7896_106# a_8342_304# 0.00412f
C4217 a_8204_212# a_8153_304# 2.13e-19
C4218 a_7663_n62# a_8623_220# 1.21e-20
C4219 a_3420_212# a_3893_122# 0.159f
C4220 a_3112_106# VSS_SW_b[6] 0.00322f
C4221 a_3421_n88# a_3625_n88# 0.117f
C4222 VSS_SW[6] a_3369_304# 8.28e-20
C4223 check[6] a_1971_1642# 0.00688f
C4224 x17.X m1_95_1942# 2.51e-20
C4225 x2.X a_10215_601# 0.2f
C4226 a_15907_627# a_15585_n88# 7.32e-20
C4227 a_14825_993# m1_95_2154# 1.86e-20
C4228 a_15767_895# a_15721_n62# 1.65e-20
C4229 a_12038_90# a_12134_n88# 0.0967f
C4230 VDD_SW[7] VSS_SW[6] 0.412f
C4231 a_14545_627# a_14999_601# 0.117f
C4232 VDD_SW_b[5] a_6730_n62# 0.0145f
C4233 check[0] a_14379_627# 0.00121f
C4234 a_13461_1642# check[0] 2.07e-21
C4235 x18.X a_14096_627# 0.0285f
C4236 check[5] a_3947_627# 4.06e-19
C4237 a_305_2457# a_473_993# 4.56e-21
C4238 x3.X a_647_601# 3.71e-19
C4239 a_9742_n88# VSS_SW[2] 4.18e-21
C4240 a_11069_122# a_11514_n62# 0.0369f
C4241 x10.X D[6] 9.68e-19
C4242 a_29_2457# VSS_SW[7] 0.0221f
C4243 VDD a_10532_n62# 7.87e-19
C4244 x2.X a_16298_n62# 1.24e-19
C4245 a_10041_993# a_9742_n88# 8.71e-20
C4246 VDD_SW[6] a_5165_627# 6.11e-20
C4247 VSS_SW[1] a_14839_n62# 3.44e-19
C4248 VSS_SW[3] a_10801_n88# 9.92e-21
C4249 VDD check[4] 2f
C4250 a_8204_212# a_10161_n62# 1.09e-19
C4251 D[2] a_15380_212# 5.78e-20
C4252 x30.A D[5] 1.01e-19
C4253 VDD a_8432_993# 0.227f
C4254 x10.X m1_95_1942# 1.18e-19
C4255 a_11325_1642# a_10983_895# 0.00232f
C4256 x8.X a_1757_1315# 1.78e-20
C4257 a_8205_n88# VSS_SW[3] 9.23e-19
C4258 a_8409_n88# a_8545_n62# 0.0697f
C4259 a_3648_993# VDD_SW_b[6] 4.99e-20
C4260 VSS_SW_b[4] a_8140_n62# 1.68e-19
C4261 D[6] D[5] 0.00189f
C4262 x3.X x9.A1 9e-19
C4263 a_11325_1642# D[3] 0.0604f
C4264 a_7369_627# a_7823_601# 0.117f
C4265 VDD a_15799_220# 0.00984f
C4266 a_8205_n88# m1_95_1942# 1.16e-21
C4267 a_7252_1467# m1_95_2154# 8.35e-20
C4268 VDD a_10103_1642# 8.63e-19
C4269 D[5] m1_95_1942# 0.0335f
C4270 check[0] a_15072_106# 8.65e-22
C4271 ready D[7] 0.038f
C4272 D[1] VSS_SW_b[1] 4.85e-19
C4273 x2.X VSS_SW_b[4] 0.0279f
C4274 a_12036_1467# check[1] 0.318f
C4275 x14.X m1_95_2154# 3.72e-20
C4276 a_5813_n88# a_6231_220# 0.00276f
C4277 a_6017_n88# a_5950_304# 9.46e-19
C4278 a_4958_n88# a_5377_n62# 0.0383f
C4279 a_5271_n62# a_7254_90# 3.67e-21
C4280 VSS_SW_b[5] a_5462_220# 5.33e-20
C4281 a_5812_212# a_6529_304# 4.45e-20
C4282 a_1029_n88# a_1501_122# 0.15f
C4283 VSS_SW[7] a_1447_220# 6.42e-21
C4284 VDD_SW_b[4] a_10597_n88# 2.44e-21
C4285 a_1028_212# VSS_SW_b[7] 0.00119f
C4286 x3.X a_505_1289# 2.51e-20
C4287 a_9646_90# a_10597_n88# 9.87e-21
C4288 x11.X a_7663_n62# 4.73e-20
C4289 VDD a_7769_n62# 0.0133f
C4290 x7.X a_941_601# 1.26e-19
C4291 a_7823_601# a_7967_627# 0.0697f
C4292 a_8117_601# a_8288_909# 0.00652f
C4293 a_1971_1642# D[7] 0.00163f
C4294 check[6] a_1256_993# 3.41e-19
C4295 x10.X a_5725_601# 5e-20
C4296 D[6] VSS_SW_b[6] 5.32e-19
C4297 VDD_SW_b[3] a_10937_n62# 0.00179f
C4298 ready a_2419_627# 1.4e-20
C4299 x9.X a_5812_212# 8.4e-22
C4300 x18.X check[0] 0.009f
C4301 a_10215_601# VDD_SW_b[3] 1.75e-20
C4302 a_10824_993# a_10359_627# 0.00316f
C4303 a_10509_601# a_10727_627# 3.73e-19
C4304 a_11123_627# a_11069_122# 2.54e-20
C4305 x16.X a_12399_1315# 2.4e-19
C4306 a_9595_627# VSS_SW[2] 4.66e-21
C4307 VDD a_13461_122# 0.313f
C4308 a_9761_627# a_10824_993# 0.0334f
C4309 a_15381_n88# a_15853_122# 0.15f
C4310 a_15380_212# VSS_SW_b[1] 0.00119f
C4311 a_9595_627# a_10041_993# 0.159f
C4312 VSS_SW[1] a_15518_304# 1.97e-20
C4313 a_4363_1642# D[6] 0.00163f
C4314 x9.X a_4149_1315# 2.08e-19
C4315 ready m1_95_2154# 1.91e-19
C4316 VDD a_1555_627# 6.99e-19
C4317 a_939_2457# m1_95_1942# 0.00139f
C4318 D[5] a_5725_601# 0.0192f
C4319 a_2610_1642# VSS_SW[6] 0.00105f
C4320 a_4811_627# a_6199_895# 0.0321f
C4321 VDD_SW_b[6] a_4137_n62# 5.22e-19
C4322 VDD a_381_627# 0.125f
C4323 a_13515_627# a_13193_n88# 7.32e-20
C4324 VDD_SW[2] a_12988_212# 4.35e-19
C4325 x9.A1 a_13216_993# 4.84e-21
C4326 a_8067_909# VDD_SW_b[4] 3.61e-21
C4327 a_12153_627# a_12851_909# 0.00276f
C4328 a_12901_601# a_13216_993# 0.13f
C4329 a_12433_993# a_12341_627# 0.0369f
C4330 a_12607_601# a_12517_993# 6.69e-20
C4331 a_8117_601# VSS_SW[3] 2.9e-20
C4332 a_8591_895# a_8545_n62# 1.65e-20
C4333 a_8731_627# a_8677_122# 2.54e-20
C4334 x9.A1 a_6539_1315# 0.00496f
C4335 a_2585_627# VDD_SW[6] 1.96e-20
C4336 a_7896_106# a_9742_n88# 1.86e-21
C4337 x6.X a_381_627# 6.12e-19
C4338 a_3333_601# a_4528_627# 5.73e-19
C4339 a_8591_895# m1_95_2154# 5.86e-20
C4340 VSS_SW_b[6] a_3839_220# 1.12e-20
C4341 a_3625_n88# a_4338_n62# 8.07e-20
C4342 a_3112_106# a_3356_n62# 0.00707f
C4343 a_3893_122# a_4137_304# 0.00972f
C4344 a_8117_601# m1_95_1942# 4.09e-20
C4345 a_3421_n88# a_4862_90# 5.39e-19
C4346 a_2879_n62# a_3535_n62# 3.73e-19
C4347 VDD_SW[5] D[4] 4.55e-19
C4348 VDD_SW_b[5] a_8204_212# 2.29e-22
C4349 a_14545_627# m1_95_1942# 3.82e-20
C4350 VDD_SW[5] VSS_SW[4] 0.396f
C4351 VDD a_3761_n62# 0.0321f
C4352 x9.A1 a_7823_601# 2.81e-20
C4353 x2.X a_7557_627# 0.0014f
C4354 x9.A1 a_16037_1642# 5.26e-19
C4355 a_10055_n62# a_10711_n62# 3.73e-19
C4356 a_4811_627# VDD_SW_b[5] 1.12e-19
C4357 D[5] a_6456_909# 8.07e-19
C4358 a_10288_106# a_10532_n62# 0.00707f
C4359 check[1] a_12495_1642# 0.00526f
C4360 D[7] a_2136_627# 0.00238f
C4361 check[5] a_3112_106# 8.68e-22
C4362 a_487_n62# a_678_220# 3.24e-19
C4363 a_7711_1642# D[4] 5.72e-19
C4364 check[3] a_7203_627# 0.0012f
C4365 x11.X a_7369_627# 1.68e-19
C4366 VDD_SW_b[4] a_8545_n62# 0.00179f
C4367 D[7] a_1256_993# 0.00608f
C4368 a_27_627# a_381_627# 0.0455f
C4369 x30.A a_4860_1467# 6.58e-20
C4370 a_9122_n62# VSS_SW[3] 6.09e-20
C4371 ready a_4149_1642# 6.63e-21
C4372 x2.X a_13375_895# 0.148f
C4373 VSS_SW_b[2] a_13103_n62# 5.23e-19
C4374 a_13193_n88# VSS_SW[1] 8.41e-20
C4375 a_13461_122# a_13329_n62# 0.025f
C4376 a_4860_1467# D[6] 2.91e-19
C4377 VDD_SW_b[4] m1_95_2154# 1.43e-20
C4378 x8.X a_647_601# 1.98e-20
C4379 x27.A x9.A1 1.25e-19
C4380 x2.X check[2] 0.148f
C4381 D[2] VSS_SW_b[2] 5.22e-19
C4382 x2.X a_5223_1315# 3.19e-19
C4383 check[6] VSS_SW[7] 0.0441f
C4384 a_4860_1467# a_5002_1642# 0.00557f
C4385 VDD a_6124_993# 0.00439f
C4386 a_14999_601# VDD_SW_b[1] 2.14e-20
C4387 a_15608_993# a_15143_627# 0.00316f
C4388 check[4] a_5431_601# 0.00262f
C4389 a_15293_601# a_15511_627# 3.73e-19
C4390 a_2773_627# VSS_SW[6] 0.00595f
C4391 a_6199_895# a_7649_993# 8e-21
C4392 a_4977_627# a_7557_627# 3.67e-21
C4393 a_5725_601# a_8117_601# 9.37e-21
C4394 a_4860_1467# m1_95_1942# 1.97e-19
C4395 x12.X a_7681_1289# 1.51e-19
C4396 a_2136_627# a_2419_627# 0.0011f
C4397 a_2468_1467# x7.X 4.97e-19
C4398 x2.X a_8140_n62# 3.68e-20
C4399 VDD a_12433_993# 0.211f
C4400 a_15380_212# a_15495_n62# 0.00272f
C4401 a_15072_106# a_15721_n62# 0.00316f
C4402 a_15853_122# a_16298_n62# 0.0369f
C4403 x9.A1 x8.X 9.17e-19
C4404 a_5812_212# a_7896_106# 5.96e-20
C4405 a_5813_n88# a_7663_n62# 4.56e-21
C4406 a_1415_895# D[6] 2.13e-19
C4407 a_1256_993# a_2419_627# 7.46e-20
C4408 VDD a_9147_1642# 0.00244f
C4409 a_720_106# a_1369_n62# 0.00316f
C4410 x2.X a_14887_1642# 2.63e-19
C4411 a_1028_212# a_1143_n62# 0.00272f
C4412 a_487_n62# VSS_SW[6] 1.64e-20
C4413 x2.X a_15243_909# 0.00138f
C4414 VDD_SW[3] m1_95_2154# 0.0327f
C4415 x9.A1 a_16109_1642# 0.195f
C4416 D[5] a_5271_n62# 0.00258f
C4417 x17.X a_12988_212# 0.245f
C4418 a_4811_627# a_5504_106# 3.88e-21
C4419 a_2136_627# m1_95_2154# 1.66e-20
C4420 a_193_627# a_941_601# 0.126f
C4421 a_647_601# a_473_993# 0.206f
C4422 a_8432_993# a_8731_627# 0.0256f
C4423 a_8117_601# VDD_SW[4] 1.83e-19
C4424 a_1415_895# m1_95_1942# 8.62e-20
C4425 a_1256_993# m1_95_2154# 4.11e-21
C4426 a_4413_2457# x2.X 0.00426f
C4427 x2.X a_3070_220# 0.0028f
C4428 a_4689_2457# x30.A 0.236f
C4429 VDD a_15855_1642# 0.196f
C4430 VDD a_14733_627# 0.125f
C4431 x2.X a_1363_627# 0.00111f
C4432 a_4689_2457# D[6] 0.00292f
C4433 a_12447_n62# a_12680_106# 0.124f
C4434 VDD_SW_b[5] a_7649_993# 8.18e-21
C4435 a_12134_n88# a_12988_212# 0.0319f
C4436 a_14428_1467# a_14887_1642# 6.64e-19
C4437 x9.A1 a_473_993# 1.02e-19
C4438 x2.X a_557_993# 5.31e-19
C4439 a_5927_n62# a_6153_n62# 3.34e-19
C4440 a_9644_1467# D[4] 2.78e-19
C4441 VDD_SW_b[7] D[6] 1.53e-19
C4442 a_10055_n62# VSS_SW_b[2] 9.32e-21
C4443 x9.A1 VDD_SW[1] 0.0323f
C4444 a_10597_n88# a_12989_n88# 1.33e-19
C4445 VDD_SW[2] a_15293_601# 2.55e-20
C4446 a_10215_601# a_10509_601# 0.199f
C4447 x16.X a_11546_1315# 5.02e-20
C4448 a_4689_2457# m1_95_1942# 3.15e-19
C4449 a_11069_122# VSS_SW_b[3] 7.15e-19
C4450 a_473_993# a_581_627# 0.00807f
C4451 a_1256_993# a_1112_909# 0.00412f
C4452 a_647_601# a_1159_627# 9.75e-19
C4453 a_193_627# a_1672_909# 7.17e-20
C4454 a_941_601# a_791_627# 0.00926f
C4455 x2.X a_14428_1467# 2.88e-19
C4456 check[5] D[6] 0.456f
C4457 a_8848_909# VDD_SW[4] 2.12e-20
C4458 a_14430_90# VSS_SW[1] 0.0819f
C4459 VDD_SW_b[7] m1_95_1942# 1.44e-20
C4460 x2.X a_4977_627# 0.0537f
C4461 D[7] VSS_SW[7] 0.118f
C4462 x2.X VSS_SW[5] 0.078f
C4463 a_6285_1642# m1_95_1942# 2.26e-19
C4464 x9.A1 D[2] 0.267f
C4465 a_4413_2457# VSS_SW[5] 3.26e-20
C4466 a_11987_627# a_13375_895# 0.0321f
C4467 a_2879_n62# VSS_SW_b[5] 1.09e-20
C4468 D[2] a_12901_601# 0.0191f
C4469 a_3421_n88# a_5813_n88# 1.33e-19
C4470 a_6539_1642# x12.X 7.67e-19
C4471 a_505_1289# a_473_993# 4.54e-19
C4472 check[2] VDD_SW_b[3] 0.00208f
C4473 check[5] m1_95_1942# 0.034f
C4474 x9.A1 x11.X 6.93e-19
C4475 VDD a_12036_1467# 0.153f
C4476 a_2585_627# a_3421_n88# 1.27e-19
C4477 a_3333_601# a_2879_n62# 3.74e-20
C4478 a_11253_1642# D[3] 5.74e-19
C4479 a_2865_993# a_3112_106# 4.96e-20
C4480 a_3039_601# a_3420_212# 4.51e-19
C4481 x2.X a_9312_627# 3.88e-19
C4482 x2.X a_15715_627# 0.00111f
C4483 x2.X a_16109_1315# 2.32e-19
C4484 a_14857_1289# VSS_SW[1] 0.00186f
C4485 VDD a_3807_895# 0.689f
C4486 x9.A1 a_1503_1642# 0.101f
C4487 a_11071_1642# m1_95_2154# 1.04e-19
C4488 VDD reset 0.158f
C4489 x2.X a_5575_627# 0.0388f
C4490 a_12851_909# VDD_SW_b[2] 2.4e-21
C4491 x9.A1 a_5165_627# 4.11e-19
C4492 a_4977_627# VSS_SW[5] 0.0232f
C4493 reset x6.X 1.55e-19
C4494 D[4] a_9761_627# 5.14e-21
C4495 x2.X a_12924_n62# 3.67e-20
C4496 VDD a_16488_627# 0.193f
C4497 VDD a_14570_1315# 0.0017f
C4498 VSS_SW[7] m1_95_2154# 0.0294f
C4499 x2.X a_11987_627# 0.354f
C4500 a_12988_212# a_12937_304# 2.13e-19
C4501 a_12989_n88# a_12638_220# 4.71e-20
C4502 a_12447_n62# a_13407_220# 1.21e-20
C4503 a_12680_106# a_13126_304# 0.00412f
C4504 VDD_SW_b[1] m1_95_1942# 2.05e-20
C4505 x2.X VDD_SW_b[3] 7.33e-19
C4506 x20.X m1_95_1942# 2.53e-20
C4507 VDD_SW_b[6] a_2566_n88# 3.21e-19
C4508 a_6285_1642# a_5725_601# 0.00263f
C4509 a_5323_2457# x11.X 3.01e-19
C4510 a_6920_627# a_7369_627# 5.39e-19
C4511 a_505_1289# a_1503_1642# 0.0146f
C4512 check[0] a_15855_1642# 0.257f
C4513 a_14379_627# a_14933_627# 0.00206f
C4514 D[3] VSS_SW_b[2] 2.05e-19
C4515 x17.X a_15293_601# 4.31e-21
C4516 a_7254_90# a_7350_n88# 0.0967f
C4517 VSS_SW_b[5] a_6529_n62# 6.93e-20
C4518 VDD VDD_SW_b[6] 0.157f
C4519 a_1028_212# VSS_SW_b[6] 0.00377f
C4520 a_1447_220# VSS_SW[6] 1.57e-20
C4521 D[7] a_3333_601# 2.67e-21
C4522 VDD_SW[4] a_10125_993# 6.61e-21
C4523 a_5725_601# a_5675_909# 1.21e-20
C4524 VDD a_10727_627# 6.2e-19
C4525 a_4977_627# a_5575_627# 6.04e-20
C4526 reset a_27_627# 7.49e-21
C4527 a_5575_627# VSS_SW[5] 0.0012f
C4528 VDD check[3] 1.92f
C4529 D[5] a_5950_304# 9.69e-19
C4530 x9.A1 VSS_SW_b[1] 1.46e-19
C4531 VDD a_2831_1315# 0.00162f
C4532 a_13715_1642# D[2] 0.0607f
C4533 x12.X m1_95_1942# 1.18e-19
C4534 VDD_SW[5] a_8067_909# 2.16e-20
C4535 a_7203_627# VSS_SW_b[4] 6.02e-20
C4536 D[4] a_8677_122# 0.00928f
C4537 VDD a_12495_1642# 0.00166f
C4538 VSS_SW[4] a_8677_122# 2.79e-21
C4539 a_2419_627# a_3333_601# 0.14f
C4540 D[6] a_2865_993# 0.00884f
C4541 x16.X m1_95_2154# 3.81e-20
C4542 a_13632_909# VDD_SW[2] 2.12e-20
C4543 x13.X a_7663_n62# 0.00192f
C4544 a_2865_993# m1_95_1942# 2.74e-20
C4545 a_3333_601# m1_95_2154# 2.82e-20
C4546 x2.X a_15853_122# 0.00427f
C4547 a_9742_n88# a_10055_n62# 0.245f
C4548 x9.A1 a_5813_n88# 7.54e-21
C4549 VDD_SW[6] a_4811_627# 0.0865f
C4550 a_4862_90# a_5812_212# 1.66e-20
C4551 x2.X a_76_1467# 2.67e-19
C4552 a_4338_n62# a_5813_n88# 3.67e-21
C4553 a_3558_304# VSS_SW_b[5] 9.9e-21
C4554 x12.X a_5725_601# 0.00124f
C4555 x9.A1 a_2585_627# 2.67e-19
C4556 x2.X a_3648_993# 0.187f
C4557 x11.X a_5812_212# 0.245f
C4558 a_11325_1642# a_10596_212# 1.17e-22
C4559 a_11123_627# a_10931_627# 4.19e-20
C4560 a_11704_627# VDD_SW[3] 0.0729f
C4561 D[6] a_3551_627# 6.12e-19
C4562 VDD_SW_b[3] a_11987_627# 5.95e-19
C4563 VDD a_5927_n62# 0.0074f
C4564 x9.A1 a_10983_895# 2.64e-19
C4565 x3.A ready 0.038f
C4566 a_10983_895# a_12901_601# 1.38e-20
C4567 VDD_SW[5] m1_95_2154# 0.0327f
C4568 VDD a_15381_n88# 0.673f
C4569 x9.A1 D[3] 0.254f
C4570 D[3] a_12901_601# 2.67e-21
C4571 VDD_SW[7] a_3807_895# 1.27e-20
C4572 check[2] a_10509_601# 1.88e-19
C4573 a_7681_1289# a_8679_1642# 0.0146f
C4574 a_9595_627# D[2] 1.19e-20
C4575 x2.X a_174_n88# 0.178f
C4576 x9.A1 a_3895_1642# 0.101f
C4577 x9.X a_3625_n88# 1.8e-19
C4578 D[1] VSS_SW[1] 0.118f
C4579 x9.A1 a_6920_627# 2.14e-20
C4580 a_12153_627# m1_95_2154# 2.61e-20
C4581 a_6199_895# a_6017_n88# 4.26e-19
C4582 a_5725_601# a_6285_122# 2.7e-19
C4583 a_1415_895# a_1028_212# 0.00165f
C4584 VDD a_977_304# 0.00318f
C4585 a_193_627# VSS_SW_b[7] 1.51e-20
C4586 a_941_601# a_1029_n88# 3.89e-19
C4587 check[1] a_13375_895# 0.00226f
C4588 a_13643_1642# D[2] 5.74e-19
C4589 x9.A1 a_8933_1315# 0.00499f
C4590 check[2] check[1] 0.0052f
C4591 check[6] VSS_SW[6] 1.39e-19
C4592 a_3333_601# a_5257_993# 1.11e-20
C4593 a_4149_1642# a_3333_601# 7.12e-21
C4594 a_3648_993# a_4977_627# 3.63e-21
C4595 check[4] D[4] 3.66e-20
C4596 check[4] VSS_SW[4] 1.4e-19
C4597 a_7203_627# a_7557_627# 0.0455f
C4598 D[4] a_8432_993# 0.00608f
C4599 a_15767_895# m1_95_2154# 5.86e-20
C4600 x2.X a_10509_601# 0.119f
C4601 a_7350_n88# a_8205_n88# 0.0477f
C4602 a_7663_n62# a_8204_212# 0.138f
C4603 a_11514_n62# a_12988_212# 5.58e-22
C4604 x9.A1 a_1501_122# 4.39e-20
C4605 VDD_SW_b[7] a_3283_909# 2.1e-21
C4606 VSS_SW[6] a_2879_n62# 3.44e-19
C4607 a_1946_n62# VSS_SW_b[6] 2.63e-19
C4608 a_14545_627# a_15293_601# 0.126f
C4609 a_14999_601# a_14825_993# 0.206f
C4610 a_5725_601# a_6147_627# 1.96e-20
C4611 x27.A x9.X 9.96e-20
C4612 a_6199_895# a_6339_627# 0.0383f
C4613 a_5257_993# VDD_SW[5] 4.17e-21
C4614 x2.X a_2897_1289# 0.0112f
C4615 VDD_SW_b[5] a_6017_n88# 0.00133f
C4616 D[5] a_7350_n88# 4.26e-19
C4617 a_12465_1289# x17.X 1.79e-20
C4618 VDD a_10937_n62# 0.0301f
C4619 VDD_SW_b[7] a_1028_212# 0.0416f
C4620 x2.X a_15316_n62# 3.67e-20
C4621 a_9761_627# a_10597_n88# 1.27e-19
C4622 x13.X a_7369_627# 1.02e-20
C4623 VSS_SW[1] a_15380_212# 1.18e-21
C4624 a_12680_106# m1_95_1942# 4.96e-22
C4625 a_5323_2457# a_6920_627# 3.86e-19
C4626 a_9595_627# a_10055_n62# 7.27e-19
C4627 VSS_SW[3] VSS_SW_b[3] 0.0075f
C4628 D[3] a_9742_n88# 0.0042f
C4629 VDD a_8921_n62# 7.11e-19
C4630 VDD a_10215_601# 0.313f
C4631 D[7] a_678_220# 1.98e-20
C4632 VDD_SW_b[6] a_5431_601# 2.23e-20
C4633 x2.X check[1] 0.149f
C4634 VDD a_1978_1315# 3.89e-19
C4635 x2.X a_7615_1315# 3.2e-19
C4636 a_12465_1289# a_12134_n88# 5.67e-21
C4637 a_1503_1642# a_1233_n88# 4.63e-19
C4638 VDD a_16298_n62# 0.109f
C4639 a_6467_1642# D[5] 5.74e-19
C4640 a_8933_1642# a_8117_601# 7.12e-21
C4641 a_9644_1467# m1_95_2154# 8.35e-20
C4642 VDD a_11539_1642# 0.00246f
C4643 check[0] a_15381_n88# 2.51e-20
C4644 x17.X a_14839_n62# 4.41e-20
C4645 check[3] a_8731_627# 1.35e-19
C4646 a_14428_1467# check[1] 1.57e-19
C4647 x2.X a_7203_627# 0.354f
C4648 D[7] VSS_SW[6] 4.85e-19
C4649 a_11325_1642# x15.X 0.0847f
C4650 a_9312_627# a_10509_601# 1.84e-20
C4651 x9.A1 a_6730_n62# 1.56e-20
C4652 a_5504_106# a_6017_n88# 0.00189f
C4653 a_4958_n88# VSS_SW_b[5] 0.134f
C4654 a_5271_n62# a_6285_122# 0.0633f
C4655 a_5812_212# a_5813_n88# 0.784f
C4656 VSS_SW[7] a_720_106# 4.63e-19
C4657 a_78_90# a_1028_212# 1.66e-20
C4658 a_12447_n62# a_14526_n88# 5.13e-21
C4659 VDD VSS_SW_b[4] 0.0971f
C4660 D[2] VSS_SW[2] 0.119f
C4661 a_7649_993# a_7663_n62# 2.63e-19
C4662 a_7823_601# a_7896_106# 1.01e-19
C4663 a_8117_601# a_7350_n88# 0.00259f
C4664 a_7369_627# a_8204_212# 1.02e-19
C4665 a_10509_601# a_11987_627# 3.81e-19
C4666 x2.X a_1166_304# 0.00334f
C4667 a_10983_895# a_11240_909# 0.00869f
C4668 a_10824_993# a_10727_627# 0.00386f
C4669 a_2419_627# VSS_SW[6] 0.0576f
C4670 a_9949_627# a_10149_627# 3.81e-19
C4671 a_10509_601# VDD_SW_b[3] 0.00636f
C4672 x9.X a_4862_90# 0.0273f
C4673 D[3] a_11240_909# 8.07e-19
C4674 a_4977_627# a_7203_627# 1.36e-20
C4675 a_4811_627# a_7369_627# 1.09e-20
C4676 a_15585_n88# VSS_SW_b[1] 9.21e-19
C4677 a_6920_627# a_5812_212# 6.63e-19
C4678 a_9595_627# a_10983_895# 0.0321f
C4679 a_6539_1642# a_7252_1467# 0.00957f
C4680 a_473_993# a_593_n62# 6.88e-22
C4681 a_9595_627# D[3] 0.138f
C4682 a_1415_895# a_1946_n62# 4.06e-19
C4683 x7.X VSS_SW_b[6] 0.0172f
C4684 a_939_2457# x7.X 2.37e-19
C4685 a_8679_1642# m1_95_1942# 2.26e-19
C4686 VSS_SW[6] m1_95_2154# 0.0337f
C4687 check[1] a_11987_627# 0.00121f
C4688 a_12607_601# a_13072_909# 9.46e-19
C4689 a_9761_627# m1_95_2154# 2.61e-20
C4690 x16.X a_11704_627# 0.0286f
C4691 x9.A1 x13.X 6.75e-19
C4692 a_7203_627# a_9312_627# 1.75e-19
C4693 a_8204_212# a_8342_304# 1.09e-19
C4694 a_3039_601# a_3504_909# 9.46e-19
C4695 a_3420_212# VSS_SW_b[6] 0.00119f
C4696 a_3421_n88# a_3893_122# 0.15f
C4697 VSS_SW[6] a_3558_304# 1.97e-20
C4698 a_14825_993# m1_95_1942# 2.74e-20
C4699 x2.X a_10246_220# 0.00279f
C4700 a_76_1467# a_174_n88# 6.87e-20
C4701 a_14379_627# m1_95_2154# 3.53e-20
C4702 VDD_SW_b[5] a_7254_90# 0.00346f
C4703 a_13461_1642# m1_95_2154# 1.04e-19
C4704 VDD_SW_b[2] m1_95_2154# 1.95e-20
C4705 a_10288_106# a_10937_n62# 0.00316f
C4706 VDD_SW_b[7] a_1946_n62# 0.0144f
C4707 a_10055_n62# VSS_SW[2] 1.46e-20
C4708 x3.X a_473_993# 4.27e-21
C4709 a_10596_212# a_10711_n62# 0.00272f
C4710 x3.A VSS_SW[7] 0.0165f
C4711 check[1] a_13929_1642# 0.00688f
C4712 a_10041_993# a_10055_n62# 2.63e-19
C4713 a_10215_601# a_10288_106# 1.01e-19
C4714 VDD_SW[6] a_5341_993# 6.61e-21
C4715 a_9147_1642# D[4] 0.00163f
C4716 a_12988_212# a_13705_n62# 0.00206f
C4717 x2.X a_12341_627# 0.00141f
C4718 VDD a_7557_627# 0.109f
C4719 a_8409_n88# VSS_SW[3] 8.81e-20
C4720 VSS_SW_b[4] a_8319_n62# 5.24e-19
C4721 a_8677_122# a_8545_n62# 0.025f
C4722 a_11704_627# a_12153_627# 5.39e-19
C4723 a_7369_627# a_7649_993# 0.15f
C4724 a_2468_1467# a_2610_1315# 0.00783f
C4725 a_15608_993# a_15511_627# 0.00386f
C4726 a_15293_601# VDD_SW_b[1] 0.00622f
C4727 x20.X a_15293_601# 1.31e-19
C4728 a_15767_895# a_16024_909# 0.00869f
C4729 a_14733_627# a_14933_627# 3.81e-19
C4730 a_11071_1642# a_11069_122# 1.57e-21
C4731 a_7252_1467# m1_95_1942# 1.97e-19
C4732 VSS_SW_b[1] a_14945_n62# 0.00335f
C4733 a_15381_n88# a_15721_n62# 6.04e-20
C4734 a_15380_212# a_16097_n62# 0.00206f
C4735 VDD a_13375_895# 0.672f
C4736 a_15585_n88# a_15495_n62# 9.75e-19
C4737 x13.X a_9742_n88# 0.00862f
C4738 x14.X VSS_SW[3] 0.251f
C4739 VDD check[2] 1.74f
C4740 VDD a_5223_1315# 9.5e-20
C4741 x9.A1 a_8204_212# 5.79e-21
C4742 a_14545_627# a_14839_n62# 2.38e-19
C4743 a_14999_601# a_14526_n88# 4.37e-19
C4744 x2.X a_15692_993# 4.67e-19
C4745 x14.X m1_95_1942# 6.49e-20
C4746 a_5812_212# a_6730_n62# 0.0453f
C4747 a_6017_n88# a_6231_220# 0.0104f
C4748 a_5813_n88# a_6529_304# 0.0018f
C4749 a_5271_n62# a_5377_n62# 0.0526f
C4750 a_1233_n88# a_1501_122# 0.206f
C4751 a_1029_n88# VSS_SW_b[7] 7.59e-19
C4752 x9.A1 a_13515_627# 5.03e-20
C4753 a_13375_895# a_14096_627# 0.0967f
C4754 a_12607_601# VDD_SW[2] 2.07e-20
C4755 x17.X a_13193_n88# 1.81e-19
C4756 a_12901_601# a_13515_627# 0.0526f
C4757 x9.A1 a_4811_627# 7.9e-19
C4758 VDD a_8140_n62# 7.87e-19
C4759 check[6] a_1555_627# 4.05e-19
C4760 x7.X a_1415_895# 0.00659f
C4761 a_7649_993# a_7967_627# 0.025f
C4762 a_7557_627# a_7733_993# 8.99e-19
C4763 a_8117_601# a_8516_993# 9.41e-19
C4764 a_7369_627# a_8335_627# 2.14e-20
C4765 VDD a_15243_909# 0.0144f
C4766 VDD a_14887_1642# 0.00172f
C4767 ready x30.A 0.00174f
C4768 a_2468_1467# a_2470_90# 1e-19
C4769 a_12680_106# a_12988_212# 0.14f
C4770 a_12447_n62# a_12989_n88# 0.125f
C4771 x2.X a_2566_n88# 0.178f
C4772 a_2566_n88# a_3070_220# 0.00869f
C4773 ready D[6] 0.0519f
C4774 x18.X m1_95_2154# 3.24e-20
C4775 reset a_29_2457# 0.201f
C4776 a_16109_1642# a_16037_1642# 6.64e-19
C4777 a_10596_212# VSS_SW_b[2] 0.0038f
C4778 a_10983_895# VSS_SW[2] 7.52e-21
C4779 VDD x2.X 9.8f
C4780 VDD_SW[2] a_15608_993# 1.08e-20
C4781 D[3] VSS_SW[2] 4.86e-19
C4782 VDD a_4413_2457# 0.228f
C4783 VDD a_3070_220# 0.00671f
C4784 a_10215_601# a_10824_993# 0.00189f
C4785 a_939_2457# a_193_627# 2.84e-21
C4786 x9.X a_2585_627# 1.07e-20
C4787 D[3] a_10041_993# 0.00884f
C4788 x2.X x6.X 2.59e-20
C4789 ready m1_95_1942# 8.93e-20
C4790 a_4811_627# a_6040_993# 0.14f
C4791 D[5] a_6199_895# 0.0296f
C4792 x9.A1 VSS_SW[1] 0.102f
C4793 VDD a_557_993# 0.00586f
C4794 x2.X a_14096_627# 3.85e-19
C4795 a_12901_601# VSS_SW[1] 2.72e-20
C4796 a_13375_895# a_13329_n62# 1.65e-20
C4797 x7.X VDD_SW_b[7] 0.242f
C4798 a_8288_909# VDD_SW_b[4] 9.38e-21
C4799 a_7967_627# a_8335_627# 3.34e-19
C4800 a_5323_2457# a_4811_627# 4.8e-19
C4801 a_3895_1642# x9.X 1.34e-19
C4802 a_8591_895# VSS_SW[3] 7.03e-21
C4803 check[4] m1_95_2154# 0.0352f
C4804 a_11987_627# a_12341_627# 0.0455f
C4805 D[2] a_13216_993# 0.00608f
C4806 a_8204_212# a_9742_n88# 6.15e-19
C4807 a_3333_601# a_3947_627# 0.0526f
C4808 a_3807_895# a_4528_627# 0.0967f
C4809 x9.A1 a_3893_122# 2.28e-20
C4810 VDD_SW_b[3] a_12341_627# 9.3e-21
C4811 a_3039_601# VDD_SW[6] 2.07e-20
C4812 a_15464_909# VDD_SW[1] 2.82e-20
C4813 a_2879_n62# a_3761_n62# 0.00926f
C4814 a_8432_993# m1_95_2154# 4.11e-21
C4815 a_3893_122# a_4338_n62# 0.0369f
C4816 a_3112_106# a_3535_n62# 0.00386f
C4817 a_2566_n88# VSS_SW[5] 4.18e-21
C4818 a_8591_895# m1_95_1942# 8.62e-20
C4819 VDD a_14428_1467# 0.154f
C4820 x7.X check[5] 5.61e-19
C4821 VDD_SW_b[5] a_8205_n88# 2.44e-21
C4822 x11.X a_6539_1315# 1.97e-19
C4823 VDD a_4977_627# 0.694f
C4824 VDD_SW_b[7] a_3420_212# 4.59e-22
C4825 VDD VSS_SW[5] 0.691f
C4826 x14.X VDD_SW[4] 0.308f
C4827 x13.X a_9595_627# 0.00295f
C4828 x2.X a_27_627# 0.352f
C4829 x2.X a_7733_993# 5.31e-19
C4830 x9.A1 a_7649_993# 9.51e-20
C4831 a_14570_1642# VSS_SW[1] 0.00105f
C4832 D[5] VDD_SW_b[5] 0.453f
C4833 VDD_SW_b[4] a_10459_909# 3.15e-21
C4834 x17.X a_14430_90# 0.0273f
C4835 D[7] a_1555_627# 0.00431f
C4836 x9.A1 a_11325_1315# 0.00496f
C4837 check[5] a_3420_212# 3.24e-20
C4838 a_7369_627# a_9949_627# 3.67e-21
C4839 check[3] D[4] 0.462f
C4840 D[7] a_381_627# 0.161f
C4841 a_27_627# a_557_993# 4.45e-20
C4842 VDD_SW_b[4] VSS_SW[3] 0.00248f
C4843 VDD a_9312_627# 0.216f
C4844 check[3] VSS_SW[4] 0.0367f
C4845 a_9646_90# VSS_SW[3] 0.082f
C4846 VDD_SW_b[6] a_4528_627# 0.186f
C4847 a_218_1315# VSS_SW[7] 7.95e-19
C4848 VDD a_15715_627# 1.09e-19
C4849 VDD_SW_b[4] m1_95_1942# 2.11e-20
C4850 x8.X a_473_993# 1.55e-20
C4851 a_12989_n88# a_13126_304# 0.00907f
C4852 a_12447_n62# a_13906_n62# 3.79e-20
C4853 a_12988_212# a_13407_220# 2.46e-19
C4854 a_12153_627# a_12447_n62# 2.38e-19
C4855 a_12607_601# a_12134_n88# 4.37e-19
C4856 a_16109_1642# a_16330_1315# 0.00783f
C4857 a_4149_1642# check[4] 1.58e-19
C4858 a_16109_1642# VDD_SW[1] 0.00494f
C4859 VDD a_5575_627# 0.0101f
C4860 check[4] a_5257_993# 6.52e-20
C4861 a_1757_1642# a_1978_1315# 0.00783f
C4862 a_10459_909# VDD_SW[3] 1.01e-20
C4863 check[0] a_14887_1642# 0.00526f
C4864 x9.A1 a_10596_212# 1.41e-20
C4865 D[1] a_15511_627# 6.11e-19
C4866 a_6199_895# a_8117_601# 1.38e-20
C4867 VDD a_12924_n62# 7.87e-19
C4868 a_9761_627# a_11704_627# 2e-20
C4869 a_2136_627# D[6] 4.35e-19
C4870 check[2] a_10288_106# 8.14e-22
C4871 a_1555_627# a_2419_627# 1.09e-19
C4872 a_6285_122# a_7350_n88# 8e-21
C4873 a_6529_304# a_6730_n62# 8.99e-19
C4874 VDD a_11987_627# 0.448f
C4875 a_5813_n88# a_7896_106# 1.67e-21
C4876 a_5812_212# a_8204_212# 9.5e-22
C4877 VDD_SW[4] a_10680_909# 2.77e-20
C4878 VDD VDD_SW_b[3] 0.266f
C4879 a_720_106# VSS_SW[6] 9.06e-21
C4880 a_1029_n88# a_1143_n62# 2.14e-20
C4881 a_1028_212# a_1369_n62# 0.00134f
C4882 VDD_SW[3] m1_95_1942# 0.0331f
C4883 x2.X check[0] 0.142f
C4884 VDD a_4370_1315# 3.89e-19
C4885 x2.X a_10007_1315# 3.2e-19
C4886 D[5] a_5504_106# 8.77e-19
C4887 a_4811_627# a_5812_212# 6.99e-20
C4888 a_647_601# a_941_601# 0.199f
C4889 a_193_627# a_1415_895# 0.0494f
C4890 a_2136_627# m1_95_1942# 2.45e-20
C4891 a_11987_627# a_14096_627# 1.75e-19
C4892 a_8432_993# a_8539_627# 0.00707f
C4893 a_8591_895# VDD_SW[4] 0.00356f
C4894 x15.X VSS_SW_b[2] 0.0171f
C4895 a_1256_993# m1_95_1942# 5.78e-21
C4896 x14.X a_10073_1289# 1.5e-19
C4897 x2.X a_3369_304# 0.00168f
C4898 a_1503_1642# x8.X 1.14e-20
C4899 x2.X VDD_SW[7] 0.0768f
C4900 VDD a_13929_1642# 0.00177f
C4901 VDD_SW_b[5] a_8117_601# 5.19e-20
C4902 x9.A1 a_941_601# 0.00103f
C4903 x2.X a_891_909# 0.00138f
C4904 x2.X a_10288_106# 0.0385f
C4905 x20.X a_14839_n62# 0.002f
C4906 VDD_SW_b[1] a_14839_n62# 5.21e-19
C4907 a_14428_1467# check[0] 0.318f
C4908 VDD_SW[2] D[1] 4.41e-19
C4909 a_193_627# VDD_SW_b[7] 0.0022f
C4910 a_1256_993# a_1340_993# 0.00857f
C4911 check[4] a_5289_1289# 0.247f
C4912 a_9742_n88# a_10596_212# 0.0319f
C4913 VDD_SW_b[4] VDD_SW[4] 3.64e-19
C4914 a_12924_n62# a_13329_n62# 2.46e-21
C4915 reset check[6] 1.32e-20
C4916 x2.X a_5431_601# 0.2f
C4917 x9.A1 a_11313_n62# 5.47e-21
C4918 x9.A1 a_9949_627# 4.11e-19
C4919 a_10983_895# a_13216_993# 1.86e-21
C4920 a_10509_601# a_12341_627# 2.42e-20
C4921 VDD a_15853_122# 0.313f
C4922 x18.X a_13936_1315# 3.11e-20
C4923 a_2585_627# a_3625_n88# 8.75e-19
C4924 check[2] a_10824_993# 2.78e-19
C4925 a_3333_601# a_3112_106# 3.46e-19
C4926 a_3039_601# a_3421_n88# 0.00322f
C4927 a_3807_895# a_2879_n62# 0.00219f
C4928 check[4] a_4958_n88# 5.26e-19
C4929 VDD a_76_1467# 0.153f
C4930 x2.X a_8731_627# 0.0151f
C4931 x9.A1 a_2927_1642# 5.26e-19
C4932 VDD a_3648_993# 0.219f
C4933 x9.A1 a_16097_n62# 5.47e-21
C4934 a_76_1467# x6.X 0.0876f
C4935 a_12433_993# m1_95_2154# 1.86e-20
C4936 a_11071_1642# m1_95_1942# 2.26e-19
C4937 a_3895_1642# a_3625_n88# 4.63e-19
C4938 x2.X a_5365_627# 3.94e-19
C4939 a_4977_627# a_5431_601# 0.117f
C4940 a_12178_1315# VSS_SW[2] 7.96e-19
C4941 a_5431_601# VSS_SW[5] 6.28e-19
C4942 x9.A1 x15.X 6.84e-19
C4943 x15.X a_12901_601# 4.02e-21
C4944 VDD a_174_n88# 0.722f
C4945 VSS_SW[7] m1_95_1942# 0.0287f
C4946 VDD_SW_b[6] a_2879_n62# 5.22e-19
C4947 a_6285_1642# a_6199_895# 5.55e-19
C4948 a_15855_1642# m1_95_2154# 1.04e-19
C4949 x2.X a_10824_993# 0.187f
C4950 a_12038_90# a_12989_n88# 9.87e-21
C4951 a_11015_220# VSS_SW_b[2] 4.16e-21
C4952 a_10596_212# a_12553_n62# 1.09e-19
C4953 a_76_1467# a_27_627# 5.32e-19
C4954 a_14825_993# a_15293_601# 0.0633f
C4955 a_14857_1289# a_14545_627# 0.00323f
C4956 a_7254_90# a_7663_n62# 4.24e-20
C4957 a_14545_627# a_15608_993# 0.0334f
C4958 x17.X D[1] 2.04e-19
C4959 a_6539_1642# VDD_SW[5] 0.00492f
C4960 a_1745_304# VSS_SW[6] 6.59e-21
C4961 VDD_SW_b[3] a_10288_106# 5.24e-19
C4962 a_1029_n88# VSS_SW_b[6] 0.00485f
C4963 a_593_n62# a_964_n62# 4.19e-20
C4964 a_5725_601# a_5896_909# 0.00652f
C4965 a_14526_n88# a_15030_220# 0.00869f
C4966 a_5431_601# a_5575_627# 0.0697f
C4967 a_9949_627# a_9742_n88# 3.32e-19
C4968 a_5365_627# VSS_SW[5] 3.8e-19
C4969 VSS_SW[1] a_15585_n88# 9.92e-21
C4970 a_12989_n88# m1_95_1942# 1.16e-21
C4971 D[5] a_6231_220# 7.13e-19
C4972 a_9595_627# a_10596_212# 6.99e-20
C4973 x8.X a_2585_627# 0.00315f
C4974 VDD a_10509_601# 0.481f
C4975 a_2897_1289# a_2566_n88# 5.67e-21
C4976 x9.A1 a_2468_1467# 0.197f
C4977 D[2] VSS_SW_b[1] 2.02e-19
C4978 a_27_627# a_174_n88# 0.00176f
C4979 a_12465_1289# a_12680_106# 5.3e-21
C4980 a_7252_1467# a_7394_1642# 0.00557f
C4981 VDD_SW_b[2] a_12447_n62# 5.22e-19
C4982 VDD a_2897_1289# 0.221f
C4983 D[6] VSS_SW_b[5] 2.03e-19
C4984 x16.X a_12038_90# 0.00259f
C4985 x8.X a_3895_1642# 1.98e-20
C4986 VDD a_15316_n62# 9.38e-19
C4987 VDD_SW[5] a_8288_909# 2.77e-20
C4988 D[4] VSS_SW_b[4] 5.32e-19
C4989 VSS_SW[4] VSS_SW_b[4] 0.0072f
C4990 D[6] a_3333_601# 0.019f
C4991 VDD check[1] 1.75f
C4992 a_2419_627# a_3807_895# 0.0321f
C4993 x15.X a_9742_n88# 1.53e-21
C4994 x10.X VDD_SW[6] 0.305f
C4995 x9.X a_4811_627# 0.00299f
C4996 a_12036_1467# m1_95_2154# 8.35e-20
C4997 x16.X m1_95_1942# 6.66e-20
C4998 a_5675_909# VDD_SW_b[5] 3.01e-21
C4999 check[0] a_15853_122# 6.43e-20
C5000 a_76_1467# a_218_1642# 0.00557f
C5001 x17.X a_15380_212# 1.68e-21
C5002 x13.X a_7896_106# 2.38e-20
C5003 a_3333_601# m1_95_1942# 4.09e-20
C5004 a_3807_895# m1_95_2154# 5.86e-20
C5005 reset m1_95_2154# 5.5e-20
C5006 x9.A1 a_6017_n88# 1.66e-20
C5007 VDD_SW[6] D[5] 4.59e-19
C5008 x2.X a_1757_1642# 5.76e-19
C5009 a_3839_220# VSS_SW_b[5] 3.96e-21
C5010 a_4862_90# a_5813_n88# 9.87e-21
C5011 a_3420_212# a_5377_n62# 1.09e-19
C5012 a_12988_212# a_14526_n88# 6.15e-19
C5013 x12.X a_6199_895# 0.00864f
C5014 x2.X a_2773_627# 0.0014f
C5015 VDD a_7203_627# 0.405f
C5016 x9.A1 a_3039_601# 2.81e-20
C5017 a_16488_627# m1_95_2154# 1.66e-20
C5018 x11.X a_5813_n88# 0.0189f
C5019 VDD a_6153_n62# 0.0323f
C5020 D[6] a_4064_909# 8.06e-19
C5021 a_2419_627# VDD_SW_b[6] 1.12e-19
C5022 VDD_SW[5] m1_95_1942# 0.0331f
C5023 a_10983_895# D[2] 2.17e-19
C5024 a_10824_993# a_11987_627# 7.46e-20
C5025 VDD_SW[7] a_3648_993# 1.08e-20
C5026 D[3] D[2] 0.00189f
C5027 a_10824_993# VDD_SW_b[3] 5e-20
C5028 x2.X a_487_n62# 0.374f
C5029 x9.X a_3893_122# 2.77e-19
C5030 VDD_SW_b[6] m1_95_2154# 1.35e-20
C5031 a_9595_627# a_9949_627# 0.0455f
C5032 x9.A1 a_6339_627# 4.53e-20
C5033 a_12153_627# m1_95_1942# 3.82e-20
C5034 check[3] a_8545_n62# 5.64e-21
C5035 a_2136_627# a_1028_212# 6.63e-19
C5036 a_6040_993# a_6017_n88# 1.86e-19
C5037 a_6199_895# a_6285_122# 4.53e-22
C5038 check[1] a_13329_n62# 5.49e-21
C5039 a_1415_895# a_1029_n88# 6.35e-19
C5040 VDD a_1166_304# 0.0164f
C5041 a_941_601# a_1233_n88# 0.00251f
C5042 a_1256_993# a_1028_212# 8.94e-21
C5043 check[3] m1_95_2154# 0.0352f
C5044 a_8933_1642# x14.X 8.08e-19
C5045 a_12607_601# a_12751_627# 0.0697f
C5046 a_12901_601# a_13072_909# 0.00652f
C5047 x12.X VDD_SW_b[5] 7.21e-19
C5048 x11.X a_6920_627# 0.0338f
C5049 a_4149_1642# a_3807_895# 0.00232f
C5050 a_3333_601# a_5725_601# 9.37e-21
C5051 a_2585_627# a_5165_627# 3.67e-21
C5052 a_3807_895# a_5257_993# 8e-21
C5053 a_10073_1289# a_11071_1642# 0.0146f
C5054 a_9786_1315# D[3] 7.54e-19
C5055 a_7203_627# a_7733_993# 4.45e-20
C5056 D[4] a_7557_627# 0.161f
C5057 a_7557_627# VSS_SW[4] 0.00595f
C5058 x15.X a_9595_627# 2.67e-20
C5059 x2.X a_10734_304# 0.00334f
C5060 a_7896_106# a_8204_212# 0.14f
C5061 a_7663_n62# a_8205_n88# 0.125f
C5062 a_15767_895# m1_95_1942# 8.62e-20
C5063 x9.A1 VSS_SW_b[7] 1.46e-19
C5064 VDD_SW_b[7] a_3504_909# 1.97e-21
C5065 a_4363_1642# VDD_SW[6] 5.38e-19
C5066 a_2470_90# VSS_SW_b[6] 0.19f
C5067 VSS_SW[6] a_3112_106# 4.63e-19
C5068 D[1] a_14545_627# 0.168f
C5069 x9.A1 a_13715_1315# 0.00499f
C5070 a_5725_601# VDD_SW[5] 1.79e-19
C5071 a_14379_627# a_14999_601# 0.149f
C5072 a_6040_993# a_6339_627# 0.0256f
C5073 a_7252_1467# a_7350_n88# 6.87e-20
C5074 VSS_SW_b[3] a_10161_n62# 0.00335f
C5075 a_10596_212# VSS_SW[2] 0.0872f
C5076 check[1] check[0] 0.00509f
C5077 a_10801_n88# a_10711_n62# 9.75e-19
C5078 a_10597_n88# a_10937_n62# 6.04e-20
C5079 VDD_SW_b[5] a_6285_122# 0.00447f
C5080 VDD_SW_b[2] a_14999_601# 1.99e-20
C5081 check[2] D[4] 6.03e-20
C5082 a_10215_601# a_10597_n88# 0.00322f
C5083 VDD_SW_b[7] a_1029_n88# 0.0406f
C5084 a_10509_601# a_10288_106# 3.46e-19
C5085 a_10983_895# a_10055_n62# 0.00219f
C5086 D[3] a_10055_n62# 0.00258f
C5087 VDD a_10246_220# 0.00412f
C5088 a_4149_1642# VDD_SW_b[6] 1.79e-19
C5089 x2.X a_5462_220# 0.00279f
C5090 VDD_SW_b[6] a_5257_993# 8.2e-21
C5091 x2.X a_12851_909# 0.00138f
C5092 a_1503_1642# a_1501_122# 1.57e-21
C5093 a_6539_1642# a_6753_1642# 0.00557f
C5094 a_29_2457# x2.X 3.13e-19
C5095 a_14857_1289# x20.X 1.7e-20
C5096 a_305_2457# a_939_2457# 8.52e-20
C5097 a_9644_1467# VSS_SW[3] 0.0274f
C5098 a_15608_993# VDD_SW_b[1] 5.61e-20
C5099 a_8933_1642# a_8591_895# 0.00232f
C5100 a_6456_909# VDD_SW[5] 2.12e-20
C5101 a_9644_1467# m1_95_1942# 1.97e-19
C5102 VDD a_12341_627# 0.125f
C5103 VSS_SW_b[1] a_15495_n62# 5.24e-19
C5104 a_15853_122# a_15721_n62# 0.025f
C5105 VDD a_6760_1315# 0.00108f
C5106 x2.X a_14933_627# 3.94e-19
C5107 a_14545_627# a_15380_212# 1.02e-19
C5108 x2.X a_12399_1315# 3.21e-19
C5109 a_14999_601# a_15072_106# 1.01e-19
C5110 a_15293_601# a_14526_n88# 0.00259f
C5111 a_14825_993# a_14839_n62# 2.63e-19
C5112 x2.X D[4] 0.185f
C5113 x9.A1 VDD_SW[2] 0.0329f
C5114 x2.X VSS_SW[4] 0.0643f
C5115 a_4860_1467# VDD_SW[6] 0.00487f
C5116 a_12901_601# VDD_SW[2] 1.75e-19
C5117 VSS_SW[5] a_5462_220# 4.26e-19
C5118 a_5812_212# a_6017_n88# 0.15f
C5119 a_5271_n62# VSS_SW_b[5] 0.0142f
C5120 a_13216_993# a_13515_627# 0.0256f
C5121 a_78_90# a_1029_n88# 9.87e-21
C5122 a_1978_1315# D[7] 0.0012f
C5123 VSS_SW[7] a_1028_212# 5.9e-22
C5124 x2.X a_4528_627# 3.85e-19
C5125 a_4413_2457# a_4528_627# 1.19e-21
C5126 x11.X a_6730_n62# 0.00162f
C5127 VDD a_15692_993# 0.00308f
C5128 VDD a_16323_1642# 0.00177f
C5129 a_12988_212# a_12989_n88# 0.785f
C5130 a_12134_n88# VSS_SW_b[2] 0.135f
C5131 a_12447_n62# a_13461_122# 0.0633f
C5132 a_8933_1642# VDD_SW_b[4] 1.9e-19
C5133 a_12680_106# a_13193_n88# 0.00189f
C5134 a_7649_993# a_7896_106# 4.96e-20
C5135 a_7369_627# a_8205_n88# 1.27e-19
C5136 a_8117_601# a_7663_n62# 3.74e-20
C5137 a_7823_601# a_8204_212# 4.51e-19
C5138 x2.X a_1447_220# 9.51e-19
C5139 a_10801_n88# VSS_SW_b[2] 5.04e-20
C5140 D[6] VSS_SW[6] 0.118f
C5141 VDD_SW[2] a_14909_993# 6.61e-21
C5142 x18.X a_14999_601# 2.4e-20
C5143 D[5] a_7369_627# 6.4e-21
C5144 a_9761_627# a_10459_909# 0.00276f
C5145 a_10509_601# a_10824_993# 0.13f
C5146 a_10041_993# a_9949_627# 0.0369f
C5147 a_4977_627# VSS_SW[4] 5.07e-21
C5148 check[4] a_7681_1289# 4.13e-21
C5149 a_6339_627# a_5812_212# 7.07e-21
C5150 D[3] a_10983_895# 0.0294f
C5151 a_10359_627# VSS_SW[3] 0.0012f
C5152 VDD a_2566_n88# 0.72f
C5153 ready x7.X 3.39e-21
C5154 a_9761_627# VSS_SW[3] 0.023f
C5155 x2.X a_13323_627# 0.00111f
C5156 VSS_SW[6] m1_95_1942# 0.033f
C5157 a_4528_627# a_4977_627# 5.39e-19
C5158 a_9761_627# m1_95_1942# 3.82e-20
C5159 a_10215_601# m1_95_2154# 2.34e-20
C5160 a_4528_627# VSS_SW[5] 0.00162f
C5161 VDD_SW_b[6] a_4958_n88# 5.91e-19
C5162 a_4689_2457# VDD_SW[6] 0.0305f
C5163 a_11987_627# a_12851_909# 2.46e-19
C5164 D[2] a_12517_993# 8.11e-19
C5165 D[4] a_9312_627# 0.00232f
C5166 x15.X VSS_SW[2] 0.138f
C5167 VDD_SW_b[3] a_12851_909# 2.62e-21
C5168 VDD_SW_b[4] a_7350_n88# 3.21e-19
C5169 a_9644_1467# VDD_SW[4] 0.00484f
C5170 a_2585_627# a_3183_627# 6.04e-20
C5171 a_8204_212# a_8623_220# 2.46e-19
C5172 a_7663_n62# a_9122_n62# 3.79e-20
C5173 VDD x6.X 0.428f
C5174 a_3333_601# a_3283_909# 1.21e-20
C5175 a_8205_n88# a_8342_304# 0.00907f
C5176 VDD a_14096_627# 0.196f
C5177 a_3421_n88# VSS_SW_b[6] 7.59e-19
C5178 VSS_SW[6] a_3839_220# 6.42e-21
C5179 a_3625_n88# a_3893_122# 0.206f
C5180 a_15316_n62# a_15721_n62# 2.46e-21
C5181 a_14379_627# m1_95_1942# 5.19e-20
C5182 VDD_SW_b[2] m1_95_1942# 2.87e-20
C5183 VDD_SW_b[5] a_5377_n62# 4.78e-19
C5184 a_13461_1642# m1_95_1942# 2.26e-19
C5185 check[5] VDD_SW[6] 0.00393f
C5186 x3.X a_941_601# 6.38e-19
C5187 a_13715_1642# VDD_SW[2] 0.00502f
C5188 VDD_SW_b[7] a_2470_90# 0.00345f
C5189 a_12178_1315# D[2] 7.54e-19
C5190 x9.A1 x17.X 6.87e-19
C5191 x17.X a_12901_601# 1.26e-19
C5192 VDD_SW[6] a_5675_909# 2.16e-20
C5193 check[5] a_2470_90# 2.5e-20
C5194 a_174_n88# a_487_n62# 0.245f
C5195 VDD a_27_627# 0.461f
C5196 VDD a_7733_993# 0.00422f
C5197 a_8677_122# VSS_SW[3] 6.66e-20
C5198 VSS_SW_b[4] a_8545_n62# 5.35e-19
C5199 a_13193_n88# a_13407_220# 0.0104f
C5200 a_12989_n88# a_13705_304# 0.0018f
C5201 a_12988_212# a_13906_n62# 0.0453f
C5202 x9.A1 a_12134_n88# 7.34e-19
C5203 a_12901_601# a_12134_n88# 0.00259f
C5204 a_12153_627# a_12988_212# 1.02e-19
C5205 a_12433_993# a_12447_n62# 2.63e-19
C5206 a_12607_601# a_12680_106# 1.01e-19
C5207 a_7823_601# a_7649_993# 0.206f
C5208 x6.X a_27_627# 0.236f
C5209 a_7369_627# a_8117_601# 0.126f
C5210 a_6539_1642# check[4] 0.318f
C5211 a_10359_627# a_10931_627# 2.46e-21
C5212 check[0] a_16323_1642# 0.00688f
C5213 D[1] VDD_SW_b[1] 0.454f
C5214 x9.A1 a_10801_n88# 3.88e-20
C5215 x20.X D[1] 0.086f
C5216 x9.A1 x10.X 9.2e-19
C5217 VDD a_13329_n62# 0.0301f
C5218 check[2] a_10597_n88# 1.93e-20
C5219 a_15072_106# m1_95_1942# 4.96e-22
C5220 x13.X a_10055_n62# 4.41e-20
C5221 x10.X a_5002_1315# 8.34e-19
C5222 x9.A1 a_8205_n88# 5.63e-21
C5223 VSS_SW_b[5] a_5950_304# 3.57e-20
C5224 a_5813_n88# a_6730_n62# 0.189f
C5225 a_5812_212# a_7254_90# 0.00102f
C5226 a_6017_n88# a_6529_304# 6.69e-20
C5227 a_5271_n62# a_5748_n62# 1.96e-20
C5228 a_5504_106# a_5377_n62# 0.0256f
C5229 x2.X check[6] 0.193f
C5230 VDD_SW[4] a_9761_627# 9.25e-19
C5231 a_1233_n88# VSS_SW_b[7] 9.21e-19
C5232 x9.A1 D[5] 0.309f
C5233 x7.X a_2136_627# 0.0338f
C5234 D[2] a_13515_627# 0.00431f
C5235 VDD a_8319_n62# 0.00521f
C5236 x11.X a_8204_212# 8.4e-22
C5237 a_4811_627# a_4862_90# 6.13e-19
C5238 a_5002_1315# D[5] 7.54e-19
C5239 a_7823_601# a_8335_627# 9.75e-19
C5240 a_7649_993# a_7757_627# 0.00807f
C5241 a_29_2457# a_76_1467# 1.6e-20
C5242 a_8117_601# a_7967_627# 0.00926f
C5243 a_8432_993# a_8288_909# 0.00412f
C5244 a_7369_627# a_8848_909# 7.17e-20
C5245 VDD a_218_1642# 0.00433f
C5246 x11.X a_4811_627# 2.67e-20
C5247 VDD check[0] 1.69f
C5248 x2.X a_2879_n62# 0.371f
C5249 a_2879_n62# a_3070_220# 3.3e-19
C5250 reset x3.A 0.00421f
C5251 x18.X m1_95_1942# 5.57e-20
C5252 x2.X a_10597_n88# 0.0213f
C5253 VDD_SW_b[1] a_15380_212# 0.0417f
C5254 x20.X a_15380_212# 0.245f
C5255 x30.A check[4] 0.00702f
C5256 a_11015_220# VSS_SW[2] 1.76e-20
C5257 a_13715_1642# x17.X 0.0841f
C5258 VDD a_3369_304# 0.00298f
C5259 a_939_2457# a_647_601# 2.7e-21
C5260 ready a_193_627# 6.76e-21
C5261 check[4] D[6] 5.94e-20
C5262 VDD VDD_SW[7] 0.474f
C5263 D[5] a_6040_993# 0.00609f
C5264 a_4811_627# a_5165_627# 0.0455f
C5265 a_14526_n88# a_14839_n62# 0.245f
C5266 check[4] a_5002_1642# 0.00688f
C5267 VDD a_891_909# 0.0143f
C5268 VDD a_10288_106# 0.356f
C5269 a_5323_2457# D[5] 0.038f
C5270 a_13705_304# a_13906_n62# 8.99e-19
C5271 D[2] VSS_SW[1] 4.85e-19
C5272 check[4] m1_95_1942# 0.034f
C5273 x9.A1 VSS_SW_b[6] 2.15e-19
C5274 a_2865_993# VDD_SW[6] 4.17e-21
C5275 a_8205_n88# a_9742_n88# 1.98e-19
C5276 a_3807_895# a_3947_627# 0.0383f
C5277 a_8204_212# a_10055_n62# 2.62e-19
C5278 a_3333_601# a_3755_627# 1.96e-20
C5279 a_939_2457# x9.A1 0.00366f
C5280 a_3420_212# a_3535_n62# 0.00272f
C5281 a_8432_993# m1_95_1942# 5.78e-21
C5282 a_3112_106# a_3761_n62# 0.00316f
C5283 a_2879_n62# VSS_SW[5] 1.64e-20
C5284 a_10073_1289# a_9761_627# 0.00323f
C5285 VDD a_5431_601# 0.343f
C5286 x13.X D[3] 2.06e-19
C5287 VDD_SW_b[7] a_3421_n88# 2.44e-21
C5288 x2.X D[7] 0.238f
C5289 x9.A1 a_8117_601# 9.51e-19
C5290 x2.X a_8067_909# 0.00138f
C5291 a_13375_895# m1_95_2154# 5.86e-20
C5292 m1_95_1942# VSS 1.29f $ **FLOATING
C5293 m1_95_2154# VSS 1.43f $ **FLOATING
C5294 a_16097_n62# VSS 0.00289f
C5295 a_15721_n62# VSS 0.189f
C5296 a_15495_n62# VSS 0.0154f
C5297 a_15316_n62# VSS 0.00254f
C5298 a_14945_n62# VSS 0.175f
C5299 a_16298_n62# VSS 0.106f
C5300 a_16097_304# VSS 0.00178f
C5301 a_15799_220# VSS 0.00285f
C5302 a_15518_304# VSS 0.00171f
C5303 a_15329_304# VSS 3.26e-21
C5304 a_15030_220# VSS 0.00102f
C5305 a_13705_n62# VSS 0.00323f
C5306 VSS_SW_b[1] VSS 0.416f
C5307 a_15853_122# VSS 0.298f
C5308 a_15585_n88# VSS 0.315f
C5309 a_15381_n88# VSS 0.398f
C5310 a_15380_212# VSS 0.86f
C5311 a_15072_106# VSS 0.261f
C5312 a_14839_n62# VSS 0.405f
C5313 a_14526_n88# VSS 0.483f
C5314 VSS_SW[1] VSS 0.617f
C5315 a_13329_n62# VSS 0.188f
C5316 a_13103_n62# VSS 0.0145f
C5317 a_12924_n62# VSS 0.00268f
C5318 a_12553_n62# VSS 0.176f
C5319 a_14430_90# VSS 0.244f
C5320 a_13906_n62# VSS 0.108f
C5321 a_13705_304# VSS 0.00223f
C5322 a_13407_220# VSS 0.00199f
C5323 a_13126_304# VSS 0.00612f
C5324 a_12937_304# VSS 5.68e-19
C5325 a_12638_220# VSS 5.97e-19
C5326 a_11313_n62# VSS 0.00265f
C5327 VSS_SW_b[2] VSS 0.422f
C5328 a_13461_122# VSS 0.304f
C5329 a_13193_n88# VSS 0.324f
C5330 a_12989_n88# VSS 0.412f
C5331 a_12988_212# VSS 0.808f
C5332 a_12680_106# VSS 0.272f
C5333 a_12447_n62# VSS 0.42f
C5334 a_12134_n88# VSS 0.489f
C5335 VSS_SW[2] VSS 0.631f
C5336 a_10937_n62# VSS 0.186f
C5337 a_10711_n62# VSS 0.0147f
C5338 a_10532_n62# VSS 0.00271f
C5339 a_10161_n62# VSS 0.179f
C5340 a_12038_90# VSS 0.241f
C5341 a_11514_n62# VSS 0.105f
C5342 a_11313_304# VSS 6.83e-19
C5343 a_11015_220# VSS 0.00377f
C5344 a_10734_304# VSS 0.00775f
C5345 a_10545_304# VSS 5.65e-19
C5346 a_10246_220# VSS 0.00255f
C5347 a_8921_n62# VSS 0.00232f
C5348 VSS_SW_b[3] VSS 0.435f
C5349 a_11069_122# VSS 0.292f
C5350 a_10801_n88# VSS 0.326f
C5351 a_10597_n88# VSS 0.384f
C5352 a_10596_212# VSS 0.793f
C5353 a_10288_106# VSS 0.275f
C5354 a_10055_n62# VSS 0.439f
C5355 a_9742_n88# VSS 0.506f
C5356 VSS_SW[3] VSS 0.705f
C5357 a_8545_n62# VSS 0.184f
C5358 a_8319_n62# VSS 0.0133f
C5359 a_8140_n62# VSS 0.00268f
C5360 a_7769_n62# VSS 0.18f
C5361 a_9646_90# VSS 0.246f
C5362 a_9122_n62# VSS 0.103f
C5363 a_8921_304# VSS 9.36e-20
C5364 a_8623_220# VSS 0.00162f
C5365 a_8342_304# VSS 0.00491f
C5366 a_8153_304# VSS 4.85e-19
C5367 a_7854_220# VSS 0.00297f
C5368 a_6529_n62# VSS 0.0024f
C5369 VSS_SW_b[4] VSS 0.45f
C5370 a_8677_122# VSS 0.283f
C5371 a_8409_n88# VSS 0.309f
C5372 a_8205_n88# VSS 0.362f
C5373 a_8204_212# VSS 0.784f
C5374 a_7896_106# VSS 0.275f
C5375 a_7663_n62# VSS 0.427f
C5376 a_7350_n88# VSS 0.502f
C5377 VSS_SW[4] VSS 0.863f
C5378 a_6153_n62# VSS 0.184f
C5379 a_5927_n62# VSS 0.0128f
C5380 a_5748_n62# VSS 0.00239f
C5381 a_5377_n62# VSS 0.176f
C5382 a_7254_90# VSS 0.253f
C5383 a_6730_n62# VSS 0.103f
C5384 a_6529_304# VSS 1.67e-19
C5385 a_6231_220# VSS 0.00134f
C5386 a_5950_304# VSS 0.00146f
C5387 a_5761_304# VSS 4.44e-20
C5388 a_5462_220# VSS 0.00158f
C5389 a_4137_n62# VSS 0.00302f
C5390 VSS_SW_b[5] VSS 0.453f
C5391 a_6285_122# VSS 0.286f
C5392 a_6017_n88# VSS 0.308f
C5393 a_5813_n88# VSS 0.361f
C5394 a_5812_212# VSS 0.789f
C5395 a_5504_106# VSS 0.263f
C5396 a_5271_n62# VSS 0.409f
C5397 a_4958_n88# VSS 0.486f
C5398 VSS_SW[5] VSS 0.898f
C5399 a_3761_n62# VSS 0.184f
C5400 a_3535_n62# VSS 0.013f
C5401 a_3356_n62# VSS 0.00239f
C5402 a_2985_n62# VSS 0.175f
C5403 a_4862_90# VSS 0.261f
C5404 a_4338_n62# VSS 0.107f
C5405 a_4137_304# VSS 0.00202f
C5406 a_3839_220# VSS 0.00123f
C5407 a_3558_304# VSS 0.00178f
C5408 a_3369_304# VSS 2.18e-20
C5409 a_3070_220# VSS 9.42e-19
C5410 a_1745_n62# VSS 0.00344f
C5411 VSS_SW_b[6] VSS 0.419f
C5412 a_3893_122# VSS 0.298f
C5413 a_3625_n88# VSS 0.316f
C5414 a_3421_n88# VSS 0.385f
C5415 a_3420_212# VSS 0.802f
C5416 a_3112_106# VSS 0.264f
C5417 a_2879_n62# VSS 0.402f
C5418 a_2566_n88# VSS 0.479f
C5419 VSS_SW[6] VSS 0.656f
C5420 a_1369_n62# VSS 0.187f
C5421 a_1143_n62# VSS 0.0143f
C5422 a_964_n62# VSS 0.00251f
C5423 a_593_n62# VSS 0.177f
C5424 a_2470_90# VSS 0.249f
C5425 a_1946_n62# VSS 0.11f
C5426 a_1745_304# VSS 0.00198f
C5427 a_1447_220# VSS 0.00335f
C5428 a_1166_304# VSS 0.00824f
C5429 a_977_304# VSS 1.42e-19
C5430 a_678_220# VSS 4.32e-19
C5431 VSS_SW_b[7] VSS 0.453f
C5432 a_1501_122# VSS 0.301f
C5433 a_1233_n88# VSS 0.325f
C5434 a_1029_n88# VSS 0.4f
C5435 a_1028_212# VSS 0.812f
C5436 a_720_106# VSS 0.264f
C5437 a_487_n62# VSS 0.416f
C5438 a_174_n88# VSS 0.479f
C5439 VSS_SW[7] VSS 0.939f
C5440 a_78_90# VSS 0.25f
C5441 VDD_SW[1] VSS 1.04f
C5442 a_15715_627# VSS 0.00255f
C5443 a_15907_627# VSS 0.178f
C5444 a_16488_627# VSS 0.267f
C5445 VDD_SW_b[1] VSS 0.56f
C5446 a_16024_909# VSS 0.00378f
C5447 a_15511_627# VSS 0.011f
C5448 a_14933_627# VSS 0.00175f
C5449 a_15143_627# VSS 0.176f
C5450 a_15692_993# VSS 6.43e-19
C5451 a_15464_909# VSS 8.85e-19
C5452 a_14909_993# VSS 8.26e-21
C5453 a_14733_627# VSS 0.101f
C5454 a_15608_993# VSS 0.263f
C5455 a_15767_895# VSS 0.501f
C5456 a_15293_601# VSS 0.415f
C5457 a_14825_993# VSS 0.258f
C5458 a_14999_601# VSS 0.278f
C5459 a_14545_627# VSS 0.316f
C5460 D[1] VSS 1.98f
C5461 a_14379_627# VSS 0.708f
C5462 VDD_SW[2] VSS 0.444f
C5463 a_13323_627# VSS 0.00318f
C5464 a_13515_627# VSS 0.182f
C5465 a_14096_627# VSS 0.256f
C5466 VDD_SW_b[2] VSS 0.561f
C5467 a_13632_909# VSS 0.00125f
C5468 a_13119_627# VSS 0.0165f
C5469 a_12541_627# VSS 0.00181f
C5470 a_12751_627# VSS 0.186f
C5471 a_13300_993# VSS 0.00208f
C5472 a_13072_909# VSS 0.00954f
C5473 a_12851_909# VSS 0.00313f
C5474 a_12517_993# VSS 6.46e-20
C5475 a_12341_627# VSS 0.1f
C5476 a_13216_993# VSS 0.28f
C5477 a_13375_895# VSS 0.484f
C5478 a_12901_601# VSS 0.439f
C5479 a_12433_993# VSS 0.263f
C5480 a_12607_601# VSS 0.302f
C5481 a_12153_627# VSS 0.339f
C5482 D[2] VSS 1.98f
C5483 a_11987_627# VSS 0.733f
C5484 VDD_SW[3] VSS 0.389f
C5485 a_10931_627# VSS 0.00328f
C5486 a_11123_627# VSS 0.177f
C5487 a_11704_627# VSS 0.222f
C5488 VDD_SW_b[3] VSS 0.463f
C5489 a_11240_909# VSS 0.00216f
C5490 a_10727_627# VSS 0.0173f
C5491 a_10149_627# VSS 0.00288f
C5492 a_10359_627# VSS 0.187f
C5493 a_10908_993# VSS 0.00101f
C5494 a_10680_909# VSS 0.00839f
C5495 a_10459_909# VSS 0.00373f
C5496 a_10125_993# VSS 0.00144f
C5497 a_9949_627# VSS 0.111f
C5498 a_10824_993# VSS 0.282f
C5499 a_10983_895# VSS 0.48f
C5500 a_10509_601# VSS 0.411f
C5501 a_10041_993# VSS 0.294f
C5502 a_10215_601# VSS 0.314f
C5503 a_9761_627# VSS 0.374f
C5504 D[3] VSS 1.84f
C5505 a_9595_627# VSS 0.764f
C5506 VDD_SW[4] VSS 0.388f
C5507 a_8539_627# VSS 0.00192f
C5508 a_8731_627# VSS 0.166f
C5509 a_9312_627# VSS 0.224f
C5510 VDD_SW_b[4] VSS 0.457f
C5511 a_8848_909# VSS 3.03e-19
C5512 a_8335_627# VSS 0.0129f
C5513 a_7757_627# VSS 0.00266f
C5514 a_7967_627# VSS 0.186f
C5515 a_8288_909# VSS 0.0032f
C5516 a_8067_909# VSS 0.00505f
C5517 a_7733_993# VSS 0.00136f
C5518 a_7557_627# VSS 0.116f
C5519 a_8432_993# VSS 0.243f
C5520 a_8591_895# VSS 0.442f
C5521 a_8117_601# VSS 0.377f
C5522 a_7649_993# VSS 0.297f
C5523 a_7823_601# VSS 0.314f
C5524 a_7369_627# VSS 0.384f
C5525 D[4] VSS 1.77f
C5526 a_7203_627# VSS 0.772f
C5527 VDD_SW[5] VSS 0.537f
C5528 a_6147_627# VSS 0.00193f
C5529 a_6339_627# VSS 0.166f
C5530 a_6920_627# VSS 0.236f
C5531 VDD_SW_b[5] VSS 0.463f
C5532 a_6456_909# VSS 3.6e-20
C5533 a_5943_627# VSS 0.0108f
C5534 a_5365_627# VSS 0.00259f
C5535 a_5575_627# VSS 0.177f
C5536 a_6124_993# VSS 5.98e-20
C5537 a_5896_909# VSS 6.28e-19
C5538 a_5341_993# VSS 0.00132f
C5539 a_5165_627# VSS 0.116f
C5540 a_6040_993# VSS 0.24f
C5541 a_6199_895# VSS 0.439f
C5542 a_5725_601# VSS 0.359f
C5543 a_5257_993# VSS 0.278f
C5544 a_5431_601# VSS 0.281f
C5545 a_4977_627# VSS 0.363f
C5546 D[5] VSS 1.69f
C5547 a_4811_627# VSS 0.751f
C5548 VDD_SW[6] VSS 0.55f
C5549 a_3755_627# VSS 0.00192f
C5550 a_3947_627# VSS 0.175f
C5551 a_4528_627# VSS 0.256f
C5552 VDD_SW_b[6] VSS 0.558f
C5553 a_4064_909# VSS 0.00152f
C5554 a_3551_627# VSS 0.0108f
C5555 a_2973_627# VSS 0.00172f
C5556 a_3183_627# VSS 0.176f
C5557 a_3732_993# VSS 4.7e-20
C5558 a_3504_909# VSS 5.82e-19
C5559 a_2949_993# VSS 3.19e-21
C5560 a_2773_627# VSS 0.0997f
C5561 a_3648_993# VSS 0.245f
C5562 a_3807_895# VSS 0.466f
C5563 a_3333_601# VSS 0.396f
C5564 a_2865_993# VSS 0.258f
C5565 a_3039_601# VSS 0.278f
C5566 a_2585_627# VSS 0.314f
C5567 D[6] VSS 1.91f
C5568 a_2419_627# VSS 0.713f
C5569 VDD_SW[7] VSS 0.505f
C5570 a_1363_627# VSS 0.00292f
C5571 a_1555_627# VSS 0.177f
C5572 a_2136_627# VSS 0.244f
C5573 VDD_SW_b[7] VSS 0.526f
C5574 a_1672_909# VSS 0.00333f
C5575 a_1159_627# VSS 0.0166f
C5576 a_581_627# VSS 0.00202f
C5577 a_791_627# VSS 0.177f
C5578 a_1340_993# VSS 8.02e-19
C5579 a_1112_909# VSS 0.00617f
C5580 a_891_909# VSS 6.69e-21
C5581 a_557_993# VSS 1.71e-19
C5582 a_381_627# VSS 0.101f
C5583 a_1256_993# VSS 0.28f
C5584 a_1415_895# VSS 0.496f
C5585 a_941_601# VSS 0.422f
C5586 a_473_993# VSS 0.261f
C5587 a_647_601# VSS 0.283f
C5588 a_193_627# VSS 0.337f
C5589 D[7] VSS 1.99f
C5590 a_27_627# VSS 0.778f
C5591 a_16330_1315# VSS 0.00466f
C5592 a_16109_1315# VSS 0.00881f
C5593 a_14791_1315# VSS 0.00733f
C5594 a_14570_1315# VSS 0.00339f
C5595 x20.X VSS 0.952f
C5596 a_13936_1315# VSS 0.00405f
C5597 a_13715_1315# VSS 0.00855f
C5598 a_12399_1315# VSS 0.00726f
C5599 a_12178_1315# VSS 0.00335f
C5600 a_16323_1642# VSS 0.00103f
C5601 a_16037_1642# VSS 0.00133f
C5602 a_14887_1642# VSS 2.7e-19
C5603 a_14570_1642# VSS 7.29e-19
C5604 a_15855_1642# VSS 0.369f
C5605 a_14857_1289# VSS 0.34f
C5606 check[0] VSS 1.09f
C5607 x18.X VSS 0.326f
C5608 x17.X VSS 0.682f
C5609 a_11546_1315# VSS 0.00336f
C5610 a_11325_1315# VSS 0.0077f
C5611 a_10007_1315# VSS 0.00863f
C5612 a_9786_1315# VSS 0.0035f
C5613 a_13929_1642# VSS 0.00102f
C5614 a_13643_1642# VSS 7.44e-19
C5615 a_12495_1642# VSS 2.7e-19
C5616 a_12178_1642# VSS 7.29e-19
C5617 a_13461_1642# VSS 0.366f
C5618 a_12465_1289# VSS 0.345f
C5619 check[1] VSS 1.13f
C5620 x16.X VSS 0.325f
C5621 x15.X VSS 0.519f
C5622 a_9154_1315# VSS 0.00335f
C5623 a_8933_1315# VSS 0.00727f
C5624 a_7615_1315# VSS 0.00869f
C5625 a_7394_1315# VSS 0.00455f
C5626 a_11539_1642# VSS 4e-19
C5627 a_11253_1642# VSS 7.89e-19
C5628 a_10103_1642# VSS 0.00113f
C5629 a_9786_1642# VSS 8.8e-19
C5630 a_11071_1642# VSS 0.367f
C5631 a_10073_1289# VSS 0.372f
C5632 check[2] VSS 1.13f
C5633 x14.X VSS 0.325f
C5634 x13.X VSS 0.519f
C5635 a_6760_1315# VSS 0.00335f
C5636 a_6539_1315# VSS 0.00726f
C5637 a_5223_1315# VSS 0.00867f
C5638 a_5002_1315# VSS 0.00473f
C5639 a_9147_1642# VSS 4e-19
C5640 a_8861_1642# VSS 2.7e-19
C5641 a_7711_1642# VSS 0.0012f
C5642 a_7394_1642# VSS 0.00235f
C5643 a_8679_1642# VSS 0.343f
C5644 a_7681_1289# VSS 0.366f
C5645 check[3] VSS 1.01f
C5646 x12.X VSS 0.392f
C5647 x11.X VSS 0.626f
C5648 a_4370_1315# VSS 0.00407f
C5649 a_4149_1315# VSS 0.00876f
C5650 a_2831_1315# VSS 0.00726f
C5651 a_2610_1315# VSS 0.0034f
C5652 a_6753_1642# VSS 3.84e-19
C5653 a_6467_1642# VSS 2.7e-19
C5654 a_5319_1642# VSS 0.00166f
C5655 a_5002_1642# VSS 0.00261f
C5656 a_6285_1642# VSS 0.338f
C5657 a_5289_1289# VSS 0.346f
C5658 check[4] VSS 0.864f
C5659 x10.X VSS 0.39f
C5660 x9.X VSS 0.736f
C5661 a_1978_1315# VSS 0.00431f
C5662 a_1757_1315# VSS 0.00815f
C5663 a_439_1315# VSS 0.00729f
C5664 a_218_1315# VSS 0.00335f
C5665 a_4363_1642# VSS 0.00108f
C5666 a_4077_1642# VSS 8.72e-19
C5667 a_2927_1642# VSS 2.7e-19
C5668 a_2610_1642# VSS 7.29e-19
C5669 a_3895_1642# VSS 0.344f
C5670 a_2897_1289# VSS 0.339f
C5671 check[5] VSS 0.99f
C5672 x8.X VSS 0.376f
C5673 x7.X VSS 0.688f
C5674 a_1971_1642# VSS 0.00118f
C5675 a_1685_1642# VSS 0.00141f
C5676 a_535_1642# VSS 2.7e-19
C5677 a_218_1642# VSS 7.29e-19
C5678 a_1503_1642# VSS 0.368f
C5679 a_505_1289# VSS 0.341f
C5680 check[6] VSS 1.06f
C5681 x6.X VSS 0.582f
C5682 a_16109_1642# VSS 0.373f
C5683 a_14428_1467# VSS 0.331f
C5684 a_13715_1642# VSS 0.356f
C5685 a_12036_1467# VSS 0.331f
C5686 a_11325_1642# VSS 0.327f
C5687 a_9644_1467# VSS 0.339f
C5688 a_8933_1642# VSS 0.327f
C5689 a_7252_1467# VSS 0.365f
C5690 a_6539_1642# VSS 0.329f
C5691 a_4860_1467# VSS 0.365f
C5692 a_4149_1642# VSS 0.355f
C5693 a_2468_1467# VSS 0.334f
C5694 a_1757_1642# VSS 0.356f
C5695 a_76_1467# VSS 0.343f
C5696 x9.A1 VSS 11.9f
C5697 x2.X VSS 18.3f
C5698 a_5323_2457# VSS 2.14f
C5699 x30.A VSS 0.991f
C5700 a_4689_2457# VSS 0.558f
C5701 x27.A VSS 0.212f
C5702 a_4413_2457# VSS 0.296f
C5703 ready VSS 2.39f
C5704 a_939_2457# VSS 2.1f
C5705 x3.X VSS 0.93f
C5706 a_305_2457# VSS 0.509f
C5707 x3.A VSS 0.196f
C5708 a_29_2457# VSS 0.274f
C5709 reset VSS 0.22f
C5710 VDD VSS 0.132p
C5711 x9.A1.n0 VSS 0.021f
C5712 x9.A1.n1 VSS 0.021f
C5713 x9.A1.n2 VSS 0.021f
C5714 x9.A1.n3 VSS 0.021f
C5715 x9.A1.n4 VSS 0.021f
C5716 x9.A1.n5 VSS 0.021f
C5717 x9.A1.n6 VSS 0.021f
C5718 x9.A1.t8 VSS 0.0273f
C5719 x9.A1.t2 VSS 0.0273f
C5720 x9.A1.n7 VSS 0.0674f
C5721 x9.A1.t12 VSS 0.0273f
C5722 x9.A1.t4 VSS 0.0273f
C5723 x9.A1.n8 VSS 0.104f
C5724 x9.A1.t11 VSS 0.0273f
C5725 x9.A1.t6 VSS 0.0273f
C5726 x9.A1.n9 VSS 0.0674f
C5727 x9.A1.n10 VSS 0.262f
C5728 x9.A1.t14 VSS 0.0273f
C5729 x9.A1.t0 VSS 0.0273f
C5730 x9.A1.n11 VSS 0.0674f
C5731 x9.A1.n12 VSS 0.158f
C5732 x9.A1.t9 VSS 0.0273f
C5733 x9.A1.t1 VSS 0.0273f
C5734 x9.A1.n13 VSS 0.0674f
C5735 x9.A1.n14 VSS 0.158f
C5736 x9.A1.t10 VSS 0.0273f
C5737 x9.A1.t3 VSS 0.0273f
C5738 x9.A1.n15 VSS 0.0674f
C5739 x9.A1.n16 VSS 0.158f
C5740 x9.A1.t13 VSS 0.0273f
C5741 x9.A1.t5 VSS 0.0273f
C5742 x9.A1.n17 VSS 0.0674f
C5743 x9.A1.n18 VSS 0.158f
C5744 x9.A1.t15 VSS 0.0273f
C5745 x9.A1.t7 VSS 0.0273f
C5746 x9.A1.n19 VSS 0.0674f
C5747 x9.A1.n20 VSS 0.158f
C5748 x9.A1.n21 VSS 0.151f
C5749 x9.A1.n22 VSS 0.0159f
C5750 x9.A1.t42 VSS 0.0747f
C5751 x9.A1.n23 VSS 0.123f
C5752 x9.A1.t55 VSS 0.0213f
C5753 x9.A1.n24 VSS 0.0625f
C5754 x9.A1.n25 VSS 0.00787f
C5755 x9.A1.n26 VSS 0.00438f
C5756 x9.A1.n27 VSS 0.00456f
C5757 x9.A1.n28 VSS 0.0141f
C5758 x9.A1.n29 VSS 0.0238f
C5759 x9.A1.n30 VSS 0.181f
C5760 x9.A1.n31 VSS 0.0136f
C5761 x9.A1.t32 VSS 0.0214f
C5762 x9.A1.n32 VSS 0.0615f
C5763 x9.A1.n33 VSS 0.00798f
C5764 x9.A1.t43 VSS 0.0749f
C5765 x9.A1.n34 VSS 0.124f
C5766 x9.A1.n35 VSS 0.00455f
C5767 x9.A1.n36 VSS 0.0238f
C5768 x9.A1.n37 VSS 0.159f
C5769 x9.A1.n38 VSS 0.487f
C5770 x9.A1.n39 VSS 0.0159f
C5771 x9.A1.t53 VSS 0.0748f
C5772 x9.A1.n40 VSS 0.123f
C5773 x9.A1.t40 VSS 0.0213f
C5774 x9.A1.n41 VSS 0.0614f
C5775 x9.A1.n42 VSS 0.00863f
C5776 x9.A1.n43 VSS 0.00438f
C5777 x9.A1.n44 VSS 0.00456f
C5778 x9.A1.n45 VSS 0.0141f
C5779 x9.A1.n46 VSS 0.0238f
C5780 x9.A1.n47 VSS 0.159f
C5781 x9.A1.n48 VSS 0.468f
C5782 x9.A1.n49 VSS 0.0136f
C5783 x9.A1.t44 VSS 0.0215f
C5784 x9.A1.n50 VSS 0.0613f
C5785 x9.A1.n51 VSS 0.00818f
C5786 x9.A1.t56 VSS 0.0749f
C5787 x9.A1.n52 VSS 0.124f
C5788 x9.A1.n53 VSS 0.00464f
C5789 x9.A1.n54 VSS 0.0238f
C5790 x9.A1.n55 VSS 0.159f
C5791 x9.A1.n56 VSS 0.468f
C5792 x9.A1.n57 VSS 0.0159f
C5793 x9.A1.t48 VSS 0.0747f
C5794 x9.A1.n58 VSS 0.123f
C5795 x9.A1.t35 VSS 0.0213f
C5796 x9.A1.n59 VSS 0.0625f
C5797 x9.A1.n60 VSS 0.00787f
C5798 x9.A1.n61 VSS 0.00438f
C5799 x9.A1.n62 VSS 0.00456f
C5800 x9.A1.n63 VSS 0.0141f
C5801 x9.A1.n64 VSS 0.0238f
C5802 x9.A1.n65 VSS 0.159f
C5803 x9.A1.n66 VSS 0.468f
C5804 x9.A1.n67 VSS 0.0136f
C5805 x9.A1.t57 VSS 0.0214f
C5806 x9.A1.n68 VSS 0.0615f
C5807 x9.A1.n69 VSS 0.00798f
C5808 x9.A1.t58 VSS 0.0749f
C5809 x9.A1.n70 VSS 0.124f
C5810 x9.A1.n71 VSS 0.00455f
C5811 x9.A1.n72 VSS 0.0238f
C5812 x9.A1.n73 VSS 0.159f
C5813 x9.A1.n74 VSS 0.469f
C5814 x9.A1.n75 VSS 0.0159f
C5815 x9.A1.t34 VSS 0.0748f
C5816 x9.A1.n76 VSS 0.123f
C5817 x9.A1.t33 VSS 0.0213f
C5818 x9.A1.n77 VSS 0.0614f
C5819 x9.A1.n78 VSS 0.00863f
C5820 x9.A1.n79 VSS 0.00438f
C5821 x9.A1.n80 VSS 0.00456f
C5822 x9.A1.n81 VSS 0.0141f
C5823 x9.A1.n82 VSS 0.0238f
C5824 x9.A1.n83 VSS 0.159f
C5825 x9.A1.n84 VSS 0.468f
C5826 x9.A1.n85 VSS 0.0136f
C5827 x9.A1.t59 VSS 0.0214f
C5828 x9.A1.n86 VSS 0.0595f
C5829 x9.A1.n87 VSS 0.00963f
C5830 x9.A1.t41 VSS 0.075f
C5831 x9.A1.n88 VSS 0.124f
C5832 x9.A1.n89 VSS 0.00447f
C5833 x9.A1.n90 VSS 0.0238f
C5834 x9.A1.n91 VSS 0.159f
C5835 x9.A1.n92 VSS 0.312f
C5836 x9.A1.n93 VSS 0.0159f
C5837 x9.A1.t51 VSS 0.0747f
C5838 x9.A1.n94 VSS 0.123f
C5839 x9.A1.t54 VSS 0.0213f
C5840 x9.A1.n95 VSS 0.0625f
C5841 x9.A1.n96 VSS 0.00787f
C5842 x9.A1.n97 VSS 0.00438f
C5843 x9.A1.n98 VSS 0.00456f
C5844 x9.A1.n99 VSS 0.0141f
C5845 x9.A1.n100 VSS 0.0238f
C5846 x9.A1.n101 VSS 0.157f
C5847 x9.A1.n102 VSS 0.0136f
C5848 x9.A1.t36 VSS 0.0214f
C5849 x9.A1.n103 VSS 0.0598f
C5850 x9.A1.n104 VSS 0.00934f
C5851 x9.A1.t45 VSS 0.075f
C5852 x9.A1.n105 VSS 0.124f
C5853 x9.A1.n106 VSS 0.00455f
C5854 x9.A1.n107 VSS 0.0238f
C5855 x9.A1.n108 VSS 0.159f
C5856 x9.A1.n109 VSS 0.0159f
C5857 x9.A1.t46 VSS 0.0748f
C5858 x9.A1.n110 VSS 0.123f
C5859 x9.A1.t49 VSS 0.0214f
C5860 x9.A1.n111 VSS 0.0612f
C5861 x9.A1.n112 VSS 0.00885f
C5862 x9.A1.n113 VSS 0.00447f
C5863 x9.A1.n114 VSS 0.00456f
C5864 x9.A1.n115 VSS 0.0141f
C5865 x9.A1.n116 VSS 0.0238f
C5866 x9.A1.n117 VSS 0.159f
C5867 x9.A1.n118 VSS 0.0136f
C5868 x9.A1.t37 VSS 0.0214f
C5869 x9.A1.n119 VSS 0.0598f
C5870 x9.A1.n120 VSS 0.00934f
C5871 x9.A1.t47 VSS 0.075f
C5872 x9.A1.n121 VSS 0.124f
C5873 x9.A1.n122 VSS 0.00455f
C5874 x9.A1.n123 VSS 0.0238f
C5875 x9.A1.n124 VSS 0.159f
C5876 x9.A1.n125 VSS 0.0159f
C5877 x9.A1.t39 VSS 0.0748f
C5878 x9.A1.n126 VSS 0.123f
C5879 x9.A1.t50 VSS 0.0214f
C5880 x9.A1.n127 VSS 0.0612f
C5881 x9.A1.n128 VSS 0.00885f
C5882 x9.A1.n129 VSS 0.00447f
C5883 x9.A1.n130 VSS 0.00456f
C5884 x9.A1.n131 VSS 0.0141f
C5885 x9.A1.n132 VSS 0.0238f
C5886 x9.A1.n133 VSS 0.159f
C5887 x9.A1.n134 VSS 0.0136f
C5888 x9.A1.t52 VSS 0.0214f
C5889 x9.A1.n135 VSS 0.0612f
C5890 x9.A1.n136 VSS 0.00834f
C5891 x9.A1.t38 VSS 0.0749f
C5892 x9.A1.n137 VSS 0.123f
C5893 x9.A1.n138 VSS 0.00447f
C5894 x9.A1.n139 VSS 0.0238f
C5895 x9.A1.n140 VSS 0.245f
C5896 x9.A1.n141 VSS 0.54f
C5897 x9.A1.n142 VSS 0.468f
C5898 x9.A1.n143 VSS 0.468f
C5899 x9.A1.n144 VSS 0.468f
C5900 x9.A1.n145 VSS 0.429f
C5901 x9.A1.n146 VSS 0.529f
C5902 x9.A1.n147 VSS 0.199f
C5903 x9.A1.t20 VSS 0.0177f
C5904 x9.A1.t28 VSS 0.0177f
C5905 x9.A1.n148 VSS 0.0842f
C5906 x9.A1.t19 VSS 0.0177f
C5907 x9.A1.t30 VSS 0.0177f
C5908 x9.A1.n149 VSS 0.0444f
C5909 x9.A1.n150 VSS 0.166f
C5910 x9.A1.t22 VSS 0.0177f
C5911 x9.A1.t24 VSS 0.0177f
C5912 x9.A1.n151 VSS 0.0444f
C5913 x9.A1.n152 VSS 0.112f
C5914 x9.A1.t17 VSS 0.0177f
C5915 x9.A1.t25 VSS 0.0177f
C5916 x9.A1.n153 VSS 0.0445f
C5917 x9.A1.n154 VSS 0.112f
C5918 x9.A1.t18 VSS 0.0177f
C5919 x9.A1.t27 VSS 0.0177f
C5920 x9.A1.n155 VSS 0.0445f
C5921 x9.A1.n156 VSS 0.112f
C5922 x9.A1.t21 VSS 0.0177f
C5923 x9.A1.t29 VSS 0.0177f
C5924 x9.A1.n157 VSS 0.0445f
C5925 x9.A1.n158 VSS 0.112f
C5926 x9.A1.t23 VSS 0.0177f
C5927 x9.A1.t31 VSS 0.0177f
C5928 x9.A1.n159 VSS 0.0445f
C5929 x9.A1.n160 VSS 0.112f
C5930 x9.A1.t16 VSS 0.0177f
C5931 x9.A1.t26 VSS 0.0177f
C5932 x9.A1.n161 VSS 0.0445f
C5933 x9.A1.n162 VSS 0.111f
C5934 x2.X.n0 VSS 0.0087f
C5935 x2.X.n1 VSS 0.0087f
C5936 x2.X.n2 VSS 0.0087f
C5937 x2.X.n3 VSS 0.0087f
C5938 x2.X.n4 VSS 0.0087f
C5939 x2.X.n5 VSS 0.0087f
C5940 x2.X.n6 VSS 0.0087f
C5941 x2.X.n7 VSS 0.00408f
C5942 x2.X.t69 VSS 0.0299f
C5943 x2.X.n8 VSS 0.0415f
C5944 x2.X.t55 VSS 0.0131f
C5945 x2.X.n9 VSS 0.0173f
C5946 x2.X.n10 VSS 0.0173f
C5947 x2.X.n11 VSS 0.0135f
C5948 x2.X.n12 VSS 0.0826f
C5949 x2.X.t52 VSS 0.031f
C5950 x2.X.t51 VSS 0.0131f
C5951 x2.X.n13 VSS 0.0592f
C5952 x2.X.n14 VSS 0.0171f
C5953 x2.X.n15 VSS 0.00673f
C5954 x2.X.n16 VSS 0.00355f
C5955 x2.X.n17 VSS 0.00485f
C5956 x2.X.n18 VSS 0.0322f
C5957 x2.X.n19 VSS 0.091f
C5958 x2.X.n20 VSS 0.0126f
C5959 x2.X.n21 VSS 0.00384f
C5960 x2.X.n22 VSS 0.00284f
C5961 x2.X.t65 VSS 0.0207f
C5962 x2.X.t50 VSS 0.0175f
C5963 x2.X.n23 VSS 0.0279f
C5964 x2.X.n24 VSS 0.0308f
C5965 x2.X.n25 VSS 0.119f
C5966 x2.X.n26 VSS 0.61f
C5967 x2.X.n27 VSS 0.00408f
C5968 x2.X.t72 VSS 0.0299f
C5969 x2.X.n28 VSS 0.0415f
C5970 x2.X.t57 VSS 0.0131f
C5971 x2.X.n29 VSS 0.0173f
C5972 x2.X.n30 VSS 0.0173f
C5973 x2.X.n31 VSS 0.0135f
C5974 x2.X.n32 VSS 0.0826f
C5975 x2.X.t66 VSS 0.031f
C5976 x2.X.t63 VSS 0.0131f
C5977 x2.X.n33 VSS 0.0592f
C5978 x2.X.n34 VSS 0.0171f
C5979 x2.X.n35 VSS 0.00673f
C5980 x2.X.n36 VSS 0.00355f
C5981 x2.X.n37 VSS 0.00485f
C5982 x2.X.n38 VSS 0.0322f
C5983 x2.X.n39 VSS 0.091f
C5984 x2.X.n40 VSS 0.0126f
C5985 x2.X.n41 VSS 0.00384f
C5986 x2.X.n42 VSS 0.00284f
C5987 x2.X.t70 VSS 0.0207f
C5988 x2.X.t54 VSS 0.0175f
C5989 x2.X.n43 VSS 0.0279f
C5990 x2.X.n44 VSS 0.0308f
C5991 x2.X.n45 VSS 0.119f
C5992 x2.X.n46 VSS 0.47f
C5993 x2.X.n47 VSS 0.925f
C5994 x2.X.n48 VSS 0.00408f
C5995 x2.X.t39 VSS 0.0299f
C5996 x2.X.n49 VSS 0.0415f
C5997 x2.X.t59 VSS 0.0131f
C5998 x2.X.n50 VSS 0.0173f
C5999 x2.X.n51 VSS 0.0173f
C6000 x2.X.n52 VSS 0.0135f
C6001 x2.X.n53 VSS 0.0828f
C6002 x2.X.t68 VSS 0.031f
C6003 x2.X.t67 VSS 0.0131f
C6004 x2.X.n54 VSS 0.0592f
C6005 x2.X.n55 VSS 0.0171f
C6006 x2.X.n56 VSS 0.00673f
C6007 x2.X.n57 VSS 0.00355f
C6008 x2.X.n58 VSS 0.00485f
C6009 x2.X.n59 VSS 0.0322f
C6010 x2.X.n60 VSS 0.0931f
C6011 x2.X.n61 VSS 0.0129f
C6012 x2.X.n62 VSS 0.00384f
C6013 x2.X.n63 VSS 0.00284f
C6014 x2.X.t73 VSS 0.0207f
C6015 x2.X.t56 VSS 0.0175f
C6016 x2.X.n64 VSS 0.0279f
C6017 x2.X.n65 VSS 0.0308f
C6018 x2.X.n66 VSS 0.119f
C6019 x2.X.n67 VSS 0.47f
C6020 x2.X.n68 VSS 0.852f
C6021 x2.X.n69 VSS 0.00408f
C6022 x2.X.t58 VSS 0.0299f
C6023 x2.X.n70 VSS 0.0415f
C6024 x2.X.t38 VSS 0.0131f
C6025 x2.X.n71 VSS 0.0173f
C6026 x2.X.n72 VSS 0.0173f
C6027 x2.X.n73 VSS 0.0135f
C6028 x2.X.n74 VSS 0.0826f
C6029 x2.X.t37 VSS 0.031f
C6030 x2.X.t36 VSS 0.0131f
C6031 x2.X.n75 VSS 0.0592f
C6032 x2.X.n76 VSS 0.0171f
C6033 x2.X.n77 VSS 0.00673f
C6034 x2.X.n78 VSS 0.00355f
C6035 x2.X.n79 VSS 0.00485f
C6036 x2.X.n80 VSS 0.0324f
C6037 x2.X.n81 VSS 0.0913f
C6038 x2.X.n82 VSS 0.0126f
C6039 x2.X.n83 VSS 0.00384f
C6040 x2.X.n84 VSS 0.00284f
C6041 x2.X.t41 VSS 0.0207f
C6042 x2.X.t71 VSS 0.0175f
C6043 x2.X.n85 VSS 0.0279f
C6044 x2.X.n86 VSS 0.0308f
C6045 x2.X.n87 VSS 0.119f
C6046 x2.X.n88 VSS 0.47f
C6047 x2.X.n89 VSS 0.853f
C6048 x2.X.n90 VSS 0.00408f
C6049 x2.X.t60 VSS 0.0299f
C6050 x2.X.n91 VSS 0.0415f
C6051 x2.X.t46 VSS 0.0131f
C6052 x2.X.n92 VSS 0.0173f
C6053 x2.X.n93 VSS 0.0173f
C6054 x2.X.n94 VSS 0.0135f
C6055 x2.X.n95 VSS 0.0826f
C6056 x2.X.t42 VSS 0.031f
C6057 x2.X.t40 VSS 0.0131f
C6058 x2.X.n96 VSS 0.0592f
C6059 x2.X.n97 VSS 0.0171f
C6060 x2.X.n98 VSS 0.00673f
C6061 x2.X.n99 VSS 0.00355f
C6062 x2.X.n100 VSS 0.00485f
C6063 x2.X.n101 VSS 0.0324f
C6064 x2.X.n102 VSS 0.0913f
C6065 x2.X.n103 VSS 0.0126f
C6066 x2.X.n104 VSS 0.00384f
C6067 x2.X.n105 VSS 0.00284f
C6068 x2.X.t48 VSS 0.0207f
C6069 x2.X.t32 VSS 0.0175f
C6070 x2.X.n106 VSS 0.0279f
C6071 x2.X.n107 VSS 0.0308f
C6072 x2.X.n108 VSS 0.119f
C6073 x2.X.n109 VSS 0.47f
C6074 x2.X.n110 VSS 0.852f
C6075 x2.X.n111 VSS 0.00408f
C6076 x2.X.t33 VSS 0.0299f
C6077 x2.X.n112 VSS 0.0415f
C6078 x2.X.t61 VSS 0.0131f
C6079 x2.X.n113 VSS 0.0173f
C6080 x2.X.n114 VSS 0.0173f
C6081 x2.X.n115 VSS 0.0135f
C6082 x2.X.n116 VSS 0.0826f
C6083 x2.X.t49 VSS 0.031f
C6084 x2.X.t45 VSS 0.0131f
C6085 x2.X.n117 VSS 0.0592f
C6086 x2.X.n118 VSS 0.0171f
C6087 x2.X.n119 VSS 0.00673f
C6088 x2.X.n120 VSS 0.00355f
C6089 x2.X.n121 VSS 0.00485f
C6090 x2.X.n122 VSS 0.0324f
C6091 x2.X.n123 VSS 0.0913f
C6092 x2.X.n124 VSS 0.0126f
C6093 x2.X.n125 VSS 0.00384f
C6094 x2.X.n126 VSS 0.00284f
C6095 x2.X.t62 VSS 0.0207f
C6096 x2.X.t44 VSS 0.0175f
C6097 x2.X.n127 VSS 0.0279f
C6098 x2.X.n128 VSS 0.0308f
C6099 x2.X.n129 VSS 0.121f
C6100 x2.X.n130 VSS 0.468f
C6101 x2.X.n131 VSS 0.625f
C6102 x2.X.n132 VSS 0.00408f
C6103 x2.X.t35 VSS 0.0299f
C6104 x2.X.n133 VSS 0.0415f
C6105 x2.X.t64 VSS 0.0131f
C6106 x2.X.n134 VSS 0.0173f
C6107 x2.X.n135 VSS 0.0173f
C6108 x2.X.n136 VSS 0.0135f
C6109 x2.X.n137 VSS 0.0826f
C6110 x2.X.t47 VSS 0.031f
C6111 x2.X.t43 VSS 0.0131f
C6112 x2.X.n138 VSS 0.0592f
C6113 x2.X.n139 VSS 0.0171f
C6114 x2.X.n140 VSS 0.00673f
C6115 x2.X.n141 VSS 0.00355f
C6116 x2.X.n142 VSS 0.00485f
C6117 x2.X.n143 VSS 0.0322f
C6118 x2.X.n144 VSS 0.091f
C6119 x2.X.n145 VSS 0.0126f
C6120 x2.X.n146 VSS 0.00384f
C6121 x2.X.n147 VSS 0.00284f
C6122 x2.X.t53 VSS 0.0208f
C6123 x2.X.t34 VSS 0.0175f
C6124 x2.X.n148 VSS 0.0272f
C6125 x2.X.n149 VSS 0.0314f
C6126 x2.X.n150 VSS 0.118f
C6127 x2.X.n151 VSS 0.631f
C6128 x2.X.n152 VSS 0.595f
C6129 x2.X.t3 VSS 0.0196f
C6130 x2.X.t14 VSS 0.0196f
C6131 x2.X.n153 VSS 0.0485f
C6132 x2.X.t8 VSS 0.0196f
C6133 x2.X.t13 VSS 0.0196f
C6134 x2.X.n154 VSS 0.0485f
C6135 x2.X.t6 VSS 0.0196f
C6136 x2.X.t11 VSS 0.0196f
C6137 x2.X.n155 VSS 0.0485f
C6138 x2.X.t4 VSS 0.0196f
C6139 x2.X.t10 VSS 0.0196f
C6140 x2.X.n156 VSS 0.0485f
C6141 x2.X.t2 VSS 0.0196f
C6142 x2.X.t1 VSS 0.0196f
C6143 x2.X.n157 VSS 0.0485f
C6144 x2.X.t9 VSS 0.0196f
C6145 x2.X.t0 VSS 0.0196f
C6146 x2.X.n158 VSS 0.0485f
C6147 x2.X.t7 VSS 0.0196f
C6148 x2.X.t12 VSS 0.0196f
C6149 x2.X.n159 VSS 0.0485f
C6150 x2.X.t5 VSS 0.0196f
C6151 x2.X.t15 VSS 0.0196f
C6152 x2.X.n160 VSS 0.0749f
C6153 x2.X.n161 VSS 0.189f
C6154 x2.X.n162 VSS 0.114f
C6155 x2.X.n163 VSS 0.114f
C6156 x2.X.n164 VSS 0.114f
C6157 x2.X.n165 VSS 0.114f
C6158 x2.X.n166 VSS 0.114f
C6159 x2.X.n167 VSS 0.108f
C6160 x2.X.n168 VSS 0.0499f
C6161 x2.X.t27 VSS 0.0128f
C6162 x2.X.t21 VSS 0.0128f
C6163 x2.X.n169 VSS 0.0605f
C6164 x2.X.t29 VSS 0.0128f
C6165 x2.X.t18 VSS 0.0128f
C6166 x2.X.n170 VSS 0.0319f
C6167 x2.X.n171 VSS 0.12f
C6168 x2.X.t31 VSS 0.0128f
C6169 x2.X.t22 VSS 0.0128f
C6170 x2.X.n172 VSS 0.0319f
C6171 x2.X.n173 VSS 0.0804f
C6172 x2.X.t24 VSS 0.0128f
C6173 x2.X.t23 VSS 0.0128f
C6174 x2.X.n174 VSS 0.0319f
C6175 x2.X.n175 VSS 0.0806f
C6176 x2.X.t26 VSS 0.0128f
C6177 x2.X.t16 VSS 0.0128f
C6178 x2.X.n176 VSS 0.0319f
C6179 x2.X.n177 VSS 0.0806f
C6180 x2.X.t28 VSS 0.0128f
C6181 x2.X.t17 VSS 0.0128f
C6182 x2.X.n178 VSS 0.0319f
C6183 x2.X.n179 VSS 0.0806f
C6184 x2.X.t30 VSS 0.0128f
C6185 x2.X.t19 VSS 0.0128f
C6186 x2.X.n180 VSS 0.0319f
C6187 x2.X.n181 VSS 0.0806f
C6188 x2.X.t25 VSS 0.0128f
C6189 x2.X.t20 VSS 0.0128f
C6190 x2.X.n182 VSS 0.0319f
C6191 x2.X.n183 VSS 0.0795f
C6192 VDD.n0 VSS 0.0517f
C6193 VDD.n1 VSS 0.00158f
C6194 VDD.t532 VSS 0.00349f
C6195 VDD.n2 VSS 0.00297f
C6196 VDD.t531 VSS 0.00616f
C6197 VDD.n3 VSS 0.00867f
C6198 VDD.n4 VSS 0.00109f
C6199 VDD.n5 VSS 0.00103f
C6200 VDD.n6 VSS 0.00302f
C6201 VDD.n7 VSS 0.0176f
C6202 VDD.n8 VSS 0.276f
C6203 VDD.n9 VSS 0.0114f
C6204 VDD.n10 VSS 0.00148f
C6205 VDD.n11 VSS 8.1e-19
C6206 VDD.n12 VSS 0.0114f
C6207 VDD.n13 VSS 0.0307f
C6208 VDD.n14 VSS 4.84e-19
C6209 VDD.n15 VSS 4.84e-19
C6210 VDD.n16 VSS 0.00653f
C6211 VDD.n17 VSS 0.00158f
C6212 VDD.n18 VSS 6.05e-19
C6213 VDD.n19 VSS 5.07e-19
C6214 VDD.t527 VSS 0.00578f
C6215 VDD.n20 VSS 0.00528f
C6216 VDD.n21 VSS 0.00109f
C6217 VDD.n22 VSS 0.00147f
C6218 VDD.n23 VSS 0.00243f
C6219 VDD.n24 VSS 0.00112f
C6220 VDD.n25 VSS 0.00154f
C6221 VDD.n26 VSS 9.31e-19
C6222 VDD.t539 VSS 0.00578f
C6223 VDD.n27 VSS 0.00528f
C6224 VDD.n28 VSS 0.00109f
C6225 VDD.n29 VSS 1.72e-19
C6226 VDD.n30 VSS 2.85e-19
C6227 VDD.t528 VSS 9.42e-19
C6228 VDD.t540 VSS 9.42e-19
C6229 VDD.n31 VSS 0.00214f
C6230 VDD.n32 VSS 0.0025f
C6231 VDD.n33 VSS 3.44e-19
C6232 VDD.n34 VSS 4.19e-19
C6233 VDD.n35 VSS 4.35e-19
C6234 VDD.n36 VSS 3.36e-19
C6235 VDD.n37 VSS 8.11e-19
C6236 VDD.n38 VSS 0.00148f
C6237 VDD.n39 VSS 0.00653f
C6238 VDD.n40 VSS 4.95e-19
C6239 VDD.t524 VSS 9.42e-19
C6240 VDD.t663 VSS 9.42e-19
C6241 VDD.n41 VSS 0.00214f
C6242 VDD.n42 VSS 0.00258f
C6243 VDD.t523 VSS 0.0106f
C6244 VDD.n43 VSS 0.00109f
C6245 VDD.n44 VSS 0.00126f
C6246 VDD.n45 VSS 0.00251f
C6247 VDD.n46 VSS 0.00142f
C6248 VDD.t657 VSS 9.42e-19
C6249 VDD.t661 VSS 9.42e-19
C6250 VDD.n47 VSS 0.00214f
C6251 VDD.n48 VSS 0.00244f
C6252 VDD.t656 VSS 0.00578f
C6253 VDD.n49 VSS 0.00528f
C6254 VDD.n50 VSS 0.00109f
C6255 VDD.n51 VSS 0.00119f
C6256 VDD.n52 VSS 0.00256f
C6257 VDD.n53 VSS 0.00154f
C6258 VDD.t662 VSS 0.00578f
C6259 VDD.n54 VSS 0.00528f
C6260 VDD.n55 VSS 0.00109f
C6261 VDD.n56 VSS 0.00144f
C6262 VDD.n57 VSS 4.19e-19
C6263 VDD.n58 VSS 4.19e-19
C6264 VDD.n59 VSS 3.1e-19
C6265 VDD.n60 VSS 3.23e-19
C6266 VDD.n61 VSS 3.23e-19
C6267 VDD.n62 VSS 0.00149f
C6268 VDD.n63 VSS 8.1e-19
C6269 VDD.n64 VSS 0.00157f
C6270 VDD.n65 VSS 6.73e-19
C6271 VDD.t518 VSS 9.42e-19
C6272 VDD.t544 VSS 9.42e-19
C6273 VDD.n66 VSS 0.00214f
C6274 VDD.n67 VSS 0.00258f
C6275 VDD.t517 VSS 0.00578f
C6276 VDD.t543 VSS 0.00578f
C6277 VDD.n68 VSS 0.00528f
C6278 VDD.n69 VSS 0.00109f
C6279 VDD.n70 VSS 9.51e-19
C6280 VDD.n71 VSS 0.00308f
C6281 VDD.t515 VSS 0.00578f
C6282 VDD.n72 VSS 0.00528f
C6283 VDD.n73 VSS 0.00109f
C6284 VDD.n74 VSS 0.00168f
C6285 VDD.n75 VSS 0.00245f
C6286 VDD.n76 VSS 9.71e-19
C6287 VDD.n77 VSS 0.00154f
C6288 VDD.n78 VSS 9.31e-19
C6289 VDD.t537 VSS 0.00578f
C6290 VDD.n79 VSS 0.00528f
C6291 VDD.n80 VSS 0.00109f
C6292 VDD.n81 VSS 1.72e-19
C6293 VDD.n82 VSS 2.85e-19
C6294 VDD.t516 VSS 9.42e-19
C6295 VDD.t538 VSS 9.42e-19
C6296 VDD.n83 VSS 0.00214f
C6297 VDD.n84 VSS 0.00246f
C6298 VDD.n85 VSS 1.82e-19
C6299 VDD.n86 VSS 5.7e-19
C6300 VDD.n87 VSS 4.35e-19
C6301 VDD.n88 VSS 4.39e-19
C6302 VDD.n89 VSS 3.36e-19
C6303 VDD.n90 VSS 0.00149f
C6304 VDD.n91 VSS 8.1e-19
C6305 VDD.n92 VSS 0.00157f
C6306 VDD.n93 VSS 4.86e-19
C6307 VDD.n94 VSS 0.00149f
C6308 VDD.n95 VSS 6.98e-19
C6309 VDD.n96 VSS 4.13e-19
C6310 VDD.t529 VSS 0.00553f
C6311 VDD.n97 VSS 0.00528f
C6312 VDD.n98 VSS 0.00109f
C6313 VDD.n99 VSS 0.0014f
C6314 VDD.n100 VSS 0.00308f
C6315 VDD.t530 VSS 9.42e-19
C6316 VDD.t542 VSS 9.42e-19
C6317 VDD.n101 VSS 0.00214f
C6318 VDD.n102 VSS 0.00258f
C6319 VDD.t541 VSS 0.00553f
C6320 VDD.n103 VSS 0.00528f
C6321 VDD.n104 VSS 0.00109f
C6322 VDD.n105 VSS 0.0014f
C6323 VDD.n106 VSS 0.00236f
C6324 VDD.n107 VSS 0.00154f
C6325 VDD.t525 VSS 0.00578f
C6326 VDD.n108 VSS 0.00528f
C6327 VDD.n109 VSS 0.00109f
C6328 VDD.t526 VSS 9.42e-19
C6329 VDD.t536 VSS 9.42e-19
C6330 VDD.n110 VSS 0.00214f
C6331 VDD.n111 VSS 0.00258f
C6332 VDD.n112 VSS 0.00123f
C6333 VDD.n113 VSS 0.00226f
C6334 VDD.t535 VSS 0.00578f
C6335 VDD.n114 VSS 0.00528f
C6336 VDD.n115 VSS 0.00109f
C6337 VDD.n116 VSS 0.00142f
C6338 VDD.n117 VSS 0.00241f
C6339 VDD.n118 VSS 9.04e-19
C6340 VDD.t533 VSS 0.00578f
C6341 VDD.n119 VSS 0.00528f
C6342 VDD.n120 VSS 0.00109f
C6343 VDD.n121 VSS 0.0017f
C6344 VDD.n122 VSS 0.00303f
C6345 VDD.n123 VSS 0.00154f
C6346 VDD.t522 VSS 9.42e-19
C6347 VDD.t534 VSS 9.42e-19
C6348 VDD.n124 VSS 0.00214f
C6349 VDD.n125 VSS 0.00255f
C6350 VDD.n126 VSS 1.42e-19
C6351 VDD.t521 VSS 0.00578f
C6352 VDD.n127 VSS 0.00528f
C6353 VDD.n128 VSS 0.00109f
C6354 VDD.n129 VSS 1.72e-19
C6355 VDD.n130 VSS 2.85e-19
C6356 VDD.n131 VSS 9.31e-19
C6357 VDD.n132 VSS 6.37e-19
C6358 VDD.n133 VSS 4.35e-19
C6359 VDD.n134 VSS 3.36e-19
C6360 VDD.n135 VSS 8.1e-19
C6361 VDD.n136 VSS 0.00157f
C6362 VDD.n137 VSS 4.85e-19
C6363 VDD.n138 VSS 5.59e-19
C6364 VDD.n139 VSS 0.00154f
C6365 VDD.n140 VSS 6.68e-19
C6366 VDD.t660 VSS 0.00578f
C6367 VDD.n141 VSS 0.00528f
C6368 VDD.n142 VSS 0.00109f
C6369 VDD.n143 VSS 1.72e-19
C6370 VDD.n144 VSS 2.85e-19
C6371 VDD.n145 VSS 9.31e-19
C6372 VDD.n146 VSS 2.85e-19
C6373 VDD.n147 VSS 0.00126f
C6374 VDD.n148 VSS 4.35e-19
C6375 VDD.n149 VSS 5.54e-19
C6376 VDD.n150 VSS 3.36e-19
C6377 VDD.n151 VSS 0.00149f
C6378 VDD.n152 VSS 8.1e-19
C6379 VDD.n153 VSS 0.00157f
C6380 VDD.n154 VSS 4.84e-19
C6381 VDD.n155 VSS 0.00158f
C6382 VDD.n156 VSS 8.1e-19
C6383 VDD.n157 VSS 0.00144f
C6384 VDD.n158 VSS 0.00148f
C6385 VDD.n159 VSS 0.00654f
C6386 VDD.n160 VSS 0.00653f
C6387 VDD.n161 VSS 4.84e-19
C6388 VDD.n162 VSS 4.84e-19
C6389 VDD.n163 VSS 4.84e-19
C6390 VDD.n164 VSS 0.00846f
C6391 VDD.n165 VSS 0.00157f
C6392 VDD.n166 VSS 0.00158f
C6393 VDD.n167 VSS 8.1e-19
C6394 VDD.n168 VSS 0.00148f
C6395 VDD.n169 VSS 0.0058f
C6396 VDD.n170 VSS 0.00158f
C6397 VDD.n171 VSS 6.05e-19
C6398 VDD.t298 VSS 7.73e-19
C6399 VDD.t336 VSS 2.51e-19
C6400 VDD.n172 VSS 0.00395f
C6401 VDD.n173 VSS 0.00308f
C6402 VDD.n174 VSS 0.00149f
C6403 VDD.n175 VSS 0.0148f
C6404 VDD.n176 VSS 0.00158f
C6405 VDD.n177 VSS 0.00149f
C6406 VDD.n178 VSS 4.52e-19
C6407 VDD.n179 VSS 6.55e-19
C6408 VDD.t258 VSS 6.03e-19
C6409 VDD.t597 VSS 6.03e-19
C6410 VDD.n180 VSS 0.0013f
C6411 VDD.n181 VSS 0.00882f
C6412 VDD.n182 VSS 5.77e-19
C6413 VDD.n183 VSS 2.18e-19
C6414 VDD.n184 VSS 6.55e-19
C6415 VDD.n185 VSS 0.00158f
C6416 VDD.n186 VSS 0.0256f
C6417 VDD.n187 VSS 0.0148f
C6418 VDD.n188 VSS 0.00158f
C6419 VDD.n189 VSS 6.93e-19
C6420 VDD.n190 VSS 5.86e-19
C6421 VDD.n191 VSS 0.00127f
C6422 VDD.n192 VSS 7.49e-19
C6423 VDD.n193 VSS 7.49e-19
C6424 VDD.n194 VSS 1.72e-19
C6425 VDD.n195 VSS 5.4e-19
C6426 VDD.n196 VSS 1.01e-19
C6427 VDD.t398 VSS 0.00476f
C6428 VDD.n197 VSS 0.0047f
C6429 VDD.n198 VSS 0.00108f
C6430 VDD.n199 VSS 0.00184f
C6431 VDD.n200 VSS 4.51e-19
C6432 VDD.n201 VSS 2.02e-20
C6433 VDD.n202 VSS 1.72e-19
C6434 VDD.n203 VSS 2.85e-19
C6435 VDD.n204 VSS 0.00151f
C6436 VDD.n205 VSS 0.00126f
C6437 VDD.n206 VSS 3.35e-20
C6438 VDD.n207 VSS 2.68e-19
C6439 VDD.n208 VSS 5.97e-19
C6440 VDD.t399 VSS 7.73e-19
C6441 VDD.t18 VSS 2.51e-19
C6442 VDD.n209 VSS 0.00395f
C6443 VDD.n210 VSS 7.49e-19
C6444 VDD.n211 VSS 1.72e-19
C6445 VDD.n212 VSS 5.4e-19
C6446 VDD.n213 VSS 1.01e-19
C6447 VDD.n214 VSS 5.4e-19
C6448 VDD.n215 VSS 1.01e-19
C6449 VDD.n216 VSS 8.97e-19
C6450 VDD.n217 VSS 4.35e-19
C6451 VDD.n218 VSS 0.0116f
C6452 VDD.n219 VSS 0.00109f
C6453 VDD.n220 VSS 0.0014f
C6454 VDD.t444 VSS 7.73e-19
C6455 VDD.t624 VSS 2.51e-19
C6456 VDD.n221 VSS 0.00395f
C6457 VDD.n222 VSS 7.29e-19
C6458 VDD.n223 VSS 0.00149f
C6459 VDD.n224 VSS 2.68e-19
C6460 VDD.n225 VSS 5.03e-20
C6461 VDD.n226 VSS 2.51e-19
C6462 VDD.n227 VSS 1.62e-19
C6463 VDD.n228 VSS 3.04e-20
C6464 VDD.n229 VSS 5.4e-19
C6465 VDD.n230 VSS 1.01e-19
C6466 VDD.t566 VSS 0.00476f
C6467 VDD.n231 VSS 0.00578f
C6468 VDD.n232 VSS 0.00108f
C6469 VDD.n233 VSS 0.00114f
C6470 VDD.n234 VSS 4.51e-19
C6471 VDD.n235 VSS 2.02e-20
C6472 VDD.n236 VSS 1.42e-19
C6473 VDD.n237 VSS 6.17e-19
C6474 VDD.n238 VSS 1.62e-19
C6475 VDD.n239 VSS 6.37e-19
C6476 VDD.n240 VSS 4.13e-19
C6477 VDD.n241 VSS 0.00158f
C6478 VDD.n242 VSS 0.00542f
C6479 VDD.n243 VSS 0.00158f
C6480 VDD.n244 VSS 6.55e-19
C6481 VDD.t616 VSS 0.00578f
C6482 VDD.n245 VSS 0.00754f
C6483 VDD.n246 VSS 0.00109f
C6484 VDD.n247 VSS 0.00177f
C6485 VDD.n248 VSS 0.00253f
C6486 VDD.n249 VSS 0.00139f
C6487 VDD.n250 VSS 5.03e-19
C6488 VDD.n251 VSS 6.05e-19
C6489 VDD.n252 VSS 0.00158f
C6490 VDD.n253 VSS 0.00149f
C6491 VDD.n254 VSS 0.0108f
C6492 VDD.n255 VSS 0.00158f
C6493 VDD.n256 VSS 0.00149f
C6494 VDD.n257 VSS 5.16e-19
C6495 VDD.n258 VSS 5.92e-19
C6496 VDD.n259 VSS 0.00124f
C6497 VDD.t163 VSS 7.73e-19
C6498 VDD.t268 VSS 2.51e-19
C6499 VDD.n260 VSS 0.00395f
C6500 VDD.n261 VSS 0.00276f
C6501 VDD.n262 VSS 6.07e-19
C6502 VDD.n263 VSS 1.72e-19
C6503 VDD.n264 VSS 4.57e-19
C6504 VDD.n265 VSS 1.01e-19
C6505 VDD.n266 VSS 4.57e-19
C6506 VDD.n267 VSS 1.01e-19
C6507 VDD.n268 VSS 6.41e-19
C6508 VDD.n269 VSS 2.35e-19
C6509 VDD.n270 VSS 6.48e-19
C6510 VDD.n271 VSS 1.72e-19
C6511 VDD.n272 VSS 1.01e-19
C6512 VDD.n273 VSS 0.00273f
C6513 VDD.n274 VSS 0.00108f
C6514 VDD.n275 VSS 4.81e-19
C6515 VDD.n276 VSS 1.01e-19
C6516 VDD.n277 VSS 6.48e-19
C6517 VDD.n278 VSS 1.72e-19
C6518 VDD.t711 VSS 7.73e-19
C6519 VDD.t676 VSS 2.51e-19
C6520 VDD.n279 VSS 0.00395f
C6521 VDD.n280 VSS 6.27e-19
C6522 VDD.n281 VSS 0.00221f
C6523 VDD.n282 VSS 0.00144f
C6524 VDD.n283 VSS 5.66e-19
C6525 VDD.n284 VSS 0.00158f
C6526 VDD.n285 VSS 0.0148f
C6527 VDD.n286 VSS 0.00158f
C6528 VDD.n287 VSS 0.00149f
C6529 VDD.n288 VSS 6.3e-19
C6530 VDD.t567 VSS 0.00578f
C6531 VDD.n289 VSS 0.00154f
C6532 VDD.n290 VSS 2.85e-19
C6533 VDD.t58 VSS 0.00578f
C6534 VDD.n291 VSS 0.00854f
C6535 VDD.n292 VSS 0.00111f
C6536 VDD.n293 VSS 0.002f
C6537 VDD.t59 VSS 0.00141f
C6538 VDD.n294 VSS 0.00295f
C6539 VDD.n295 VSS 2.1e-19
C6540 VDD.n296 VSS 5.86e-19
C6541 VDD.n297 VSS 4.39e-19
C6542 VDD.n298 VSS 0.00158f
C6543 VDD.n299 VSS 0.0571f
C6544 VDD.n300 VSS 0.00158f
C6545 VDD.n301 VSS 0.00149f
C6546 VDD.n302 VSS 6.93e-19
C6547 VDD.n303 VSS 0.0026f
C6548 VDD.n304 VSS 1.72e-19
C6549 VDD.n305 VSS 5.97e-19
C6550 VDD.n306 VSS 5.97e-19
C6551 VDD.n307 VSS 0.00124f
C6552 VDD.n308 VSS 2.02e-20
C6553 VDD.n309 VSS 5.97e-19
C6554 VDD.n310 VSS 1.72e-19
C6555 VDD.n311 VSS 4.51e-19
C6556 VDD.n312 VSS 1.01e-19
C6557 VDD.t602 VSS 7.73e-19
C6558 VDD.t232 VSS 2.51e-19
C6559 VDD.n313 VSS 0.00395f
C6560 VDD.n314 VSS 0.00274f
C6561 VDD.n315 VSS 5.87e-19
C6562 VDD.n316 VSS 1.72e-19
C6563 VDD.n317 VSS 0.00889f
C6564 VDD.n318 VSS 4.51e-19
C6565 VDD.n319 VSS 1.01e-19
C6566 VDD.n320 VSS 0.00558f
C6567 VDD.n321 VSS 0.00461f
C6568 VDD.t231 VSS 0.00184f
C6569 VDD.n322 VSS 0.0021f
C6570 VDD.n323 VSS 0.00108f
C6571 VDD.n324 VSS 0.00394f
C6572 VDD.n325 VSS 5.4e-19
C6573 VDD.n326 VSS 3.24e-19
C6574 VDD.n327 VSS 1.72e-19
C6575 VDD.n328 VSS 2.85e-19
C6576 VDD.n329 VSS 0.00152f
C6577 VDD.n330 VSS 0.00127f
C6578 VDD.n331 VSS 5.97e-19
C6579 VDD.n332 VSS 5.97e-19
C6580 VDD.n333 VSS 1.72e-19
C6581 VDD.n334 VSS 4.51e-19
C6582 VDD.n335 VSS 1.01e-19
C6583 VDD.t601 VSS 0.00476f
C6584 VDD.n336 VSS 0.00279f
C6585 VDD.n337 VSS 0.00108f
C6586 VDD.n338 VSS 0.00375f
C6587 VDD.n339 VSS 5.4e-19
C6588 VDD.n340 VSS 3.24e-19
C6589 VDD.n341 VSS 1.72e-19
C6590 VDD.n342 VSS 2.85e-19
C6591 VDD.n343 VSS 0.00152f
C6592 VDD.n344 VSS 0.00127f
C6593 VDD.n345 VSS 5.97e-19
C6594 VDD.n346 VSS 5.97e-19
C6595 VDD.n347 VSS 1.72e-19
C6596 VDD.n348 VSS 4.51e-19
C6597 VDD.n349 VSS 1.01e-19
C6598 VDD.t564 VSS 0.00476f
C6599 VDD.n350 VSS 0.00483f
C6600 VDD.n351 VSS 0.00108f
C6601 VDD.n352 VSS 0.00305f
C6602 VDD.n353 VSS 5.4e-19
C6603 VDD.n354 VSS 3.24e-19
C6604 VDD.n355 VSS 1.72e-19
C6605 VDD.n356 VSS 2.85e-19
C6606 VDD.n357 VSS 0.00152f
C6607 VDD.n358 VSS 0.00127f
C6608 VDD.n359 VSS 5.97e-19
C6609 VDD.n360 VSS 5.97e-19
C6610 VDD.n361 VSS 1.72e-19
C6611 VDD.n362 VSS 4.51e-19
C6612 VDD.n363 VSS 1.01e-19
C6613 VDD.n364 VSS 0.0047f
C6614 VDD.n365 VSS 0.00108f
C6615 VDD.n366 VSS 0.00578f
C6616 VDD.n367 VSS 5.4e-19
C6617 VDD.n368 VSS 3.24e-19
C6618 VDD.n369 VSS 1.72e-19
C6619 VDD.n370 VSS 2.85e-19
C6620 VDD.n371 VSS 0.00152f
C6621 VDD.n372 VSS 0.00127f
C6622 VDD.n373 VSS 5.97e-19
C6623 VDD.n374 VSS 5.97e-19
C6624 VDD.n375 VSS 1.72e-19
C6625 VDD.n376 VSS 4.51e-19
C6626 VDD.n377 VSS 1.01e-19
C6627 VDD.t281 VSS 0.00476f
C6628 VDD.n378 VSS 0.00343f
C6629 VDD.n379 VSS 0.00108f
C6630 VDD.n380 VSS 0.00114f
C6631 VDD.n381 VSS 5.4e-19
C6632 VDD.n382 VSS 3.24e-19
C6633 VDD.n383 VSS 1.72e-19
C6634 VDD.n384 VSS 2.85e-19
C6635 VDD.n385 VSS 0.00152f
C6636 VDD.n386 VSS 0.00127f
C6637 VDD.n387 VSS 5.97e-19
C6638 VDD.n388 VSS 1.42e-19
C6639 VDD.n389 VSS 1.72e-19
C6640 VDD.n390 VSS 4.51e-19
C6641 VDD.n391 VSS 1.01e-19
C6642 VDD.t323 VSS 0.00476f
C6643 VDD.n392 VSS 0.00368f
C6644 VDD.n393 VSS 0.00108f
C6645 VDD.n394 VSS 0.00241f
C6646 VDD.n395 VSS 5.4e-19
C6647 VDD.n396 VSS 3.24e-19
C6648 VDD.n397 VSS 1.72e-19
C6649 VDD.n398 VSS 2.85e-19
C6650 VDD.n399 VSS 0.00152f
C6651 VDD.n400 VSS 0.00127f
C6652 VDD.t324 VSS 5.42e-19
C6653 VDD.t175 VSS 4.25e-19
C6654 VDD.n401 VSS 0.00111f
C6655 VDD.n402 VSS 0.00224f
C6656 VDD.n403 VSS 4.66e-19
C6657 VDD.n404 VSS 4.51e-19
C6658 VDD.n405 VSS 1.01e-19
C6659 VDD.t174 VSS 0.00476f
C6660 VDD.n406 VSS 0.00483f
C6661 VDD.n407 VSS 0.00108f
C6662 VDD.n408 VSS 0.00216f
C6663 VDD.n409 VSS 5.4e-19
C6664 VDD.n410 VSS 3.24e-19
C6665 VDD.n411 VSS 1.72e-19
C6666 VDD.n412 VSS 2.85e-19
C6667 VDD.n413 VSS 0.00152f
C6668 VDD.n414 VSS 0.00127f
C6669 VDD.n415 VSS 0.00158f
C6670 VDD.n416 VSS 0.0921f
C6671 VDD.n417 VSS 0.0123f
C6672 VDD.n418 VSS 0.00158f
C6673 VDD.n419 VSS 0.00149f
C6674 VDD.n420 VSS 5.03e-19
C6675 VDD.n421 VSS 0.0138f
C6676 VDD.n422 VSS 0.00196f
C6677 VDD.t15 VSS -2.71e-19
C6678 VDD.t312 VSS 8.49e-19
C6679 VDD.n423 VSS 0.00391f
C6680 VDD.n424 VSS 0.00413f
C6681 VDD.t14 VSS 0.00663f
C6682 VDD.n425 VSS 0.00597f
C6683 VDD.n426 VSS 0.00109f
C6684 VDD.n427 VSS 9.92e-19
C6685 VDD.n428 VSS 0.00727f
C6686 VDD.t311 VSS 0.00578f
C6687 VDD.n429 VSS 0.00835f
C6688 VDD.n430 VSS 0.00109f
C6689 VDD.n431 VSS 0.00186f
C6690 VDD.n432 VSS 0.00308f
C6691 VDD.t315 VSS 0.00955f
C6692 VDD.n433 VSS 0.00923f
C6693 VDD.n434 VSS 6.76e-19
C6694 VDD.n435 VSS 0.00179f
C6695 VDD.n436 VSS 0.00308f
C6696 VDD.t316 VSS -5.07e-19
C6697 VDD.t107 VSS 9.16e-19
C6698 VDD.n437 VSS 0.00359f
C6699 VDD.n438 VSS 0.002f
C6700 VDD.n439 VSS 0.00187f
C6701 VDD.n440 VSS 0.00281f
C6702 VDD.n441 VSS 0.00152f
C6703 VDD.t768 VSS 8.67e-19
C6704 VDD.n442 VSS 0.00281f
C6705 VDD.t105 VSS 0.00159f
C6706 VDD.n443 VSS 0.0034f
C6707 VDD.n444 VSS 7.55e-19
C6708 VDD.n445 VSS 0.00215f
C6709 VDD.n446 VSS 3.97e-19
C6710 VDD.n447 VSS 2.85e-19
C6711 VDD.n448 VSS 0.00154f
C6712 VDD.t503 VSS 0.00262f
C6713 VDD.n449 VSS 0.00271f
C6714 VDD.t106 VSS 0.0139f
C6715 VDD.n450 VSS 0.0119f
C6716 VDD.n451 VSS 7.81e-19
C6717 VDD.n452 VSS 0.00267f
C6718 VDD.n453 VSS 0.00307f
C6719 VDD.t502 VSS 0.00578f
C6720 VDD.t647 VSS 0.00578f
C6721 VDD.n454 VSS 0.00452f
C6722 VDD.n455 VSS 0.00109f
C6723 VDD.n456 VSS 0.00172f
C6724 VDD.n457 VSS 0.00308f
C6725 VDD.n458 VSS 0.00666f
C6726 VDD.n459 VSS 0.00109f
C6727 VDD.n460 VSS 0.00164f
C6728 VDD.n461 VSS 0.00308f
C6729 VDD.t580 VSS 5.72e-19
C6730 VDD.t314 VSS 7.62e-19
C6731 VDD.n462 VSS 0.0014f
C6732 VDD.t579 VSS 0.00578f
C6733 VDD.n463 VSS 0.0076f
C6734 VDD.n464 VSS 0.00111f
C6735 VDD.n465 VSS 0.00204f
C6736 VDD.n466 VSS 0.00252f
C6737 VDD.n467 VSS 0.00308f
C6738 VDD.t313 VSS 0.00578f
C6739 VDD.n468 VSS 0.00603f
C6740 VDD.n469 VSS 0.00109f
C6741 VDD.n470 VSS 0.00132f
C6742 VDD.n471 VSS 0.00308f
C6743 VDD.t625 VSS 0.00578f
C6744 VDD.n472 VSS 0.00634f
C6745 VDD.n473 VSS 0.00109f
C6746 VDD.n474 VSS 0.00178f
C6747 VDD.n475 VSS 0.00295f
C6748 VDD.n476 VSS 0.00154f
C6749 VDD.n477 VSS 9.31e-19
C6750 VDD.t638 VSS 0.00578f
C6751 VDD.n478 VSS 0.00528f
C6752 VDD.n479 VSS 0.00109f
C6753 VDD.n480 VSS 1.72e-19
C6754 VDD.n481 VSS 2.85e-19
C6755 VDD.n482 VSS 9.31e-19
C6756 VDD.n483 VSS 4.35e-19
C6757 VDD.n484 VSS 0.00905f
C6758 VDD.n485 VSS 0.00109f
C6759 VDD.n486 VSS 0.00177f
C6760 VDD.n487 VSS 0.0025f
C6761 VDD.n488 VSS 0.00111f
C6762 VDD.n489 VSS 4.35e-19
C6763 VDD.n490 VSS 6.05e-19
C6764 VDD.n491 VSS 3.36e-19
C6765 VDD.n492 VSS 8.1e-19
C6766 VDD.n493 VSS 0.00158f
C6767 VDD.n494 VSS 0.00149f
C6768 VDD.n495 VSS 4.77e-19
C6769 VDD.t642 VSS 6.03e-19
C6770 VDD.t240 VSS 6.03e-19
C6771 VDD.n496 VSS 0.0013f
C6772 VDD.n497 VSS 0.00153f
C6773 VDD.n498 VSS 0.00109f
C6774 VDD.t641 VSS 0.00472f
C6775 VDD.t239 VSS 0.00579f
C6776 VDD.n499 VSS 0.00529f
C6777 VDD.n500 VSS 0.00111f
C6778 VDD.n501 VSS 0.00202f
C6779 VDD.n502 VSS 0.0027f
C6780 VDD.n503 VSS 0.0028f
C6781 VDD.n504 VSS 0.00907f
C6782 VDD.n505 VSS 0.00109f
C6783 VDD.n506 VSS 0.00118f
C6784 VDD.n507 VSS 0.00308f
C6785 VDD.t165 VSS 0.00142f
C6786 VDD.t164 VSS 0.00579f
C6787 VDD.n508 VSS 0.00857f
C6788 VDD.n509 VSS 0.00111f
C6789 VDD.n510 VSS 0.00203f
C6790 VDD.n511 VSS 0.00312f
C6791 VDD.n512 VSS 0.00308f
C6792 VDD.t241 VSS 0.00579f
C6793 VDD.n513 VSS 0.00579f
C6794 VDD.n514 VSS 0.00109f
C6795 VDD.n515 VSS 0.00151f
C6796 VDD.n516 VSS 0.00308f
C6797 VDD.t690 VSS 0.00579f
C6798 VDD.n517 VSS 0.00529f
C6799 VDD.n518 VSS 0.00109f
C6800 VDD.n519 VSS 0.00186f
C6801 VDD.n520 VSS 0.00308f
C6802 VDD.t666 VSS 0.0107f
C6803 VDD.n521 VSS 0.00756f
C6804 VDD.n522 VSS 0.00191f
C6805 VDD.n523 VSS 0.00177f
C6806 VDD.n524 VSS 0.00308f
C6807 VDD.n525 VSS 0.00198f
C6808 VDD.t667 VSS 5.42e-19
C6809 VDD.t101 VSS 5.72e-19
C6810 VDD.n526 VSS 0.00119f
C6811 VDD.n527 VSS 0.00282f
C6812 VDD.n528 VSS 0.00296f
C6813 VDD.n529 VSS 0.0015f
C6814 VDD.n530 VSS 1.36e-19
C6815 VDD.t135 VSS 0.00149f
C6816 VDD.t759 VSS 6.37e-19
C6817 VDD.n531 VSS 0.00279f
C6818 VDD.n532 VSS 2.33e-19
C6819 VDD.n533 VSS 6.77e-19
C6820 VDD.n534 VSS 0.00141f
C6821 VDD.n535 VSS 2.33e-19
C6822 VDD.n536 VSS 0.00388f
C6823 VDD.n537 VSS 5.31e-19
C6824 VDD.n538 VSS 0.00105f
C6825 VDD.t766 VSS 6.29e-19
C6826 VDD.n539 VSS 0.00315f
C6827 VDD.t99 VSS 0.00188f
C6828 VDD.n540 VSS 0.00172f
C6829 VDD.n541 VSS 2.3e-19
C6830 VDD.n542 VSS 9.31e-19
C6831 VDD.n543 VSS 1.72e-19
C6832 VDD.n544 VSS 2.85e-19
C6833 VDD.n545 VSS 0.00154f
C6834 VDD.t100 VSS 0.0134f
C6835 VDD.t600 VSS 0.00542f
C6836 VDD.n546 VSS 0.0068f
C6837 VDD.n547 VSS 0.00115f
C6838 VDD.n548 VSS 0.00176f
C6839 VDD.n549 VSS 0.00291f
C6840 VDD.t7 VSS 9.67e-19
C6841 VDD.t665 VSS 0.00217f
C6842 VDD.n550 VSS 0.00349f
C6843 VDD.n551 VSS 0.00457f
C6844 VDD.t6 VSS 0.00567f
C6845 VDD.n552 VSS 0.00617f
C6846 VDD.n553 VSS 0.00109f
C6847 VDD.n554 VSS 0.00102f
C6848 VDD.n555 VSS 0.00308f
C6849 VDD.t664 VSS 0.00579f
C6850 VDD.n556 VSS 0.00825f
C6851 VDD.n557 VSS 0.00109f
C6852 VDD.n558 VSS 0.00103f
C6853 VDD.n559 VSS 0.00296f
C6854 VDD.n560 VSS 0.00154f
C6855 VDD.n561 VSS 9.31e-19
C6856 VDD.n562 VSS 0.00907f
C6857 VDD.n563 VSS 0.00109f
C6858 VDD.n564 VSS 1.72e-19
C6859 VDD.n565 VSS 2.85e-19
C6860 VDD.n566 VSS 9.31e-19
C6861 VDD.n567 VSS 4.86e-19
C6862 VDD.t242 VSS 0.00579f
C6863 VDD.n568 VSS 0.00636f
C6864 VDD.n569 VSS 0.00109f
C6865 VDD.n570 VSS 0.00186f
C6866 VDD.n571 VSS 0.00308f
C6867 VDD.t691 VSS 0.00579f
C6868 VDD.n572 VSS 0.00529f
C6869 VDD.n573 VSS 0.00109f
C6870 VDD.n574 VSS 0.00176f
C6871 VDD.n575 VSS 0.00248f
C6872 VDD.n576 VSS 0.00106f
C6873 VDD.n577 VSS 4.35e-19
C6874 VDD.n578 VSS 6.3e-19
C6875 VDD.n579 VSS 3.36e-19
C6876 VDD.n580 VSS 8.1e-19
C6877 VDD.n581 VSS 0.00158f
C6878 VDD.n582 VSS 0.00717f
C6879 VDD.n583 VSS 0.00144f
C6880 VDD.n584 VSS 0.00148f
C6881 VDD.n585 VSS 8.1e-19
C6882 VDD.n586 VSS 0.00158f
C6883 VDD.n587 VSS 0.00149f
C6884 VDD.n588 VSS 4.77e-19
C6885 VDD.t747 VSS 0.00578f
C6886 VDD.n589 VSS 0.00823f
C6887 VDD.n590 VSS 0.00109f
C6888 VDD.n591 VSS 0.0011f
C6889 VDD.n592 VSS 0.00298f
C6890 VDD.n593 VSS 0.00154f
C6891 VDD.t748 VSS 0.00217f
C6892 VDD.t501 VSS 9.67e-19
C6893 VDD.n594 VSS 0.00349f
C6894 VDD.n595 VSS 0.0045f
C6895 VDD.n596 VSS 9.11e-20
C6896 VDD.t500 VSS 0.00565f
C6897 VDD.n597 VSS 0.00616f
C6898 VDD.n598 VSS 0.00109f
C6899 VDD.n599 VSS 1.72e-19
C6900 VDD.n600 VSS 2.85e-19
C6901 VDD.n601 VSS 9.31e-19
C6902 VDD.n602 VSS 5.03e-19
C6903 VDD.t581 VSS 0.0054f
C6904 VDD.n603 VSS 0.0059f
C6905 VDD.n604 VSS 0.00109f
C6906 VDD.n605 VSS 0.00175f
C6907 VDD.n606 VSS 0.00246f
C6908 VDD.n607 VSS 0.00104f
C6909 VDD.n608 VSS 4.35e-19
C6910 VDD.n609 VSS 6.3e-19
C6911 VDD.n610 VSS 3.36e-19
C6912 VDD.n611 VSS 8.1e-19
C6913 VDD.n612 VSS 0.00158f
C6914 VDD.n613 VSS 0.00144f
C6915 VDD.n614 VSS 0.00148f
C6916 VDD.n615 VSS 8.1e-19
C6917 VDD.n616 VSS 0.00158f
C6918 VDD.n617 VSS 0.00149f
C6919 VDD.n618 VSS 6.8e-19
C6920 VDD.t0 VSS 0.00578f
C6921 VDD.n619 VSS 0.00666f
C6922 VDD.n620 VSS 0.00109f
C6923 VDD.n621 VSS 0.00118f
C6924 VDD.n622 VSS 0.00241f
C6925 VDD.n623 VSS 9.21e-19
C6926 VDD.n624 VSS 0.00154f
C6927 VDD.n625 VSS 2.85e-19
C6928 VDD.t745 VSS 0.00578f
C6929 VDD.n626 VSS 0.00666f
C6930 VDD.n627 VSS 0.00111f
C6931 VDD.n628 VSS 0.00201f
C6932 VDD.t1 VSS 5.72e-19
C6933 VDD.t746 VSS 5.42e-19
C6934 VDD.n629 VSS 0.00118f
C6935 VDD.n630 VSS 0.0026f
C6936 VDD.n631 VSS 2.25e-19
C6937 VDD.n632 VSS 6.2e-19
C6938 VDD.n633 VSS 4.35e-19
C6939 VDD.n634 VSS 4.26e-19
C6940 VDD.n635 VSS 3.36e-19
C6941 VDD.n636 VSS 8.1e-19
C6942 VDD.n637 VSS 0.00158f
C6943 VDD.n638 VSS 0.00149f
C6944 VDD.n639 VSS 4.9e-19
C6945 VDD.n640 VSS 3.23e-19
C6946 VDD.n641 VSS 3.23e-19
C6947 VDD.n642 VSS 3.1e-19
C6948 VDD.n643 VSS 8.1e-19
C6949 VDD.n644 VSS 0.00158f
C6950 VDD.n645 VSS 0.00144f
C6951 VDD.n646 VSS 0.00148f
C6952 VDD.n647 VSS 8.1e-19
C6953 VDD.n648 VSS 0.00158f
C6954 VDD.n649 VSS 0.00149f
C6955 VDD.n650 VSS 5.41e-19
C6956 VDD.n651 VSS 5.66e-19
C6957 VDD.n652 VSS 0.00754f
C6958 VDD.n653 VSS 0.00109f
C6959 VDD.n654 VSS 0.00175f
C6960 VDD.n655 VSS 0.00256f
C6961 VDD.n656 VSS 0.00131f
C6962 VDD.t628 VSS 0.00578f
C6963 VDD.n657 VSS 0.00578f
C6964 VDD.n658 VSS 0.00109f
C6965 VDD.n659 VSS 0.00136f
C6966 VDD.n660 VSS 0.00276f
C6967 VDD.n661 VSS 0.00154f
C6968 VDD.t637 VSS 0.00578f
C6969 VDD.n662 VSS 0.00528f
C6970 VDD.n663 VSS 0.00109f
C6971 VDD.n664 VSS 9.31e-19
C6972 VDD.n665 VSS 1.72e-19
C6973 VDD.n666 VSS 2.85e-19
C6974 VDD.n667 VSS 9.31e-19
C6975 VDD.n668 VSS 2.35e-19
C6976 VDD.n669 VSS 4.35e-19
C6977 VDD.n670 VSS 3.36e-19
C6978 VDD.n671 VSS 8.1e-19
C6979 VDD.n672 VSS 0.00158f
C6980 VDD.n673 VSS 0.00149f
C6981 VDD.n674 VSS 4.52e-19
C6982 VDD.t44 VSS 0.00579f
C6983 VDD.n675 VSS 0.00605f
C6984 VDD.n676 VSS 0.00109f
C6985 VDD.n677 VSS 0.00132f
C6986 VDD.n678 VSS 0.00236f
C6987 VDD.n679 VSS 0.00154f
C6988 VDD.t45 VSS 7.62e-19
C6989 VDD.t137 VSS 5.72e-19
C6990 VDD.n680 VSS 0.0014f
C6991 VDD.t136 VSS 0.00579f
C6992 VDD.n681 VSS 0.00762f
C6993 VDD.n682 VSS 0.00111f
C6994 VDD.n683 VSS 0.00204f
C6995 VDD.n684 VSS 0.00252f
C6996 VDD.n685 VSS 0.00226f
C6997 VDD.n686 VSS 0.00668f
C6998 VDD.n687 VSS 0.00109f
C6999 VDD.n688 VSS 0.00164f
C7000 VDD.n689 VSS 0.00268f
C7001 VDD.n690 VSS 0.00144f
C7002 VDD.n691 VSS 4.02e-19
C7003 VDD.t648 VSS 0.00579f
C7004 VDD.t4 VSS 0.00579f
C7005 VDD.n692 VSS 0.00453f
C7006 VDD.n693 VSS 0.00109f
C7007 VDD.n694 VSS 0.00172f
C7008 VDD.n695 VSS 4.19e-19
C7009 VDD.n696 VSS 0.00154f
C7010 VDD.t5 VSS 0.00262f
C7011 VDD.n697 VSS 0.00271f
C7012 VDD.n698 VSS 0.00882f
C7013 VDD.n699 VSS 9.91e-19
C7014 VDD.n700 VSS 0.00229f
C7015 VDD.n701 VSS 0.00241f
C7016 VDD.n702 VSS 0.00154f
C7017 VDD.t46 VSS 0.00579f
C7018 VDD.n703 VSS 0.00838f
C7019 VDD.n704 VSS 0.00109f
C7020 VDD.n705 VSS 0.00182f
C7021 VDD.n706 VSS 0.00258f
C7022 VDD.n707 VSS 0.00127f
C7023 VDD.n708 VSS 4.35e-19
C7024 VDD.n709 VSS 9.31e-19
C7025 VDD.n710 VSS 2.68e-19
C7026 VDD.n711 VSS 7.06e-19
C7027 VDD.n712 VSS 0.00926f
C7028 VDD.n713 VSS 9.85e-19
C7029 VDD.n714 VSS 1.72e-19
C7030 VDD.n715 VSS 2.85e-19
C7031 VDD.n716 VSS 0.00152f
C7032 VDD.n717 VSS 0.00132f
C7033 VDD.n718 VSS 0.00164f
C7034 VDD.t270 VSS 9.16e-19
C7035 VDD.t43 VSS -5.07e-19
C7036 VDD.n719 VSS 0.00359f
C7037 VDD.n720 VSS 6.69e-19
C7038 VDD.n721 VSS 0.00132f
C7039 VDD.n722 VSS 5.4e-19
C7040 VDD.t42 VSS 0.00466f
C7041 VDD.n723 VSS 0.00227f
C7042 VDD.n724 VSS 0.00491f
C7043 VDD.n725 VSS 6.53e-19
C7044 VDD.n726 VSS 4.21e-19
C7045 VDD.n727 VSS 1.4e-19
C7046 VDD.n728 VSS 2.85e-19
C7047 VDD.n729 VSS 0.00117f
C7048 VDD.n730 VSS 9.88e-19
C7049 VDD.n731 VSS 3.68e-19
C7050 VDD.n732 VSS 0.00213f
C7051 VDD.n733 VSS 3.97e-19
C7052 VDD.n734 VSS 0.00178f
C7053 VDD.n735 VSS 5.4e-19
C7054 VDD.n736 VSS 1.01e-19
C7055 VDD.n737 VSS 0.00573f
C7056 VDD.n738 VSS 0.00107f
C7057 VDD.t269 VSS 0.00586f
C7058 VDD.n739 VSS 0.00208f
C7059 VDD.n740 VSS 5.58e-19
C7060 VDD.n741 VSS 4.21e-19
C7061 VDD.n742 VSS 6.37e-19
C7062 VDD.n743 VSS 4.39e-19
C7063 VDD.n744 VSS 5.55e-19
C7064 VDD.n745 VSS 8.1e-19
C7065 VDD.n746 VSS 0.0493f
C7066 VDD.n747 VSS 0.0148f
C7067 VDD.n748 VSS 0.0148f
C7068 VDD.n749 VSS 0.0148f
C7069 VDD.n750 VSS 0.0148f
C7070 VDD.n751 VSS 0.0399f
C7071 VDD.n752 VSS 0.0478f
C7072 VDD.n753 VSS 0.0241f
C7073 VDD.n754 VSS 0.0148f
C7074 VDD.n755 VSS 0.0148f
C7075 VDD.n756 VSS 0.00985f
C7076 VDD.n757 VSS 0.0148f
C7077 VDD.n758 VSS 0.0148f
C7078 VDD.n759 VSS 0.0153f
C7079 VDD.n760 VSS 0.0788f
C7080 VDD.n761 VSS 0.0734f
C7081 VDD.n762 VSS 0.00985f
C7082 VDD.n763 VSS 0.00542f
C7083 VDD.n764 VSS 0.0143f
C7084 VDD.n765 VSS 0.00985f
C7085 VDD.n766 VSS 0.00542f
C7086 VDD.n767 VSS 0.0143f
C7087 VDD.n768 VSS 0.00985f
C7088 VDD.n769 VSS 0.107f
C7089 VDD.n770 VSS 0.108f
C7090 VDD.n771 VSS 0.00394f
C7091 VDD.n772 VSS 0.0133f
C7092 VDD.n773 VSS 0.0123f
C7093 VDD.n774 VSS 0.00394f
C7094 VDD.n775 VSS 0.0133f
C7095 VDD.n776 VSS 8.1e-19
C7096 VDD.n777 VSS 0.00148f
C7097 VDD.n778 VSS 0.00144f
C7098 VDD.n779 VSS 0.00832f
C7099 VDD.n780 VSS 7.71e-19
C7100 VDD.n781 VSS 2.85e-19
C7101 VDD.n782 VSS 1.72e-19
C7102 VDD.n783 VSS 5.46e-19
C7103 VDD.n784 VSS 1.01e-19
C7104 VDD.n785 VSS 0.00584f
C7105 VDD.n786 VSS 0.00108f
C7106 VDD.n787 VSS 0.00578f
C7107 VDD.n788 VSS 5.4e-19
C7108 VDD.n789 VSS 3.24e-19
C7109 VDD.n790 VSS 1.72e-19
C7110 VDD.n791 VSS 8.42e-19
C7111 VDD.n792 VSS 0.0116f
C7112 VDD.n793 VSS 0.00109f
C7113 VDD.n794 VSS 0.00155f
C7114 VDD.n795 VSS 0.0117f
C7115 VDD.n796 VSS 0.00109f
C7116 VDD.n797 VSS 0.00157f
C7117 VDD.n798 VSS 0.0117f
C7118 VDD.n799 VSS 0.00109f
C7119 VDD.n800 VSS 0.00157f
C7120 VDD.n801 VSS 0.0117f
C7121 VDD.n802 VSS 0.00109f
C7122 VDD.n803 VSS 0.00157f
C7123 VDD.n804 VSS 0.0117f
C7124 VDD.n805 VSS 0.00109f
C7125 VDD.n806 VSS 0.00157f
C7126 VDD.n807 VSS 0.0113f
C7127 VDD.n808 VSS 0.00106f
C7128 VDD.n809 VSS 0.00151f
C7129 VDD.n810 VSS 8.67e-19
C7130 VDD.n811 VSS 1.72e-19
C7131 VDD.n812 VSS 5.46e-19
C7132 VDD.n813 VSS 1.01e-19
C7133 VDD.n814 VSS 0.00584f
C7134 VDD.n815 VSS 0.00108f
C7135 VDD.n816 VSS 0.00546f
C7136 VDD.n817 VSS 5.1e-19
C7137 VDD.n818 VSS 2.23e-19
C7138 VDD.n819 VSS 6.48e-19
C7139 VDD.n820 VSS 1.72e-19
C7140 VDD.n821 VSS 2.85e-19
C7141 VDD.n822 VSS 0.00136f
C7142 VDD.n823 VSS 0.00144f
C7143 VDD.n824 VSS 6.48e-19
C7144 VDD.n825 VSS 1.72e-19
C7145 VDD.n826 VSS 4.81e-19
C7146 VDD.n827 VSS 1.01e-19
C7147 VDD.n828 VSS 0.00514f
C7148 VDD.n829 VSS 0.00108f
C7149 VDD.t639 VSS 0.00476f
C7150 VDD.n830 VSS 0.00152f
C7151 VDD.n831 VSS 5.1e-19
C7152 VDD.n832 VSS 2.23e-19
C7153 VDD.n833 VSS 4.66e-19
C7154 VDD.n834 VSS 1.72e-19
C7155 VDD.n835 VSS 2.85e-19
C7156 VDD.n836 VSS 7.2e-19
C7157 VDD.n837 VSS 0.00126f
C7158 VDD.n838 VSS 8.21e-19
C7159 VDD.t640 VSS 4.25e-19
C7160 VDD.t393 VSS 5.42e-19
C7161 VDD.n839 VSS 0.00111f
C7162 VDD.n840 VSS 0.00224f
C7163 VDD.n841 VSS 2.43e-19
C7164 VDD.n842 VSS 1.72e-19
C7165 VDD.n843 VSS 4.81e-19
C7166 VDD.n844 VSS 1.01e-19
C7167 VDD.n845 VSS 0.00432f
C7168 VDD.n846 VSS 0.00108f
C7169 VDD.t392 VSS 0.00476f
C7170 VDD.n847 VSS 0.00178f
C7171 VDD.n848 VSS 5.1e-19
C7172 VDD.n849 VSS 2.23e-19
C7173 VDD.n850 VSS 6.48e-19
C7174 VDD.n851 VSS 1.72e-19
C7175 VDD.n852 VSS 2.85e-19
C7176 VDD.n853 VSS 0.00136f
C7177 VDD.n854 VSS 0.00144f
C7178 VDD.n855 VSS 6.48e-19
C7179 VDD.n856 VSS 1.72e-19
C7180 VDD.n857 VSS 4.81e-19
C7181 VDD.n858 VSS 1.01e-19
C7182 VDD.n859 VSS 0.00406f
C7183 VDD.n860 VSS 8.89e-19
C7184 VDD.t34 VSS 6.99e-19
C7185 VDD.n861 VSS 0.00495f
C7186 VDD.n862 VSS 5.1e-19
C7187 VDD.n863 VSS 2.23e-19
C7188 VDD.n864 VSS 6.48e-19
C7189 VDD.n865 VSS 1.72e-19
C7190 VDD.n866 VSS 2.85e-19
C7191 VDD.n867 VSS 0.00136f
C7192 VDD.n868 VSS 0.00144f
C7193 VDD.n869 VSS 6.48e-19
C7194 VDD.n870 VSS 1.72e-19
C7195 VDD.n871 VSS 4.81e-19
C7196 VDD.n872 VSS 1.01e-19
C7197 VDD.n873 VSS 0.00514f
C7198 VDD.n874 VSS 0.00108f
C7199 VDD.n875 VSS 0.00546f
C7200 VDD.n876 VSS 5.1e-19
C7201 VDD.n877 VSS 2.23e-19
C7202 VDD.n878 VSS 6.48e-19
C7203 VDD.n879 VSS 1.72e-19
C7204 VDD.n880 VSS 2.85e-19
C7205 VDD.n881 VSS 8.71e-19
C7206 VDD.n882 VSS 8.04e-19
C7207 VDD.n883 VSS 0.00136f
C7208 VDD.n884 VSS 6.48e-19
C7209 VDD.n885 VSS 1.72e-19
C7210 VDD.n886 VSS 4.81e-19
C7211 VDD.n887 VSS 1.01e-19
C7212 VDD.n888 VSS 0.00343f
C7213 VDD.n889 VSS 0.00108f
C7214 VDD.t710 VSS 0.00476f
C7215 VDD.n890 VSS 0.00311f
C7216 VDD.n891 VSS 5.1e-19
C7217 VDD.n892 VSS 2.23e-19
C7218 VDD.n893 VSS 6.48e-19
C7219 VDD.n894 VSS 1.72e-19
C7220 VDD.n895 VSS 2.85e-19
C7221 VDD.n896 VSS 0.00144f
C7222 VDD.n897 VSS 0.00131f
C7223 VDD.n898 VSS 1.01e-19
C7224 VDD.n899 VSS 2.35e-19
C7225 VDD.n900 VSS 2.35e-19
C7226 VDD.n901 VSS 6.48e-19
C7227 VDD.n902 VSS 1.42e-19
C7228 VDD.n903 VSS 6.17e-19
C7229 VDD.n904 VSS 6.07e-20
C7230 VDD.n905 VSS 1.42e-19
C7231 VDD.n906 VSS 4.81e-19
C7232 VDD.n907 VSS 1.01e-19
C7233 VDD.n908 VSS 0.00514f
C7234 VDD.n909 VSS 0.00108f
C7235 VDD.t557 VSS 0.00476f
C7236 VDD.n910 VSS 0.00241f
C7237 VDD.n911 VSS 5.1e-19
C7238 VDD.n912 VSS 1.42e-19
C7239 VDD.n913 VSS 1.11e-19
C7240 VDD.n914 VSS 4.52e-19
C7241 VDD.n915 VSS 4.35e-19
C7242 VDD.n916 VSS 4.13e-19
C7243 VDD.n917 VSS 3.36e-19
C7244 VDD.n918 VSS 8.1e-19
C7245 VDD.n919 VSS 0.0266f
C7246 VDD.n920 VSS 0.0148f
C7247 VDD.n921 VSS 0.00936f
C7248 VDD.n922 VSS 0.0118f
C7249 VDD.n923 VSS 0.00158f
C7250 VDD.n924 VSS 0.00149f
C7251 VDD.n925 VSS 5.66e-19
C7252 VDD.n926 VSS 5.41e-19
C7253 VDD.n927 VSS 3.36e-19
C7254 VDD.n928 VSS 8.1e-19
C7255 VDD.n929 VSS 0.0148f
C7256 VDD.n930 VSS 0.0803f
C7257 VDD.n931 VSS 0.0892f
C7258 VDD.n932 VSS 0.0148f
C7259 VDD.n933 VSS 0.0148f
C7260 VDD.n934 VSS 0.00149f
C7261 VDD.n935 VSS 8.1e-19
C7262 VDD.n936 VSS 6.68e-19
C7263 VDD.n937 VSS 3.36e-19
C7264 VDD.n938 VSS 4.35e-19
C7265 VDD.n939 VSS 9.55e-19
C7266 VDD.n940 VSS 0.00905f
C7267 VDD.n941 VSS 0.00109f
C7268 VDD.n942 VSS 0.00118f
C7269 VDD.n943 VSS 0.00243f
C7270 VDD.t627 VSS 6.03e-19
C7271 VDD.t568 VSS 6.03e-19
C7272 VDD.n944 VSS 0.0013f
C7273 VDD.t626 VSS 0.00578f
C7274 VDD.n945 VSS 0.00528f
C7275 VDD.n946 VSS 0.00111f
C7276 VDD.n947 VSS 0.00202f
C7277 VDD.n948 VSS 0.0027f
C7278 VDD.n949 VSS 0.00308f
C7279 VDD.n950 VSS 0.00183f
C7280 VDD.n951 VSS 0.00151f
C7281 VDD.n952 VSS 0.00109f
C7282 VDD.n953 VSS 0.00773f
C7283 VDD.n954 VSS 0.00109f
C7284 VDD.n955 VSS 0.0018f
C7285 VDD.n956 VSS 0.00231f
C7286 VDD.t713 VSS -2.71e-19
C7287 VDD.t464 VSS 8.49e-19
C7288 VDD.n957 VSS 0.00391f
C7289 VDD.n958 VSS 0.00413f
C7290 VDD.t712 VSS 0.00578f
C7291 VDD.n959 VSS 0.00597f
C7292 VDD.n960 VSS 0.00109f
C7293 VDD.n961 VSS 9.92e-19
C7294 VDD.n962 VSS 0.00308f
C7295 VDD.t463 VSS 0.00578f
C7296 VDD.n963 VSS 0.00835f
C7297 VDD.n964 VSS 0.00109f
C7298 VDD.n965 VSS 0.00186f
C7299 VDD.n966 VSS 0.00308f
C7300 VDD.t461 VSS 0.00955f
C7301 VDD.n967 VSS 0.00923f
C7302 VDD.n968 VSS 6.76e-19
C7303 VDD.n969 VSS 0.00179f
C7304 VDD.n970 VSS 0.00308f
C7305 VDD.t462 VSS -5.07e-19
C7306 VDD.t95 VSS 9.16e-19
C7307 VDD.n971 VSS 0.00359f
C7308 VDD.n972 VSS 0.00204f
C7309 VDD.n973 VSS 0.00187f
C7310 VDD.n974 VSS 0.00281f
C7311 VDD.n975 VSS 0.00154f
C7312 VDD.t773 VSS 8.67e-19
C7313 VDD.n976 VSS 0.00281f
C7314 VDD.t93 VSS 0.00159f
C7315 VDD.n977 VSS 0.00354f
C7316 VDD.n978 VSS 7.59e-19
C7317 VDD.n979 VSS 0.00215f
C7318 VDD.n980 VSS 3.97e-19
C7319 VDD.n981 VSS 2.85e-19
C7320 VDD.n982 VSS 0.00154f
C7321 VDD.t202 VSS 0.00262f
C7322 VDD.n983 VSS 0.00271f
C7323 VDD.t94 VSS 0.0139f
C7324 VDD.n984 VSS 0.0119f
C7325 VDD.n985 VSS 7.81e-19
C7326 VDD.n986 VSS 0.00267f
C7327 VDD.n987 VSS 0.00307f
C7328 VDD.t201 VSS 0.00578f
C7329 VDD.t328 VSS 0.00578f
C7330 VDD.n988 VSS 0.00452f
C7331 VDD.n989 VSS 0.00109f
C7332 VDD.n990 VSS 0.00172f
C7333 VDD.n991 VSS 0.00308f
C7334 VDD.n992 VSS 0.00666f
C7335 VDD.n993 VSS 0.00109f
C7336 VDD.n994 VSS 0.00164f
C7337 VDD.n995 VSS 0.00308f
C7338 VDD.t723 VSS 5.72e-19
C7339 VDD.t460 VSS 7.62e-19
C7340 VDD.n996 VSS 0.0014f
C7341 VDD.t722 VSS 0.00578f
C7342 VDD.n997 VSS 0.0076f
C7343 VDD.n998 VSS 0.00111f
C7344 VDD.n999 VSS 0.00204f
C7345 VDD.n1000 VSS 0.00252f
C7346 VDD.n1001 VSS 0.00308f
C7347 VDD.t459 VSS 0.00578f
C7348 VDD.n1002 VSS 0.00603f
C7349 VDD.n1003 VSS 0.00109f
C7350 VDD.n1004 VSS 0.00132f
C7351 VDD.n1005 VSS 0.00308f
C7352 VDD.t585 VSS 0.00578f
C7353 VDD.n1006 VSS 0.00634f
C7354 VDD.n1007 VSS 0.00109f
C7355 VDD.n1008 VSS 0.00186f
C7356 VDD.n1009 VSS 0.00308f
C7357 VDD.t81 VSS 0.00578f
C7358 VDD.n1010 VSS 0.00528f
C7359 VDD.n1011 VSS 0.00109f
C7360 VDD.n1012 VSS 0.00186f
C7361 VDD.n1013 VSS 0.00308f
C7362 VDD.n1014 VSS 0.00905f
C7363 VDD.n1015 VSS 0.00109f
C7364 VDD.n1016 VSS 0.00186f
C7365 VDD.n1017 VSS 0.00308f
C7366 VDD.t369 VSS 0.00578f
C7367 VDD.n1018 VSS 0.00823f
C7368 VDD.n1019 VSS 0.00109f
C7369 VDD.n1020 VSS 0.0011f
C7370 VDD.n1021 VSS 0.00308f
C7371 VDD.t370 VSS 0.00217f
C7372 VDD.t200 VSS 9.67e-19
C7373 VDD.n1022 VSS 0.00349f
C7374 VDD.n1023 VSS 0.00457f
C7375 VDD.t199 VSS 0.00565f
C7376 VDD.n1024 VSS 0.00616f
C7377 VDD.n1025 VSS 0.00109f
C7378 VDD.n1026 VSS 0.00102f
C7379 VDD.n1027 VSS 0.00308f
C7380 VDD.t317 VSS 0.0054f
C7381 VDD.n1028 VSS 0.0059f
C7382 VDD.n1029 VSS 0.00109f
C7383 VDD.n1030 VSS 0.00186f
C7384 VDD.n1031 VSS 0.00308f
C7385 VDD.t271 VSS 0.00578f
C7386 VDD.n1032 VSS 0.00666f
C7387 VDD.n1033 VSS 0.00109f
C7388 VDD.n1034 VSS 0.00118f
C7389 VDD.n1035 VSS 0.00248f
C7390 VDD.n1036 VSS 0.00106f
C7391 VDD.n1037 VSS 0.00154f
C7392 VDD.n1038 VSS 2.85e-19
C7393 VDD.t371 VSS 0.00578f
C7394 VDD.n1039 VSS 0.00666f
C7395 VDD.n1040 VSS 0.00111f
C7396 VDD.n1041 VSS 0.00201f
C7397 VDD.t272 VSS 5.72e-19
C7398 VDD.t372 VSS 5.42e-19
C7399 VDD.n1042 VSS 0.00118f
C7400 VDD.n1043 VSS 0.0026f
C7401 VDD.n1044 VSS 2.25e-19
C7402 VDD.n1045 VSS 4.86e-19
C7403 VDD.n1046 VSS 4.35e-19
C7404 VDD.n1047 VSS 4.77e-19
C7405 VDD.n1048 VSS 3.36e-19
C7406 VDD.n1049 VSS 8.1e-19
C7407 VDD.n1050 VSS 0.0133f
C7408 VDD.n1051 VSS 0.00542f
C7409 VDD.n1052 VSS 0.0108f
C7410 VDD.n1053 VSS 0.0241f
C7411 VDD.n1054 VSS 0.0389f
C7412 VDD.n1055 VSS 0.388f
C7413 VDD.n1056 VSS 3.58f
C7414 VDD.n1057 VSS 0.0409f
C7415 VDD.n1058 VSS 0.0148f
C7416 VDD.n1059 VSS 0.00158f
C7417 VDD.n1060 VSS 5.66e-19
C7418 VDD.t47 VSS 8.49e-19
C7419 VDD.t499 VSS -2.71e-19
C7420 VDD.n1061 VSS 0.00391f
C7421 VDD.n1062 VSS 0.00409f
C7422 VDD.t498 VSS 0.00579f
C7423 VDD.n1063 VSS 0.00598f
C7424 VDD.n1064 VSS 0.00109f
C7425 VDD.n1065 VSS 9.92e-19
C7426 VDD.n1066 VSS 0.00258f
C7427 VDD.n1067 VSS 0.00124f
C7428 VDD.n1068 VSS 7.71e-19
C7429 VDD.n1069 VSS 9.31e-19
C7430 VDD.t365 VSS 0.00472f
C7431 VDD.t249 VSS 0.00579f
C7432 VDD.n1070 VSS 0.00529f
C7433 VDD.n1071 VSS 0.00111f
C7434 VDD.n1072 VSS 0.00202f
C7435 VDD.t366 VSS 6.03e-19
C7436 VDD.t250 VSS 6.03e-19
C7437 VDD.n1073 VSS 0.0013f
C7438 VDD.n1074 VSS 0.0027f
C7439 VDD.t346 VSS 0.00262f
C7440 VDD.n1075 VSS 0.0026f
C7441 VDD.n1076 VSS 0.00995f
C7442 VDD.n1077 VSS 0.0011f
C7443 VDD.n1078 VSS 0.00231f
C7444 VDD.n1079 VSS 0.00228f
C7445 VDD.n1080 VSS 0.00121f
C7446 VDD.n1081 VSS 5.41e-19
C7447 VDD.n1082 VSS 5.66e-19
C7448 VDD.n1083 VSS 0.00158f
C7449 VDD.n1084 VSS 0.00149f
C7450 VDD.n1085 VSS 8.1e-19
C7451 VDD.n1086 VSS 3.36e-19
C7452 VDD.n1087 VSS 4.35e-19
C7453 VDD.n1088 VSS 8.45e-19
C7454 VDD.n1089 VSS 3.35e-19
C7455 VDD.n1090 VSS 9.31e-19
C7456 VDD.t310 VSS 0.00579f
C7457 VDD.t345 VSS 0.00579f
C7458 VDD.n1091 VSS 0.00453f
C7459 VDD.n1092 VSS 0.00109f
C7460 VDD.n1093 VSS 1.72e-19
C7461 VDD.n1094 VSS 2.85e-19
C7462 VDD.n1095 VSS 0.00154f
C7463 VDD.n1096 VSS 0.00668f
C7464 VDD.n1097 VSS 0.00109f
C7465 VDD.n1098 VSS 0.00153f
C7466 VDD.n1099 VSS 0.0029f
C7467 VDD.t717 VSS 7.62e-19
C7468 VDD.t116 VSS 5.72e-19
C7469 VDD.n1100 VSS 0.0014f
C7470 VDD.t115 VSS 0.00579f
C7471 VDD.n1101 VSS 0.00762f
C7472 VDD.n1102 VSS 0.00111f
C7473 VDD.n1103 VSS 0.00204f
C7474 VDD.n1104 VSS 0.00252f
C7475 VDD.n1105 VSS 0.00308f
C7476 VDD.t716 VSS 0.00579f
C7477 VDD.n1106 VSS 0.00605f
C7478 VDD.n1107 VSS 0.00109f
C7479 VDD.n1108 VSS 0.00132f
C7480 VDD.n1109 VSS 0.00308f
C7481 VDD.t252 VSS 0.00579f
C7482 VDD.n1110 VSS 0.00636f
C7483 VDD.n1111 VSS 0.00109f
C7484 VDD.n1112 VSS 0.00186f
C7485 VDD.n1113 VSS 0.00308f
C7486 VDD.t395 VSS 0.00579f
C7487 VDD.n1114 VSS 0.00529f
C7488 VDD.n1115 VSS 0.00109f
C7489 VDD.n1116 VSS 0.00186f
C7490 VDD.n1117 VSS 0.00308f
C7491 VDD.n1118 VSS 0.00907f
C7492 VDD.n1119 VSS 0.00109f
C7493 VDD.n1120 VSS 0.00186f
C7494 VDD.n1121 VSS 0.00308f
C7495 VDD.t205 VSS 0.00579f
C7496 VDD.n1122 VSS 0.00825f
C7497 VDD.n1123 VSS 0.00109f
C7498 VDD.n1124 VSS 0.0011f
C7499 VDD.n1125 VSS 0.00308f
C7500 VDD.t348 VSS 9.67e-19
C7501 VDD.t206 VSS 0.00217f
C7502 VDD.n1126 VSS 0.00349f
C7503 VDD.n1127 VSS 0.00457f
C7504 VDD.t347 VSS 0.00567f
C7505 VDD.n1128 VSS 0.00617f
C7506 VDD.n1129 VSS 0.00109f
C7507 VDD.n1130 VSS 0.00102f
C7508 VDD.n1131 VSS 0.00308f
C7509 VDD.t97 VSS 0.0134f
C7510 VDD.t744 VSS 0.00542f
C7511 VDD.n1132 VSS 0.0068f
C7512 VDD.n1133 VSS 0.00103f
C7513 VDD.n1134 VSS 0.00176f
C7514 VDD.n1135 VSS 0.00291f
C7515 VDD.n1136 VSS 0.00154f
C7516 VDD.n1137 VSS 1.36e-19
C7517 VDD.t114 VSS 0.00149f
C7518 VDD.t767 VSS 6.37e-19
C7519 VDD.n1138 VSS 0.00279f
C7520 VDD.n1139 VSS 2.33e-19
C7521 VDD.n1140 VSS 6.77e-19
C7522 VDD.n1141 VSS 0.00141f
C7523 VDD.n1142 VSS 2.33e-19
C7524 VDD.n1143 VSS 0.00388f
C7525 VDD.n1144 VSS 5.31e-19
C7526 VDD.n1145 VSS 0.00105f
C7527 VDD.t769 VSS 6.29e-19
C7528 VDD.n1146 VSS 0.00315f
C7529 VDD.t96 VSS 0.00189f
C7530 VDD.n1147 VSS 0.00174f
C7531 VDD.n1148 VSS 2.32e-19
C7532 VDD.n1149 VSS 9.31e-19
C7533 VDD.n1150 VSS 1.72e-19
C7534 VDD.n1151 VSS 2.85e-19
C7535 VDD.n1152 VSS 0.00146f
C7536 VDD.n1153 VSS 0.00198f
C7537 VDD.t204 VSS 5.42e-19
C7538 VDD.t98 VSS 5.72e-19
C7539 VDD.n1154 VSS 0.00119f
C7540 VDD.n1155 VSS 0.00282f
C7541 VDD.n1156 VSS 0.00296f
C7542 VDD.t203 VSS 0.0107f
C7543 VDD.n1157 VSS 0.00756f
C7544 VDD.n1158 VSS 0.00191f
C7545 VDD.n1159 VSS 0.00177f
C7546 VDD.n1160 VSS 0.00308f
C7547 VDD.t394 VSS 0.00579f
C7548 VDD.n1161 VSS 0.00529f
C7549 VDD.n1162 VSS 0.00109f
C7550 VDD.n1163 VSS 0.00186f
C7551 VDD.n1164 VSS 0.00308f
C7552 VDD.t251 VSS 0.00579f
C7553 VDD.n1165 VSS 0.00579f
C7554 VDD.n1166 VSS 0.00109f
C7555 VDD.n1167 VSS 0.00151f
C7556 VDD.n1168 VSS 0.00308f
C7557 VDD.t216 VSS 0.00142f
C7558 VDD.t215 VSS 0.00579f
C7559 VDD.n1169 VSS 0.00857f
C7560 VDD.n1170 VSS 0.00111f
C7561 VDD.n1171 VSS 0.00203f
C7562 VDD.n1172 VSS 0.00312f
C7563 VDD.n1173 VSS 0.00308f
C7564 VDD.n1174 VSS 0.00907f
C7565 VDD.n1175 VSS 0.00109f
C7566 VDD.n1176 VSS 0.00118f
C7567 VDD.n1177 VSS 0.00308f
C7568 VDD.n1178 VSS 0.0028f
C7569 VDD.n1179 VSS 0.00106f
C7570 VDD.n1180 VSS 0.00138f
C7571 VDD.n1181 VSS 0.00109f
C7572 VDD.n1182 VSS 0.00882f
C7573 VDD.n1183 VSS 0.00109f
C7574 VDD.n1184 VSS 1.72e-19
C7575 VDD.n1185 VSS 2.85e-19
C7576 VDD.n1186 VSS 8.7e-19
C7577 VDD.n1187 VSS 3.01e-19
C7578 VDD.n1188 VSS 4.35e-19
C7579 VDD.n1189 VSS 5.41e-19
C7580 VDD.n1190 VSS 3.36e-19
C7581 VDD.n1191 VSS 0.00149f
C7582 VDD.n1192 VSS 8.1e-19
C7583 VDD.n1193 VSS 0.0148f
C7584 VDD.n1194 VSS 0.0148f
C7585 VDD.n1195 VSS 0.00149f
C7586 VDD.n1196 VSS 8.1e-19
C7587 VDD.n1197 VSS 5.41e-19
C7588 VDD.n1198 VSS 3.36e-19
C7589 VDD.n1199 VSS 3.35e-19
C7590 VDD.n1200 VSS 0.00112f
C7591 VDD.n1201 VSS 0.00102f
C7592 VDD.n1202 VSS 2.85e-19
C7593 VDD.n1203 VSS 1.32e-19
C7594 VDD.n1204 VSS 2.23e-19
C7595 VDD.n1205 VSS 5.1e-19
C7596 VDD.n1206 VSS 0.00419f
C7597 VDD.t675 VSS 0.00476f
C7598 VDD.n1207 VSS 4.81e-19
C7599 VDD.n1208 VSS 0.00108f
C7600 VDD.n1209 VSS 0.00584f
C7601 VDD.n1210 VSS 5.46e-19
C7602 VDD.n1211 VSS 1.72e-19
C7603 VDD.n1212 VSS 0.0107f
C7604 VDD.n1213 VSS 0.001f
C7605 VDD.n1214 VSS 0.00133f
C7606 VDD.n1215 VSS 0.011f
C7607 VDD.n1216 VSS 0.00103f
C7608 VDD.n1217 VSS 0.00129f
C7609 VDD.n1218 VSS 6.55e-19
C7610 VDD.n1219 VSS 1.21e-19
C7611 VDD.n1220 VSS 1.11e-19
C7612 VDD.n1221 VSS 1.11e-19
C7613 VDD.n1222 VSS 1.84e-19
C7614 VDD.n1223 VSS 1.84e-19
C7615 VDD.n1224 VSS 2.01e-19
C7616 VDD.n1225 VSS 1.68e-19
C7617 VDD.n1226 VSS 0.00298f
C7618 VDD.n1227 VSS 3.01e-19
C7619 VDD.n1228 VSS 2.85e-19
C7620 VDD.n1229 VSS 1.72e-19
C7621 VDD.n1230 VSS 6.07e-19
C7622 VDD.n1231 VSS 1.72e-19
C7623 VDD.n1232 VSS 3.04e-19
C7624 VDD.n1233 VSS 5.46e-19
C7625 VDD.n1234 VSS 0.00584f
C7626 VDD.n1235 VSS 0.00108f
C7627 VDD.n1236 VSS 0.00114f
C7628 VDD.t267 VSS 0.00191f
C7629 VDD.n1237 VSS 0.00222f
C7630 VDD.n1238 VSS 0.00108f
C7631 VDD.n1239 VSS 0.00381f
C7632 VDD.n1240 VSS 5.34e-19
C7633 VDD.n1241 VSS 3.04e-19
C7634 VDD.n1242 VSS 1.72e-19
C7635 VDD.n1243 VSS 2.85e-19
C7636 VDD.n1244 VSS 0.00151f
C7637 VDD.n1245 VSS 0.00129f
C7638 VDD.n1246 VSS 6.07e-19
C7639 VDD.n1247 VSS 6.07e-19
C7640 VDD.n1248 VSS 1.72e-19
C7641 VDD.n1249 VSS 4.57e-19
C7642 VDD.n1250 VSS 1.01e-19
C7643 VDD.t162 VSS 0.00476f
C7644 VDD.n1251 VSS 0.00292f
C7645 VDD.n1252 VSS 0.00108f
C7646 VDD.n1253 VSS 0.00362f
C7647 VDD.n1254 VSS 5.34e-19
C7648 VDD.n1255 VSS 3.04e-19
C7649 VDD.n1256 VSS 1.72e-19
C7650 VDD.n1257 VSS 2.85e-19
C7651 VDD.n1258 VSS 0.00151f
C7652 VDD.n1259 VSS 0.00129f
C7653 VDD.n1260 VSS 6.07e-19
C7654 VDD.n1261 VSS 6.07e-19
C7655 VDD.n1262 VSS 1.72e-19
C7656 VDD.n1263 VSS 4.57e-19
C7657 VDD.n1264 VSS 1.01e-19
C7658 VDD.t561 VSS 0.00476f
C7659 VDD.n1265 VSS 0.00489f
C7660 VDD.n1266 VSS 0.00108f
C7661 VDD.n1267 VSS 0.00292f
C7662 VDD.n1268 VSS 5.34e-19
C7663 VDD.n1269 VSS 3.04e-19
C7664 VDD.n1270 VSS 1.72e-19
C7665 VDD.n1271 VSS 2.85e-19
C7666 VDD.n1272 VSS 0.00151f
C7667 VDD.n1273 VSS 0.00129f
C7668 VDD.n1274 VSS 6.07e-19
C7669 VDD.n1275 VSS 6.07e-19
C7670 VDD.n1276 VSS 1.72e-19
C7671 VDD.n1277 VSS 4.57e-19
C7672 VDD.n1278 VSS 1.01e-19
C7673 VDD.n1279 VSS 0.00483f
C7674 VDD.n1280 VSS 0.00108f
C7675 VDD.n1281 VSS 0.00572f
C7676 VDD.n1282 VSS 5.34e-19
C7677 VDD.n1283 VSS 3.04e-19
C7678 VDD.n1284 VSS 1.72e-19
C7679 VDD.n1285 VSS 2.85e-19
C7680 VDD.n1286 VSS 0.00151f
C7681 VDD.n1287 VSS 0.00129f
C7682 VDD.n1288 VSS 6.07e-19
C7683 VDD.n1289 VSS 6.07e-19
C7684 VDD.n1290 VSS 1.72e-19
C7685 VDD.n1291 VSS 4.57e-19
C7686 VDD.n1292 VSS 1.01e-19
C7687 VDD.t618 VSS 0.00476f
C7688 VDD.n1293 VSS 0.00356f
C7689 VDD.n1294 VSS 0.00108f
C7690 VDD.n1295 VSS 0.00102f
C7691 VDD.n1296 VSS 5.34e-19
C7692 VDD.n1297 VSS 3.04e-19
C7693 VDD.n1298 VSS 1.72e-19
C7694 VDD.n1299 VSS 2.85e-19
C7695 VDD.n1300 VSS 0.00151f
C7696 VDD.n1301 VSS 0.00129f
C7697 VDD.n1302 VSS 6.07e-19
C7698 VDD.t514 VSS 5.42e-19
C7699 VDD.t218 VSS 4.25e-19
C7700 VDD.n1303 VSS 0.00111f
C7701 VDD.n1304 VSS 0.00224f
C7702 VDD.n1305 VSS 1.62e-19
C7703 VDD.n1306 VSS 1.72e-19
C7704 VDD.n1307 VSS 4.57e-19
C7705 VDD.n1308 VSS 1.01e-19
C7706 VDD.t513 VSS 0.00476f
C7707 VDD.n1309 VSS 0.00381f
C7708 VDD.n1310 VSS 0.00108f
C7709 VDD.n1311 VSS 0.00229f
C7710 VDD.n1312 VSS 5.34e-19
C7711 VDD.n1313 VSS 3.04e-19
C7712 VDD.n1314 VSS 1.72e-19
C7713 VDD.n1315 VSS 2.85e-19
C7714 VDD.n1316 VSS 0.00151f
C7715 VDD.n1317 VSS 0.00129f
C7716 VDD.n1318 VSS 4.66e-19
C7717 VDD.n1319 VSS 6.07e-19
C7718 VDD.n1320 VSS 1.72e-19
C7719 VDD.n1321 VSS 4.57e-19
C7720 VDD.n1322 VSS 1.01e-19
C7721 VDD.t217 VSS 0.00476f
C7722 VDD.n1323 VSS 0.00489f
C7723 VDD.n1324 VSS 0.00108f
C7724 VDD.n1325 VSS 0.00203f
C7725 VDD.n1326 VSS 5.34e-19
C7726 VDD.n1327 VSS 3.04e-19
C7727 VDD.n1328 VSS 1.72e-19
C7728 VDD.n1329 VSS 2.85e-19
C7729 VDD.n1330 VSS 0.00151f
C7730 VDD.n1331 VSS 0.00129f
C7731 VDD.n1332 VSS 6.07e-19
C7732 VDD.n1333 VSS 0.0116f
C7733 VDD.n1334 VSS 0.00108f
C7734 VDD.n1335 VSS 0.00154f
C7735 VDD.n1336 VSS 8.47e-19
C7736 VDD.n1337 VSS 1.72e-19
C7737 VDD.n1338 VSS 5.46e-19
C7738 VDD.n1339 VSS 1.01e-19
C7739 VDD.n1340 VSS 0.00584f
C7740 VDD.n1341 VSS 0.00108f
C7741 VDD.n1342 VSS 0.00572f
C7742 VDD.n1343 VSS 5.34e-19
C7743 VDD.n1344 VSS 3.04e-19
C7744 VDD.n1345 VSS 1.72e-19
C7745 VDD.n1346 VSS 2.85e-19
C7746 VDD.n1347 VSS 7.71e-19
C7747 VDD.n1348 VSS 0.0109f
C7748 VDD.n1349 VSS 0.0117f
C7749 VDD.n1350 VSS 0.00109f
C7750 VDD.n1351 VSS 0.00157f
C7751 VDD.n1352 VSS 0.0117f
C7752 VDD.n1353 VSS 0.00109f
C7753 VDD.n1354 VSS 0.00157f
C7754 VDD.n1355 VSS 0.0117f
C7755 VDD.n1356 VSS 0.00109f
C7756 VDD.n1357 VSS 0.00157f
C7757 VDD.n1358 VSS 0.0117f
C7758 VDD.n1359 VSS 0.00109f
C7759 VDD.n1360 VSS 0.00157f
C7760 VDD.n1361 VSS 0.0113f
C7761 VDD.n1362 VSS 0.00106f
C7762 VDD.n1363 VSS 0.00151f
C7763 VDD.n1364 VSS 8.67e-19
C7764 VDD.n1365 VSS 1.72e-19
C7765 VDD.n1366 VSS 5.46e-19
C7766 VDD.n1367 VSS 1.01e-19
C7767 VDD.n1368 VSS 0.00584f
C7768 VDD.n1369 VSS 0.00108f
C7769 VDD.n1370 VSS 0.00546f
C7770 VDD.n1371 VSS 5.1e-19
C7771 VDD.n1372 VSS 2.23e-19
C7772 VDD.n1373 VSS 6.48e-19
C7773 VDD.n1374 VSS 1.72e-19
C7774 VDD.n1375 VSS 2.85e-19
C7775 VDD.n1376 VSS 0.00136f
C7776 VDD.n1377 VSS 0.00127f
C7777 VDD.n1378 VSS 1.84e-19
C7778 VDD.n1379 VSS 2.68e-19
C7779 VDD.n1380 VSS 1.17e-19
C7780 VDD.n1381 VSS 6.48e-19
C7781 VDD.n1382 VSS 1.72e-19
C7782 VDD.n1383 VSS 4.81e-19
C7783 VDD.n1384 VSS 1.01e-19
C7784 VDD.n1385 VSS 0.00514f
C7785 VDD.n1386 VSS 0.00108f
C7786 VDD.t382 VSS 0.00476f
C7787 VDD.n1387 VSS 0.00152f
C7788 VDD.n1388 VSS 5.1e-19
C7789 VDD.n1389 VSS 1.21e-19
C7790 VDD.n1390 VSS 1.11e-19
C7791 VDD.n1391 VSS 1.62e-19
C7792 VDD.n1392 VSS 7.08e-20
C7793 VDD.t383 VSS 4.25e-19
C7794 VDD.t511 VSS 5.42e-19
C7795 VDD.n1393 VSS 0.00111f
C7796 VDD.n1394 VSS 0.00223f
C7797 VDD.n1395 VSS 4.05e-19
C7798 VDD.n1396 VSS 2.85e-19
C7799 VDD.n1397 VSS 0.00144f
C7800 VDD.n1398 VSS 0.00136f
C7801 VDD.n1399 VSS 2.43e-19
C7802 VDD.n1400 VSS 1.72e-19
C7803 VDD.n1401 VSS 4.81e-19
C7804 VDD.n1402 VSS 1.01e-19
C7805 VDD.n1403 VSS 0.00432f
C7806 VDD.n1404 VSS 0.00108f
C7807 VDD.t510 VSS 0.00476f
C7808 VDD.n1405 VSS 0.00178f
C7809 VDD.n1406 VSS 5.1e-19
C7810 VDD.n1407 VSS 2.23e-19
C7811 VDD.n1408 VSS 6.48e-19
C7812 VDD.n1409 VSS 1.72e-19
C7813 VDD.n1410 VSS 2.85e-19
C7814 VDD.n1411 VSS 9.88e-19
C7815 VDD.n1412 VSS 9.71e-19
C7816 VDD.n1413 VSS 4.35e-19
C7817 VDD.n1414 VSS 3.36e-19
C7818 VDD.n1415 VSS 8.1e-19
C7819 VDD.n1416 VSS 0.0148f
C7820 VDD.n1417 VSS 0.0148f
C7821 VDD.n1418 VSS 0.0468f
C7822 VDD.n1419 VSS 0.0601f
C7823 VDD.n1420 VSS 0.00158f
C7824 VDD.n1421 VSS 0.00149f
C7825 VDD.n1422 VSS 8.1e-19
C7826 VDD.n1423 VSS 0.00158f
C7827 VDD.n1424 VSS 0.00144f
C7828 VDD.n1425 VSS 0.00148f
C7829 VDD.n1426 VSS 8.1e-19
C7830 VDD.n1427 VSS 0.00158f
C7831 VDD.n1428 VSS 0.00149f
C7832 VDD.n1429 VSS 6.05e-19
C7833 VDD.n1430 VSS 0.00104f
C7834 VDD.n1431 VSS 3.01e-19
C7835 VDD.n1432 VSS 8.97e-19
C7836 VDD.n1433 VSS 1.72e-19
C7837 VDD.n1434 VSS 5.4e-19
C7838 VDD.n1435 VSS 1.01e-19
C7839 VDD.n1436 VSS 0.004f
C7840 VDD.n1437 VSS 0.00108f
C7841 VDD.n1438 VSS 5.4e-19
C7842 VDD.n1439 VSS 1.01e-19
C7843 VDD.t406 VSS 7.73e-19
C7844 VDD.t320 VSS 2.51e-19
C7845 VDD.n1440 VSS 0.00395f
C7846 VDD.n1441 VSS 7.49e-19
C7847 VDD.n1442 VSS 5.97e-19
C7848 VDD.n1443 VSS 1.42e-19
C7849 VDD.n1444 VSS 0.0023f
C7850 VDD.n1445 VSS 3.04e-20
C7851 VDD.n1446 VSS 7.49e-19
C7852 VDD.n1447 VSS 9.88e-19
C7853 VDD.n1448 VSS 2.68e-19
C7854 VDD.n1449 VSS 2.68e-19
C7855 VDD.n1450 VSS 3.35e-20
C7856 VDD.n1451 VSS 0.00127f
C7857 VDD.n1452 VSS 7.49e-19
C7858 VDD.n1453 VSS 7.49e-19
C7859 VDD.n1454 VSS 1.72e-19
C7860 VDD.n1455 VSS 5.4e-19
C7861 VDD.n1456 VSS 1.01e-19
C7862 VDD.t405 VSS 0.00476f
C7863 VDD.n1457 VSS 0.0047f
C7864 VDD.n1458 VSS 0.00108f
C7865 VDD.n1459 VSS 0.00184f
C7866 VDD.n1460 VSS 4.51e-19
C7867 VDD.n1461 VSS 2.02e-20
C7868 VDD.n1462 VSS 1.72e-19
C7869 VDD.n1463 VSS 2.85e-19
C7870 VDD.n1464 VSS 0.00107f
C7871 VDD.n1465 VSS 0.00106f
C7872 VDD.n1466 VSS 5.79e-19
C7873 VDD.n1467 VSS 5.28e-19
C7874 VDD.n1468 VSS 0.00158f
C7875 VDD.n1469 VSS 0.00149f
C7876 VDD.n1470 VSS 8.1e-19
C7877 VDD.n1471 VSS 3.36e-19
C7878 VDD.n1472 VSS 4.35e-19
C7879 VDD.n1473 VSS 2.01e-19
C7880 VDD.n1474 VSS 1.72e-19
C7881 VDD.n1475 VSS 2.02e-20
C7882 VDD.n1476 VSS 4.51e-19
C7883 VDD.n1477 VSS 0.00203f
C7884 VDD.t319 VSS 0.00279f
C7885 VDD.n1478 VSS 0.00292f
C7886 VDD.n1479 VSS 0.00108f
C7887 VDD.n1480 VSS 0.00584f
C7888 VDD.n1481 VSS 5.46e-19
C7889 VDD.n1482 VSS 2.02e-20
C7890 VDD.n1483 VSS 1.72e-19
C7891 VDD.n1484 VSS 2.85e-19
C7892 VDD.n1485 VSS 0.00295f
C7893 VDD.n1486 VSS 1.68e-19
C7894 VDD.n1487 VSS 1.68e-19
C7895 VDD.n1488 VSS 2.18e-19
C7896 VDD.n1489 VSS 6.48e-19
C7897 VDD.n1490 VSS 1.72e-19
C7898 VDD.n1491 VSS 1.01e-19
C7899 VDD.n1492 VSS 0.00273f
C7900 VDD.n1493 VSS 0.00108f
C7901 VDD.n1494 VSS 4.81e-19
C7902 VDD.n1495 VSS 1.01e-19
C7903 VDD.n1496 VSS 6.48e-19
C7904 VDD.n1497 VSS 1.72e-19
C7905 VDD.t636 VSS 7.73e-19
C7906 VDD.t208 VSS 2.51e-19
C7907 VDD.n1498 VSS 0.00395f
C7908 VDD.n1499 VSS 6.27e-19
C7909 VDD.n1500 VSS 0.00221f
C7910 VDD.n1501 VSS 0.00144f
C7911 VDD.n1502 VSS 9.88e-19
C7912 VDD.n1503 VSS 2.85e-19
C7913 VDD.n1504 VSS 1.32e-19
C7914 VDD.n1505 VSS 2.23e-19
C7915 VDD.n1506 VSS 5.1e-19
C7916 VDD.n1507 VSS 0.00419f
C7917 VDD.t207 VSS 0.00476f
C7918 VDD.n1508 VSS 4.81e-19
C7919 VDD.n1509 VSS 0.00108f
C7920 VDD.n1510 VSS 0.00978f
C7921 VDD.n1511 VSS 8.64e-19
C7922 VDD.n1512 VSS 1.52e-19
C7923 VDD.n1513 VSS 0.0149f
C7924 VDD.n1514 VSS 0.00135f
C7925 VDD.n1515 VSS 0.00165f
C7926 VDD.n1516 VSS 0.00122f
C7927 VDD.n1517 VSS 1.01e-19
C7928 VDD.n1518 VSS 1.32e-19
C7929 VDD.n1519 VSS 1.11e-19
C7930 VDD.n1520 VSS 1.84e-19
C7931 VDD.n1521 VSS 2.85e-19
C7932 VDD.n1522 VSS 3.68e-19
C7933 VDD.n1523 VSS 5.03e-19
C7934 VDD.n1524 VSS 3.36e-19
C7935 VDD.n1525 VSS 8.1e-19
C7936 VDD.n1526 VSS 0.00158f
C7937 VDD.n1527 VSS 0.00149f
C7938 VDD.n1528 VSS 8.1e-19
C7939 VDD.n1529 VSS 0.00158f
C7940 VDD.n1530 VSS 0.00149f
C7941 VDD.n1531 VSS 5.54e-19
C7942 VDD.n1532 VSS 5.54e-19
C7943 VDD.t191 VSS 6.03e-19
C7944 VDD.t296 VSS 6.03e-19
C7945 VDD.n1533 VSS 0.0013f
C7946 VDD.n1534 VSS 0.00882f
C7947 VDD.n1535 VSS 5.77e-19
C7948 VDD.n1536 VSS 0.00129f
C7949 VDD.n1537 VSS 0.00898f
C7950 VDD.n1538 VSS 2.54e-19
C7951 VDD.n1539 VSS 3.35e-20
C7952 VDD.n1540 VSS 2.7e-19
C7953 VDD.n1541 VSS 0.00213f
C7954 VDD.n1542 VSS 3.74e-19
C7955 VDD.n1543 VSS 4.68e-20
C7956 VDD.n1544 VSS 5.4e-19
C7957 VDD.t720 VSS 0.00466f
C7958 VDD.n1545 VSS 0.00195f
C7959 VDD.n1546 VSS 0.00693f
C7960 VDD.n1547 VSS 6.53e-19
C7961 VDD.n1548 VSS 3.74e-19
C7962 VDD.n1549 VSS 0.00166f
C7963 VDD.n1550 VSS 3.97e-19
C7964 VDD.n1551 VSS 6.6e-19
C7965 VDD.n1552 VSS 4.13e-19
C7966 VDD.n1553 VSS 6.93e-19
C7967 VDD.n1554 VSS 3.36e-19
C7968 VDD.n1555 VSS 4.4e-19
C7969 VDD.n1556 VSS 7.11e-19
C7970 VDD.n1557 VSS 0.00802f
C7971 VDD.t721 VSS 9.16e-19
C7972 VDD.t719 VSS -5.07e-19
C7973 VDD.n1558 VSS 0.00359f
C7974 VDD.n1559 VSS 0.00203f
C7975 VDD.t718 VSS 0.00579f
C7976 VDD.n1560 VSS 0.00611f
C7977 VDD.n1561 VSS 9.85e-19
C7978 VDD.n1562 VSS 0.00187f
C7979 VDD.n1563 VSS 0.00171f
C7980 VDD.n1564 VSS 0.00926f
C7981 VDD.n1565 VSS 0.00109f
C7982 VDD.n1566 VSS 0.00179f
C7983 VDD.n1567 VSS 0.00231f
C7984 VDD.n1568 VSS 0.00154f
C7985 VDD.t714 VSS 0.00579f
C7986 VDD.n1569 VSS 0.00838f
C7987 VDD.n1570 VSS 0.00109f
C7988 VDD.n1571 VSS 0.00186f
C7989 VDD.n1572 VSS 0.00231f
C7990 VDD.t715 VSS 8.49e-19
C7991 VDD.t151 VSS -2.71e-19
C7992 VDD.n1573 VSS 0.00391f
C7993 VDD.n1574 VSS 0.00413f
C7994 VDD.t150 VSS 0.00579f
C7995 VDD.n1575 VSS 0.00598f
C7996 VDD.n1576 VSS 0.00109f
C7997 VDD.n1577 VSS 9.92e-19
C7998 VDD.n1578 VSS 0.00308f
C7999 VDD.n1579 VSS 0.00109f
C8000 VDD.n1580 VSS 0.00168f
C8001 VDD.n1581 VSS 0.00231f
C8002 VDD.n1582 VSS 2.18e-19
C8003 VDD.n1583 VSS 6.55e-19
C8004 VDD.n1584 VSS 4.52e-19
C8005 VDD.n1585 VSS 3.36e-19
C8006 VDD.n1586 VSS 4.35e-19
C8007 VDD.n1587 VSS 9.31e-19
C8008 VDD.n1588 VSS 5.53e-19
C8009 VDD.n1589 VSS 2.85e-19
C8010 VDD.n1590 VSS 2.85e-19
C8011 VDD.n1591 VSS 1.72e-19
C8012 VDD.n1592 VSS 0.00109f
C8013 VDD.t190 VSS 0.00472f
C8014 VDD.t295 VSS 0.00579f
C8015 VDD.n1593 VSS 0.00529f
C8016 VDD.n1594 VSS 0.00111f
C8017 VDD.n1595 VSS 0.00185f
C8018 VDD.n1596 VSS 0.0027f
C8019 VDD.n1597 VSS 0.0026f
C8020 VDD.n1598 VSS 0.00154f
C8021 VDD.n1599 VSS 6.17e-19
C8022 VDD.n1600 VSS 0.00907f
C8023 VDD.n1601 VSS 0.00109f
C8024 VDD.n1602 VSS 1.72e-19
C8025 VDD.n1603 VSS 2.85e-19
C8026 VDD.n1604 VSS 5.67e-19
C8027 VDD.n1605 VSS 3.01e-19
C8028 VDD.t77 VSS 0.00142f
C8029 VDD.t76 VSS 0.00579f
C8030 VDD.n1606 VSS 0.00857f
C8031 VDD.n1607 VSS 0.00111f
C8032 VDD.n1608 VSS 0.00198f
C8033 VDD.n1609 VSS 0.00312f
C8034 VDD.n1610 VSS 0.00256f
C8035 VDD.n1611 VSS 0.00124f
C8036 VDD.n1612 VSS 4.35e-19
C8037 VDD.n1613 VSS 3.36e-19
C8038 VDD.n1614 VSS 8.1e-19
C8039 VDD.n1615 VSS 0.0108f
C8040 VDD.n1616 VSS 0.0133f
C8041 VDD.n1617 VSS 0.00542f
C8042 VDD.n1618 VSS 0.0163f
C8043 VDD.n1619 VSS 0.101f
C8044 VDD.n1620 VSS 0.101f
C8045 VDD.n1621 VSS 0.0296f
C8046 VDD.n1622 VSS 0.0261f
C8047 VDD.n1623 VSS 0.0261f
C8048 VDD.n1624 VSS 0.0296f
C8049 VDD.n1625 VSS 0.0867f
C8050 VDD.n1626 VSS 0.0867f
C8051 VDD.n1627 VSS 0.00149f
C8052 VDD.n1628 VSS 0.00144f
C8053 VDD.n1629 VSS 0.00157f
C8054 VDD.n1630 VSS 8.1e-19
C8055 VDD.n1631 VSS 0.0296f
C8056 VDD.n1632 VSS 0.0217f
C8057 VDD.n1633 VSS 0.0217f
C8058 VDD.n1634 VSS 0.00158f
C8059 VDD.n1635 VSS 6.3e-19
C8060 VDD.n1636 VSS 6.48e-19
C8061 VDD.n1637 VSS 1.72e-19
C8062 VDD.n1638 VSS 4.81e-19
C8063 VDD.n1639 VSS 1.01e-19
C8064 VDD.n1640 VSS 0.00406f
C8065 VDD.n1641 VSS 8.89e-19
C8066 VDD.t497 VSS 6.99e-19
C8067 VDD.n1642 VSS 0.00495f
C8068 VDD.n1643 VSS 5.1e-19
C8069 VDD.n1644 VSS 2.23e-19
C8070 VDD.n1645 VSS 6.48e-19
C8071 VDD.n1646 VSS 1.72e-19
C8072 VDD.n1647 VSS 2.85e-19
C8073 VDD.n1648 VSS 0.00136f
C8074 VDD.n1649 VSS 0.00144f
C8075 VDD.n1650 VSS 6.48e-19
C8076 VDD.n1651 VSS 1.72e-19
C8077 VDD.n1652 VSS 4.81e-19
C8078 VDD.n1653 VSS 1.01e-19
C8079 VDD.n1654 VSS 0.00514f
C8080 VDD.n1655 VSS 0.00108f
C8081 VDD.n1656 VSS 0.00546f
C8082 VDD.n1657 VSS 5.1e-19
C8083 VDD.n1658 VSS 2.23e-19
C8084 VDD.n1659 VSS 6.48e-19
C8085 VDD.n1660 VSS 1.72e-19
C8086 VDD.n1661 VSS 2.85e-19
C8087 VDD.n1662 VSS 9.55e-19
C8088 VDD.n1663 VSS 9.71e-19
C8089 VDD.n1664 VSS 0.00136f
C8090 VDD.n1665 VSS 6.27e-19
C8091 VDD.n1666 VSS 1.72e-19
C8092 VDD.n1667 VSS 4.81e-19
C8093 VDD.n1668 VSS 1.01e-19
C8094 VDD.n1669 VSS 0.00343f
C8095 VDD.n1670 VSS 0.00108f
C8096 VDD.t635 VSS 0.00476f
C8097 VDD.n1671 VSS 0.00311f
C8098 VDD.n1672 VSS 5.1e-19
C8099 VDD.n1673 VSS 2.23e-19
C8100 VDD.n1674 VSS 6.48e-19
C8101 VDD.n1675 VSS 1.72e-19
C8102 VDD.n1676 VSS 2.85e-19
C8103 VDD.n1677 VSS 0.00141f
C8104 VDD.n1678 VSS 0.00126f
C8105 VDD.n1679 VSS 1.34e-19
C8106 VDD.n1680 VSS 2.51e-19
C8107 VDD.n1681 VSS 6.48e-19
C8108 VDD.n1682 VSS 1.72e-19
C8109 VDD.n1683 VSS 4.81e-19
C8110 VDD.n1684 VSS 1.01e-19
C8111 VDD.n1685 VSS 0.00514f
C8112 VDD.n1686 VSS 0.00108f
C8113 VDD.t562 VSS 0.00476f
C8114 VDD.n1687 VSS 0.00241f
C8115 VDD.n1688 VSS 5.1e-19
C8116 VDD.n1689 VSS 1.32e-19
C8117 VDD.n1690 VSS 5.87e-19
C8118 VDD.n1691 VSS 8.1e-20
C8119 VDD.n1692 VSS 1.52e-19
C8120 VDD.n1693 VSS 1.11e-19
C8121 VDD.n1694 VSS 1.84e-19
C8122 VDD.n1695 VSS 3.18e-19
C8123 VDD.n1696 VSS 4.02e-19
C8124 VDD.n1697 VSS 4.77e-19
C8125 VDD.n1698 VSS 3.36e-19
C8126 VDD.n1699 VSS 0.00149f
C8127 VDD.n1700 VSS 8.1e-19
C8128 VDD.n1701 VSS 0.0296f
C8129 VDD.n1702 VSS 0.0424f
C8130 VDD.n1703 VSS 0.0424f
C8131 VDD.n1704 VSS 0.0241f
C8132 VDD.n1705 VSS 0.0148f
C8133 VDD.n1706 VSS 0.0148f
C8134 VDD.n1707 VSS 0.0241f
C8135 VDD.n1708 VSS 8.1e-19
C8136 VDD.n1709 VSS 3.36e-19
C8137 VDD.n1710 VSS 4.35e-19
C8138 VDD.t80 VSS 0.00578f
C8139 VDD.n1711 VSS 0.00528f
C8140 VDD.n1712 VSS 0.00109f
C8141 VDD.n1713 VSS 0.00186f
C8142 VDD.n1714 VSS 0.00169f
C8143 VDD.t582 VSS 0.00578f
C8144 VDD.n1715 VSS 0.00578f
C8145 VDD.n1716 VSS 0.00109f
C8146 VDD.n1717 VSS 0.00151f
C8147 VDD.n1718 VSS 0.00308f
C8148 VDD.t67 VSS 0.00142f
C8149 VDD.t66 VSS 0.00578f
C8150 VDD.n1719 VSS 0.00854f
C8151 VDD.n1720 VSS 0.00111f
C8152 VDD.n1721 VSS 0.00203f
C8153 VDD.n1722 VSS 0.00312f
C8154 VDD.n1723 VSS 0.00231f
C8155 VDD.n1724 VSS 0.00154f
C8156 VDD.n1725 VSS 0.00905f
C8157 VDD.n1726 VSS 0.00109f
C8158 VDD.n1727 VSS 0.00118f
C8159 VDD.n1728 VSS 0.00231f
C8160 VDD.t584 VSS 6.03e-19
C8161 VDD.t617 VSS 6.03e-19
C8162 VDD.n1729 VSS 0.0013f
C8163 VDD.t583 VSS 0.00578f
C8164 VDD.n1730 VSS 0.00528f
C8165 VDD.n1731 VSS 0.00111f
C8166 VDD.n1732 VSS 0.00202f
C8167 VDD.n1733 VSS 0.0027f
C8168 VDD.n1734 VSS 0.00308f
C8169 VDD.n1735 VSS 0.00183f
C8170 VDD.n1736 VSS 0.00151f
C8171 VDD.n1737 VSS 0.00109f
C8172 VDD.n1738 VSS 0.00773f
C8173 VDD.n1739 VSS 0.00109f
C8174 VDD.n1740 VSS 0.0018f
C8175 VDD.n1741 VSS 0.00231f
C8176 VDD.t644 VSS -2.71e-19
C8177 VDD.t472 VSS 8.49e-19
C8178 VDD.n1742 VSS 0.00391f
C8179 VDD.n1743 VSS 0.00413f
C8180 VDD.t643 VSS 0.00578f
C8181 VDD.n1744 VSS 0.00597f
C8182 VDD.n1745 VSS 0.00109f
C8183 VDD.n1746 VSS 9.92e-19
C8184 VDD.n1747 VSS 0.00308f
C8185 VDD.t471 VSS 0.00578f
C8186 VDD.n1748 VSS 0.00835f
C8187 VDD.n1749 VSS 0.00109f
C8188 VDD.n1750 VSS 0.00174f
C8189 VDD.n1751 VSS 0.00245f
C8190 VDD.n1752 VSS 9.88e-19
C8191 VDD.n1753 VSS 0.00154f
C8192 VDD.t469 VSS 0.00955f
C8193 VDD.n1754 VSS 0.00923f
C8194 VDD.n1755 VSS 6.76e-19
C8195 VDD.n1756 VSS 8.61e-19
C8196 VDD.n1757 VSS 1.72e-19
C8197 VDD.n1758 VSS 2.85e-19
C8198 VDD.n1759 VSS 9.31e-19
C8199 VDD.n1760 VSS 5.53e-19
C8200 VDD.n1761 VSS 4.35e-19
C8201 VDD.n1762 VSS 4.52e-19
C8202 VDD.n1763 VSS 3.36e-19
C8203 VDD.n1764 VSS 0.00149f
C8204 VDD.n1765 VSS 8.1e-19
C8205 VDD.n1766 VSS 0.0148f
C8206 VDD.n1767 VSS 0.0148f
C8207 VDD.n1768 VSS 0.0739f
C8208 VDD.n1769 VSS 0.0709f
C8209 VDD.n1770 VSS 0.0064f
C8210 VDD.n1771 VSS 0.0138f
C8211 VDD.n1772 VSS 0.00158f
C8212 VDD.n1773 VSS 0.00149f
C8213 VDD.n1774 VSS 5.28e-19
C8214 VDD.t470 VSS -5.07e-19
C8215 VDD.t149 VSS 9.16e-19
C8216 VDD.n1775 VSS 0.00359f
C8217 VDD.n1776 VSS 0.00204f
C8218 VDD.n1777 VSS 0.00181f
C8219 VDD.n1778 VSS 0.00253f
C8220 VDD.n1779 VSS 0.00127f
C8221 VDD.n1780 VSS 2.51e-19
C8222 VDD.t381 VSS 5.72e-19
C8223 VDD.t468 VSS 7.62e-19
C8224 VDD.n1781 VSS 0.0014f
C8225 VDD.t380 VSS 0.00578f
C8226 VDD.n1782 VSS 0.0076f
C8227 VDD.n1783 VSS 0.00111f
C8228 VDD.n1784 VSS 0.00204f
C8229 VDD.n1785 VSS 0.00252f
C8230 VDD.t578 VSS 5.72e-19
C8231 VDD.t364 VSS 5.42e-19
C8232 VDD.n1786 VSS 0.00119f
C8233 VDD.t363 VSS 0.00578f
C8234 VDD.n1787 VSS 0.00666f
C8235 VDD.n1788 VSS 0.00111f
C8236 VDD.n1789 VSS 0.00204f
C8237 VDD.n1790 VSS 0.00278f
C8238 VDD.t75 VSS 0.00142f
C8239 VDD.t74 VSS 0.00578f
C8240 VDD.n1791 VSS 0.00854f
C8241 VDD.n1792 VSS 0.00111f
C8242 VDD.n1793 VSS 0.00203f
C8243 VDD.n1794 VSS 0.00312f
C8244 VDD.t265 VSS 6.03e-19
C8245 VDD.t450 VSS 6.03e-19
C8246 VDD.n1795 VSS 0.0013f
C8247 VDD.n1796 VSS 0.0027f
C8248 VDD.t264 VSS 0.00578f
C8249 VDD.n1797 VSS 0.00202f
C8250 VDD.n1798 VSS 0.00111f
C8251 VDD.n1799 VSS 0.00528f
C8252 VDD.t449 VSS 0.00578f
C8253 VDD.t234 VSS -5.07e-19
C8254 VDD.t140 VSS 9.16e-19
C8255 VDD.n1800 VSS 0.00359f
C8256 VDD.n1801 VSS 0.00204f
C8257 VDD.n1802 VSS 0.00183f
C8258 VDD.n1803 VSS 0.00276f
C8259 VDD.n1804 VSS 0.00154f
C8260 VDD.n1805 VSS 8.58e-19
C8261 VDD.t233 VSS 0.00955f
C8262 VDD.n1806 VSS 0.00923f
C8263 VDD.n1807 VSS 6.76e-19
C8264 VDD.n1808 VSS 1.72e-19
C8265 VDD.n1809 VSS 2.85e-19
C8266 VDD.n1810 VSS 9.31e-19
C8267 VDD.n1811 VSS 6.37e-19
C8268 VDD.n1812 VSS 6.93e-19
C8269 VDD.n1813 VSS 0.00158f
C8270 VDD.n1814 VSS 0.0148f
C8271 VDD.n1815 VSS 0.00158f
C8272 VDD.n1816 VSS 0.00149f
C8273 VDD.n1817 VSS 4.64e-19
C8274 VDD.n1818 VSS 0.00154f
C8275 VDD.t756 VSS 8.67e-19
C8276 VDD.n1819 VSS 0.00281f
C8277 VDD.t138 VSS 0.0016f
C8278 VDD.n1820 VSS 0.00355f
C8279 VDD.n1821 VSS 7.59e-19
C8280 VDD.n1822 VSS 0.00215f
C8281 VDD.n1823 VSS 3.97e-19
C8282 VDD.n1824 VSS 2.85e-19
C8283 VDD.n1825 VSS 0.00116f
C8284 VDD.n1826 VSS 0.00147f
C8285 VDD.t696 VSS 0.00578f
C8286 VDD.t16 VSS 0.00578f
C8287 VDD.n1827 VSS 0.00452f
C8288 VDD.n1828 VSS 0.00109f
C8289 VDD.n1829 VSS 0.00172f
C8290 VDD.n1830 VSS 0.00245f
C8291 VDD.n1831 VSS 0.00154f
C8292 VDD.t697 VSS 0.00262f
C8293 VDD.n1832 VSS 0.00271f
C8294 VDD.t139 VSS 0.0139f
C8295 VDD.n1833 VSS 0.0119f
C8296 VDD.n1834 VSS 7.6e-19
C8297 VDD.n1835 VSS 0.00267f
C8298 VDD.n1836 VSS 3.85e-19
C8299 VDD.n1837 VSS 3.85e-19
C8300 VDD.n1838 VSS 3.87e-19
C8301 VDD.n1839 VSS 2.97e-19
C8302 VDD.n1840 VSS 2.97e-19
C8303 VDD.n1841 VSS 8.1e-19
C8304 VDD.n1842 VSS 0.0148f
C8305 VDD.n1843 VSS 0.0177f
C8306 VDD.n1844 VSS 0.0261f
C8307 VDD.n1845 VSS 0.0261f
C8308 VDD.n1846 VSS 0.00158f
C8309 VDD.n1847 VSS 6.55e-19
C8310 VDD.n1848 VSS 0.00152f
C8311 VDD.n1849 VSS 7.49e-19
C8312 VDD.n1850 VSS 7.49e-19
C8313 VDD.n1851 VSS 1.72e-19
C8314 VDD.n1852 VSS 5.4e-19
C8315 VDD.n1853 VSS 1.01e-19
C8316 VDD.t559 VSS 0.00476f
C8317 VDD.n1854 VSS 0.00578f
C8318 VDD.n1855 VSS 0.00108f
C8319 VDD.n1856 VSS 0.00114f
C8320 VDD.n1857 VSS 4.51e-19
C8321 VDD.n1858 VSS 2.02e-20
C8322 VDD.n1859 VSS 1.72e-19
C8323 VDD.n1860 VSS 2.85e-19
C8324 VDD.n1861 VSS 9.21e-19
C8325 VDD.n1862 VSS 9.88e-19
C8326 VDD.n1863 VSS 0.00126f
C8327 VDD.n1864 VSS 1.01e-19
C8328 VDD.n1865 VSS 2.01e-19
C8329 VDD.n1866 VSS 6.38e-19
C8330 VDD.n1867 VSS 7.08e-19
C8331 VDD.n1868 VSS 1.62e-19
C8332 VDD.n1869 VSS 5.06e-20
C8333 VDD.n1870 VSS 5.4e-19
C8334 VDD.n1871 VSS 1.01e-19
C8335 VDD.n1872 VSS 0.00578f
C8336 VDD.n1873 VSS 0.00108f
C8337 VDD.n1874 VSS 0.00483f
C8338 VDD.n1875 VSS 4.51e-19
C8339 VDD.n1876 VSS 2.02e-20
C8340 VDD.n1877 VSS 1.21e-19
C8341 VDD.n1878 VSS 1.62e-19
C8342 VDD.n1879 VSS 2.68e-19
C8343 VDD.n1880 VSS 3.52e-19
C8344 VDD.n1881 VSS 3.52e-19
C8345 VDD.n1882 VSS 4.52e-19
C8346 VDD.n1883 VSS 3.36e-19
C8347 VDD.n1884 VSS 0.00149f
C8348 VDD.n1885 VSS 8.1e-19
C8349 VDD.n1886 VSS 0.0296f
C8350 VDD.n1887 VSS 0.0975f
C8351 VDD.n1888 VSS 0.0975f
C8352 VDD.n1889 VSS 0.0271f
C8353 VDD.n1890 VSS 0.00149f
C8354 VDD.n1891 VSS 8.1e-19
C8355 VDD.n1892 VSS 4.13e-19
C8356 VDD.n1893 VSS 3.36e-19
C8357 VDD.n1894 VSS 4.35e-19
C8358 VDD.n1895 VSS 9.04e-19
C8359 VDD.t235 VSS 0.00578f
C8360 VDD.n1896 VSS 0.00835f
C8361 VDD.n1897 VSS 0.00109f
C8362 VDD.n1898 VSS 0.00172f
C8363 VDD.n1899 VSS 0.00241f
C8364 VDD.t9 VSS -2.71e-19
C8365 VDD.t236 VSS 8.49e-19
C8366 VDD.n1900 VSS 0.00391f
C8367 VDD.n1901 VSS 0.00413f
C8368 VDD.t8 VSS 0.00578f
C8369 VDD.n1902 VSS 0.00597f
C8370 VDD.n1903 VSS 0.00109f
C8371 VDD.n1904 VSS 9.92e-19
C8372 VDD.n1905 VSS 0.00308f
C8373 VDD.n1906 VSS 0.00231f
C8374 VDD.n1907 VSS 0.0018f
C8375 VDD.n1908 VSS 0.00109f
C8376 VDD.n1909 VSS 0.00773f
C8377 VDD.n1910 VSS 0.00109f
C8378 VDD.n1911 VSS 0.00151f
C8379 VDD.n1912 VSS 0.00183f
C8380 VDD.n1913 VSS 0.00308f
C8381 VDD.n1914 VSS 0.00905f
C8382 VDD.n1915 VSS 0.00109f
C8383 VDD.n1916 VSS 0.00118f
C8384 VDD.n1917 VSS 0.00308f
C8385 VDD.n1918 VSS 0.00308f
C8386 VDD.t266 VSS 0.00578f
C8387 VDD.n1919 VSS 0.00578f
C8388 VDD.n1920 VSS 0.00109f
C8389 VDD.n1921 VSS 0.00151f
C8390 VDD.n1922 VSS 0.00308f
C8391 VDD.t481 VSS 0.00578f
C8392 VDD.n1923 VSS 0.00528f
C8393 VDD.n1924 VSS 0.00109f
C8394 VDD.n1925 VSS 0.00186f
C8395 VDD.n1926 VSS 0.00308f
C8396 VDD.n1927 VSS 0.00754f
C8397 VDD.n1928 VSS 0.00109f
C8398 VDD.n1929 VSS 0.00177f
C8399 VDD.n1930 VSS 0.00308f
C8400 VDD.n1931 VSS 0.00308f
C8401 VDD.t577 VSS 0.00578f
C8402 VDD.n1932 VSS 0.00666f
C8403 VDD.n1933 VSS 0.00109f
C8404 VDD.n1934 VSS 0.00118f
C8405 VDD.n1935 VSS 0.00308f
C8406 VDD.t318 VSS 0.0054f
C8407 VDD.n1936 VSS 0.0059f
C8408 VDD.n1937 VSS 0.00109f
C8409 VDD.n1938 VSS 0.00186f
C8410 VDD.n1939 VSS 0.00308f
C8411 VDD.t362 VSS 0.00217f
C8412 VDD.t284 VSS 9.67e-19
C8413 VDD.n1940 VSS 0.00349f
C8414 VDD.n1941 VSS 0.00457f
C8415 VDD.t283 VSS 0.00565f
C8416 VDD.n1942 VSS 0.00616f
C8417 VDD.n1943 VSS 0.00109f
C8418 VDD.n1944 VSS 0.00102f
C8419 VDD.n1945 VSS 0.00308f
C8420 VDD.t361 VSS 0.00578f
C8421 VDD.n1946 VSS 0.00823f
C8422 VDD.n1947 VSS 0.00109f
C8423 VDD.n1948 VSS 0.0011f
C8424 VDD.n1949 VSS 0.00308f
C8425 VDD.n1950 VSS 0.00905f
C8426 VDD.n1951 VSS 0.00109f
C8427 VDD.n1952 VSS 0.00186f
C8428 VDD.n1953 VSS 0.00308f
C8429 VDD.t482 VSS 0.00578f
C8430 VDD.n1954 VSS 0.00528f
C8431 VDD.n1955 VSS 0.00109f
C8432 VDD.n1956 VSS 0.00186f
C8433 VDD.n1957 VSS 0.00308f
C8434 VDD.t263 VSS 0.00578f
C8435 VDD.n1958 VSS 0.00634f
C8436 VDD.n1959 VSS 0.00109f
C8437 VDD.n1960 VSS 0.00186f
C8438 VDD.n1961 VSS 0.00308f
C8439 VDD.t467 VSS 0.00578f
C8440 VDD.n1962 VSS 0.00603f
C8441 VDD.n1963 VSS 0.00109f
C8442 VDD.n1964 VSS 0.00132f
C8443 VDD.n1965 VSS 0.00308f
C8444 VDD.n1966 VSS 0.00308f
C8445 VDD.n1967 VSS 0.00666f
C8446 VDD.n1968 VSS 0.00109f
C8447 VDD.n1969 VSS 0.00164f
C8448 VDD.n1970 VSS 0.00308f
C8449 VDD.t285 VSS 0.00578f
C8450 VDD.t23 VSS 0.00578f
C8451 VDD.n1971 VSS 0.00452f
C8452 VDD.n1972 VSS 0.00109f
C8453 VDD.n1973 VSS 0.00172f
C8454 VDD.n1974 VSS 0.00308f
C8455 VDD.t286 VSS 0.00262f
C8456 VDD.n1975 VSS 0.00271f
C8457 VDD.t148 VSS 0.0139f
C8458 VDD.n1976 VSS 0.0119f
C8459 VDD.n1977 VSS 7.81e-19
C8460 VDD.n1978 VSS 0.00234f
C8461 VDD.n1979 VSS 0.00283f
C8462 VDD.n1980 VSS 0.00152f
C8463 VDD.n1981 VSS 2.51e-19
C8464 VDD.n1982 VSS 5.03e-20
C8465 VDD.t753 VSS 8.67e-19
C8466 VDD.n1983 VSS 0.00281f
C8467 VDD.t147 VSS 0.0016f
C8468 VDD.n1984 VSS 0.00355f
C8469 VDD.n1985 VSS 7.12e-19
C8470 VDD.n1986 VSS 0.00213f
C8471 VDD.n1987 VSS 3.51e-19
C8472 VDD.n1988 VSS 7.01e-20
C8473 VDD.n1989 VSS 3.74e-19
C8474 VDD.n1990 VSS 2.18e-19
C8475 VDD.n1991 VSS 2.35e-19
C8476 VDD.n1992 VSS 5.79e-19
C8477 VDD.n1993 VSS 3.36e-19
C8478 VDD.n1994 VSS 8.1e-19
C8479 VDD.n1995 VSS 0.00158f
C8480 VDD.n1996 VSS 0.00149f
C8481 VDD.n1997 VSS 4.64e-19
C8482 VDD.n1998 VSS 4e-19
C8483 VDD.n1999 VSS 2.97e-19
C8484 VDD.t293 VSS 0.00579f
C8485 VDD.n2000 VSS 0.00579f
C8486 VDD.n2001 VSS 0.00109f
C8487 VDD.n2002 VSS 0.00151f
C8488 VDD.n2003 VSS 0.00271f
C8489 VDD.n2004 VSS 0.00151f
C8490 VDD.t480 VSS 7.62e-19
C8491 VDD.t110 VSS 5.72e-19
C8492 VDD.n2005 VSS 0.0014f
C8493 VDD.t109 VSS 0.00579f
C8494 VDD.n2006 VSS 0.00762f
C8495 VDD.n2007 VSS 0.00111f
C8496 VDD.n2008 VSS 0.00204f
C8497 VDD.n2009 VSS 0.00252f
C8498 VDD.n2010 VSS 0.00109f
C8499 VDD.n2011 VSS 0.00168f
C8500 VDD.n2012 VSS 0.00231f
C8501 VDD.t476 VSS 8.49e-19
C8502 VDD.t334 VSS -2.71e-19
C8503 VDD.n2013 VSS 0.00391f
C8504 VDD.n2014 VSS 0.00413f
C8505 VDD.t333 VSS 0.00579f
C8506 VDD.n2015 VSS 0.00598f
C8507 VDD.n2016 VSS 0.00109f
C8508 VDD.n2017 VSS 9.92e-19
C8509 VDD.n2018 VSS 0.00308f
C8510 VDD.t475 VSS 0.00579f
C8511 VDD.n2019 VSS 0.00838f
C8512 VDD.n2020 VSS 0.00109f
C8513 VDD.n2021 VSS 0.00186f
C8514 VDD.n2022 VSS 0.00308f
C8515 VDD.n2023 VSS 0.00926f
C8516 VDD.n2024 VSS 9.85e-19
C8517 VDD.n2025 VSS 0.00163f
C8518 VDD.n2026 VSS 0.00307f
C8519 VDD.n2027 VSS 0.00154f
C8520 VDD.n2028 VSS 0.00164f
C8521 VDD.t607 VSS 9.16e-19
C8522 VDD.t478 VSS -5.07e-19
C8523 VDD.n2029 VSS 0.00359f
C8524 VDD.n2030 VSS 6.69e-19
C8525 VDD.n2031 VSS 0.00143f
C8526 VDD.n2032 VSS 3.97e-19
C8527 VDD.n2033 VSS 5.34e-19
C8528 VDD.n2034 VSS 1.01e-19
C8529 VDD.t477 VSS 0.00466f
C8530 VDD.n2035 VSS 0.0022f
C8531 VDD.n2036 VSS 0.00107f
C8532 VDD.n2037 VSS 0.0039f
C8533 VDD.n2038 VSS 5.58e-19
C8534 VDD.n2039 VSS 4.68e-20
C8535 VDD.n2040 VSS 1.4e-19
C8536 VDD.n2041 VSS 2.85e-19
C8537 VDD.n2042 VSS 0.00126f
C8538 VDD.n2043 VSS 0.00127f
C8539 VDD.n2044 VSS 0.00213f
C8540 VDD.n2045 VSS 3.97e-19
C8541 VDD.n2046 VSS 0.00178f
C8542 VDD.n2047 VSS 5.4e-19
C8543 VDD.n2048 VSS 1.01e-19
C8544 VDD.n2049 VSS 0.00573f
C8545 VDD.n2050 VSS 0.00107f
C8546 VDD.t606 VSS 0.00586f
C8547 VDD.n2051 VSS 0.00208f
C8548 VDD.n2052 VSS 5.58e-19
C8549 VDD.n2053 VSS 4.21e-19
C8550 VDD.n2054 VSS 0.00183f
C8551 VDD.t49 VSS 0.00262f
C8552 VDD.n2055 VSS 0.00271f
C8553 VDD.n2056 VSS 0.00882f
C8554 VDD.n2057 VSS 9.91e-19
C8555 VDD.n2058 VSS 0.00229f
C8556 VDD.n2059 VSS 0.00308f
C8557 VDD.t325 VSS 0.00579f
C8558 VDD.t48 VSS 0.00579f
C8559 VDD.n2060 VSS 0.00453f
C8560 VDD.n2061 VSS 0.00109f
C8561 VDD.n2062 VSS 0.00172f
C8562 VDD.n2063 VSS 0.00308f
C8563 VDD.n2064 VSS 0.00668f
C8564 VDD.n2065 VSS 0.00109f
C8565 VDD.n2066 VSS 0.00164f
C8566 VDD.n2067 VSS 0.00308f
C8567 VDD.n2068 VSS 0.00308f
C8568 VDD.t479 VSS 0.00579f
C8569 VDD.n2069 VSS 0.00605f
C8570 VDD.n2070 VSS 0.00109f
C8571 VDD.n2071 VSS 0.00132f
C8572 VDD.n2072 VSS 0.00308f
C8573 VDD.t294 VSS 0.00579f
C8574 VDD.n2073 VSS 0.00636f
C8575 VDD.n2074 VSS 0.00109f
C8576 VDD.n2075 VSS 0.00186f
C8577 VDD.n2076 VSS 0.00308f
C8578 VDD.t72 VSS 0.00579f
C8579 VDD.n2077 VSS 0.00529f
C8580 VDD.n2078 VSS 0.00109f
C8581 VDD.n2079 VSS 0.00186f
C8582 VDD.n2080 VSS 0.00308f
C8583 VDD.n2081 VSS 0.00907f
C8584 VDD.n2082 VSS 0.00109f
C8585 VDD.n2083 VSS 0.00186f
C8586 VDD.n2084 VSS 0.00308f
C8587 VDD.t21 VSS 0.00579f
C8588 VDD.n2085 VSS 0.00825f
C8589 VDD.n2086 VSS 0.00109f
C8590 VDD.n2087 VSS 0.0011f
C8591 VDD.n2088 VSS 0.00308f
C8592 VDD.t51 VSS 9.67e-19
C8593 VDD.t22 VSS 0.00217f
C8594 VDD.n2089 VSS 0.00349f
C8595 VDD.n2090 VSS 0.00457f
C8596 VDD.t50 VSS 0.00567f
C8597 VDD.n2091 VSS 0.00617f
C8598 VDD.n2092 VSS 0.00109f
C8599 VDD.n2093 VSS 0.00102f
C8600 VDD.n2094 VSS 0.00308f
C8601 VDD.t88 VSS 0.0134f
C8602 VDD.t248 VSS 0.00542f
C8603 VDD.n2095 VSS 0.0068f
C8604 VDD.n2096 VSS 0.00103f
C8605 VDD.n2097 VSS 0.00176f
C8606 VDD.n2098 VSS 0.00291f
C8607 VDD.n2099 VSS 0.00154f
C8608 VDD.n2100 VSS 1.36e-19
C8609 VDD.t108 VSS 0.00149f
C8610 VDD.t772 VSS 6.37e-19
C8611 VDD.n2101 VSS 0.00279f
C8612 VDD.n2102 VSS 2.33e-19
C8613 VDD.n2103 VSS 6.77e-19
C8614 VDD.n2104 VSS 0.00141f
C8615 VDD.n2105 VSS 2.33e-19
C8616 VDD.n2106 VSS 0.00388f
C8617 VDD.n2107 VSS 5.31e-19
C8618 VDD.n2108 VSS 0.00105f
C8619 VDD.t770 VSS 6.29e-19
C8620 VDD.n2109 VSS 0.00315f
C8621 VDD.t87 VSS 0.00189f
C8622 VDD.n2110 VSS 0.00174f
C8623 VDD.n2111 VSS 2.32e-19
C8624 VDD.n2112 VSS 9.31e-19
C8625 VDD.n2113 VSS 1.72e-19
C8626 VDD.n2114 VSS 2.85e-19
C8627 VDD.n2115 VSS 0.00146f
C8628 VDD.n2116 VSS 0.00198f
C8629 VDD.t20 VSS 5.42e-19
C8630 VDD.t89 VSS 5.72e-19
C8631 VDD.n2117 VSS 0.00119f
C8632 VDD.n2118 VSS 0.00282f
C8633 VDD.n2119 VSS 0.00296f
C8634 VDD.t19 VSS 0.0107f
C8635 VDD.n2120 VSS 0.00756f
C8636 VDD.n2121 VSS 0.0011f
C8637 VDD.n2122 VSS 0.00177f
C8638 VDD.n2123 VSS 0.00273f
C8639 VDD.n2124 VSS 0.00154f
C8640 VDD.t73 VSS 0.00579f
C8641 VDD.n2125 VSS 0.00529f
C8642 VDD.n2126 VSS 0.00109f
C8643 VDD.n2127 VSS 0.00186f
C8644 VDD.n2128 VSS 3.85e-19
C8645 VDD.n2129 VSS 3.68e-19
C8646 VDD.n2130 VSS 2.84e-19
C8647 VDD.n2131 VSS 8.1e-19
C8648 VDD.n2132 VSS 0.00158f
C8649 VDD.n2133 VSS 0.00149f
C8650 VDD.n2134 VSS 5.92e-19
C8651 VDD.n2135 VSS 5.16e-19
C8652 VDD.n2136 VSS 3.36e-19
C8653 VDD.n2137 VSS 8.1e-19
C8654 VDD.n2138 VSS 0.0256f
C8655 VDD.n2139 VSS 0.0296f
C8656 VDD.n2140 VSS 0.0931f
C8657 VDD.n2141 VSS 0.29f
C8658 VDD.n2142 VSS 2.12f
C8659 VDD.n2143 VSS 0.032f
C8660 VDD.n2144 VSS 0.0064f
C8661 VDD.n2145 VSS 0.00936f
C8662 VDD.n2146 VSS 0.0138f
C8663 VDD.n2147 VSS 0.0064f
C8664 VDD.n2148 VSS 0.00936f
C8665 VDD.n2149 VSS 0.00149f
C8666 VDD.n2150 VSS 8.1e-19
C8667 VDD.n2151 VSS 6.93e-19
C8668 VDD.n2152 VSS 3.36e-19
C8669 VDD.n2153 VSS 4.35e-19
C8670 VDD.n2154 VSS 6.2e-19
C8671 VDD.n2155 VSS 8.54e-19
C8672 VDD.n2156 VSS 7.49e-19
C8673 VDD.n2157 VSS 7.49e-19
C8674 VDD.n2158 VSS 1.72e-19
C8675 VDD.n2159 VSS 5.4e-19
C8676 VDD.n2160 VSS 1.01e-19
C8677 VDD.n2161 VSS 0.00578f
C8678 VDD.n2162 VSS 0.00108f
C8679 VDD.n2163 VSS 0.00483f
C8680 VDD.n2164 VSS 4.51e-19
C8681 VDD.n2165 VSS 2.02e-20
C8682 VDD.n2166 VSS 1.72e-19
C8683 VDD.n2167 VSS 2.85e-19
C8684 VDD.n2168 VSS 0.00127f
C8685 VDD.n2169 VSS 0.00152f
C8686 VDD.n2170 VSS 7.49e-19
C8687 VDD.n2171 VSS 7.49e-19
C8688 VDD.n2172 VSS 1.72e-19
C8689 VDD.n2173 VSS 5.4e-19
C8690 VDD.n2174 VSS 1.01e-19
C8691 VDD.n2175 VSS 0.00457f
C8692 VDD.t255 VSS 0.00102f
C8693 VDD.n2176 VSS 8.26e-19
C8694 VDD.n2177 VSS 0.00483f
C8695 VDD.n2178 VSS 4.51e-19
C8696 VDD.n2179 VSS 2.02e-20
C8697 VDD.n2180 VSS 1.72e-19
C8698 VDD.n2181 VSS 2.85e-19
C8699 VDD.n2182 VSS 0.00127f
C8700 VDD.n2183 VSS 0.00152f
C8701 VDD.n2184 VSS 7.49e-19
C8702 VDD.t599 VSS 5.42e-19
C8703 VDD.t171 VSS 4.25e-19
C8704 VDD.n2185 VSS 0.00111f
C8705 VDD.n2186 VSS 0.00224f
C8706 VDD.n2187 VSS 4.45e-19
C8707 VDD.n2188 VSS 1.72e-19
C8708 VDD.n2189 VSS 5.4e-19
C8709 VDD.n2190 VSS 1.01e-19
C8710 VDD.t598 VSS 0.00476f
C8711 VDD.n2191 VSS 0.00559f
C8712 VDD.n2192 VSS 0.00108f
C8713 VDD.n2193 VSS 5.08e-19
C8714 VDD.n2194 VSS 4.51e-19
C8715 VDD.n2195 VSS 2.02e-20
C8716 VDD.n2196 VSS 1.72e-19
C8717 VDD.n2197 VSS 2.85e-19
C8718 VDD.n2198 VSS 0.00127f
C8719 VDD.n2199 VSS 0.00152f
C8720 VDD.n2200 VSS 4.66e-19
C8721 VDD.n2201 VSS 7.49e-19
C8722 VDD.n2202 VSS 1.72e-19
C8723 VDD.n2203 VSS 5.4e-19
C8724 VDD.n2204 VSS 1.01e-19
C8725 VDD.t170 VSS 0.00476f
C8726 VDD.n2205 VSS 0.00578f
C8727 VDD.n2206 VSS 0.00108f
C8728 VDD.n2207 VSS 2.54e-19
C8729 VDD.n2208 VSS 4.51e-19
C8730 VDD.n2209 VSS 2.02e-20
C8731 VDD.n2210 VSS 1.72e-19
C8732 VDD.n2211 VSS 2.85e-19
C8733 VDD.n2212 VSS 0.00127f
C8734 VDD.n2213 VSS 0.00152f
C8735 VDD.n2214 VSS 7.49e-19
C8736 VDD.n2215 VSS 0.0117f
C8737 VDD.n2216 VSS 0.00109f
C8738 VDD.n2217 VSS 0.00157f
C8739 VDD.n2218 VSS 0.0117f
C8740 VDD.n2219 VSS 0.00109f
C8741 VDD.n2220 VSS 0.00157f
C8742 VDD.n2221 VSS 0.0107f
C8743 VDD.n2222 VSS 9.97e-19
C8744 VDD.n2223 VSS 0.00143f
C8745 VDD.n2224 VSS 9.1e-19
C8746 VDD.n2225 VSS 1.72e-19
C8747 VDD.n2226 VSS 5.46e-19
C8748 VDD.n2227 VSS 1.01e-19
C8749 VDD.n2228 VSS 0.00584f
C8750 VDD.n2229 VSS 0.00108f
C8751 VDD.n2230 VSS 0.00483f
C8752 VDD.n2231 VSS 4.51e-19
C8753 VDD.n2232 VSS 2.02e-20
C8754 VDD.n2233 VSS 1.72e-19
C8755 VDD.n2234 VSS 2.85e-19
C8756 VDD.n2235 VSS 7.71e-19
C8757 VDD.n2236 VSS 0.0117f
C8758 VDD.n2237 VSS 0.00109f
C8759 VDD.n2238 VSS 0.00157f
C8760 VDD.n2239 VSS 0.0117f
C8761 VDD.n2240 VSS 0.00109f
C8762 VDD.n2241 VSS 0.00157f
C8763 VDD.n2242 VSS 0.0117f
C8764 VDD.n2243 VSS 0.00109f
C8765 VDD.n2244 VSS 0.00157f
C8766 VDD.n2245 VSS 0.0117f
C8767 VDD.n2246 VSS 0.00109f
C8768 VDD.n2247 VSS 0.00129f
C8769 VDD.n2248 VSS 0.00927f
C8770 VDD.n2249 VSS 0.00109f
C8771 VDD.n2250 VSS 9.31e-19
C8772 VDD.n2251 VSS 9.39e-19
C8773 VDD.n2252 VSS 0.0125f
C8774 VDD.t441 VSS 0.00584f
C8775 VDD.n2253 VSS 0.0061f
C8776 VDD.n2254 VSS 0.00109f
C8777 VDD.n2255 VSS 4.66e-19
C8778 VDD.n2256 VSS 9.31e-19
C8779 VDD.n2257 VSS 0.00308f
C8780 VDD.t442 VSS 4.25e-19
C8781 VDD.t69 VSS 5.42e-19
C8782 VDD.n2258 VSS 0.00111f
C8783 VDD.n2259 VSS 0.00218f
C8784 VDD.t68 VSS 0.00584f
C8785 VDD.t282 VSS 0.00584f
C8786 VDD.n2260 VSS 0.00457f
C8787 VDD.n2261 VSS 0.00109f
C8788 VDD.n2262 VSS 9.31e-19
C8789 VDD.n2263 VSS 8.7e-19
C8790 VDD.n2264 VSS 0.00308f
C8791 VDD.n2265 VSS 0.00927f
C8792 VDD.n2266 VSS 0.00109f
C8793 VDD.n2267 VSS 9.31e-19
C8794 VDD.n2268 VSS 9.31e-19
C8795 VDD.n2269 VSS 0.00308f
C8796 VDD.n2270 VSS 0.0102f
C8797 VDD.n2271 VSS 0.00109f
C8798 VDD.n2272 VSS 9.31e-19
C8799 VDD.n2273 VSS 9.31e-19
C8800 VDD.n2274 VSS 0.00308f
C8801 VDD.t563 VSS 0.00584f
C8802 VDD.n2275 VSS 0.00654f
C8803 VDD.n2276 VSS 0.00109f
C8804 VDD.n2277 VSS 9.31e-19
C8805 VDD.n2278 VSS 9.31e-19
C8806 VDD.n2279 VSS 0.00308f
C8807 VDD.t443 VSS 0.00584f
C8808 VDD.n2280 VSS 0.00667f
C8809 VDD.n2281 VSS 0.00109f
C8810 VDD.n2282 VSS 9.31e-19
C8811 VDD.n2283 VSS 9.31e-19
C8812 VDD.n2284 VSS 0.00308f
C8813 VDD.n2285 VSS 0.00116f
C8814 VDD.n2286 VSS 0.00253f
C8815 VDD.n2287 VSS 5.46e-19
C8816 VDD.n2288 VSS 0.00255f
C8817 VDD.n2289 VSS 8.4e-19
C8818 VDD.n2290 VSS 0.00109f
C8819 VDD.n2291 VSS 0.0061f
C8820 VDD.t623 VSS 0.00152f
C8821 VDD.n2292 VSS 0.0102f
C8822 VDD.n2293 VSS 0.00109f
C8823 VDD.n2294 VSS 0.00112f
C8824 VDD.n2295 VSS 4.05e-19
C8825 VDD.n2296 VSS 1.72e-19
C8826 VDD.n2297 VSS 5.26e-19
C8827 VDD.n2298 VSS 3.85e-19
C8828 VDD.n2299 VSS 2.85e-19
C8829 VDD.n2300 VSS 2.68e-19
C8830 VDD.n2301 VSS 0.00295f
C8831 VDD.n2302 VSS 3.01e-19
C8832 VDD.n2303 VSS 2.85e-19
C8833 VDD.n2304 VSS 1.72e-19
C8834 VDD.n2305 VSS 7.49e-19
C8835 VDD.n2306 VSS 1.72e-19
C8836 VDD.n2307 VSS 2.02e-20
C8837 VDD.n2308 VSS 5.46e-19
C8838 VDD.n2309 VSS 0.00584f
C8839 VDD.n2310 VSS 0.00108f
C8840 VDD.n2311 VSS 0.00292f
C8841 VDD.t17 VSS 0.00279f
C8842 VDD.n2312 VSS 0.004f
C8843 VDD.n2313 VSS 0.00108f
C8844 VDD.n2314 VSS 0.00203f
C8845 VDD.n2315 VSS 4.51e-19
C8846 VDD.n2316 VSS 2.02e-20
C8847 VDD.n2317 VSS 3.04e-20
C8848 VDD.n2318 VSS 0.0023f
C8849 VDD.n2319 VSS 1.42e-19
C8850 VDD.n2320 VSS 2.68e-19
C8851 VDD.n2321 VSS 4.02e-19
C8852 VDD.n2322 VSS 4.19e-19
C8853 VDD.n2323 VSS 4.13e-19
C8854 VDD.n2324 VSS 3.36e-19
C8855 VDD.n2325 VSS 0.00149f
C8856 VDD.n2326 VSS 8.1e-19
C8857 VDD.n2327 VSS 0.0271f
C8858 VDD.n2328 VSS 0.0916f
C8859 VDD.n2329 VSS 0.0916f
C8860 VDD.n2330 VSS 0.0296f
C8861 VDD.n2331 VSS 0.00149f
C8862 VDD.n2332 VSS 8.1e-19
C8863 VDD.n2333 VSS 4.52e-19
C8864 VDD.n2334 VSS 3.36e-19
C8865 VDD.n2335 VSS 4.35e-19
C8866 VDD.n2336 VSS 9.31e-19
C8867 VDD.n2337 VSS 5.53e-19
C8868 VDD.n2338 VSS 2.85e-19
C8869 VDD.n2339 VSS 2.85e-19
C8870 VDD.n2340 VSS 1.72e-19
C8871 VDD.n2341 VSS 0.00109f
C8872 VDD.t257 VSS 0.00472f
C8873 VDD.t596 VSS 0.00579f
C8874 VDD.n2342 VSS 0.00529f
C8875 VDD.n2343 VSS 0.00111f
C8876 VDD.n2344 VSS 0.00197f
C8877 VDD.n2345 VSS 0.0027f
C8878 VDD.n2346 VSS 0.0028f
C8879 VDD.n2347 VSS 0.00907f
C8880 VDD.n2348 VSS 0.00109f
C8881 VDD.n2349 VSS 0.00118f
C8882 VDD.n2350 VSS 0.00308f
C8883 VDD.t340 VSS 0.00142f
C8884 VDD.t339 VSS 0.00579f
C8885 VDD.n2351 VSS 0.00857f
C8886 VDD.n2352 VSS 0.00111f
C8887 VDD.n2353 VSS 0.00203f
C8888 VDD.n2354 VSS 0.00312f
C8889 VDD.n2355 VSS 0.00308f
C8890 VDD.t594 VSS 0.00579f
C8891 VDD.n2356 VSS 0.00579f
C8892 VDD.n2357 VSS 0.00109f
C8893 VDD.n2358 VSS 0.00151f
C8894 VDD.n2359 VSS 0.00308f
C8895 VDD.t167 VSS 0.00579f
C8896 VDD.n2360 VSS 0.00529f
C8897 VDD.n2361 VSS 0.00109f
C8898 VDD.n2362 VSS 0.00181f
C8899 VDD.n2363 VSS 0.003f
C8900 VDD.n2364 VSS 0.00154f
C8901 VDD.n2365 VSS 9.31e-19
C8902 VDD.t302 VSS 0.0107f
C8903 VDD.n2366 VSS 0.00756f
C8904 VDD.n2367 VSS 0.00103f
C8905 VDD.n2368 VSS 1.72e-19
C8906 VDD.n2369 VSS 2.85e-19
C8907 VDD.n2370 VSS 8.4e-19
C8908 VDD.n2371 VSS 5.53e-19
C8909 VDD.n2372 VSS 9.88e-19
C8910 VDD.n2373 VSS 4.35e-19
C8911 VDD.n2374 VSS 3.36e-19
C8912 VDD.n2375 VSS 8.1e-19
C8913 VDD.n2376 VSS 0.0177f
C8914 VDD.n2377 VSS 0.0281f
C8915 VDD.n2378 VSS 0.0281f
C8916 VDD.n2379 VSS 0.00158f
C8917 VDD.n2380 VSS 0.00149f
C8918 VDD.n2381 VSS 5.16e-19
C8919 VDD.n2382 VSS 0.00144f
C8920 VDD.n2383 VSS 7.49e-19
C8921 VDD.n2384 VSS 7.49e-19
C8922 VDD.n2385 VSS 1.72e-19
C8923 VDD.n2386 VSS 5.4e-19
C8924 VDD.n2387 VSS 1.01e-19
C8925 VDD.n2388 VSS 0.00457f
C8926 VDD.t35 VSS 0.00102f
C8927 VDD.n2389 VSS 8.26e-19
C8928 VDD.n2390 VSS 0.00483f
C8929 VDD.n2391 VSS 4.51e-19
C8930 VDD.n2392 VSS 2.02e-20
C8931 VDD.n2393 VSS 1.72e-19
C8932 VDD.n2394 VSS 2.85e-19
C8933 VDD.n2395 VSS 0.00111f
C8934 VDD.n2396 VSS 0.00126f
C8935 VDD.n2397 VSS 2.68e-19
C8936 VDD.n2398 VSS 7.71e-19
C8937 VDD.n2399 VSS 7.49e-19
C8938 VDD.n2400 VSS 0.0117f
C8939 VDD.n2401 VSS 0.00109f
C8940 VDD.n2402 VSS 0.00157f
C8941 VDD.n2403 VSS 0.0117f
C8942 VDD.n2404 VSS 0.00109f
C8943 VDD.n2405 VSS 0.00157f
C8944 VDD.n2406 VSS 0.0107f
C8945 VDD.n2407 VSS 9.97e-19
C8946 VDD.n2408 VSS 0.00143f
C8947 VDD.n2409 VSS 9.1e-19
C8948 VDD.n2410 VSS 1.72e-19
C8949 VDD.n2411 VSS 5.46e-19
C8950 VDD.n2412 VSS 1.01e-19
C8951 VDD.n2413 VSS 0.00584f
C8952 VDD.n2414 VSS 0.00108f
C8953 VDD.n2415 VSS 0.00483f
C8954 VDD.n2416 VSS 4.51e-19
C8955 VDD.n2417 VSS 2.02e-20
C8956 VDD.n2418 VSS 1.72e-19
C8957 VDD.n2419 VSS 2.85e-19
C8958 VDD.n2420 VSS 0.00152f
C8959 VDD.n2421 VSS 0.00127f
C8960 VDD.n2422 VSS 4.66e-19
C8961 VDD.n2423 VSS 7.49e-19
C8962 VDD.n2424 VSS 1.72e-19
C8963 VDD.n2425 VSS 5.4e-19
C8964 VDD.n2426 VSS 1.01e-19
C8965 VDD.t78 VSS 0.00476f
C8966 VDD.n2427 VSS 0.00578f
C8967 VDD.n2428 VSS 0.00108f
C8968 VDD.n2429 VSS 2.54e-19
C8969 VDD.n2430 VSS 4.51e-19
C8970 VDD.n2431 VSS 2.02e-20
C8971 VDD.n2432 VSS 1.72e-19
C8972 VDD.n2433 VSS 2.85e-19
C8973 VDD.n2434 VSS 0.00126f
C8974 VDD.n2435 VSS 0.00126f
C8975 VDD.n2436 VSS 2.85e-19
C8976 VDD.n2437 VSS 7.49e-19
C8977 VDD.t368 VSS 5.42e-19
C8978 VDD.t79 VSS 4.25e-19
C8979 VDD.n2438 VSS 0.00111f
C8980 VDD.n2439 VSS 0.00224f
C8981 VDD.n2440 VSS 2.93e-19
C8982 VDD.n2441 VSS 1.62e-19
C8983 VDD.n2442 VSS 1.62e-19
C8984 VDD.n2443 VSS 5.4e-19
C8985 VDD.n2444 VSS 1.01e-19
C8986 VDD.t367 VSS 0.00476f
C8987 VDD.n2445 VSS 0.00559f
C8988 VDD.n2446 VSS 0.00108f
C8989 VDD.n2447 VSS 5.08e-19
C8990 VDD.n2448 VSS 4.51e-19
C8991 VDD.n2449 VSS 2.02e-20
C8992 VDD.n2450 VSS 1.72e-19
C8993 VDD.n2451 VSS 1.84e-19
C8994 VDD.n2452 VSS 2.68e-19
C8995 VDD.n2453 VSS 5.92e-19
C8996 VDD.n2454 VSS 3.36e-19
C8997 VDD.n2455 VSS 8.1e-19
C8998 VDD.n2456 VSS 0.0296f
C8999 VDD.n2457 VSS 0.0202f
C9000 VDD.n2458 VSS 0.0202f
C9001 VDD.n2459 VSS 0.00158f
C9002 VDD.n2460 VSS 3.1e-19
C9003 VDD.n2461 VSS 3.23e-19
C9004 VDD.n2462 VSS 0.00154f
C9005 VDD.n2463 VSS 0.00666f
C9006 VDD.n2464 VSS 0.00109f
C9007 VDD.n2465 VSS 0.00164f
C9008 VDD.n2466 VSS 4.19e-19
C9009 VDD.t25 VSS 5.72e-19
C9010 VDD.t238 VSS 7.62e-19
C9011 VDD.n2467 VSS 0.0014f
C9012 VDD.t24 VSS 0.00578f
C9013 VDD.n2468 VSS 0.0076f
C9014 VDD.n2469 VSS 0.00111f
C9015 VDD.n2470 VSS 0.00189f
C9016 VDD.n2471 VSS 0.00252f
C9017 VDD.n2472 VSS 0.00241f
C9018 VDD.n2473 VSS 0.00142f
C9019 VDD.n2474 VSS 4.19e-19
C9020 VDD.n2475 VSS 4.9e-19
C9021 VDD.n2476 VSS 3.23e-19
C9022 VDD.n2477 VSS 0.00149f
C9023 VDD.n2478 VSS 8.1e-19
C9024 VDD.n2479 VSS 0.0207f
C9025 VDD.n2480 VSS 0.0148f
C9026 VDD.n2481 VSS 0.0148f
C9027 VDD.n2482 VSS 0.00149f
C9028 VDD.n2483 VSS 0.00186f
C9029 VDD.t303 VSS 5.42e-19
C9030 VDD.t131 VSS 5.72e-19
C9031 VDD.n2484 VSS 0.00119f
C9032 VDD.n2485 VSS 0.00282f
C9033 VDD.n2486 VSS 0.00232f
C9034 VDD.n2487 VSS 0.00146f
C9035 VDD.n2488 VSS 1.36e-19
C9036 VDD.t90 VSS 0.00149f
C9037 VDD.t754 VSS 6.37e-19
C9038 VDD.n2489 VSS 0.00279f
C9039 VDD.n2490 VSS 2.33e-19
C9040 VDD.n2491 VSS 6.77e-19
C9041 VDD.n2492 VSS 0.00141f
C9042 VDD.n2493 VSS 2.33e-19
C9043 VDD.n2494 VSS 0.00388f
C9044 VDD.n2495 VSS 5.31e-19
C9045 VDD.n2496 VSS 0.00105f
C9046 VDD.t755 VSS 6.29e-19
C9047 VDD.n2497 VSS 0.00315f
C9048 VDD.t129 VSS 0.00189f
C9049 VDD.n2498 VSS 0.00174f
C9050 VDD.n2499 VSS 2.32e-19
C9051 VDD.n2500 VSS 9.31e-19
C9052 VDD.n2501 VSS 1.72e-19
C9053 VDD.n2502 VSS 2.85e-19
C9054 VDD.n2503 VSS 8.21e-19
C9055 VDD.t403 VSS 0.00567f
C9056 VDD.n2504 VSS 0.00617f
C9057 VDD.n2505 VSS 0.00109f
C9058 VDD.t404 VSS 9.67e-19
C9059 VDD.t301 VSS 0.00217f
C9060 VDD.n2506 VSS 0.00349f
C9061 VDD.n2507 VSS 0.00443f
C9062 VDD.n2508 VSS 0.00102f
C9063 VDD.n2509 VSS 0.00243f
C9064 VDD.t130 VSS 0.0134f
C9065 VDD.t668 VSS 0.00542f
C9066 VDD.n2510 VSS 0.0068f
C9067 VDD.n2511 VSS 0.00115f
C9068 VDD.n2512 VSS 0.00176f
C9069 VDD.n2513 VSS 0.00226f
C9070 VDD.n2514 VSS 0.00137f
C9071 VDD.n2515 VSS 0.00144f
C9072 VDD.n2516 VSS 0.00157f
C9073 VDD.n2517 VSS 8.1e-19
C9074 VDD.n2518 VSS 0.0207f
C9075 VDD.n2519 VSS 0.0537f
C9076 VDD.n2520 VSS 0.0434f
C9077 VDD.n2521 VSS 0.0148f
C9078 VDD.n2522 VSS 0.00158f
C9079 VDD.n2523 VSS 0.00149f
C9080 VDD.n2524 VSS 8.1e-19
C9081 VDD.n2525 VSS 0.00158f
C9082 VDD.n2526 VSS 0.00149f
C9083 VDD.n2527 VSS 6.68e-19
C9084 VDD.n2528 VSS 4.39e-19
C9085 VDD.n2529 VSS 9.55e-19
C9086 VDD.n2530 VSS 0.00109f
C9087 VDD.n2531 VSS 0.00109f
C9088 VDD.n2532 VSS 0.00882f
C9089 VDD.t547 VSS 0.00472f
C9090 VDD.t221 VSS 0.00579f
C9091 VDD.n2533 VSS 0.00529f
C9092 VDD.n2534 VSS 0.00111f
C9093 VDD.n2535 VSS 0.00202f
C9094 VDD.t751 VSS 0.0107f
C9095 VDD.n2536 VSS 0.00756f
C9096 VDD.n2537 VSS 0.00126f
C9097 VDD.n2538 VSS 0.00176f
C9098 VDD.n2539 VSS 0.00269f
C9099 VDD.n2540 VSS 0.00137f
C9100 VDD.n2541 VSS 6.05e-19
C9101 VDD.n2542 VSS 0.00158f
C9102 VDD.n2543 VSS 4.95e-19
C9103 VDD.n2544 VSS 0.00198f
C9104 VDD.t752 VSS 5.42e-19
C9105 VDD.t122 VSS 5.72e-19
C9106 VDD.n2545 VSS 0.00119f
C9107 VDD.n2546 VSS 0.00282f
C9108 VDD.n2547 VSS 0.00154f
C9109 VDD.n2548 VSS 5.38e-19
C9110 VDD.n2549 VSS 0.00154f
C9111 VDD.n2550 VSS 1.36e-19
C9112 VDD.t132 VSS 0.00149f
C9113 VDD.t760 VSS 6.37e-19
C9114 VDD.n2551 VSS 0.00279f
C9115 VDD.n2552 VSS 2.33e-19
C9116 VDD.n2553 VSS 6.77e-19
C9117 VDD.n2554 VSS 0.00141f
C9118 VDD.n2555 VSS 2.33e-19
C9119 VDD.n2556 VSS 0.00388f
C9120 VDD.n2557 VSS 5.31e-19
C9121 VDD.n2558 VSS 0.00105f
C9122 VDD.t758 VSS 6.29e-19
C9123 VDD.n2559 VSS 0.00315f
C9124 VDD.t120 VSS 0.00189f
C9125 VDD.n2560 VSS 0.00174f
C9126 VDD.n2561 VSS 2.32e-19
C9127 VDD.n2562 VSS 9.31e-19
C9128 VDD.n2563 VSS 1.72e-19
C9129 VDD.n2564 VSS 2.85e-19
C9130 VDD.n2565 VSS 8.76e-19
C9131 VDD.n2566 VSS 9.59e-19
C9132 VDD.n2567 VSS 4.35e-19
C9133 VDD.n2568 VSS 6.17e-19
C9134 VDD.n2569 VSS 3.36e-19
C9135 VDD.n2570 VSS 0.00149f
C9136 VDD.n2571 VSS 8.1e-19
C9137 VDD.n2572 VSS 0.00157f
C9138 VDD.n2573 VSS 0.0058f
C9139 VDD.n2574 VSS 0.00158f
C9140 VDD.n2575 VSS 6.55e-19
C9141 VDD.t452 VSS 0.00579f
C9142 VDD.n2576 VSS 0.00529f
C9143 VDD.n2577 VSS 0.00109f
C9144 VDD.n2578 VSS 0.00172f
C9145 VDD.n2579 VSS 0.00241f
C9146 VDD.t224 VSS 0.00579f
C9147 VDD.n2580 VSS 0.00636f
C9148 VDD.n2581 VSS 0.00109f
C9149 VDD.n2582 VSS 0.00186f
C9150 VDD.n2583 VSS 0.00308f
C9151 VDD.t60 VSS 0.00579f
C9152 VDD.n2584 VSS 0.00605f
C9153 VDD.n2585 VSS 0.00109f
C9154 VDD.n2586 VSS 0.00132f
C9155 VDD.n2587 VSS 0.00246f
C9156 VDD.n2588 VSS 0.00101f
C9157 VDD.t321 VSS 0.00472f
C9158 VDD.t83 VSS 0.00579f
C9159 VDD.n2589 VSS 0.00529f
C9160 VDD.n2590 VSS 0.00111f
C9161 VDD.n2591 VSS 0.00202f
C9162 VDD.t322 VSS 6.03e-19
C9163 VDD.t84 VSS 6.03e-19
C9164 VDD.n2592 VSS 0.0013f
C9165 VDD.n2593 VSS 0.0027f
C9166 VDD.t674 VSS 0.00142f
C9167 VDD.t673 VSS 0.00579f
C9168 VDD.n2594 VSS 0.00857f
C9169 VDD.n2595 VSS 0.00111f
C9170 VDD.n2596 VSS 0.00203f
C9171 VDD.n2597 VSS 0.00312f
C9172 VDD.n2598 VSS 0.00154f
C9173 VDD.n2599 VSS 0.00907f
C9174 VDD.n2600 VSS 0.00109f
C9175 VDD.n2601 VSS 0.00186f
C9176 VDD.n2602 VSS 0.00231f
C9177 VDD.t386 VSS 0.00579f
C9178 VDD.n2603 VSS 0.00825f
C9179 VDD.n2604 VSS 0.00109f
C9180 VDD.n2605 VSS 0.0011f
C9181 VDD.n2606 VSS 0.00266f
C9182 VDD.n2607 VSS 0.00144f
C9183 VDD.n2608 VSS 3.36e-19
C9184 VDD.n2609 VSS 3.1e-19
C9185 VDD.n2610 VSS 4.82e-19
C9186 VDD.n2611 VSS 0.00158f
C9187 VDD.n2612 VSS 0.00605f
C9188 VDD.n2613 VSS 0.00158f
C9189 VDD.n2614 VSS 4.26e-19
C9190 VDD.n2615 VSS 6.85e-19
C9191 VDD.n2616 VSS 0.00127f
C9192 VDD.n2617 VSS 7.18e-19
C9193 VDD.n2618 VSS 0.00926f
C9194 VDD.n2619 VSS 0.0011f
C9195 VDD.n2620 VSS 1.72e-19
C9196 VDD.n2621 VSS 2.85e-19
C9197 VDD.n2622 VSS 9.31e-19
C9198 VDD.n2623 VSS 6.37e-19
C9199 VDD.t343 VSS 0.00472f
C9200 VDD.t731 VSS 0.00579f
C9201 VDD.n2624 VSS 0.00529f
C9202 VDD.n2625 VSS 0.00111f
C9203 VDD.n2626 VSS 0.00202f
C9204 VDD.t344 VSS 6.03e-19
C9205 VDD.t732 VSS 6.03e-19
C9206 VDD.n2627 VSS 0.0013f
C9207 VDD.n2628 VSS 0.0027f
C9208 VDD.t177 VSS 0.00142f
C9209 VDD.t176 VSS 0.00579f
C9210 VDD.n2629 VSS 0.00857f
C9211 VDD.n2630 VSS 0.00111f
C9212 VDD.n2631 VSS 0.00203f
C9213 VDD.n2632 VSS 0.00312f
C9214 VDD.n2633 VSS 0.00154f
C9215 VDD.n2634 VSS 0.00668f
C9216 VDD.n2635 VSS 0.00109f
C9217 VDD.n2636 VSS 0.00164f
C9218 VDD.n2637 VSS 0.00226f
C9219 VDD.t307 VSS 7.62e-19
C9220 VDD.t128 VSS 5.72e-19
C9221 VDD.n2638 VSS 0.0014f
C9222 VDD.t127 VSS 0.00579f
C9223 VDD.n2639 VSS 0.00762f
C9224 VDD.n2640 VSS 0.00111f
C9225 VDD.n2641 VSS 0.00203f
C9226 VDD.n2642 VSS 0.00252f
C9227 VDD.n2643 VSS 0.00263f
C9228 VDD.n2644 VSS 0.00136f
C9229 VDD.n2645 VSS 5.97e-19
C9230 VDD.n2646 VSS 5.16e-19
C9231 VDD.n2647 VSS 0.00158f
C9232 VDD.n2648 VSS 5.79e-19
C9233 VDD.n2649 VSS 0.00154f
C9234 VDD.n2650 VSS 9.31e-19
C9235 VDD.t724 VSS 0.00578f
C9236 VDD.n2651 VSS 0.00528f
C9237 VDD.n2652 VSS 0.00109f
C9238 VDD.n2653 VSS 1.72e-19
C9239 VDD.n2654 VSS 2.85e-19
C9240 VDD.n2655 VSS 9.31e-19
C9241 VDD.n2656 VSS 2.18e-19
C9242 VDD.t549 VSS 0.00578f
C9243 VDD.n2657 VSS 0.00578f
C9244 VDD.n2658 VSS 0.00109f
C9245 VDD.n2659 VSS 0.00149f
C9246 VDD.n2660 VSS 0.00251f
C9247 VDD.n2661 VSS 0.00132f
C9248 VDD.n2662 VSS 4.35e-19
C9249 VDD.n2663 VSS 5.33e-19
C9250 VDD.n2664 VSS 3.36e-19
C9251 VDD.n2665 VSS 8.1e-19
C9252 VDD.n2666 VSS 0.00148f
C9253 VDD.n2667 VSS 0.00123f
C9254 VDD.n2668 VSS 0.00158f
C9255 VDD.n2669 VSS 6.8e-19
C9256 VDD.n2670 VSS 4.3e-19
C9257 VDD.t160 VSS 0.00578f
C9258 VDD.n2671 VSS 0.00154f
C9259 VDD.n2672 VSS 2.85e-19
C9260 VDD.t671 VSS 0.00578f
C9261 VDD.n2673 VSS 0.00854f
C9262 VDD.n2674 VSS 0.00111f
C9263 VDD.n2675 VSS 0.002f
C9264 VDD.t672 VSS 0.00141f
C9265 VDD.n2676 VSS 0.00295f
C9266 VDD.n2677 VSS 2.1e-19
C9267 VDD.n2678 VSS 5.7e-19
C9268 VDD.n2679 VSS 4.52e-19
C9269 VDD.n2680 VSS 0.00158f
C9270 VDD.n2681 VSS 0.00158f
C9271 VDD.n2682 VSS 4.9e-19
C9272 VDD.n2683 VSS 0.00693f
C9273 VDD.n2684 VSS 0.0117f
C9274 VDD.n2685 VSS 0.00109f
C9275 VDD.n2686 VSS 0.00157f
C9276 VDD.n2687 VSS 0.0117f
C9277 VDD.n2688 VSS 0.00109f
C9278 VDD.n2689 VSS 0.00157f
C9279 VDD.n2690 VSS 0.0117f
C9280 VDD.n2691 VSS 0.00109f
C9281 VDD.n2692 VSS 0.00157f
C9282 VDD.n2693 VSS 0.0117f
C9283 VDD.n2694 VSS 0.00109f
C9284 VDD.n2695 VSS 0.00179f
C9285 VDD.n2696 VSS 0.0039f
C9286 VDD.n2697 VSS 0.00154f
C9287 VDD.n2698 VSS 9.31e-19
C9288 VDD.t396 VSS 0.00584f
C9289 VDD.n2699 VSS 0.00597f
C9290 VDD.n2700 VSS 0.00109f
C9291 VDD.n2701 VSS 1.72e-19
C9292 VDD.n2702 VSS 2.85e-19
C9293 VDD.t397 VSS 4.25e-19
C9294 VDD.t591 VSS 5.42e-19
C9295 VDD.n2703 VSS 0.00111f
C9296 VDD.n2704 VSS 0.00249f
C9297 VDD.n2705 VSS 4.66e-19
C9298 VDD.n2706 VSS 4.69e-19
C9299 VDD.t453 VSS 0.00546f
C9300 VDD.n2707 VSS 0.00673f
C9301 VDD.n2708 VSS 0.00109f
C9302 VDD.n2709 VSS 0.00186f
C9303 VDD.n2710 VSS 0.00308f
C9304 VDD.t590 VSS 0.00495f
C9305 VDD.n2711 VSS 0.0061f
C9306 VDD.n2712 VSS 0.00109f
C9307 VDD.n2713 VSS 0.0014f
C9308 VDD.n2714 VSS 0.00248f
C9309 VDD.n2715 VSS 0.00107f
C9310 VDD.n2716 VSS 4.35e-19
C9311 VDD.n2717 VSS 6.22e-19
C9312 VDD.n2718 VSS 3.36e-19
C9313 VDD.n2719 VSS 8.1e-19
C9314 VDD.n2720 VSS 0.00148f
C9315 VDD.n2721 VSS 0.00144f
C9316 VDD.n2722 VSS 0.00148f
C9317 VDD.n2723 VSS 8.1e-19
C9318 VDD.n2724 VSS 0.00157f
C9319 VDD.n2725 VSS 0.00727f
C9320 VDD.n2726 VSS 0.00149f
C9321 VDD.n2727 VSS 5.46e-19
C9322 VDD.n2728 VSS 5.66e-19
C9323 VDD.n2729 VSS 0.0117f
C9324 VDD.n2730 VSS 0.00109f
C9325 VDD.n2731 VSS 0.00183f
C9326 VDD.n2732 VSS 0.0026f
C9327 VDD.n2733 VSS 0.00129f
C9328 VDD.n2734 VSS 0.00181f
C9329 VDD.t374 VSS 7.73e-19
C9330 VDD.t274 VSS 2.51e-19
C9331 VDD.n2735 VSS 0.00395f
C9332 VDD.n2736 VSS 0.00308f
C9333 VDD.n2737 VSS 9.11e-19
C9334 VDD.n2738 VSS 0.0117f
C9335 VDD.n2739 VSS 0.00109f
C9336 VDD.n2740 VSS 0.00157f
C9337 VDD.n2741 VSS 0.0117f
C9338 VDD.n2742 VSS 0.00109f
C9339 VDD.n2743 VSS 0.00157f
C9340 VDD.n2744 VSS 0.0117f
C9341 VDD.n2745 VSS 0.00109f
C9342 VDD.n2746 VSS 0.00157f
C9343 VDD.n2747 VSS 0.0117f
C9344 VDD.n2748 VSS 0.00109f
C9345 VDD.n2749 VSS 0.00157f
C9346 VDD.n2750 VSS 0.0117f
C9347 VDD.n2751 VSS 0.00109f
C9348 VDD.n2752 VSS 0.00157f
C9349 VDD.n2753 VSS 0.0117f
C9350 VDD.n2754 VSS 0.00109f
C9351 VDD.n2755 VSS 0.00186f
C9352 VDD.n2756 VSS 0.00226f
C9353 VDD.n2757 VSS 0.00346f
C9354 VDD.n2758 VSS 0.0246f
C9355 VDD.n2759 VSS 0.00615f
C9356 VDD.n2760 VSS 0.00158f
C9357 VDD.n2761 VSS 5.41e-19
C9358 VDD.n2762 VSS 5.71e-19
C9359 VDD.n2763 VSS 3.36e-19
C9360 VDD.n2764 VSS 8.1e-19
C9361 VDD.n2765 VSS 0.00148f
C9362 VDD.n2766 VSS 0.00158f
C9363 VDD.n2767 VSS 8.1e-19
C9364 VDD.n2768 VSS 0.00144f
C9365 VDD.n2769 VSS 0.00148f
C9366 VDD.n2770 VSS 0.00615f
C9367 VDD.n2771 VSS 0.00148f
C9368 VDD.n2772 VSS 0.00158f
C9369 VDD.n2773 VSS 6.05e-19
C9370 VDD.n2774 VSS 2.53e-19
C9371 VDD.t486 VSS 0.00394f
C9372 VDD.n2775 VSS 0.00642f
C9373 VDD.n2776 VSS 9.31e-19
C9374 VDD.t683 VSS 0.00578f
C9375 VDD.n2777 VSS 0.00528f
C9376 VDD.n2778 VSS 0.00109f
C9377 VDD.t684 VSS 9.42e-19
C9378 VDD.t678 VSS 9.42e-19
C9379 VDD.n2779 VSS 0.00214f
C9380 VDD.n2780 VSS 0.00258f
C9381 VDD.n2781 VSS 0.00119f
C9382 VDD.n2782 VSS 0.00233f
C9383 VDD.t677 VSS 0.00578f
C9384 VDD.n2783 VSS 0.00528f
C9385 VDD.n2784 VSS 0.00109f
C9386 VDD.n2785 VSS 0.00149f
C9387 VDD.n2786 VSS 0.00246f
C9388 VDD.n2787 VSS 0.00101f
C9389 VDD.n2788 VSS 6.55e-19
C9390 VDD.n2789 VSS 4.52e-19
C9391 VDD.n2790 VSS 0.00158f
C9392 VDD.n2791 VSS 0.00149f
C9393 VDD.n2792 VSS 0.00943f
C9394 VDD.n2793 VSS 0.00725f
C9395 VDD.n2794 VSS 0.252f
C9396 VDD.n2795 VSS 0.0155f
C9397 VDD.n2796 VSS 0.00158f
C9398 VDD.n2797 VSS 0.00149f
C9399 VDD.n2798 VSS 5.92e-19
C9400 VDD.n2799 VSS 0.00154f
C9401 VDD.n2800 VSS 4.15e-19
C9402 VDD.t154 VSS 0.00578f
C9403 VDD.n2801 VSS 0.00528f
C9404 VDD.n2802 VSS 0.00109f
C9405 VDD.n2803 VSS 1.72e-19
C9406 VDD.n2804 VSS 2.85e-19
C9407 VDD.n2805 VSS 8.8e-19
C9408 VDD.n2806 VSS 6.37e-19
C9409 VDD.n2807 VSS 4.26e-19
C9410 VDD.n2808 VSS 0.00158f
C9411 VDD.n2809 VSS 0.0106f
C9412 VDD.n2810 VSS 0.00158f
C9413 VDD.n2811 VSS 0.00149f
C9414 VDD.n2812 VSS 5.28e-19
C9415 VDD.n2813 VSS 9.31e-19
C9416 VDD.t654 VSS 0.00578f
C9417 VDD.n2814 VSS 0.00528f
C9418 VDD.n2815 VSS 0.00109f
C9419 VDD.t655 VSS 9.42e-19
C9420 VDD.t659 VSS 9.42e-19
C9421 VDD.n2816 VSS 0.00214f
C9422 VDD.n2817 VSS 0.00258f
C9423 VDD.n2818 VSS 9.92e-19
C9424 VDD.n2819 VSS 0.00258f
C9425 VDD.t658 VSS 0.00578f
C9426 VDD.t652 VSS 0.00578f
C9427 VDD.n2820 VSS 0.00528f
C9428 VDD.n2821 VSS 0.00109f
C9429 VDD.n2822 VSS 0.0017f
C9430 VDD.n2823 VSS 0.00261f
C9431 VDD.n2824 VSS 0.00132f
C9432 VDD.n2825 VSS 5.28e-19
C9433 VDD.n2826 VSS 5.79e-19
C9434 VDD.n2827 VSS 0.00158f
C9435 VDD.n2828 VSS 0.0121f
C9436 VDD.n2829 VSS 0.0106f
C9437 VDD.n2830 VSS 0.00335f
C9438 VDD.n2831 VSS 0.00149f
C9439 VDD.n2832 VSS 8.1e-19
C9440 VDD.n2833 VSS 3.36e-19
C9441 VDD.n2834 VSS 4.35e-19
C9442 VDD.t653 VSS 0.00374f
C9443 VDD.n2835 VSS 0.00362f
C9444 VDD.n2836 VSS 6.07e-20
C9445 VDD.n2837 VSS 2.18e-19
C9446 VDD.n2838 VSS 2.68e-19
C9447 VDD.n2839 VSS 2.85e-19
C9448 VDD.n2840 VSS 1.72e-19
C9449 VDD.n2841 VSS 0.00109f
C9450 VDD.n2842 VSS 0.00402f
C9451 VDD.n2843 VSS 0.00955f
C9452 VDD.n2844 VSS 0.00109f
C9453 VDD.n2845 VSS 2.53e-19
C9454 VDD.t153 VSS 0.00394f
C9455 VDD.n2846 VSS 0.00648f
C9456 VDD.n2847 VSS 7.89e-19
C9457 VDD.n2848 VSS 0.00214f
C9458 VDD.n2849 VSS 0.00154f
C9459 VDD.t152 VSS 0.00578f
C9460 VDD.n2850 VSS 0.00528f
C9461 VDD.n2851 VSS 0.00109f
C9462 VDD.n2852 VSS 1.72e-19
C9463 VDD.n2853 VSS 2.85e-19
C9464 VDD.n2854 VSS 7.79e-19
C9465 VDD.n2855 VSS 3.68e-19
C9466 VDD.t157 VSS 9.42e-19
C9467 VDD.t155 VSS 9.42e-19
C9468 VDD.n2856 VSS 0.00224f
C9469 VDD.t156 VSS 0.00578f
C9470 VDD.n2857 VSS 0.00528f
C9471 VDD.n2858 VSS 0.00111f
C9472 VDD.n2859 VSS 0.00193f
C9473 VDD.n2860 VSS 0.00383f
C9474 VDD.n2861 VSS 0.0025f
C9475 VDD.n2862 VSS 0.00117f
C9476 VDD.n2863 VSS 4.35e-19
C9477 VDD.n2864 VSS 5.79e-19
C9478 VDD.n2865 VSS 3.36e-19
C9479 VDD.n2866 VSS 8.1e-19
C9480 VDD.n2867 VSS 0.00335f
C9481 VDD.n2868 VSS 0.00949f
C9482 VDD.n2869 VSS 0.00949f
C9483 VDD.n2870 VSS 0.0155f
C9484 VDD.n2871 VSS 0.00335f
C9485 VDD.n2872 VSS 0.00149f
C9486 VDD.n2873 VSS 8.1e-19
C9487 VDD.n2874 VSS 6.8e-19
C9488 VDD.n2875 VSS 3.36e-19
C9489 VDD.n2876 VSS 4.35e-19
C9490 VDD.n2877 VSS 9.04e-19
C9491 VDD.t159 VSS 9.42e-19
C9492 VDD.t262 VSS 9.42e-19
C9493 VDD.n2878 VSS 0.00215f
C9494 VDD.n2879 VSS 0.00319f
C9495 VDD.t158 VSS 0.00578f
C9496 VDD.t261 VSS 0.00578f
C9497 VDD.n2880 VSS 0.00528f
C9498 VDD.n2881 VSS 0.00109f
C9499 VDD.n2882 VSS 9.82e-19
C9500 VDD.n2883 VSS 0.0024f
C9501 VDD.n2884 VSS 0.00181f
C9502 VDD.n2885 VSS 0.00186f
C9503 VDD.n2886 VSS 0.00109f
C9504 VDD.n2887 VSS 0.00402f
C9505 VDD.n2888 VSS 0.00779f
C9506 VDD.n2889 VSS 0.00109f
C9507 VDD.n2890 VSS 0.00153f
C9508 VDD.n2891 VSS 0.00178f
C9509 VDD.n2892 VSS 0.00117f
C9510 VDD.n2893 VSS 9.04e-19
C9511 VDD.n2894 VSS 4.26e-19
C9512 VDD.n2895 VSS 6.8e-19
C9513 VDD.n2896 VSS 0.00158f
C9514 VDD.n2897 VSS 0.00725f
C9515 VDD.n2898 VSS 0.00149f
C9516 VDD.n2899 VSS 8.23e-19
C9517 VDD.n2900 VSS 0.00144f
C9518 VDD.n2901 VSS 0.00157f
C9519 VDD.n2902 VSS 0.00726f
C9520 VDD.n2903 VSS 0.00726f
C9521 VDD.n2904 VSS 0.037f
C9522 VDD.n2905 VSS 0.00149f
C9523 VDD.n2906 VSS 8.11e-19
C9524 VDD.n2907 VSS 3.36e-19
C9525 VDD.n2908 VSS 4.35e-19
C9526 VDD.n2909 VSS 9.31e-19
C9527 VDD.n2910 VSS 6.37e-19
C9528 VDD.t416 VSS 0.00349f
C9529 VDD.n2911 VSS 0.00294f
C9530 VDD.n2912 VSS 1.42e-19
C9531 VDD.t415 VSS 0.00616f
C9532 VDD.n2913 VSS 0.00867f
C9533 VDD.n2914 VSS 0.00109f
C9534 VDD.n2915 VSS 1.72e-19
C9535 VDD.n2916 VSS 2.85e-19
C9536 VDD.n2917 VSS 0.00154f
C9537 VDD.n2918 VSS 0.0176f
C9538 VDD.n2919 VSS 0.00322f
C9539 VDD.n2920 VSS 0.0264f
C9540 VDD.n2921 VSS 0.00408f
C9541 VDD.n2922 VSS 0.00109f
C9542 VDD.n2923 VSS 0.00153f
C9543 VDD.n2924 VSS 0.00164f
C9544 VDD.n2925 VSS 0.00154f
C9545 VDD.n2926 VSS 2.85e-19
C9546 VDD.t38 VSS 0.00578f
C9547 VDD.t326 VSS 0.00578f
C9548 VDD.n2927 VSS 0.00553f
C9549 VDD.n2928 VSS 0.00111f
C9550 VDD.n2929 VSS 0.00199f
C9551 VDD.t39 VSS 7.99e-19
C9552 VDD.t327 VSS 7.99e-19
C9553 VDD.n2930 VSS 0.00191f
C9554 VDD.n2931 VSS 0.00352f
C9555 VDD.n2932 VSS 1.96e-19
C9556 VDD.n2933 VSS 3.68e-19
C9557 VDD.n2934 VSS 4.35e-19
C9558 VDD.n2935 VSS 5.16e-19
C9559 VDD.n2936 VSS 3.36e-19
C9560 VDD.n2937 VSS 8.1e-19
C9561 VDD.n2938 VSS 0.00335f
C9562 VDD.n2939 VSS 0.0326f
C9563 VDD.n2940 VSS 0.297f
C9564 VDD.n2941 VSS 0.00676f
C9565 VDD.n2942 VSS 0.00158f
C9566 VDD.n2943 VSS 5.41e-19
C9567 VDD.t437 VSS 0.00578f
C9568 VDD.n2944 VSS 0.00528f
C9569 VDD.n2945 VSS 0.00109f
C9570 VDD.n2946 VSS 0.00141f
C9571 VDD.n2947 VSS 0.0024f
C9572 VDD.t438 VSS 9.42e-19
C9573 VDD.t426 VSS 9.42e-19
C9574 VDD.n2948 VSS 0.00214f
C9575 VDD.n2949 VSS 0.00258f
C9576 VDD.t425 VSS 0.00578f
C9577 VDD.n2950 VSS 0.00528f
C9578 VDD.n2951 VSS 0.00109f
C9579 VDD.n2952 VSS 0.0012f
C9580 VDD.n2953 VSS 0.0026f
C9581 VDD.n2954 VSS 0.00129f
C9582 VDD.t436 VSS 9.42e-19
C9583 VDD.t422 VSS 9.42e-19
C9584 VDD.n2955 VSS 0.00214f
C9585 VDD.n2956 VSS 0.00243f
C9586 VDD.t421 VSS 0.00553f
C9587 VDD.n2957 VSS 0.00528f
C9588 VDD.n2958 VSS 0.00109f
C9589 VDD.n2959 VSS 0.0014f
C9590 VDD.n2960 VSS 0.00285f
C9591 VDD.n2961 VSS 0.00154f
C9592 VDD.n2962 VSS 4.66e-19
C9593 VDD.t435 VSS 0.00553f
C9594 VDD.n2963 VSS 0.00528f
C9595 VDD.n2964 VSS 0.00109f
C9596 VDD.n2965 VSS 1.72e-19
C9597 VDD.n2966 VSS 2.85e-19
C9598 VDD.n2967 VSS 9.31e-19
C9599 VDD.n2968 VSS 2.51e-19
C9600 VDD.n2969 VSS 4.35e-19
C9601 VDD.n2970 VSS 5.66e-19
C9602 VDD.n2971 VSS 3.36e-19
C9603 VDD.n2972 VSS 0.00149f
C9604 VDD.n2973 VSS 8.1e-19
C9605 VDD.n2974 VSS 0.00335f
C9606 VDD.n2975 VSS 0.0138f
C9607 VDD.n2976 VSS 0.0138f
C9608 VDD.n2977 VSS 0.00158f
C9609 VDD.n2978 VSS 5.41e-19
C9610 VDD.t432 VSS 9.42e-19
C9611 VDD.t418 VSS 9.42e-19
C9612 VDD.n2979 VSS 0.00214f
C9613 VDD.n2980 VSS 0.00256f
C9614 VDD.t431 VSS 0.00578f
C9615 VDD.n2981 VSS 0.00528f
C9616 VDD.n2982 VSS 0.00109f
C9617 VDD.n2983 VSS 0.00123f
C9618 VDD.n2984 VSS 0.00261f
C9619 VDD.n2985 VSS 0.00131f
C9620 VDD.t430 VSS 9.42e-19
C9621 VDD.t414 VSS 9.42e-19
C9622 VDD.n2986 VSS 0.00214f
C9623 VDD.n2987 VSS 0.00258f
C9624 VDD.t429 VSS 0.00578f
C9625 VDD.n2988 VSS 0.00528f
C9626 VDD.n2989 VSS 0.00109f
C9627 VDD.n2990 VSS 9.21e-19
C9628 VDD.n2991 VSS 0.00283f
C9629 VDD.n2992 VSS 0.00154f
C9630 VDD.n2993 VSS 9.31e-19
C9631 VDD.t417 VSS 0.00578f
C9632 VDD.n2994 VSS 0.00528f
C9633 VDD.n2995 VSS 0.00109f
C9634 VDD.n2996 VSS 1.72e-19
C9635 VDD.n2997 VSS 2.85e-19
C9636 VDD.n2998 VSS 6.27e-19
C9637 VDD.n2999 VSS 2.35e-19
C9638 VDD.n3000 VSS 4.35e-19
C9639 VDD.n3001 VSS 5.66e-19
C9640 VDD.n3002 VSS 3.36e-19
C9641 VDD.n3003 VSS 0.00149f
C9642 VDD.n3004 VSS 8.1e-19
C9643 VDD.n3005 VSS 0.00335f
C9644 VDD.n3006 VSS 0.0136f
C9645 VDD.n3007 VSS 0.0136f
C9646 VDD.n3008 VSS 0.00158f
C9647 VDD.n3009 VSS 5.54e-19
C9648 VDD.n3010 VSS 5.54e-19
C9649 VDD.t413 VSS 0.00578f
C9650 VDD.n3011 VSS 0.00528f
C9651 VDD.n3012 VSS 0.00109f
C9652 VDD.n3013 VSS 0.00169f
C9653 VDD.n3014 VSS 0.0026f
C9654 VDD.n3015 VSS 0.00127f
C9655 VDD.t409 VSS 0.00578f
C9656 VDD.n3016 VSS 0.00528f
C9657 VDD.n3017 VSS 0.00109f
C9658 VDD.n3018 VSS 0.00154f
C9659 VDD.n3019 VSS 0.00263f
C9660 VDD.n3020 VSS 0.00154f
C9661 VDD.n3021 VSS 9.31e-19
C9662 VDD.t411 VSS 0.00578f
C9663 VDD.t427 VSS 0.00578f
C9664 VDD.n3022 VSS 0.00528f
C9665 VDD.n3023 VSS 0.00109f
C9666 VDD.n3024 VSS 1.62e-19
C9667 VDD.n3025 VSS 2.85e-19
C9668 VDD.t412 VSS 9.42e-19
C9669 VDD.t428 VSS 9.42e-19
C9670 VDD.n3026 VSS 0.00214f
C9671 VDD.n3027 VSS 0.00168f
C9672 VDD.n3028 VSS 9.11e-19
C9673 VDD.n3029 VSS 2.68e-19
C9674 VDD.n3030 VSS 4.35e-19
C9675 VDD.n3031 VSS 3.36e-19
C9676 VDD.n3032 VSS 0.00149f
C9677 VDD.n3033 VSS 8.1e-19
C9678 VDD.n3034 VSS 0.00335f
C9679 VDD.n3035 VSS 0.0104f
C9680 VDD.n3036 VSS 0.0104f
C9681 VDD.n3037 VSS 0.00158f
C9682 VDD.n3038 VSS 0.00149f
C9683 VDD.n3039 VSS 5.54e-19
C9684 VDD.n3040 VSS 0.00154f
C9685 VDD.t410 VSS 9.42e-19
C9686 VDD.t424 VSS 9.42e-19
C9687 VDD.n3041 VSS 0.00214f
C9688 VDD.n3042 VSS 0.00244f
C9689 VDD.n3043 VSS 1.82e-19
C9690 VDD.t423 VSS 0.00578f
C9691 VDD.n3044 VSS 0.00528f
C9692 VDD.n3045 VSS 0.00109f
C9693 VDD.n3046 VSS 1.72e-19
C9694 VDD.n3047 VSS 2.85e-19
C9695 VDD.n3048 VSS 9.31e-19
C9696 VDD.n3049 VSS 2.85e-19
C9697 VDD.t433 VSS 0.00578f
C9698 VDD.n3050 VSS 0.00528f
C9699 VDD.n3051 VSS 0.00109f
C9700 VDD.n3052 VSS 0.00148f
C9701 VDD.n3053 VSS 0.00251f
C9702 VDD.n3054 VSS 0.00126f
C9703 VDD.n3055 VSS 4.35e-19
C9704 VDD.n3056 VSS 5.54e-19
C9705 VDD.n3057 VSS 3.36e-19
C9706 VDD.n3058 VSS 8.1e-19
C9707 VDD.n3059 VSS 0.00335f
C9708 VDD.n3060 VSS 0.00955f
C9709 VDD.n3061 VSS 0.00955f
C9710 VDD.n3062 VSS 0.00158f
C9711 VDD.n3063 VSS 0.00149f
C9712 VDD.n3064 VSS 4.52e-19
C9713 VDD.n3065 VSS 0.00154f
C9714 VDD.t434 VSS 9.42e-19
C9715 VDD.t420 VSS 9.42e-19
C9716 VDD.n3066 VSS 0.00214f
C9717 VDD.n3067 VSS 0.00254f
C9718 VDD.n3068 VSS 3.44e-19
C9719 VDD.t419 VSS 0.00578f
C9720 VDD.n3069 VSS 0.00528f
C9721 VDD.n3070 VSS 0.00109f
C9722 VDD.n3071 VSS 1.72e-19
C9723 VDD.n3072 VSS 2.85e-19
C9724 VDD.n3073 VSS 9.31e-19
C9725 VDD.n3074 VSS 5.7e-19
C9726 VDD.n3075 VSS 0.00154f
C9727 VDD.t679 VSS 0.00578f
C9728 VDD.n3076 VSS 0.00528f
C9729 VDD.n3077 VSS 0.00109f
C9730 VDD.n3078 VSS 0.00144f
C9731 VDD.n3079 VSS 0.00229f
C9732 VDD.t440 VSS 9.42e-19
C9733 VDD.t680 VSS 9.42e-19
C9734 VDD.n3080 VSS 0.00214f
C9735 VDD.n3081 VSS 0.00258f
C9736 VDD.t439 VSS 0.0106f
C9737 VDD.n3082 VSS 0.00109f
C9738 VDD.n3083 VSS 0.00122f
C9739 VDD.n3084 VSS 0.00243f
C9740 VDD.n3085 VSS 9.71e-19
C9741 VDD.n3086 VSS 4.35e-19
C9742 VDD.n3087 VSS 6.55e-19
C9743 VDD.n3088 VSS 3.36e-19
C9744 VDD.n3089 VSS 8.1e-19
C9745 VDD.n3090 VSS 0.00335f
C9746 VDD.n3091 VSS 0.00921f
C9747 VDD.n3092 VSS 0.00921f
C9748 VDD.n3093 VSS 0.00158f
C9749 VDD.n3094 VSS 0.00144f
C9750 VDD.n3095 VSS 0.00148f
C9751 VDD.n3096 VSS 8.1e-19
C9752 VDD.n3097 VSS 0.00335f
C9753 VDD.n3098 VSS 0.00944f
C9754 VDD.n3099 VSS 0.00944f
C9755 VDD.n3100 VSS 0.00335f
C9756 VDD.n3101 VSS 8.1e-19
C9757 VDD.n3102 VSS 3.36e-19
C9758 VDD.n3103 VSS 4.35e-19
C9759 VDD.n3104 VSS 9.31e-19
C9760 VDD.n3105 VSS 5.36e-19
C9761 VDD.t681 VSS 0.00578f
C9762 VDD.n3106 VSS 0.00528f
C9763 VDD.n3107 VSS 0.00109f
C9764 VDD.t682 VSS 9.42e-19
C9765 VDD.t688 VSS 9.42e-19
C9766 VDD.n3108 VSS 0.00214f
C9767 VDD.n3109 VSS 0.00252f
C9768 VDD.n3110 VSS 1.01e-19
C9769 VDD.n3111 VSS 1.72e-19
C9770 VDD.n3112 VSS 2.85e-19
C9771 VDD.n3113 VSS 0.00154f
C9772 VDD.t687 VSS 0.00578f
C9773 VDD.t685 VSS 0.00578f
C9774 VDD.n3114 VSS 0.00528f
C9775 VDD.n3115 VSS 0.00109f
C9776 VDD.n3116 VSS 0.0017f
C9777 VDD.n3117 VSS 0.00251f
C9778 VDD.n3118 VSS 0.00131f
C9779 VDD.n3119 VSS 4.35e-19
C9780 VDD.t686 VSS 0.00374f
C9781 VDD.n3120 VSS 0.00362f
C9782 VDD.n3121 VSS 6.07e-20
C9783 VDD.n3122 VSS 2.35e-19
C9784 VDD.n3123 VSS 2.68e-19
C9785 VDD.n3124 VSS 2.85e-19
C9786 VDD.n3125 VSS 1.72e-19
C9787 VDD.n3126 VSS 0.00109f
C9788 VDD.n3127 VSS 0.00402f
C9789 VDD.n3128 VSS 0.00955f
C9790 VDD.n3129 VSS 0.00109f
C9791 VDD.n3130 VSS 7.89e-19
C9792 VDD.n3131 VSS 0.00204f
C9793 VDD.n3132 VSS 0.00154f
C9794 VDD.t485 VSS 0.00578f
C9795 VDD.n3133 VSS 0.00528f
C9796 VDD.n3134 VSS 0.00109f
C9797 VDD.n3135 VSS 1.72e-19
C9798 VDD.n3136 VSS 2.85e-19
C9799 VDD.n3137 VSS 7.79e-19
C9800 VDD.n3138 VSS 1.68e-19
C9801 VDD.t484 VSS 9.42e-19
C9802 VDD.t488 VSS 9.42e-19
C9803 VDD.n3139 VSS 0.00224f
C9804 VDD.t483 VSS 0.00578f
C9805 VDD.n3140 VSS 0.00528f
C9806 VDD.n3141 VSS 0.00111f
C9807 VDD.n3142 VSS 0.00188f
C9808 VDD.n3143 VSS 0.00383f
C9809 VDD.n3144 VSS 0.00241f
C9810 VDD.n3145 VSS 0.00137f
C9811 VDD.n3146 VSS 4.35e-19
C9812 VDD.n3147 VSS 5.07e-19
C9813 VDD.n3148 VSS 3.36e-19
C9814 VDD.n3149 VSS 8.1e-19
C9815 VDD.n3150 VSS 0.00148f
C9816 VDD.n3151 VSS 5.72e-19
C9817 VDD.n3152 VSS 0.00154f
C9818 VDD.n3153 VSS 4.15e-19
C9819 VDD.t487 VSS 0.00578f
C9820 VDD.n3154 VSS 0.00528f
C9821 VDD.n3155 VSS 0.00109f
C9822 VDD.n3156 VSS 1.72e-19
C9823 VDD.n3157 VSS 2.85e-19
C9824 VDD.n3158 VSS 8.8e-19
C9825 VDD.n3159 VSS 2.68e-19
C9826 VDD.n3160 VSS 7.71e-19
C9827 VDD.n3161 VSS 1.72e-19
C9828 VDD.n3162 VSS 0.00408f
C9829 VDD.n3163 VSS 0.00109f
C9830 VDD.n3164 VSS 1.72e-19
C9831 VDD.n3165 VSS 7.71e-19
C9832 VDD.n3166 VSS 2.85e-19
C9833 VDD.n3167 VSS 5.97e-19
C9834 VDD.n3168 VSS 5.19e-19
C9835 VDD.n3169 VSS 6.43e-19
C9836 VDD.n3170 VSS 4.69e-19
C9837 VDD.n3171 VSS 0.00158f
C9838 VDD.n3172 VSS 8.1e-19
C9839 VDD.n3173 VSS 3.36e-19
C9840 VDD.n3174 VSS 4.35e-19
C9841 VDD.n3175 VSS 0.00102f
C9842 VDD.t13 VSS 7.99e-19
C9843 VDD.t574 VSS 7.99e-19
C9844 VDD.n3176 VSS 0.00194f
C9845 VDD.t12 VSS 0.00578f
C9846 VDD.t573 VSS 0.00578f
C9847 VDD.n3177 VSS 0.00553f
C9848 VDD.n3178 VSS 0.00111f
C9849 VDD.n3179 VSS 0.00191f
C9850 VDD.n3180 VSS 0.00366f
C9851 VDD.n3181 VSS 0.00246f
C9852 VDD.n3182 VSS 0.00231f
C9853 VDD.n3183 VSS 0.00137f
C9854 VDD.n3184 VSS 0.00109f
C9855 VDD.n3185 VSS 0.00779f
C9856 VDD.n3186 VSS 0.00402f
C9857 VDD.n3187 VSS 0.00109f
C9858 VDD.n3188 VSS 0.00109f
C9859 VDD.n3189 VSS 0.00226f
C9860 VDD.t490 VSS 9.42e-19
C9861 VDD.t342 VSS 9.42e-19
C9862 VDD.n3190 VSS 0.00215f
C9863 VDD.n3191 VSS 0.0033f
C9864 VDD.t489 VSS 0.00578f
C9865 VDD.t341 VSS 0.00578f
C9866 VDD.n3192 VSS 0.00528f
C9867 VDD.n3193 VSS 0.00109f
C9868 VDD.n3194 VSS 9.82e-19
C9869 VDD.n3195 VSS 0.00258f
C9870 VDD.n3196 VSS 0.00127f
C9871 VDD.n3197 VSS 4.35e-19
C9872 VDD.n3198 VSS 5.41e-19
C9873 VDD.n3199 VSS 3.36e-19
C9874 VDD.n3200 VSS 0.00149f
C9875 VDD.n3201 VSS 8.1e-19
C9876 VDD.n3202 VSS 0.00157f
C9877 VDD.n3203 VSS 0.00615f
C9878 VDD.n3204 VSS 0.00615f
C9879 VDD.n3205 VSS 0.0084f
C9880 VDD.n3206 VSS 0.224f
C9881 VDD.n3207 VSS 0.214f
C9882 VDD.n3208 VSS 6.15e-19
C9883 VDD.n3209 VSS 0.00574f
C9884 VDD.n3210 VSS 0.00158f
C9885 VDD.n3211 VSS 4.26e-19
C9886 VDD.n3212 VSS 2.84e-19
C9887 VDD.n3213 VSS 0.00154f
C9888 VDD.t743 VSS 7.73e-19
C9889 VDD.t245 VSS 2.51e-19
C9890 VDD.n3214 VSS 0.00395f
C9891 VDD.n3215 VSS 0.00308f
C9892 VDD.n3216 VSS 0.00273f
C9893 VDD.n3217 VSS 9.51e-19
C9894 VDD.n3218 VSS 0.00109f
C9895 VDD.n3219 VSS 0.00692f
C9896 VDD.t244 VSS 0.00406f
C9897 VDD.n3220 VSS 0.0127f
C9898 VDD.n3221 VSS 0.00184f
C9899 VDD.n3222 VSS 3.68e-19
C9900 VDD.n3223 VSS 2.68e-19
C9901 VDD.n3224 VSS 5.03e-19
C9902 VDD.n3225 VSS 4.56e-19
C9903 VDD.n3226 VSS 2.84e-19
C9904 VDD.n3227 VSS 8.1e-19
C9905 VDD.n3228 VSS 0.00148f
C9906 VDD.n3229 VSS 0.00594f
C9907 VDD.n3230 VSS 0.00158f
C9908 VDD.n3231 VSS 5.03e-19
C9909 VDD.n3232 VSS 6.09e-19
C9910 VDD.n3233 VSS 3.36e-19
C9911 VDD.n3234 VSS 8.1e-19
C9912 VDD.n3235 VSS 0.00148f
C9913 VDD.n3236 VSS 0.00158f
C9914 VDD.n3237 VSS 4.64e-19
C9915 VDD.n3238 VSS 6.47e-19
C9916 VDD.n3239 VSS 0.00154f
C9917 VDD.n3240 VSS 2.85e-19
C9918 VDD.t70 VSS 0.00578f
C9919 VDD.n3241 VSS 0.00854f
C9920 VDD.n3242 VSS 0.00111f
C9921 VDD.n3243 VSS 0.002f
C9922 VDD.t71 VSS 0.00141f
C9923 VDD.n3244 VSS 0.00295f
C9924 VDD.n3245 VSS 2.1e-19
C9925 VDD.n3246 VSS 5.19e-19
C9926 VDD.t551 VSS 6.03e-19
C9927 VDD.t737 VSS 6.03e-19
C9928 VDD.n3247 VSS 0.0013f
C9929 VDD.n3248 VSS 0.0027f
C9930 VDD.t550 VSS 0.00578f
C9931 VDD.n3249 VSS 0.00202f
C9932 VDD.n3250 VSS 0.00111f
C9933 VDD.n3251 VSS 0.00528f
C9934 VDD.t736 VSS 0.00578f
C9935 VDD.n3252 VSS 0.00106f
C9936 VDD.n3253 VSS 0.00151f
C9937 VDD.n3254 VSS 0.00183f
C9938 VDD.n3255 VSS 0.00308f
C9939 VDD.n3256 VSS 0.00905f
C9940 VDD.n3257 VSS 0.00109f
C9941 VDD.n3258 VSS 0.00118f
C9942 VDD.n3259 VSS 0.00246f
C9943 VDD.n3260 VSS 0.00102f
C9944 VDD.n3261 VSS 4.35e-19
C9945 VDD.n3262 VSS 3.36e-19
C9946 VDD.n3263 VSS 8.1e-19
C9947 VDD.n3264 VSS 0.00148f
C9948 VDD.n3265 VSS 0.00553f
C9949 VDD.n3266 VSS 0.00492f
C9950 VDD.n3267 VSS 6.15e-19
C9951 VDD.n3268 VSS 0.00123f
C9952 VDD.n3269 VSS 0.128f
C9953 VDD.n3270 VSS 0.127f
C9954 VDD.n3271 VSS 6.15e-19
C9955 VDD.n3272 VSS 0.00594f
C9956 VDD.n3273 VSS 0.00574f
C9957 VDD.n3274 VSS 0.00149f
C9958 VDD.n3275 VSS 4.31e-19
C9959 VDD.n3276 VSS 6.8e-19
C9960 VDD.t375 VSS 0.00584f
C9961 VDD.n3277 VSS 0.00597f
C9962 VDD.n3278 VSS 0.00109f
C9963 VDD.n3279 VSS 0.0014f
C9964 VDD.n3280 VSS 0.00265f
C9965 VDD.n3281 VSS 0.00139f
C9966 VDD.n3282 VSS 4.35e-19
C9967 VDD.t376 VSS 4.25e-19
C9968 VDD.t448 VSS 5.42e-19
C9969 VDD.n3283 VSS 0.00111f
C9970 VDD.n3284 VSS 0.00259f
C9971 VDD.t447 VSS 0.00495f
C9972 VDD.n3285 VSS 0.0061f
C9973 VDD.n3286 VSS 0.00109f
C9974 VDD.n3287 VSS 0.0014f
C9975 VDD.n3288 VSS 0.00169f
C9976 VDD.t178 VSS 0.00546f
C9977 VDD.n3289 VSS 0.00673f
C9978 VDD.n3290 VSS 0.00109f
C9979 VDD.n3291 VSS 0.00186f
C9980 VDD.n3292 VSS 0.00308f
C9981 VDD.n3293 VSS 0.0117f
C9982 VDD.n3294 VSS 0.00109f
C9983 VDD.n3295 VSS 0.00183f
C9984 VDD.n3296 VSS 0.00303f
C9985 VDD.n3297 VSS 0.00154f
C9986 VDD.n3298 VSS 9.31e-19
C9987 VDD.t558 VSS 0.00584f
C9988 VDD.n3299 VSS 0.00686f
C9989 VDD.n3300 VSS 0.00109f
C9990 VDD.n3301 VSS 1.72e-19
C9991 VDD.n3302 VSS 2.85e-19
C9992 VDD.n3303 VSS 9.31e-19
C9993 VDD.n3304 VSS 6.2e-19
C9994 VDD.t742 VSS 0.00584f
C9995 VDD.n3305 VSS 0.00654f
C9996 VDD.n3306 VSS 0.00109f
C9997 VDD.n3307 VSS 0.00172f
C9998 VDD.n3308 VSS 0.00241f
C9999 VDD.n3309 VSS 9.21e-19
C10000 VDD.n3310 VSS 4.35e-19
C10001 VDD.n3311 VSS 3.36e-19
C10002 VDD.n3312 VSS 8.1e-19
C10003 VDD.n3313 VSS 0.00157f
C10004 VDD.n3314 VSS 6.23e-19
C10005 VDD.n3315 VSS 0.00157f
C10006 VDD.n3316 VSS 8.1e-19
C10007 VDD.n3317 VSS 0.00148f
C10008 VDD.n3318 VSS 0.00144f
C10009 VDD.n3319 VSS 0.0109f
C10010 VDD.n3320 VSS 0.0094f
C10011 VDD.n3321 VSS 0.00109f
C10012 VDD.n3322 VSS 9.31e-19
C10013 VDD.n3323 VSS 0.0117f
C10014 VDD.n3324 VSS 0.00109f
C10015 VDD.n3325 VSS 0.00157f
C10016 VDD.n3326 VSS 0.0117f
C10017 VDD.n3327 VSS 0.00109f
C10018 VDD.n3328 VSS 0.0013f
C10019 VDD.n3329 VSS 9.41e-19
C10020 VDD.n3330 VSS 0.00231f
C10021 VDD.t32 VSS 0.00584f
C10022 VDD.n3331 VSS 0.0061f
C10023 VDD.n3332 VSS 0.00109f
C10024 VDD.n3333 VSS 4.66e-19
C10025 VDD.n3334 VSS 9.31e-19
C10026 VDD.n3335 VSS 0.00308f
C10027 VDD.t605 VSS 0.00584f
C10028 VDD.t10 VSS 0.00584f
C10029 VDD.n3336 VSS 0.00457f
C10030 VDD.n3337 VSS 0.00109f
C10031 VDD.n3338 VSS 9.31e-19
C10032 VDD.t11 VSS 5.42e-19
C10033 VDD.t33 VSS 4.25e-19
C10034 VDD.n3339 VSS 0.00111f
C10035 VDD.n3340 VSS 0.0022f
C10036 VDD.n3341 VSS 8.5e-19
C10037 VDD.n3342 VSS 0.00308f
C10038 VDD.n3343 VSS 0.00915f
C10039 VDD.n3344 VSS 0.00109f
C10040 VDD.n3345 VSS 9.31e-19
C10041 VDD.n3346 VSS 9.31e-19
C10042 VDD.n3347 VSS 0.00308f
C10043 VDD.n3348 VSS 0.0103f
C10044 VDD.n3349 VSS 0.00109f
C10045 VDD.n3350 VSS 9.31e-19
C10046 VDD.n3351 VSS 9.31e-19
C10047 VDD.n3352 VSS 0.00308f
C10048 VDD.t553 VSS 0.00584f
C10049 VDD.n3353 VSS 0.00654f
C10050 VDD.n3354 VSS 0.00109f
C10051 VDD.n3355 VSS 9.31e-19
C10052 VDD.n3356 VSS 9.31e-19
C10053 VDD.n3357 VSS 0.00308f
C10054 VDD.n3358 VSS 9.31e-19
C10055 VDD.n3359 VSS 0.00308f
C10056 VDD.t646 VSS 7.73e-19
C10057 VDD.t693 VSS 2.51e-19
C10058 VDD.n3360 VSS 0.00395f
C10059 VDD.n3361 VSS 0.00253f
C10060 VDD.t692 VSS 0.00584f
C10061 VDD.n3362 VSS 0.00109f
C10062 VDD.n3363 VSS 8.89e-19
C10063 VDD.t645 VSS 0.00584f
C10064 VDD.n3364 VSS 0.00603f
C10065 VDD.n3365 VSS 0.00109f
C10066 VDD.n3366 VSS 9.31e-19
C10067 VDD.n3367 VSS 5.67e-19
C10068 VDD.n3368 VSS 0.00278f
C10069 VDD.n3369 VSS 0.00325f
C10070 VDD.n3370 VSS 9.31e-19
C10071 VDD.n3371 VSS 0.0113f
C10072 VDD.n3372 VSS 0.00109f
C10073 VDD.n3373 VSS 0.00121f
C10074 VDD.n3374 VSS 0.0117f
C10075 VDD.n3375 VSS 0.00109f
C10076 VDD.n3376 VSS 0.00156f
C10077 VDD.n3377 VSS 0.00184f
C10078 VDD.n3378 VSS 0.00109f
C10079 VDD.n3379 VSS 0.00762f
C10080 VDD.t273 VSS 0.00406f
C10081 VDD.n3380 VSS 0.00692f
C10082 VDD.n3381 VSS 0.00109f
C10083 VDD.n3382 VSS 9.51e-19
C10084 VDD.n3383 VSS 0.00308f
C10085 VDD.t373 VSS 0.00584f
C10086 VDD.n3384 VSS 0.00654f
C10087 VDD.n3385 VSS 0.00109f
C10088 VDD.n3386 VSS 0.00172f
C10089 VDD.n3387 VSS 0.00285f
C10090 VDD.n3388 VSS 0.00154f
C10091 VDD.t555 VSS 0.00584f
C10092 VDD.n3389 VSS 0.00686f
C10093 VDD.n3390 VSS 0.00109f
C10094 VDD.n3391 VSS 9.31e-19
C10095 VDD.n3392 VSS 1.72e-19
C10096 VDD.n3393 VSS 2.85e-19
C10097 VDD.n3394 VSS 9.31e-19
C10098 VDD.n3395 VSS 2.51e-19
C10099 VDD.n3396 VSS 4.35e-19
C10100 VDD.n3397 VSS 3.36e-19
C10101 VDD.n3398 VSS 8.1e-19
C10102 VDD.n3399 VSS 0.00157f
C10103 VDD.n3400 VSS 0.00278f
C10104 VDD.t407 VSS 0.00584f
C10105 VDD.n3401 VSS 0.0113f
C10106 VDD.n3402 VSS 0.00109f
C10107 VDD.n3403 VSS 0.00121f
C10108 VDD.n3404 VSS 0.00144f
C10109 VDD.n3405 VSS 0.00707f
C10110 VDD.n3406 VSS 0.0442f
C10111 VDD.n3407 VSS 0.00377f
C10112 VDD.n3408 VSS 0.00582f
C10113 VDD.n3409 VSS 0.0117f
C10114 VDD.n3410 VSS 0.00109f
C10115 VDD.n3411 VSS 0.00186f
C10116 VDD.n3412 VSS 0.00248f
C10117 VDD.t391 VSS 4.25e-19
C10118 VDD.t466 VSS 5.42e-19
C10119 VDD.n3413 VSS 0.00111f
C10120 VDD.n3414 VSS 0.00259f
C10121 VDD.t390 VSS 0.00584f
C10122 VDD.n3415 VSS 0.00597f
C10123 VDD.n3416 VSS 0.00109f
C10124 VDD.n3417 VSS 0.0014f
C10125 VDD.n3418 VSS 0.00308f
C10126 VDD.t465 VSS 0.00495f
C10127 VDD.n3419 VSS 0.0061f
C10128 VDD.n3420 VSS 0.00109f
C10129 VDD.n3421 VSS 0.0014f
C10130 VDD.n3422 VSS 0.00308f
C10131 VDD.t256 VSS 0.00546f
C10132 VDD.n3423 VSS 0.00673f
C10133 VDD.n3424 VSS 0.00109f
C10134 VDD.n3425 VSS 0.00186f
C10135 VDD.n3426 VSS 0.00308f
C10136 VDD.n3427 VSS 0.0117f
C10137 VDD.n3428 VSS 0.00109f
C10138 VDD.n3429 VSS 0.00186f
C10139 VDD.n3430 VSS 0.00308f
C10140 VDD.t556 VSS 0.00584f
C10141 VDD.n3431 VSS 0.00686f
C10142 VDD.n3432 VSS 0.00109f
C10143 VDD.n3433 VSS 0.00186f
C10144 VDD.n3434 VSS 0.00308f
C10145 VDD.t702 VSS 0.00584f
C10146 VDD.n3435 VSS 0.00654f
C10147 VDD.n3436 VSS 0.00109f
C10148 VDD.n3437 VSS 0.00186f
C10149 VDD.n3438 VSS 0.00308f
C10150 VDD.n3439 VSS 0.00308f
C10151 VDD.n3440 VSS 0.0117f
C10152 VDD.n3441 VSS 0.00109f
C10153 VDD.n3442 VSS 0.00156f
C10154 VDD.t703 VSS 7.73e-19
C10155 VDD.t41 VSS 2.51e-19
C10156 VDD.n3443 VSS 0.00395f
C10157 VDD.n3444 VSS 0.00308f
C10158 VDD.n3445 VSS 9.51e-19
C10159 VDD.n3446 VSS 0.00109f
C10160 VDD.n3447 VSS 0.00692f
C10161 VDD.t40 VSS 0.00406f
C10162 VDD.n3448 VSS 0.00762f
C10163 VDD.n3449 VSS 0.00109f
C10164 VDD.n3450 VSS 0.00184f
C10165 VDD.n3451 VSS 0.00181f
C10166 VDD.n3452 VSS 0.00325f
C10167 VDD.n3453 VSS 9.31e-19
C10168 VDD.t741 VSS 7.73e-19
C10169 VDD.t408 VSS 2.51e-19
C10170 VDD.n3454 VSS 0.00395f
C10171 VDD.n3455 VSS 5.67e-19
C10172 VDD.n3456 VSS 0.00253f
C10173 VDD.n3457 VSS 9.11e-19
C10174 VDD.n3458 VSS 0.00109f
C10175 VDD.n3459 VSS 8.89e-19
C10176 VDD.t740 VSS 0.00584f
C10177 VDD.n3460 VSS 0.00603f
C10178 VDD.n3461 VSS 0.00109f
C10179 VDD.n3462 VSS 9.31e-19
C10180 VDD.n3463 VSS 9.31e-19
C10181 VDD.n3464 VSS 0.00308f
C10182 VDD.t554 VSS 0.00584f
C10183 VDD.n3465 VSS 0.00654f
C10184 VDD.n3466 VSS 0.00109f
C10185 VDD.n3467 VSS 9.31e-19
C10186 VDD.n3468 VSS 9.31e-19
C10187 VDD.n3469 VSS 0.00308f
C10188 VDD.n3470 VSS 0.0103f
C10189 VDD.n3471 VSS 0.00109f
C10190 VDD.n3472 VSS 9.31e-19
C10191 VDD.n3473 VSS 9.31e-19
C10192 VDD.n3474 VSS 0.00308f
C10193 VDD.n3475 VSS 0.00915f
C10194 VDD.n3476 VSS 0.00109f
C10195 VDD.n3477 VSS 9.31e-19
C10196 VDD.n3478 VSS 9.31e-19
C10197 VDD.n3479 VSS 0.00308f
C10198 VDD.t604 VSS 0.00584f
C10199 VDD.t219 VSS 0.00584f
C10200 VDD.n3480 VSS 0.00457f
C10201 VDD.n3481 VSS 0.00109f
C10202 VDD.n3482 VSS 9.31e-19
C10203 VDD.n3483 VSS 8.5e-19
C10204 VDD.n3484 VSS 0.00308f
C10205 VDD.t220 VSS 5.42e-19
C10206 VDD.t173 VSS 4.25e-19
C10207 VDD.n3485 VSS 0.00111f
C10208 VDD.n3486 VSS 0.0022f
C10209 VDD.t172 VSS 0.00584f
C10210 VDD.n3487 VSS 0.0061f
C10211 VDD.n3488 VSS 0.00109f
C10212 VDD.n3489 VSS 4.66e-19
C10213 VDD.n3490 VSS 9.31e-19
C10214 VDD.n3491 VSS 0.00308f
C10215 VDD.n3492 VSS 0.0094f
C10216 VDD.n3493 VSS 0.00109f
C10217 VDD.n3494 VSS 9.31e-19
C10218 VDD.n3495 VSS 0.0117f
C10219 VDD.n3496 VSS 0.00109f
C10220 VDD.n3497 VSS 0.00157f
C10221 VDD.n3498 VSS 0.0117f
C10222 VDD.n3499 VSS 0.00107f
C10223 VDD.n3500 VSS 0.00157f
C10224 VDD.n3501 VSS 0.0117f
C10225 VDD.n3502 VSS 0.00141f
C10226 VDD.n3503 VSS 0.00157f
C10227 VDD.n3504 VSS 0.0117f
C10228 VDD.n3505 VSS 0.00107f
C10229 VDD.n3506 VSS 0.0013f
C10230 VDD.n3507 VSS 9.41e-19
C10231 VDD.n3508 VSS 0.00228f
C10232 VDD.n3509 VSS 0.00158f
C10233 VDD.n3510 VSS 8.1e-19
C10234 VDD.n3511 VSS 0.00148f
C10235 VDD.n3512 VSS 0.00144f
C10236 VDD.n3513 VSS 0.00844f
C10237 VDD.n3514 VSS 7.71e-19
C10238 VDD.n3515 VSS 0.00144f
C10239 VDD.n3516 VSS 0.00148f
C10240 VDD.n3517 VSS 8.1e-19
C10241 VDD.n3518 VSS 0.00157f
C10242 VDD.n3519 VSS 0.00726f
C10243 VDD.n3520 VSS 0.00725f
C10244 VDD.n3521 VSS 0.151f
C10245 VDD.n3522 VSS 0.151f
C10246 VDD.n3523 VSS 9.67e-19
C10247 VDD.n3524 VSS 0.00121f
C10248 VDD.n3525 VSS 0.00145f
C10249 VDD.n3526 VSS 0.00556f
C10250 VDD.n3527 VSS 0.00149f
C10251 VDD.n3528 VSS 5.97e-19
C10252 VDD.n3529 VSS 5.16e-19
C10253 VDD.t611 VSS 0.00217f
C10254 VDD.t228 VSS 9.67e-19
C10255 VDD.n3530 VSS 0.00349f
C10256 VDD.n3531 VSS 0.00457f
C10257 VDD.t227 VSS 0.00565f
C10258 VDD.n3532 VSS 0.00616f
C10259 VDD.n3533 VSS 0.00109f
C10260 VDD.n3534 VSS 9.61e-19
C10261 VDD.n3535 VSS 0.00255f
C10262 VDD.n3536 VSS 0.00117f
C10263 VDD.n3537 VSS 4.35e-19
C10264 VDD.n3538 VSS 0.00136f
C10265 VDD.t495 VSS 0.00578f
C10266 VDD.n3539 VSS 0.00666f
C10267 VDD.n3540 VSS 0.00109f
C10268 VDD.n3541 VSS 0.00107f
C10269 VDD.n3542 VSS 0.00245f
C10270 VDD.n3543 VSS 0.00154f
C10271 VDD.n3544 VSS 9.31e-19
C10272 VDD.t512 VSS 0.0054f
C10273 VDD.n3545 VSS 0.0059f
C10274 VDD.n3546 VSS 0.00109f
C10275 VDD.n3547 VSS 1.72e-19
C10276 VDD.n3548 VSS 2.85e-19
C10277 VDD.n3549 VSS 9.31e-19
C10278 VDD.n3550 VSS 3.68e-19
C10279 VDD.n3551 VSS 4.35e-19
C10280 VDD.n3552 VSS 3.36e-19
C10281 VDD.n3553 VSS 8.1e-19
C10282 VDD.n3554 VSS 0.00157f
C10283 VDD.n3555 VSS 0.00532f
C10284 VDD.n3556 VSS 0.00158f
C10285 VDD.n3557 VSS 6.17e-19
C10286 VDD.t193 VSS 0.00578f
C10287 VDD.n3558 VSS 0.00528f
C10288 VDD.n3559 VSS 0.00109f
C10289 VDD.n3560 VSS 0.00178f
C10290 VDD.n3561 VSS 0.00251f
C10291 VDD.n3562 VSS 0.00111f
C10292 VDD.t610 VSS 0.00578f
C10293 VDD.n3563 VSS 0.00823f
C10294 VDD.n3564 VSS 0.00109f
C10295 VDD.n3565 VSS 0.00101f
C10296 VDD.n3566 VSS 0.00293f
C10297 VDD.n3567 VSS 0.00154f
C10298 VDD.n3568 VSS 0.00905f
C10299 VDD.n3569 VSS 0.00109f
C10300 VDD.n3570 VSS 9.31e-19
C10301 VDD.n3571 VSS 1.72e-19
C10302 VDD.n3572 VSS 2.85e-19
C10303 VDD.n3573 VSS 9.31e-19
C10304 VDD.n3574 VSS 4.35e-19
C10305 VDD.n3575 VSS 4.35e-19
C10306 VDD.n3576 VSS 4.94e-19
C10307 VDD.n3577 VSS 3.36e-19
C10308 VDD.n3578 VSS 8.1e-19
C10309 VDD.n3579 VSS 0.00148f
C10310 VDD.n3580 VSS 9.68e-19
C10311 VDD.n3581 VSS 0.00193f
C10312 VDD.n3582 VSS 0.151f
C10313 VDD.n3583 VSS 0.15f
C10314 VDD.n3584 VSS 0.00145f
C10315 VDD.n3585 VSS 0.00121f
C10316 VDD.n3586 VSS 9.67e-19
C10317 VDD.n3587 VSS 0.00532f
C10318 VDD.n3588 VSS 0.00158f
C10319 VDD.n3589 VSS 5.16e-19
C10320 VDD.n3590 VSS 5.96e-19
C10321 VDD.n3591 VSS 3.36e-19
C10322 VDD.n3592 VSS 8.1e-19
C10323 VDD.n3593 VSS 0.00148f
C10324 VDD.n3594 VSS 0.00556f
C10325 VDD.n3595 VSS 0.00158f
C10326 VDD.n3596 VSS 3.87e-19
C10327 VDD.n3597 VSS 2.97e-19
C10328 VDD.n3598 VSS 4.69e-19
C10329 VDD.t496 VSS 5.72e-19
C10330 VDD.t609 VSS 5.42e-19
C10331 VDD.n3599 VSS 0.00118f
C10332 VDD.n3600 VSS 0.00258f
C10333 VDD.n3601 VSS 2.25e-19
C10334 VDD.n3602 VSS 1.84e-19
C10335 VDD.n3603 VSS 8.4e-19
C10336 VDD.n3604 VSS 5.49e-19
C10337 VDD.t608 VSS 0.00578f
C10338 VDD.n3605 VSS 0.00666f
C10339 VDD.n3606 VSS 0.0011f
C10340 VDD.n3607 VSS 6.6e-19
C10341 VDD.n3608 VSS 3.28e-19
C10342 VDD.n3609 VSS 0.00154f
C10343 VDD.n3610 VSS 0.00754f
C10344 VDD.n3611 VSS 0.00109f
C10345 VDD.n3612 VSS 0.0017f
C10346 VDD.n3613 VSS 0.00248f
C10347 VDD.n3614 VSS 0.00154f
C10348 VDD.t192 VSS 0.00578f
C10349 VDD.n3615 VSS 0.00528f
C10350 VDD.n3616 VSS 0.00109f
C10351 VDD.n3617 VSS 0.00186f
C10352 VDD.n3618 VSS 3.85e-19
C10353 VDD.t180 VSS 0.00578f
C10354 VDD.n3619 VSS 0.00578f
C10355 VDD.n3620 VSS 0.00109f
C10356 VDD.n3621 VSS 0.00151f
C10357 VDD.n3622 VSS 0.00263f
C10358 VDD.n3623 VSS 0.00149f
C10359 VDD.n3624 VSS 3.85e-19
C10360 VDD.n3625 VSS 2.97e-19
C10361 VDD.n3626 VSS 8.1e-19
C10362 VDD.n3627 VSS 0.00148f
C10363 VDD.n3628 VSS 0.00145f
C10364 VDD.n3629 VSS 4.69e-19
C10365 VDD.t738 VSS 0.00578f
C10366 VDD.n3630 VSS 0.00151f
C10367 VDD.t708 VSS 0.00578f
C10368 VDD.n3631 VSS 0.00154f
C10369 VDD.n3632 VSS 3.85e-19
C10370 VDD.t237 VSS 0.00578f
C10371 VDD.n3633 VSS 0.00603f
C10372 VDD.n3634 VSS 0.00109f
C10373 VDD.n3635 VSS 1.72e-19
C10374 VDD.n3636 VSS 2.85e-19
C10375 VDD.n3637 VSS 9.31e-19
C10376 VDD.n3638 VSS 2.18e-19
C10377 VDD.n3639 VSS 5.79e-19
C10378 VDD.n3640 VSS 5.28e-19
C10379 VDD.n3641 VSS 3.36e-19
C10380 VDD.n3642 VSS 4.35e-19
C10381 VDD.n3643 VSS 0.00132f
C10382 VDD.t706 VSS 0.00578f
C10383 VDD.n3644 VSS 0.00634f
C10384 VDD.n3645 VSS 0.00109f
C10385 VDD.n3646 VSS 0.00184f
C10386 VDD.n3647 VSS 0.00261f
C10387 VDD.t225 VSS 0.00578f
C10388 VDD.n3648 VSS 0.00528f
C10389 VDD.n3649 VSS 0.00109f
C10390 VDD.n3650 VSS 0.00186f
C10391 VDD.n3651 VSS 0.00308f
C10392 VDD.n3652 VSS 0.00905f
C10393 VDD.n3653 VSS 0.00109f
C10394 VDD.n3654 VSS 0.00186f
C10395 VDD.n3655 VSS 0.00308f
C10396 VDD.t194 VSS 0.00578f
C10397 VDD.n3656 VSS 0.00823f
C10398 VDD.n3657 VSS 0.00109f
C10399 VDD.n3658 VSS 0.0011f
C10400 VDD.n3659 VSS 0.00308f
C10401 VDD.t195 VSS 0.00217f
C10402 VDD.t695 VSS 9.67e-19
C10403 VDD.n3660 VSS 0.00349f
C10404 VDD.n3661 VSS 0.00457f
C10405 VDD.t694 VSS 0.00565f
C10406 VDD.n3662 VSS 0.00616f
C10407 VDD.n3663 VSS 0.00109f
C10408 VDD.n3664 VSS 0.00102f
C10409 VDD.n3665 VSS 0.00308f
C10410 VDD.t704 VSS 0.0054f
C10411 VDD.n3666 VSS 0.0059f
C10412 VDD.n3667 VSS 0.00109f
C10413 VDD.n3668 VSS 0.00186f
C10414 VDD.n3669 VSS 0.00308f
C10415 VDD.t378 VSS 0.00578f
C10416 VDD.n3670 VSS 0.00666f
C10417 VDD.n3671 VSS 0.00109f
C10418 VDD.n3672 VSS 0.00118f
C10419 VDD.n3673 VSS 0.00308f
C10420 VDD.t379 VSS 5.72e-19
C10421 VDD.t197 VSS 5.42e-19
C10422 VDD.n3674 VSS 0.00119f
C10423 VDD.t196 VSS 0.00578f
C10424 VDD.n3675 VSS 0.00666f
C10425 VDD.n3676 VSS 0.00111f
C10426 VDD.n3677 VSS 0.00204f
C10427 VDD.n3678 VSS 0.00278f
C10428 VDD.n3679 VSS 0.00308f
C10429 VDD.n3680 VSS 0.00754f
C10430 VDD.n3681 VSS 0.00109f
C10431 VDD.n3682 VSS 0.00177f
C10432 VDD.n3683 VSS 0.00308f
C10433 VDD.t226 VSS 0.00578f
C10434 VDD.n3684 VSS 0.00528f
C10435 VDD.n3685 VSS 0.00109f
C10436 VDD.n3686 VSS 0.00186f
C10437 VDD.n3687 VSS 0.00308f
C10438 VDD.t707 VSS 0.00578f
C10439 VDD.n3688 VSS 0.00578f
C10440 VDD.n3689 VSS 0.00109f
C10441 VDD.n3690 VSS 0.00151f
C10442 VDD.n3691 VSS 0.00308f
C10443 VDD.t338 VSS 0.00142f
C10444 VDD.t337 VSS 0.00578f
C10445 VDD.n3692 VSS 0.00854f
C10446 VDD.n3693 VSS 0.00111f
C10447 VDD.n3694 VSS 0.00203f
C10448 VDD.n3695 VSS 0.00312f
C10449 VDD.n3696 VSS 0.00308f
C10450 VDD.n3697 VSS 0.00905f
C10451 VDD.n3698 VSS 0.00109f
C10452 VDD.n3699 VSS 0.00118f
C10453 VDD.n3700 VSS 0.00308f
C10454 VDD.n3701 VSS 0.00183f
C10455 VDD.n3702 VSS 0.00308f
C10456 VDD.t709 VSS 6.03e-19
C10457 VDD.t292 VSS 6.03e-19
C10458 VDD.n3703 VSS 0.0013f
C10459 VDD.n3704 VSS 0.0027f
C10460 VDD.n3705 VSS 0.00202f
C10461 VDD.n3706 VSS 0.00111f
C10462 VDD.n3707 VSS 0.00528f
C10463 VDD.t291 VSS 0.00578f
C10464 VDD.n3708 VSS 0.00109f
C10465 VDD.n3709 VSS 0.00773f
C10466 VDD.n3710 VSS 0.00109f
C10467 VDD.n3711 VSS 0.0018f
C10468 VDD.n3712 VSS 0.00231f
C10469 VDD.t260 VSS -2.71e-19
C10470 VDD.t187 VSS 8.49e-19
C10471 VDD.n3713 VSS 0.00391f
C10472 VDD.n3714 VSS 0.00413f
C10473 VDD.t259 VSS 0.00578f
C10474 VDD.n3715 VSS 0.00597f
C10475 VDD.n3716 VSS 0.00109f
C10476 VDD.n3717 VSS 9.92e-19
C10477 VDD.n3718 VSS 0.00308f
C10478 VDD.t186 VSS 0.00578f
C10479 VDD.n3719 VSS 0.00835f
C10480 VDD.n3720 VSS 0.00109f
C10481 VDD.n3721 VSS 0.00186f
C10482 VDD.n3722 VSS 0.00308f
C10483 VDD.t184 VSS 0.00955f
C10484 VDD.n3723 VSS 0.00923f
C10485 VDD.n3724 VSS 6.76e-19
C10486 VDD.n3725 VSS 0.00179f
C10487 VDD.n3726 VSS 0.00308f
C10488 VDD.t185 VSS -5.07e-19
C10489 VDD.t119 VSS 9.16e-19
C10490 VDD.n3727 VSS 0.00359f
C10491 VDD.n3728 VSS 0.00204f
C10492 VDD.n3729 VSS 0.00187f
C10493 VDD.n3730 VSS 0.00281f
C10494 VDD.n3731 VSS 0.00154f
C10495 VDD.t763 VSS 8.67e-19
C10496 VDD.n3732 VSS 0.00281f
C10497 VDD.t117 VSS 0.00159f
C10498 VDD.n3733 VSS 0.00354f
C10499 VDD.n3734 VSS 7.59e-19
C10500 VDD.n3735 VSS 0.00206f
C10501 VDD.n3736 VSS 3.97e-19
C10502 VDD.n3737 VSS 2.85e-19
C10503 VDD.n3738 VSS 0.00147f
C10504 VDD.n3739 VSS 0.00152f
C10505 VDD.n3740 VSS 0.00213f
C10506 VDD.t118 VSS 0.0139f
C10507 VDD.n3741 VSS 0.0119f
C10508 VDD.n3742 VSS 7.81e-19
C10509 VDD.n3743 VSS 3.97e-19
C10510 VDD.n3744 VSS 2.85e-19
C10511 VDD.t288 VSS 0.00262f
C10512 VDD.n3745 VSS 0.0024f
C10513 VDD.n3746 VSS 5.38e-19
C10514 VDD.n3747 VSS 5.7e-19
C10515 VDD.n3748 VSS 4.52e-19
C10516 VDD.n3749 VSS 0.00158f
C10517 VDD.n3750 VSS 0.00218f
C10518 VDD.n3751 VSS 0.152f
C10519 VDD.n3752 VSS 0.151f
C10520 VDD.n3753 VSS 9.67e-19
C10521 VDD.n3754 VSS 0.00121f
C10522 VDD.n3755 VSS 0.00121f
C10523 VDD.n3756 VSS 0.00556f
C10524 VDD.n3757 VSS 0.00556f
C10525 VDD.n3758 VSS 9.67e-19
C10526 VDD.n3759 VSS 9.67e-19
C10527 VDD.n3760 VSS 0.00121f
C10528 VDD.n3761 VSS 0.15f
C10529 VDD.n3762 VSS 0.15f
C10530 VDD.n3763 VSS 0.00121f
C10531 VDD.n3764 VSS 0.00121f
C10532 VDD.n3765 VSS 9.67e-19
C10533 VDD.n3766 VSS 0.00556f
C10534 VDD.n3767 VSS 0.00556f
C10535 VDD.n3768 VSS 0.00121f
C10536 VDD.n3769 VSS 0.00122f
C10537 VDD.n3770 VSS 9.68e-19
C10538 VDD.n3771 VSS 0.00556f
C10539 VDD.n3772 VSS 0.00148f
C10540 VDD.n3773 VSS 8.1e-19
C10541 VDD.n3774 VSS 6.6e-19
C10542 VDD.n3775 VSS 3.36e-19
C10543 VDD.n3776 VSS 4.35e-19
C10544 VDD.n3777 VSS 9.71e-19
C10545 VDD.t287 VSS 0.00578f
C10546 VDD.t651 VSS 0.00578f
C10547 VDD.n3778 VSS 0.00452f
C10548 VDD.n3779 VSS 0.00109f
C10549 VDD.n3780 VSS 0.00171f
C10550 VDD.n3781 VSS 0.00241f
C10551 VDD.n3782 VSS 0.00154f
C10552 VDD.n3783 VSS 9.31e-19
C10553 VDD.n3784 VSS 0.00666f
C10554 VDD.n3785 VSS 0.00109f
C10555 VDD.n3786 VSS 1.72e-19
C10556 VDD.n3787 VSS 2.85e-19
C10557 VDD.n3788 VSS 7.08e-19
C10558 VDD.n3789 VSS 6.87e-19
C10559 VDD.n3790 VSS 4.05e-19
C10560 VDD.n3791 VSS 7.06e-19
C10561 VDD.n3792 VSS 0.00157f
C10562 VDD.n3793 VSS 0.00149f
C10563 VDD.n3794 VSS 8.1e-19
C10564 VDD.n3795 VSS 3.36e-19
C10565 VDD.n3796 VSS 4.35e-19
C10566 VDD.n3797 VSS 8.54e-19
C10567 VDD.t27 VSS 5.72e-19
C10568 VDD.t189 VSS 7.62e-19
C10569 VDD.n3798 VSS 0.0014f
C10570 VDD.t26 VSS 0.00578f
C10571 VDD.n3799 VSS 0.0076f
C10572 VDD.n3800 VSS 0.00111f
C10573 VDD.n3801 VSS 0.00188f
C10574 VDD.n3802 VSS 0.00252f
C10575 VDD.n3803 VSS 0.00238f
C10576 VDD.t188 VSS 0.00578f
C10577 VDD.n3804 VSS 0.00603f
C10578 VDD.n3805 VSS 0.00109f
C10579 VDD.n3806 VSS 0.00121f
C10580 VDD.n3807 VSS 0.00248f
C10581 VDD.n3808 VSS 0.00104f
C10582 VDD.n3809 VSS 6.43e-19
C10583 VDD.n3810 VSS 4.69e-19
C10584 VDD.n3811 VSS 0.00158f
C10585 VDD.n3812 VSS 0.00148f
C10586 VDD.n3813 VSS 8.1e-19
C10587 VDD.n3814 VSS 3.36e-19
C10588 VDD.n3815 VSS 4.35e-19
C10589 VDD.n3816 VSS 9.31e-19
C10590 VDD.n3817 VSS 5.03e-19
C10591 VDD.n3818 VSS 9.31e-19
C10592 VDD.t331 VSS 0.00578f
C10593 VDD.n3819 VSS 0.00634f
C10594 VDD.n3820 VSS 0.00109f
C10595 VDD.n3821 VSS 1.72e-19
C10596 VDD.n3822 VSS 2.85e-19
C10597 VDD.n3823 VSS 0.00154f
C10598 VDD.t355 VSS 0.00578f
C10599 VDD.n3824 VSS 0.00528f
C10600 VDD.n3825 VSS 0.00109f
C10601 VDD.n3826 VSS 0.00171f
C10602 VDD.n3827 VSS 0.0024f
C10603 VDD.n3828 VSS 0.00112f
C10604 VDD.n3829 VSS 6.1e-19
C10605 VDD.n3830 VSS 5.03e-19
C10606 VDD.n3831 VSS 0.00157f
C10607 VDD.n3832 VSS 0.00149f
C10608 VDD.n3833 VSS 8.1e-19
C10609 VDD.n3834 VSS 3.36e-19
C10610 VDD.n3835 VSS 4.35e-19
C10611 VDD.n3836 VSS 9.31e-19
C10612 VDD.n3837 VSS 4.19e-19
C10613 VDD.n3838 VSS 0.00905f
C10614 VDD.n3839 VSS 0.00109f
C10615 VDD.n3840 VSS 9.31e-19
C10616 VDD.n3841 VSS 1.72e-19
C10617 VDD.n3842 VSS 2.85e-19
C10618 VDD.n3843 VSS 0.00154f
C10619 VDD.t588 VSS 0.00578f
C10620 VDD.n3844 VSS 0.00823f
C10621 VDD.n3845 VSS 0.00109f
C10622 VDD.n3846 VSS 0.00101f
C10623 VDD.n3847 VSS 0.00293f
C10624 VDD.t589 VSS 0.00217f
C10625 VDD.t290 VSS 9.67e-19
C10626 VDD.n3848 VSS 0.00349f
C10627 VDD.n3849 VSS 0.00457f
C10628 VDD.t289 VSS 0.00565f
C10629 VDD.n3850 VSS 0.00616f
C10630 VDD.n3851 VSS 0.00109f
C10631 VDD.n3852 VSS 0.00102f
C10632 VDD.n3853 VSS 0.00308f
C10633 VDD.t735 VSS 0.0054f
C10634 VDD.n3854 VSS 0.0059f
C10635 VDD.n3855 VSS 0.00109f
C10636 VDD.n3856 VSS 0.0017f
C10637 VDD.n3857 VSS 0.00238f
C10638 VDD.n3858 VSS 0.00148f
C10639 VDD.n3859 VSS 8.1e-19
C10640 VDD.n3860 VSS 0.00157f
C10641 VDD.n3861 VSS 3.92e-19
C10642 VDD.n3862 VSS 0.00105f
C10643 VDD.n3863 VSS 0.00127f
C10644 VDD.n3864 VSS 9.31e-19
C10645 VDD.n3865 VSS 7.03e-19
C10646 VDD.t508 VSS 0.00578f
C10647 VDD.n3866 VSS 0.00666f
C10648 VDD.n3867 VSS 0.00109f
C10649 VDD.n3868 VSS 2.53e-19
C10650 VDD.n3869 VSS 1.72e-19
C10651 VDD.n3870 VSS 2.85e-19
C10652 VDD.n3871 VSS 0.00154f
C10653 VDD.t509 VSS 5.72e-19
C10654 VDD.t587 VSS 5.42e-19
C10655 VDD.n3872 VSS 0.00119f
C10656 VDD.t586 VSS 0.00578f
C10657 VDD.n3873 VSS 0.00666f
C10658 VDD.n3874 VSS 0.00111f
C10659 VDD.n3875 VSS 0.00203f
C10660 VDD.n3876 VSS 0.00278f
C10661 VDD.n3877 VSS 0.00307f
C10662 VDD.n3878 VSS 0.00754f
C10663 VDD.n3879 VSS 0.00109f
C10664 VDD.n3880 VSS 0.00177f
C10665 VDD.n3881 VSS 0.00308f
C10666 VDD.t356 VSS 0.00578f
C10667 VDD.n3882 VSS 0.00528f
C10668 VDD.n3883 VSS 0.00109f
C10669 VDD.n3884 VSS 0.00186f
C10670 VDD.n3885 VSS 0.00308f
C10671 VDD.t332 VSS 0.00578f
C10672 VDD.n3886 VSS 0.00578f
C10673 VDD.n3887 VSS 0.00109f
C10674 VDD.n3888 VSS 0.00151f
C10675 VDD.n3889 VSS 0.00308f
C10676 VDD.t570 VSS 0.00142f
C10677 VDD.t569 VSS 0.00578f
C10678 VDD.n3890 VSS 0.00854f
C10679 VDD.n3891 VSS 0.00111f
C10680 VDD.n3892 VSS 0.00203f
C10681 VDD.n3893 VSS 0.00312f
C10682 VDD.n3894 VSS 0.00308f
C10683 VDD.n3895 VSS 0.00905f
C10684 VDD.n3896 VSS 0.00109f
C10685 VDD.n3897 VSS 0.00118f
C10686 VDD.n3898 VSS 0.00308f
C10687 VDD.t330 VSS 6.03e-19
C10688 VDD.t739 VSS 6.03e-19
C10689 VDD.n3899 VSS 0.0013f
C10690 VDD.t329 VSS 0.00578f
C10691 VDD.n3900 VSS 0.00528f
C10692 VDD.n3901 VSS 0.00111f
C10693 VDD.n3902 VSS 0.00202f
C10694 VDD.n3903 VSS 0.0027f
C10695 VDD.n3904 VSS 0.00308f
C10696 VDD.n3905 VSS 0.00183f
C10697 VDD.n3906 VSS 0.00151f
C10698 VDD.n3907 VSS 0.00109f
C10699 VDD.n3908 VSS 0.00773f
C10700 VDD.n3909 VSS 0.00109f
C10701 VDD.n3910 VSS 0.0018f
C10702 VDD.n3911 VSS 0.00231f
C10703 VDD.t37 VSS -2.71e-19
C10704 VDD.t350 VSS 8.49e-19
C10705 VDD.n3912 VSS 0.00391f
C10706 VDD.n3913 VSS 0.00413f
C10707 VDD.t36 VSS 0.00578f
C10708 VDD.n3914 VSS 0.00597f
C10709 VDD.n3915 VSS 0.00109f
C10710 VDD.n3916 VSS 9.92e-19
C10711 VDD.n3917 VSS 0.00308f
C10712 VDD.t349 VSS 0.00578f
C10713 VDD.n3918 VSS 0.00835f
C10714 VDD.n3919 VSS 0.00109f
C10715 VDD.n3920 VSS 0.00186f
C10716 VDD.n3921 VSS 0.00308f
C10717 VDD.t353 VSS 0.00955f
C10718 VDD.n3922 VSS 0.00923f
C10719 VDD.n3923 VSS 6.76e-19
C10720 VDD.n3924 VSS 0.00179f
C10721 VDD.n3925 VSS 0.00308f
C10722 VDD.t354 VSS -5.07e-19
C10723 VDD.t113 VSS 9.16e-19
C10724 VDD.n3926 VSS 0.00359f
C10725 VDD.n3927 VSS 0.00204f
C10726 VDD.n3928 VSS 0.00187f
C10727 VDD.n3929 VSS 0.00281f
C10728 VDD.n3930 VSS 0.00154f
C10729 VDD.t765 VSS 8.67e-19
C10730 VDD.n3931 VSS 0.00281f
C10731 VDD.t111 VSS 0.00159f
C10732 VDD.n3932 VSS 0.00354f
C10733 VDD.n3933 VSS 7.59e-19
C10734 VDD.n3934 VSS 0.00215f
C10735 VDD.n3935 VSS 3.97e-19
C10736 VDD.n3936 VSS 2.85e-19
C10737 VDD.n3937 VSS 0.00154f
C10738 VDD.t112 VSS 0.0139f
C10739 VDD.n3938 VSS 0.0119f
C10740 VDD.n3939 VSS 7.5e-19
C10741 VDD.t230 VSS 0.00262f
C10742 VDD.n3940 VSS 0.00271f
C10743 VDD.n3941 VSS 0.00267f
C10744 VDD.n3942 VSS 0.00307f
C10745 VDD.t229 VSS 0.00578f
C10746 VDD.t299 VSS 0.00578f
C10747 VDD.n3943 VSS 0.00452f
C10748 VDD.n3944 VSS 0.00109f
C10749 VDD.n3945 VSS 0.00172f
C10750 VDD.n3946 VSS 0.00308f
C10751 VDD.n3947 VSS 0.00666f
C10752 VDD.n3948 VSS 0.00109f
C10753 VDD.n3949 VSS 0.00164f
C10754 VDD.n3950 VSS 0.00308f
C10755 VDD.t169 VSS 5.72e-19
C10756 VDD.t352 VSS 7.62e-19
C10757 VDD.n3951 VSS 0.0014f
C10758 VDD.t168 VSS 0.00578f
C10759 VDD.n3952 VSS 0.0076f
C10760 VDD.n3953 VSS 0.00111f
C10761 VDD.n3954 VSS 0.00198f
C10762 VDD.n3955 VSS 0.00252f
C10763 VDD.n3956 VSS 0.00298f
C10764 VDD.n3957 VSS 0.00154f
C10765 VDD.n3958 VSS 3.85e-19
C10766 VDD.t351 VSS 0.00578f
C10767 VDD.n3959 VSS 0.00603f
C10768 VDD.n3960 VSS 0.00109f
C10769 VDD.n3961 VSS 1.72e-19
C10770 VDD.n3962 VSS 2.85e-19
C10771 VDD.n3963 VSS 9.31e-19
C10772 VDD.n3964 VSS 5.19e-19
C10773 VDD.t183 VSS 0.00578f
C10774 VDD.n3965 VSS 0.00634f
C10775 VDD.n3966 VSS 0.00109f
C10776 VDD.n3967 VSS 0.00175f
C10777 VDD.n3968 VSS 0.00246f
C10778 VDD.n3969 VSS 0.00102f
C10779 VDD.n3970 VSS 4.35e-19
C10780 VDD.n3971 VSS 6.43e-19
C10781 VDD.n3972 VSS 3.36e-19
C10782 VDD.n3973 VSS 0.00149f
C10783 VDD.n3974 VSS 8.1e-19
C10784 VDD.n3975 VSS 0.00157f
C10785 VDD.n3976 VSS 0.00121f
C10786 VDD.n3977 VSS 0.00148f
C10787 VDD.n3978 VSS 8.1e-19
C10788 VDD.n3979 VSS 6.6e-19
C10789 VDD.n3980 VSS 3.36e-19
C10790 VDD.n3981 VSS 4.35e-19
C10791 VDD.n3982 VSS 9.71e-19
C10792 VDD.n3983 VSS 0.00905f
C10793 VDD.n3984 VSS 0.00109f
C10794 VDD.n3985 VSS 0.00118f
C10795 VDD.n3986 VSS 0.00243f
C10796 VDD.t182 VSS 6.03e-19
C10797 VDD.t161 VSS 6.03e-19
C10798 VDD.n3987 VSS 0.0013f
C10799 VDD.t181 VSS 0.00578f
C10800 VDD.n3988 VSS 0.00528f
C10801 VDD.n3989 VSS 0.00111f
C10802 VDD.n3990 VSS 0.00202f
C10803 VDD.n3991 VSS 0.0027f
C10804 VDD.n3992 VSS 0.00308f
C10805 VDD.n3993 VSS 0.00183f
C10806 VDD.n3994 VSS 0.00151f
C10807 VDD.n3995 VSS 0.00109f
C10808 VDD.n3996 VSS 0.00773f
C10809 VDD.n3997 VSS 0.00109f
C10810 VDD.n3998 VSS 0.0018f
C10811 VDD.n3999 VSS 0.00231f
C10812 VDD.t446 VSS -2.71e-19
C10813 VDD.t280 VSS 8.49e-19
C10814 VDD.n4000 VSS 0.00391f
C10815 VDD.n4001 VSS 0.00413f
C10816 VDD.t445 VSS 0.00578f
C10817 VDD.n4002 VSS 0.00597f
C10818 VDD.n4003 VSS 0.00109f
C10819 VDD.n4004 VSS 9.92e-19
C10820 VDD.n4005 VSS 0.00308f
C10821 VDD.t279 VSS 0.00578f
C10822 VDD.n4006 VSS 0.00835f
C10823 VDD.n4007 VSS 0.00109f
C10824 VDD.n4008 VSS 0.00186f
C10825 VDD.n4009 VSS 0.00308f
C10826 VDD.t277 VSS 0.00955f
C10827 VDD.n4010 VSS 0.00923f
C10828 VDD.n4011 VSS 6.76e-19
C10829 VDD.n4012 VSS 0.00179f
C10830 VDD.n4013 VSS 0.00308f
C10831 VDD.t278 VSS -5.07e-19
C10832 VDD.t143 VSS 9.16e-19
C10833 VDD.n4014 VSS 0.00359f
C10834 VDD.n4015 VSS 0.00204f
C10835 VDD.n4016 VSS 0.00187f
C10836 VDD.n4017 VSS 0.00281f
C10837 VDD.n4018 VSS 0.00154f
C10838 VDD.t757 VSS 8.67e-19
C10839 VDD.n4019 VSS 0.00281f
C10840 VDD.t141 VSS 0.0016f
C10841 VDD.n4020 VSS 0.00355f
C10842 VDD.n4021 VSS 7.59e-19
C10843 VDD.n4022 VSS 0.00215f
C10844 VDD.n4023 VSS 3.97e-19
C10845 VDD.n4024 VSS 2.85e-19
C10846 VDD.n4025 VSS 0.00154f
C10847 VDD.t699 VSS 0.00262f
C10848 VDD.n4026 VSS 0.00271f
C10849 VDD.t142 VSS 0.0139f
C10850 VDD.n4027 VSS 0.0119f
C10851 VDD.n4028 VSS 9.48e-19
C10852 VDD.n4029 VSS 0.00267f
C10853 VDD.n4030 VSS 0.00307f
C10854 VDD.t698 VSS 0.00578f
C10855 VDD.t705 VSS 0.00578f
C10856 VDD.n4031 VSS 0.00452f
C10857 VDD.n4032 VSS 0.00109f
C10858 VDD.n4033 VSS 0.00172f
C10859 VDD.n4034 VSS 0.00308f
C10860 VDD.n4035 VSS 0.00666f
C10861 VDD.n4036 VSS 0.00109f
C10862 VDD.n4037 VSS 0.00164f
C10863 VDD.n4038 VSS 0.00308f
C10864 VDD.t505 VSS 5.72e-19
C10865 VDD.t276 VSS 7.62e-19
C10866 VDD.n4039 VSS 0.0014f
C10867 VDD.t504 VSS 0.00578f
C10868 VDD.n4040 VSS 0.0076f
C10869 VDD.n4041 VSS 0.00111f
C10870 VDD.n4042 VSS 0.00204f
C10871 VDD.n4043 VSS 0.00252f
C10872 VDD.n4044 VSS 0.00308f
C10873 VDD.t275 VSS 0.00578f
C10874 VDD.n4045 VSS 0.00603f
C10875 VDD.n4046 VSS 0.00109f
C10876 VDD.n4047 VSS 0.00132f
C10877 VDD.n4048 VSS 0.00308f
C10878 VDD.t552 VSS 0.00578f
C10879 VDD.n4049 VSS 0.00634f
C10880 VDD.n4050 VSS 0.00109f
C10881 VDD.n4051 VSS 0.00186f
C10882 VDD.n4052 VSS 0.00308f
C10883 VDD.t725 VSS 0.00578f
C10884 VDD.n4053 VSS 0.00528f
C10885 VDD.n4054 VSS 0.00109f
C10886 VDD.n4055 VSS 0.00186f
C10887 VDD.n4056 VSS 0.00308f
C10888 VDD.n4057 VSS 0.00905f
C10889 VDD.n4058 VSS 0.00109f
C10890 VDD.n4059 VSS 0.00186f
C10891 VDD.n4060 VSS 0.00308f
C10892 VDD.t614 VSS 0.00578f
C10893 VDD.n4061 VSS 0.00823f
C10894 VDD.n4062 VSS 0.00109f
C10895 VDD.n4063 VSS 0.0011f
C10896 VDD.n4064 VSS 0.00308f
C10897 VDD.t615 VSS 0.00217f
C10898 VDD.t701 VSS 9.67e-19
C10899 VDD.n4065 VSS 0.00349f
C10900 VDD.n4066 VSS 0.00457f
C10901 VDD.t700 VSS 0.00565f
C10902 VDD.n4067 VSS 0.00616f
C10903 VDD.n4068 VSS 0.00109f
C10904 VDD.n4069 VSS 8.8e-19
C10905 VDD.n4070 VSS 0.00241f
C10906 VDD.n4071 VSS 9.21e-19
C10907 VDD.n4072 VSS 0.00154f
C10908 VDD.n4073 VSS 9.31e-19
C10909 VDD.t82 VSS 0.0054f
C10910 VDD.n4074 VSS 0.0059f
C10911 VDD.n4075 VSS 0.00109f
C10912 VDD.n4076 VSS 1.72e-19
C10913 VDD.n4077 VSS 2.85e-19
C10914 VDD.n4078 VSS 9.31e-19
C10915 VDD.n4079 VSS 6.2e-19
C10916 VDD.n4080 VSS 4.35e-19
C10917 VDD.n4081 VSS 3.36e-19
C10918 VDD.n4082 VSS 8.1e-19
C10919 VDD.n4083 VSS 0.00148f
C10920 VDD.n4084 VSS 6.16e-19
C10921 VDD.n4085 VSS 0.00158f
C10922 VDD.n4086 VSS 2.97e-19
C10923 VDD.n4087 VSS 3.23e-19
C10924 VDD.t28 VSS 0.00578f
C10925 VDD.n4088 VSS 0.00666f
C10926 VDD.n4089 VSS 0.00109f
C10927 VDD.n4090 VSS 0.00115f
C10928 VDD.n4091 VSS 0.00275f
C10929 VDD.n4092 VSS 0.00154f
C10930 VDD.t29 VSS 5.72e-19
C10931 VDD.t613 VSS 5.42e-19
C10932 VDD.n4093 VSS 0.00119f
C10933 VDD.t612 VSS 0.00578f
C10934 VDD.n4094 VSS 0.00666f
C10935 VDD.n4095 VSS 0.00111f
C10936 VDD.n4096 VSS 0.00203f
C10937 VDD.n4097 VSS 0.00279f
C10938 VDD.n4098 VSS 4.19e-19
C10939 VDD.n4099 VSS 0.00754f
C10940 VDD.n4100 VSS 0.00109f
C10941 VDD.n4101 VSS 0.00162f
C10942 VDD.n4102 VSS 0.0024f
C10943 VDD.n4103 VSS 0.00141f
C10944 VDD.n4104 VSS 4.35e-19
C10945 VDD.n4105 VSS 4.94e-19
C10946 VDD.n4106 VSS 3.36e-19
C10947 VDD.n4107 VSS 8.1e-19
C10948 VDD.n4108 VSS 0.00148f
C10949 VDD.n4109 VSS 0.00492f
C10950 VDD.n4110 VSS 0.00553f
C10951 VDD.n4111 VSS 0.00123f
C10952 VDD.n4112 VSS 6.15e-19
C10953 VDD.n4113 VSS 0.128f
C10954 VDD.n4114 VSS 0.128f
C10955 VDD.n4115 VSS 6.15e-19
C10956 VDD.n4116 VSS 0.00102f
C10957 VDD.n4117 VSS 0.00553f
C10958 VDD.n4118 VSS 0.00149f
C10959 VDD.n4119 VSS 5.46e-19
C10960 VDD.n4120 VSS 5.66e-19
C10961 VDD.t198 VSS 0.00579f
C10962 VDD.t728 VSS 0.00579f
C10963 VDD.n4121 VSS 0.00453f
C10964 VDD.n4122 VSS 0.00109f
C10965 VDD.n4123 VSS 0.00119f
C10966 VDD.n4124 VSS 0.00236f
C10967 VDD.t729 VSS 0.00265f
C10968 VDD.n4125 VSS 0.00411f
C10969 VDD.n4126 VSS 0.00863f
C10970 VDD.n4127 VSS 9.9e-19
C10971 VDD.n4128 VSS 0.00143f
C10972 VDD.n4129 VSS 5.17e-19
C10973 VDD.n4130 VSS 0.0026f
C10974 VDD.n4131 VSS 0.00129f
C10975 VDD.n4132 VSS 4.35e-19
C10976 VDD.n4133 VSS 9.47e-19
C10977 VDD.n4134 VSS 2.68e-19
C10978 VDD.n4135 VSS 7.11e-19
C10979 VDD.n4136 VSS 0.00926f
C10980 VDD.n4137 VSS 0.00101f
C10981 VDD.n4138 VSS 1.75e-19
C10982 VDD.n4139 VSS 2.85e-19
C10983 VDD.n4140 VSS 0.00151f
C10984 VDD.n4141 VSS 0.00132f
C10985 VDD.n4142 VSS 0.00172f
C10986 VDD.t3 VSS 9.16e-19
C10987 VDD.t309 VSS -5.07e-19
C10988 VDD.n4143 VSS 0.00359f
C10989 VDD.n4144 VSS 6.49e-19
C10990 VDD.n4145 VSS 0.00127f
C10991 VDD.n4146 VSS 4e-19
C10992 VDD.n4147 VSS 5.43e-19
C10993 VDD.n4148 VSS 1.04e-19
C10994 VDD.t308 VSS 0.0046f
C10995 VDD.n4149 VSS 0.00214f
C10996 VDD.n4150 VSS 0.00107f
C10997 VDD.n4151 VSS 0.00397f
C10998 VDD.n4152 VSS 5.98e-19
C10999 VDD.n4153 VSS 7.05e-20
C11000 VDD.n4154 VSS 1.65e-19
C11001 VDD.n4155 VSS 2.85e-19
C11002 VDD.n4156 VSS 0.00131f
C11003 VDD.n4157 VSS 0.00129f
C11004 VDD.n4158 VSS 2.85e-19
C11005 VDD.n4159 VSS 0.00137f
C11006 VDD.n4160 VSS 4e-19
C11007 VDD.n4161 VSS 0.00181f
C11008 VDD.n4162 VSS 4e-19
C11009 VDD.n4163 VSS 5.2e-19
C11010 VDD.n4164 VSS 1.04e-19
C11011 VDD.n4165 VSS 0.00535f
C11012 VDD.n4166 VSS 0.00107f
C11013 VDD.t2 VSS 0.00611f
C11014 VDD.n4167 VSS 0.00246f
C11015 VDD.n4168 VSS 6.17e-19
C11016 VDD.n4169 VSS 1.65e-19
C11017 VDD.n4170 VSS 2.51e-19
C11018 VDD.n4171 VSS 4.35e-19
C11019 VDD.n4172 VSS 3.36e-19
C11020 VDD.n4173 VSS 8.1e-19
C11021 VDD.n4174 VSS 0.00157f
C11022 VDD.n4175 VSS 0.00512f
C11023 VDD.n4176 VSS 0.00158f
C11024 VDD.n4177 VSS 6.17e-19
C11025 VDD.n4178 VSS 0.00127f
C11026 VDD.t304 VSS 0.00579f
C11027 VDD.n4179 VSS 0.00838f
C11028 VDD.n4180 VSS 0.00112f
C11029 VDD.n4181 VSS 0.00185f
C11030 VDD.n4182 VSS 0.00258f
C11031 VDD.t305 VSS 8.49e-19
C11032 VDD.t358 VSS -2.71e-19
C11033 VDD.n4183 VSS 0.00391f
C11034 VDD.n4184 VSS 0.00405f
C11035 VDD.t357 VSS 0.00665f
C11036 VDD.n4185 VSS 0.00598f
C11037 VDD.n4186 VSS 0.00112f
C11038 VDD.n4187 VSS 0.00101f
C11039 VDD.n4188 VSS 0.0025f
C11040 VDD.n4189 VSS 0.00109f
C11041 VDD.n4190 VSS 0.0139f
C11042 VDD.n4191 VSS 9.04e-19
C11043 VDD.n4192 VSS 0.001f
C11044 VDD.n4193 VSS 8.85e-19
C11045 VDD.n4194 VSS 5.19e-19
C11046 VDD.n4195 VSS 4.35e-19
C11047 VDD.n4196 VSS 4.94e-19
C11048 VDD.n4197 VSS 3.36e-19
C11049 VDD.n4198 VSS 8.1e-19
C11050 VDD.n4199 VSS 0.00148f
C11051 VDD.n4200 VSS 0.00149f
C11052 VDD.n4201 VSS 5.71e-19
C11053 VDD.n4202 VSS 5.41e-19
C11054 VDD.n4203 VSS 3.36e-19
C11055 VDD.n4204 VSS 8.14e-19
C11056 VDD.n4205 VSS 0.00157f
C11057 VDD.n4206 VSS 0.0842f
C11058 VDD.n4207 VSS 6.15e-19
C11059 VDD.n4208 VSS 0.00512f
C11060 VDD.n4209 VSS 0.00553f
C11061 VDD.n4210 VSS 0.00144f
C11062 VDD.n4211 VSS 0.00148f
C11063 VDD.n4212 VSS 8.1e-19
C11064 VDD.n4213 VSS 0.00157f
C11065 VDD.n4214 VSS 0.00103f
C11066 VDD.n4215 VSS 6.16e-19
C11067 VDD.n4216 VSS 0.00157f
C11068 VDD.n4217 VSS 0.00149f
C11069 VDD.n4218 VSS 8.1e-19
C11070 VDD.n4219 VSS 3.36e-19
C11071 VDD.n4220 VSS 4.35e-19
C11072 VDD.n4221 VSS 3.85e-19
C11073 VDD.n4222 VSS 1.84e-19
C11074 VDD.n4223 VSS 9.31e-19
C11075 VDD.t306 VSS 0.00579f
C11076 VDD.n4224 VSS 0.00605f
C11077 VDD.n4225 VSS 0.00109f
C11078 VDD.n4226 VSS 1.72e-19
C11079 VDD.n4227 VSS 2.85e-19
C11080 VDD.n4228 VSS 0.00154f
C11081 VDD.t733 VSS 0.00579f
C11082 VDD.n4229 VSS 0.00636f
C11083 VDD.n4230 VSS 0.00109f
C11084 VDD.n4231 VSS 0.0017f
C11085 VDD.n4232 VSS 0.00281f
C11086 VDD.t473 VSS 0.00579f
C11087 VDD.n4233 VSS 0.00529f
C11088 VDD.n4234 VSS 0.00109f
C11089 VDD.n4235 VSS 0.00186f
C11090 VDD.n4236 VSS 0.00308f
C11091 VDD.n4237 VSS 0.00907f
C11092 VDD.n4238 VSS 0.00109f
C11093 VDD.n4239 VSS 0.00186f
C11094 VDD.n4240 VSS 0.00308f
C11095 VDD.t454 VSS 0.00579f
C11096 VDD.n4241 VSS 0.00825f
C11097 VDD.n4242 VSS 0.00109f
C11098 VDD.n4243 VSS 0.0011f
C11099 VDD.n4244 VSS 0.00308f
C11100 VDD.t727 VSS 9.67e-19
C11101 VDD.t455 VSS 0.00217f
C11102 VDD.n4245 VSS 0.00349f
C11103 VDD.n4246 VSS 0.00457f
C11104 VDD.t726 VSS 0.00567f
C11105 VDD.n4247 VSS 0.00617f
C11106 VDD.n4248 VSS 0.00109f
C11107 VDD.n4249 VSS 0.00102f
C11108 VDD.n4250 VSS 0.00308f
C11109 VDD.t145 VSS 0.0134f
C11110 VDD.t400 VSS 0.00542f
C11111 VDD.n4251 VSS 0.0068f
C11112 VDD.n4252 VSS 0.00103f
C11113 VDD.n4253 VSS 0.00176f
C11114 VDD.n4254 VSS 0.00291f
C11115 VDD.n4255 VSS 0.00154f
C11116 VDD.n4256 VSS 1.36e-19
C11117 VDD.t126 VSS 0.00149f
C11118 VDD.t761 VSS 6.37e-19
C11119 VDD.n4257 VSS 0.00279f
C11120 VDD.n4258 VSS 2.33e-19
C11121 VDD.n4259 VSS 6.77e-19
C11122 VDD.n4260 VSS 0.00141f
C11123 VDD.n4261 VSS 2.33e-19
C11124 VDD.n4262 VSS 0.00388f
C11125 VDD.n4263 VSS 5.31e-19
C11126 VDD.n4264 VSS 0.00105f
C11127 VDD.t771 VSS 6.29e-19
C11128 VDD.n4265 VSS 0.00315f
C11129 VDD.t144 VSS 0.00189f
C11130 VDD.n4266 VSS 0.00174f
C11131 VDD.n4267 VSS 2.32e-19
C11132 VDD.n4268 VSS 9.31e-19
C11133 VDD.n4269 VSS 1.72e-19
C11134 VDD.n4270 VSS 2.85e-19
C11135 VDD.n4271 VSS 0.00146f
C11136 VDD.n4272 VSS 0.00198f
C11137 VDD.t457 VSS 5.42e-19
C11138 VDD.t146 VSS 5.72e-19
C11139 VDD.n4273 VSS 0.00119f
C11140 VDD.n4274 VSS 0.00282f
C11141 VDD.n4275 VSS 0.00296f
C11142 VDD.t456 VSS 0.0107f
C11143 VDD.n4276 VSS 0.00756f
C11144 VDD.n4277 VSS 0.00103f
C11145 VDD.n4278 VSS 0.00177f
C11146 VDD.n4279 VSS 0.00308f
C11147 VDD.t474 VSS 0.00579f
C11148 VDD.n4280 VSS 0.00529f
C11149 VDD.n4281 VSS 0.00109f
C11150 VDD.n4282 VSS 0.00186f
C11151 VDD.n4283 VSS 0.00308f
C11152 VDD.t730 VSS 0.00579f
C11153 VDD.n4284 VSS 0.00579f
C11154 VDD.n4285 VSS 0.00109f
C11155 VDD.n4286 VSS 0.00151f
C11156 VDD.n4287 VSS 0.00308f
C11157 VDD.n4288 VSS 0.00308f
C11158 VDD.n4289 VSS 0.00907f
C11159 VDD.n4290 VSS 0.00109f
C11160 VDD.n4291 VSS 0.00118f
C11161 VDD.n4292 VSS 0.00308f
C11162 VDD.n4293 VSS 0.0028f
C11163 VDD.n4294 VSS 0.00106f
C11164 VDD.n4295 VSS 0.00151f
C11165 VDD.n4296 VSS 0.00109f
C11166 VDD.n4297 VSS 0.00882f
C11167 VDD.n4298 VSS 0.00109f
C11168 VDD.n4299 VSS 0.0018f
C11169 VDD.n4300 VSS 0.00231f
C11170 VDD.t214 VSS 8.49e-19
C11171 VDD.t360 VSS -2.71e-19
C11172 VDD.n4301 VSS 0.00391f
C11173 VDD.n4302 VSS 0.00413f
C11174 VDD.t359 VSS 0.00579f
C11175 VDD.n4303 VSS 0.00598f
C11176 VDD.n4304 VSS 0.00109f
C11177 VDD.n4305 VSS 9.92e-19
C11178 VDD.n4306 VSS 0.00308f
C11179 VDD.t213 VSS 0.00579f
C11180 VDD.n4307 VSS 0.00838f
C11181 VDD.n4308 VSS 0.00109f
C11182 VDD.n4309 VSS 0.00171f
C11183 VDD.n4310 VSS 0.0024f
C11184 VDD.n4311 VSS 9.04e-19
C11185 VDD.n4312 VSS 4.35e-19
C11186 VDD.n4313 VSS 3.36e-19
C11187 VDD.n4314 VSS 8.1e-19
C11188 VDD.n4315 VSS 0.00148f
C11189 VDD.n4316 VSS 0.0984f
C11190 VDD.n4317 VSS 0.00193f
C11191 VDD.n4318 VSS 0.00653f
C11192 VDD.n4319 VSS 0.00158f
C11193 VDD.n4320 VSS 6.17e-19
C11194 VDD.t254 VSS 0.00579f
C11195 VDD.n4321 VSS 0.00529f
C11196 VDD.n4322 VSS 0.00109f
C11197 VDD.n4323 VSS 0.00186f
C11198 VDD.n4324 VSS 0.00231f
C11199 VDD.t86 VSS 0.00579f
C11200 VDD.n4325 VSS 0.00636f
C11201 VDD.n4326 VSS 0.00109f
C11202 VDD.n4327 VSS 0.00186f
C11203 VDD.n4328 VSS 0.00308f
C11204 VDD.t211 VSS 0.00579f
C11205 VDD.n4329 VSS 0.00605f
C11206 VDD.n4330 VSS 0.00109f
C11207 VDD.n4331 VSS 0.00132f
C11208 VDD.n4332 VSS 0.0025f
C11209 VDD.n4333 VSS 0.00109f
C11210 VDD.n4334 VSS 0.00154f
C11211 VDD.n4335 VSS 2.85e-19
C11212 VDD.t124 VSS 0.00579f
C11213 VDD.n4336 VSS 0.00762f
C11214 VDD.n4337 VSS 0.00111f
C11215 VDD.n4338 VSS 0.00201f
C11216 VDD.t212 VSS 7.62e-19
C11217 VDD.t125 VSS 5.72e-19
C11218 VDD.n4339 VSS 0.00139f
C11219 VDD.n4340 VSS 0.00235f
C11220 VDD.n4341 VSS 2.25e-19
C11221 VDD.n4342 VSS 4.52e-19
C11222 VDD.n4343 VSS 4.35e-19
C11223 VDD.n4344 VSS 4.94e-19
C11224 VDD.n4345 VSS 3.36e-19
C11225 VDD.n4346 VSS 8.1e-19
C11226 VDD.n4347 VSS 0.00148f
C11227 VDD.n4348 VSS 4.69e-19
C11228 VDD.n4349 VSS 0.00154f
C11229 VDD.n4350 VSS 0.00203f
C11230 VDD.n4351 VSS 3.74e-19
C11231 VDD.n4352 VSS 1.17e-19
C11232 VDD.n4353 VSS 5.4e-19
C11233 VDD.n4354 VSS 1.01e-19
C11234 VDD.n4355 VSS 0.00573f
C11235 VDD.n4356 VSS 0.00107f
C11236 VDD.t592 VSS 0.00466f
C11237 VDD.n4357 VSS 0.00208f
C11238 VDD.n4358 VSS 4.45e-19
C11239 VDD.n4359 VSS 3.04e-19
C11240 VDD.n4360 VSS 2.85e-19
C11241 VDD.n4361 VSS 0.00145f
C11242 VDD.n4362 VSS 3.97e-19
C11243 VDD.n4363 VSS 2.85e-19
C11244 VDD.n4364 VSS 3.35e-19
C11245 VDD.n4365 VSS 0.00151f
C11246 VDD.n4366 VSS 0.00164f
C11247 VDD.t593 VSS 9.16e-19
C11248 VDD.t210 VSS -5.07e-19
C11249 VDD.n4367 VSS 0.00359f
C11250 VDD.n4368 VSS 6.69e-19
C11251 VDD.n4369 VSS 9.35e-20
C11252 VDD.n4370 VSS 5.34e-19
C11253 VDD.n4371 VSS 1.01e-19
C11254 VDD.n4372 VSS 0.00365f
C11255 VDD.n4373 VSS 0.00107f
C11256 VDD.t209 VSS 0.00586f
C11257 VDD.n4374 VSS 0.00246f
C11258 VDD.n4375 VSS 5.58e-19
C11259 VDD.n4376 VSS 4.68e-20
C11260 VDD.n4377 VSS 0.00149f
C11261 VDD.n4378 VSS 3.97e-19
C11262 VDD.n4379 VSS 2.85e-19
C11263 VDD.n4380 VSS 9.04e-19
C11264 VDD.n4381 VSS 9.88e-19
C11265 VDD.n4382 VSS 3.52e-19
C11266 VDD.n4383 VSS 6.43e-19
C11267 VDD.n4384 VSS 3.36e-19
C11268 VDD.n4385 VSS 0.00149f
C11269 VDD.n4386 VSS 8.1e-19
C11270 VDD.n4387 VSS 0.00157f
C11271 VDD.n4388 VSS 0.00605f
C11272 VDD.n4389 VSS 0.00158f
C11273 VDD.n4390 VSS 3.36e-19
C11274 VDD.n4391 VSS 3.1e-19
C11275 VDD.n4392 VSS 4.82e-19
C11276 VDD.n4393 VSS 0.00668f
C11277 VDD.n4394 VSS 0.00109f
C11278 VDD.n4395 VSS 0.00164f
C11279 VDD.n4396 VSS 0.00265f
C11280 VDD.n4397 VSS 0.00154f
C11281 VDD.t734 VSS 0.00579f
C11282 VDD.t621 VSS 0.00579f
C11283 VDD.n4398 VSS 0.00453f
C11284 VDD.n4399 VSS 0.00109f
C11285 VDD.n4400 VSS 0.00172f
C11286 VDD.n4401 VSS 4.02e-19
C11287 VDD.t622 VSS 0.00262f
C11288 VDD.n4402 VSS 0.00271f
C11289 VDD.n4403 VSS 0.00882f
C11290 VDD.n4404 VSS 9.91e-19
C11291 VDD.n4405 VSS 0.00229f
C11292 VDD.n4406 VSS 0.00258f
C11293 VDD.n4407 VSS 0.00144f
C11294 VDD.n4408 VSS 4.19e-19
C11295 VDD.n4409 VSS 3.23e-19
C11296 VDD.n4410 VSS 8.1e-19
C11297 VDD.n4411 VSS 0.00148f
C11298 VDD.n4412 VSS 0.00149f
C11299 VDD.n4413 VSS 8.1e-19
C11300 VDD.n4414 VSS 0.00144f
C11301 VDD.n4415 VSS 0.00157f
C11302 VDD.n4416 VSS 0.00194f
C11303 VDD.n4417 VSS 0.00653f
C11304 VDD.n4418 VSS 0.00148f
C11305 VDD.n4419 VSS 8.1e-19
C11306 VDD.n4420 VSS 3.23e-19
C11307 VDD.n4421 VSS 4.19e-19
C11308 VDD.t620 VSS 9.67e-19
C11309 VDD.t387 VSS 0.00217f
C11310 VDD.n4422 VSS 0.00349f
C11311 VDD.n4423 VSS 0.00457f
C11312 VDD.t619 VSS 0.00567f
C11313 VDD.n4424 VSS 0.00617f
C11314 VDD.n4425 VSS 0.00109f
C11315 VDD.n4426 VSS 0.00102f
C11316 VDD.n4427 VSS 4.02e-19
C11317 VDD.n4428 VSS 0.00154f
C11318 VDD.t103 VSS 0.0134f
C11319 VDD.t243 VSS 0.00542f
C11320 VDD.n4429 VSS 0.0068f
C11321 VDD.n4430 VSS 0.00108f
C11322 VDD.n4431 VSS 0.00176f
C11323 VDD.n4432 VSS 0.00261f
C11324 VDD.n4433 VSS 0.00154f
C11325 VDD.n4434 VSS 1.36e-19
C11326 VDD.t123 VSS 0.00149f
C11327 VDD.t762 VSS 6.37e-19
C11328 VDD.n4435 VSS 0.00279f
C11329 VDD.n4436 VSS 2.33e-19
C11330 VDD.n4437 VSS 6.77e-19
C11331 VDD.n4438 VSS 0.00141f
C11332 VDD.n4439 VSS 2.33e-19
C11333 VDD.n4440 VSS 0.00388f
C11334 VDD.n4441 VSS 5.31e-19
C11335 VDD.n4442 VSS 0.00105f
C11336 VDD.t764 VSS 6.29e-19
C11337 VDD.n4443 VSS 0.00315f
C11338 VDD.t102 VSS 0.00189f
C11339 VDD.n4444 VSS 0.00174f
C11340 VDD.n4445 VSS 2.32e-19
C11341 VDD.n4446 VSS 9.31e-19
C11342 VDD.n4447 VSS 1.72e-19
C11343 VDD.n4448 VSS 2.85e-19
C11344 VDD.n4449 VSS 0.00146f
C11345 VDD.n4450 VSS 0.00198f
C11346 VDD.t389 VSS 5.42e-19
C11347 VDD.t104 VSS 5.72e-19
C11348 VDD.n4451 VSS 0.00119f
C11349 VDD.n4452 VSS 0.00282f
C11350 VDD.n4453 VSS 0.00296f
C11351 VDD.t388 VSS 0.0107f
C11352 VDD.n4454 VSS 0.00756f
C11353 VDD.n4455 VSS 0.00103f
C11354 VDD.n4456 VSS 0.00177f
C11355 VDD.n4457 VSS 0.00308f
C11356 VDD.t253 VSS 0.00579f
C11357 VDD.n4458 VSS 0.00529f
C11358 VDD.n4459 VSS 0.00109f
C11359 VDD.n4460 VSS 0.00186f
C11360 VDD.n4461 VSS 0.00308f
C11361 VDD.t85 VSS 0.00579f
C11362 VDD.n4462 VSS 0.00579f
C11363 VDD.n4463 VSS 0.00109f
C11364 VDD.n4464 VSS 0.00151f
C11365 VDD.n4465 VSS 0.00308f
C11366 VDD.n4466 VSS 0.00308f
C11367 VDD.n4467 VSS 0.00907f
C11368 VDD.n4468 VSS 0.00109f
C11369 VDD.n4469 VSS 0.00118f
C11370 VDD.n4470 VSS 0.00308f
C11371 VDD.n4471 VSS 0.0028f
C11372 VDD.n4472 VSS 0.00106f
C11373 VDD.n4473 VSS 0.00151f
C11374 VDD.n4474 VSS 0.00109f
C11375 VDD.n4475 VSS 0.00882f
C11376 VDD.n4476 VSS 0.00109f
C11377 VDD.n4477 VSS 0.0018f
C11378 VDD.n4478 VSS 0.00231f
C11379 VDD.t65 VSS 8.49e-19
C11380 VDD.t53 VSS -2.71e-19
C11381 VDD.n4479 VSS 0.00391f
C11382 VDD.n4480 VSS 0.00413f
C11383 VDD.t52 VSS 0.00579f
C11384 VDD.n4481 VSS 0.00598f
C11385 VDD.n4482 VSS 0.00109f
C11386 VDD.n4483 VSS 9.92e-19
C11387 VDD.n4484 VSS 0.00308f
C11388 VDD.t64 VSS 0.00579f
C11389 VDD.n4485 VSS 0.00838f
C11390 VDD.n4486 VSS 0.00109f
C11391 VDD.n4487 VSS 0.00186f
C11392 VDD.n4488 VSS 0.00308f
C11393 VDD.n4489 VSS 0.00926f
C11394 VDD.n4490 VSS 9.85e-19
C11395 VDD.n4491 VSS 0.00163f
C11396 VDD.n4492 VSS 0.00307f
C11397 VDD.n4493 VSS 0.00154f
C11398 VDD.n4494 VSS 0.00203f
C11399 VDD.t31 VSS 9.16e-19
C11400 VDD.t63 VSS -5.07e-19
C11401 VDD.n4495 VSS 0.00359f
C11402 VDD.n4496 VSS 6.69e-19
C11403 VDD.n4497 VSS 0.00143f
C11404 VDD.n4498 VSS 3.97e-19
C11405 VDD.n4499 VSS 5.34e-19
C11406 VDD.n4500 VSS 1.01e-19
C11407 VDD.t62 VSS 0.00466f
C11408 VDD.n4501 VSS 0.0022f
C11409 VDD.n4502 VSS 0.00107f
C11410 VDD.n4503 VSS 0.0039f
C11411 VDD.n4504 VSS 5.58e-19
C11412 VDD.n4505 VSS 4.68e-20
C11413 VDD.n4506 VSS 1.4e-19
C11414 VDD.n4507 VSS 2.85e-19
C11415 VDD.n4508 VSS 0.00154f
C11416 VDD.t30 VSS 0.00586f
C11417 VDD.n4509 VSS 0.00781f
C11418 VDD.n4510 VSS 0.0011f
C11419 VDD.n4511 VSS 0.00393f
C11420 VDD.n4512 VSS 0.00281f
C11421 VDD.t494 VSS 0.00262f
C11422 VDD.n4513 VSS 0.00271f
C11423 VDD.n4514 VSS 0.00989f
C11424 VDD.n4515 VSS 0.00109f
C11425 VDD.n4516 VSS 0.00269f
C11426 VDD.n4517 VSS 0.00308f
C11427 VDD.t377 VSS 0.00579f
C11428 VDD.t493 VSS 0.00579f
C11429 VDD.n4518 VSS 0.00453f
C11430 VDD.n4519 VSS 0.00109f
C11431 VDD.n4520 VSS 0.00172f
C11432 VDD.n4521 VSS 0.00308f
C11433 VDD.n4522 VSS 0.00668f
C11434 VDD.n4523 VSS 0.00109f
C11435 VDD.n4524 VSS 0.00164f
C11436 VDD.n4525 VSS 0.00298f
C11437 VDD.n4526 VSS 0.00154f
C11438 VDD.n4527 VSS 2.85e-19
C11439 VDD.t133 VSS 0.00579f
C11440 VDD.n4528 VSS 0.00762f
C11441 VDD.n4529 VSS 0.00111f
C11442 VDD.n4530 VSS 0.00201f
C11443 VDD.t61 VSS 7.62e-19
C11444 VDD.t134 VSS 5.72e-19
C11445 VDD.n4531 VSS 0.00139f
C11446 VDD.n4532 VSS 0.00235f
C11447 VDD.n4533 VSS 2.25e-19
C11448 VDD.n4534 VSS 5.36e-19
C11449 VDD.n4535 VSS 4.35e-19
C11450 VDD.n4536 VSS 4.56e-19
C11451 VDD.n4537 VSS 3.36e-19
C11452 VDD.n4538 VSS 8.1e-19
C11453 VDD.n4539 VSS 0.00148f
C11454 VDD.n4540 VSS 0.0991f
C11455 VDD.n4541 VSS 9.67e-19
C11456 VDD.n4542 VSS 0.00121f
C11457 VDD.n4543 VSS 0.0058f
C11458 VDD.n4544 VSS 0.00149f
C11459 VDD.n4545 VSS 4.44e-19
C11460 VDD.n4546 VSS 6.68e-19
C11461 VDD.n4547 VSS 3.36e-19
C11462 VDD.n4548 VSS 8.12e-19
C11463 VDD.n4549 VSS 0.00157f
C11464 VDD.n4550 VSS 0.00556f
C11465 VDD.n4551 VSS 9.68e-19
C11466 VDD.n4552 VSS 6.6e-19
C11467 VDD.t121 VSS 0.0134f
C11468 VDD.t458 VSS 0.00542f
C11469 VDD.n4553 VSS 0.0068f
C11470 VDD.n4554 VSS 0.00115f
C11471 VDD.n4555 VSS 0.00165f
C11472 VDD.n4556 VSS 0.00229f
C11473 VDD.n4557 VSS 0.00101f
C11474 VDD.n4558 VSS 9.38e-19
C11475 VDD.n4559 VSS 4.35e-19
C11476 VDD.n4560 VSS 9.31e-19
C11477 VDD.n4561 VSS 6.03e-19
C11478 VDD.n4562 VSS 9.31e-19
C11479 VDD.n4563 VSS 0.00907f
C11480 VDD.n4564 VSS 0.00109f
C11481 VDD.n4565 VSS 1.72e-19
C11482 VDD.n4566 VSS 2.85e-19
C11483 VDD.n4567 VSS 0.00154f
C11484 VDD.t749 VSS 0.00579f
C11485 VDD.n4568 VSS 0.00825f
C11486 VDD.n4569 VSS 0.00109f
C11487 VDD.n4570 VSS 0.00107f
C11488 VDD.n4571 VSS 0.00293f
C11489 VDD.n4572 VSS 0.00154f
C11490 VDD.t491 VSS 0.00567f
C11491 VDD.n4573 VSS 0.00617f
C11492 VDD.n4574 VSS 0.00109f
C11493 VDD.t492 VSS 9.67e-19
C11494 VDD.t750 VSS 0.00217f
C11495 VDD.n4575 VSS 0.00349f
C11496 VDD.n4576 VSS 0.0045f
C11497 VDD.n4577 VSS 9.11e-20
C11498 VDD.n4578 VSS 1.72e-19
C11499 VDD.n4579 VSS 2.85e-19
C11500 VDD.n4580 VSS 9.31e-19
C11501 VDD.n4581 VSS 5.36e-19
C11502 VDD.n4582 VSS 4.35e-19
C11503 VDD.n4583 VSS 4.52e-19
C11504 VDD.n4584 VSS 3.36e-19
C11505 VDD.n4585 VSS 0.00149f
C11506 VDD.n4586 VSS 8.1e-19
C11507 VDD.n4587 VSS 0.00157f
C11508 VDD.n4588 VSS 9.68e-19
C11509 VDD.n4589 VSS 0.00121f
C11510 VDD.n4590 VSS 0.00148f
C11511 VDD.n4591 VSS 8.1e-19
C11512 VDD.n4592 VSS 5.07e-19
C11513 VDD.n4593 VSS 3.36e-19
C11514 VDD.n4594 VSS 4.35e-19
C11515 VDD.n4595 VSS 9.31e-19
C11516 VDD.n4596 VSS 1.68e-19
C11517 VDD.n4597 VSS 9.31e-19
C11518 VDD.t451 VSS 0.00579f
C11519 VDD.n4598 VSS 0.00529f
C11520 VDD.n4599 VSS 0.00109f
C11521 VDD.n4600 VSS 1.72e-19
C11522 VDD.n4601 VSS 2.85e-19
C11523 VDD.n4602 VSS 0.00154f
C11524 VDD.t223 VSS 0.00579f
C11525 VDD.n4603 VSS 0.00579f
C11526 VDD.n4604 VSS 0.00109f
C11527 VDD.n4605 VSS 0.00135f
C11528 VDD.n4606 VSS 0.00281f
C11529 VDD.t572 VSS 0.00142f
C11530 VDD.t571 VSS 0.00579f
C11531 VDD.n4607 VSS 0.00857f
C11532 VDD.n4608 VSS 0.00111f
C11533 VDD.n4609 VSS 0.00203f
C11534 VDD.n4610 VSS 0.00312f
C11535 VDD.n4611 VSS 0.00308f
C11536 VDD.n4612 VSS 0.00907f
C11537 VDD.n4613 VSS 0.00109f
C11538 VDD.n4614 VSS 0.00118f
C11539 VDD.n4615 VSS 0.00308f
C11540 VDD.t548 VSS 6.03e-19
C11541 VDD.t222 VSS 6.03e-19
C11542 VDD.n4616 VSS 0.0013f
C11543 VDD.n4617 VSS 0.0027f
C11544 VDD.n4618 VSS 0.0028f
C11545 VDD.n4619 VSS 0.00106f
C11546 VDD.n4620 VSS 0.00151f
C11547 VDD.n4621 VSS 0.0018f
C11548 VDD.n4622 VSS 0.00231f
C11549 VDD.t649 VSS 0.00579f
C11550 VDD.n4623 VSS 0.00598f
C11551 VDD.n4624 VSS 0.00109f
C11552 VDD.t630 VSS 8.49e-19
C11553 VDD.t650 VSS -2.71e-19
C11554 VDD.n4625 VSS 0.00391f
C11555 VDD.n4626 VSS 0.00413f
C11556 VDD.n4627 VSS 9.92e-19
C11557 VDD.n4628 VSS 0.00308f
C11558 VDD.t629 VSS 0.00579f
C11559 VDD.n4629 VSS 0.00838f
C11560 VDD.n4630 VSS 0.00109f
C11561 VDD.n4631 VSS 0.00186f
C11562 VDD.n4632 VSS 0.00308f
C11563 VDD.n4633 VSS 0.00926f
C11564 VDD.n4634 VSS 0.00109f
C11565 VDD.n4635 VSS 0.00164f
C11566 VDD.n4636 VSS 0.0028f
C11567 VDD.n4637 VSS 0.00154f
C11568 VDD.n4638 VSS 0.00203f
C11569 VDD.t507 VSS 9.16e-19
C11570 VDD.t632 VSS -5.07e-19
C11571 VDD.n4639 VSS 0.00359f
C11572 VDD.n4640 VSS 6.69e-19
C11573 VDD.n4641 VSS 1.17e-19
C11574 VDD.n4642 VSS 5.4e-19
C11575 VDD.n4643 VSS 1.01e-19
C11576 VDD.n4644 VSS 0.00372f
C11577 VDD.n4645 VSS 0.00107f
C11578 VDD.t631 VSS 0.00579f
C11579 VDD.n4646 VSS 0.00239f
C11580 VDD.n4647 VSS 5.52e-19
C11581 VDD.n4648 VSS 0.0015f
C11582 VDD.n4649 VSS 4.21e-19
C11583 VDD.n4650 VSS 0.00183f
C11584 VDD.t506 VSS 0.00472f
C11585 VDD.n4651 VSS 0.00781f
C11586 VDD.n4652 VSS 9.91e-19
C11587 VDD.n4653 VSS 0.0039f
C11588 VDD.n4654 VSS 0.00308f
C11589 VDD.t402 VSS 0.00262f
C11590 VDD.n4655 VSS 0.00271f
C11591 VDD.n4656 VSS 0.00989f
C11592 VDD.n4657 VSS 0.00109f
C11593 VDD.n4658 VSS 0.00269f
C11594 VDD.n4659 VSS 0.00308f
C11595 VDD.t689 VSS 0.00579f
C11596 VDD.t401 VSS 0.00579f
C11597 VDD.n4660 VSS 0.00453f
C11598 VDD.n4661 VSS 0.00109f
C11599 VDD.n4662 VSS 0.00172f
C11600 VDD.n4663 VSS 0.00308f
C11601 VDD.n4664 VSS 0.00668f
C11602 VDD.n4665 VSS 0.00109f
C11603 VDD.n4666 VSS 0.00164f
C11604 VDD.n4667 VSS 0.00308f
C11605 VDD.t634 VSS 7.62e-19
C11606 VDD.t92 VSS 5.72e-19
C11607 VDD.n4668 VSS 0.0014f
C11608 VDD.t91 VSS 0.00579f
C11609 VDD.n4669 VSS 0.00762f
C11610 VDD.n4670 VSS 0.00111f
C11611 VDD.n4671 VSS 0.00204f
C11612 VDD.n4672 VSS 0.00252f
C11613 VDD.n4673 VSS 0.00308f
C11614 VDD.t633 VSS 0.00579f
C11615 VDD.n4674 VSS 0.00605f
C11616 VDD.n4675 VSS 0.00109f
C11617 VDD.n4676 VSS 0.00132f
C11618 VDD.n4677 VSS 0.00308f
C11619 VDD.t595 VSS 0.00579f
C11620 VDD.n4678 VSS 0.00636f
C11621 VDD.n4679 VSS 0.00109f
C11622 VDD.n4680 VSS 0.00186f
C11623 VDD.n4681 VSS 0.00308f
C11624 VDD.t166 VSS 0.00579f
C11625 VDD.n4682 VSS 0.00529f
C11626 VDD.n4683 VSS 0.00109f
C11627 VDD.n4684 VSS 0.00186f
C11628 VDD.n4685 VSS 0.00308f
C11629 VDD.n4686 VSS 0.00907f
C11630 VDD.n4687 VSS 0.00109f
C11631 VDD.n4688 VSS 0.00182f
C11632 VDD.n4689 VSS 0.00302f
C11633 VDD.n4690 VSS 0.00154f
C11634 VDD.t300 VSS 0.00579f
C11635 VDD.n4691 VSS 0.00825f
C11636 VDD.n4692 VSS 0.00109f
C11637 VDD.n4693 VSS 9.31e-19
C11638 VDD.n4694 VSS 1.72e-19
C11639 VDD.n4695 VSS 2.85e-19
C11640 VDD.n4696 VSS 1.72e-19
C11641 VDD.n4697 VSS 5.86e-19
C11642 VDD.n4698 VSS 4.35e-19
C11643 VDD.n4699 VSS 3.36e-19
C11644 VDD.n4700 VSS 8.1e-19
C11645 VDD.n4701 VSS 0.0217f
C11646 VDD.n4702 VSS 0.0113f
C11647 VDD.n4703 VSS 0.00788f
C11648 VDD.n4704 VSS 0.0103f
C11649 VDD.n4705 VSS 0.0113f
C11650 VDD.n4706 VSS 0.0148f
C11651 VDD.n4707 VSS 8.1e-19
C11652 VDD.n4708 VSS 0.00157f
C11653 VDD.n4709 VSS 0.00144f
C11654 VDD.n4710 VSS 0.0109f
C11655 VDD.n4711 VSS 0.0117f
C11656 VDD.n4712 VSS 0.00109f
C11657 VDD.n4713 VSS 0.00157f
C11658 VDD.n4714 VSS 0.0117f
C11659 VDD.n4715 VSS 0.00109f
C11660 VDD.n4716 VSS 0.00157f
C11661 VDD.n4717 VSS 0.0117f
C11662 VDD.n4718 VSS 0.00109f
C11663 VDD.n4719 VSS 0.00157f
C11664 VDD.n4720 VSS 0.0117f
C11665 VDD.n4721 VSS 0.00109f
C11666 VDD.n4722 VSS 0.00129f
C11667 VDD.n4723 VSS 0.00927f
C11668 VDD.n4724 VSS 0.00109f
C11669 VDD.n4725 VSS 9.31e-19
C11670 VDD.n4726 VSS 9.39e-19
C11671 VDD.n4727 VSS 0.0123f
C11672 VDD.t670 VSS 4.25e-19
C11673 VDD.t247 VSS 5.42e-19
C11674 VDD.n4728 VSS 0.00111f
C11675 VDD.n4729 VSS 0.00218f
C11676 VDD.t669 VSS 0.00584f
C11677 VDD.n4730 VSS 0.0061f
C11678 VDD.n4731 VSS 0.00109f
C11679 VDD.n4732 VSS 4.66e-19
C11680 VDD.n4733 VSS 9.31e-19
C11681 VDD.n4734 VSS 0.00308f
C11682 VDD.t246 VSS 0.00584f
C11683 VDD.t603 VSS 0.00584f
C11684 VDD.n4735 VSS 0.00457f
C11685 VDD.n4736 VSS 0.00109f
C11686 VDD.n4737 VSS 9.31e-19
C11687 VDD.n4738 VSS 8.7e-19
C11688 VDD.n4739 VSS 0.00308f
C11689 VDD.n4740 VSS 0.00927f
C11690 VDD.n4741 VSS 0.00109f
C11691 VDD.n4742 VSS 9.31e-19
C11692 VDD.n4743 VSS 9.31e-19
C11693 VDD.n4744 VSS 0.00308f
C11694 VDD.n4745 VSS 0.0102f
C11695 VDD.n4746 VSS 0.00109f
C11696 VDD.n4747 VSS 9.31e-19
C11697 VDD.n4748 VSS 9.31e-19
C11698 VDD.n4749 VSS 0.00308f
C11699 VDD.t560 VSS 0.00584f
C11700 VDD.n4750 VSS 0.00654f
C11701 VDD.n4751 VSS 0.00109f
C11702 VDD.n4752 VSS 9.31e-19
C11703 VDD.n4753 VSS 9.31e-19
C11704 VDD.n4754 VSS 0.00308f
C11705 VDD.t575 VSS 0.00584f
C11706 VDD.n4755 VSS 0.00667f
C11707 VDD.n4756 VSS 0.00109f
C11708 VDD.n4757 VSS 9.31e-19
C11709 VDD.n4758 VSS 9.31e-19
C11710 VDD.n4759 VSS 0.00308f
C11711 VDD.n4760 VSS 0.00308f
C11712 VDD.n4761 VSS 0.0117f
C11713 VDD.n4762 VSS 0.00109f
C11714 VDD.n4763 VSS 0.00157f
C11715 VDD.t576 VSS 7.73e-19
C11716 VDD.t55 VSS 2.51e-19
C11717 VDD.n4764 VSS 0.00395f
C11718 VDD.n4765 VSS 5.46e-19
C11719 VDD.n4766 VSS 0.00255f
C11720 VDD.n4767 VSS 9.11e-19
C11721 VDD.n4768 VSS 0.00109f
C11722 VDD.n4769 VSS 0.0061f
C11723 VDD.t54 VSS 0.00152f
C11724 VDD.n4770 VSS 0.0102f
C11725 VDD.n4771 VSS 0.00109f
C11726 VDD.n4772 VSS 0.00122f
C11727 VDD.n4773 VSS 9.31e-19
C11728 VDD.n4774 VSS 0.00181f
C11729 VDD.n4775 VSS 0.00328f
C11730 VDD.n4776 VSS 0.00184f
C11731 VDD.n4777 VSS 0.00109f
C11732 VDD.n4778 VSS 0.00889f
C11733 VDD.t335 VSS 0.00394f
C11734 VDD.n4779 VSS 0.00603f
C11735 VDD.n4780 VSS 0.00109f
C11736 VDD.n4781 VSS 9.51e-19
C11737 VDD.n4782 VSS 0.00278f
C11738 VDD.t297 VSS 0.00584f
C11739 VDD.n4783 VSS 0.00654f
C11740 VDD.n4784 VSS 0.00109f
C11741 VDD.n4785 VSS 0.00186f
C11742 VDD.n4786 VSS 0.00308f
C11743 VDD.t565 VSS 0.00584f
C11744 VDD.n4787 VSS 0.00686f
C11745 VDD.n4788 VSS 0.00109f
C11746 VDD.n4789 VSS 0.00178f
C11747 VDD.n4790 VSS 0.00251f
C11748 VDD.n4791 VSS 0.00112f
C11749 VDD.t384 VSS 0.00495f
C11750 VDD.n4792 VSS 0.0061f
C11751 VDD.n4793 VSS 0.00109f
C11752 VDD.n4794 VSS 0.0014f
C11753 VDD.n4795 VSS 0.00308f
C11754 VDD.t179 VSS 0.00546f
C11755 VDD.n4796 VSS 0.00673f
C11756 VDD.n4797 VSS 0.00109f
C11757 VDD.n4798 VSS 0.00177f
C11758 VDD.n4799 VSS 0.00293f
C11759 VDD.n4800 VSS 0.00154f
C11760 VDD.n4801 VSS 9.31e-19
C11761 VDD.n4802 VSS 0.0117f
C11762 VDD.n4803 VSS 0.00109f
C11763 VDD.n4804 VSS 1.72e-19
C11764 VDD.n4805 VSS 2.85e-19
C11765 VDD.n4806 VSS 9.31e-19
C11766 VDD.n4807 VSS 4.19e-19
C11767 VDD.n4808 VSS 4.35e-19
C11768 VDD.n4809 VSS 5.07e-19
C11769 VDD.n4810 VSS 3.36e-19
C11770 VDD.n4811 VSS 8.1e-19
C11771 VDD.n4812 VSS 0.00148f
C11772 VDD.n4813 VSS 0.00653f
C11773 VDD.n4814 VSS 0.00218f
C11774 VDD.t385 VSS 5.42e-19
C11775 VDD.t57 VSS 4.25e-19
C11776 VDD.n4815 VSS 0.00111f
C11777 VDD.n4816 VSS 0.00259f
C11778 VDD.t56 VSS 0.00584f
C11779 VDD.n4817 VSS 0.00597f
C11780 VDD.n4818 VSS 0.00109f
C11781 VDD.n4819 VSS 0.00134f
C11782 VDD.n4820 VSS 0.00298f
C11783 VDD.n4821 VSS 0.00154f
C11784 VDD.n4822 VSS 9.31e-19
C11785 VDD.n4823 VSS 0.0442f
C11786 VDD.n4824 VSS 0.00377f
C11787 VDD.n4825 VSS 1.72e-19
C11788 VDD.n4826 VSS 2.85e-19
C11789 VDD.n4827 VSS 0.00533f
C11790 VDD.n4828 VSS 5.03e-19
C11791 VDD.n4829 VSS 4.82e-19
C11792 VDD.n4830 VSS 0.00149f
C11793 VDD.n4831 VSS 8.1e-19
C11794 VDD.n4832 VSS 6.3e-19
C11795 VDD.n4833 VSS 3.36e-19
C11796 VDD.n4834 VSS 4.35e-19
C11797 VDD.n4835 VSS 2.68e-19
C11798 VDD.n4836 VSS 0.00995f
C11799 VDD.n4837 VSS 0.00144f
C11800 VDD.n4838 VSS 0.00148f
C11801 VDD.n4839 VSS 8.1e-19
C11802 VDD.n4840 VSS 0.00157f
C11803 VDD.n4841 VSS 0.00581f
C11804 VDD.n4842 VSS 0.00653f
C11805 VDD.n4843 VSS 0.00218f
C11806 VDD.n4844 VSS 0.252f
C11807 VDD.n4845 VSS 0.263f
C11808 VDD.n4846 VSS 0.00441f
C11809 VDD.n4847 VSS 0.00158f
C11810 VDD.n4848 VSS 4.39e-19
C11811 VDD.n4849 VSS 0.00154f
C11812 VDD.n4850 VSS 9.31e-19
C11813 VDD.t519 VSS 0.00578f
C11814 VDD.n4851 VSS 0.00528f
C11815 VDD.n4852 VSS 0.00109f
C11816 VDD.n4853 VSS 1.72e-19
C11817 VDD.n4854 VSS 2.85e-19
C11818 VDD.n4855 VSS 6.27e-19
C11819 VDD.n4856 VSS 5.86e-19
C11820 VDD.t520 VSS 9.42e-19
C11821 VDD.t546 VSS 9.42e-19
C11822 VDD.n4857 VSS 0.00214f
C11823 VDD.n4858 VSS 0.00244f
C11824 VDD.t545 VSS 0.00578f
C11825 VDD.n4859 VSS 0.00528f
C11826 VDD.n4860 VSS 0.00109f
C11827 VDD.n4861 VSS 0.00123f
C11828 VDD.n4862 VSS 0.00243f
C11829 VDD.n4863 VSS 9.55e-19
C11830 VDD.n4864 VSS 4.35e-19
C11831 VDD.n4865 VSS 6.68e-19
C11832 VDD.n4866 VSS 3.36e-19
C11833 VDD.n4867 VSS 0.00149f
C11834 VDD.n4868 VSS 8.1e-19
C11835 VDD.n4869 VSS 0.00335f
C11836 VDD.n4870 VSS 0.0136f
C11837 VDD.n4871 VSS 0.0136f
C11838 VDD.n4872 VSS 0.00335f
C11839 VDD.n4873 VSS 0.00179f
C11840 VDD.n4874 VSS 0.67f
.ends

