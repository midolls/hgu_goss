* NGSPICE file created from hgu_comp_flat.ext - technology: sky130A

.subckt hgu_comp ready cdac_vn comp_outp comp_outn cdac_vp clk VDD VSS
X0 Q cdac_vn.t0 a_582_n702# VSS.t65 sky130_fd_pr__nfet_01v8_lvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1 ready.t1 a_564_n1721# VDD.t2 VDD.t1 sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0.244 ps=2.26 w=0.84 l=0.15
X2 a_564_n1721# a_476_n1721# a_564_n1266# VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.15
X3 comp_outn.t5 a_1950_n1721# VDD.t14 VDD.t13 sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.3 as=0.139 ps=1.17 w=0.84 l=0.15
X4 a_582_n702# cdac_vn.t1 Q VSS.t64 sky130_fd_pr__nfet_01v8_lvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X5 a_1950_n1721# RS_n VDD.t8 VDD.t7 sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0.244 ps=2.26 w=0.84 l=0.15
X6 a_482_n1818# a_1716_n1348# VSS.t43 VSS.t42 sky130_fd_pr__nfet_01v8 ad=0.0759 pd=0.79 as=0.143 ps=1.54 w=0.46 l=0.15
X7 a_564_n1721# a_482_n1818# a_476_n1721# VDD.t49 sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.15
X8 VDD.t32 a_1026_n1747# comp_outp.t5 VDD.t31 sky130_fd_pr__pfet_01v8 ad=0.139 pd=1.17 as=0.26 ps=2.3 w=0.84 l=0.15
X9 VSS.t53 RS_p a_1026_n1747# VSS.t52 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X10 VDD.t22 clk.t0 a_1248_n288# VDD.t21 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X11 a_674_n702# cdac_vp.t0 a_582_n702# VSS.t26 sky130_fd_pr__nfet_01v8_lvt ad=0.165 pd=1.33 as=0.31 ps=2.62 w=1 l=0.15
X12 VDD.t20 a_852_n296# a_476_n1721# VDD.t19 sky130_fd_pr__pfet_01v8 ad=0.139 pd=1.17 as=0.26 ps=2.3 w=0.84 l=0.15
X13 comp_outp.t4 a_1026_n1747# VDD.t30 VDD.t29 sky130_fd_pr__pfet_01v8 ad=0.139 pd=1.17 as=0.139 ps=1.17 w=0.84 l=0.15
X14 a_476_n1721# a_852_n296# VDD.t18 VDD.t17 sky130_fd_pr__pfet_01v8 ad=0.139 pd=1.17 as=0.139 ps=1.17 w=0.84 l=0.15
X15 a_582_n702# cdac_vn.t2 Q VSS.t63 sky130_fd_pr__nfet_01v8_lvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X16 a_582_n702# cdac_vp.t1 a_674_n702# VSS.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X17 comp_outn.t2 a_1950_n1721# VSS.t15 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.54 as=0.0759 ps=0.79 w=0.46 l=0.15
X18 VDD.t48 RS_p a_1026_n1747# VDD.t47 sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0.244 ps=2.26 w=0.84 l=0.15
X19 VDD.t16 a_852_n296# a_476_n1721# VDD.t15 sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.3 as=0.139 ps=1.17 w=0.84 l=0.15
X20 a_674_n702# cdac_vp.t2 a_582_n702# VSS.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X21 Q cdac_vn.t3 a_582_n702# VSS.t62 sky130_fd_pr__nfet_01v8_lvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X22 a_564_n1266# a_482_n1818# VSS.t55 VSS.t54 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.15
X23 VSS.t36 a_1026_n1747# comp_outp.t2 VSS.t35 sky130_fd_pr__nfet_01v8 ad=0.0759 pd=0.79 as=0.143 ps=1.54 w=0.46 l=0.15
X24 a_1950_n1721# RS_n VSS.t9 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X25 a_1566_n378# clk.t1 VDD.t40 VDD.t39 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X26 VSS.t25 a_852_n296# a_476_n1721# VSS.t24 sky130_fd_pr__nfet_01v8 ad=0.0759 pd=0.79 as=0.143 ps=1.54 w=0.46 l=0.15
X27 VDD.t26 a_1248_n288# a_852_n296# VDD.t25 sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0.244 ps=2.26 w=0.84 l=0.15
X28 a_482_n1818# a_1716_n1348# VSS.t41 VSS.t40 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.54 as=0.0759 ps=0.79 w=0.46 l=0.15
X29 a_582_n702# clk.t2 VSS.t17 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X30 comp_outp.t1 a_1026_n1747# VSS.t34 VSS.t33 sky130_fd_pr__nfet_01v8 ad=0.0759 pd=0.79 as=0.0759 ps=0.79 w=0.46 l=0.15
X31 VSS.t30 a_1248_n288# a_852_n296# VSS.t29 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X32 a_674_n702# cdac_vp.t3 a_582_n702# VSS.t47 sky130_fd_pr__nfet_01v8_lvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X33 a_582_n702# cdac_vn.t4 Q VSS.t61 sky130_fd_pr__nfet_01v8_lvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X34 a_1248_n288# a_1566_n378# VDD.t44 VDD.t43 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X35 Q clk.t3 VDD.t51 VDD.t50 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X36 a_582_n702# cdac_vp.t4 a_674_n702# VSS.t27 sky130_fd_pr__nfet_01v8_lvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X37 VDD.t28 a_1026_n1747# comp_outp.t3 VDD.t27 sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.3 as=0.139 ps=1.17 w=0.84 l=0.15
X38 RS_n a_1716_n1348# VSS.t39 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.15
X39 comp_outn.t4 a_1950_n1721# VDD.t12 VDD.t11 sky130_fd_pr__pfet_01v8 ad=0.139 pd=1.17 as=0.26 ps=2.3 w=0.84 l=0.15
X40 a_1716_n1348# a_1566_n378# VSS.t51 VSS.t50 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X41 VSS.t38 a_1716_n1348# a_482_n1818# VSS.t37 sky130_fd_pr__nfet_01v8 ad=0.0759 pd=0.79 as=0.0759 ps=0.79 w=0.46 l=0.15
X42 VSS.t57 clk.t4 a_582_n702# VSS.t56 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.31 ps=2.62 w=1 l=0.15
X43 a_582_n702# cdac_vn.t5 Q VSS.t60 sky130_fd_pr__nfet_01v8_lvt ad=0.31 pd=2.62 as=0.165 ps=1.33 w=1 l=0.15
X44 VSS.t23 a_852_n296# a_476_n1721# VSS.t22 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.54 as=0.0759 ps=0.79 w=0.46 l=0.15
X45 Q a_1566_n378# a_1248_n288# VSS.t49 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X46 Q cdac_vn.t6 a_582_n702# VSS.t59 sky130_fd_pr__nfet_01v8_lvt ad=0.165 pd=1.33 as=0.31 ps=2.62 w=1 l=0.15
X47 RS_n RS_p VDD.t46 VDD.t45 sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.15
X48 VDD.t10 a_1950_n1721# comp_outn.t3 VDD.t9 sky130_fd_pr__pfet_01v8 ad=0.139 pd=1.17 as=0.139 ps=1.17 w=0.84 l=0.15
X49 a_1716_n1348# a_1566_n378# VDD.t42 VDD.t41 sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0.244 ps=2.26 w=0.84 l=0.15
X50 a_582_n702# clk.t5 VSS.t46 VSS.t45 sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.165 ps=1.33 w=1 l=0.15
X51 VDD.t4 clk.t6 a_674_n702# VDD.t3 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X52 a_674_n702# cdac_vp.t5 a_582_n702# VSS.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X53 VSS.t32 a_1026_n1747# comp_outp.t0 VSS.t31 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.54 as=0.0759 ps=0.79 w=0.46 l=0.15
X54 comp_outn.t1 a_1950_n1721# VSS.t13 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0.0759 pd=0.79 as=0.143 ps=1.54 w=0.46 l=0.15
X55 a_482_n1818# a_1716_n1348# VDD.t38 VDD.t37 sky130_fd_pr__pfet_01v8 ad=0.139 pd=1.17 as=0.26 ps=2.3 w=0.84 l=0.15
X56 a_482_n1818# a_1716_n1348# VDD.t36 VDD.t35 sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.3 as=0.139 ps=1.17 w=0.84 l=0.15
X57 a_582_n702# cdac_vp.t6 a_674_n702# VSS.t48 sky130_fd_pr__nfet_01v8_lvt ad=0.31 pd=2.62 as=0.165 ps=1.33 w=1 l=0.15
X58 VSS.t21 a_852_n296# RS_p VSS.t20 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.15
X59 VDD.t34 a_1716_n1348# a_482_n1818# VDD.t33 sky130_fd_pr__pfet_01v8 ad=0.139 pd=1.17 as=0.139 ps=1.17 w=0.84 l=0.15
X60 Q cdac_vn.t7 a_582_n702# VSS.t58 sky130_fd_pr__nfet_01v8_lvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X61 ready.t0 a_564_n1721# VSS.t3 VSS.t2 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X62 a_482_n1818# a_476_n1721# a_564_n1721# VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.15
X63 VSS.t11 a_1950_n1721# comp_outn.t0 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0.0759 pd=0.79 as=0.0759 ps=0.79 w=0.46 l=0.15
X64 a_476_n1721# a_852_n296# VSS.t19 VSS.t18 sky130_fd_pr__nfet_01v8 ad=0.0759 pd=0.79 as=0.0759 ps=0.79 w=0.46 l=0.15
X65 VDD.t24 a_1248_n288# a_1566_n378# VDD.t23 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X66 a_1566_n378# a_1248_n288# a_674_n702# VSS.t28 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X67 a_582_n702# cdac_vp.t7 a_674_n702# VSS.t44 sky130_fd_pr__nfet_01v8_lvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X68 VSS.t6 clk.t7 a_582_n702# VSS.t5 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X69 VDD.t6 RS_n RS_p VDD.t5 sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.15
R0 cdac_vn.n0 cdac_vn.t6 340.613
R1 cdac_vn.n6 cdac_vn.t5 186.374
R2 cdac_vn.n0 cdac_vn.t2 186.374
R3 cdac_vn.n1 cdac_vn.t0 186.374
R4 cdac_vn.n2 cdac_vn.t4 186.374
R5 cdac_vn.n3 cdac_vn.t3 186.374
R6 cdac_vn.n4 cdac_vn.t1 186.374
R7 cdac_vn.n5 cdac_vn.t7 186.374
R8 cdac_vn.n6 cdac_vn.n5 154.24
R9 cdac_vn.n5 cdac_vn.n4 154.24
R10 cdac_vn.n4 cdac_vn.n3 154.24
R11 cdac_vn.n3 cdac_vn.n2 154.24
R12 cdac_vn.n2 cdac_vn.n1 154.24
R13 cdac_vn.n1 cdac_vn.n0 154.24
R14 cdac_vn cdac_vn.n6 106.293
R15 VSS.n108 VSS.t59 179.739
R16 VSS.n102 VSS.t8 179.739
R17 VSS.n118 VSS.t10 175.16
R18 VSS.n78 VSS.t52 172.549
R19 VSS.n65 VSS.t31 172.549
R20 VSS.n69 VSS.t48 165.359
R21 VSS.n65 VSS.t27 165.359
R22 VSS.n91 VSS.t5 165.359
R23 VSS.n113 VSS.t12 161.147
R24 VSS.n91 VSS.t20 150.981
R25 VSS.n112 VSS.t65 140.127
R26 VSS.n31 VSS.t54 129.412
R27 VSS.n85 VSS.t28 122.222
R28 VSS.n97 VSS.t49 107.844
R29 VSS.n39 VSS.t44 107.844
R30 VSS.t29 VSS.t7 100.654
R31 VSS.n61 VSS.t22 93.4646
R32 VSS.n35 VSS.t26 93.4646
R33 VSS.n160 VSS.t58 91.0833
R34 VSS.n143 VSS.t51 86.7771
R35 VSS.n9 VSS.t30 85.4529
R36 VSS.n30 VSS.t55 83.725
R37 VSS.n13 VSS.t23 80.7031
R38 VSS.n139 VSS.t43 80.7031
R39 VSS.n71 VSS.t32 80.7031
R40 VSS.n106 VSS.t13 80.7031
R41 VSS.n43 VSS.t3 80.5977
R42 VSS.n80 VSS.t53 80.5977
R43 VSS.n3 VSS.t9 80.5977
R44 VSS.n69 VSS.t29 79.0855
R45 VSS.n55 VSS.t18 79.0855
R46 VSS.t26 VSS.t0 79.0855
R47 VSS.t50 VSS.t63 79.0708
R48 VSS.n164 VSS.t60 77.0706
R49 VSS.n96 VSS.n95 71.5328
R50 VSS.n84 VSS.n83 71.5328
R51 VSS.n117 VSS.t42 70.0642
R52 VSS.n50 VSS.t24 64.7064
R53 VSS.n107 VSS.t50 57.5168
R54 VSS.t22 VSS.t1 57.5168
R55 VSS.t18 VSS.t4 57.5168
R56 VSS.t24 VSS.t47 57.5168
R57 VSS.t40 VSS.t64 56.0515
R58 VSS.t37 VSS.t62 56.0515
R59 VSS.n124 VSS.t37 56.0515
R60 VSS.t42 VSS.t61 56.0515
R61 VSS.n90 VSS.n89 51.9572
R62 VSS.t47 VSS.t2 50.3273
R63 VSS.t49 VSS.t45 43.1378
R64 VSS.t28 VSS.t56 43.1378
R65 VSS.n21 VSS.t19 43.044
R66 VSS.n21 VSS.t25 43.044
R67 VSS.n135 VSS.t41 43.044
R68 VSS.n135 VSS.t38 43.044
R69 VSS.n59 VSS.t34 43.044
R70 VSS.n59 VSS.t36 43.044
R71 VSS.n120 VSS.t15 43.044
R72 VSS.n120 VSS.t11 43.044
R73 VSS.n130 VSS.t40 42.0387
R74 VSS.n22 VSS.n21 37.6596
R75 VSS.n136 VSS.n135 37.6596
R76 VSS.n60 VSS.n59 37.6596
R77 VSS.n121 VSS.n120 37.6596
R78 VSS.t20 VSS.t16 28.7587
R79 VSS.n45 VSS.n44 28.7587
R80 VSS.t61 VSS.t14 28.026
R81 VSS.n89 VSS.t39 20.7148
R82 VSS.n89 VSS.t21 20.7148
R83 VSS.n95 VSS.t46 19.8005
R84 VSS.n95 VSS.t6 19.8005
R85 VSS.n83 VSS.t17 19.8005
R86 VSS.n83 VSS.t57 19.8005
R87 VSS.n141 VSS.n140 9.15497
R88 VSS.n145 VSS.n144 9.15497
R89 VSS.n138 VSS.n137 9.15497
R90 VSS.n149 VSS.n148 9.15497
R91 VSS.n24 VSS.n23 9.15497
R92 VSS.n11 VSS.n10 9.15497
R93 VSS.n15 VSS.n14 9.15497
R94 VSS.n18 VSS.n17 9.15497
R95 VSS.n143 VSS.n142 9.15497
R96 VSS.n9 VSS.n8 9.15497
R97 VSS.n30 VSS.n29 9.15497
R98 VSS.n47 VSS.n46 9.15497
R99 VSS.n46 VSS.n45 9.15497
R100 VSS.n41 VSS.n40 9.15497
R101 VSS.n40 VSS.n39 9.15497
R102 VSS.n138 VSS.n136 7.94533
R103 VSS.n108 VSS.n107 7.19004
R104 VSS.t27 VSS.t33 7.19004
R105 VSS.t1 VSS.t35 7.19004
R106 VSS.n131 VSS.n130 7.00687
R107 VSS.n125 VSS.n124 7.00687
R108 VSS.n118 VSS.n117 7.00687
R109 VSS.n113 VSS.n112 7.00687
R110 VSS.n24 VSS.n22 6.62119
R111 VSS.n141 VSS.n139 6.17981
R112 VSS.n15 VSS.n13 4.85567
R113 VSS.n147 VSS.n141 4.6505
R114 VSS.n150 VSS.n149 4.6505
R115 VSS.n19 VSS.n18 4.6505
R116 VSS.n16 VSS.n15 4.6505
R117 VSS.n48 VSS.n47 4.6505
R118 VSS.n42 VSS.n41 4.6505
R119 VSS.n6 VSS.n5 4.57773
R120 VSS.n5 VSS.n4 4.57773
R121 VSS.n33 VSS.n32 4.57773
R122 VSS.n32 VSS.n31 4.57773
R123 VSS.n37 VSS.n36 4.57773
R124 VSS.n36 VSS.n35 4.57773
R125 VSS.n81 VSS.n79 4.57773
R126 VSS.n79 VSS.n78 4.57773
R127 VSS.n76 VSS.n75 4.57773
R128 VSS.n75 VSS.n74 4.57773
R129 VSS.n72 VSS.n70 4.57773
R130 VSS.n70 VSS.n69 4.57773
R131 VSS.n67 VSS.n66 4.57773
R132 VSS.n66 VSS.n65 4.57773
R133 VSS.n63 VSS.n62 4.57773
R134 VSS.n62 VSS.n61 4.57773
R135 VSS.n57 VSS.n56 4.57773
R136 VSS.n56 VSS.n55 4.57773
R137 VSS.n52 VSS.n51 4.57773
R138 VSS.n51 VSS.n50 4.57773
R139 VSS.n99 VSS.n98 4.57773
R140 VSS.n98 VSS.n97 4.57773
R141 VSS.n93 VSS.n92 4.57773
R142 VSS.n92 VSS.n91 4.57773
R143 VSS.n87 VSS.n86 4.57773
R144 VSS.n86 VSS.n85 4.57773
R145 VSS.n2 VSS.n1 4.57773
R146 VSS.n1 VSS.n0 4.57773
R147 VSS.n166 VSS.n165 4.57773
R148 VSS.n165 VSS.n164 4.57773
R149 VSS.n162 VSS.n161 4.57773
R150 VSS.n161 VSS.n160 4.57773
R151 VSS.n133 VSS.n132 4.57773
R152 VSS.n132 VSS.n131 4.57773
R153 VSS.n127 VSS.n126 4.57773
R154 VSS.n126 VSS.n125 4.57773
R155 VSS.n122 VSS.n119 4.57773
R156 VSS.n119 VSS.n118 4.57773
R157 VSS.n115 VSS.n114 4.57773
R158 VSS.n114 VSS.n113 4.57773
R159 VSS.n110 VSS.n109 4.57773
R160 VSS.n109 VSS.n108 4.57773
R161 VSS.n104 VSS.n103 4.57773
R162 VSS.n103 VSS.n102 4.57773
R163 VSS.n12 VSS.n9 3.40067
R164 VSS.n146 VSS.n143 3.40067
R165 VSS.n12 VSS.n11 3.25009
R166 VSS.n146 VSS.n145 3.25009
R167 VSS.n153 VSS.n138 3.03426
R168 VSS.n25 VSS.n24 3.03311
R169 VSS.n168 VSS.n2 2.34608
R170 VSS.n38 VSS.n37 2.3255
R171 VSS.n82 VSS.n81 2.3255
R172 VSS.n77 VSS.n76 2.3255
R173 VSS.n73 VSS.n72 2.3255
R174 VSS.n68 VSS.n67 2.3255
R175 VSS.n64 VSS.n63 2.3255
R176 VSS.n58 VSS.n57 2.3255
R177 VSS.n100 VSS.n99 2.3255
R178 VSS.n94 VSS.n93 2.3255
R179 VSS.n88 VSS.n87 2.3255
R180 VSS.n101 VSS.n6 2.3255
R181 VSS.n167 VSS.n166 2.3255
R182 VSS.n163 VSS.n162 2.3255
R183 VSS.n128 VSS.n127 2.3255
R184 VSS.n123 VSS.n122 2.3255
R185 VSS.n116 VSS.n115 2.3255
R186 VSS.n111 VSS.n110 2.3255
R187 VSS.n105 VSS.n104 2.3255
R188 VSS.n158 VSS.n157 2.2505
R189 VSS.n27 VSS.n26 2.24128
R190 VSS.n28 VSS.n27 1.84746
R191 VSS.n156 VSS.n155 1.84746
R192 VSS.n53 VSS.n52 1.83603
R193 VSS.n134 VSS.n133 1.83603
R194 VSS.n154 VSS.n153 1.50988
R195 VSS.n38 VSS.n34 1.24353
R196 VSS.n54 VSS.n28 1.16147
R197 VSS.n34 VSS.n30 1.11176
R198 VSS.n16 VSS.n12 0.932839
R199 VSS.n147 VSS.n146 0.932839
R200 VSS.n34 VSS.n33 0.548326
R201 VSS.n99 VSS.n96 0.312695
R202 VSS.n47 VSS.n43 0.234646
R203 VSS.n110 VSS.n106 0.234646
R204 VSS.n6 VSS.n3 0.234646
R205 VSS VSS.n168 0.231462
R206 VSS.n19 VSS.n16 0.216017
R207 VSS.n150 VSS.n147 0.216017
R208 VSS.n20 VSS.n19 0.187208
R209 VSS.n151 VSS.n150 0.166381
R210 VSS.n81 VSS.n80 0.156598
R211 VSS.n72 VSS.n71 0.156598
R212 VSS.n63 VSS.n60 0.156598
R213 VSS.n93 VSS.n90 0.104565
R214 VSS.n87 VSS.n84 0.104565
R215 VSS.n122 VSS.n121 0.0785488
R216 VSS.n100 VSS.n94 0.051313
R217 VSS.n94 VSS.n88 0.051313
R218 VSS.n42 VSS.n38 0.0493088
R219 VSS.n101 VSS.n100 0.0481372
R220 VSS.n88 VSS.n82 0.047375
R221 VSS.n152 VSS.n151 0.0415156
R222 VSS.n82 VSS.n77 0.0386098
R223 VSS.n77 VSS.n73 0.0386098
R224 VSS.n73 VSS.n68 0.0386098
R225 VSS.n68 VSS.n64 0.0386098
R226 VSS.n64 VSS.n58 0.0386098
R227 VSS.n167 VSS.n163 0.0386098
R228 VSS.n128 VSS.n123 0.0386098
R229 VSS.n123 VSS.n116 0.0386098
R230 VSS.n116 VSS.n111 0.0386098
R231 VSS.n111 VSS.n105 0.0386098
R232 VSS.n105 VSS.n101 0.0386098
R233 VSS.n58 VSS.n54 0.0382053
R234 VSS.n157 VSS.n156 0.0356562
R235 VSS.n129 VSS.n128 0.0351228
R236 VSS.n163 VSS.n159 0.0302256
R237 VSS.n49 VSS.n48 0.0298445
R238 VSS.n27 VSS.n7 0.0263062
R239 VSS.n155 VSS.n154 0.0263062
R240 VSS.n26 VSS.n20 0.0215034
R241 VSS.n168 VSS.n167 0.0180305
R242 VSS.n53 VSS.n49 0.00850305
R243 VSS.n159 VSS.n158 0.00850305
R244 VSS.n134 VSS.n129 0.00497985
R245 VSS.n54 VSS.n53 0.00389195
R246 VSS.n26 VSS.n25 0.00245312
R247 VSS.n153 VSS.n152 0.0023033
R248 VSS.n48 VSS.n42 0.00126219
R249 VSS.n158 VSS.n134 0.000881098
R250 VDD.n241 VDD.t0 425.812
R251 VDD.t0 VDD.t49 183.923
R252 VDD.n243 VDD.t2 122.26
R253 VDD.n262 VDD.t48 113.861
R254 VDD.n173 VDD.t37 112.871
R255 VDD.n16 VDD.t15 112.871
R256 VDD.n330 VDD.t11 112.871
R257 VDD.n50 VDD.t26 112.731
R258 VDD.n137 VDD.t42 112.731
R259 VDD.n313 VDD.t8 112.356
R260 VDD.n234 VDD.t31 103.466
R261 VDD.n277 VDD.t5 97.2098
R262 VDD.n18 VDD.t16 91.0302
R263 VDD.n154 VDD.t38 91.0302
R264 VDD.n329 VDD.t12 91.0302
R265 VDD.n203 VDD.t28 91.0302
R266 VDD.n99 VDD.t21 89.3422
R267 VDD.n201 VDD.t27 84.654
R268 VDD.n33 VDD.t19 84.1029
R269 VDD.n361 VDD.t13 84.1029
R270 VDD.n85 VDD.t39 71.4739
R271 VDD.n187 VDD.t35 65.291
R272 VDD.n85 VDD.t23 59.5616
R273 VDD.n68 VDD.n67 58.3564
R274 VDD.n102 VDD.n101 58.3564
R275 VDD.n122 VDD.n121 58.3564
R276 VDD.n135 VDD.t41 53.6055
R277 VDD.n294 VDD.t45 53.5216
R278 VDD.n28 VDD.n27 52.3338
R279 VDD.n172 VDD.n171 52.3338
R280 VDD.n347 VDD.n346 52.3338
R281 VDD.n226 VDD.n225 52.3338
R282 VDD.n99 VDD.t43 41.6933
R283 VDD.n311 VDD.t7 39.1171
R284 VDD.n27 VDD.t18 38.6969
R285 VDD.n27 VDD.t20 38.6969
R286 VDD.n171 VDD.t36 38.6969
R287 VDD.n171 VDD.t34 38.6969
R288 VDD.n346 VDD.t14 38.6969
R289 VDD.n346 VDD.t10 38.6969
R290 VDD.n225 VDD.t30 38.6969
R291 VDD.n225 VDD.t32 38.6969
R292 VDD.n173 VDD.t33 37.6243
R293 VDD.n51 VDD.t25 35.7372
R294 VDD.n297 VDD.n296 35.0339
R295 VDD.n296 VDD.t46 34.0065
R296 VDD.n296 VDD.t6 34.0065
R297 VDD.n69 VDD.t3 29.7811
R298 VDD.n67 VDD.t40 28.5655
R299 VDD.n67 VDD.t4 28.5655
R300 VDD.n101 VDD.t44 28.5655
R301 VDD.n101 VDD.t24 28.5655
R302 VDD.n121 VDD.t51 28.5655
R303 VDD.n121 VDD.t22 28.5655
R304 VDD.n25 VDD.t17 18.8124
R305 VDD.n348 VDD.t9 18.8124
R306 VDD.n175 VDD.n172 14.4005
R307 VDD.n103 VDD.n102 14.4005
R308 VDD.n298 VDD.n297 13.6005
R309 VDD.n71 VDD.n68 12.8005
R310 VDD.n29 VDD.n28 12.0005
R311 VDD.n350 VDD.n347 12.0005
R312 VDD.n119 VDD.t50 11.9127
R313 VDD.n264 VDD.n263 10.6304
R314 VDD.n123 VDD.n122 10.4005
R315 VDD.n242 VDD.n241 9.92059
R316 VDD.n227 VDD.t29 9.40644
R317 VDD.n29 VDD.n26 8.85536
R318 VDD.n26 VDD.n25 8.85536
R319 VDD.n19 VDD.n17 8.85536
R320 VDD.n17 VDD.n16 8.85536
R321 VDD.n53 VDD.n52 8.85536
R322 VDD.n52 VDD.n51 8.85536
R323 VDD.n71 VDD.n70 8.85536
R324 VDD.n70 VDD.n69 8.85536
R325 VDD.n87 VDD.n86 8.85536
R326 VDD.n86 VDD.n85 8.85536
R327 VDD.n103 VDD.n100 8.85536
R328 VDD.n100 VDD.n99 8.85536
R329 VDD.n123 VDD.n120 8.85536
R330 VDD.n120 VDD.n119 8.85536
R331 VDD.n138 VDD.n136 8.85536
R332 VDD.n136 VDD.n135 8.85536
R333 VDD.n188 VDD.n187 8.85536
R334 VDD.n175 VDD.n174 8.85536
R335 VDD.n174 VDD.n173 8.85536
R336 VDD.n157 VDD.n156 8.85536
R337 VDD.n156 VDD.n155 8.85536
R338 VDD.n34 VDD.n33 8.85536
R339 VDD.n332 VDD.n331 8.85536
R340 VDD.n331 VDD.n330 8.85536
R341 VDD.n229 VDD.n228 8.85536
R342 VDD.n228 VDD.n227 8.85536
R343 VDD.n204 VDD.n202 8.85536
R344 VDD.n202 VDD.n201 8.85536
R345 VDD.n265 VDD.n264 8.85536
R346 VDD.n279 VDD.n278 8.85536
R347 VDD.n278 VDD.n277 8.85536
R348 VDD.n298 VDD.n295 8.85536
R349 VDD.n295 VDD.n294 8.85536
R350 VDD.n314 VDD.n312 8.85536
R351 VDD.n312 VDD.n311 8.85536
R352 VDD.n236 VDD.n235 8.85536
R353 VDD.n235 VDD.n234 8.85536
R354 VDD.n243 VDD.n242 8.85536
R355 VDD.n362 VDD.n361 8.85536
R356 VDD.n350 VDD.n349 8.85536
R357 VDD.n349 VDD.n348 8.85536
R358 VDD.n229 VDD.n226 8.4005
R359 VDD.n265 VDD.n262 7.6005
R360 VDD.n157 VDD.n154 7.2005
R361 VDD.n263 VDD.t47 5.50293
R362 VDD.n19 VDD.n18 4.8005
R363 VDD.n332 VDD.n329 4.8005
R364 VDD.n53 VDD.n50 4.0005
R365 VDD.n314 VDD.n313 4.0005
R366 VDD.n35 VDD.n34 3.03483
R367 VDD.n30 VDD.n29 3.03311
R368 VDD.n88 VDD.n87 3.03311
R369 VDD.n104 VDD.n103 3.03311
R370 VDD.n124 VDD.n123 3.03311
R371 VDD.n139 VDD.n138 3.03311
R372 VDD.n176 VDD.n175 3.03311
R373 VDD.n189 VDD.n188 3.03311
R374 VDD.n20 VDD.n19 3.03311
R375 VDD.n54 VDD.n53 3.03311
R376 VDD.n72 VDD.n71 3.03311
R377 VDD.n158 VDD.n157 3.03311
R378 VDD.n230 VDD.n229 3.03311
R379 VDD.n363 VDD.n362 3.03311
R380 VDD.n244 VDD.n243 3.03311
R381 VDD.n205 VDD.n204 3.03311
R382 VDD.n266 VDD.n265 3.03311
R383 VDD.n280 VDD.n279 3.03311
R384 VDD.n299 VDD.n298 3.03311
R385 VDD.n315 VDD.n314 3.03311
R386 VDD.n333 VDD.n332 3.03311
R387 VDD.n237 VDD.n236 3.03311
R388 VDD.n351 VDD.n350 3.03311
R389 VDD.n241 VDD.t1 1.83498
R390 VDD.n58 VDD.n57 1.7055
R391 VDD.n76 VDD.n75 1.7055
R392 VDD.n162 VDD.n161 1.7055
R393 VDD.n193 VDD.n192 1.7055
R394 VDD.n180 VDD.n179 1.7055
R395 VDD.n145 VDD.n144 1.7055
R396 VDD.n128 VDD.n127 1.7055
R397 VDD.n110 VDD.n109 1.7055
R398 VDD.n92 VDD.n91 1.7055
R399 VDD.n356 VDD.n355 1.7055
R400 VDD.n338 VDD.n337 1.7055
R401 VDD.n321 VDD.n320 1.7055
R402 VDD.n304 VDD.n303 1.7055
R403 VDD.n286 VDD.n285 1.7055
R404 VDD.n270 VDD.n269 1.7055
R405 VDD.n368 VDD.n367 1.7055
R406 VDD.n138 VDD.n137 1.6005
R407 VDD.n56 VDD.n55 1.35607
R408 VDD.n74 VDD.n73 1.35607
R409 VDD.n160 VDD.n159 1.35607
R410 VDD.n191 VDD.n190 1.35607
R411 VDD.n178 VDD.n177 1.35607
R412 VDD.n142 VDD.n141 1.35607
R413 VDD.n126 VDD.n125 1.35607
R414 VDD.n107 VDD.n106 1.35607
R415 VDD.n90 VDD.n89 1.35607
R416 VDD.n204 VDD.n203 1.2005
R417 VDD.n37 VDD.n36 1.14764
R418 VDD.n366 VDD.n365 1.04225
R419 VDD.n207 VDD.n206 1.04225
R420 VDD.n268 VDD.n267 1.04225
R421 VDD.n283 VDD.n282 1.04225
R422 VDD.n302 VDD.n301 1.04225
R423 VDD.n318 VDD.n317 1.04225
R424 VDD.n336 VDD.n335 1.04225
R425 VDD.n354 VDD.n353 1.04225
R426 VDD.n246 VDD.n245 0.866746
R427 VDD.n36 VDD.n35 0.850734
R428 VDD.n370 VDD.n194 0.731708
R429 VDD.n245 VDD.n244 0.715888
R430 VDD.n370 VDD.n369 0.43282
R431 VDD.n15 VDD.n14 0.225109
R432 VDD.n32 VDD.n31 0.223156
R433 VDD.n224 VDD.n223 0.221203
R434 VDD.n233 VDD.n232 0.221203
R435 VDD.n23 VDD.n22 0.217297
R436 VDD.n240 VDD.n239 0.189953
R437 VDD.n196 VDD.n195 0.117957
R438 VDD.n209 VDD.n208 0.115802
R439 VDD.n215 VDD.n214 0.115802
R440 VDD.n12 VDD.n11 0.113847
R441 VDD.n6 VDD.n5 0.10961
R442 VDD.n221 VDD.n220 0.0996379
R443 VDD.n256 VDD.n255 0.0539828
R444 VDD.n340 VDD.n339 0.0531724
R445 VDD.n306 VDD.n305 0.0531724
R446 VDD.n147 VDD.n146 0.0530763
R447 VDD.n44 VDD.n43 0.0530763
R448 VDD.n253 VDD.n252 0.0523621
R449 VDD.n250 VDD.n249 0.0523621
R450 VDD.n112 VDD.n111 0.0522797
R451 VDD.n38 VDD.n37 0.0522797
R452 VDD.n358 VDD.n357 0.0515517
R453 VDD.n288 VDD.n287 0.0515517
R454 VDD.n182 VDD.n181 0.0514831
R455 VDD.n78 VDD.n77 0.0514831
R456 VDD.n323 VDD.n322 0.0507414
R457 VDD.n272 VDD.n271 0.0507414
R458 VDD.n164 VDD.n163 0.0506864
R459 VDD.n130 VDD.n129 0.0506864
R460 VDD.n94 VDD.n93 0.0506864
R461 VDD.n60 VDD.n59 0.0506864
R462 VDD.n41 VDD.n40 0.0498898
R463 VDD.n247 VDD.n246 0.0462845
R464 VDD.n35 VDD.n32 0.0427461
R465 VDD.n189 VDD.n186 0.0415156
R466 VDD.n177 VDD.n169 0.0415156
R467 VDD.n176 VDD.n170 0.0415156
R468 VDD.n139 VDD.n134 0.0415156
R469 VDD.n141 VDD.n140 0.0415156
R470 VDD.n125 VDD.n117 0.0415156
R471 VDD.n124 VDD.n118 0.0415156
R472 VDD.n104 VDD.n98 0.0415156
R473 VDD.n106 VDD.n105 0.0415156
R474 VDD.n89 VDD.n83 0.0415156
R475 VDD.n88 VDD.n84 0.0415156
R476 VDD.n73 VDD.n65 0.0415156
R477 VDD.n72 VDD.n66 0.0415156
R478 VDD.n20 VDD.n15 0.0415156
R479 VDD.n22 VDD.n21 0.0415156
R480 VDD.n315 VDD.n310 0.0415156
R481 VDD.n317 VDD.n316 0.0415156
R482 VDD.n280 VDD.n276 0.0415156
R483 VDD.n282 VDD.n281 0.0415156
R484 VDD.n205 VDD.n200 0.0415156
R485 VDD.n230 VDD.n224 0.0415156
R486 VDD.n232 VDD.n231 0.0415156
R487 VDD.n237 VDD.n233 0.0415156
R488 VDD.n239 VDD.n238 0.0415156
R489 VDD.n244 VDD.n240 0.0415156
R490 VDD.n159 VDD.n152 0.0395625
R491 VDD.n158 VDD.n153 0.0395625
R492 VDD.n55 VDD.n49 0.0395625
R493 VDD.n24 VDD.n23 0.0395625
R494 VDD.n31 VDD.n30 0.0395625
R495 VDD.n351 VDD.n345 0.0395625
R496 VDD.n353 VDD.n352 0.0395625
R497 VDD.n299 VDD.n293 0.0395625
R498 VDD.n301 VDD.n300 0.0395625
R499 VDD.n267 VDD.n260 0.0395625
R500 VDD.n266 VDD.n261 0.0395625
R501 VDD.n365 VDD.n364 0.0376094
R502 VDD.n333 VDD.n328 0.0376094
R503 VDD.n335 VDD.n334 0.0376094
R504 VDD.n245 VDD.n222 0.0259356
R505 VDD.n318 VDD.n309 0.0231293
R506 VDD.n283 VDD.n275 0.0231293
R507 VDD.n208 VDD.n207 0.0231293
R508 VDD.n214 VDD.n213 0.0231293
R509 VDD.n220 VDD.n219 0.0231293
R510 VDD.n185 VDD.n184 0.0227458
R511 VDD.n168 VDD.n167 0.0227458
R512 VDD.n142 VDD.n133 0.0227458
R513 VDD.n116 VDD.n115 0.0227458
R514 VDD.n107 VDD.n97 0.0227458
R515 VDD.n82 VDD.n81 0.0227458
R516 VDD.n64 VDD.n63 0.0227458
R517 VDD.n5 VDD.n4 0.0227458
R518 VDD.n343 VDD.n342 0.0220517
R519 VDD.n354 VDD.n344 0.0220517
R520 VDD.n320 VDD.n308 0.0220517
R521 VDD.n291 VDD.n290 0.0220517
R522 VDD.n302 VDD.n292 0.0220517
R523 VDD.n285 VDD.n274 0.0220517
R524 VDD.n198 VDD.n197 0.0220517
R525 VDD.n211 VDD.n210 0.0220517
R526 VDD.n217 VDD.n216 0.0220517
R527 VDD.n36 VDD.n13 0.0218329
R528 VDD.n151 VDD.n150 0.0216864
R529 VDD.n144 VDD.n132 0.0216864
R530 VDD.n109 VDD.n96 0.0216864
R531 VDD.n48 VDD.n47 0.0216864
R532 VDD.n2 VDD.n1 0.0216864
R533 VDD.n11 VDD.n10 0.0216864
R534 VDD.n366 VDD.n360 0.0209741
R535 VDD.n326 VDD.n325 0.0209741
R536 VDD.n336 VDD.n327 0.0209741
R537 VDD.n192 VDD.n183 0.0206271
R538 VDD.n179 VDD.n166 0.0206271
R539 VDD.n127 VDD.n114 0.0206271
R540 VDD.n91 VDD.n80 0.0206271
R541 VDD.n75 VDD.n62 0.0206271
R542 VDD.n269 VDD.n258 0.0198966
R543 VDD.n161 VDD.n149 0.0195678
R544 VDD.n57 VDD.n46 0.0195678
R545 VDD.n8 VDD.n7 0.0195678
R546 VDD VDD.n370 0.0161119
R547 VDD.n367 VDD.n359 0.0144047
R548 VDD.n369 VDD.n368 0.0110345
R549 VDD.n357 VDD.n356 0.0110345
R550 VDD.n339 VDD.n338 0.0110345
R551 VDD.n322 VDD.n321 0.0110345
R552 VDD.n305 VDD.n304 0.0110345
R553 VDD.n287 VDD.n286 0.0110345
R554 VDD.n271 VDD.n270 0.0110345
R555 VDD.n255 VDD.n254 0.0110345
R556 VDD.n252 VDD.n251 0.0110345
R557 VDD.n249 VDD.n248 0.0110345
R558 VDD.n194 VDD.n193 0.0108559
R559 VDD.n181 VDD.n180 0.0108559
R560 VDD.n163 VDD.n162 0.0108559
R561 VDD.n146 VDD.n145 0.0108559
R562 VDD.n129 VDD.n128 0.0108559
R563 VDD.n111 VDD.n110 0.0108559
R564 VDD.n93 VDD.n92 0.0108559
R565 VDD.n77 VDD.n76 0.0108559
R566 VDD.n59 VDD.n58 0.0108559
R567 VDD.n43 VDD.n42 0.0108559
R568 VDD.n40 VDD.n39 0.0108559
R569 VDD.n365 VDD.n363 0.0102656
R570 VDD.n335 VDD.n333 0.0102656
R571 VDD.n258 VDD.n257 0.00912069
R572 VDD.n149 VDD.n148 0.00897458
R573 VDD.n46 VDD.n45 0.00897458
R574 VDD.n7 VDD.n6 0.00897458
R575 VDD.n166 VDD.n165 0.00791525
R576 VDD.n114 VDD.n113 0.00791525
R577 VDD.n80 VDD.n79 0.00791525
R578 VDD.n62 VDD.n61 0.00791525
R579 VDD.n13 VDD.n12 0.00791525
R580 VDD.n308 VDD.n307 0.00696552
R581 VDD.n274 VDD.n273 0.00696552
R582 VDD.n197 VDD.n196 0.00696552
R583 VDD.n210 VDD.n209 0.00696552
R584 VDD.n216 VDD.n215 0.00696552
R585 VDD.n132 VDD.n131 0.00685593
R586 VDD.n96 VDD.n95 0.00685593
R587 VDD.n1 VDD.n0 0.00685593
R588 VDD.n159 VDD.n158 0.00635938
R589 VDD.n55 VDD.n54 0.00635938
R590 VDD.n30 VDD.n24 0.00635938
R591 VDD.n353 VDD.n351 0.00635938
R592 VDD.n301 VDD.n299 0.00635938
R593 VDD.n267 VDD.n266 0.00635938
R594 VDD.n342 VDD.n341 0.00588793
R595 VDD.n290 VDD.n289 0.00588793
R596 VDD.n222 VDD.n221 0.00588793
R597 VDD.n325 VDD.n324 0.00481034
R598 VDD.n337 VDD.n326 0.00373276
R599 VDD.n268 VDD.n259 0.00373276
R600 VDD.n160 VDD.n151 0.00367797
R601 VDD.n56 VDD.n48 0.00367797
R602 VDD.n10 VDD.n9 0.00367797
R603 VDD.n367 VDD.n366 0.00265517
R604 VDD.n355 VDD.n354 0.00265517
R605 VDD.n337 VDD.n336 0.00265517
R606 VDD.n303 VDD.n302 0.00265517
R607 VDD.n269 VDD.n268 0.00265517
R608 VDD.n192 VDD.n191 0.00261864
R609 VDD.n179 VDD.n178 0.00261864
R610 VDD.n161 VDD.n160 0.00261864
R611 VDD.n127 VDD.n126 0.00261864
R612 VDD.n91 VDD.n90 0.00261864
R613 VDD.n75 VDD.n74 0.00261864
R614 VDD.n57 VDD.n56 0.00261864
R615 VDD.n9 VDD.n8 0.00261864
R616 VDD.n190 VDD.n189 0.00245312
R617 VDD.n177 VDD.n176 0.00245312
R618 VDD.n141 VDD.n139 0.00245312
R619 VDD.n125 VDD.n124 0.00245312
R620 VDD.n106 VDD.n104 0.00245312
R621 VDD.n89 VDD.n88 0.00245312
R622 VDD.n73 VDD.n72 0.00245312
R623 VDD.n21 VDD.n20 0.00245312
R624 VDD.n317 VDD.n315 0.00245312
R625 VDD.n282 VDD.n280 0.00245312
R626 VDD.n206 VDD.n205 0.00245312
R627 VDD.n231 VDD.n230 0.00245312
R628 VDD.n238 VDD.n237 0.00245312
R629 VDD.n355 VDD.n343 0.00157759
R630 VDD.n320 VDD.n319 0.00157759
R631 VDD.n319 VDD.n318 0.00157759
R632 VDD.n303 VDD.n291 0.00157759
R633 VDD.n285 VDD.n284 0.00157759
R634 VDD.n284 VDD.n283 0.00157759
R635 VDD.n199 VDD.n198 0.00157759
R636 VDD.n207 VDD.n199 0.00157759
R637 VDD.n212 VDD.n211 0.00157759
R638 VDD.n213 VDD.n212 0.00157759
R639 VDD.n218 VDD.n217 0.00157759
R640 VDD.n219 VDD.n218 0.00157759
R641 VDD.n191 VDD.n185 0.00155932
R642 VDD.n178 VDD.n168 0.00155932
R643 VDD.n144 VDD.n143 0.00155932
R644 VDD.n143 VDD.n142 0.00155932
R645 VDD.n126 VDD.n116 0.00155932
R646 VDD.n109 VDD.n108 0.00155932
R647 VDD.n108 VDD.n107 0.00155932
R648 VDD.n90 VDD.n82 0.00155932
R649 VDD.n74 VDD.n64 0.00155932
R650 VDD.n3 VDD.n2 0.00155932
R651 VDD.n4 VDD.n3 0.00155932
R652 VDD.n368 VDD.n358 0.00131035
R653 VDD.n356 VDD.n340 0.00131035
R654 VDD.n338 VDD.n323 0.00131035
R655 VDD.n321 VDD.n306 0.00131035
R656 VDD.n304 VDD.n288 0.00131035
R657 VDD.n286 VDD.n272 0.00131035
R658 VDD.n270 VDD.n256 0.00131035
R659 VDD.n254 VDD.n253 0.00131035
R660 VDD.n251 VDD.n250 0.00131035
R661 VDD.n248 VDD.n247 0.00131035
R662 VDD.n193 VDD.n182 0.00129661
R663 VDD.n180 VDD.n164 0.00129661
R664 VDD.n162 VDD.n147 0.00129661
R665 VDD.n145 VDD.n130 0.00129661
R666 VDD.n128 VDD.n112 0.00129661
R667 VDD.n110 VDD.n94 0.00129661
R668 VDD.n92 VDD.n78 0.00129661
R669 VDD.n76 VDD.n60 0.00129661
R670 VDD.n58 VDD.n44 0.00129661
R671 VDD.n42 VDD.n41 0.00129661
R672 VDD.n39 VDD.n38 0.00129661
R673 ready.n0 ready.t1 77.6295
R674 ready.n0 ready.t0 42.3121
R675 ready ready.n0 14.5094
R676 comp_outn.n0 comp_outn.t2 43.1877
R677 comp_outn.n1 comp_outn.t0 43.044
R678 comp_outn.n1 comp_outn.t1 43.044
R679 comp_outn comp_outn.t5 38.7789
R680 comp_outn.n4 comp_outn.t3 38.6969
R681 comp_outn.n4 comp_outn.t4 38.6969
R682 comp_outn.n2 comp_outn 1.15859
R683 comp_outn comp_outn.n4 0.984675
R684 comp_outn.n0 comp_outn 0.932565
R685 comp_outn.n5 comp_outn.n3 0.596088
R686 comp_outn.n5 comp_outn 0.438
R687 comp_outn.n2 comp_outn.n1 0.247153
R688 comp_outn comp_outn.n6 0.206382
R689 comp_outn.n3 comp_outn 0.15592
R690 comp_outn.n6 comp_outn 0.152674
R691 comp_outn.n6 comp_outn.n5 0.107118
R692 comp_outn.n2 comp_outn.n0 0.103441
R693 comp_outn.n5 comp_outn 0.063
R694 comp_outn.n3 comp_outn.n2 0.0193053
R695 comp_outp.n1 comp_outp.t2 43.3421
R696 comp_outp.n0 comp_outp.t0 43.044
R697 comp_outp.n0 comp_outp.t1 43.044
R698 comp_outp.n3 comp_outp.t5 39.1234
R699 comp_outp.n2 comp_outp.t3 38.6969
R700 comp_outp.n2 comp_outp.t4 38.6969
R701 comp_outp comp_outp.n4 14.0184
R702 comp_outp.n3 comp_outp.n2 1.09812
R703 comp_outp.n1 comp_outp.n0 1.00398
R704 comp_outp.n4 comp_outp.n3 0.449029
R705 comp_outp.n4 comp_outp.n1 0.294618
R706 clk.n4 clk.t4 356.68
R707 clk.n3 clk.t5 356.68
R708 clk.n1 clk.t1 269.921
R709 clk.n0 clk.t0 269.921
R710 clk.n4 clk.t2 202.44
R711 clk.n3 clk.t7 202.44
R712 clk.n1 clk.t6 195.721
R713 clk.n0 clk.t3 195.721
R714 clk.n5 clk.n4 41.3896
R715 clk.n5 clk.n3 41.3896
R716 clk.n2 clk.n0 38.0628
R717 clk.n2 clk.n1 38.0536
R718 clk.n6 clk.n5 12.3898
R719 clk clk.n6 8.69013
R720 clk.n6 clk.n2 3.40229
R721 cdac_vp.n0 cdac_vp.t6 340.613
R722 cdac_vp.n6 cdac_vp.t0 186.374
R723 cdac_vp.n5 cdac_vp.t7 186.374
R724 cdac_vp.n4 cdac_vp.t3 186.374
R725 cdac_vp.n3 cdac_vp.t1 186.374
R726 cdac_vp.n2 cdac_vp.t5 186.374
R727 cdac_vp.n1 cdac_vp.t4 186.374
R728 cdac_vp.n0 cdac_vp.t2 186.374
R729 cdac_vp.n1 cdac_vp.n0 154.24
R730 cdac_vp.n2 cdac_vp.n1 154.24
R731 cdac_vp.n3 cdac_vp.n2 154.24
R732 cdac_vp.n4 cdac_vp.n3 154.24
R733 cdac_vp.n5 cdac_vp.n4 154.24
R734 cdac_vp.n6 cdac_vp.n5 154.24
R735 cdac_vp cdac_vp.n6 102.329
C0 clk a_482_n1818# 0.171f
C1 a_582_n702# RS_p 2.32e-19
C2 Q cdac_vp 0.0548f
C3 a_1716_n1348# a_476_n1721# 0.0571f
C4 VDD RS_n 0.589f
C5 a_476_n1721# a_852_n296# 0.311f
C6 a_1566_n378# a_1248_n288# 0.406f
C7 a_1026_n1747# a_1716_n1348# 2.23e-21
C8 a_1566_n378# a_674_n702# 0.194f
C9 comp_outp a_1248_n288# 4.23e-21
C10 a_1026_n1747# a_852_n296# 0.0112f
C11 comp_outp a_674_n702# 1.74e-19
C12 a_1566_n378# VDD 0.804f
C13 a_564_n1266# cdac_vp 6.99e-19
C14 comp_outn RS_n 1.85e-19
C15 comp_outp VDD 0.67f
C16 VDD a_564_n1721# 0.159f
C17 a_582_n702# a_482_n1818# 0.0103f
C18 clk a_582_n702# 0.0987f
C19 Q a_1248_n288# 0.195f
C20 VDD a_1950_n1721# 0.771f
C21 cdac_vn a_476_n1721# 0.0373f
C22 Q a_674_n702# 0.00486f
C23 comp_outp comp_outn 0.053f
C24 comp_outn a_564_n1721# 8.24e-22
C25 Q VDD 0.368f
C26 a_1716_n1348# RS_n 0.133f
C27 a_852_n296# RS_n 0.0212f
C28 a_1026_n1747# cdac_vn 0.00935f
C29 ready a_476_n1721# 0.0403f
C30 cdac_vp a_1248_n288# 0.0204f
C31 comp_outn a_1950_n1721# 0.116f
C32 a_674_n702# cdac_vp 0.185f
C33 a_1026_n1747# ready 0.0571f
C34 a_1716_n1348# a_1566_n378# 0.137f
C35 VDD cdac_vp 0.0207f
C36 a_564_n1266# VDD 5.28e-20
C37 a_1566_n378# a_852_n296# 0.011f
C38 a_1716_n1348# comp_outp 0.0993f
C39 comp_outp a_852_n296# 0.105f
C40 a_476_n1721# RS_p 0.00222f
C41 a_1716_n1348# a_564_n1721# 1.33e-20
C42 a_852_n296# a_564_n1721# 0.00163f
C43 a_1026_n1747# RS_p 0.15f
C44 a_1716_n1348# a_1950_n1721# 0.011f
C45 cdac_vn RS_n 0.0068f
C46 a_1716_n1348# Q 0.141f
C47 a_674_n702# a_1248_n288# 0.133f
C48 Q a_852_n296# 0.00112f
C49 ready RS_n 0.0795f
C50 VDD a_1248_n288# 0.854f
C51 cdac_vn a_1566_n378# 0.00873f
C52 VDD a_674_n702# 0.368f
C53 cdac_vn comp_outp 0.0114f
C54 a_476_n1721# a_482_n1818# 1.63f
C55 a_1716_n1348# cdac_vp 0.0379f
C56 cdac_vp a_852_n296# 0.0836f
C57 a_476_n1721# clk 0.459f
C58 a_564_n1266# a_852_n296# 2.36e-21
C59 cdac_vn a_564_n1721# 0.00591f
C60 ready a_1566_n378# 6.39e-21
C61 ready comp_outp 1.69f
C62 a_1026_n1747# a_482_n1818# 4.38e-19
C63 RS_n RS_p 0.317f
C64 cdac_vn a_1950_n1721# 0.0164f
C65 ready a_564_n1721# 0.072f
C66 comp_outn VDD 0.608f
C67 cdac_vn Q 0.186f
C68 ready a_1950_n1721# 0.0553f
C69 a_1566_n378# RS_p 4.77e-20
C70 comp_outp RS_p 0.0757f
C71 a_564_n1721# RS_p 0.00308f
C72 a_1716_n1348# a_1248_n288# 0.00907f
C73 a_852_n296# a_1248_n288# 0.136f
C74 cdac_vn cdac_vp 0.574f
C75 a_1716_n1348# a_674_n702# 0.00112f
C76 cdac_vn a_564_n1266# 0.00183f
C77 a_674_n702# a_852_n296# 0.142f
C78 RS_n a_482_n1818# 6.34e-20
C79 a_476_n1721# a_582_n702# 0.0586f
C80 a_1950_n1721# RS_p 1.26e-19
C81 a_1716_n1348# VDD 0.791f
C82 VDD a_852_n296# 0.785f
C83 clk RS_n 0.00117f
C84 ready cdac_vp 8.68e-19
C85 a_1026_n1747# a_582_n702# 6e-19
C86 a_1566_n378# a_482_n1818# 0.0257f
C87 comp_outp a_482_n1818# 0.00372f
C88 a_1716_n1348# comp_outn 0.00481f
C89 a_1566_n378# clk 0.524f
C90 comp_outp clk 0.00305f
C91 a_564_n1721# a_482_n1818# 0.211f
C92 cdac_vp RS_p 5.9e-20
C93 cdac_vn a_1248_n288# 8.75e-19
C94 cdac_vn a_674_n702# 0.033f
C95 a_1950_n1721# a_482_n1818# 2.63e-20
C96 cdac_vn VDD 0.193f
C97 ready a_1248_n288# 3.55e-21
C98 ready a_674_n702# 1.77e-19
C99 Q a_482_n1818# 0.0238f
C100 a_582_n702# RS_n 1.86e-19
C101 a_1716_n1348# a_852_n296# 0.215f
C102 Q clk 0.113f
C103 ready VDD 0.616f
C104 cdac_vn comp_outn 0.00607f
C105 cdac_vp a_482_n1818# 0.224f
C106 a_1566_n378# a_582_n702# 0.00927f
C107 a_1248_n288# RS_p 2.46e-19
C108 a_564_n1266# a_482_n1818# 0.0165f
C109 a_674_n702# RS_p 1e-19
C110 comp_outp a_582_n702# 0.00255f
C111 clk cdac_vp 0.615f
C112 ready comp_outn 0.0692f
C113 VDD RS_p 0.544f
C114 a_582_n702# a_564_n1721# 3.35e-19
C115 a_582_n702# a_1950_n1721# 5.99e-19
C116 a_1026_n1747# a_476_n1721# 0.00775f
C117 a_1716_n1348# cdac_vn 0.0917f
C118 cdac_vn a_852_n296# 0.0564f
C119 Q a_582_n702# 1.53f
C120 comp_outn RS_p 8.63e-21
C121 ready a_852_n296# 5.96e-19
C122 a_1248_n288# a_482_n1818# 0.0534f
C123 a_674_n702# a_482_n1818# 0.0145f
C124 clk a_1248_n288# 0.601f
C125 clk a_674_n702# 0.0975f
C126 VDD a_482_n1818# 1.47f
C127 cdac_vp a_582_n702# 0.237f
C128 clk VDD 0.777f
C129 a_1716_n1348# RS_p 0.0744f
C130 a_852_n296# RS_p 0.158f
C131 a_476_n1721# RS_n 0.00191f
C132 comp_outn a_482_n1818# 1.01e-21
C133 a_1026_n1747# RS_n 7.23e-19
C134 ready cdac_vn 0.00511f
C135 a_1566_n378# a_476_n1721# 0.116f
C136 comp_outp a_476_n1721# 0.0165f
C137 a_582_n702# a_1248_n288# 0.00778f
C138 a_674_n702# a_582_n702# 1.53f
C139 a_476_n1721# a_564_n1721# 0.389f
C140 a_1026_n1747# comp_outp 0.17f
C141 a_1716_n1348# a_482_n1818# 0.197f
C142 VDD a_582_n702# 0.0163f
C143 a_852_n296# a_482_n1818# 0.042f
C144 a_476_n1721# a_1950_n1721# 5.72e-19
C145 cdac_vn RS_p 0.00689f
C146 a_1026_n1747# a_564_n1721# 0.0216f
C147 a_1716_n1348# clk 0.112f
C148 clk a_852_n296# 0.0265f
C149 Q a_476_n1721# 0.00925f
C150 a_1026_n1747# a_1950_n1721# 1.46e-19
C151 ready RS_p 0.0657f
C152 a_476_n1721# cdac_vp 0.541f
C153 a_1566_n378# RS_n 1.34e-19
C154 a_564_n1266# a_476_n1721# 0.0214f
C155 comp_outp RS_n 0.0437f
C156 cdac_vn a_482_n1818# 0.0389f
C157 a_1026_n1747# cdac_vp 0.00723f
C158 a_564_n1721# RS_n 3.53e-20
C159 a_1026_n1747# a_564_n1266# 1.65e-20
C160 cdac_vn clk 0.0627f
C161 a_1716_n1348# a_582_n702# 0.0741f
C162 a_582_n702# a_852_n296# 0.0742f
C163 ready a_482_n1818# 8.24e-20
C164 a_1950_n1721# RS_n 0.149f
C165 a_1566_n378# comp_outp 6.13e-21
C166 ready clk 2.93e-20
C167 Q RS_n 7.8e-20
C168 comp_outp a_564_n1721# 0.00587f
C169 a_476_n1721# a_1248_n288# 0.109f
C170 a_476_n1721# a_674_n702# 0.0774f
C171 comp_outp a_1950_n1721# 0.0559f
C172 RS_p a_482_n1818# 8.41e-20
C173 a_1566_n378# Q 0.156f
C174 a_476_n1721# VDD 0.799f
C175 cdac_vp RS_n 6.35e-20
C176 clk RS_p 0.00116f
C177 a_1950_n1721# a_564_n1721# 3.46e-21
C178 a_1026_n1747# a_674_n702# 3.37e-19
C179 Q comp_outp 7.85e-19
C180 cdac_vn a_582_n702# 0.379f
C181 a_1026_n1747# VDD 0.767f
C182 a_1566_n378# cdac_vp 0.019f
C183 a_476_n1721# comp_outn 1.55e-19
C184 Q a_1950_n1721# 3.37e-19
C185 ready a_582_n702# 2.06e-19
C186 comp_outp cdac_vp 0.00134f
C187 cdac_vp a_564_n1721# 0.00284f
C188 a_564_n1266# a_564_n1721# 0.161f
.ends

