* NGSPICE file created from hgu_comp_flat.ext - technology: sky130A

.subckt hgu_comp ready cdac_vn comp_outp comp_outn cdac_vp clk VDD VSS
X0 Q cdac_vn.t0 a_582_n702# VSS.t42 sky130_fd_pr__nfet_01v8_lvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1 ready.t0 a_564_n1721# VDD.t39 VDD.t38 sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0.244 ps=2.26 w=0.84 l=0.15
X2 a_564_n1721# a_476_n1721# a_564_n1266# VSS.t12 sky130_fd_pr__nfet_01v8 ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.15
X3 comp_outn.t2 a_1950_n1721# VDD.t25 VDD.t24 sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.3 as=0.139 ps=1.17 w=0.84 l=0.15
X4 a_582_n702# cdac_vn.t1 Q VSS.t41 sky130_fd_pr__nfet_01v8_lvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X5 a_1950_n1721# RS_n VDD.t3 VDD.t2 sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0.244 ps=2.26 w=0.84 l=0.15
X6 a_482_n1818# a_1716_n1348# VSS.t62 VSS.t61 sky130_fd_pr__nfet_01v8 ad=0.0759 pd=0.79 as=0.143 ps=1.54 w=0.46 l=0.15
X7 a_564_n1721# a_482_n1818# a_476_n1721# VDD.t13 sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.15
X8 VDD.t19 a_1026_n1747# comp_outp.t2 VDD.t18 sky130_fd_pr__pfet_01v8 ad=0.139 pd=1.17 as=0.26 ps=2.3 w=0.84 l=0.15
X9 VSS.t65 RS_p a_1026_n1747# VSS.t64 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X10 VDD.t5 clk.t0 a_1248_n288# VDD.t4 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X11 a_674_n702# cdac_vp.t0 a_582_n702# VSS.t63 sky130_fd_pr__nfet_01v8_lvt ad=0.165 pd=1.33 as=0.31 ps=2.62 w=1 l=0.15
X12 VDD.t31 a_852_n296# a_476_n1721# VDD.t30 sky130_fd_pr__pfet_01v8 ad=0.139 pd=1.17 as=0.26 ps=2.3 w=0.84 l=0.15
X13 comp_outp.t1 a_1026_n1747# VDD.t17 VDD.t16 sky130_fd_pr__pfet_01v8 ad=0.139 pd=1.17 as=0.139 ps=1.17 w=0.84 l=0.15
X14 a_476_n1721# a_852_n296# VDD.t29 VDD.t28 sky130_fd_pr__pfet_01v8 ad=0.139 pd=1.17 as=0.139 ps=1.17 w=0.84 l=0.15
X15 a_582_n702# cdac_vn.t2 Q VSS.t40 sky130_fd_pr__nfet_01v8_lvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X16 a_582_n702# cdac_vp.t1 a_674_n702# VSS.t54 sky130_fd_pr__nfet_01v8_lvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X17 comp_outn.t5 a_1950_n1721# VSS.t26 VSS.t25 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.54 as=0.0759 ps=0.79 w=0.46 l=0.15
X18 VDD.t51 RS_p a_1026_n1747# VDD.t50 sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0.244 ps=2.26 w=0.84 l=0.15
X19 VDD.t27 a_852_n296# a_476_n1721# VDD.t26 sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.3 as=0.139 ps=1.17 w=0.84 l=0.15
X20 a_674_n702# cdac_vp.t2 a_582_n702# VSS.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X21 Q cdac_vn.t3 a_582_n702# VSS.t39 sky130_fd_pr__nfet_01v8_lvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X22 a_564_n1266# a_482_n1818# VSS.t14 VSS.t13 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.15
X23 VSS.t20 a_1026_n1747# comp_outp.t5 VSS.t19 sky130_fd_pr__nfet_01v8 ad=0.0759 pd=0.79 as=0.143 ps=1.54 w=0.46 l=0.15
X24 a_1950_n1721# RS_n VSS.t3 VSS.t2 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X25 a_1566_n378# clk.t1 VDD.t37 VDD.t36 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X26 VSS.t34 a_852_n296# a_476_n1721# VSS.t33 sky130_fd_pr__nfet_01v8 ad=0.0759 pd=0.79 as=0.143 ps=1.54 w=0.46 l=0.15
X27 VDD.t11 a_1248_n288# a_852_n296# VDD.t10 sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0.244 ps=2.26 w=0.84 l=0.15
X28 a_482_n1818# a_1716_n1348# VSS.t60 VSS.t59 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.54 as=0.0759 ps=0.79 w=0.46 l=0.15
X29 a_582_n702# clk.t2 VSS.t50 VSS.t49 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X30 comp_outp.t4 a_1026_n1747# VSS.t18 VSS.t17 sky130_fd_pr__nfet_01v8 ad=0.0759 pd=0.79 as=0.0759 ps=0.79 w=0.46 l=0.15
X31 VSS.t11 a_1248_n288# a_852_n296# VSS.t10 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X32 a_674_n702# cdac_vp.t3 a_582_n702# VSS.t48 sky130_fd_pr__nfet_01v8_lvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X33 a_582_n702# cdac_vn.t4 Q VSS.t38 sky130_fd_pr__nfet_01v8_lvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X34 a_1248_n288# a_1566_n378# VDD.t35 VDD.t34 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X35 Q clk.t3 VDD.t7 VDD.t6 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X36 a_582_n702# cdac_vp.t4 a_674_n702# VSS.t51 sky130_fd_pr__nfet_01v8_lvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X37 VDD.t15 a_1026_n1747# comp_outp.t0 VDD.t14 sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.3 as=0.139 ps=1.17 w=0.84 l=0.15
X38 RS_n a_1716_n1348# VSS.t58 VSS.t46 sky130_fd_pr__nfet_01v8 ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.15
X39 comp_outn.t1 a_1950_n1721# VDD.t23 VDD.t22 sky130_fd_pr__pfet_01v8 ad=0.139 pd=1.17 as=0.26 ps=2.3 w=0.84 l=0.15
X40 a_1716_n1348# a_1566_n378# VSS.t45 VSS.t44 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X41 VSS.t57 a_1716_n1348# a_482_n1818# VSS.t56 sky130_fd_pr__nfet_01v8 ad=0.0759 pd=0.79 as=0.0759 ps=0.79 w=0.46 l=0.15
X42 VSS.t8 clk.t4 a_582_n702# VSS.t7 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.31 ps=2.62 w=1 l=0.15
X43 a_582_n702# cdac_vn.t5 Q VSS.t37 sky130_fd_pr__nfet_01v8_lvt ad=0.31 pd=2.62 as=0.165 ps=1.33 w=1 l=0.15
X44 VSS.t32 a_852_n296# a_476_n1721# VSS.t31 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.54 as=0.0759 ps=0.79 w=0.46 l=0.15
X45 Q a_1566_n378# a_1248_n288# VSS.t43 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X46 Q cdac_vn.t6 a_582_n702# VSS.t36 sky130_fd_pr__nfet_01v8_lvt ad=0.165 pd=1.33 as=0.31 ps=2.62 w=1 l=0.15
X47 RS_n RS_p VDD.t49 VDD.t48 sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.15
X48 VDD.t21 a_1950_n1721# comp_outn.t0 VDD.t20 sky130_fd_pr__pfet_01v8 ad=0.139 pd=1.17 as=0.139 ps=1.17 w=0.84 l=0.15
X49 a_1716_n1348# a_1566_n378# VDD.t33 VDD.t32 sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0.244 ps=2.26 w=0.84 l=0.15
X50 a_582_n702# clk.t5 VSS.t1 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.165 ps=1.33 w=1 l=0.15
X51 VDD.t47 clk.t6 a_674_n702# VDD.t46 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X52 a_674_n702# cdac_vp.t5 a_582_n702# VSS.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X53 VSS.t16 a_1026_n1747# comp_outp.t3 VSS.t15 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.54 as=0.0759 ps=0.79 w=0.46 l=0.15
X54 comp_outn.t4 a_1950_n1721# VSS.t24 VSS.t23 sky130_fd_pr__nfet_01v8 ad=0.0759 pd=0.79 as=0.143 ps=1.54 w=0.46 l=0.15
X55 a_482_n1818# a_1716_n1348# VDD.t45 VDD.t44 sky130_fd_pr__pfet_01v8 ad=0.139 pd=1.17 as=0.26 ps=2.3 w=0.84 l=0.15
X56 a_482_n1818# a_1716_n1348# VDD.t43 VDD.t42 sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.3 as=0.139 ps=1.17 w=0.84 l=0.15
X57 a_582_n702# cdac_vp.t6 a_674_n702# VSS.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.31 pd=2.62 as=0.165 ps=1.33 w=1 l=0.15
X58 VSS.t30 a_852_n296# RS_p VSS.t29 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.15
X59 VDD.t41 a_1716_n1348# a_482_n1818# VDD.t40 sky130_fd_pr__pfet_01v8 ad=0.139 pd=1.17 as=0.139 ps=1.17 w=0.84 l=0.15
X60 Q cdac_vn.t7 a_582_n702# VSS.t35 sky130_fd_pr__nfet_01v8_lvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X61 ready.t1 a_564_n1721# VSS.t53 VSS.t52 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X62 a_482_n1818# a_476_n1721# a_564_n1721# VDD.t12 sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.15
X63 VSS.t22 a_1950_n1721# comp_outn.t3 VSS.t21 sky130_fd_pr__nfet_01v8 ad=0.0759 pd=0.79 as=0.0759 ps=0.79 w=0.46 l=0.15
X64 a_476_n1721# a_852_n296# VSS.t28 VSS.t27 sky130_fd_pr__nfet_01v8 ad=0.0759 pd=0.79 as=0.0759 ps=0.79 w=0.46 l=0.15
X65 VDD.t9 a_1248_n288# a_1566_n378# VDD.t8 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X66 a_1566_n378# a_1248_n288# a_674_n702# VSS.t9 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X67 a_582_n702# cdac_vp.t7 a_674_n702# VSS.t55 sky130_fd_pr__nfet_01v8_lvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X68 VSS.t47 clk.t7 a_582_n702# VSS.t46 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X69 VDD.t1 RS_n RS_p VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.15
R0 cdac_vn.n0 cdac_vn.t6 340.613
R1 cdac_vn.n6 cdac_vn.t5 186.374
R2 cdac_vn.n0 cdac_vn.t2 186.374
R3 cdac_vn.n1 cdac_vn.t0 186.374
R4 cdac_vn.n2 cdac_vn.t4 186.374
R5 cdac_vn.n3 cdac_vn.t3 186.374
R6 cdac_vn.n4 cdac_vn.t1 186.374
R7 cdac_vn.n5 cdac_vn.t7 186.374
R8 cdac_vn.n6 cdac_vn.n5 154.24
R9 cdac_vn.n5 cdac_vn.n4 154.24
R10 cdac_vn.n4 cdac_vn.n3 154.24
R11 cdac_vn.n3 cdac_vn.n2 154.24
R12 cdac_vn.n2 cdac_vn.n1 154.24
R13 cdac_vn.n1 cdac_vn.n0 154.24
R14 cdac_vn cdac_vn.n6 102.109
R15 VSS.n63 VSS.t36 179.739
R16 VSS.n68 VSS.t2 179.739
R17 VSS.n87 VSS.t49 179.739
R18 VSS.n92 VSS.t64 172.549
R19 VSS.n106 VSS.t15 172.549
R20 VSS.n53 VSS.t23 165.359
R21 VSS.n101 VSS.t5 165.359
R22 VSS.n106 VSS.t51 165.359
R23 VSS.n81 VSS.t46 165.359
R24 VSS.n81 VSS.t29 150.981
R25 VSS.n52 VSS.t42 143.792
R26 VSS.n156 VSS.t13 129.412
R27 VSS.n87 VSS.t9 122.222
R28 VSS.n75 VSS.t43 107.844
R29 VSS.n160 VSS.t55 107.844
R30 VSS.t44 VSS.t40 100.654
R31 VSS.n5 VSS.t35 93.4646
R32 VSS.n112 VSS.t31 93.4646
R33 VSS.n163 VSS.t63 93.4646
R34 VSS.n18 VSS.t45 86.7771
R35 VSS.n122 VSS.t11 85.4529
R36 VSS.n155 VSS.t14 83.725
R37 VSS.n14 VSS.t62 80.7031
R38 VSS.n126 VSS.t32 80.7031
R39 VSS.n103 VSS.t16 80.7031
R40 VSS.n57 VSS.t24 80.7031
R41 VSS.n148 VSS.t53 80.5977
R42 VSS.n94 VSS.t65 80.5977
R43 VSS.n67 VSS.t3 80.5977
R44 VSS.n0 VSS.t37 79.0855
R45 VSS.n101 VSS.t10 79.0855
R46 VSS.n116 VSS.t27 79.0855
R47 VSS.t63 VSS.t12 79.0855
R48 VSS.n45 VSS.t61 71.8959
R49 VSS.n74 VSS.n73 71.5328
R50 VSS.n86 VSS.n85 71.5328
R51 VSS.n143 VSS.t33 64.7064
R52 VSS.t59 VSS.t41 57.5168
R53 VSS.t56 VSS.t39 57.5168
R54 VSS.n40 VSS.t56 57.5168
R55 VSS.t61 VSS.t38 57.5168
R56 VSS.n58 VSS.t44 57.5168
R57 VSS.t31 VSS.t4 57.5168
R58 VSS.t27 VSS.t54 57.5168
R59 VSS.t33 VSS.t48 57.5168
R60 VSS.n80 VSS.n79 51.9572
R61 VSS.t48 VSS.t52 50.3273
R62 VSS.n34 VSS.t59 43.1378
R63 VSS.t43 VSS.t0 43.1378
R64 VSS.t9 VSS.t7 43.1378
R65 VSS.n10 VSS.t60 43.044
R66 VSS.n10 VSS.t57 43.044
R67 VSS.n134 VSS.t28 43.044
R68 VSS.n134 VSS.t34 43.044
R69 VSS.n110 VSS.t18 43.044
R70 VSS.n110 VSS.t20 43.044
R71 VSS.n48 VSS.t26 43.044
R72 VSS.n48 VSS.t22 43.044
R73 VSS.n11 VSS.n10 37.6596
R74 VSS.n135 VSS.n134 37.6596
R75 VSS.n111 VSS.n110 37.6596
R76 VSS.n49 VSS.n48 37.6596
R77 VSS.t38 VSS.t25 28.7587
R78 VSS.t42 VSS.t21 28.7587
R79 VSS.n79 VSS.t58 20.7148
R80 VSS.n79 VSS.t30 20.7148
R81 VSS.n73 VSS.t1 19.8005
R82 VSS.n73 VSS.t47 19.8005
R83 VSS.n85 VSS.t50 19.8005
R84 VSS.n85 VSS.t8 19.8005
R85 VSS.n137 VSS.n136 9.15497
R86 VSS.n124 VSS.n123 9.15497
R87 VSS.n128 VSS.n127 9.15497
R88 VSS.n131 VSS.n130 9.15497
R89 VSS.n16 VSS.n15 9.15497
R90 VSS.n20 VSS.n19 9.15497
R91 VSS.n18 VSS.n17 9.15497
R92 VSS.n13 VSS.n12 9.15497
R93 VSS.n24 VSS.n23 9.15497
R94 VSS.n122 VSS.n121 9.15497
R95 VSS.n155 VSS.n154 9.15497
R96 VSS.n151 VSS.n150 9.15497
R97 VSS.n150 VSS.n149 9.15497
R98 VSS.n162 VSS.n161 9.15497
R99 VSS.n161 VSS.n160 9.15497
R100 VSS.n13 VSS.n11 7.94533
R101 VSS.n35 VSS.n34 7.19004
R102 VSS.n41 VSS.n40 7.19004
R103 VSS.n46 VSS.n45 7.19004
R104 VSS.n53 VSS.n52 7.19004
R105 VSS.n59 VSS.n58 7.19004
R106 VSS.t15 VSS.t6 7.19004
R107 VSS.t51 VSS.t17 7.19004
R108 VSS.t4 VSS.t19 7.19004
R109 VSS.n137 VSS.n135 6.62119
R110 VSS.n16 VSS.n14 6.17981
R111 VSS.n4 VSS.n3 5.65173
R112 VSS.n165 VSS.n162 4.99852
R113 VSS.n128 VSS.n126 4.85567
R114 VSS.n22 VSS.n16 4.6505
R115 VSS.n132 VSS.n131 4.6505
R116 VSS.n129 VSS.n128 4.6505
R117 VSS.n25 VSS.n24 4.6505
R118 VSS.n152 VSS.n151 4.6505
R119 VSS.n162 VSS.n153 4.6505
R120 VSS.n2 VSS.n1 4.57773
R121 VSS.n1 VSS.n0 4.57773
R122 VSS.n7 VSS.n6 4.57773
R123 VSS.n6 VSS.n5 4.57773
R124 VSS.n37 VSS.n36 4.57773
R125 VSS.n36 VSS.n35 4.57773
R126 VSS.n43 VSS.n42 4.57773
R127 VSS.n42 VSS.n41 4.57773
R128 VSS.n50 VSS.n47 4.57773
R129 VSS.n47 VSS.n46 4.57773
R130 VSS.n55 VSS.n54 4.57773
R131 VSS.n54 VSS.n53 4.57773
R132 VSS.n61 VSS.n60 4.57773
R133 VSS.n60 VSS.n59 4.57773
R134 VSS.n65 VSS.n64 4.57773
R135 VSS.n64 VSS.n63 4.57773
R136 VSS.n70 VSS.n69 4.57773
R137 VSS.n69 VSS.n68 4.57773
R138 VSS.n77 VSS.n76 4.57773
R139 VSS.n76 VSS.n75 4.57773
R140 VSS.n83 VSS.n82 4.57773
R141 VSS.n82 VSS.n81 4.57773
R142 VSS.n89 VSS.n88 4.57773
R143 VSS.n88 VSS.n87 4.57773
R144 VSS.n95 VSS.n93 4.57773
R145 VSS.n93 VSS.n92 4.57773
R146 VSS.n99 VSS.n98 4.57773
R147 VSS.n98 VSS.n97 4.57773
R148 VSS.n104 VSS.n102 4.57773
R149 VSS.n102 VSS.n101 4.57773
R150 VSS.n108 VSS.n107 4.57773
R151 VSS.n107 VSS.n106 4.57773
R152 VSS.n114 VSS.n113 4.57773
R153 VSS.n113 VSS.n112 4.57773
R154 VSS.n118 VSS.n117 4.57773
R155 VSS.n117 VSS.n116 4.57773
R156 VSS.n145 VSS.n144 4.57773
R157 VSS.n144 VSS.n143 4.57773
R158 VSS.n158 VSS.n157 4.57773
R159 VSS.n157 VSS.n156 4.57773
R160 VSS.n165 VSS.n164 4.57773
R161 VSS.n164 VSS.n163 4.57773
R162 VSS.n21 VSS.n18 3.40067
R163 VSS.n125 VSS.n122 3.40067
R164 VSS.n125 VSS.n124 3.25009
R165 VSS.n21 VSS.n20 3.25009
R166 VSS.n28 VSS.n13 3.03426
R167 VSS.n138 VSS.n137 3.03311
R168 VSS.n8 VSS.n7 2.3255
R169 VSS.n44 VSS.n43 2.3255
R170 VSS.n51 VSS.n50 2.3255
R171 VSS.n56 VSS.n55 2.3255
R172 VSS.n62 VSS.n61 2.3255
R173 VSS.n66 VSS.n65 2.3255
R174 VSS.n71 VSS.n70 2.3255
R175 VSS.n78 VSS.n77 2.3255
R176 VSS.n84 VSS.n83 2.3255
R177 VSS.n90 VSS.n89 2.3255
R178 VSS.n96 VSS.n95 2.3255
R179 VSS.n100 VSS.n99 2.3255
R180 VSS.n105 VSS.n104 2.3255
R181 VSS.n109 VSS.n108 2.3255
R182 VSS.n115 VSS.n114 2.3255
R183 VSS.n119 VSS.n118 2.3255
R184 VSS.n166 VSS.n165 2.3255
R185 VSS.n33 VSS.n32 2.2505
R186 VSS.n140 VSS.n139 2.24128
R187 VSS.n31 VSS.n30 1.84746
R188 VSS.n141 VSS.n140 1.84746
R189 VSS.n38 VSS.n37 1.83603
R190 VSS.n146 VSS.n145 1.83603
R191 VSS.n29 VSS.n28 1.50988
R192 VSS.n166 VSS.n159 1.24358
R193 VSS.n142 VSS.n141 1.16147
R194 VSS.n159 VSS.n155 1.11247
R195 VSS.n4 VSS.n2 1.05718
R196 VSS.n22 VSS.n21 0.932839
R197 VSS.n129 VSS.n125 0.932839
R198 VSS.n8 VSS.n4 0.678677
R199 VSS.n159 VSS.n158 0.548468
R200 VSS.n72 VSS 0.441811
R201 VSS.n91 VSS 0.414118
R202 VSS.n77 VSS.n74 0.312695
R203 VSS.n151 VSS.n148 0.234646
R204 VSS.n61 VSS.n57 0.234646
R205 VSS.n70 VSS.n67 0.234646
R206 VSS.n25 VSS.n22 0.216017
R207 VSS.n132 VSS.n129 0.216017
R208 VSS.n133 VSS.n132 0.187208
R209 VSS.n26 VSS.n25 0.166381
R210 VSS.n95 VSS.n94 0.156598
R211 VSS.n104 VSS.n103 0.156598
R212 VSS.n114 VSS.n111 0.156598
R213 VSS.n83 VSS.n80 0.104565
R214 VSS.n89 VSS.n86 0.104565
R215 VSS.n50 VSS.n49 0.0785488
R216 VSS.n84 VSS.n78 0.051313
R217 VSS.n90 VSS.n84 0.051313
R218 VSS.n27 VSS.n26 0.0415156
R219 VSS.n51 VSS.n44 0.0386098
R220 VSS.n56 VSS.n51 0.0386098
R221 VSS.n62 VSS.n56 0.0386098
R222 VSS.n66 VSS.n62 0.0386098
R223 VSS.n71 VSS.n66 0.0386098
R224 VSS.n78 VSS.n72 0.0386098
R225 VSS.n100 VSS.n96 0.0386098
R226 VSS.n105 VSS.n100 0.0386098
R227 VSS.n109 VSS.n105 0.0386098
R228 VSS.n115 VSS.n109 0.0386098
R229 VSS.n119 VSS.n115 0.0386098
R230 VSS.n142 VSS.n119 0.0382053
R231 VSS.n32 VSS.n31 0.0356562
R232 VSS.n91 VSS.n90 0.035561
R233 VSS.n44 VSS.n39 0.0351228
R234 VSS.n167 VSS 0.0325248
R235 VSS.n9 VSS.n8 0.0302256
R236 VSS.n152 VSS.n147 0.0298445
R237 VSS.n30 VSS.n29 0.0263062
R238 VSS.n140 VSS.n120 0.0263062
R239 VSS VSS.n167 0.024128
R240 VSS.n139 VSS.n133 0.0215034
R241 VSS.n96 VSS.n91 0.012314
R242 VSS.n72 VSS.n71 0.0100274
R243 VSS VSS.n166 0.00928099
R244 VSS.n33 VSS.n9 0.00850305
R245 VSS.n147 VSS.n146 0.00850305
R246 VSS.n167 VSS.n153 0.00850305
R247 VSS.n39 VSS.n38 0.00497985
R248 VSS.n146 VSS.n142 0.00389195
R249 VSS.n139 VSS.n138 0.00245312
R250 VSS.n28 VSS.n27 0.0023033
R251 VSS.n153 VSS.n152 0.00126219
R252 VSS.n38 VSS.n33 0.000881098
R253 VDD.n0 VDD.t12 378.817
R254 VDD.t12 VDD.t13 163.237
R255 VDD.n99 VDD.t26 112.871
R256 VDD.n57 VDD.t44 112.871
R257 VDD.n39 VDD.t22 112.871
R258 VDD.n3 VDD.t18 103.466
R259 VDD.n2 VDD.t39 96.2456
R260 VDD.n98 VDD.t27 91.0302
R261 VDD.n61 VDD.t45 91.0302
R262 VDD.n38 VDD.t23 91.0302
R263 VDD.n13 VDD.t15 91.0302
R264 VDD.n79 VDD.t4 89.3422
R265 VDD.n18 VDD.t51 87.8456
R266 VDD.n23 VDD.t0 86.3641
R267 VDD.n93 VDD.t11 86.3397
R268 VDD.n66 VDD.t33 86.3397
R269 VDD.n33 VDD.t3 86.3397
R270 VDD.n14 VDD.t14 84.654
R271 VDD.n109 VDD.t30 84.1029
R272 VDD.n49 VDD.t24 84.1029
R273 VDD.n83 VDD.t36 71.4739
R274 VDD.n52 VDD.t42 65.291
R275 VDD.n83 VDD.t8 59.5616
R276 VDD.n88 VDD.n87 58.3564
R277 VDD.n78 VDD.n77 58.3564
R278 VDD.n74 VDD.n73 58.3564
R279 VDD.n67 VDD.t32 53.6055
R280 VDD.n106 VDD.n105 52.3338
R281 VDD.n56 VDD.n55 52.3338
R282 VDD.n44 VDD.n43 52.3338
R283 VDD.n28 VDD.n27 52.3338
R284 VDD.n8 VDD.n7 52.3338
R285 VDD.n29 VDD.t48 47.5005
R286 VDD.n79 VDD.t34 41.6933
R287 VDD.n105 VDD.t29 38.6969
R288 VDD.n105 VDD.t31 38.6969
R289 VDD.n55 VDD.t43 38.6969
R290 VDD.n55 VDD.t41 38.6969
R291 VDD.n43 VDD.t25 38.6969
R292 VDD.n43 VDD.t21 38.6969
R293 VDD.n7 VDD.t17 38.6969
R294 VDD.n7 VDD.t19 38.6969
R295 VDD.n57 VDD.t40 37.6243
R296 VDD.n94 VDD.t10 35.7372
R297 VDD.n34 VDD.t2 35.3521
R298 VDD.n27 VDD.t49 34.0065
R299 VDD.n27 VDD.t1 34.0065
R300 VDD.n89 VDD.t46 29.7811
R301 VDD.n87 VDD.t37 28.5655
R302 VDD.n87 VDD.t47 28.5655
R303 VDD.n77 VDD.t35 28.5655
R304 VDD.n77 VDD.t9 28.5655
R305 VDD.n73 VDD.t7 28.5655
R306 VDD.n73 VDD.t5 28.5655
R307 VDD.n103 VDD.t28 18.8124
R308 VDD.n45 VDD.t20 18.8124
R309 VDD.n54 VDD.n51 15.515
R310 VDD.n59 VDD.n56 14.4005
R311 VDD.n81 VDD.n78 14.4005
R312 VDD.n31 VDD.n28 13.6005
R313 VDD.n91 VDD.n88 12.8005
R314 VDD.n107 VDD.n106 12.0005
R315 VDD.n47 VDD.n44 12.0005
R316 VDD.n71 VDD.t6 11.9127
R317 VDD.n20 VDD.n19 10.7543
R318 VDD.n75 VDD.n74 10.4005
R319 VDD.n1 VDD.n0 9.99493
R320 VDD.n9 VDD.t16 9.40644
R321 VDD.n53 VDD.n52 8.85536
R322 VDD.n47 VDD.n46 8.85536
R323 VDD.n46 VDD.n45 8.85536
R324 VDD.n2 VDD.n1 8.85536
R325 VDD.n41 VDD.n40 8.85536
R326 VDD.n40 VDD.n39 8.85536
R327 VDD.n36 VDD.n35 8.85536
R328 VDD.n35 VDD.n34 8.85536
R329 VDD.n31 VDD.n30 8.85536
R330 VDD.n30 VDD.n29 8.85536
R331 VDD.n25 VDD.n24 8.85536
R332 VDD.n24 VDD.n23 8.85536
R333 VDD.n21 VDD.n20 8.85536
R334 VDD.n16 VDD.n15 8.85536
R335 VDD.n15 VDD.n14 8.85536
R336 VDD.n11 VDD.n10 8.85536
R337 VDD.n10 VDD.n9 8.85536
R338 VDD.n5 VDD.n4 8.85536
R339 VDD.n4 VDD.n3 8.85536
R340 VDD.n50 VDD.n49 8.85536
R341 VDD.n59 VDD.n58 8.85536
R342 VDD.n58 VDD.n57 8.85536
R343 VDD.n64 VDD.n63 8.85536
R344 VDD.n63 VDD.n62 8.85536
R345 VDD.n69 VDD.n68 8.85536
R346 VDD.n68 VDD.n67 8.85536
R347 VDD.n75 VDD.n72 8.85536
R348 VDD.n72 VDD.n71 8.85536
R349 VDD.n81 VDD.n80 8.85536
R350 VDD.n80 VDD.n79 8.85536
R351 VDD.n85 VDD.n84 8.85536
R352 VDD.n84 VDD.n83 8.85536
R353 VDD.n91 VDD.n90 8.85536
R354 VDD.n90 VDD.n89 8.85536
R355 VDD.n96 VDD.n95 8.85536
R356 VDD.n95 VDD.n94 8.85536
R357 VDD.n101 VDD.n100 8.85536
R358 VDD.n100 VDD.n99 8.85536
R359 VDD.n107 VDD.n104 8.85536
R360 VDD.n104 VDD.n103 8.85536
R361 VDD.n110 VDD.n109 8.85536
R362 VDD.n11 VDD.n8 8.4005
R363 VDD.n21 VDD.n18 7.6005
R364 VDD.n64 VDD.n61 7.2005
R365 VDD.n19 VDD.t50 5.23036
R366 VDD.n101 VDD.n98 4.8005
R367 VDD.n41 VDD.n38 4.8005
R368 VDD VDD.n110 4.6837
R369 VDD.n48 VDD.n47 4.6505
R370 VDD.n42 VDD.n41 4.6505
R371 VDD.n37 VDD.n36 4.6505
R372 VDD.n32 VDD.n31 4.6505
R373 VDD.n26 VDD.n25 4.6505
R374 VDD.n22 VDD.n21 4.6505
R375 VDD.n17 VDD.n16 4.6505
R376 VDD.n12 VDD.n11 4.6505
R377 VDD.n51 VDD.n50 4.6505
R378 VDD.n54 VDD.n53 4.6505
R379 VDD.n60 VDD.n59 4.6505
R380 VDD.n65 VDD.n64 4.6505
R381 VDD.n70 VDD.n69 4.6505
R382 VDD.n76 VDD.n75 4.6505
R383 VDD.n82 VDD.n81 4.6505
R384 VDD.n86 VDD.n85 4.6505
R385 VDD.n92 VDD.n91 4.6505
R386 VDD.n97 VDD.n96 4.6505
R387 VDD.n102 VDD.n101 4.6505
R388 VDD.n108 VDD.n107 4.6505
R389 VDD.n96 VDD.n93 4.0005
R390 VDD.n36 VDD.n33 4.0005
R391 VDD.n6 VDD.n2 3.66998
R392 VDD.n6 VDD.n5 3.46621
R393 VDD.n0 VDD.t38 1.74412
R394 VDD.n69 VDD.n66 1.6005
R395 VDD.n16 VDD.n13 1.2005
R396 VDD.n12 VDD.n6 0.915
R397 VDD.n51 VDD.n48 0.305188
R398 VDD.n48 VDD.n42 0.305188
R399 VDD.n42 VDD.n37 0.305188
R400 VDD.n37 VDD.n32 0.305188
R401 VDD.n32 VDD.n26 0.305188
R402 VDD.n26 VDD.n22 0.305188
R403 VDD.n22 VDD.n17 0.305188
R404 VDD.n17 VDD.n12 0.305188
R405 VDD.n60 VDD.n54 0.305188
R406 VDD.n65 VDD.n60 0.305188
R407 VDD.n70 VDD.n65 0.305188
R408 VDD.n76 VDD.n70 0.305188
R409 VDD.n82 VDD.n76 0.305188
R410 VDD.n86 VDD.n82 0.305188
R411 VDD.n92 VDD.n86 0.305188
R412 VDD.n97 VDD.n92 0.305188
R413 VDD.n102 VDD.n97 0.305188
R414 VDD.n108 VDD.n102 0.305188
R415 VDD VDD.n108 0.271984
R416 ready.n0 ready.t1 41.5677
R417 ready ready.t0 34.2053
R418 ready.n1 ready.n0 1.04094
R419 ready.n0 ready 0.804848
R420 ready ready.n1 0.0482941
R421 ready.n1 ready 0.0358261
R422 comp_outn.n0 comp_outn.t5 43.1877
R423 comp_outn.n1 comp_outn.t3 43.044
R424 comp_outn.n1 comp_outn.t4 43.044
R425 comp_outn comp_outn.t2 38.7789
R426 comp_outn.n4 comp_outn.t0 38.6969
R427 comp_outn.n4 comp_outn.t1 38.6969
R428 comp_outn.n2 comp_outn 1.15859
R429 comp_outn comp_outn.n4 0.984675
R430 comp_outn.n0 comp_outn 0.932565
R431 comp_outn.n5 comp_outn.n3 0.596088
R432 comp_outn.n5 comp_outn 0.438
R433 comp_outn.n2 comp_outn.n1 0.247153
R434 comp_outn comp_outn.n6 0.206382
R435 comp_outn.n3 comp_outn 0.15592
R436 comp_outn.n6 comp_outn 0.152674
R437 comp_outn.n6 comp_outn.n5 0.107118
R438 comp_outn.n2 comp_outn.n0 0.103441
R439 comp_outn.n5 comp_outn 0.063
R440 comp_outn.n3 comp_outn.n2 0.0193053
R441 comp_outp.n1 comp_outp.t5 43.1877
R442 comp_outp.n0 comp_outp.t3 43.044
R443 comp_outp.n0 comp_outp.t4 43.044
R444 comp_outp comp_outp.t2 38.7789
R445 comp_outp.n4 comp_outp.t0 38.6969
R446 comp_outp.n4 comp_outp.t1 38.6969
R447 comp_outp.n2 comp_outp 1.15859
R448 comp_outp.n5 comp_outp.n4 1.04718
R449 comp_outp.n1 comp_outp 0.932565
R450 comp_outp.n5 comp_outp.n3 0.596088
R451 comp_outp.n5 comp_outp 0.438
R452 comp_outp.n2 comp_outp.n0 0.247153
R453 comp_outp comp_outp.n6 0.206382
R454 comp_outp.n3 comp_outp 0.15592
R455 comp_outp.n6 comp_outp 0.152674
R456 comp_outp.n6 comp_outp.n5 0.107118
R457 comp_outp.n2 comp_outp.n1 0.103441
R458 comp_outp.n5 comp_outp 0.063
R459 comp_outp.n3 comp_outp.n2 0.0193053
R460 clk.n6 clk.t4 356.68
R461 clk.n5 clk.t5 356.68
R462 clk.n1 clk.t1 269.921
R463 clk.n0 clk.t0 269.921
R464 clk.n6 clk.t2 202.44
R465 clk.n5 clk.t7 202.44
R466 clk.n1 clk.t6 195.721
R467 clk.n0 clk.t3 195.721
R468 clk.n7 clk.n6 41.3896
R469 clk.n7 clk.n5 41.3896
R470 clk.n2 clk.n0 38.0628
R471 clk.n2 clk.n1 38.0536
R472 clk.n8 clk.n7 11.7969
R473 clk.n9 clk.n2 4.144
R474 clk.n10 clk.n9 1.12115
R475 clk.n11 clk.n10 0.0415156
R476 clk.n8 clk.n4 0.0415156
R477 clk.n9 clk.n8 0.012434
R478 clk clk.n11 0.0102656
R479 clk.n4 clk.n3 0.0083125
R480 cdac_vp.n0 cdac_vp.t6 340.613
R481 cdac_vp.n6 cdac_vp.t0 186.374
R482 cdac_vp.n5 cdac_vp.t7 186.374
R483 cdac_vp.n4 cdac_vp.t3 186.374
R484 cdac_vp.n3 cdac_vp.t1 186.374
R485 cdac_vp.n2 cdac_vp.t5 186.374
R486 cdac_vp.n1 cdac_vp.t4 186.374
R487 cdac_vp.n0 cdac_vp.t2 186.374
R488 cdac_vp.n1 cdac_vp.n0 154.24
R489 cdac_vp.n2 cdac_vp.n1 154.24
R490 cdac_vp.n3 cdac_vp.n2 154.24
R491 cdac_vp.n4 cdac_vp.n3 154.24
R492 cdac_vp.n5 cdac_vp.n4 154.24
R493 cdac_vp.n6 cdac_vp.n5 154.24
R494 cdac_vp cdac_vp.n6 102.168
C0 a_1026_n1747# a_476_n1721# 0.0123f
C1 Q cdac_vp 7.66e-20
C2 VDD a_582_n702# 0.0559f
C3 a_852_n296# VDD 0.755f
C4 comp_outn cdac_vn 3.55e-19
C5 a_1950_n1721# a_1026_n1747# 1.46e-19
C6 a_482_n1818# a_1716_n1348# 0.197f
C7 clk a_476_n1721# 0.0394f
C8 ready a_476_n1721# 0.0265f
C9 RS_n a_476_n1721# 0.00497f
C10 RS_n a_1950_n1721# 0.148f
C11 a_564_n1721# cdac_vp 0.00237f
C12 a_582_n702# a_482_n1818# 0.0247f
C13 a_852_n296# a_482_n1818# 0.0421f
C14 a_674_n702# a_1026_n1747# 3.37e-19
C15 clk a_1566_n378# 0.45f
C16 RS_n a_1566_n378# 1.34e-19
C17 VDD cdac_vn 0.0492f
C18 a_1950_n1721# a_476_n1721# 0.00449f
C19 a_564_n1266# cdac_vp 2.39e-20
C20 clk a_674_n702# 0.0918f
C21 a_564_n1721# a_564_n1266# 0.161f
C22 a_1566_n378# a_476_n1721# 0.119f
C23 a_1248_n288# VDD 0.814f
C24 RS_p a_564_n1721# 0.00308f
C25 a_482_n1818# cdac_vn 0.00294f
C26 a_1716_n1348# a_1026_n1747# 2.23e-21
C27 a_674_n702# a_476_n1721# 0.0934f
C28 VDD comp_outp 0.563f
C29 a_1248_n288# a_482_n1818# 0.0534f
C30 a_582_n702# a_1026_n1747# 6e-19
C31 clk a_1716_n1348# 0.0172f
C32 RS_n a_1716_n1348# 0.138f
C33 a_852_n296# a_1026_n1747# 0.015f
C34 a_674_n702# a_1566_n378# 0.194f
C35 clk a_582_n702# 0.0964f
C36 a_482_n1818# comp_outp 6.02e-19
C37 RS_n a_582_n702# 1.86e-19
C38 a_852_n296# ready 3.31e-19
C39 a_852_n296# clk 0.0178f
C40 a_852_n296# RS_n 0.025f
C41 a_1716_n1348# a_476_n1721# 0.067f
C42 a_1716_n1348# a_1950_n1721# 0.0147f
C43 a_582_n702# a_476_n1721# 0.0955f
C44 a_852_n296# a_476_n1721# 0.314f
C45 a_564_n1721# comp_outn 8.24e-22
C46 a_1716_n1348# a_1566_n378# 0.136f
C47 a_582_n702# a_1950_n1721# 5.99e-19
C48 VDD Q 0.366f
C49 clk cdac_vn 0.00752f
C50 a_582_n702# a_1566_n378# 0.00935f
C51 a_674_n702# a_1716_n1348# 0.00133f
C52 a_852_n296# a_1566_n378# 0.0115f
C53 RS_p comp_outn 8.63e-21
C54 a_1248_n288# clk 0.575f
C55 VDD cdac_vp 0.0153f
C56 comp_outp a_1026_n1747# 0.116f
C57 a_582_n702# a_674_n702# 1.53f
C58 a_482_n1818# Q 0.0238f
C59 VDD a_564_n1721# 0.165f
C60 a_852_n296# a_674_n702# 0.142f
C61 cdac_vn a_476_n1721# 0.0116f
C62 comp_outp ready 0.261f
C63 RS_n comp_outp 1.57e-19
C64 a_1950_n1721# cdac_vn 0.00709f
C65 a_1248_n288# a_476_n1721# 0.114f
C66 a_482_n1818# cdac_vp 0.016f
C67 VDD a_564_n1266# 2.11e-19
C68 a_564_n1721# a_482_n1818# 0.209f
C69 a_1566_n378# cdac_vn 0.00729f
C70 VDD RS_p 0.556f
C71 a_582_n702# a_1716_n1348# 0.0741f
C72 comp_outp a_476_n1721# 0.00983f
C73 a_852_n296# a_1716_n1348# 0.218f
C74 a_1248_n288# a_1566_n378# 0.406f
C75 a_674_n702# cdac_vn 7.65e-20
C76 a_564_n1266# a_482_n1818# 0.0165f
C77 a_852_n296# a_582_n702# 0.0742f
C78 RS_p a_482_n1818# 8.41e-20
C79 a_1248_n288# a_674_n702# 0.133f
C80 clk Q 0.0916f
C81 RS_n Q 7.8e-20
C82 a_1716_n1348# cdac_vn 0.0363f
C83 a_1026_n1747# cdac_vp 0.00723f
C84 a_564_n1721# a_1026_n1747# 0.0216f
C85 a_1248_n288# a_1716_n1348# 0.00935f
C86 a_582_n702# cdac_vn 0.129f
C87 a_852_n296# cdac_vn 0.00105f
C88 ready cdac_vp 2.7e-19
C89 Q a_476_n1721# 0.0281f
C90 clk cdac_vp 0.00752f
C91 VDD comp_outn 0.578f
C92 a_564_n1721# ready 0.068f
C93 RS_n a_564_n1721# 3.53e-20
C94 a_1248_n288# a_582_n702# 0.00778f
C95 a_564_n1266# a_1026_n1747# 1.65e-20
C96 Q a_1950_n1721# 3.37e-19
C97 a_852_n296# a_1248_n288# 0.135f
C98 RS_p a_1026_n1747# 0.149f
C99 Q a_1566_n378# 0.156f
C100 cdac_vp a_476_n1721# 0.0581f
C101 a_482_n1818# comp_outn 1.01e-21
C102 a_564_n1721# a_476_n1721# 0.388f
C103 a_852_n296# comp_outp 0.00587f
C104 clk RS_p 0.00119f
C105 RS_p ready 9.49e-21
C106 RS_n RS_p 0.314f
C107 Q a_674_n702# 0.00486f
C108 a_564_n1721# a_1950_n1721# 3.46e-21
C109 a_1566_n378# cdac_vp 1.93e-20
C110 a_564_n1266# a_476_n1721# 0.0219f
C111 a_1248_n288# cdac_vn 1.93e-20
C112 RS_p a_476_n1721# 0.00555f
C113 a_674_n702# cdac_vp 0.126f
C114 VDD a_482_n1818# 1.11f
C115 RS_p a_1950_n1721# 1.26e-19
C116 Q a_1716_n1348# 0.141f
C117 RS_p a_1566_n378# 4.77e-20
C118 a_582_n702# Q 1.53f
C119 a_852_n296# Q 0.00133f
C120 RS_p a_674_n702# 1e-19
C121 a_1716_n1348# cdac_vp 0.00105f
C122 a_564_n1721# a_1716_n1348# 1.33e-20
C123 RS_n comp_outn 1.85e-19
C124 a_582_n702# cdac_vp 0.129f
C125 a_852_n296# cdac_vp 0.0363f
C126 a_564_n1721# a_582_n702# 3.35e-19
C127 a_852_n296# a_564_n1721# 0.00163f
C128 VDD a_1026_n1747# 0.734f
C129 comp_outn a_476_n1721# 0.00199f
C130 RS_p a_1716_n1348# 0.0811f
C131 Q cdac_vn 0.126f
C132 comp_outn a_1950_n1721# 0.116f
C133 VDD ready 0.198f
C134 clk VDD 0.53f
C135 VDD RS_n 0.61f
C136 a_852_n296# a_564_n1266# 2.36e-21
C137 RS_p a_582_n702# 2.32e-19
C138 a_1248_n288# Q 0.195f
C139 a_482_n1818# a_1026_n1747# 4.38e-19
C140 a_852_n296# RS_p 0.166f
C141 VDD a_476_n1721# 0.811f
C142 a_482_n1818# ready 5.82e-20
C143 clk a_482_n1818# 0.113f
C144 RS_n a_482_n1818# 6.34e-20
C145 a_1248_n288# cdac_vp 0.00652f
C146 VDD a_1950_n1721# 0.743f
C147 VDD a_1566_n378# 0.767f
C148 comp_outp cdac_vp 3.55e-19
C149 a_482_n1818# a_476_n1721# 1.73f
C150 a_564_n1721# comp_outp 0.00514f
C151 a_1716_n1348# comp_outn 0.0058f
C152 a_482_n1818# a_1950_n1721# 2.63e-20
C153 VDD a_674_n702# 0.355f
C154 a_1248_n288# RS_p 2.46e-19
C155 a_482_n1818# a_1566_n378# 0.0258f
C156 RS_p comp_outp 1.16e-19
C157 ready a_1026_n1747# 0.00146f
C158 RS_n a_1026_n1747# 7.23e-19
C159 a_482_n1818# a_674_n702# 0.0145f
C160 VDD a_1716_n1348# 0.827f
C161 RS_n ready 2.19e-20
C162 clk RS_n 0.00115f
.ends

