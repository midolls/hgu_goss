magic
tech sky130A
timestamp 1698229845
<< nwell >>
rect -21 763 8335 930
<< metal1 >>
rect -299 1216 8722 1264
rect -299 944 8722 992
rect -299 882 8722 930
rect -299 610 8722 658
rect -299 548 883 596
rect -299 276 8722 324
rect -299 214 8722 262
rect -299 -58 8722 -10
use sky130_fd_sc_hd__buf_1  x1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1697295826
transform 1 0 0 0 1 968
box -19 -24 157 296
use sky130_fd_sc_hd__buf_16  x2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 414 0 1 968
box -19 -24 1031 296
use sky130_fd_sc_hd__buf_4  x3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1697295826
transform 1 0 138 0 1 968
box -19 -24 295 296
use sky130_fd_sc_hd__dfbbn_1  x4 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 0 0 1 300
box -19 -24 1215 296
use sky130_fd_sc_hd__dfbbn_1  x5
timestamp 1683767628
transform -1 0 1196 0 1 -34
box -19 -24 1215 296
use sky130_fd_sc_hd__mux2_1  x6 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 0 0 1 634
box -19 -24 433 296
use sky130_fd_sc_hd__mux2_1  x7
timestamp 1683767628
transform -1 0 1138 0 1 634
box -19 -24 433 296
use sky130_fd_sc_hd__mux2_1  x8
timestamp 1683767628
transform 1 0 1196 0 1 634
box -19 -24 433 296
use sky130_fd_sc_hd__mux2_1  x9
timestamp 1683767628
transform -1 0 2334 0 1 634
box -19 -24 433 296
use sky130_fd_sc_hd__mux2_1  x10
timestamp 1683767628
transform 1 0 2392 0 1 634
box -19 -24 433 296
use sky130_fd_sc_hd__mux2_1  x11
timestamp 1683767628
transform -1 0 3529 0 1 634
box -19 -24 433 296
use sky130_fd_sc_hd__mux2_1  x12
timestamp 1683767628
transform 1 0 3588 0 1 634
box -19 -24 433 296
use sky130_fd_sc_hd__mux2_1  x13
timestamp 1683767628
transform -1 0 4726 0 1 634
box -19 -24 433 296
use sky130_fd_sc_hd__mux2_1  x14
timestamp 1683767628
transform 1 0 4784 0 1 634
box -19 -24 433 296
use sky130_fd_sc_hd__mux2_1  x15
timestamp 1683767628
transform -1 0 5922 0 1 634
box -19 -24 433 296
use sky130_fd_sc_hd__mux2_1  x16
timestamp 1683767628
transform 1 0 5980 0 1 634
box -19 -24 433 296
use sky130_fd_sc_hd__mux2_1  x17
timestamp 1683767628
transform -1 0 7117 0 1 634
box -19 -24 433 296
use sky130_fd_sc_hd__mux2_1  x18
timestamp 1683767628
transform 1 0 7176 0 1 634
box -19 -24 433 296
use sky130_fd_sc_hd__dfbbn_1  x19
timestamp 1683767628
transform 1 0 1196 0 1 300
box -19 -24 1215 296
use sky130_fd_sc_hd__mux2_1  x20
timestamp 1683767628
transform -1 0 8314 0 1 634
box -19 -24 433 296
use sky130_fd_sc_hd__dfbbn_1  x21
timestamp 1683767628
transform -1 0 2392 0 1 -34
box -19 -24 1215 296
use sky130_fd_sc_hd__dfbbn_1  x23
timestamp 1683767628
transform 1 0 2392 0 1 300
box -19 -24 1215 296
use sky130_fd_sc_hd__dfbbn_1  x24
timestamp 1683767628
transform -1 0 3588 0 1 -34
box -19 -24 1215 296
use sky130_fd_sc_hd__dfbbn_1  x25
timestamp 1683767628
transform 1 0 3588 0 1 300
box -19 -24 1215 296
use sky130_fd_sc_hd__dfbbn_1  x26
timestamp 1683767628
transform -1 0 4784 0 1 -34
box -19 -24 1215 296
use sky130_fd_sc_hd__dfbbn_1  x28
timestamp 1683767628
transform 1 0 4784 0 1 300
box -19 -24 1215 296
use sky130_fd_sc_hd__dfbbn_1  x29
timestamp 1683767628
transform -1 0 5980 0 1 -34
box -19 -24 1215 296
use sky130_fd_sc_hd__dfbbn_1  x31
timestamp 1683767628
transform 1 0 5980 0 1 300
box -19 -24 1215 296
use sky130_fd_sc_hd__dfbbn_1  x32
timestamp 1683767628
transform -1 0 7176 0 1 -34
box -19 -24 1215 296
use sky130_fd_sc_hd__dfbbn_1  x34
timestamp 1683767628
transform 1 0 7176 0 1 300
box -19 -24 1215 296
use sky130_fd_sc_hd__dfbbn_1  x35
timestamp 1683767628
transform -1 0 8372 0 1 -34
box -19 -24 1215 296
<< end >>
