magic
tech sky130A
magscale 1 2
timestamp 1697888221
<< nwell >>
rect 652 -78 2714 528
rect 1252 -110 2114 -78
rect 338 -1940 2546 -1334
<< nmos >>
rect 852 -270 882 -178
rect 948 -270 978 -178
rect 1044 -270 1074 -178
rect 1248 -262 1278 -178
rect 1536 -378 1566 -178
rect 1800 -378 1830 -178
rect 2088 -262 2118 -178
rect 2292 -270 2322 -178
rect 2388 -270 2418 -178
rect 2484 -270 2514 -178
rect 1524 -702 1554 -502
rect 1620 -702 1650 -502
rect 1716 -702 1746 -502
rect 1812 -702 1842 -502
rect 534 -1266 564 -1098
rect 622 -1266 652 -1098
rect 822 -1266 852 -1182
rect 1026 -1266 1056 -1174
rect 1122 -1266 1152 -1174
rect 1218 -1266 1248 -1174
rect 1422 -1266 1452 -1182
rect 1628 -1260 1658 -1092
rect 1716 -1260 1746 -1092
rect 1920 -1266 1950 -1182
rect 2124 -1266 2154 -1174
rect 2220 -1266 2250 -1174
rect 2316 -1266 2346 -1174
<< pmos >>
rect 852 141 882 309
rect 948 141 978 309
rect 1044 141 1074 309
rect 1248 141 1278 309
rect 1448 109 1478 309
rect 1536 109 1566 309
rect 1624 109 1654 309
rect 1712 109 1742 309
rect 1800 109 1830 309
rect 1888 109 1918 309
rect 2088 141 2118 309
rect 2292 141 2322 309
rect 2388 141 2418 309
rect 2484 141 2514 309
rect 534 -1721 564 -1553
rect 622 -1721 652 -1553
rect 822 -1721 852 -1553
rect 1026 -1721 1056 -1553
rect 1122 -1721 1152 -1553
rect 1218 -1721 1248 -1553
rect 1422 -1721 1452 -1553
rect 1628 -1721 1658 -1553
rect 1716 -1721 1746 -1553
rect 1920 -1721 1950 -1553
rect 2124 -1721 2154 -1553
rect 2220 -1721 2250 -1553
rect 2316 -1721 2346 -1553
<< nmoslvt >>
rect 644 -702 674 -502
rect 740 -702 770 -502
rect 836 -702 866 -502
rect 932 -702 962 -502
rect 1028 -702 1058 -502
rect 1124 -702 1154 -502
rect 1220 -702 1250 -502
rect 1316 -702 1346 -502
rect 2020 -702 2050 -502
rect 2116 -702 2146 -502
rect 2212 -702 2242 -502
rect 2308 -702 2338 -502
rect 2404 -702 2434 -502
rect 2500 -702 2530 -502
rect 2596 -702 2626 -502
rect 2692 -702 2722 -502
<< ndiff >>
rect 790 -190 852 -178
rect 790 -258 802 -190
rect 836 -258 852 -190
rect 790 -270 852 -258
rect 882 -190 948 -178
rect 882 -258 898 -190
rect 932 -258 948 -190
rect 882 -270 948 -258
rect 978 -190 1044 -178
rect 978 -258 994 -190
rect 1028 -258 1044 -190
rect 978 -270 1044 -258
rect 1074 -190 1136 -178
rect 1074 -258 1090 -190
rect 1124 -258 1136 -190
rect 1074 -270 1136 -258
rect 1190 -190 1248 -178
rect 1190 -250 1202 -190
rect 1236 -250 1248 -190
rect 1190 -262 1248 -250
rect 1278 -190 1336 -178
rect 1278 -250 1290 -190
rect 1324 -250 1336 -190
rect 1278 -262 1336 -250
rect 1478 -190 1536 -178
rect 1478 -366 1490 -190
rect 1524 -366 1536 -190
rect 1478 -378 1536 -366
rect 1566 -190 1624 -178
rect 1566 -366 1578 -190
rect 1612 -366 1624 -190
rect 1566 -378 1624 -366
rect 1742 -190 1800 -178
rect 1742 -366 1754 -190
rect 1788 -366 1800 -190
rect 1742 -378 1800 -366
rect 1830 -190 1888 -178
rect 1830 -366 1842 -190
rect 1876 -366 1888 -190
rect 1830 -378 1888 -366
rect 2030 -190 2088 -178
rect 2030 -250 2042 -190
rect 2076 -250 2088 -190
rect 2030 -262 2088 -250
rect 2118 -190 2176 -178
rect 2118 -250 2130 -190
rect 2164 -250 2176 -190
rect 2118 -262 2176 -250
rect 2230 -190 2292 -178
rect 2230 -258 2242 -190
rect 2276 -258 2292 -190
rect 2230 -270 2292 -258
rect 2322 -190 2388 -178
rect 2322 -258 2338 -190
rect 2372 -258 2388 -190
rect 2322 -270 2388 -258
rect 2418 -190 2484 -178
rect 2418 -258 2434 -190
rect 2468 -258 2484 -190
rect 2418 -270 2484 -258
rect 2514 -190 2576 -178
rect 2514 -258 2530 -190
rect 2564 -258 2576 -190
rect 2514 -270 2576 -258
rect 582 -514 644 -502
rect 582 -690 594 -514
rect 628 -690 644 -514
rect 582 -702 644 -690
rect 674 -514 740 -502
rect 674 -690 690 -514
rect 724 -690 740 -514
rect 674 -702 740 -690
rect 770 -514 836 -502
rect 770 -690 786 -514
rect 820 -690 836 -514
rect 770 -702 836 -690
rect 866 -514 932 -502
rect 866 -690 882 -514
rect 916 -690 932 -514
rect 866 -702 932 -690
rect 962 -514 1028 -502
rect 962 -690 978 -514
rect 1012 -690 1028 -514
rect 962 -702 1028 -690
rect 1058 -514 1124 -502
rect 1058 -690 1074 -514
rect 1108 -690 1124 -514
rect 1058 -702 1124 -690
rect 1154 -514 1220 -502
rect 1154 -690 1170 -514
rect 1204 -690 1220 -514
rect 1154 -702 1220 -690
rect 1250 -514 1316 -502
rect 1250 -690 1266 -514
rect 1300 -690 1316 -514
rect 1250 -702 1316 -690
rect 1346 -514 1408 -502
rect 1346 -690 1362 -514
rect 1396 -690 1408 -514
rect 1346 -702 1408 -690
rect 1462 -514 1524 -502
rect 1462 -690 1474 -514
rect 1508 -690 1524 -514
rect 1462 -702 1524 -690
rect 1554 -514 1620 -502
rect 1554 -690 1570 -514
rect 1604 -690 1620 -514
rect 1554 -702 1620 -690
rect 1650 -514 1716 -502
rect 1650 -690 1666 -514
rect 1700 -690 1716 -514
rect 1650 -702 1716 -690
rect 1746 -514 1812 -502
rect 1746 -690 1762 -514
rect 1796 -690 1812 -514
rect 1746 -702 1812 -690
rect 1842 -514 1904 -502
rect 1842 -690 1858 -514
rect 1892 -690 1904 -514
rect 1842 -702 1904 -690
rect 1958 -514 2020 -502
rect 1958 -690 1970 -514
rect 2004 -690 2020 -514
rect 1958 -702 2020 -690
rect 2050 -514 2116 -502
rect 2050 -690 2066 -514
rect 2100 -690 2116 -514
rect 2050 -702 2116 -690
rect 2146 -514 2212 -502
rect 2146 -690 2162 -514
rect 2196 -690 2212 -514
rect 2146 -702 2212 -690
rect 2242 -514 2308 -502
rect 2242 -690 2258 -514
rect 2292 -690 2308 -514
rect 2242 -702 2308 -690
rect 2338 -514 2404 -502
rect 2338 -690 2354 -514
rect 2388 -690 2404 -514
rect 2338 -702 2404 -690
rect 2434 -514 2500 -502
rect 2434 -690 2450 -514
rect 2484 -690 2500 -514
rect 2434 -702 2500 -690
rect 2530 -514 2596 -502
rect 2530 -690 2546 -514
rect 2580 -690 2596 -514
rect 2530 -702 2596 -690
rect 2626 -514 2692 -502
rect 2626 -690 2642 -514
rect 2676 -690 2692 -514
rect 2626 -702 2692 -690
rect 2722 -514 2784 -502
rect 2722 -690 2738 -514
rect 2772 -690 2784 -514
rect 2722 -702 2784 -690
rect 476 -1110 534 -1098
rect 476 -1254 488 -1110
rect 522 -1254 534 -1110
rect 476 -1266 534 -1254
rect 564 -1110 622 -1098
rect 564 -1254 576 -1110
rect 610 -1254 622 -1110
rect 564 -1266 622 -1254
rect 652 -1110 710 -1098
rect 652 -1254 664 -1110
rect 698 -1254 710 -1110
rect 1570 -1104 1628 -1092
rect 652 -1266 710 -1254
rect 764 -1194 822 -1182
rect 764 -1254 776 -1194
rect 810 -1254 822 -1194
rect 764 -1266 822 -1254
rect 852 -1194 910 -1182
rect 852 -1254 864 -1194
rect 898 -1254 910 -1194
rect 852 -1266 910 -1254
rect 964 -1186 1026 -1174
rect 964 -1254 976 -1186
rect 1010 -1254 1026 -1186
rect 964 -1266 1026 -1254
rect 1056 -1186 1122 -1174
rect 1056 -1254 1072 -1186
rect 1106 -1254 1122 -1186
rect 1056 -1266 1122 -1254
rect 1152 -1186 1218 -1174
rect 1152 -1254 1168 -1186
rect 1202 -1254 1218 -1186
rect 1152 -1266 1218 -1254
rect 1248 -1186 1310 -1174
rect 1248 -1254 1264 -1186
rect 1298 -1254 1310 -1186
rect 1248 -1266 1310 -1254
rect 1364 -1194 1422 -1182
rect 1364 -1254 1376 -1194
rect 1410 -1254 1422 -1194
rect 1364 -1266 1422 -1254
rect 1452 -1194 1510 -1182
rect 1452 -1254 1464 -1194
rect 1498 -1254 1510 -1194
rect 1452 -1266 1510 -1254
rect 1570 -1248 1582 -1104
rect 1616 -1248 1628 -1104
rect 1570 -1260 1628 -1248
rect 1658 -1104 1716 -1092
rect 1658 -1248 1670 -1104
rect 1704 -1248 1716 -1104
rect 1658 -1260 1716 -1248
rect 1746 -1104 1804 -1092
rect 1746 -1248 1758 -1104
rect 1792 -1248 1804 -1104
rect 1746 -1260 1804 -1248
rect 1862 -1194 1920 -1182
rect 1862 -1254 1874 -1194
rect 1908 -1254 1920 -1194
rect 1862 -1266 1920 -1254
rect 1950 -1194 2008 -1182
rect 1950 -1254 1962 -1194
rect 1996 -1254 2008 -1194
rect 1950 -1266 2008 -1254
rect 2062 -1186 2124 -1174
rect 2062 -1254 2074 -1186
rect 2108 -1254 2124 -1186
rect 2062 -1266 2124 -1254
rect 2154 -1186 2220 -1174
rect 2154 -1254 2170 -1186
rect 2204 -1254 2220 -1186
rect 2154 -1266 2220 -1254
rect 2250 -1186 2316 -1174
rect 2250 -1254 2266 -1186
rect 2300 -1254 2316 -1186
rect 2250 -1266 2316 -1254
rect 2346 -1186 2408 -1174
rect 2346 -1254 2362 -1186
rect 2396 -1254 2408 -1186
rect 2346 -1266 2408 -1254
<< pdiff >>
rect 790 297 852 309
rect 790 153 802 297
rect 836 153 852 297
rect 790 141 852 153
rect 882 297 948 309
rect 882 153 898 297
rect 932 153 948 297
rect 882 141 948 153
rect 978 297 1044 309
rect 978 153 994 297
rect 1028 153 1044 297
rect 978 141 1044 153
rect 1074 297 1136 309
rect 1074 153 1090 297
rect 1124 153 1136 297
rect 1074 141 1136 153
rect 1190 297 1248 309
rect 1190 153 1202 297
rect 1236 153 1248 297
rect 1190 141 1248 153
rect 1278 297 1336 309
rect 1278 153 1290 297
rect 1324 153 1336 297
rect 1278 141 1336 153
rect 1390 297 1448 309
rect 1390 121 1402 297
rect 1436 121 1448 297
rect 1390 109 1448 121
rect 1478 297 1536 309
rect 1478 121 1490 297
rect 1524 121 1536 297
rect 1478 109 1536 121
rect 1566 297 1624 309
rect 1566 121 1578 297
rect 1612 121 1624 297
rect 1566 109 1624 121
rect 1654 297 1712 309
rect 1654 121 1666 297
rect 1700 121 1712 297
rect 1654 109 1712 121
rect 1742 297 1800 309
rect 1742 121 1754 297
rect 1788 121 1800 297
rect 1742 109 1800 121
rect 1830 297 1888 309
rect 1830 121 1842 297
rect 1876 121 1888 297
rect 1830 109 1888 121
rect 1918 297 1976 309
rect 1918 121 1930 297
rect 1964 121 1976 297
rect 2030 297 2088 309
rect 2030 153 2042 297
rect 2076 153 2088 297
rect 2030 141 2088 153
rect 2118 297 2176 309
rect 2118 153 2130 297
rect 2164 153 2176 297
rect 2118 141 2176 153
rect 2230 297 2292 309
rect 2230 153 2242 297
rect 2276 153 2292 297
rect 2230 141 2292 153
rect 2322 297 2388 309
rect 2322 153 2338 297
rect 2372 153 2388 297
rect 2322 141 2388 153
rect 2418 297 2484 309
rect 2418 153 2434 297
rect 2468 153 2484 297
rect 2418 141 2484 153
rect 2514 297 2576 309
rect 2514 153 2530 297
rect 2564 153 2576 297
rect 2514 141 2576 153
rect 1918 109 1976 121
rect 476 -1565 534 -1553
rect 476 -1709 488 -1565
rect 522 -1709 534 -1565
rect 476 -1721 534 -1709
rect 564 -1565 622 -1553
rect 564 -1709 576 -1565
rect 610 -1709 622 -1565
rect 564 -1721 622 -1709
rect 652 -1565 710 -1553
rect 652 -1709 664 -1565
rect 698 -1709 710 -1565
rect 652 -1721 710 -1709
rect 764 -1565 822 -1553
rect 764 -1709 776 -1565
rect 810 -1709 822 -1565
rect 764 -1721 822 -1709
rect 852 -1565 910 -1553
rect 852 -1709 864 -1565
rect 898 -1709 910 -1565
rect 852 -1721 910 -1709
rect 964 -1565 1026 -1553
rect 964 -1709 976 -1565
rect 1010 -1709 1026 -1565
rect 964 -1721 1026 -1709
rect 1056 -1565 1122 -1553
rect 1056 -1709 1072 -1565
rect 1106 -1709 1122 -1565
rect 1056 -1721 1122 -1709
rect 1152 -1565 1218 -1553
rect 1152 -1709 1168 -1565
rect 1202 -1709 1218 -1565
rect 1152 -1721 1218 -1709
rect 1248 -1565 1310 -1553
rect 1248 -1709 1264 -1565
rect 1298 -1709 1310 -1565
rect 1248 -1721 1310 -1709
rect 1364 -1565 1422 -1553
rect 1364 -1709 1376 -1565
rect 1410 -1709 1422 -1565
rect 1364 -1721 1422 -1709
rect 1452 -1565 1510 -1553
rect 1452 -1709 1464 -1565
rect 1498 -1709 1510 -1565
rect 1452 -1721 1510 -1709
rect 1570 -1565 1628 -1553
rect 1570 -1709 1582 -1565
rect 1616 -1709 1628 -1565
rect 1570 -1721 1628 -1709
rect 1658 -1565 1716 -1553
rect 1658 -1709 1670 -1565
rect 1704 -1709 1716 -1565
rect 1658 -1721 1716 -1709
rect 1746 -1565 1804 -1553
rect 1746 -1709 1758 -1565
rect 1792 -1709 1804 -1565
rect 1746 -1721 1804 -1709
rect 1862 -1565 1920 -1553
rect 1862 -1709 1874 -1565
rect 1908 -1709 1920 -1565
rect 1862 -1721 1920 -1709
rect 1950 -1565 2008 -1553
rect 1950 -1709 1962 -1565
rect 1996 -1709 2008 -1565
rect 1950 -1721 2008 -1709
rect 2062 -1565 2124 -1553
rect 2062 -1709 2074 -1565
rect 2108 -1709 2124 -1565
rect 2062 -1721 2124 -1709
rect 2154 -1565 2220 -1553
rect 2154 -1709 2170 -1565
rect 2204 -1709 2220 -1565
rect 2154 -1721 2220 -1709
rect 2250 -1565 2316 -1553
rect 2250 -1709 2266 -1565
rect 2300 -1709 2316 -1565
rect 2250 -1721 2316 -1709
rect 2346 -1565 2408 -1553
rect 2346 -1709 2362 -1565
rect 2396 -1709 2408 -1565
rect 2346 -1721 2408 -1709
<< ndiffc >>
rect 802 -258 836 -190
rect 898 -258 932 -190
rect 994 -258 1028 -190
rect 1090 -258 1124 -190
rect 1202 -250 1236 -190
rect 1290 -250 1324 -190
rect 1490 -366 1524 -190
rect 1578 -366 1612 -190
rect 1754 -366 1788 -190
rect 1842 -366 1876 -190
rect 2042 -250 2076 -190
rect 2130 -250 2164 -190
rect 2242 -258 2276 -190
rect 2338 -258 2372 -190
rect 2434 -258 2468 -190
rect 2530 -258 2564 -190
rect 594 -690 628 -514
rect 690 -690 724 -514
rect 786 -690 820 -514
rect 882 -690 916 -514
rect 978 -690 1012 -514
rect 1074 -690 1108 -514
rect 1170 -690 1204 -514
rect 1266 -690 1300 -514
rect 1362 -690 1396 -514
rect 1474 -690 1508 -514
rect 1570 -690 1604 -514
rect 1666 -690 1700 -514
rect 1762 -690 1796 -514
rect 1858 -690 1892 -514
rect 1970 -690 2004 -514
rect 2066 -690 2100 -514
rect 2162 -690 2196 -514
rect 2258 -690 2292 -514
rect 2354 -690 2388 -514
rect 2450 -690 2484 -514
rect 2546 -690 2580 -514
rect 2642 -690 2676 -514
rect 2738 -690 2772 -514
rect 488 -1254 522 -1110
rect 576 -1254 610 -1110
rect 664 -1254 698 -1110
rect 776 -1254 810 -1194
rect 864 -1254 898 -1194
rect 976 -1254 1010 -1186
rect 1072 -1254 1106 -1186
rect 1168 -1254 1202 -1186
rect 1264 -1254 1298 -1186
rect 1376 -1254 1410 -1194
rect 1464 -1254 1498 -1194
rect 1582 -1248 1616 -1104
rect 1670 -1248 1704 -1104
rect 1758 -1248 1792 -1104
rect 1874 -1254 1908 -1194
rect 1962 -1254 1996 -1194
rect 2074 -1254 2108 -1186
rect 2170 -1254 2204 -1186
rect 2266 -1254 2300 -1186
rect 2362 -1254 2396 -1186
<< pdiffc >>
rect 802 153 836 297
rect 898 153 932 297
rect 994 153 1028 297
rect 1090 153 1124 297
rect 1202 153 1236 297
rect 1290 153 1324 297
rect 1402 121 1436 297
rect 1490 121 1524 297
rect 1578 121 1612 297
rect 1666 121 1700 297
rect 1754 121 1788 297
rect 1842 121 1876 297
rect 1930 121 1964 297
rect 2042 153 2076 297
rect 2130 153 2164 297
rect 2242 153 2276 297
rect 2338 153 2372 297
rect 2434 153 2468 297
rect 2530 153 2564 297
rect 488 -1709 522 -1565
rect 576 -1709 610 -1565
rect 664 -1709 698 -1565
rect 776 -1709 810 -1565
rect 864 -1709 898 -1565
rect 976 -1709 1010 -1565
rect 1072 -1709 1106 -1565
rect 1168 -1709 1202 -1565
rect 1264 -1709 1298 -1565
rect 1376 -1709 1410 -1565
rect 1464 -1709 1498 -1565
rect 1582 -1709 1616 -1565
rect 1670 -1709 1704 -1565
rect 1758 -1709 1792 -1565
rect 1874 -1709 1908 -1565
rect 1962 -1709 1996 -1565
rect 2074 -1709 2108 -1565
rect 2170 -1709 2204 -1565
rect 2266 -1709 2300 -1565
rect 2362 -1709 2396 -1565
<< psubdiff >>
rect 826 -336 1338 -324
rect 826 -370 868 -336
rect 902 -370 968 -336
rect 1002 -370 1068 -336
rect 1102 -370 1168 -336
rect 1202 -370 1268 -336
rect 1302 -370 1338 -336
rect 826 -382 1338 -370
rect 2028 -336 2540 -324
rect 2028 -370 2070 -336
rect 2104 -370 2170 -336
rect 2204 -370 2270 -336
rect 2304 -370 2370 -336
rect 2404 -370 2470 -336
rect 2504 -370 2540 -336
rect 2028 -382 2540 -370
rect 544 -816 2834 -792
rect 544 -850 568 -816
rect 602 -850 668 -816
rect 702 -850 768 -816
rect 802 -850 868 -816
rect 902 -850 968 -816
rect 1002 -850 1068 -816
rect 1102 -850 1168 -816
rect 1202 -850 1268 -816
rect 1302 -850 1368 -816
rect 1402 -850 1468 -816
rect 1502 -850 1568 -816
rect 1602 -850 1668 -816
rect 1702 -850 1768 -816
rect 1802 -850 1868 -816
rect 1902 -850 1968 -816
rect 2002 -850 2068 -816
rect 2102 -850 2168 -816
rect 2202 -850 2268 -816
rect 2302 -850 2368 -816
rect 2402 -850 2468 -816
rect 2502 -850 2568 -816
rect 2602 -850 2668 -816
rect 2702 -850 2768 -816
rect 2802 -850 2834 -816
rect 544 -976 2834 -850
rect 544 -1010 568 -976
rect 602 -1010 668 -976
rect 702 -980 2834 -976
rect 702 -1010 1568 -980
rect 544 -1014 1568 -1010
rect 1602 -1014 1668 -980
rect 1702 -1014 1768 -980
rect 1802 -1014 2834 -980
rect 544 -1034 2834 -1014
rect 764 -1038 2834 -1034
rect 764 -1062 1516 -1038
rect 764 -1096 770 -1062
rect 804 -1096 868 -1062
rect 902 -1096 968 -1062
rect 1002 -1096 1068 -1062
rect 1102 -1096 1168 -1062
rect 1202 -1096 1268 -1062
rect 1302 -1096 1368 -1062
rect 1402 -1096 1468 -1062
rect 1502 -1096 1516 -1062
rect 1860 -1062 2834 -1038
rect 764 -1120 1516 -1096
rect 1860 -1096 1868 -1062
rect 1902 -1096 1968 -1062
rect 2002 -1096 2068 -1062
rect 2102 -1096 2168 -1062
rect 2202 -1096 2268 -1062
rect 2302 -1096 2368 -1062
rect 2402 -1096 2468 -1062
rect 2502 -1096 2568 -1062
rect 2602 -1096 2668 -1062
rect 2702 -1096 2768 -1062
rect 2802 -1096 2834 -1062
rect 1860 -1120 2834 -1096
<< nsubdiff >>
rect 762 412 2624 428
rect 762 378 802 412
rect 836 378 958 412
rect 992 378 1114 412
rect 1148 378 1270 412
rect 1304 378 1426 412
rect 1460 378 1582 412
rect 1616 378 1738 412
rect 1772 378 1894 412
rect 1928 378 2050 412
rect 2084 378 2206 412
rect 2240 378 2362 412
rect 2396 378 2518 412
rect 2552 378 2624 412
rect 762 364 2624 378
rect 758 -1792 2440 -1776
rect 758 -1826 818 -1792
rect 852 -1826 958 -1792
rect 992 -1826 1114 -1792
rect 1148 -1826 1270 -1792
rect 1304 -1826 1426 -1792
rect 1460 -1826 1582 -1792
rect 1616 -1826 1738 -1792
rect 1772 -1826 1894 -1792
rect 1928 -1826 2050 -1792
rect 2084 -1826 2206 -1792
rect 2240 -1826 2362 -1792
rect 2396 -1826 2440 -1792
rect 758 -1840 2440 -1826
<< psubdiffcont >>
rect 868 -370 902 -336
rect 968 -370 1002 -336
rect 1068 -370 1102 -336
rect 1168 -370 1202 -336
rect 1268 -370 1302 -336
rect 2070 -370 2104 -336
rect 2170 -370 2204 -336
rect 2270 -370 2304 -336
rect 2370 -370 2404 -336
rect 2470 -370 2504 -336
rect 568 -850 602 -816
rect 668 -850 702 -816
rect 768 -850 802 -816
rect 868 -850 902 -816
rect 968 -850 1002 -816
rect 1068 -850 1102 -816
rect 1168 -850 1202 -816
rect 1268 -850 1302 -816
rect 1368 -850 1402 -816
rect 1468 -850 1502 -816
rect 1568 -850 1602 -816
rect 1668 -850 1702 -816
rect 1768 -850 1802 -816
rect 1868 -850 1902 -816
rect 1968 -850 2002 -816
rect 2068 -850 2102 -816
rect 2168 -850 2202 -816
rect 2268 -850 2302 -816
rect 2368 -850 2402 -816
rect 2468 -850 2502 -816
rect 2568 -850 2602 -816
rect 2668 -850 2702 -816
rect 2768 -850 2802 -816
rect 568 -1010 602 -976
rect 668 -1010 702 -976
rect 1568 -1014 1602 -980
rect 1668 -1014 1702 -980
rect 1768 -1014 1802 -980
rect 770 -1096 804 -1062
rect 868 -1096 902 -1062
rect 968 -1096 1002 -1062
rect 1068 -1096 1102 -1062
rect 1168 -1096 1202 -1062
rect 1268 -1096 1302 -1062
rect 1368 -1096 1402 -1062
rect 1468 -1096 1502 -1062
rect 1868 -1096 1902 -1062
rect 1968 -1096 2002 -1062
rect 2068 -1096 2102 -1062
rect 2168 -1096 2202 -1062
rect 2268 -1096 2302 -1062
rect 2368 -1096 2402 -1062
rect 2468 -1096 2502 -1062
rect 2568 -1096 2602 -1062
rect 2668 -1096 2702 -1062
rect 2768 -1096 2802 -1062
<< nsubdiffcont >>
rect 802 378 836 412
rect 958 378 992 412
rect 1114 378 1148 412
rect 1270 378 1304 412
rect 1426 378 1460 412
rect 1582 378 1616 412
rect 1738 378 1772 412
rect 1894 378 1928 412
rect 2050 378 2084 412
rect 2206 378 2240 412
rect 2362 378 2396 412
rect 2518 378 2552 412
rect 818 -1826 852 -1792
rect 958 -1826 992 -1792
rect 1114 -1826 1148 -1792
rect 1270 -1826 1304 -1792
rect 1426 -1826 1460 -1792
rect 1582 -1826 1616 -1792
rect 1738 -1826 1772 -1792
rect 1894 -1826 1928 -1792
rect 2050 -1826 2084 -1792
rect 2206 -1826 2240 -1792
rect 2362 -1826 2396 -1792
<< poly >>
rect 852 309 882 335
rect 948 309 978 340
rect 1044 309 1074 335
rect 1248 309 1278 340
rect 1448 309 1478 340
rect 1536 309 1566 340
rect 1624 309 1654 340
rect 1712 309 1742 340
rect 1800 309 1830 340
rect 1888 309 1918 340
rect 2088 309 2118 340
rect 2292 309 2322 335
rect 2388 309 2418 340
rect 2484 309 2514 335
rect 852 126 882 141
rect 948 126 978 141
rect 1044 126 1074 141
rect 852 96 1074 126
rect 1040 24 1074 96
rect 1040 8 1106 24
rect 1040 -26 1056 8
rect 1090 -26 1106 8
rect 1040 -42 1106 -26
rect 1248 -22 1278 141
rect 1448 94 1478 109
rect 1536 94 1566 109
rect 1416 64 1566 94
rect 1248 -38 1328 -22
rect 1040 -132 1074 -42
rect 852 -162 1074 -132
rect 852 -178 882 -162
rect 948 -178 978 -162
rect 1044 -178 1074 -162
rect 1248 -72 1278 -38
rect 1312 -72 1328 -38
rect 1248 -88 1328 -72
rect 1248 -178 1278 -88
rect 852 -296 882 -270
rect 948 -296 978 -270
rect 1044 -296 1074 -270
rect 1248 -288 1278 -262
rect 578 -430 674 -414
rect 578 -464 594 -430
rect 628 -456 674 -430
rect 1416 -446 1446 64
rect 1624 22 1654 109
rect 1536 -8 1654 22
rect 1712 22 1742 109
rect 1800 94 1830 109
rect 1888 94 1918 109
rect 1800 64 1950 94
rect 1712 -8 1830 22
rect 1536 -26 1566 -8
rect 1488 -38 1566 -26
rect 1488 -72 1504 -38
rect 1538 -72 1566 -38
rect 1488 -84 1566 -72
rect 1536 -178 1566 -84
rect 1800 -94 1830 -8
rect 1800 -106 1878 -94
rect 1800 -140 1828 -106
rect 1862 -140 1878 -106
rect 1800 -152 1878 -140
rect 1800 -178 1830 -152
rect 1536 -404 1566 -378
rect 1650 -398 1716 -384
rect 1650 -432 1666 -398
rect 1700 -432 1716 -398
rect 1800 -404 1830 -378
rect 1650 -446 1716 -432
rect 1920 -446 1950 64
rect 2088 -86 2118 141
rect 2292 126 2322 141
rect 2388 126 2418 141
rect 2484 126 2514 141
rect 2292 96 2514 126
rect 2292 24 2322 96
rect 2256 8 2322 24
rect 2256 -26 2272 8
rect 2306 -26 2322 8
rect 2256 -42 2322 -26
rect 2036 -102 2118 -86
rect 2036 -136 2052 -102
rect 2086 -136 2118 -102
rect 2036 -152 2118 -136
rect 2088 -178 2118 -152
rect 2292 -132 2322 -42
rect 2292 -162 2514 -132
rect 2292 -178 2322 -162
rect 2388 -178 2418 -162
rect 2484 -178 2514 -162
rect 2088 -288 2118 -262
rect 2292 -296 2322 -270
rect 2388 -296 2418 -270
rect 2484 -296 2514 -270
rect 628 -464 1346 -456
rect 578 -476 1346 -464
rect 1416 -476 1950 -446
rect 2692 -430 2788 -414
rect 2692 -456 2738 -430
rect 2020 -464 2738 -456
rect 2772 -464 2788 -430
rect 2020 -476 2788 -464
rect 644 -486 1346 -476
rect 644 -502 674 -486
rect 740 -502 770 -486
rect 836 -502 866 -486
rect 932 -502 962 -486
rect 1028 -502 1058 -486
rect 1124 -502 1154 -486
rect 1220 -502 1250 -486
rect 1316 -502 1346 -486
rect 1524 -502 1554 -476
rect 1620 -502 1650 -476
rect 1716 -502 1746 -476
rect 1812 -502 1842 -476
rect 2020 -486 2722 -476
rect 2020 -502 2050 -486
rect 2116 -502 2146 -486
rect 2212 -502 2242 -486
rect 2308 -502 2338 -486
rect 2404 -502 2434 -486
rect 2500 -502 2530 -486
rect 2596 -502 2626 -486
rect 2692 -502 2722 -486
rect 644 -728 674 -702
rect 740 -728 770 -702
rect 836 -728 866 -702
rect 932 -728 962 -702
rect 1028 -728 1058 -702
rect 1124 -728 1154 -702
rect 1220 -728 1250 -702
rect 1316 -728 1346 -702
rect 1524 -728 1554 -702
rect 1620 -728 1650 -702
rect 1716 -728 1746 -702
rect 1812 -728 1842 -702
rect 2020 -728 2050 -702
rect 2116 -728 2146 -702
rect 2212 -728 2242 -702
rect 2308 -728 2338 -702
rect 2404 -728 2434 -702
rect 2500 -728 2530 -702
rect 2596 -728 2626 -702
rect 2692 -728 2722 -702
rect 534 -1098 564 -1072
rect 622 -1098 652 -1072
rect 1628 -1092 1658 -1066
rect 1716 -1092 1746 -1066
rect 822 -1182 852 -1156
rect 1026 -1174 1056 -1148
rect 1122 -1174 1152 -1148
rect 1218 -1174 1248 -1148
rect 1422 -1182 1452 -1156
rect 1920 -1182 1950 -1156
rect 2124 -1174 2154 -1148
rect 2220 -1174 2250 -1148
rect 2316 -1174 2346 -1148
rect 534 -1553 564 -1266
rect 622 -1456 652 -1266
rect 822 -1290 852 -1266
rect 768 -1306 852 -1290
rect 768 -1340 784 -1306
rect 818 -1340 852 -1306
rect 1026 -1282 1056 -1266
rect 1122 -1282 1152 -1266
rect 1218 -1282 1248 -1266
rect 1026 -1312 1248 -1282
rect 768 -1356 852 -1340
rect 622 -1472 704 -1456
rect 622 -1506 654 -1472
rect 688 -1506 704 -1472
rect 622 -1522 704 -1506
rect 622 -1553 652 -1522
rect 822 -1553 852 -1356
rect 1216 -1394 1248 -1312
rect 1422 -1394 1452 -1266
rect 1628 -1286 1658 -1260
rect 1592 -1300 1658 -1286
rect 1592 -1334 1608 -1300
rect 1642 -1334 1658 -1300
rect 1592 -1348 1658 -1334
rect 1716 -1286 1746 -1260
rect 1716 -1300 1782 -1286
rect 1716 -1334 1732 -1300
rect 1766 -1334 1782 -1300
rect 1716 -1348 1782 -1334
rect 1216 -1408 1314 -1394
rect 1216 -1442 1264 -1408
rect 1298 -1442 1314 -1408
rect 1216 -1456 1314 -1442
rect 1422 -1408 1506 -1394
rect 1422 -1442 1456 -1408
rect 1490 -1442 1506 -1408
rect 1422 -1456 1506 -1442
rect 1716 -1404 1782 -1390
rect 1920 -1394 1950 -1266
rect 2124 -1282 2154 -1266
rect 2220 -1282 2250 -1266
rect 2316 -1282 2346 -1266
rect 2124 -1312 2346 -1282
rect 2124 -1394 2156 -1312
rect 1716 -1438 1732 -1404
rect 1766 -1438 1782 -1404
rect 1716 -1452 1782 -1438
rect 1872 -1408 1950 -1394
rect 1872 -1442 1888 -1408
rect 1922 -1442 1950 -1408
rect 1216 -1508 1248 -1456
rect 1026 -1538 1248 -1508
rect 1026 -1553 1056 -1538
rect 1122 -1553 1152 -1538
rect 1218 -1553 1248 -1538
rect 1422 -1553 1452 -1456
rect 1592 -1472 1658 -1458
rect 1592 -1506 1608 -1472
rect 1642 -1506 1658 -1472
rect 1592 -1520 1658 -1506
rect 1628 -1553 1658 -1520
rect 1716 -1553 1746 -1452
rect 1872 -1456 1950 -1442
rect 2060 -1408 2156 -1394
rect 2060 -1442 2076 -1408
rect 2110 -1442 2156 -1408
rect 2060 -1456 2156 -1442
rect 1920 -1553 1950 -1456
rect 2124 -1508 2156 -1456
rect 2124 -1538 2346 -1508
rect 2124 -1553 2154 -1538
rect 2220 -1553 2250 -1538
rect 2316 -1553 2346 -1538
rect 534 -1752 564 -1721
rect 622 -1752 652 -1721
rect 822 -1752 852 -1721
rect 1026 -1747 1056 -1721
rect 1122 -1752 1152 -1721
rect 1218 -1747 1248 -1721
rect 1422 -1752 1452 -1721
rect 1628 -1752 1658 -1721
rect 1716 -1752 1746 -1721
rect 1920 -1752 1950 -1721
rect 2124 -1747 2154 -1721
rect 2220 -1752 2250 -1721
rect 2316 -1747 2346 -1721
rect 482 -1768 564 -1752
rect 482 -1802 498 -1768
rect 532 -1802 564 -1768
rect 482 -1818 564 -1802
<< polycont >>
rect 1056 -26 1090 8
rect 1278 -72 1312 -38
rect 594 -464 628 -430
rect 1504 -72 1538 -38
rect 1828 -140 1862 -106
rect 1666 -432 1700 -398
rect 2272 -26 2306 8
rect 2052 -136 2086 -102
rect 2738 -464 2772 -430
rect 784 -1340 818 -1306
rect 654 -1506 688 -1472
rect 1608 -1334 1642 -1300
rect 1732 -1334 1766 -1300
rect 1264 -1442 1298 -1408
rect 1456 -1442 1490 -1408
rect 1732 -1438 1766 -1404
rect 1888 -1442 1922 -1408
rect 1608 -1506 1642 -1472
rect 2076 -1442 2110 -1408
rect 498 -1802 532 -1768
<< locali >>
rect 762 412 2624 428
rect 762 378 802 412
rect 836 378 958 412
rect 992 378 1114 412
rect 1148 378 1270 412
rect 1304 378 1426 412
rect 1460 378 1582 412
rect 1616 378 1738 412
rect 1772 378 1894 412
rect 1928 378 2050 412
rect 2084 378 2206 412
rect 2240 378 2362 412
rect 2396 378 2518 412
rect 2552 378 2624 412
rect 762 364 2624 378
rect 802 297 836 313
rect 802 137 836 153
rect 898 297 932 364
rect 898 137 932 153
rect 994 297 1028 313
rect 994 137 1028 153
rect 1090 297 1124 364
rect 1090 137 1124 153
rect 1202 297 1236 313
rect 1202 137 1236 153
rect 1290 297 1324 364
rect 1290 137 1324 153
rect 1402 297 1436 313
rect 1402 105 1436 121
rect 1490 297 1524 364
rect 1490 105 1524 121
rect 1578 297 1612 313
rect 1578 105 1612 121
rect 1666 297 1700 364
rect 1666 105 1700 121
rect 1754 297 1788 313
rect 1754 105 1788 121
rect 1842 297 1876 364
rect 1842 105 1876 121
rect 1930 297 1964 313
rect 2042 297 2076 364
rect 2042 137 2076 153
rect 2130 297 2164 313
rect 2130 137 2164 153
rect 2242 297 2276 364
rect 2242 137 2276 153
rect 2338 297 2372 313
rect 2338 137 2372 153
rect 2434 297 2468 364
rect 2434 137 2468 153
rect 2530 297 2564 313
rect 2530 137 2564 153
rect 1930 105 1964 121
rect 1040 -26 1056 8
rect 1090 -26 1106 8
rect 2256 -26 2272 8
rect 2306 -26 2322 8
rect 1262 -72 1278 -38
rect 1312 -72 1328 -38
rect 1488 -72 1504 -38
rect 1538 -72 1554 -38
rect 1812 -140 1828 -106
rect 1862 -140 1878 -106
rect 2036 -136 2052 -102
rect 2086 -136 2102 -102
rect 802 -190 836 -174
rect 802 -274 836 -258
rect 898 -190 932 -174
rect 898 -324 932 -258
rect 994 -190 1028 -174
rect 994 -274 1028 -258
rect 1090 -190 1124 -174
rect 1090 -324 1124 -258
rect 1202 -190 1236 -174
rect 1202 -266 1236 -250
rect 1290 -190 1324 -174
rect 1290 -324 1324 -250
rect 1490 -190 1524 -174
rect 826 -336 1338 -324
rect 826 -370 868 -336
rect 902 -370 968 -336
rect 1002 -370 1068 -336
rect 1102 -370 1168 -336
rect 1202 -370 1268 -336
rect 1302 -370 1338 -336
rect 826 -382 1338 -370
rect 1490 -382 1524 -366
rect 1578 -190 1612 -174
rect 1578 -382 1612 -366
rect 1754 -190 1788 -174
rect 1754 -382 1788 -366
rect 1842 -190 1876 -174
rect 2042 -190 2076 -174
rect 2042 -324 2076 -250
rect 2130 -190 2164 -174
rect 2130 -266 2164 -250
rect 2242 -190 2276 -174
rect 2242 -324 2276 -258
rect 2338 -190 2372 -174
rect 2338 -274 2372 -258
rect 2434 -190 2468 -174
rect 2434 -324 2468 -258
rect 2530 -190 2564 -174
rect 2530 -274 2564 -258
rect 1842 -382 1876 -366
rect 2028 -336 2540 -324
rect 2028 -370 2070 -336
rect 2104 -370 2170 -336
rect 2204 -370 2270 -336
rect 2304 -370 2370 -336
rect 2404 -370 2470 -336
rect 2504 -370 2540 -336
rect 2028 -382 2540 -370
rect 578 -464 594 -430
rect 628 -464 644 -430
rect 1650 -432 1666 -398
rect 1700 -432 1716 -398
rect 2722 -464 2738 -430
rect 2772 -464 2788 -430
rect 594 -514 628 -498
rect 594 -706 628 -690
rect 690 -514 724 -498
rect 690 -706 724 -690
rect 786 -514 820 -498
rect 786 -706 820 -690
rect 882 -514 916 -498
rect 882 -706 916 -690
rect 978 -514 1012 -498
rect 978 -706 1012 -690
rect 1074 -514 1108 -498
rect 1074 -706 1108 -690
rect 1170 -514 1204 -498
rect 1170 -706 1204 -690
rect 1266 -514 1300 -498
rect 1266 -706 1300 -690
rect 1362 -514 1396 -498
rect 1362 -706 1396 -690
rect 1474 -514 1508 -498
rect 1474 -706 1508 -690
rect 1570 -514 1604 -498
rect 1570 -792 1604 -690
rect 1666 -514 1700 -498
rect 1666 -706 1700 -690
rect 1762 -514 1796 -498
rect 1762 -792 1796 -690
rect 1858 -514 1892 -498
rect 1858 -706 1892 -690
rect 1970 -514 2004 -498
rect 1970 -706 2004 -690
rect 2066 -514 2100 -498
rect 2066 -706 2100 -690
rect 2162 -514 2196 -498
rect 2162 -706 2196 -690
rect 2258 -514 2292 -498
rect 2258 -706 2292 -690
rect 2354 -514 2388 -498
rect 2354 -706 2388 -690
rect 2450 -514 2484 -498
rect 2450 -706 2484 -690
rect 2546 -514 2580 -498
rect 2546 -706 2580 -690
rect 2642 -514 2676 -498
rect 2642 -706 2676 -690
rect 2738 -514 2772 -498
rect 2738 -706 2772 -690
rect 544 -816 2834 -792
rect 544 -850 568 -816
rect 602 -850 668 -816
rect 702 -850 768 -816
rect 802 -850 868 -816
rect 902 -850 968 -816
rect 1002 -850 1068 -816
rect 1102 -850 1168 -816
rect 1202 -850 1268 -816
rect 1302 -850 1368 -816
rect 1402 -850 1468 -816
rect 1502 -850 1568 -816
rect 1602 -850 1668 -816
rect 1702 -850 1768 -816
rect 1802 -850 1868 -816
rect 1902 -850 1968 -816
rect 2002 -850 2068 -816
rect 2102 -850 2168 -816
rect 2202 -850 2268 -816
rect 2302 -850 2368 -816
rect 2402 -850 2468 -816
rect 2502 -850 2568 -816
rect 2602 -850 2668 -816
rect 2702 -850 2768 -816
rect 2802 -850 2834 -816
rect 544 -976 2834 -850
rect 544 -1010 568 -976
rect 602 -1010 668 -976
rect 702 -980 2834 -976
rect 702 -1010 1568 -980
rect 544 -1014 1568 -1010
rect 1602 -1014 1668 -980
rect 1702 -1014 1768 -980
rect 1802 -1014 2834 -980
rect 544 -1034 2834 -1014
rect 488 -1110 522 -1094
rect 488 -1270 522 -1254
rect 576 -1110 610 -1094
rect 576 -1270 610 -1254
rect 664 -1110 698 -1034
rect 764 -1038 2834 -1034
rect 764 -1062 1516 -1038
rect 764 -1096 770 -1062
rect 804 -1096 868 -1062
rect 902 -1096 968 -1062
rect 1002 -1096 1068 -1062
rect 1102 -1096 1168 -1062
rect 1202 -1096 1268 -1062
rect 1302 -1096 1368 -1062
rect 1402 -1096 1468 -1062
rect 1502 -1096 1516 -1062
rect 764 -1120 1516 -1096
rect 1582 -1104 1616 -1088
rect 664 -1270 698 -1254
rect 776 -1194 810 -1120
rect 776 -1270 810 -1254
rect 864 -1194 898 -1178
rect 864 -1270 898 -1254
rect 976 -1186 1010 -1170
rect 976 -1270 1010 -1254
rect 1072 -1186 1106 -1120
rect 1072 -1270 1106 -1254
rect 1168 -1186 1202 -1170
rect 1168 -1270 1202 -1254
rect 1264 -1186 1298 -1120
rect 1264 -1270 1298 -1254
rect 1376 -1194 1410 -1178
rect 1376 -1270 1410 -1254
rect 1464 -1194 1498 -1120
rect 1464 -1270 1498 -1254
rect 1582 -1264 1616 -1248
rect 1670 -1104 1704 -1038
rect 1860 -1062 2834 -1038
rect 1670 -1264 1704 -1248
rect 1758 -1104 1792 -1088
rect 1860 -1096 1868 -1062
rect 1902 -1096 1968 -1062
rect 2002 -1096 2068 -1062
rect 2102 -1096 2168 -1062
rect 2202 -1096 2268 -1062
rect 2302 -1096 2368 -1062
rect 2402 -1096 2468 -1062
rect 2502 -1096 2568 -1062
rect 2602 -1096 2668 -1062
rect 2702 -1096 2768 -1062
rect 2802 -1096 2834 -1062
rect 1860 -1120 2834 -1096
rect 1758 -1264 1792 -1248
rect 1874 -1194 1908 -1120
rect 1874 -1270 1908 -1254
rect 1962 -1194 1996 -1178
rect 1962 -1270 1996 -1254
rect 2074 -1186 2108 -1120
rect 2074 -1270 2108 -1254
rect 2170 -1186 2204 -1170
rect 2170 -1270 2204 -1254
rect 2266 -1186 2300 -1120
rect 2266 -1270 2300 -1254
rect 2362 -1186 2396 -1170
rect 2362 -1270 2396 -1254
rect 768 -1340 784 -1306
rect 818 -1340 834 -1306
rect 1592 -1334 1608 -1300
rect 1642 -1334 1658 -1300
rect 1716 -1334 1732 -1300
rect 1766 -1334 1782 -1300
rect 1248 -1442 1264 -1408
rect 1298 -1442 1314 -1408
rect 1440 -1442 1456 -1408
rect 1490 -1442 1506 -1408
rect 1716 -1438 1732 -1404
rect 1766 -1438 1782 -1404
rect 1872 -1442 1888 -1408
rect 1922 -1442 1938 -1408
rect 2060 -1442 2076 -1408
rect 2110 -1442 2126 -1408
rect 488 -1506 654 -1472
rect 688 -1506 704 -1472
rect 1592 -1506 1608 -1472
rect 1642 -1506 1658 -1472
rect 488 -1565 522 -1506
rect 488 -1725 522 -1709
rect 576 -1565 610 -1549
rect 576 -1725 610 -1709
rect 664 -1565 698 -1549
rect 664 -1725 698 -1709
rect 776 -1565 810 -1549
rect 482 -1802 498 -1768
rect 532 -1802 548 -1768
rect 776 -1776 810 -1709
rect 864 -1565 898 -1549
rect 864 -1725 898 -1709
rect 976 -1565 1010 -1549
rect 976 -1725 1010 -1709
rect 1072 -1565 1106 -1549
rect 1072 -1776 1106 -1709
rect 1168 -1565 1202 -1549
rect 1168 -1725 1202 -1709
rect 1264 -1565 1298 -1549
rect 1264 -1776 1298 -1709
rect 1376 -1565 1410 -1549
rect 1376 -1725 1410 -1709
rect 1464 -1565 1498 -1549
rect 1464 -1776 1498 -1709
rect 1582 -1565 1616 -1549
rect 1582 -1725 1616 -1709
rect 1670 -1565 1704 -1549
rect 1670 -1776 1704 -1709
rect 1758 -1565 1792 -1549
rect 1758 -1725 1792 -1709
rect 1874 -1565 1908 -1549
rect 1874 -1776 1908 -1709
rect 1962 -1565 1996 -1549
rect 1962 -1725 1996 -1709
rect 2074 -1565 2108 -1549
rect 2074 -1776 2108 -1709
rect 2170 -1565 2204 -1549
rect 2170 -1725 2204 -1709
rect 2266 -1565 2300 -1549
rect 2266 -1776 2300 -1709
rect 2362 -1565 2396 -1549
rect 2362 -1725 2396 -1709
rect 758 -1792 2440 -1776
rect 758 -1826 818 -1792
rect 852 -1826 958 -1792
rect 992 -1826 1114 -1792
rect 1148 -1826 1270 -1792
rect 1304 -1826 1426 -1792
rect 1460 -1826 1582 -1792
rect 1616 -1826 1738 -1792
rect 1772 -1826 1894 -1792
rect 1928 -1826 2050 -1792
rect 2084 -1826 2206 -1792
rect 2240 -1826 2362 -1792
rect 2396 -1826 2440 -1792
rect 758 -1840 2440 -1826
<< viali >>
rect 802 378 836 412
rect 958 378 992 412
rect 1114 378 1148 412
rect 1270 378 1304 412
rect 1426 378 1460 412
rect 1582 378 1616 412
rect 1738 378 1772 412
rect 1894 378 1928 412
rect 2050 378 2084 412
rect 2206 378 2240 412
rect 2362 378 2396 412
rect 2518 378 2552 412
rect 802 153 836 297
rect 898 153 932 297
rect 994 153 1028 297
rect 1090 153 1124 297
rect 1202 153 1236 297
rect 1290 153 1324 297
rect 1402 121 1436 297
rect 1490 121 1524 297
rect 1578 121 1612 297
rect 1666 121 1700 297
rect 1754 121 1788 297
rect 1842 121 1876 297
rect 1930 121 1964 297
rect 2042 153 2076 297
rect 2130 153 2164 297
rect 2242 153 2276 297
rect 2338 153 2372 297
rect 2434 153 2468 297
rect 2530 153 2564 297
rect 1056 -26 1090 8
rect 2272 -26 2306 8
rect 1278 -72 1312 -38
rect 1504 -72 1538 -38
rect 1828 -140 1862 -106
rect 2052 -136 2086 -102
rect 802 -258 836 -190
rect 898 -258 932 -190
rect 994 -258 1028 -190
rect 1090 -258 1124 -190
rect 1202 -250 1236 -190
rect 1290 -250 1324 -190
rect 868 -370 902 -336
rect 968 -370 1002 -336
rect 1068 -370 1102 -336
rect 1168 -370 1202 -336
rect 1268 -370 1302 -336
rect 1490 -366 1524 -190
rect 1578 -366 1612 -190
rect 1754 -366 1788 -190
rect 1842 -366 1876 -190
rect 2042 -250 2076 -190
rect 2130 -250 2164 -190
rect 2242 -258 2276 -190
rect 2338 -258 2372 -190
rect 2434 -258 2468 -190
rect 2530 -258 2564 -190
rect 2070 -370 2104 -336
rect 2170 -370 2204 -336
rect 2270 -370 2304 -336
rect 2370 -370 2404 -336
rect 2470 -370 2504 -336
rect 594 -464 628 -430
rect 1666 -432 1700 -398
rect 2738 -464 2772 -430
rect 594 -690 628 -514
rect 690 -690 724 -514
rect 786 -690 820 -514
rect 882 -690 916 -514
rect 978 -690 1012 -514
rect 1074 -690 1108 -514
rect 1170 -690 1204 -514
rect 1266 -690 1300 -514
rect 1362 -690 1396 -514
rect 1474 -690 1508 -514
rect 1570 -690 1604 -514
rect 1666 -690 1700 -514
rect 1762 -690 1796 -514
rect 1858 -690 1892 -514
rect 1970 -690 2004 -514
rect 2066 -690 2100 -514
rect 2162 -690 2196 -514
rect 2258 -690 2292 -514
rect 2354 -690 2388 -514
rect 2450 -690 2484 -514
rect 2546 -690 2580 -514
rect 2642 -690 2676 -514
rect 2738 -690 2772 -514
rect 568 -850 602 -816
rect 668 -850 702 -816
rect 768 -850 802 -816
rect 868 -850 902 -816
rect 968 -850 1002 -816
rect 1068 -850 1102 -816
rect 1168 -850 1202 -816
rect 1268 -850 1302 -816
rect 1368 -850 1402 -816
rect 1468 -850 1502 -816
rect 1568 -850 1602 -816
rect 1668 -850 1702 -816
rect 1768 -850 1802 -816
rect 1868 -850 1902 -816
rect 1968 -850 2002 -816
rect 2068 -850 2102 -816
rect 2168 -850 2202 -816
rect 2268 -850 2302 -816
rect 2368 -850 2402 -816
rect 2468 -850 2502 -816
rect 2568 -850 2602 -816
rect 2668 -850 2702 -816
rect 2768 -850 2802 -816
rect 568 -1010 602 -976
rect 668 -1010 702 -976
rect 1568 -1014 1602 -980
rect 1668 -1014 1702 -980
rect 1768 -1014 1802 -980
rect 488 -1254 522 -1110
rect 576 -1254 610 -1110
rect 664 -1254 698 -1110
rect 770 -1096 804 -1062
rect 868 -1096 902 -1062
rect 968 -1096 1002 -1062
rect 1068 -1096 1102 -1062
rect 1168 -1096 1202 -1062
rect 1268 -1096 1302 -1062
rect 1368 -1096 1402 -1062
rect 1468 -1096 1502 -1062
rect 776 -1254 810 -1194
rect 864 -1254 898 -1194
rect 976 -1254 1010 -1186
rect 1072 -1254 1106 -1186
rect 1168 -1254 1202 -1186
rect 1264 -1254 1298 -1186
rect 1376 -1254 1410 -1194
rect 1464 -1254 1498 -1194
rect 1582 -1248 1616 -1104
rect 1670 -1248 1704 -1104
rect 1758 -1248 1792 -1104
rect 1868 -1096 1902 -1062
rect 1968 -1096 2002 -1062
rect 2068 -1096 2102 -1062
rect 2168 -1096 2202 -1062
rect 2268 -1096 2302 -1062
rect 2368 -1096 2402 -1062
rect 2468 -1096 2502 -1062
rect 2568 -1096 2602 -1062
rect 2668 -1096 2702 -1062
rect 2768 -1096 2802 -1062
rect 1874 -1254 1908 -1194
rect 1962 -1254 1996 -1194
rect 2074 -1254 2108 -1186
rect 2170 -1254 2204 -1186
rect 2266 -1254 2300 -1186
rect 2362 -1254 2396 -1186
rect 784 -1340 818 -1306
rect 1608 -1334 1642 -1300
rect 1732 -1334 1766 -1300
rect 1264 -1442 1298 -1408
rect 1456 -1442 1490 -1408
rect 1732 -1438 1766 -1404
rect 1888 -1442 1922 -1408
rect 2076 -1442 2110 -1408
rect 654 -1506 688 -1472
rect 1608 -1506 1642 -1472
rect 488 -1709 522 -1565
rect 576 -1709 610 -1565
rect 664 -1709 698 -1565
rect 776 -1709 810 -1565
rect 498 -1802 532 -1768
rect 864 -1709 898 -1565
rect 976 -1709 1010 -1565
rect 1072 -1709 1106 -1565
rect 1168 -1709 1202 -1565
rect 1264 -1709 1298 -1565
rect 1376 -1709 1410 -1565
rect 1464 -1709 1498 -1565
rect 1582 -1709 1616 -1565
rect 1670 -1709 1704 -1565
rect 1758 -1709 1792 -1565
rect 1874 -1709 1908 -1565
rect 1962 -1709 1996 -1565
rect 2074 -1709 2108 -1565
rect 2170 -1709 2204 -1565
rect 2266 -1709 2300 -1565
rect 2362 -1709 2396 -1565
rect 818 -1826 852 -1792
rect 958 -1826 992 -1792
rect 1114 -1826 1148 -1792
rect 1270 -1826 1304 -1792
rect 1426 -1826 1460 -1792
rect 1582 -1826 1616 -1792
rect 1738 -1826 1772 -1792
rect 1894 -1826 1928 -1792
rect 2050 -1826 2084 -1792
rect 2206 -1826 2240 -1792
rect 2362 -1826 2396 -1792
<< metal1 >>
rect 762 422 2834 428
rect 762 412 2776 422
rect 762 378 802 412
rect 836 378 958 412
rect 992 378 1114 412
rect 1148 378 1270 412
rect 1304 378 1426 412
rect 1460 378 1582 412
rect 1616 378 1738 412
rect 1772 378 1894 412
rect 1928 378 2050 412
rect 2084 378 2206 412
rect 2240 378 2362 412
rect 2396 378 2518 412
rect 2552 378 2776 412
rect 762 370 2776 378
rect 2828 370 2834 422
rect 762 364 2834 370
rect 796 297 842 309
rect 796 153 802 297
rect 836 153 842 297
rect 796 141 842 153
rect 892 297 938 309
rect 892 153 898 297
rect 932 153 938 297
rect 892 141 938 153
rect 988 297 1034 309
rect 988 153 994 297
rect 1028 153 1034 297
rect 988 141 1034 153
rect 1084 297 1130 309
rect 1084 153 1090 297
rect 1124 153 1130 297
rect 1084 141 1130 153
rect 1196 297 1242 309
rect 1196 153 1202 297
rect 1236 153 1242 297
rect 1196 141 1242 153
rect 1284 297 1330 309
rect 1284 153 1290 297
rect 1324 153 1330 297
rect 1284 141 1330 153
rect 1396 297 1442 309
rect 802 100 836 141
rect 994 100 1028 141
rect 802 66 1028 100
rect 802 -60 836 66
rect 1042 16 1106 22
rect 1042 -36 1048 16
rect 1100 8 1106 16
rect 1202 8 1236 141
rect 1396 121 1402 297
rect 1436 121 1442 297
rect 1396 109 1442 121
rect 1484 297 1530 309
rect 1484 121 1490 297
rect 1524 121 1530 297
rect 1484 109 1530 121
rect 1572 297 1618 309
rect 1572 121 1578 297
rect 1612 121 1618 297
rect 1572 109 1618 121
rect 1660 297 1706 309
rect 1660 121 1666 297
rect 1700 121 1706 297
rect 1660 109 1706 121
rect 1748 297 1794 309
rect 1748 121 1754 297
rect 1788 121 1794 297
rect 1748 109 1794 121
rect 1836 297 1882 309
rect 1836 121 1842 297
rect 1876 121 1882 297
rect 1836 109 1882 121
rect 1924 297 1970 309
rect 1924 121 1930 297
rect 1964 121 1970 297
rect 2036 297 2082 309
rect 2036 153 2042 297
rect 2076 153 2082 297
rect 2036 141 2082 153
rect 2124 297 2170 309
rect 2124 153 2130 297
rect 2164 153 2170 297
rect 2124 141 2170 153
rect 2236 297 2282 309
rect 2236 153 2242 297
rect 2276 153 2282 297
rect 2236 141 2282 153
rect 2332 297 2378 309
rect 2332 153 2338 297
rect 2372 153 2378 297
rect 2332 141 2378 153
rect 2428 297 2474 309
rect 2428 153 2434 297
rect 2468 153 2474 297
rect 2428 141 2474 153
rect 2524 297 2570 309
rect 2524 153 2530 297
rect 2564 153 2570 297
rect 2524 141 2570 153
rect 1924 109 1970 121
rect 1100 -26 1236 8
rect 1100 -36 1106 -26
rect 1042 -42 1106 -36
rect 802 -72 878 -60
rect 802 -124 814 -72
rect 866 -102 878 -72
rect 866 -124 1028 -102
rect 802 -136 1028 -124
rect 802 -178 836 -136
rect 994 -178 1028 -136
rect 1202 -178 1236 -26
rect 1264 -28 1328 -22
rect 1264 -80 1270 -28
rect 1322 -80 1328 -28
rect 1264 -86 1328 -80
rect 1486 -28 1550 -22
rect 1486 -80 1492 -28
rect 1544 -80 1550 -28
rect 1486 -86 1550 -80
rect 1578 -86 1612 109
rect 1754 -18 1788 109
rect 1724 -24 1788 -18
rect 1724 -76 1730 -24
rect 1782 -76 1788 -24
rect 1724 -82 1788 -76
rect 1578 -92 1642 -86
rect 1578 -144 1584 -92
rect 1636 -144 1642 -92
rect 1578 -150 1642 -144
rect 1578 -178 1612 -150
rect 1754 -178 1788 -82
rect 2130 8 2164 141
rect 2338 100 2372 141
rect 2530 112 2564 141
rect 2530 100 2608 112
rect 2338 66 2544 100
rect 2530 48 2544 66
rect 2596 48 2608 100
rect 2530 36 2608 48
rect 2256 16 2320 22
rect 2256 8 2262 16
rect 2130 -26 2262 8
rect 1816 -92 1880 -86
rect 1816 -144 1822 -92
rect 1874 -144 1880 -92
rect 1816 -150 1880 -144
rect 2036 -92 2100 -86
rect 2036 -144 2042 -92
rect 2094 -144 2100 -92
rect 2036 -150 2100 -144
rect 2130 -178 2164 -26
rect 2256 -36 2262 -26
rect 2314 -36 2320 16
rect 2256 -42 2320 -36
rect 2530 -102 2564 36
rect 2338 -136 2564 -102
rect 2338 -178 2372 -136
rect 2530 -178 2564 -136
rect 796 -190 842 -178
rect 796 -258 802 -190
rect 836 -258 842 -190
rect 796 -270 842 -258
rect 892 -190 938 -178
rect 892 -258 898 -190
rect 932 -258 938 -190
rect 892 -270 938 -258
rect 988 -190 1034 -178
rect 988 -258 994 -190
rect 1028 -258 1034 -190
rect 988 -270 1034 -258
rect 1084 -190 1130 -178
rect 1084 -258 1090 -190
rect 1124 -258 1130 -190
rect 1084 -270 1130 -258
rect 1196 -190 1242 -178
rect 1196 -250 1202 -190
rect 1236 -250 1242 -190
rect 1196 -262 1242 -250
rect 1284 -190 1330 -178
rect 1284 -250 1290 -190
rect 1324 -250 1330 -190
rect 1284 -262 1330 -250
rect 1484 -190 1530 -178
rect 826 -336 1338 -324
rect 826 -370 868 -336
rect 902 -370 968 -336
rect 1002 -370 1068 -336
rect 1102 -370 1168 -336
rect 1202 -370 1268 -336
rect 1302 -370 1338 -336
rect 548 -430 640 -380
rect 826 -382 1338 -370
rect 1484 -366 1490 -190
rect 1524 -366 1530 -190
rect 1484 -378 1530 -366
rect 1572 -190 1618 -178
rect 1572 -366 1578 -190
rect 1612 -366 1618 -190
rect 1572 -378 1618 -366
rect 1748 -190 1794 -178
rect 1748 -366 1754 -190
rect 1788 -366 1794 -190
rect 1748 -378 1794 -366
rect 1836 -190 1882 -178
rect 1836 -366 1842 -190
rect 1876 -366 1882 -190
rect 2036 -190 2082 -178
rect 2036 -250 2042 -190
rect 2076 -250 2082 -190
rect 2036 -262 2082 -250
rect 2124 -190 2170 -178
rect 2124 -250 2130 -190
rect 2164 -250 2170 -190
rect 2124 -262 2170 -250
rect 2236 -190 2282 -178
rect 2236 -258 2242 -190
rect 2276 -258 2282 -190
rect 2236 -270 2282 -258
rect 2332 -190 2378 -178
rect 2332 -258 2338 -190
rect 2372 -258 2378 -190
rect 2332 -270 2378 -258
rect 2428 -190 2474 -178
rect 2428 -258 2434 -190
rect 2468 -258 2474 -190
rect 2428 -270 2474 -258
rect 2524 -190 2570 -178
rect 2524 -258 2530 -190
rect 2564 -258 2570 -190
rect 2524 -270 2570 -258
rect 1836 -378 1882 -366
rect 2028 -336 2540 -324
rect 2028 -370 2070 -336
rect 2104 -370 2170 -336
rect 2204 -370 2270 -336
rect 2304 -370 2370 -336
rect 2404 -370 2470 -336
rect 2504 -370 2540 -336
rect 548 -464 594 -430
rect 628 -464 640 -430
rect 1490 -440 1524 -378
rect 548 -470 640 -464
rect 690 -474 1524 -440
rect 1650 -388 1714 -382
rect 1650 -440 1656 -388
rect 1708 -440 1714 -388
rect 1650 -446 1714 -440
rect 1842 -440 1876 -378
rect 2028 -382 2540 -370
rect 2726 -430 2818 -378
rect 1842 -474 2676 -440
rect 2726 -464 2738 -430
rect 2772 -464 2818 -430
rect 2726 -468 2818 -464
rect 2726 -470 2784 -468
rect 690 -502 724 -474
rect 882 -502 916 -474
rect 1074 -502 1108 -474
rect 1266 -502 1300 -474
rect 2066 -502 2100 -474
rect 2258 -502 2292 -474
rect 2450 -502 2484 -474
rect 2642 -502 2676 -474
rect 588 -514 634 -502
rect 588 -690 594 -514
rect 628 -690 634 -514
rect 588 -702 634 -690
rect 684 -514 730 -502
rect 684 -690 690 -514
rect 724 -690 730 -514
rect 684 -702 730 -690
rect 780 -514 826 -502
rect 780 -690 786 -514
rect 820 -690 826 -514
rect 780 -702 826 -690
rect 876 -514 922 -502
rect 876 -690 882 -514
rect 916 -690 922 -514
rect 876 -702 922 -690
rect 972 -514 1018 -502
rect 972 -690 978 -514
rect 1012 -690 1018 -514
rect 972 -702 1018 -690
rect 1068 -514 1114 -502
rect 1068 -690 1074 -514
rect 1108 -690 1114 -514
rect 1068 -702 1114 -690
rect 1164 -514 1210 -502
rect 1164 -690 1170 -514
rect 1204 -690 1210 -514
rect 1164 -702 1210 -690
rect 1260 -514 1306 -502
rect 1260 -690 1266 -514
rect 1300 -690 1306 -514
rect 1260 -702 1306 -690
rect 1356 -514 1402 -502
rect 1356 -690 1362 -514
rect 1396 -690 1402 -514
rect 1356 -702 1402 -690
rect 1468 -514 1514 -502
rect 1468 -690 1474 -514
rect 1508 -690 1514 -514
rect 1468 -702 1514 -690
rect 1564 -514 1610 -502
rect 1564 -690 1570 -514
rect 1604 -690 1610 -514
rect 1564 -702 1610 -690
rect 1660 -514 1706 -502
rect 1660 -690 1666 -514
rect 1700 -690 1706 -514
rect 1660 -702 1706 -690
rect 1756 -514 1802 -502
rect 1756 -690 1762 -514
rect 1796 -690 1802 -514
rect 1756 -702 1802 -690
rect 1852 -514 1898 -502
rect 1852 -690 1858 -514
rect 1892 -690 1898 -514
rect 1852 -702 1898 -690
rect 1964 -514 2010 -502
rect 1964 -690 1970 -514
rect 2004 -690 2010 -514
rect 1964 -702 2010 -690
rect 2060 -514 2106 -502
rect 2060 -690 2066 -514
rect 2100 -690 2106 -514
rect 2060 -702 2106 -690
rect 2156 -514 2202 -502
rect 2156 -690 2162 -514
rect 2196 -690 2202 -514
rect 2156 -702 2202 -690
rect 2252 -514 2298 -502
rect 2252 -690 2258 -514
rect 2292 -690 2298 -514
rect 2252 -702 2298 -690
rect 2348 -514 2394 -502
rect 2348 -690 2354 -514
rect 2388 -690 2394 -514
rect 2348 -702 2394 -690
rect 2444 -514 2490 -502
rect 2444 -690 2450 -514
rect 2484 -690 2490 -514
rect 2444 -702 2490 -690
rect 2540 -514 2586 -502
rect 2540 -690 2546 -514
rect 2580 -690 2586 -514
rect 2540 -702 2586 -690
rect 2636 -514 2682 -502
rect 2636 -690 2642 -514
rect 2676 -690 2682 -514
rect 2636 -702 2682 -690
rect 2732 -514 2778 -502
rect 2732 -690 2738 -514
rect 2772 -690 2778 -514
rect 2732 -702 2778 -690
rect 594 -730 628 -702
rect 786 -730 820 -702
rect 978 -730 1012 -702
rect 1170 -730 1204 -702
rect 1362 -730 1396 -702
rect 1474 -730 1508 -702
rect 1666 -730 1700 -702
rect 1970 -730 2004 -702
rect 2162 -730 2196 -702
rect 2354 -730 2388 -702
rect 2546 -730 2580 -702
rect 2738 -730 2772 -702
rect 594 -764 2772 -730
rect 544 -816 2834 -792
rect 544 -850 568 -816
rect 602 -850 668 -816
rect 702 -850 768 -816
rect 802 -850 868 -816
rect 902 -850 968 -816
rect 1002 -850 1068 -816
rect 1102 -850 1168 -816
rect 1202 -850 1268 -816
rect 1302 -850 1368 -816
rect 1402 -850 1468 -816
rect 1502 -850 1568 -816
rect 1602 -850 1668 -816
rect 1702 -850 1768 -816
rect 1802 -850 1868 -816
rect 1902 -850 1968 -816
rect 2002 -850 2068 -816
rect 2102 -850 2168 -816
rect 2202 -850 2268 -816
rect 2302 -850 2368 -816
rect 2402 -850 2468 -816
rect 2502 -850 2568 -816
rect 2602 -850 2668 -816
rect 2702 -850 2768 -816
rect 2802 -850 2834 -816
rect 544 -976 2834 -850
rect 544 -1010 568 -976
rect 602 -1010 668 -976
rect 702 -980 2834 -976
rect 702 -1010 1568 -980
rect 544 -1014 1568 -1010
rect 1602 -1014 1668 -980
rect 1702 -1014 1768 -980
rect 1802 -1014 2834 -980
rect 544 -1034 2834 -1014
rect 764 -1038 2834 -1034
rect 764 -1062 1516 -1038
rect 764 -1096 770 -1062
rect 804 -1096 868 -1062
rect 902 -1096 968 -1062
rect 1002 -1096 1068 -1062
rect 1102 -1096 1168 -1062
rect 1202 -1096 1268 -1062
rect 1302 -1096 1368 -1062
rect 1402 -1096 1468 -1062
rect 1502 -1096 1516 -1062
rect 1860 -1062 2834 -1038
rect 482 -1110 528 -1098
rect 482 -1254 488 -1110
rect 522 -1254 528 -1110
rect 482 -1266 528 -1254
rect 570 -1110 616 -1098
rect 570 -1254 576 -1110
rect 610 -1254 616 -1110
rect 570 -1266 616 -1254
rect 658 -1110 704 -1098
rect 658 -1254 664 -1110
rect 698 -1254 704 -1110
rect 764 -1120 1516 -1096
rect 1576 -1104 1622 -1092
rect 658 -1266 704 -1254
rect 770 -1194 816 -1182
rect 770 -1254 776 -1194
rect 810 -1254 816 -1194
rect 770 -1266 816 -1254
rect 858 -1194 904 -1182
rect 858 -1254 864 -1194
rect 898 -1254 904 -1194
rect 858 -1266 904 -1254
rect 970 -1186 1016 -1174
rect 970 -1254 976 -1186
rect 1010 -1254 1016 -1186
rect 970 -1266 1016 -1254
rect 1066 -1186 1112 -1174
rect 1066 -1254 1072 -1186
rect 1106 -1254 1112 -1186
rect 1066 -1266 1112 -1254
rect 1162 -1186 1208 -1174
rect 1162 -1254 1168 -1186
rect 1202 -1254 1208 -1186
rect 1162 -1266 1208 -1254
rect 1258 -1186 1304 -1174
rect 1258 -1254 1264 -1186
rect 1298 -1254 1304 -1186
rect 1258 -1266 1304 -1254
rect 1370 -1194 1416 -1182
rect 1370 -1254 1376 -1194
rect 1410 -1254 1416 -1194
rect 1370 -1266 1416 -1254
rect 1458 -1194 1504 -1182
rect 1458 -1254 1464 -1194
rect 1498 -1254 1504 -1194
rect 1576 -1232 1582 -1104
rect 1458 -1266 1504 -1254
rect 1532 -1248 1582 -1232
rect 1616 -1248 1622 -1104
rect 1532 -1260 1622 -1248
rect 1664 -1104 1710 -1092
rect 1664 -1248 1670 -1104
rect 1704 -1248 1710 -1104
rect 1664 -1260 1710 -1248
rect 1752 -1104 1798 -1092
rect 1752 -1248 1758 -1104
rect 1792 -1232 1798 -1104
rect 1860 -1096 1868 -1062
rect 1902 -1096 1968 -1062
rect 2002 -1096 2068 -1062
rect 2102 -1096 2168 -1062
rect 2202 -1096 2268 -1062
rect 2302 -1096 2368 -1062
rect 2402 -1096 2468 -1062
rect 2502 -1096 2568 -1062
rect 2602 -1096 2668 -1062
rect 2702 -1096 2768 -1062
rect 2802 -1096 2834 -1062
rect 1860 -1120 2834 -1096
rect 1868 -1194 1914 -1182
rect 1792 -1248 1840 -1232
rect 1752 -1260 1840 -1248
rect 488 -1306 522 -1266
rect 768 -1306 830 -1300
rect 488 -1340 784 -1306
rect 818 -1340 830 -1306
rect 576 -1553 610 -1340
rect 768 -1346 830 -1340
rect 864 -1438 898 -1266
rect 976 -1294 1010 -1266
rect 1168 -1294 1202 -1266
rect 976 -1328 1202 -1294
rect 864 -1444 928 -1438
rect 640 -1458 704 -1456
rect 638 -1462 704 -1458
rect 638 -1512 646 -1462
rect 640 -1514 646 -1512
rect 698 -1514 704 -1462
rect 640 -1520 704 -1514
rect 864 -1496 870 -1444
rect 922 -1496 928 -1444
rect 864 -1502 928 -1496
rect 976 -1490 1010 -1328
rect 1252 -1408 1310 -1402
rect 1382 -1408 1416 -1266
rect 1252 -1442 1264 -1408
rect 1298 -1442 1416 -1408
rect 1252 -1448 1310 -1442
rect 864 -1553 898 -1502
rect 976 -1524 1202 -1490
rect 976 -1553 1010 -1524
rect 1168 -1553 1202 -1524
rect 1382 -1553 1416 -1442
rect 1444 -1408 1502 -1402
rect 1532 -1404 1566 -1260
rect 1594 -1294 1658 -1288
rect 1594 -1346 1600 -1294
rect 1652 -1346 1658 -1294
rect 1594 -1352 1658 -1346
rect 1714 -1294 1778 -1288
rect 1714 -1346 1720 -1294
rect 1772 -1346 1778 -1294
rect 1714 -1352 1778 -1346
rect 1720 -1404 1778 -1398
rect 1532 -1408 1732 -1404
rect 1444 -1442 1456 -1408
rect 1490 -1438 1732 -1408
rect 1766 -1438 1778 -1404
rect 1490 -1442 1566 -1438
rect 1444 -1448 1502 -1442
rect 1532 -1552 1566 -1442
rect 1720 -1444 1778 -1438
rect 1806 -1408 1840 -1260
rect 1868 -1254 1874 -1194
rect 1908 -1254 1914 -1194
rect 1868 -1266 1914 -1254
rect 1956 -1194 2002 -1182
rect 1956 -1254 1962 -1194
rect 1996 -1254 2002 -1194
rect 1956 -1266 2002 -1254
rect 2068 -1186 2114 -1174
rect 2068 -1254 2074 -1186
rect 2108 -1254 2114 -1186
rect 2068 -1266 2114 -1254
rect 2164 -1186 2210 -1174
rect 2164 -1254 2170 -1186
rect 2204 -1254 2210 -1186
rect 2164 -1266 2210 -1254
rect 2260 -1186 2306 -1174
rect 2260 -1254 2266 -1186
rect 2300 -1254 2306 -1186
rect 2260 -1266 2306 -1254
rect 2356 -1186 2402 -1174
rect 2356 -1254 2362 -1186
rect 2396 -1254 2402 -1186
rect 2356 -1266 2402 -1254
rect 1876 -1408 1934 -1402
rect 1806 -1442 1888 -1408
rect 1922 -1442 1934 -1408
rect 1596 -1472 1654 -1466
rect 1806 -1472 1840 -1442
rect 1876 -1448 1934 -1442
rect 1962 -1408 1996 -1266
rect 2170 -1294 2204 -1266
rect 2362 -1294 2396 -1266
rect 2170 -1328 2396 -1294
rect 2064 -1408 2122 -1402
rect 1962 -1442 2076 -1408
rect 2110 -1442 2122 -1408
rect 1596 -1506 1608 -1472
rect 1642 -1506 1840 -1472
rect 1596 -1512 1654 -1506
rect 1806 -1552 1840 -1506
rect 1532 -1553 1616 -1552
rect 482 -1565 528 -1553
rect 482 -1709 488 -1565
rect 522 -1709 528 -1565
rect 482 -1721 528 -1709
rect 570 -1565 616 -1553
rect 570 -1709 576 -1565
rect 610 -1709 616 -1565
rect 570 -1721 616 -1709
rect 658 -1565 704 -1553
rect 658 -1709 664 -1565
rect 698 -1709 704 -1565
rect 658 -1721 704 -1709
rect 770 -1565 816 -1553
rect 770 -1709 776 -1565
rect 810 -1709 816 -1565
rect 770 -1721 816 -1709
rect 858 -1565 904 -1553
rect 858 -1709 864 -1565
rect 898 -1709 904 -1565
rect 858 -1721 904 -1709
rect 970 -1565 1016 -1553
rect 970 -1709 976 -1565
rect 1010 -1709 1016 -1565
rect 970 -1721 1016 -1709
rect 1066 -1565 1112 -1553
rect 1066 -1709 1072 -1565
rect 1106 -1709 1112 -1565
rect 1066 -1721 1112 -1709
rect 1162 -1565 1208 -1553
rect 1162 -1709 1168 -1565
rect 1202 -1709 1208 -1565
rect 1162 -1721 1208 -1709
rect 1258 -1565 1304 -1553
rect 1258 -1709 1264 -1565
rect 1298 -1709 1304 -1565
rect 1258 -1721 1304 -1709
rect 1370 -1565 1416 -1553
rect 1370 -1709 1376 -1565
rect 1410 -1709 1416 -1565
rect 1370 -1721 1416 -1709
rect 1458 -1565 1504 -1553
rect 1458 -1709 1464 -1565
rect 1498 -1709 1504 -1565
rect 1532 -1565 1622 -1553
rect 1532 -1586 1582 -1565
rect 1458 -1721 1504 -1709
rect 1576 -1709 1582 -1586
rect 1616 -1709 1622 -1565
rect 1576 -1721 1622 -1709
rect 1664 -1565 1710 -1553
rect 1664 -1709 1670 -1565
rect 1704 -1709 1710 -1565
rect 1664 -1721 1710 -1709
rect 1752 -1565 1840 -1552
rect 1962 -1553 1996 -1442
rect 2064 -1448 2122 -1442
rect 2362 -1490 2396 -1328
rect 2170 -1524 2396 -1490
rect 2170 -1553 2204 -1524
rect 2362 -1553 2396 -1524
rect 1752 -1709 1758 -1565
rect 1792 -1586 1840 -1565
rect 1868 -1565 1914 -1553
rect 1792 -1709 1798 -1586
rect 1752 -1721 1798 -1709
rect 1868 -1709 1874 -1565
rect 1908 -1709 1914 -1565
rect 1868 -1721 1914 -1709
rect 1956 -1565 2002 -1553
rect 1956 -1709 1962 -1565
rect 1996 -1709 2002 -1565
rect 1956 -1721 2002 -1709
rect 2068 -1565 2114 -1553
rect 2068 -1709 2074 -1565
rect 2108 -1709 2114 -1565
rect 2068 -1721 2114 -1709
rect 2164 -1565 2210 -1553
rect 2164 -1709 2170 -1565
rect 2204 -1709 2210 -1565
rect 2164 -1721 2210 -1709
rect 2260 -1565 2306 -1553
rect 2260 -1709 2266 -1565
rect 2300 -1709 2306 -1565
rect 2260 -1721 2306 -1709
rect 2356 -1565 2402 -1553
rect 2356 -1709 2362 -1565
rect 2396 -1709 2402 -1565
rect 2356 -1721 2402 -1709
rect 482 -1758 546 -1752
rect 482 -1810 488 -1758
rect 540 -1768 546 -1758
rect 664 -1768 698 -1721
rect 540 -1802 698 -1768
rect 758 -1782 2828 -1776
rect 758 -1792 2770 -1782
rect 540 -1810 546 -1802
rect 482 -1816 546 -1810
rect 758 -1826 818 -1792
rect 852 -1826 958 -1792
rect 992 -1826 1114 -1792
rect 1148 -1826 1270 -1792
rect 1304 -1826 1426 -1792
rect 1460 -1826 1582 -1792
rect 1616 -1826 1738 -1792
rect 1772 -1826 1894 -1792
rect 1928 -1826 2050 -1792
rect 2084 -1826 2206 -1792
rect 2240 -1826 2362 -1792
rect 2396 -1826 2770 -1792
rect 758 -1834 2770 -1826
rect 2822 -1834 2828 -1782
rect 758 -1840 2828 -1834
<< via1 >>
rect 2776 370 2828 422
rect 1048 8 1100 16
rect 1048 -26 1056 8
rect 1056 -26 1090 8
rect 1090 -26 1100 8
rect 1048 -36 1100 -26
rect 814 -124 866 -72
rect 1270 -38 1322 -28
rect 1270 -72 1278 -38
rect 1278 -72 1312 -38
rect 1312 -72 1322 -38
rect 1270 -80 1322 -72
rect 1492 -38 1544 -28
rect 1492 -72 1504 -38
rect 1504 -72 1538 -38
rect 1538 -72 1544 -38
rect 1492 -80 1544 -72
rect 1730 -76 1782 -24
rect 1584 -144 1636 -92
rect 2544 48 2596 100
rect 2262 8 2314 16
rect 2262 -26 2272 8
rect 2272 -26 2306 8
rect 2306 -26 2314 8
rect 1822 -106 1874 -92
rect 1822 -140 1828 -106
rect 1828 -140 1862 -106
rect 1862 -140 1874 -106
rect 1822 -144 1874 -140
rect 2042 -102 2094 -92
rect 2042 -136 2052 -102
rect 2052 -136 2086 -102
rect 2086 -136 2094 -102
rect 2042 -144 2094 -136
rect 2262 -36 2314 -26
rect 1656 -398 1708 -388
rect 1656 -432 1666 -398
rect 1666 -432 1700 -398
rect 1700 -432 1708 -398
rect 1656 -440 1708 -432
rect 646 -1472 698 -1462
rect 646 -1506 654 -1472
rect 654 -1506 688 -1472
rect 688 -1506 698 -1472
rect 646 -1514 698 -1506
rect 870 -1496 922 -1444
rect 1600 -1300 1652 -1294
rect 1600 -1334 1608 -1300
rect 1608 -1334 1642 -1300
rect 1642 -1334 1652 -1300
rect 1600 -1346 1652 -1334
rect 1720 -1300 1772 -1294
rect 1720 -1334 1732 -1300
rect 1732 -1334 1766 -1300
rect 1766 -1334 1772 -1300
rect 1720 -1346 1772 -1334
rect 488 -1768 540 -1758
rect 488 -1802 498 -1768
rect 498 -1802 532 -1768
rect 532 -1802 540 -1768
rect 488 -1810 540 -1802
rect 2770 -1834 2822 -1782
<< metal2 >>
rect 2770 422 2834 428
rect 2770 370 2776 422
rect 2828 370 2834 422
rect 2770 364 2834 370
rect 488 102 564 112
rect 488 46 498 102
rect 554 46 564 102
rect 488 36 564 46
rect 488 -1752 516 36
rect 670 -60 698 112
rect 2532 102 2608 112
rect 2532 46 2542 102
rect 2598 46 2608 102
rect 2532 36 2608 46
rect 1042 16 1106 22
rect 1042 -36 1048 16
rect 1100 -36 1106 16
rect 2256 16 2320 22
rect 1042 -42 1106 -36
rect 1264 -24 1550 -22
rect 1724 -24 1788 -18
rect 1264 -28 1730 -24
rect 658 -70 734 -60
rect 658 -126 668 -70
rect 724 -126 734 -70
rect 658 -136 734 -126
rect 802 -70 878 -60
rect 802 -126 812 -70
rect 868 -126 878 -70
rect 802 -136 878 -126
rect 670 -1456 698 -136
rect 1062 -982 1090 -42
rect 1264 -80 1270 -28
rect 1322 -56 1492 -28
rect 1322 -80 1328 -56
rect 1264 -86 1328 -80
rect 1486 -80 1492 -56
rect 1544 -58 1730 -28
rect 1544 -80 1550 -58
rect 1486 -86 1550 -80
rect 1724 -76 1730 -58
rect 1782 -76 1788 -24
rect 2256 -36 2262 16
rect 2314 -36 2320 16
rect 2256 -42 2320 -36
rect 1724 -82 1788 -76
rect 1578 -92 1642 -86
rect 1578 -144 1584 -92
rect 1636 -116 1642 -92
rect 1816 -92 1880 -86
rect 1816 -116 1822 -92
rect 1636 -144 1822 -116
rect 1874 -116 1880 -92
rect 2036 -92 2100 -86
rect 2036 -116 2042 -92
rect 1874 -144 2042 -116
rect 2094 -144 2100 -92
rect 1578 -150 2100 -144
rect 1650 -388 1714 -382
rect 1650 -440 1656 -388
rect 1708 -440 1714 -388
rect 1650 -446 1714 -440
rect 2272 -982 2300 -42
rect 1062 -1010 1618 -982
rect 1590 -1288 1618 -1010
rect 1744 -1012 2300 -982
rect 1744 -1288 1772 -1012
rect 1590 -1294 1658 -1288
rect 1590 -1346 1600 -1294
rect 1652 -1346 1658 -1294
rect 1590 -1352 1658 -1346
rect 1714 -1294 1784 -1288
rect 1714 -1346 1720 -1294
rect 1772 -1346 1784 -1294
rect 1714 -1352 1784 -1346
rect 864 -1444 928 -1438
rect 640 -1462 704 -1456
rect 640 -1514 646 -1462
rect 698 -1514 704 -1462
rect 864 -1496 870 -1444
rect 922 -1496 928 -1444
rect 864 -1502 928 -1496
rect 640 -1520 704 -1514
rect 482 -1758 546 -1752
rect 482 -1810 488 -1758
rect 540 -1810 546 -1758
rect 482 -1816 546 -1810
rect 670 -1816 698 -1520
rect 2800 -1776 2828 364
rect 2764 -1782 2828 -1776
rect 2764 -1834 2770 -1782
rect 2822 -1834 2828 -1782
rect 2764 -1840 2828 -1834
<< via2 >>
rect 498 46 554 102
rect 2542 100 2598 102
rect 2542 48 2544 100
rect 2544 48 2596 100
rect 2596 48 2598 100
rect 2542 46 2598 48
rect 668 -126 724 -70
rect 812 -72 868 -70
rect 812 -124 814 -72
rect 814 -124 866 -72
rect 866 -124 868 -72
rect 812 -126 868 -124
<< metal3 >>
rect 488 104 564 112
rect 2532 104 2608 112
rect 488 102 2608 104
rect 488 46 498 102
rect 554 46 2542 102
rect 2598 46 2608 102
rect 488 44 2608 46
rect 488 36 564 44
rect 2532 36 2608 44
rect 658 -66 734 -60
rect 802 -66 878 -60
rect 488 -70 2608 -66
rect 488 -126 668 -70
rect 724 -126 812 -70
rect 868 -126 2608 -70
rect 658 -136 734 -126
rect 802 -136 878 -126
<< labels >>
flabel space 1578 -92 1612 121 0 FreeSans 288 0 0 0 X
flabel space 1754 -24 1788 121 0 FreeSans 288 0 0 0 Y
flabel space 2130 -190 2164 153 0 FreeSans 288 0 0 0 X_inv
flabel space 2530 -190 2564 48 0 FreeSans 288 0 0 0 X_drive
flabel metal1 2726 -468 2818 -378 0 FreeSans 288 0 0 0 cdac_vn
port 1 nsew
flabel metal1 548 -470 640 -380 0 FreeSans 288 0 0 0 cdac_vp
port 2 nsew
flabel space 1202 -220 1236 153 0 FreeSans 240 0 0 0 Y_inv
flabel space 802 -72 836 153 0 FreeSans 240 0 0 0 Y_drive
flabel space 864 -1444 898 -1254 0 FreeSans 240 0 0 0 ready
port 3 nsew
flabel metal1 2362 -1609 2396 -1254 0 FreeSans 240 0 0 0 comp_outp
port 5 nsew
flabel metal1 976 -1609 1010 -1254 0 FreeSans 240 0 0 0 comp_outn
port 6 nsew
flabel metal1 1806 -1586 1840 -1232 0 FreeSans 240 0 0 0 RS_p
flabel metal1 1532 -1586 1566 -1232 0 FreeSans 240 0 0 0 RS_n
flabel via1 1656 -440 1708 -388 0 FreeSans 240 0 0 0 clk
port 7 nsew
flabel metal1 836 364 958 428 0 FreeSans 240 0 0 0 VDD
port 8 nsew
flabel metal1 702 -980 2834 -850 0 FreeSans 240 0 0 0 VSS
port 9 nsew
<< end >>
