magic
tech sky130A
magscale 1 2
timestamp 1701018915
<< nwell >>
rect 2877 38830 2941 38831
rect 1279 38265 3154 38830
rect 1279 38264 1569 38265
rect 1629 37421 3020 37437
rect 1463 37186 3020 37421
rect 1463 37177 2960 37186
rect 1463 37176 1925 37177
<< psubdiff >>
rect 924 39679 5204 39727
rect 924 39519 1306 39679
rect 1466 39519 1706 39679
rect 1866 39519 2106 39679
rect 2266 39519 2506 39679
rect 2666 39519 2906 39679
rect 3066 39519 3306 39679
rect 3466 39519 3706 39679
rect 3866 39519 4106 39679
rect 4266 39519 4506 39679
rect 4666 39519 5204 39679
rect 924 39496 5204 39519
rect 924 39336 980 39496
rect 1140 39476 4983 39496
rect 1140 39336 1187 39476
rect 924 39096 1187 39336
rect 924 38936 980 39096
rect 1140 38936 1187 39096
rect 4915 39336 4983 39476
rect 5143 39476 5204 39496
rect 5143 39336 5203 39476
rect 4915 39096 5203 39336
rect 924 38696 1187 38936
rect 4915 38936 4983 39096
rect 5143 38936 5203 39096
rect 924 38536 980 38696
rect 1140 38536 1187 38696
rect 924 38296 1187 38536
rect 924 38136 980 38296
rect 1140 38136 1187 38296
rect 924 37896 1187 38136
rect 924 37736 980 37896
rect 1140 37736 1187 37896
rect 924 37496 1187 37736
rect 924 37336 980 37496
rect 1140 37336 1187 37496
rect 924 37096 1187 37336
rect 4915 38696 5203 38936
rect 4915 38536 4983 38696
rect 5143 38536 5203 38696
rect 4915 38296 5203 38536
rect 4915 38136 4983 38296
rect 5143 38136 5203 38296
rect 4915 37896 5203 38136
rect 4915 37736 4983 37896
rect 5143 37736 5203 37896
rect 4915 37496 5203 37736
rect 4915 37336 4983 37496
rect 5143 37336 5203 37496
rect 924 36936 980 37096
rect 1140 36936 1187 37096
rect 4915 37096 5203 37336
rect 924 36650 1187 36936
rect 4915 36936 4983 37096
rect 5143 36936 5203 37096
rect 4915 36732 5203 36936
rect 4915 36650 5204 36732
rect 924 36649 2538 36650
rect 2685 36649 5204 36650
rect 924 36614 5204 36649
rect 924 36454 980 36614
rect 1140 36454 1408 36614
rect 1568 36454 1808 36614
rect 1968 36454 2208 36614
rect 2368 36609 3408 36614
rect 2368 36454 2742 36609
rect 924 36449 2742 36454
rect 2902 36449 3069 36609
rect 3229 36454 3408 36609
rect 3568 36454 3808 36614
rect 3968 36454 4208 36614
rect 4368 36454 4608 36614
rect 4768 36454 4983 36614
rect 5143 36454 5204 36614
rect 3229 36449 5204 36454
rect 924 36411 5203 36449
<< psubdiffcont >>
rect 1306 39519 1466 39679
rect 1706 39519 1866 39679
rect 2106 39519 2266 39679
rect 2506 39519 2666 39679
rect 2906 39519 3066 39679
rect 3306 39519 3466 39679
rect 3706 39519 3866 39679
rect 4106 39519 4266 39679
rect 4506 39519 4666 39679
rect 980 39336 1140 39496
rect 980 38936 1140 39096
rect 4983 39336 5143 39496
rect 4983 38936 5143 39096
rect 980 38536 1140 38696
rect 980 38136 1140 38296
rect 980 37736 1140 37896
rect 980 37336 1140 37496
rect 4983 38536 5143 38696
rect 4983 38136 5143 38296
rect 4983 37736 5143 37896
rect 4983 37336 5143 37496
rect 980 36936 1140 37096
rect 4983 36936 5143 37096
rect 980 36454 1140 36614
rect 1408 36454 1568 36614
rect 1808 36454 1968 36614
rect 2208 36454 2368 36614
rect 2742 36449 2902 36609
rect 3069 36449 3229 36609
rect 3408 36454 3568 36614
rect 3808 36454 3968 36614
rect 4208 36454 4368 36614
rect 4608 36454 4768 36614
rect 4983 36454 5143 36614
<< poly >>
rect 2885 38981 2951 38994
rect 2885 38966 2901 38981
rect 2039 38964 2901 38966
rect 1650 38947 2901 38964
rect 2935 38947 2951 38981
rect 1650 38934 2951 38947
rect 1650 38870 2965 38892
rect 1650 38862 2921 38870
rect 1650 38819 1750 38862
rect 1808 38819 1908 38862
rect 2081 38816 2181 38862
rect 2239 38817 2339 38862
rect 2526 38817 2626 38862
rect 2684 38817 2784 38862
rect 2911 38836 2921 38862
rect 2955 38836 2965 38870
rect 2911 38820 2965 38836
rect 2526 38816 2538 38817
rect 2003 37144 2103 37197
rect 2161 37144 2261 37198
rect 2483 37144 2583 37198
rect 2641 37144 2741 37197
rect 2884 37172 2952 37182
rect 2884 37144 2902 37172
rect 2003 37138 2902 37144
rect 2936 37138 2952 37172
rect 2003 37114 2952 37138
rect 2003 37040 2969 37070
rect 2900 37038 2969 37040
rect 2900 37003 2916 37038
rect 2953 37003 2969 37038
rect 2900 36992 2969 37003
<< polycont >>
rect 2901 38947 2935 38981
rect 2921 38836 2955 38870
rect 2902 37138 2936 37172
rect 2916 37003 2953 37038
<< locali >>
rect 463 75060 946 75109
rect 463 74984 504 75060
rect 576 74984 626 75060
rect 698 74984 752 75060
rect 824 74984 946 75060
rect 463 74913 946 74984
rect 463 74837 504 74913
rect 576 74837 626 74913
rect 698 74837 752 74913
rect 824 74837 946 74913
rect 463 74776 946 74837
rect 463 74700 504 74776
rect 576 74700 626 74776
rect 698 74700 752 74776
rect 824 74700 946 74776
rect 463 74650 946 74700
rect 463 73300 946 73349
rect 463 73224 504 73300
rect 576 73224 626 73300
rect 698 73224 752 73300
rect 824 73224 946 73300
rect 463 73153 946 73224
rect 463 73077 504 73153
rect 576 73077 626 73153
rect 698 73077 752 73153
rect 824 73077 946 73153
rect 463 73016 946 73077
rect 463 72940 504 73016
rect 576 72940 626 73016
rect 698 72940 752 73016
rect 824 72940 946 73016
rect 463 72890 946 72940
rect 463 71060 946 71109
rect 463 70984 504 71060
rect 576 70984 626 71060
rect 698 70984 752 71060
rect 824 70984 946 71060
rect 463 70913 946 70984
rect 463 70837 504 70913
rect 576 70837 626 70913
rect 698 70837 752 70913
rect 824 70837 946 70913
rect 463 70776 946 70837
rect 463 70700 504 70776
rect 576 70700 626 70776
rect 698 70700 752 70776
rect 824 70700 946 70776
rect 463 70650 946 70700
rect 463 69300 946 69349
rect 463 69224 504 69300
rect 576 69224 626 69300
rect 698 69224 752 69300
rect 824 69224 946 69300
rect 463 69153 946 69224
rect 463 69077 504 69153
rect 576 69077 626 69153
rect 698 69077 752 69153
rect 824 69077 946 69153
rect 463 69016 946 69077
rect 463 68940 504 69016
rect 576 68940 626 69016
rect 698 68940 752 69016
rect 824 68940 946 69016
rect 463 68890 946 68940
rect 463 67060 946 67109
rect 463 66984 504 67060
rect 576 66984 626 67060
rect 698 66984 752 67060
rect 824 66984 946 67060
rect 463 66913 946 66984
rect 463 66837 504 66913
rect 576 66837 626 66913
rect 698 66837 752 66913
rect 824 66837 946 66913
rect 463 66776 946 66837
rect 463 66700 504 66776
rect 576 66700 626 66776
rect 698 66700 752 66776
rect 824 66700 946 66776
rect 463 66650 946 66700
rect 463 65301 946 65350
rect 463 65225 504 65301
rect 576 65225 626 65301
rect 698 65225 752 65301
rect 824 65225 946 65301
rect 463 65154 946 65225
rect 463 65078 504 65154
rect 576 65078 626 65154
rect 698 65078 752 65154
rect 824 65078 946 65154
rect 463 65017 946 65078
rect 463 64941 504 65017
rect 576 64941 626 65017
rect 698 64941 752 65017
rect 824 64941 946 65017
rect 463 64891 946 64941
rect 464 63068 947 63109
rect 463 63060 947 63068
rect 463 62984 504 63060
rect 576 62984 626 63060
rect 698 62984 752 63060
rect 824 62984 947 63060
rect 463 62913 947 62984
rect 463 62837 504 62913
rect 576 62837 626 62913
rect 698 62837 752 62913
rect 824 62837 947 62913
rect 463 62776 947 62837
rect 463 62700 504 62776
rect 576 62700 626 62776
rect 698 62700 752 62776
rect 824 62700 947 62776
rect 463 62650 947 62700
rect 463 61301 946 61350
rect 463 61225 504 61301
rect 576 61225 626 61301
rect 698 61225 752 61301
rect 824 61225 946 61301
rect 463 61154 946 61225
rect 463 61078 504 61154
rect 576 61078 626 61154
rect 698 61078 752 61154
rect 824 61078 946 61154
rect 463 61017 946 61078
rect 463 60941 504 61017
rect 576 60941 626 61017
rect 698 60941 752 61017
rect 824 60941 946 61017
rect 463 60891 946 60941
rect 464 59068 947 59109
rect 463 59060 947 59068
rect 463 58984 504 59060
rect 576 58984 626 59060
rect 698 58984 752 59060
rect 824 58984 947 59060
rect 463 58913 947 58984
rect 463 58837 504 58913
rect 576 58837 626 58913
rect 698 58837 752 58913
rect 824 58837 947 58913
rect 463 58776 947 58837
rect 463 58700 504 58776
rect 576 58700 626 58776
rect 698 58700 752 58776
rect 824 58700 947 58776
rect 463 58650 947 58700
rect 463 57299 946 57348
rect 463 57223 504 57299
rect 576 57223 626 57299
rect 698 57223 752 57299
rect 824 57223 946 57299
rect 463 57152 946 57223
rect 463 57076 504 57152
rect 576 57076 626 57152
rect 698 57076 752 57152
rect 824 57076 946 57152
rect 463 57015 946 57076
rect 463 56939 504 57015
rect 576 56939 626 57015
rect 698 56939 752 57015
rect 824 56939 946 57015
rect 463 56889 946 56939
rect 463 55060 946 55109
rect 463 54984 504 55060
rect 576 54984 626 55060
rect 698 54984 752 55060
rect 824 54984 946 55060
rect 463 54913 946 54984
rect 463 54837 504 54913
rect 576 54837 626 54913
rect 698 54837 752 54913
rect 824 54837 946 54913
rect 463 54776 946 54837
rect 463 54700 504 54776
rect 576 54700 626 54776
rect 698 54700 752 54776
rect 824 54700 946 54776
rect 463 54650 946 54700
rect 463 53301 946 53350
rect 463 53225 504 53301
rect 576 53225 626 53301
rect 698 53225 752 53301
rect 824 53225 946 53301
rect 463 53154 946 53225
rect 463 53078 504 53154
rect 576 53078 626 53154
rect 698 53078 752 53154
rect 824 53078 946 53154
rect 463 53017 946 53078
rect 463 52941 504 53017
rect 576 52941 626 53017
rect 698 52941 752 53017
rect 824 52941 946 53017
rect 463 52891 946 52941
rect 463 51060 946 51109
rect 463 50984 504 51060
rect 576 50984 626 51060
rect 698 50984 752 51060
rect 824 50984 946 51060
rect 463 50913 946 50984
rect 463 50837 504 50913
rect 576 50837 626 50913
rect 698 50837 752 50913
rect 824 50837 946 50913
rect 463 50776 946 50837
rect 463 50700 504 50776
rect 576 50700 626 50776
rect 698 50700 752 50776
rect 824 50700 946 50776
rect 463 50650 946 50700
rect 463 49301 946 49350
rect 463 49225 504 49301
rect 576 49225 626 49301
rect 698 49225 752 49301
rect 824 49225 946 49301
rect 463 49154 946 49225
rect 463 49078 504 49154
rect 576 49078 626 49154
rect 698 49078 752 49154
rect 824 49078 946 49154
rect 463 49017 946 49078
rect 463 48941 504 49017
rect 576 48941 626 49017
rect 698 48941 752 49017
rect 824 48941 946 49017
rect 463 48891 946 48941
rect 463 47060 946 47109
rect 463 46984 504 47060
rect 576 46984 626 47060
rect 698 46984 752 47060
rect 824 46984 946 47060
rect 463 46913 946 46984
rect 463 46837 504 46913
rect 576 46837 626 46913
rect 698 46837 752 46913
rect 824 46837 946 46913
rect 463 46776 946 46837
rect 463 46700 504 46776
rect 576 46700 626 46776
rect 698 46700 752 46776
rect 824 46700 946 46776
rect 463 46650 946 46700
rect 463 45300 946 45350
rect 463 45224 504 45300
rect 576 45224 626 45300
rect 698 45224 752 45300
rect 824 45224 946 45300
rect 463 45153 946 45224
rect 463 45077 504 45153
rect 576 45077 626 45153
rect 698 45077 752 45153
rect 824 45077 946 45153
rect 463 45016 946 45077
rect 463 44940 504 45016
rect 576 44940 626 45016
rect 698 44940 752 45016
rect 824 44940 946 45016
rect 463 44891 946 44940
rect 463 44890 836 44891
rect 924 39679 5204 39727
rect 924 39519 1306 39679
rect 1466 39519 1706 39679
rect 1866 39519 2106 39679
rect 2266 39519 2506 39679
rect 2666 39519 2906 39679
rect 3066 39519 3306 39679
rect 3466 39519 3706 39679
rect 3866 39519 4106 39679
rect 4266 39519 4506 39679
rect 4666 39519 5204 39679
rect 924 39496 5204 39519
rect 924 39336 980 39496
rect 1140 39476 4983 39496
rect 1140 39336 1188 39476
rect 924 39138 1188 39336
rect 1868 39395 2503 39410
rect 1650 39321 1796 39329
rect 1650 39279 1662 39321
rect 1704 39279 1742 39321
rect 1784 39279 1796 39321
rect 1650 39241 1796 39279
rect 1868 39281 1885 39395
rect 2003 39281 2041 39395
rect 2159 39281 2197 39395
rect 2315 39281 2503 39395
rect 4914 39336 4983 39476
rect 5143 39336 5204 39496
rect 1868 39271 2503 39281
rect 1868 39270 2009 39271
rect 1650 39199 1662 39241
rect 1704 39199 1742 39241
rect 1784 39223 1796 39241
rect 2192 39230 2227 39237
rect 1784 39199 2192 39223
rect 1650 39191 2192 39199
rect 1650 39189 2227 39191
rect 924 39137 1098 39138
rect 924 39062 941 39137
rect 1013 39096 1098 39137
rect 1165 39063 1188 39138
rect 924 39021 980 39062
rect 1140 39024 1188 39063
rect 1604 39125 1638 39139
rect 1919 39124 1954 39139
rect 1604 39052 1638 39059
rect 924 38946 944 39021
rect 1165 38949 1188 39024
rect 1762 38999 1796 39090
rect 1919 39069 1920 39124
rect 2192 39078 2227 39189
rect 2351 39085 2503 39271
rect 2539 39328 2685 39336
rect 2539 39286 2551 39328
rect 2593 39286 2631 39328
rect 2673 39286 2685 39328
rect 2539 39248 2685 39286
rect 2539 39206 2551 39248
rect 2593 39206 2631 39248
rect 2673 39206 2685 39248
rect 2539 39196 2685 39206
rect 2638 39085 2672 39196
rect 4914 39108 5204 39336
rect 4721 39096 5204 39108
rect 1919 39058 1953 39069
rect 924 38936 980 38946
rect 1140 38936 1188 38949
rect 924 38696 1188 38936
rect 1604 38944 1638 38989
rect 1604 38797 1638 38889
rect 1762 38798 1796 38977
rect 1920 38944 1954 38989
rect 1920 38797 1954 38889
rect 2035 38944 2069 38997
rect 2035 38796 2069 38889
rect 2193 38795 2227 38988
rect 2351 38977 2514 39085
rect 2793 38977 2831 39085
rect 4721 39074 4983 39096
rect 2351 38944 2385 38977
rect 2351 38796 2385 38889
rect 2479 38949 2514 38977
rect 2479 38851 2514 38889
rect 2480 38797 2514 38851
rect 2638 38797 2672 38977
rect 2796 38949 2831 38977
rect 2796 38890 2797 38949
rect 2885 38981 2951 38982
rect 2885 38947 2901 38981
rect 2935 38947 2951 38981
rect 2885 38946 2951 38947
rect 4914 38936 4983 39074
rect 5143 38936 5204 39096
rect 2796 38851 2831 38890
rect 4315 38870 4557 38876
rect 2796 38797 2830 38851
rect 2900 38836 2921 38870
rect 2955 38836 2973 38870
rect 4315 38836 4339 38870
rect 4373 38836 4557 38870
rect 4315 38828 4557 38836
rect 4591 38871 4663 38876
rect 4591 38836 4615 38871
rect 4650 38836 4663 38871
rect 4591 38829 4663 38836
rect 4591 38828 4638 38829
rect 924 38536 980 38696
rect 1140 38536 1188 38696
rect 924 38296 1188 38536
rect 4914 38696 5204 38936
rect 4914 38536 4983 38696
rect 5143 38536 5204 38696
rect 924 38136 980 38296
rect 1140 38136 1188 38296
rect 1339 38260 1523 38269
rect 1339 38225 1479 38260
rect 1515 38225 1523 38260
rect 1339 38217 1523 38225
rect 2818 38202 2942 38343
rect 3740 38202 3864 38343
rect 4914 38296 5204 38536
rect 4632 38258 4704 38262
rect 4632 38224 4662 38258
rect 4696 38224 4704 38258
rect 4632 38207 4704 38224
rect 924 37896 1188 38136
rect 4914 38136 4983 38296
rect 5143 38136 5204 38296
rect 4914 38020 5204 38136
rect 4812 37986 5204 38020
rect 924 37736 980 37896
rect 1140 37736 1188 37896
rect 4914 37896 5204 37986
rect 1573 37745 1769 37788
rect 924 37496 1188 37736
rect 2818 37663 2942 37804
rect 3740 37663 3864 37804
rect 4696 37748 4704 37780
rect 4675 37745 4704 37748
rect 4914 37736 4983 37896
rect 5143 37736 5204 37896
rect 924 37336 980 37496
rect 1140 37336 1188 37496
rect 4914 37496 5204 37736
rect 1963 37442 1997 37465
rect 924 37096 1188 37336
rect 1680 37358 1739 37375
rect 1680 37310 1686 37358
rect 1732 37310 1739 37358
rect 2114 37312 2149 37451
rect 4914 37336 4983 37496
rect 5143 37336 5204 37496
rect 1680 37245 1739 37310
rect 1680 37200 1686 37245
rect 1732 37200 1739 37245
rect 1680 37187 1739 37200
rect 924 37079 980 37096
rect 1140 37079 1188 37096
rect 924 36991 947 37079
rect 1165 36991 1188 37079
rect 1957 37144 1991 37257
rect 1957 37029 1991 37090
rect 2115 37029 2149 37256
rect 2273 37143 2307 37257
rect 2273 37029 2307 37089
rect 2436 37146 2471 37255
rect 2436 37029 2471 37095
rect 2595 37029 2629 37258
rect 2753 37143 2787 37267
rect 2884 37138 2902 37172
rect 2936 37138 2952 37172
rect 4315 37170 4557 37178
rect 4315 37136 4523 37170
rect 4315 37130 4557 37136
rect 4591 37170 4661 37178
rect 4591 37136 4615 37170
rect 4649 37136 4661 37170
rect 4591 37131 4661 37136
rect 4591 37130 4657 37131
rect 2753 37029 2787 37092
rect 4914 37096 5204 37336
rect 2913 37038 2956 37058
rect 924 36949 980 36991
rect 1140 36949 1188 36991
rect 924 36861 947 36949
rect 1042 36861 1081 36936
rect 1165 36861 1188 36949
rect 1946 36921 1991 37029
rect 2273 36921 2318 37029
rect 2423 36921 2471 37029
rect 2753 36928 2800 37029
rect 2913 37003 2916 37038
rect 2953 37003 2956 37038
rect 2913 36987 2956 37003
rect 4914 36936 4983 37096
rect 5143 36936 5204 37096
rect 4914 36932 5204 36936
rect 924 36650 1188 36861
rect 2595 36838 2629 36921
rect 2753 36838 2879 36928
rect 4721 36898 5204 36932
rect 2538 36830 2685 36838
rect 2538 36788 2551 36830
rect 2593 36788 2631 36830
rect 2673 36788 2685 36830
rect 2538 36750 2685 36788
rect 2538 36711 2551 36750
rect 2593 36711 2631 36750
rect 2673 36711 2685 36750
rect 2538 36703 2685 36711
rect 2752 36830 2899 36838
rect 2752 36788 2765 36830
rect 2807 36788 2845 36830
rect 2887 36788 2899 36830
rect 2752 36747 2899 36788
rect 2752 36713 2765 36747
rect 2807 36713 2845 36747
rect 2887 36713 2899 36747
rect 2752 36707 2899 36713
rect 4914 36650 5204 36898
rect 924 36614 5204 36650
rect 924 36454 980 36614
rect 1140 36454 1408 36614
rect 1568 36454 1808 36614
rect 1968 36454 2208 36614
rect 2368 36609 3408 36614
rect 2368 36454 2742 36609
rect 924 36449 2742 36454
rect 2902 36449 3069 36609
rect 3229 36454 3408 36609
rect 3568 36454 3808 36614
rect 3968 36454 4208 36614
rect 4368 36454 4608 36614
rect 4768 36454 4983 36614
rect 5143 36454 5204 36614
rect 3229 36449 5204 36454
rect 924 36411 5203 36449
rect 20526 35592 21428 35642
rect 20526 35516 21069 35592
rect 21141 35516 21191 35592
rect 21263 35516 21317 35592
rect 21389 35516 21428 35592
rect 20526 35445 21428 35516
rect 20526 35369 21069 35445
rect 21141 35369 21191 35445
rect 21263 35369 21317 35445
rect 21389 35369 21428 35445
rect 20526 35308 21428 35369
rect 20526 35232 21069 35308
rect 21141 35232 21191 35308
rect 21263 35232 21317 35308
rect 21389 35232 21428 35308
rect 20526 35183 21428 35232
rect 20526 35182 21401 35183
rect 20526 33832 21428 33882
rect 20526 33756 21069 33832
rect 21141 33756 21191 33832
rect 21263 33756 21317 33832
rect 21389 33756 21428 33832
rect 20526 33685 21428 33756
rect 20526 33609 21069 33685
rect 21141 33609 21191 33685
rect 21263 33609 21317 33685
rect 21389 33609 21428 33685
rect 20526 33548 21428 33609
rect 20526 33472 21069 33548
rect 21141 33472 21191 33548
rect 21263 33472 21317 33548
rect 21389 33472 21428 33548
rect 20526 33423 21428 33472
rect 20526 33422 21401 33423
rect 485 31110 847 31111
rect 463 31061 1116 31110
rect 463 30985 504 31061
rect 576 30985 626 31061
rect 698 30985 752 31061
rect 824 30985 1116 31061
rect 463 30914 1116 30985
rect 463 30838 504 30914
rect 576 30838 626 30914
rect 698 30838 752 30914
rect 824 30838 1116 30914
rect 463 30777 1116 30838
rect 463 30701 504 30777
rect 576 30701 626 30777
rect 698 30701 752 30777
rect 824 30701 1116 30777
rect 463 30652 1116 30701
rect 463 30651 946 30652
rect 463 29294 1026 29350
rect 463 29218 504 29294
rect 576 29218 626 29294
rect 698 29218 752 29294
rect 824 29218 1026 29294
rect 463 29147 1026 29218
rect 463 29071 504 29147
rect 576 29071 626 29147
rect 698 29071 752 29147
rect 824 29071 1026 29147
rect 463 29010 1026 29071
rect 463 28934 504 29010
rect 576 28934 626 29010
rect 698 28934 752 29010
rect 824 28934 1026 29010
rect 463 28890 1026 28934
rect 463 27060 946 27109
rect 463 26984 504 27060
rect 576 26984 626 27060
rect 698 26984 752 27060
rect 824 26984 946 27060
rect 463 26913 946 26984
rect 463 26837 504 26913
rect 576 26837 626 26913
rect 698 26837 752 26913
rect 824 26837 946 26913
rect 463 26776 946 26837
rect 463 26700 504 26776
rect 576 26700 626 26776
rect 698 26700 752 26776
rect 824 26700 946 26776
rect 463 26650 946 26700
rect 463 25300 946 25349
rect 463 25224 504 25300
rect 576 25224 626 25300
rect 698 25224 752 25300
rect 824 25224 946 25300
rect 463 25153 946 25224
rect 463 25077 504 25153
rect 576 25077 626 25153
rect 698 25077 752 25153
rect 824 25077 946 25153
rect 463 25016 946 25077
rect 463 24940 504 25016
rect 576 24940 626 25016
rect 698 24940 752 25016
rect 824 24940 946 25016
rect 463 24890 946 24940
rect 463 23060 946 23109
rect 463 22984 504 23060
rect 576 22984 626 23060
rect 698 22984 752 23060
rect 824 22984 946 23060
rect 463 22913 946 22984
rect 463 22837 504 22913
rect 576 22837 626 22913
rect 698 22837 752 22913
rect 824 22837 946 22913
rect 463 22776 946 22837
rect 463 22700 504 22776
rect 576 22700 626 22776
rect 698 22700 752 22776
rect 824 22700 946 22776
rect 463 22650 946 22700
rect 463 21301 946 21350
rect 463 21225 504 21301
rect 576 21225 626 21301
rect 698 21225 752 21301
rect 824 21225 946 21301
rect 463 21154 946 21225
rect 463 21078 504 21154
rect 576 21078 626 21154
rect 698 21078 752 21154
rect 824 21078 946 21154
rect 463 21017 946 21078
rect 463 20941 504 21017
rect 576 20941 626 21017
rect 698 20941 752 21017
rect 824 20941 946 21017
rect 463 20891 946 20941
rect 463 19060 946 19109
rect 463 18984 504 19060
rect 576 18984 626 19060
rect 698 18984 752 19060
rect 824 18984 946 19060
rect 463 18913 946 18984
rect 463 18837 504 18913
rect 576 18837 626 18913
rect 698 18837 752 18913
rect 824 18837 946 18913
rect 463 18776 946 18837
rect 463 18700 504 18776
rect 576 18700 626 18776
rect 698 18700 752 18776
rect 824 18700 946 18776
rect 463 18650 946 18700
rect 463 17300 946 17349
rect 463 17224 504 17300
rect 576 17224 626 17300
rect 698 17224 752 17300
rect 824 17224 946 17300
rect 463 17153 946 17224
rect 463 17077 504 17153
rect 576 17077 626 17153
rect 698 17077 752 17153
rect 824 17077 946 17153
rect 463 17016 946 17077
rect 463 16940 504 17016
rect 576 16940 626 17016
rect 698 16940 752 17016
rect 824 16940 946 17016
rect 463 16890 946 16940
rect 463 15060 946 15109
rect 463 14984 504 15060
rect 576 14984 626 15060
rect 698 14984 752 15060
rect 824 14984 946 15060
rect 463 14913 946 14984
rect 463 14837 504 14913
rect 576 14837 626 14913
rect 698 14837 752 14913
rect 824 14837 946 14913
rect 463 14776 946 14837
rect 463 14700 504 14776
rect 576 14700 626 14776
rect 698 14700 752 14776
rect 824 14700 946 14776
rect 463 14650 946 14700
rect 463 13300 946 13349
rect 463 13224 504 13300
rect 576 13224 626 13300
rect 698 13224 752 13300
rect 824 13224 946 13300
rect 463 13153 946 13224
rect 463 13077 504 13153
rect 576 13077 626 13153
rect 698 13077 752 13153
rect 824 13077 946 13153
rect 463 13016 946 13077
rect 463 12940 504 13016
rect 576 12940 626 13016
rect 698 12940 752 13016
rect 824 12940 946 13016
rect 463 12890 946 12940
rect 463 11061 946 11110
rect 463 10985 504 11061
rect 576 10985 626 11061
rect 698 10985 752 11061
rect 824 10985 946 11061
rect 463 10914 946 10985
rect 463 10838 504 10914
rect 576 10838 626 10914
rect 698 10838 752 10914
rect 824 10838 946 10914
rect 463 10777 946 10838
rect 463 10701 504 10777
rect 576 10701 626 10777
rect 698 10701 752 10777
rect 824 10701 946 10777
rect 463 10651 946 10701
rect 463 9299 946 9348
rect 463 9223 504 9299
rect 576 9223 626 9299
rect 698 9223 752 9299
rect 824 9223 946 9299
rect 463 9152 946 9223
rect 463 9076 504 9152
rect 576 9076 626 9152
rect 698 9076 752 9152
rect 824 9076 946 9152
rect 463 9015 946 9076
rect 463 8939 504 9015
rect 576 8939 626 9015
rect 698 8939 752 9015
rect 824 8939 946 9015
rect 463 8889 946 8939
rect 463 7061 946 7110
rect 463 6985 504 7061
rect 576 6985 626 7061
rect 698 6985 752 7061
rect 824 6985 946 7061
rect 463 6914 946 6985
rect 463 6838 504 6914
rect 576 6838 626 6914
rect 698 6838 752 6914
rect 824 6838 946 6914
rect 463 6777 946 6838
rect 463 6701 504 6777
rect 576 6701 626 6777
rect 698 6701 752 6777
rect 824 6701 946 6777
rect 463 6651 946 6701
rect 463 5300 946 5349
rect 463 5224 504 5300
rect 576 5224 626 5300
rect 698 5224 752 5300
rect 824 5224 946 5300
rect 463 5153 946 5224
rect 463 5077 504 5153
rect 576 5077 626 5153
rect 698 5077 752 5153
rect 824 5077 946 5153
rect 463 5016 946 5077
rect 463 4940 504 5016
rect 576 4940 626 5016
rect 698 4940 752 5016
rect 824 4940 946 5016
rect 463 4890 946 4940
rect 463 3061 946 3110
rect 463 2985 504 3061
rect 576 2985 626 3061
rect 698 2985 752 3061
rect 824 2985 946 3061
rect 463 2914 946 2985
rect 463 2838 504 2914
rect 576 2838 626 2914
rect 698 2838 752 2914
rect 824 2838 946 2914
rect 463 2777 946 2838
rect 463 2701 504 2777
rect 576 2701 626 2777
rect 698 2701 752 2777
rect 824 2701 946 2777
rect 463 2651 946 2701
rect 463 1300 946 1349
rect 463 1224 504 1300
rect 576 1224 626 1300
rect 698 1224 752 1300
rect 824 1224 946 1300
rect 463 1153 946 1224
rect 463 1077 504 1153
rect 576 1077 626 1153
rect 698 1077 752 1153
rect 824 1077 946 1153
rect 463 1016 946 1077
rect 463 940 504 1016
rect 576 940 626 1016
rect 698 940 752 1016
rect 824 940 946 1016
rect 463 890 946 940
<< viali >>
rect 503 75376 575 75452
rect 629 75376 701 75452
rect 749 75376 821 75452
rect 21068 75416 21140 75492
rect 21194 75416 21266 75492
rect 21314 75416 21386 75492
rect 503 75258 575 75334
rect 629 75258 701 75334
rect 749 75258 821 75334
rect 21068 75298 21140 75374
rect 21194 75298 21266 75374
rect 21314 75298 21386 75374
rect 504 74984 576 75060
rect 626 74984 698 75060
rect 752 74984 824 75060
rect 504 74837 576 74913
rect 626 74837 698 74913
rect 752 74837 824 74913
rect 504 74700 576 74776
rect 626 74700 698 74776
rect 752 74700 824 74776
rect 22010 73995 22082 74071
rect 22136 73995 22208 74071
rect 22256 73995 22328 74071
rect 22010 73877 22082 73953
rect 22136 73877 22208 73953
rect 22256 73877 22328 73953
rect 504 73224 576 73300
rect 626 73224 698 73300
rect 752 73224 824 73300
rect 504 73077 576 73153
rect 626 73077 698 73153
rect 752 73077 824 73153
rect 504 72940 576 73016
rect 626 72940 698 73016
rect 752 72940 824 73016
rect 503 72703 575 72779
rect 629 72703 701 72779
rect 749 72703 821 72779
rect 503 72585 575 72661
rect 629 72585 701 72661
rect 749 72585 821 72661
rect 21068 72619 21140 72695
rect 21194 72619 21266 72695
rect 21314 72619 21386 72695
rect 21068 72501 21140 72577
rect 21194 72501 21266 72577
rect 21314 72501 21386 72577
rect 503 71376 575 71452
rect 629 71376 701 71452
rect 749 71376 821 71452
rect 21068 71416 21140 71492
rect 21194 71416 21266 71492
rect 21314 71416 21386 71492
rect 503 71258 575 71334
rect 629 71258 701 71334
rect 749 71258 821 71334
rect 21068 71298 21140 71374
rect 21194 71298 21266 71374
rect 21314 71298 21386 71374
rect 504 70984 576 71060
rect 626 70984 698 71060
rect 752 70984 824 71060
rect 504 70837 576 70913
rect 626 70837 698 70913
rect 752 70837 824 70913
rect 504 70700 576 70776
rect 626 70700 698 70776
rect 752 70700 824 70776
rect 22010 69995 22082 70071
rect 22136 69995 22208 70071
rect 22256 69995 22328 70071
rect 22010 69877 22082 69953
rect 22136 69877 22208 69953
rect 22256 69877 22328 69953
rect 504 69224 576 69300
rect 626 69224 698 69300
rect 752 69224 824 69300
rect 504 69077 576 69153
rect 626 69077 698 69153
rect 752 69077 824 69153
rect 504 68940 576 69016
rect 626 68940 698 69016
rect 752 68940 824 69016
rect 503 68703 575 68779
rect 629 68703 701 68779
rect 749 68703 821 68779
rect 503 68585 575 68661
rect 629 68585 701 68661
rect 749 68585 821 68661
rect 21068 68619 21140 68695
rect 21194 68619 21266 68695
rect 21314 68619 21386 68695
rect 21068 68501 21140 68577
rect 21194 68501 21266 68577
rect 21314 68501 21386 68577
rect 503 67374 575 67450
rect 629 67374 701 67450
rect 749 67374 821 67450
rect 21068 67416 21140 67492
rect 21194 67416 21266 67492
rect 21314 67416 21386 67492
rect 503 67256 575 67332
rect 629 67256 701 67332
rect 749 67256 821 67332
rect 21068 67298 21140 67374
rect 21194 67298 21266 67374
rect 21314 67298 21386 67374
rect 504 66984 576 67060
rect 626 66984 698 67060
rect 752 66984 824 67060
rect 504 66837 576 66913
rect 626 66837 698 66913
rect 752 66837 824 66913
rect 504 66700 576 66776
rect 626 66700 698 66776
rect 752 66700 824 66776
rect 22010 65982 22082 66058
rect 22136 65982 22208 66058
rect 22256 65982 22328 66058
rect 22010 65864 22082 65940
rect 22136 65864 22208 65940
rect 22256 65864 22328 65940
rect 504 65225 576 65301
rect 626 65225 698 65301
rect 752 65225 824 65301
rect 504 65078 576 65154
rect 626 65078 698 65154
rect 752 65078 824 65154
rect 504 64941 576 65017
rect 626 64941 698 65017
rect 752 64941 824 65017
rect 503 64634 575 64710
rect 629 64634 701 64710
rect 749 64634 821 64710
rect 21068 64619 21140 64695
rect 21194 64619 21266 64695
rect 21314 64619 21386 64695
rect 503 64516 575 64592
rect 629 64516 701 64592
rect 749 64516 821 64592
rect 21068 64501 21140 64577
rect 21194 64501 21266 64577
rect 21314 64501 21386 64577
rect 503 63456 575 63532
rect 629 63456 701 63532
rect 749 63456 821 63532
rect 21068 63416 21140 63492
rect 21194 63416 21266 63492
rect 21314 63416 21386 63492
rect 503 63338 575 63414
rect 629 63338 701 63414
rect 749 63338 821 63414
rect 21068 63298 21140 63374
rect 21194 63298 21266 63374
rect 21314 63298 21386 63374
rect 504 62984 576 63060
rect 626 62984 698 63060
rect 752 62984 824 63060
rect 504 62837 576 62913
rect 626 62837 698 62913
rect 752 62837 824 62913
rect 504 62700 576 62776
rect 626 62700 698 62776
rect 752 62700 824 62776
rect 22010 61981 22082 62057
rect 22136 61981 22208 62057
rect 22256 61981 22328 62057
rect 22010 61863 22082 61939
rect 22136 61863 22208 61939
rect 22256 61863 22328 61939
rect 504 61225 576 61301
rect 626 61225 698 61301
rect 752 61225 824 61301
rect 504 61078 576 61154
rect 626 61078 698 61154
rect 752 61078 824 61154
rect 504 60941 576 61017
rect 626 60941 698 61017
rect 752 60941 824 61017
rect 503 60608 575 60684
rect 629 60608 701 60684
rect 749 60608 821 60684
rect 21068 60619 21140 60695
rect 21194 60619 21266 60695
rect 21314 60619 21386 60695
rect 503 60490 575 60566
rect 629 60490 701 60566
rect 749 60490 821 60566
rect 21068 60501 21140 60577
rect 21194 60501 21266 60577
rect 21314 60501 21386 60577
rect 503 59405 575 59481
rect 629 59405 701 59481
rect 749 59405 821 59481
rect 21068 59470 21140 59546
rect 21194 59470 21266 59546
rect 21314 59470 21386 59546
rect 503 59287 575 59363
rect 629 59287 701 59363
rect 749 59287 821 59363
rect 21068 59352 21140 59428
rect 21194 59352 21266 59428
rect 21314 59352 21386 59428
rect 504 58984 576 59060
rect 626 58984 698 59060
rect 752 58984 824 59060
rect 504 58837 576 58913
rect 626 58837 698 58913
rect 752 58837 824 58913
rect 504 58700 576 58776
rect 626 58700 698 58776
rect 752 58700 824 58776
rect 22010 58020 22082 58096
rect 22136 58020 22208 58096
rect 22256 58020 22328 58096
rect 22010 57902 22082 57978
rect 22136 57902 22208 57978
rect 22256 57902 22328 57978
rect 504 57223 576 57299
rect 626 57223 698 57299
rect 752 57223 824 57299
rect 504 57076 576 57152
rect 626 57076 698 57152
rect 752 57076 824 57152
rect 504 56939 576 57015
rect 626 56939 698 57015
rect 752 56939 824 57015
rect 503 56628 575 56704
rect 629 56628 701 56704
rect 749 56628 821 56704
rect 503 56510 575 56586
rect 629 56510 701 56586
rect 749 56510 821 56586
rect 21068 56554 21140 56630
rect 21194 56554 21266 56630
rect 21314 56554 21386 56630
rect 21068 56436 21140 56512
rect 21194 56436 21266 56512
rect 21314 56436 21386 56512
rect 503 55421 575 55497
rect 629 55421 701 55497
rect 749 55421 821 55497
rect 503 55303 575 55379
rect 629 55303 701 55379
rect 749 55303 821 55379
rect 21068 55371 21140 55447
rect 21194 55371 21266 55447
rect 21314 55371 21386 55447
rect 21068 55253 21140 55329
rect 21194 55253 21266 55329
rect 21314 55253 21386 55329
rect 504 54984 576 55060
rect 626 54984 698 55060
rect 752 54984 824 55060
rect 504 54837 576 54913
rect 626 54837 698 54913
rect 752 54837 824 54913
rect 504 54700 576 54776
rect 626 54700 698 54776
rect 752 54700 824 54776
rect 22010 54003 22082 54079
rect 22136 54003 22208 54079
rect 22256 54003 22328 54079
rect 22010 53885 22082 53961
rect 22136 53885 22208 53961
rect 22256 53885 22328 53961
rect 504 53225 576 53301
rect 626 53225 698 53301
rect 752 53225 824 53301
rect 504 53078 576 53154
rect 626 53078 698 53154
rect 752 53078 824 53154
rect 504 52941 576 53017
rect 626 52941 698 53017
rect 752 52941 824 53017
rect 503 52655 575 52731
rect 629 52655 701 52731
rect 749 52655 821 52731
rect 503 52537 575 52613
rect 629 52537 701 52613
rect 749 52537 821 52613
rect 21068 52499 21140 52575
rect 21194 52499 21266 52575
rect 21314 52499 21386 52575
rect 21068 52381 21140 52457
rect 21194 52381 21266 52457
rect 21314 52381 21386 52457
rect 503 51468 575 51544
rect 629 51468 701 51544
rect 749 51468 821 51544
rect 503 51350 575 51426
rect 629 51350 701 51426
rect 749 51350 821 51426
rect 21068 51364 21140 51440
rect 21194 51364 21266 51440
rect 21314 51364 21386 51440
rect 21068 51246 21140 51322
rect 21194 51246 21266 51322
rect 21314 51246 21386 51322
rect 504 50984 576 51060
rect 626 50984 698 51060
rect 752 50984 824 51060
rect 504 50837 576 50913
rect 626 50837 698 50913
rect 752 50837 824 50913
rect 504 50700 576 50776
rect 626 50700 698 50776
rect 752 50700 824 50776
rect 22010 50082 22082 50158
rect 22136 50082 22208 50158
rect 22256 50082 22328 50158
rect 22010 49964 22082 50040
rect 22136 49964 22208 50040
rect 22256 49964 22328 50040
rect 504 49225 576 49301
rect 626 49225 698 49301
rect 752 49225 824 49301
rect 504 49078 576 49154
rect 626 49078 698 49154
rect 752 49078 824 49154
rect 504 48941 576 49017
rect 626 48941 698 49017
rect 752 48941 824 49017
rect 503 48646 575 48722
rect 629 48646 701 48722
rect 749 48646 821 48722
rect 21068 48605 21140 48681
rect 21194 48605 21266 48681
rect 21314 48605 21386 48681
rect 503 48528 575 48604
rect 629 48528 701 48604
rect 749 48528 821 48604
rect 21068 48487 21140 48563
rect 21194 48487 21266 48563
rect 21314 48487 21386 48563
rect 503 47493 575 47569
rect 629 47493 701 47569
rect 749 47493 821 47569
rect 21068 47452 21140 47528
rect 21194 47452 21266 47528
rect 21314 47452 21386 47528
rect 503 47375 575 47451
rect 629 47375 701 47451
rect 749 47375 821 47451
rect 21068 47334 21140 47410
rect 21194 47334 21266 47410
rect 21314 47334 21386 47410
rect 504 46984 576 47060
rect 626 46984 698 47060
rect 752 46984 824 47060
rect 504 46837 576 46913
rect 626 46837 698 46913
rect 752 46837 824 46913
rect 504 46700 576 46776
rect 626 46700 698 46776
rect 752 46700 824 46776
rect 22010 45824 22082 45900
rect 22136 45824 22208 45900
rect 22256 45824 22328 45900
rect 22010 45706 22082 45782
rect 22136 45706 22208 45782
rect 22256 45706 22328 45782
rect 504 45224 576 45300
rect 626 45224 698 45300
rect 752 45224 824 45300
rect 504 45077 576 45153
rect 626 45077 698 45153
rect 752 45077 824 45153
rect 504 44940 576 45016
rect 626 44940 698 45016
rect 752 44940 824 45016
rect 503 44433 575 44509
rect 629 44433 701 44509
rect 749 44433 821 44509
rect 503 44315 575 44391
rect 629 44315 701 44391
rect 749 44315 821 44391
rect 21068 44336 21140 44412
rect 21194 44336 21266 44412
rect 21314 44336 21386 44412
rect 21068 44218 21140 44294
rect 21194 44218 21266 44294
rect 21314 44218 21386 44294
rect 1662 39279 1704 39321
rect 1742 39279 1784 39321
rect 1885 39281 2003 39395
rect 2041 39281 2159 39395
rect 2197 39281 2315 39395
rect 1662 39199 1704 39241
rect 1742 39199 1784 39241
rect 2192 39191 2227 39230
rect 941 39096 1013 39137
rect 1098 39096 1165 39138
rect 941 39062 980 39096
rect 980 39062 1013 39096
rect 1098 39063 1140 39096
rect 1140 39063 1165 39096
rect 1604 39059 1638 39125
rect 944 38946 980 39021
rect 980 38946 1016 39021
rect 1098 38949 1140 39024
rect 1140 38949 1165 39024
rect 1920 39069 1954 39124
rect 2551 39286 2593 39328
rect 2631 39286 2673 39328
rect 2551 39206 2593 39248
rect 2631 39206 2673 39248
rect 1604 38889 1638 38944
rect 1920 38889 1954 38944
rect 2035 38889 2069 38944
rect 2351 38889 2385 38944
rect 2479 38889 2514 38949
rect 2797 38890 2831 38949
rect 2901 38947 2935 38981
rect 4251 38926 4285 38960
rect 2921 38836 2955 38870
rect 3253 38836 3288 38870
rect 3553 38836 3587 38870
rect 4105 38836 4139 38870
rect 4339 38836 4373 38870
rect 4615 38836 4650 38871
rect 1762 38706 1796 38782
rect 3800 38779 3835 38813
rect 1479 38225 1515 38260
rect 1715 38224 1749 38258
rect 1807 38227 1841 38261
rect 1899 38224 1933 38258
rect 2029 38218 2063 38252
rect 4662 38224 4696 38258
rect 1481 37748 1515 37782
rect 1805 37753 1839 37787
rect 1889 37754 1923 37788
rect 1986 37748 2020 37782
rect 4662 37748 4696 37782
rect 1686 37310 1732 37358
rect 1686 37200 1732 37245
rect 947 36991 980 37079
rect 980 36991 1042 37079
rect 1080 36991 1140 37079
rect 1140 36991 1165 37079
rect 1957 37090 1991 37144
rect 2273 37089 2307 37143
rect 2436 37095 2471 37146
rect 3807 37193 3841 37227
rect 2753 37092 2787 37143
rect 2902 37138 2936 37172
rect 3237 37137 3271 37171
rect 3553 37136 3587 37170
rect 4105 37136 4139 37170
rect 4523 37136 4557 37170
rect 4615 37136 4649 37170
rect 4251 37046 4285 37080
rect 947 36936 980 36949
rect 980 36936 1042 36949
rect 1081 36936 1140 36949
rect 1140 36936 1165 36949
rect 947 36861 1042 36936
rect 1081 36861 1165 36936
rect 2916 37003 2953 37038
rect 2551 36788 2593 36830
rect 2631 36788 2673 36830
rect 2551 36711 2593 36750
rect 2631 36711 2673 36750
rect 2765 36788 2807 36830
rect 2845 36788 2887 36830
rect 2765 36713 2807 36747
rect 2845 36713 2887 36747
rect 21069 35516 21141 35592
rect 21191 35516 21263 35592
rect 21317 35516 21389 35592
rect 21069 35369 21141 35445
rect 21191 35369 21263 35445
rect 21317 35369 21389 35445
rect 21069 35232 21141 35308
rect 21191 35232 21263 35308
rect 21317 35232 21389 35308
rect 21069 33756 21141 33832
rect 21191 33756 21263 33832
rect 21317 33756 21389 33832
rect 21069 33609 21141 33685
rect 21191 33609 21263 33685
rect 21317 33609 21389 33685
rect 21069 33472 21141 33548
rect 21191 33472 21263 33548
rect 21317 33472 21389 33548
rect 503 32226 575 32302
rect 629 32226 701 32302
rect 749 32226 821 32302
rect 21068 32226 21140 32302
rect 21194 32226 21266 32302
rect 21314 32226 21386 32302
rect 503 32108 575 32184
rect 629 32108 701 32184
rect 749 32108 821 32184
rect 21068 32108 21140 32184
rect 21194 32108 21266 32184
rect 21314 32108 21386 32184
rect 503 31444 575 31520
rect 629 31444 701 31520
rect 749 31444 821 31520
rect 21068 31444 21140 31520
rect 21194 31444 21266 31520
rect 21314 31444 21386 31520
rect 503 31326 575 31402
rect 629 31326 701 31402
rect 749 31326 821 31402
rect 21068 31326 21140 31402
rect 21194 31326 21266 31402
rect 21314 31326 21386 31402
rect 504 30985 576 31061
rect 626 30985 698 31061
rect 752 30985 824 31061
rect 504 30838 576 30914
rect 626 30838 698 30914
rect 752 30838 824 30914
rect 504 30701 576 30777
rect 626 30701 698 30777
rect 752 30701 824 30777
rect 22010 30054 22082 30130
rect 22136 30054 22208 30130
rect 22256 30054 22328 30130
rect 22010 29936 22082 30012
rect 22136 29936 22208 30012
rect 22256 29936 22328 30012
rect 504 29218 576 29294
rect 626 29218 698 29294
rect 752 29218 824 29294
rect 504 29071 576 29147
rect 626 29071 698 29147
rect 752 29071 824 29147
rect 504 28934 576 29010
rect 626 28934 698 29010
rect 752 28934 824 29010
rect 503 28532 575 28608
rect 629 28532 701 28608
rect 749 28532 821 28608
rect 503 28414 575 28490
rect 629 28414 701 28490
rect 749 28414 821 28490
rect 21068 28483 21140 28559
rect 21194 28483 21266 28559
rect 21314 28483 21386 28559
rect 21068 28365 21140 28441
rect 21194 28365 21266 28441
rect 21314 28365 21386 28441
rect 503 27528 575 27604
rect 629 27528 701 27604
rect 749 27528 821 27604
rect 503 27410 575 27486
rect 629 27410 701 27486
rect 749 27410 821 27486
rect 21068 27366 21140 27442
rect 21194 27366 21266 27442
rect 21314 27366 21386 27442
rect 21068 27248 21140 27324
rect 21194 27248 21266 27324
rect 21314 27248 21386 27324
rect 504 26984 576 27060
rect 626 26984 698 27060
rect 752 26984 824 27060
rect 504 26837 576 26913
rect 626 26837 698 26913
rect 752 26837 824 26913
rect 504 26700 576 26776
rect 626 26700 698 26776
rect 752 26700 824 26776
rect 22010 25895 22082 25971
rect 22136 25895 22208 25971
rect 22256 25895 22328 25971
rect 22010 25777 22082 25853
rect 22136 25777 22208 25853
rect 22256 25777 22328 25853
rect 504 25224 576 25300
rect 626 25224 698 25300
rect 752 25224 824 25300
rect 504 25077 576 25153
rect 626 25077 698 25153
rect 752 25077 824 25153
rect 504 24940 576 25016
rect 626 24940 698 25016
rect 752 24940 824 25016
rect 503 24550 575 24626
rect 629 24550 701 24626
rect 749 24550 821 24626
rect 21068 24523 21140 24599
rect 21194 24523 21266 24599
rect 21314 24523 21386 24599
rect 503 24432 575 24508
rect 629 24432 701 24508
rect 749 24432 821 24508
rect 21068 24405 21140 24481
rect 21194 24405 21266 24481
rect 21314 24405 21386 24481
rect 503 23468 575 23544
rect 629 23468 701 23544
rect 749 23468 821 23544
rect 503 23350 575 23426
rect 629 23350 701 23426
rect 749 23350 821 23426
rect 21068 23348 21140 23424
rect 21194 23348 21266 23424
rect 21314 23348 21386 23424
rect 21068 23230 21140 23306
rect 21194 23230 21266 23306
rect 21314 23230 21386 23306
rect 504 22984 576 23060
rect 626 22984 698 23060
rect 752 22984 824 23060
rect 504 22837 576 22913
rect 626 22837 698 22913
rect 752 22837 824 22913
rect 504 22700 576 22776
rect 626 22700 698 22776
rect 752 22700 824 22776
rect 22010 22105 22082 22181
rect 22136 22105 22208 22181
rect 22256 22105 22328 22181
rect 22010 21987 22082 22063
rect 22136 21987 22208 22063
rect 22256 21987 22328 22063
rect 504 21225 576 21301
rect 626 21225 698 21301
rect 752 21225 824 21301
rect 504 21078 576 21154
rect 626 21078 698 21154
rect 752 21078 824 21154
rect 504 20941 576 21017
rect 626 20941 698 21017
rect 752 20941 824 21017
rect 503 20593 575 20669
rect 629 20593 701 20669
rect 749 20593 821 20669
rect 503 20475 575 20551
rect 629 20475 701 20551
rect 749 20475 821 20551
rect 21068 20507 21140 20583
rect 21194 20507 21266 20583
rect 21314 20507 21386 20583
rect 21068 20389 21140 20465
rect 21194 20389 21266 20465
rect 21314 20389 21386 20465
rect 503 19492 575 19568
rect 629 19492 701 19568
rect 749 19492 821 19568
rect 503 19374 575 19450
rect 629 19374 701 19450
rect 749 19374 821 19450
rect 21068 19336 21140 19412
rect 21194 19336 21266 19412
rect 21314 19336 21386 19412
rect 21068 19218 21140 19294
rect 21194 19218 21266 19294
rect 21314 19218 21386 19294
rect 504 18984 576 19060
rect 626 18984 698 19060
rect 752 18984 824 19060
rect 504 18837 576 18913
rect 626 18837 698 18913
rect 752 18837 824 18913
rect 504 18700 576 18776
rect 626 18700 698 18776
rect 752 18700 824 18776
rect 22010 17998 22082 18074
rect 22136 17998 22208 18074
rect 22256 17998 22328 18074
rect 22010 17880 22082 17956
rect 22136 17880 22208 17956
rect 22256 17880 22328 17956
rect 504 17224 576 17300
rect 626 17224 698 17300
rect 752 17224 824 17300
rect 504 17077 576 17153
rect 626 17077 698 17153
rect 752 17077 824 17153
rect 504 16940 576 17016
rect 626 16940 698 17016
rect 752 16940 824 17016
rect 503 16626 575 16702
rect 629 16626 701 16702
rect 749 16626 821 16702
rect 503 16508 575 16584
rect 629 16508 701 16584
rect 749 16508 821 16584
rect 21068 16575 21140 16651
rect 21194 16575 21266 16651
rect 21314 16575 21386 16651
rect 21068 16457 21140 16533
rect 21194 16457 21266 16533
rect 21314 16457 21386 16533
rect 503 15410 575 15486
rect 629 15410 701 15486
rect 749 15410 821 15486
rect 503 15292 575 15368
rect 629 15292 701 15368
rect 749 15292 821 15368
rect 21068 15361 21140 15437
rect 21194 15361 21266 15437
rect 21314 15361 21386 15437
rect 21068 15243 21140 15319
rect 21194 15243 21266 15319
rect 21314 15243 21386 15319
rect 504 14984 576 15060
rect 626 14984 698 15060
rect 752 14984 824 15060
rect 504 14837 576 14913
rect 626 14837 698 14913
rect 752 14837 824 14913
rect 504 14700 576 14776
rect 626 14700 698 14776
rect 752 14700 824 14776
rect 22010 14180 22082 14256
rect 22136 14180 22208 14256
rect 22256 14180 22328 14256
rect 22010 14062 22082 14138
rect 22136 14062 22208 14138
rect 22256 14062 22328 14138
rect 504 13224 576 13300
rect 626 13224 698 13300
rect 752 13224 824 13300
rect 504 13077 576 13153
rect 626 13077 698 13153
rect 752 13077 824 13153
rect 504 12940 576 13016
rect 626 12940 698 13016
rect 752 12940 824 13016
rect 503 12545 575 12621
rect 629 12545 701 12621
rect 749 12545 821 12621
rect 21068 12518 21140 12594
rect 21194 12518 21266 12594
rect 21314 12518 21386 12594
rect 503 12427 575 12503
rect 629 12427 701 12503
rect 749 12427 821 12503
rect 21068 12400 21140 12476
rect 21194 12400 21266 12476
rect 21314 12400 21386 12476
rect 503 11423 575 11499
rect 629 11423 701 11499
rect 749 11423 821 11499
rect 503 11305 575 11381
rect 629 11305 701 11381
rect 749 11305 821 11381
rect 21068 11361 21140 11437
rect 21194 11361 21266 11437
rect 21314 11361 21386 11437
rect 21068 11243 21140 11319
rect 21194 11243 21266 11319
rect 21314 11243 21386 11319
rect 504 10985 576 11061
rect 626 10985 698 11061
rect 752 10985 824 11061
rect 504 10838 576 10914
rect 626 10838 698 10914
rect 752 10838 824 10914
rect 504 10701 576 10777
rect 626 10701 698 10777
rect 752 10701 824 10777
rect 22010 10216 22082 10292
rect 22136 10216 22208 10292
rect 22256 10216 22328 10292
rect 22010 10098 22082 10174
rect 22136 10098 22208 10174
rect 22256 10098 22328 10174
rect 504 9223 576 9299
rect 626 9223 698 9299
rect 752 9223 824 9299
rect 504 9076 576 9152
rect 626 9076 698 9152
rect 752 9076 824 9152
rect 504 8939 576 9015
rect 626 8939 698 9015
rect 752 8939 824 9015
rect 503 8563 575 8639
rect 629 8563 701 8639
rect 749 8563 821 8639
rect 503 8445 575 8521
rect 629 8445 701 8521
rect 749 8445 821 8521
rect 21068 8518 21140 8594
rect 21194 8518 21266 8594
rect 21314 8518 21386 8594
rect 21068 8400 21140 8476
rect 21194 8400 21266 8476
rect 21314 8400 21386 8476
rect 503 7452 575 7528
rect 629 7452 701 7528
rect 749 7452 821 7528
rect 503 7334 575 7410
rect 629 7334 701 7410
rect 749 7334 821 7410
rect 21068 7361 21140 7437
rect 21194 7361 21266 7437
rect 21314 7361 21386 7437
rect 21068 7243 21140 7319
rect 21194 7243 21266 7319
rect 21314 7243 21386 7319
rect 504 6985 576 7061
rect 626 6985 698 7061
rect 752 6985 824 7061
rect 504 6838 576 6914
rect 626 6838 698 6914
rect 752 6838 824 6914
rect 504 6701 576 6777
rect 626 6701 698 6777
rect 752 6701 824 6777
rect 22010 6204 22082 6280
rect 22136 6204 22208 6280
rect 22256 6204 22328 6280
rect 22010 6086 22082 6162
rect 22136 6086 22208 6162
rect 22256 6086 22328 6162
rect 504 5224 576 5300
rect 626 5224 698 5300
rect 752 5224 824 5300
rect 504 5077 576 5153
rect 626 5077 698 5153
rect 752 5077 824 5153
rect 504 4940 576 5016
rect 626 4940 698 5016
rect 752 4940 824 5016
rect 503 4629 575 4705
rect 629 4629 701 4705
rect 749 4629 821 4705
rect 503 4511 575 4587
rect 629 4511 701 4587
rect 749 4511 821 4587
rect 21068 4518 21140 4594
rect 21194 4518 21266 4594
rect 21314 4518 21386 4594
rect 21068 4400 21140 4476
rect 21194 4400 21266 4476
rect 21314 4400 21386 4476
rect 503 3452 575 3528
rect 629 3452 701 3528
rect 749 3452 821 3528
rect 503 3334 575 3410
rect 629 3334 701 3410
rect 749 3334 821 3410
rect 21068 3361 21140 3437
rect 21194 3361 21266 3437
rect 21314 3361 21386 3437
rect 21068 3243 21140 3319
rect 21194 3243 21266 3319
rect 21314 3243 21386 3319
rect 504 2985 576 3061
rect 626 2985 698 3061
rect 752 2985 824 3061
rect 504 2838 576 2914
rect 626 2838 698 2914
rect 752 2838 824 2914
rect 504 2701 576 2777
rect 626 2701 698 2777
rect 752 2701 824 2777
rect 22010 2204 22082 2280
rect 22136 2204 22208 2280
rect 22256 2204 22328 2280
rect 22010 2086 22082 2162
rect 22136 2086 22208 2162
rect 22256 2086 22328 2162
rect 504 1224 576 1300
rect 626 1224 698 1300
rect 752 1224 824 1300
rect 504 1077 576 1153
rect 626 1077 698 1153
rect 752 1077 824 1153
rect 504 940 576 1016
rect 626 940 698 1016
rect 752 940 824 1016
rect 503 629 575 705
rect 629 629 701 705
rect 749 629 821 705
rect 503 511 575 587
rect 629 511 701 587
rect 749 511 821 587
rect 21068 518 21140 594
rect 21194 518 21266 594
rect 21314 518 21386 594
rect 21068 400 21140 476
rect 21194 400 21266 476
rect 21314 400 21386 476
<< metal1 >>
rect 20946 75492 21426 75517
rect 463 75452 946 75477
rect 463 75376 503 75452
rect 575 75376 629 75452
rect 701 75376 749 75452
rect 821 75376 946 75452
rect 463 75334 946 75376
rect 463 75258 503 75334
rect 575 75258 629 75334
rect 701 75258 749 75334
rect 821 75258 946 75334
rect 20946 75416 21068 75492
rect 21140 75416 21194 75492
rect 21266 75416 21314 75492
rect 21386 75416 21426 75492
rect 20946 75374 21426 75416
rect 20946 75298 21068 75374
rect 21140 75298 21194 75374
rect 21266 75298 21314 75374
rect 21386 75298 21426 75374
rect 20946 75262 21426 75298
rect 463 75222 946 75258
rect 463 75060 863 75109
rect 463 74984 504 75060
rect 576 74984 626 75060
rect 698 74984 752 75060
rect 824 74984 863 75060
rect 463 74913 863 74984
rect 463 74837 504 74913
rect 576 74837 626 74913
rect 698 74837 752 74913
rect 824 74837 863 74913
rect 463 74776 863 74837
rect 463 74700 504 74776
rect 576 74700 626 74776
rect 698 74700 752 74776
rect 824 74700 863 74776
rect 463 74650 863 74700
rect 20946 74071 22370 74096
rect 20946 73995 22010 74071
rect 22082 73995 22136 74071
rect 22208 73995 22256 74071
rect 22328 73995 22370 74071
rect 20946 73953 22370 73995
rect 20946 73877 22010 73953
rect 22082 73877 22136 73953
rect 22208 73877 22256 73953
rect 22328 73877 22370 73953
rect 20946 73841 22370 73877
rect 463 73300 863 73349
rect 463 73224 504 73300
rect 576 73224 626 73300
rect 698 73224 752 73300
rect 824 73224 863 73300
rect 463 73153 863 73224
rect 463 73077 504 73153
rect 576 73077 626 73153
rect 698 73077 752 73153
rect 824 73077 863 73153
rect 463 73016 863 73077
rect 463 72940 504 73016
rect 576 72940 626 73016
rect 698 72940 752 73016
rect 824 72940 863 73016
rect 463 72890 863 72940
rect 463 72779 946 72804
rect 463 72703 503 72779
rect 575 72703 629 72779
rect 701 72703 749 72779
rect 821 72703 946 72779
rect 463 72661 946 72703
rect 463 72585 503 72661
rect 575 72585 629 72661
rect 701 72585 749 72661
rect 821 72585 946 72661
rect 463 72549 946 72585
rect 20946 72695 21428 72720
rect 20946 72619 21068 72695
rect 21140 72619 21194 72695
rect 21266 72619 21314 72695
rect 21386 72619 21428 72695
rect 20946 72577 21428 72619
rect 20946 72501 21068 72577
rect 21140 72501 21194 72577
rect 21266 72501 21314 72577
rect 21386 72501 21428 72577
rect 20946 72465 21428 72501
rect 20946 71492 21426 71517
rect 463 71452 947 71477
rect 463 71376 503 71452
rect 575 71376 629 71452
rect 701 71376 749 71452
rect 821 71376 947 71452
rect 463 71334 947 71376
rect 463 71258 503 71334
rect 575 71258 629 71334
rect 701 71258 749 71334
rect 821 71258 947 71334
rect 20946 71416 21068 71492
rect 21140 71416 21194 71492
rect 21266 71416 21314 71492
rect 21386 71416 21426 71492
rect 20946 71374 21426 71416
rect 20946 71298 21068 71374
rect 21140 71298 21194 71374
rect 21266 71298 21314 71374
rect 21386 71298 21426 71374
rect 20946 71262 21426 71298
rect 463 71222 947 71258
rect 463 71060 863 71109
rect 463 70984 504 71060
rect 576 70984 626 71060
rect 698 70984 752 71060
rect 824 70984 863 71060
rect 463 70913 863 70984
rect 463 70837 504 70913
rect 576 70837 626 70913
rect 698 70837 752 70913
rect 824 70837 863 70913
rect 463 70776 863 70837
rect 463 70700 504 70776
rect 576 70700 626 70776
rect 698 70700 752 70776
rect 824 70700 863 70776
rect 463 70650 863 70700
rect 20946 70071 22370 70096
rect 20946 69995 22010 70071
rect 22082 69995 22136 70071
rect 22208 69995 22256 70071
rect 22328 69995 22370 70071
rect 20946 69953 22370 69995
rect 20946 69877 22010 69953
rect 22082 69877 22136 69953
rect 22208 69877 22256 69953
rect 22328 69877 22370 69953
rect 20946 69841 22370 69877
rect 463 69300 863 69349
rect 463 69224 504 69300
rect 576 69224 626 69300
rect 698 69224 752 69300
rect 824 69224 863 69300
rect 463 69153 863 69224
rect 463 69077 504 69153
rect 576 69077 626 69153
rect 698 69077 752 69153
rect 824 69077 863 69153
rect 463 69016 863 69077
rect 463 68940 504 69016
rect 576 68940 626 69016
rect 698 68940 752 69016
rect 824 68940 863 69016
rect 463 68890 863 68940
rect 463 68779 947 68804
rect 463 68703 503 68779
rect 575 68703 629 68779
rect 701 68703 749 68779
rect 821 68703 947 68779
rect 463 68661 947 68703
rect 463 68585 503 68661
rect 575 68585 629 68661
rect 701 68585 749 68661
rect 821 68585 947 68661
rect 463 68549 947 68585
rect 20946 68695 21428 68720
rect 20946 68619 21068 68695
rect 21140 68619 21194 68695
rect 21266 68619 21314 68695
rect 21386 68619 21428 68695
rect 20946 68577 21428 68619
rect 20946 68501 21068 68577
rect 21140 68501 21194 68577
rect 21266 68501 21314 68577
rect 21386 68501 21428 68577
rect 20946 68465 21428 68501
rect 20945 67517 20946 67530
rect 20945 67492 21426 67517
rect 463 67450 947 67475
rect 463 67374 503 67450
rect 575 67374 629 67450
rect 701 67374 749 67450
rect 821 67374 947 67450
rect 463 67332 947 67374
rect 463 67256 503 67332
rect 575 67256 629 67332
rect 701 67256 749 67332
rect 821 67256 947 67332
rect 20945 67416 21068 67492
rect 21140 67416 21194 67492
rect 21266 67416 21314 67492
rect 21386 67416 21426 67492
rect 20945 67374 21426 67416
rect 20945 67298 21068 67374
rect 21140 67298 21194 67374
rect 21266 67298 21314 67374
rect 21386 67298 21426 67374
rect 20945 67275 21426 67298
rect 20946 67262 21426 67275
rect 463 67220 947 67256
rect 463 67060 863 67109
rect 463 66984 504 67060
rect 576 66984 626 67060
rect 698 66984 752 67060
rect 824 66984 863 67060
rect 463 66913 863 66984
rect 463 66837 504 66913
rect 576 66837 626 66913
rect 698 66837 752 66913
rect 824 66837 863 66913
rect 463 66776 863 66837
rect 463 66700 504 66776
rect 576 66700 626 66776
rect 698 66700 752 66776
rect 824 66700 863 66776
rect 463 66650 863 66700
rect 20946 66058 22370 66083
rect 20946 65982 22010 66058
rect 22082 65982 22136 66058
rect 22208 65982 22256 66058
rect 22328 65982 22370 66058
rect 20946 65940 22370 65982
rect 20946 65864 22010 65940
rect 22082 65864 22136 65940
rect 22208 65864 22256 65940
rect 22328 65864 22370 65940
rect 20946 65828 22370 65864
rect 463 65301 863 65350
rect 463 65225 504 65301
rect 576 65225 626 65301
rect 698 65225 752 65301
rect 824 65225 863 65301
rect 463 65154 863 65225
rect 463 65078 504 65154
rect 576 65078 626 65154
rect 698 65078 752 65154
rect 824 65078 863 65154
rect 463 65017 863 65078
rect 463 64941 504 65017
rect 576 64941 626 65017
rect 698 64941 752 65017
rect 824 64941 863 65017
rect 463 64891 863 64941
rect 463 64710 947 64735
rect 463 64634 503 64710
rect 575 64634 629 64710
rect 701 64634 749 64710
rect 821 64634 947 64710
rect 463 64592 947 64634
rect 463 64516 503 64592
rect 575 64516 629 64592
rect 701 64516 749 64592
rect 821 64516 947 64592
rect 463 64480 947 64516
rect 20945 64720 20946 64760
rect 20945 64695 21428 64720
rect 20945 64619 21068 64695
rect 21140 64619 21194 64695
rect 21266 64619 21314 64695
rect 21386 64619 21428 64695
rect 20945 64577 21428 64619
rect 20945 64505 21068 64577
rect 20946 64501 21068 64505
rect 21140 64501 21194 64577
rect 21266 64501 21314 64577
rect 21386 64501 21428 64577
rect 20946 64465 21428 64501
rect 463 63532 947 63557
rect 463 63456 503 63532
rect 575 63456 629 63532
rect 701 63456 749 63532
rect 821 63456 947 63532
rect 463 63414 947 63456
rect 463 63338 503 63414
rect 575 63338 629 63414
rect 701 63338 749 63414
rect 821 63338 947 63414
rect 463 63302 947 63338
rect 20944 63492 21426 63517
rect 20944 63416 21068 63492
rect 21140 63416 21194 63492
rect 21266 63416 21314 63492
rect 21386 63416 21426 63492
rect 20944 63374 21426 63416
rect 20944 63298 21068 63374
rect 21140 63298 21194 63374
rect 21266 63298 21314 63374
rect 21386 63298 21426 63374
rect 20944 63262 21426 63298
rect 464 63068 864 63109
rect 463 63060 864 63068
rect 463 62984 504 63060
rect 576 62984 626 63060
rect 698 62984 752 63060
rect 824 62984 864 63060
rect 463 62913 864 62984
rect 463 62837 504 62913
rect 576 62837 626 62913
rect 698 62837 752 62913
rect 824 62837 864 62913
rect 463 62776 864 62837
rect 463 62700 504 62776
rect 576 62700 626 62776
rect 698 62700 752 62776
rect 824 62700 864 62776
rect 463 62650 864 62700
rect 20946 62057 22370 62082
rect 20946 61981 22010 62057
rect 22082 61981 22136 62057
rect 22208 61981 22256 62057
rect 22328 61981 22370 62057
rect 20946 61939 22370 61981
rect 20946 61863 22010 61939
rect 22082 61863 22136 61939
rect 22208 61863 22256 61939
rect 22328 61863 22370 61939
rect 20946 61827 22370 61863
rect 463 61301 863 61350
rect 463 61225 504 61301
rect 576 61225 626 61301
rect 698 61225 752 61301
rect 824 61225 863 61301
rect 463 61154 863 61225
rect 463 61078 504 61154
rect 576 61078 626 61154
rect 698 61078 752 61154
rect 824 61078 863 61154
rect 463 61017 863 61078
rect 463 60941 504 61017
rect 576 60941 626 61017
rect 698 60941 752 61017
rect 824 60941 863 61017
rect 463 60891 863 60941
rect 463 60684 949 60709
rect 463 60608 503 60684
rect 575 60608 629 60684
rect 701 60608 749 60684
rect 821 60608 949 60684
rect 463 60566 949 60608
rect 463 60490 503 60566
rect 575 60490 629 60566
rect 701 60490 749 60566
rect 821 60490 949 60566
rect 463 60454 949 60490
rect 20946 60695 21428 60720
rect 20946 60619 21068 60695
rect 21140 60619 21194 60695
rect 21266 60619 21314 60695
rect 21386 60619 21428 60695
rect 20946 60577 21428 60619
rect 20946 60501 21068 60577
rect 21140 60501 21194 60577
rect 21266 60501 21314 60577
rect 21386 60501 21428 60577
rect 20946 60465 21428 60501
rect 20945 59546 21427 59571
rect 463 59481 947 59506
rect 463 59405 503 59481
rect 575 59405 629 59481
rect 701 59405 749 59481
rect 821 59405 947 59481
rect 463 59363 947 59405
rect 463 59287 503 59363
rect 575 59287 629 59363
rect 701 59287 749 59363
rect 821 59287 947 59363
rect 20945 59470 21068 59546
rect 21140 59470 21194 59546
rect 21266 59470 21314 59546
rect 21386 59470 21427 59546
rect 20945 59428 21427 59470
rect 20945 59352 21068 59428
rect 21140 59352 21194 59428
rect 21266 59352 21314 59428
rect 21386 59352 21427 59428
rect 20945 59316 21427 59352
rect 463 59251 947 59287
rect 464 59068 864 59109
rect 463 59060 864 59068
rect 463 58984 504 59060
rect 576 58984 626 59060
rect 698 58984 752 59060
rect 824 58984 864 59060
rect 463 58913 864 58984
rect 463 58837 504 58913
rect 576 58837 626 58913
rect 698 58837 752 58913
rect 824 58837 864 58913
rect 463 58776 864 58837
rect 463 58700 504 58776
rect 576 58700 626 58776
rect 698 58700 752 58776
rect 824 58700 864 58776
rect 463 58650 864 58700
rect 20946 58096 22370 58121
rect 20946 58020 22010 58096
rect 22082 58020 22136 58096
rect 22208 58020 22256 58096
rect 22328 58020 22370 58096
rect 20946 57978 22370 58020
rect 20946 57902 22010 57978
rect 22082 57902 22136 57978
rect 22208 57902 22256 57978
rect 22328 57902 22370 57978
rect 20946 57866 22370 57902
rect 463 57299 863 57348
rect 463 57223 504 57299
rect 576 57223 626 57299
rect 698 57223 752 57299
rect 824 57223 863 57299
rect 463 57152 863 57223
rect 463 57076 504 57152
rect 576 57076 626 57152
rect 698 57076 752 57152
rect 824 57076 863 57152
rect 463 57015 863 57076
rect 463 56939 504 57015
rect 576 56939 626 57015
rect 698 56939 752 57015
rect 824 56939 863 57015
rect 463 56889 863 56939
rect 463 56704 947 56729
rect 463 56628 503 56704
rect 575 56628 629 56704
rect 701 56628 749 56704
rect 821 56628 947 56704
rect 463 56586 947 56628
rect 463 56510 503 56586
rect 575 56510 629 56586
rect 701 56510 749 56586
rect 821 56510 947 56586
rect 463 56474 947 56510
rect 20946 56630 21428 56655
rect 20946 56554 21068 56630
rect 21140 56554 21194 56630
rect 21266 56554 21314 56630
rect 21386 56554 21428 56630
rect 20946 56512 21428 56554
rect 20946 56436 21068 56512
rect 21140 56436 21194 56512
rect 21266 56436 21314 56512
rect 21386 56436 21428 56512
rect 20946 56400 21428 56436
rect 463 55497 949 55522
rect 463 55421 503 55497
rect 575 55421 629 55497
rect 701 55421 749 55497
rect 821 55421 949 55497
rect 463 55379 949 55421
rect 463 55303 503 55379
rect 575 55303 629 55379
rect 701 55303 749 55379
rect 821 55303 949 55379
rect 463 55267 949 55303
rect 20945 55447 21427 55472
rect 20945 55371 21068 55447
rect 21140 55371 21194 55447
rect 21266 55371 21314 55447
rect 21386 55371 21427 55447
rect 20945 55329 21427 55371
rect 20945 55253 21068 55329
rect 21140 55253 21194 55329
rect 21266 55253 21314 55329
rect 21386 55253 21427 55329
rect 20945 55217 21427 55253
rect 463 55060 863 55109
rect 463 54984 504 55060
rect 576 54984 626 55060
rect 698 54984 752 55060
rect 824 54984 863 55060
rect 463 54913 863 54984
rect 463 54837 504 54913
rect 576 54837 626 54913
rect 698 54837 752 54913
rect 824 54837 863 54913
rect 463 54776 863 54837
rect 463 54700 504 54776
rect 576 54700 626 54776
rect 698 54700 752 54776
rect 824 54700 863 54776
rect 463 54650 863 54700
rect 20946 54079 22370 54104
rect 20946 54003 22010 54079
rect 22082 54003 22136 54079
rect 22208 54003 22256 54079
rect 22328 54003 22370 54079
rect 20946 53961 22370 54003
rect 20946 53885 22010 53961
rect 22082 53885 22136 53961
rect 22208 53885 22256 53961
rect 22328 53885 22370 53961
rect 20946 53849 22370 53885
rect 463 53301 863 53350
rect 463 53225 504 53301
rect 576 53225 626 53301
rect 698 53225 752 53301
rect 824 53225 863 53301
rect 463 53154 863 53225
rect 463 53078 504 53154
rect 576 53078 626 53154
rect 698 53078 752 53154
rect 824 53078 863 53154
rect 463 53017 863 53078
rect 463 52941 504 53017
rect 576 52941 626 53017
rect 698 52941 752 53017
rect 824 52941 863 53017
rect 463 52891 863 52941
rect 463 52731 947 52756
rect 463 52655 503 52731
rect 575 52655 629 52731
rect 701 52655 749 52731
rect 821 52655 947 52731
rect 463 52613 947 52655
rect 463 52537 503 52613
rect 575 52537 629 52613
rect 701 52537 749 52613
rect 821 52537 947 52613
rect 463 52501 947 52537
rect 20946 52575 21428 52600
rect 20946 52499 21068 52575
rect 21140 52499 21194 52575
rect 21266 52499 21314 52575
rect 21386 52499 21428 52575
rect 20946 52457 21428 52499
rect 20946 52381 21068 52457
rect 21140 52381 21194 52457
rect 21266 52381 21314 52457
rect 21386 52381 21428 52457
rect 20946 52345 21428 52381
rect 463 51544 947 51569
rect 463 51468 503 51544
rect 575 51468 629 51544
rect 701 51468 749 51544
rect 821 51468 947 51544
rect 463 51426 947 51468
rect 463 51350 503 51426
rect 575 51350 629 51426
rect 701 51350 749 51426
rect 821 51350 947 51426
rect 463 51314 947 51350
rect 20946 51440 21428 51465
rect 20946 51364 21068 51440
rect 21140 51364 21194 51440
rect 21266 51364 21314 51440
rect 21386 51364 21428 51440
rect 20946 51322 21428 51364
rect 20946 51246 21068 51322
rect 21140 51246 21194 51322
rect 21266 51246 21314 51322
rect 21386 51246 21428 51322
rect 20946 51210 21428 51246
rect 463 51060 863 51109
rect 463 50984 504 51060
rect 576 50984 626 51060
rect 698 50984 752 51060
rect 824 50984 863 51060
rect 463 50913 863 50984
rect 463 50837 504 50913
rect 576 50837 626 50913
rect 698 50837 752 50913
rect 824 50837 863 50913
rect 463 50776 863 50837
rect 463 50700 504 50776
rect 576 50700 626 50776
rect 698 50700 752 50776
rect 824 50700 863 50776
rect 463 50650 863 50700
rect 20946 50158 22370 50183
rect 20946 50082 22010 50158
rect 22082 50082 22136 50158
rect 22208 50082 22256 50158
rect 22328 50082 22370 50158
rect 20946 50040 22370 50082
rect 20946 49964 22010 50040
rect 22082 49964 22136 50040
rect 22208 49964 22256 50040
rect 22328 49964 22370 50040
rect 20946 49928 22370 49964
rect 463 49301 863 49350
rect 463 49225 504 49301
rect 576 49225 626 49301
rect 698 49225 752 49301
rect 824 49225 863 49301
rect 463 49154 863 49225
rect 463 49078 504 49154
rect 576 49078 626 49154
rect 698 49078 752 49154
rect 824 49078 863 49154
rect 463 49017 863 49078
rect 463 48941 504 49017
rect 576 48941 626 49017
rect 698 48941 752 49017
rect 824 48941 863 49017
rect 463 48891 863 48941
rect 463 48722 947 48747
rect 463 48646 503 48722
rect 575 48646 629 48722
rect 701 48646 749 48722
rect 821 48646 947 48722
rect 463 48604 947 48646
rect 463 48528 503 48604
rect 575 48528 629 48604
rect 701 48528 749 48604
rect 821 48528 947 48604
rect 463 48492 947 48528
rect 20946 48681 21428 48706
rect 20946 48605 21068 48681
rect 21140 48605 21194 48681
rect 21266 48605 21314 48681
rect 21386 48605 21428 48681
rect 20946 48563 21428 48605
rect 20946 48487 21068 48563
rect 21140 48487 21194 48563
rect 21266 48487 21314 48563
rect 21386 48487 21428 48563
rect 20946 48451 21428 48487
rect 463 47569 947 47594
rect 463 47493 503 47569
rect 575 47493 629 47569
rect 701 47493 749 47569
rect 821 47493 947 47569
rect 463 47451 947 47493
rect 463 47375 503 47451
rect 575 47375 629 47451
rect 701 47375 749 47451
rect 821 47375 947 47451
rect 463 47339 947 47375
rect 20946 47528 21428 47553
rect 20946 47452 21068 47528
rect 21140 47452 21194 47528
rect 21266 47452 21314 47528
rect 21386 47452 21428 47528
rect 20946 47410 21428 47452
rect 20946 47334 21068 47410
rect 21140 47334 21194 47410
rect 21266 47334 21314 47410
rect 21386 47334 21428 47410
rect 20946 47298 21428 47334
rect 463 47060 863 47109
rect 463 46984 504 47060
rect 576 46984 626 47060
rect 698 46984 752 47060
rect 824 46984 863 47060
rect 463 46913 863 46984
rect 463 46837 504 46913
rect 576 46837 626 46913
rect 698 46837 752 46913
rect 824 46837 863 46913
rect 463 46776 863 46837
rect 463 46700 504 46776
rect 576 46700 626 46776
rect 698 46700 752 46776
rect 824 46700 863 46776
rect 463 46650 863 46700
rect 20946 45900 22370 45925
rect 20946 45824 22010 45900
rect 22082 45824 22136 45900
rect 22208 45824 22256 45900
rect 22328 45824 22370 45900
rect 20946 45782 22370 45824
rect 20946 45706 22010 45782
rect 22082 45706 22136 45782
rect 22208 45706 22256 45782
rect 22328 45706 22370 45782
rect 20946 45670 22370 45706
rect 463 45300 863 45350
rect 463 45224 504 45300
rect 576 45224 626 45300
rect 698 45224 752 45300
rect 824 45224 863 45300
rect 463 45153 863 45224
rect 463 45077 504 45153
rect 576 45077 626 45153
rect 698 45077 752 45153
rect 824 45077 863 45153
rect 463 45016 863 45077
rect 463 44940 504 45016
rect 576 44940 626 45016
rect 698 44940 752 45016
rect 824 44940 863 45016
rect 463 44891 863 44940
rect 463 44890 836 44891
rect 463 44509 946 44534
rect 463 44433 503 44509
rect 575 44433 629 44509
rect 701 44433 749 44509
rect 821 44433 946 44509
rect 463 44391 946 44433
rect 463 44315 503 44391
rect 575 44315 629 44391
rect 701 44315 749 44391
rect 821 44315 946 44391
rect 463 44279 946 44315
rect 20946 44412 21428 44437
rect 20946 44336 21068 44412
rect 21140 44336 21194 44412
rect 21266 44336 21314 44412
rect 21386 44336 21428 44412
rect 20946 44294 21428 44336
rect 20946 44218 21068 44294
rect 21140 44218 21194 44294
rect 21266 44218 21314 44294
rect 21386 44218 21428 44294
rect 20946 44182 21428 44218
rect 3287 39752 4421 39753
rect 0 39741 21902 39752
rect 0 39661 32 39741
rect 112 39661 157 39741
rect 237 39661 282 39741
rect 362 39726 21902 39741
rect 362 39661 21535 39726
rect 0 39646 21535 39661
rect 21615 39646 21660 39726
rect 21740 39646 21785 39726
rect 21865 39646 21902 39726
rect 0 39635 21902 39646
rect 0 39555 32 39635
rect 112 39555 157 39635
rect 237 39555 282 39635
rect 362 39606 21902 39635
rect 362 39555 21534 39606
rect 0 39526 21534 39555
rect 21614 39526 21659 39606
rect 21739 39526 21784 39606
rect 21864 39526 21902 39606
rect 0 39497 21902 39526
rect 1868 39395 2335 39410
rect 1650 39321 1796 39329
rect 1650 39269 1662 39321
rect 1714 39269 1732 39321
rect 1784 39269 1796 39321
rect 1868 39281 1885 39395
rect 2003 39281 2041 39395
rect 2159 39281 2197 39395
rect 2315 39281 2335 39395
rect 1868 39270 2335 39281
rect 2539 39328 2685 39336
rect 2539 39276 2551 39328
rect 2603 39276 2621 39328
rect 2673 39276 2685 39328
rect 1650 39251 1796 39269
rect 1650 39199 1662 39251
rect 1714 39199 1732 39251
rect 1784 39233 1796 39251
rect 2539 39258 2685 39276
rect 2167 39233 2239 39236
rect 1784 39230 2239 39233
rect 1784 39199 2192 39230
rect 1650 39191 2192 39199
rect 2227 39191 2239 39230
rect 2539 39206 2551 39258
rect 2603 39206 2621 39258
rect 2673 39206 2685 39258
rect 2539 39196 2685 39206
rect 1650 39189 2239 39191
rect 2167 39185 2239 39189
rect 924 39139 1188 39173
rect 463 39138 2973 39139
rect 463 39137 1098 39138
rect 463 39130 941 39137
rect 463 39052 479 39130
rect 561 39052 593 39130
rect 675 39052 707 39130
rect 789 39062 941 39130
rect 1013 39063 1098 39137
rect 1165 39125 2973 39138
rect 1165 39063 1604 39125
rect 1013 39062 1604 39063
rect 789 39059 1604 39062
rect 1638 39124 2973 39125
rect 1638 39069 1920 39124
rect 1954 39069 2973 39124
rect 1638 39059 2973 39069
rect 789 39052 2973 39059
rect 463 39043 2973 39052
rect 924 39024 1188 39043
rect 924 39021 1098 39024
rect 924 38946 944 39021
rect 1016 38949 1098 39021
rect 1165 38949 1188 39024
rect 2889 38982 2950 38987
rect 2889 38981 3370 38982
rect 1016 38946 1188 38949
rect 924 38923 1188 38946
rect 1592 38944 1966 38954
rect 1592 38889 1604 38944
rect 1638 38889 1920 38944
rect 1954 38889 1966 38944
rect 1592 38882 1966 38889
rect 2022 38944 2397 38954
rect 2022 38889 2035 38944
rect 2069 38889 2351 38944
rect 2385 38889 2397 38944
rect 2022 38882 2397 38889
rect 2467 38949 2843 38955
rect 2467 38889 2479 38949
rect 2514 38890 2797 38949
rect 2831 38890 2843 38949
rect 2889 38947 2901 38981
rect 2935 38947 3370 38981
rect 2889 38946 3370 38947
rect 2889 38941 2950 38946
rect 2514 38889 2843 38890
rect 2467 38883 2843 38889
rect 2900 38870 3301 38876
rect 2900 38836 2921 38870
rect 2955 38836 3253 38870
rect 3288 38836 3301 38870
rect 2900 38829 3301 38836
rect 1755 38782 1802 38794
rect 1495 38774 1569 38781
rect 1495 38722 1503 38774
rect 1563 38770 1569 38774
rect 1755 38770 1762 38782
rect 1563 38722 1762 38770
rect 1495 38717 1762 38722
rect 1755 38706 1762 38717
rect 1796 38706 1802 38782
rect 3342 38772 3370 38946
rect 3615 38960 4297 38966
rect 3615 38926 4251 38960
rect 4285 38926 4297 38960
rect 3615 38920 4297 38926
rect 3523 38828 3529 38880
rect 3581 38876 3587 38880
rect 3615 38876 3650 38920
rect 4610 38879 4662 38885
rect 4092 38876 4156 38878
rect 3581 38870 3650 38876
rect 3587 38836 3650 38870
rect 3581 38830 3650 38836
rect 4075 38870 4385 38876
rect 4075 38836 4105 38870
rect 4139 38836 4339 38870
rect 4373 38836 4385 38870
rect 4075 38830 4385 38836
rect 3581 38828 3587 38830
rect 4092 38826 4156 38830
rect 4608 38829 4610 38877
rect 3792 38813 3841 38825
rect 4610 38821 4662 38827
rect 3792 38779 3800 38813
rect 3835 38779 3841 38813
rect 3792 38772 3841 38779
rect 3341 38737 3841 38772
rect 1755 38694 1802 38706
rect 0 38586 1593 38595
rect 0 38508 16 38586
rect 98 38508 130 38586
rect 212 38508 244 38586
rect 326 38508 1593 38586
rect 0 38499 1593 38508
rect 3608 38348 3660 38354
rect 1893 38305 3608 38334
rect 1465 38217 1471 38269
rect 1523 38268 1529 38269
rect 1523 38258 1773 38268
rect 1523 38224 1715 38258
rect 1749 38224 1773 38258
rect 1523 38218 1773 38224
rect 1801 38261 1847 38275
rect 1801 38227 1807 38261
rect 1841 38227 1847 38261
rect 1523 38217 1529 38218
rect 1801 38210 1847 38227
rect 1893 38258 1941 38305
rect 3608 38290 3660 38296
rect 1893 38224 1899 38258
rect 1933 38224 1941 38258
rect 1893 38212 1941 38224
rect 2019 38252 2076 38275
rect 2019 38218 2029 38252
rect 2063 38218 2076 38252
rect 1805 38184 1847 38210
rect 2019 38202 2076 38218
rect 4652 38267 4704 38273
rect 4652 38209 4704 38215
rect 2019 38184 2063 38202
rect 1805 38155 2063 38184
rect 463 38042 2056 38051
rect 463 37964 479 38042
rect 561 37964 593 38042
rect 675 37964 707 38042
rect 789 37964 2056 38042
rect 463 37955 2056 37964
rect 3517 37889 3523 37897
rect 1874 37854 3523 37889
rect 1457 37738 1463 37790
rect 1515 37738 1539 37790
rect 1799 37787 1845 37851
rect 1799 37753 1805 37787
rect 1839 37753 1845 37787
rect 1799 37708 1845 37753
rect 1874 37788 1940 37854
rect 3517 37845 3523 37854
rect 3575 37845 3581 37897
rect 1874 37754 1889 37788
rect 1923 37754 1940 37788
rect 1874 37738 1940 37754
rect 1980 37782 2032 37795
rect 1980 37748 1986 37782
rect 2020 37748 2032 37782
rect 1980 37708 2032 37748
rect 4652 37791 4704 37797
rect 4652 37733 4704 37739
rect 1799 37680 2032 37708
rect 0 37498 1317 37507
rect 0 37420 16 37498
rect 98 37420 130 37498
rect 212 37420 244 37498
rect 326 37420 1317 37498
rect 0 37411 1317 37420
rect 1680 37358 1739 37375
rect 1680 37306 1683 37358
rect 1735 37306 1739 37358
rect 1680 37252 1739 37306
rect 1680 37200 1683 37252
rect 1735 37200 1739 37252
rect 1680 37150 1739 37200
rect 3332 37265 3841 37300
rect 2867 37172 3295 37178
rect 1680 37144 2320 37150
rect 924 37079 1188 37111
rect 1680 37090 1957 37144
rect 1991 37143 2320 37144
rect 1991 37090 2273 37143
rect 1680 37089 2273 37090
rect 2307 37089 2320 37143
rect 1680 37084 2320 37089
rect 2416 37146 2804 37152
rect 2416 37095 2436 37146
rect 2471 37143 2804 37146
rect 2471 37095 2753 37143
rect 2416 37092 2753 37095
rect 2787 37092 2804 37143
rect 2867 37138 2902 37172
rect 2936 37171 3295 37172
rect 2936 37138 3237 37171
rect 2867 37137 3237 37138
rect 3271 37137 3295 37171
rect 2867 37131 3295 37137
rect 2416 37085 2804 37092
rect 1680 37083 1739 37084
rect 1945 37083 2320 37084
rect 924 36991 947 37079
rect 1042 36991 1080 37079
rect 1165 36991 1188 37079
rect 3332 37069 3375 37265
rect 3806 37233 3841 37265
rect 3801 37227 3848 37233
rect 3801 37193 3807 37227
rect 3841 37193 3848 37227
rect 3547 37176 3553 37182
rect 3523 37130 3553 37176
rect 3605 37130 3646 37182
rect 3801 37181 3848 37193
rect 4609 37181 4661 37187
rect 2969 37058 3375 37069
rect 2910 37038 3375 37058
rect 3610 37086 3646 37130
rect 4075 37178 4156 37180
rect 4075 37170 4569 37178
rect 4075 37136 4105 37170
rect 4139 37136 4523 37170
rect 4557 37136 4569 37170
rect 4075 37130 4569 37136
rect 4075 37128 4156 37130
rect 4609 37123 4661 37129
rect 3610 37080 4297 37086
rect 3610 37046 4251 37080
rect 4285 37046 4297 37080
rect 3610 37038 4297 37046
rect 2910 37003 2916 37038
rect 2953 37034 3375 37038
rect 2953 37023 2987 37034
rect 2953 37003 2959 37023
rect 2910 36991 2959 37003
rect 924 36963 1188 36991
rect 463 36954 2973 36963
rect 463 36876 479 36954
rect 561 36876 593 36954
rect 675 36876 707 36954
rect 789 36949 2973 36954
rect 789 36876 947 36949
rect 463 36867 947 36876
rect 924 36861 947 36867
rect 1042 36861 1081 36949
rect 1165 36867 2973 36949
rect 1165 36861 1188 36867
rect 924 36835 1188 36861
rect 2538 36830 2685 36838
rect 2538 36778 2551 36830
rect 2603 36778 2621 36830
rect 2673 36778 2685 36830
rect 2538 36763 2685 36778
rect 2538 36711 2551 36763
rect 2603 36711 2621 36763
rect 2673 36711 2685 36763
rect 2538 36649 2685 36711
rect 2752 36830 2899 36838
rect 2752 36778 2765 36830
rect 2817 36778 2835 36830
rect 2887 36778 2899 36830
rect 2752 36765 2899 36778
rect 2752 36713 2765 36765
rect 2817 36713 2835 36765
rect 2887 36713 2899 36765
rect 2752 36707 2899 36713
rect 20527 36172 21428 36198
rect 20527 36092 21061 36172
rect 21141 36092 21186 36172
rect 21266 36092 21311 36172
rect 21391 36092 21428 36172
rect 20527 36052 21428 36092
rect 20527 35972 21060 36052
rect 21140 35972 21185 36052
rect 21265 35972 21310 36052
rect 21390 35972 21428 36052
rect 20527 35943 21428 35972
rect 21028 35592 21428 35642
rect 21028 35516 21069 35592
rect 21141 35516 21191 35592
rect 21263 35516 21317 35592
rect 21389 35516 21428 35592
rect 21028 35445 21428 35516
rect 21028 35369 21069 35445
rect 21141 35369 21191 35445
rect 21263 35369 21317 35445
rect 21389 35369 21428 35445
rect 21028 35308 21428 35369
rect 21028 35232 21069 35308
rect 21141 35232 21191 35308
rect 21263 35232 21317 35308
rect 21389 35232 21428 35308
rect 21028 35183 21428 35232
rect 21028 35182 21401 35183
rect 20526 34676 21902 34702
rect 20526 34596 20560 34676
rect 20640 34596 20685 34676
rect 20765 34596 20810 34676
rect 20890 34596 21535 34676
rect 21615 34596 21660 34676
rect 21740 34596 21785 34676
rect 21865 34596 21902 34676
rect 20526 34556 21902 34596
rect 20526 34476 20559 34556
rect 20639 34476 20684 34556
rect 20764 34476 20809 34556
rect 20889 34476 21534 34556
rect 21614 34476 21659 34556
rect 21739 34476 21784 34556
rect 21864 34476 21902 34556
rect 20526 34447 21902 34476
rect 21028 33832 21428 33882
rect 21028 33756 21069 33832
rect 21141 33756 21191 33832
rect 21263 33756 21317 33832
rect 21389 33756 21428 33832
rect 21028 33685 21428 33756
rect 21028 33609 21069 33685
rect 21141 33609 21191 33685
rect 21263 33609 21317 33685
rect 21389 33609 21428 33685
rect 21028 33548 21428 33609
rect 21028 33472 21069 33548
rect 21141 33472 21191 33548
rect 21263 33472 21317 33548
rect 21389 33472 21428 33548
rect 21028 33423 21428 33472
rect 21028 33422 21401 33423
rect 20514 33117 21427 33143
rect 20514 33037 21060 33117
rect 21140 33037 21185 33117
rect 21265 33037 21310 33117
rect 21390 33037 21427 33117
rect 20514 32997 21427 33037
rect 20514 32917 21059 32997
rect 21139 32917 21184 32997
rect 21264 32917 21309 32997
rect 21389 32917 21427 32997
rect 20514 32888 21427 32917
rect 463 32302 21428 32360
rect 463 32226 503 32302
rect 575 32226 629 32302
rect 701 32226 749 32302
rect 821 32226 21068 32302
rect 21140 32226 21194 32302
rect 21266 32226 21314 32302
rect 21386 32226 21428 32302
rect 463 32184 21428 32226
rect 463 32108 503 32184
rect 575 32108 629 32184
rect 701 32108 749 32184
rect 821 32108 21068 32184
rect 21140 32108 21194 32184
rect 21266 32108 21314 32184
rect 21386 32108 21428 32184
rect 463 32073 21428 32108
rect 463 32072 1825 32073
rect 2313 32072 21428 32073
rect 463 31520 946 31545
rect 463 31444 503 31520
rect 575 31444 629 31520
rect 701 31444 749 31520
rect 821 31444 946 31520
rect 463 31402 946 31444
rect 463 31326 503 31402
rect 575 31326 629 31402
rect 701 31326 749 31402
rect 821 31326 946 31402
rect 463 31290 946 31326
rect 20946 31520 21428 31545
rect 20946 31444 21068 31520
rect 21140 31444 21194 31520
rect 21266 31444 21314 31520
rect 21386 31444 21428 31520
rect 20946 31402 21428 31444
rect 20946 31326 21068 31402
rect 21140 31326 21194 31402
rect 21266 31326 21314 31402
rect 21386 31326 21428 31402
rect 20946 31290 21428 31326
rect 463 31061 863 31111
rect 463 30985 504 31061
rect 576 30985 626 31061
rect 698 30985 752 31061
rect 824 30985 863 31061
rect 463 30914 863 30985
rect 463 30838 504 30914
rect 576 30838 626 30914
rect 698 30838 752 30914
rect 824 30838 863 30914
rect 463 30777 863 30838
rect 463 30701 504 30777
rect 576 30701 626 30777
rect 698 30701 752 30777
rect 824 30701 863 30777
rect 463 30651 863 30701
rect 20946 30130 22370 30155
rect 20946 30054 22010 30130
rect 22082 30054 22136 30130
rect 22208 30054 22256 30130
rect 22328 30054 22370 30130
rect 20946 30012 22370 30054
rect 20946 29936 22010 30012
rect 22082 29936 22136 30012
rect 22208 29936 22256 30012
rect 22328 29936 22370 30012
rect 20946 29900 22370 29936
rect 463 29294 863 29350
rect 463 29218 504 29294
rect 576 29218 626 29294
rect 698 29218 752 29294
rect 824 29218 863 29294
rect 463 29147 863 29218
rect 463 29071 504 29147
rect 576 29071 626 29147
rect 698 29071 752 29147
rect 824 29071 863 29147
rect 463 29010 863 29071
rect 463 28934 504 29010
rect 576 28934 626 29010
rect 698 28934 752 29010
rect 824 28934 863 29010
rect 463 28890 863 28934
rect 463 28608 946 28633
rect 463 28532 503 28608
rect 575 28532 629 28608
rect 701 28532 749 28608
rect 821 28532 946 28608
rect 463 28490 946 28532
rect 463 28414 503 28490
rect 575 28414 629 28490
rect 701 28414 749 28490
rect 821 28414 946 28490
rect 463 28378 946 28414
rect 20946 28559 21428 28584
rect 20946 28483 21068 28559
rect 21140 28483 21194 28559
rect 21266 28483 21314 28559
rect 21386 28483 21428 28559
rect 20946 28441 21428 28483
rect 20946 28365 21068 28441
rect 21140 28365 21194 28441
rect 21266 28365 21314 28441
rect 21386 28365 21428 28441
rect 20946 28329 21428 28365
rect 463 27604 946 27629
rect 463 27528 503 27604
rect 575 27528 629 27604
rect 701 27528 749 27604
rect 821 27528 946 27604
rect 463 27486 946 27528
rect 463 27410 503 27486
rect 575 27410 629 27486
rect 701 27410 749 27486
rect 821 27410 946 27486
rect 463 27374 946 27410
rect 20945 27442 21427 27467
rect 20945 27366 21068 27442
rect 21140 27366 21194 27442
rect 21266 27366 21314 27442
rect 21386 27366 21427 27442
rect 20945 27324 21427 27366
rect 20945 27248 21068 27324
rect 21140 27248 21194 27324
rect 21266 27248 21314 27324
rect 21386 27248 21427 27324
rect 20945 27212 21427 27248
rect 463 27060 863 27109
rect 463 26984 504 27060
rect 576 26984 626 27060
rect 698 26984 752 27060
rect 824 26984 863 27060
rect 463 26913 863 26984
rect 463 26837 504 26913
rect 576 26837 626 26913
rect 698 26837 752 26913
rect 824 26837 863 26913
rect 463 26776 863 26837
rect 463 26700 504 26776
rect 576 26700 626 26776
rect 698 26700 752 26776
rect 824 26700 863 26776
rect 463 26650 863 26700
rect 20946 25971 22370 25996
rect 20946 25895 22010 25971
rect 22082 25895 22136 25971
rect 22208 25895 22256 25971
rect 22328 25895 22370 25971
rect 20946 25853 22370 25895
rect 20946 25777 22010 25853
rect 22082 25777 22136 25853
rect 22208 25777 22256 25853
rect 22328 25777 22370 25853
rect 20946 25741 22370 25777
rect 463 25300 863 25349
rect 463 25224 504 25300
rect 576 25224 626 25300
rect 698 25224 752 25300
rect 824 25224 863 25300
rect 463 25153 863 25224
rect 463 25077 504 25153
rect 576 25077 626 25153
rect 698 25077 752 25153
rect 824 25077 863 25153
rect 463 25016 863 25077
rect 463 24940 504 25016
rect 576 24940 626 25016
rect 698 24940 752 25016
rect 824 24940 863 25016
rect 463 24890 863 24940
rect 463 24626 947 24651
rect 463 24550 503 24626
rect 575 24550 629 24626
rect 701 24550 749 24626
rect 821 24550 947 24626
rect 463 24508 947 24550
rect 463 24432 503 24508
rect 575 24432 629 24508
rect 701 24432 749 24508
rect 821 24432 947 24508
rect 463 24396 947 24432
rect 20946 24599 21428 24624
rect 20946 24523 21068 24599
rect 21140 24523 21194 24599
rect 21266 24523 21314 24599
rect 21386 24523 21428 24599
rect 20946 24481 21428 24523
rect 20946 24405 21068 24481
rect 21140 24405 21194 24481
rect 21266 24405 21314 24481
rect 21386 24405 21428 24481
rect 20946 24369 21428 24405
rect 463 23544 947 23569
rect 463 23468 503 23544
rect 575 23468 629 23544
rect 701 23468 749 23544
rect 821 23468 947 23544
rect 463 23426 947 23468
rect 463 23350 503 23426
rect 575 23350 629 23426
rect 701 23350 749 23426
rect 821 23350 947 23426
rect 463 23314 947 23350
rect 20946 23424 21428 23449
rect 20946 23348 21068 23424
rect 21140 23348 21194 23424
rect 21266 23348 21314 23424
rect 21386 23348 21428 23424
rect 20946 23306 21428 23348
rect 20946 23230 21068 23306
rect 21140 23230 21194 23306
rect 21266 23230 21314 23306
rect 21386 23230 21428 23306
rect 20946 23194 21428 23230
rect 463 23060 863 23109
rect 463 22984 504 23060
rect 576 22984 626 23060
rect 698 22984 752 23060
rect 824 22984 863 23060
rect 463 22913 863 22984
rect 463 22837 504 22913
rect 576 22837 626 22913
rect 698 22837 752 22913
rect 824 22837 863 22913
rect 463 22776 863 22837
rect 463 22700 504 22776
rect 576 22700 626 22776
rect 698 22700 752 22776
rect 824 22700 863 22776
rect 463 22650 863 22700
rect 20946 22181 22370 22206
rect 20946 22105 22010 22181
rect 22082 22105 22136 22181
rect 22208 22105 22256 22181
rect 22328 22105 22370 22181
rect 20946 22063 22370 22105
rect 20946 21987 22010 22063
rect 22082 21987 22136 22063
rect 22208 21987 22256 22063
rect 22328 21987 22370 22063
rect 20946 21951 22370 21987
rect 463 21301 863 21350
rect 463 21225 504 21301
rect 576 21225 626 21301
rect 698 21225 752 21301
rect 824 21225 863 21301
rect 463 21154 863 21225
rect 463 21078 504 21154
rect 576 21078 626 21154
rect 698 21078 752 21154
rect 824 21078 863 21154
rect 463 21017 863 21078
rect 463 20941 504 21017
rect 576 20941 626 21017
rect 698 20941 752 21017
rect 824 20941 863 21017
rect 463 20891 863 20941
rect 463 20669 947 20694
rect 463 20593 503 20669
rect 575 20593 629 20669
rect 701 20593 749 20669
rect 821 20593 947 20669
rect 463 20551 947 20593
rect 463 20475 503 20551
rect 575 20475 629 20551
rect 701 20475 749 20551
rect 821 20475 947 20551
rect 463 20439 947 20475
rect 20945 20583 21427 20608
rect 20945 20507 21068 20583
rect 21140 20507 21194 20583
rect 21266 20507 21314 20583
rect 21386 20507 21427 20583
rect 20945 20465 21427 20507
rect 20945 20389 21068 20465
rect 21140 20389 21194 20465
rect 21266 20389 21314 20465
rect 21386 20389 21427 20465
rect 20945 20353 21427 20389
rect 463 19568 947 19593
rect 463 19492 503 19568
rect 575 19492 629 19568
rect 701 19492 749 19568
rect 821 19492 947 19568
rect 463 19450 947 19492
rect 463 19374 503 19450
rect 575 19374 629 19450
rect 701 19374 749 19450
rect 821 19374 947 19450
rect 463 19338 947 19374
rect 20945 19412 21427 19437
rect 20945 19336 21068 19412
rect 21140 19336 21194 19412
rect 21266 19336 21314 19412
rect 21386 19336 21427 19412
rect 20945 19294 21427 19336
rect 20945 19218 21068 19294
rect 21140 19218 21194 19294
rect 21266 19218 21314 19294
rect 21386 19218 21427 19294
rect 20945 19182 21427 19218
rect 463 19060 863 19109
rect 463 18984 504 19060
rect 576 18984 626 19060
rect 698 18984 752 19060
rect 824 18984 863 19060
rect 463 18913 863 18984
rect 463 18837 504 18913
rect 576 18837 626 18913
rect 698 18837 752 18913
rect 824 18837 863 18913
rect 463 18776 863 18837
rect 463 18700 504 18776
rect 576 18700 626 18776
rect 698 18700 752 18776
rect 824 18700 863 18776
rect 463 18650 863 18700
rect 20946 18074 22370 18099
rect 20946 17998 22010 18074
rect 22082 17998 22136 18074
rect 22208 17998 22256 18074
rect 22328 17998 22370 18074
rect 20946 17956 22370 17998
rect 20946 17880 22010 17956
rect 22082 17880 22136 17956
rect 22208 17880 22256 17956
rect 22328 17880 22370 17956
rect 20946 17844 22370 17880
rect 463 17300 863 17349
rect 463 17224 504 17300
rect 576 17224 626 17300
rect 698 17224 752 17300
rect 824 17224 863 17300
rect 463 17153 863 17224
rect 463 17077 504 17153
rect 576 17077 626 17153
rect 698 17077 752 17153
rect 824 17077 863 17153
rect 463 17016 863 17077
rect 463 16940 504 17016
rect 576 16940 626 17016
rect 698 16940 752 17016
rect 824 16940 863 17016
rect 463 16890 863 16940
rect 463 16702 948 16727
rect 463 16626 503 16702
rect 575 16626 629 16702
rect 701 16626 749 16702
rect 821 16626 948 16702
rect 463 16584 948 16626
rect 463 16508 503 16584
rect 575 16508 629 16584
rect 701 16508 749 16584
rect 821 16508 948 16584
rect 463 16472 948 16508
rect 20945 16651 21427 16676
rect 20945 16575 21068 16651
rect 21140 16575 21194 16651
rect 21266 16575 21314 16651
rect 21386 16575 21427 16651
rect 20945 16533 21427 16575
rect 20945 16457 21068 16533
rect 21140 16457 21194 16533
rect 21266 16457 21314 16533
rect 21386 16457 21427 16533
rect 20945 16421 21427 16457
rect 463 15486 949 15511
rect 463 15410 503 15486
rect 575 15410 629 15486
rect 701 15410 749 15486
rect 821 15410 949 15486
rect 463 15368 949 15410
rect 463 15292 503 15368
rect 575 15292 629 15368
rect 701 15292 749 15368
rect 821 15292 949 15368
rect 463 15256 949 15292
rect 20945 15437 21427 15462
rect 20945 15361 21068 15437
rect 21140 15361 21194 15437
rect 21266 15361 21314 15437
rect 21386 15361 21427 15437
rect 20945 15319 21427 15361
rect 20945 15243 21068 15319
rect 21140 15243 21194 15319
rect 21266 15243 21314 15319
rect 21386 15243 21427 15319
rect 20945 15207 21427 15243
rect 463 15060 863 15109
rect 463 14984 504 15060
rect 576 14984 626 15060
rect 698 14984 752 15060
rect 824 14984 863 15060
rect 463 14913 863 14984
rect 463 14837 504 14913
rect 576 14837 626 14913
rect 698 14837 752 14913
rect 824 14837 863 14913
rect 463 14776 863 14837
rect 463 14700 504 14776
rect 576 14700 626 14776
rect 698 14700 752 14776
rect 824 14700 863 14776
rect 463 14650 863 14700
rect 20946 14256 22370 14281
rect 20946 14180 22010 14256
rect 22082 14180 22136 14256
rect 22208 14180 22256 14256
rect 22328 14180 22370 14256
rect 20946 14138 22370 14180
rect 20946 14062 22010 14138
rect 22082 14062 22136 14138
rect 22208 14062 22256 14138
rect 22328 14062 22370 14138
rect 20946 14026 22370 14062
rect 463 13300 863 13349
rect 463 13224 504 13300
rect 576 13224 626 13300
rect 698 13224 752 13300
rect 824 13224 863 13300
rect 463 13153 863 13224
rect 463 13077 504 13153
rect 576 13077 626 13153
rect 698 13077 752 13153
rect 824 13077 863 13153
rect 463 13016 863 13077
rect 463 12940 504 13016
rect 576 12940 626 13016
rect 698 12940 752 13016
rect 824 12940 863 13016
rect 463 12890 863 12940
rect 463 12621 947 12646
rect 463 12545 503 12621
rect 575 12545 629 12621
rect 701 12545 749 12621
rect 821 12545 947 12621
rect 463 12503 947 12545
rect 463 12427 503 12503
rect 575 12427 629 12503
rect 701 12427 749 12503
rect 821 12427 947 12503
rect 463 12391 947 12427
rect 20946 12594 21428 12619
rect 20946 12518 21068 12594
rect 21140 12518 21194 12594
rect 21266 12518 21314 12594
rect 21386 12518 21428 12594
rect 20946 12476 21428 12518
rect 20946 12400 21068 12476
rect 21140 12400 21194 12476
rect 21266 12400 21314 12476
rect 21386 12400 21428 12476
rect 20946 12364 21428 12400
rect 463 11499 947 11524
rect 463 11423 503 11499
rect 575 11423 629 11499
rect 701 11423 749 11499
rect 821 11423 947 11499
rect 463 11381 947 11423
rect 463 11305 503 11381
rect 575 11305 629 11381
rect 701 11305 749 11381
rect 821 11305 947 11381
rect 463 11269 947 11305
rect 20946 11437 21427 11462
rect 20946 11361 21068 11437
rect 21140 11361 21194 11437
rect 21266 11361 21314 11437
rect 21386 11361 21427 11437
rect 20946 11319 21427 11361
rect 20946 11243 21068 11319
rect 21140 11243 21194 11319
rect 21266 11243 21314 11319
rect 21386 11243 21427 11319
rect 20946 11207 21427 11243
rect 463 11061 863 11110
rect 463 10985 504 11061
rect 576 10985 626 11061
rect 698 10985 752 11061
rect 824 10985 863 11061
rect 463 10914 863 10985
rect 463 10838 504 10914
rect 576 10838 626 10914
rect 698 10838 752 10914
rect 824 10838 863 10914
rect 463 10777 863 10838
rect 463 10701 504 10777
rect 576 10701 626 10777
rect 698 10701 752 10777
rect 824 10701 863 10777
rect 463 10651 863 10701
rect 20946 10292 22370 10317
rect 20946 10216 22010 10292
rect 22082 10216 22136 10292
rect 22208 10216 22256 10292
rect 22328 10216 22370 10292
rect 20946 10174 22370 10216
rect 20946 10098 22010 10174
rect 22082 10098 22136 10174
rect 22208 10098 22256 10174
rect 22328 10098 22370 10174
rect 20946 10062 22370 10098
rect 463 9299 863 9348
rect 463 9223 504 9299
rect 576 9223 626 9299
rect 698 9223 752 9299
rect 824 9223 863 9299
rect 463 9152 863 9223
rect 463 9076 504 9152
rect 576 9076 626 9152
rect 698 9076 752 9152
rect 824 9076 863 9152
rect 463 9015 863 9076
rect 463 8939 504 9015
rect 576 8939 626 9015
rect 698 8939 752 9015
rect 824 8939 863 9015
rect 463 8889 863 8939
rect 463 8639 946 8664
rect 463 8563 503 8639
rect 575 8563 629 8639
rect 701 8563 749 8639
rect 821 8563 946 8639
rect 463 8521 946 8563
rect 463 8445 503 8521
rect 575 8445 629 8521
rect 701 8445 749 8521
rect 821 8445 946 8521
rect 463 8409 946 8445
rect 20946 8594 21428 8619
rect 20946 8518 21068 8594
rect 21140 8518 21194 8594
rect 21266 8518 21314 8594
rect 21386 8518 21428 8594
rect 20946 8476 21428 8518
rect 20946 8400 21068 8476
rect 21140 8400 21194 8476
rect 21266 8400 21314 8476
rect 21386 8400 21428 8476
rect 20946 8364 21428 8400
rect 463 7528 946 7553
rect 463 7452 503 7528
rect 575 7452 629 7528
rect 701 7452 749 7528
rect 821 7452 946 7528
rect 463 7410 946 7452
rect 463 7334 503 7410
rect 575 7334 629 7410
rect 701 7334 749 7410
rect 821 7334 946 7410
rect 463 7298 946 7334
rect 20946 7437 21427 7462
rect 20946 7361 21068 7437
rect 21140 7361 21194 7437
rect 21266 7361 21314 7437
rect 21386 7361 21427 7437
rect 20946 7319 21427 7361
rect 20946 7243 21068 7319
rect 21140 7243 21194 7319
rect 21266 7243 21314 7319
rect 21386 7243 21427 7319
rect 20946 7207 21427 7243
rect 463 7061 863 7110
rect 463 6985 504 7061
rect 576 6985 626 7061
rect 698 6985 752 7061
rect 824 6985 863 7061
rect 463 6914 863 6985
rect 463 6838 504 6914
rect 576 6838 626 6914
rect 698 6838 752 6914
rect 824 6838 863 6914
rect 463 6777 863 6838
rect 463 6701 504 6777
rect 576 6701 626 6777
rect 698 6701 752 6777
rect 824 6701 863 6777
rect 463 6651 863 6701
rect 20946 6280 22370 6305
rect 20946 6204 22010 6280
rect 22082 6204 22136 6280
rect 22208 6204 22256 6280
rect 22328 6204 22370 6280
rect 20946 6162 22370 6204
rect 20946 6086 22010 6162
rect 22082 6086 22136 6162
rect 22208 6086 22256 6162
rect 22328 6086 22370 6162
rect 20946 6050 22370 6086
rect 463 5300 863 5349
rect 463 5224 504 5300
rect 576 5224 626 5300
rect 698 5224 752 5300
rect 824 5224 863 5300
rect 463 5153 863 5224
rect 463 5077 504 5153
rect 576 5077 626 5153
rect 698 5077 752 5153
rect 824 5077 863 5153
rect 463 5016 863 5077
rect 463 4940 504 5016
rect 576 4940 626 5016
rect 698 4940 752 5016
rect 824 4940 863 5016
rect 463 4890 863 4940
rect 463 4705 948 4730
rect 463 4629 503 4705
rect 575 4629 629 4705
rect 701 4629 749 4705
rect 821 4629 948 4705
rect 463 4587 948 4629
rect 463 4511 503 4587
rect 575 4511 629 4587
rect 701 4511 749 4587
rect 821 4511 948 4587
rect 463 4475 948 4511
rect 20946 4594 21428 4619
rect 20946 4518 21068 4594
rect 21140 4518 21194 4594
rect 21266 4518 21314 4594
rect 21386 4518 21428 4594
rect 20946 4476 21428 4518
rect 20946 4400 21068 4476
rect 21140 4400 21194 4476
rect 21266 4400 21314 4476
rect 21386 4400 21428 4476
rect 20946 4364 21428 4400
rect 463 3528 946 3553
rect 463 3452 503 3528
rect 575 3452 629 3528
rect 701 3452 749 3528
rect 821 3452 946 3528
rect 463 3410 946 3452
rect 463 3334 503 3410
rect 575 3334 629 3410
rect 701 3334 749 3410
rect 821 3334 946 3410
rect 463 3298 946 3334
rect 20946 3437 21427 3462
rect 20946 3361 21068 3437
rect 21140 3361 21194 3437
rect 21266 3361 21314 3437
rect 21386 3361 21427 3437
rect 20946 3319 21427 3361
rect 20946 3243 21068 3319
rect 21140 3243 21194 3319
rect 21266 3243 21314 3319
rect 21386 3243 21427 3319
rect 20946 3207 21427 3243
rect 463 3061 863 3110
rect 463 2985 504 3061
rect 576 2985 626 3061
rect 698 2985 752 3061
rect 824 2985 863 3061
rect 463 2914 863 2985
rect 463 2838 504 2914
rect 576 2838 626 2914
rect 698 2838 752 2914
rect 824 2838 863 2914
rect 463 2777 863 2838
rect 463 2701 504 2777
rect 576 2701 626 2777
rect 698 2701 752 2777
rect 824 2701 863 2777
rect 463 2651 863 2701
rect 20946 2280 22370 2305
rect 20946 2204 22010 2280
rect 22082 2204 22136 2280
rect 22208 2204 22256 2280
rect 22328 2204 22370 2280
rect 20946 2162 22370 2204
rect 20946 2086 22010 2162
rect 22082 2086 22136 2162
rect 22208 2086 22256 2162
rect 22328 2086 22370 2162
rect 20946 2050 22370 2086
rect 463 1300 863 1349
rect 463 1224 504 1300
rect 576 1224 626 1300
rect 698 1224 752 1300
rect 824 1224 863 1300
rect 463 1153 863 1224
rect 463 1077 504 1153
rect 576 1077 626 1153
rect 698 1077 752 1153
rect 824 1077 863 1153
rect 463 1016 863 1077
rect 463 940 504 1016
rect 576 940 626 1016
rect 698 940 752 1016
rect 824 940 863 1016
rect 463 890 863 940
rect 463 705 946 730
rect 463 629 503 705
rect 575 629 629 705
rect 701 629 749 705
rect 821 629 946 705
rect 463 587 946 629
rect 463 511 503 587
rect 575 511 629 587
rect 701 511 749 587
rect 821 511 946 587
rect 463 475 946 511
rect 20946 594 21428 619
rect 20946 518 21068 594
rect 21140 518 21194 594
rect 21266 518 21314 594
rect 21386 518 21428 594
rect 20946 476 21428 518
rect 20946 400 21068 476
rect 21140 400 21194 476
rect 21266 400 21314 476
rect 21386 400 21428 476
rect 20946 364 21428 400
<< via1 >>
rect 503 75376 575 75452
rect 629 75376 701 75452
rect 749 75376 821 75452
rect 503 75258 575 75334
rect 629 75258 701 75334
rect 749 75258 821 75334
rect 21068 75416 21140 75492
rect 21194 75416 21266 75492
rect 21314 75416 21386 75492
rect 21068 75298 21140 75374
rect 21194 75298 21266 75374
rect 21314 75298 21386 75374
rect 504 74984 576 75060
rect 626 74984 698 75060
rect 752 74984 824 75060
rect 504 74837 576 74913
rect 626 74837 698 74913
rect 752 74837 824 74913
rect 504 74700 576 74776
rect 626 74700 698 74776
rect 752 74700 824 74776
rect 22010 73995 22082 74071
rect 22136 73995 22208 74071
rect 22256 73995 22328 74071
rect 22010 73877 22082 73953
rect 22136 73877 22208 73953
rect 22256 73877 22328 73953
rect 504 73224 576 73300
rect 626 73224 698 73300
rect 752 73224 824 73300
rect 504 73077 576 73153
rect 626 73077 698 73153
rect 752 73077 824 73153
rect 504 72940 576 73016
rect 626 72940 698 73016
rect 752 72940 824 73016
rect 503 72703 575 72779
rect 629 72703 701 72779
rect 749 72703 821 72779
rect 503 72585 575 72661
rect 629 72585 701 72661
rect 749 72585 821 72661
rect 21068 72619 21140 72695
rect 21194 72619 21266 72695
rect 21314 72619 21386 72695
rect 21068 72501 21140 72577
rect 21194 72501 21266 72577
rect 21314 72501 21386 72577
rect 503 71376 575 71452
rect 629 71376 701 71452
rect 749 71376 821 71452
rect 503 71258 575 71334
rect 629 71258 701 71334
rect 749 71258 821 71334
rect 21068 71416 21140 71492
rect 21194 71416 21266 71492
rect 21314 71416 21386 71492
rect 21068 71298 21140 71374
rect 21194 71298 21266 71374
rect 21314 71298 21386 71374
rect 504 70984 576 71060
rect 626 70984 698 71060
rect 752 70984 824 71060
rect 504 70837 576 70913
rect 626 70837 698 70913
rect 752 70837 824 70913
rect 504 70700 576 70776
rect 626 70700 698 70776
rect 752 70700 824 70776
rect 22010 69995 22082 70071
rect 22136 69995 22208 70071
rect 22256 69995 22328 70071
rect 22010 69877 22082 69953
rect 22136 69877 22208 69953
rect 22256 69877 22328 69953
rect 504 69224 576 69300
rect 626 69224 698 69300
rect 752 69224 824 69300
rect 504 69077 576 69153
rect 626 69077 698 69153
rect 752 69077 824 69153
rect 504 68940 576 69016
rect 626 68940 698 69016
rect 752 68940 824 69016
rect 503 68703 575 68779
rect 629 68703 701 68779
rect 749 68703 821 68779
rect 503 68585 575 68661
rect 629 68585 701 68661
rect 749 68585 821 68661
rect 21068 68619 21140 68695
rect 21194 68619 21266 68695
rect 21314 68619 21386 68695
rect 21068 68501 21140 68577
rect 21194 68501 21266 68577
rect 21314 68501 21386 68577
rect 503 67374 575 67450
rect 629 67374 701 67450
rect 749 67374 821 67450
rect 503 67256 575 67332
rect 629 67256 701 67332
rect 749 67256 821 67332
rect 21068 67416 21140 67492
rect 21194 67416 21266 67492
rect 21314 67416 21386 67492
rect 21068 67298 21140 67374
rect 21194 67298 21266 67374
rect 21314 67298 21386 67374
rect 504 66984 576 67060
rect 626 66984 698 67060
rect 752 66984 824 67060
rect 504 66837 576 66913
rect 626 66837 698 66913
rect 752 66837 824 66913
rect 504 66700 576 66776
rect 626 66700 698 66776
rect 752 66700 824 66776
rect 22010 65982 22082 66058
rect 22136 65982 22208 66058
rect 22256 65982 22328 66058
rect 22010 65864 22082 65940
rect 22136 65864 22208 65940
rect 22256 65864 22328 65940
rect 504 65225 576 65301
rect 626 65225 698 65301
rect 752 65225 824 65301
rect 504 65078 576 65154
rect 626 65078 698 65154
rect 752 65078 824 65154
rect 504 64941 576 65017
rect 626 64941 698 65017
rect 752 64941 824 65017
rect 503 64634 575 64710
rect 629 64634 701 64710
rect 749 64634 821 64710
rect 503 64516 575 64592
rect 629 64516 701 64592
rect 749 64516 821 64592
rect 21068 64619 21140 64695
rect 21194 64619 21266 64695
rect 21314 64619 21386 64695
rect 21068 64501 21140 64577
rect 21194 64501 21266 64577
rect 21314 64501 21386 64577
rect 503 63456 575 63532
rect 629 63456 701 63532
rect 749 63456 821 63532
rect 503 63338 575 63414
rect 629 63338 701 63414
rect 749 63338 821 63414
rect 21068 63416 21140 63492
rect 21194 63416 21266 63492
rect 21314 63416 21386 63492
rect 21068 63298 21140 63374
rect 21194 63298 21266 63374
rect 21314 63298 21386 63374
rect 504 62984 576 63060
rect 626 62984 698 63060
rect 752 62984 824 63060
rect 504 62837 576 62913
rect 626 62837 698 62913
rect 752 62837 824 62913
rect 504 62700 576 62776
rect 626 62700 698 62776
rect 752 62700 824 62776
rect 22010 61981 22082 62057
rect 22136 61981 22208 62057
rect 22256 61981 22328 62057
rect 22010 61863 22082 61939
rect 22136 61863 22208 61939
rect 22256 61863 22328 61939
rect 504 61225 576 61301
rect 626 61225 698 61301
rect 752 61225 824 61301
rect 504 61078 576 61154
rect 626 61078 698 61154
rect 752 61078 824 61154
rect 504 60941 576 61017
rect 626 60941 698 61017
rect 752 60941 824 61017
rect 503 60608 575 60684
rect 629 60608 701 60684
rect 749 60608 821 60684
rect 503 60490 575 60566
rect 629 60490 701 60566
rect 749 60490 821 60566
rect 21068 60619 21140 60695
rect 21194 60619 21266 60695
rect 21314 60619 21386 60695
rect 21068 60501 21140 60577
rect 21194 60501 21266 60577
rect 21314 60501 21386 60577
rect 503 59405 575 59481
rect 629 59405 701 59481
rect 749 59405 821 59481
rect 503 59287 575 59363
rect 629 59287 701 59363
rect 749 59287 821 59363
rect 21068 59470 21140 59546
rect 21194 59470 21266 59546
rect 21314 59470 21386 59546
rect 21068 59352 21140 59428
rect 21194 59352 21266 59428
rect 21314 59352 21386 59428
rect 504 58984 576 59060
rect 626 58984 698 59060
rect 752 58984 824 59060
rect 504 58837 576 58913
rect 626 58837 698 58913
rect 752 58837 824 58913
rect 504 58700 576 58776
rect 626 58700 698 58776
rect 752 58700 824 58776
rect 22010 58020 22082 58096
rect 22136 58020 22208 58096
rect 22256 58020 22328 58096
rect 22010 57902 22082 57978
rect 22136 57902 22208 57978
rect 22256 57902 22328 57978
rect 504 57223 576 57299
rect 626 57223 698 57299
rect 752 57223 824 57299
rect 504 57076 576 57152
rect 626 57076 698 57152
rect 752 57076 824 57152
rect 504 56939 576 57015
rect 626 56939 698 57015
rect 752 56939 824 57015
rect 503 56628 575 56704
rect 629 56628 701 56704
rect 749 56628 821 56704
rect 503 56510 575 56586
rect 629 56510 701 56586
rect 749 56510 821 56586
rect 21068 56554 21140 56630
rect 21194 56554 21266 56630
rect 21314 56554 21386 56630
rect 21068 56436 21140 56512
rect 21194 56436 21266 56512
rect 21314 56436 21386 56512
rect 503 55421 575 55497
rect 629 55421 701 55497
rect 749 55421 821 55497
rect 503 55303 575 55379
rect 629 55303 701 55379
rect 749 55303 821 55379
rect 21068 55371 21140 55447
rect 21194 55371 21266 55447
rect 21314 55371 21386 55447
rect 21068 55253 21140 55329
rect 21194 55253 21266 55329
rect 21314 55253 21386 55329
rect 504 54984 576 55060
rect 626 54984 698 55060
rect 752 54984 824 55060
rect 504 54837 576 54913
rect 626 54837 698 54913
rect 752 54837 824 54913
rect 504 54700 576 54776
rect 626 54700 698 54776
rect 752 54700 824 54776
rect 22010 54003 22082 54079
rect 22136 54003 22208 54079
rect 22256 54003 22328 54079
rect 22010 53885 22082 53961
rect 22136 53885 22208 53961
rect 22256 53885 22328 53961
rect 504 53225 576 53301
rect 626 53225 698 53301
rect 752 53225 824 53301
rect 504 53078 576 53154
rect 626 53078 698 53154
rect 752 53078 824 53154
rect 504 52941 576 53017
rect 626 52941 698 53017
rect 752 52941 824 53017
rect 503 52655 575 52731
rect 629 52655 701 52731
rect 749 52655 821 52731
rect 503 52537 575 52613
rect 629 52537 701 52613
rect 749 52537 821 52613
rect 21068 52499 21140 52575
rect 21194 52499 21266 52575
rect 21314 52499 21386 52575
rect 21068 52381 21140 52457
rect 21194 52381 21266 52457
rect 21314 52381 21386 52457
rect 503 51468 575 51544
rect 629 51468 701 51544
rect 749 51468 821 51544
rect 503 51350 575 51426
rect 629 51350 701 51426
rect 749 51350 821 51426
rect 21068 51364 21140 51440
rect 21194 51364 21266 51440
rect 21314 51364 21386 51440
rect 21068 51246 21140 51322
rect 21194 51246 21266 51322
rect 21314 51246 21386 51322
rect 504 50984 576 51060
rect 626 50984 698 51060
rect 752 50984 824 51060
rect 504 50837 576 50913
rect 626 50837 698 50913
rect 752 50837 824 50913
rect 504 50700 576 50776
rect 626 50700 698 50776
rect 752 50700 824 50776
rect 22010 50082 22082 50158
rect 22136 50082 22208 50158
rect 22256 50082 22328 50158
rect 22010 49964 22082 50040
rect 22136 49964 22208 50040
rect 22256 49964 22328 50040
rect 504 49225 576 49301
rect 626 49225 698 49301
rect 752 49225 824 49301
rect 504 49078 576 49154
rect 626 49078 698 49154
rect 752 49078 824 49154
rect 504 48941 576 49017
rect 626 48941 698 49017
rect 752 48941 824 49017
rect 503 48646 575 48722
rect 629 48646 701 48722
rect 749 48646 821 48722
rect 503 48528 575 48604
rect 629 48528 701 48604
rect 749 48528 821 48604
rect 21068 48605 21140 48681
rect 21194 48605 21266 48681
rect 21314 48605 21386 48681
rect 21068 48487 21140 48563
rect 21194 48487 21266 48563
rect 21314 48487 21386 48563
rect 503 47493 575 47569
rect 629 47493 701 47569
rect 749 47493 821 47569
rect 503 47375 575 47451
rect 629 47375 701 47451
rect 749 47375 821 47451
rect 21068 47452 21140 47528
rect 21194 47452 21266 47528
rect 21314 47452 21386 47528
rect 21068 47334 21140 47410
rect 21194 47334 21266 47410
rect 21314 47334 21386 47410
rect 504 46984 576 47060
rect 626 46984 698 47060
rect 752 46984 824 47060
rect 504 46837 576 46913
rect 626 46837 698 46913
rect 752 46837 824 46913
rect 504 46700 576 46776
rect 626 46700 698 46776
rect 752 46700 824 46776
rect 22010 45824 22082 45900
rect 22136 45824 22208 45900
rect 22256 45824 22328 45900
rect 22010 45706 22082 45782
rect 22136 45706 22208 45782
rect 22256 45706 22328 45782
rect 504 45224 576 45300
rect 626 45224 698 45300
rect 752 45224 824 45300
rect 504 45077 576 45153
rect 626 45077 698 45153
rect 752 45077 824 45153
rect 504 44940 576 45016
rect 626 44940 698 45016
rect 752 44940 824 45016
rect 503 44433 575 44509
rect 629 44433 701 44509
rect 749 44433 821 44509
rect 503 44315 575 44391
rect 629 44315 701 44391
rect 749 44315 821 44391
rect 21068 44336 21140 44412
rect 21194 44336 21266 44412
rect 21314 44336 21386 44412
rect 21068 44218 21140 44294
rect 21194 44218 21266 44294
rect 21314 44218 21386 44294
rect 32 39661 112 39741
rect 157 39661 237 39741
rect 282 39661 362 39741
rect 21535 39646 21615 39726
rect 21660 39646 21740 39726
rect 21785 39646 21865 39726
rect 32 39555 112 39635
rect 157 39555 237 39635
rect 282 39555 362 39635
rect 21534 39526 21614 39606
rect 21659 39526 21739 39606
rect 21784 39526 21864 39606
rect 1662 39279 1704 39321
rect 1704 39279 1714 39321
rect 1662 39269 1714 39279
rect 1732 39279 1742 39321
rect 1742 39279 1784 39321
rect 1732 39269 1784 39279
rect 1885 39281 2003 39395
rect 2041 39281 2159 39395
rect 2197 39281 2315 39395
rect 2551 39286 2593 39328
rect 2593 39286 2603 39328
rect 2551 39276 2603 39286
rect 2621 39286 2631 39328
rect 2631 39286 2673 39328
rect 2621 39276 2673 39286
rect 1662 39241 1714 39251
rect 1662 39199 1704 39241
rect 1704 39199 1714 39241
rect 1732 39241 1784 39251
rect 1732 39199 1742 39241
rect 1742 39199 1784 39241
rect 2551 39248 2603 39258
rect 2551 39206 2593 39248
rect 2593 39206 2603 39248
rect 2621 39248 2673 39258
rect 2621 39206 2631 39248
rect 2631 39206 2673 39248
rect 479 39052 561 39130
rect 593 39052 675 39130
rect 707 39052 789 39130
rect 1503 38722 1563 38774
rect 3529 38870 3581 38880
rect 3529 38836 3553 38870
rect 3553 38836 3581 38870
rect 3529 38828 3581 38836
rect 4610 38871 4662 38879
rect 4610 38836 4615 38871
rect 4615 38836 4650 38871
rect 4650 38836 4662 38871
rect 4610 38827 4662 38836
rect 16 38508 98 38586
rect 130 38508 212 38586
rect 244 38508 326 38586
rect 1471 38260 1523 38269
rect 1471 38225 1479 38260
rect 1479 38225 1515 38260
rect 1515 38225 1523 38260
rect 1471 38217 1523 38225
rect 3608 38296 3660 38348
rect 4652 38258 4704 38267
rect 4652 38224 4662 38258
rect 4662 38224 4696 38258
rect 4696 38224 4704 38258
rect 4652 38215 4704 38224
rect 479 37964 561 38042
rect 593 37964 675 38042
rect 707 37964 789 38042
rect 1463 37782 1515 37790
rect 1463 37748 1481 37782
rect 1481 37748 1515 37782
rect 1463 37738 1515 37748
rect 3523 37845 3575 37897
rect 4652 37782 4704 37791
rect 4652 37748 4662 37782
rect 4662 37748 4696 37782
rect 4696 37748 4704 37782
rect 4652 37739 4704 37748
rect 16 37420 98 37498
rect 130 37420 212 37498
rect 244 37420 326 37498
rect 1683 37310 1686 37358
rect 1686 37310 1732 37358
rect 1732 37310 1735 37358
rect 1683 37306 1735 37310
rect 1683 37245 1735 37252
rect 1683 37200 1686 37245
rect 1686 37200 1732 37245
rect 1732 37200 1735 37245
rect 3553 37170 3605 37182
rect 3553 37136 3587 37170
rect 3587 37136 3605 37170
rect 3553 37130 3605 37136
rect 4609 37170 4661 37181
rect 4609 37136 4615 37170
rect 4615 37136 4649 37170
rect 4649 37136 4661 37170
rect 4609 37129 4661 37136
rect 479 36876 561 36954
rect 593 36876 675 36954
rect 707 36876 789 36954
rect 2551 36788 2593 36830
rect 2593 36788 2603 36830
rect 2551 36778 2603 36788
rect 2621 36788 2631 36830
rect 2631 36788 2673 36830
rect 2621 36778 2673 36788
rect 2551 36750 2603 36763
rect 2551 36711 2593 36750
rect 2593 36711 2603 36750
rect 2621 36750 2673 36763
rect 2621 36711 2631 36750
rect 2631 36711 2673 36750
rect 2765 36788 2807 36830
rect 2807 36788 2817 36830
rect 2765 36778 2817 36788
rect 2835 36788 2845 36830
rect 2845 36788 2887 36830
rect 2835 36778 2887 36788
rect 2765 36747 2817 36765
rect 2765 36713 2807 36747
rect 2807 36713 2817 36747
rect 2835 36747 2887 36765
rect 2835 36713 2845 36747
rect 2845 36713 2887 36747
rect 21061 36092 21141 36172
rect 21186 36092 21266 36172
rect 21311 36092 21391 36172
rect 21060 35972 21140 36052
rect 21185 35972 21265 36052
rect 21310 35972 21390 36052
rect 21069 35516 21141 35592
rect 21191 35516 21263 35592
rect 21317 35516 21389 35592
rect 21069 35369 21141 35445
rect 21191 35369 21263 35445
rect 21317 35369 21389 35445
rect 21069 35232 21141 35308
rect 21191 35232 21263 35308
rect 21317 35232 21389 35308
rect 20560 34596 20640 34676
rect 20685 34596 20765 34676
rect 20810 34596 20890 34676
rect 21535 34596 21615 34676
rect 21660 34596 21740 34676
rect 21785 34596 21865 34676
rect 20559 34476 20639 34556
rect 20684 34476 20764 34556
rect 20809 34476 20889 34556
rect 21534 34476 21614 34556
rect 21659 34476 21739 34556
rect 21784 34476 21864 34556
rect 21069 33756 21141 33832
rect 21191 33756 21263 33832
rect 21317 33756 21389 33832
rect 21069 33609 21141 33685
rect 21191 33609 21263 33685
rect 21317 33609 21389 33685
rect 21069 33472 21141 33548
rect 21191 33472 21263 33548
rect 21317 33472 21389 33548
rect 21060 33037 21140 33117
rect 21185 33037 21265 33117
rect 21310 33037 21390 33117
rect 21059 32917 21139 32997
rect 21184 32917 21264 32997
rect 21309 32917 21389 32997
rect 503 32226 575 32302
rect 629 32226 701 32302
rect 749 32226 821 32302
rect 21068 32226 21140 32302
rect 21194 32226 21266 32302
rect 21314 32226 21386 32302
rect 503 32108 575 32184
rect 629 32108 701 32184
rect 749 32108 821 32184
rect 21068 32108 21140 32184
rect 21194 32108 21266 32184
rect 21314 32108 21386 32184
rect 503 31444 575 31520
rect 629 31444 701 31520
rect 749 31444 821 31520
rect 503 31326 575 31402
rect 629 31326 701 31402
rect 749 31326 821 31402
rect 21068 31444 21140 31520
rect 21194 31444 21266 31520
rect 21314 31444 21386 31520
rect 21068 31326 21140 31402
rect 21194 31326 21266 31402
rect 21314 31326 21386 31402
rect 504 30985 576 31061
rect 626 30985 698 31061
rect 752 30985 824 31061
rect 504 30838 576 30914
rect 626 30838 698 30914
rect 752 30838 824 30914
rect 504 30701 576 30777
rect 626 30701 698 30777
rect 752 30701 824 30777
rect 22010 30054 22082 30130
rect 22136 30054 22208 30130
rect 22256 30054 22328 30130
rect 22010 29936 22082 30012
rect 22136 29936 22208 30012
rect 22256 29936 22328 30012
rect 504 29218 576 29294
rect 626 29218 698 29294
rect 752 29218 824 29294
rect 504 29071 576 29147
rect 626 29071 698 29147
rect 752 29071 824 29147
rect 504 28934 576 29010
rect 626 28934 698 29010
rect 752 28934 824 29010
rect 503 28532 575 28608
rect 629 28532 701 28608
rect 749 28532 821 28608
rect 503 28414 575 28490
rect 629 28414 701 28490
rect 749 28414 821 28490
rect 21068 28483 21140 28559
rect 21194 28483 21266 28559
rect 21314 28483 21386 28559
rect 21068 28365 21140 28441
rect 21194 28365 21266 28441
rect 21314 28365 21386 28441
rect 503 27528 575 27604
rect 629 27528 701 27604
rect 749 27528 821 27604
rect 503 27410 575 27486
rect 629 27410 701 27486
rect 749 27410 821 27486
rect 21068 27366 21140 27442
rect 21194 27366 21266 27442
rect 21314 27366 21386 27442
rect 21068 27248 21140 27324
rect 21194 27248 21266 27324
rect 21314 27248 21386 27324
rect 504 26984 576 27060
rect 626 26984 698 27060
rect 752 26984 824 27060
rect 504 26837 576 26913
rect 626 26837 698 26913
rect 752 26837 824 26913
rect 504 26700 576 26776
rect 626 26700 698 26776
rect 752 26700 824 26776
rect 22010 25895 22082 25971
rect 22136 25895 22208 25971
rect 22256 25895 22328 25971
rect 22010 25777 22082 25853
rect 22136 25777 22208 25853
rect 22256 25777 22328 25853
rect 504 25224 576 25300
rect 626 25224 698 25300
rect 752 25224 824 25300
rect 504 25077 576 25153
rect 626 25077 698 25153
rect 752 25077 824 25153
rect 504 24940 576 25016
rect 626 24940 698 25016
rect 752 24940 824 25016
rect 503 24550 575 24626
rect 629 24550 701 24626
rect 749 24550 821 24626
rect 503 24432 575 24508
rect 629 24432 701 24508
rect 749 24432 821 24508
rect 21068 24523 21140 24599
rect 21194 24523 21266 24599
rect 21314 24523 21386 24599
rect 21068 24405 21140 24481
rect 21194 24405 21266 24481
rect 21314 24405 21386 24481
rect 503 23468 575 23544
rect 629 23468 701 23544
rect 749 23468 821 23544
rect 503 23350 575 23426
rect 629 23350 701 23426
rect 749 23350 821 23426
rect 21068 23348 21140 23424
rect 21194 23348 21266 23424
rect 21314 23348 21386 23424
rect 21068 23230 21140 23306
rect 21194 23230 21266 23306
rect 21314 23230 21386 23306
rect 504 22984 576 23060
rect 626 22984 698 23060
rect 752 22984 824 23060
rect 504 22837 576 22913
rect 626 22837 698 22913
rect 752 22837 824 22913
rect 504 22700 576 22776
rect 626 22700 698 22776
rect 752 22700 824 22776
rect 22010 22105 22082 22181
rect 22136 22105 22208 22181
rect 22256 22105 22328 22181
rect 22010 21987 22082 22063
rect 22136 21987 22208 22063
rect 22256 21987 22328 22063
rect 504 21225 576 21301
rect 626 21225 698 21301
rect 752 21225 824 21301
rect 504 21078 576 21154
rect 626 21078 698 21154
rect 752 21078 824 21154
rect 504 20941 576 21017
rect 626 20941 698 21017
rect 752 20941 824 21017
rect 503 20593 575 20669
rect 629 20593 701 20669
rect 749 20593 821 20669
rect 503 20475 575 20551
rect 629 20475 701 20551
rect 749 20475 821 20551
rect 21068 20507 21140 20583
rect 21194 20507 21266 20583
rect 21314 20507 21386 20583
rect 21068 20389 21140 20465
rect 21194 20389 21266 20465
rect 21314 20389 21386 20465
rect 503 19492 575 19568
rect 629 19492 701 19568
rect 749 19492 821 19568
rect 503 19374 575 19450
rect 629 19374 701 19450
rect 749 19374 821 19450
rect 21068 19336 21140 19412
rect 21194 19336 21266 19412
rect 21314 19336 21386 19412
rect 21068 19218 21140 19294
rect 21194 19218 21266 19294
rect 21314 19218 21386 19294
rect 504 18984 576 19060
rect 626 18984 698 19060
rect 752 18984 824 19060
rect 504 18837 576 18913
rect 626 18837 698 18913
rect 752 18837 824 18913
rect 504 18700 576 18776
rect 626 18700 698 18776
rect 752 18700 824 18776
rect 22010 17998 22082 18074
rect 22136 17998 22208 18074
rect 22256 17998 22328 18074
rect 22010 17880 22082 17956
rect 22136 17880 22208 17956
rect 22256 17880 22328 17956
rect 504 17224 576 17300
rect 626 17224 698 17300
rect 752 17224 824 17300
rect 504 17077 576 17153
rect 626 17077 698 17153
rect 752 17077 824 17153
rect 504 16940 576 17016
rect 626 16940 698 17016
rect 752 16940 824 17016
rect 503 16626 575 16702
rect 629 16626 701 16702
rect 749 16626 821 16702
rect 503 16508 575 16584
rect 629 16508 701 16584
rect 749 16508 821 16584
rect 21068 16575 21140 16651
rect 21194 16575 21266 16651
rect 21314 16575 21386 16651
rect 21068 16457 21140 16533
rect 21194 16457 21266 16533
rect 21314 16457 21386 16533
rect 503 15410 575 15486
rect 629 15410 701 15486
rect 749 15410 821 15486
rect 503 15292 575 15368
rect 629 15292 701 15368
rect 749 15292 821 15368
rect 21068 15361 21140 15437
rect 21194 15361 21266 15437
rect 21314 15361 21386 15437
rect 21068 15243 21140 15319
rect 21194 15243 21266 15319
rect 21314 15243 21386 15319
rect 504 14984 576 15060
rect 626 14984 698 15060
rect 752 14984 824 15060
rect 504 14837 576 14913
rect 626 14837 698 14913
rect 752 14837 824 14913
rect 504 14700 576 14776
rect 626 14700 698 14776
rect 752 14700 824 14776
rect 22010 14180 22082 14256
rect 22136 14180 22208 14256
rect 22256 14180 22328 14256
rect 22010 14062 22082 14138
rect 22136 14062 22208 14138
rect 22256 14062 22328 14138
rect 504 13224 576 13300
rect 626 13224 698 13300
rect 752 13224 824 13300
rect 504 13077 576 13153
rect 626 13077 698 13153
rect 752 13077 824 13153
rect 504 12940 576 13016
rect 626 12940 698 13016
rect 752 12940 824 13016
rect 503 12545 575 12621
rect 629 12545 701 12621
rect 749 12545 821 12621
rect 503 12427 575 12503
rect 629 12427 701 12503
rect 749 12427 821 12503
rect 21068 12518 21140 12594
rect 21194 12518 21266 12594
rect 21314 12518 21386 12594
rect 21068 12400 21140 12476
rect 21194 12400 21266 12476
rect 21314 12400 21386 12476
rect 503 11423 575 11499
rect 629 11423 701 11499
rect 749 11423 821 11499
rect 503 11305 575 11381
rect 629 11305 701 11381
rect 749 11305 821 11381
rect 21068 11361 21140 11437
rect 21194 11361 21266 11437
rect 21314 11361 21386 11437
rect 21068 11243 21140 11319
rect 21194 11243 21266 11319
rect 21314 11243 21386 11319
rect 504 10985 576 11061
rect 626 10985 698 11061
rect 752 10985 824 11061
rect 504 10838 576 10914
rect 626 10838 698 10914
rect 752 10838 824 10914
rect 504 10701 576 10777
rect 626 10701 698 10777
rect 752 10701 824 10777
rect 22010 10216 22082 10292
rect 22136 10216 22208 10292
rect 22256 10216 22328 10292
rect 22010 10098 22082 10174
rect 22136 10098 22208 10174
rect 22256 10098 22328 10174
rect 504 9223 576 9299
rect 626 9223 698 9299
rect 752 9223 824 9299
rect 504 9076 576 9152
rect 626 9076 698 9152
rect 752 9076 824 9152
rect 504 8939 576 9015
rect 626 8939 698 9015
rect 752 8939 824 9015
rect 503 8563 575 8639
rect 629 8563 701 8639
rect 749 8563 821 8639
rect 503 8445 575 8521
rect 629 8445 701 8521
rect 749 8445 821 8521
rect 21068 8518 21140 8594
rect 21194 8518 21266 8594
rect 21314 8518 21386 8594
rect 21068 8400 21140 8476
rect 21194 8400 21266 8476
rect 21314 8400 21386 8476
rect 503 7452 575 7528
rect 629 7452 701 7528
rect 749 7452 821 7528
rect 503 7334 575 7410
rect 629 7334 701 7410
rect 749 7334 821 7410
rect 21068 7361 21140 7437
rect 21194 7361 21266 7437
rect 21314 7361 21386 7437
rect 21068 7243 21140 7319
rect 21194 7243 21266 7319
rect 21314 7243 21386 7319
rect 504 6985 576 7061
rect 626 6985 698 7061
rect 752 6985 824 7061
rect 504 6838 576 6914
rect 626 6838 698 6914
rect 752 6838 824 6914
rect 504 6701 576 6777
rect 626 6701 698 6777
rect 752 6701 824 6777
rect 22010 6204 22082 6280
rect 22136 6204 22208 6280
rect 22256 6204 22328 6280
rect 22010 6086 22082 6162
rect 22136 6086 22208 6162
rect 22256 6086 22328 6162
rect 504 5224 576 5300
rect 626 5224 698 5300
rect 752 5224 824 5300
rect 504 5077 576 5153
rect 626 5077 698 5153
rect 752 5077 824 5153
rect 504 4940 576 5016
rect 626 4940 698 5016
rect 752 4940 824 5016
rect 503 4629 575 4705
rect 629 4629 701 4705
rect 749 4629 821 4705
rect 503 4511 575 4587
rect 629 4511 701 4587
rect 749 4511 821 4587
rect 21068 4518 21140 4594
rect 21194 4518 21266 4594
rect 21314 4518 21386 4594
rect 21068 4400 21140 4476
rect 21194 4400 21266 4476
rect 21314 4400 21386 4476
rect 503 3452 575 3528
rect 629 3452 701 3528
rect 749 3452 821 3528
rect 503 3334 575 3410
rect 629 3334 701 3410
rect 749 3334 821 3410
rect 21068 3361 21140 3437
rect 21194 3361 21266 3437
rect 21314 3361 21386 3437
rect 21068 3243 21140 3319
rect 21194 3243 21266 3319
rect 21314 3243 21386 3319
rect 504 2985 576 3061
rect 626 2985 698 3061
rect 752 2985 824 3061
rect 504 2838 576 2914
rect 626 2838 698 2914
rect 752 2838 824 2914
rect 504 2701 576 2777
rect 626 2701 698 2777
rect 752 2701 824 2777
rect 22010 2204 22082 2280
rect 22136 2204 22208 2280
rect 22256 2204 22328 2280
rect 22010 2086 22082 2162
rect 22136 2086 22208 2162
rect 22256 2086 22328 2162
rect 504 1224 576 1300
rect 626 1224 698 1300
rect 752 1224 824 1300
rect 504 1077 576 1153
rect 626 1077 698 1153
rect 752 1077 824 1153
rect 504 940 576 1016
rect 626 940 698 1016
rect 752 940 824 1016
rect 503 629 575 705
rect 629 629 701 705
rect 749 629 821 705
rect 503 511 575 587
rect 629 511 701 587
rect 749 511 821 587
rect 21068 518 21140 594
rect 21194 518 21266 594
rect 21314 518 21386 594
rect 21068 400 21140 476
rect 21194 400 21266 476
rect 21314 400 21386 476
<< metal2 >>
rect 21026 75492 21426 75517
rect 463 75452 864 75477
rect 463 75376 503 75452
rect 575 75376 629 75452
rect 701 75376 749 75452
rect 821 75376 864 75452
rect 463 75334 864 75376
rect 463 75258 503 75334
rect 575 75258 629 75334
rect 701 75258 749 75334
rect 821 75258 864 75334
rect 21026 75416 21068 75492
rect 21140 75416 21194 75492
rect 21266 75416 21314 75492
rect 21386 75416 21426 75492
rect 21026 75374 21426 75416
rect 21026 75298 21068 75374
rect 21140 75298 21194 75374
rect 21266 75298 21314 75374
rect 21386 75298 21426 75374
rect 21026 75262 21426 75298
rect 463 75222 864 75258
rect 463 75060 863 75109
rect 463 74984 504 75060
rect 576 74984 626 75060
rect 698 74984 752 75060
rect 824 74984 863 75060
rect 463 74913 863 74984
rect 463 74837 504 74913
rect 576 74837 626 74913
rect 698 74837 752 74913
rect 824 74837 863 74913
rect 463 74776 863 74837
rect 463 74700 504 74776
rect 576 74700 626 74776
rect 698 74700 752 74776
rect 824 74700 863 74776
rect 463 74650 863 74700
rect 21970 74071 22370 74096
rect 21970 73995 22010 74071
rect 22082 73995 22136 74071
rect 22208 73995 22256 74071
rect 22328 73995 22370 74071
rect 21970 73953 22370 73995
rect 21970 73877 22010 73953
rect 22082 73877 22136 73953
rect 22208 73877 22256 73953
rect 22328 73877 22370 73953
rect 21970 73841 22370 73877
rect 463 73300 863 73349
rect 463 73224 504 73300
rect 576 73224 626 73300
rect 698 73224 752 73300
rect 824 73224 863 73300
rect 463 73153 863 73224
rect 463 73077 504 73153
rect 576 73077 626 73153
rect 698 73077 752 73153
rect 824 73077 863 73153
rect 463 73016 863 73077
rect 463 72940 504 73016
rect 576 72940 626 73016
rect 698 72940 752 73016
rect 824 72940 863 73016
rect 463 72890 863 72940
rect 463 72779 864 72804
rect 463 72703 503 72779
rect 575 72703 629 72779
rect 701 72703 749 72779
rect 821 72703 864 72779
rect 463 72661 864 72703
rect 463 72585 503 72661
rect 575 72585 629 72661
rect 701 72585 749 72661
rect 821 72585 864 72661
rect 463 72549 864 72585
rect 21028 72695 21428 72720
rect 21028 72619 21068 72695
rect 21140 72619 21194 72695
rect 21266 72619 21314 72695
rect 21386 72619 21428 72695
rect 21028 72577 21428 72619
rect 21028 72501 21068 72577
rect 21140 72501 21194 72577
rect 21266 72501 21314 72577
rect 21386 72501 21428 72577
rect 21028 72465 21428 72501
rect 21026 71492 21426 71517
rect 463 71452 864 71477
rect 463 71376 503 71452
rect 575 71376 629 71452
rect 701 71376 749 71452
rect 821 71376 864 71452
rect 463 71334 864 71376
rect 463 71258 503 71334
rect 575 71258 629 71334
rect 701 71258 749 71334
rect 821 71258 864 71334
rect 21026 71416 21068 71492
rect 21140 71416 21194 71492
rect 21266 71416 21314 71492
rect 21386 71416 21426 71492
rect 21026 71374 21426 71416
rect 21026 71298 21068 71374
rect 21140 71298 21194 71374
rect 21266 71298 21314 71374
rect 21386 71298 21426 71374
rect 21026 71262 21426 71298
rect 463 71222 864 71258
rect 463 71060 863 71109
rect 463 70984 504 71060
rect 576 70984 626 71060
rect 698 70984 752 71060
rect 824 70984 863 71060
rect 463 70913 863 70984
rect 463 70837 504 70913
rect 576 70837 626 70913
rect 698 70837 752 70913
rect 824 70837 863 70913
rect 463 70776 863 70837
rect 463 70700 504 70776
rect 576 70700 626 70776
rect 698 70700 752 70776
rect 824 70700 863 70776
rect 463 70650 863 70700
rect 21970 70071 22370 70096
rect 21970 69995 22010 70071
rect 22082 69995 22136 70071
rect 22208 69995 22256 70071
rect 22328 69995 22370 70071
rect 21970 69953 22370 69995
rect 21970 69877 22010 69953
rect 22082 69877 22136 69953
rect 22208 69877 22256 69953
rect 22328 69877 22370 69953
rect 21970 69841 22370 69877
rect 463 69300 863 69349
rect 463 69224 504 69300
rect 576 69224 626 69300
rect 698 69224 752 69300
rect 824 69224 863 69300
rect 463 69153 863 69224
rect 463 69077 504 69153
rect 576 69077 626 69153
rect 698 69077 752 69153
rect 824 69077 863 69153
rect 463 69016 863 69077
rect 463 68940 504 69016
rect 576 68940 626 69016
rect 698 68940 752 69016
rect 824 68940 863 69016
rect 463 68890 863 68940
rect 463 68779 864 68804
rect 463 68703 503 68779
rect 575 68703 629 68779
rect 701 68703 749 68779
rect 821 68703 864 68779
rect 463 68661 864 68703
rect 463 68585 503 68661
rect 575 68585 629 68661
rect 701 68585 749 68661
rect 821 68585 864 68661
rect 463 68549 864 68585
rect 21028 68695 21428 68720
rect 21028 68619 21068 68695
rect 21140 68619 21194 68695
rect 21266 68619 21314 68695
rect 21386 68619 21428 68695
rect 21028 68577 21428 68619
rect 21028 68501 21068 68577
rect 21140 68501 21194 68577
rect 21266 68501 21314 68577
rect 21386 68501 21428 68577
rect 21028 68465 21428 68501
rect 21026 67492 21426 67517
rect 463 67450 864 67475
rect 463 67374 503 67450
rect 575 67374 629 67450
rect 701 67374 749 67450
rect 821 67374 864 67450
rect 463 67332 864 67374
rect 463 67256 503 67332
rect 575 67256 629 67332
rect 701 67256 749 67332
rect 821 67256 864 67332
rect 21026 67416 21068 67492
rect 21140 67416 21194 67492
rect 21266 67416 21314 67492
rect 21386 67416 21426 67492
rect 21026 67374 21426 67416
rect 21026 67298 21068 67374
rect 21140 67298 21194 67374
rect 21266 67298 21314 67374
rect 21386 67298 21426 67374
rect 21026 67262 21426 67298
rect 463 67220 864 67256
rect 463 67060 863 67109
rect 463 66984 504 67060
rect 576 66984 626 67060
rect 698 66984 752 67060
rect 824 66984 863 67060
rect 463 66913 863 66984
rect 463 66837 504 66913
rect 576 66837 626 66913
rect 698 66837 752 66913
rect 824 66837 863 66913
rect 463 66776 863 66837
rect 463 66700 504 66776
rect 576 66700 626 66776
rect 698 66700 752 66776
rect 824 66700 863 66776
rect 463 66650 863 66700
rect 21970 66058 22370 66083
rect 21970 65982 22010 66058
rect 22082 65982 22136 66058
rect 22208 65982 22256 66058
rect 22328 65982 22370 66058
rect 21970 65940 22370 65982
rect 21970 65864 22010 65940
rect 22082 65864 22136 65940
rect 22208 65864 22256 65940
rect 22328 65864 22370 65940
rect 21970 65828 22370 65864
rect 463 65301 863 65350
rect 463 65225 504 65301
rect 576 65225 626 65301
rect 698 65225 752 65301
rect 824 65225 863 65301
rect 463 65154 863 65225
rect 463 65078 504 65154
rect 576 65078 626 65154
rect 698 65078 752 65154
rect 824 65078 863 65154
rect 463 65017 863 65078
rect 463 64941 504 65017
rect 576 64941 626 65017
rect 698 64941 752 65017
rect 824 64941 863 65017
rect 463 64891 863 64941
rect 463 64710 864 64735
rect 463 64634 503 64710
rect 575 64634 629 64710
rect 701 64634 749 64710
rect 821 64634 864 64710
rect 463 64592 864 64634
rect 463 64516 503 64592
rect 575 64516 629 64592
rect 701 64516 749 64592
rect 821 64516 864 64592
rect 463 64480 864 64516
rect 21028 64695 21428 64720
rect 21028 64619 21068 64695
rect 21140 64619 21194 64695
rect 21266 64619 21314 64695
rect 21386 64619 21428 64695
rect 21028 64577 21428 64619
rect 21028 64501 21068 64577
rect 21140 64501 21194 64577
rect 21266 64501 21314 64577
rect 21386 64501 21428 64577
rect 21028 64465 21428 64501
rect 463 63532 864 63557
rect 463 63456 503 63532
rect 575 63456 629 63532
rect 701 63456 749 63532
rect 821 63456 864 63532
rect 463 63414 864 63456
rect 463 63338 503 63414
rect 575 63338 629 63414
rect 701 63338 749 63414
rect 821 63338 864 63414
rect 463 63302 864 63338
rect 21026 63492 21426 63517
rect 21026 63416 21068 63492
rect 21140 63416 21194 63492
rect 21266 63416 21314 63492
rect 21386 63416 21426 63492
rect 21026 63374 21426 63416
rect 21026 63298 21068 63374
rect 21140 63298 21194 63374
rect 21266 63298 21314 63374
rect 21386 63298 21426 63374
rect 21026 63262 21426 63298
rect 464 63068 864 63109
rect 463 63060 864 63068
rect 463 62984 504 63060
rect 576 62984 626 63060
rect 698 62984 752 63060
rect 824 62984 864 63060
rect 463 62913 864 62984
rect 463 62837 504 62913
rect 576 62837 626 62913
rect 698 62837 752 62913
rect 824 62837 864 62913
rect 463 62776 864 62837
rect 463 62700 504 62776
rect 576 62700 626 62776
rect 698 62700 752 62776
rect 824 62700 864 62776
rect 463 62650 864 62700
rect 21970 62057 22370 62082
rect 21970 61981 22010 62057
rect 22082 61981 22136 62057
rect 22208 61981 22256 62057
rect 22328 61981 22370 62057
rect 21970 61939 22370 61981
rect 21970 61863 22010 61939
rect 22082 61863 22136 61939
rect 22208 61863 22256 61939
rect 22328 61863 22370 61939
rect 21970 61827 22370 61863
rect 463 61301 863 61350
rect 463 61225 504 61301
rect 576 61225 626 61301
rect 698 61225 752 61301
rect 824 61225 863 61301
rect 463 61154 863 61225
rect 463 61078 504 61154
rect 576 61078 626 61154
rect 698 61078 752 61154
rect 824 61078 863 61154
rect 463 61017 863 61078
rect 463 60941 504 61017
rect 576 60941 626 61017
rect 698 60941 752 61017
rect 824 60941 863 61017
rect 463 60891 863 60941
rect 463 60684 866 60709
rect 463 60608 503 60684
rect 575 60608 629 60684
rect 701 60608 749 60684
rect 821 60608 866 60684
rect 463 60566 866 60608
rect 463 60490 503 60566
rect 575 60490 629 60566
rect 701 60490 749 60566
rect 821 60490 866 60566
rect 463 60454 866 60490
rect 21028 60695 21428 60720
rect 21028 60619 21068 60695
rect 21140 60619 21194 60695
rect 21266 60619 21314 60695
rect 21386 60619 21428 60695
rect 21028 60577 21428 60619
rect 21028 60501 21068 60577
rect 21140 60501 21194 60577
rect 21266 60501 21314 60577
rect 21386 60501 21428 60577
rect 21028 60465 21428 60501
rect 21027 59546 21427 59571
rect 463 59481 864 59506
rect 463 59405 503 59481
rect 575 59405 629 59481
rect 701 59405 749 59481
rect 821 59405 864 59481
rect 463 59363 864 59405
rect 463 59287 503 59363
rect 575 59287 629 59363
rect 701 59287 749 59363
rect 821 59287 864 59363
rect 21027 59470 21068 59546
rect 21140 59470 21194 59546
rect 21266 59470 21314 59546
rect 21386 59470 21427 59546
rect 21027 59428 21427 59470
rect 21027 59352 21068 59428
rect 21140 59352 21194 59428
rect 21266 59352 21314 59428
rect 21386 59352 21427 59428
rect 21027 59316 21427 59352
rect 463 59251 864 59287
rect 464 59068 864 59109
rect 463 59060 864 59068
rect 463 58984 504 59060
rect 576 58984 626 59060
rect 698 58984 752 59060
rect 824 58984 864 59060
rect 463 58913 864 58984
rect 463 58837 504 58913
rect 576 58837 626 58913
rect 698 58837 752 58913
rect 824 58837 864 58913
rect 463 58776 864 58837
rect 463 58700 504 58776
rect 576 58700 626 58776
rect 698 58700 752 58776
rect 824 58700 864 58776
rect 463 58650 864 58700
rect 21970 58096 22370 58121
rect 21970 58020 22010 58096
rect 22082 58020 22136 58096
rect 22208 58020 22256 58096
rect 22328 58020 22370 58096
rect 21970 57978 22370 58020
rect 21970 57902 22010 57978
rect 22082 57902 22136 57978
rect 22208 57902 22256 57978
rect 22328 57902 22370 57978
rect 21970 57866 22370 57902
rect 463 57299 863 57348
rect 463 57223 504 57299
rect 576 57223 626 57299
rect 698 57223 752 57299
rect 824 57223 863 57299
rect 463 57152 863 57223
rect 463 57076 504 57152
rect 576 57076 626 57152
rect 698 57076 752 57152
rect 824 57076 863 57152
rect 463 57015 863 57076
rect 463 56939 504 57015
rect 576 56939 626 57015
rect 698 56939 752 57015
rect 824 56939 863 57015
rect 463 56889 863 56939
rect 463 56704 864 56729
rect 463 56628 503 56704
rect 575 56628 629 56704
rect 701 56628 749 56704
rect 821 56628 864 56704
rect 463 56586 864 56628
rect 463 56510 503 56586
rect 575 56510 629 56586
rect 701 56510 749 56586
rect 821 56510 864 56586
rect 463 56474 864 56510
rect 21028 56630 21428 56655
rect 21028 56554 21068 56630
rect 21140 56554 21194 56630
rect 21266 56554 21314 56630
rect 21386 56554 21428 56630
rect 21028 56512 21428 56554
rect 21028 56436 21068 56512
rect 21140 56436 21194 56512
rect 21266 56436 21314 56512
rect 21386 56436 21428 56512
rect 21028 56400 21428 56436
rect 463 55497 866 55522
rect 463 55421 503 55497
rect 575 55421 629 55497
rect 701 55421 749 55497
rect 821 55421 866 55497
rect 463 55379 866 55421
rect 463 55303 503 55379
rect 575 55303 629 55379
rect 701 55303 749 55379
rect 821 55303 866 55379
rect 463 55267 866 55303
rect 21027 55447 21427 55472
rect 21027 55371 21068 55447
rect 21140 55371 21194 55447
rect 21266 55371 21314 55447
rect 21386 55371 21427 55447
rect 21027 55329 21427 55371
rect 21027 55253 21068 55329
rect 21140 55253 21194 55329
rect 21266 55253 21314 55329
rect 21386 55253 21427 55329
rect 21027 55217 21427 55253
rect 463 55060 863 55109
rect 463 54984 504 55060
rect 576 54984 626 55060
rect 698 54984 752 55060
rect 824 54984 863 55060
rect 463 54913 863 54984
rect 463 54837 504 54913
rect 576 54837 626 54913
rect 698 54837 752 54913
rect 824 54837 863 54913
rect 463 54776 863 54837
rect 463 54700 504 54776
rect 576 54700 626 54776
rect 698 54700 752 54776
rect 824 54700 863 54776
rect 463 54650 863 54700
rect 21970 54079 22370 54104
rect 21970 54003 22010 54079
rect 22082 54003 22136 54079
rect 22208 54003 22256 54079
rect 22328 54003 22370 54079
rect 21970 53961 22370 54003
rect 21970 53885 22010 53961
rect 22082 53885 22136 53961
rect 22208 53885 22256 53961
rect 22328 53885 22370 53961
rect 21970 53849 22370 53885
rect 463 53301 863 53350
rect 463 53225 504 53301
rect 576 53225 626 53301
rect 698 53225 752 53301
rect 824 53225 863 53301
rect 463 53154 863 53225
rect 463 53078 504 53154
rect 576 53078 626 53154
rect 698 53078 752 53154
rect 824 53078 863 53154
rect 463 53017 863 53078
rect 463 52941 504 53017
rect 576 52941 626 53017
rect 698 52941 752 53017
rect 824 52941 863 53017
rect 463 52891 863 52941
rect 463 52731 864 52756
rect 463 52655 503 52731
rect 575 52655 629 52731
rect 701 52655 749 52731
rect 821 52655 864 52731
rect 463 52613 864 52655
rect 463 52537 503 52613
rect 575 52537 629 52613
rect 701 52537 749 52613
rect 821 52537 864 52613
rect 463 52501 864 52537
rect 21028 52575 21428 52600
rect 21028 52499 21068 52575
rect 21140 52499 21194 52575
rect 21266 52499 21314 52575
rect 21386 52499 21428 52575
rect 21028 52457 21428 52499
rect 21028 52381 21068 52457
rect 21140 52381 21194 52457
rect 21266 52381 21314 52457
rect 21386 52381 21428 52457
rect 21028 52345 21428 52381
rect 463 51544 864 51569
rect 463 51468 503 51544
rect 575 51468 629 51544
rect 701 51468 749 51544
rect 821 51468 864 51544
rect 463 51426 864 51468
rect 463 51350 503 51426
rect 575 51350 629 51426
rect 701 51350 749 51426
rect 821 51350 864 51426
rect 463 51314 864 51350
rect 21028 51440 21428 51465
rect 21028 51364 21068 51440
rect 21140 51364 21194 51440
rect 21266 51364 21314 51440
rect 21386 51364 21428 51440
rect 21028 51322 21428 51364
rect 21028 51246 21068 51322
rect 21140 51246 21194 51322
rect 21266 51246 21314 51322
rect 21386 51246 21428 51322
rect 21028 51210 21428 51246
rect 463 51060 863 51109
rect 463 50984 504 51060
rect 576 50984 626 51060
rect 698 50984 752 51060
rect 824 50984 863 51060
rect 463 50913 863 50984
rect 463 50837 504 50913
rect 576 50837 626 50913
rect 698 50837 752 50913
rect 824 50837 863 50913
rect 463 50776 863 50837
rect 463 50700 504 50776
rect 576 50700 626 50776
rect 698 50700 752 50776
rect 824 50700 863 50776
rect 463 50650 863 50700
rect 21970 50158 22370 50183
rect 21970 50082 22010 50158
rect 22082 50082 22136 50158
rect 22208 50082 22256 50158
rect 22328 50082 22370 50158
rect 21970 50040 22370 50082
rect 21970 49964 22010 50040
rect 22082 49964 22136 50040
rect 22208 49964 22256 50040
rect 22328 49964 22370 50040
rect 21970 49928 22370 49964
rect 463 49301 863 49350
rect 463 49225 504 49301
rect 576 49225 626 49301
rect 698 49225 752 49301
rect 824 49225 863 49301
rect 463 49154 863 49225
rect 463 49078 504 49154
rect 576 49078 626 49154
rect 698 49078 752 49154
rect 824 49078 863 49154
rect 463 49017 863 49078
rect 463 48941 504 49017
rect 576 48941 626 49017
rect 698 48941 752 49017
rect 824 48941 863 49017
rect 463 48891 863 48941
rect 463 48722 864 48747
rect 463 48646 503 48722
rect 575 48646 629 48722
rect 701 48646 749 48722
rect 821 48646 864 48722
rect 463 48604 864 48646
rect 463 48528 503 48604
rect 575 48528 629 48604
rect 701 48528 749 48604
rect 821 48528 864 48604
rect 463 48492 864 48528
rect 21028 48681 21428 48706
rect 21028 48605 21068 48681
rect 21140 48605 21194 48681
rect 21266 48605 21314 48681
rect 21386 48605 21428 48681
rect 21028 48563 21428 48605
rect 21028 48487 21068 48563
rect 21140 48487 21194 48563
rect 21266 48487 21314 48563
rect 21386 48487 21428 48563
rect 21028 48451 21428 48487
rect 463 47569 864 47594
rect 463 47493 503 47569
rect 575 47493 629 47569
rect 701 47493 749 47569
rect 821 47493 864 47569
rect 463 47451 864 47493
rect 463 47375 503 47451
rect 575 47375 629 47451
rect 701 47375 749 47451
rect 821 47375 864 47451
rect 463 47339 864 47375
rect 21028 47528 21428 47553
rect 21028 47452 21068 47528
rect 21140 47452 21194 47528
rect 21266 47452 21314 47528
rect 21386 47452 21428 47528
rect 21028 47410 21428 47452
rect 21028 47334 21068 47410
rect 21140 47334 21194 47410
rect 21266 47334 21314 47410
rect 21386 47334 21428 47410
rect 21028 47298 21428 47334
rect 463 47060 863 47109
rect 463 46984 504 47060
rect 576 46984 626 47060
rect 698 46984 752 47060
rect 824 46984 863 47060
rect 463 46913 863 46984
rect 463 46837 504 46913
rect 576 46837 626 46913
rect 698 46837 752 46913
rect 824 46837 863 46913
rect 463 46776 863 46837
rect 463 46700 504 46776
rect 576 46700 626 46776
rect 698 46700 752 46776
rect 824 46700 863 46776
rect 463 46650 863 46700
rect 21970 45900 22370 45925
rect 21970 45824 22010 45900
rect 22082 45824 22136 45900
rect 22208 45824 22256 45900
rect 22328 45824 22370 45900
rect 21970 45782 22370 45824
rect 21970 45706 22010 45782
rect 22082 45706 22136 45782
rect 22208 45706 22256 45782
rect 22328 45706 22370 45782
rect 21970 45670 22370 45706
rect 463 45300 863 45350
rect 463 45224 504 45300
rect 576 45224 626 45300
rect 698 45224 752 45300
rect 824 45224 863 45300
rect 463 45153 863 45224
rect 463 45077 504 45153
rect 576 45077 626 45153
rect 698 45077 752 45153
rect 824 45077 863 45153
rect 463 45016 863 45077
rect 463 44940 504 45016
rect 576 44940 626 45016
rect 698 44940 752 45016
rect 824 44940 863 45016
rect 463 44891 863 44940
rect 463 44890 836 44891
rect 463 44509 863 44534
rect 463 44433 503 44509
rect 575 44433 629 44509
rect 701 44433 749 44509
rect 821 44433 863 44509
rect 463 44391 863 44433
rect 463 44315 503 44391
rect 575 44315 629 44391
rect 701 44315 749 44391
rect 821 44315 863 44391
rect 463 44279 863 44315
rect 21028 44412 21428 44437
rect 21028 44336 21068 44412
rect 21140 44336 21194 44412
rect 21266 44336 21314 44412
rect 21386 44336 21428 44412
rect 21028 44294 21428 44336
rect 21028 44218 21068 44294
rect 21140 44218 21194 44294
rect 21266 44218 21314 44294
rect 21386 44218 21428 44294
rect 21028 44182 21428 44218
rect 1650 39925 2398 39940
rect 1650 39869 2257 39925
rect 2313 39869 2337 39925
rect 2393 39869 2398 39925
rect 1650 39845 2398 39869
rect 1650 39789 2257 39845
rect 2313 39789 2337 39845
rect 2393 39789 2398 39845
rect 1650 39776 2398 39789
rect 1650 39774 2396 39776
rect 0 39741 400 39752
rect 0 39661 32 39741
rect 112 39661 157 39741
rect 237 39661 282 39741
rect 362 39661 400 39741
rect 0 39635 400 39661
rect 0 39555 32 39635
rect 112 39555 157 39635
rect 237 39555 282 39635
rect 362 39555 400 39635
rect 0 39528 400 39555
rect 1411 39320 1569 39333
rect 1411 39319 1498 39320
rect 1411 39263 1416 39319
rect 1472 39264 1498 39319
rect 1554 39264 1569 39320
rect 1472 39263 1569 39264
rect 1411 39240 1569 39263
rect 1411 39239 1499 39240
rect 1411 39183 1417 39239
rect 1473 39184 1499 39239
rect 1555 39184 1569 39240
rect 1650 39321 1796 39774
rect 2468 39711 2867 44000
rect 21970 43838 22370 43870
rect 21970 43514 22006 43838
rect 22298 43514 22370 43838
rect 21970 43480 22370 43514
rect 3352 39904 3502 39919
rect 3352 39848 3361 39904
rect 3417 39848 3441 39904
rect 3497 39848 3502 39904
rect 3352 39824 3502 39848
rect 3352 39768 3361 39824
rect 3417 39768 3441 39824
rect 3497 39768 3502 39824
rect 3352 39755 3502 39768
rect 3352 39754 3500 39755
rect 1867 39438 2868 39711
rect 1650 39269 1662 39321
rect 1714 39269 1732 39321
rect 1784 39269 1796 39321
rect 1650 39251 1796 39269
rect 1650 39199 1662 39251
rect 1714 39199 1732 39251
rect 1784 39199 1796 39251
rect 1650 39189 1796 39199
rect 1868 39410 2267 39438
rect 1868 39395 2335 39410
rect 1868 39281 1885 39395
rect 2003 39281 2041 39395
rect 2159 39281 2197 39395
rect 2315 39281 2335 39395
rect 1868 39270 2335 39281
rect 2538 39328 2685 39336
rect 2538 39276 2551 39328
rect 2603 39276 2621 39328
rect 2673 39276 2685 39328
rect 1473 39183 1569 39184
rect 1411 39169 1569 39183
rect 463 39130 805 39139
rect 463 39052 479 39130
rect 561 39052 593 39130
rect 675 39052 707 39130
rect 789 39052 805 39130
rect 463 39043 805 39052
rect 1495 38774 1569 39169
rect 1495 38722 1503 38774
rect 1563 38722 1569 38774
rect 1495 38717 1569 38722
rect 0 38586 342 38595
rect 0 38508 16 38586
rect 98 38508 130 38586
rect 212 38508 244 38586
rect 326 38508 342 38586
rect 0 38499 342 38508
rect 1471 38269 1523 38275
rect 1471 38211 1523 38217
rect 463 38042 805 38051
rect 463 37964 479 38042
rect 561 37964 593 38042
rect 675 37964 707 38042
rect 789 37964 805 38042
rect 463 37955 805 37964
rect 1471 37797 1504 38211
rect 1463 37790 1515 37797
rect 1463 37732 1515 37738
rect 0 37498 342 37507
rect 0 37420 16 37498
rect 98 37420 130 37498
rect 212 37420 244 37498
rect 326 37420 342 37498
rect 0 37411 342 37420
rect 1680 37358 1739 39189
rect 1680 37306 1683 37358
rect 1735 37306 1739 37358
rect 1680 37252 1739 37306
rect 1680 37200 1683 37252
rect 1735 37200 1739 37252
rect 1680 37187 1739 37200
rect 463 36954 805 36963
rect 463 36876 479 36954
rect 561 36876 593 36954
rect 675 36876 707 36954
rect 789 36876 805 36954
rect 463 36867 805 36876
rect 1868 32936 2267 39270
rect 2538 39258 2685 39276
rect 2538 39206 2551 39258
rect 2603 39206 2621 39258
rect 2673 39206 2685 39258
rect 2751 39318 2899 39332
rect 2751 39262 2760 39318
rect 2816 39317 2899 39318
rect 2816 39262 2840 39317
rect 2751 39261 2840 39262
rect 2896 39261 2899 39317
rect 2751 39253 2899 39261
rect 2538 36830 2685 39206
rect 2538 36778 2551 36830
rect 2603 36778 2621 36830
rect 2673 36778 2685 36830
rect 2538 36763 2685 36778
rect 2538 36711 2551 36763
rect 2603 36711 2621 36763
rect 2673 36711 2685 36763
rect 2538 36476 2685 36711
rect 2752 39237 2899 39253
rect 2752 39181 2761 39237
rect 2817 39181 2841 39237
rect 2897 39181 2899 39237
rect 2752 36830 2899 39181
rect 3352 39317 3499 39754
rect 21502 39726 21902 39752
rect 21502 39646 21535 39726
rect 21615 39646 21660 39726
rect 21740 39646 21785 39726
rect 21865 39646 21902 39726
rect 21502 39606 21902 39646
rect 21502 39526 21534 39606
rect 21614 39526 21659 39606
rect 21739 39526 21784 39606
rect 21864 39526 21902 39606
rect 21502 39497 21902 39526
rect 3352 39261 3360 39317
rect 3416 39316 3499 39317
rect 3416 39261 3440 39316
rect 3352 39260 3440 39261
rect 3496 39260 3499 39316
rect 3352 39236 3499 39260
rect 3352 39180 3361 39236
rect 3417 39180 3441 39236
rect 3497 39180 3499 39236
rect 3352 39169 3499 39180
rect 3523 38828 3529 38880
rect 3581 38828 3587 38880
rect 4610 38879 4704 38885
rect 3537 37897 3568 38828
rect 4662 38827 4704 38879
rect 4610 38821 4704 38827
rect 3608 38348 3660 38354
rect 3608 38290 3660 38296
rect 3517 37845 3523 37897
rect 3575 37845 3581 37897
rect 3620 37185 3649 38290
rect 4652 38267 4704 38821
rect 4652 38209 4704 38215
rect 4652 37791 4704 37797
rect 4652 37187 4704 37739
rect 3536 37182 3649 37185
rect 3536 37130 3553 37182
rect 3605 37130 3649 37182
rect 3536 37126 3649 37130
rect 4609 37181 4704 37187
rect 4661 37129 4704 37181
rect 4609 37123 4704 37129
rect 2752 36778 2765 36830
rect 2817 36778 2835 36830
rect 2887 36778 2899 36830
rect 2752 36765 2899 36778
rect 2752 36713 2765 36765
rect 2817 36713 2835 36765
rect 2887 36713 2899 36765
rect 2752 36707 2899 36713
rect 21970 36954 22370 36986
rect 21970 36630 22006 36954
rect 22298 36630 22370 36954
rect 21970 36596 22370 36630
rect 2535 36475 2685 36476
rect 2535 36463 2689 36475
rect 2535 36401 2544 36463
rect 2600 36401 2624 36463
rect 2680 36401 2689 36463
rect 2535 36391 2689 36401
rect 21028 36172 21428 36198
rect 21028 36092 21061 36172
rect 21141 36092 21186 36172
rect 21266 36092 21311 36172
rect 21391 36092 21428 36172
rect 21028 36052 21428 36092
rect 21028 35972 21060 36052
rect 21140 35972 21185 36052
rect 21265 35972 21310 36052
rect 21390 35972 21428 36052
rect 21028 35943 21428 35972
rect 21028 35592 21428 35642
rect 21028 35516 21069 35592
rect 21141 35516 21191 35592
rect 21263 35516 21317 35592
rect 21389 35516 21428 35592
rect 21028 35445 21428 35516
rect 21028 35369 21069 35445
rect 21141 35369 21191 35445
rect 21263 35369 21317 35445
rect 21389 35369 21428 35445
rect 21028 35308 21428 35369
rect 21028 35232 21069 35308
rect 21141 35232 21191 35308
rect 21263 35232 21317 35308
rect 21389 35232 21428 35308
rect 21028 35183 21428 35232
rect 21028 35182 21401 35183
rect 20527 34676 20927 34702
rect 20527 34596 20560 34676
rect 20640 34596 20685 34676
rect 20765 34596 20810 34676
rect 20890 34596 20927 34676
rect 20527 34556 20927 34596
rect 20527 34476 20559 34556
rect 20639 34476 20684 34556
rect 20764 34476 20809 34556
rect 20889 34476 20927 34556
rect 20527 34447 20927 34476
rect 21502 34676 21902 34702
rect 21502 34596 21535 34676
rect 21615 34596 21660 34676
rect 21740 34596 21785 34676
rect 21865 34596 21902 34676
rect 21502 34556 21902 34596
rect 21502 34476 21534 34556
rect 21614 34476 21659 34556
rect 21739 34476 21784 34556
rect 21864 34476 21902 34556
rect 21502 34447 21902 34476
rect 21028 33832 21428 33882
rect 21028 33756 21069 33832
rect 21141 33756 21191 33832
rect 21263 33756 21317 33832
rect 21389 33756 21428 33832
rect 21028 33685 21428 33756
rect 21028 33609 21069 33685
rect 21141 33609 21191 33685
rect 21263 33609 21317 33685
rect 21389 33609 21428 33685
rect 21028 33548 21428 33609
rect 21028 33472 21069 33548
rect 21141 33472 21191 33548
rect 21263 33472 21317 33548
rect 21389 33472 21428 33548
rect 21028 33423 21428 33472
rect 21028 33422 21401 33423
rect 21027 33117 21427 33143
rect 21027 33037 21060 33117
rect 21140 33037 21185 33117
rect 21265 33037 21310 33117
rect 21390 33037 21427 33117
rect 21027 32997 21427 33037
rect 1868 32710 2742 32936
rect 21027 32917 21059 32997
rect 21139 32917 21184 32997
rect 21264 32917 21309 32997
rect 21389 32917 21427 32997
rect 21027 32888 21427 32917
rect 1866 32485 2742 32710
rect 463 32302 866 32360
rect 463 32226 503 32302
rect 575 32226 629 32302
rect 701 32226 749 32302
rect 821 32226 866 32302
rect 463 32184 866 32226
rect 463 32108 503 32184
rect 575 32108 629 32184
rect 701 32108 749 32184
rect 821 32108 866 32184
rect 463 32072 866 32108
rect 2306 31967 2742 32485
rect 21025 32302 21428 32360
rect 21025 32226 21068 32302
rect 21140 32226 21194 32302
rect 21266 32226 21314 32302
rect 21386 32226 21428 32302
rect 21025 32184 21428 32226
rect 21025 32108 21068 32184
rect 21140 32108 21194 32184
rect 21266 32108 21314 32184
rect 21386 32108 21428 32184
rect 21025 32072 21428 32108
rect 463 31520 863 31545
rect 463 31444 503 31520
rect 575 31444 629 31520
rect 701 31444 749 31520
rect 821 31444 863 31520
rect 463 31402 863 31444
rect 463 31326 503 31402
rect 575 31326 629 31402
rect 701 31326 749 31402
rect 821 31326 863 31402
rect 463 31290 863 31326
rect 21028 31520 21428 31545
rect 21028 31444 21068 31520
rect 21140 31444 21194 31520
rect 21266 31444 21314 31520
rect 21386 31444 21428 31520
rect 21028 31402 21428 31444
rect 21028 31326 21068 31402
rect 21140 31326 21194 31402
rect 21266 31326 21314 31402
rect 21386 31326 21428 31402
rect 21028 31290 21428 31326
rect 463 31061 863 31111
rect 463 30985 504 31061
rect 576 30985 626 31061
rect 698 30985 752 31061
rect 824 30985 863 31061
rect 463 30914 863 30985
rect 463 30838 504 30914
rect 576 30838 626 30914
rect 698 30838 752 30914
rect 824 30838 863 30914
rect 463 30777 863 30838
rect 463 30701 504 30777
rect 576 30701 626 30777
rect 698 30701 752 30777
rect 824 30701 863 30777
rect 463 30651 863 30701
rect 21970 30130 22370 30155
rect 21970 30054 22010 30130
rect 22082 30054 22136 30130
rect 22208 30054 22256 30130
rect 22328 30054 22370 30130
rect 21970 30012 22370 30054
rect 21970 29936 22010 30012
rect 22082 29936 22136 30012
rect 22208 29936 22256 30012
rect 22328 29936 22370 30012
rect 21970 29900 22370 29936
rect 463 29294 863 29349
rect 463 29218 504 29294
rect 576 29218 626 29294
rect 698 29218 752 29294
rect 824 29218 863 29294
rect 463 29147 863 29218
rect 463 29071 504 29147
rect 576 29071 626 29147
rect 698 29071 752 29147
rect 824 29071 863 29147
rect 463 29010 863 29071
rect 463 28934 504 29010
rect 576 28934 626 29010
rect 698 28934 752 29010
rect 824 28934 863 29010
rect 463 28890 863 28934
rect 463 28608 863 28633
rect 463 28532 503 28608
rect 575 28532 629 28608
rect 701 28532 749 28608
rect 821 28532 863 28608
rect 463 28490 863 28532
rect 463 28414 503 28490
rect 575 28414 629 28490
rect 701 28414 749 28490
rect 821 28414 863 28490
rect 463 28378 863 28414
rect 21028 28559 21428 28584
rect 21028 28483 21068 28559
rect 21140 28483 21194 28559
rect 21266 28483 21314 28559
rect 21386 28483 21428 28559
rect 21028 28441 21428 28483
rect 21028 28365 21068 28441
rect 21140 28365 21194 28441
rect 21266 28365 21314 28441
rect 21386 28365 21428 28441
rect 21028 28329 21428 28365
rect 463 27604 863 27629
rect 463 27528 503 27604
rect 575 27528 629 27604
rect 701 27528 749 27604
rect 821 27528 863 27604
rect 463 27486 863 27528
rect 463 27410 503 27486
rect 575 27410 629 27486
rect 701 27410 749 27486
rect 821 27410 863 27486
rect 463 27374 863 27410
rect 21027 27442 21427 27467
rect 21027 27366 21068 27442
rect 21140 27366 21194 27442
rect 21266 27366 21314 27442
rect 21386 27366 21427 27442
rect 21027 27324 21427 27366
rect 21027 27248 21068 27324
rect 21140 27248 21194 27324
rect 21266 27248 21314 27324
rect 21386 27248 21427 27324
rect 21027 27212 21427 27248
rect 463 27060 863 27109
rect 463 26984 504 27060
rect 576 26984 626 27060
rect 698 26984 752 27060
rect 824 26984 863 27060
rect 463 26913 863 26984
rect 463 26837 504 26913
rect 576 26837 626 26913
rect 698 26837 752 26913
rect 824 26837 863 26913
rect 463 26776 863 26837
rect 463 26700 504 26776
rect 576 26700 626 26776
rect 698 26700 752 26776
rect 824 26700 863 26776
rect 463 26650 863 26700
rect 21970 25971 22370 25996
rect 21970 25895 22010 25971
rect 22082 25895 22136 25971
rect 22208 25895 22256 25971
rect 22328 25895 22370 25971
rect 21970 25853 22370 25895
rect 21970 25777 22010 25853
rect 22082 25777 22136 25853
rect 22208 25777 22256 25853
rect 22328 25777 22370 25853
rect 21970 25741 22370 25777
rect 463 25300 863 25349
rect 463 25224 504 25300
rect 576 25224 626 25300
rect 698 25224 752 25300
rect 824 25224 863 25300
rect 463 25153 863 25224
rect 463 25077 504 25153
rect 576 25077 626 25153
rect 698 25077 752 25153
rect 824 25077 863 25153
rect 463 25016 863 25077
rect 463 24940 504 25016
rect 576 24940 626 25016
rect 698 24940 752 25016
rect 824 24940 863 25016
rect 463 24890 863 24940
rect 463 24626 864 24651
rect 463 24550 503 24626
rect 575 24550 629 24626
rect 701 24550 749 24626
rect 821 24550 864 24626
rect 463 24508 864 24550
rect 463 24432 503 24508
rect 575 24432 629 24508
rect 701 24432 749 24508
rect 821 24432 864 24508
rect 463 24396 864 24432
rect 21028 24599 21428 24624
rect 21028 24523 21068 24599
rect 21140 24523 21194 24599
rect 21266 24523 21314 24599
rect 21386 24523 21428 24599
rect 21028 24481 21428 24523
rect 21028 24405 21068 24481
rect 21140 24405 21194 24481
rect 21266 24405 21314 24481
rect 21386 24405 21428 24481
rect 21028 24369 21428 24405
rect 463 23544 864 23569
rect 463 23468 503 23544
rect 575 23468 629 23544
rect 701 23468 749 23544
rect 821 23468 864 23544
rect 463 23426 864 23468
rect 463 23350 503 23426
rect 575 23350 629 23426
rect 701 23350 749 23426
rect 821 23350 864 23426
rect 463 23314 864 23350
rect 21028 23424 21428 23449
rect 21028 23348 21068 23424
rect 21140 23348 21194 23424
rect 21266 23348 21314 23424
rect 21386 23348 21428 23424
rect 21028 23306 21428 23348
rect 21028 23230 21068 23306
rect 21140 23230 21194 23306
rect 21266 23230 21314 23306
rect 21386 23230 21428 23306
rect 21028 23194 21428 23230
rect 463 23060 863 23109
rect 463 22984 504 23060
rect 576 22984 626 23060
rect 698 22984 752 23060
rect 824 22984 863 23060
rect 463 22913 863 22984
rect 463 22837 504 22913
rect 576 22837 626 22913
rect 698 22837 752 22913
rect 824 22837 863 22913
rect 463 22776 863 22837
rect 463 22700 504 22776
rect 576 22700 626 22776
rect 698 22700 752 22776
rect 824 22700 863 22776
rect 463 22650 863 22700
rect 21970 22181 22370 22206
rect 21970 22105 22010 22181
rect 22082 22105 22136 22181
rect 22208 22105 22256 22181
rect 22328 22105 22370 22181
rect 21970 22063 22370 22105
rect 21970 21987 22010 22063
rect 22082 21987 22136 22063
rect 22208 21987 22256 22063
rect 22328 21987 22370 22063
rect 21970 21951 22370 21987
rect 463 21301 863 21350
rect 463 21225 504 21301
rect 576 21225 626 21301
rect 698 21225 752 21301
rect 824 21225 863 21301
rect 463 21154 863 21225
rect 463 21078 504 21154
rect 576 21078 626 21154
rect 698 21078 752 21154
rect 824 21078 863 21154
rect 463 21017 863 21078
rect 463 20941 504 21017
rect 576 20941 626 21017
rect 698 20941 752 21017
rect 824 20941 863 21017
rect 463 20891 863 20941
rect 463 20669 864 20694
rect 463 20593 503 20669
rect 575 20593 629 20669
rect 701 20593 749 20669
rect 821 20593 864 20669
rect 463 20551 864 20593
rect 463 20475 503 20551
rect 575 20475 629 20551
rect 701 20475 749 20551
rect 821 20475 864 20551
rect 463 20439 864 20475
rect 21027 20583 21427 20608
rect 21027 20507 21068 20583
rect 21140 20507 21194 20583
rect 21266 20507 21314 20583
rect 21386 20507 21427 20583
rect 21027 20465 21427 20507
rect 21027 20389 21068 20465
rect 21140 20389 21194 20465
rect 21266 20389 21314 20465
rect 21386 20389 21427 20465
rect 21027 20353 21427 20389
rect 463 19568 864 19593
rect 463 19492 503 19568
rect 575 19492 629 19568
rect 701 19492 749 19568
rect 821 19492 864 19568
rect 463 19450 864 19492
rect 463 19374 503 19450
rect 575 19374 629 19450
rect 701 19374 749 19450
rect 821 19374 864 19450
rect 463 19338 864 19374
rect 21027 19412 21427 19437
rect 21027 19336 21068 19412
rect 21140 19336 21194 19412
rect 21266 19336 21314 19412
rect 21386 19336 21427 19412
rect 21027 19294 21427 19336
rect 21027 19218 21068 19294
rect 21140 19218 21194 19294
rect 21266 19218 21314 19294
rect 21386 19218 21427 19294
rect 21027 19182 21427 19218
rect 463 19060 863 19109
rect 463 18984 504 19060
rect 576 18984 626 19060
rect 698 18984 752 19060
rect 824 18984 863 19060
rect 463 18913 863 18984
rect 463 18837 504 18913
rect 576 18837 626 18913
rect 698 18837 752 18913
rect 824 18837 863 18913
rect 463 18776 863 18837
rect 463 18700 504 18776
rect 576 18700 626 18776
rect 698 18700 752 18776
rect 824 18700 863 18776
rect 463 18650 863 18700
rect 21970 18074 22370 18099
rect 21970 17998 22010 18074
rect 22082 17998 22136 18074
rect 22208 17998 22256 18074
rect 22328 17998 22370 18074
rect 21970 17956 22370 17998
rect 21970 17880 22010 17956
rect 22082 17880 22136 17956
rect 22208 17880 22256 17956
rect 22328 17880 22370 17956
rect 21970 17844 22370 17880
rect 463 17300 863 17349
rect 463 17224 504 17300
rect 576 17224 626 17300
rect 698 17224 752 17300
rect 824 17224 863 17300
rect 463 17153 863 17224
rect 463 17077 504 17153
rect 576 17077 626 17153
rect 698 17077 752 17153
rect 824 17077 863 17153
rect 463 17016 863 17077
rect 463 16940 504 17016
rect 576 16940 626 17016
rect 698 16940 752 17016
rect 824 16940 863 17016
rect 463 16890 863 16940
rect 463 16702 865 16727
rect 463 16626 503 16702
rect 575 16626 629 16702
rect 701 16626 749 16702
rect 821 16626 865 16702
rect 463 16584 865 16626
rect 463 16508 503 16584
rect 575 16508 629 16584
rect 701 16508 749 16584
rect 821 16508 865 16584
rect 463 16472 865 16508
rect 21027 16651 21427 16676
rect 21027 16575 21068 16651
rect 21140 16575 21194 16651
rect 21266 16575 21314 16651
rect 21386 16575 21427 16651
rect 21027 16533 21427 16575
rect 21027 16457 21068 16533
rect 21140 16457 21194 16533
rect 21266 16457 21314 16533
rect 21386 16457 21427 16533
rect 21027 16421 21427 16457
rect 463 15486 866 15511
rect 463 15410 503 15486
rect 575 15410 629 15486
rect 701 15410 749 15486
rect 821 15410 866 15486
rect 463 15368 866 15410
rect 463 15292 503 15368
rect 575 15292 629 15368
rect 701 15292 749 15368
rect 821 15292 866 15368
rect 463 15256 866 15292
rect 21027 15437 21427 15462
rect 21027 15361 21068 15437
rect 21140 15361 21194 15437
rect 21266 15361 21314 15437
rect 21386 15361 21427 15437
rect 21027 15319 21427 15361
rect 21027 15243 21068 15319
rect 21140 15243 21194 15319
rect 21266 15243 21314 15319
rect 21386 15243 21427 15319
rect 21027 15207 21427 15243
rect 463 15060 863 15109
rect 463 14984 504 15060
rect 576 14984 626 15060
rect 698 14984 752 15060
rect 824 14984 863 15060
rect 463 14913 863 14984
rect 463 14837 504 14913
rect 576 14837 626 14913
rect 698 14837 752 14913
rect 824 14837 863 14913
rect 463 14776 863 14837
rect 463 14700 504 14776
rect 576 14700 626 14776
rect 698 14700 752 14776
rect 824 14700 863 14776
rect 463 14650 863 14700
rect 21970 14256 22370 14281
rect 21970 14180 22010 14256
rect 22082 14180 22136 14256
rect 22208 14180 22256 14256
rect 22328 14180 22370 14256
rect 21970 14138 22370 14180
rect 21970 14062 22010 14138
rect 22082 14062 22136 14138
rect 22208 14062 22256 14138
rect 22328 14062 22370 14138
rect 21970 14026 22370 14062
rect 463 13300 863 13349
rect 463 13224 504 13300
rect 576 13224 626 13300
rect 698 13224 752 13300
rect 824 13224 863 13300
rect 463 13153 863 13224
rect 463 13077 504 13153
rect 576 13077 626 13153
rect 698 13077 752 13153
rect 824 13077 863 13153
rect 463 13016 863 13077
rect 463 12940 504 13016
rect 576 12940 626 13016
rect 698 12940 752 13016
rect 824 12940 863 13016
rect 463 12890 863 12940
rect 463 12621 864 12646
rect 463 12545 503 12621
rect 575 12545 629 12621
rect 701 12545 749 12621
rect 821 12545 864 12621
rect 463 12503 864 12545
rect 463 12427 503 12503
rect 575 12427 629 12503
rect 701 12427 749 12503
rect 821 12427 864 12503
rect 463 12391 864 12427
rect 21028 12594 21428 12619
rect 21028 12518 21068 12594
rect 21140 12518 21194 12594
rect 21266 12518 21314 12594
rect 21386 12518 21428 12594
rect 21028 12476 21428 12518
rect 21028 12400 21068 12476
rect 21140 12400 21194 12476
rect 21266 12400 21314 12476
rect 21386 12400 21428 12476
rect 21028 12364 21428 12400
rect 463 11499 864 11524
rect 463 11423 503 11499
rect 575 11423 629 11499
rect 701 11423 749 11499
rect 821 11423 864 11499
rect 463 11381 864 11423
rect 463 11305 503 11381
rect 575 11305 629 11381
rect 701 11305 749 11381
rect 821 11305 864 11381
rect 463 11269 864 11305
rect 21027 11437 21427 11462
rect 21027 11361 21068 11437
rect 21140 11361 21194 11437
rect 21266 11361 21314 11437
rect 21386 11361 21427 11437
rect 21027 11319 21427 11361
rect 21027 11243 21068 11319
rect 21140 11243 21194 11319
rect 21266 11243 21314 11319
rect 21386 11243 21427 11319
rect 21027 11207 21427 11243
rect 463 11061 863 11110
rect 463 10985 504 11061
rect 576 10985 626 11061
rect 698 10985 752 11061
rect 824 10985 863 11061
rect 463 10914 863 10985
rect 463 10838 504 10914
rect 576 10838 626 10914
rect 698 10838 752 10914
rect 824 10838 863 10914
rect 463 10777 863 10838
rect 463 10701 504 10777
rect 576 10701 626 10777
rect 698 10701 752 10777
rect 824 10701 863 10777
rect 463 10651 863 10701
rect 21970 10292 22370 10317
rect 21970 10216 22010 10292
rect 22082 10216 22136 10292
rect 22208 10216 22256 10292
rect 22328 10216 22370 10292
rect 21970 10174 22370 10216
rect 21970 10098 22010 10174
rect 22082 10098 22136 10174
rect 22208 10098 22256 10174
rect 22328 10098 22370 10174
rect 21970 10062 22370 10098
rect 463 9299 863 9348
rect 463 9223 504 9299
rect 576 9223 626 9299
rect 698 9223 752 9299
rect 824 9223 863 9299
rect 463 9152 863 9223
rect 463 9076 504 9152
rect 576 9076 626 9152
rect 698 9076 752 9152
rect 824 9076 863 9152
rect 463 9015 863 9076
rect 463 8939 504 9015
rect 576 8939 626 9015
rect 698 8939 752 9015
rect 824 8939 863 9015
rect 463 8889 863 8939
rect 463 8639 863 8664
rect 463 8563 503 8639
rect 575 8563 629 8639
rect 701 8563 749 8639
rect 821 8563 863 8639
rect 463 8521 863 8563
rect 463 8445 503 8521
rect 575 8445 629 8521
rect 701 8445 749 8521
rect 821 8445 863 8521
rect 463 8409 863 8445
rect 21028 8594 21428 8619
rect 21028 8518 21068 8594
rect 21140 8518 21194 8594
rect 21266 8518 21314 8594
rect 21386 8518 21428 8594
rect 21028 8476 21428 8518
rect 21028 8400 21068 8476
rect 21140 8400 21194 8476
rect 21266 8400 21314 8476
rect 21386 8400 21428 8476
rect 21028 8364 21428 8400
rect 463 7528 863 7553
rect 463 7452 503 7528
rect 575 7452 629 7528
rect 701 7452 749 7528
rect 821 7452 863 7528
rect 463 7410 863 7452
rect 463 7334 503 7410
rect 575 7334 629 7410
rect 701 7334 749 7410
rect 821 7334 863 7410
rect 463 7298 863 7334
rect 21027 7437 21427 7462
rect 21027 7361 21068 7437
rect 21140 7361 21194 7437
rect 21266 7361 21314 7437
rect 21386 7361 21427 7437
rect 21027 7319 21427 7361
rect 21027 7243 21068 7319
rect 21140 7243 21194 7319
rect 21266 7243 21314 7319
rect 21386 7243 21427 7319
rect 21027 7207 21427 7243
rect 463 7061 863 7110
rect 463 6985 504 7061
rect 576 6985 626 7061
rect 698 6985 752 7061
rect 824 6985 863 7061
rect 463 6914 863 6985
rect 463 6838 504 6914
rect 576 6838 626 6914
rect 698 6838 752 6914
rect 824 6838 863 6914
rect 463 6777 863 6838
rect 463 6701 504 6777
rect 576 6701 626 6777
rect 698 6701 752 6777
rect 824 6701 863 6777
rect 463 6651 863 6701
rect 21970 6280 22370 6305
rect 21970 6204 22010 6280
rect 22082 6204 22136 6280
rect 22208 6204 22256 6280
rect 22328 6204 22370 6280
rect 21970 6162 22370 6204
rect 21970 6086 22010 6162
rect 22082 6086 22136 6162
rect 22208 6086 22256 6162
rect 22328 6086 22370 6162
rect 21970 6050 22370 6086
rect 463 5300 863 5349
rect 463 5224 504 5300
rect 576 5224 626 5300
rect 698 5224 752 5300
rect 824 5224 863 5300
rect 463 5153 863 5224
rect 463 5077 504 5153
rect 576 5077 626 5153
rect 698 5077 752 5153
rect 824 5077 863 5153
rect 463 5016 863 5077
rect 463 4940 504 5016
rect 576 4940 626 5016
rect 698 4940 752 5016
rect 824 4940 863 5016
rect 463 4890 863 4940
rect 463 4705 865 4730
rect 463 4629 503 4705
rect 575 4629 629 4705
rect 701 4629 749 4705
rect 821 4629 865 4705
rect 463 4587 865 4629
rect 463 4511 503 4587
rect 575 4511 629 4587
rect 701 4511 749 4587
rect 821 4511 865 4587
rect 463 4475 865 4511
rect 21028 4594 21428 4619
rect 21028 4518 21068 4594
rect 21140 4518 21194 4594
rect 21266 4518 21314 4594
rect 21386 4518 21428 4594
rect 21028 4476 21428 4518
rect 21028 4400 21068 4476
rect 21140 4400 21194 4476
rect 21266 4400 21314 4476
rect 21386 4400 21428 4476
rect 21028 4364 21428 4400
rect 463 3528 863 3553
rect 463 3452 503 3528
rect 575 3452 629 3528
rect 701 3452 749 3528
rect 821 3452 863 3528
rect 463 3410 863 3452
rect 463 3334 503 3410
rect 575 3334 629 3410
rect 701 3334 749 3410
rect 821 3334 863 3410
rect 463 3298 863 3334
rect 21027 3437 21427 3462
rect 21027 3361 21068 3437
rect 21140 3361 21194 3437
rect 21266 3361 21314 3437
rect 21386 3361 21427 3437
rect 21027 3319 21427 3361
rect 21027 3243 21068 3319
rect 21140 3243 21194 3319
rect 21266 3243 21314 3319
rect 21386 3243 21427 3319
rect 21027 3207 21427 3243
rect 463 3061 863 3110
rect 463 2985 504 3061
rect 576 2985 626 3061
rect 698 2985 752 3061
rect 824 2985 863 3061
rect 463 2914 863 2985
rect 463 2838 504 2914
rect 576 2838 626 2914
rect 698 2838 752 2914
rect 824 2838 863 2914
rect 463 2777 863 2838
rect 463 2701 504 2777
rect 576 2701 626 2777
rect 698 2701 752 2777
rect 824 2701 863 2777
rect 463 2651 863 2701
rect 21970 2280 22370 2305
rect 21970 2204 22010 2280
rect 22082 2204 22136 2280
rect 22208 2204 22256 2280
rect 22328 2204 22370 2280
rect 21970 2162 22370 2204
rect 21970 2086 22010 2162
rect 22082 2086 22136 2162
rect 22208 2086 22256 2162
rect 22328 2086 22370 2162
rect 21970 2050 22370 2086
rect 463 1300 863 1349
rect 463 1224 504 1300
rect 576 1224 626 1300
rect 698 1224 752 1300
rect 824 1224 863 1300
rect 463 1153 863 1224
rect 463 1077 504 1153
rect 576 1077 626 1153
rect 698 1077 752 1153
rect 824 1077 863 1153
rect 463 1016 863 1077
rect 463 940 504 1016
rect 576 940 626 1016
rect 698 940 752 1016
rect 824 940 863 1016
rect 463 890 863 940
rect 463 705 865 730
rect 463 629 503 705
rect 575 629 629 705
rect 701 629 749 705
rect 821 629 865 705
rect 463 587 865 629
rect 463 511 503 587
rect 575 511 629 587
rect 701 511 749 587
rect 821 511 865 587
rect 463 475 865 511
rect 21028 594 21428 619
rect 21028 518 21068 594
rect 21140 518 21194 594
rect 21266 518 21314 594
rect 21386 518 21428 594
rect 21028 476 21428 518
rect 21028 400 21068 476
rect 21140 400 21194 476
rect 21266 400 21314 476
rect 21386 400 21428 476
rect 21028 364 21428 400
<< via2 >>
rect 503 75376 575 75452
rect 629 75376 701 75452
rect 749 75376 821 75452
rect 503 75258 575 75334
rect 629 75258 701 75334
rect 749 75258 821 75334
rect 21068 75416 21140 75492
rect 21194 75416 21266 75492
rect 21314 75416 21386 75492
rect 21068 75298 21140 75374
rect 21194 75298 21266 75374
rect 21314 75298 21386 75374
rect 504 74984 576 75060
rect 626 74984 698 75060
rect 752 74984 824 75060
rect 504 74837 576 74913
rect 626 74837 698 74913
rect 752 74837 824 74913
rect 504 74700 576 74776
rect 626 74700 698 74776
rect 752 74700 824 74776
rect 22010 73995 22082 74071
rect 22136 73995 22208 74071
rect 22256 73995 22328 74071
rect 22010 73877 22082 73953
rect 22136 73877 22208 73953
rect 22256 73877 22328 73953
rect 504 73224 576 73300
rect 626 73224 698 73300
rect 752 73224 824 73300
rect 504 73077 576 73153
rect 626 73077 698 73153
rect 752 73077 824 73153
rect 504 72940 576 73016
rect 626 72940 698 73016
rect 752 72940 824 73016
rect 503 72703 575 72779
rect 629 72703 701 72779
rect 749 72703 821 72779
rect 503 72585 575 72661
rect 629 72585 701 72661
rect 749 72585 821 72661
rect 21068 72619 21140 72695
rect 21194 72619 21266 72695
rect 21314 72619 21386 72695
rect 21068 72501 21140 72577
rect 21194 72501 21266 72577
rect 21314 72501 21386 72577
rect 503 71376 575 71452
rect 629 71376 701 71452
rect 749 71376 821 71452
rect 503 71258 575 71334
rect 629 71258 701 71334
rect 749 71258 821 71334
rect 21068 71416 21140 71492
rect 21194 71416 21266 71492
rect 21314 71416 21386 71492
rect 21068 71298 21140 71374
rect 21194 71298 21266 71374
rect 21314 71298 21386 71374
rect 504 70984 576 71060
rect 626 70984 698 71060
rect 752 70984 824 71060
rect 504 70837 576 70913
rect 626 70837 698 70913
rect 752 70837 824 70913
rect 504 70700 576 70776
rect 626 70700 698 70776
rect 752 70700 824 70776
rect 22010 69995 22082 70071
rect 22136 69995 22208 70071
rect 22256 69995 22328 70071
rect 22010 69877 22082 69953
rect 22136 69877 22208 69953
rect 22256 69877 22328 69953
rect 504 69224 576 69300
rect 626 69224 698 69300
rect 752 69224 824 69300
rect 504 69077 576 69153
rect 626 69077 698 69153
rect 752 69077 824 69153
rect 504 68940 576 69016
rect 626 68940 698 69016
rect 752 68940 824 69016
rect 503 68703 575 68779
rect 629 68703 701 68779
rect 749 68703 821 68779
rect 503 68585 575 68661
rect 629 68585 701 68661
rect 749 68585 821 68661
rect 21068 68619 21140 68695
rect 21194 68619 21266 68695
rect 21314 68619 21386 68695
rect 21068 68501 21140 68577
rect 21194 68501 21266 68577
rect 21314 68501 21386 68577
rect 503 67374 575 67450
rect 629 67374 701 67450
rect 749 67374 821 67450
rect 503 67256 575 67332
rect 629 67256 701 67332
rect 749 67256 821 67332
rect 21068 67416 21140 67492
rect 21194 67416 21266 67492
rect 21314 67416 21386 67492
rect 21068 67298 21140 67374
rect 21194 67298 21266 67374
rect 21314 67298 21386 67374
rect 504 66984 576 67060
rect 626 66984 698 67060
rect 752 66984 824 67060
rect 504 66837 576 66913
rect 626 66837 698 66913
rect 752 66837 824 66913
rect 504 66700 576 66776
rect 626 66700 698 66776
rect 752 66700 824 66776
rect 22010 65982 22082 66058
rect 22136 65982 22208 66058
rect 22256 65982 22328 66058
rect 22010 65864 22082 65940
rect 22136 65864 22208 65940
rect 22256 65864 22328 65940
rect 504 65225 576 65301
rect 626 65225 698 65301
rect 752 65225 824 65301
rect 504 65078 576 65154
rect 626 65078 698 65154
rect 752 65078 824 65154
rect 504 64941 576 65017
rect 626 64941 698 65017
rect 752 64941 824 65017
rect 503 64634 575 64710
rect 629 64634 701 64710
rect 749 64634 821 64710
rect 503 64516 575 64592
rect 629 64516 701 64592
rect 749 64516 821 64592
rect 21068 64619 21140 64695
rect 21194 64619 21266 64695
rect 21314 64619 21386 64695
rect 21068 64501 21140 64577
rect 21194 64501 21266 64577
rect 21314 64501 21386 64577
rect 503 63456 575 63532
rect 629 63456 701 63532
rect 749 63456 821 63532
rect 503 63338 575 63414
rect 629 63338 701 63414
rect 749 63338 821 63414
rect 21068 63416 21140 63492
rect 21194 63416 21266 63492
rect 21314 63416 21386 63492
rect 21068 63298 21140 63374
rect 21194 63298 21266 63374
rect 21314 63298 21386 63374
rect 504 62984 576 63060
rect 626 62984 698 63060
rect 752 62984 824 63060
rect 504 62837 576 62913
rect 626 62837 698 62913
rect 752 62837 824 62913
rect 504 62700 576 62776
rect 626 62700 698 62776
rect 752 62700 824 62776
rect 22010 61981 22082 62057
rect 22136 61981 22208 62057
rect 22256 61981 22328 62057
rect 22010 61863 22082 61939
rect 22136 61863 22208 61939
rect 22256 61863 22328 61939
rect 504 61225 576 61301
rect 626 61225 698 61301
rect 752 61225 824 61301
rect 504 61078 576 61154
rect 626 61078 698 61154
rect 752 61078 824 61154
rect 504 60941 576 61017
rect 626 60941 698 61017
rect 752 60941 824 61017
rect 503 60608 575 60684
rect 629 60608 701 60684
rect 749 60608 821 60684
rect 503 60490 575 60566
rect 629 60490 701 60566
rect 749 60490 821 60566
rect 21068 60619 21140 60695
rect 21194 60619 21266 60695
rect 21314 60619 21386 60695
rect 21068 60501 21140 60577
rect 21194 60501 21266 60577
rect 21314 60501 21386 60577
rect 503 59405 575 59481
rect 629 59405 701 59481
rect 749 59405 821 59481
rect 503 59287 575 59363
rect 629 59287 701 59363
rect 749 59287 821 59363
rect 21068 59470 21140 59546
rect 21194 59470 21266 59546
rect 21314 59470 21386 59546
rect 21068 59352 21140 59428
rect 21194 59352 21266 59428
rect 21314 59352 21386 59428
rect 504 58984 576 59060
rect 626 58984 698 59060
rect 752 58984 824 59060
rect 504 58837 576 58913
rect 626 58837 698 58913
rect 752 58837 824 58913
rect 504 58700 576 58776
rect 626 58700 698 58776
rect 752 58700 824 58776
rect 22010 58020 22082 58096
rect 22136 58020 22208 58096
rect 22256 58020 22328 58096
rect 22010 57902 22082 57978
rect 22136 57902 22208 57978
rect 22256 57902 22328 57978
rect 504 57223 576 57299
rect 626 57223 698 57299
rect 752 57223 824 57299
rect 504 57076 576 57152
rect 626 57076 698 57152
rect 752 57076 824 57152
rect 504 56939 576 57015
rect 626 56939 698 57015
rect 752 56939 824 57015
rect 503 56628 575 56704
rect 629 56628 701 56704
rect 749 56628 821 56704
rect 503 56510 575 56586
rect 629 56510 701 56586
rect 749 56510 821 56586
rect 21068 56554 21140 56630
rect 21194 56554 21266 56630
rect 21314 56554 21386 56630
rect 21068 56436 21140 56512
rect 21194 56436 21266 56512
rect 21314 56436 21386 56512
rect 503 55421 575 55497
rect 629 55421 701 55497
rect 749 55421 821 55497
rect 503 55303 575 55379
rect 629 55303 701 55379
rect 749 55303 821 55379
rect 21068 55371 21140 55447
rect 21194 55371 21266 55447
rect 21314 55371 21386 55447
rect 21068 55253 21140 55329
rect 21194 55253 21266 55329
rect 21314 55253 21386 55329
rect 504 54984 576 55060
rect 626 54984 698 55060
rect 752 54984 824 55060
rect 504 54837 576 54913
rect 626 54837 698 54913
rect 752 54837 824 54913
rect 504 54700 576 54776
rect 626 54700 698 54776
rect 752 54700 824 54776
rect 22010 54003 22082 54079
rect 22136 54003 22208 54079
rect 22256 54003 22328 54079
rect 22010 53885 22082 53961
rect 22136 53885 22208 53961
rect 22256 53885 22328 53961
rect 504 53225 576 53301
rect 626 53225 698 53301
rect 752 53225 824 53301
rect 504 53078 576 53154
rect 626 53078 698 53154
rect 752 53078 824 53154
rect 504 52941 576 53017
rect 626 52941 698 53017
rect 752 52941 824 53017
rect 503 52655 575 52731
rect 629 52655 701 52731
rect 749 52655 821 52731
rect 503 52537 575 52613
rect 629 52537 701 52613
rect 749 52537 821 52613
rect 21068 52499 21140 52575
rect 21194 52499 21266 52575
rect 21314 52499 21386 52575
rect 21068 52381 21140 52457
rect 21194 52381 21266 52457
rect 21314 52381 21386 52457
rect 503 51468 575 51544
rect 629 51468 701 51544
rect 749 51468 821 51544
rect 503 51350 575 51426
rect 629 51350 701 51426
rect 749 51350 821 51426
rect 21068 51364 21140 51440
rect 21194 51364 21266 51440
rect 21314 51364 21386 51440
rect 21068 51246 21140 51322
rect 21194 51246 21266 51322
rect 21314 51246 21386 51322
rect 504 50984 576 51060
rect 626 50984 698 51060
rect 752 50984 824 51060
rect 504 50837 576 50913
rect 626 50837 698 50913
rect 752 50837 824 50913
rect 504 50700 576 50776
rect 626 50700 698 50776
rect 752 50700 824 50776
rect 22010 50082 22082 50158
rect 22136 50082 22208 50158
rect 22256 50082 22328 50158
rect 22010 49964 22082 50040
rect 22136 49964 22208 50040
rect 22256 49964 22328 50040
rect 504 49225 576 49301
rect 626 49225 698 49301
rect 752 49225 824 49301
rect 504 49078 576 49154
rect 626 49078 698 49154
rect 752 49078 824 49154
rect 504 48941 576 49017
rect 626 48941 698 49017
rect 752 48941 824 49017
rect 503 48646 575 48722
rect 629 48646 701 48722
rect 749 48646 821 48722
rect 503 48528 575 48604
rect 629 48528 701 48604
rect 749 48528 821 48604
rect 21068 48605 21140 48681
rect 21194 48605 21266 48681
rect 21314 48605 21386 48681
rect 21068 48487 21140 48563
rect 21194 48487 21266 48563
rect 21314 48487 21386 48563
rect 503 47493 575 47569
rect 629 47493 701 47569
rect 749 47493 821 47569
rect 503 47375 575 47451
rect 629 47375 701 47451
rect 749 47375 821 47451
rect 21068 47452 21140 47528
rect 21194 47452 21266 47528
rect 21314 47452 21386 47528
rect 21068 47334 21140 47410
rect 21194 47334 21266 47410
rect 21314 47334 21386 47410
rect 504 46984 576 47060
rect 626 46984 698 47060
rect 752 46984 824 47060
rect 504 46837 576 46913
rect 626 46837 698 46913
rect 752 46837 824 46913
rect 504 46700 576 46776
rect 626 46700 698 46776
rect 752 46700 824 46776
rect 22010 45824 22082 45900
rect 22136 45824 22208 45900
rect 22256 45824 22328 45900
rect 22010 45706 22082 45782
rect 22136 45706 22208 45782
rect 22256 45706 22328 45782
rect 504 45224 576 45300
rect 626 45224 698 45300
rect 752 45224 824 45300
rect 504 45077 576 45153
rect 626 45077 698 45153
rect 752 45077 824 45153
rect 504 44940 576 45016
rect 626 44940 698 45016
rect 752 44940 824 45016
rect 503 44433 575 44509
rect 629 44433 701 44509
rect 749 44433 821 44509
rect 503 44315 575 44391
rect 629 44315 701 44391
rect 749 44315 821 44391
rect 21068 44336 21140 44412
rect 21194 44336 21266 44412
rect 21314 44336 21386 44412
rect 21068 44218 21140 44294
rect 21194 44218 21266 44294
rect 21314 44218 21386 44294
rect 2257 39869 2313 39925
rect 2337 39869 2393 39925
rect 2257 39789 2313 39845
rect 2337 39789 2393 39845
rect 32 39661 112 39741
rect 157 39661 237 39741
rect 282 39661 362 39741
rect 32 39555 112 39635
rect 157 39555 237 39635
rect 282 39555 362 39635
rect 1416 39263 1472 39319
rect 1498 39264 1554 39320
rect 1417 39183 1473 39239
rect 1499 39184 1555 39240
rect 22006 43514 22298 43838
rect 3361 39848 3417 39904
rect 3441 39848 3497 39904
rect 3361 39768 3417 39824
rect 3441 39768 3497 39824
rect 479 39052 561 39130
rect 593 39052 675 39130
rect 707 39052 789 39130
rect 16 38508 98 38586
rect 130 38508 212 38586
rect 244 38508 326 38586
rect 479 37964 561 38042
rect 593 37964 675 38042
rect 707 37964 789 38042
rect 16 37420 98 37498
rect 130 37420 212 37498
rect 244 37420 326 37498
rect 479 36876 561 36954
rect 593 36876 675 36954
rect 707 36876 789 36954
rect 2760 39262 2816 39318
rect 2840 39261 2896 39317
rect 2761 39181 2817 39237
rect 2841 39181 2897 39237
rect 21535 39646 21615 39726
rect 21660 39646 21740 39726
rect 21785 39646 21865 39726
rect 21534 39526 21614 39606
rect 21659 39526 21739 39606
rect 21784 39526 21864 39606
rect 3360 39261 3416 39317
rect 3440 39260 3496 39316
rect 3361 39180 3417 39236
rect 3441 39180 3497 39236
rect 22006 36630 22298 36954
rect 2544 36401 2600 36463
rect 2624 36401 2680 36463
rect 21061 36092 21141 36172
rect 21186 36092 21266 36172
rect 21311 36092 21391 36172
rect 21060 35972 21140 36052
rect 21185 35972 21265 36052
rect 21310 35972 21390 36052
rect 21069 35516 21141 35592
rect 21191 35516 21263 35592
rect 21317 35516 21389 35592
rect 21069 35369 21141 35445
rect 21191 35369 21263 35445
rect 21317 35369 21389 35445
rect 21069 35232 21141 35308
rect 21191 35232 21263 35308
rect 21317 35232 21389 35308
rect 20560 34596 20640 34676
rect 20685 34596 20765 34676
rect 20810 34596 20890 34676
rect 20559 34476 20639 34556
rect 20684 34476 20764 34556
rect 20809 34476 20889 34556
rect 21535 34596 21615 34676
rect 21660 34596 21740 34676
rect 21785 34596 21865 34676
rect 21534 34476 21614 34556
rect 21659 34476 21739 34556
rect 21784 34476 21864 34556
rect 21069 33756 21141 33832
rect 21191 33756 21263 33832
rect 21317 33756 21389 33832
rect 21069 33609 21141 33685
rect 21191 33609 21263 33685
rect 21317 33609 21389 33685
rect 21069 33472 21141 33548
rect 21191 33472 21263 33548
rect 21317 33472 21389 33548
rect 21060 33037 21140 33117
rect 21185 33037 21265 33117
rect 21310 33037 21390 33117
rect 21059 32917 21139 32997
rect 21184 32917 21264 32997
rect 21309 32917 21389 32997
rect 503 32226 575 32302
rect 629 32226 701 32302
rect 749 32226 821 32302
rect 503 32108 575 32184
rect 629 32108 701 32184
rect 749 32108 821 32184
rect 21068 32226 21140 32302
rect 21194 32226 21266 32302
rect 21314 32226 21386 32302
rect 21068 32108 21140 32184
rect 21194 32108 21266 32184
rect 21314 32108 21386 32184
rect 503 31444 575 31520
rect 629 31444 701 31520
rect 749 31444 821 31520
rect 503 31326 575 31402
rect 629 31326 701 31402
rect 749 31326 821 31402
rect 21068 31444 21140 31520
rect 21194 31444 21266 31520
rect 21314 31444 21386 31520
rect 21068 31326 21140 31402
rect 21194 31326 21266 31402
rect 21314 31326 21386 31402
rect 504 30985 576 31061
rect 626 30985 698 31061
rect 752 30985 824 31061
rect 504 30838 576 30914
rect 626 30838 698 30914
rect 752 30838 824 30914
rect 504 30701 576 30777
rect 626 30701 698 30777
rect 752 30701 824 30777
rect 22010 30054 22082 30130
rect 22136 30054 22208 30130
rect 22256 30054 22328 30130
rect 22010 29936 22082 30012
rect 22136 29936 22208 30012
rect 22256 29936 22328 30012
rect 504 29218 576 29294
rect 626 29218 698 29294
rect 752 29218 824 29294
rect 504 29071 576 29147
rect 626 29071 698 29147
rect 752 29071 824 29147
rect 504 28934 576 29010
rect 626 28934 698 29010
rect 752 28934 824 29010
rect 503 28532 575 28608
rect 629 28532 701 28608
rect 749 28532 821 28608
rect 503 28414 575 28490
rect 629 28414 701 28490
rect 749 28414 821 28490
rect 21068 28483 21140 28559
rect 21194 28483 21266 28559
rect 21314 28483 21386 28559
rect 21068 28365 21140 28441
rect 21194 28365 21266 28441
rect 21314 28365 21386 28441
rect 503 27528 575 27604
rect 629 27528 701 27604
rect 749 27528 821 27604
rect 503 27410 575 27486
rect 629 27410 701 27486
rect 749 27410 821 27486
rect 21068 27366 21140 27442
rect 21194 27366 21266 27442
rect 21314 27366 21386 27442
rect 21068 27248 21140 27324
rect 21194 27248 21266 27324
rect 21314 27248 21386 27324
rect 504 26984 576 27060
rect 626 26984 698 27060
rect 752 26984 824 27060
rect 504 26837 576 26913
rect 626 26837 698 26913
rect 752 26837 824 26913
rect 504 26700 576 26776
rect 626 26700 698 26776
rect 752 26700 824 26776
rect 22010 25895 22082 25971
rect 22136 25895 22208 25971
rect 22256 25895 22328 25971
rect 22010 25777 22082 25853
rect 22136 25777 22208 25853
rect 22256 25777 22328 25853
rect 504 25224 576 25300
rect 626 25224 698 25300
rect 752 25224 824 25300
rect 504 25077 576 25153
rect 626 25077 698 25153
rect 752 25077 824 25153
rect 504 24940 576 25016
rect 626 24940 698 25016
rect 752 24940 824 25016
rect 503 24550 575 24626
rect 629 24550 701 24626
rect 749 24550 821 24626
rect 503 24432 575 24508
rect 629 24432 701 24508
rect 749 24432 821 24508
rect 21068 24523 21140 24599
rect 21194 24523 21266 24599
rect 21314 24523 21386 24599
rect 21068 24405 21140 24481
rect 21194 24405 21266 24481
rect 21314 24405 21386 24481
rect 503 23468 575 23544
rect 629 23468 701 23544
rect 749 23468 821 23544
rect 503 23350 575 23426
rect 629 23350 701 23426
rect 749 23350 821 23426
rect 21068 23348 21140 23424
rect 21194 23348 21266 23424
rect 21314 23348 21386 23424
rect 21068 23230 21140 23306
rect 21194 23230 21266 23306
rect 21314 23230 21386 23306
rect 504 22984 576 23060
rect 626 22984 698 23060
rect 752 22984 824 23060
rect 504 22837 576 22913
rect 626 22837 698 22913
rect 752 22837 824 22913
rect 504 22700 576 22776
rect 626 22700 698 22776
rect 752 22700 824 22776
rect 22010 22105 22082 22181
rect 22136 22105 22208 22181
rect 22256 22105 22328 22181
rect 22010 21987 22082 22063
rect 22136 21987 22208 22063
rect 22256 21987 22328 22063
rect 504 21225 576 21301
rect 626 21225 698 21301
rect 752 21225 824 21301
rect 504 21078 576 21154
rect 626 21078 698 21154
rect 752 21078 824 21154
rect 504 20941 576 21017
rect 626 20941 698 21017
rect 752 20941 824 21017
rect 503 20593 575 20669
rect 629 20593 701 20669
rect 749 20593 821 20669
rect 503 20475 575 20551
rect 629 20475 701 20551
rect 749 20475 821 20551
rect 21068 20507 21140 20583
rect 21194 20507 21266 20583
rect 21314 20507 21386 20583
rect 21068 20389 21140 20465
rect 21194 20389 21266 20465
rect 21314 20389 21386 20465
rect 503 19492 575 19568
rect 629 19492 701 19568
rect 749 19492 821 19568
rect 503 19374 575 19450
rect 629 19374 701 19450
rect 749 19374 821 19450
rect 21068 19336 21140 19412
rect 21194 19336 21266 19412
rect 21314 19336 21386 19412
rect 21068 19218 21140 19294
rect 21194 19218 21266 19294
rect 21314 19218 21386 19294
rect 504 18984 576 19060
rect 626 18984 698 19060
rect 752 18984 824 19060
rect 504 18837 576 18913
rect 626 18837 698 18913
rect 752 18837 824 18913
rect 504 18700 576 18776
rect 626 18700 698 18776
rect 752 18700 824 18776
rect 22010 17998 22082 18074
rect 22136 17998 22208 18074
rect 22256 17998 22328 18074
rect 22010 17880 22082 17956
rect 22136 17880 22208 17956
rect 22256 17880 22328 17956
rect 504 17224 576 17300
rect 626 17224 698 17300
rect 752 17224 824 17300
rect 504 17077 576 17153
rect 626 17077 698 17153
rect 752 17077 824 17153
rect 504 16940 576 17016
rect 626 16940 698 17016
rect 752 16940 824 17016
rect 503 16626 575 16702
rect 629 16626 701 16702
rect 749 16626 821 16702
rect 503 16508 575 16584
rect 629 16508 701 16584
rect 749 16508 821 16584
rect 21068 16575 21140 16651
rect 21194 16575 21266 16651
rect 21314 16575 21386 16651
rect 21068 16457 21140 16533
rect 21194 16457 21266 16533
rect 21314 16457 21386 16533
rect 503 15410 575 15486
rect 629 15410 701 15486
rect 749 15410 821 15486
rect 503 15292 575 15368
rect 629 15292 701 15368
rect 749 15292 821 15368
rect 21068 15361 21140 15437
rect 21194 15361 21266 15437
rect 21314 15361 21386 15437
rect 21068 15243 21140 15319
rect 21194 15243 21266 15319
rect 21314 15243 21386 15319
rect 504 14984 576 15060
rect 626 14984 698 15060
rect 752 14984 824 15060
rect 504 14837 576 14913
rect 626 14837 698 14913
rect 752 14837 824 14913
rect 504 14700 576 14776
rect 626 14700 698 14776
rect 752 14700 824 14776
rect 22010 14180 22082 14256
rect 22136 14180 22208 14256
rect 22256 14180 22328 14256
rect 22010 14062 22082 14138
rect 22136 14062 22208 14138
rect 22256 14062 22328 14138
rect 504 13224 576 13300
rect 626 13224 698 13300
rect 752 13224 824 13300
rect 504 13077 576 13153
rect 626 13077 698 13153
rect 752 13077 824 13153
rect 504 12940 576 13016
rect 626 12940 698 13016
rect 752 12940 824 13016
rect 503 12545 575 12621
rect 629 12545 701 12621
rect 749 12545 821 12621
rect 503 12427 575 12503
rect 629 12427 701 12503
rect 749 12427 821 12503
rect 21068 12518 21140 12594
rect 21194 12518 21266 12594
rect 21314 12518 21386 12594
rect 21068 12400 21140 12476
rect 21194 12400 21266 12476
rect 21314 12400 21386 12476
rect 503 11423 575 11499
rect 629 11423 701 11499
rect 749 11423 821 11499
rect 503 11305 575 11381
rect 629 11305 701 11381
rect 749 11305 821 11381
rect 21068 11361 21140 11437
rect 21194 11361 21266 11437
rect 21314 11361 21386 11437
rect 21068 11243 21140 11319
rect 21194 11243 21266 11319
rect 21314 11243 21386 11319
rect 504 10985 576 11061
rect 626 10985 698 11061
rect 752 10985 824 11061
rect 504 10838 576 10914
rect 626 10838 698 10914
rect 752 10838 824 10914
rect 504 10701 576 10777
rect 626 10701 698 10777
rect 752 10701 824 10777
rect 22010 10216 22082 10292
rect 22136 10216 22208 10292
rect 22256 10216 22328 10292
rect 22010 10098 22082 10174
rect 22136 10098 22208 10174
rect 22256 10098 22328 10174
rect 504 9223 576 9299
rect 626 9223 698 9299
rect 752 9223 824 9299
rect 504 9076 576 9152
rect 626 9076 698 9152
rect 752 9076 824 9152
rect 504 8939 576 9015
rect 626 8939 698 9015
rect 752 8939 824 9015
rect 503 8563 575 8639
rect 629 8563 701 8639
rect 749 8563 821 8639
rect 503 8445 575 8521
rect 629 8445 701 8521
rect 749 8445 821 8521
rect 21068 8518 21140 8594
rect 21194 8518 21266 8594
rect 21314 8518 21386 8594
rect 21068 8400 21140 8476
rect 21194 8400 21266 8476
rect 21314 8400 21386 8476
rect 503 7452 575 7528
rect 629 7452 701 7528
rect 749 7452 821 7528
rect 503 7334 575 7410
rect 629 7334 701 7410
rect 749 7334 821 7410
rect 21068 7361 21140 7437
rect 21194 7361 21266 7437
rect 21314 7361 21386 7437
rect 21068 7243 21140 7319
rect 21194 7243 21266 7319
rect 21314 7243 21386 7319
rect 504 6985 576 7061
rect 626 6985 698 7061
rect 752 6985 824 7061
rect 504 6838 576 6914
rect 626 6838 698 6914
rect 752 6838 824 6914
rect 504 6701 576 6777
rect 626 6701 698 6777
rect 752 6701 824 6777
rect 22010 6204 22082 6280
rect 22136 6204 22208 6280
rect 22256 6204 22328 6280
rect 22010 6086 22082 6162
rect 22136 6086 22208 6162
rect 22256 6086 22328 6162
rect 504 5224 576 5300
rect 626 5224 698 5300
rect 752 5224 824 5300
rect 504 5077 576 5153
rect 626 5077 698 5153
rect 752 5077 824 5153
rect 504 4940 576 5016
rect 626 4940 698 5016
rect 752 4940 824 5016
rect 503 4629 575 4705
rect 629 4629 701 4705
rect 749 4629 821 4705
rect 503 4511 575 4587
rect 629 4511 701 4587
rect 749 4511 821 4587
rect 21068 4518 21140 4594
rect 21194 4518 21266 4594
rect 21314 4518 21386 4594
rect 21068 4400 21140 4476
rect 21194 4400 21266 4476
rect 21314 4400 21386 4476
rect 503 3452 575 3528
rect 629 3452 701 3528
rect 749 3452 821 3528
rect 503 3334 575 3410
rect 629 3334 701 3410
rect 749 3334 821 3410
rect 21068 3361 21140 3437
rect 21194 3361 21266 3437
rect 21314 3361 21386 3437
rect 21068 3243 21140 3319
rect 21194 3243 21266 3319
rect 21314 3243 21386 3319
rect 504 2985 576 3061
rect 626 2985 698 3061
rect 752 2985 824 3061
rect 504 2838 576 2914
rect 626 2838 698 2914
rect 752 2838 824 2914
rect 504 2701 576 2777
rect 626 2701 698 2777
rect 752 2701 824 2777
rect 22010 2204 22082 2280
rect 22136 2204 22208 2280
rect 22256 2204 22328 2280
rect 22010 2086 22082 2162
rect 22136 2086 22208 2162
rect 22256 2086 22328 2162
rect 504 1224 576 1300
rect 626 1224 698 1300
rect 752 1224 824 1300
rect 504 1077 576 1153
rect 626 1077 698 1153
rect 752 1077 824 1153
rect 504 940 576 1016
rect 626 940 698 1016
rect 752 940 824 1016
rect 503 629 575 705
rect 629 629 701 705
rect 749 629 821 705
rect 503 511 575 587
rect 629 511 701 587
rect 749 511 821 587
rect 21068 518 21140 594
rect 21194 518 21266 594
rect 21314 518 21386 594
rect 21068 400 21140 476
rect 21194 400 21266 476
rect 21314 400 21386 476
<< metal3 >>
rect 21026 75492 21426 75517
rect 463 75452 864 75477
rect 463 75376 503 75452
rect 575 75376 629 75452
rect 701 75376 749 75452
rect 821 75376 864 75452
rect 463 75334 864 75376
rect 463 75258 503 75334
rect 575 75258 629 75334
rect 701 75258 749 75334
rect 821 75258 864 75334
rect 21026 75416 21068 75492
rect 21140 75416 21194 75492
rect 21266 75416 21314 75492
rect 21386 75416 21426 75492
rect 21026 75374 21426 75416
rect 21026 75298 21068 75374
rect 21140 75298 21194 75374
rect 21266 75298 21314 75374
rect 21386 75298 21426 75374
rect 21026 75262 21426 75298
rect 463 75222 864 75258
rect 463 75060 863 75109
rect 463 74984 504 75060
rect 576 74984 626 75060
rect 698 74984 752 75060
rect 824 74984 863 75060
rect 463 74913 863 74984
rect 463 74837 504 74913
rect 576 74837 626 74913
rect 698 74837 752 74913
rect 824 74837 863 74913
rect 463 74776 863 74837
rect 463 74700 504 74776
rect 576 74700 626 74776
rect 698 74700 752 74776
rect 824 74700 863 74776
rect 463 74650 863 74700
rect 21970 74071 22370 74096
rect 21970 73995 22010 74071
rect 22082 73995 22136 74071
rect 22208 73995 22256 74071
rect 22328 73995 22370 74071
rect 21970 73953 22370 73995
rect 21970 73877 22010 73953
rect 22082 73877 22136 73953
rect 22208 73877 22256 73953
rect 22328 73877 22370 73953
rect 21970 73841 22370 73877
rect 463 73300 863 73349
rect 463 73224 504 73300
rect 576 73224 626 73300
rect 698 73224 752 73300
rect 824 73224 863 73300
rect 463 73153 863 73224
rect 463 73077 504 73153
rect 576 73077 626 73153
rect 698 73077 752 73153
rect 824 73077 863 73153
rect 463 73016 863 73077
rect 463 72940 504 73016
rect 576 72940 626 73016
rect 698 72940 752 73016
rect 824 72940 863 73016
rect 463 72890 863 72940
rect 463 72779 864 72804
rect 463 72703 503 72779
rect 575 72703 629 72779
rect 701 72703 749 72779
rect 821 72703 864 72779
rect 463 72661 864 72703
rect 463 72585 503 72661
rect 575 72585 629 72661
rect 701 72585 749 72661
rect 821 72585 864 72661
rect 463 72549 864 72585
rect 21028 72695 21428 72720
rect 21028 72619 21068 72695
rect 21140 72619 21194 72695
rect 21266 72619 21314 72695
rect 21386 72619 21428 72695
rect 21028 72577 21428 72619
rect 21028 72501 21068 72577
rect 21140 72501 21194 72577
rect 21266 72501 21314 72577
rect 21386 72501 21428 72577
rect 21028 72465 21428 72501
rect 21026 71492 21426 71517
rect 463 71452 864 71477
rect 463 71376 503 71452
rect 575 71376 629 71452
rect 701 71376 749 71452
rect 821 71376 864 71452
rect 463 71334 864 71376
rect 463 71258 503 71334
rect 575 71258 629 71334
rect 701 71258 749 71334
rect 821 71258 864 71334
rect 21026 71416 21068 71492
rect 21140 71416 21194 71492
rect 21266 71416 21314 71492
rect 21386 71416 21426 71492
rect 21026 71374 21426 71416
rect 21026 71298 21068 71374
rect 21140 71298 21194 71374
rect 21266 71298 21314 71374
rect 21386 71298 21426 71374
rect 21026 71262 21426 71298
rect 463 71222 864 71258
rect 463 71060 863 71109
rect 463 70984 504 71060
rect 576 70984 626 71060
rect 698 70984 752 71060
rect 824 70984 863 71060
rect 463 70913 863 70984
rect 463 70837 504 70913
rect 576 70837 626 70913
rect 698 70837 752 70913
rect 824 70837 863 70913
rect 463 70776 863 70837
rect 463 70700 504 70776
rect 576 70700 626 70776
rect 698 70700 752 70776
rect 824 70700 863 70776
rect 463 70650 863 70700
rect 21970 70071 22370 70096
rect 21970 69995 22010 70071
rect 22082 69995 22136 70071
rect 22208 69995 22256 70071
rect 22328 69995 22370 70071
rect 21970 69953 22370 69995
rect 21970 69877 22010 69953
rect 22082 69877 22136 69953
rect 22208 69877 22256 69953
rect 22328 69877 22370 69953
rect 21970 69841 22370 69877
rect 463 69300 863 69349
rect 463 69224 504 69300
rect 576 69224 626 69300
rect 698 69224 752 69300
rect 824 69224 863 69300
rect 463 69153 863 69224
rect 463 69077 504 69153
rect 576 69077 626 69153
rect 698 69077 752 69153
rect 824 69077 863 69153
rect 463 69016 863 69077
rect 463 68940 504 69016
rect 576 68940 626 69016
rect 698 68940 752 69016
rect 824 68940 863 69016
rect 463 68890 863 68940
rect 463 68779 864 68804
rect 463 68703 503 68779
rect 575 68703 629 68779
rect 701 68703 749 68779
rect 821 68703 864 68779
rect 463 68661 864 68703
rect 463 68585 503 68661
rect 575 68585 629 68661
rect 701 68585 749 68661
rect 821 68585 864 68661
rect 463 68549 864 68585
rect 21028 68695 21428 68720
rect 21028 68619 21068 68695
rect 21140 68619 21194 68695
rect 21266 68619 21314 68695
rect 21386 68619 21428 68695
rect 21028 68577 21428 68619
rect 21028 68501 21068 68577
rect 21140 68501 21194 68577
rect 21266 68501 21314 68577
rect 21386 68501 21428 68577
rect 21028 68465 21428 68501
rect 21026 67492 21426 67517
rect 463 67450 864 67475
rect 463 67374 503 67450
rect 575 67374 629 67450
rect 701 67374 749 67450
rect 821 67374 864 67450
rect 463 67332 864 67374
rect 463 67256 503 67332
rect 575 67256 629 67332
rect 701 67256 749 67332
rect 821 67256 864 67332
rect 21026 67416 21068 67492
rect 21140 67416 21194 67492
rect 21266 67416 21314 67492
rect 21386 67416 21426 67492
rect 21026 67374 21426 67416
rect 21026 67298 21068 67374
rect 21140 67298 21194 67374
rect 21266 67298 21314 67374
rect 21386 67298 21426 67374
rect 21026 67262 21426 67298
rect 463 67220 864 67256
rect 463 67060 863 67109
rect 463 66984 504 67060
rect 576 66984 626 67060
rect 698 66984 752 67060
rect 824 66984 863 67060
rect 463 66913 863 66984
rect 463 66837 504 66913
rect 576 66837 626 66913
rect 698 66837 752 66913
rect 824 66837 863 66913
rect 463 66776 863 66837
rect 463 66700 504 66776
rect 576 66700 626 66776
rect 698 66700 752 66776
rect 824 66700 863 66776
rect 463 66650 863 66700
rect 21970 66058 22370 66083
rect 21970 65982 22010 66058
rect 22082 65982 22136 66058
rect 22208 65982 22256 66058
rect 22328 65982 22370 66058
rect 21970 65940 22370 65982
rect 21970 65864 22010 65940
rect 22082 65864 22136 65940
rect 22208 65864 22256 65940
rect 22328 65864 22370 65940
rect 21970 65828 22370 65864
rect 463 65301 863 65350
rect 463 65225 504 65301
rect 576 65225 626 65301
rect 698 65225 752 65301
rect 824 65225 863 65301
rect 463 65154 863 65225
rect 463 65078 504 65154
rect 576 65078 626 65154
rect 698 65078 752 65154
rect 824 65078 863 65154
rect 463 65017 863 65078
rect 463 64941 504 65017
rect 576 64941 626 65017
rect 698 64941 752 65017
rect 824 64941 863 65017
rect 463 64891 863 64941
rect 463 64710 864 64735
rect 463 64634 503 64710
rect 575 64634 629 64710
rect 701 64634 749 64710
rect 821 64634 864 64710
rect 463 64592 864 64634
rect 463 64516 503 64592
rect 575 64516 629 64592
rect 701 64516 749 64592
rect 821 64516 864 64592
rect 463 64480 864 64516
rect 21028 64695 21428 64720
rect 21028 64619 21068 64695
rect 21140 64619 21194 64695
rect 21266 64619 21314 64695
rect 21386 64619 21428 64695
rect 21028 64577 21428 64619
rect 21028 64501 21068 64577
rect 21140 64501 21194 64577
rect 21266 64501 21314 64577
rect 21386 64501 21428 64577
rect 21028 64465 21428 64501
rect 463 63532 864 63557
rect 463 63456 503 63532
rect 575 63456 629 63532
rect 701 63456 749 63532
rect 821 63456 864 63532
rect 463 63414 864 63456
rect 463 63338 503 63414
rect 575 63338 629 63414
rect 701 63338 749 63414
rect 821 63338 864 63414
rect 463 63302 864 63338
rect 21026 63492 21426 63517
rect 21026 63416 21068 63492
rect 21140 63416 21194 63492
rect 21266 63416 21314 63492
rect 21386 63416 21426 63492
rect 21026 63374 21426 63416
rect 21026 63298 21068 63374
rect 21140 63298 21194 63374
rect 21266 63298 21314 63374
rect 21386 63298 21426 63374
rect 21026 63262 21426 63298
rect 464 63068 864 63109
rect 463 63060 864 63068
rect 463 62984 504 63060
rect 576 62984 626 63060
rect 698 62984 752 63060
rect 824 62984 864 63060
rect 463 62913 864 62984
rect 463 62837 504 62913
rect 576 62837 626 62913
rect 698 62837 752 62913
rect 824 62837 864 62913
rect 463 62776 864 62837
rect 463 62700 504 62776
rect 576 62700 626 62776
rect 698 62700 752 62776
rect 824 62700 864 62776
rect 463 62650 864 62700
rect 21970 62057 22370 62082
rect 21970 61981 22010 62057
rect 22082 61981 22136 62057
rect 22208 61981 22256 62057
rect 22328 61981 22370 62057
rect 21970 61939 22370 61981
rect 21970 61863 22010 61939
rect 22082 61863 22136 61939
rect 22208 61863 22256 61939
rect 22328 61863 22370 61939
rect 21970 61827 22370 61863
rect 463 61301 863 61350
rect 463 61225 504 61301
rect 576 61225 626 61301
rect 698 61225 752 61301
rect 824 61225 863 61301
rect 463 61154 863 61225
rect 463 61078 504 61154
rect 576 61078 626 61154
rect 698 61078 752 61154
rect 824 61078 863 61154
rect 463 61017 863 61078
rect 463 60941 504 61017
rect 576 60941 626 61017
rect 698 60941 752 61017
rect 824 60941 863 61017
rect 463 60891 863 60941
rect 463 60684 866 60709
rect 463 60608 503 60684
rect 575 60608 629 60684
rect 701 60608 749 60684
rect 821 60608 866 60684
rect 463 60566 866 60608
rect 463 60490 503 60566
rect 575 60490 629 60566
rect 701 60490 749 60566
rect 821 60490 866 60566
rect 463 60454 866 60490
rect 21028 60695 21428 60720
rect 21028 60619 21068 60695
rect 21140 60619 21194 60695
rect 21266 60619 21314 60695
rect 21386 60619 21428 60695
rect 21028 60577 21428 60619
rect 21028 60501 21068 60577
rect 21140 60501 21194 60577
rect 21266 60501 21314 60577
rect 21386 60501 21428 60577
rect 21028 60465 21428 60501
rect 21027 59546 21427 59571
rect 463 59481 864 59506
rect 463 59405 503 59481
rect 575 59405 629 59481
rect 701 59405 749 59481
rect 821 59405 864 59481
rect 463 59363 864 59405
rect 463 59287 503 59363
rect 575 59287 629 59363
rect 701 59287 749 59363
rect 821 59287 864 59363
rect 21027 59470 21068 59546
rect 21140 59470 21194 59546
rect 21266 59470 21314 59546
rect 21386 59470 21427 59546
rect 21027 59428 21427 59470
rect 21027 59352 21068 59428
rect 21140 59352 21194 59428
rect 21266 59352 21314 59428
rect 21386 59352 21427 59428
rect 21027 59316 21427 59352
rect 463 59251 864 59287
rect 464 59068 864 59109
rect 463 59060 864 59068
rect 463 58984 504 59060
rect 576 58984 626 59060
rect 698 58984 752 59060
rect 824 58984 864 59060
rect 463 58913 864 58984
rect 463 58837 504 58913
rect 576 58837 626 58913
rect 698 58837 752 58913
rect 824 58837 864 58913
rect 463 58776 864 58837
rect 463 58700 504 58776
rect 576 58700 626 58776
rect 698 58700 752 58776
rect 824 58700 864 58776
rect 463 58650 864 58700
rect 21970 58096 22370 58121
rect 21970 58020 22010 58096
rect 22082 58020 22136 58096
rect 22208 58020 22256 58096
rect 22328 58020 22370 58096
rect 21970 57978 22370 58020
rect 21970 57902 22010 57978
rect 22082 57902 22136 57978
rect 22208 57902 22256 57978
rect 22328 57902 22370 57978
rect 21970 57866 22370 57902
rect 463 57299 863 57348
rect 463 57223 504 57299
rect 576 57223 626 57299
rect 698 57223 752 57299
rect 824 57223 863 57299
rect 463 57152 863 57223
rect 463 57076 504 57152
rect 576 57076 626 57152
rect 698 57076 752 57152
rect 824 57076 863 57152
rect 463 57015 863 57076
rect 463 56939 504 57015
rect 576 56939 626 57015
rect 698 56939 752 57015
rect 824 56939 863 57015
rect 463 56889 863 56939
rect 463 56704 864 56729
rect 463 56628 503 56704
rect 575 56628 629 56704
rect 701 56628 749 56704
rect 821 56628 864 56704
rect 463 56586 864 56628
rect 463 56510 503 56586
rect 575 56510 629 56586
rect 701 56510 749 56586
rect 821 56510 864 56586
rect 463 56474 864 56510
rect 21028 56630 21428 56655
rect 21028 56554 21068 56630
rect 21140 56554 21194 56630
rect 21266 56554 21314 56630
rect 21386 56554 21428 56630
rect 21028 56512 21428 56554
rect 21028 56436 21068 56512
rect 21140 56436 21194 56512
rect 21266 56436 21314 56512
rect 21386 56436 21428 56512
rect 21028 56400 21428 56436
rect 463 55497 866 55522
rect 463 55421 503 55497
rect 575 55421 629 55497
rect 701 55421 749 55497
rect 821 55421 866 55497
rect 463 55379 866 55421
rect 463 55303 503 55379
rect 575 55303 629 55379
rect 701 55303 749 55379
rect 821 55303 866 55379
rect 463 55267 866 55303
rect 21027 55447 21427 55472
rect 21027 55371 21068 55447
rect 21140 55371 21194 55447
rect 21266 55371 21314 55447
rect 21386 55371 21427 55447
rect 21027 55329 21427 55371
rect 21027 55253 21068 55329
rect 21140 55253 21194 55329
rect 21266 55253 21314 55329
rect 21386 55253 21427 55329
rect 21027 55217 21427 55253
rect 463 55060 863 55109
rect 463 54984 504 55060
rect 576 54984 626 55060
rect 698 54984 752 55060
rect 824 54984 863 55060
rect 463 54913 863 54984
rect 463 54837 504 54913
rect 576 54837 626 54913
rect 698 54837 752 54913
rect 824 54837 863 54913
rect 463 54776 863 54837
rect 463 54700 504 54776
rect 576 54700 626 54776
rect 698 54700 752 54776
rect 824 54700 863 54776
rect 463 54650 863 54700
rect 21970 54079 22370 54104
rect 21970 54003 22010 54079
rect 22082 54003 22136 54079
rect 22208 54003 22256 54079
rect 22328 54003 22370 54079
rect 21970 53961 22370 54003
rect 21970 53885 22010 53961
rect 22082 53885 22136 53961
rect 22208 53885 22256 53961
rect 22328 53885 22370 53961
rect 21970 53849 22370 53885
rect 463 53301 863 53350
rect 463 53225 504 53301
rect 576 53225 626 53301
rect 698 53225 752 53301
rect 824 53225 863 53301
rect 463 53154 863 53225
rect 463 53078 504 53154
rect 576 53078 626 53154
rect 698 53078 752 53154
rect 824 53078 863 53154
rect 463 53017 863 53078
rect 463 52941 504 53017
rect 576 52941 626 53017
rect 698 52941 752 53017
rect 824 52941 863 53017
rect 463 52891 863 52941
rect 463 52731 864 52756
rect 463 52655 503 52731
rect 575 52655 629 52731
rect 701 52655 749 52731
rect 821 52655 864 52731
rect 463 52613 864 52655
rect 463 52537 503 52613
rect 575 52537 629 52613
rect 701 52537 749 52613
rect 821 52537 864 52613
rect 463 52501 864 52537
rect 21028 52575 21428 52600
rect 21028 52499 21068 52575
rect 21140 52499 21194 52575
rect 21266 52499 21314 52575
rect 21386 52499 21428 52575
rect 21028 52457 21428 52499
rect 21028 52381 21068 52457
rect 21140 52381 21194 52457
rect 21266 52381 21314 52457
rect 21386 52381 21428 52457
rect 21028 52345 21428 52381
rect 463 51544 864 51569
rect 463 51468 503 51544
rect 575 51468 629 51544
rect 701 51468 749 51544
rect 821 51468 864 51544
rect 463 51426 864 51468
rect 463 51350 503 51426
rect 575 51350 629 51426
rect 701 51350 749 51426
rect 821 51350 864 51426
rect 463 51314 864 51350
rect 21028 51440 21428 51465
rect 21028 51364 21068 51440
rect 21140 51364 21194 51440
rect 21266 51364 21314 51440
rect 21386 51364 21428 51440
rect 21028 51322 21428 51364
rect 21028 51246 21068 51322
rect 21140 51246 21194 51322
rect 21266 51246 21314 51322
rect 21386 51246 21428 51322
rect 21028 51210 21428 51246
rect 463 51060 863 51109
rect 463 50984 504 51060
rect 576 50984 626 51060
rect 698 50984 752 51060
rect 824 50984 863 51060
rect 463 50913 863 50984
rect 463 50837 504 50913
rect 576 50837 626 50913
rect 698 50837 752 50913
rect 824 50837 863 50913
rect 463 50776 863 50837
rect 463 50700 504 50776
rect 576 50700 626 50776
rect 698 50700 752 50776
rect 824 50700 863 50776
rect 463 50650 863 50700
rect 21970 50158 22370 50183
rect 21970 50082 22010 50158
rect 22082 50082 22136 50158
rect 22208 50082 22256 50158
rect 22328 50082 22370 50158
rect 21970 50040 22370 50082
rect 21970 49964 22010 50040
rect 22082 49964 22136 50040
rect 22208 49964 22256 50040
rect 22328 49964 22370 50040
rect 21970 49928 22370 49964
rect 463 49301 863 49350
rect 463 49225 504 49301
rect 576 49225 626 49301
rect 698 49225 752 49301
rect 824 49225 863 49301
rect 463 49154 863 49225
rect 463 49078 504 49154
rect 576 49078 626 49154
rect 698 49078 752 49154
rect 824 49078 863 49154
rect 463 49017 863 49078
rect 463 48941 504 49017
rect 576 48941 626 49017
rect 698 48941 752 49017
rect 824 48941 863 49017
rect 463 48891 863 48941
rect 463 48722 864 48747
rect 463 48646 503 48722
rect 575 48646 629 48722
rect 701 48646 749 48722
rect 821 48646 864 48722
rect 463 48604 864 48646
rect 463 48528 503 48604
rect 575 48528 629 48604
rect 701 48528 749 48604
rect 821 48528 864 48604
rect 463 48492 864 48528
rect 21028 48681 21428 48706
rect 21028 48605 21068 48681
rect 21140 48605 21194 48681
rect 21266 48605 21314 48681
rect 21386 48605 21428 48681
rect 21028 48563 21428 48605
rect 21028 48487 21068 48563
rect 21140 48487 21194 48563
rect 21266 48487 21314 48563
rect 21386 48487 21428 48563
rect 21028 48451 21428 48487
rect 463 47569 864 47594
rect 463 47493 503 47569
rect 575 47493 629 47569
rect 701 47493 749 47569
rect 821 47493 864 47569
rect 463 47451 864 47493
rect 463 47375 503 47451
rect 575 47375 629 47451
rect 701 47375 749 47451
rect 821 47375 864 47451
rect 463 47339 864 47375
rect 21028 47528 21428 47553
rect 21028 47452 21068 47528
rect 21140 47452 21194 47528
rect 21266 47452 21314 47528
rect 21386 47452 21428 47528
rect 21028 47410 21428 47452
rect 21028 47334 21068 47410
rect 21140 47334 21194 47410
rect 21266 47334 21314 47410
rect 21386 47334 21428 47410
rect 21028 47298 21428 47334
rect 463 47060 863 47109
rect 463 46984 504 47060
rect 576 46984 626 47060
rect 698 46984 752 47060
rect 824 46984 863 47060
rect 463 46913 863 46984
rect 463 46837 504 46913
rect 576 46837 626 46913
rect 698 46837 752 46913
rect 824 46837 863 46913
rect 463 46776 863 46837
rect 463 46700 504 46776
rect 576 46700 626 46776
rect 698 46700 752 46776
rect 824 46700 863 46776
rect 463 46650 863 46700
rect 21970 45900 22370 45925
rect 21970 45824 22010 45900
rect 22082 45824 22136 45900
rect 22208 45824 22256 45900
rect 22328 45824 22370 45900
rect 21970 45782 22370 45824
rect 21970 45706 22010 45782
rect 22082 45706 22136 45782
rect 22208 45706 22256 45782
rect 22328 45706 22370 45782
rect 21970 45670 22370 45706
rect 463 45300 863 45350
rect 463 45224 504 45300
rect 576 45224 626 45300
rect 698 45224 752 45300
rect 824 45224 863 45300
rect 463 45153 863 45224
rect 463 45077 504 45153
rect 576 45077 626 45153
rect 698 45077 752 45153
rect 824 45077 863 45153
rect 463 45016 863 45077
rect 463 44940 504 45016
rect 576 44940 626 45016
rect 698 44940 752 45016
rect 824 44940 863 45016
rect 463 44891 863 44940
rect 463 44890 836 44891
rect 463 44509 863 44534
rect 463 44433 503 44509
rect 575 44433 629 44509
rect 701 44433 749 44509
rect 821 44433 863 44509
rect 463 44391 863 44433
rect 463 44315 503 44391
rect 575 44315 629 44391
rect 701 44315 749 44391
rect 821 44315 863 44391
rect 463 44279 863 44315
rect 21028 44412 21428 44437
rect 21028 44336 21068 44412
rect 21140 44336 21194 44412
rect 21266 44336 21314 44412
rect 21386 44336 21428 44412
rect 21028 44294 21428 44336
rect 21028 44218 21068 44294
rect 21140 44218 21194 44294
rect 21266 44218 21314 44294
rect 21386 44218 21428 44294
rect 21028 44182 21428 44218
rect 21970 43838 22370 43870
rect 21970 43514 22006 43838
rect 22298 43514 22370 43838
rect 21970 43480 22370 43514
rect 2248 39925 2401 39940
rect 2248 39861 2249 39925
rect 2313 39861 2337 39925
rect 2248 39845 2401 39861
rect 2248 39781 2249 39845
rect 2313 39781 2337 39845
rect 2248 39775 2401 39781
rect 3352 39905 4345 39920
rect 3352 39904 4192 39905
rect 3352 39848 3361 39904
rect 3417 39848 3441 39904
rect 3497 39848 4192 39904
rect 3352 39841 4192 39848
rect 4256 39841 4280 39905
rect 4344 39841 4345 39905
rect 3352 39825 4345 39841
rect 3352 39824 4192 39825
rect 3352 39768 3361 39824
rect 3417 39768 3441 39824
rect 3497 39768 4192 39824
rect 3352 39761 4192 39768
rect 4256 39761 4280 39825
rect 4344 39761 4345 39825
rect 3352 39754 4345 39761
rect 0 39741 400 39752
rect 0 39661 32 39741
rect 112 39661 156 39741
rect 237 39661 282 39741
rect 362 39661 400 39741
rect 0 39635 400 39661
rect 0 39555 32 39635
rect 112 39555 156 39635
rect 237 39555 282 39635
rect 362 39555 400 39635
rect 0 39528 400 39555
rect 21502 39726 21902 39752
rect 21502 39646 21535 39726
rect 21615 39646 21660 39726
rect 21740 39646 21785 39726
rect 21865 39646 21902 39726
rect 21502 39606 21902 39646
rect 21502 39526 21534 39606
rect 21614 39526 21659 39606
rect 21739 39526 21784 39606
rect 21864 39526 21902 39606
rect 21502 39497 21902 39526
rect 2689 39333 3502 39334
rect 1411 39320 3502 39333
rect 1411 39319 1498 39320
rect 1411 39263 1416 39319
rect 1472 39264 1498 39319
rect 1554 39318 3502 39320
rect 1554 39264 2760 39318
rect 1472 39263 2760 39264
rect 1411 39262 2760 39263
rect 2816 39317 3502 39318
rect 2816 39262 2840 39317
rect 1411 39261 2840 39262
rect 2896 39261 3360 39317
rect 3416 39316 3502 39317
rect 3416 39261 3440 39316
rect 1411 39260 3440 39261
rect 3496 39260 3502 39316
rect 1411 39240 3502 39260
rect 1411 39239 1499 39240
rect 1411 39183 1417 39239
rect 1473 39184 1499 39239
rect 1555 39237 3502 39240
rect 1555 39184 2761 39237
rect 1473 39183 2761 39184
rect 1411 39181 2761 39183
rect 2817 39181 2841 39237
rect 2897 39236 3502 39237
rect 2897 39181 3361 39236
rect 1411 39180 3361 39181
rect 3417 39180 3441 39236
rect 3497 39180 3502 39236
rect 1411 39169 3502 39180
rect 463 39131 805 39139
rect 463 39051 478 39131
rect 562 39051 592 39131
rect 676 39051 706 39131
rect 790 39051 805 39131
rect 463 39043 805 39051
rect 0 38587 342 38595
rect 0 38507 15 38587
rect 99 38507 129 38587
rect 213 38507 243 38587
rect 327 38507 342 38587
rect 0 38499 342 38507
rect 463 38043 805 38051
rect 463 37963 478 38043
rect 562 37963 592 38043
rect 676 37963 706 38043
rect 790 37963 805 38043
rect 463 37955 805 37963
rect 0 37499 342 37507
rect 0 37419 15 37499
rect 99 37419 129 37499
rect 213 37419 243 37499
rect 327 37419 342 37499
rect 0 37411 342 37419
rect 463 36955 805 36963
rect 463 36875 478 36955
rect 562 36875 592 36955
rect 676 36875 706 36955
rect 790 36875 805 36955
rect 463 36867 805 36875
rect 21970 36954 22370 36986
rect 21970 36630 22006 36954
rect 22298 36630 22370 36954
rect 21970 36596 22370 36630
rect 2535 36475 2688 36476
rect 2535 36463 2689 36475
rect 2535 36399 2536 36463
rect 2600 36399 2624 36463
rect 2688 36399 2689 36463
rect 2535 36391 2689 36399
rect 21028 36172 21428 36198
rect 21028 36092 21061 36172
rect 21141 36092 21186 36172
rect 21266 36092 21311 36172
rect 21391 36092 21428 36172
rect 21028 36052 21428 36092
rect 21028 35972 21060 36052
rect 21140 35972 21185 36052
rect 21265 35972 21310 36052
rect 21390 35972 21428 36052
rect 21028 35943 21428 35972
rect 21028 35592 21428 35642
rect 21028 35516 21069 35592
rect 21141 35516 21191 35592
rect 21263 35516 21317 35592
rect 21389 35516 21428 35592
rect 21028 35445 21428 35516
rect 21028 35369 21069 35445
rect 21141 35369 21191 35445
rect 21263 35369 21317 35445
rect 21389 35369 21428 35445
rect 21028 35308 21428 35369
rect 21028 35232 21069 35308
rect 21141 35232 21191 35308
rect 21263 35232 21317 35308
rect 21389 35232 21428 35308
rect 21028 35183 21428 35232
rect 21028 35182 21401 35183
rect 20527 34676 20927 34702
rect 20527 34596 20560 34676
rect 20640 34596 20685 34676
rect 20765 34596 20810 34676
rect 20890 34596 20927 34676
rect 20527 34556 20927 34596
rect 20527 34476 20559 34556
rect 20639 34476 20684 34556
rect 20764 34476 20809 34556
rect 20889 34476 20927 34556
rect 20527 34447 20927 34476
rect 21502 34676 21902 34702
rect 21502 34596 21535 34676
rect 21615 34596 21660 34676
rect 21740 34596 21785 34676
rect 21865 34596 21902 34676
rect 21502 34556 21902 34596
rect 21502 34476 21534 34556
rect 21614 34476 21659 34556
rect 21739 34476 21784 34556
rect 21864 34476 21902 34556
rect 21502 34447 21902 34476
rect 21028 33832 21428 33882
rect 21028 33756 21069 33832
rect 21141 33756 21191 33832
rect 21263 33756 21317 33832
rect 21389 33756 21428 33832
rect 21028 33685 21428 33756
rect 21028 33609 21069 33685
rect 21141 33609 21191 33685
rect 21263 33609 21317 33685
rect 21389 33609 21428 33685
rect 21028 33548 21428 33609
rect 21028 33472 21069 33548
rect 21141 33472 21191 33548
rect 21263 33472 21317 33548
rect 21389 33472 21428 33548
rect 21028 33423 21428 33472
rect 21028 33422 21401 33423
rect 21027 33117 21427 33143
rect 21027 33037 21060 33117
rect 21140 33037 21185 33117
rect 21265 33037 21310 33117
rect 21390 33037 21427 33117
rect 21027 32997 21427 33037
rect 21027 32917 21059 32997
rect 21139 32917 21184 32997
rect 21264 32917 21309 32997
rect 21389 32917 21427 32997
rect 21027 32888 21427 32917
rect 463 32302 866 32360
rect 463 32226 503 32302
rect 575 32226 629 32302
rect 701 32226 749 32302
rect 821 32226 866 32302
rect 463 32184 866 32226
rect 463 32108 503 32184
rect 575 32108 629 32184
rect 701 32108 749 32184
rect 821 32108 866 32184
rect 463 32072 866 32108
rect 21025 32302 21428 32360
rect 21025 32226 21068 32302
rect 21140 32226 21194 32302
rect 21266 32226 21314 32302
rect 21386 32226 21428 32302
rect 21025 32184 21428 32226
rect 21025 32108 21068 32184
rect 21140 32108 21194 32184
rect 21266 32108 21314 32184
rect 21386 32108 21428 32184
rect 21025 32072 21428 32108
rect 463 31520 863 31545
rect 463 31444 503 31520
rect 575 31444 629 31520
rect 701 31444 749 31520
rect 821 31444 863 31520
rect 463 31402 863 31444
rect 463 31326 503 31402
rect 575 31326 629 31402
rect 701 31326 749 31402
rect 821 31326 863 31402
rect 463 31290 863 31326
rect 21028 31520 21428 31545
rect 21028 31444 21068 31520
rect 21140 31444 21194 31520
rect 21266 31444 21314 31520
rect 21386 31444 21428 31520
rect 21028 31402 21428 31444
rect 21028 31326 21068 31402
rect 21140 31326 21194 31402
rect 21266 31326 21314 31402
rect 21386 31326 21428 31402
rect 21028 31290 21428 31326
rect 463 31061 863 31111
rect 463 30985 504 31061
rect 576 30985 626 31061
rect 698 30985 752 31061
rect 824 30985 863 31061
rect 463 30914 863 30985
rect 463 30838 504 30914
rect 576 30838 626 30914
rect 698 30838 752 30914
rect 824 30838 863 30914
rect 463 30777 863 30838
rect 463 30701 504 30777
rect 576 30701 626 30777
rect 698 30701 752 30777
rect 824 30701 863 30777
rect 463 30651 863 30701
rect 21970 30130 22370 30155
rect 21970 30054 22010 30130
rect 22082 30054 22136 30130
rect 22208 30054 22256 30130
rect 22328 30054 22370 30130
rect 21970 30012 22370 30054
rect 21970 29936 22010 30012
rect 22082 29936 22136 30012
rect 22208 29936 22256 30012
rect 22328 29936 22370 30012
rect 21970 29900 22370 29936
rect 463 29294 863 29349
rect 463 29218 504 29294
rect 576 29218 626 29294
rect 698 29218 752 29294
rect 824 29218 863 29294
rect 463 29147 863 29218
rect 463 29071 504 29147
rect 576 29071 626 29147
rect 698 29071 752 29147
rect 824 29071 863 29147
rect 463 29010 863 29071
rect 463 28934 504 29010
rect 576 28934 626 29010
rect 698 28934 752 29010
rect 824 28934 863 29010
rect 463 28890 863 28934
rect 463 28608 863 28633
rect 463 28532 503 28608
rect 575 28532 629 28608
rect 701 28532 749 28608
rect 821 28532 863 28608
rect 463 28490 863 28532
rect 463 28414 503 28490
rect 575 28414 629 28490
rect 701 28414 749 28490
rect 821 28414 863 28490
rect 463 28378 863 28414
rect 21028 28559 21428 28584
rect 21028 28483 21068 28559
rect 21140 28483 21194 28559
rect 21266 28483 21314 28559
rect 21386 28483 21428 28559
rect 21028 28441 21428 28483
rect 21028 28365 21068 28441
rect 21140 28365 21194 28441
rect 21266 28365 21314 28441
rect 21386 28365 21428 28441
rect 21028 28329 21428 28365
rect 463 27604 863 27629
rect 463 27528 503 27604
rect 575 27528 629 27604
rect 701 27528 749 27604
rect 821 27528 863 27604
rect 463 27486 863 27528
rect 463 27410 503 27486
rect 575 27410 629 27486
rect 701 27410 749 27486
rect 821 27410 863 27486
rect 463 27374 863 27410
rect 21027 27442 21427 27467
rect 21027 27366 21068 27442
rect 21140 27366 21194 27442
rect 21266 27366 21314 27442
rect 21386 27366 21427 27442
rect 21027 27324 21427 27366
rect 21027 27248 21068 27324
rect 21140 27248 21194 27324
rect 21266 27248 21314 27324
rect 21386 27248 21427 27324
rect 21027 27212 21427 27248
rect 463 27060 863 27109
rect 463 26984 504 27060
rect 576 26984 626 27060
rect 698 26984 752 27060
rect 824 26984 863 27060
rect 463 26913 863 26984
rect 463 26837 504 26913
rect 576 26837 626 26913
rect 698 26837 752 26913
rect 824 26837 863 26913
rect 463 26776 863 26837
rect 463 26700 504 26776
rect 576 26700 626 26776
rect 698 26700 752 26776
rect 824 26700 863 26776
rect 463 26650 863 26700
rect 21970 25971 22370 25996
rect 21970 25895 22010 25971
rect 22082 25895 22136 25971
rect 22208 25895 22256 25971
rect 22328 25895 22370 25971
rect 21970 25853 22370 25895
rect 21970 25777 22010 25853
rect 22082 25777 22136 25853
rect 22208 25777 22256 25853
rect 22328 25777 22370 25853
rect 21970 25741 22370 25777
rect 463 25300 863 25349
rect 463 25224 504 25300
rect 576 25224 626 25300
rect 698 25224 752 25300
rect 824 25224 863 25300
rect 463 25153 863 25224
rect 463 25077 504 25153
rect 576 25077 626 25153
rect 698 25077 752 25153
rect 824 25077 863 25153
rect 463 25016 863 25077
rect 463 24940 504 25016
rect 576 24940 626 25016
rect 698 24940 752 25016
rect 824 24940 863 25016
rect 463 24890 863 24940
rect 463 24626 864 24651
rect 463 24550 503 24626
rect 575 24550 629 24626
rect 701 24550 749 24626
rect 821 24550 864 24626
rect 463 24508 864 24550
rect 463 24432 503 24508
rect 575 24432 629 24508
rect 701 24432 749 24508
rect 821 24432 864 24508
rect 463 24396 864 24432
rect 21028 24599 21428 24624
rect 21028 24523 21068 24599
rect 21140 24523 21194 24599
rect 21266 24523 21314 24599
rect 21386 24523 21428 24599
rect 21028 24481 21428 24523
rect 21028 24405 21068 24481
rect 21140 24405 21194 24481
rect 21266 24405 21314 24481
rect 21386 24405 21428 24481
rect 21028 24369 21428 24405
rect 463 23544 864 23569
rect 463 23468 503 23544
rect 575 23468 629 23544
rect 701 23468 749 23544
rect 821 23468 864 23544
rect 463 23426 864 23468
rect 463 23350 503 23426
rect 575 23350 629 23426
rect 701 23350 749 23426
rect 821 23350 864 23426
rect 463 23314 864 23350
rect 21028 23424 21428 23449
rect 21028 23348 21068 23424
rect 21140 23348 21194 23424
rect 21266 23348 21314 23424
rect 21386 23348 21428 23424
rect 21028 23306 21428 23348
rect 21028 23230 21068 23306
rect 21140 23230 21194 23306
rect 21266 23230 21314 23306
rect 21386 23230 21428 23306
rect 21028 23194 21428 23230
rect 463 23060 863 23109
rect 463 22984 504 23060
rect 576 22984 626 23060
rect 698 22984 752 23060
rect 824 22984 863 23060
rect 463 22913 863 22984
rect 463 22837 504 22913
rect 576 22837 626 22913
rect 698 22837 752 22913
rect 824 22837 863 22913
rect 463 22776 863 22837
rect 463 22700 504 22776
rect 576 22700 626 22776
rect 698 22700 752 22776
rect 824 22700 863 22776
rect 463 22650 863 22700
rect 21970 22181 22370 22206
rect 21970 22105 22010 22181
rect 22082 22105 22136 22181
rect 22208 22105 22256 22181
rect 22328 22105 22370 22181
rect 21970 22063 22370 22105
rect 21970 21987 22010 22063
rect 22082 21987 22136 22063
rect 22208 21987 22256 22063
rect 22328 21987 22370 22063
rect 21970 21951 22370 21987
rect 463 21301 863 21350
rect 463 21225 504 21301
rect 576 21225 626 21301
rect 698 21225 752 21301
rect 824 21225 863 21301
rect 463 21154 863 21225
rect 463 21078 504 21154
rect 576 21078 626 21154
rect 698 21078 752 21154
rect 824 21078 863 21154
rect 463 21017 863 21078
rect 463 20941 504 21017
rect 576 20941 626 21017
rect 698 20941 752 21017
rect 824 20941 863 21017
rect 463 20891 863 20941
rect 463 20669 864 20694
rect 463 20593 503 20669
rect 575 20593 629 20669
rect 701 20593 749 20669
rect 821 20593 864 20669
rect 463 20551 864 20593
rect 463 20475 503 20551
rect 575 20475 629 20551
rect 701 20475 749 20551
rect 821 20475 864 20551
rect 463 20439 864 20475
rect 21027 20583 21427 20608
rect 21027 20507 21068 20583
rect 21140 20507 21194 20583
rect 21266 20507 21314 20583
rect 21386 20507 21427 20583
rect 21027 20465 21427 20507
rect 21027 20389 21068 20465
rect 21140 20389 21194 20465
rect 21266 20389 21314 20465
rect 21386 20389 21427 20465
rect 21027 20353 21427 20389
rect 463 19568 864 19593
rect 463 19492 503 19568
rect 575 19492 629 19568
rect 701 19492 749 19568
rect 821 19492 864 19568
rect 463 19450 864 19492
rect 463 19374 503 19450
rect 575 19374 629 19450
rect 701 19374 749 19450
rect 821 19374 864 19450
rect 463 19338 864 19374
rect 21027 19412 21427 19437
rect 21027 19336 21068 19412
rect 21140 19336 21194 19412
rect 21266 19336 21314 19412
rect 21386 19336 21427 19412
rect 21027 19294 21427 19336
rect 21027 19218 21068 19294
rect 21140 19218 21194 19294
rect 21266 19218 21314 19294
rect 21386 19218 21427 19294
rect 21027 19182 21427 19218
rect 463 19060 863 19109
rect 463 18984 504 19060
rect 576 18984 626 19060
rect 698 18984 752 19060
rect 824 18984 863 19060
rect 463 18913 863 18984
rect 463 18837 504 18913
rect 576 18837 626 18913
rect 698 18837 752 18913
rect 824 18837 863 18913
rect 463 18776 863 18837
rect 463 18700 504 18776
rect 576 18700 626 18776
rect 698 18700 752 18776
rect 824 18700 863 18776
rect 463 18650 863 18700
rect 21970 18074 22370 18099
rect 21970 17998 22010 18074
rect 22082 17998 22136 18074
rect 22208 17998 22256 18074
rect 22328 17998 22370 18074
rect 21970 17956 22370 17998
rect 21970 17880 22010 17956
rect 22082 17880 22136 17956
rect 22208 17880 22256 17956
rect 22328 17880 22370 17956
rect 21970 17844 22370 17880
rect 463 17300 863 17349
rect 463 17224 504 17300
rect 576 17224 626 17300
rect 698 17224 752 17300
rect 824 17224 863 17300
rect 463 17153 863 17224
rect 463 17077 504 17153
rect 576 17077 626 17153
rect 698 17077 752 17153
rect 824 17077 863 17153
rect 463 17016 863 17077
rect 463 16940 504 17016
rect 576 16940 626 17016
rect 698 16940 752 17016
rect 824 16940 863 17016
rect 463 16890 863 16940
rect 463 16702 865 16727
rect 463 16626 503 16702
rect 575 16626 629 16702
rect 701 16626 749 16702
rect 821 16626 865 16702
rect 463 16584 865 16626
rect 463 16508 503 16584
rect 575 16508 629 16584
rect 701 16508 749 16584
rect 821 16508 865 16584
rect 463 16472 865 16508
rect 21027 16651 21427 16676
rect 21027 16575 21068 16651
rect 21140 16575 21194 16651
rect 21266 16575 21314 16651
rect 21386 16575 21427 16651
rect 21027 16533 21427 16575
rect 21027 16457 21068 16533
rect 21140 16457 21194 16533
rect 21266 16457 21314 16533
rect 21386 16457 21427 16533
rect 21027 16421 21427 16457
rect 463 15486 866 15511
rect 463 15410 503 15486
rect 575 15410 629 15486
rect 701 15410 749 15486
rect 821 15410 866 15486
rect 463 15368 866 15410
rect 463 15292 503 15368
rect 575 15292 629 15368
rect 701 15292 749 15368
rect 821 15292 866 15368
rect 463 15256 866 15292
rect 21027 15437 21427 15462
rect 21027 15361 21068 15437
rect 21140 15361 21194 15437
rect 21266 15361 21314 15437
rect 21386 15361 21427 15437
rect 21027 15319 21427 15361
rect 21027 15243 21068 15319
rect 21140 15243 21194 15319
rect 21266 15243 21314 15319
rect 21386 15243 21427 15319
rect 21027 15207 21427 15243
rect 463 15060 863 15109
rect 463 14984 504 15060
rect 576 14984 626 15060
rect 698 14984 752 15060
rect 824 14984 863 15060
rect 463 14913 863 14984
rect 463 14837 504 14913
rect 576 14837 626 14913
rect 698 14837 752 14913
rect 824 14837 863 14913
rect 463 14776 863 14837
rect 463 14700 504 14776
rect 576 14700 626 14776
rect 698 14700 752 14776
rect 824 14700 863 14776
rect 463 14650 863 14700
rect 21970 14256 22370 14281
rect 21970 14180 22010 14256
rect 22082 14180 22136 14256
rect 22208 14180 22256 14256
rect 22328 14180 22370 14256
rect 21970 14138 22370 14180
rect 21970 14062 22010 14138
rect 22082 14062 22136 14138
rect 22208 14062 22256 14138
rect 22328 14062 22370 14138
rect 21970 14026 22370 14062
rect 463 13300 863 13349
rect 463 13224 504 13300
rect 576 13224 626 13300
rect 698 13224 752 13300
rect 824 13224 863 13300
rect 463 13153 863 13224
rect 463 13077 504 13153
rect 576 13077 626 13153
rect 698 13077 752 13153
rect 824 13077 863 13153
rect 463 13016 863 13077
rect 463 12940 504 13016
rect 576 12940 626 13016
rect 698 12940 752 13016
rect 824 12940 863 13016
rect 463 12890 863 12940
rect 463 12621 864 12646
rect 463 12545 503 12621
rect 575 12545 629 12621
rect 701 12545 749 12621
rect 821 12545 864 12621
rect 463 12503 864 12545
rect 463 12427 503 12503
rect 575 12427 629 12503
rect 701 12427 749 12503
rect 821 12427 864 12503
rect 463 12391 864 12427
rect 21028 12594 21428 12619
rect 21028 12518 21068 12594
rect 21140 12518 21194 12594
rect 21266 12518 21314 12594
rect 21386 12518 21428 12594
rect 21028 12476 21428 12518
rect 21028 12400 21068 12476
rect 21140 12400 21194 12476
rect 21266 12400 21314 12476
rect 21386 12400 21428 12476
rect 21028 12364 21428 12400
rect 463 11499 864 11524
rect 463 11423 503 11499
rect 575 11423 629 11499
rect 701 11423 749 11499
rect 821 11423 864 11499
rect 463 11381 864 11423
rect 463 11305 503 11381
rect 575 11305 629 11381
rect 701 11305 749 11381
rect 821 11305 864 11381
rect 463 11269 864 11305
rect 21027 11437 21427 11462
rect 21027 11361 21068 11437
rect 21140 11361 21194 11437
rect 21266 11361 21314 11437
rect 21386 11361 21427 11437
rect 21027 11319 21427 11361
rect 21027 11243 21068 11319
rect 21140 11243 21194 11319
rect 21266 11243 21314 11319
rect 21386 11243 21427 11319
rect 21027 11207 21427 11243
rect 463 11061 863 11110
rect 463 10985 504 11061
rect 576 10985 626 11061
rect 698 10985 752 11061
rect 824 10985 863 11061
rect 463 10914 863 10985
rect 463 10838 504 10914
rect 576 10838 626 10914
rect 698 10838 752 10914
rect 824 10838 863 10914
rect 463 10777 863 10838
rect 463 10701 504 10777
rect 576 10701 626 10777
rect 698 10701 752 10777
rect 824 10701 863 10777
rect 463 10651 863 10701
rect 21970 10292 22370 10317
rect 21970 10216 22010 10292
rect 22082 10216 22136 10292
rect 22208 10216 22256 10292
rect 22328 10216 22370 10292
rect 21970 10174 22370 10216
rect 21970 10098 22010 10174
rect 22082 10098 22136 10174
rect 22208 10098 22256 10174
rect 22328 10098 22370 10174
rect 21970 10062 22370 10098
rect 463 9299 863 9348
rect 463 9223 504 9299
rect 576 9223 626 9299
rect 698 9223 752 9299
rect 824 9223 863 9299
rect 463 9152 863 9223
rect 463 9076 504 9152
rect 576 9076 626 9152
rect 698 9076 752 9152
rect 824 9076 863 9152
rect 463 9015 863 9076
rect 463 8939 504 9015
rect 576 8939 626 9015
rect 698 8939 752 9015
rect 824 8939 863 9015
rect 463 8889 863 8939
rect 463 8639 863 8664
rect 463 8563 503 8639
rect 575 8563 629 8639
rect 701 8563 749 8639
rect 821 8563 863 8639
rect 463 8521 863 8563
rect 463 8445 503 8521
rect 575 8445 629 8521
rect 701 8445 749 8521
rect 821 8445 863 8521
rect 463 8409 863 8445
rect 21028 8594 21428 8619
rect 21028 8518 21068 8594
rect 21140 8518 21194 8594
rect 21266 8518 21314 8594
rect 21386 8518 21428 8594
rect 21028 8476 21428 8518
rect 21028 8400 21068 8476
rect 21140 8400 21194 8476
rect 21266 8400 21314 8476
rect 21386 8400 21428 8476
rect 21028 8364 21428 8400
rect 463 7528 863 7553
rect 463 7452 503 7528
rect 575 7452 629 7528
rect 701 7452 749 7528
rect 821 7452 863 7528
rect 463 7410 863 7452
rect 463 7334 503 7410
rect 575 7334 629 7410
rect 701 7334 749 7410
rect 821 7334 863 7410
rect 463 7298 863 7334
rect 21027 7437 21427 7462
rect 21027 7361 21068 7437
rect 21140 7361 21194 7437
rect 21266 7361 21314 7437
rect 21386 7361 21427 7437
rect 21027 7319 21427 7361
rect 21027 7243 21068 7319
rect 21140 7243 21194 7319
rect 21266 7243 21314 7319
rect 21386 7243 21427 7319
rect 21027 7207 21427 7243
rect 463 7061 863 7110
rect 463 6985 504 7061
rect 576 6985 626 7061
rect 698 6985 752 7061
rect 824 6985 863 7061
rect 463 6914 863 6985
rect 463 6838 504 6914
rect 576 6838 626 6914
rect 698 6838 752 6914
rect 824 6838 863 6914
rect 463 6777 863 6838
rect 463 6701 504 6777
rect 576 6701 626 6777
rect 698 6701 752 6777
rect 824 6701 863 6777
rect 463 6651 863 6701
rect 21970 6280 22370 6305
rect 21970 6204 22010 6280
rect 22082 6204 22136 6280
rect 22208 6204 22256 6280
rect 22328 6204 22370 6280
rect 21970 6162 22370 6204
rect 21970 6086 22010 6162
rect 22082 6086 22136 6162
rect 22208 6086 22256 6162
rect 22328 6086 22370 6162
rect 21970 6050 22370 6086
rect 463 5300 863 5349
rect 463 5224 504 5300
rect 576 5224 626 5300
rect 698 5224 752 5300
rect 824 5224 863 5300
rect 463 5153 863 5224
rect 463 5077 504 5153
rect 576 5077 626 5153
rect 698 5077 752 5153
rect 824 5077 863 5153
rect 463 5016 863 5077
rect 463 4940 504 5016
rect 576 4940 626 5016
rect 698 4940 752 5016
rect 824 4940 863 5016
rect 463 4890 863 4940
rect 463 4705 865 4730
rect 463 4629 503 4705
rect 575 4629 629 4705
rect 701 4629 749 4705
rect 821 4629 865 4705
rect 463 4587 865 4629
rect 463 4511 503 4587
rect 575 4511 629 4587
rect 701 4511 749 4587
rect 821 4511 865 4587
rect 463 4475 865 4511
rect 21028 4594 21428 4619
rect 21028 4518 21068 4594
rect 21140 4518 21194 4594
rect 21266 4518 21314 4594
rect 21386 4518 21428 4594
rect 21028 4476 21428 4518
rect 21028 4400 21068 4476
rect 21140 4400 21194 4476
rect 21266 4400 21314 4476
rect 21386 4400 21428 4476
rect 21028 4364 21428 4400
rect 463 3528 863 3553
rect 463 3452 503 3528
rect 575 3452 629 3528
rect 701 3452 749 3528
rect 821 3452 863 3528
rect 463 3410 863 3452
rect 463 3334 503 3410
rect 575 3334 629 3410
rect 701 3334 749 3410
rect 821 3334 863 3410
rect 463 3298 863 3334
rect 21027 3437 21427 3462
rect 21027 3361 21068 3437
rect 21140 3361 21194 3437
rect 21266 3361 21314 3437
rect 21386 3361 21427 3437
rect 21027 3319 21427 3361
rect 21027 3243 21068 3319
rect 21140 3243 21194 3319
rect 21266 3243 21314 3319
rect 21386 3243 21427 3319
rect 21027 3207 21427 3243
rect 463 3061 863 3110
rect 463 2985 504 3061
rect 576 2985 626 3061
rect 698 2985 752 3061
rect 824 2985 863 3061
rect 463 2914 863 2985
rect 463 2838 504 2914
rect 576 2838 626 2914
rect 698 2838 752 2914
rect 824 2838 863 2914
rect 463 2777 863 2838
rect 463 2701 504 2777
rect 576 2701 626 2777
rect 698 2701 752 2777
rect 824 2701 863 2777
rect 463 2651 863 2701
rect 21970 2280 22370 2305
rect 21970 2204 22010 2280
rect 22082 2204 22136 2280
rect 22208 2204 22256 2280
rect 22328 2204 22370 2280
rect 21970 2162 22370 2204
rect 21970 2086 22010 2162
rect 22082 2086 22136 2162
rect 22208 2086 22256 2162
rect 22328 2086 22370 2162
rect 21970 2050 22370 2086
rect 463 1300 863 1349
rect 463 1224 504 1300
rect 576 1224 626 1300
rect 698 1224 752 1300
rect 824 1224 863 1300
rect 463 1153 863 1224
rect 463 1077 504 1153
rect 576 1077 626 1153
rect 698 1077 752 1153
rect 824 1077 863 1153
rect 463 1016 863 1077
rect 463 940 504 1016
rect 576 940 626 1016
rect 698 940 752 1016
rect 824 940 863 1016
rect 463 890 863 940
rect 463 705 865 730
rect 463 629 503 705
rect 575 629 629 705
rect 701 629 749 705
rect 821 629 865 705
rect 463 587 865 629
rect 463 511 503 587
rect 575 511 629 587
rect 701 511 749 587
rect 821 511 865 587
rect 463 475 865 511
rect 21028 594 21428 619
rect 21028 518 21068 594
rect 21140 518 21194 594
rect 21266 518 21314 594
rect 21386 518 21428 594
rect 21028 476 21428 518
rect 21028 400 21068 476
rect 21140 400 21194 476
rect 21266 400 21314 476
rect 21386 400 21428 476
rect 21028 364 21428 400
<< via3 >>
rect 503 75376 575 75452
rect 629 75376 701 75452
rect 749 75376 821 75452
rect 503 75258 575 75334
rect 629 75258 701 75334
rect 749 75258 821 75334
rect 21068 75416 21140 75492
rect 21194 75416 21266 75492
rect 21314 75416 21386 75492
rect 21068 75298 21140 75374
rect 21194 75298 21266 75374
rect 21314 75298 21386 75374
rect 504 74984 576 75060
rect 626 74984 698 75060
rect 752 74984 824 75060
rect 504 74837 576 74913
rect 626 74837 698 74913
rect 752 74837 824 74913
rect 504 74700 576 74776
rect 626 74700 698 74776
rect 752 74700 824 74776
rect 22010 73995 22082 74071
rect 22136 73995 22208 74071
rect 22256 73995 22328 74071
rect 22010 73877 22082 73953
rect 22136 73877 22208 73953
rect 22256 73877 22328 73953
rect 504 73224 576 73300
rect 626 73224 698 73300
rect 752 73224 824 73300
rect 504 73077 576 73153
rect 626 73077 698 73153
rect 752 73077 824 73153
rect 504 72940 576 73016
rect 626 72940 698 73016
rect 752 72940 824 73016
rect 503 72703 575 72779
rect 629 72703 701 72779
rect 749 72703 821 72779
rect 503 72585 575 72661
rect 629 72585 701 72661
rect 749 72585 821 72661
rect 21068 72619 21140 72695
rect 21194 72619 21266 72695
rect 21314 72619 21386 72695
rect 21068 72501 21140 72577
rect 21194 72501 21266 72577
rect 21314 72501 21386 72577
rect 503 71376 575 71452
rect 629 71376 701 71452
rect 749 71376 821 71452
rect 503 71258 575 71334
rect 629 71258 701 71334
rect 749 71258 821 71334
rect 21068 71416 21140 71492
rect 21194 71416 21266 71492
rect 21314 71416 21386 71492
rect 21068 71298 21140 71374
rect 21194 71298 21266 71374
rect 21314 71298 21386 71374
rect 504 70984 576 71060
rect 626 70984 698 71060
rect 752 70984 824 71060
rect 504 70837 576 70913
rect 626 70837 698 70913
rect 752 70837 824 70913
rect 504 70700 576 70776
rect 626 70700 698 70776
rect 752 70700 824 70776
rect 22010 69995 22082 70071
rect 22136 69995 22208 70071
rect 22256 69995 22328 70071
rect 22010 69877 22082 69953
rect 22136 69877 22208 69953
rect 22256 69877 22328 69953
rect 504 69224 576 69300
rect 626 69224 698 69300
rect 752 69224 824 69300
rect 504 69077 576 69153
rect 626 69077 698 69153
rect 752 69077 824 69153
rect 504 68940 576 69016
rect 626 68940 698 69016
rect 752 68940 824 69016
rect 503 68703 575 68779
rect 629 68703 701 68779
rect 749 68703 821 68779
rect 503 68585 575 68661
rect 629 68585 701 68661
rect 749 68585 821 68661
rect 21068 68619 21140 68695
rect 21194 68619 21266 68695
rect 21314 68619 21386 68695
rect 21068 68501 21140 68577
rect 21194 68501 21266 68577
rect 21314 68501 21386 68577
rect 503 67374 575 67450
rect 629 67374 701 67450
rect 749 67374 821 67450
rect 503 67256 575 67332
rect 629 67256 701 67332
rect 749 67256 821 67332
rect 21068 67416 21140 67492
rect 21194 67416 21266 67492
rect 21314 67416 21386 67492
rect 21068 67298 21140 67374
rect 21194 67298 21266 67374
rect 21314 67298 21386 67374
rect 504 66984 576 67060
rect 626 66984 698 67060
rect 752 66984 824 67060
rect 504 66837 576 66913
rect 626 66837 698 66913
rect 752 66837 824 66913
rect 504 66700 576 66776
rect 626 66700 698 66776
rect 752 66700 824 66776
rect 22010 65982 22082 66058
rect 22136 65982 22208 66058
rect 22256 65982 22328 66058
rect 22010 65864 22082 65940
rect 22136 65864 22208 65940
rect 22256 65864 22328 65940
rect 504 65225 576 65301
rect 626 65225 698 65301
rect 752 65225 824 65301
rect 504 65078 576 65154
rect 626 65078 698 65154
rect 752 65078 824 65154
rect 504 64941 576 65017
rect 626 64941 698 65017
rect 752 64941 824 65017
rect 503 64634 575 64710
rect 629 64634 701 64710
rect 749 64634 821 64710
rect 503 64516 575 64592
rect 629 64516 701 64592
rect 749 64516 821 64592
rect 21068 64619 21140 64695
rect 21194 64619 21266 64695
rect 21314 64619 21386 64695
rect 21068 64501 21140 64577
rect 21194 64501 21266 64577
rect 21314 64501 21386 64577
rect 503 63456 575 63532
rect 629 63456 701 63532
rect 749 63456 821 63532
rect 503 63338 575 63414
rect 629 63338 701 63414
rect 749 63338 821 63414
rect 21068 63416 21140 63492
rect 21194 63416 21266 63492
rect 21314 63416 21386 63492
rect 21068 63298 21140 63374
rect 21194 63298 21266 63374
rect 21314 63298 21386 63374
rect 504 62984 576 63060
rect 626 62984 698 63060
rect 752 62984 824 63060
rect 504 62837 576 62913
rect 626 62837 698 62913
rect 752 62837 824 62913
rect 504 62700 576 62776
rect 626 62700 698 62776
rect 752 62700 824 62776
rect 22010 61981 22082 62057
rect 22136 61981 22208 62057
rect 22256 61981 22328 62057
rect 22010 61863 22082 61939
rect 22136 61863 22208 61939
rect 22256 61863 22328 61939
rect 504 61225 576 61301
rect 626 61225 698 61301
rect 752 61225 824 61301
rect 504 61078 576 61154
rect 626 61078 698 61154
rect 752 61078 824 61154
rect 504 60941 576 61017
rect 626 60941 698 61017
rect 752 60941 824 61017
rect 503 60608 575 60684
rect 629 60608 701 60684
rect 749 60608 821 60684
rect 503 60490 575 60566
rect 629 60490 701 60566
rect 749 60490 821 60566
rect 21068 60619 21140 60695
rect 21194 60619 21266 60695
rect 21314 60619 21386 60695
rect 21068 60501 21140 60577
rect 21194 60501 21266 60577
rect 21314 60501 21386 60577
rect 503 59405 575 59481
rect 629 59405 701 59481
rect 749 59405 821 59481
rect 503 59287 575 59363
rect 629 59287 701 59363
rect 749 59287 821 59363
rect 21068 59470 21140 59546
rect 21194 59470 21266 59546
rect 21314 59470 21386 59546
rect 21068 59352 21140 59428
rect 21194 59352 21266 59428
rect 21314 59352 21386 59428
rect 504 58984 576 59060
rect 626 58984 698 59060
rect 752 58984 824 59060
rect 504 58837 576 58913
rect 626 58837 698 58913
rect 752 58837 824 58913
rect 504 58700 576 58776
rect 626 58700 698 58776
rect 752 58700 824 58776
rect 22010 58020 22082 58096
rect 22136 58020 22208 58096
rect 22256 58020 22328 58096
rect 22010 57902 22082 57978
rect 22136 57902 22208 57978
rect 22256 57902 22328 57978
rect 504 57223 576 57299
rect 626 57223 698 57299
rect 752 57223 824 57299
rect 504 57076 576 57152
rect 626 57076 698 57152
rect 752 57076 824 57152
rect 504 56939 576 57015
rect 626 56939 698 57015
rect 752 56939 824 57015
rect 503 56628 575 56704
rect 629 56628 701 56704
rect 749 56628 821 56704
rect 503 56510 575 56586
rect 629 56510 701 56586
rect 749 56510 821 56586
rect 21068 56554 21140 56630
rect 21194 56554 21266 56630
rect 21314 56554 21386 56630
rect 21068 56436 21140 56512
rect 21194 56436 21266 56512
rect 21314 56436 21386 56512
rect 503 55421 575 55497
rect 629 55421 701 55497
rect 749 55421 821 55497
rect 503 55303 575 55379
rect 629 55303 701 55379
rect 749 55303 821 55379
rect 21068 55371 21140 55447
rect 21194 55371 21266 55447
rect 21314 55371 21386 55447
rect 21068 55253 21140 55329
rect 21194 55253 21266 55329
rect 21314 55253 21386 55329
rect 504 54984 576 55060
rect 626 54984 698 55060
rect 752 54984 824 55060
rect 504 54837 576 54913
rect 626 54837 698 54913
rect 752 54837 824 54913
rect 504 54700 576 54776
rect 626 54700 698 54776
rect 752 54700 824 54776
rect 22010 54003 22082 54079
rect 22136 54003 22208 54079
rect 22256 54003 22328 54079
rect 22010 53885 22082 53961
rect 22136 53885 22208 53961
rect 22256 53885 22328 53961
rect 504 53225 576 53301
rect 626 53225 698 53301
rect 752 53225 824 53301
rect 504 53078 576 53154
rect 626 53078 698 53154
rect 752 53078 824 53154
rect 504 52941 576 53017
rect 626 52941 698 53017
rect 752 52941 824 53017
rect 503 52655 575 52731
rect 629 52655 701 52731
rect 749 52655 821 52731
rect 503 52537 575 52613
rect 629 52537 701 52613
rect 749 52537 821 52613
rect 21068 52499 21140 52575
rect 21194 52499 21266 52575
rect 21314 52499 21386 52575
rect 21068 52381 21140 52457
rect 21194 52381 21266 52457
rect 21314 52381 21386 52457
rect 503 51468 575 51544
rect 629 51468 701 51544
rect 749 51468 821 51544
rect 503 51350 575 51426
rect 629 51350 701 51426
rect 749 51350 821 51426
rect 21068 51364 21140 51440
rect 21194 51364 21266 51440
rect 21314 51364 21386 51440
rect 21068 51246 21140 51322
rect 21194 51246 21266 51322
rect 21314 51246 21386 51322
rect 504 50984 576 51060
rect 626 50984 698 51060
rect 752 50984 824 51060
rect 504 50837 576 50913
rect 626 50837 698 50913
rect 752 50837 824 50913
rect 504 50700 576 50776
rect 626 50700 698 50776
rect 752 50700 824 50776
rect 22010 50082 22082 50158
rect 22136 50082 22208 50158
rect 22256 50082 22328 50158
rect 22010 49964 22082 50040
rect 22136 49964 22208 50040
rect 22256 49964 22328 50040
rect 504 49225 576 49301
rect 626 49225 698 49301
rect 752 49225 824 49301
rect 504 49078 576 49154
rect 626 49078 698 49154
rect 752 49078 824 49154
rect 504 48941 576 49017
rect 626 48941 698 49017
rect 752 48941 824 49017
rect 503 48646 575 48722
rect 629 48646 701 48722
rect 749 48646 821 48722
rect 503 48528 575 48604
rect 629 48528 701 48604
rect 749 48528 821 48604
rect 21068 48605 21140 48681
rect 21194 48605 21266 48681
rect 21314 48605 21386 48681
rect 21068 48487 21140 48563
rect 21194 48487 21266 48563
rect 21314 48487 21386 48563
rect 503 47493 575 47569
rect 629 47493 701 47569
rect 749 47493 821 47569
rect 503 47375 575 47451
rect 629 47375 701 47451
rect 749 47375 821 47451
rect 21068 47452 21140 47528
rect 21194 47452 21266 47528
rect 21314 47452 21386 47528
rect 21068 47334 21140 47410
rect 21194 47334 21266 47410
rect 21314 47334 21386 47410
rect 504 46984 576 47060
rect 626 46984 698 47060
rect 752 46984 824 47060
rect 504 46837 576 46913
rect 626 46837 698 46913
rect 752 46837 824 46913
rect 504 46700 576 46776
rect 626 46700 698 46776
rect 752 46700 824 46776
rect 22010 45824 22082 45900
rect 22136 45824 22208 45900
rect 22256 45824 22328 45900
rect 22010 45706 22082 45782
rect 22136 45706 22208 45782
rect 22256 45706 22328 45782
rect 504 45224 576 45300
rect 626 45224 698 45300
rect 752 45224 824 45300
rect 504 45077 576 45153
rect 626 45077 698 45153
rect 752 45077 824 45153
rect 504 44940 576 45016
rect 626 44940 698 45016
rect 752 44940 824 45016
rect 503 44433 575 44509
rect 629 44433 701 44509
rect 749 44433 821 44509
rect 503 44315 575 44391
rect 629 44315 701 44391
rect 749 44315 821 44391
rect 21068 44336 21140 44412
rect 21194 44336 21266 44412
rect 21314 44336 21386 44412
rect 21068 44218 21140 44294
rect 21194 44218 21266 44294
rect 21314 44218 21386 44294
rect 22006 43514 22298 43838
rect 2249 39869 2257 39925
rect 2257 39869 2313 39925
rect 2249 39861 2313 39869
rect 2337 39869 2393 39925
rect 2393 39869 2401 39925
rect 2337 39861 2401 39869
rect 2249 39789 2257 39845
rect 2257 39789 2313 39845
rect 2249 39781 2313 39789
rect 2337 39789 2393 39845
rect 2393 39789 2401 39845
rect 2337 39781 2401 39789
rect 4192 39841 4256 39905
rect 4280 39841 4344 39905
rect 4192 39761 4256 39825
rect 4280 39761 4344 39825
rect 32 39661 111 39741
rect 156 39661 157 39741
rect 157 39661 236 39741
rect 282 39661 362 39741
rect 32 39555 111 39635
rect 156 39555 157 39635
rect 157 39555 236 39635
rect 282 39555 362 39635
rect 21535 39646 21615 39726
rect 21660 39646 21740 39726
rect 21785 39646 21865 39726
rect 21534 39526 21614 39606
rect 21659 39526 21739 39606
rect 21784 39526 21864 39606
rect 478 39130 562 39131
rect 478 39052 479 39130
rect 479 39052 561 39130
rect 561 39052 562 39130
rect 478 39051 562 39052
rect 592 39130 676 39131
rect 592 39052 593 39130
rect 593 39052 675 39130
rect 675 39052 676 39130
rect 592 39051 676 39052
rect 706 39130 790 39131
rect 706 39052 707 39130
rect 707 39052 789 39130
rect 789 39052 790 39130
rect 706 39051 790 39052
rect 15 38586 99 38587
rect 15 38508 16 38586
rect 16 38508 98 38586
rect 98 38508 99 38586
rect 15 38507 99 38508
rect 129 38586 213 38587
rect 129 38508 130 38586
rect 130 38508 212 38586
rect 212 38508 213 38586
rect 129 38507 213 38508
rect 243 38586 327 38587
rect 243 38508 244 38586
rect 244 38508 326 38586
rect 326 38508 327 38586
rect 243 38507 327 38508
rect 478 38042 562 38043
rect 478 37964 479 38042
rect 479 37964 561 38042
rect 561 37964 562 38042
rect 478 37963 562 37964
rect 592 38042 676 38043
rect 592 37964 593 38042
rect 593 37964 675 38042
rect 675 37964 676 38042
rect 592 37963 676 37964
rect 706 38042 790 38043
rect 706 37964 707 38042
rect 707 37964 789 38042
rect 789 37964 790 38042
rect 706 37963 790 37964
rect 15 37498 99 37499
rect 15 37420 16 37498
rect 16 37420 98 37498
rect 98 37420 99 37498
rect 15 37419 99 37420
rect 129 37498 213 37499
rect 129 37420 130 37498
rect 130 37420 212 37498
rect 212 37420 213 37498
rect 129 37419 213 37420
rect 243 37498 327 37499
rect 243 37420 244 37498
rect 244 37420 326 37498
rect 326 37420 327 37498
rect 243 37419 327 37420
rect 478 36954 562 36955
rect 478 36876 479 36954
rect 479 36876 561 36954
rect 561 36876 562 36954
rect 478 36875 562 36876
rect 592 36954 676 36955
rect 592 36876 593 36954
rect 593 36876 675 36954
rect 675 36876 676 36954
rect 592 36875 676 36876
rect 706 36954 790 36955
rect 706 36876 707 36954
rect 707 36876 789 36954
rect 789 36876 790 36954
rect 706 36875 790 36876
rect 22006 36630 22298 36954
rect 2536 36401 2544 36463
rect 2544 36401 2600 36463
rect 2536 36399 2600 36401
rect 2624 36401 2680 36463
rect 2680 36401 2688 36463
rect 2624 36399 2688 36401
rect 21061 36092 21141 36172
rect 21186 36092 21266 36172
rect 21311 36092 21391 36172
rect 21060 35972 21140 36052
rect 21185 35972 21265 36052
rect 21310 35972 21390 36052
rect 21069 35516 21141 35592
rect 21191 35516 21263 35592
rect 21317 35516 21389 35592
rect 21069 35369 21141 35445
rect 21191 35369 21263 35445
rect 21317 35369 21389 35445
rect 21069 35232 21141 35308
rect 21191 35232 21263 35308
rect 21317 35232 21389 35308
rect 20560 34596 20640 34676
rect 20685 34596 20765 34676
rect 20810 34596 20890 34676
rect 20559 34476 20639 34556
rect 20684 34476 20764 34556
rect 20809 34476 20889 34556
rect 21535 34596 21615 34676
rect 21660 34596 21740 34676
rect 21785 34596 21865 34676
rect 21534 34476 21614 34556
rect 21659 34476 21739 34556
rect 21784 34476 21864 34556
rect 21069 33756 21141 33832
rect 21191 33756 21263 33832
rect 21317 33756 21389 33832
rect 21069 33609 21141 33685
rect 21191 33609 21263 33685
rect 21317 33609 21389 33685
rect 21069 33472 21141 33548
rect 21191 33472 21263 33548
rect 21317 33472 21389 33548
rect 21060 33037 21140 33117
rect 21185 33037 21265 33117
rect 21310 33037 21390 33117
rect 21059 32917 21139 32997
rect 21184 32917 21264 32997
rect 21309 32917 21389 32997
rect 503 32226 575 32302
rect 629 32226 701 32302
rect 749 32226 821 32302
rect 503 32108 575 32184
rect 629 32108 701 32184
rect 749 32108 821 32184
rect 21068 32226 21140 32302
rect 21194 32226 21266 32302
rect 21314 32226 21386 32302
rect 21068 32108 21140 32184
rect 21194 32108 21266 32184
rect 21314 32108 21386 32184
rect 503 31444 575 31520
rect 629 31444 701 31520
rect 749 31444 821 31520
rect 503 31326 575 31402
rect 629 31326 701 31402
rect 749 31326 821 31402
rect 21068 31444 21140 31520
rect 21194 31444 21266 31520
rect 21314 31444 21386 31520
rect 21068 31326 21140 31402
rect 21194 31326 21266 31402
rect 21314 31326 21386 31402
rect 504 30985 576 31061
rect 626 30985 698 31061
rect 752 30985 824 31061
rect 504 30838 576 30914
rect 626 30838 698 30914
rect 752 30838 824 30914
rect 504 30701 576 30777
rect 626 30701 698 30777
rect 752 30701 824 30777
rect 22010 30054 22082 30130
rect 22136 30054 22208 30130
rect 22256 30054 22328 30130
rect 22010 29936 22082 30012
rect 22136 29936 22208 30012
rect 22256 29936 22328 30012
rect 504 29218 576 29294
rect 626 29218 698 29294
rect 752 29218 824 29294
rect 504 29071 576 29147
rect 626 29071 698 29147
rect 752 29071 824 29147
rect 504 28934 576 29010
rect 626 28934 698 29010
rect 752 28934 824 29010
rect 503 28532 575 28608
rect 629 28532 701 28608
rect 749 28532 821 28608
rect 503 28414 575 28490
rect 629 28414 701 28490
rect 749 28414 821 28490
rect 21068 28483 21140 28559
rect 21194 28483 21266 28559
rect 21314 28483 21386 28559
rect 21068 28365 21140 28441
rect 21194 28365 21266 28441
rect 21314 28365 21386 28441
rect 503 27528 575 27604
rect 629 27528 701 27604
rect 749 27528 821 27604
rect 503 27410 575 27486
rect 629 27410 701 27486
rect 749 27410 821 27486
rect 21068 27366 21140 27442
rect 21194 27366 21266 27442
rect 21314 27366 21386 27442
rect 21068 27248 21140 27324
rect 21194 27248 21266 27324
rect 21314 27248 21386 27324
rect 504 26984 576 27060
rect 626 26984 698 27060
rect 752 26984 824 27060
rect 504 26837 576 26913
rect 626 26837 698 26913
rect 752 26837 824 26913
rect 504 26700 576 26776
rect 626 26700 698 26776
rect 752 26700 824 26776
rect 22010 25895 22082 25971
rect 22136 25895 22208 25971
rect 22256 25895 22328 25971
rect 22010 25777 22082 25853
rect 22136 25777 22208 25853
rect 22256 25777 22328 25853
rect 504 25224 576 25300
rect 626 25224 698 25300
rect 752 25224 824 25300
rect 504 25077 576 25153
rect 626 25077 698 25153
rect 752 25077 824 25153
rect 504 24940 576 25016
rect 626 24940 698 25016
rect 752 24940 824 25016
rect 503 24550 575 24626
rect 629 24550 701 24626
rect 749 24550 821 24626
rect 503 24432 575 24508
rect 629 24432 701 24508
rect 749 24432 821 24508
rect 21068 24523 21140 24599
rect 21194 24523 21266 24599
rect 21314 24523 21386 24599
rect 21068 24405 21140 24481
rect 21194 24405 21266 24481
rect 21314 24405 21386 24481
rect 503 23468 575 23544
rect 629 23468 701 23544
rect 749 23468 821 23544
rect 503 23350 575 23426
rect 629 23350 701 23426
rect 749 23350 821 23426
rect 21068 23348 21140 23424
rect 21194 23348 21266 23424
rect 21314 23348 21386 23424
rect 21068 23230 21140 23306
rect 21194 23230 21266 23306
rect 21314 23230 21386 23306
rect 504 22984 576 23060
rect 626 22984 698 23060
rect 752 22984 824 23060
rect 504 22837 576 22913
rect 626 22837 698 22913
rect 752 22837 824 22913
rect 504 22700 576 22776
rect 626 22700 698 22776
rect 752 22700 824 22776
rect 22010 22105 22082 22181
rect 22136 22105 22208 22181
rect 22256 22105 22328 22181
rect 22010 21987 22082 22063
rect 22136 21987 22208 22063
rect 22256 21987 22328 22063
rect 504 21225 576 21301
rect 626 21225 698 21301
rect 752 21225 824 21301
rect 504 21078 576 21154
rect 626 21078 698 21154
rect 752 21078 824 21154
rect 504 20941 576 21017
rect 626 20941 698 21017
rect 752 20941 824 21017
rect 503 20593 575 20669
rect 629 20593 701 20669
rect 749 20593 821 20669
rect 503 20475 575 20551
rect 629 20475 701 20551
rect 749 20475 821 20551
rect 21068 20507 21140 20583
rect 21194 20507 21266 20583
rect 21314 20507 21386 20583
rect 21068 20389 21140 20465
rect 21194 20389 21266 20465
rect 21314 20389 21386 20465
rect 503 19492 575 19568
rect 629 19492 701 19568
rect 749 19492 821 19568
rect 503 19374 575 19450
rect 629 19374 701 19450
rect 749 19374 821 19450
rect 21068 19336 21140 19412
rect 21194 19336 21266 19412
rect 21314 19336 21386 19412
rect 21068 19218 21140 19294
rect 21194 19218 21266 19294
rect 21314 19218 21386 19294
rect 504 18984 576 19060
rect 626 18984 698 19060
rect 752 18984 824 19060
rect 504 18837 576 18913
rect 626 18837 698 18913
rect 752 18837 824 18913
rect 504 18700 576 18776
rect 626 18700 698 18776
rect 752 18700 824 18776
rect 22010 17998 22082 18074
rect 22136 17998 22208 18074
rect 22256 17998 22328 18074
rect 22010 17880 22082 17956
rect 22136 17880 22208 17956
rect 22256 17880 22328 17956
rect 504 17224 576 17300
rect 626 17224 698 17300
rect 752 17224 824 17300
rect 504 17077 576 17153
rect 626 17077 698 17153
rect 752 17077 824 17153
rect 504 16940 576 17016
rect 626 16940 698 17016
rect 752 16940 824 17016
rect 503 16626 575 16702
rect 629 16626 701 16702
rect 749 16626 821 16702
rect 503 16508 575 16584
rect 629 16508 701 16584
rect 749 16508 821 16584
rect 21068 16575 21140 16651
rect 21194 16575 21266 16651
rect 21314 16575 21386 16651
rect 21068 16457 21140 16533
rect 21194 16457 21266 16533
rect 21314 16457 21386 16533
rect 503 15410 575 15486
rect 629 15410 701 15486
rect 749 15410 821 15486
rect 503 15292 575 15368
rect 629 15292 701 15368
rect 749 15292 821 15368
rect 21068 15361 21140 15437
rect 21194 15361 21266 15437
rect 21314 15361 21386 15437
rect 21068 15243 21140 15319
rect 21194 15243 21266 15319
rect 21314 15243 21386 15319
rect 504 14984 576 15060
rect 626 14984 698 15060
rect 752 14984 824 15060
rect 504 14837 576 14913
rect 626 14837 698 14913
rect 752 14837 824 14913
rect 504 14700 576 14776
rect 626 14700 698 14776
rect 752 14700 824 14776
rect 22010 14180 22082 14256
rect 22136 14180 22208 14256
rect 22256 14180 22328 14256
rect 22010 14062 22082 14138
rect 22136 14062 22208 14138
rect 22256 14062 22328 14138
rect 504 13224 576 13300
rect 626 13224 698 13300
rect 752 13224 824 13300
rect 504 13077 576 13153
rect 626 13077 698 13153
rect 752 13077 824 13153
rect 504 12940 576 13016
rect 626 12940 698 13016
rect 752 12940 824 13016
rect 503 12545 575 12621
rect 629 12545 701 12621
rect 749 12545 821 12621
rect 503 12427 575 12503
rect 629 12427 701 12503
rect 749 12427 821 12503
rect 21068 12518 21140 12594
rect 21194 12518 21266 12594
rect 21314 12518 21386 12594
rect 21068 12400 21140 12476
rect 21194 12400 21266 12476
rect 21314 12400 21386 12476
rect 503 11423 575 11499
rect 629 11423 701 11499
rect 749 11423 821 11499
rect 503 11305 575 11381
rect 629 11305 701 11381
rect 749 11305 821 11381
rect 21068 11361 21140 11437
rect 21194 11361 21266 11437
rect 21314 11361 21386 11437
rect 21068 11243 21140 11319
rect 21194 11243 21266 11319
rect 21314 11243 21386 11319
rect 504 10985 576 11061
rect 626 10985 698 11061
rect 752 10985 824 11061
rect 504 10838 576 10914
rect 626 10838 698 10914
rect 752 10838 824 10914
rect 504 10701 576 10777
rect 626 10701 698 10777
rect 752 10701 824 10777
rect 22010 10216 22082 10292
rect 22136 10216 22208 10292
rect 22256 10216 22328 10292
rect 22010 10098 22082 10174
rect 22136 10098 22208 10174
rect 22256 10098 22328 10174
rect 504 9223 576 9299
rect 626 9223 698 9299
rect 752 9223 824 9299
rect 504 9076 576 9152
rect 626 9076 698 9152
rect 752 9076 824 9152
rect 504 8939 576 9015
rect 626 8939 698 9015
rect 752 8939 824 9015
rect 503 8563 575 8639
rect 629 8563 701 8639
rect 749 8563 821 8639
rect 503 8445 575 8521
rect 629 8445 701 8521
rect 749 8445 821 8521
rect 21068 8518 21140 8594
rect 21194 8518 21266 8594
rect 21314 8518 21386 8594
rect 21068 8400 21140 8476
rect 21194 8400 21266 8476
rect 21314 8400 21386 8476
rect 503 7452 575 7528
rect 629 7452 701 7528
rect 749 7452 821 7528
rect 503 7334 575 7410
rect 629 7334 701 7410
rect 749 7334 821 7410
rect 21068 7361 21140 7437
rect 21194 7361 21266 7437
rect 21314 7361 21386 7437
rect 21068 7243 21140 7319
rect 21194 7243 21266 7319
rect 21314 7243 21386 7319
rect 504 6985 576 7061
rect 626 6985 698 7061
rect 752 6985 824 7061
rect 504 6838 576 6914
rect 626 6838 698 6914
rect 752 6838 824 6914
rect 504 6701 576 6777
rect 626 6701 698 6777
rect 752 6701 824 6777
rect 22010 6204 22082 6280
rect 22136 6204 22208 6280
rect 22256 6204 22328 6280
rect 22010 6086 22082 6162
rect 22136 6086 22208 6162
rect 22256 6086 22328 6162
rect 504 5224 576 5300
rect 626 5224 698 5300
rect 752 5224 824 5300
rect 504 5077 576 5153
rect 626 5077 698 5153
rect 752 5077 824 5153
rect 504 4940 576 5016
rect 626 4940 698 5016
rect 752 4940 824 5016
rect 503 4629 575 4705
rect 629 4629 701 4705
rect 749 4629 821 4705
rect 503 4511 575 4587
rect 629 4511 701 4587
rect 749 4511 821 4587
rect 21068 4518 21140 4594
rect 21194 4518 21266 4594
rect 21314 4518 21386 4594
rect 21068 4400 21140 4476
rect 21194 4400 21266 4476
rect 21314 4400 21386 4476
rect 503 3452 575 3528
rect 629 3452 701 3528
rect 749 3452 821 3528
rect 503 3334 575 3410
rect 629 3334 701 3410
rect 749 3334 821 3410
rect 21068 3361 21140 3437
rect 21194 3361 21266 3437
rect 21314 3361 21386 3437
rect 21068 3243 21140 3319
rect 21194 3243 21266 3319
rect 21314 3243 21386 3319
rect 504 2985 576 3061
rect 626 2985 698 3061
rect 752 2985 824 3061
rect 504 2838 576 2914
rect 626 2838 698 2914
rect 752 2838 824 2914
rect 504 2701 576 2777
rect 626 2701 698 2777
rect 752 2701 824 2777
rect 22010 2204 22082 2280
rect 22136 2204 22208 2280
rect 22256 2204 22328 2280
rect 22010 2086 22082 2162
rect 22136 2086 22208 2162
rect 22256 2086 22328 2162
rect 504 1224 576 1300
rect 626 1224 698 1300
rect 752 1224 824 1300
rect 504 1077 576 1153
rect 626 1077 698 1153
rect 752 1077 824 1153
rect 504 940 576 1016
rect 626 940 698 1016
rect 752 940 824 1016
rect 503 629 575 705
rect 629 629 701 705
rect 749 629 821 705
rect 503 511 575 587
rect 629 511 701 587
rect 749 511 821 587
rect 21068 518 21140 594
rect 21194 518 21266 594
rect 21314 518 21386 594
rect 21068 400 21140 476
rect 21194 400 21266 476
rect 21314 400 21386 476
<< metal4 >>
rect 0 39741 400 76000
rect 0 39661 32 39741
rect 111 39661 156 39741
rect 236 39661 282 39741
rect 362 39661 400 39741
rect 0 39635 400 39661
rect 0 39555 32 39635
rect 111 39555 156 39635
rect 236 39555 282 39635
rect 362 39555 400 39635
rect 0 38587 400 39555
rect 0 38507 15 38587
rect 99 38507 129 38587
rect 213 38507 243 38587
rect 327 38507 400 38587
rect 0 37499 400 38507
rect 0 37419 15 37499
rect 99 37419 129 37499
rect 213 37419 243 37499
rect 327 37419 400 37499
rect 0 0 400 37419
rect 463 75477 863 76000
rect 21028 75517 21428 76000
rect 21026 75492 21428 75517
rect 463 75452 864 75477
rect 463 75376 503 75452
rect 575 75376 629 75452
rect 701 75376 749 75452
rect 821 75376 864 75452
rect 463 75334 864 75376
rect 463 75258 503 75334
rect 575 75258 629 75334
rect 701 75258 749 75334
rect 821 75258 864 75334
rect 21026 75416 21068 75492
rect 21140 75416 21194 75492
rect 21266 75416 21314 75492
rect 21386 75416 21428 75492
rect 21026 75374 21428 75416
rect 21026 75298 21068 75374
rect 21140 75298 21194 75374
rect 21266 75298 21314 75374
rect 21386 75298 21428 75374
rect 21026 75262 21428 75298
rect 463 75222 864 75258
rect 463 75060 863 75222
rect 463 74984 504 75060
rect 576 74984 626 75060
rect 698 74984 752 75060
rect 824 74984 863 75060
rect 463 74913 863 74984
rect 463 74837 504 74913
rect 576 74837 626 74913
rect 698 74837 752 74913
rect 824 74837 863 74913
rect 463 74776 863 74837
rect 463 74700 504 74776
rect 576 74700 626 74776
rect 698 74700 752 74776
rect 824 74700 863 74776
rect 463 73300 863 74700
rect 463 73224 504 73300
rect 576 73224 626 73300
rect 698 73224 752 73300
rect 824 73224 863 73300
rect 463 73153 863 73224
rect 463 73077 504 73153
rect 576 73077 626 73153
rect 698 73077 752 73153
rect 824 73077 863 73153
rect 463 73016 863 73077
rect 463 72940 504 73016
rect 576 72940 626 73016
rect 698 72940 752 73016
rect 824 72940 863 73016
rect 463 72804 863 72940
rect 463 72779 864 72804
rect 463 72703 503 72779
rect 575 72703 629 72779
rect 701 72703 749 72779
rect 821 72703 864 72779
rect 463 72661 864 72703
rect 463 72585 503 72661
rect 575 72585 629 72661
rect 701 72585 749 72661
rect 821 72585 864 72661
rect 463 72549 864 72585
rect 21028 72695 21428 75262
rect 21028 72619 21068 72695
rect 21140 72619 21194 72695
rect 21266 72619 21314 72695
rect 21386 72619 21428 72695
rect 21028 72577 21428 72619
rect 463 71477 863 72549
rect 21028 72501 21068 72577
rect 21140 72501 21194 72577
rect 21266 72501 21314 72577
rect 21386 72501 21428 72577
rect 21028 71517 21428 72501
rect 21026 71492 21428 71517
rect 463 71452 864 71477
rect 463 71376 503 71452
rect 575 71376 629 71452
rect 701 71376 749 71452
rect 821 71376 864 71452
rect 463 71334 864 71376
rect 463 71258 503 71334
rect 575 71258 629 71334
rect 701 71258 749 71334
rect 821 71258 864 71334
rect 21026 71416 21068 71492
rect 21140 71416 21194 71492
rect 21266 71416 21314 71492
rect 21386 71416 21428 71492
rect 21026 71374 21428 71416
rect 21026 71298 21068 71374
rect 21140 71298 21194 71374
rect 21266 71298 21314 71374
rect 21386 71298 21428 71374
rect 21026 71262 21428 71298
rect 463 71222 864 71258
rect 463 71060 863 71222
rect 463 70984 504 71060
rect 576 70984 626 71060
rect 698 70984 752 71060
rect 824 70984 863 71060
rect 463 70913 863 70984
rect 463 70837 504 70913
rect 576 70837 626 70913
rect 698 70837 752 70913
rect 824 70837 863 70913
rect 463 70776 863 70837
rect 463 70700 504 70776
rect 576 70700 626 70776
rect 698 70700 752 70776
rect 824 70700 863 70776
rect 463 69300 863 70700
rect 463 69224 504 69300
rect 576 69224 626 69300
rect 698 69224 752 69300
rect 824 69224 863 69300
rect 463 69153 863 69224
rect 463 69077 504 69153
rect 576 69077 626 69153
rect 698 69077 752 69153
rect 824 69077 863 69153
rect 463 69016 863 69077
rect 463 68940 504 69016
rect 576 68940 626 69016
rect 698 68940 752 69016
rect 824 68940 863 69016
rect 463 68804 863 68940
rect 463 68779 864 68804
rect 463 68703 503 68779
rect 575 68703 629 68779
rect 701 68703 749 68779
rect 821 68703 864 68779
rect 463 68661 864 68703
rect 463 68585 503 68661
rect 575 68585 629 68661
rect 701 68585 749 68661
rect 821 68585 864 68661
rect 463 68549 864 68585
rect 21028 68695 21428 71262
rect 21028 68619 21068 68695
rect 21140 68619 21194 68695
rect 21266 68619 21314 68695
rect 21386 68619 21428 68695
rect 21028 68577 21428 68619
rect 463 67475 863 68549
rect 21028 68501 21068 68577
rect 21140 68501 21194 68577
rect 21266 68501 21314 68577
rect 21386 68501 21428 68577
rect 21028 67517 21428 68501
rect 21026 67492 21428 67517
rect 463 67450 864 67475
rect 463 67374 503 67450
rect 575 67374 629 67450
rect 701 67374 749 67450
rect 821 67374 864 67450
rect 463 67332 864 67374
rect 463 67256 503 67332
rect 575 67256 629 67332
rect 701 67256 749 67332
rect 821 67256 864 67332
rect 21026 67416 21068 67492
rect 21140 67416 21194 67492
rect 21266 67416 21314 67492
rect 21386 67416 21428 67492
rect 21026 67374 21428 67416
rect 21026 67298 21068 67374
rect 21140 67298 21194 67374
rect 21266 67298 21314 67374
rect 21386 67298 21428 67374
rect 21026 67262 21428 67298
rect 463 67220 864 67256
rect 463 67060 863 67220
rect 463 66984 504 67060
rect 576 66984 626 67060
rect 698 66984 752 67060
rect 824 66984 863 67060
rect 463 66913 863 66984
rect 463 66837 504 66913
rect 576 66837 626 66913
rect 698 66837 752 66913
rect 824 66837 863 66913
rect 463 66776 863 66837
rect 463 66700 504 66776
rect 576 66700 626 66776
rect 698 66700 752 66776
rect 824 66700 863 66776
rect 463 65301 863 66700
rect 463 65225 504 65301
rect 576 65225 626 65301
rect 698 65225 752 65301
rect 824 65225 863 65301
rect 463 65154 863 65225
rect 463 65078 504 65154
rect 576 65078 626 65154
rect 698 65078 752 65154
rect 824 65078 863 65154
rect 463 65017 863 65078
rect 463 64941 504 65017
rect 576 64941 626 65017
rect 698 64941 752 65017
rect 824 64941 863 65017
rect 463 64735 863 64941
rect 463 64710 864 64735
rect 463 64634 503 64710
rect 575 64634 629 64710
rect 701 64634 749 64710
rect 821 64634 864 64710
rect 463 64592 864 64634
rect 463 64516 503 64592
rect 575 64516 629 64592
rect 701 64516 749 64592
rect 821 64516 864 64592
rect 463 64480 864 64516
rect 21028 64695 21428 67262
rect 21028 64619 21068 64695
rect 21140 64619 21194 64695
rect 21266 64619 21314 64695
rect 21386 64619 21428 64695
rect 21028 64577 21428 64619
rect 21028 64501 21068 64577
rect 21140 64501 21194 64577
rect 21266 64501 21314 64577
rect 21386 64501 21428 64577
rect 463 63557 863 64480
rect 463 63532 864 63557
rect 463 63456 503 63532
rect 575 63456 629 63532
rect 701 63456 749 63532
rect 821 63456 864 63532
rect 21028 63517 21428 64501
rect 463 63414 864 63456
rect 463 63338 503 63414
rect 575 63338 629 63414
rect 701 63338 749 63414
rect 821 63338 864 63414
rect 463 63302 864 63338
rect 21026 63492 21428 63517
rect 21026 63416 21068 63492
rect 21140 63416 21194 63492
rect 21266 63416 21314 63492
rect 21386 63416 21428 63492
rect 21026 63374 21428 63416
rect 463 63109 863 63302
rect 21026 63298 21068 63374
rect 21140 63298 21194 63374
rect 21266 63298 21314 63374
rect 21386 63298 21428 63374
rect 21026 63262 21428 63298
rect 463 63060 864 63109
rect 463 62984 504 63060
rect 576 62984 626 63060
rect 698 62984 752 63060
rect 824 62984 864 63060
rect 463 62913 864 62984
rect 463 62837 504 62913
rect 576 62837 626 62913
rect 698 62837 752 62913
rect 824 62837 864 62913
rect 463 62776 864 62837
rect 463 62700 504 62776
rect 576 62700 626 62776
rect 698 62700 752 62776
rect 824 62700 864 62776
rect 463 62650 864 62700
rect 463 61301 863 62650
rect 463 61225 504 61301
rect 576 61225 626 61301
rect 698 61225 752 61301
rect 824 61225 863 61301
rect 463 61154 863 61225
rect 463 61078 504 61154
rect 576 61078 626 61154
rect 698 61078 752 61154
rect 824 61078 863 61154
rect 463 61017 863 61078
rect 463 60941 504 61017
rect 576 60941 626 61017
rect 698 60941 752 61017
rect 824 60941 863 61017
rect 463 60709 863 60941
rect 463 60684 866 60709
rect 463 60608 503 60684
rect 575 60608 629 60684
rect 701 60608 749 60684
rect 821 60608 866 60684
rect 463 60566 866 60608
rect 463 60490 503 60566
rect 575 60490 629 60566
rect 701 60490 749 60566
rect 821 60490 866 60566
rect 463 60454 866 60490
rect 21028 60695 21428 63262
rect 21028 60619 21068 60695
rect 21140 60619 21194 60695
rect 21266 60619 21314 60695
rect 21386 60619 21428 60695
rect 21028 60577 21428 60619
rect 21028 60501 21068 60577
rect 21140 60501 21194 60577
rect 21266 60501 21314 60577
rect 21386 60501 21428 60577
rect 463 59506 863 60454
rect 21028 59571 21428 60501
rect 21027 59546 21428 59571
rect 463 59481 864 59506
rect 463 59405 503 59481
rect 575 59405 629 59481
rect 701 59405 749 59481
rect 821 59405 864 59481
rect 463 59363 864 59405
rect 463 59287 503 59363
rect 575 59287 629 59363
rect 701 59287 749 59363
rect 821 59287 864 59363
rect 21027 59470 21068 59546
rect 21140 59470 21194 59546
rect 21266 59470 21314 59546
rect 21386 59470 21428 59546
rect 21027 59428 21428 59470
rect 21027 59352 21068 59428
rect 21140 59352 21194 59428
rect 21266 59352 21314 59428
rect 21386 59352 21428 59428
rect 21027 59316 21428 59352
rect 463 59251 864 59287
rect 463 59109 863 59251
rect 463 59060 864 59109
rect 463 58984 504 59060
rect 576 58984 626 59060
rect 698 58984 752 59060
rect 824 58984 864 59060
rect 463 58913 864 58984
rect 463 58837 504 58913
rect 576 58837 626 58913
rect 698 58837 752 58913
rect 824 58837 864 58913
rect 463 58776 864 58837
rect 463 58700 504 58776
rect 576 58700 626 58776
rect 698 58700 752 58776
rect 824 58700 864 58776
rect 463 58650 864 58700
rect 463 57299 863 58650
rect 463 57223 504 57299
rect 576 57223 626 57299
rect 698 57223 752 57299
rect 824 57223 863 57299
rect 463 57152 863 57223
rect 463 57076 504 57152
rect 576 57076 626 57152
rect 698 57076 752 57152
rect 824 57076 863 57152
rect 463 57015 863 57076
rect 463 56939 504 57015
rect 576 56939 626 57015
rect 698 56939 752 57015
rect 824 56939 863 57015
rect 463 56729 863 56939
rect 463 56704 864 56729
rect 463 56628 503 56704
rect 575 56628 629 56704
rect 701 56628 749 56704
rect 821 56628 864 56704
rect 463 56586 864 56628
rect 463 56510 503 56586
rect 575 56510 629 56586
rect 701 56510 749 56586
rect 821 56510 864 56586
rect 463 56474 864 56510
rect 21028 56630 21428 59316
rect 21028 56554 21068 56630
rect 21140 56554 21194 56630
rect 21266 56554 21314 56630
rect 21386 56554 21428 56630
rect 21028 56512 21428 56554
rect 463 55522 863 56474
rect 21028 56436 21068 56512
rect 21140 56436 21194 56512
rect 21266 56436 21314 56512
rect 21386 56436 21428 56512
rect 463 55497 866 55522
rect 463 55421 503 55497
rect 575 55421 629 55497
rect 701 55421 749 55497
rect 821 55421 866 55497
rect 21028 55472 21428 56436
rect 463 55379 866 55421
rect 463 55303 503 55379
rect 575 55303 629 55379
rect 701 55303 749 55379
rect 821 55303 866 55379
rect 463 55267 866 55303
rect 21027 55447 21428 55472
rect 21027 55371 21068 55447
rect 21140 55371 21194 55447
rect 21266 55371 21314 55447
rect 21386 55371 21428 55447
rect 21027 55329 21428 55371
rect 463 55060 863 55267
rect 21027 55253 21068 55329
rect 21140 55253 21194 55329
rect 21266 55253 21314 55329
rect 21386 55253 21428 55329
rect 21027 55217 21428 55253
rect 463 54984 504 55060
rect 576 54984 626 55060
rect 698 54984 752 55060
rect 824 54984 863 55060
rect 463 54913 863 54984
rect 463 54837 504 54913
rect 576 54837 626 54913
rect 698 54837 752 54913
rect 824 54837 863 54913
rect 463 54776 863 54837
rect 463 54700 504 54776
rect 576 54700 626 54776
rect 698 54700 752 54776
rect 824 54700 863 54776
rect 463 53301 863 54700
rect 463 53225 504 53301
rect 576 53225 626 53301
rect 698 53225 752 53301
rect 824 53225 863 53301
rect 463 53154 863 53225
rect 463 53078 504 53154
rect 576 53078 626 53154
rect 698 53078 752 53154
rect 824 53078 863 53154
rect 463 53017 863 53078
rect 463 52941 504 53017
rect 576 52941 626 53017
rect 698 52941 752 53017
rect 824 52941 863 53017
rect 463 52756 863 52941
rect 463 52731 864 52756
rect 463 52655 503 52731
rect 575 52655 629 52731
rect 701 52655 749 52731
rect 821 52655 864 52731
rect 463 52613 864 52655
rect 463 52537 503 52613
rect 575 52537 629 52613
rect 701 52537 749 52613
rect 821 52537 864 52613
rect 463 52501 864 52537
rect 21028 52575 21428 55217
rect 463 51569 863 52501
rect 21028 52499 21068 52575
rect 21140 52499 21194 52575
rect 21266 52499 21314 52575
rect 21386 52499 21428 52575
rect 21028 52457 21428 52499
rect 21028 52381 21068 52457
rect 21140 52381 21194 52457
rect 21266 52381 21314 52457
rect 21386 52381 21428 52457
rect 463 51544 864 51569
rect 463 51468 503 51544
rect 575 51468 629 51544
rect 701 51468 749 51544
rect 821 51468 864 51544
rect 463 51426 864 51468
rect 463 51350 503 51426
rect 575 51350 629 51426
rect 701 51350 749 51426
rect 821 51350 864 51426
rect 463 51314 864 51350
rect 21028 51440 21428 52381
rect 21028 51364 21068 51440
rect 21140 51364 21194 51440
rect 21266 51364 21314 51440
rect 21386 51364 21428 51440
rect 21028 51322 21428 51364
rect 463 51060 863 51314
rect 463 50984 504 51060
rect 576 50984 626 51060
rect 698 50984 752 51060
rect 824 50984 863 51060
rect 463 50913 863 50984
rect 463 50837 504 50913
rect 576 50837 626 50913
rect 698 50837 752 50913
rect 824 50837 863 50913
rect 463 50776 863 50837
rect 463 50700 504 50776
rect 576 50700 626 50776
rect 698 50700 752 50776
rect 824 50700 863 50776
rect 463 49301 863 50700
rect 463 49225 504 49301
rect 576 49225 626 49301
rect 698 49225 752 49301
rect 824 49225 863 49301
rect 463 49154 863 49225
rect 463 49078 504 49154
rect 576 49078 626 49154
rect 698 49078 752 49154
rect 824 49078 863 49154
rect 463 49017 863 49078
rect 463 48941 504 49017
rect 576 48941 626 49017
rect 698 48941 752 49017
rect 824 48941 863 49017
rect 463 48747 863 48941
rect 21028 51246 21068 51322
rect 21140 51246 21194 51322
rect 21266 51246 21314 51322
rect 21386 51246 21428 51322
rect 463 48722 864 48747
rect 463 48646 503 48722
rect 575 48646 629 48722
rect 701 48646 749 48722
rect 821 48646 864 48722
rect 463 48604 864 48646
rect 463 48528 503 48604
rect 575 48528 629 48604
rect 701 48528 749 48604
rect 821 48528 864 48604
rect 463 48492 864 48528
rect 21028 48681 21428 51246
rect 21028 48605 21068 48681
rect 21140 48605 21194 48681
rect 21266 48605 21314 48681
rect 21386 48605 21428 48681
rect 21028 48563 21428 48605
rect 463 47594 863 48492
rect 21028 48487 21068 48563
rect 21140 48487 21194 48563
rect 21266 48487 21314 48563
rect 21386 48487 21428 48563
rect 463 47569 864 47594
rect 463 47493 503 47569
rect 575 47493 629 47569
rect 701 47493 749 47569
rect 821 47493 864 47569
rect 463 47451 864 47493
rect 463 47375 503 47451
rect 575 47375 629 47451
rect 701 47375 749 47451
rect 821 47375 864 47451
rect 463 47339 864 47375
rect 21028 47528 21428 48487
rect 21028 47452 21068 47528
rect 21140 47452 21194 47528
rect 21266 47452 21314 47528
rect 21386 47452 21428 47528
rect 21028 47410 21428 47452
rect 463 47060 863 47339
rect 463 46984 504 47060
rect 576 46984 626 47060
rect 698 46984 752 47060
rect 824 46984 863 47060
rect 463 46913 863 46984
rect 463 46837 504 46913
rect 576 46837 626 46913
rect 698 46837 752 46913
rect 824 46837 863 46913
rect 463 46776 863 46837
rect 463 46700 504 46776
rect 576 46700 626 46776
rect 698 46700 752 46776
rect 824 46700 863 46776
rect 463 45300 863 46700
rect 463 45224 504 45300
rect 576 45224 626 45300
rect 698 45224 752 45300
rect 824 45224 863 45300
rect 463 45153 863 45224
rect 463 45077 504 45153
rect 576 45077 626 45153
rect 698 45077 752 45153
rect 824 45077 863 45153
rect 463 45016 863 45077
rect 463 44940 504 45016
rect 576 44940 626 45016
rect 698 44940 752 45016
rect 824 44940 863 45016
rect 463 44509 863 44940
rect 463 44433 503 44509
rect 575 44433 629 44509
rect 701 44433 749 44509
rect 821 44433 863 44509
rect 463 44391 863 44433
rect 463 44315 503 44391
rect 575 44315 629 44391
rect 701 44315 749 44391
rect 821 44315 863 44391
rect 463 39131 863 44315
rect 21028 47334 21068 47410
rect 21140 47334 21194 47410
rect 21266 47334 21314 47410
rect 21386 47334 21428 47410
rect 21028 44412 21428 47334
rect 21028 44336 21068 44412
rect 21140 44336 21194 44412
rect 21266 44336 21314 44412
rect 21386 44336 21428 44412
rect 21028 44294 21428 44336
rect 21028 44218 21068 44294
rect 21140 44218 21194 44294
rect 21266 44218 21314 44294
rect 21386 44218 21428 44294
rect 2306 39942 2868 44002
rect 2246 39925 2868 39942
rect 2246 39861 2249 39925
rect 2313 39861 2337 39925
rect 2401 39861 2868 39925
rect 2246 39845 2868 39861
rect 2246 39781 2249 39845
rect 2313 39781 2337 39845
rect 2401 39781 2868 39845
rect 2246 39775 2868 39781
rect 2306 39774 2868 39775
rect 4119 39905 4490 44000
rect 4119 39841 4192 39905
rect 4256 39841 4280 39905
rect 4344 39841 4490 39905
rect 4119 39825 4490 39841
rect 4119 39761 4192 39825
rect 4256 39761 4280 39825
rect 4344 39761 4490 39825
rect 4119 39754 4490 39761
rect 463 39051 478 39131
rect 562 39051 592 39131
rect 676 39051 706 39131
rect 790 39051 863 39131
rect 463 38043 863 39051
rect 463 37963 478 38043
rect 562 37963 592 38043
rect 676 37963 706 38043
rect 790 37963 863 38043
rect 463 36955 863 37963
rect 463 36875 478 36955
rect 562 36875 592 36955
rect 676 36875 706 36955
rect 790 36875 863 36955
rect 463 32360 863 36875
rect 2306 36463 2738 36476
rect 2306 36399 2536 36463
rect 2600 36399 2624 36463
rect 2688 36399 2738 36463
rect 463 32302 866 32360
rect 463 32226 503 32302
rect 575 32226 629 32302
rect 701 32226 749 32302
rect 821 32226 866 32302
rect 463 32184 866 32226
rect 463 32108 503 32184
rect 575 32108 629 32184
rect 701 32108 749 32184
rect 821 32108 866 32184
rect 463 32072 866 32108
rect 463 32000 863 32072
rect 2306 32000 2738 36399
rect 21028 36198 21428 44218
rect 20527 36172 21428 36198
rect 20527 36092 21061 36172
rect 21141 36092 21186 36172
rect 21266 36092 21311 36172
rect 21391 36092 21428 36172
rect 20527 36052 21428 36092
rect 20527 35972 21060 36052
rect 21140 35972 21185 36052
rect 21265 35972 21310 36052
rect 21390 35972 21428 36052
rect 20527 35943 21428 35972
rect 21028 35592 21428 35943
rect 21028 35516 21069 35592
rect 21141 35516 21191 35592
rect 21263 35516 21317 35592
rect 21389 35516 21428 35592
rect 21028 35445 21428 35516
rect 21028 35369 21069 35445
rect 21141 35369 21191 35445
rect 21263 35369 21317 35445
rect 21389 35369 21428 35445
rect 21028 35308 21428 35369
rect 21028 35232 21069 35308
rect 21141 35232 21191 35308
rect 21263 35232 21317 35308
rect 21389 35232 21428 35308
rect 20527 34676 20927 34702
rect 20527 34596 20560 34676
rect 20640 34596 20685 34676
rect 20765 34596 20810 34676
rect 20890 34596 20927 34676
rect 20527 34556 20927 34596
rect 20527 34476 20559 34556
rect 20639 34476 20684 34556
rect 20764 34476 20809 34556
rect 20889 34476 20927 34556
rect 20527 34447 20927 34476
rect 21028 33832 21428 35232
rect 21028 33756 21069 33832
rect 21141 33756 21191 33832
rect 21263 33756 21317 33832
rect 21389 33756 21428 33832
rect 21028 33685 21428 33756
rect 21028 33609 21069 33685
rect 21141 33609 21191 33685
rect 21263 33609 21317 33685
rect 21389 33609 21428 33685
rect 21028 33548 21428 33609
rect 21028 33472 21069 33548
rect 21141 33472 21191 33548
rect 21263 33472 21317 33548
rect 21389 33472 21428 33548
rect 21028 33143 21428 33472
rect 20514 33117 21428 33143
rect 20514 33037 21060 33117
rect 21140 33037 21185 33117
rect 21265 33037 21310 33117
rect 21390 33037 21428 33117
rect 20514 32997 21428 33037
rect 20514 32917 21059 32997
rect 21139 32917 21184 32997
rect 21264 32917 21309 32997
rect 21389 32917 21428 32997
rect 20514 32888 21428 32917
rect 21028 32360 21428 32888
rect 21025 32302 21428 32360
rect 21025 32226 21068 32302
rect 21140 32226 21194 32302
rect 21266 32226 21314 32302
rect 21386 32226 21428 32302
rect 21025 32184 21428 32226
rect 21025 32108 21068 32184
rect 21140 32108 21194 32184
rect 21266 32108 21314 32184
rect 21386 32108 21428 32184
rect 21025 32072 21428 32108
rect 463 31760 946 32000
rect 463 31520 863 31760
rect 463 31444 503 31520
rect 575 31444 629 31520
rect 701 31444 749 31520
rect 821 31444 863 31520
rect 463 31402 863 31444
rect 463 31326 503 31402
rect 575 31326 629 31402
rect 701 31326 749 31402
rect 821 31326 863 31402
rect 463 31061 863 31326
rect 21028 31520 21428 32072
rect 21028 31444 21068 31520
rect 21140 31444 21194 31520
rect 21266 31444 21314 31520
rect 21386 31444 21428 31520
rect 21028 31402 21428 31444
rect 21028 31326 21068 31402
rect 21140 31326 21194 31402
rect 21266 31326 21314 31402
rect 21386 31326 21428 31402
rect 953 31120 1155 31121
rect 463 30985 504 31061
rect 576 30985 626 31061
rect 698 30985 752 31061
rect 824 30985 863 31061
rect 463 30914 863 30985
rect 463 30838 504 30914
rect 576 30838 626 30914
rect 698 30838 752 30914
rect 824 30838 863 30914
rect 463 30777 863 30838
rect 463 30701 504 30777
rect 576 30701 626 30777
rect 698 30701 752 30777
rect 824 30701 863 30777
rect 463 29294 863 30701
rect 463 29218 504 29294
rect 576 29218 626 29294
rect 698 29218 752 29294
rect 824 29218 863 29294
rect 463 29147 863 29218
rect 463 29071 504 29147
rect 576 29071 626 29147
rect 698 29071 752 29147
rect 824 29071 863 29147
rect 463 29010 863 29071
rect 463 28934 504 29010
rect 576 28934 626 29010
rect 698 28934 752 29010
rect 824 28934 863 29010
rect 463 28608 863 28934
rect 463 28532 503 28608
rect 575 28532 629 28608
rect 701 28532 749 28608
rect 821 28532 863 28608
rect 463 28490 863 28532
rect 463 28414 503 28490
rect 575 28414 629 28490
rect 701 28414 749 28490
rect 821 28414 863 28490
rect 463 28238 863 28414
rect 21028 28559 21428 31326
rect 21028 28483 21068 28559
rect 21140 28483 21194 28559
rect 21266 28483 21314 28559
rect 21386 28483 21428 28559
rect 21028 28441 21428 28483
rect 21028 28365 21068 28441
rect 21140 28365 21194 28441
rect 21266 28365 21314 28441
rect 21386 28365 21428 28441
rect 463 28209 946 28238
rect 21028 28232 21428 28365
rect 462 27979 946 28209
rect 463 27760 946 27979
rect 20946 27766 21428 28232
rect 463 27604 863 27760
rect 463 27528 503 27604
rect 575 27528 629 27604
rect 701 27528 749 27604
rect 821 27528 863 27604
rect 463 27486 863 27528
rect 463 27410 503 27486
rect 575 27410 629 27486
rect 701 27410 749 27486
rect 821 27410 863 27486
rect 21028 27467 21428 27766
rect 463 27060 863 27410
rect 21027 27442 21428 27467
rect 21027 27366 21068 27442
rect 21140 27366 21194 27442
rect 21266 27366 21314 27442
rect 21386 27366 21428 27442
rect 21027 27324 21428 27366
rect 21027 27248 21068 27324
rect 21140 27248 21194 27324
rect 21266 27248 21314 27324
rect 21386 27248 21428 27324
rect 21027 27212 21428 27248
rect 463 26984 504 27060
rect 576 26984 626 27060
rect 698 26984 752 27060
rect 824 26984 863 27060
rect 463 26913 863 26984
rect 463 26837 504 26913
rect 576 26837 626 26913
rect 698 26837 752 26913
rect 824 26837 863 26913
rect 463 26776 863 26837
rect 463 26700 504 26776
rect 576 26700 626 26776
rect 698 26700 752 26776
rect 824 26700 863 26776
rect 463 25300 863 26700
rect 463 25224 504 25300
rect 576 25224 626 25300
rect 698 25224 752 25300
rect 824 25224 863 25300
rect 463 25153 863 25224
rect 463 25077 504 25153
rect 576 25077 626 25153
rect 698 25077 752 25153
rect 824 25077 863 25153
rect 463 25016 863 25077
rect 463 24940 504 25016
rect 576 24940 626 25016
rect 698 24940 752 25016
rect 824 24940 863 25016
rect 463 24651 863 24940
rect 463 24626 864 24651
rect 463 24550 503 24626
rect 575 24550 629 24626
rect 701 24550 749 24626
rect 821 24550 864 24626
rect 463 24508 864 24550
rect 463 24432 503 24508
rect 575 24432 629 24508
rect 701 24432 749 24508
rect 821 24432 864 24508
rect 463 24396 864 24432
rect 21028 24599 21428 27212
rect 21028 24523 21068 24599
rect 21140 24523 21194 24599
rect 21266 24523 21314 24599
rect 21386 24523 21428 24599
rect 21028 24481 21428 24523
rect 21028 24405 21068 24481
rect 21140 24405 21194 24481
rect 21266 24405 21314 24481
rect 21386 24405 21428 24481
rect 463 24239 863 24396
rect 463 23759 947 24239
rect 21028 24232 21428 24405
rect 20946 23767 21428 24232
rect 463 23569 863 23759
rect 463 23544 864 23569
rect 463 23468 503 23544
rect 575 23468 629 23544
rect 701 23468 749 23544
rect 821 23468 864 23544
rect 463 23426 864 23468
rect 463 23350 503 23426
rect 575 23350 629 23426
rect 701 23350 749 23426
rect 821 23350 864 23426
rect 463 23314 864 23350
rect 21028 23424 21428 23767
rect 21028 23348 21068 23424
rect 21140 23348 21194 23424
rect 21266 23348 21314 23424
rect 21386 23348 21428 23424
rect 463 23060 863 23314
rect 463 22984 504 23060
rect 576 22984 626 23060
rect 698 22984 752 23060
rect 824 22984 863 23060
rect 463 22913 863 22984
rect 463 22837 504 22913
rect 576 22837 626 22913
rect 698 22837 752 22913
rect 824 22837 863 22913
rect 463 22776 863 22837
rect 463 22700 504 22776
rect 576 22700 626 22776
rect 698 22700 752 22776
rect 824 22700 863 22776
rect 463 21301 863 22700
rect 463 21225 504 21301
rect 576 21225 626 21301
rect 698 21225 752 21301
rect 824 21225 863 21301
rect 463 21154 863 21225
rect 463 21078 504 21154
rect 576 21078 626 21154
rect 698 21078 752 21154
rect 824 21078 863 21154
rect 463 21017 863 21078
rect 463 20941 504 21017
rect 576 20941 626 21017
rect 698 20941 752 21017
rect 824 20941 863 21017
rect 463 20694 863 20941
rect 21028 23306 21428 23348
rect 21028 23230 21068 23306
rect 21140 23230 21194 23306
rect 21266 23230 21314 23306
rect 21386 23230 21428 23306
rect 463 20669 864 20694
rect 463 20593 503 20669
rect 575 20593 629 20669
rect 701 20593 749 20669
rect 821 20593 864 20669
rect 21028 20608 21428 23230
rect 463 20551 864 20593
rect 463 20475 503 20551
rect 575 20475 629 20551
rect 701 20475 749 20551
rect 821 20475 864 20551
rect 463 20439 864 20475
rect 21027 20583 21428 20608
rect 21027 20507 21068 20583
rect 21140 20507 21194 20583
rect 21266 20507 21314 20583
rect 21386 20507 21428 20583
rect 21027 20465 21428 20507
rect 463 20240 863 20439
rect 21027 20389 21068 20465
rect 21140 20389 21194 20465
rect 21266 20389 21314 20465
rect 21386 20389 21428 20465
rect 21027 20353 21428 20389
rect 463 19760 946 20240
rect 21028 20233 21428 20353
rect 20946 19768 21428 20233
rect 463 19593 863 19760
rect 463 19568 864 19593
rect 463 19492 503 19568
rect 575 19492 629 19568
rect 701 19492 749 19568
rect 821 19492 864 19568
rect 463 19450 864 19492
rect 463 19374 503 19450
rect 575 19374 629 19450
rect 701 19374 749 19450
rect 821 19374 864 19450
rect 21028 19437 21428 19768
rect 463 19338 864 19374
rect 21027 19412 21428 19437
rect 463 19060 863 19338
rect 21027 19336 21068 19412
rect 21140 19336 21194 19412
rect 21266 19336 21314 19412
rect 21386 19336 21428 19412
rect 21027 19294 21428 19336
rect 21027 19218 21068 19294
rect 21140 19218 21194 19294
rect 21266 19218 21314 19294
rect 21386 19218 21428 19294
rect 21027 19182 21428 19218
rect 463 18984 504 19060
rect 576 18984 626 19060
rect 698 18984 752 19060
rect 824 18984 863 19060
rect 463 18913 863 18984
rect 463 18837 504 18913
rect 576 18837 626 18913
rect 698 18837 752 18913
rect 824 18837 863 18913
rect 463 18776 863 18837
rect 463 18700 504 18776
rect 576 18700 626 18776
rect 698 18700 752 18776
rect 824 18700 863 18776
rect 463 17300 863 18700
rect 463 17224 504 17300
rect 576 17224 626 17300
rect 698 17224 752 17300
rect 824 17224 863 17300
rect 463 17153 863 17224
rect 463 17077 504 17153
rect 576 17077 626 17153
rect 698 17077 752 17153
rect 824 17077 863 17153
rect 463 17016 863 17077
rect 463 16940 504 17016
rect 576 16940 626 17016
rect 698 16940 752 17016
rect 824 16940 863 17016
rect 463 16727 863 16940
rect 463 16702 865 16727
rect 463 16626 503 16702
rect 575 16626 629 16702
rect 701 16626 749 16702
rect 821 16626 865 16702
rect 21028 16676 21428 19182
rect 463 16584 865 16626
rect 463 16508 503 16584
rect 575 16508 629 16584
rect 701 16508 749 16584
rect 821 16508 865 16584
rect 463 16472 865 16508
rect 21027 16651 21428 16676
rect 21027 16575 21068 16651
rect 21140 16575 21194 16651
rect 21266 16575 21314 16651
rect 21386 16575 21428 16651
rect 21027 16533 21428 16575
rect 463 16239 863 16472
rect 21027 16457 21068 16533
rect 21140 16457 21194 16533
rect 21266 16457 21314 16533
rect 21386 16457 21428 16533
rect 21027 16421 21428 16457
rect 463 15759 946 16239
rect 21028 16232 21428 16421
rect 20946 15766 21428 16232
rect 463 15511 863 15759
rect 463 15486 866 15511
rect 463 15410 503 15486
rect 575 15410 629 15486
rect 701 15410 749 15486
rect 821 15410 866 15486
rect 21028 15462 21428 15766
rect 463 15368 866 15410
rect 463 15292 503 15368
rect 575 15292 629 15368
rect 701 15292 749 15368
rect 821 15292 866 15368
rect 463 15256 866 15292
rect 21027 15437 21428 15462
rect 21027 15361 21068 15437
rect 21140 15361 21194 15437
rect 21266 15361 21314 15437
rect 21386 15361 21428 15437
rect 21027 15319 21428 15361
rect 463 15060 863 15256
rect 21027 15243 21068 15319
rect 21140 15243 21194 15319
rect 21266 15243 21314 15319
rect 21386 15243 21428 15319
rect 21027 15207 21428 15243
rect 463 14984 504 15060
rect 576 14984 626 15060
rect 698 14984 752 15060
rect 824 14984 863 15060
rect 463 14913 863 14984
rect 463 14837 504 14913
rect 576 14837 626 14913
rect 698 14837 752 14913
rect 824 14837 863 14913
rect 463 14776 863 14837
rect 463 14700 504 14776
rect 576 14700 626 14776
rect 698 14700 752 14776
rect 824 14700 863 14776
rect 463 13300 863 14700
rect 463 13224 504 13300
rect 576 13224 626 13300
rect 698 13224 752 13300
rect 824 13224 863 13300
rect 463 13153 863 13224
rect 463 13077 504 13153
rect 576 13077 626 13153
rect 698 13077 752 13153
rect 824 13077 863 13153
rect 463 13016 863 13077
rect 463 12940 504 13016
rect 576 12940 626 13016
rect 698 12940 752 13016
rect 824 12940 863 13016
rect 463 12646 863 12940
rect 463 12621 864 12646
rect 463 12545 503 12621
rect 575 12545 629 12621
rect 701 12545 749 12621
rect 821 12545 864 12621
rect 463 12503 864 12545
rect 463 12427 503 12503
rect 575 12427 629 12503
rect 701 12427 749 12503
rect 821 12427 864 12503
rect 463 12391 864 12427
rect 21028 12594 21428 15207
rect 21028 12518 21068 12594
rect 21140 12518 21194 12594
rect 21266 12518 21314 12594
rect 21386 12518 21428 12594
rect 21028 12476 21428 12518
rect 21028 12400 21068 12476
rect 21140 12400 21194 12476
rect 21266 12400 21314 12476
rect 21386 12400 21428 12476
rect 463 12238 863 12391
rect 463 11998 947 12238
rect 21028 12233 21428 12400
rect 463 11758 946 11998
rect 20946 11766 21428 12233
rect 463 11524 863 11758
rect 463 11499 864 11524
rect 463 11423 503 11499
rect 575 11423 629 11499
rect 701 11423 749 11499
rect 821 11423 864 11499
rect 21028 11462 21428 11766
rect 463 11381 864 11423
rect 463 11305 503 11381
rect 575 11305 629 11381
rect 701 11305 749 11381
rect 821 11305 864 11381
rect 463 11269 864 11305
rect 21027 11437 21428 11462
rect 21027 11361 21068 11437
rect 21140 11361 21194 11437
rect 21266 11361 21314 11437
rect 21386 11361 21428 11437
rect 21027 11319 21428 11361
rect 463 11061 863 11269
rect 21027 11243 21068 11319
rect 21140 11243 21194 11319
rect 21266 11243 21314 11319
rect 21386 11243 21428 11319
rect 21027 11207 21428 11243
rect 463 10985 504 11061
rect 576 10985 626 11061
rect 698 10985 752 11061
rect 824 10985 863 11061
rect 463 10914 863 10985
rect 463 10838 504 10914
rect 576 10838 626 10914
rect 698 10838 752 10914
rect 824 10838 863 10914
rect 463 10777 863 10838
rect 463 10701 504 10777
rect 576 10701 626 10777
rect 698 10701 752 10777
rect 824 10701 863 10777
rect 463 9299 863 10701
rect 463 9223 504 9299
rect 576 9223 626 9299
rect 698 9223 752 9299
rect 824 9223 863 9299
rect 463 9152 863 9223
rect 463 9076 504 9152
rect 576 9076 626 9152
rect 698 9076 752 9152
rect 824 9076 863 9152
rect 463 9015 863 9076
rect 463 8939 504 9015
rect 576 8939 626 9015
rect 698 8939 752 9015
rect 824 8939 863 9015
rect 463 8639 863 8939
rect 463 8563 503 8639
rect 575 8563 629 8639
rect 701 8563 749 8639
rect 821 8563 863 8639
rect 463 8521 863 8563
rect 463 8445 503 8521
rect 575 8445 629 8521
rect 701 8445 749 8521
rect 821 8445 863 8521
rect 463 8238 863 8445
rect 21028 8594 21428 11207
rect 21028 8518 21068 8594
rect 21140 8518 21194 8594
rect 21266 8518 21314 8594
rect 21386 8518 21428 8594
rect 21028 8476 21428 8518
rect 21028 8400 21068 8476
rect 21140 8400 21194 8476
rect 21266 8400 21314 8476
rect 21386 8400 21428 8476
rect 463 8000 946 8238
rect 21028 8233 21428 8400
rect 463 7760 947 8000
rect 20946 7766 21428 8233
rect 463 7528 863 7760
rect 463 7452 503 7528
rect 575 7452 629 7528
rect 701 7452 749 7528
rect 821 7452 863 7528
rect 21028 7462 21428 7766
rect 463 7410 863 7452
rect 463 7334 503 7410
rect 575 7334 629 7410
rect 701 7334 749 7410
rect 821 7334 863 7410
rect 463 7061 863 7334
rect 21027 7437 21428 7462
rect 21027 7361 21068 7437
rect 21140 7361 21194 7437
rect 21266 7361 21314 7437
rect 21386 7361 21428 7437
rect 21027 7319 21428 7361
rect 21027 7243 21068 7319
rect 21140 7243 21194 7319
rect 21266 7243 21314 7319
rect 21386 7243 21428 7319
rect 21027 7207 21428 7243
rect 463 6985 504 7061
rect 576 6985 626 7061
rect 698 6985 752 7061
rect 824 6985 863 7061
rect 463 6914 863 6985
rect 463 6838 504 6914
rect 576 6838 626 6914
rect 698 6838 752 6914
rect 824 6838 863 6914
rect 463 6777 863 6838
rect 463 6701 504 6777
rect 576 6701 626 6777
rect 698 6701 752 6777
rect 824 6701 863 6777
rect 463 5300 863 6701
rect 463 5224 504 5300
rect 576 5224 626 5300
rect 698 5224 752 5300
rect 824 5224 863 5300
rect 463 5153 863 5224
rect 463 5077 504 5153
rect 576 5077 626 5153
rect 698 5077 752 5153
rect 824 5077 863 5153
rect 463 5016 863 5077
rect 463 4940 504 5016
rect 576 4940 626 5016
rect 698 4940 752 5016
rect 824 4940 863 5016
rect 463 4730 863 4940
rect 463 4705 865 4730
rect 463 4629 503 4705
rect 575 4629 629 4705
rect 701 4629 749 4705
rect 821 4629 865 4705
rect 463 4587 865 4629
rect 463 4511 503 4587
rect 575 4511 629 4587
rect 701 4511 749 4587
rect 821 4511 865 4587
rect 463 4475 865 4511
rect 21028 4594 21428 7207
rect 21028 4518 21068 4594
rect 21140 4518 21194 4594
rect 21266 4518 21314 4594
rect 21386 4518 21428 4594
rect 21028 4476 21428 4518
rect 463 4239 863 4475
rect 21028 4400 21068 4476
rect 21140 4400 21194 4476
rect 21266 4400 21314 4476
rect 21386 4400 21428 4476
rect 463 4000 947 4239
rect 21028 4233 21428 4400
rect 463 3760 946 4000
rect 20946 3766 21428 4233
rect 463 3528 863 3760
rect 463 3452 503 3528
rect 575 3452 629 3528
rect 701 3452 749 3528
rect 821 3452 863 3528
rect 21028 3462 21428 3766
rect 463 3410 863 3452
rect 463 3334 503 3410
rect 575 3334 629 3410
rect 701 3334 749 3410
rect 821 3334 863 3410
rect 463 3061 863 3334
rect 21027 3437 21428 3462
rect 21027 3361 21068 3437
rect 21140 3361 21194 3437
rect 21266 3361 21314 3437
rect 21386 3361 21428 3437
rect 21027 3319 21428 3361
rect 21027 3243 21068 3319
rect 21140 3243 21194 3319
rect 21266 3243 21314 3319
rect 21386 3243 21428 3319
rect 21027 3207 21428 3243
rect 463 2985 504 3061
rect 576 2985 626 3061
rect 698 2985 752 3061
rect 824 2985 863 3061
rect 463 2914 863 2985
rect 463 2838 504 2914
rect 576 2838 626 2914
rect 698 2838 752 2914
rect 824 2838 863 2914
rect 463 2777 863 2838
rect 463 2701 504 2777
rect 576 2701 626 2777
rect 698 2701 752 2777
rect 824 2701 863 2777
rect 463 1300 863 2701
rect 463 1224 504 1300
rect 576 1224 626 1300
rect 698 1224 752 1300
rect 824 1224 863 1300
rect 463 1153 863 1224
rect 463 1077 504 1153
rect 576 1077 626 1153
rect 698 1077 752 1153
rect 824 1077 863 1153
rect 463 1016 863 1077
rect 463 940 504 1016
rect 576 940 626 1016
rect 698 940 752 1016
rect 824 940 863 1016
rect 463 730 863 940
rect 463 705 865 730
rect 463 629 503 705
rect 575 629 629 705
rect 701 629 749 705
rect 821 629 865 705
rect 463 587 865 629
rect 463 511 503 587
rect 575 511 629 587
rect 701 511 749 587
rect 821 511 865 587
rect 463 475 865 511
rect 21028 594 21428 3207
rect 21028 518 21068 594
rect 21140 518 21194 594
rect 21266 518 21314 594
rect 21386 518 21428 594
rect 21028 476 21428 518
rect 463 239 863 475
rect 21028 400 21068 476
rect 21140 400 21194 476
rect 21266 400 21314 476
rect 21386 400 21428 476
rect 463 0 946 239
rect 21028 233 21428 400
rect 20946 0 21428 233
rect 21502 39726 21902 76000
rect 21502 39646 21535 39726
rect 21615 39646 21660 39726
rect 21740 39646 21785 39726
rect 21865 39646 21902 39726
rect 21502 39606 21902 39646
rect 21502 39526 21534 39606
rect 21614 39526 21659 39606
rect 21739 39526 21784 39606
rect 21864 39526 21902 39606
rect 21502 34676 21902 39526
rect 21502 34596 21535 34676
rect 21615 34596 21660 34676
rect 21740 34596 21785 34676
rect 21865 34596 21902 34676
rect 21502 34556 21902 34596
rect 21502 34476 21534 34556
rect 21614 34476 21659 34556
rect 21739 34476 21784 34556
rect 21864 34476 21902 34556
rect 21502 0 21902 34476
rect 21970 74071 22370 76000
rect 21970 73995 22010 74071
rect 22082 73995 22136 74071
rect 22208 73995 22256 74071
rect 22328 73995 22370 74071
rect 21970 73953 22370 73995
rect 21970 73877 22010 73953
rect 22082 73877 22136 73953
rect 22208 73877 22256 73953
rect 22328 73877 22370 73953
rect 21970 70071 22370 73877
rect 21970 69995 22010 70071
rect 22082 69995 22136 70071
rect 22208 69995 22256 70071
rect 22328 69995 22370 70071
rect 21970 69953 22370 69995
rect 21970 69877 22010 69953
rect 22082 69877 22136 69953
rect 22208 69877 22256 69953
rect 22328 69877 22370 69953
rect 21970 66058 22370 69877
rect 21970 65982 22010 66058
rect 22082 65982 22136 66058
rect 22208 65982 22256 66058
rect 22328 65982 22370 66058
rect 21970 65940 22370 65982
rect 21970 65864 22010 65940
rect 22082 65864 22136 65940
rect 22208 65864 22256 65940
rect 22328 65864 22370 65940
rect 21970 62057 22370 65864
rect 21970 61981 22010 62057
rect 22082 61981 22136 62057
rect 22208 61981 22256 62057
rect 22328 61981 22370 62057
rect 21970 61939 22370 61981
rect 21970 61863 22010 61939
rect 22082 61863 22136 61939
rect 22208 61863 22256 61939
rect 22328 61863 22370 61939
rect 21970 58096 22370 61863
rect 21970 58020 22010 58096
rect 22082 58020 22136 58096
rect 22208 58020 22256 58096
rect 22328 58020 22370 58096
rect 21970 57978 22370 58020
rect 21970 57902 22010 57978
rect 22082 57902 22136 57978
rect 22208 57902 22256 57978
rect 22328 57902 22370 57978
rect 21970 54079 22370 57902
rect 21970 54003 22010 54079
rect 22082 54003 22136 54079
rect 22208 54003 22256 54079
rect 22328 54003 22370 54079
rect 21970 53961 22370 54003
rect 21970 53885 22010 53961
rect 22082 53885 22136 53961
rect 22208 53885 22256 53961
rect 22328 53885 22370 53961
rect 21970 50158 22370 53885
rect 21970 50082 22010 50158
rect 22082 50082 22136 50158
rect 22208 50082 22256 50158
rect 22328 50082 22370 50158
rect 21970 50040 22370 50082
rect 21970 49964 22010 50040
rect 22082 49964 22136 50040
rect 22208 49964 22256 50040
rect 22328 49964 22370 50040
rect 21970 45900 22370 49964
rect 21970 45824 22010 45900
rect 22082 45824 22136 45900
rect 22208 45824 22256 45900
rect 22328 45824 22370 45900
rect 21970 45782 22370 45824
rect 21970 45706 22010 45782
rect 22082 45706 22136 45782
rect 22208 45706 22256 45782
rect 22328 45706 22370 45782
rect 21970 43838 22370 45706
rect 21970 43514 22006 43838
rect 22298 43514 22370 43838
rect 21970 36954 22370 43514
rect 21970 36630 22006 36954
rect 22298 36630 22370 36954
rect 21970 30130 22370 36630
rect 21970 30054 22010 30130
rect 22082 30054 22136 30130
rect 22208 30054 22256 30130
rect 22328 30054 22370 30130
rect 21970 30012 22370 30054
rect 21970 29936 22010 30012
rect 22082 29936 22136 30012
rect 22208 29936 22256 30012
rect 22328 29936 22370 30012
rect 21970 25971 22370 29936
rect 21970 25895 22010 25971
rect 22082 25895 22136 25971
rect 22208 25895 22256 25971
rect 22328 25895 22370 25971
rect 21970 25853 22370 25895
rect 21970 25777 22010 25853
rect 22082 25777 22136 25853
rect 22208 25777 22256 25853
rect 22328 25777 22370 25853
rect 21970 22181 22370 25777
rect 21970 22105 22010 22181
rect 22082 22105 22136 22181
rect 22208 22105 22256 22181
rect 22328 22105 22370 22181
rect 21970 22063 22370 22105
rect 21970 21987 22010 22063
rect 22082 21987 22136 22063
rect 22208 21987 22256 22063
rect 22328 21987 22370 22063
rect 21970 18074 22370 21987
rect 21970 17998 22010 18074
rect 22082 17998 22136 18074
rect 22208 17998 22256 18074
rect 22328 17998 22370 18074
rect 21970 17956 22370 17998
rect 21970 17880 22010 17956
rect 22082 17880 22136 17956
rect 22208 17880 22256 17956
rect 22328 17880 22370 17956
rect 21970 14256 22370 17880
rect 21970 14180 22010 14256
rect 22082 14180 22136 14256
rect 22208 14180 22256 14256
rect 22328 14180 22370 14256
rect 21970 14138 22370 14180
rect 21970 14062 22010 14138
rect 22082 14062 22136 14138
rect 22208 14062 22256 14138
rect 22328 14062 22370 14138
rect 21970 10292 22370 14062
rect 21970 10216 22010 10292
rect 22082 10216 22136 10292
rect 22208 10216 22256 10292
rect 22328 10216 22370 10292
rect 21970 10174 22370 10216
rect 21970 10098 22010 10174
rect 22082 10098 22136 10174
rect 22208 10098 22256 10174
rect 22328 10098 22370 10174
rect 21970 6280 22370 10098
rect 21970 6204 22010 6280
rect 22082 6204 22136 6280
rect 22208 6204 22256 6280
rect 22328 6204 22370 6280
rect 21970 6162 22370 6204
rect 21970 6086 22010 6162
rect 22082 6086 22136 6162
rect 22208 6086 22256 6162
rect 22328 6086 22370 6162
rect 21970 2280 22370 6086
rect 21970 2204 22010 2280
rect 22082 2204 22136 2280
rect 22208 2204 22256 2280
rect 22328 2204 22370 2280
rect 21970 2162 22370 2204
rect 21970 2086 22010 2162
rect 22082 2086 22136 2162
rect 22208 2086 22256 2162
rect 22328 2086 22370 2162
rect 21970 0 22370 2086
use adc_noise_decoup_cell1  adc_noise_decoup_cell1_0
array 0 2 4000 0 0 4000
timestamp 1681461446
transform 1 0 8527 0 1 32532
box 0 0 4000 4000
use adc_noise_decoup_cell1  adc_noise_decoup_cell1_1
array 0 4 4000 0 7 4000
timestamp 1681461446
transform 1 0 946 0 1 0
box 0 0 4000 4000
use adc_noise_decoup_cell1  adc_noise_decoup_cell1_3
array 0 4 4000 0 7 4000
timestamp 1681461446
transform 1 0 946 0 1 44000
box 0 0 4000 4000
use nfet_01v8_w500_l500_nf2  nfet_01v8_w500_l500_nf2_0
timestamp 1663599054
transform 1 0 2655 0 1 39031
box -187 -76 187 76
use nfet_01v8_w500_l500_nf2  nfet_01v8_w500_l500_nf2_1
timestamp 1663599054
transform 1 0 2210 0 1 39031
box -187 -76 187 76
use nfet_01v8_w500_l500_nf2  nfet_01v8_w500_l500_nf2_2
timestamp 1663599054
transform 1 0 2612 0 1 36975
box -187 -76 187 76
use nfet_01v8_w500_l500_nf2  nfet_01v8_w500_l500_nf2_3
timestamp 1663599054
transform 1 0 2132 0 1 36975
box -187 -76 187 76
use nfet_01v8_w500_l500_nf2  nfet_01v8_w500_l500_nf2_4
timestamp 1663599054
transform 1 0 1779 0 -1 39031
box -187 -76 187 76
use pfet_01v8_w500_l500_nf2  pfet_01v8_w500_l500_nf2_0
timestamp 1664545144
transform 1 0 2655 0 1 38693
box -224 -36 223 138
use pfet_01v8_w500_l500_nf2  pfet_01v8_w500_l500_nf2_1
timestamp 1664545144
transform 1 0 2210 0 1 38692
box -224 -36 223 138
use pfet_01v8_w500_l500_nf2  pfet_01v8_w500_l500_nf2_2
timestamp 1664545144
transform 1 0 2612 0 1 37213
box -224 -36 223 138
use pfet_01v8_w500_l500_nf2  pfet_01v8_w500_l500_nf2_3
timestamp 1664545144
transform 1 0 2132 0 1 37213
box -224 -36 223 138
use pfet_01v8_w500_l500_nf2  pfet_01v8_w500_l500_nf2_4
timestamp 1664545144
transform 1 0 1779 0 -1 38794
box -224 -36 223 138
use sky130_fd_sc_hd__buf_4  sky130_fd_sc_hd__buf_4_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform -1 0 4169 0 -1 39091
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  sky130_fd_sc_hd__buf_4_1
timestamp 1683767628
transform -1 0 3617 0 -1 39091
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  sky130_fd_sc_hd__buf_4_2
timestamp 1683767628
transform -1 0 4169 0 1 36915
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  sky130_fd_sc_hd__buf_4_3
timestamp 1683767628
transform -1 0 3617 0 1 36915
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s6s_1  sky130_fd_sc_hd__dlymetal6s6s_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 1961 0 1 38003
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s6s_1  sky130_fd_sc_hd__dlymetal6s6s_1_1
timestamp 1683767628
transform 1 0 1961 0 -1 38003
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s6s_1  sky130_fd_sc_hd__dlymetal6s6s_1_2
timestamp 1683767628
transform 1 0 2881 0 1 38003
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s6s_1  sky130_fd_sc_hd__dlymetal6s6s_1_3
timestamp 1683767628
transform 1 0 3801 0 1 38003
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s6s_1  sky130_fd_sc_hd__dlymetal6s6s_1_4
timestamp 1683767628
transform 1 0 2881 0 -1 38003
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s6s_1  sky130_fd_sc_hd__dlymetal6s6s_1_5
timestamp 1683767628
transform 1 0 3801 0 -1 38003
box -38 -48 958 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform -1 0 4721 0 -1 39091
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_1
timestamp 1683767628
transform -1 0 4721 0 1 36915
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_2
timestamp 1683767628
transform -1 0 4445 0 -1 39091
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_3
timestamp 1683767628
transform -1 0 4445 0 1 36915
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_4
timestamp 1683767628
transform 1 0 1409 0 -1 38003
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform -1 0 1961 0 1 38003
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_1
timestamp 1683767628
transform 1 0 1685 0 -1 38003
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 1593 0 1 38003
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1
timestamp 1683767628
transform -1 0 3065 0 -1 39091
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_2
timestamp 1683767628
transform -1 0 3065 0 1 36915
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_3
timestamp 1683767628
transform 1 0 1317 0 -1 38003
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_4
timestamp 1683767628
transform 1 0 1501 0 1 36915
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_5
timestamp 1683767628
transform 1 0 1388 0 -1 39092
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_6
timestamp 1683767628
transform 1 0 4721 0 1 38003
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_7
timestamp 1683767628
transform 1 0 4721 0 -1 38003
box -38 -48 130 592
<< labels >>
flabel metal4 s 0 0 400 76000 0 FreeSans 1600 90 0 0 VDD
port 1 nsew power bidirectional
flabel metal4 s 463 0 863 76000 0 FreeSans 1600 90 0 0 VSS
port 2 nsew ground bidirectional
flabel metal4 2306 39775 2467 40000 0 FreeSans 480 90 0 0 mimtop1
flabel locali 1339 38217 1373 38269 0 FreeSans 800 0 0 0 clk
port 3 nsew signal input
flabel metal1 2919 37023 2956 37058 0 FreeSans 320 180 0 0 phi2
flabel metal1 2900 38829 2937 38876 0 FreeSans 320 180 0 0 phi1_n
flabel metal1 2899 38946 2935 38981 0 FreeSans 320 180 0 0 phi1
flabel metal4 2493 32001 2737 32321 0 FreeSans 480 90 0 0 mimtop2
flabel metal4 4189 39754 4348 40000 0 FreeSans 480 90 0 0 mimbot1
flabel metal4 21028 0 21428 76000 0 FreeSans 1600 90 0 0 VSS
port 2 nsew ground bidirectional
flabel metal4 21502 0 21902 76000 0 FreeSans 1600 90 0 0 VDD
port 1 nsew power bidirectional
rlabel metal2 22306 36596 22370 36986 3 vcm
port 4 nsew signal output
flabel metal1 2867 37131 2904 37178 0 FreeSans 320 180 0 0 phi2_n
<< properties >>
string LEFclass BLOCK
string LEForigin 0 0
string LEFsource USER
<< end >>
