../mag/hgu_sarlogic.spice