* NGSPICE file created from hgu_sw_cap.ext - technology: sky130A

.subckt hgu_sw_cap SW CTOP delay_signal
X0 delay_signal SW x2.CBOT VSUBS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
.ends

