magic
tech sky130A
magscale 1 2
timestamp 1698248449
<< psubdiff >>
rect 356 204 706 208
rect 356 166 398 204
rect 436 166 474 204
rect 512 166 550 204
rect 588 166 626 204
rect 664 166 706 204
rect 356 162 706 166
<< nsubdiff >>
rect 356 784 706 788
rect 356 746 398 784
rect 436 746 474 784
rect 512 746 550 784
rect 588 746 626 784
rect 664 746 706 784
rect 356 742 706 746
<< psubdiffcont >>
rect 398 166 436 204
rect 474 166 512 204
rect 550 166 588 204
rect 626 166 664 204
<< nsubdiffcont >>
rect 398 746 436 784
rect 474 746 512 784
rect 550 746 588 784
rect 626 746 664 784
<< poly >>
rect 516 435 546 451
rect 450 419 546 435
rect 450 385 466 419
rect 500 385 546 419
rect 450 372 546 385
rect 450 369 516 372
<< polycont >>
rect 466 385 500 419
<< locali >>
rect 320 784 742 788
rect 320 746 398 784
rect 436 746 474 784
rect 512 746 550 784
rect 588 746 626 784
rect 664 746 742 784
rect 320 742 742 746
rect 450 385 466 419
rect 500 385 516 419
rect 558 334 592 537
rect 470 208 504 258
rect 320 204 742 208
rect 320 166 398 204
rect 436 166 474 204
rect 512 166 550 204
rect 588 166 626 204
rect 664 166 742 204
rect 320 162 742 166
<< viali >>
rect 398 746 436 784
rect 474 746 512 784
rect 550 746 588 784
rect 626 746 664 784
rect 466 385 500 419
rect 398 166 436 204
rect 474 166 512 204
rect 550 166 588 204
rect 626 166 664 204
<< metal1 >>
rect 320 784 742 790
rect 320 746 398 784
rect 436 746 474 784
rect 512 746 550 784
rect 588 746 626 784
rect 664 746 742 784
rect 320 740 742 746
rect 320 679 742 711
rect 470 646 504 679
rect 450 419 516 429
rect 450 385 466 419
rect 500 385 516 419
rect 450 375 516 385
rect 320 204 742 210
rect 320 166 398 204
rect 436 166 474 204
rect 512 166 550 204
rect 588 166 626 204
rect 664 166 742 204
rect 320 160 742 166
use sky130_fd_pr__nfet_01v8_L8T3GD  sky130_fd_pr__nfet_01v8_L8T3GD_0 /foss/designs/hgu_goss/hgu/mag
timestamp 1697868789
transform 1 0 531 0 1 264
box -73 -28 73 108
use sky130_fd_pr__pfet_01v8_MQX2PY  XM2
timestamp 1697875053
transform 1 0 531 0 1 592
box -211 -153 211 233
<< labels >>
flabel metal1 334 164 360 206 0 FreeSans 160 0 0 0 VSS
port 11 nsew
flabel poly 472 373 494 429 0 FreeSans 160 0 0 0 IN
port 4 nsew
flabel locali 566 388 586 424 0 FreeSans 160 0 0 0 OUT
port 15 nsew
flabel metal1 429 689 456 704 0 FreeSans 160 0 0 0 VREF
port 19 nsew
flabel metal1 330 749 366 776 0 FreeSans 160 0 0 0 VDD
port 17 nsew
<< end >>
