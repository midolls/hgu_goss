* NGSPICE file created from hgu_sarlogic_retimer_flat.ext - technology: sky130A

.subckt hgu_sarlogic_retimer_flat eob delay_code[2] delay_code[1] delay_code[3] sar_logic[1]
+ sar_logic[2] sar_logic[5] sar_logic[4] sar_retimer[1] sar_retimer[0] sar_retimer[3]
+ sar_retimer[2] sar_retimer[5] sar_retimer[4] sar_retimer[6] sar_retimer[7] sar_logic[3]
+ delay_code[0] VSS VDD
X0 a_14018_6401# a_13844_6793# a_14158_6427# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X1 sar_retimer[3] a_17898_6427# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X2 a_16654_5787# a_16236_5787# a_16410_5761# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X3 a_16410_7041# a_16236_7067# a_16550_7433# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X4 VSS a_17191_5121# a_17126_5147# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X5 a_13751_5147# sar_retimer[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X6 a_16922_6109# a_16410_5761# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X7 VSS a_16410_5121# a_16344_5147# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X8 VSS eob a_12385_8002# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X9 a_14530_7389# a_14018_7041# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X10 sar_retimer[2] a_15506_6427# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X11 a_14483_5787# a_14018_5761# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X12 a_16410_5761# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X13 a_18195_9356# x2.x9.output_stack VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X14 x3.X a_18499_9105# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X15 VDD a_16704_7267# a_16654_7067# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X16 VDD a_17191_7041# a_17898_7083# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X17 x2.x3[1].floating delay_code[1] x2.x9.output_stack VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X18 VSS x3.X a_13397_7073# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X19 x1[0].Q_N a_14799_7041# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X20 VDD VDD a_14312_6401# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X21 a_16236_5787# a_15955_5793# a_16143_5787# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X22 VDD x3.X a_13397_5147# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X23 a_14262_7067# a_13844_7067# a_14018_7041# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X24 a_16143_6427# sar_logic[3] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X25 a_14734_7445# a_13397_7073# a_14625_7445# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X26 a_14915_6153# a_14312_5987# a_14799_5761# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X27 a_13928_5513# a_13397_5147# a_13844_5513# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X28 VSS a_14018_7041# a_13952_7445# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X29 a_16236_7067# a_15789_7073# a_16143_7067# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X30 VSS a_14799_5761# a_14734_6165# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X31 a_13844_5787# a_13563_5793# a_13751_5787# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X32 VDD VDD a_16704_7267# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X33 VDD a_17191_5761# a_17898_5803# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X34 a_14018_7041# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X35 a_13751_6427# sar_logic[2] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X36 a_16654_6709# a_16236_6793# a_16410_6401# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X37 VDD a_17191_6401# a_17103_6793# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X38 VSS x3.X a_13397_5147# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X39 a_14018_7041# a_13844_7067# a_14158_7433# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X40 a_15033_7067# a_14625_7445# a_14799_7041# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X41 VDD a_16410_6401# a_16320_6793# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X42 VDD x3.X a_15789_5793# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X43 a_16410_5761# a_16236_5787# a_16550_6153# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X44 a_16875_5429# a_16410_5121# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X45 a_13844_7067# a_13397_7073# a_13751_7067# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X46 VSS VDD a_16704_7267# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X47 sar_retimer[1] a_17898_7083# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X48 a_14483_6709# a_14018_6401# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X49 a_17103_5787# a_15955_5793# a_17017_6165# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X50 VDD a_16704_7267# a_17425_7067# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X51 a_14530_6109# a_14018_5761# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X52 a_17307_6153# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X53 VSS a_14018_5121# a_13952_5147# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X54 a_16550_6427# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X55 VDD a_14799_7041# a_15506_7083# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X56 a_15955_7073# a_15789_7073# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X57 a_16922_5147# a_16410_5121# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X58 VDD a_14312_5121# a_14262_5429# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X59 sar_retimer[0] a_15506_7083# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X60 a_17191_6401# a_17017_6427# a_17307_6427# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X61 a_14711_5787# a_13563_5793# a_14625_6165# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X62 x2.x9.output_stack x2.x10.Y x2.x5[7].floating VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X63 a_12385_8278# eob a_12297_8278# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X64 a_14915_6153# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X65 VSS VDD a_16704_5121# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X66 VDD VDD a_14312_5121# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X67 VSS VDD a_14312_6401# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X68 VSS a_17191_6401# a_17898_6427# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X69 a_16143_5147# sar_retimer[7] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X70 a_17017_6165# a_15789_5793# a_16875_5787# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X71 a_18195_9015# x2.x9.output_stack VSS VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X72 a_16320_6793# a_15789_6427# a_16236_6793# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X73 VDD a_14799_5761# a_15506_5803# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X74 x1[7].Q_N a_17191_5121# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X75 VDD a_17191_5121# a_17103_5513# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X76 a_14915_5147# a_14312_5121# a_14799_5121# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X77 a_13751_5147# sar_retimer[6] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X78 a_17191_7041# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X79 VDD a_14018_6401# a_13928_6793# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X80 x1[2].Q_N a_14799_6401# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X81 VDD x3.X a_13397_5793# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X82 a_14018_5761# a_13844_5787# a_14158_6153# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X83 VDD a_16410_5121# a_16320_5513# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X84 a_16550_6427# a_16704_6401# a_16410_6401# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X85 x2.x10.Y delay_code[3] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X86 a_14158_6427# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X87 a_16410_5121# a_16236_5513# a_16550_5147# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X88 VDD a_14312_5121# a_15033_5429# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X89 a_17017_7445# a_15955_7073# a_16922_7389# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X90 a_16344_5147# a_15955_5147# a_16236_5513# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X91 a_18195_9356# x2.x9.output_stack x3.A VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.122 ps=1.42 w=0.42 l=0.15
X92 a_14625_7445# a_13397_7073# a_14483_7067# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X93 VDD a_14799_7041# a_14711_7067# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X94 a_14530_5147# a_14018_5121# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X95 a_12385_8692# eob a_12297_8554# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X96 a_15955_7073# a_15789_7073# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X97 a_17191_7041# a_17017_7445# a_17307_7433# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X98 a_14799_6401# a_14625_6427# a_14915_6427# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X99 x1[6].Q_N a_14799_5121# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X100 a_13952_5147# a_13563_5147# a_13844_5513# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X101 x1[1].Q_N a_17191_7041# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X102 VSS a_14799_6401# a_15506_6427# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X103 a_14799_5761# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X104 sar_retimer[3] a_17898_6427# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X105 VSS x3.X a_15789_5793# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X106 a_16143_5787# sar_logic[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X107 a_15955_5147# a_15789_5147# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X108 a_17425_5787# a_17017_6165# a_17191_5761# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X109 x2.x9.output_stack x2.x10.Y x2.x5[7].floating VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X110 x2.x9.output_stack delay_code[2] x2.x4[3].floating VSS sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X111 a_14625_5147# a_13563_5147# a_14530_5147# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X112 a_12385_8968# eob a_12297_8830# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X113 a_12457_8140# eob a_12385_8278# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X114 a_17126_7445# a_15789_7073# a_17017_7445# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X115 a_13563_6427# a_13397_6427# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X116 a_13751_5787# sar_logic[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X117 VSS a_17191_5761# a_17126_6165# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X118 a_16320_5513# a_15789_5147# a_16236_5513# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X119 x2.x9.output_stack x2.x7.SW x2.x7.floating VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X120 a_18195_9015# x3.A VDD VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X121 sar_retimer[2] a_15506_6427# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X122 VDD a_14018_5121# a_13928_5513# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X123 a_16410_6401# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X124 VSS a_16410_5761# a_16344_6165# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X125 a_15955_5147# a_15789_5147# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X126 x3.X a_18499_9105# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X127 a_16550_7433# a_16704_7267# a_16410_7041# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X128 VDD a_16704_5987# a_16654_5787# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X129 x2.x9.output_stack x2.x10.Y x2.x5[7].floating VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X130 a_13563_6427# a_13397_6427# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X131 x1[4].Q_N a_14799_5761# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X132 sar_retimer[7] a_17898_5147# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X133 a_14018_5121# a_13844_5513# a_14158_5147# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X134 a_16236_6793# a_15955_6427# a_16143_6427# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X135 a_16875_7067# a_16410_7041# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X136 a_14262_5787# a_13844_5787# a_14018_5761# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X137 a_13928_7067# a_13397_7073# a_13844_7067# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X138 sar_retimer[6] a_15506_5147# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X139 a_17191_5761# a_17017_6165# a_17307_6153# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X140 VDD x2.x7.SW x2.x6.SW VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X141 a_14799_7041# a_14625_7445# a_14915_7433# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X142 VDD eob a_12322_10357# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X143 a_13844_6793# a_13563_6427# a_13751_6427# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X144 a_17425_6709# a_17017_6427# a_17191_6401# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X145 VDD VDD a_16704_5987# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X146 x1[5].Q_N a_17191_5761# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X147 VDD a_14312_7267# a_14262_7067# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X148 VSS x3.X a_13397_5793# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X149 a_14018_5761# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X150 x2.x9.output_stack delay_code[1] x2.x3[1].floating VSS sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X151 a_14734_6427# a_13397_6427# a_14625_6427# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X152 a_15033_5787# a_14625_6165# a_14799_5761# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X153 a_12457_8692# eob a_12385_8692# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X154 a_16236_6793# a_15789_6427# a_16143_6427# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X155 sar_retimer[5] a_17898_5803# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X156 a_12410_9943# eob a_12322_9805# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X157 VDD a_16704_6401# a_16654_6709# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X158 a_17103_6793# a_15955_6427# a_17017_6427# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X159 a_14734_6165# a_13397_5793# a_14625_6165# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X160 VDD a_16704_5987# a_17425_5787# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X161 a_16550_7433# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X162 VSS a_14799_6401# a_14734_6427# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X163 VSS a_14018_5761# a_13952_6165# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X164 a_16236_5787# a_15789_5793# a_16143_5787# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X165 a_16410_5121# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X166 a_13844_6793# a_13397_6427# a_13751_6427# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X167 VDD a_17191_6401# a_17898_6427# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X168 a_15955_5793# a_15789_5793# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X169 a_16550_6153# a_16704_5987# a_16410_5761# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X170 a_16654_5429# a_16236_5513# a_16410_5121# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X171 x2.x9.output_stack eob a_12385_8968# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X172 a_14711_6793# a_13563_6427# a_14625_6427# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X173 sar_retimer[4] a_15506_5803# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X174 VDD VDD a_14312_7267# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X175 a_13844_5787# a_13397_5793# a_13751_5787# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X176 VSS VDD a_16704_5987# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X177 a_14262_6709# a_13844_6793# a_14018_6401# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X178 a_16236_5513# a_15955_5147# a_16143_5147# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X179 a_16143_7067# sar_logic[1] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X180 VSS a_17191_7041# a_17898_7083# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X181 a_14483_5429# a_14018_5121# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X182 VSS VDD a_14312_7267# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X183 a_16550_5147# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X184 a_12385_8554# eob a_12297_8554# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X185 a_17307_6427# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X186 a_17307_6427# a_16704_6401# a_17191_6401# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X187 a_14799_5761# a_14625_6165# a_14915_6153# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X188 a_13844_5513# a_13563_5147# a_13751_5147# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X189 a_13751_7067# x1[0].D VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X190 VDD a_14312_7267# a_15033_7067# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X191 VDD a_17191_7041# a_17103_7067# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X192 a_15033_6709# a_14625_6427# a_14799_6401# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X193 a_17017_6427# a_15789_6427# a_16875_6709# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X194 a_13563_7073# a_13397_7073# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X195 a_17191_5121# a_17017_5147# a_17307_5147# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X196 a_17191_5761# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X197 VDD a_16410_7041# a_16320_7067# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X198 a_14915_6427# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X199 VSS a_17191_5121# a_17898_5147# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X200 VDD a_16704_6401# a_17425_6709# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X201 a_17103_5513# a_15955_5147# a_17017_5147# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X202 VSS VDD a_14312_5121# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X203 x2.x5[7].floating x2.x10.Y x2.x9.output_stack VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X204 VDD x3.A a_18499_9105# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X205 VDD x3.A a_18195_9015# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0651 ps=0.73 w=0.42 l=0.15
X206 a_14158_7433# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X207 VSS x3.A a_18499_9105# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X208 VDD a_14799_6401# a_15506_6427# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X209 x2.x5[7].floating x2.x10.Y x2.x9.output_stack VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X210 x1[3].Q_N a_17191_6401# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X211 a_14625_6165# a_13397_5793# a_14483_5787# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X212 x1[6].Q_N a_14799_5121# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X213 a_14711_5513# a_13563_5147# a_14625_5147# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X214 a_12410_9943# eob a_12322_10081# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X215 a_16344_7445# a_15955_7073# a_16236_7067# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X216 VDD a_14799_5761# a_14711_5787# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X217 a_16550_5147# a_16704_5121# a_16410_5121# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X218 a_18195_9356# x3.A VSS VDD sky130_fd_pr__pfet_01v8_hvt ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X219 a_17017_6427# a_15955_6427# a_16922_6427# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X220 VSS a_14799_7041# a_15506_7083# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X221 a_14799_6401# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X222 a_14158_6427# a_14312_6401# a_14018_6401# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X223 a_14158_5147# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X224 a_12410_10219# eob a_12322_10357# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X225 a_13952_7445# a_13563_7073# a_13844_7067# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X226 a_16320_7067# a_15789_7073# a_16236_7067# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X227 a_17307_7433# a_16704_7267# a_17191_7041# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X228 a_17017_6165# a_15955_5793# a_16922_6109# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X229 a_17017_5147# a_15789_5147# a_16875_5429# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X230 VDD x3.X a_15789_6427# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X231 x2.x5[7].floating x2.x10.Y x2.x9.output_stack VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X232 a_14625_7445# a_13563_7073# a_14530_7389# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X233 VDD a_14018_7041# a_13928_7067# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X234 a_15955_5793# a_15789_5793# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X235 a_14799_5121# a_14625_5147# a_14915_5147# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X236 VDD a_18499_9105# x3.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X237 a_12457_8416# eob a_12385_8554# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X238 a_17126_6427# a_15789_6427# a_17017_6427# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X239 VSS a_14799_5121# a_15506_5147# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X240 a_13563_7073# a_13397_7073# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X241 a_16143_6427# sar_logic[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X242 sar_retimer[7] a_17898_5147# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X243 x2.x9.output_stack eob a_12322_9805# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X244 x1[0].Q_N a_14799_7041# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X245 VSS x3.X a_15789_6427# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X246 a_17126_6165# a_15789_5793# a_17017_6165# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X247 a_13563_5147# a_13397_5147# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X248 a_16875_5787# a_16410_5761# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X249 sar_retimer[6] a_15506_5147# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X250 a_12385_8140# eob a_12297_8002# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X251 a_13751_6427# sar_logic[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X252 VSS a_17191_6401# a_17126_6427# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X253 a_13928_5787# a_13397_5793# a_13844_5787# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X254 VSS a_16410_6401# a_16344_6427# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X255 x1[1].Q_N a_17191_7041# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X256 a_13563_5147# a_13397_5147# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X257 a_14018_6401# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X258 VDD VDD a_16704_6401# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X259 a_14799_5121# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X260 a_12385_8416# eob a_12297_8278# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X261 a_14158_7433# a_14312_7267# a_14018_7041# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X262 a_16654_7067# a_16236_7067# a_16410_7041# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X263 VDD a_14312_5987# a_14262_5787# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X264 a_17307_6153# a_16704_5987# a_17191_5761# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X265 VDD x3.X a_13397_6427# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X266 a_14483_7067# a_14018_7041# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X267 sar_retimer[1] a_17898_7083# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X268 x2.x9.output_stack x2.x10.Y x2.x5[7].floating VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X269 VSS a_14799_7041# a_14734_7445# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X270 a_16410_7041# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X271 a_17425_5429# a_17017_5147# a_17191_5121# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X272 sar_retimer[0] a_15506_7083# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X273 VSS x3.X a_13397_6427# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X274 a_16875_6709# a_16410_6401# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X275 x1[4].Q_N a_14799_5761# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X276 VDD VDD a_14312_5987# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X277 a_14734_5147# a_13397_5147# a_14625_5147# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X278 x2.x10.Y delay_code[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X279 a_16236_7067# a_15955_7073# a_16143_7067# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X280 a_16236_5513# a_15789_5147# a_16143_5147# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X281 a_16143_5787# sar_logic[5] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X282 x2.x2.floating delay_code[0] x2.x9.output_stack VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.124 ps=1.43 w=0.42 l=0.15
X283 a_16550_6153# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X284 VDD a_16704_5121# a_16654_5429# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X285 VSS a_14799_5121# a_14734_5147# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X286 a_13844_7067# a_13563_7073# a_13751_7067# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X287 a_17307_7433# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X288 VSS a_14018_6401# a_13952_6427# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X289 VSS x3.A a_18195_9356# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0651 ps=0.73 w=0.42 l=0.15
X290 VDD a_14312_6401# a_14262_6709# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X291 a_13751_5787# sar_logic[4] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X292 VDD a_14312_5987# a_15033_5787# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X293 VDD a_17191_5121# a_17898_5147# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X294 a_13844_5513# a_13397_5147# a_13751_5147# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X295 VDD a_17191_5761# a_17103_5787# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X296 a_17191_6401# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X297 a_16922_6427# a_16410_6401# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X298 VDD VDD a_16704_5121# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X299 a_14018_5121# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X300 a_14915_7433# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X301 VDD x3.X a_15789_7073# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X302 VSS VDD a_16704_6401# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X303 a_13563_5793# a_13397_5793# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X304 a_14158_6153# a_14312_5987# a_14018_5761# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X305 VDD a_16410_5761# a_16320_5787# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X306 a_14262_5429# a_13844_5513# a_14018_5121# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X307 a_12410_10219# eob a_12322_10081# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X308 x2.x9.output_stack x2.x6.SW x2.x6.floating VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X309 x2.x4[3].floating delay_code[2] x2.x9.output_stack VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X310 a_12385_8830# eob a_12297_8830# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X311 a_12457_8140# eob a_12385_8140# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X312 VSS a_17191_5761# a_17898_5803# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X313 a_17103_7067# a_15955_7073# a_17017_7445# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X314 VSS VDD a_14312_5987# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X315 a_17307_5147# a_16704_5121# a_17191_5121# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X316 a_17307_5147# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X317 sar_retimer[5] a_17898_5803# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X318 a_12457_8416# eob a_12385_8416# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X319 x1[3].Q_N a_17191_6401# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X320 a_15033_5429# a_14625_5147# a_14799_5121# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X321 a_14711_7067# a_13563_7073# a_14625_7445# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X322 a_14915_6427# a_14312_6401# a_14799_6401# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X323 sar_retimer[4] a_15506_5803# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X324 a_14625_6427# a_13397_6427# a_14483_6709# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X325 VDD a_14799_6401# a_14711_6793# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X326 a_14915_5147# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X327 VDD a_16704_5121# a_17425_5429# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X328 a_12385_8002# eob a_12297_8002# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X329 a_16410_6401# a_16236_6793# a_16550_6427# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X330 a_14158_6153# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X331 a_17017_7445# a_15789_7073# a_16875_7067# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X332 VDD a_14312_6401# a_15033_6709# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X333 a_16344_6427# a_15955_6427# a_16236_6793# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X334 a_16320_5787# a_15789_5793# a_16236_5787# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X335 VDD a_14799_5121# a_15506_5147# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X336 x1[7].Q_N a_17191_5121# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X337 VSS x2.x7.SW x2.x6.SW VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X338 x2.x9.output_stack delay_code[2] x2.x4[3].floating VSS sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X339 a_16922_7389# a_16410_7041# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X340 a_14530_6427# a_14018_6401# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X341 VDD a_14018_5761# a_13928_5787# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X342 a_17191_5121# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X343 VSS a_18499_9105# x3.X VSS sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X344 VDD x3.X a_13397_7073# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X345 a_16344_6165# a_15955_5793# a_16236_5787# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X346 x2.x5[7].floating x2.x10.Y x2.x9.output_stack VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X347 a_13952_6427# a_13563_6427# a_13844_6793# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X348 x1[2].Q_N a_14799_6401# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X349 VSS a_14799_5761# a_15506_5803# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X350 a_17017_5147# a_15955_5147# a_16922_5147# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X351 a_16143_7067# sar_logic[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X352 a_15955_6427# a_15789_6427# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X353 a_14158_5147# a_14312_5121# a_14018_5121# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X354 x2.x4[3].floating delay_code[2] x2.x9.output_stack VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X355 VSS x3.X a_15789_7073# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X356 a_14625_6427# a_13563_6427# a_14530_6427# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X357 a_13952_6165# a_13563_5793# a_13844_5787# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X358 VDD x3.X a_15789_5147# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X359 a_12457_8692# eob a_12385_8830# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X360 a_13751_7067# x1[0].D VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X361 a_14915_7433# a_14312_7267# a_14799_7041# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X362 VSS a_17191_7041# a_17126_7445# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X363 a_13928_6793# a_13397_6427# a_13844_6793# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X364 a_14625_6165# a_13563_5793# a_14530_6109# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X365 a_14625_5147# a_13397_5147# a_14483_5429# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X366 VSS a_16410_7041# a_16344_7445# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X367 a_15955_6427# a_15789_6427# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X368 a_17126_5147# a_15789_5147# a_17017_5147# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X369 VDD a_14799_5121# a_14711_5513# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X370 a_14799_7041# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X371 x1[5].Q_N a_17191_5761# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X372 a_18195_9015# x2.x9.output_stack x3.A VSS sky130_fd_pr__nfet_01v8 ad=0.0651 pd=0.73 as=0.122 ps=1.42 w=0.42 l=0.15
X373 a_17425_7067# a_17017_7445# a_17191_7041# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X374 a_13563_5793# a_13397_5793# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X375 a_16143_5147# sar_retimer[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X376 VSS x3.X a_15789_5147# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

