magic
tech sky130A
magscale 1 2
timestamp 1698486619
<< pwell >>
rect 1006 4372 1032 4404
rect 1612 4372 1638 4404
rect 1006 3212 1032 3244
rect 1612 3212 1638 3244
<< metal3 >>
rect 686 5182 1964 5184
rect 686 5118 790 5182
rect 854 5118 870 5182
rect 934 5118 950 5182
rect 1014 5118 1030 5182
rect 1094 5118 1110 5182
rect 1174 5118 1190 5182
rect 1254 5118 1396 5182
rect 1460 5118 1476 5182
rect 1540 5118 1556 5182
rect 1620 5118 1636 5182
rect 1700 5118 1716 5182
rect 1780 5118 1796 5182
rect 1860 5118 1964 5182
rect 686 5116 1964 5118
rect 686 4962 752 5116
rect 686 4898 687 4962
rect 751 4898 752 4962
rect 686 4882 752 4898
rect 686 4818 687 4882
rect 751 4818 752 4882
rect 686 4802 752 4818
rect 686 4738 687 4802
rect 751 4738 752 4802
rect 686 4722 752 4738
rect 686 4658 687 4722
rect 751 4658 752 4722
rect 686 4642 752 4658
rect 686 4578 687 4642
rect 751 4578 752 4642
rect 686 4562 752 4578
rect 686 4498 687 4562
rect 751 4498 752 4562
rect 686 4482 752 4498
rect 686 4418 687 4482
rect 751 4418 752 4482
rect 686 4402 752 4418
rect 686 4338 687 4402
rect 751 4338 752 4402
rect 686 4322 752 4338
rect 686 4258 687 4322
rect 751 4258 752 4322
rect 686 4242 752 4258
rect 686 4178 687 4242
rect 751 4178 752 4242
rect 686 4088 752 4178
rect 812 4084 872 5116
rect 932 4024 992 5054
rect 1052 4084 1112 5116
rect 1172 4024 1232 5054
rect 1292 4962 1358 5116
rect 1292 4898 1293 4962
rect 1357 4898 1358 4962
rect 1292 4882 1358 4898
rect 1292 4818 1293 4882
rect 1357 4818 1358 4882
rect 1292 4802 1358 4818
rect 1292 4738 1293 4802
rect 1357 4738 1358 4802
rect 1292 4722 1358 4738
rect 1292 4658 1293 4722
rect 1357 4658 1358 4722
rect 1292 4642 1358 4658
rect 1292 4578 1293 4642
rect 1357 4578 1358 4642
rect 1292 4562 1358 4578
rect 1292 4498 1293 4562
rect 1357 4498 1358 4562
rect 1292 4482 1358 4498
rect 1292 4418 1293 4482
rect 1357 4418 1358 4482
rect 1292 4402 1358 4418
rect 1292 4338 1293 4402
rect 1357 4338 1358 4402
rect 1292 4322 1358 4338
rect 1292 4258 1293 4322
rect 1357 4258 1358 4322
rect 1292 4242 1358 4258
rect 1292 4178 1293 4242
rect 1357 4178 1358 4242
rect 1292 4088 1358 4178
rect 1418 4084 1478 5116
rect 1538 4024 1598 5054
rect 1658 4084 1718 5116
rect 1778 4024 1838 5054
rect 1898 4962 1964 5116
rect 1898 4898 1899 4962
rect 1963 4898 1964 4962
rect 1898 4882 1964 4898
rect 1898 4818 1899 4882
rect 1963 4818 1964 4882
rect 1898 4802 1964 4818
rect 1898 4738 1899 4802
rect 1963 4738 1964 4802
rect 1898 4722 1964 4738
rect 1898 4658 1899 4722
rect 1963 4658 1964 4722
rect 1898 4642 1964 4658
rect 1898 4578 1899 4642
rect 1963 4578 1964 4642
rect 1898 4562 1964 4578
rect 1898 4498 1899 4562
rect 1963 4498 1964 4562
rect 1898 4482 1964 4498
rect 1898 4418 1899 4482
rect 1963 4418 1964 4482
rect 1898 4402 1964 4418
rect 1898 4338 1899 4402
rect 1963 4338 1964 4402
rect 1898 4322 1964 4338
rect 1898 4258 1899 4322
rect 1963 4258 1964 4322
rect 1898 4242 1964 4258
rect 1898 4178 1899 4242
rect 1963 4178 1964 4242
rect 1898 4088 1964 4178
rect 686 4022 1964 4024
rect 686 3958 790 4022
rect 854 3958 870 4022
rect 934 3958 950 4022
rect 1014 3958 1030 4022
rect 1094 3958 1110 4022
rect 1174 3958 1190 4022
rect 1254 3958 1396 4022
rect 1460 3958 1476 4022
rect 1540 3958 1556 4022
rect 1620 3958 1636 4022
rect 1700 3958 1716 4022
rect 1780 3958 1796 4022
rect 1860 3958 1964 4022
rect 686 3956 1964 3958
rect 686 3802 752 3956
rect 686 3738 687 3802
rect 751 3738 752 3802
rect 686 3722 752 3738
rect 686 3658 687 3722
rect 751 3658 752 3722
rect 686 3642 752 3658
rect 686 3578 687 3642
rect 751 3578 752 3642
rect 686 3562 752 3578
rect 686 3498 687 3562
rect 751 3498 752 3562
rect 686 3482 752 3498
rect 686 3418 687 3482
rect 751 3418 752 3482
rect 686 3402 752 3418
rect 686 3338 687 3402
rect 751 3338 752 3402
rect 686 3322 752 3338
rect 686 3258 687 3322
rect 751 3258 752 3322
rect 686 3242 752 3258
rect 686 3178 687 3242
rect 751 3178 752 3242
rect 686 3162 752 3178
rect 686 3098 687 3162
rect 751 3098 752 3162
rect 686 3082 752 3098
rect 686 3018 687 3082
rect 751 3018 752 3082
rect 686 2928 752 3018
rect 812 2924 872 3956
rect 932 2864 992 3894
rect 1052 2924 1112 3956
rect 1172 2864 1232 3894
rect 1292 3802 1358 3956
rect 1292 3738 1293 3802
rect 1357 3738 1358 3802
rect 1292 3722 1358 3738
rect 1292 3658 1293 3722
rect 1357 3658 1358 3722
rect 1292 3642 1358 3658
rect 1292 3578 1293 3642
rect 1357 3578 1358 3642
rect 1292 3562 1358 3578
rect 1292 3498 1293 3562
rect 1357 3498 1358 3562
rect 1292 3482 1358 3498
rect 1292 3418 1293 3482
rect 1357 3418 1358 3482
rect 1292 3402 1358 3418
rect 1292 3338 1293 3402
rect 1357 3338 1358 3402
rect 1292 3322 1358 3338
rect 1292 3258 1293 3322
rect 1357 3258 1358 3322
rect 1292 3242 1358 3258
rect 1292 3178 1293 3242
rect 1357 3178 1358 3242
rect 1292 3162 1358 3178
rect 1292 3098 1293 3162
rect 1357 3098 1358 3162
rect 1292 3082 1358 3098
rect 1292 3018 1293 3082
rect 1357 3018 1358 3082
rect 1292 2928 1358 3018
rect 1418 2924 1478 3956
rect 1538 2864 1598 3894
rect 1658 2924 1718 3956
rect 1778 2864 1838 3894
rect 1898 3802 1964 3956
rect 1898 3738 1899 3802
rect 1963 3738 1964 3802
rect 1898 3722 1964 3738
rect 1898 3658 1899 3722
rect 1963 3658 1964 3722
rect 1898 3642 1964 3658
rect 1898 3578 1899 3642
rect 1963 3578 1964 3642
rect 1898 3562 1964 3578
rect 1898 3498 1899 3562
rect 1963 3498 1964 3562
rect 1898 3482 1964 3498
rect 1898 3418 1899 3482
rect 1963 3418 1964 3482
rect 1898 3402 1964 3418
rect 1898 3338 1899 3402
rect 1963 3338 1964 3402
rect 1898 3322 1964 3338
rect 1898 3258 1899 3322
rect 1963 3258 1964 3322
rect 1898 3242 1964 3258
rect 1898 3178 1899 3242
rect 1963 3178 1964 3242
rect 1898 3162 1964 3178
rect 1898 3098 1899 3162
rect 1963 3098 1964 3162
rect 1898 3082 1964 3098
rect 1898 3018 1899 3082
rect 1963 3018 1964 3082
rect 1898 2928 1964 3018
rect 686 2862 1964 2864
rect 686 2798 790 2862
rect 854 2798 870 2862
rect 934 2798 950 2862
rect 1014 2798 1030 2862
rect 1094 2798 1110 2862
rect 1174 2798 1190 2862
rect 1254 2798 1396 2862
rect 1460 2798 1476 2862
rect 1540 2798 1556 2862
rect 1620 2798 1636 2862
rect 1700 2798 1716 2862
rect 1780 2798 1796 2862
rect 1860 2798 1964 2862
rect 686 2796 1964 2798
<< via3 >>
rect 790 5118 854 5182
rect 870 5118 934 5182
rect 950 5118 1014 5182
rect 1030 5118 1094 5182
rect 1110 5118 1174 5182
rect 1190 5118 1254 5182
rect 1396 5118 1460 5182
rect 1476 5118 1540 5182
rect 1556 5118 1620 5182
rect 1636 5118 1700 5182
rect 1716 5118 1780 5182
rect 1796 5118 1860 5182
rect 687 4898 751 4962
rect 687 4818 751 4882
rect 687 4738 751 4802
rect 687 4658 751 4722
rect 687 4578 751 4642
rect 687 4498 751 4562
rect 687 4418 751 4482
rect 687 4338 751 4402
rect 687 4258 751 4322
rect 687 4178 751 4242
rect 1293 4898 1357 4962
rect 1293 4818 1357 4882
rect 1293 4738 1357 4802
rect 1293 4658 1357 4722
rect 1293 4578 1357 4642
rect 1293 4498 1357 4562
rect 1293 4418 1357 4482
rect 1293 4338 1357 4402
rect 1293 4258 1357 4322
rect 1293 4178 1357 4242
rect 1899 4898 1963 4962
rect 1899 4818 1963 4882
rect 1899 4738 1963 4802
rect 1899 4658 1963 4722
rect 1899 4578 1963 4642
rect 1899 4498 1963 4562
rect 1899 4418 1963 4482
rect 1899 4338 1963 4402
rect 1899 4258 1963 4322
rect 1899 4178 1963 4242
rect 790 3958 854 4022
rect 870 3958 934 4022
rect 950 3958 1014 4022
rect 1030 3958 1094 4022
rect 1110 3958 1174 4022
rect 1190 3958 1254 4022
rect 1396 3958 1460 4022
rect 1476 3958 1540 4022
rect 1556 3958 1620 4022
rect 1636 3958 1700 4022
rect 1716 3958 1780 4022
rect 1796 3958 1860 4022
rect 687 3738 751 3802
rect 687 3658 751 3722
rect 687 3578 751 3642
rect 687 3498 751 3562
rect 687 3418 751 3482
rect 687 3338 751 3402
rect 687 3258 751 3322
rect 687 3178 751 3242
rect 687 3098 751 3162
rect 687 3018 751 3082
rect 1293 3738 1357 3802
rect 1293 3658 1357 3722
rect 1293 3578 1357 3642
rect 1293 3498 1357 3562
rect 1293 3418 1357 3482
rect 1293 3338 1357 3402
rect 1293 3258 1357 3322
rect 1293 3178 1357 3242
rect 1293 3098 1357 3162
rect 1293 3018 1357 3082
rect 1899 3738 1963 3802
rect 1899 3658 1963 3722
rect 1899 3578 1963 3642
rect 1899 3498 1963 3562
rect 1899 3418 1963 3482
rect 1899 3338 1963 3402
rect 1899 3258 1963 3322
rect 1899 3178 1963 3242
rect 1899 3098 1963 3162
rect 1899 3018 1963 3082
rect 790 2798 854 2862
rect 870 2798 934 2862
rect 950 2798 1014 2862
rect 1030 2798 1094 2862
rect 1110 2798 1174 2862
rect 1190 2798 1254 2862
rect 1396 2798 1460 2862
rect 1476 2798 1540 2862
rect 1556 2798 1620 2862
rect 1636 2798 1700 2862
rect 1716 2798 1780 2862
rect 1796 2798 1860 2862
<< metal4 >>
rect 686 5182 1964 5184
rect 686 5118 790 5182
rect 854 5118 870 5182
rect 934 5118 950 5182
rect 1014 5118 1030 5182
rect 1094 5118 1110 5182
rect 1174 5118 1190 5182
rect 1254 5118 1396 5182
rect 1460 5118 1476 5182
rect 1540 5118 1556 5182
rect 1620 5118 1636 5182
rect 1700 5118 1716 5182
rect 1780 5118 1796 5182
rect 1860 5118 1964 5182
rect 686 5116 1964 5118
rect 686 4962 752 5116
rect 686 4898 687 4962
rect 751 4898 752 4962
rect 686 4882 752 4898
rect 686 4818 687 4882
rect 751 4818 752 4882
rect 686 4802 752 4818
rect 686 4738 687 4802
rect 751 4738 752 4802
rect 686 4722 752 4738
rect 686 4658 687 4722
rect 751 4658 752 4722
rect 686 4642 752 4658
rect 686 4578 687 4642
rect 751 4578 752 4642
rect 686 4562 752 4578
rect 686 4498 687 4562
rect 751 4498 752 4562
rect 686 4482 752 4498
rect 686 4418 687 4482
rect 751 4418 752 4482
rect 686 4402 752 4418
rect 686 4338 687 4402
rect 751 4338 752 4402
rect 686 4322 752 4338
rect 686 4258 687 4322
rect 751 4258 752 4322
rect 686 4242 752 4258
rect 686 4178 687 4242
rect 751 4178 752 4242
rect 686 4088 752 4178
rect 812 4024 872 5054
rect 932 4084 992 5116
rect 1052 4024 1112 5054
rect 1172 4084 1232 5116
rect 1292 4962 1358 5116
rect 1292 4898 1293 4962
rect 1357 4898 1358 4962
rect 1292 4882 1358 4898
rect 1292 4818 1293 4882
rect 1357 4818 1358 4882
rect 1292 4802 1358 4818
rect 1292 4738 1293 4802
rect 1357 4738 1358 4802
rect 1292 4722 1358 4738
rect 1292 4658 1293 4722
rect 1357 4658 1358 4722
rect 1292 4642 1358 4658
rect 1292 4578 1293 4642
rect 1357 4578 1358 4642
rect 1292 4562 1358 4578
rect 1292 4498 1293 4562
rect 1357 4498 1358 4562
rect 1292 4482 1358 4498
rect 1292 4418 1293 4482
rect 1357 4418 1358 4482
rect 1292 4402 1358 4418
rect 1292 4338 1293 4402
rect 1357 4338 1358 4402
rect 1292 4322 1358 4338
rect 1292 4258 1293 4322
rect 1357 4258 1358 4322
rect 1292 4242 1358 4258
rect 1292 4178 1293 4242
rect 1357 4178 1358 4242
rect 1292 4088 1358 4178
rect 1418 4024 1478 5054
rect 1538 4084 1598 5116
rect 1658 4024 1718 5054
rect 1778 4084 1838 5116
rect 1898 4962 1964 5116
rect 1898 4898 1899 4962
rect 1963 4898 1964 4962
rect 1898 4882 1964 4898
rect 1898 4818 1899 4882
rect 1963 4818 1964 4882
rect 1898 4802 1964 4818
rect 1898 4738 1899 4802
rect 1963 4738 1964 4802
rect 1898 4722 1964 4738
rect 1898 4658 1899 4722
rect 1963 4658 1964 4722
rect 1898 4642 1964 4658
rect 1898 4578 1899 4642
rect 1963 4578 1964 4642
rect 1898 4562 1964 4578
rect 1898 4498 1899 4562
rect 1963 4498 1964 4562
rect 1898 4482 1964 4498
rect 1898 4418 1899 4482
rect 1963 4418 1964 4482
rect 1898 4402 1964 4418
rect 1898 4338 1899 4402
rect 1963 4338 1964 4402
rect 1898 4322 1964 4338
rect 1898 4258 1899 4322
rect 1963 4258 1964 4322
rect 1898 4242 1964 4258
rect 1898 4178 1899 4242
rect 1963 4178 1964 4242
rect 1898 4088 1964 4178
rect 686 4022 1964 4024
rect 686 3958 790 4022
rect 854 3958 870 4022
rect 934 3958 950 4022
rect 1014 3958 1030 4022
rect 1094 3958 1110 4022
rect 1174 3958 1190 4022
rect 1254 3958 1396 4022
rect 1460 3958 1476 4022
rect 1540 3958 1556 4022
rect 1620 3958 1636 4022
rect 1700 3958 1716 4022
rect 1780 3958 1796 4022
rect 1860 3958 1964 4022
rect 686 3956 1964 3958
rect 686 3802 752 3956
rect 686 3738 687 3802
rect 751 3738 752 3802
rect 686 3722 752 3738
rect 686 3658 687 3722
rect 751 3658 752 3722
rect 686 3642 752 3658
rect 686 3578 687 3642
rect 751 3578 752 3642
rect 686 3562 752 3578
rect 686 3498 687 3562
rect 751 3498 752 3562
rect 686 3482 752 3498
rect 686 3418 687 3482
rect 751 3418 752 3482
rect 686 3402 752 3418
rect 686 3338 687 3402
rect 751 3338 752 3402
rect 686 3322 752 3338
rect 686 3258 687 3322
rect 751 3258 752 3322
rect 686 3242 752 3258
rect 686 3178 687 3242
rect 751 3178 752 3242
rect 686 3162 752 3178
rect 686 3098 687 3162
rect 751 3098 752 3162
rect 686 3082 752 3098
rect 686 3018 687 3082
rect 751 3018 752 3082
rect 686 2928 752 3018
rect 812 2864 872 3894
rect 932 2924 992 3956
rect 1052 2864 1112 3894
rect 1172 2924 1232 3956
rect 1292 3802 1358 3956
rect 1292 3738 1293 3802
rect 1357 3738 1358 3802
rect 1292 3722 1358 3738
rect 1292 3658 1293 3722
rect 1357 3658 1358 3722
rect 1292 3642 1358 3658
rect 1292 3578 1293 3642
rect 1357 3578 1358 3642
rect 1292 3562 1358 3578
rect 1292 3498 1293 3562
rect 1357 3498 1358 3562
rect 1292 3482 1358 3498
rect 1292 3418 1293 3482
rect 1357 3418 1358 3482
rect 1292 3402 1358 3418
rect 1292 3338 1293 3402
rect 1357 3338 1358 3402
rect 1292 3322 1358 3338
rect 1292 3258 1293 3322
rect 1357 3258 1358 3322
rect 1292 3242 1358 3258
rect 1292 3178 1293 3242
rect 1357 3178 1358 3242
rect 1292 3162 1358 3178
rect 1292 3098 1293 3162
rect 1357 3098 1358 3162
rect 1292 3082 1358 3098
rect 1292 3018 1293 3082
rect 1357 3018 1358 3082
rect 1292 2928 1358 3018
rect 1418 2864 1478 3894
rect 1538 2924 1598 3956
rect 1658 2864 1718 3894
rect 1778 2924 1838 3956
rect 1898 3802 1964 3956
rect 1898 3738 1899 3802
rect 1963 3738 1964 3802
rect 1898 3722 1964 3738
rect 1898 3658 1899 3722
rect 1963 3658 1964 3722
rect 1898 3642 1964 3658
rect 1898 3578 1899 3642
rect 1963 3578 1964 3642
rect 1898 3562 1964 3578
rect 1898 3498 1899 3562
rect 1963 3498 1964 3562
rect 1898 3482 1964 3498
rect 1898 3418 1899 3482
rect 1963 3418 1964 3482
rect 1898 3402 1964 3418
rect 1898 3338 1899 3402
rect 1963 3338 1964 3402
rect 1898 3322 1964 3338
rect 1898 3258 1899 3322
rect 1963 3258 1964 3322
rect 1898 3242 1964 3258
rect 1898 3178 1899 3242
rect 1963 3178 1964 3242
rect 1898 3162 1964 3178
rect 1898 3098 1899 3162
rect 1963 3098 1964 3162
rect 1898 3082 1964 3098
rect 1898 3018 1899 3082
rect 1963 3018 1964 3082
rect 1898 2928 1964 3018
rect 686 2862 1964 2864
rect 686 2798 790 2862
rect 854 2798 870 2862
rect 934 2798 950 2862
rect 1014 2798 1030 2862
rect 1094 2798 1110 2862
rect 1174 2798 1190 2862
rect 1254 2798 1396 2862
rect 1460 2798 1476 2862
rect 1540 2798 1556 2862
rect 1620 2798 1636 2862
rect 1700 2798 1716 2862
rect 1780 2798 1796 2862
rect 1860 2798 1964 2862
rect 686 2796 1964 2798
<< labels >>
flabel pwell 1612 3212 1638 3244 0 FreeSans 160 0 0 0 x1[2].SUB
flabel metal4 1554 3546 1580 3578 0 FreeSans 320 0 0 0 x1[2].CBOT
flabel metal4 1672 2956 1698 2988 0 FreeSans 320 0 0 0 x1[2].CTOP
flabel pwell 1006 3212 1032 3244 0 FreeSans 160 0 0 0 x1[0].SUB
flabel metal4 948 3546 974 3578 0 FreeSans 320 0 0 0 x1[0].CBOT
flabel metal4 1066 2956 1092 2988 0 FreeSans 320 0 0 0 x1[0].CTOP
flabel pwell 1006 4372 1032 4404 0 FreeSans 160 0 0 0 x1[1].SUB
flabel metal4 948 4706 974 4738 0 FreeSans 320 0 0 0 x1[1].CBOT
flabel metal4 1066 4116 1092 4148 0 FreeSans 320 0 0 0 x1[1].CTOP
flabel pwell 1612 4372 1638 4404 0 FreeSans 160 0 0 0 x1[3].SUB
flabel metal4 1554 4706 1580 4738 0 FreeSans 320 0 0 0 x1[3].CBOT
flabel metal4 1672 4116 1698 4148 0 FreeSans 320 0 0 0 x1[3].CTOP
<< end >>
