magic
tech sky130A
magscale 1 2
timestamp 1702253744
<< nwell >>
rect 984 3863 1018 3872
rect 984 3845 1039 3863
rect 984 3838 1018 3845
<< psubdiff >>
rect 1806 1934 1822 1982
<< nsubdiff >>
rect 984 3863 1018 3872
rect 984 3845 1039 3863
rect 984 3838 1018 3845
<< poly >>
rect 1148 5162 1466 5192
rect 1532 5162 1658 5192
rect 1148 3979 1475 4010
rect 1440 3966 1475 3979
rect 1628 3989 1694 4010
rect 1440 3950 1507 3966
rect 1440 3916 1457 3950
rect 1491 3916 1507 3950
rect 1628 3955 1644 3989
rect 1678 3955 1694 3989
rect 1628 3943 1694 3955
rect 1440 3900 1507 3916
rect 1476 3631 1543 3647
rect 1476 3611 1493 3631
rect 1436 3597 1493 3611
rect 1527 3597 1543 3631
rect 1436 3581 1543 3597
rect 1617 3626 1684 3642
rect 1617 3592 1633 3626
rect 1667 3592 1684 3626
rect 1436 3568 1466 3581
rect 1617 3576 1684 3592
rect 1148 3537 1466 3568
rect 1628 3536 1658 3576
rect 1532 2905 1658 2935
rect 1532 2717 1658 2747
rect 1148 2084 1466 2115
rect 1436 2071 1466 2084
rect 1628 2076 1658 2116
rect 1436 2055 1543 2071
rect 1436 2041 1493 2055
rect 1476 2021 1493 2041
rect 1527 2021 1543 2055
rect 1476 2005 1543 2021
rect 1617 2060 1684 2076
rect 1617 2026 1633 2060
rect 1667 2026 1684 2060
rect 1617 2010 1684 2026
rect 1440 1736 1507 1752
rect 1440 1702 1457 1736
rect 1491 1702 1507 1736
rect 1440 1686 1507 1702
rect 1628 1697 1694 1709
rect 1440 1673 1475 1686
rect 1148 1642 1475 1673
rect 1628 1663 1644 1697
rect 1678 1663 1694 1697
rect 1628 1642 1694 1663
rect 1148 460 1466 491
rect 1532 460 1658 490
<< polycont >>
rect 1457 3916 1491 3950
rect 1644 3955 1678 3989
rect 1493 3597 1527 3631
rect 1633 3592 1667 3626
rect 1493 2021 1527 2055
rect 1633 2026 1667 2060
rect 1457 1702 1491 1736
rect 1644 1663 1678 1697
<< locali >>
rect 1628 3955 1644 3989
rect 1678 3955 1694 3989
rect 1441 3916 1457 3950
rect 1491 3916 1507 3950
rect 1018 3845 1039 3863
rect 1477 3597 1493 3631
rect 1527 3597 1543 3631
rect 1633 3626 1667 3642
rect 1633 3576 1667 3592
rect 995 2819 1026 2838
rect 1633 2060 1667 2076
rect 1477 2021 1493 2055
rect 1527 2021 1543 2055
rect 1633 2010 1667 2026
rect 1806 1934 1822 1982
rect 1441 1702 1457 1736
rect 1491 1702 1507 1736
rect 1628 1663 1644 1697
rect 1678 1663 1694 1697
<< viali >>
rect 1644 3955 1678 3989
rect 1457 3916 1491 3950
rect 984 3838 1018 3872
rect 1493 3597 1527 3631
rect 1633 3592 1667 3626
rect 1493 2021 1527 2055
rect 1633 2026 1667 2060
rect 984 1783 1018 1817
rect 1457 1702 1491 1736
rect 1644 1663 1678 1697
<< metal1 >>
rect 51660 8985 51724 8991
rect 51660 8933 51666 8985
rect 51718 8977 51724 8985
rect 53592 8985 53656 8991
rect 53592 8977 53598 8985
rect 51718 8940 53598 8977
rect 51718 8933 51724 8940
rect 51660 8927 51724 8933
rect 53592 8933 53598 8940
rect 53650 8933 53656 8985
rect 53592 8927 53656 8933
rect 51551 7952 51615 7958
rect 51551 7900 51557 7952
rect 51609 7945 51615 7952
rect 53481 7954 53545 7960
rect 53481 7945 53487 7954
rect 51609 7908 53487 7945
rect 51609 7900 51615 7908
rect 51551 7894 51615 7900
rect 53481 7902 53487 7908
rect 53539 7902 53545 7954
rect 53481 7896 53545 7902
rect 53589 7109 53653 7115
rect 53589 7057 53595 7109
rect 53647 7057 53653 7109
rect 53589 7051 53653 7057
rect 53492 6079 53556 6085
rect 1611 6035 1723 6042
rect 1611 5933 1617 6035
rect 1716 5933 1723 6035
rect 53492 6027 53498 6079
rect 53550 6074 53556 6079
rect 53550 6037 53595 6074
rect 53550 6027 53556 6037
rect 53492 6021 53556 6027
rect 1611 5928 1723 5933
rect 1627 5209 1708 5928
rect 1098 5175 1708 5209
rect 1098 5124 1132 5175
rect 1290 5124 1324 5175
rect 1482 5124 1516 5175
rect 1578 5124 1612 5175
rect 1674 5124 1708 5175
rect 1709 4036 1799 4070
rect 1635 4002 1687 4008
rect 1289 3975 1323 3980
rect 379 3903 505 3913
rect 379 3797 389 3903
rect 495 3879 505 3903
rect 495 3872 1030 3879
rect 495 3838 984 3872
rect 1018 3838 1030 3872
rect 495 3831 1030 3838
rect 495 3797 505 3831
rect 379 3787 505 3797
rect 918 3701 1044 3711
rect 918 3595 928 3701
rect 1034 3668 1044 3701
rect 1289 3668 1323 3974
rect 1448 3959 1500 3965
rect 1631 3955 1635 3989
rect 1687 3955 1691 3989
rect 1444 3916 1448 3950
rect 1500 3916 1504 3950
rect 1635 3944 1687 3950
rect 1448 3901 1500 3907
rect 1034 3634 1323 3668
rect 1034 3595 1044 3634
rect 918 3585 1044 3595
rect 1289 3573 1323 3634
rect 1484 3640 1536 3646
rect 1633 3635 1667 3639
rect 1480 3597 1484 3631
rect 1536 3597 1540 3631
rect 1484 3582 1536 3588
rect 1618 3583 1624 3635
rect 1676 3583 1682 3635
rect 1633 3579 1667 3583
rect 1194 3539 1420 3573
rect 1765 3511 1799 4036
rect 1708 3477 1799 3511
rect 1714 3476 1799 3477
rect 1578 2888 1612 2973
rect 1674 2888 1708 2973
rect 1578 2679 1612 2764
rect 1674 2679 1708 2764
rect 1708 2141 1785 2175
rect 1194 2079 1420 2113
rect 918 2047 1044 2057
rect 918 1941 928 2047
rect 1034 2018 1044 2047
rect 1289 2018 1323 2079
rect 1484 2064 1536 2070
rect 1633 2069 1667 2073
rect 1480 2021 1484 2055
rect 1536 2021 1540 2055
rect 1034 1984 1323 2018
rect 1618 2017 1624 2069
rect 1676 2017 1682 2069
rect 1633 2013 1667 2017
rect 1484 2006 1536 2012
rect 1034 1941 1044 1984
rect 918 1931 1044 1941
rect 376 1847 502 1857
rect 376 1741 386 1847
rect 492 1829 502 1847
rect 492 1817 1030 1829
rect 492 1783 984 1817
rect 1018 1783 1030 1817
rect 492 1771 1030 1783
rect 492 1741 502 1771
rect 376 1731 502 1741
rect 1289 1678 1323 1984
rect 1448 1745 1500 1751
rect 1444 1702 1448 1736
rect 1500 1702 1504 1736
rect 1635 1702 1687 1708
rect 1448 1687 1500 1693
rect 1289 1672 1323 1677
rect 1631 1663 1635 1697
rect 1687 1663 1691 1697
rect 1635 1644 1687 1650
rect 1751 1616 1785 2141
rect 1714 1582 1785 1616
rect 1098 477 1132 528
rect 1290 477 1324 528
rect 1482 477 1516 528
rect 1578 477 1612 528
rect 1674 477 1708 529
rect 1098 443 1708 477
rect 1627 -241 1708 443
rect 1612 -246 1724 -241
rect 1612 -348 1619 -246
rect 1718 -348 1724 -246
rect 1612 -355 1724 -348
<< via1 >>
rect 51666 8933 51718 8985
rect 53598 8933 53650 8985
rect 51557 7900 51609 7952
rect 53487 7902 53539 7954
rect 53595 7057 53647 7109
rect 1617 5933 1716 6035
rect 53498 6027 53550 6079
rect 1635 3989 1687 4002
rect 389 3797 495 3903
rect 928 3595 1034 3701
rect 1448 3950 1500 3959
rect 1635 3955 1644 3989
rect 1644 3955 1678 3989
rect 1678 3955 1687 3989
rect 1635 3950 1687 3955
rect 1448 3916 1457 3950
rect 1457 3916 1491 3950
rect 1491 3916 1500 3950
rect 1448 3907 1500 3916
rect 1484 3631 1536 3640
rect 1484 3597 1493 3631
rect 1493 3597 1527 3631
rect 1527 3597 1536 3631
rect 1484 3588 1536 3597
rect 1624 3626 1676 3635
rect 1624 3592 1633 3626
rect 1633 3592 1667 3626
rect 1667 3592 1676 3626
rect 1624 3583 1676 3592
rect 928 1941 1034 2047
rect 1484 2055 1536 2064
rect 1484 2021 1493 2055
rect 1493 2021 1527 2055
rect 1527 2021 1536 2055
rect 1484 2012 1536 2021
rect 1624 2060 1676 2069
rect 1624 2026 1633 2060
rect 1633 2026 1667 2060
rect 1667 2026 1676 2060
rect 1624 2017 1676 2026
rect 386 1741 492 1847
rect 1448 1736 1500 1745
rect 1448 1702 1457 1736
rect 1457 1702 1491 1736
rect 1491 1702 1500 1736
rect 1448 1693 1500 1702
rect 1635 1697 1687 1702
rect 1635 1663 1644 1697
rect 1644 1663 1678 1697
rect 1678 1663 1687 1697
rect 1635 1650 1687 1663
rect 1619 -348 1718 -246
<< metal2 >>
rect 51390 13547 51587 13556
rect 1880 13507 2046 13516
rect 1880 13363 1889 13507
rect 2037 13363 2046 13507
rect 1880 13353 2046 13363
rect 51390 13362 51398 13547
rect 51578 13467 51587 13547
rect 51578 13434 51712 13467
rect 51578 13362 51587 13434
rect 51390 13353 51587 13362
rect 1939 13336 1984 13353
rect 1722 12519 1888 12528
rect 1722 12375 1731 12519
rect 1879 12375 1888 12519
rect 1722 12365 1888 12375
rect 1789 12348 1862 12365
rect 1829 9815 1862 12348
rect 1597 6044 1736 6054
rect 1597 5923 1607 6044
rect 1727 5923 1736 6044
rect 1597 5913 1736 5923
rect 1629 4002 1694 4009
rect 1442 3959 1506 3965
rect 369 3787 379 3913
rect 505 3787 515 3913
rect 1442 3907 1448 3959
rect 1500 3907 1506 3959
rect 1629 3950 1635 4002
rect 1687 3972 1694 4002
rect 1687 3950 1701 3972
rect 1629 3944 1701 3950
rect 1442 3901 1506 3907
rect 1442 3738 1476 3901
rect 1667 3873 1701 3944
rect 1508 3864 1564 3873
rect 1508 3799 1564 3808
rect 1673 3864 1729 3873
rect 1673 3799 1729 3808
rect 908 3585 918 3711
rect 1044 3585 1054 3711
rect 1406 3682 1415 3738
rect 1471 3682 1480 3738
rect 1508 3646 1542 3799
rect 1829 3740 1863 9815
rect 1939 3880 1973 13336
rect 51279 12547 51476 12556
rect 51279 12362 51287 12547
rect 51467 12467 51476 12547
rect 51467 12434 51601 12467
rect 51467 12362 51476 12434
rect 51279 12353 51476 12362
rect 51564 7958 51601 12434
rect 51675 8991 51712 13434
rect 51660 8985 51724 8991
rect 51660 8933 51666 8985
rect 51718 8933 51724 8985
rect 51660 8927 51724 8933
rect 53592 8985 53656 8991
rect 53592 8933 53598 8985
rect 53650 8933 53656 8985
rect 53592 8927 53656 8933
rect 51551 7952 51615 7958
rect 51551 7900 51557 7952
rect 51609 7900 51615 7952
rect 51551 7894 51615 7900
rect 53481 7954 53545 7960
rect 53481 7902 53487 7954
rect 53539 7902 53545 7954
rect 53481 7896 53545 7902
rect 53495 6085 53532 7896
rect 53606 7115 53643 8927
rect 53589 7109 53653 7115
rect 53589 7057 53595 7109
rect 53647 7057 53653 7109
rect 53589 7051 53653 7057
rect 53492 6079 53556 6085
rect 53492 6027 53498 6079
rect 53550 6027 53556 6079
rect 53492 6021 53556 6027
rect 1915 3871 1989 3880
rect 1915 3815 1924 3871
rect 1980 3815 1989 3871
rect 1915 3806 1989 3815
rect 1570 3682 1580 3738
rect 1636 3721 1645 3738
rect 1812 3731 1887 3740
rect 1636 3682 1660 3721
rect 1478 3640 1542 3646
rect 1626 3641 1660 3682
rect 1812 3675 1822 3731
rect 1878 3675 1887 3731
rect 1812 3666 1887 3675
rect 1478 3588 1484 3640
rect 1536 3588 1542 3640
rect 1478 3582 1542 3588
rect 1618 3635 1682 3641
rect 1618 3583 1624 3635
rect 1676 3583 1682 3635
rect 1618 3577 1682 3583
rect 1478 2064 1542 2070
rect 908 1931 918 2057
rect 1044 1931 1054 2057
rect 1478 2012 1484 2064
rect 1536 2012 1542 2064
rect 1478 2006 1542 2012
rect 1618 2069 1682 2075
rect 1618 2017 1624 2069
rect 1676 2017 1682 2069
rect 1618 2011 1682 2017
rect 1406 1915 1415 1971
rect 1471 1915 1480 1971
rect 366 1731 376 1857
rect 502 1731 512 1857
rect 1442 1751 1476 1915
rect 1508 1853 1542 2006
rect 1626 1971 1660 2011
rect 1830 1982 1864 3666
rect 1570 1915 1580 1971
rect 1636 1934 1660 1971
rect 1806 1973 1888 1982
rect 1636 1915 1645 1934
rect 1806 1917 1815 1973
rect 1878 1917 1888 1973
rect 1806 1908 1888 1917
rect 1508 1844 1564 1853
rect 1508 1779 1564 1788
rect 1673 1844 1729 1853
rect 1939 1848 1973 3806
rect 1673 1779 1729 1788
rect 1906 1839 1980 1848
rect 1906 1783 1915 1839
rect 1971 1783 1980 1839
rect 1442 1745 1506 1751
rect 1442 1693 1448 1745
rect 1500 1693 1506 1745
rect 1667 1708 1701 1779
rect 1906 1774 1980 1783
rect 1442 1687 1506 1693
rect 1629 1702 1701 1708
rect 1629 1650 1635 1702
rect 1687 1680 1701 1702
rect 1687 1650 1694 1680
rect 1629 1643 1694 1650
rect 1599 -236 1738 -226
rect 1599 -357 1608 -236
rect 1728 -357 1738 -236
rect 1599 -367 1738 -357
<< via2 >>
rect 1889 13363 2037 13507
rect 51398 13362 51578 13547
rect 1731 12375 1879 12519
rect 1607 6035 1727 6044
rect 1607 5933 1617 6035
rect 1617 5933 1716 6035
rect 1716 5933 1727 6035
rect 1607 5923 1727 5933
rect 379 3903 505 3913
rect 379 3797 389 3903
rect 389 3797 495 3903
rect 495 3797 505 3903
rect 379 3787 505 3797
rect 1508 3808 1564 3864
rect 1673 3808 1729 3864
rect 918 3701 1044 3711
rect 918 3595 928 3701
rect 928 3595 1034 3701
rect 1034 3595 1044 3701
rect 918 3585 1044 3595
rect 1415 3682 1471 3738
rect 51287 12362 51467 12547
rect 1924 3815 1980 3871
rect 1580 3682 1636 3738
rect 1822 3675 1878 3731
rect 918 2047 1044 2057
rect 918 1941 928 2047
rect 928 1941 1034 2047
rect 1034 1941 1044 2047
rect 918 1931 1044 1941
rect 1415 1915 1471 1971
rect 376 1847 502 1857
rect 376 1741 386 1847
rect 386 1741 492 1847
rect 492 1741 502 1847
rect 376 1731 502 1741
rect 1580 1915 1636 1971
rect 1815 1917 1878 1973
rect 1508 1788 1564 1844
rect 1673 1788 1729 1844
rect 1915 1783 1971 1839
rect 1608 -246 1728 -236
rect 1608 -348 1619 -246
rect 1619 -348 1718 -246
rect 1718 -348 1728 -246
rect 1608 -357 1728 -348
<< metal3 >>
rect 51368 13561 51604 13562
rect 1861 13533 2066 13539
rect 1861 13336 1867 13533
rect 2060 13336 2066 13533
rect 51368 13348 51381 13561
rect 51592 13348 51604 13561
rect 1861 13330 2066 13336
rect 51257 12561 51493 12562
rect 1703 12545 1908 12551
rect 1703 12348 1709 12545
rect 1902 12348 1908 12545
rect 51257 12348 51270 12561
rect 51481 12348 51493 12561
rect 1703 12342 1908 12348
rect 1573 6071 1761 6078
rect 1573 5895 1579 6071
rect 1756 5895 1761 6071
rect 1573 5889 1761 5895
rect 363 3780 369 3920
rect 515 3780 521 3920
rect 1915 3871 1989 3880
rect 1503 3866 1734 3869
rect 1915 3866 1924 3871
rect 1503 3864 1924 3866
rect 1503 3808 1508 3864
rect 1564 3808 1673 3864
rect 1729 3815 1924 3864
rect 1980 3815 1989 3871
rect 1729 3808 1989 3815
rect 1503 3806 1989 3808
rect 1503 3803 1734 3806
rect 1406 3740 1641 3743
rect 1406 3738 1887 3740
rect 902 3578 908 3718
rect 1054 3578 1060 3718
rect 1406 3682 1415 3738
rect 1471 3682 1580 3738
rect 1636 3731 1887 3738
rect 1636 3682 1822 3731
rect 1406 3680 1822 3682
rect 1406 3677 1641 3680
rect 1812 3675 1822 3680
rect 1878 3675 1887 3731
rect 1812 3666 1887 3675
rect 902 1924 908 2064
rect 1054 1924 1060 2064
rect 1410 1971 1641 1977
rect 1410 1915 1415 1971
rect 1471 1915 1580 1971
rect 1636 1969 1641 1971
rect 1806 1973 1888 1982
rect 1806 1969 1815 1973
rect 1636 1917 1815 1969
rect 1878 1917 1888 1973
rect 1636 1915 1888 1917
rect 1410 1909 1888 1915
rect 1806 1908 1888 1909
rect 360 1724 366 1864
rect 512 1724 518 1864
rect 1503 1848 1734 1849
rect 1503 1844 1980 1848
rect 1503 1788 1508 1844
rect 1564 1788 1673 1844
rect 1729 1839 1980 1844
rect 1729 1788 1915 1839
rect 1503 1783 1734 1788
rect 1906 1783 1915 1788
rect 1971 1783 1980 1839
rect 1906 1774 1980 1783
rect 1574 -208 1762 -202
rect 1574 -384 1579 -208
rect 1756 -384 1762 -208
rect 1574 -391 1762 -384
<< via3 >>
rect 1867 13507 2060 13533
rect 1867 13363 1889 13507
rect 1889 13363 2037 13507
rect 2037 13363 2060 13507
rect 1867 13336 2060 13363
rect 51381 13547 51592 13561
rect 51381 13362 51398 13547
rect 51398 13362 51578 13547
rect 51578 13362 51592 13547
rect 51381 13348 51592 13362
rect 1709 12519 1902 12545
rect 1709 12375 1731 12519
rect 1731 12375 1879 12519
rect 1879 12375 1902 12519
rect 1709 12348 1902 12375
rect 51270 12547 51481 12561
rect 51270 12362 51287 12547
rect 51287 12362 51467 12547
rect 51467 12362 51481 12547
rect 51270 12348 51481 12362
rect 1579 6044 1756 6071
rect 1579 5923 1607 6044
rect 1607 5923 1727 6044
rect 1727 5923 1756 6044
rect 1579 5895 1756 5923
rect 369 3913 515 3920
rect 369 3787 379 3913
rect 379 3787 505 3913
rect 505 3787 515 3913
rect 369 3780 515 3787
rect 908 3711 1054 3718
rect 908 3585 918 3711
rect 918 3585 1044 3711
rect 1044 3585 1054 3711
rect 908 3578 1054 3585
rect 908 2057 1054 2064
rect 908 1931 918 2057
rect 918 1931 1044 2057
rect 1044 1931 1054 2057
rect 908 1924 1054 1931
rect 366 1857 512 1864
rect 366 1731 376 1857
rect 376 1731 502 1857
rect 502 1731 512 1857
rect 366 1724 512 1731
rect 1579 -236 1756 -208
rect 1579 -357 1608 -236
rect 1608 -357 1728 -236
rect 1728 -357 1756 -236
rect 1579 -384 1756 -357
<< metal4 >>
rect 51253 12572 51505 12573
rect 51253 12336 51257 12572
rect 51493 12336 51505 12572
rect 1622 7512 2241 7580
rect 1622 6102 1700 7512
rect 339 3920 545 3935
rect 339 3780 369 3920
rect 515 3780 545 3920
rect 339 1864 545 3780
rect 339 1724 366 1864
rect 512 1724 545 1864
rect 339 1688 545 1724
rect 1622 -1830 1700 -415
rect 1622 -1898 2241 -1830
<< via4 >>
rect 51368 13561 51604 13572
rect 1838 13533 2092 13557
rect 1838 13336 1867 13533
rect 1867 13336 2060 13533
rect 2060 13336 2092 13533
rect 51368 13348 51381 13561
rect 51381 13348 51592 13561
rect 51592 13348 51604 13561
rect 51368 13336 51604 13348
rect 1838 13308 2092 13336
rect 1680 12545 1934 12569
rect 1680 12348 1709 12545
rect 1709 12348 1902 12545
rect 1902 12348 1934 12545
rect 1680 12320 1934 12348
rect 51257 12561 51493 12572
rect 51257 12348 51270 12561
rect 51270 12348 51481 12561
rect 51481 12348 51493 12561
rect 51257 12336 51493 12348
rect 1549 6071 1786 6102
rect 1549 5895 1579 6071
rect 1579 5895 1756 6071
rect 1756 5895 1786 6071
rect 1549 5866 1786 5895
rect 806 3718 1060 3816
rect 806 3578 908 3718
rect 908 3578 1054 3718
rect 1054 3578 1060 3718
rect 806 3560 1060 3578
rect 806 2064 1060 2094
rect 806 1924 908 2064
rect 908 1924 1054 2064
rect 1054 1924 1060 2064
rect 806 1838 1060 1924
rect 1549 -208 1786 -179
rect 1549 -384 1579 -208
rect 1579 -384 1756 -208
rect 1756 -384 1786 -208
rect 1549 -415 1786 -384
<< metal5 >>
rect 1812 13572 51630 13597
rect 1812 13557 51368 13572
rect 1812 13308 1838 13557
rect 2092 13336 51368 13557
rect 51604 13336 51630 13572
rect 2092 13308 51630 13336
rect 1812 13277 51630 13308
rect 1655 12572 51519 12604
rect 1655 12569 51257 12572
rect 1655 12320 1680 12569
rect 1934 12336 51257 12569
rect 51493 12336 51519 12572
rect 1934 12320 51519 12336
rect 1655 12284 51519 12320
rect 1503 6102 42326 6145
rect 1503 5866 1549 6102
rect 1786 5866 42326 6102
rect 1503 5813 42326 5866
rect 554 3816 1110 3852
rect 554 3560 806 3816
rect 1060 3560 1110 3816
rect 554 3530 1110 3560
rect 554 2094 1110 2130
rect 554 1838 806 2094
rect 1060 1838 1110 2094
rect 554 1808 1110 1838
rect 1504 -179 42326 -131
rect 1504 -415 1549 -179
rect 1786 -415 42326 -179
rect 1504 -463 42326 -415
rect 1504 -465 2198 -463
use sky130_fd_pr__nfet_01v8_5AY3TR  sky130_fd_pr__nfet_01v8_5AY3TR_0
timestamp 1699633464
transform 1 0 1595 0 1 3236
box -145 -427 227 482
use sky130_fd_pr__nfet_01v8_5AY3TR  sky130_fd_pr__nfet_01v8_5AY3TR_1
timestamp 1699633464
transform 1 0 1595 0 -1 2416
box -145 -427 227 482
use sky130_fd_pr__nfet_01v8_YCY3T5  sky130_fd_pr__nfet_01v8_YCY3T5_0
timestamp 1699707102
transform 1 0 1307 0 -1 2416
box -323 -427 401 482
use sky130_fd_pr__nfet_01v8_YCY3T5  sky130_fd_pr__nfet_01v8_YCY3T5_1
timestamp 1699707102
transform 1 0 1307 0 1 3236
box -323 -427 401 482
use sky130_fd_pr__pfet_01v8_UJB66J  sky130_fd_pr__pfet_01v8_UJB66J_0
timestamp 1699707026
transform 1 0 1595 0 -1 1066
box -263 -787 263 769
use sky130_fd_pr__pfet_01v8_UJB66J  sky130_fd_pr__pfet_01v8_UJB66J_1
timestamp 1699707026
transform 1 0 1595 0 1 4586
box -263 -787 263 769
use sky130_fd_pr__pfet_01v8_UJKTUG  sky130_fd_pr__pfet_01v8_UJKTUG_0
timestamp 1699600097
transform 1 0 1307 0 1 4586
box -359 -787 359 769
use sky130_fd_pr__pfet_01v8_UJKTUG  sky130_fd_pr__pfet_01v8_UJKTUG_1
timestamp 1699600097
transform 1 0 1307 0 -1 1066
box -359 -787 359 769
<< labels >>
flabel metal1 1292 1862 1320 1901 0 FreeSans 320 0 0 0 vin
port 16 nsew
flabel locali 995 2819 1026 2838 0 FreeSans 320 0 0 0 VSS
port 35 nsew
flabel metal4 372 2724 509 2933 0 FreeSans 640 0 0 0 VDD
port 24 nsew
flabel metal1 1293 3796 1316 3825 0 FreeSans 320 0 0 0 vip
port 3 nsew
flabel metal5 41990 5874 42264 6088 0 FreeSans 1600 0 0 0 tah_vp
port 37 nsew
flabel metal5 42026 -392 42274 -192 0 FreeSans 1600 0 0 0 tah_vn
port 39 nsew
flabel via1 53595 7057 53647 7109 0 FreeSans 320 0 0 0 sw
port 42 nsew
flabel via1 53498 6027 53550 6079 0 FreeSans 320 0 0 0 sw_n
port 44 nsew
flabel metal2 1939 1839 1973 3815 0 FreeSans 320 0 0 0 sw
flabel metal2 1830 1973 1864 3675 0 FreeSans 320 0 0 0 sw_n
<< end >>
