magic
tech sky130A
magscale 1 2
timestamp 1697713470
<< nmos >>
rect -205 -138 205 138
<< ndiff >>
rect -263 126 -205 138
rect -263 -126 -251 126
rect -217 -126 -205 126
rect -263 -138 -205 -126
rect 205 126 263 138
rect 205 -126 217 126
rect 251 -126 263 126
rect 205 -138 263 -126
<< ndiffc >>
rect -251 -126 -217 126
rect 217 -126 251 126
<< poly >>
rect -205 138 205 164
rect -205 -164 205 -138
<< locali >>
rect -251 126 -217 142
rect -251 -142 -217 -126
rect 217 126 251 142
rect 217 -142 251 -126
<< properties >>
string FIXED_BBOX -348 -295 348 295
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.375 l 2.045 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
