magic
tech sky130A
magscale 1 2
timestamp 1698614885
use hgu_inverter  x1[0]
timestamp 1698608947
transform 1 0 53 0 1 2200
box 372 160 690 825
use hgu_inverter  x1[1]
timestamp 1698608947
transform -1 0 1203 0 1 2200
box 372 160 690 825
use hgu_inverter  x1[2]
timestamp 1698608947
transform 1 0 229 0 1 2200
box 372 160 690 825
use hgu_inverter  x1[3]
timestamp 1698608947
transform -1 0 1379 0 1 2200
box 372 160 690 825
use hgu_inverter  x1[4]
timestamp 1698608947
transform 1 0 405 0 1 2200
box 372 160 690 825
use hgu_inverter  x1[5]
timestamp 1698608947
transform -1 0 1555 0 1 2200
box 372 160 690 825
use hgu_inverter  x1[6]
timestamp 1698608947
transform 1 0 581 0 1 2200
box 372 160 690 825
use hgu_inverter  x1[7]
timestamp 1698608947
transform -1 0 1731 0 1 2200
box 372 160 690 825
<< end >>
