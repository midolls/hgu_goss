* NGSPICE file created from hgu_delay_flat.ext - technology: sky130A

.subckt hgu_delay_flat out sample_delay_offset in sample_code2[3] sample_code3[3]
+ sample_code1[1] sample_code1[0] sample_code3[0] sample_code3[1] sample_code3[2]
+ sample_code2[1] sample_code2[2] sample_code1[2] sample_code0[2] sample_code0[1]
+ sample_code0[0] sample_code0[3] sample_code1[3] sample_code2[0] VSS VDD
X0 x2.x6.SW sample_delay_offset.t0 VDD.t49 VDD.t48 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1 VSS.t47 x3.IN a_6749_n1239# VDD.t37 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2 a_7436_1812# x1.IN a_7364_1812# VSS.t15 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 x2.x9.output_stack x2.x10.Y.t2 x2.x5[7].floating.t7 VDD.t53 sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X4 a_6465_2476# x4.x9.output_stack x1.IN VDD.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.122 ps=1.42 w=0.42 l=0.15
X5 a_727_1536# in.t0 a_655_1674# VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 a_655_1122# in.t1 a_567_1122# VSS.t4 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X7 x1.x9.output_stack sample_code1[1].t0 x1.x3[1].floating VSS.t32 sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X8 a_7389_3063# x1.IN a_7301_2925# VDD.t17 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X9 a_6058_n161# x3.IN a_5970_n161# VSS.t42 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X10 VDD.t76 sample_code2[3].t0 x2.x10.Y.t1 VDD.t75 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X11 a_12767_n299# x2.IN a_12679_n437# VSS.t24 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X12 VSS.t63 sample_delay_offset.t1 x4.x6.SW VSS.t62 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X13 x4.x9.output_stack x4.x10.Y.t2 x4.x5[7].floating.t7 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X14 a_12839_n851# x2.IN a_12767_n713# VSS.t25 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X15 a_7389_3339# x1.IN a_7301_3201# VDD.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X16 x2.x3[1].floating sample_code2[1].t0 x2.x9.output_stack VSS.t81 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X17 x3.x4[3].floating sample_code3[2].t0 x3.x9.output_stack VSS.t77 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X18 a_6058_n437# x3.IN a_5970_n437# VSS.t42 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X19 a_6465_2135# x1.IN VDD.t15 VSS.t20 sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X20 a_6749_n1036# x3.IN VDD.t36 VSS.t46 sky130_fd_pr__nfet_01v8 ad=0.0651 pd=0.73 as=0.0693 ps=0.75 w=0.42 l=0.15
X21 x4.x9.output_stack sample_delay_offset.t2 x4.x7.floating VSS.t61 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X22 out.t1 x3.x9.output_stack a_40_n1239# VDD.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.0651 ps=0.73 w=0.42 l=0.15
X23 x3.x4[3].floating sample_code3[2].t1 x3.x9.output_stack VSS.t51 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X24 a_7436_1260# x1.IN a_7364_1398# VSS.t15 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X25 x1.x9.output_stack sample_delay_offset.t3 x1.x7.floating VSS.t60 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X26 a_6105_n2378# x3.IN VDD.t35 VDD.t32 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X27 a_680_3063# in.t2 a_592_3201# VDD.t57 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X28 x1.x9.output_stack x1.x10.Y.t2 x1.x5[7].floating.t7 VDD.t21 sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X29 x4.x3[1].floating sample_code0[1].t0 x4.x9.output_stack VSS.t38 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X30 VDD.t27 x2.IN a_13174_2135# VSS.t29 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0651 ps=0.73 w=0.42 l=0.15
X31 x3.x9.output_stack x3.x10.Y.t2 x3.x5[7].floating.t7 VDD.t2 sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X32 x1.x5[7].floating.t6 x1.x10.Y.t3 x1.x9.output_stack VDD.t21 sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X33 x4.x9.output_stack sample_code0[1].t1 x4.x3[1].floating VSS.t79 sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X34 a_7364_2088# x1.IN a_7276_1950# VSS.t14 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X35 a_655_1812# in.t3 a_567_1674# VSS.t4 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X36 a_6058_n851# x3.IN x3.x9.output_stack VSS.t42 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X37 a_12839_n299# x2.IN a_12767_n299# VSS.t25 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X38 x1.x5[7].floating.t5 x1.x10.Y.t4 x1.x9.output_stack VDD.t21 sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X39 x1.x9.output_stack x1.IN a_7301_2925# VDD.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X40 a_727_1260# in.t4 a_655_1260# VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X41 x3.x6.floating x3.x6.SW x3.x9.output_stack VDD.t56 sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X42 a_13174_2476# x2.IN VSS.t28 VDD.t26 sky130_fd_pr__pfet_01v8_hvt ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X43 a_727_1536# in.t5 a_655_1536# VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X44 x3.x9.output_stack sample_code3[2].t2 x3.x4[3].floating VSS.t70 sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X45 x4.x10.Y.t0 sample_code0[3].t0 VSS.t65 VSS.t64 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X46 x2.x9.output_stack x2.x10.Y.t3 x2.x5[7].floating.t6 VDD.t65 sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X47 x3.x5[7].floating.t6 x3.x10.Y.t3 x3.x9.output_stack VDD.t64 sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X48 a_6130_n575# x3.IN a_6058_n575# VSS.t41 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X49 a_6105_n2102# x3.IN a_6017_n1964# VDD.t32 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X50 x3.x9.output_stack sample_code3[2].t3 x3.x4[3].floating VSS.t10 sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X51 x1.x10.Y.t1 sample_code1[3].t0 VDD.t51 VDD.t50 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X52 a_655_1398# in.t6 a_567_1398# VSS.t4 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X53 x3.x6.SW sample_delay_offset.t4 VSS.t59 VSS.t58 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X54 x3.x5[7].floating.t5 x3.x10.Y.t4 x3.x9.output_stack VDD.t41 sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X55 VDD.t13 x1.IN a_6465_2135# VSS.t19 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0651 ps=0.73 w=0.42 l=0.15
X56 x3.x5[7].floating.t4 x3.x10.Y.t5 x3.x9.output_stack VDD.t69 sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X57 x3.IN x2.x9.output_stack a_6749_n1036# VSS.t34 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0651 ps=0.73 w=0.42 l=0.15
X58 a_7364_1674# x1.IN a_7276_1674# VSS.t14 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X59 x4.x9.output_stack sample_code0[2].t0 x4.x4[3].floating VSS.t1 sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X60 x1.x9.output_stack x1.IN a_7364_2088# VSS.t15 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X61 x4.x5[7].floating.t6 x4.x10.Y.t3 x4.x9.output_stack VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X62 a_6465_2476# x1.IN VSS.t18 VDD.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X63 a_727_1812# in.t7 a_655_1950# VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X64 VDD.t30 x2.x9.output_stack a_6749_n1239# VDD.t29 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X65 a_6749_n1239# x3.IN VSS.t45 VDD.t34 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.0693 ps=0.75 w=0.42 l=0.15
X66 x3.x5[7].floating.t3 x3.x10.Y.t6 x3.x9.output_stack VDD.t73 sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X67 VSS.t76 sample_code3[3].t0 x3.x10.Y.t1 VSS.t75 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X68 x1.x9.output_stack sample_code1[2].t0 x1.x4[3].floating VSS.t7 sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X69 a_12814_n2102# x2.IN a_12726_n2240# VDD.t23 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X70 a_6105_n2378# x3.IN a_6017_n2240# VDD.t32 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X71 a_12767_n575# x2.IN a_12679_n713# VSS.t24 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X72 VDD.t12 x1.IN a_7301_3477# VDD.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X73 x2.x4[3].floating sample_code2[2].t0 x2.x9.output_stack VSS.t67 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X74 a_6058_n713# x3.IN a_5970_n713# VSS.t42 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X75 VSS.t3 in.t8 a_655_1122# VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X76 x1.x5[7].floating.t4 x1.x10.Y.t5 x1.x9.output_stack VDD.t21 sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X77 a_680_3339# in.t9 a_592_3477# VDD.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X78 a_13174_2476# x1.x9.output_stack VDD.t63 VDD.t62 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X79 VSS.t27 x2.IN a_13174_2476# VDD.t26 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0651 ps=0.73 w=0.42 l=0.15
X80 a_12814_n1826# x2.IN x2.x9.output_stack VDD.t23 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X81 x2.x4[3].floating sample_code2[2].t1 x2.x9.output_stack VSS.t83 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X82 a_6130_n299# x3.IN a_6058_n161# VSS.t41 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X83 x1.x4[3].floating sample_code1[2].t1 x1.x9.output_stack VSS.t80 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X84 VDD.t47 sample_delay_offset.t5 x1.x6.SW VDD.t46 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X85 x4.x9.output_stack x4.x10.Y.t4 x4.x5[7].floating.t5 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X86 a_7436_1536# x1.IN a_7364_1674# VSS.t15 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X87 a_6130_n23# x3.IN a_6058_n23# VSS.t41 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X88 a_6130_n575# x3.IN a_6058_n437# VSS.t41 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X89 x2.x7.floating sample_delay_offset.t6 x2.x9.output_stack VSS.t57 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X90 x3.x9.output_stack sample_code3[0].t0 x3.x2.floating VSS.t33 sky130_fd_pr__nfet_01v8 ad=0.124 pd=1.43 as=0.122 ps=1.42 w=0.42 l=0.15
X91 a_655_2088# in.t10 a_567_1950# VSS.t4 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X92 a_7364_1260# x1.IN a_7276_1122# VSS.t14 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X93 a_12839_n23# x2.IN a_12767_n23# VSS.t25 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X94 a_6105_n1826# x3.IN a_6017_n1964# VDD.t32 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X95 a_12839_n575# x2.IN a_12767_n575# VSS.t25 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X96 a_7364_1536# x1.IN a_7276_1398# VSS.t14 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X97 VDD.t39 out.t2 a_40_n1036# VSS.t48 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X98 a_6058_n299# x3.IN a_5970_n437# VSS.t42 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X99 x1.x9.output_stack x1.x10.Y.t6 x1.x5[7].floating.t3 VDD.t21 sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X100 a_40_n1036# out.t3 VDD.t52 VSS.t66 sky130_fd_pr__nfet_01v8 ad=0.0651 pd=0.73 as=0.0693 ps=0.75 w=0.42 l=0.15
X101 x1.x9.output_stack x1.x10.Y.t7 x1.x5[7].floating.t2 VDD.t21 sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X102 a_6130_n23# x3.IN a_6058_115# VSS.t41 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X103 x3.x3[1].floating sample_code3[1].t0 x3.x9.output_stack VSS.t71 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X104 x4.x5[7].floating.t4 x4.x10.Y.t5 x4.x9.output_stack VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X105 a_727_1812# in.t11 a_655_1812# VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X106 a_12767_n161# x2.IN a_12679_n161# VSS.t24 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X107 a_6465_2476# x4.x9.output_stack VDD.t19 VDD.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X108 VSS.t17 x1.IN a_6465_2476# VDD.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0651 ps=0.73 w=0.42 l=0.15
X109 x2.x6.floating x2.x6.SW x2.x9.output_stack VDD.t31 sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X110 x3.IN x2.x9.output_stack a_6749_n1239# VDD.t29 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.0651 ps=0.73 w=0.42 l=0.15
X111 a_12839_n23# x2.IN a_12767_115# VSS.t25 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X112 x2.x9.output_stack sample_code2[2].t2 x2.x4[3].floating VSS.t49 sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X113 x2.x9.output_stack sample_code2[0].t0 x2.x2.floating VSS.t31 sky130_fd_pr__nfet_01v8 ad=0.124 pd=1.43 as=0.122 ps=1.42 w=0.42 l=0.15
X114 a_7389_3063# x1.IN a_7301_3201# VDD.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X115 x4.x4[3].floating sample_code0[2].t1 x4.x9.output_stack VSS.t36 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X116 x2.x5[7].floating.t5 x2.x10.Y.t4 x2.x9.output_stack VDD.t72 sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X117 x3.x9.output_stack x3.x10.Y.t7 x3.x5[7].floating.t2 VDD.t68 sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X118 a_6130_n851# x3.IN a_6058_n851# VSS.t41 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X119 x1.x10.Y.t0 sample_code1[3].t1 VSS.t6 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X120 a_12767_n437# x2.IN a_12679_n437# VSS.t24 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X121 a_680_3063# in.t12 a_592_2925# VDD.t40 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X122 a_13174_2135# x1.x9.output_stack x2.IN VSS.t73 sky130_fd_pr__nfet_01v8 ad=0.0651 pd=0.73 as=0.122 ps=1.42 w=0.42 l=0.15
X123 x3.x6.SW sample_delay_offset.t7 VDD.t45 VDD.t44 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X124 a_655_1674# in.t13 a_567_1674# VSS.t4 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X125 x2.x5[7].floating.t4 x2.x10.Y.t5 x2.x9.output_stack VDD.t20 sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X126 a_7436_1260# x1.IN a_7364_1260# VSS.t15 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X127 x2.x5[7].floating.t3 x2.x10.Y.t6 x2.x9.output_stack VDD.t28 sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X128 x3.x9.output_stack x3.x10.Y.t8 x3.x5[7].floating.t1 VDD.t74 sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X129 x1.x9.output_stack x1.x6.SW x1.x6.floating VDD.t22 sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X130 a_7364_1950# x1.IN a_7276_1950# VSS.t14 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X131 a_12814_n2378# x2.IN VDD.t25 VDD.t23 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X132 a_680_3339# in.t14 a_592_3201# VDD.t71 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X133 x1.x2.floating sample_code1[0].t0 x1.x9.output_stack VSS.t82 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.124 ps=1.43 w=0.42 l=0.15
X134 a_7436_1536# x1.IN a_7364_1536# VSS.t15 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X135 x2.x6.SW sample_delay_offset.t8 VSS.t56 VSS.t55 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X136 x2.x5[7].floating.t2 x2.x10.Y.t7 x2.x9.output_stack VDD.t66 sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X137 a_12767_n23# x2.IN a_12679_n161# VSS.t24 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X138 x3.x9.output_stack x3.x10.Y.t9 x3.x5[7].floating.t0 VDD.t70 sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X139 x1.x3[1].floating sample_code1[1].t1 x1.x9.output_stack VSS.t30 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X140 a_6058_n23# x3.IN a_5970_n161# VSS.t42 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X141 VDD.t59 sample_code3[3].t1 x3.x10.Y.t0 VDD.t58 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X142 a_727_1260# in.t15 a_655_1398# VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X143 a_7364_1122# x1.IN a_7276_1122# VSS.t14 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X144 a_12767_n851# x2.IN x2.x9.output_stack VSS.t24 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X145 a_12839_n299# x2.IN a_12767_n161# VSS.t25 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X146 VSS.t13 x3.x9.output_stack a_40_n1036# VSS.t12 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X147 x4.x5[7].floating.t3 x4.x10.Y.t6 x4.x9.output_stack VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X148 VSS.t40 sample_code2[3].t1 x2.x10.Y.t0 VSS.t39 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X149 x2.x9.output_stack sample_code2[2].t3 x2.x4[3].floating VSS.t78 sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X150 VDD.t33 x3.IN a_6749_n1036# VSS.t44 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X151 x3.x9.output_stack sample_code3[1].t1 x3.x3[1].floating VSS.t68 sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X152 a_12839_n575# x2.IN a_12767_n437# VSS.t25 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X153 VSS.t54 sample_delay_offset.t9 x1.x6.SW VSS.t53 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X154 x3.x7.floating sample_delay_offset.t10 x3.x9.output_stack VSS.t52 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X155 a_6465_2135# x4.x9.output_stack x1.IN VSS.t21 sky130_fd_pr__nfet_01v8 ad=0.0651 pd=0.73 as=0.122 ps=1.42 w=0.42 l=0.15
X156 a_12767_115# x2.IN VSS.t26 VSS.t24 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X157 x1.x4[3].floating sample_code1[2].t2 x1.x9.output_stack VSS.t72 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X158 VDD.t43 sample_delay_offset.t11 x4.x6.SW VDD.t42 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X159 a_6058_115# x3.IN VSS.t43 VSS.t42 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X160 a_12814_n2102# x2.IN a_12726_n1964# VDD.t23 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X161 x4.x9.output_stack in.t16 a_592_2925# VDD.t77 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X162 a_7436_1812# x1.IN a_7364_1950# VSS.t15 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X163 x1.x9.output_stack sample_code1[2].t3 x1.x4[3].floating VSS.t37 sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X164 VSS.t11 out.t4 a_40_n1239# VDD.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X165 x4.x2.floating sample_code0[0].t0 x4.x9.output_stack VSS.t69 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.124 ps=1.43 w=0.42 l=0.15
X166 VSS.t35 x2.x9.output_stack a_6749_n1036# VSS.t34 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X167 x1.x5[7].floating.t1 x1.x10.Y.t8 x1.x9.output_stack VDD.t21 sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X168 a_40_n1239# out.t5 VSS.t8 VDD.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.0693 ps=0.75 w=0.42 l=0.15
X169 a_6130_n851# x3.IN a_6058_n713# VSS.t41 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X170 a_655_1260# in.t17 a_567_1122# VSS.t4 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X171 x4.x9.output_stack x4.x10.Y.t7 x4.x5[7].floating.t2 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X172 a_13174_2135# x1.x9.output_stack VSS.t74 VSS.t73 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X173 x4.x9.output_stack x4.x6.SW x4.x6.floating VDD.t7 sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X174 a_655_1536# in.t18 a_567_1398# VSS.t4 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X175 out.t0 x3.x9.output_stack a_40_n1036# VSS.t12 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0651 ps=0.73 w=0.42 l=0.15
X176 a_7364_1812# x1.IN a_7276_1674# VSS.t14 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X177 VSS.t16 x1.IN a_7364_1122# VSS.t15 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X178 a_12814_n2378# x2.IN a_12726_n2240# VDD.t23 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X179 a_12839_n851# x2.IN a_12767_n851# VSS.t25 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X180 a_6058_n575# x3.IN a_5970_n713# VSS.t42 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X181 a_7389_3339# x1.IN a_7301_3477# VDD.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X182 a_13174_2476# x1.x9.output_stack x2.IN VDD.t26 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.122 ps=1.42 w=0.42 l=0.15
X183 a_6105_n2102# x3.IN a_6017_n2240# VDD.t32 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X184 x4.x9.output_stack in.t19 a_655_2088# VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X185 VDD.t6 x3.x9.output_stack a_40_n1239# VDD.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X186 x2.x9.output_stack sample_code2[1].t1 x2.x3[1].floating VSS.t9 sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X187 x1.x9.output_stack x1.x10.Y.t9 x1.x5[7].floating.t0 VDD.t21 sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X188 a_12767_n713# x2.IN a_12679_n713# VSS.t24 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X189 x4.x9.output_stack sample_code0[2].t2 x4.x4[3].floating VSS.t50 sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X190 a_6130_n299# x3.IN a_6058_n299# VSS.t41 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X191 x4.x9.output_stack x4.x10.Y.t8 x4.x5[7].floating.t1 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X192 x4.x5[7].floating.t0 x4.x10.Y.t9 x4.x9.output_stack VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X193 a_13174_2135# x2.IN VDD.t24 VSS.t23 sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X194 x4.x10.Y.t1 sample_code0[3].t1 VDD.t55 VDD.t54 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X195 a_655_1950# in.t20 a_567_1950# VSS.t4 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X196 x2.x9.output_stack x2.x10.Y.t8 x2.x5[7].floating.t1 VDD.t67 sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X197 a_6105_n1826# x3.IN x3.x9.output_stack VDD.t32 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X198 x2.x9.output_stack x2.x10.Y.t9 x2.x5[7].floating.t0 VDD.t38 sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X199 x4.x4[3].floating sample_code0[2].t3 x4.x9.output_stack VSS.t2 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X200 VDD.t61 in.t21 a_592_3477# VDD.t60 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X201 a_6465_2135# x4.x9.output_stack VSS.t22 VSS.t21 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X202 a_7364_1398# x1.IN a_7276_1398# VSS.t14 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X203 a_12814_n1826# x2.IN a_12726_n1964# VDD.t23 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
R0 sample_delay_offset.n30 sample_delay_offset.t11 230.016
R1 sample_delay_offset.n2 sample_delay_offset.t5 230.016
R2 sample_delay_offset.n18 sample_delay_offset.t7 229.971
R3 sample_delay_offset.n7 sample_delay_offset.t0 229.971
R4 sample_delay_offset.n18 sample_delay_offset.t4 158.351
R5 sample_delay_offset.n7 sample_delay_offset.t8 158.351
R6 sample_delay_offset.n29 sample_delay_offset.t1 153.665
R7 sample_delay_offset.n1 sample_delay_offset.t9 153.665
R8 sample_delay_offset.n30 sample_delay_offset 153.601
R9 sample_delay_offset.n2 sample_delay_offset 153.601
R10 sample_delay_offset sample_delay_offset.t2 140.379
R11 sample_delay_offset sample_delay_offset.t3 140.379
R12 sample_delay_offset.n26 sample_delay_offset.t10 140.34
R13 sample_delay_offset.n15 sample_delay_offset.t6 140.34
R14 sample_delay_offset.n31 sample_delay_offset.n30 9.3005
R15 sample_delay_offset.n3 sample_delay_offset.n2 9.3005
R16 sample_delay_offset.n38 sample_delay_offset.n16 9.14466
R17 sample_delay_offset.n19 sample_delay_offset.n18 7.39809
R18 sample_delay_offset.n8 sample_delay_offset.n7 7.39809
R19 sample_delay_offset.n36 sample_delay_offset.n35 5.90325
R20 sample_delay_offset.n37 sample_delay_offset.n36 5.46925
R21 sample_delay_offset.n30 sample_delay_offset.n29 4.91671
R22 sample_delay_offset.n2 sample_delay_offset.n1 4.91671
R23 sample_delay_offset.n5 sample_delay_offset.n3 4.90192
R24 sample_delay_offset.n33 sample_delay_offset.n31 4.9013
R25 sample_delay_offset.n27 sample_delay_offset.n26 4.18104
R26 sample_delay_offset.n16 sample_delay_offset.n15 4.18104
R27 sample_delay_offset.n35 sample_delay_offset 4.14309
R28 sample_delay_offset.n39 sample_delay_offset 4.14309
R29 sample_delay_offset.n21 sample_delay_offset.n20 4.0005
R30 sample_delay_offset.n10 sample_delay_offset.n9 4.0005
R31 sample_delay_offset.n39 sample_delay_offset.n38 3.76287
R32 sample_delay_offset.n37 sample_delay_offset.n27 3.75602
R33 sample_delay_offset.n22 sample_delay_offset.n21 3.03311
R34 sample_delay_offset.n11 sample_delay_offset.n10 3.03311
R35 sample_delay_offset sample_delay_offset.n28 2.4005
R36 sample_delay_offset sample_delay_offset.n0 2.4005
R37 sample_delay_offset.n38 sample_delay_offset.n37 2.01947
R38 sample_delay_offset.n25 sample_delay_offset.n24 1.87694
R39 sample_delay_offset.n14 sample_delay_offset.n13 1.87694
R40 sample_delay_offset.n20 sample_delay_offset 1.6005
R41 sample_delay_offset.n9 sample_delay_offset 1.6005
R42 sample_delay_offset.n25 sample_delay_offset 1.43349
R43 sample_delay_offset.n14 sample_delay_offset 1.43349
R44 sample_delay_offset.n24 sample_delay_offset.n23 1.12626
R45 sample_delay_offset.n13 sample_delay_offset.n12 1.12626
R46 sample_delay_offset.n34 sample_delay_offset 1.01229
R47 sample_delay_offset sample_delay_offset.n40 1.01229
R48 sample_delay_offset.n34 sample_delay_offset.n33 0.726043
R49 sample_delay_offset.n27 sample_delay_offset.n25 0.726043
R50 sample_delay_offset.n16 sample_delay_offset.n14 0.726043
R51 sample_delay_offset.n40 sample_delay_offset.n5 0.726043
R52 sample_delay_offset.n36 sample_delay_offset 0.718134
R53 sample_delay_offset.n31 sample_delay_offset.n28 0.533833
R54 sample_delay_offset.n21 sample_delay_offset.n19 0.533833
R55 sample_delay_offset.n10 sample_delay_offset.n8 0.533833
R56 sample_delay_offset.n3 sample_delay_offset.n0 0.533833
R57 sample_delay_offset.n33 sample_delay_offset.n32 0.421696
R58 sample_delay_offset.n5 sample_delay_offset.n4 0.421696
R59 sample_delay_offset.n35 sample_delay_offset.n34 0.0783302
R60 sample_delay_offset.n40 sample_delay_offset.n39 0.0783302
R61 sample_delay_offset.n27 sample_delay_offset 0.0447308
R62 sample_delay_offset.n16 sample_delay_offset 0.0447308
R63 sample_delay_offset.n26 sample_delay_offset 0.0384464
R64 sample_delay_offset.n15 sample_delay_offset 0.0384464
R65 sample_delay_offset.n32 sample_delay_offset 0.0195217
R66 sample_delay_offset.n27 sample_delay_offset 0.0195217
R67 sample_delay_offset.n16 sample_delay_offset 0.0195217
R68 sample_delay_offset.n4 sample_delay_offset 0.0195217
R69 sample_delay_offset.n22 sample_delay_offset.n17 0.0179598
R70 sample_delay_offset.n11 sample_delay_offset.n6 0.0179598
R71 sample_delay_offset.n32 sample_delay_offset 0.0170094
R72 sample_delay_offset.n4 sample_delay_offset 0.0170094
R73 sample_delay_offset.n23 sample_delay_offset.n22 0.00504545
R74 sample_delay_offset.n12 sample_delay_offset.n11 0.00504545
R75 VDD.n2595 VDD.n2564 76633.3
R76 VDD.n4990 VDD.n641 3782.21
R77 VDD.n2540 VDD.t37 1820.83
R78 VDD.t4 VDD.n3823 1820.83
R79 VDD.n6147 VDD.n12 1116.08
R80 VDD.n6095 VDD.n606 426
R81 VDD.n2621 VDD.n2455 423
R82 VDD.n4966 VDD.n4932 423
R83 VDD.n2599 VDD.n2485 354
R84 VDD.n4970 VDD.n1238 354
R85 VDD.n6128 VDD.n604 351
R86 VDD.n7273 VDD.t42 258.856
R87 VDD.n4967 VDD.t48 256.267
R88 VDD.n6159 VDD 242.981
R89 VDD VDD.t23 237.195
R90 VDD.n2539 VDD.n2538 198.234
R91 VDD.n1393 VDD.n1379 198.234
R92 VDD.n3822 VDD.n3821 198.234
R93 VDD.n2759 VDD.n2758 198.234
R94 VDD.n6842 VDD.n6841 198.118
R95 VDD.n6616 VDD.n6615 198.118
R96 VDD.n6390 VDD.n6389 198.118
R97 VDD.n7225 VDD.n7224 198.118
R98 VDD.n6075 VDD.n6074 198.118
R99 VDD.n5706 VDD.n5705 198.118
R100 VDD.n5478 VDD.n5477 198.118
R101 VDD.n5250 VDD.n5249 198.118
R102 VDD.n6392 VDD.n6391 198.118
R103 VDD.n6618 VDD.n6617 198.118
R104 VDD.n6844 VDD.n6843 198.118
R105 VDD.n4969 VDD.t75 191.554
R106 VDD.n7271 VDD.t54 188.965
R107 VDD.n2755 VDD.n2753 185
R108 VDD.n2772 VDD.n2755 185
R109 VDD.n4317 VDD.n4316 185
R110 VDD.n4318 VDD.n4317 185
R111 VDD.n2826 VDD.n2825 185
R112 VDD.n2825 VDD.n2824 185
R113 VDD.n2816 VDD.n2814 185
R114 VDD.n2836 VDD.n2816 185
R115 VDD.n2839 VDD.n2817 185
R116 VDD.n4292 VDD.n2817 185
R117 VDD.n4273 VDD.n4272 185
R118 VDD.n4274 VDD.n4273 185
R119 VDD.n2923 VDD.n2922 185
R120 VDD.n2924 VDD.n2923 185
R121 VDD.n2913 VDD.n2911 185
R122 VDD.n4254 VDD.n2913 185
R123 VDD.n2966 VDD.n2965 185
R124 VDD.n2967 VDD.n2966 185
R125 VDD.n2956 VDD.n2954 185
R126 VDD.n4233 VDD.n2956 185
R127 VDD.n3012 VDD.n3011 185
R128 VDD.n3013 VDD.n3012 185
R129 VDD.n4206 VDD.n4205 185
R130 VDD.n4207 VDD.n4206 185
R131 VDD.n3068 VDD.n3067 185
R132 VDD.n3067 VDD.n3066 185
R133 VDD.n3058 VDD.n3056 185
R134 VDD.n3078 VDD.n3058 185
R135 VDD.n4179 VDD.n4178 185
R136 VDD.n4180 VDD.n4179 185
R137 VDD.n3132 VDD.n3131 185
R138 VDD.n3131 VDD.n3130 185
R139 VDD.n4154 VDD.n4153 185
R140 VDD.n4155 VDD.n4154 185
R141 VDD.n3189 VDD.n3188 185
R142 VDD.n3190 VDD.n3189 185
R143 VDD.n3179 VDD.n3177 185
R144 VDD.n4135 VDD.n3179 185
R145 VDD.n3232 VDD.n3231 185
R146 VDD.n3233 VDD.n3232 185
R147 VDD.n3222 VDD.n3220 185
R148 VDD.n4114 VDD.n3222 185
R149 VDD.n3278 VDD.n3277 185
R150 VDD.n3279 VDD.n3278 185
R151 VDD.n4087 VDD.n4086 185
R152 VDD.n4088 VDD.n4087 185
R153 VDD.n3334 VDD.n3333 185
R154 VDD.n3333 VDD.n3332 185
R155 VDD.n3324 VDD.n3322 185
R156 VDD.n3344 VDD.n3324 185
R157 VDD.n4060 VDD.n4059 185
R158 VDD.n4061 VDD.n4060 185
R159 VDD.n3398 VDD.n3397 185
R160 VDD.n3397 VDD.n3396 185
R161 VDD.n4035 VDD.n4034 185
R162 VDD.n4036 VDD.n4035 185
R163 VDD.n3455 VDD.n3454 185
R164 VDD.n3456 VDD.n3455 185
R165 VDD.n3445 VDD.n3443 185
R166 VDD.n4016 VDD.n3445 185
R167 VDD.n3498 VDD.n3497 185
R168 VDD.n3499 VDD.n3498 185
R169 VDD.n3488 VDD.n3486 185
R170 VDD.n3995 VDD.n3488 185
R171 VDD.n3544 VDD.n3543 185
R172 VDD.n3545 VDD.n3544 185
R173 VDD.n3968 VDD.n3967 185
R174 VDD.n3969 VDD.n3968 185
R175 VDD.n3600 VDD.n3599 185
R176 VDD.n3599 VDD.n3598 185
R177 VDD.n3590 VDD.n3588 185
R178 VDD.n3610 VDD.n3590 185
R179 VDD.n3941 VDD.n3940 185
R180 VDD.n3942 VDD.n3941 185
R181 VDD.n3664 VDD.n3663 185
R182 VDD.n3663 VDD.n3662 185
R183 VDD.n3916 VDD.n3915 185
R184 VDD.n3917 VDD.n3916 185
R185 VDD.n3721 VDD.n3720 185
R186 VDD.n3722 VDD.n3721 185
R187 VDD.n3711 VDD.n3709 185
R188 VDD.n3897 VDD.n3711 185
R189 VDD.n3764 VDD.n3763 185
R190 VDD.n3765 VDD.n3764 185
R191 VDD.n3754 VDD.n3752 185
R192 VDD.n3876 VDD.n3754 185
R193 VDD.n3874 VDD.n3873 185
R194 VDD.n3875 VDD.n3874 185
R195 VDD.n3762 VDD.n3753 185
R196 VDD.n3766 VDD.n3753 185
R197 VDD.n3895 VDD.n3894 185
R198 VDD.n3896 VDD.n3895 185
R199 VDD.n3719 VDD.n3710 185
R200 VDD.n3723 VDD.n3710 185
R201 VDD.n3819 VDD.n3818 185
R202 VDD.n3658 VDD.n3657 185
R203 VDD.n3918 VDD.n3658 185
R204 VDD.n3613 VDD.n3591 185
R205 VDD.n3943 VDD.n3591 185
R206 VDD.n3608 VDD.n3607 185
R207 VDD.n3609 VDD.n3608 185
R208 VDD.n3596 VDD.n3595 185
R209 VDD.n3597 VDD.n3596 185
R210 VDD.n3549 VDD.n3535 185
R211 VDD.n3970 VDD.n3535 185
R212 VDD.n3665 VDD.n3660 185
R213 VDD.n3660 VDD.n3659 185
R214 VDD.n3534 VDD.n3532 185
R215 VDD.n3546 VDD.n3534 185
R216 VDD.n3993 VDD.n3992 185
R217 VDD.n3994 VDD.n3993 185
R218 VDD.n3496 VDD.n3487 185
R219 VDD.n3500 VDD.n3487 185
R220 VDD.n4014 VDD.n4013 185
R221 VDD.n4015 VDD.n4014 185
R222 VDD.n3453 VDD.n3444 185
R223 VDD.n3457 VDD.n3444 185
R224 VDD.n3542 VDD.n3541 185
R225 VDD.n3541 VDD.n3540 185
R226 VDD.n3538 VDD.n3537 185
R227 VDD.n3539 VDD.n3538 185
R228 VDD.n3392 VDD.n3391 185
R229 VDD.n4037 VDD.n3392 185
R230 VDD.n3347 VDD.n3325 185
R231 VDD.n4062 VDD.n3325 185
R232 VDD.n3342 VDD.n3341 185
R233 VDD.n3343 VDD.n3342 185
R234 VDD.n3330 VDD.n3329 185
R235 VDD.n3331 VDD.n3330 185
R236 VDD.n3283 VDD.n3269 185
R237 VDD.n4089 VDD.n3269 185
R238 VDD.n3399 VDD.n3394 185
R239 VDD.n3394 VDD.n3393 185
R240 VDD.n3268 VDD.n3266 185
R241 VDD.n3280 VDD.n3268 185
R242 VDD.n4112 VDD.n4111 185
R243 VDD.n4113 VDD.n4112 185
R244 VDD.n3230 VDD.n3221 185
R245 VDD.n3234 VDD.n3221 185
R246 VDD.n4133 VDD.n4132 185
R247 VDD.n4134 VDD.n4133 185
R248 VDD.n3187 VDD.n3178 185
R249 VDD.n3191 VDD.n3178 185
R250 VDD.n3276 VDD.n3275 185
R251 VDD.n3275 VDD.n3274 185
R252 VDD.n3272 VDD.n3271 185
R253 VDD.n3273 VDD.n3272 185
R254 VDD.n3126 VDD.n3125 185
R255 VDD.n4156 VDD.n3126 185
R256 VDD.n3081 VDD.n3059 185
R257 VDD.n4181 VDD.n3059 185
R258 VDD.n3076 VDD.n3075 185
R259 VDD.n3077 VDD.n3076 185
R260 VDD.n3064 VDD.n3063 185
R261 VDD.n3065 VDD.n3064 185
R262 VDD.n3017 VDD.n3003 185
R263 VDD.n4208 VDD.n3003 185
R264 VDD.n3133 VDD.n3128 185
R265 VDD.n3128 VDD.n3127 185
R266 VDD.n3002 VDD.n3000 185
R267 VDD.n3014 VDD.n3002 185
R268 VDD.n4231 VDD.n4230 185
R269 VDD.n4232 VDD.n4231 185
R270 VDD.n2964 VDD.n2955 185
R271 VDD.n2968 VDD.n2955 185
R272 VDD.n4252 VDD.n4251 185
R273 VDD.n4253 VDD.n4252 185
R274 VDD.n2921 VDD.n2912 185
R275 VDD.n2925 VDD.n2912 185
R276 VDD.n3010 VDD.n3009 185
R277 VDD.n3009 VDD.n3008 185
R278 VDD.n3006 VDD.n3005 185
R279 VDD.n3007 VDD.n3006 185
R280 VDD.n2849 VDD.n2847 185
R281 VDD.n4275 VDD.n2849 185
R282 VDD.n2834 VDD.n2833 185
R283 VDD.n2835 VDD.n2834 185
R284 VDD.n2822 VDD.n2821 185
R285 VDD.n2823 VDD.n2822 185
R286 VDD.n2770 VDD.n2769 185
R287 VDD.n2771 VDD.n2770 185
R288 VDD.n2775 VDD.n2756 185
R289 VDD.n4319 VDD.n2756 185
R290 VDD.n4290 VDD.n4289 185
R291 VDD.n4291 VDD.n4290 185
R292 VDD.n2761 VDD.n2760 185
R293 VDD.n2454 VDD.n2453 185
R294 VDD.n2627 VDD.n2454 185
R295 VDD.n2639 VDD.n2638 185
R296 VDD.n2640 VDD.n2639 185
R297 VDD.n2644 VDD.n2448 185
R298 VDD.n4372 VDD.n2448 185
R299 VDD.n2696 VDD.n2695 185
R300 VDD.n2697 VDD.n2696 185
R301 VDD.n2708 VDD.n2707 185
R302 VDD.n2709 VDD.n2708 185
R303 VDD.n2713 VDD.n2691 185
R304 VDD.n4345 VDD.n2691 185
R305 VDD.n2630 VDD.n2629 185
R306 VDD.n2629 VDD.n2628 185
R307 VDD.n2447 VDD.n2445 185
R308 VDD.n2641 VDD.n2447 185
R309 VDD.n4370 VDD.n4369 185
R310 VDD.n4371 VDD.n4370 185
R311 VDD.n2700 VDD.n2699 185
R312 VDD.n2699 VDD.n2698 185
R313 VDD.n2690 VDD.n2688 185
R314 VDD.n2710 VDD.n2690 185
R315 VDD.n4343 VDD.n4342 185
R316 VDD.n4344 VDD.n4343 185
R317 VDD.n2600 VDD.n2599 185
R318 VDD.n2599 VDD.n2598 185
R319 VDD.n4868 VDD.n4867 185
R320 VDD.n4869 VDD.n4868 185
R321 VDD.n1452 VDD.n1451 185
R322 VDD.n1451 VDD.n1450 185
R323 VDD.n1442 VDD.n1440 185
R324 VDD.n1462 VDD.n1442 185
R325 VDD.n4841 VDD.n4840 185
R326 VDD.n4842 VDD.n4841 185
R327 VDD.n1516 VDD.n1515 185
R328 VDD.n1515 VDD.n1514 185
R329 VDD.n4816 VDD.n4815 185
R330 VDD.n4817 VDD.n4816 185
R331 VDD.n1572 VDD.n1571 185
R332 VDD.n1573 VDD.n1572 185
R333 VDD.n1561 VDD.n1559 185
R334 VDD.n4796 VDD.n1561 185
R335 VDD.n1614 VDD.n1613 185
R336 VDD.n1615 VDD.n1614 185
R337 VDD.n1603 VDD.n1601 185
R338 VDD.n4774 VDD.n1603 185
R339 VDD.n1660 VDD.n1659 185
R340 VDD.n1661 VDD.n1660 185
R341 VDD.n4747 VDD.n4746 185
R342 VDD.n4748 VDD.n4747 185
R343 VDD.n1716 VDD.n1715 185
R344 VDD.n1715 VDD.n1714 185
R345 VDD.n1706 VDD.n1704 185
R346 VDD.n1726 VDD.n1706 185
R347 VDD.n4720 VDD.n4719 185
R348 VDD.n4721 VDD.n4720 185
R349 VDD.n1780 VDD.n1779 185
R350 VDD.n1779 VDD.n1778 185
R351 VDD.n4695 VDD.n4694 185
R352 VDD.n4696 VDD.n4695 185
R353 VDD.n1836 VDD.n1835 185
R354 VDD.n1837 VDD.n1836 185
R355 VDD.n1825 VDD.n1823 185
R356 VDD.n4675 VDD.n1825 185
R357 VDD.n1878 VDD.n1877 185
R358 VDD.n1879 VDD.n1878 185
R359 VDD.n1867 VDD.n1865 185
R360 VDD.n4653 VDD.n1867 185
R361 VDD.n1924 VDD.n1923 185
R362 VDD.n1925 VDD.n1924 185
R363 VDD.n4626 VDD.n4625 185
R364 VDD.n4627 VDD.n4626 185
R365 VDD.n1980 VDD.n1979 185
R366 VDD.n1979 VDD.n1978 185
R367 VDD.n1970 VDD.n1968 185
R368 VDD.n1990 VDD.n1970 185
R369 VDD.n4599 VDD.n4598 185
R370 VDD.n4600 VDD.n4599 185
R371 VDD.n2044 VDD.n2043 185
R372 VDD.n2043 VDD.n2042 185
R373 VDD.n4574 VDD.n4573 185
R374 VDD.n4575 VDD.n4574 185
R375 VDD.n2100 VDD.n2099 185
R376 VDD.n2101 VDD.n2100 185
R377 VDD.n2089 VDD.n2087 185
R378 VDD.n4554 VDD.n2089 185
R379 VDD.n2142 VDD.n2141 185
R380 VDD.n2143 VDD.n2142 185
R381 VDD.n2131 VDD.n2129 185
R382 VDD.n4532 VDD.n2131 185
R383 VDD.n2188 VDD.n2187 185
R384 VDD.n2189 VDD.n2188 185
R385 VDD.n4505 VDD.n4504 185
R386 VDD.n4506 VDD.n4505 185
R387 VDD.n2244 VDD.n2243 185
R388 VDD.n2243 VDD.n2242 185
R389 VDD.n2234 VDD.n2232 185
R390 VDD.n2254 VDD.n2234 185
R391 VDD.n4478 VDD.n4477 185
R392 VDD.n4479 VDD.n4478 185
R393 VDD.n2308 VDD.n2307 185
R394 VDD.n2307 VDD.n2306 185
R395 VDD.n4453 VDD.n4452 185
R396 VDD.n4454 VDD.n4453 185
R397 VDD.n2364 VDD.n2363 185
R398 VDD.n2365 VDD.n2364 185
R399 VDD.n2353 VDD.n2351 185
R400 VDD.n4433 VDD.n2353 185
R401 VDD.n2406 VDD.n2405 185
R402 VDD.n2407 VDD.n2406 185
R403 VDD.n2395 VDD.n2393 185
R404 VDD.n4411 VDD.n2395 185
R405 VDD.n4409 VDD.n4408 185
R406 VDD.n4410 VDD.n4409 185
R407 VDD.n2404 VDD.n2394 185
R408 VDD.n2408 VDD.n2394 185
R409 VDD.n4431 VDD.n4430 185
R410 VDD.n4432 VDD.n4431 185
R411 VDD.n2362 VDD.n2352 185
R412 VDD.n2366 VDD.n2352 185
R413 VDD.n2536 VDD.n2535 185
R414 VDD.n2302 VDD.n2301 185
R415 VDD.n4455 VDD.n2302 185
R416 VDD.n2257 VDD.n2235 185
R417 VDD.n4480 VDD.n2235 185
R418 VDD.n2252 VDD.n2251 185
R419 VDD.n2253 VDD.n2252 185
R420 VDD.n2240 VDD.n2239 185
R421 VDD.n2241 VDD.n2240 185
R422 VDD.n2193 VDD.n2179 185
R423 VDD.n4507 VDD.n2179 185
R424 VDD.n2309 VDD.n2304 185
R425 VDD.n2304 VDD.n2303 185
R426 VDD.n2178 VDD.n2176 185
R427 VDD.n2190 VDD.n2178 185
R428 VDD.n4530 VDD.n4529 185
R429 VDD.n4531 VDD.n4530 185
R430 VDD.n2140 VDD.n2130 185
R431 VDD.n2144 VDD.n2130 185
R432 VDD.n4552 VDD.n4551 185
R433 VDD.n4553 VDD.n4552 185
R434 VDD.n2098 VDD.n2088 185
R435 VDD.n2102 VDD.n2088 185
R436 VDD.n2186 VDD.n2185 185
R437 VDD.n2185 VDD.n2184 185
R438 VDD.n2182 VDD.n2181 185
R439 VDD.n2183 VDD.n2182 185
R440 VDD.n2038 VDD.n2037 185
R441 VDD.n4576 VDD.n2038 185
R442 VDD.n1993 VDD.n1971 185
R443 VDD.n4601 VDD.n1971 185
R444 VDD.n1988 VDD.n1987 185
R445 VDD.n1989 VDD.n1988 185
R446 VDD.n1976 VDD.n1975 185
R447 VDD.n1977 VDD.n1976 185
R448 VDD.n1929 VDD.n1915 185
R449 VDD.n4628 VDD.n1915 185
R450 VDD.n2045 VDD.n2040 185
R451 VDD.n2040 VDD.n2039 185
R452 VDD.n1914 VDD.n1912 185
R453 VDD.n1926 VDD.n1914 185
R454 VDD.n4651 VDD.n4650 185
R455 VDD.n4652 VDD.n4651 185
R456 VDD.n1876 VDD.n1866 185
R457 VDD.n1880 VDD.n1866 185
R458 VDD.n4673 VDD.n4672 185
R459 VDD.n4674 VDD.n4673 185
R460 VDD.n1834 VDD.n1824 185
R461 VDD.n1838 VDD.n1824 185
R462 VDD.n1922 VDD.n1921 185
R463 VDD.n1921 VDD.n1920 185
R464 VDD.n1918 VDD.n1917 185
R465 VDD.n1919 VDD.n1918 185
R466 VDD.n1774 VDD.n1773 185
R467 VDD.n4697 VDD.n1774 185
R468 VDD.n1729 VDD.n1707 185
R469 VDD.n4722 VDD.n1707 185
R470 VDD.n1724 VDD.n1723 185
R471 VDD.n1725 VDD.n1724 185
R472 VDD.n1712 VDD.n1711 185
R473 VDD.n1713 VDD.n1712 185
R474 VDD.n1665 VDD.n1651 185
R475 VDD.n4749 VDD.n1651 185
R476 VDD.n1781 VDD.n1776 185
R477 VDD.n1776 VDD.n1775 185
R478 VDD.n1650 VDD.n1648 185
R479 VDD.n1662 VDD.n1650 185
R480 VDD.n4772 VDD.n4771 185
R481 VDD.n4773 VDD.n4772 185
R482 VDD.n1612 VDD.n1602 185
R483 VDD.n1616 VDD.n1602 185
R484 VDD.n4794 VDD.n4793 185
R485 VDD.n4795 VDD.n4794 185
R486 VDD.n1570 VDD.n1560 185
R487 VDD.n1574 VDD.n1560 185
R488 VDD.n1658 VDD.n1657 185
R489 VDD.n1657 VDD.n1656 185
R490 VDD.n1654 VDD.n1653 185
R491 VDD.n1655 VDD.n1654 185
R492 VDD.n1510 VDD.n1509 185
R493 VDD.n4818 VDD.n1510 185
R494 VDD.n1465 VDD.n1443 185
R495 VDD.n4843 VDD.n1443 185
R496 VDD.n1460 VDD.n1459 185
R497 VDD.n1461 VDD.n1460 185
R498 VDD.n1397 VDD.n1382 185
R499 VDD.n4870 VDD.n1382 185
R500 VDD.n1448 VDD.n1447 185
R501 VDD.n1449 VDD.n1448 185
R502 VDD.n1517 VDD.n1512 185
R503 VDD.n1512 VDD.n1511 185
R504 VDD.n1394 VDD.n1381 185
R505 VDD.n4928 VDD.n4927 185
R506 VDD.n4929 VDD.n4928 185
R507 VDD.n1249 VDD.n1246 185
R508 VDD.n4922 VDD.n1246 185
R509 VDD.n1321 VDD.n1320 185
R510 VDD.n1322 VDD.n1321 185
R511 VDD.n1333 VDD.n1332 185
R512 VDD.n1334 VDD.n1333 185
R513 VDD.n1338 VDD.n1316 185
R514 VDD.n4895 VDD.n1316 185
R515 VDD.n1388 VDD.n1387 185
R516 VDD.n1387 VDD.n1386 185
R517 VDD.n4926 VDD.n1243 185
R518 VDD.n1243 VDD.n1242 185
R519 VDD.n4920 VDD.n4919 185
R520 VDD.n4921 VDD.n4920 185
R521 VDD.n1325 VDD.n1324 185
R522 VDD.n1324 VDD.n1323 185
R523 VDD.n1315 VDD.n1313 185
R524 VDD.n1335 VDD.n1315 185
R525 VDD.n4893 VDD.n4892 185
R526 VDD.n4894 VDD.n4893 185
R527 VDD.n1389 VDD.n1384 185
R528 VDD.n1384 VDD.n1383 185
R529 VDD.n4971 VDD.n4970 185
R530 VDD.n4970 VDD.n4969 185
R531 VDD.n5043 VDD.n1188 185
R532 VDD.n5072 VDD.n5071 185
R533 VDD.n1161 VDD.n1160 185
R534 VDD.n5106 VDD.n5105 185
R535 VDD.n5124 VDD.n5123 185
R536 VDD.n1134 VDD.n1116 185
R537 VDD.n5155 VDD.n1115 185
R538 VDD.n5185 VDD.n5184 185
R539 VDD.n1083 VDD.n1082 185
R540 VDD.n5213 VDD.n5212 185
R541 VDD.n5271 VDD.n1053 185
R542 VDD.n5300 VDD.n5299 185
R543 VDD.n1026 VDD.n1025 185
R544 VDD.n5334 VDD.n5333 185
R545 VDD.n5352 VDD.n5351 185
R546 VDD.n999 VDD.n981 185
R547 VDD.n5383 VDD.n980 185
R548 VDD.n5413 VDD.n5412 185
R549 VDD.n948 VDD.n947 185
R550 VDD.n5441 VDD.n5440 185
R551 VDD.n5499 VDD.n918 185
R552 VDD.n5528 VDD.n5527 185
R553 VDD.n891 VDD.n890 185
R554 VDD.n5562 VDD.n5561 185
R555 VDD.n5580 VDD.n5579 185
R556 VDD.n864 VDD.n846 185
R557 VDD.n5611 VDD.n845 185
R558 VDD.n5641 VDD.n5640 185
R559 VDD.n813 VDD.n812 185
R560 VDD.n5669 VDD.n5668 185
R561 VDD.n5727 VDD.n783 185
R562 VDD.n5756 VDD.n5755 185
R563 VDD.n756 VDD.n755 185
R564 VDD.n5790 VDD.n5789 185
R565 VDD.n5807 VDD.n5806 185
R566 VDD.n5829 VDD.n715 185
R567 VDD.n5849 VDD.n714 185
R568 VDD.n713 VDD.n711 185
R569 VDD.n5884 VDD.n694 185
R570 VDD.n5918 VDD.n5917 185
R571 VDD.n5920 VDD.n674 185
R572 VDD.n5887 VDD.n5886 185
R573 VDD.n710 VDD.n695 185
R574 VDD.n5850 VDD.n709 185
R575 VDD.n5828 VDD.n5827 185
R576 VDD.n5787 VDD.n754 185
R577 VDD.n5761 VDD.n5760 185
R578 VDD.n5754 VDD.n771 185
R579 VDD.n5725 VDD.n5724 185
R580 VDD.n5809 VDD.n734 185
R581 VDD.n5708 VDD.n5707 185
R582 VDD.n5670 VDD.n795 185
R583 VDD.n5664 VDD.n5663 185
R584 VDD.n5643 VDD.n827 185
R585 VDD.n5614 VDD.n5613 185
R586 VDD.n5704 VDD.n5703 185
R587 VDD.n5703 VDD.n641 185
R588 VDD.n5702 VDD.n794 185
R589 VDD.n867 VDD.n865 185
R590 VDD.n5559 VDD.n889 185
R591 VDD.n5533 VDD.n5532 185
R592 VDD.n5526 VDD.n906 185
R593 VDD.n5497 VDD.n5496 185
R594 VDD.n5582 VDD.n860 185
R595 VDD.n5480 VDD.n5479 185
R596 VDD.n5442 VDD.n930 185
R597 VDD.n5436 VDD.n5435 185
R598 VDD.n5415 VDD.n962 185
R599 VDD.n5386 VDD.n5385 185
R600 VDD.n5476 VDD.n5475 185
R601 VDD.n5475 VDD.n641 185
R602 VDD.n5474 VDD.n929 185
R603 VDD.n1002 VDD.n1000 185
R604 VDD.n5331 VDD.n1024 185
R605 VDD.n5305 VDD.n5304 185
R606 VDD.n5298 VDD.n1041 185
R607 VDD.n5269 VDD.n5268 185
R608 VDD.n5354 VDD.n995 185
R609 VDD.n5252 VDD.n5251 185
R610 VDD.n5214 VDD.n1065 185
R611 VDD.n5208 VDD.n5207 185
R612 VDD.n5187 VDD.n1097 185
R613 VDD.n5158 VDD.n5157 185
R614 VDD.n5248 VDD.n5247 185
R615 VDD.n5247 VDD.n641 185
R616 VDD.n5246 VDD.n1064 185
R617 VDD.n1137 VDD.n1135 185
R618 VDD.n5103 VDD.n1159 185
R619 VDD.n5077 VDD.n5076 185
R620 VDD.n5041 VDD.n5040 185
R621 VDD.n5070 VDD.n1176 185
R622 VDD.n5126 VDD.n1130 185
R623 VDD.n6069 VDD.n6068 185
R624 VDD.n656 VDD.n655 185
R625 VDD.n5967 VDD.n5966 185
R626 VDD.n6044 VDD.n6043 185
R627 VDD.n6014 VDD.n6013 185
R628 VDD.n6016 VDD.n6015 185
R629 VDD.n6042 VDD.n644 185
R630 VDD.n6073 VDD.n644 185
R631 VDD.n5968 VDD.n648 185
R632 VDD.n6073 VDD.n648 185
R633 VDD.n5958 VDD.n642 185
R634 VDD.n6073 VDD.n642 185
R635 VDD.n640 VDD.n639 185
R636 VDD.n6070 VDD.n651 185
R637 VDD.n6122 VDD.n604 185
R638 VDD.n6126 VDD.n604 185
R639 VDD.n7219 VDD.n7218 185
R640 VDD.n27 VDD.n26 185
R641 VDD.n7117 VDD.n7116 185
R642 VDD.n7194 VDD.n7193 185
R643 VDD.n7164 VDD.n7163 185
R644 VDD.n7108 VDD.n13 185
R645 VDD.n7223 VDD.n13 185
R646 VDD.n7118 VDD.n19 185
R647 VDD.n7223 VDD.n19 185
R648 VDD.n7192 VDD.n15 185
R649 VDD.n7223 VDD.n15 185
R650 VDD.n7166 VDD.n7165 185
R651 VDD.n11 VDD.n10 185
R652 VDD.n7220 VDD.n22 185
R653 VDD.n6195 VDD.n6194 185
R654 VDD.n540 VDD.n539 185
R655 VDD.n6244 VDD.n6243 185
R656 VDD.n6263 VDD.n527 185
R657 VDD.n6281 VDD.n6280 185
R658 VDD.n6300 VDD.n492 185
R659 VDD.n6299 VDD.n495 185
R660 VDD.n6303 VDD.n494 185
R661 VDD.n493 VDD.n478 185
R662 VDD.n6339 VDD.n6338 185
R663 VDD.n6336 VDD.n477 185
R664 VDD.n6366 VDD.n6365 185
R665 VDD.n6368 VDD.n459 185
R666 VDD.n6387 VDD.n6386 185
R667 VDD.n449 VDD.n448 185
R668 VDD.n6393 VDD.n447 185
R669 VDD.n421 VDD.n420 185
R670 VDD.n406 VDD.n405 185
R671 VDD.n6470 VDD.n6469 185
R672 VDD.n6489 VDD.n393 185
R673 VDD.n6507 VDD.n6506 185
R674 VDD.n6526 VDD.n358 185
R675 VDD.n6525 VDD.n361 185
R676 VDD.n6529 VDD.n360 185
R677 VDD.n359 VDD.n344 185
R678 VDD.n6565 VDD.n6564 185
R679 VDD.n6562 VDD.n343 185
R680 VDD.n6592 VDD.n6591 185
R681 VDD.n6594 VDD.n325 185
R682 VDD.n6613 VDD.n6612 185
R683 VDD.n315 VDD.n314 185
R684 VDD.n6619 VDD.n313 185
R685 VDD.n287 VDD.n286 185
R686 VDD.n272 VDD.n271 185
R687 VDD.n6696 VDD.n6695 185
R688 VDD.n6715 VDD.n259 185
R689 VDD.n6733 VDD.n6732 185
R690 VDD.n6752 VDD.n224 185
R691 VDD.n6751 VDD.n227 185
R692 VDD.n6755 VDD.n226 185
R693 VDD.n225 VDD.n210 185
R694 VDD.n6791 VDD.n6790 185
R695 VDD.n6788 VDD.n209 185
R696 VDD.n6818 VDD.n6817 185
R697 VDD.n6820 VDD.n191 185
R698 VDD.n6839 VDD.n6838 185
R699 VDD.n181 VDD.n180 185
R700 VDD.n6845 VDD.n179 185
R701 VDD.n153 VDD.n152 185
R702 VDD.n138 VDD.n137 185
R703 VDD.n6922 VDD.n6921 185
R704 VDD.n6941 VDD.n125 185
R705 VDD.n6959 VDD.n6958 185
R706 VDD.n6978 VDD.n90 185
R707 VDD.n6977 VDD.n93 185
R708 VDD.n6981 VDD.n92 185
R709 VDD.n91 VDD.n76 185
R710 VDD.n7017 VDD.n7016 185
R711 VDD.n7014 VDD.n75 185
R712 VDD.n7044 VDD.n7043 185
R713 VDD.n7046 VDD.n57 185
R714 VDD.n7070 VDD.n7069 185
R715 VDD.n46 VDD.n45 185
R716 VDD.n6939 VDD.n6938 185
R717 VDD.n6919 VDD.n136 185
R718 VDD.n6894 VDD.n6893 185
R719 VDD.n6873 VDD.n6872 185
R720 VDD.n6960 VDD.n105 185
R721 VDD.n164 VDD.n163 185
R722 VDD.n6713 VDD.n6712 185
R723 VDD.n6693 VDD.n270 185
R724 VDD.n6668 VDD.n6667 185
R725 VDD.n6647 VDD.n6646 185
R726 VDD.n6734 VDD.n239 185
R727 VDD.n298 VDD.n297 185
R728 VDD.n6487 VDD.n6486 185
R729 VDD.n6467 VDD.n404 185
R730 VDD.n6442 VDD.n6441 185
R731 VDD.n6421 VDD.n6420 185
R732 VDD.n6508 VDD.n373 185
R733 VDD.n432 VDD.n431 185
R734 VDD.n6261 VDD.n6260 185
R735 VDD.n6241 VDD.n538 185
R736 VDD.n6216 VDD.n6215 185
R737 VDD.n6282 VDD.n507 185
R738 VDD.n6193 VDD.n555 185
R739 VDD.n4931 VDD 165.668
R740 VDD.n7251 VDD 160.49
R741 VDD.n6130 VDD.t51 152.88
R742 VDD.n7254 VDD.t55 152.88
R743 VDD.n630 VDD.t47 152.879
R744 VDD.n2472 VDD.t59 152.879
R745 VDD.n2619 VDD.t45 152.879
R746 VDD.n1235 VDD.t76 152.879
R747 VDD.n4956 VDD.t49 152.879
R748 VDD.n0 VDD.t43 152.879
R749 VDD.t32 VDD 141.034
R750 VDD.n2759 VDD 131.415
R751 VDD.n1393 VDD 131.415
R752 VDD.t75 VDD.n1240 113.897
R753 VDD.n5921 VDD.n5920 111.234
R754 VDD.n5041 VDD.n1189 111.234
R755 VDD.n7012 VDD.n76 111.177
R756 VDD.n7048 VDD.n7046 111.177
R757 VDD.n6872 VDD.n6870 111.177
R758 VDD.n6893 VDD.n6891 111.177
R759 VDD.n6919 VDD.n6918 111.177
R760 VDD.n6939 VDD.n126 111.177
R761 VDD.n6786 VDD.n210 111.177
R762 VDD.n6822 VDD.n6820 111.177
R763 VDD.n6646 VDD.n6644 111.177
R764 VDD.n6667 VDD.n6665 111.177
R765 VDD.n6693 VDD.n6692 111.177
R766 VDD.n6713 VDD.n260 111.177
R767 VDD.n6560 VDD.n344 111.177
R768 VDD.n6596 VDD.n6594 111.177
R769 VDD.n6420 VDD.n6418 111.177
R770 VDD.n6441 VDD.n6439 111.177
R771 VDD.n6467 VDD.n6466 111.177
R772 VDD.n6487 VDD.n394 111.177
R773 VDD.n6334 VDD.n478 111.177
R774 VDD.n6370 VDD.n6368 111.177
R775 VDD.n6215 VDD.n6213 111.177
R776 VDD.n6241 VDD.n6240 111.177
R777 VDD.n6261 VDD.n528 111.177
R778 VDD.n7218 VDD.n7217 111.177
R779 VDD.n7114 VDD.n13 111.177
R780 VDD.n7195 VDD.n19 111.177
R781 VDD.n7161 VDD.n15 111.177
R782 VDD.n6068 VDD.n6067 111.177
R783 VDD.n5964 VDD.n642 111.177
R784 VDD.n6045 VDD.n648 111.177
R785 VDD.n6011 VDD.n644 111.177
R786 VDD.n5847 VDD.n715 111.177
R787 VDD.n5882 VDD.n695 111.177
R788 VDD.n5725 VDD.n784 111.177
R789 VDD.n5760 VDD.n5758 111.177
R790 VDD.n5807 VDD.n744 111.177
R791 VDD.n5609 VDD.n846 111.177
R792 VDD.n5645 VDD.n5643 111.177
R793 VDD.n5700 VDD.n795 111.177
R794 VDD.n5497 VDD.n919 111.177
R795 VDD.n5532 VDD.n5530 111.177
R796 VDD.n5580 VDD.n879 111.177
R797 VDD.n5381 VDD.n981 111.177
R798 VDD.n5417 VDD.n5415 111.177
R799 VDD.n5472 VDD.n930 111.177
R800 VDD.n5269 VDD.n1054 111.177
R801 VDD.n5304 VDD.n5302 111.177
R802 VDD.n5352 VDD.n1014 111.177
R803 VDD.n5153 VDD.n1116 111.177
R804 VDD.n5189 VDD.n5187 111.177
R805 VDD.n5244 VDD.n1065 111.177
R806 VDD.n5076 VDD.n5074 111.177
R807 VDD.n5124 VDD.n1149 111.177
R808 VDD.n4924 VDD.n1246 111.177
R809 VDD.n1321 VDD.n1248 111.177
R810 VDD.n1333 VDD.n1318 111.177
R811 VDD.n4897 VDD.n1316 111.177
R812 VDD.n1387 VDD.n1337 111.177
R813 VDD.n4453 VDD.n2326 111.177
R814 VDD.n4435 VDD.n2352 111.177
R815 VDD.n4431 VDD.n2368 111.177
R816 VDD.n4413 VDD.n2394 111.177
R817 VDD.n4409 VDD.n2410 111.177
R818 VDD.n4509 VDD.n2179 111.177
R819 VDD.n2240 VDD.n2192 111.177
R820 VDD.n2252 VDD.n2237 111.177
R821 VDD.n4482 VDD.n2235 111.177
R822 VDD.n2307 VDD.n2256 111.177
R823 VDD.n4574 VDD.n2062 111.177
R824 VDD.n4556 VDD.n2088 111.177
R825 VDD.n4552 VDD.n2104 111.177
R826 VDD.n4534 VDD.n2130 111.177
R827 VDD.n4530 VDD.n2146 111.177
R828 VDD.n4630 VDD.n1915 111.177
R829 VDD.n1976 VDD.n1928 111.177
R830 VDD.n1988 VDD.n1973 111.177
R831 VDD.n4603 VDD.n1971 111.177
R832 VDD.n2043 VDD.n1992 111.177
R833 VDD.n4695 VDD.n1798 111.177
R834 VDD.n4677 VDD.n1824 111.177
R835 VDD.n4673 VDD.n1840 111.177
R836 VDD.n4655 VDD.n1866 111.177
R837 VDD.n4651 VDD.n1882 111.177
R838 VDD.n4751 VDD.n1651 111.177
R839 VDD.n1712 VDD.n1664 111.177
R840 VDD.n1724 VDD.n1709 111.177
R841 VDD.n4724 VDD.n1707 111.177
R842 VDD.n1779 VDD.n1728 111.177
R843 VDD.n4816 VDD.n1534 111.177
R844 VDD.n4798 VDD.n1560 111.177
R845 VDD.n4794 VDD.n1576 111.177
R846 VDD.n4776 VDD.n1602 111.177
R847 VDD.n4772 VDD.n1618 111.177
R848 VDD.n4872 VDD.n1382 111.177
R849 VDD.n1448 VDD.n1396 111.177
R850 VDD.n1460 VDD.n1445 111.177
R851 VDD.n4845 VDD.n1443 111.177
R852 VDD.n1515 VDD.n1464 111.177
R853 VDD.n2639 VDD.n2450 111.177
R854 VDD.n4374 VDD.n2448 111.177
R855 VDD.n2696 VDD.n2643 111.177
R856 VDD.n2708 VDD.n2693 111.177
R857 VDD.n4347 VDD.n2691 111.177
R858 VDD.n3916 VDD.n3682 111.177
R859 VDD.n3899 VDD.n3710 111.177
R860 VDD.n3895 VDD.n3725 111.177
R861 VDD.n3878 VDD.n3753 111.177
R862 VDD.n3874 VDD.n3768 111.177
R863 VDD.n3972 VDD.n3535 111.177
R864 VDD.n3596 VDD.n3548 111.177
R865 VDD.n3608 VDD.n3593 111.177
R866 VDD.n3945 VDD.n3591 111.177
R867 VDD.n3663 VDD.n3612 111.177
R868 VDD.n4035 VDD.n3416 111.177
R869 VDD.n4018 VDD.n3444 111.177
R870 VDD.n4014 VDD.n3459 111.177
R871 VDD.n3997 VDD.n3487 111.177
R872 VDD.n3993 VDD.n3502 111.177
R873 VDD.n4091 VDD.n3269 111.177
R874 VDD.n3330 VDD.n3282 111.177
R875 VDD.n3342 VDD.n3327 111.177
R876 VDD.n4064 VDD.n3325 111.177
R877 VDD.n3397 VDD.n3346 111.177
R878 VDD.n4154 VDD.n3150 111.177
R879 VDD.n4137 VDD.n3178 111.177
R880 VDD.n4133 VDD.n3193 111.177
R881 VDD.n4116 VDD.n3221 111.177
R882 VDD.n4112 VDD.n3236 111.177
R883 VDD.n4210 VDD.n3003 111.177
R884 VDD.n3064 VDD.n3016 111.177
R885 VDD.n3076 VDD.n3061 111.177
R886 VDD.n4183 VDD.n3059 111.177
R887 VDD.n3131 VDD.n3080 111.177
R888 VDD.n4273 VDD.n2852 111.177
R889 VDD.n4256 VDD.n2912 111.177
R890 VDD.n4252 VDD.n2927 111.177
R891 VDD.n4235 VDD.n2955 111.177
R892 VDD.n4231 VDD.n2970 111.177
R893 VDD.n2770 VDD.n2762 111.177
R894 VDD.n4321 VDD.n2756 111.177
R895 VDD.n2822 VDD.n2774 111.177
R896 VDD.n2834 VDD.n2819 111.177
R897 VDD.n4294 VDD.n2817 111.177
R898 VDD.n4931 VDD.t48 108.719
R899 VDD.n2486 VDD.n2484 92.5005
R900 VDD.n2597 VDD.n2486 92.5005
R901 VDD.n2621 VDD.n2620 92.5005
R902 VDD.n2622 VDD.n2621 92.5005
R903 VDD.n2485 VDD.n2473 92.5005
R904 VDD.n2563 VDD.n2485 92.5005
R905 VDD.n1238 VDD.n1236 92.5005
R906 VDD.n1240 VDD.n1238 92.5005
R907 VDD.n4968 VDD.n1239 92.5005
R908 VDD.n1239 VDD.n1237 92.5005
R909 VDD.n4957 VDD.n4932 92.5005
R910 VDD.n4932 VDD.n4931 92.5005
R911 VDD.n6124 VDD.n6123 92.5005
R912 VDD.n6125 VDD.n6124 92.5005
R913 VDD.n6129 VDD.n6128 92.5005
R914 VDD.n6128 VDD.n6127 92.5005
R915 VDD.n6095 VDD.n6094 92.5005
R916 VDD.n6096 VDD.n6095 92.5005
R917 VDD.n7253 VDD.n7252 92.5005
R918 VDD.n7252 VDD.n7251 92.5005
R919 VDD.n6157 VDD.n6156 92.5005
R920 VDD.n6158 VDD.n6157 92.5005
R921 VDD.n4990 VDD 89.6591
R922 VDD.n2564 VDD.n2562 88.3561
R923 VDD.n4873 VDD.n1379 86.9025
R924 VDD.n2538 VDD.n2537 86.9025
R925 VDD.n2758 VDD.n2739 86.9025
R926 VDD.n3821 VDD.n3820 86.9025
R927 VDD.n5125 VDD.n641 85.9427
R928 VDD.n1136 VDD.n641 85.9427
R929 VDD.n5186 VDD.n641 85.9427
R930 VDD.n5211 VDD.n641 85.9427
R931 VDD.n5250 VDD.n641 85.9427
R932 VDD.n5353 VDD.n641 85.9427
R933 VDD.n1001 VDD.n641 85.9427
R934 VDD.n5414 VDD.n641 85.9427
R935 VDD.n5439 VDD.n641 85.9427
R936 VDD.n5478 VDD.n641 85.9427
R937 VDD.n5581 VDD.n641 85.9427
R938 VDD.n866 VDD.n641 85.9427
R939 VDD.n5642 VDD.n641 85.9427
R940 VDD.n5667 VDD.n641 85.9427
R941 VDD.n5706 VDD.n641 85.9427
R942 VDD.n5808 VDD.n641 85.9427
R943 VDD.n5826 VDD.n641 85.9427
R944 VDD.n712 VDD.n641 85.9427
R945 VDD.n5919 VDD.n641 85.9427
R946 VDD.n5759 VDD.n641 85.9427
R947 VDD.n5726 VDD.n641 85.9427
R948 VDD.n5531 VDD.n641 85.9427
R949 VDD.n5498 VDD.n641 85.9427
R950 VDD.n5303 VDD.n641 85.9427
R951 VDD.n5270 VDD.n641 85.9427
R952 VDD.n5075 VDD.n641 85.9427
R953 VDD.n5042 VDD.n641 85.9427
R954 VDD.n6073 VDD.n650 85.9427
R955 VDD.n6074 VDD.n6073 85.9427
R956 VDD.n7223 VDD.n21 85.9427
R957 VDD.n7224 VDD.n7223 85.9427
R958 VDD.n6214 VDD.n12 85.9427
R959 VDD.n6242 VDD.n12 85.9427
R960 VDD.n6262 VDD.n12 85.9427
R961 VDD.n6302 VDD.n12 85.9427
R962 VDD.n6367 VDD.n12 85.9427
R963 VDD.n6392 VDD.n12 85.9427
R964 VDD.n6389 VDD.n12 85.9427
R965 VDD.n6419 VDD.n12 85.9427
R966 VDD.n6440 VDD.n12 85.9427
R967 VDD.n6468 VDD.n12 85.9427
R968 VDD.n6488 VDD.n12 85.9427
R969 VDD.n6528 VDD.n12 85.9427
R970 VDD.n6593 VDD.n12 85.9427
R971 VDD.n6618 VDD.n12 85.9427
R972 VDD.n6615 VDD.n12 85.9427
R973 VDD.n6645 VDD.n12 85.9427
R974 VDD.n6666 VDD.n12 85.9427
R975 VDD.n6694 VDD.n12 85.9427
R976 VDD.n6714 VDD.n12 85.9427
R977 VDD.n6754 VDD.n12 85.9427
R978 VDD.n6819 VDD.n12 85.9427
R979 VDD.n6844 VDD.n12 85.9427
R980 VDD.n6841 VDD.n12 85.9427
R981 VDD.n6871 VDD.n12 85.9427
R982 VDD.n6892 VDD.n12 85.9427
R983 VDD.n6920 VDD.n12 85.9427
R984 VDD.n6940 VDD.n12 85.9427
R985 VDD.n6980 VDD.n12 85.9427
R986 VDD.n7045 VDD.n12 85.9427
R987 VDD.n3008 VDD 85.8969
R988 VDD.n3274 VDD 85.8969
R989 VDD.n3540 VDD 85.8969
R990 VDD VDD.n3822 85.8969
R991 VDD.n1656 VDD 85.8969
R992 VDD.n1920 VDD 85.8969
R993 VDD.n2184 VDD 85.8969
R994 VDD VDD.n2539 85.8969
R995 VDD.n2594 VDD.t44 85.2946
R996 VDD.n2626 VDD 79.2895
R997 VDD VDD.n4930 79.2895
R998 VDD VDD.n6158 77.6572
R999 VDD.n2564 VDD 73.5299
R1000 VDD.n2598 VDD.t58 72.5495
R1001 VDD.n1240 VDD 72.4801
R1002 VDD VDD.t56 71.2138
R1003 VDD VDD.t31 71.2138
R1004 VDD.n6177 VDD.t19 70.3649
R1005 VDD.n5016 VDD.t63 70.3649
R1006 VDD.n3831 VDD.t6 70.3628
R1007 VDD.n2507 VDD.t30 70.3628
R1008 VDD.t50 VDD.n6126 69.629
R1009 VDD.n6077 VDD.t12 68.0287
R1010 VDD.n7227 VDD.t61 68.0287
R1011 VDD.n2624 VDD.t35 68.0287
R1012 VDD.n1267 VDD.t25 68.0287
R1013 VDD.n1532 VDD.t66 67.9081
R1014 VDD.n1796 VDD.t20 67.9081
R1015 VDD.n2060 VDD.t72 67.9081
R1016 VDD.n2324 VDD.t28 67.9081
R1017 VDD.n2850 VDD.t41 67.9081
R1018 VDD.n3148 VDD.t64 67.9081
R1019 VDD.n3414 VDD.t69 67.9081
R1020 VDD.n3680 VDD.t73 67.9081
R1021 VDD.n6194 VDD.n6192 67.5405
R1022 VDD.n7071 VDD.n7070 67.5405
R1023 VDD.n6959 VDD.n115 67.3307
R1024 VDD.n6733 VDD.n249 67.3307
R1025 VDD.n6507 VDD.n383 67.3307
R1026 VDD.n6281 VDD.n517 67.3307
R1027 VDD.n7165 VDD.n17 67.3307
R1028 VDD.n6015 VDD.n646 67.3307
R1029 VDD.n5851 VDD.n5850 67.3307
R1030 VDD.n5886 VDD.n5885 67.3307
R1031 VDD.n5613 VDD.n5612 67.3307
R1032 VDD.n5665 VDD.n5664 67.3307
R1033 VDD.n5385 VDD.n5384 67.3307
R1034 VDD.n5437 VDD.n5436 67.3307
R1035 VDD.n5157 VDD.n5156 67.3307
R1036 VDD.n5209 VDD.n5208 67.3307
R1037 VDD.n5787 VDD.n5786 67.3307
R1038 VDD.n5728 VDD.n771 67.3307
R1039 VDD.n5559 VDD.n5558 67.3307
R1040 VDD.n5500 VDD.n906 67.3307
R1041 VDD.n5331 VDD.n5330 67.3307
R1042 VDD.n5272 VDD.n1041 67.3307
R1043 VDD.n5103 VDD.n5102 67.3307
R1044 VDD.n5044 VDD.n1176 67.3307
R1045 VDD.n6301 VDD.n6300 67.3307
R1046 VDD.n6338 VDD.n6337 67.3307
R1047 VDD.n6388 VDD.n6387 67.3307
R1048 VDD.n6527 VDD.n6526 67.3307
R1049 VDD.n6564 VDD.n6563 67.3307
R1050 VDD.n6614 VDD.n6613 67.3307
R1051 VDD.n6753 VDD.n6752 67.3307
R1052 VDD.n6790 VDD.n6789 67.3307
R1053 VDD.n6840 VDD.n6839 67.3307
R1054 VDD.n6979 VDD.n6978 67.3307
R1055 VDD.n7016 VDD.n7015 67.3307
R1056 VDD.t3 VDD.t5 65.1272
R1057 VDD.t34 VDD.t29 65.1272
R1058 VDD VDD.n2622 62.7456
R1059 VDD.n6127 VDD 59.137
R1060 VDD.t5 VDD 55.7965
R1061 VDD.t29 VDD 55.7965
R1062 VDD.n619 VDD.n605 48.6451
R1063 VDD.t14 VDD.t62 47.6077
R1064 VDD.t77 VDD.t18 47.6077
R1065 VDD.n594 VDD.t15 47.1434
R1066 VDD.n594 VDD.t13 47.1434
R1067 VDD.n3838 VDD.t52 47.1434
R1068 VDD.n3838 VDD.t39 47.1434
R1069 VDD.n2514 VDD.t36 47.1434
R1070 VDD.n2514 VDD.t33 47.1434
R1071 VDD.n1224 VDD.t24 47.1434
R1072 VDD.n1224 VDD.t27 47.1434
R1073 VDD.n2640 VDD.n2449 46.2524
R1074 VDD.n4373 VDD.n4372 46.2524
R1075 VDD.n2697 VDD.n2642 46.2524
R1076 VDD.n2709 VDD.n2692 46.2524
R1077 VDD.n4346 VDD.n4345 46.2524
R1078 VDD.n2771 VDD.n2757 46.2524
R1079 VDD.n4320 VDD.n4319 46.2524
R1080 VDD.n2823 VDD.n2773 46.2524
R1081 VDD.n2835 VDD.n2818 46.2524
R1082 VDD.n4293 VDD.n4292 46.2524
R1083 VDD.n4274 VDD.n2851 46.2524
R1084 VDD.n4255 VDD.n2925 46.2524
R1085 VDD.n4253 VDD.n2926 46.2524
R1086 VDD.n4234 VDD.n2968 46.2524
R1087 VDD.n4232 VDD.n2969 46.2524
R1088 VDD.n4209 VDD.n4208 46.2524
R1089 VDD.n3065 VDD.n3015 46.2524
R1090 VDD.n3077 VDD.n3060 46.2524
R1091 VDD.n4182 VDD.n4181 46.2524
R1092 VDD.n3130 VDD.n3079 46.2524
R1093 VDD.n4155 VDD.n3149 46.2524
R1094 VDD.n4136 VDD.n3191 46.2524
R1095 VDD.n4134 VDD.n3192 46.2524
R1096 VDD.n4115 VDD.n3234 46.2524
R1097 VDD.n4113 VDD.n3235 46.2524
R1098 VDD.n4090 VDD.n4089 46.2524
R1099 VDD.n3331 VDD.n3281 46.2524
R1100 VDD.n3343 VDD.n3326 46.2524
R1101 VDD.n4063 VDD.n4062 46.2524
R1102 VDD.n3396 VDD.n3345 46.2524
R1103 VDD.n4036 VDD.n3415 46.2524
R1104 VDD.n4017 VDD.n3457 46.2524
R1105 VDD.n4015 VDD.n3458 46.2524
R1106 VDD.n3996 VDD.n3500 46.2524
R1107 VDD.n3994 VDD.n3501 46.2524
R1108 VDD.n3971 VDD.n3970 46.2524
R1109 VDD.n3597 VDD.n3547 46.2524
R1110 VDD.n3609 VDD.n3592 46.2524
R1111 VDD.n3944 VDD.n3943 46.2524
R1112 VDD.n3662 VDD.n3611 46.2524
R1113 VDD.n3917 VDD.n3681 46.2524
R1114 VDD.n3898 VDD.n3723 46.2524
R1115 VDD.n3896 VDD.n3724 46.2524
R1116 VDD.n3877 VDD.n3766 46.2524
R1117 VDD.n3875 VDD.n3767 46.2524
R1118 VDD.n4923 VDD.n4922 46.2524
R1119 VDD.n1322 VDD.n1247 46.2524
R1120 VDD.n1334 VDD.n1317 46.2524
R1121 VDD.n4896 VDD.n4895 46.2524
R1122 VDD.n1386 VDD.n1336 46.2524
R1123 VDD.n4871 VDD.n4870 46.2524
R1124 VDD.n1449 VDD.n1395 46.2524
R1125 VDD.n1461 VDD.n1444 46.2524
R1126 VDD.n4844 VDD.n4843 46.2524
R1127 VDD.n1514 VDD.n1463 46.2524
R1128 VDD.n4817 VDD.n1533 46.2524
R1129 VDD.n4797 VDD.n1574 46.2524
R1130 VDD.n4795 VDD.n1575 46.2524
R1131 VDD.n4775 VDD.n1616 46.2524
R1132 VDD.n4773 VDD.n1617 46.2524
R1133 VDD.n4750 VDD.n4749 46.2524
R1134 VDD.n1713 VDD.n1663 46.2524
R1135 VDD.n1725 VDD.n1708 46.2524
R1136 VDD.n4723 VDD.n4722 46.2524
R1137 VDD.n1778 VDD.n1727 46.2524
R1138 VDD.n4696 VDD.n1797 46.2524
R1139 VDD.n4676 VDD.n1838 46.2524
R1140 VDD.n4674 VDD.n1839 46.2524
R1141 VDD.n4654 VDD.n1880 46.2524
R1142 VDD.n4652 VDD.n1881 46.2524
R1143 VDD.n4629 VDD.n4628 46.2524
R1144 VDD.n1977 VDD.n1927 46.2524
R1145 VDD.n1989 VDD.n1972 46.2524
R1146 VDD.n4602 VDD.n4601 46.2524
R1147 VDD.n2042 VDD.n1991 46.2524
R1148 VDD.n4575 VDD.n2061 46.2524
R1149 VDD.n4555 VDD.n2102 46.2524
R1150 VDD.n4553 VDD.n2103 46.2524
R1151 VDD.n4533 VDD.n2144 46.2524
R1152 VDD.n4531 VDD.n2145 46.2524
R1153 VDD.n4508 VDD.n4507 46.2524
R1154 VDD.n2241 VDD.n2191 46.2524
R1155 VDD.n2253 VDD.n2236 46.2524
R1156 VDD.n4481 VDD.n4480 46.2524
R1157 VDD.n2306 VDD.n2255 46.2524
R1158 VDD.n4454 VDD.n2325 46.2524
R1159 VDD.n4434 VDD.n2366 46.2524
R1160 VDD.n4432 VDD.n2367 46.2524
R1161 VDD.n4412 VDD.n2408 46.2524
R1162 VDD.n4410 VDD.n2409 46.2524
R1163 VDD VDD.t32 44.7841
R1164 VDD.t23 VDD 44.7841
R1165 VDD.n2563 VDD.t58 43.1378
R1166 VDD.n6127 VDD.t50 41.9684
R1167 VDD.n3013 VDD 41.8475
R1168 VDD.n3279 VDD 41.8475
R1169 VDD.n3545 VDD 41.8475
R1170 VDD.n1661 VDD 41.8475
R1171 VDD.n1925 VDD 41.8475
R1172 VDD.n2189 VDD 41.8475
R1173 VDD.n2622 VDD.t44 41.177
R1174 VDD.t46 VDD.n6096 40.0607
R1175 VDD.n6147 VDD 39.1069
R1176 VDD.n6124 VDD.n604 39.0005
R1177 VDD.n7270 VDD.n7269 39.0005
R1178 VDD.n3824 VDD.t4 37.4425
R1179 VDD.n2562 VDD.n2561 37.3561
R1180 VDD.n6097 VDD.t46 36.2455
R1181 VDD.n2599 VDD.n2486 36.0005
R1182 VDD.n4970 VDD.n1239 36.0005
R1183 VDD.n6391 VDD.n6390 33.746
R1184 VDD.n6617 VDD.n6616 33.746
R1185 VDD.n6843 VDD.n6842 33.746
R1186 VDD.n1659 VDD.n1658 33.746
R1187 VDD.n1923 VDD.n1922 33.746
R1188 VDD.n2187 VDD.n2186 33.746
R1189 VDD.n3011 VDD.n3010 33.746
R1190 VDD.n3277 VDD.n3276 33.746
R1191 VDD.n3543 VDD.n3542 33.746
R1192 VDD.n5249 VDD.n5248 33.746
R1193 VDD.n5477 VDD.n5476 33.746
R1194 VDD.n5705 VDD.n5704 33.746
R1195 VDD.n7272 VDD.n7271 33.6517
R1196 VDD.n515 VDD.n508 32.9702
R1197 VDD.n381 VDD.n374 32.9702
R1198 VDD.n247 VDD.n240 32.9702
R1199 VDD.n113 VDD.n106 32.9702
R1200 VDD.n1521 VDD.n1518 32.9702
R1201 VDD.n1785 VDD.n1782 32.9702
R1202 VDD.n2049 VDD.n2046 32.9702
R1203 VDD.n2313 VDD.n2310 32.9702
R1204 VDD.n4280 VDD.n2846 32.9702
R1205 VDD.n3137 VDD.n3134 32.9702
R1206 VDD.n3403 VDD.n3400 32.9702
R1207 VDD.n3669 VDD.n3666 32.9702
R1208 VDD.n1147 VDD.n1131 32.9702
R1209 VDD.n1012 VDD.n996 32.9702
R1210 VDD.n877 VDD.n861 32.9702
R1211 VDD.n742 VDD.n735 32.9702
R1212 VDD.n4969 VDD.n4968 31.0632
R1213 VDD.n6076 VDD.n638 29.4128
R1214 VDD.n7226 VDD.n9 29.4128
R1215 VDD.n2626 VDD.n2625 29.2586
R1216 VDD.n4930 VDD.n1241 29.2586
R1217 VDD.t56 VDD.n2711 28.6326
R1218 VDD.t41 VDD.n2837 28.6326
R1219 VDD.n4276 VDD.t68 28.6326
R1220 VDD.t64 VDD.n3147 28.6326
R1221 VDD.n4157 VDD.t74 28.6326
R1222 VDD.t69 VDD.n3413 28.6326
R1223 VDD.n4038 VDD.t70 28.6326
R1224 VDD.t73 VDD.n3679 28.6326
R1225 VDD.n3919 VDD.t2 28.6326
R1226 VDD.t31 VDD.n1392 28.6326
R1227 VDD.t66 VDD.n1531 28.6326
R1228 VDD.n4819 VDD.t67 28.6326
R1229 VDD.t20 VDD.n1795 28.6326
R1230 VDD.n4698 VDD.t53 28.6326
R1231 VDD.t72 VDD.n2059 28.6326
R1232 VDD.n4577 VDD.t38 28.6326
R1233 VDD.t28 VDD.n2323 28.6326
R1234 VDD.n4456 VDD.t65 28.6326
R1235 VDD.n6096 VDD 28.615
R1236 VDD.n6978 VDD.n6977 28.2358
R1237 VDD.n7016 VDD.n7014 28.2358
R1238 VDD.n7070 VDD.n45 28.2358
R1239 VDD.n6960 VDD.n6959 28.2358
R1240 VDD.n6752 VDD.n6751 28.2358
R1241 VDD.n6790 VDD.n6788 28.2358
R1242 VDD.n6839 VDD.n180 28.2358
R1243 VDD.n6734 VDD.n6733 28.2358
R1244 VDD.n6526 VDD.n6525 28.2358
R1245 VDD.n6564 VDD.n6562 28.2358
R1246 VDD.n6613 VDD.n314 28.2358
R1247 VDD.n6508 VDD.n6507 28.2358
R1248 VDD.n6300 VDD.n6299 28.2358
R1249 VDD.n6338 VDD.n6336 28.2358
R1250 VDD.n6387 VDD.n448 28.2358
R1251 VDD.n6194 VDD.n6193 28.2358
R1252 VDD.n6282 VDD.n6281 28.2358
R1253 VDD.n26 VDD.n13 28.2358
R1254 VDD.n7116 VDD.n19 28.2358
R1255 VDD.n7193 VDD.n15 28.2358
R1256 VDD.n7165 VDD.n7164 28.2358
R1257 VDD.n655 VDD.n642 28.2358
R1258 VDD.n5966 VDD.n648 28.2358
R1259 VDD.n6043 VDD.n644 28.2358
R1260 VDD.n6015 VDD.n6014 28.2358
R1261 VDD.n5850 VDD.n5849 28.2358
R1262 VDD.n5886 VDD.n5884 28.2358
R1263 VDD.n5756 VDD.n771 28.2358
R1264 VDD.n5789 VDD.n5787 28.2358
R1265 VDD.n5613 VDD.n5611 28.2358
R1266 VDD.n5664 VDD.n812 28.2358
R1267 VDD.n5703 VDD.n5702 28.2358
R1268 VDD.n5528 VDD.n906 28.2358
R1269 VDD.n5561 VDD.n5559 28.2358
R1270 VDD.n5385 VDD.n5383 28.2358
R1271 VDD.n5436 VDD.n947 28.2358
R1272 VDD.n5475 VDD.n5474 28.2358
R1273 VDD.n5300 VDD.n1041 28.2358
R1274 VDD.n5333 VDD.n5331 28.2358
R1275 VDD.n5157 VDD.n5155 28.2358
R1276 VDD.n5208 VDD.n1082 28.2358
R1277 VDD.n5247 VDD.n5246 28.2358
R1278 VDD.n5072 VDD.n1176 28.2358
R1279 VDD.n5105 VDD.n5103 28.2358
R1280 VDD.n4928 VDD.n1243 28.2358
R1281 VDD.n4920 VDD.n1246 28.2358
R1282 VDD.n1324 VDD.n1321 28.2358
R1283 VDD.n1333 VDD.n1315 28.2358
R1284 VDD.n4893 VDD.n1316 28.2358
R1285 VDD.n1387 VDD.n1384 28.2358
R1286 VDD.n4453 VDD.n2302 28.2358
R1287 VDD.n2364 VDD.n2352 28.2358
R1288 VDD.n4431 VDD.n2353 28.2358
R1289 VDD.n2406 VDD.n2394 28.2358
R1290 VDD.n4409 VDD.n2395 28.2358
R1291 VDD.n2188 VDD.n2178 28.2358
R1292 VDD.n4505 VDD.n2179 28.2358
R1293 VDD.n2243 VDD.n2240 28.2358
R1294 VDD.n2252 VDD.n2234 28.2358
R1295 VDD.n4478 VDD.n2235 28.2358
R1296 VDD.n2307 VDD.n2304 28.2358
R1297 VDD.n4574 VDD.n2038 28.2358
R1298 VDD.n2100 VDD.n2088 28.2358
R1299 VDD.n4552 VDD.n2089 28.2358
R1300 VDD.n2142 VDD.n2130 28.2358
R1301 VDD.n4530 VDD.n2131 28.2358
R1302 VDD.n2185 VDD.n2182 28.2358
R1303 VDD.n1924 VDD.n1914 28.2358
R1304 VDD.n4626 VDD.n1915 28.2358
R1305 VDD.n1979 VDD.n1976 28.2358
R1306 VDD.n1988 VDD.n1970 28.2358
R1307 VDD.n4599 VDD.n1971 28.2358
R1308 VDD.n2043 VDD.n2040 28.2358
R1309 VDD.n4695 VDD.n1774 28.2358
R1310 VDD.n1836 VDD.n1824 28.2358
R1311 VDD.n4673 VDD.n1825 28.2358
R1312 VDD.n1878 VDD.n1866 28.2358
R1313 VDD.n4651 VDD.n1867 28.2358
R1314 VDD.n1921 VDD.n1918 28.2358
R1315 VDD.n1660 VDD.n1650 28.2358
R1316 VDD.n4747 VDD.n1651 28.2358
R1317 VDD.n1715 VDD.n1712 28.2358
R1318 VDD.n1724 VDD.n1706 28.2358
R1319 VDD.n4720 VDD.n1707 28.2358
R1320 VDD.n1779 VDD.n1776 28.2358
R1321 VDD.n4816 VDD.n1510 28.2358
R1322 VDD.n1572 VDD.n1560 28.2358
R1323 VDD.n4794 VDD.n1561 28.2358
R1324 VDD.n1614 VDD.n1602 28.2358
R1325 VDD.n4772 VDD.n1603 28.2358
R1326 VDD.n1657 VDD.n1654 28.2358
R1327 VDD.n4868 VDD.n1382 28.2358
R1328 VDD.n1451 VDD.n1448 28.2358
R1329 VDD.n1460 VDD.n1442 28.2358
R1330 VDD.n4841 VDD.n1443 28.2358
R1331 VDD.n1515 VDD.n1512 28.2358
R1332 VDD.n2629 VDD.n2454 28.2358
R1333 VDD.n2639 VDD.n2447 28.2358
R1334 VDD.n4370 VDD.n2448 28.2358
R1335 VDD.n2699 VDD.n2696 28.2358
R1336 VDD.n2708 VDD.n2690 28.2358
R1337 VDD.n4343 VDD.n2691 28.2358
R1338 VDD.n3916 VDD.n3658 28.2358
R1339 VDD.n3721 VDD.n3710 28.2358
R1340 VDD.n3895 VDD.n3711 28.2358
R1341 VDD.n3764 VDD.n3753 28.2358
R1342 VDD.n3874 VDD.n3754 28.2358
R1343 VDD.n3544 VDD.n3534 28.2358
R1344 VDD.n3968 VDD.n3535 28.2358
R1345 VDD.n3599 VDD.n3596 28.2358
R1346 VDD.n3608 VDD.n3590 28.2358
R1347 VDD.n3941 VDD.n3591 28.2358
R1348 VDD.n3663 VDD.n3660 28.2358
R1349 VDD.n4035 VDD.n3392 28.2358
R1350 VDD.n3455 VDD.n3444 28.2358
R1351 VDD.n4014 VDD.n3445 28.2358
R1352 VDD.n3498 VDD.n3487 28.2358
R1353 VDD.n3993 VDD.n3488 28.2358
R1354 VDD.n3541 VDD.n3538 28.2358
R1355 VDD.n3278 VDD.n3268 28.2358
R1356 VDD.n4087 VDD.n3269 28.2358
R1357 VDD.n3333 VDD.n3330 28.2358
R1358 VDD.n3342 VDD.n3324 28.2358
R1359 VDD.n4060 VDD.n3325 28.2358
R1360 VDD.n3397 VDD.n3394 28.2358
R1361 VDD.n4154 VDD.n3126 28.2358
R1362 VDD.n3189 VDD.n3178 28.2358
R1363 VDD.n4133 VDD.n3179 28.2358
R1364 VDD.n3232 VDD.n3221 28.2358
R1365 VDD.n4112 VDD.n3222 28.2358
R1366 VDD.n3275 VDD.n3272 28.2358
R1367 VDD.n3012 VDD.n3002 28.2358
R1368 VDD.n4206 VDD.n3003 28.2358
R1369 VDD.n3067 VDD.n3064 28.2358
R1370 VDD.n3076 VDD.n3058 28.2358
R1371 VDD.n4179 VDD.n3059 28.2358
R1372 VDD.n3131 VDD.n3128 28.2358
R1373 VDD.n4273 VDD.n2849 28.2358
R1374 VDD.n2923 VDD.n2912 28.2358
R1375 VDD.n4252 VDD.n2913 28.2358
R1376 VDD.n2966 VDD.n2955 28.2358
R1377 VDD.n4231 VDD.n2956 28.2358
R1378 VDD.n3009 VDD.n3006 28.2358
R1379 VDD.n2770 VDD.n2755 28.2358
R1380 VDD.n4317 VDD.n2756 28.2358
R1381 VDD.n2825 VDD.n2822 28.2358
R1382 VDD.n2834 VDD.n2816 28.2358
R1383 VDD.n4290 VDD.n2817 28.2358
R1384 VDD VDD.n2563 27.4515
R1385 VDD.n6093 VDD.n631 27.3454
R1386 VDD.n2476 VDD.n2456 27.1422
R1387 VDD.n4958 VDD.n4954 27.1422
R1388 VDD.n3823 VDD.n3808 25.696
R1389 VDD.n2541 VDD.n2540 25.696
R1390 VDD.n2601 VDD.n2600 23.0907
R1391 VDD.n4972 VDD.n4971 23.0907
R1392 VDD.n6122 VDD.n603 22.8875
R1393 VDD.t62 VDD.t26 21.1252
R1394 VDD.t18 VDD.t10 21.1252
R1395 VDD.n3808 VDD.n3807 20.7428
R1396 VDD.n3825 VDD.n3811 20.7428
R1397 VDD.n3824 VDD.n3817 20.7428
R1398 VDD.n3824 VDD.n3814 20.7428
R1399 VDD.n3826 VDD.n3825 20.7428
R1400 VDD.n2594 VDD.n2593 20.7428
R1401 VDD.n2594 VDD.n2566 20.7428
R1402 VDD.n2594 VDD.n2565 20.7428
R1403 VDD.n2550 VDD.n2487 20.7428
R1404 VDD.n2561 VDD.n2560 20.7428
R1405 VDD.n2561 VDD.n2488 20.7428
R1406 VDD.n2502 VDD.n2487 20.7428
R1407 VDD.n2542 VDD.n2541 20.7428
R1408 VDD.n1218 VDD.n1217 20.7428
R1409 VDD.n4989 VDD.n4988 20.7428
R1410 VDD.n5002 VDD.n5000 20.7428
R1411 VDD.n4999 VDD.n4997 20.7428
R1412 VDD.n5010 VDD.n1203 20.7428
R1413 VDD.n6099 VDD.n6097 20.7428
R1414 VDD.n623 VDD.n619 20.7428
R1415 VDD.n6107 VDD.n619 20.7428
R1416 VDD.n6171 VDD.n573 20.7428
R1417 VDD.n588 VDD.n587 20.7428
R1418 VDD.n6146 VDD.n6145 20.7428
R1419 VDD.n6163 VDD.n6161 20.7428
R1420 VDD.n6160 VDD.n6154 20.7428
R1421 VDD.t68 VDD.n2850 20.3031
R1422 VDD.t74 VDD.n3148 20.3031
R1423 VDD.t70 VDD.n3414 20.3031
R1424 VDD.t2 VDD.n3680 20.3031
R1425 VDD.t67 VDD.n1532 20.3031
R1426 VDD.t53 VDD.n1796 20.3031
R1427 VDD.t38 VDD.n2060 20.3031
R1428 VDD.t65 VDD.n2324 20.3031
R1429 VDD.t16 VDD.n1218 18.5229
R1430 VDD.t71 VDD.n588 18.5229
R1431 VDD VDD.t8 16.5329
R1432 VDD VDD.t1 16.5329
R1433 VDD.n2472 VDD 15.4887
R1434 VDD.n1235 VDD 15.4887
R1435 VDD.n6131 VDD.n6130 15.4666
R1436 VDD.n7255 VDD.n7254 15.4666
R1437 VDD VDD.n630 15.1421
R1438 VDD VDD.n0 15.1421
R1439 VDD.n2619 VDD.n2618 15.12
R1440 VDD.n4956 VDD.n4955 15.12
R1441 VDD.n2486 VDD.n2455 15.0005
R1442 VDD.n4966 VDD.n1239 15.0005
R1443 VDD.n2625 VDD.n2624 13.7917
R1444 VDD.n1267 VDD.n1241 13.7917
R1445 VDD.n6077 VDD.n6076 13.3673
R1446 VDD.n7227 VDD.n7226 13.3673
R1447 VDD.n6981 VDD.n6980 13.1177
R1448 VDD.n7045 VDD.n7044 13.1177
R1449 VDD.n6871 VDD.n152 13.1177
R1450 VDD.n6892 VDD.n137 13.1177
R1451 VDD.n6921 VDD.n6920 13.1177
R1452 VDD.n6941 VDD.n6940 13.1177
R1453 VDD.n6755 VDD.n6754 13.1177
R1454 VDD.n6819 VDD.n6818 13.1177
R1455 VDD.n6845 VDD.n6844 13.1177
R1456 VDD.n6645 VDD.n286 13.1177
R1457 VDD.n6666 VDD.n271 13.1177
R1458 VDD.n6695 VDD.n6694 13.1177
R1459 VDD.n6715 VDD.n6714 13.1177
R1460 VDD.n6529 VDD.n6528 13.1177
R1461 VDD.n6593 VDD.n6592 13.1177
R1462 VDD.n6619 VDD.n6618 13.1177
R1463 VDD.n6419 VDD.n420 13.1177
R1464 VDD.n6440 VDD.n405 13.1177
R1465 VDD.n6469 VDD.n6468 13.1177
R1466 VDD.n6489 VDD.n6488 13.1177
R1467 VDD.n6303 VDD.n6302 13.1177
R1468 VDD.n6367 VDD.n6366 13.1177
R1469 VDD.n6393 VDD.n6392 13.1177
R1470 VDD.n6214 VDD.n539 13.1177
R1471 VDD.n6243 VDD.n6242 13.1177
R1472 VDD.n6263 VDD.n6262 13.1177
R1473 VDD.n7218 VDD.n21 13.1177
R1474 VDD.n6068 VDD.n650 13.1177
R1475 VDD.n5826 VDD.n715 13.1177
R1476 VDD.n713 VDD.n712 13.1177
R1477 VDD.n5919 VDD.n5918 13.1177
R1478 VDD.n5726 VDD.n5725 13.1177
R1479 VDD.n5760 VDD.n5759 13.1177
R1480 VDD.n5808 VDD.n5807 13.1177
R1481 VDD.n866 VDD.n846 13.1177
R1482 VDD.n5642 VDD.n5641 13.1177
R1483 VDD.n5668 VDD.n5667 13.1177
R1484 VDD.n5498 VDD.n5497 13.1177
R1485 VDD.n5532 VDD.n5531 13.1177
R1486 VDD.n5581 VDD.n5580 13.1177
R1487 VDD.n1001 VDD.n981 13.1177
R1488 VDD.n5414 VDD.n5413 13.1177
R1489 VDD.n5440 VDD.n5439 13.1177
R1490 VDD.n5270 VDD.n5269 13.1177
R1491 VDD.n5304 VDD.n5303 13.1177
R1492 VDD.n5353 VDD.n5352 13.1177
R1493 VDD.n1136 VDD.n1116 13.1177
R1494 VDD.n5186 VDD.n5185 13.1177
R1495 VDD.n5212 VDD.n5211 13.1177
R1496 VDD.n5042 VDD.n5041 13.1177
R1497 VDD.n5076 VDD.n5075 13.1177
R1498 VDD.n5125 VDD.n5124 13.1177
R1499 VDD.n5043 VDD.n5042 13.1177
R1500 VDD.n5075 VDD.n1160 13.1177
R1501 VDD.n5271 VDD.n5270 13.1177
R1502 VDD.n5303 VDD.n1025 13.1177
R1503 VDD.n5499 VDD.n5498 13.1177
R1504 VDD.n5531 VDD.n890 13.1177
R1505 VDD.n5727 VDD.n5726 13.1177
R1506 VDD.n5759 VDD.n755 13.1177
R1507 VDD.n5920 VDD.n5919 13.1177
R1508 VDD.n712 VDD.n695 13.1177
R1509 VDD.n5827 VDD.n5826 13.1177
R1510 VDD.n5809 VDD.n5808 13.1177
R1511 VDD.n5707 VDD.n5706 13.1177
R1512 VDD.n5667 VDD.n795 13.1177
R1513 VDD.n5643 VDD.n5642 13.1177
R1514 VDD.n867 VDD.n866 13.1177
R1515 VDD.n5582 VDD.n5581 13.1177
R1516 VDD.n5479 VDD.n5478 13.1177
R1517 VDD.n5439 VDD.n930 13.1177
R1518 VDD.n5415 VDD.n5414 13.1177
R1519 VDD.n1002 VDD.n1001 13.1177
R1520 VDD.n5354 VDD.n5353 13.1177
R1521 VDD.n5251 VDD.n5250 13.1177
R1522 VDD.n5211 VDD.n1065 13.1177
R1523 VDD.n5187 VDD.n5186 13.1177
R1524 VDD.n1137 VDD.n1136 13.1177
R1525 VDD.n5126 VDD.n5125 13.1177
R1526 VDD.n6074 VDD.n640 13.1177
R1527 VDD.n651 VDD.n650 13.1177
R1528 VDD.n7224 VDD.n11 13.1177
R1529 VDD.n22 VDD.n21 13.1177
R1530 VDD.n6302 VDD.n478 13.1177
R1531 VDD.n6368 VDD.n6367 13.1177
R1532 VDD.n6528 VDD.n344 13.1177
R1533 VDD.n6594 VDD.n6593 13.1177
R1534 VDD.n6754 VDD.n210 13.1177
R1535 VDD.n6820 VDD.n6819 13.1177
R1536 VDD.n6980 VDD.n76 13.1177
R1537 VDD.n7046 VDD.n7045 13.1177
R1538 VDD.n6940 VDD.n6939 13.1177
R1539 VDD.n6920 VDD.n6919 13.1177
R1540 VDD.n6893 VDD.n6892 13.1177
R1541 VDD.n6872 VDD.n6871 13.1177
R1542 VDD.n6841 VDD.n163 13.1177
R1543 VDD.n6714 VDD.n6713 13.1177
R1544 VDD.n6694 VDD.n6693 13.1177
R1545 VDD.n6667 VDD.n6666 13.1177
R1546 VDD.n6646 VDD.n6645 13.1177
R1547 VDD.n6615 VDD.n297 13.1177
R1548 VDD.n6488 VDD.n6487 13.1177
R1549 VDD.n6468 VDD.n6467 13.1177
R1550 VDD.n6441 VDD.n6440 13.1177
R1551 VDD.n6420 VDD.n6419 13.1177
R1552 VDD.n6389 VDD.n431 13.1177
R1553 VDD.n6262 VDD.n6261 13.1177
R1554 VDD.n6242 VDD.n6241 13.1177
R1555 VDD.n6215 VDD.n6214 13.1177
R1556 VDD.n3821 VDD.n3819 13.0163
R1557 VDD.n2761 VDD.n2758 13.0163
R1558 VDD.n2538 VDD.n2536 13.0163
R1559 VDD.n1381 VDD.n1379 13.0163
R1560 VDD.n4968 VDD.n4967 12.9433
R1561 VDD.t17 VDD.n4999 12.5529
R1562 VDD.t40 VDD.n6160 12.5529
R1563 VDD.n2627 VDD.n2626 12.4812
R1564 VDD.n4930 VDD.n4929 12.4812
R1565 VDD.n6126 VDD.n6125 12.4001
R1566 VDD.n6124 VDD.n606 12.0005
R1567 VDD.n7274 VDD.n7270 12.0005
R1568 VDD.n6129 VDD.n603 11.9758
R1569 VDD.n2601 VDD.n2473 11.9758
R1570 VDD.n4972 VDD.n1236 11.9758
R1571 VDD.n2598 VDD.n2597 11.7652
R1572 VDD.n2628 VDD.n2627 11.747
R1573 VDD.n2641 VDD.n2640 11.747
R1574 VDD.n4372 VDD.n4371 11.747
R1575 VDD.n2698 VDD.n2697 11.747
R1576 VDD.n2710 VDD.n2709 11.747
R1577 VDD.n4345 VDD.n4344 11.747
R1578 VDD.n2760 VDD.n2759 11.747
R1579 VDD.n2772 VDD.n2771 11.747
R1580 VDD.n4319 VDD.n4318 11.747
R1581 VDD.n2824 VDD.n2823 11.747
R1582 VDD.n2836 VDD.n2835 11.747
R1583 VDD.n4292 VDD.n4291 11.747
R1584 VDD.n4275 VDD.n4274 11.747
R1585 VDD.n2925 VDD.n2924 11.747
R1586 VDD.n4254 VDD.n4253 11.747
R1587 VDD.n2968 VDD.n2967 11.747
R1588 VDD.n4233 VDD.n4232 11.747
R1589 VDD.n3008 VDD.n3007 11.747
R1590 VDD.n3014 VDD.n3013 11.747
R1591 VDD.n4208 VDD.n4207 11.747
R1592 VDD.n3066 VDD.n3065 11.747
R1593 VDD.n3078 VDD.n3077 11.747
R1594 VDD.n4181 VDD.n4180 11.747
R1595 VDD.n3130 VDD.n3127 11.747
R1596 VDD.n4156 VDD.n4155 11.747
R1597 VDD.n3191 VDD.n3190 11.747
R1598 VDD.n4135 VDD.n4134 11.747
R1599 VDD.n3234 VDD.n3233 11.747
R1600 VDD.n4114 VDD.n4113 11.747
R1601 VDD.n3274 VDD.n3273 11.747
R1602 VDD.n3280 VDD.n3279 11.747
R1603 VDD.n4089 VDD.n4088 11.747
R1604 VDD.n3332 VDD.n3331 11.747
R1605 VDD.n3344 VDD.n3343 11.747
R1606 VDD.n4062 VDD.n4061 11.747
R1607 VDD.n3396 VDD.n3393 11.747
R1608 VDD.n4037 VDD.n4036 11.747
R1609 VDD.n3457 VDD.n3456 11.747
R1610 VDD.n4016 VDD.n4015 11.747
R1611 VDD.n3500 VDD.n3499 11.747
R1612 VDD.n3995 VDD.n3994 11.747
R1613 VDD.n3540 VDD.n3539 11.747
R1614 VDD.n3546 VDD.n3545 11.747
R1615 VDD.n3970 VDD.n3969 11.747
R1616 VDD.n3598 VDD.n3597 11.747
R1617 VDD.n3610 VDD.n3609 11.747
R1618 VDD.n3943 VDD.n3942 11.747
R1619 VDD.n3662 VDD.n3659 11.747
R1620 VDD.n3918 VDD.n3917 11.747
R1621 VDD.n3723 VDD.n3722 11.747
R1622 VDD.n3897 VDD.n3896 11.747
R1623 VDD.n3766 VDD.n3765 11.747
R1624 VDD.n3876 VDD.n3875 11.747
R1625 VDD.n3822 VDD.n3818 11.747
R1626 VDD.n4929 VDD.n1242 11.747
R1627 VDD.n4922 VDD.n4921 11.747
R1628 VDD.n1323 VDD.n1322 11.747
R1629 VDD.n1335 VDD.n1334 11.747
R1630 VDD.n4895 VDD.n4894 11.747
R1631 VDD.n1386 VDD.n1383 11.747
R1632 VDD.n1394 VDD.n1393 11.747
R1633 VDD.n4870 VDD.n4869 11.747
R1634 VDD.n1450 VDD.n1449 11.747
R1635 VDD.n1462 VDD.n1461 11.747
R1636 VDD.n4843 VDD.n4842 11.747
R1637 VDD.n1514 VDD.n1511 11.747
R1638 VDD.n4818 VDD.n4817 11.747
R1639 VDD.n1574 VDD.n1573 11.747
R1640 VDD.n4796 VDD.n4795 11.747
R1641 VDD.n1616 VDD.n1615 11.747
R1642 VDD.n4774 VDD.n4773 11.747
R1643 VDD.n1656 VDD.n1655 11.747
R1644 VDD.n1662 VDD.n1661 11.747
R1645 VDD.n4749 VDD.n4748 11.747
R1646 VDD.n1714 VDD.n1713 11.747
R1647 VDD.n1726 VDD.n1725 11.747
R1648 VDD.n4722 VDD.n4721 11.747
R1649 VDD.n1778 VDD.n1775 11.747
R1650 VDD.n4697 VDD.n4696 11.747
R1651 VDD.n1838 VDD.n1837 11.747
R1652 VDD.n4675 VDD.n4674 11.747
R1653 VDD.n1880 VDD.n1879 11.747
R1654 VDD.n4653 VDD.n4652 11.747
R1655 VDD.n1920 VDD.n1919 11.747
R1656 VDD.n1926 VDD.n1925 11.747
R1657 VDD.n4628 VDD.n4627 11.747
R1658 VDD.n1978 VDD.n1977 11.747
R1659 VDD.n1990 VDD.n1989 11.747
R1660 VDD.n4601 VDD.n4600 11.747
R1661 VDD.n2042 VDD.n2039 11.747
R1662 VDD.n4576 VDD.n4575 11.747
R1663 VDD.n2102 VDD.n2101 11.747
R1664 VDD.n4554 VDD.n4553 11.747
R1665 VDD.n2144 VDD.n2143 11.747
R1666 VDD.n4532 VDD.n4531 11.747
R1667 VDD.n2184 VDD.n2183 11.747
R1668 VDD.n2190 VDD.n2189 11.747
R1669 VDD.n4507 VDD.n4506 11.747
R1670 VDD.n2242 VDD.n2241 11.747
R1671 VDD.n2254 VDD.n2253 11.747
R1672 VDD.n4480 VDD.n4479 11.747
R1673 VDD.n2306 VDD.n2303 11.747
R1674 VDD.n4455 VDD.n4454 11.747
R1675 VDD.n2366 VDD.n2365 11.747
R1676 VDD.n4433 VDD.n4432 11.747
R1677 VDD.n2408 VDD.n2407 11.747
R1678 VDD.n4411 VDD.n4410 11.747
R1679 VDD.n2539 VDD.n2535 11.747
R1680 VDD.n7072 VDD.n7071 11.5452
R1681 VDD.n6192 VDD.n6191 11.5452
R1682 VDD.n5000 VDD.t17 11.4813
R1683 VDD.n6161 VDD.t40 11.4813
R1684 VDD.n6094 VDD.n6093 11.2229
R1685 VDD.n2620 VDD.n2456 11.2229
R1686 VDD.n4958 VDD.n4957 11.2229
R1687 VDD.n6097 VDD.n619 10.4925
R1688 VDD.n7273 VDD.n7272 10.3547
R1689 VDD.n5000 VDD.t9 9.64439
R1690 VDD.n6161 VDD.t57 9.64439
R1691 VDD.n6976 VDD.n6975 9.38471
R1692 VDD.n6962 VDD.n6961 9.38471
R1693 VDD.n6750 VDD.n6749 9.38471
R1694 VDD.n6736 VDD.n6735 9.38471
R1695 VDD.n6524 VDD.n6523 9.38471
R1696 VDD.n6510 VDD.n6509 9.38471
R1697 VDD.n6298 VDD.n6297 9.38471
R1698 VDD.n6284 VDD.n6283 9.38471
R1699 VDD.n6023 VDD.n6022 9.3005
R1700 VDD.n6041 VDD.n6040 9.3005
R1701 VDD.n5969 VDD.n5955 9.3005
R1702 VDD.n5933 VDD.n653 9.3005
R1703 VDD.n5960 VDD.n5959 9.3005
R1704 VDD.n6089 VDD.n631 9.3005
R1705 VDD.n515 VDD.n514 9.3005
R1706 VDD.n6385 VDD.n6384 9.3005
R1707 VDD.n6341 VDD.n6340 9.3005
R1708 VDD.n6308 VDD.n6307 9.3005
R1709 VDD.n509 VDD.n508 9.3005
R1710 VDD.n480 VDD.n479 9.3005
R1711 VDD.n465 VDD.n464 9.3005
R1712 VDD.n381 VDD.n380 9.3005
R1713 VDD.n6611 VDD.n6610 9.3005
R1714 VDD.n6567 VDD.n6566 9.3005
R1715 VDD.n6534 VDD.n6533 9.3005
R1716 VDD.n375 VDD.n374 9.3005
R1717 VDD.n346 VDD.n345 9.3005
R1718 VDD.n331 VDD.n330 9.3005
R1719 VDD.n247 VDD.n246 9.3005
R1720 VDD.n6837 VDD.n6836 9.3005
R1721 VDD.n6793 VDD.n6792 9.3005
R1722 VDD.n6760 VDD.n6759 9.3005
R1723 VDD.n241 VDD.n240 9.3005
R1724 VDD.n212 VDD.n211 9.3005
R1725 VDD.n197 VDD.n196 9.3005
R1726 VDD.n113 VDD.n112 9.3005
R1727 VDD.n7068 VDD.n7067 9.3005
R1728 VDD.n7019 VDD.n7018 9.3005
R1729 VDD.n6986 VDD.n6985 9.3005
R1730 VDD.n107 VDD.n106 9.3005
R1731 VDD.n78 VDD.n77 9.3005
R1732 VDD.n63 VDD.n62 9.3005
R1733 VDD.n6957 VDD.n6956 9.3005
R1734 VDD.n6937 VDD.n6936 9.3005
R1735 VDD.n143 VDD.n142 9.3005
R1736 VDD.n6896 VDD.n6895 9.3005
R1737 VDD.n6875 VDD.n6874 9.3005
R1738 VDD.n6731 VDD.n6730 9.3005
R1739 VDD.n6711 VDD.n6710 9.3005
R1740 VDD.n277 VDD.n276 9.3005
R1741 VDD.n6670 VDD.n6669 9.3005
R1742 VDD.n6649 VDD.n6648 9.3005
R1743 VDD.n6505 VDD.n6504 9.3005
R1744 VDD.n6485 VDD.n6484 9.3005
R1745 VDD.n411 VDD.n410 9.3005
R1746 VDD.n6444 VDD.n6443 9.3005
R1747 VDD.n6423 VDD.n6422 9.3005
R1748 VDD.n6279 VDD.n6278 9.3005
R1749 VDD.n6259 VDD.n6258 9.3005
R1750 VDD.n545 VDD.n544 9.3005
R1751 VDD.n6197 VDD.n6196 9.3005
R1752 VDD.n6218 VDD.n6217 9.3005
R1753 VDD.n7083 VDD.n24 9.3005
R1754 VDD.n7110 VDD.n7109 9.3005
R1755 VDD.n7119 VDD.n7105 9.3005
R1756 VDD.n7191 VDD.n7190 9.3005
R1757 VDD.n7173 VDD.n7172 9.3005
R1758 VDD.n2637 VDD.n2636 9.3005
R1759 VDD.n2664 VDD.n2663 9.3005
R1760 VDD.n2694 VDD.n2648 9.3005
R1761 VDD.n2706 VDD.n2705 9.3005
R1762 VDD.n2727 VDD.n2726 9.3005
R1763 VDD.n1519 VDD.n1518 9.3005
R1764 VDD.n1522 VDD.n1521 9.3005
R1765 VDD.n4770 VDD.n4769 9.3005
R1766 VDD.n1783 VDD.n1782 9.3005
R1767 VDD.n1786 VDD.n1785 9.3005
R1768 VDD.n4649 VDD.n4648 9.3005
R1769 VDD.n2047 VDD.n2046 9.3005
R1770 VDD.n2050 VDD.n2049 9.3005
R1771 VDD.n4528 VDD.n4527 9.3005
R1772 VDD.n2311 VDD.n2310 9.3005
R1773 VDD.n2314 VDD.n2313 9.3005
R1774 VDD.n4407 VDD.n4406 9.3005
R1775 VDD.n2403 VDD.n2402 9.3005
R1776 VDD.n4429 VDD.n4428 9.3005
R1777 VDD.n2361 VDD.n2360 9.3005
R1778 VDD.n4451 VDD.n4450 9.3005
R1779 VDD.n2305 VDD.n2261 9.3005
R1780 VDD.n2277 VDD.n2276 9.3005
R1781 VDD.n2250 VDD.n2249 9.3005
R1782 VDD.n2238 VDD.n2197 9.3005
R1783 VDD.n2208 VDD.n2207 9.3005
R1784 VDD.n2139 VDD.n2138 9.3005
R1785 VDD.n4550 VDD.n4549 9.3005
R1786 VDD.n2097 VDD.n2096 9.3005
R1787 VDD.n4572 VDD.n4571 9.3005
R1788 VDD.n2041 VDD.n1997 9.3005
R1789 VDD.n2013 VDD.n2012 9.3005
R1790 VDD.n1986 VDD.n1985 9.3005
R1791 VDD.n1974 VDD.n1933 9.3005
R1792 VDD.n1944 VDD.n1943 9.3005
R1793 VDD.n1875 VDD.n1874 9.3005
R1794 VDD.n4671 VDD.n4670 9.3005
R1795 VDD.n1833 VDD.n1832 9.3005
R1796 VDD.n4693 VDD.n4692 9.3005
R1797 VDD.n1777 VDD.n1733 9.3005
R1798 VDD.n1749 VDD.n1748 9.3005
R1799 VDD.n1722 VDD.n1721 9.3005
R1800 VDD.n1710 VDD.n1669 9.3005
R1801 VDD.n1680 VDD.n1679 9.3005
R1802 VDD.n1611 VDD.n1610 9.3005
R1803 VDD.n4792 VDD.n4791 9.3005
R1804 VDD.n1569 VDD.n1568 9.3005
R1805 VDD.n4814 VDD.n4813 9.3005
R1806 VDD.n1513 VDD.n1469 9.3005
R1807 VDD.n1485 VDD.n1484 9.3005
R1808 VDD.n1446 VDD.n1401 9.3005
R1809 VDD.n1458 VDD.n1457 9.3005
R1810 VDD.n1416 VDD.n1415 9.3005
R1811 VDD.n1289 VDD.n1288 9.3005
R1812 VDD.n1319 VDD.n1253 9.3005
R1813 VDD.n1331 VDD.n1330 9.3005
R1814 VDD.n1358 VDD.n1357 9.3005
R1815 VDD.n1385 VDD.n1342 9.3005
R1816 VDD.n2477 VDD.n2476 9.3005
R1817 VDD.n2846 VDD.n2843 9.3005
R1818 VDD.n4281 VDD.n4280 9.3005
R1819 VDD.n4229 VDD.n4228 9.3005
R1820 VDD.n3135 VDD.n3134 9.3005
R1821 VDD.n3138 VDD.n3137 9.3005
R1822 VDD.n4110 VDD.n4109 9.3005
R1823 VDD.n3401 VDD.n3400 9.3005
R1824 VDD.n3404 VDD.n3403 9.3005
R1825 VDD.n3991 VDD.n3990 9.3005
R1826 VDD.n3667 VDD.n3666 9.3005
R1827 VDD.n3670 VDD.n3669 9.3005
R1828 VDD.n3872 VDD.n3871 9.3005
R1829 VDD.n3761 VDD.n3760 9.3005
R1830 VDD.n3893 VDD.n3892 9.3005
R1831 VDD.n3718 VDD.n3717 9.3005
R1832 VDD.n3914 VDD.n3913 9.3005
R1833 VDD.n3661 VDD.n3617 9.3005
R1834 VDD.n3633 VDD.n3632 9.3005
R1835 VDD.n3606 VDD.n3605 9.3005
R1836 VDD.n3594 VDD.n3553 9.3005
R1837 VDD.n3564 VDD.n3563 9.3005
R1838 VDD.n3495 VDD.n3494 9.3005
R1839 VDD.n4012 VDD.n4011 9.3005
R1840 VDD.n3452 VDD.n3451 9.3005
R1841 VDD.n4033 VDD.n4032 9.3005
R1842 VDD.n3395 VDD.n3351 9.3005
R1843 VDD.n3367 VDD.n3366 9.3005
R1844 VDD.n3340 VDD.n3339 9.3005
R1845 VDD.n3328 VDD.n3287 9.3005
R1846 VDD.n3298 VDD.n3297 9.3005
R1847 VDD.n3229 VDD.n3228 9.3005
R1848 VDD.n4131 VDD.n4130 9.3005
R1849 VDD.n3186 VDD.n3185 9.3005
R1850 VDD.n4152 VDD.n4151 9.3005
R1851 VDD.n3129 VDD.n3085 9.3005
R1852 VDD.n3101 VDD.n3100 9.3005
R1853 VDD.n3074 VDD.n3073 9.3005
R1854 VDD.n3062 VDD.n3021 9.3005
R1855 VDD.n3032 VDD.n3031 9.3005
R1856 VDD.n2963 VDD.n2962 9.3005
R1857 VDD.n4250 VDD.n4249 9.3005
R1858 VDD.n2920 VDD.n2919 9.3005
R1859 VDD.n4271 VDD.n4270 9.3005
R1860 VDD.n2878 VDD.n2877 9.3005
R1861 VDD.n2832 VDD.n2831 9.3005
R1862 VDD.n2790 VDD.n2789 9.3005
R1863 VDD.n2820 VDD.n2779 9.3005
R1864 VDD.n2768 VDD.n2767 9.3005
R1865 VDD.n3880 VDD.n3879 9.3005
R1866 VDD.n3879 VDD.n3878 9.3005
R1867 VDD.n3878 VDD.n3877 9.3005
R1868 VDD.n3755 VDD.n3728 9.3005
R1869 VDD.n3755 VDD.n3725 9.3005
R1870 VDD.n3725 VDD.n3724 9.3005
R1871 VDD.n3901 VDD.n3900 9.3005
R1872 VDD.n3900 VDD.n3899 9.3005
R1873 VDD.n3899 VDD.n3898 9.3005
R1874 VDD.n3712 VDD.n3685 9.3005
R1875 VDD.n3712 VDD.n3682 9.3005
R1876 VDD.n3682 VDD.n3681 9.3005
R1877 VDD.n3820 VDD.n3771 9.3005
R1878 VDD.n3820 VDD.n3768 9.3005
R1879 VDD.n3768 VDD.n3767 9.3005
R1880 VDD.n3922 VDD.n3921 9.3005
R1881 VDD.n3921 VDD.n3920 9.3005
R1882 VDD.n3920 VDD.n3919 9.3005
R1883 VDD.n3939 VDD.n3938 9.3005
R1884 VDD.n3939 VDD.n3612 9.3005
R1885 VDD.n3612 VDD.n3611 9.3005
R1886 VDD.n3947 VDD.n3946 9.3005
R1887 VDD.n3946 VDD.n3945 9.3005
R1888 VDD.n3945 VDD.n3944 9.3005
R1889 VDD.n3601 VDD.n3555 9.3005
R1890 VDD.n3601 VDD.n3593 9.3005
R1891 VDD.n3593 VDD.n3592 9.3005
R1892 VDD.n3966 VDD.n3965 9.3005
R1893 VDD.n3966 VDD.n3548 9.3005
R1894 VDD.n3548 VDD.n3547 9.3005
R1895 VDD.n3677 VDD.n3619 9.3005
R1896 VDD.n3678 VDD.n3677 9.3005
R1897 VDD.n3679 VDD.n3678 9.3005
R1898 VDD.n3974 VDD.n3973 9.3005
R1899 VDD.n3973 VDD.n3972 9.3005
R1900 VDD.n3972 VDD.n3971 9.3005
R1901 VDD.n3999 VDD.n3998 9.3005
R1902 VDD.n3998 VDD.n3997 9.3005
R1903 VDD.n3997 VDD.n3996 9.3005
R1904 VDD.n3489 VDD.n3462 9.3005
R1905 VDD.n3489 VDD.n3459 9.3005
R1906 VDD.n3459 VDD.n3458 9.3005
R1907 VDD.n4020 VDD.n4019 9.3005
R1908 VDD.n4019 VDD.n4018 9.3005
R1909 VDD.n4018 VDD.n4017 9.3005
R1910 VDD.n3446 VDD.n3419 9.3005
R1911 VDD.n3446 VDD.n3416 9.3005
R1912 VDD.n3416 VDD.n3415 9.3005
R1913 VDD.n3536 VDD.n3505 9.3005
R1914 VDD.n3536 VDD.n3502 9.3005
R1915 VDD.n3502 VDD.n3501 9.3005
R1916 VDD.n4041 VDD.n4040 9.3005
R1917 VDD.n4040 VDD.n4039 9.3005
R1918 VDD.n4039 VDD.n4038 9.3005
R1919 VDD.n4058 VDD.n4057 9.3005
R1920 VDD.n4058 VDD.n3346 9.3005
R1921 VDD.n3346 VDD.n3345 9.3005
R1922 VDD.n4066 VDD.n4065 9.3005
R1923 VDD.n4065 VDD.n4064 9.3005
R1924 VDD.n4064 VDD.n4063 9.3005
R1925 VDD.n3335 VDD.n3289 9.3005
R1926 VDD.n3335 VDD.n3327 9.3005
R1927 VDD.n3327 VDD.n3326 9.3005
R1928 VDD.n4085 VDD.n4084 9.3005
R1929 VDD.n4085 VDD.n3282 9.3005
R1930 VDD.n3282 VDD.n3281 9.3005
R1931 VDD.n3411 VDD.n3353 9.3005
R1932 VDD.n3412 VDD.n3411 9.3005
R1933 VDD.n3413 VDD.n3412 9.3005
R1934 VDD.n4093 VDD.n4092 9.3005
R1935 VDD.n4092 VDD.n4091 9.3005
R1936 VDD.n4091 VDD.n4090 9.3005
R1937 VDD.n4118 VDD.n4117 9.3005
R1938 VDD.n4117 VDD.n4116 9.3005
R1939 VDD.n4116 VDD.n4115 9.3005
R1940 VDD.n3223 VDD.n3196 9.3005
R1941 VDD.n3223 VDD.n3193 9.3005
R1942 VDD.n3193 VDD.n3192 9.3005
R1943 VDD.n4139 VDD.n4138 9.3005
R1944 VDD.n4138 VDD.n4137 9.3005
R1945 VDD.n4137 VDD.n4136 9.3005
R1946 VDD.n3180 VDD.n3153 9.3005
R1947 VDD.n3180 VDD.n3150 9.3005
R1948 VDD.n3150 VDD.n3149 9.3005
R1949 VDD.n3270 VDD.n3239 9.3005
R1950 VDD.n3270 VDD.n3236 9.3005
R1951 VDD.n3236 VDD.n3235 9.3005
R1952 VDD.n4160 VDD.n4159 9.3005
R1953 VDD.n4159 VDD.n4158 9.3005
R1954 VDD.n4158 VDD.n4157 9.3005
R1955 VDD.n4177 VDD.n4176 9.3005
R1956 VDD.n4177 VDD.n3080 9.3005
R1957 VDD.n3080 VDD.n3079 9.3005
R1958 VDD.n4185 VDD.n4184 9.3005
R1959 VDD.n4184 VDD.n4183 9.3005
R1960 VDD.n4183 VDD.n4182 9.3005
R1961 VDD.n3069 VDD.n3023 9.3005
R1962 VDD.n3069 VDD.n3061 9.3005
R1963 VDD.n3061 VDD.n3060 9.3005
R1964 VDD.n4204 VDD.n4203 9.3005
R1965 VDD.n4204 VDD.n3016 9.3005
R1966 VDD.n3016 VDD.n3015 9.3005
R1967 VDD.n3145 VDD.n3087 9.3005
R1968 VDD.n3146 VDD.n3145 9.3005
R1969 VDD.n3147 VDD.n3146 9.3005
R1970 VDD.n4212 VDD.n4211 9.3005
R1971 VDD.n4211 VDD.n4210 9.3005
R1972 VDD.n4210 VDD.n4209 9.3005
R1973 VDD.n4237 VDD.n4236 9.3005
R1974 VDD.n4236 VDD.n4235 9.3005
R1975 VDD.n4235 VDD.n4234 9.3005
R1976 VDD.n2957 VDD.n2930 9.3005
R1977 VDD.n2957 VDD.n2927 9.3005
R1978 VDD.n2927 VDD.n2926 9.3005
R1979 VDD.n4258 VDD.n4257 9.3005
R1980 VDD.n4257 VDD.n4256 9.3005
R1981 VDD.n4256 VDD.n4255 9.3005
R1982 VDD.n2914 VDD.n2855 9.3005
R1983 VDD.n2914 VDD.n2852 9.3005
R1984 VDD.n2852 VDD.n2851 9.3005
R1985 VDD.n3004 VDD.n2973 9.3005
R1986 VDD.n3004 VDD.n2970 9.3005
R1987 VDD.n2970 VDD.n2969 9.3005
R1988 VDD.n4278 VDD.n2848 9.3005
R1989 VDD.n4278 VDD.n4277 9.3005
R1990 VDD.n4277 VDD.n4276 9.3005
R1991 VDD.n4296 VDD.n4295 9.3005
R1992 VDD.n4295 VDD.n4294 9.3005
R1993 VDD.n4294 VDD.n4293 9.3005
R1994 VDD.n2827 VDD.n2781 9.3005
R1995 VDD.n2827 VDD.n2819 9.3005
R1996 VDD.n2819 VDD.n2818 9.3005
R1997 VDD.n4323 VDD.n4322 9.3005
R1998 VDD.n4322 VDD.n4321 9.3005
R1999 VDD.n4321 VDD.n4320 9.3005
R2000 VDD.n4315 VDD.n4314 9.3005
R2001 VDD.n4315 VDD.n2774 9.3005
R2002 VDD.n2774 VDD.n2773 9.3005
R2003 VDD.n4288 VDD.n4287 9.3005
R2004 VDD.n4288 VDD.n2838 9.3005
R2005 VDD.n2838 VDD.n2837 9.3005
R2006 VDD.n4333 VDD.n2739 9.3005
R2007 VDD.n2762 VDD.n2739 9.3005
R2008 VDD.n2762 VDD.n2757 9.3005
R2009 VDD.n2632 VDD.n2631 9.3005
R2010 VDD.n2631 VDD.n2450 9.3005
R2011 VDD.n2450 VDD.n2449 9.3005
R2012 VDD.n4376 VDD.n4375 9.3005
R2013 VDD.n4375 VDD.n4374 9.3005
R2014 VDD.n4374 VDD.n4373 9.3005
R2015 VDD.n4368 VDD.n4367 9.3005
R2016 VDD.n4368 VDD.n2643 9.3005
R2017 VDD.n2643 VDD.n2642 9.3005
R2018 VDD.n2701 VDD.n2650 9.3005
R2019 VDD.n2701 VDD.n2693 9.3005
R2020 VDD.n2693 VDD.n2692 9.3005
R2021 VDD.n4349 VDD.n4348 9.3005
R2022 VDD.n4348 VDD.n4347 9.3005
R2023 VDD.n4347 VDD.n4346 9.3005
R2024 VDD.n4341 VDD.n2712 9.3005
R2025 VDD.n2712 VDD.n2711 9.3005
R2026 VDD.n2483 VDD.n2482 9.3005
R2027 VDD.n2483 VDD.n2455 9.3005
R2028 VDD.n2596 VDD.n2455 9.3005
R2029 VDD.n4415 VDD.n4414 9.3005
R2030 VDD.n4414 VDD.n4413 9.3005
R2031 VDD.n4413 VDD.n4412 9.3005
R2032 VDD.n2396 VDD.n2371 9.3005
R2033 VDD.n2396 VDD.n2368 9.3005
R2034 VDD.n2368 VDD.n2367 9.3005
R2035 VDD.n4437 VDD.n4436 9.3005
R2036 VDD.n4436 VDD.n4435 9.3005
R2037 VDD.n4435 VDD.n4434 9.3005
R2038 VDD.n2354 VDD.n2329 9.3005
R2039 VDD.n2354 VDD.n2326 9.3005
R2040 VDD.n2326 VDD.n2325 9.3005
R2041 VDD.n2537 VDD.n2413 9.3005
R2042 VDD.n2537 VDD.n2410 9.3005
R2043 VDD.n2410 VDD.n2409 9.3005
R2044 VDD.n4459 VDD.n4458 9.3005
R2045 VDD.n4458 VDD.n4457 9.3005
R2046 VDD.n4457 VDD.n4456 9.3005
R2047 VDD.n4476 VDD.n4475 9.3005
R2048 VDD.n4476 VDD.n2256 9.3005
R2049 VDD.n2256 VDD.n2255 9.3005
R2050 VDD.n4484 VDD.n4483 9.3005
R2051 VDD.n4483 VDD.n4482 9.3005
R2052 VDD.n4482 VDD.n4481 9.3005
R2053 VDD.n2245 VDD.n2199 9.3005
R2054 VDD.n2245 VDD.n2237 9.3005
R2055 VDD.n2237 VDD.n2236 9.3005
R2056 VDD.n4503 VDD.n4502 9.3005
R2057 VDD.n4503 VDD.n2192 9.3005
R2058 VDD.n2192 VDD.n2191 9.3005
R2059 VDD.n2321 VDD.n2263 9.3005
R2060 VDD.n2322 VDD.n2321 9.3005
R2061 VDD.n2323 VDD.n2322 9.3005
R2062 VDD.n4511 VDD.n4510 9.3005
R2063 VDD.n4510 VDD.n4509 9.3005
R2064 VDD.n4509 VDD.n4508 9.3005
R2065 VDD.n4536 VDD.n4535 9.3005
R2066 VDD.n4535 VDD.n4534 9.3005
R2067 VDD.n4534 VDD.n4533 9.3005
R2068 VDD.n2132 VDD.n2107 9.3005
R2069 VDD.n2132 VDD.n2104 9.3005
R2070 VDD.n2104 VDD.n2103 9.3005
R2071 VDD.n4558 VDD.n4557 9.3005
R2072 VDD.n4557 VDD.n4556 9.3005
R2073 VDD.n4556 VDD.n4555 9.3005
R2074 VDD.n2090 VDD.n2065 9.3005
R2075 VDD.n2090 VDD.n2062 9.3005
R2076 VDD.n2062 VDD.n2061 9.3005
R2077 VDD.n2180 VDD.n2149 9.3005
R2078 VDD.n2180 VDD.n2146 9.3005
R2079 VDD.n2146 VDD.n2145 9.3005
R2080 VDD.n4580 VDD.n4579 9.3005
R2081 VDD.n4579 VDD.n4578 9.3005
R2082 VDD.n4578 VDD.n4577 9.3005
R2083 VDD.n4597 VDD.n4596 9.3005
R2084 VDD.n4597 VDD.n1992 9.3005
R2085 VDD.n1992 VDD.n1991 9.3005
R2086 VDD.n4605 VDD.n4604 9.3005
R2087 VDD.n4604 VDD.n4603 9.3005
R2088 VDD.n4603 VDD.n4602 9.3005
R2089 VDD.n1981 VDD.n1935 9.3005
R2090 VDD.n1981 VDD.n1973 9.3005
R2091 VDD.n1973 VDD.n1972 9.3005
R2092 VDD.n4624 VDD.n4623 9.3005
R2093 VDD.n4624 VDD.n1928 9.3005
R2094 VDD.n1928 VDD.n1927 9.3005
R2095 VDD.n2057 VDD.n1999 9.3005
R2096 VDD.n2058 VDD.n2057 9.3005
R2097 VDD.n2059 VDD.n2058 9.3005
R2098 VDD.n4632 VDD.n4631 9.3005
R2099 VDD.n4631 VDD.n4630 9.3005
R2100 VDD.n4630 VDD.n4629 9.3005
R2101 VDD.n4657 VDD.n4656 9.3005
R2102 VDD.n4656 VDD.n4655 9.3005
R2103 VDD.n4655 VDD.n4654 9.3005
R2104 VDD.n1868 VDD.n1843 9.3005
R2105 VDD.n1868 VDD.n1840 9.3005
R2106 VDD.n1840 VDD.n1839 9.3005
R2107 VDD.n4679 VDD.n4678 9.3005
R2108 VDD.n4678 VDD.n4677 9.3005
R2109 VDD.n4677 VDD.n4676 9.3005
R2110 VDD.n1826 VDD.n1801 9.3005
R2111 VDD.n1826 VDD.n1798 9.3005
R2112 VDD.n1798 VDD.n1797 9.3005
R2113 VDD.n1916 VDD.n1885 9.3005
R2114 VDD.n1916 VDD.n1882 9.3005
R2115 VDD.n1882 VDD.n1881 9.3005
R2116 VDD.n4701 VDD.n4700 9.3005
R2117 VDD.n4700 VDD.n4699 9.3005
R2118 VDD.n4699 VDD.n4698 9.3005
R2119 VDD.n4718 VDD.n4717 9.3005
R2120 VDD.n4718 VDD.n1728 9.3005
R2121 VDD.n1728 VDD.n1727 9.3005
R2122 VDD.n4726 VDD.n4725 9.3005
R2123 VDD.n4725 VDD.n4724 9.3005
R2124 VDD.n4724 VDD.n4723 9.3005
R2125 VDD.n1717 VDD.n1671 9.3005
R2126 VDD.n1717 VDD.n1709 9.3005
R2127 VDD.n1709 VDD.n1708 9.3005
R2128 VDD.n4745 VDD.n4744 9.3005
R2129 VDD.n4745 VDD.n1664 9.3005
R2130 VDD.n1664 VDD.n1663 9.3005
R2131 VDD.n1793 VDD.n1735 9.3005
R2132 VDD.n1794 VDD.n1793 9.3005
R2133 VDD.n1795 VDD.n1794 9.3005
R2134 VDD.n4753 VDD.n4752 9.3005
R2135 VDD.n4752 VDD.n4751 9.3005
R2136 VDD.n4751 VDD.n4750 9.3005
R2137 VDD.n4778 VDD.n4777 9.3005
R2138 VDD.n4777 VDD.n4776 9.3005
R2139 VDD.n4776 VDD.n4775 9.3005
R2140 VDD.n1604 VDD.n1579 9.3005
R2141 VDD.n1604 VDD.n1576 9.3005
R2142 VDD.n1576 VDD.n1575 9.3005
R2143 VDD.n4800 VDD.n4799 9.3005
R2144 VDD.n4799 VDD.n4798 9.3005
R2145 VDD.n4798 VDD.n4797 9.3005
R2146 VDD.n1562 VDD.n1537 9.3005
R2147 VDD.n1562 VDD.n1534 9.3005
R2148 VDD.n1534 VDD.n1533 9.3005
R2149 VDD.n1652 VDD.n1621 9.3005
R2150 VDD.n1652 VDD.n1618 9.3005
R2151 VDD.n1618 VDD.n1617 9.3005
R2152 VDD.n4822 VDD.n4821 9.3005
R2153 VDD.n4821 VDD.n4820 9.3005
R2154 VDD.n4820 VDD.n4819 9.3005
R2155 VDD.n4839 VDD.n4838 9.3005
R2156 VDD.n4839 VDD.n1464 9.3005
R2157 VDD.n1464 VDD.n1463 9.3005
R2158 VDD.n4847 VDD.n4846 9.3005
R2159 VDD.n4846 VDD.n4845 9.3005
R2160 VDD.n4845 VDD.n4844 9.3005
R2161 VDD.n4866 VDD.n4865 9.3005
R2162 VDD.n4866 VDD.n1396 9.3005
R2163 VDD.n1396 VDD.n1395 9.3005
R2164 VDD.n1453 VDD.n1403 9.3005
R2165 VDD.n1453 VDD.n1445 9.3005
R2166 VDD.n1445 VDD.n1444 9.3005
R2167 VDD.n1529 VDD.n1471 9.3005
R2168 VDD.n1530 VDD.n1529 9.3005
R2169 VDD.n1531 VDD.n1530 9.3005
R2170 VDD.n4874 VDD.n4873 9.3005
R2171 VDD.n4873 VDD.n4872 9.3005
R2172 VDD.n4872 VDD.n4871 9.3005
R2173 VDD.n4925 VDD.n1245 9.3005
R2174 VDD.n4925 VDD.n4924 9.3005
R2175 VDD.n4924 VDD.n4923 9.3005
R2176 VDD.n4918 VDD.n4917 9.3005
R2177 VDD.n4918 VDD.n1248 9.3005
R2178 VDD.n1248 VDD.n1247 9.3005
R2179 VDD.n1326 VDD.n1255 9.3005
R2180 VDD.n1326 VDD.n1318 9.3005
R2181 VDD.n1318 VDD.n1317 9.3005
R2182 VDD.n4899 VDD.n4898 9.3005
R2183 VDD.n4898 VDD.n4897 9.3005
R2184 VDD.n4897 VDD.n4896 9.3005
R2185 VDD.n4891 VDD.n4890 9.3005
R2186 VDD.n4891 VDD.n1337 9.3005
R2187 VDD.n1337 VDD.n1336 9.3005
R2188 VDD.n1391 VDD.n1390 9.3005
R2189 VDD.n1392 VDD.n1391 9.3005
R2190 VDD.n4965 VDD.n4964 9.3005
R2191 VDD.n4966 VDD.n4965 9.3005
R2192 VDD.n4967 VDD.n4966 9.3005
R2193 VDD.n4954 VDD.n4935 9.3005
R2194 VDD.n1147 VDD.n1146 9.3005
R2195 VDD.n1133 VDD.n1131 9.3005
R2196 VDD.n5216 VDD.n5215 9.3005
R2197 VDD.n1012 VDD.n1011 9.3005
R2198 VDD.n998 VDD.n996 9.3005
R2199 VDD.n5444 VDD.n5443 9.3005
R2200 VDD.n877 VDD.n876 9.3005
R2201 VDD.n863 VDD.n861 9.3005
R2202 VDD.n5672 VDD.n5671 9.3005
R2203 VDD.n742 VDD.n741 9.3005
R2204 VDD.n736 VDD.n735 9.3005
R2205 VDD.n680 VDD.n679 9.3005
R2206 VDD.n5889 VDD.n5888 9.3005
R2207 VDD.n697 VDD.n696 9.3005
R2208 VDD.n5856 VDD.n5855 9.3005
R2209 VDD.n5831 VDD.n5830 9.3005
R2210 VDD.n5805 VDD.n5804 9.3005
R2211 VDD.n761 VDD.n760 9.3005
R2212 VDD.n5763 VDD.n5762 9.3005
R2213 VDD.n5753 VDD.n5752 9.3005
R2214 VDD.n5723 VDD.n5722 9.3005
R2215 VDD.n5662 VDD.n5661 9.3005
R2216 VDD.n833 VDD.n832 9.3005
R2217 VDD.n5616 VDD.n5615 9.3005
R2218 VDD.n848 VDD.n847 9.3005
R2219 VDD.n5578 VDD.n5577 9.3005
R2220 VDD.n896 VDD.n895 9.3005
R2221 VDD.n5535 VDD.n5534 9.3005
R2222 VDD.n5525 VDD.n5524 9.3005
R2223 VDD.n5495 VDD.n5494 9.3005
R2224 VDD.n5434 VDD.n5433 9.3005
R2225 VDD.n968 VDD.n967 9.3005
R2226 VDD.n5388 VDD.n5387 9.3005
R2227 VDD.n983 VDD.n982 9.3005
R2228 VDD.n5350 VDD.n5349 9.3005
R2229 VDD.n1031 VDD.n1030 9.3005
R2230 VDD.n5307 VDD.n5306 9.3005
R2231 VDD.n5297 VDD.n5296 9.3005
R2232 VDD.n5267 VDD.n5266 9.3005
R2233 VDD.n5206 VDD.n5205 9.3005
R2234 VDD.n1103 VDD.n1102 9.3005
R2235 VDD.n5160 VDD.n5159 9.3005
R2236 VDD.n1118 VDD.n1117 9.3005
R2237 VDD.n5122 VDD.n5121 9.3005
R2238 VDD.n1166 VDD.n1165 9.3005
R2239 VDD.n5069 VDD.n5068 9.3005
R2240 VDD.n5079 VDD.n5078 9.3005
R2241 VDD.n5039 VDD.n5038 9.3005
R2242 VDD.n5916 VDD.n5915 9.3005
R2243 VDD.n5916 VDD.n675 9.3005
R2244 VDD.n5881 VDD.n693 9.3005
R2245 VDD.n5882 VDD.n5881 9.3005
R2246 VDD.n5853 VDD.n699 9.3005
R2247 VDD.n5853 VDD.n5852 9.3005
R2248 VDD.n5846 VDD.n5845 9.3005
R2249 VDD.n5847 VDD.n5846 9.3005
R2250 VDD.n5923 VDD.n5922 9.3005
R2251 VDD.n5824 VDD.n5823 9.3005
R2252 VDD.n5825 VDD.n5824 9.3005
R2253 VDD.n5825 VDD.n641 9.3005
R2254 VDD.n5792 VDD.n5791 9.3005
R2255 VDD.n5791 VDD.n744 9.3005
R2256 VDD.n5784 VDD.n5783 9.3005
R2257 VDD.n5785 VDD.n5784 9.3005
R2258 VDD.n5744 VDD.n770 9.3005
R2259 VDD.n5758 VDD.n770 9.3005
R2260 VDD.n5731 VDD.n5730 9.3005
R2261 VDD.n5730 VDD.n5729 9.3005
R2262 VDD.n5812 VDD.n5811 9.3005
R2263 VDD.n5811 VDD.n5810 9.3005
R2264 VDD.n5810 VDD.n641 9.3005
R2265 VDD.n5710 VDD.n5709 9.3005
R2266 VDD.n5709 VDD.n784 9.3005
R2267 VDD.n784 VDD.n641 9.3005
R2268 VDD.n811 VDD.n810 9.3005
R2269 VDD.n5666 VDD.n811 9.3005
R2270 VDD.n5647 VDD.n5646 9.3005
R2271 VDD.n5646 VDD.n5645 9.3005
R2272 VDD.n5639 VDD.n5638 9.3005
R2273 VDD.n5639 VDD.n828 9.3005
R2274 VDD.n5608 VDD.n844 9.3005
R2275 VDD.n5609 VDD.n5608 9.3005
R2276 VDD.n5699 VDD.n5698 9.3005
R2277 VDD.n5700 VDD.n5699 9.3005
R2278 VDD.n869 VDD.n850 9.3005
R2279 VDD.n869 VDD.n868 9.3005
R2280 VDD.n868 VDD.n641 9.3005
R2281 VDD.n5564 VDD.n5563 9.3005
R2282 VDD.n5563 VDD.n879 9.3005
R2283 VDD.n5556 VDD.n5555 9.3005
R2284 VDD.n5557 VDD.n5556 9.3005
R2285 VDD.n5516 VDD.n905 9.3005
R2286 VDD.n5530 VDD.n905 9.3005
R2287 VDD.n5503 VDD.n5502 9.3005
R2288 VDD.n5502 VDD.n5501 9.3005
R2289 VDD.n5585 VDD.n5584 9.3005
R2290 VDD.n5584 VDD.n5583 9.3005
R2291 VDD.n5583 VDD.n641 9.3005
R2292 VDD.n5482 VDD.n5481 9.3005
R2293 VDD.n5481 VDD.n919 9.3005
R2294 VDD.n919 VDD.n641 9.3005
R2295 VDD.n946 VDD.n945 9.3005
R2296 VDD.n5438 VDD.n946 9.3005
R2297 VDD.n5419 VDD.n5418 9.3005
R2298 VDD.n5418 VDD.n5417 9.3005
R2299 VDD.n5411 VDD.n5410 9.3005
R2300 VDD.n5411 VDD.n963 9.3005
R2301 VDD.n5380 VDD.n979 9.3005
R2302 VDD.n5381 VDD.n5380 9.3005
R2303 VDD.n5471 VDD.n5470 9.3005
R2304 VDD.n5472 VDD.n5471 9.3005
R2305 VDD.n1004 VDD.n985 9.3005
R2306 VDD.n1004 VDD.n1003 9.3005
R2307 VDD.n1003 VDD.n641 9.3005
R2308 VDD.n5336 VDD.n5335 9.3005
R2309 VDD.n5335 VDD.n1014 9.3005
R2310 VDD.n5328 VDD.n5327 9.3005
R2311 VDD.n5329 VDD.n5328 9.3005
R2312 VDD.n5288 VDD.n1040 9.3005
R2313 VDD.n5302 VDD.n1040 9.3005
R2314 VDD.n5275 VDD.n5274 9.3005
R2315 VDD.n5274 VDD.n5273 9.3005
R2316 VDD.n5357 VDD.n5356 9.3005
R2317 VDD.n5356 VDD.n5355 9.3005
R2318 VDD.n5355 VDD.n641 9.3005
R2319 VDD.n5254 VDD.n5253 9.3005
R2320 VDD.n5253 VDD.n1054 9.3005
R2321 VDD.n1054 VDD.n641 9.3005
R2322 VDD.n1081 VDD.n1080 9.3005
R2323 VDD.n5210 VDD.n1081 9.3005
R2324 VDD.n5191 VDD.n5190 9.3005
R2325 VDD.n5190 VDD.n5189 9.3005
R2326 VDD.n5183 VDD.n5182 9.3005
R2327 VDD.n5183 VDD.n1098 9.3005
R2328 VDD.n5152 VDD.n1114 9.3005
R2329 VDD.n5153 VDD.n5152 9.3005
R2330 VDD.n5243 VDD.n5242 9.3005
R2331 VDD.n5244 VDD.n5243 9.3005
R2332 VDD.n1139 VDD.n1120 9.3005
R2333 VDD.n1139 VDD.n1138 9.3005
R2334 VDD.n1138 VDD.n641 9.3005
R2335 VDD.n5108 VDD.n5107 9.3005
R2336 VDD.n5107 VDD.n1149 9.3005
R2337 VDD.n5100 VDD.n5099 9.3005
R2338 VDD.n5101 VDD.n5100 9.3005
R2339 VDD.n5047 VDD.n5046 9.3005
R2340 VDD.n5046 VDD.n5045 9.3005
R2341 VDD.n5060 VDD.n1175 9.3005
R2342 VDD.n5074 VDD.n1175 9.3005
R2343 VDD.n5129 VDD.n5128 9.3005
R2344 VDD.n5128 VDD.n5127 9.3005
R2345 VDD.n5127 VDD.n641 9.3005
R2346 VDD.n5026 VDD.n5025 9.3005
R2347 VDD.n6012 VDD.n5972 9.3005
R2348 VDD.n6012 VDD.n6011 9.3005
R2349 VDD.n6046 VDD.n5957 9.3005
R2350 VDD.n6046 VDD.n6045 9.3005
R2351 VDD.n6066 VDD.n6065 9.3005
R2352 VDD.n6067 VDD.n6066 9.3005
R2353 VDD.n5965 VDD.n5954 9.3005
R2354 VDD.n5965 VDD.n5964 9.3005
R2355 VDD.n6027 VDD.n6026 9.3005
R2356 VDD.n6026 VDD.n6025 9.3005
R2357 VDD.n6072 VDD.n6071 9.3005
R2358 VDD.n6073 VDD.n6072 9.3005
R2359 VDD.n6121 VDD.n6120 9.3005
R2360 VDD.n6121 VDD.n606 9.3005
R2361 VDD.n606 VDD.n605 9.3005
R2362 VDD.n7216 VDD.n7215 9.3005
R2363 VDD.n7217 VDD.n7216 9.3005
R2364 VDD.n7115 VDD.n7104 9.3005
R2365 VDD.n7115 VDD.n7114 9.3005
R2366 VDD.n7196 VDD.n7107 9.3005
R2367 VDD.n7196 VDD.n7195 9.3005
R2368 VDD.n7162 VDD.n7122 9.3005
R2369 VDD.n7162 VDD.n7161 9.3005
R2370 VDD.n7177 VDD.n7176 9.3005
R2371 VDD.n7176 VDD.n7175 9.3005
R2372 VDD.n7222 VDD.n7221 9.3005
R2373 VDD.n7223 VDD.n7222 9.3005
R2374 VDD.n6396 VDD.n6395 9.3005
R2375 VDD.n6395 VDD.n6394 9.3005
R2376 VDD.n6364 VDD.n6363 9.3005
R2377 VDD.n6364 VDD.n460 9.3005
R2378 VDD.n6305 VDD.n482 9.3005
R2379 VDD.n6305 VDD.n6304 9.3005
R2380 VDD.n6297 VDD.n6296 9.3005
R2381 VDD.n6333 VDD.n476 9.3005
R2382 VDD.n6334 VDD.n6333 9.3005
R2383 VDD.n6372 VDD.n6371 9.3005
R2384 VDD.n6371 VDD.n6370 9.3005
R2385 VDD.n6622 VDD.n6621 9.3005
R2386 VDD.n6621 VDD.n6620 9.3005
R2387 VDD.n6590 VDD.n6589 9.3005
R2388 VDD.n6590 VDD.n326 9.3005
R2389 VDD.n6531 VDD.n348 9.3005
R2390 VDD.n6531 VDD.n6530 9.3005
R2391 VDD.n6523 VDD.n6522 9.3005
R2392 VDD.n6559 VDD.n342 9.3005
R2393 VDD.n6560 VDD.n6559 9.3005
R2394 VDD.n6598 VDD.n6597 9.3005
R2395 VDD.n6597 VDD.n6596 9.3005
R2396 VDD.n6848 VDD.n6847 9.3005
R2397 VDD.n6847 VDD.n6846 9.3005
R2398 VDD.n6816 VDD.n6815 9.3005
R2399 VDD.n6816 VDD.n192 9.3005
R2400 VDD.n6757 VDD.n214 9.3005
R2401 VDD.n6757 VDD.n6756 9.3005
R2402 VDD.n6749 VDD.n6748 9.3005
R2403 VDD.n6785 VDD.n208 9.3005
R2404 VDD.n6786 VDD.n6785 9.3005
R2405 VDD.n6824 VDD.n6823 9.3005
R2406 VDD.n6823 VDD.n6822 9.3005
R2407 VDD.n7042 VDD.n7041 9.3005
R2408 VDD.n7042 VDD.n58 9.3005
R2409 VDD.n6983 VDD.n80 9.3005
R2410 VDD.n6983 VDD.n6982 9.3005
R2411 VDD.n6975 VDD.n6974 9.3005
R2412 VDD.n7011 VDD.n74 9.3005
R2413 VDD.n7012 VDD.n7011 9.3005
R2414 VDD.n7050 VDD.n7049 9.3005
R2415 VDD.n7049 VDD.n7048 9.3005
R2416 VDD.n7073 VDD.n7072 9.3005
R2417 VDD.n6944 VDD.n6943 9.3005
R2418 VDD.n6943 VDD.n6942 9.3005
R2419 VDD.n6924 VDD.n6923 9.3005
R2420 VDD.n6923 VDD.n126 9.3005
R2421 VDD.n126 VDD.n12 9.3005
R2422 VDD.n6917 VDD.n6916 9.3005
R2423 VDD.n6918 VDD.n6917 9.3005
R2424 VDD.n6918 VDD.n12 9.3005
R2425 VDD.n6890 VDD.n6889 9.3005
R2426 VDD.n6891 VDD.n6890 9.3005
R2427 VDD.n6891 VDD.n12 9.3005
R2428 VDD.n6963 VDD.n6962 9.3005
R2429 VDD.n6869 VDD.n6868 9.3005
R2430 VDD.n6870 VDD.n6869 9.3005
R2431 VDD.n6870 VDD.n12 9.3005
R2432 VDD.n6718 VDD.n6717 9.3005
R2433 VDD.n6717 VDD.n6716 9.3005
R2434 VDD.n6698 VDD.n6697 9.3005
R2435 VDD.n6697 VDD.n260 9.3005
R2436 VDD.n260 VDD.n12 9.3005
R2437 VDD.n6691 VDD.n6690 9.3005
R2438 VDD.n6692 VDD.n6691 9.3005
R2439 VDD.n6692 VDD.n12 9.3005
R2440 VDD.n6664 VDD.n6663 9.3005
R2441 VDD.n6665 VDD.n6664 9.3005
R2442 VDD.n6665 VDD.n12 9.3005
R2443 VDD.n6737 VDD.n6736 9.3005
R2444 VDD.n6643 VDD.n6642 9.3005
R2445 VDD.n6644 VDD.n6643 9.3005
R2446 VDD.n6644 VDD.n12 9.3005
R2447 VDD.n6492 VDD.n6491 9.3005
R2448 VDD.n6491 VDD.n6490 9.3005
R2449 VDD.n6472 VDD.n6471 9.3005
R2450 VDD.n6471 VDD.n394 9.3005
R2451 VDD.n394 VDD.n12 9.3005
R2452 VDD.n6465 VDD.n6464 9.3005
R2453 VDD.n6466 VDD.n6465 9.3005
R2454 VDD.n6466 VDD.n12 9.3005
R2455 VDD.n6438 VDD.n6437 9.3005
R2456 VDD.n6439 VDD.n6438 9.3005
R2457 VDD.n6439 VDD.n12 9.3005
R2458 VDD.n6511 VDD.n6510 9.3005
R2459 VDD.n6417 VDD.n6416 9.3005
R2460 VDD.n6418 VDD.n6417 9.3005
R2461 VDD.n6418 VDD.n12 9.3005
R2462 VDD.n6266 VDD.n6265 9.3005
R2463 VDD.n6265 VDD.n6264 9.3005
R2464 VDD.n6246 VDD.n6245 9.3005
R2465 VDD.n6245 VDD.n528 9.3005
R2466 VDD.n528 VDD.n12 9.3005
R2467 VDD.n6239 VDD.n6238 9.3005
R2468 VDD.n6240 VDD.n6239 9.3005
R2469 VDD.n6240 VDD.n12 9.3005
R2470 VDD.n6285 VDD.n6284 9.3005
R2471 VDD.n6191 VDD.n6190 9.3005
R2472 VDD.n6212 VDD.n6211 9.3005
R2473 VDD.n6213 VDD.n6212 9.3005
R2474 VDD.n7275 VDD.n7274 9.3005
R2475 VDD.n7274 VDD.n7273 9.3005
R2476 VDD.n6069 VDD.n653 8.92171
R2477 VDD.n5959 VDD.n5958 8.92171
R2478 VDD.n5969 VDD.n5968 8.92171
R2479 VDD.n6042 VDD.n6041 8.92171
R2480 VDD.n6023 VDD.n6016 8.92171
R2481 VDD.n6196 VDD.n6195 8.92171
R2482 VDD.n6217 VDD.n6216 8.92171
R2483 VDD.n544 VDD.n538 8.92171
R2484 VDD.n6260 VDD.n6259 8.92171
R2485 VDD.n6280 VDD.n6279 8.92171
R2486 VDD.n6307 VDD.n492 8.92171
R2487 VDD.n493 VDD.n479 8.92171
R2488 VDD.n6340 VDD.n6339 8.92171
R2489 VDD.n464 VDD.n459 8.92171
R2490 VDD.n6386 VDD.n6385 8.92171
R2491 VDD.n6422 VDD.n6421 8.92171
R2492 VDD.n6443 VDD.n6442 8.92171
R2493 VDD.n410 VDD.n404 8.92171
R2494 VDD.n6486 VDD.n6485 8.92171
R2495 VDD.n6506 VDD.n6505 8.92171
R2496 VDD.n6533 VDD.n358 8.92171
R2497 VDD.n359 VDD.n345 8.92171
R2498 VDD.n6566 VDD.n6565 8.92171
R2499 VDD.n330 VDD.n325 8.92171
R2500 VDD.n6612 VDD.n6611 8.92171
R2501 VDD.n6648 VDD.n6647 8.92171
R2502 VDD.n6669 VDD.n6668 8.92171
R2503 VDD.n276 VDD.n270 8.92171
R2504 VDD.n6712 VDD.n6711 8.92171
R2505 VDD.n6732 VDD.n6731 8.92171
R2506 VDD.n6759 VDD.n224 8.92171
R2507 VDD.n225 VDD.n211 8.92171
R2508 VDD.n6792 VDD.n6791 8.92171
R2509 VDD.n196 VDD.n191 8.92171
R2510 VDD.n6838 VDD.n6837 8.92171
R2511 VDD.n6874 VDD.n6873 8.92171
R2512 VDD.n6895 VDD.n6894 8.92171
R2513 VDD.n142 VDD.n136 8.92171
R2514 VDD.n6938 VDD.n6937 8.92171
R2515 VDD.n6958 VDD.n6957 8.92171
R2516 VDD.n6985 VDD.n90 8.92171
R2517 VDD.n91 VDD.n77 8.92171
R2518 VDD.n7018 VDD.n7017 8.92171
R2519 VDD.n62 VDD.n57 8.92171
R2520 VDD.n7069 VDD.n7068 8.92171
R2521 VDD.n7219 VDD.n24 8.92171
R2522 VDD.n7109 VDD.n7108 8.92171
R2523 VDD.n7119 VDD.n7118 8.92171
R2524 VDD.n7192 VDD.n7191 8.92171
R2525 VDD.n7173 VDD.n7166 8.92171
R2526 VDD.n2638 VDD.n2637 8.92171
R2527 VDD.n2663 VDD.n2644 8.92171
R2528 VDD.n2695 VDD.n2694 8.92171
R2529 VDD.n2707 VDD.n2706 8.92171
R2530 VDD.n2726 VDD.n2713 8.92171
R2531 VDD.n1415 VDD.n1397 8.92171
R2532 VDD.n1447 VDD.n1446 8.92171
R2533 VDD.n1459 VDD.n1458 8.92171
R2534 VDD.n1484 VDD.n1465 8.92171
R2535 VDD.n1516 VDD.n1513 8.92171
R2536 VDD.n4815 VDD.n4814 8.92171
R2537 VDD.n1570 VDD.n1569 8.92171
R2538 VDD.n4793 VDD.n4792 8.92171
R2539 VDD.n1612 VDD.n1611 8.92171
R2540 VDD.n4771 VDD.n4770 8.92171
R2541 VDD.n1679 VDD.n1665 8.92171
R2542 VDD.n1711 VDD.n1710 8.92171
R2543 VDD.n1723 VDD.n1722 8.92171
R2544 VDD.n1748 VDD.n1729 8.92171
R2545 VDD.n1780 VDD.n1777 8.92171
R2546 VDD.n4694 VDD.n4693 8.92171
R2547 VDD.n1834 VDD.n1833 8.92171
R2548 VDD.n4672 VDD.n4671 8.92171
R2549 VDD.n1876 VDD.n1875 8.92171
R2550 VDD.n4650 VDD.n4649 8.92171
R2551 VDD.n1943 VDD.n1929 8.92171
R2552 VDD.n1975 VDD.n1974 8.92171
R2553 VDD.n1987 VDD.n1986 8.92171
R2554 VDD.n2012 VDD.n1993 8.92171
R2555 VDD.n2044 VDD.n2041 8.92171
R2556 VDD.n4573 VDD.n4572 8.92171
R2557 VDD.n2098 VDD.n2097 8.92171
R2558 VDD.n4551 VDD.n4550 8.92171
R2559 VDD.n2140 VDD.n2139 8.92171
R2560 VDD.n4529 VDD.n4528 8.92171
R2561 VDD.n2207 VDD.n2193 8.92171
R2562 VDD.n2239 VDD.n2238 8.92171
R2563 VDD.n2251 VDD.n2250 8.92171
R2564 VDD.n2276 VDD.n2257 8.92171
R2565 VDD.n2308 VDD.n2305 8.92171
R2566 VDD.n4452 VDD.n4451 8.92171
R2567 VDD.n2362 VDD.n2361 8.92171
R2568 VDD.n4430 VDD.n4429 8.92171
R2569 VDD.n2404 VDD.n2403 8.92171
R2570 VDD.n4408 VDD.n4407 8.92171
R2571 VDD.n1288 VDD.n1249 8.92171
R2572 VDD.n1320 VDD.n1319 8.92171
R2573 VDD.n1332 VDD.n1331 8.92171
R2574 VDD.n1357 VDD.n1338 8.92171
R2575 VDD.n1388 VDD.n1385 8.92171
R2576 VDD.n2769 VDD.n2768 8.92171
R2577 VDD.n2789 VDD.n2775 8.92171
R2578 VDD.n2821 VDD.n2820 8.92171
R2579 VDD.n2833 VDD.n2832 8.92171
R2580 VDD.n2877 VDD.n2839 8.92171
R2581 VDD.n4272 VDD.n4271 8.92171
R2582 VDD.n2921 VDD.n2920 8.92171
R2583 VDD.n4251 VDD.n4250 8.92171
R2584 VDD.n2964 VDD.n2963 8.92171
R2585 VDD.n4230 VDD.n4229 8.92171
R2586 VDD.n3031 VDD.n3017 8.92171
R2587 VDD.n3063 VDD.n3062 8.92171
R2588 VDD.n3075 VDD.n3074 8.92171
R2589 VDD.n3100 VDD.n3081 8.92171
R2590 VDD.n3132 VDD.n3129 8.92171
R2591 VDD.n4153 VDD.n4152 8.92171
R2592 VDD.n3187 VDD.n3186 8.92171
R2593 VDD.n4132 VDD.n4131 8.92171
R2594 VDD.n3230 VDD.n3229 8.92171
R2595 VDD.n4111 VDD.n4110 8.92171
R2596 VDD.n3297 VDD.n3283 8.92171
R2597 VDD.n3329 VDD.n3328 8.92171
R2598 VDD.n3341 VDD.n3340 8.92171
R2599 VDD.n3366 VDD.n3347 8.92171
R2600 VDD.n3398 VDD.n3395 8.92171
R2601 VDD.n4034 VDD.n4033 8.92171
R2602 VDD.n3453 VDD.n3452 8.92171
R2603 VDD.n4013 VDD.n4012 8.92171
R2604 VDD.n3496 VDD.n3495 8.92171
R2605 VDD.n3992 VDD.n3991 8.92171
R2606 VDD.n3563 VDD.n3549 8.92171
R2607 VDD.n3595 VDD.n3594 8.92171
R2608 VDD.n3607 VDD.n3606 8.92171
R2609 VDD.n3632 VDD.n3613 8.92171
R2610 VDD.n3664 VDD.n3661 8.92171
R2611 VDD.n3915 VDD.n3914 8.92171
R2612 VDD.n3719 VDD.n3718 8.92171
R2613 VDD.n3894 VDD.n3893 8.92171
R2614 VDD.n3762 VDD.n3761 8.92171
R2615 VDD.n3873 VDD.n3872 8.92171
R2616 VDD.n5040 VDD.n5039 8.92171
R2617 VDD.n5070 VDD.n5069 8.92171
R2618 VDD.n5078 VDD.n5077 8.92171
R2619 VDD.n1165 VDD.n1159 8.92171
R2620 VDD.n5123 VDD.n5122 8.92171
R2621 VDD.n1134 VDD.n1117 8.92171
R2622 VDD.n5159 VDD.n5158 8.92171
R2623 VDD.n1102 VDD.n1097 8.92171
R2624 VDD.n5207 VDD.n5206 8.92171
R2625 VDD.n5215 VDD.n5214 8.92171
R2626 VDD.n5268 VDD.n5267 8.92171
R2627 VDD.n5298 VDD.n5297 8.92171
R2628 VDD.n5306 VDD.n5305 8.92171
R2629 VDD.n1030 VDD.n1024 8.92171
R2630 VDD.n5351 VDD.n5350 8.92171
R2631 VDD.n999 VDD.n982 8.92171
R2632 VDD.n5387 VDD.n5386 8.92171
R2633 VDD.n967 VDD.n962 8.92171
R2634 VDD.n5435 VDD.n5434 8.92171
R2635 VDD.n5443 VDD.n5442 8.92171
R2636 VDD.n5496 VDD.n5495 8.92171
R2637 VDD.n5526 VDD.n5525 8.92171
R2638 VDD.n5534 VDD.n5533 8.92171
R2639 VDD.n895 VDD.n889 8.92171
R2640 VDD.n5579 VDD.n5578 8.92171
R2641 VDD.n864 VDD.n847 8.92171
R2642 VDD.n5615 VDD.n5614 8.92171
R2643 VDD.n832 VDD.n827 8.92171
R2644 VDD.n5663 VDD.n5662 8.92171
R2645 VDD.n5671 VDD.n5670 8.92171
R2646 VDD.n5724 VDD.n5723 8.92171
R2647 VDD.n5754 VDD.n5753 8.92171
R2648 VDD.n5762 VDD.n5761 8.92171
R2649 VDD.n760 VDD.n754 8.92171
R2650 VDD.n5806 VDD.n5805 8.92171
R2651 VDD.n5830 VDD.n5829 8.92171
R2652 VDD.n5855 VDD.n709 8.92171
R2653 VDD.n710 VDD.n696 8.92171
R2654 VDD.n5888 VDD.n5887 8.92171
R2655 VDD.n679 VDD.n674 8.92171
R2656 VDD.n5073 VDD.n641 8.77616
R2657 VDD.n5104 VDD.n641 8.77616
R2658 VDD.n5301 VDD.n641 8.77616
R2659 VDD.n5332 VDD.n641 8.77616
R2660 VDD.n5529 VDD.n641 8.77616
R2661 VDD.n5560 VDD.n641 8.77616
R2662 VDD.n5757 VDD.n641 8.77616
R2663 VDD.n5788 VDD.n641 8.77616
R2664 VDD.n5883 VDD.n641 8.77616
R2665 VDD.n5848 VDD.n641 8.77616
R2666 VDD.n5644 VDD.n641 8.77616
R2667 VDD.n5610 VDD.n641 8.77616
R2668 VDD.n5701 VDD.n641 8.77616
R2669 VDD.n5416 VDD.n641 8.77616
R2670 VDD.n5382 VDD.n641 8.77616
R2671 VDD.n5473 VDD.n641 8.77616
R2672 VDD.n5188 VDD.n641 8.77616
R2673 VDD.n5154 VDD.n641 8.77616
R2674 VDD.n5245 VDD.n641 8.77616
R2675 VDD.n6073 VDD.n649 8.77616
R2676 VDD.n6073 VDD.n643 8.77616
R2677 VDD.n6073 VDD.n647 8.77616
R2678 VDD.n6073 VDD.n645 8.77616
R2679 VDD.n7223 VDD.n20 8.77616
R2680 VDD.n7223 VDD.n14 8.77616
R2681 VDD.n7223 VDD.n18 8.77616
R2682 VDD.n7223 VDD.n16 8.77616
R2683 VDD.n6298 VDD.n12 8.77616
R2684 VDD.n6335 VDD.n12 8.77616
R2685 VDD.n6369 VDD.n12 8.77616
R2686 VDD.n6524 VDD.n12 8.77616
R2687 VDD.n6561 VDD.n12 8.77616
R2688 VDD.n6595 VDD.n12 8.77616
R2689 VDD.n6750 VDD.n12 8.77616
R2690 VDD.n6787 VDD.n12 8.77616
R2691 VDD.n6821 VDD.n12 8.77616
R2692 VDD.n6976 VDD.n12 8.77616
R2693 VDD.n7013 VDD.n12 8.77616
R2694 VDD.n7047 VDD.n12 8.77616
R2695 VDD.n6961 VDD.n12 8.77616
R2696 VDD.n6735 VDD.n12 8.77616
R2697 VDD.n6509 VDD.n12 8.77616
R2698 VDD.n6283 VDD.n12 8.77616
R2699 VDD.n554 VDD.n12 8.77616
R2700 VDD.n4999 VDD.t14 8.57285
R2701 VDD.n5025 VDD.n1189 8.45943
R2702 VDD.n5922 VDD.n5921 8.4584
R2703 VDD.n5921 VDD.n641 8.45416
R2704 VDD.n1189 VDD.n641 8.45226
R2705 VDD.t9 VDD.n4990 8.41977
R2706 VDD.t57 VDD.n6147 8.41977
R2707 VDD.n4990 VDD.n4989 7.96054
R2708 VDD.n6147 VDD.n6146 7.96054
R2709 VDD.n2595 VDD.n2594 7.84364
R2710 VDD.n5885 VDD.n641 5.63319
R2711 VDD.n5851 VDD.n641 5.63319
R2712 VDD.n5786 VDD.n641 5.63319
R2713 VDD.n5728 VDD.n641 5.63319
R2714 VDD.n5665 VDD.n641 5.63319
R2715 VDD.n5612 VDD.n641 5.63319
R2716 VDD.n5558 VDD.n641 5.63319
R2717 VDD.n5500 VDD.n641 5.63319
R2718 VDD.n5437 VDD.n641 5.63319
R2719 VDD.n5384 VDD.n641 5.63319
R2720 VDD.n5330 VDD.n641 5.63319
R2721 VDD.n5272 VDD.n641 5.63319
R2722 VDD.n5209 VDD.n641 5.63319
R2723 VDD.n5156 VDD.n641 5.63319
R2724 VDD.n5102 VDD.n641 5.63319
R2725 VDD.n5044 VDD.n641 5.63319
R2726 VDD.n6073 VDD.n646 5.63319
R2727 VDD.n7223 VDD.n17 5.63319
R2728 VDD.n517 VDD.n12 5.63319
R2729 VDD.n6388 VDD.n12 5.63319
R2730 VDD.n6337 VDD.n12 5.63319
R2731 VDD.n6301 VDD.n12 5.63319
R2732 VDD.n383 VDD.n12 5.63319
R2733 VDD.n6614 VDD.n12 5.63319
R2734 VDD.n6563 VDD.n12 5.63319
R2735 VDD.n6527 VDD.n12 5.63319
R2736 VDD.n249 VDD.n12 5.63319
R2737 VDD.n6840 VDD.n12 5.63319
R2738 VDD.n6789 VDD.n12 5.63319
R2739 VDD.n6753 VDD.n12 5.63319
R2740 VDD.n115 VDD.n12 5.63319
R2741 VDD.n7015 VDD.n12 5.63319
R2742 VDD.n6979 VDD.n12 5.63319
R2743 VDD.n6192 VDD.n12 5.1329
R2744 VDD.n7071 VDD.n12 5.1329
R2745 VDD.n4980 VDD 5.06361
R2746 VDD.n6159 VDD.t77 5.05206
R2747 VDD.n2597 VDD.n2596 4.90246
R2748 VDD.n4989 VDD.t16 4.74591
R2749 VDD.n6146 VDD.t71 4.74591
R2750 VDD.n603 VDD.n602 4.6505
R2751 VDD.n6093 VDD.n6092 4.6505
R2752 VDD.n2602 VDD.n2601 4.6505
R2753 VDD.n2457 VDD.n2456 4.6505
R2754 VDD.n4973 VDD.n4972 4.6505
R2755 VDD.n4959 VDD.n4958 4.6505
R2756 VDD.n7250 VDD.n7249 4.6505
R2757 VDD.n7281 VDD.n7280 4.6505
R2758 VDD.n5026 VDD.n5024 4.54027
R2759 VDD.n5924 VDD.n5923 4.54027
R2760 VDD.n6190 VDD.n565 4.54027
R2761 VDD.n7074 VDD.n7073 4.54027
R2762 VDD.n4334 VDD.n4333 4.54027
R2763 VDD.n3861 VDD.n3771 4.54027
R2764 VDD.n4875 VDD.n4874 4.54027
R2765 VDD.n4396 VDD.n2413 4.54027
R2766 VDD.n596 VDD.n595 4.52882
R2767 VDD.n3840 VDD.n3839 4.52882
R2768 VDD.n2516 VDD.n2515 4.52882
R2769 VDD.n1226 VDD.n1225 4.52882
R2770 VDD.n5936 VDD.n5935 4.5005
R2771 VDD.n5934 VDD.n657 4.5005
R2772 VDD.n657 VDD.n654 4.5005
R2773 VDD.n6064 VDD.n6063 4.5005
R2774 VDD.n5938 VDD.n5937 4.5005
R2775 VDD.n5998 VDD.n637 4.5005
R2776 VDD.n6018 VDD.n6017 4.5005
R2777 VDD.n5973 VDD.n5971 4.5005
R2778 VDD.n6039 VDD.n6038 4.5005
R2779 VDD.n6039 VDD.n5970 4.5005
R2780 VDD.n5988 VDD.n5987 4.5005
R2781 VDD.n6051 VDD.n6050 4.5005
R2782 VDD.n6049 VDD.n6048 4.5005
R2783 VDD.n6048 VDD.n6047 4.5005
R2784 VDD.n6053 VDD.n6052 4.5005
R2785 VDD.n661 VDD.n659 4.5005
R2786 VDD.n5962 VDD.n5961 4.5005
R2787 VDD.n5963 VDD.n5962 4.5005
R2788 VDD.n6021 VDD.n6020 4.5005
R2789 VDD.n6010 VDD.n5997 4.5005
R2790 VDD.n6024 VDD.n6010 4.5005
R2791 VDD.n6091 VDD.n6090 4.5005
R2792 VDD.n610 VDD.n608 4.5005
R2793 VDD.n611 VDD.n609 4.5005
R2794 VDD.n563 VDD.n562 4.5005
R2795 VDD.n564 VDD.n563 4.5005
R2796 VDD.n6199 VDD.n6198 4.5005
R2797 VDD.n6220 VDD.n6219 4.5005
R2798 VDD.n513 VDD.n512 4.5005
R2799 VDD.n521 VDD.n505 4.5005
R2800 VDD.n6406 VDD.n433 4.5005
R2801 VDD.n445 VDD.n438 4.5005
R2802 VDD.n6383 VDD.n6382 4.5005
R2803 VDD.n444 VDD.n442 4.5005
R2804 VDD.n446 VDD.n444 4.5005
R2805 VDD.n6362 VDD.n6361 4.5005
R2806 VDD.n6344 VDD.n6343 4.5005
R2807 VDD.n6342 VDD.n462 4.5005
R2808 VDD.n462 VDD.n461 4.5005
R2809 VDD.n6327 VDD.n6326 4.5005
R2810 VDD.n6310 VDD.n6309 4.5005
R2811 VDD.n491 VDD.n489 4.5005
R2812 VDD.n6306 VDD.n491 4.5005
R2813 VDD.n490 VDD.n488 4.5005
R2814 VDD.n511 VDD.n510 4.5005
R2815 VDD.n498 VDD.n497 4.5005
R2816 VDD.n497 VDD.n496 4.5005
R2817 VDD.n6346 VDD.n6345 4.5005
R2818 VDD.n6329 VDD.n6328 4.5005
R2819 VDD.n6331 VDD.n6330 4.5005
R2820 VDD.n6332 VDD.n6331 4.5005
R2821 VDD.n451 VDD.n450 4.5005
R2822 VDD.n468 VDD.n466 4.5005
R2823 VDD.n457 VDD.n455 4.5005
R2824 VDD.n458 VDD.n457 4.5005
R2825 VDD.n379 VDD.n378 4.5005
R2826 VDD.n387 VDD.n371 4.5005
R2827 VDD.n6632 VDD.n299 4.5005
R2828 VDD.n311 VDD.n304 4.5005
R2829 VDD.n6609 VDD.n6608 4.5005
R2830 VDD.n310 VDD.n308 4.5005
R2831 VDD.n312 VDD.n310 4.5005
R2832 VDD.n6588 VDD.n6587 4.5005
R2833 VDD.n6570 VDD.n6569 4.5005
R2834 VDD.n6568 VDD.n328 4.5005
R2835 VDD.n328 VDD.n327 4.5005
R2836 VDD.n6553 VDD.n6552 4.5005
R2837 VDD.n6536 VDD.n6535 4.5005
R2838 VDD.n357 VDD.n355 4.5005
R2839 VDD.n6532 VDD.n357 4.5005
R2840 VDD.n356 VDD.n354 4.5005
R2841 VDD.n377 VDD.n376 4.5005
R2842 VDD.n364 VDD.n363 4.5005
R2843 VDD.n363 VDD.n362 4.5005
R2844 VDD.n6572 VDD.n6571 4.5005
R2845 VDD.n6555 VDD.n6554 4.5005
R2846 VDD.n6557 VDD.n6556 4.5005
R2847 VDD.n6558 VDD.n6557 4.5005
R2848 VDD.n317 VDD.n316 4.5005
R2849 VDD.n334 VDD.n332 4.5005
R2850 VDD.n323 VDD.n321 4.5005
R2851 VDD.n324 VDD.n323 4.5005
R2852 VDD.n245 VDD.n244 4.5005
R2853 VDD.n253 VDD.n237 4.5005
R2854 VDD.n6858 VDD.n165 4.5005
R2855 VDD.n177 VDD.n170 4.5005
R2856 VDD.n6835 VDD.n6834 4.5005
R2857 VDD.n176 VDD.n174 4.5005
R2858 VDD.n178 VDD.n176 4.5005
R2859 VDD.n6814 VDD.n6813 4.5005
R2860 VDD.n6796 VDD.n6795 4.5005
R2861 VDD.n6794 VDD.n194 4.5005
R2862 VDD.n194 VDD.n193 4.5005
R2863 VDD.n6779 VDD.n6778 4.5005
R2864 VDD.n6762 VDD.n6761 4.5005
R2865 VDD.n223 VDD.n221 4.5005
R2866 VDD.n6758 VDD.n223 4.5005
R2867 VDD.n222 VDD.n220 4.5005
R2868 VDD.n243 VDD.n242 4.5005
R2869 VDD.n230 VDD.n229 4.5005
R2870 VDD.n229 VDD.n228 4.5005
R2871 VDD.n6798 VDD.n6797 4.5005
R2872 VDD.n6781 VDD.n6780 4.5005
R2873 VDD.n6783 VDD.n6782 4.5005
R2874 VDD.n6784 VDD.n6783 4.5005
R2875 VDD.n183 VDD.n182 4.5005
R2876 VDD.n200 VDD.n198 4.5005
R2877 VDD.n189 VDD.n187 4.5005
R2878 VDD.n190 VDD.n189 4.5005
R2879 VDD.n111 VDD.n110 4.5005
R2880 VDD.n119 VDD.n103 4.5005
R2881 VDD.n7066 VDD.n7065 4.5005
R2882 VDD.n7040 VDD.n7039 4.5005
R2883 VDD.n7022 VDD.n7021 4.5005
R2884 VDD.n7020 VDD.n60 4.5005
R2885 VDD.n60 VDD.n59 4.5005
R2886 VDD.n7005 VDD.n7004 4.5005
R2887 VDD.n6988 VDD.n6987 4.5005
R2888 VDD.n89 VDD.n87 4.5005
R2889 VDD.n6984 VDD.n89 4.5005
R2890 VDD.n88 VDD.n86 4.5005
R2891 VDD.n109 VDD.n108 4.5005
R2892 VDD.n96 VDD.n95 4.5005
R2893 VDD.n95 VDD.n94 4.5005
R2894 VDD.n7024 VDD.n7023 4.5005
R2895 VDD.n7007 VDD.n7006 4.5005
R2896 VDD.n7009 VDD.n7008 4.5005
R2897 VDD.n7010 VDD.n7009 4.5005
R2898 VDD.n48 VDD.n47 4.5005
R2899 VDD.n66 VDD.n64 4.5005
R2900 VDD.n55 VDD.n53 4.5005
R2901 VDD.n56 VDD.n55 4.5005
R2902 VDD.n7064 VDD.n42 4.5005
R2903 VDD.n44 VDD.n42 4.5005
R2904 VDD.n6878 VDD.n154 4.5005
R2905 VDD.n6955 VDD.n6954 4.5005
R2906 VDD.n130 VDD.n124 4.5005
R2907 VDD.n118 VDD.n117 4.5005
R2908 VDD.n117 VDD.n116 4.5005
R2909 VDD.n6935 VDD.n6934 4.5005
R2910 VDD.n144 VDD.n135 4.5005
R2911 VDD.n129 VDD.n128 4.5005
R2912 VDD.n128 VDD.n127 4.5005
R2913 VDD.n6913 VDD.n6912 4.5005
R2914 VDD.n6900 VDD.n140 4.5005
R2915 VDD.n6915 VDD.n6914 4.5005
R2916 VDD.n6915 VDD.n139 4.5005
R2917 VDD.n150 VDD.n149 4.5005
R2918 VDD.n151 VDD.n150 4.5005
R2919 VDD.n6898 VDD.n6897 4.5005
R2920 VDD.n104 VDD.n102 4.5005
R2921 VDD.n114 VDD.n104 4.5005
R2922 VDD.n161 VDD.n160 4.5005
R2923 VDD.n162 VDD.n161 4.5005
R2924 VDD.n6877 VDD.n6876 4.5005
R2925 VDD.n6652 VDD.n288 4.5005
R2926 VDD.n6729 VDD.n6728 4.5005
R2927 VDD.n264 VDD.n258 4.5005
R2928 VDD.n252 VDD.n251 4.5005
R2929 VDD.n251 VDD.n250 4.5005
R2930 VDD.n6709 VDD.n6708 4.5005
R2931 VDD.n278 VDD.n269 4.5005
R2932 VDD.n263 VDD.n262 4.5005
R2933 VDD.n262 VDD.n261 4.5005
R2934 VDD.n6687 VDD.n6686 4.5005
R2935 VDD.n6674 VDD.n274 4.5005
R2936 VDD.n6689 VDD.n6688 4.5005
R2937 VDD.n6689 VDD.n273 4.5005
R2938 VDD.n284 VDD.n283 4.5005
R2939 VDD.n285 VDD.n284 4.5005
R2940 VDD.n6672 VDD.n6671 4.5005
R2941 VDD.n238 VDD.n236 4.5005
R2942 VDD.n248 VDD.n238 4.5005
R2943 VDD.n295 VDD.n294 4.5005
R2944 VDD.n296 VDD.n295 4.5005
R2945 VDD.n6651 VDD.n6650 4.5005
R2946 VDD.n6426 VDD.n422 4.5005
R2947 VDD.n6503 VDD.n6502 4.5005
R2948 VDD.n398 VDD.n392 4.5005
R2949 VDD.n386 VDD.n385 4.5005
R2950 VDD.n385 VDD.n384 4.5005
R2951 VDD.n6483 VDD.n6482 4.5005
R2952 VDD.n412 VDD.n403 4.5005
R2953 VDD.n397 VDD.n396 4.5005
R2954 VDD.n396 VDD.n395 4.5005
R2955 VDD.n6461 VDD.n6460 4.5005
R2956 VDD.n6448 VDD.n408 4.5005
R2957 VDD.n6463 VDD.n6462 4.5005
R2958 VDD.n6463 VDD.n407 4.5005
R2959 VDD.n418 VDD.n417 4.5005
R2960 VDD.n419 VDD.n418 4.5005
R2961 VDD.n6446 VDD.n6445 4.5005
R2962 VDD.n372 VDD.n370 4.5005
R2963 VDD.n382 VDD.n372 4.5005
R2964 VDD.n429 VDD.n428 4.5005
R2965 VDD.n430 VDD.n429 4.5005
R2966 VDD.n6425 VDD.n6424 4.5005
R2967 VDD.n6222 VDD.n542 4.5005
R2968 VDD.n6277 VDD.n6276 4.5005
R2969 VDD.n532 VDD.n526 4.5005
R2970 VDD.n520 VDD.n519 4.5005
R2971 VDD.n519 VDD.n518 4.5005
R2972 VDD.n6257 VDD.n6256 4.5005
R2973 VDD.n546 VDD.n537 4.5005
R2974 VDD.n531 VDD.n530 4.5005
R2975 VDD.n530 VDD.n529 4.5005
R2976 VDD.n6237 VDD.n6236 4.5005
R2977 VDD.n6237 VDD.n541 4.5005
R2978 VDD.n6235 VDD.n6234 4.5005
R2979 VDD.n506 VDD.n504 4.5005
R2980 VDD.n516 VDD.n506 4.5005
R2981 VDD.n552 VDD.n551 4.5005
R2982 VDD.n553 VDD.n552 4.5005
R2983 VDD.n6200 VDD.n556 4.5005
R2984 VDD.n7171 VDD.n7170 4.5005
R2985 VDD.n7160 VDD.n7147 4.5005
R2986 VDD.n7174 VDD.n7160 4.5005
R2987 VDD.n7148 VDD.n8 4.5005
R2988 VDD.n7088 VDD.n7087 4.5005
R2989 VDD.n7214 VDD.n7213 4.5005
R2990 VDD.n7086 VDD.n7085 4.5005
R2991 VDD.n7084 VDD.n28 4.5005
R2992 VDD.n28 VDD.n25 4.5005
R2993 VDD.n7203 VDD.n7202 4.5005
R2994 VDD.n32 VDD.n30 4.5005
R2995 VDD.n7112 VDD.n7111 4.5005
R2996 VDD.n7113 VDD.n7112 4.5005
R2997 VDD.n7138 VDD.n7137 4.5005
R2998 VDD.n7201 VDD.n7200 4.5005
R2999 VDD.n7199 VDD.n7198 4.5005
R3000 VDD.n7198 VDD.n7197 4.5005
R3001 VDD.n7168 VDD.n7167 4.5005
R3002 VDD.n7123 VDD.n7121 4.5005
R3003 VDD.n7189 VDD.n7188 4.5005
R3004 VDD.n7189 VDD.n7120 4.5005
R3005 VDD.n2730 VDD.n2714 4.5005
R3006 VDD.n2729 VDD.n2728 4.5005
R3007 VDD.n4351 VDD.n4350 4.5005
R3008 VDD.n2725 VDD.n2687 4.5005
R3009 VDD.n2689 VDD.n2687 4.5005
R3010 VDD.n2685 VDD.n2683 4.5005
R3011 VDD.n4362 VDD.n4361 4.5005
R3012 VDD.n2704 VDD.n2703 4.5005
R3013 VDD.n2704 VDD.n2702 4.5005
R3014 VDD.n4364 VDD.n4363 4.5005
R3015 VDD.n2668 VDD.n2646 4.5005
R3016 VDD.n4366 VDD.n4365 4.5005
R3017 VDD.n4366 VDD.n2645 4.5005
R3018 VDD.n2666 VDD.n2665 4.5005
R3019 VDD.n4378 VDD.n4377 4.5005
R3020 VDD.n2662 VDD.n2444 4.5005
R3021 VDD.n2446 VDD.n2444 4.5005
R3022 VDD.n2442 VDD.n2440 4.5005
R3023 VDD.n2452 VDD.n2431 4.5005
R3024 VDD.n2635 VDD.n2634 4.5005
R3025 VDD.n2635 VDD.n2451 4.5005
R3026 VDD.n1420 VDD.n1399 4.5005
R3027 VDD.n4864 VDD.n4863 4.5005
R3028 VDD.n4864 VDD.n1398 4.5005
R3029 VDD.n4862 VDD.n4861 4.5005
R3030 VDD.n1418 VDD.n1417 4.5005
R3031 VDD.n1525 VDD.n1524 4.5005
R3032 VDD.n1523 VDD.n1520 4.5005
R3033 VDD.n1545 VDD.n1507 4.5005
R3034 VDD.n1645 VDD.n1644 4.5005
R3035 VDD.n1646 VDD.n1639 4.5005
R3036 VDD.n1682 VDD.n1681 4.5005
R3037 VDD.n1789 VDD.n1788 4.5005
R3038 VDD.n1787 VDD.n1784 4.5005
R3039 VDD.n1809 VDD.n1771 4.5005
R3040 VDD.n1909 VDD.n1908 4.5005
R3041 VDD.n1910 VDD.n1903 4.5005
R3042 VDD.n1946 VDD.n1945 4.5005
R3043 VDD.n2053 VDD.n2052 4.5005
R3044 VDD.n2051 VDD.n2048 4.5005
R3045 VDD.n2073 VDD.n2035 4.5005
R3046 VDD.n2173 VDD.n2172 4.5005
R3047 VDD.n2174 VDD.n2167 4.5005
R3048 VDD.n2210 VDD.n2209 4.5005
R3049 VDD.n2317 VDD.n2316 4.5005
R3050 VDD.n2315 VDD.n2312 4.5005
R3051 VDD.n2337 VDD.n2299 4.5005
R3052 VDD.n2421 VDD.n2391 4.5005
R3053 VDD.n2401 VDD.n2400 4.5005
R3054 VDD.n2390 VDD.n2388 4.5005
R3055 VDD.n2392 VDD.n2390 4.5005
R3056 VDD.n2398 VDD.n2397 4.5005
R3057 VDD.n2372 VDD.n2370 4.5005
R3058 VDD.n4427 VDD.n4426 4.5005
R3059 VDD.n4427 VDD.n2369 4.5005
R3060 VDD.n2379 VDD.n2349 4.5005
R3061 VDD.n2359 VDD.n2358 4.5005
R3062 VDD.n2348 VDD.n2346 4.5005
R3063 VDD.n2350 VDD.n2348 4.5005
R3064 VDD.n2356 VDD.n2355 4.5005
R3065 VDD.n2330 VDD.n2328 4.5005
R3066 VDD.n4449 VDD.n4448 4.5005
R3067 VDD.n4449 VDD.n2327 4.5005
R3068 VDD.n2414 VDD.n2412 4.5005
R3069 VDD.n4405 VDD.n4404 4.5005
R3070 VDD.n4405 VDD.n2411 4.5005
R3071 VDD.n2298 VDD.n2296 4.5005
R3072 VDD.n2300 VDD.n2298 4.5005
R3073 VDD.n4472 VDD.n4471 4.5005
R3074 VDD.n2281 VDD.n2259 4.5005
R3075 VDD.n4474 VDD.n4473 4.5005
R3076 VDD.n4474 VDD.n2258 4.5005
R3077 VDD.n2279 VDD.n2278 4.5005
R3078 VDD.n4486 VDD.n4485 4.5005
R3079 VDD.n2275 VDD.n2231 4.5005
R3080 VDD.n2233 VDD.n2231 4.5005
R3081 VDD.n2229 VDD.n2227 4.5005
R3082 VDD.n4497 VDD.n4496 4.5005
R3083 VDD.n2248 VDD.n2247 4.5005
R3084 VDD.n2248 VDD.n2246 4.5005
R3085 VDD.n4499 VDD.n4498 4.5005
R3086 VDD.n2212 VDD.n2195 4.5005
R3087 VDD.n4501 VDD.n4500 4.5005
R3088 VDD.n4501 VDD.n2194 4.5005
R3089 VDD.n4470 VDD.n4469 4.5005
R3090 VDD.n2319 VDD.n2318 4.5005
R3091 VDD.n2320 VDD.n2319 4.5005
R3092 VDD.n2175 VDD.n2168 4.5005
R3093 VDD.n2177 VDD.n2175 4.5005
R3094 VDD.n2157 VDD.n2127 4.5005
R3095 VDD.n2137 VDD.n2136 4.5005
R3096 VDD.n2126 VDD.n2124 4.5005
R3097 VDD.n2128 VDD.n2126 4.5005
R3098 VDD.n2134 VDD.n2133 4.5005
R3099 VDD.n2108 VDD.n2106 4.5005
R3100 VDD.n4548 VDD.n4547 4.5005
R3101 VDD.n4548 VDD.n2105 4.5005
R3102 VDD.n2115 VDD.n2085 4.5005
R3103 VDD.n2095 VDD.n2094 4.5005
R3104 VDD.n2084 VDD.n2082 4.5005
R3105 VDD.n2086 VDD.n2084 4.5005
R3106 VDD.n2092 VDD.n2091 4.5005
R3107 VDD.n2066 VDD.n2064 4.5005
R3108 VDD.n4570 VDD.n4569 4.5005
R3109 VDD.n4570 VDD.n2063 4.5005
R3110 VDD.n2150 VDD.n2148 4.5005
R3111 VDD.n4526 VDD.n4525 4.5005
R3112 VDD.n4526 VDD.n2147 4.5005
R3113 VDD.n2034 VDD.n2032 4.5005
R3114 VDD.n2036 VDD.n2034 4.5005
R3115 VDD.n4593 VDD.n4592 4.5005
R3116 VDD.n2017 VDD.n1995 4.5005
R3117 VDD.n4595 VDD.n4594 4.5005
R3118 VDD.n4595 VDD.n1994 4.5005
R3119 VDD.n2015 VDD.n2014 4.5005
R3120 VDD.n4607 VDD.n4606 4.5005
R3121 VDD.n2011 VDD.n1967 4.5005
R3122 VDD.n1969 VDD.n1967 4.5005
R3123 VDD.n1965 VDD.n1963 4.5005
R3124 VDD.n4618 VDD.n4617 4.5005
R3125 VDD.n1984 VDD.n1983 4.5005
R3126 VDD.n1984 VDD.n1982 4.5005
R3127 VDD.n4620 VDD.n4619 4.5005
R3128 VDD.n1948 VDD.n1931 4.5005
R3129 VDD.n4622 VDD.n4621 4.5005
R3130 VDD.n4622 VDD.n1930 4.5005
R3131 VDD.n4591 VDD.n4590 4.5005
R3132 VDD.n2055 VDD.n2054 4.5005
R3133 VDD.n2056 VDD.n2055 4.5005
R3134 VDD.n1911 VDD.n1904 4.5005
R3135 VDD.n1913 VDD.n1911 4.5005
R3136 VDD.n1893 VDD.n1863 4.5005
R3137 VDD.n1873 VDD.n1872 4.5005
R3138 VDD.n1862 VDD.n1860 4.5005
R3139 VDD.n1864 VDD.n1862 4.5005
R3140 VDD.n1870 VDD.n1869 4.5005
R3141 VDD.n1844 VDD.n1842 4.5005
R3142 VDD.n4669 VDD.n4668 4.5005
R3143 VDD.n4669 VDD.n1841 4.5005
R3144 VDD.n1851 VDD.n1821 4.5005
R3145 VDD.n1831 VDD.n1830 4.5005
R3146 VDD.n1820 VDD.n1818 4.5005
R3147 VDD.n1822 VDD.n1820 4.5005
R3148 VDD.n1828 VDD.n1827 4.5005
R3149 VDD.n1802 VDD.n1800 4.5005
R3150 VDD.n4691 VDD.n4690 4.5005
R3151 VDD.n4691 VDD.n1799 4.5005
R3152 VDD.n1886 VDD.n1884 4.5005
R3153 VDD.n4647 VDD.n4646 4.5005
R3154 VDD.n4647 VDD.n1883 4.5005
R3155 VDD.n1770 VDD.n1768 4.5005
R3156 VDD.n1772 VDD.n1770 4.5005
R3157 VDD.n4714 VDD.n4713 4.5005
R3158 VDD.n1753 VDD.n1731 4.5005
R3159 VDD.n4716 VDD.n4715 4.5005
R3160 VDD.n4716 VDD.n1730 4.5005
R3161 VDD.n1751 VDD.n1750 4.5005
R3162 VDD.n4728 VDD.n4727 4.5005
R3163 VDD.n1747 VDD.n1703 4.5005
R3164 VDD.n1705 VDD.n1703 4.5005
R3165 VDD.n1701 VDD.n1699 4.5005
R3166 VDD.n4739 VDD.n4738 4.5005
R3167 VDD.n1720 VDD.n1719 4.5005
R3168 VDD.n1720 VDD.n1718 4.5005
R3169 VDD.n4741 VDD.n4740 4.5005
R3170 VDD.n1684 VDD.n1667 4.5005
R3171 VDD.n4743 VDD.n4742 4.5005
R3172 VDD.n4743 VDD.n1666 4.5005
R3173 VDD.n4712 VDD.n4711 4.5005
R3174 VDD.n1791 VDD.n1790 4.5005
R3175 VDD.n1792 VDD.n1791 4.5005
R3176 VDD.n1647 VDD.n1640 4.5005
R3177 VDD.n1649 VDD.n1647 4.5005
R3178 VDD.n1629 VDD.n1599 4.5005
R3179 VDD.n1609 VDD.n1608 4.5005
R3180 VDD.n1598 VDD.n1596 4.5005
R3181 VDD.n1600 VDD.n1598 4.5005
R3182 VDD.n1606 VDD.n1605 4.5005
R3183 VDD.n1580 VDD.n1578 4.5005
R3184 VDD.n4790 VDD.n4789 4.5005
R3185 VDD.n4790 VDD.n1577 4.5005
R3186 VDD.n1587 VDD.n1557 4.5005
R3187 VDD.n1567 VDD.n1566 4.5005
R3188 VDD.n1556 VDD.n1554 4.5005
R3189 VDD.n1558 VDD.n1556 4.5005
R3190 VDD.n1564 VDD.n1563 4.5005
R3191 VDD.n1538 VDD.n1536 4.5005
R3192 VDD.n4812 VDD.n4811 4.5005
R3193 VDD.n4812 VDD.n1535 4.5005
R3194 VDD.n1622 VDD.n1620 4.5005
R3195 VDD.n4768 VDD.n4767 4.5005
R3196 VDD.n4768 VDD.n1619 4.5005
R3197 VDD.n1506 VDD.n1504 4.5005
R3198 VDD.n1508 VDD.n1506 4.5005
R3199 VDD.n4835 VDD.n4834 4.5005
R3200 VDD.n1489 VDD.n1467 4.5005
R3201 VDD.n4837 VDD.n4836 4.5005
R3202 VDD.n4837 VDD.n1466 4.5005
R3203 VDD.n1487 VDD.n1486 4.5005
R3204 VDD.n4849 VDD.n4848 4.5005
R3205 VDD.n1483 VDD.n1439 4.5005
R3206 VDD.n1441 VDD.n1439 4.5005
R3207 VDD.n1437 VDD.n1435 4.5005
R3208 VDD.n4860 VDD.n4859 4.5005
R3209 VDD.n1456 VDD.n1455 4.5005
R3210 VDD.n1456 VDD.n1454 4.5005
R3211 VDD.n4833 VDD.n4832 4.5005
R3212 VDD.n1527 VDD.n1526 4.5005
R3213 VDD.n1528 VDD.n1527 4.5005
R3214 VDD.n1414 VDD.n1378 4.5005
R3215 VDD.n1380 VDD.n1378 4.5005
R3216 VDD.n4885 VDD.n4884 4.5005
R3217 VDD.n4887 VDD.n4886 4.5005
R3218 VDD.n1362 VDD.n1340 4.5005
R3219 VDD.n4889 VDD.n4888 4.5005
R3220 VDD.n4889 VDD.n1339 4.5005
R3221 VDD.n1360 VDD.n1359 4.5005
R3222 VDD.n4901 VDD.n4900 4.5005
R3223 VDD.n1356 VDD.n1312 4.5005
R3224 VDD.n1314 VDD.n1312 4.5005
R3225 VDD.n1310 VDD.n1308 4.5005
R3226 VDD.n4912 VDD.n4911 4.5005
R3227 VDD.n1329 VDD.n1328 4.5005
R3228 VDD.n1329 VDD.n1327 4.5005
R3229 VDD.n4914 VDD.n4913 4.5005
R3230 VDD.n1293 VDD.n1251 4.5005
R3231 VDD.n4916 VDD.n4915 4.5005
R3232 VDD.n4916 VDD.n1250 4.5005
R3233 VDD.n1291 VDD.n1290 4.5005
R3234 VDD.n1276 VDD.n1275 4.5005
R3235 VDD.n1287 VDD.n1286 4.5005
R3236 VDD.n1287 VDD.n1244 4.5005
R3237 VDD.n2471 VDD.n2470 4.5005
R3238 VDD.n2481 VDD.n2480 4.5005
R3239 VDD.n2479 VDD.n2478 4.5005
R3240 VDD.n2751 VDD.n2748 4.5005
R3241 VDD.n2792 VDD.n2791 4.5005
R3242 VDD.n2766 VDD.n2765 4.5005
R3243 VDD.n4284 VDD.n4283 4.5005
R3244 VDD.n4282 VDD.n2844 4.5005
R3245 VDD.n2897 VDD.n2896 4.5005
R3246 VDD.n2997 VDD.n2996 4.5005
R3247 VDD.n2998 VDD.n2991 4.5005
R3248 VDD.n3034 VDD.n3033 4.5005
R3249 VDD.n3141 VDD.n3140 4.5005
R3250 VDD.n3139 VDD.n3136 4.5005
R3251 VDD.n3163 VDD.n3123 4.5005
R3252 VDD.n3263 VDD.n3262 4.5005
R3253 VDD.n3264 VDD.n3257 4.5005
R3254 VDD.n3300 VDD.n3299 4.5005
R3255 VDD.n3407 VDD.n3406 4.5005
R3256 VDD.n3405 VDD.n3402 4.5005
R3257 VDD.n3429 VDD.n3389 4.5005
R3258 VDD.n3529 VDD.n3528 4.5005
R3259 VDD.n3530 VDD.n3523 4.5005
R3260 VDD.n3566 VDD.n3565 4.5005
R3261 VDD.n3673 VDD.n3672 4.5005
R3262 VDD.n3671 VDD.n3668 4.5005
R3263 VDD.n3695 VDD.n3655 4.5005
R3264 VDD.n3779 VDD.n3750 4.5005
R3265 VDD.n3759 VDD.n3758 4.5005
R3266 VDD.n3756 VDD.n3731 4.5005
R3267 VDD.n3729 VDD.n3727 4.5005
R3268 VDD.n3738 VDD.n3707 4.5005
R3269 VDD.n3716 VDD.n3715 4.5005
R3270 VDD.n3713 VDD.n3688 4.5005
R3271 VDD.n3686 VDD.n3684 4.5005
R3272 VDD.n3772 VDD.n3770 4.5005
R3273 VDD.n3935 VDD.n3934 4.5005
R3274 VDD.n3637 VDD.n3615 4.5005
R3275 VDD.n3635 VDD.n3634 4.5005
R3276 VDD.n3949 VDD.n3948 4.5005
R3277 VDD.n3585 VDD.n3583 4.5005
R3278 VDD.n3960 VDD.n3959 4.5005
R3279 VDD.n3962 VDD.n3961 4.5005
R3280 VDD.n3568 VDD.n3551 4.5005
R3281 VDD.n3933 VDD.n3932 4.5005
R3282 VDD.n3513 VDD.n3484 4.5005
R3283 VDD.n3493 VDD.n3492 4.5005
R3284 VDD.n3490 VDD.n3465 4.5005
R3285 VDD.n3463 VDD.n3461 4.5005
R3286 VDD.n3472 VDD.n3441 4.5005
R3287 VDD.n3450 VDD.n3449 4.5005
R3288 VDD.n3447 VDD.n3422 4.5005
R3289 VDD.n3420 VDD.n3418 4.5005
R3290 VDD.n3506 VDD.n3504 4.5005
R3291 VDD.n4054 VDD.n4053 4.5005
R3292 VDD.n3371 VDD.n3349 4.5005
R3293 VDD.n3369 VDD.n3368 4.5005
R3294 VDD.n4068 VDD.n4067 4.5005
R3295 VDD.n3319 VDD.n3317 4.5005
R3296 VDD.n4079 VDD.n4078 4.5005
R3297 VDD.n4081 VDD.n4080 4.5005
R3298 VDD.n3302 VDD.n3285 4.5005
R3299 VDD.n4052 VDD.n4051 4.5005
R3300 VDD.n3247 VDD.n3218 4.5005
R3301 VDD.n3227 VDD.n3226 4.5005
R3302 VDD.n3224 VDD.n3199 4.5005
R3303 VDD.n3197 VDD.n3195 4.5005
R3304 VDD.n3206 VDD.n3175 4.5005
R3305 VDD.n3184 VDD.n3183 4.5005
R3306 VDD.n3181 VDD.n3156 4.5005
R3307 VDD.n3154 VDD.n3152 4.5005
R3308 VDD.n3240 VDD.n3238 4.5005
R3309 VDD.n4173 VDD.n4172 4.5005
R3310 VDD.n3105 VDD.n3083 4.5005
R3311 VDD.n3103 VDD.n3102 4.5005
R3312 VDD.n4187 VDD.n4186 4.5005
R3313 VDD.n3053 VDD.n3051 4.5005
R3314 VDD.n4198 VDD.n4197 4.5005
R3315 VDD.n4200 VDD.n4199 4.5005
R3316 VDD.n3036 VDD.n3019 4.5005
R3317 VDD.n4171 VDD.n4170 4.5005
R3318 VDD.n2981 VDD.n2952 4.5005
R3319 VDD.n2961 VDD.n2960 4.5005
R3320 VDD.n2958 VDD.n2933 4.5005
R3321 VDD.n2931 VDD.n2929 4.5005
R3322 VDD.n2940 VDD.n2909 4.5005
R3323 VDD.n2918 VDD.n2917 4.5005
R3324 VDD.n2915 VDD.n2858 4.5005
R3325 VDD.n2856 VDD.n2854 4.5005
R3326 VDD.n2974 VDD.n2972 4.5005
R3327 VDD.n2880 VDD.n2879 4.5005
R3328 VDD.n4298 VDD.n4297 4.5005
R3329 VDD.n2811 VDD.n2809 4.5005
R3330 VDD.n4309 VDD.n4308 4.5005
R3331 VDD.n4311 VDD.n4310 4.5005
R3332 VDD.n2794 VDD.n2777 4.5005
R3333 VDD.n2882 VDD.n2841 4.5005
R3334 VDD.n2752 VDD.n2749 4.5005
R3335 VDD.n2754 VDD.n2752 4.5005
R3336 VDD.n3749 VDD.n3747 4.5005
R3337 VDD.n3751 VDD.n3749 4.5005
R3338 VDD.n3891 VDD.n3890 4.5005
R3339 VDD.n3891 VDD.n3726 4.5005
R3340 VDD.n3706 VDD.n3704 4.5005
R3341 VDD.n3708 VDD.n3706 4.5005
R3342 VDD.n3912 VDD.n3911 4.5005
R3343 VDD.n3912 VDD.n3683 4.5005
R3344 VDD.n3870 VDD.n3869 4.5005
R3345 VDD.n3870 VDD.n3769 4.5005
R3346 VDD.n3654 VDD.n3652 4.5005
R3347 VDD.n3656 VDD.n3654 4.5005
R3348 VDD.n3937 VDD.n3936 4.5005
R3349 VDD.n3937 VDD.n3614 4.5005
R3350 VDD.n3631 VDD.n3587 4.5005
R3351 VDD.n3589 VDD.n3587 4.5005
R3352 VDD.n3604 VDD.n3603 4.5005
R3353 VDD.n3604 VDD.n3602 4.5005
R3354 VDD.n3964 VDD.n3963 4.5005
R3355 VDD.n3964 VDD.n3550 4.5005
R3356 VDD.n3675 VDD.n3674 4.5005
R3357 VDD.n3676 VDD.n3675 4.5005
R3358 VDD.n3531 VDD.n3525 4.5005
R3359 VDD.n3533 VDD.n3531 4.5005
R3360 VDD.n3483 VDD.n3481 4.5005
R3361 VDD.n3485 VDD.n3483 4.5005
R3362 VDD.n4010 VDD.n4009 4.5005
R3363 VDD.n4010 VDD.n3460 4.5005
R3364 VDD.n3440 VDD.n3438 4.5005
R3365 VDD.n3442 VDD.n3440 4.5005
R3366 VDD.n4031 VDD.n4030 4.5005
R3367 VDD.n4031 VDD.n3417 4.5005
R3368 VDD.n3989 VDD.n3988 4.5005
R3369 VDD.n3989 VDD.n3503 4.5005
R3370 VDD.n3388 VDD.n3386 4.5005
R3371 VDD.n3390 VDD.n3388 4.5005
R3372 VDD.n4056 VDD.n4055 4.5005
R3373 VDD.n4056 VDD.n3348 4.5005
R3374 VDD.n3365 VDD.n3321 4.5005
R3375 VDD.n3323 VDD.n3321 4.5005
R3376 VDD.n3338 VDD.n3337 4.5005
R3377 VDD.n3338 VDD.n3336 4.5005
R3378 VDD.n4083 VDD.n4082 4.5005
R3379 VDD.n4083 VDD.n3284 4.5005
R3380 VDD.n3409 VDD.n3408 4.5005
R3381 VDD.n3410 VDD.n3409 4.5005
R3382 VDD.n3265 VDD.n3259 4.5005
R3383 VDD.n3267 VDD.n3265 4.5005
R3384 VDD.n3217 VDD.n3215 4.5005
R3385 VDD.n3219 VDD.n3217 4.5005
R3386 VDD.n4129 VDD.n4128 4.5005
R3387 VDD.n4129 VDD.n3194 4.5005
R3388 VDD.n3174 VDD.n3172 4.5005
R3389 VDD.n3176 VDD.n3174 4.5005
R3390 VDD.n4150 VDD.n4149 4.5005
R3391 VDD.n4150 VDD.n3151 4.5005
R3392 VDD.n4108 VDD.n4107 4.5005
R3393 VDD.n4108 VDD.n3237 4.5005
R3394 VDD.n3122 VDD.n3120 4.5005
R3395 VDD.n3124 VDD.n3122 4.5005
R3396 VDD.n4175 VDD.n4174 4.5005
R3397 VDD.n4175 VDD.n3082 4.5005
R3398 VDD.n3099 VDD.n3055 4.5005
R3399 VDD.n3057 VDD.n3055 4.5005
R3400 VDD.n3072 VDD.n3071 4.5005
R3401 VDD.n3072 VDD.n3070 4.5005
R3402 VDD.n4202 VDD.n4201 4.5005
R3403 VDD.n4202 VDD.n3018 4.5005
R3404 VDD.n3143 VDD.n3142 4.5005
R3405 VDD.n3144 VDD.n3143 4.5005
R3406 VDD.n2999 VDD.n2993 4.5005
R3407 VDD.n3001 VDD.n2999 4.5005
R3408 VDD.n2951 VDD.n2949 4.5005
R3409 VDD.n2953 VDD.n2951 4.5005
R3410 VDD.n4248 VDD.n4247 4.5005
R3411 VDD.n4248 VDD.n2928 4.5005
R3412 VDD.n2908 VDD.n2906 4.5005
R3413 VDD.n2910 VDD.n2908 4.5005
R3414 VDD.n4269 VDD.n4268 4.5005
R3415 VDD.n4269 VDD.n2853 4.5005
R3416 VDD.n4227 VDD.n4226 4.5005
R3417 VDD.n4227 VDD.n2971 4.5005
R3418 VDD.n2863 VDD.n2845 4.5005
R3419 VDD.n4279 VDD.n2845 4.5005
R3420 VDD.n2876 VDD.n2813 4.5005
R3421 VDD.n2815 VDD.n2813 4.5005
R3422 VDD.n2830 VDD.n2829 4.5005
R3423 VDD.n2830 VDD.n2828 4.5005
R3424 VDD.n4313 VDD.n4312 4.5005
R3425 VDD.n4313 VDD.n2776 4.5005
R3426 VDD.n4286 VDD.n4285 4.5005
R3427 VDD.n4286 VDD.n2840 4.5005
R3428 VDD.n2741 VDD.n2740 4.5005
R3429 VDD.n2763 VDD.n2740 4.5005
R3430 VDD.n4943 VDD.n1234 4.5005
R3431 VDD.n4963 VDD.n4962 4.5005
R3432 VDD.n4961 VDD.n4960 4.5005
R3433 VDD.n1193 VDD.n1187 4.5005
R3434 VDD.n5067 VDD.n5066 4.5005
R3435 VDD.n5037 VDD.n5036 4.5005
R3436 VDD.n1145 VDD.n1144 4.5005
R3437 VDD.n1143 VDD.n1132 4.5005
R3438 VDD.n5146 VDD.n5145 4.5005
R3439 VDD.n5241 VDD.n5240 4.5005
R3440 VDD.n1070 VDD.n1063 4.5005
R3441 VDD.n5265 VDD.n5264 4.5005
R3442 VDD.n1010 VDD.n1009 4.5005
R3443 VDD.n1008 VDD.n997 4.5005
R3444 VDD.n5374 VDD.n5373 4.5005
R3445 VDD.n5469 VDD.n5468 4.5005
R3446 VDD.n935 VDD.n928 4.5005
R3447 VDD.n5493 VDD.n5492 4.5005
R3448 VDD.n875 VDD.n874 4.5005
R3449 VDD.n873 VDD.n862 4.5005
R3450 VDD.n5602 VDD.n5601 4.5005
R3451 VDD.n5697 VDD.n5696 4.5005
R3452 VDD.n800 VDD.n793 4.5005
R3453 VDD.n5721 VDD.n5720 4.5005
R3454 VDD.n740 VDD.n739 4.5005
R3455 VDD.n738 VDD.n737 4.5005
R3456 VDD.n723 VDD.n722 4.5005
R3457 VDD.n5914 VDD.n5913 4.5005
R3458 VDD.n5892 VDD.n5891 4.5005
R3459 VDD.n5894 VDD.n5893 4.5005
R3460 VDD.n5877 VDD.n5876 4.5005
R3461 VDD.n5875 VDD.n5874 4.5005
R3462 VDD.n5858 VDD.n5857 4.5005
R3463 VDD.n707 VDD.n705 4.5005
R3464 VDD.n5833 VDD.n5832 4.5005
R3465 VDD.n684 VDD.n681 4.5005
R3466 VDD.n5803 VDD.n5802 4.5005
R3467 VDD.n762 VDD.n753 4.5005
R3468 VDD.n5780 VDD.n5779 4.5005
R3469 VDD.n5767 VDD.n758 4.5005
R3470 VDD.n5765 VDD.n5764 4.5005
R3471 VDD.n776 VDD.n774 4.5005
R3472 VDD.n5751 VDD.n5750 4.5005
R3473 VDD.n788 VDD.n782 4.5005
R3474 VDD.n748 VDD.n732 4.5005
R3475 VDD.n5677 VDD.n5676 4.5005
R3476 VDD.n5658 VDD.n815 4.5005
R3477 VDD.n825 VDD.n816 4.5005
R3478 VDD.n836 VDD.n834 4.5005
R3479 VDD.n5637 VDD.n5636 4.5005
R3480 VDD.n5619 VDD.n5618 4.5005
R3481 VDD.n5621 VDD.n5620 4.5005
R3482 VDD.n5604 VDD.n5603 4.5005
R3483 VDD.n5675 VDD.n5674 4.5005
R3484 VDD.n5576 VDD.n5575 4.5005
R3485 VDD.n897 VDD.n888 4.5005
R3486 VDD.n5552 VDD.n5551 4.5005
R3487 VDD.n5539 VDD.n893 4.5005
R3488 VDD.n5537 VDD.n5536 4.5005
R3489 VDD.n911 VDD.n909 4.5005
R3490 VDD.n5523 VDD.n5522 4.5005
R3491 VDD.n923 VDD.n917 4.5005
R3492 VDD.n883 VDD.n858 4.5005
R3493 VDD.n5449 VDD.n5448 4.5005
R3494 VDD.n5430 VDD.n950 4.5005
R3495 VDD.n960 VDD.n951 4.5005
R3496 VDD.n971 VDD.n969 4.5005
R3497 VDD.n5409 VDD.n5408 4.5005
R3498 VDD.n5391 VDD.n5390 4.5005
R3499 VDD.n5393 VDD.n5392 4.5005
R3500 VDD.n5376 VDD.n5375 4.5005
R3501 VDD.n5447 VDD.n5446 4.5005
R3502 VDD.n5348 VDD.n5347 4.5005
R3503 VDD.n1032 VDD.n1023 4.5005
R3504 VDD.n5324 VDD.n5323 4.5005
R3505 VDD.n5311 VDD.n1028 4.5005
R3506 VDD.n5309 VDD.n5308 4.5005
R3507 VDD.n1046 VDD.n1044 4.5005
R3508 VDD.n5295 VDD.n5294 4.5005
R3509 VDD.n1058 VDD.n1052 4.5005
R3510 VDD.n1018 VDD.n993 4.5005
R3511 VDD.n5221 VDD.n5220 4.5005
R3512 VDD.n5202 VDD.n1085 4.5005
R3513 VDD.n1095 VDD.n1086 4.5005
R3514 VDD.n1106 VDD.n1104 4.5005
R3515 VDD.n5181 VDD.n5180 4.5005
R3516 VDD.n5163 VDD.n5162 4.5005
R3517 VDD.n5165 VDD.n5164 4.5005
R3518 VDD.n5148 VDD.n5147 4.5005
R3519 VDD.n5219 VDD.n5218 4.5005
R3520 VDD.n5120 VDD.n5119 4.5005
R3521 VDD.n1167 VDD.n1158 4.5005
R3522 VDD.n5096 VDD.n5095 4.5005
R3523 VDD.n5083 VDD.n1163 4.5005
R3524 VDD.n5081 VDD.n5080 4.5005
R3525 VDD.n1181 VDD.n1179 4.5005
R3526 VDD.n1153 VDD.n1128 4.5005
R3527 VDD.n1180 VDD.n1178 4.5005
R3528 VDD.n1178 VDD.n1177 4.5005
R3529 VDD.n5890 VDD.n677 4.5005
R3530 VDD.n677 VDD.n676 4.5005
R3531 VDD.n5879 VDD.n5878 4.5005
R3532 VDD.n5880 VDD.n5879 4.5005
R3533 VDD.n708 VDD.n706 4.5005
R3534 VDD.n5854 VDD.n708 4.5005
R3535 VDD.n718 VDD.n717 4.5005
R3536 VDD.n717 VDD.n716 4.5005
R3537 VDD.n683 VDD.n671 4.5005
R3538 VDD.n673 VDD.n671 4.5005
R3539 VDD.n726 VDD.n725 4.5005
R3540 VDD.n725 VDD.n724 4.5005
R3541 VDD.n747 VDD.n746 4.5005
R3542 VDD.n746 VDD.n745 4.5005
R3543 VDD.n5782 VDD.n5781 4.5005
R3544 VDD.n5782 VDD.n757 4.5005
R3545 VDD.n768 VDD.n767 4.5005
R3546 VDD.n769 VDD.n768 4.5005
R3547 VDD.n775 VDD.n773 4.5005
R3548 VDD.n773 VDD.n772 4.5005
R3549 VDD.n733 VDD.n731 4.5005
R3550 VDD.n743 VDD.n733 4.5005
R3551 VDD.n787 VDD.n786 4.5005
R3552 VDD.n786 VDD.n785 4.5005
R3553 VDD.n5660 VDD.n5659 4.5005
R3554 VDD.n5660 VDD.n814 4.5005
R3555 VDD.n824 VDD.n822 4.5005
R3556 VDD.n826 VDD.n824 4.5005
R3557 VDD.n5617 VDD.n830 4.5005
R3558 VDD.n830 VDD.n829 4.5005
R3559 VDD.n5606 VDD.n5605 4.5005
R3560 VDD.n5607 VDD.n5606 4.5005
R3561 VDD.n5673 VDD.n797 4.5005
R3562 VDD.n797 VDD.n796 4.5005
R3563 VDD.n872 VDD.n871 4.5005
R3564 VDD.n871 VDD.n870 4.5005
R3565 VDD.n882 VDD.n881 4.5005
R3566 VDD.n881 VDD.n880 4.5005
R3567 VDD.n5554 VDD.n5553 4.5005
R3568 VDD.n5554 VDD.n892 4.5005
R3569 VDD.n903 VDD.n902 4.5005
R3570 VDD.n904 VDD.n903 4.5005
R3571 VDD.n910 VDD.n908 4.5005
R3572 VDD.n908 VDD.n907 4.5005
R3573 VDD.n859 VDD.n857 4.5005
R3574 VDD.n878 VDD.n859 4.5005
R3575 VDD.n922 VDD.n921 4.5005
R3576 VDD.n921 VDD.n920 4.5005
R3577 VDD.n5432 VDD.n5431 4.5005
R3578 VDD.n5432 VDD.n949 4.5005
R3579 VDD.n959 VDD.n957 4.5005
R3580 VDD.n961 VDD.n959 4.5005
R3581 VDD.n5389 VDD.n965 4.5005
R3582 VDD.n965 VDD.n964 4.5005
R3583 VDD.n5378 VDD.n5377 4.5005
R3584 VDD.n5379 VDD.n5378 4.5005
R3585 VDD.n5445 VDD.n932 4.5005
R3586 VDD.n932 VDD.n931 4.5005
R3587 VDD.n1007 VDD.n1006 4.5005
R3588 VDD.n1006 VDD.n1005 4.5005
R3589 VDD.n1017 VDD.n1016 4.5005
R3590 VDD.n1016 VDD.n1015 4.5005
R3591 VDD.n5326 VDD.n5325 4.5005
R3592 VDD.n5326 VDD.n1027 4.5005
R3593 VDD.n1038 VDD.n1037 4.5005
R3594 VDD.n1039 VDD.n1038 4.5005
R3595 VDD.n1045 VDD.n1043 4.5005
R3596 VDD.n1043 VDD.n1042 4.5005
R3597 VDD.n994 VDD.n992 4.5005
R3598 VDD.n1013 VDD.n994 4.5005
R3599 VDD.n1057 VDD.n1056 4.5005
R3600 VDD.n1056 VDD.n1055 4.5005
R3601 VDD.n5204 VDD.n5203 4.5005
R3602 VDD.n5204 VDD.n1084 4.5005
R3603 VDD.n1094 VDD.n1092 4.5005
R3604 VDD.n1096 VDD.n1094 4.5005
R3605 VDD.n5161 VDD.n1100 4.5005
R3606 VDD.n1100 VDD.n1099 4.5005
R3607 VDD.n5150 VDD.n5149 4.5005
R3608 VDD.n5151 VDD.n5150 4.5005
R3609 VDD.n5217 VDD.n1067 4.5005
R3610 VDD.n1067 VDD.n1066 4.5005
R3611 VDD.n1142 VDD.n1141 4.5005
R3612 VDD.n1141 VDD.n1140 4.5005
R3613 VDD.n1152 VDD.n1151 4.5005
R3614 VDD.n1151 VDD.n1150 4.5005
R3615 VDD.n5098 VDD.n5097 4.5005
R3616 VDD.n5098 VDD.n1162 4.5005
R3617 VDD.n1173 VDD.n1172 4.5005
R3618 VDD.n1174 VDD.n1173 4.5005
R3619 VDD.n1129 VDD.n1127 4.5005
R3620 VDD.n1148 VDD.n1129 4.5005
R3621 VDD.n1192 VDD.n1191 4.5005
R3622 VDD.n1191 VDD.n1190 4.5005
R3623 VDD.n6073 VDD 4.28667
R3624 VDD.n7223 VDD 4.28667
R3625 VDD.n2596 VDD.n2595 3.92207
R3626 VDD.n6125 VDD.n605 3.81576
R3627 VDD.n3825 VDD.n3808 3.67129
R3628 VDD.n2541 VDD.n2487 3.67129
R3629 VDD.n6160 VDD.n6159 3.52129
R3630 VDD.n6087 VDD.n632 3.46788
R3631 VDD.n6134 VDD.n6133 3.46651
R3632 VDD.n2616 VDD.n2615 3.46651
R3633 VDD.n2604 VDD.n2466 3.46651
R3634 VDD.n4952 VDD.n4951 3.46651
R3635 VDD.n4975 VDD.n1232 3.46651
R3636 VDD.n3804 VDD.n3802 3.46575
R3637 VDD.n3812 VDD.n3798 3.46575
R3638 VDD.n3815 VDD.n3794 3.46575
R3639 VDD.n3809 VDD.n3790 3.46575
R3640 VDD.n3805 VDD.n3786 3.46575
R3641 VDD.n2578 VDD.n2577 3.46575
R3642 VDD.n2572 VDD.n2571 3.46575
R3643 VDD.n2589 VDD.n2567 3.46575
R3644 VDD.n2534 VDD.n2532 3.46575
R3645 VDD.n2501 VDD.n2499 3.46575
R3646 VDD.n2494 VDD.n2493 3.46575
R3647 VDD.n2556 VDD.n2489 3.46575
R3648 VDD.n2549 VDD.n2530 3.46575
R3649 VDD.n6178 VDD.n6177 3.46323
R3650 VDD.n5017 VDD.n5016 3.46323
R3651 VDD.n3832 VDD.n3831 3.46323
R3652 VDD.n2508 VDD.n2507 3.46323
R3653 VDD.n597 VDD.n591 3.46321
R3654 VDD.n3841 VDD.n3835 3.46321
R3655 VDD.n2517 VDD.n2511 3.46321
R3656 VDD.n1227 VDD.n1221 3.46321
R3657 VDD.n6109 VDD.n6108 3.45407
R3658 VDD.n624 VDD.n616 3.45407
R3659 VDD.n6101 VDD.n6100 3.45407
R3660 VDD.n6153 VDD.n6149 3.45407
R3661 VDD.n6165 VDD.n6164 3.45407
R3662 VDD.n6144 VDD.n6142 3.45407
R3663 VDD.n586 VDD.n582 3.45407
R3664 VDD.n6173 VDD.n6172 3.45407
R3665 VDD.n5012 VDD.n5011 3.45407
R3666 VDD.n4996 VDD.n4992 3.45407
R3667 VDD.n5004 VDD.n5003 3.45407
R3668 VDD.n4987 VDD.n4985 3.45407
R3669 VDD.n1216 VDD.n1212 3.45407
R3670 VDD.n6106 VDD.n6105 3.44028
R3671 VDD.n622 VDD.n621 3.44028
R3672 VDD.n6098 VDD.n628 3.44028
R3673 VDD.n6150 VDD.n6148 3.44028
R3674 VDD.n6162 VDD.n577 3.44028
R3675 VDD.n6141 VDD.n6140 3.44028
R3676 VDD.n583 VDD.n581 3.44028
R3677 VDD.n6170 VDD.n6169 3.44028
R3678 VDD.n5009 VDD.n5008 3.44028
R3679 VDD.n4993 VDD.n4991 3.44028
R3680 VDD.n5001 VDD.n1207 3.44028
R3681 VDD.n4984 VDD.n4983 3.44028
R3682 VDD.n1213 VDD.n1211 3.44028
R3683 VDD.n3828 VDD.n3827 3.4393
R3684 VDD.n3813 VDD.n3800 3.4393
R3685 VDD.n3816 VDD.n3796 3.4393
R3686 VDD.n3810 VDD.n3792 3.4393
R3687 VDD.n3806 VDD.n3788 3.4393
R3688 VDD.n2581 VDD.n2580 3.4393
R3689 VDD.n2575 VDD.n2574 3.4393
R3690 VDD.n2592 VDD.n2591 3.4393
R3691 VDD.n2544 VDD.n2543 3.4393
R3692 VDD.n2504 VDD.n2503 3.4393
R3693 VDD.n2497 VDD.n2496 3.4393
R3694 VDD.n2559 VDD.n2558 3.4393
R3695 VDD.n2552 VDD.n2551 3.4393
R3696 VDD.n4338 VDD.n4337 3.43054
R3697 VDD.n4879 VDD.n4878 3.43054
R3698 VDD.n5930 VDD.n5929 3.42985
R3699 VDD.n7080 VDD.n7079 3.42985
R3700 VDD.n2470 VDD.n2463 3.42739
R3701 VDD.n4944 VDD.n4943 3.42739
R3702 VDD.n7231 VDD.n7230 3.42653
R3703 VDD.n6116 VDD.n611 3.4257
R3704 VDD.n6176 VDD.n6175 3.42476
R3705 VDD.n5015 VDD.n5014 3.42476
R3706 VDD.n6081 VDD.n6080 3.42443
R3707 VDD.n4393 VDD.n4392 3.42443
R3708 VDD.n1272 VDD.n1229 3.42443
R3709 VDD.n6182 VDD.n565 3.42376
R3710 VDD.n7075 VDD.n7074 3.42376
R3711 VDD.n4876 VDD.n4875 3.42376
R3712 VDD.n4397 VDD.n4396 3.42376
R3713 VDD.n4335 VDD.n4334 3.42376
R3714 VDD.n3862 VDD.n3861 3.42376
R3715 VDD.n5024 VDD.n5023 3.42376
R3716 VDD.n5925 VDD.n5924 3.42376
R3717 VDD.n593 VDD.n590 3.41853
R3718 VDD.n1223 VDD.n1220 3.41853
R3719 VDD.n6090 VDD.n612 3.41388
R3720 VDD.n5926 VDD.n5925 3.41326
R3721 VDD.n7076 VDD.n7075 3.41326
R3722 VDD.n3863 VDD.n3862 3.41326
R3723 VDD.n4398 VDD.n4397 3.41326
R3724 VDD.n5023 VDD.n5020 3.41257
R3725 VDD.n6182 VDD.n6181 3.41257
R3726 VDD.n4336 VDD.n4335 3.41257
R3727 VDD.n4877 VDD.n4876 3.41257
R3728 VDD.n2479 VDD.n2461 3.41219
R3729 VDD.n4961 VDD.n4937 3.41219
R3730 VDD.n6105 VDD.n6104 3.41218
R3731 VDD.n6110 VDD.n6109 3.41218
R3732 VDD.n6104 VDD.n621 3.41218
R3733 VDD.n6110 VDD.n616 3.41218
R3734 VDD.n628 VDD.n620 3.41218
R3735 VDD.n6101 VDD.n615 3.41218
R3736 VDD.n6179 VDD.n6178 3.41218
R3737 VDD.n6150 VDD.n574 3.41218
R3738 VDD.n6149 VDD.n570 3.41218
R3739 VDD.n6139 VDD.n577 3.41218
R3740 VDD.n6165 VDD.n580 3.41218
R3741 VDD.n6140 VDD.n6139 3.41218
R3742 VDD.n6142 VDD.n580 3.41218
R3743 VDD.n583 VDD.n574 3.41218
R3744 VDD.n582 VDD.n570 3.41218
R3745 VDD.n6169 VDD.n6168 3.41218
R3746 VDD.n6174 VDD.n6173 3.41218
R3747 VDD.n5008 VDD.n5007 3.41218
R3748 VDD.n5013 VDD.n5012 3.41218
R3749 VDD.n5018 VDD.n5017 3.41218
R3750 VDD.n4993 VDD.n1204 3.41218
R3751 VDD.n4992 VDD.n1200 3.41218
R3752 VDD.n4982 VDD.n1207 3.41218
R3753 VDD.n5004 VDD.n1210 3.41218
R3754 VDD.n4983 VDD.n4982 3.41218
R3755 VDD.n4985 VDD.n1210 3.41218
R3756 VDD.n1213 VDD.n1204 3.41218
R3757 VDD.n1212 VDD.n1200 3.41218
R3758 VDD.n3832 VDD.n3829 3.41218
R3759 VDD.n3828 VDD.n3801 3.41218
R3760 VDD.n3800 VDD.n3797 3.41218
R3761 VDD.n3796 VDD.n3793 3.41218
R3762 VDD.n3792 VDD.n3789 3.41218
R3763 VDD.n3788 VDD.n3785 3.41218
R3764 VDD.n2581 VDD.n2576 3.41218
R3765 VDD.n2575 VDD.n2570 3.41218
R3766 VDD.n2591 VDD.n2590 3.41218
R3767 VDD.n2544 VDD.n2531 3.41218
R3768 VDD.n2508 VDD.n2505 3.41218
R3769 VDD.n2504 VDD.n2498 3.41218
R3770 VDD.n2497 VDD.n2492 3.41218
R3771 VDD.n2558 VDD.n2557 3.41218
R3772 VDD.n2552 VDD.n2529 3.41218
R3773 VDD.n592 VDD.n589 3.41162
R3774 VDD.n3834 VDD.n3833 3.41162
R3775 VDD.n3836 VDD.n3833 3.41162
R3776 VDD.n2510 VDD.n2509 3.41162
R3777 VDD.n2512 VDD.n2509 3.41162
R3778 VDD.n1222 VDD.n1219 3.41162
R3779 VDD.n5931 VDD.n5930 3.4105
R3780 VDD.n5932 VDD.n665 3.4105
R3781 VDD.n6062 VDD.n6061 3.4105
R3782 VDD.n5953 VDD.n5951 3.4105
R3783 VDD.n5952 VDD.n5950 3.4105
R3784 VDD.n5990 VDD.n5989 3.4105
R3785 VDD.n5978 VDD.n5956 3.4105
R3786 VDD.n6019 VDD.n5995 3.4105
R3787 VDD.n6037 VDD.n6036 3.4105
R3788 VDD.n6000 VDD.n5999 3.4105
R3789 VDD.n6029 VDD.n6028 3.4105
R3790 VDD.n5945 VDD.n658 3.4105
R3791 VDD.n6003 VDD.n636 3.4105
R3792 VDD.n6111 VDD.n614 3.4105
R3793 VDD.n6115 VDD.n6114 3.4105
R3794 VDD.n6113 VDD.n601 3.4105
R3795 VDD.n633 VDD.n613 3.4105
R3796 VDD.n6202 VDD.n6201 3.4105
R3797 VDD.n6210 VDD.n6209 3.4105
R3798 VDD.n6295 VDD.n6294 3.4105
R3799 VDD.n6314 VDD.n483 3.4105
R3800 VDD.n6319 VDD.n474 3.4105
R3801 VDD.n6353 VDD.n463 3.4105
R3802 VDD.n6374 VDD.n6373 3.4105
R3803 VDD.n6398 VDD.n6397 3.4105
R3804 VDD.n6408 VDD.n6407 3.4105
R3805 VDD.n6521 VDD.n6520 3.4105
R3806 VDD.n6540 VDD.n349 3.4105
R3807 VDD.n6545 VDD.n340 3.4105
R3808 VDD.n6579 VDD.n329 3.4105
R3809 VDD.n6600 VDD.n6599 3.4105
R3810 VDD.n6624 VDD.n6623 3.4105
R3811 VDD.n6634 VDD.n6633 3.4105
R3812 VDD.n6747 VDD.n6746 3.4105
R3813 VDD.n6766 VDD.n215 3.4105
R3814 VDD.n6771 VDD.n206 3.4105
R3815 VDD.n6805 VDD.n195 3.4105
R3816 VDD.n6826 VDD.n6825 3.4105
R3817 VDD.n6850 VDD.n6849 3.4105
R3818 VDD.n6860 VDD.n6859 3.4105
R3819 VDD.n6973 VDD.n6972 3.4105
R3820 VDD.n6992 VDD.n81 3.4105
R3821 VDD.n6997 VDD.n72 3.4105
R3822 VDD.n7031 VDD.n61 3.4105
R3823 VDD.n7052 VDD.n7051 3.4105
R3824 VDD.n7056 VDD.n43 3.4105
R3825 VDD.n7063 VDD.n7062 3.4105
R3826 VDD.n7038 VDD.n7037 3.4105
R3827 VDD.n73 VDD.n69 3.4105
R3828 VDD.n83 VDD.n79 3.4105
R3829 VDD.n6990 VDD.n6989 3.4105
R3830 VDD.n6946 VDD.n6945 3.4105
R3831 VDD.n6933 VDD.n6932 3.4105
R3832 VDD.n6926 VDD.n6925 3.4105
R3833 VDD.n6911 VDD.n6910 3.4105
R3834 VDD.n6904 VDD.n141 3.4105
R3835 VDD.n6899 VDD.n147 3.4105
R3836 VDD.n6888 VDD.n6887 3.4105
R3837 VDD.n6880 VDD.n6879 3.4105
R3838 VDD.n6953 VDD.n6952 3.4105
R3839 VDD.n6965 VDD.n6964 3.4105
R3840 VDD.n6867 VDD.n6866 3.4105
R3841 VDD.n6857 VDD.n6856 3.4105
R3842 VDD.n6833 VDD.n6832 3.4105
R3843 VDD.n6812 VDD.n6811 3.4105
R3844 VDD.n207 VDD.n203 3.4105
R3845 VDD.n217 VDD.n213 3.4105
R3846 VDD.n6764 VDD.n6763 3.4105
R3847 VDD.n6720 VDD.n6719 3.4105
R3848 VDD.n6707 VDD.n6706 3.4105
R3849 VDD.n6700 VDD.n6699 3.4105
R3850 VDD.n6685 VDD.n6684 3.4105
R3851 VDD.n6678 VDD.n275 3.4105
R3852 VDD.n6673 VDD.n281 3.4105
R3853 VDD.n6662 VDD.n6661 3.4105
R3854 VDD.n6654 VDD.n6653 3.4105
R3855 VDD.n6727 VDD.n6726 3.4105
R3856 VDD.n6739 VDD.n6738 3.4105
R3857 VDD.n6641 VDD.n6640 3.4105
R3858 VDD.n6631 VDD.n6630 3.4105
R3859 VDD.n6607 VDD.n6606 3.4105
R3860 VDD.n6586 VDD.n6585 3.4105
R3861 VDD.n341 VDD.n337 3.4105
R3862 VDD.n351 VDD.n347 3.4105
R3863 VDD.n6538 VDD.n6537 3.4105
R3864 VDD.n6494 VDD.n6493 3.4105
R3865 VDD.n6481 VDD.n6480 3.4105
R3866 VDD.n6474 VDD.n6473 3.4105
R3867 VDD.n6459 VDD.n6458 3.4105
R3868 VDD.n6452 VDD.n409 3.4105
R3869 VDD.n6447 VDD.n415 3.4105
R3870 VDD.n6436 VDD.n6435 3.4105
R3871 VDD.n6428 VDD.n6427 3.4105
R3872 VDD.n6501 VDD.n6500 3.4105
R3873 VDD.n6513 VDD.n6512 3.4105
R3874 VDD.n6415 VDD.n6414 3.4105
R3875 VDD.n6405 VDD.n6404 3.4105
R3876 VDD.n6381 VDD.n6380 3.4105
R3877 VDD.n6360 VDD.n6359 3.4105
R3878 VDD.n475 VDD.n471 3.4105
R3879 VDD.n485 VDD.n481 3.4105
R3880 VDD.n6312 VDD.n6311 3.4105
R3881 VDD.n6268 VDD.n6267 3.4105
R3882 VDD.n6255 VDD.n6254 3.4105
R3883 VDD.n6248 VDD.n6247 3.4105
R3884 VDD.n6233 VDD.n6232 3.4105
R3885 VDD.n6226 VDD.n543 3.4105
R3886 VDD.n6221 VDD.n549 3.4105
R3887 VDD.n6275 VDD.n6274 3.4105
R3888 VDD.n6287 VDD.n6286 3.4105
R3889 VDD.n6189 VDD.n6188 3.4105
R3890 VDD.n7153 VDD.n7 3.4105
R3891 VDD.n7150 VDD.n7149 3.4105
R3892 VDD.n7081 VDD.n7080 3.4105
R3893 VDD.n7082 VDD.n36 3.4105
R3894 VDD.n7169 VDD.n7145 3.4105
R3895 VDD.n7187 VDD.n7186 3.4105
R3896 VDD.n7140 VDD.n7139 3.4105
R3897 VDD.n7128 VDD.n7106 3.4105
R3898 VDD.n7103 VDD.n7101 3.4105
R3899 VDD.n7102 VDD.n7100 3.4105
R3900 VDD.n7212 VDD.n7211 3.4105
R3901 VDD.n7095 VDD.n29 3.4105
R3902 VDD.n7179 VDD.n7178 3.4105
R3903 VDD.n7156 VDD.n7155 3.4105
R3904 VDD.n7180 VDD.n7144 3.4105
R3905 VDD.n7143 VDD.n7125 3.4105
R3906 VDD.n7183 VDD.n7126 3.4105
R3907 VDD.n7182 VDD.n7181 3.4105
R3908 VDD.n7142 VDD.n7141 3.4105
R3909 VDD.n7132 VDD.n7131 3.4105
R3910 VDD.n7135 VDD.n7127 3.4105
R3911 VDD.n7208 VDD.n34 3.4105
R3912 VDD.n7205 VDD.n7099 3.4105
R3913 VDD.n7130 VDD.n7129 3.4105
R3914 VDD.n7210 VDD.n7209 3.4105
R3915 VDD.n7094 VDD.n35 3.4105
R3916 VDD.n7098 VDD.n33 3.4105
R3917 VDD.n7154 VDD.n7152 3.4105
R3918 VDD.n7091 VDD.n7090 3.4105
R3919 VDD.n7093 VDD.n7092 3.4105
R3920 VDD.n7158 VDD.n7157 3.4105
R3921 VDD.n6184 VDD.n6183 3.4105
R3922 VDD.n6187 VDD.n6186 3.4105
R3923 VDD.n6208 VDD.n6207 3.4105
R3924 VDD.n7059 VDD.n50 3.4105
R3925 VDD.n40 VDD.n39 3.4105
R3926 VDD.n7061 VDD.n7060 3.4105
R3927 VDD.n52 VDD.n51 3.4105
R3928 VDD.n7055 VDD.n49 3.4105
R3929 VDD.n7036 VDD.n7035 3.4105
R3930 VDD.n7030 VDD.n68 3.4105
R3931 VDD.n7034 VDD.n67 3.4105
R3932 VDD.n7029 VDD.n7028 3.4105
R3933 VDD.n6998 VDD.n6996 3.4105
R3934 VDD.n7027 VDD.n7026 3.4105
R3935 VDD.n7000 VDD.n6999 3.4105
R3936 VDD.n6994 VDD.n6993 3.4105
R3937 VDD.n7002 VDD.n7001 3.4105
R3938 VDD.n6991 VDD.n84 3.4105
R3939 VDD.n6968 VDD.n98 3.4105
R3940 VDD.n6969 VDD.n85 3.4105
R3941 VDD.n6886 VDD.n6885 3.4105
R3942 VDD.n159 VDD.n158 3.4105
R3943 VDD.n6882 VDD.n6881 3.4105
R3944 VDD.n6906 VDD.n6905 3.4105
R3945 VDD.n6884 VDD.n157 3.4105
R3946 VDD.n6902 VDD.n148 3.4105
R3947 VDD.n6928 VDD.n6927 3.4105
R3948 VDD.n6907 VDD.n145 3.4105
R3949 VDD.n6909 VDD.n6908 3.4105
R3950 VDD.n6948 VDD.n6947 3.4105
R3951 VDD.n6929 VDD.n131 3.4105
R3952 VDD.n6931 VDD.n6930 3.4105
R3953 VDD.n6967 VDD.n6966 3.4105
R3954 VDD.n6949 VDD.n120 3.4105
R3955 VDD.n6951 VDD.n6950 3.4105
R3956 VDD.n6865 VDD.n6864 3.4105
R3957 VDD.n169 VDD.n168 3.4105
R3958 VDD.n6862 VDD.n6861 3.4105
R3959 VDD.n6855 VDD.n6854 3.4105
R3960 VDD.n173 VDD.n172 3.4105
R3961 VDD.n6853 VDD.n171 3.4105
R3962 VDD.n6831 VDD.n6830 3.4105
R3963 VDD.n186 VDD.n185 3.4105
R3964 VDD.n6829 VDD.n184 3.4105
R3965 VDD.n6810 VDD.n6809 3.4105
R3966 VDD.n6804 VDD.n202 3.4105
R3967 VDD.n6808 VDD.n201 3.4105
R3968 VDD.n6803 VDD.n6802 3.4105
R3969 VDD.n6772 VDD.n6770 3.4105
R3970 VDD.n6801 VDD.n6800 3.4105
R3971 VDD.n6774 VDD.n6773 3.4105
R3972 VDD.n6768 VDD.n6767 3.4105
R3973 VDD.n6776 VDD.n6775 3.4105
R3974 VDD.n6765 VDD.n218 3.4105
R3975 VDD.n6742 VDD.n232 3.4105
R3976 VDD.n6743 VDD.n219 3.4105
R3977 VDD.n6660 VDD.n6659 3.4105
R3978 VDD.n293 VDD.n292 3.4105
R3979 VDD.n6656 VDD.n6655 3.4105
R3980 VDD.n6680 VDD.n6679 3.4105
R3981 VDD.n6658 VDD.n291 3.4105
R3982 VDD.n6676 VDD.n282 3.4105
R3983 VDD.n6702 VDD.n6701 3.4105
R3984 VDD.n6681 VDD.n279 3.4105
R3985 VDD.n6683 VDD.n6682 3.4105
R3986 VDD.n6722 VDD.n6721 3.4105
R3987 VDD.n6703 VDD.n265 3.4105
R3988 VDD.n6705 VDD.n6704 3.4105
R3989 VDD.n6741 VDD.n6740 3.4105
R3990 VDD.n6723 VDD.n254 3.4105
R3991 VDD.n6725 VDD.n6724 3.4105
R3992 VDD.n6639 VDD.n6638 3.4105
R3993 VDD.n303 VDD.n302 3.4105
R3994 VDD.n6636 VDD.n6635 3.4105
R3995 VDD.n6629 VDD.n6628 3.4105
R3996 VDD.n307 VDD.n306 3.4105
R3997 VDD.n6627 VDD.n305 3.4105
R3998 VDD.n6605 VDD.n6604 3.4105
R3999 VDD.n320 VDD.n319 3.4105
R4000 VDD.n6603 VDD.n318 3.4105
R4001 VDD.n6584 VDD.n6583 3.4105
R4002 VDD.n6578 VDD.n336 3.4105
R4003 VDD.n6582 VDD.n335 3.4105
R4004 VDD.n6577 VDD.n6576 3.4105
R4005 VDD.n6546 VDD.n6544 3.4105
R4006 VDD.n6575 VDD.n6574 3.4105
R4007 VDD.n6548 VDD.n6547 3.4105
R4008 VDD.n6542 VDD.n6541 3.4105
R4009 VDD.n6550 VDD.n6549 3.4105
R4010 VDD.n6539 VDD.n352 3.4105
R4011 VDD.n6516 VDD.n366 3.4105
R4012 VDD.n6517 VDD.n353 3.4105
R4013 VDD.n6434 VDD.n6433 3.4105
R4014 VDD.n427 VDD.n426 3.4105
R4015 VDD.n6430 VDD.n6429 3.4105
R4016 VDD.n6454 VDD.n6453 3.4105
R4017 VDD.n6432 VDD.n425 3.4105
R4018 VDD.n6450 VDD.n416 3.4105
R4019 VDD.n6476 VDD.n6475 3.4105
R4020 VDD.n6455 VDD.n413 3.4105
R4021 VDD.n6457 VDD.n6456 3.4105
R4022 VDD.n6496 VDD.n6495 3.4105
R4023 VDD.n6477 VDD.n399 3.4105
R4024 VDD.n6479 VDD.n6478 3.4105
R4025 VDD.n6515 VDD.n6514 3.4105
R4026 VDD.n6497 VDD.n388 3.4105
R4027 VDD.n6499 VDD.n6498 3.4105
R4028 VDD.n6413 VDD.n6412 3.4105
R4029 VDD.n437 VDD.n436 3.4105
R4030 VDD.n6410 VDD.n6409 3.4105
R4031 VDD.n6403 VDD.n6402 3.4105
R4032 VDD.n441 VDD.n440 3.4105
R4033 VDD.n6401 VDD.n439 3.4105
R4034 VDD.n6379 VDD.n6378 3.4105
R4035 VDD.n454 VDD.n453 3.4105
R4036 VDD.n6377 VDD.n452 3.4105
R4037 VDD.n6358 VDD.n6357 3.4105
R4038 VDD.n6352 VDD.n470 3.4105
R4039 VDD.n6356 VDD.n469 3.4105
R4040 VDD.n6351 VDD.n6350 3.4105
R4041 VDD.n6320 VDD.n6318 3.4105
R4042 VDD.n6349 VDD.n6348 3.4105
R4043 VDD.n6322 VDD.n6321 3.4105
R4044 VDD.n6316 VDD.n6315 3.4105
R4045 VDD.n6324 VDD.n6323 3.4105
R4046 VDD.n6313 VDD.n486 3.4105
R4047 VDD.n6290 VDD.n500 3.4105
R4048 VDD.n6291 VDD.n487 3.4105
R4049 VDD.n6228 VDD.n6227 3.4105
R4050 VDD.n6206 VDD.n559 3.4105
R4051 VDD.n6224 VDD.n550 3.4105
R4052 VDD.n6250 VDD.n6249 3.4105
R4053 VDD.n6229 VDD.n547 3.4105
R4054 VDD.n6231 VDD.n6230 3.4105
R4055 VDD.n6270 VDD.n6269 3.4105
R4056 VDD.n6251 VDD.n533 3.4105
R4057 VDD.n6253 VDD.n6252 3.4105
R4058 VDD.n6289 VDD.n6288 3.4105
R4059 VDD.n6271 VDD.n522 3.4105
R4060 VDD.n6273 VDD.n6272 3.4105
R4061 VDD.n6204 VDD.n6203 3.4105
R4062 VDD.n561 VDD.n560 3.4105
R4063 VDD.n593 VDD.n592 3.4105
R4064 VDD.n598 VDD.n597 3.4105
R4065 VDD.n6136 VDD.n6135 3.4105
R4066 VDD.n6117 VDD.n599 3.4105
R4067 VDD.n6085 VDD.n6084 3.4105
R4068 VDD.n6004 VDD.n6002 3.4105
R4069 VDD.n6008 VDD.n6007 3.4105
R4070 VDD.n5993 VDD.n5975 3.4105
R4071 VDD.n6033 VDD.n5976 3.4105
R4072 VDD.n6032 VDD.n6031 3.4105
R4073 VDD.n6030 VDD.n5994 3.4105
R4074 VDD.n5992 VDD.n5991 3.4105
R4075 VDD.n5982 VDD.n5981 3.4105
R4076 VDD.n5985 VDD.n5977 3.4105
R4077 VDD.n6058 VDD.n663 3.4105
R4078 VDD.n6055 VDD.n5949 3.4105
R4079 VDD.n5980 VDD.n5979 3.4105
R4080 VDD.n6060 VDD.n6059 3.4105
R4081 VDD.n5944 VDD.n664 3.4105
R4082 VDD.n5948 VDD.n662 3.4105
R4083 VDD.n5941 VDD.n5940 3.4105
R4084 VDD.n5943 VDD.n5942 3.4105
R4085 VDD.n6006 VDD.n6005 3.4105
R4086 VDD.n3837 VDD.n3834 3.4105
R4087 VDD.n3837 VDD.n3836 3.4105
R4088 VDD.n3859 VDD.n3858 3.4105
R4089 VDD.n3860 VDD.n3859 3.4105
R4090 VDD.n3856 VDD.n3855 3.4105
R4091 VDD.n3857 VDD.n3856 3.4105
R4092 VDD.n3853 VDD.n3852 3.4105
R4093 VDD.n3854 VDD.n3853 3.4105
R4094 VDD.n3850 VDD.n3849 3.4105
R4095 VDD.n3851 VDD.n3850 3.4105
R4096 VDD.n3847 VDD.n3846 3.4105
R4097 VDD.n3848 VDD.n3847 3.4105
R4098 VDD.n3844 VDD.n3843 3.4105
R4099 VDD.n3845 VDD.n3844 3.4105
R4100 VDD.n4388 VDD.n4387 3.4105
R4101 VDD.n2732 VDD.n2731 3.4105
R4102 VDD.n2633 VDD.n2438 3.4105
R4103 VDD.n4380 VDD.n4379 3.4105
R4104 VDD.n2660 VDD.n2443 3.4105
R4105 VDD.n2670 VDD.n2669 3.4105
R4106 VDD.n2676 VDD.n2647 3.4105
R4107 VDD.n2652 VDD.n2649 3.4105
R4108 VDD.n2681 VDD.n2651 3.4105
R4109 VDD.n4353 VDD.n4352 3.4105
R4110 VDD.n2718 VDD.n2686 3.4105
R4111 VDD.n4339 VDD.n4338 3.4105
R4112 VDD.n4390 VDD.n4389 3.4105
R4113 VDD.n1412 VDD.n1377 3.4105
R4114 VDD.n2357 VDD.n2344 3.4105
R4115 VDD.n4447 VDD.n4446 3.4105
R4116 VDD.n2381 VDD.n2380 3.4105
R4117 VDD.n4439 VDD.n4438 3.4105
R4118 VDD.n2399 VDD.n2386 3.4105
R4119 VDD.n4425 VDD.n4424 3.4105
R4120 VDD.n2423 VDD.n2422 3.4105
R4121 VDD.n4417 VDD.n4416 3.4105
R4122 VDD.n4403 VDD.n4402 3.4105
R4123 VDD.n2339 VDD.n2338 3.4105
R4124 VDD.n4461 VDD.n4460 3.4105
R4125 VDD.n2214 VDD.n2213 3.4105
R4126 VDD.n2220 VDD.n2196 3.4105
R4127 VDD.n2201 VDD.n2198 3.4105
R4128 VDD.n2225 VDD.n2200 3.4105
R4129 VDD.n4488 VDD.n4487 3.4105
R4130 VDD.n2273 VDD.n2230 3.4105
R4131 VDD.n2283 VDD.n2282 3.4105
R4132 VDD.n2289 VDD.n2260 3.4105
R4133 VDD.n2265 VDD.n2262 3.4105
R4134 VDD.n2294 VDD.n2264 3.4105
R4135 VDD.n2170 VDD.n2164 3.4105
R4136 VDD.n4512 VDD.n2169 3.4105
R4137 VDD.n2093 VDD.n2080 3.4105
R4138 VDD.n4568 VDD.n4567 3.4105
R4139 VDD.n2117 VDD.n2116 3.4105
R4140 VDD.n4560 VDD.n4559 3.4105
R4141 VDD.n2135 VDD.n2122 3.4105
R4142 VDD.n4546 VDD.n4545 3.4105
R4143 VDD.n2159 VDD.n2158 3.4105
R4144 VDD.n4538 VDD.n4537 3.4105
R4145 VDD.n2171 VDD.n2163 3.4105
R4146 VDD.n4524 VDD.n4523 3.4105
R4147 VDD.n2075 VDD.n2074 3.4105
R4148 VDD.n4582 VDD.n4581 3.4105
R4149 VDD.n1950 VDD.n1949 3.4105
R4150 VDD.n1956 VDD.n1932 3.4105
R4151 VDD.n1937 VDD.n1934 3.4105
R4152 VDD.n1961 VDD.n1936 3.4105
R4153 VDD.n4609 VDD.n4608 3.4105
R4154 VDD.n2009 VDD.n1966 3.4105
R4155 VDD.n2019 VDD.n2018 3.4105
R4156 VDD.n2025 VDD.n1996 3.4105
R4157 VDD.n2001 VDD.n1998 3.4105
R4158 VDD.n2030 VDD.n2000 3.4105
R4159 VDD.n1906 VDD.n1900 3.4105
R4160 VDD.n4633 VDD.n1905 3.4105
R4161 VDD.n1829 VDD.n1816 3.4105
R4162 VDD.n4689 VDD.n4688 3.4105
R4163 VDD.n1853 VDD.n1852 3.4105
R4164 VDD.n4681 VDD.n4680 3.4105
R4165 VDD.n1871 VDD.n1858 3.4105
R4166 VDD.n4667 VDD.n4666 3.4105
R4167 VDD.n1895 VDD.n1894 3.4105
R4168 VDD.n4659 VDD.n4658 3.4105
R4169 VDD.n1907 VDD.n1899 3.4105
R4170 VDD.n4645 VDD.n4644 3.4105
R4171 VDD.n1811 VDD.n1810 3.4105
R4172 VDD.n4703 VDD.n4702 3.4105
R4173 VDD.n1686 VDD.n1685 3.4105
R4174 VDD.n1692 VDD.n1668 3.4105
R4175 VDD.n1673 VDD.n1670 3.4105
R4176 VDD.n1697 VDD.n1672 3.4105
R4177 VDD.n4730 VDD.n4729 3.4105
R4178 VDD.n1745 VDD.n1702 3.4105
R4179 VDD.n1755 VDD.n1754 3.4105
R4180 VDD.n1761 VDD.n1732 3.4105
R4181 VDD.n1737 VDD.n1734 3.4105
R4182 VDD.n1766 VDD.n1736 3.4105
R4183 VDD.n1642 VDD.n1636 3.4105
R4184 VDD.n4754 VDD.n1641 3.4105
R4185 VDD.n1565 VDD.n1552 3.4105
R4186 VDD.n4810 VDD.n4809 3.4105
R4187 VDD.n1589 VDD.n1588 3.4105
R4188 VDD.n4802 VDD.n4801 3.4105
R4189 VDD.n1607 VDD.n1594 3.4105
R4190 VDD.n4788 VDD.n4787 3.4105
R4191 VDD.n1631 VDD.n1630 3.4105
R4192 VDD.n4780 VDD.n4779 3.4105
R4193 VDD.n1643 VDD.n1635 3.4105
R4194 VDD.n4766 VDD.n4765 3.4105
R4195 VDD.n1547 VDD.n1546 3.4105
R4196 VDD.n4824 VDD.n4823 3.4105
R4197 VDD.n1405 VDD.n1402 3.4105
R4198 VDD.n1433 VDD.n1404 3.4105
R4199 VDD.n4851 VDD.n4850 3.4105
R4200 VDD.n1481 VDD.n1438 3.4105
R4201 VDD.n1491 VDD.n1490 3.4105
R4202 VDD.n1497 VDD.n1468 3.4105
R4203 VDD.n1473 VDD.n1470 3.4105
R4204 VDD.n1502 VDD.n1472 3.4105
R4205 VDD.n1428 VDD.n1400 3.4105
R4206 VDD.n1422 VDD.n1421 3.4105
R4207 VDD.n1278 VDD.n1277 3.4105
R4208 VDD.n1346 VDD.n1343 3.4105
R4209 VDD.n1285 VDD.n1284 3.4105
R4210 VDD.n1295 VDD.n1294 3.4105
R4211 VDD.n1301 VDD.n1252 3.4105
R4212 VDD.n1257 VDD.n1254 3.4105
R4213 VDD.n1306 VDD.n1256 3.4105
R4214 VDD.n4903 VDD.n4902 3.4105
R4215 VDD.n1354 VDD.n1311 3.4105
R4216 VDD.n1364 VDD.n1363 3.4105
R4217 VDD.n1370 VDD.n1341 3.4105
R4218 VDD.n4878 VDD.n1345 3.4105
R4219 VDD.n1268 VDD.n1266 3.4105
R4220 VDD.n1373 VDD.n1372 3.4105
R4221 VDD.n4882 VDD.n4881 3.4105
R4222 VDD.n1371 VDD.n1348 3.4105
R4223 VDD.n1366 VDD.n1365 3.4105
R4224 VDD.n1367 VDD.n1349 3.4105
R4225 VDD.n1355 VDD.n1350 3.4105
R4226 VDD.n4904 VDD.n1305 3.4105
R4227 VDD.n1351 VDD.n1307 3.4105
R4228 VDD.n4906 VDD.n4905 3.4105
R4229 VDD.n1304 VDD.n1303 3.4105
R4230 VDD.n4909 VDD.n4908 3.4105
R4231 VDD.n1302 VDD.n1259 3.4105
R4232 VDD.n1297 VDD.n1296 3.4105
R4233 VDD.n1298 VDD.n1260 3.4105
R4234 VDD.n1262 VDD.n1261 3.4105
R4235 VDD.n1280 VDD.n1279 3.4105
R4236 VDD.n1281 VDD.n1264 3.4105
R4237 VDD.n1269 VDD.n1265 3.4105
R4238 VDD.n2426 VDD.n2416 3.4105
R4239 VDD.n4399 VDD.n2417 3.4105
R4240 VDD.n2425 VDD.n2424 3.4105
R4241 VDD.n4418 VDD.n2385 3.4105
R4242 VDD.n2420 VDD.n2419 3.4105
R4243 VDD.n2384 VDD.n2374 3.4105
R4244 VDD.n4421 VDD.n2375 3.4105
R4245 VDD.n4420 VDD.n4419 3.4105
R4246 VDD.n2383 VDD.n2382 3.4105
R4247 VDD.n4440 VDD.n2343 3.4105
R4248 VDD.n2378 VDD.n2377 3.4105
R4249 VDD.n2342 VDD.n2332 3.4105
R4250 VDD.n4443 VDD.n2333 3.4105
R4251 VDD.n4442 VDD.n4441 3.4105
R4252 VDD.n2341 VDD.n2340 3.4105
R4253 VDD.n4462 VDD.n2293 3.4105
R4254 VDD.n2336 VDD.n2335 3.4105
R4255 VDD.n2292 VDD.n2291 3.4105
R4256 VDD.n4467 VDD.n4466 3.4105
R4257 VDD.n4464 VDD.n4463 3.4105
R4258 VDD.n2290 VDD.n2267 3.4105
R4259 VDD.n2285 VDD.n2284 3.4105
R4260 VDD.n2286 VDD.n2268 3.4105
R4261 VDD.n4489 VDD.n2224 3.4105
R4262 VDD.n2270 VDD.n2226 3.4105
R4263 VDD.n2274 VDD.n2269 3.4105
R4264 VDD.n4491 VDD.n4490 3.4105
R4265 VDD.n2223 VDD.n2222 3.4105
R4266 VDD.n4494 VDD.n4493 3.4105
R4267 VDD.n2216 VDD.n2215 3.4105
R4268 VDD.n2217 VDD.n2204 3.4105
R4269 VDD.n2221 VDD.n2203 3.4105
R4270 VDD.n2206 VDD.n2205 3.4105
R4271 VDD.n4517 VDD.n4516 3.4105
R4272 VDD.n4515 VDD.n4514 3.4105
R4273 VDD.n2162 VDD.n2152 3.4105
R4274 VDD.n4520 VDD.n2153 3.4105
R4275 VDD.n4519 VDD.n4518 3.4105
R4276 VDD.n2161 VDD.n2160 3.4105
R4277 VDD.n4539 VDD.n2121 3.4105
R4278 VDD.n2156 VDD.n2155 3.4105
R4279 VDD.n2120 VDD.n2110 3.4105
R4280 VDD.n4542 VDD.n2111 3.4105
R4281 VDD.n4541 VDD.n4540 3.4105
R4282 VDD.n2119 VDD.n2118 3.4105
R4283 VDD.n4561 VDD.n2079 3.4105
R4284 VDD.n2114 VDD.n2113 3.4105
R4285 VDD.n2078 VDD.n2068 3.4105
R4286 VDD.n4564 VDD.n2069 3.4105
R4287 VDD.n4563 VDD.n4562 3.4105
R4288 VDD.n2077 VDD.n2076 3.4105
R4289 VDD.n4583 VDD.n2029 3.4105
R4290 VDD.n2072 VDD.n2071 3.4105
R4291 VDD.n2028 VDD.n2027 3.4105
R4292 VDD.n4588 VDD.n4587 3.4105
R4293 VDD.n4585 VDD.n4584 3.4105
R4294 VDD.n2026 VDD.n2003 3.4105
R4295 VDD.n2021 VDD.n2020 3.4105
R4296 VDD.n2022 VDD.n2004 3.4105
R4297 VDD.n4610 VDD.n1960 3.4105
R4298 VDD.n2006 VDD.n1962 3.4105
R4299 VDD.n2010 VDD.n2005 3.4105
R4300 VDD.n4612 VDD.n4611 3.4105
R4301 VDD.n1959 VDD.n1958 3.4105
R4302 VDD.n4615 VDD.n4614 3.4105
R4303 VDD.n1952 VDD.n1951 3.4105
R4304 VDD.n1953 VDD.n1940 3.4105
R4305 VDD.n1957 VDD.n1939 3.4105
R4306 VDD.n1942 VDD.n1941 3.4105
R4307 VDD.n4638 VDD.n4637 3.4105
R4308 VDD.n4636 VDD.n4635 3.4105
R4309 VDD.n1898 VDD.n1888 3.4105
R4310 VDD.n4641 VDD.n1889 3.4105
R4311 VDD.n4640 VDD.n4639 3.4105
R4312 VDD.n1897 VDD.n1896 3.4105
R4313 VDD.n4660 VDD.n1857 3.4105
R4314 VDD.n1892 VDD.n1891 3.4105
R4315 VDD.n1856 VDD.n1846 3.4105
R4316 VDD.n4663 VDD.n1847 3.4105
R4317 VDD.n4662 VDD.n4661 3.4105
R4318 VDD.n1855 VDD.n1854 3.4105
R4319 VDD.n4682 VDD.n1815 3.4105
R4320 VDD.n1850 VDD.n1849 3.4105
R4321 VDD.n1814 VDD.n1804 3.4105
R4322 VDD.n4685 VDD.n1805 3.4105
R4323 VDD.n4684 VDD.n4683 3.4105
R4324 VDD.n1813 VDD.n1812 3.4105
R4325 VDD.n4704 VDD.n1765 3.4105
R4326 VDD.n1808 VDD.n1807 3.4105
R4327 VDD.n1764 VDD.n1763 3.4105
R4328 VDD.n4709 VDD.n4708 3.4105
R4329 VDD.n4706 VDD.n4705 3.4105
R4330 VDD.n1762 VDD.n1739 3.4105
R4331 VDD.n1757 VDD.n1756 3.4105
R4332 VDD.n1758 VDD.n1740 3.4105
R4333 VDD.n4731 VDD.n1696 3.4105
R4334 VDD.n1742 VDD.n1698 3.4105
R4335 VDD.n1746 VDD.n1741 3.4105
R4336 VDD.n4733 VDD.n4732 3.4105
R4337 VDD.n1695 VDD.n1694 3.4105
R4338 VDD.n4736 VDD.n4735 3.4105
R4339 VDD.n1688 VDD.n1687 3.4105
R4340 VDD.n1689 VDD.n1676 3.4105
R4341 VDD.n1693 VDD.n1675 3.4105
R4342 VDD.n1678 VDD.n1677 3.4105
R4343 VDD.n4759 VDD.n4758 3.4105
R4344 VDD.n4757 VDD.n4756 3.4105
R4345 VDD.n1634 VDD.n1624 3.4105
R4346 VDD.n4762 VDD.n1625 3.4105
R4347 VDD.n4761 VDD.n4760 3.4105
R4348 VDD.n1633 VDD.n1632 3.4105
R4349 VDD.n4781 VDD.n1593 3.4105
R4350 VDD.n1628 VDD.n1627 3.4105
R4351 VDD.n1592 VDD.n1582 3.4105
R4352 VDD.n4784 VDD.n1583 3.4105
R4353 VDD.n4783 VDD.n4782 3.4105
R4354 VDD.n1591 VDD.n1590 3.4105
R4355 VDD.n4803 VDD.n1551 3.4105
R4356 VDD.n1586 VDD.n1585 3.4105
R4357 VDD.n1550 VDD.n1540 3.4105
R4358 VDD.n4806 VDD.n1541 3.4105
R4359 VDD.n4805 VDD.n4804 3.4105
R4360 VDD.n1549 VDD.n1548 3.4105
R4361 VDD.n4825 VDD.n1501 3.4105
R4362 VDD.n1544 VDD.n1543 3.4105
R4363 VDD.n1500 VDD.n1499 3.4105
R4364 VDD.n4830 VDD.n4829 3.4105
R4365 VDD.n4827 VDD.n4826 3.4105
R4366 VDD.n1498 VDD.n1475 3.4105
R4367 VDD.n1493 VDD.n1492 3.4105
R4368 VDD.n1494 VDD.n1476 3.4105
R4369 VDD.n4852 VDD.n1432 3.4105
R4370 VDD.n1478 VDD.n1434 3.4105
R4371 VDD.n1482 VDD.n1477 3.4105
R4372 VDD.n4854 VDD.n4853 3.4105
R4373 VDD.n1431 VDD.n1430 3.4105
R4374 VDD.n4857 VDD.n4856 3.4105
R4375 VDD.n1424 VDD.n1423 3.4105
R4376 VDD.n1425 VDD.n1408 3.4105
R4377 VDD.n1429 VDD.n1407 3.4105
R4378 VDD.n1413 VDD.n1409 3.4105
R4379 VDD.n1375 VDD.n1374 3.4105
R4380 VDD.n2513 VDD.n2510 3.4105
R4381 VDD.n2513 VDD.n2512 3.4105
R4382 VDD.n2554 VDD.n2553 3.4105
R4383 VDD.n2553 VDD.n2547 3.4105
R4384 VDD.n2528 VDD.n2491 3.4105
R4385 VDD.n2555 VDD.n2491 3.4105
R4386 VDD.n2526 VDD.n2525 3.4105
R4387 VDD.n2527 VDD.n2526 3.4105
R4388 VDD.n2523 VDD.n2522 3.4105
R4389 VDD.n2524 VDD.n2523 3.4105
R4390 VDD.n2520 VDD.n2519 3.4105
R4391 VDD.n2521 VDD.n2520 3.4105
R4392 VDD.n2546 VDD.n2545 3.4105
R4393 VDD.n2545 VDD.n2427 3.4105
R4394 VDD.n2467 VDD.n2462 3.4105
R4395 VDD.n2612 VDD.n2611 3.4105
R4396 VDD.n2469 VDD.n2468 3.4105
R4397 VDD.n2614 VDD.n2613 3.4105
R4398 VDD.n2587 VDD.n2569 3.4105
R4399 VDD.n2588 VDD.n2569 3.4105
R4400 VDD.n2585 VDD.n2584 3.4105
R4401 VDD.n2586 VDD.n2585 3.4105
R4402 VDD.n2582 VDD.n2465 3.4105
R4403 VDD.n2583 VDD.n2582 3.4105
R4404 VDD.n2607 VDD.n2459 3.4105
R4405 VDD.n2607 VDD.n2606 3.4105
R4406 VDD.n2609 VDD.n2608 3.4105
R4407 VDD.n2724 VDD.n2717 3.4105
R4408 VDD.n2734 VDD.n2733 3.4105
R4409 VDD.n2723 VDD.n2722 3.4105
R4410 VDD.n4354 VDD.n2680 3.4105
R4411 VDD.n2719 VDD.n2682 3.4105
R4412 VDD.n2679 VDD.n2678 3.4105
R4413 VDD.n4359 VDD.n4358 3.4105
R4414 VDD.n4356 VDD.n4355 3.4105
R4415 VDD.n2677 VDD.n2654 3.4105
R4416 VDD.n2672 VDD.n2671 3.4105
R4417 VDD.n2673 VDD.n2655 3.4105
R4418 VDD.n4381 VDD.n2437 3.4105
R4419 VDD.n2657 VDD.n2439 3.4105
R4420 VDD.n2661 VDD.n2656 3.4105
R4421 VDD.n4383 VDD.n4382 3.4105
R4422 VDD.n2436 VDD.n2432 3.4105
R4423 VDD.n4386 VDD.n4385 3.4105
R4424 VDD.n2435 VDD.n2430 3.4105
R4425 VDD.n3784 VDD.n3774 3.4105
R4426 VDD.n3783 VDD.n3782 3.4105
R4427 VDD.n3883 VDD.n3745 3.4105
R4428 VDD.n3885 VDD.n3884 3.4105
R4429 VDD.n3743 VDD.n3742 3.4105
R4430 VDD.n3741 VDD.n3734 3.4105
R4431 VDD.n3904 VDD.n3702 3.4105
R4432 VDD.n3906 VDD.n3905 3.4105
R4433 VDD.n3700 VDD.n3699 3.4105
R4434 VDD.n3698 VDD.n3691 3.4105
R4435 VDD.n3925 VDD.n3649 3.4105
R4436 VDD.n3927 VDD.n3926 3.4105
R4437 VDD.n3648 VDD.n3647 3.4105
R4438 VDD.n3646 VDD.n3623 3.4105
R4439 VDD.n3641 VDD.n3640 3.4105
R4440 VDD.n3630 VDD.n3625 3.4105
R4441 VDD.n3952 VDD.n3580 3.4105
R4442 VDD.n3954 VDD.n3953 3.4105
R4443 VDD.n3579 VDD.n3578 3.4105
R4444 VDD.n3577 VDD.n3559 3.4105
R4445 VDD.n3572 VDD.n3571 3.4105
R4446 VDD.n3562 VDD.n3561 3.4105
R4447 VDD.n3980 VDD.n3979 3.4105
R4448 VDD.n3982 VDD.n3981 3.4105
R4449 VDD.n3518 VDD.n3508 3.4105
R4450 VDD.n3517 VDD.n3516 3.4105
R4451 VDD.n4002 VDD.n3479 3.4105
R4452 VDD.n4004 VDD.n4003 3.4105
R4453 VDD.n3477 VDD.n3476 3.4105
R4454 VDD.n3475 VDD.n3468 3.4105
R4455 VDD.n4023 VDD.n3436 3.4105
R4456 VDD.n4025 VDD.n4024 3.4105
R4457 VDD.n3434 VDD.n3433 3.4105
R4458 VDD.n3432 VDD.n3425 3.4105
R4459 VDD.n4044 VDD.n3383 3.4105
R4460 VDD.n4046 VDD.n4045 3.4105
R4461 VDD.n3382 VDD.n3381 3.4105
R4462 VDD.n3380 VDD.n3357 3.4105
R4463 VDD.n3375 VDD.n3374 3.4105
R4464 VDD.n3364 VDD.n3359 3.4105
R4465 VDD.n4071 VDD.n3314 3.4105
R4466 VDD.n4073 VDD.n4072 3.4105
R4467 VDD.n3313 VDD.n3312 3.4105
R4468 VDD.n3311 VDD.n3293 3.4105
R4469 VDD.n3306 VDD.n3305 3.4105
R4470 VDD.n3296 VDD.n3295 3.4105
R4471 VDD.n4099 VDD.n4098 3.4105
R4472 VDD.n4101 VDD.n4100 3.4105
R4473 VDD.n3252 VDD.n3242 3.4105
R4474 VDD.n3251 VDD.n3250 3.4105
R4475 VDD.n4121 VDD.n3213 3.4105
R4476 VDD.n4123 VDD.n4122 3.4105
R4477 VDD.n3211 VDD.n3210 3.4105
R4478 VDD.n3209 VDD.n3202 3.4105
R4479 VDD.n4142 VDD.n3170 3.4105
R4480 VDD.n4144 VDD.n4143 3.4105
R4481 VDD.n3168 VDD.n3167 3.4105
R4482 VDD.n3166 VDD.n3159 3.4105
R4483 VDD.n4163 VDD.n3117 3.4105
R4484 VDD.n4165 VDD.n4164 3.4105
R4485 VDD.n3116 VDD.n3115 3.4105
R4486 VDD.n3114 VDD.n3091 3.4105
R4487 VDD.n3109 VDD.n3108 3.4105
R4488 VDD.n3098 VDD.n3093 3.4105
R4489 VDD.n4190 VDD.n3048 3.4105
R4490 VDD.n4192 VDD.n4191 3.4105
R4491 VDD.n3047 VDD.n3046 3.4105
R4492 VDD.n3045 VDD.n3027 3.4105
R4493 VDD.n3040 VDD.n3039 3.4105
R4494 VDD.n3030 VDD.n3029 3.4105
R4495 VDD.n4218 VDD.n4217 3.4105
R4496 VDD.n4220 VDD.n4219 3.4105
R4497 VDD.n2986 VDD.n2976 3.4105
R4498 VDD.n2985 VDD.n2984 3.4105
R4499 VDD.n4240 VDD.n2947 3.4105
R4500 VDD.n4242 VDD.n4241 3.4105
R4501 VDD.n2945 VDD.n2944 3.4105
R4502 VDD.n2943 VDD.n2936 3.4105
R4503 VDD.n4261 VDD.n2904 3.4105
R4504 VDD.n4263 VDD.n4262 3.4105
R4505 VDD.n2902 VDD.n2901 3.4105
R4506 VDD.n2900 VDD.n2861 3.4105
R4507 VDD.n2889 VDD.n2864 3.4105
R4508 VDD.n2888 VDD.n2887 3.4105
R4509 VDD.n2874 VDD.n2873 3.4105
R4510 VDD.n2872 VDD.n2867 3.4105
R4511 VDD.n4301 VDD.n2806 3.4105
R4512 VDD.n4303 VDD.n4302 3.4105
R4513 VDD.n2805 VDD.n2804 3.4105
R4514 VDD.n2803 VDD.n2785 3.4105
R4515 VDD.n2798 VDD.n2797 3.4105
R4516 VDD.n2788 VDD.n2787 3.4105
R4517 VDD.n4328 VDD.n2743 3.4105
R4518 VDD.n4330 VDD.n4329 3.4105
R4519 VDD.n3864 VDD.n3775 3.4105
R4520 VDD.n3778 VDD.n3777 3.4105
R4521 VDD.n3887 VDD.n3886 3.4105
R4522 VDD.n3737 VDD.n3736 3.4105
R4523 VDD.n3908 VDD.n3907 3.4105
R4524 VDD.n3694 VDD.n3693 3.4105
R4525 VDD.n3930 VDD.n3929 3.4105
R4526 VDD.n3642 VDD.n3624 3.4105
R4527 VDD.n3626 VDD.n3582 3.4105
R4528 VDD.n3957 VDD.n3956 3.4105
R4529 VDD.n3573 VDD.n3560 3.4105
R4530 VDD.n3978 VDD.n3977 3.4105
R4531 VDD.n3983 VDD.n3509 3.4105
R4532 VDD.n3512 VDD.n3511 3.4105
R4533 VDD.n4006 VDD.n4005 3.4105
R4534 VDD.n3471 VDD.n3470 3.4105
R4535 VDD.n4027 VDD.n4026 3.4105
R4536 VDD.n3428 VDD.n3427 3.4105
R4537 VDD.n4049 VDD.n4048 3.4105
R4538 VDD.n3376 VDD.n3358 3.4105
R4539 VDD.n3360 VDD.n3316 3.4105
R4540 VDD.n4076 VDD.n4075 3.4105
R4541 VDD.n3307 VDD.n3294 3.4105
R4542 VDD.n4097 VDD.n4096 3.4105
R4543 VDD.n4102 VDD.n3243 3.4105
R4544 VDD.n3246 VDD.n3245 3.4105
R4545 VDD.n4125 VDD.n4124 3.4105
R4546 VDD.n3205 VDD.n3204 3.4105
R4547 VDD.n4146 VDD.n4145 3.4105
R4548 VDD.n3162 VDD.n3161 3.4105
R4549 VDD.n4168 VDD.n4167 3.4105
R4550 VDD.n3110 VDD.n3092 3.4105
R4551 VDD.n3094 VDD.n3050 3.4105
R4552 VDD.n4195 VDD.n4194 3.4105
R4553 VDD.n3041 VDD.n3028 3.4105
R4554 VDD.n4216 VDD.n4215 3.4105
R4555 VDD.n4221 VDD.n2977 3.4105
R4556 VDD.n2980 VDD.n2979 3.4105
R4557 VDD.n4244 VDD.n4243 3.4105
R4558 VDD.n2939 VDD.n2938 3.4105
R4559 VDD.n4265 VDD.n4264 3.4105
R4560 VDD.n2890 VDD.n2862 3.4105
R4561 VDD.n2884 VDD.n2875 3.4105
R4562 VDD.n2868 VDD.n2808 3.4105
R4563 VDD.n4306 VDD.n4305 3.4105
R4564 VDD.n2799 VDD.n2786 3.4105
R4565 VDD.n4327 VDD.n4326 3.4105
R4566 VDD.n4332 VDD.n4331 3.4105
R4567 VDD.n3714 VDD.n3690 3.4105
R4568 VDD.n3910 VDD.n3687 3.4105
R4569 VDD.n3740 VDD.n3739 3.4105
R4570 VDD.n3903 VDD.n3902 3.4105
R4571 VDD.n3757 VDD.n3733 3.4105
R4572 VDD.n3889 VDD.n3730 3.4105
R4573 VDD.n3781 VDD.n3780 3.4105
R4574 VDD.n3882 VDD.n3881 3.4105
R4575 VDD.n3868 VDD.n3867 3.4105
R4576 VDD.n3697 VDD.n3696 3.4105
R4577 VDD.n3924 VDD.n3923 3.4105
R4578 VDD.n3570 VDD.n3569 3.4105
R4579 VDD.n3576 VDD.n3552 3.4105
R4580 VDD.n3557 VDD.n3554 3.4105
R4581 VDD.n3581 VDD.n3556 3.4105
R4582 VDD.n3951 VDD.n3950 3.4105
R4583 VDD.n3629 VDD.n3586 3.4105
R4584 VDD.n3639 VDD.n3638 3.4105
R4585 VDD.n3645 VDD.n3616 3.4105
R4586 VDD.n3621 VDD.n3618 3.4105
R4587 VDD.n3650 VDD.n3620 3.4105
R4588 VDD.n3526 VDD.n3520 3.4105
R4589 VDD.n3975 VDD.n3524 3.4105
R4590 VDD.n3448 VDD.n3424 3.4105
R4591 VDD.n4029 VDD.n3421 3.4105
R4592 VDD.n3474 VDD.n3473 3.4105
R4593 VDD.n4022 VDD.n4021 3.4105
R4594 VDD.n3491 VDD.n3467 3.4105
R4595 VDD.n4008 VDD.n3464 3.4105
R4596 VDD.n3515 VDD.n3514 3.4105
R4597 VDD.n4001 VDD.n4000 3.4105
R4598 VDD.n3527 VDD.n3519 3.4105
R4599 VDD.n3987 VDD.n3986 3.4105
R4600 VDD.n3431 VDD.n3430 3.4105
R4601 VDD.n4043 VDD.n4042 3.4105
R4602 VDD.n3304 VDD.n3303 3.4105
R4603 VDD.n3310 VDD.n3286 3.4105
R4604 VDD.n3291 VDD.n3288 3.4105
R4605 VDD.n3315 VDD.n3290 3.4105
R4606 VDD.n4070 VDD.n4069 3.4105
R4607 VDD.n3363 VDD.n3320 3.4105
R4608 VDD.n3373 VDD.n3372 3.4105
R4609 VDD.n3379 VDD.n3350 3.4105
R4610 VDD.n3355 VDD.n3352 3.4105
R4611 VDD.n3384 VDD.n3354 3.4105
R4612 VDD.n3260 VDD.n3254 3.4105
R4613 VDD.n4094 VDD.n3258 3.4105
R4614 VDD.n3182 VDD.n3158 3.4105
R4615 VDD.n4148 VDD.n3155 3.4105
R4616 VDD.n3208 VDD.n3207 3.4105
R4617 VDD.n4141 VDD.n4140 3.4105
R4618 VDD.n3225 VDD.n3201 3.4105
R4619 VDD.n4127 VDD.n3198 3.4105
R4620 VDD.n3249 VDD.n3248 3.4105
R4621 VDD.n4120 VDD.n4119 3.4105
R4622 VDD.n3261 VDD.n3253 3.4105
R4623 VDD.n4106 VDD.n4105 3.4105
R4624 VDD.n3165 VDD.n3164 3.4105
R4625 VDD.n4162 VDD.n4161 3.4105
R4626 VDD.n3038 VDD.n3037 3.4105
R4627 VDD.n3044 VDD.n3020 3.4105
R4628 VDD.n3025 VDD.n3022 3.4105
R4629 VDD.n3049 VDD.n3024 3.4105
R4630 VDD.n4189 VDD.n4188 3.4105
R4631 VDD.n3097 VDD.n3054 3.4105
R4632 VDD.n3107 VDD.n3106 3.4105
R4633 VDD.n3113 VDD.n3084 3.4105
R4634 VDD.n3089 VDD.n3086 3.4105
R4635 VDD.n3118 VDD.n3088 3.4105
R4636 VDD.n2994 VDD.n2988 3.4105
R4637 VDD.n4213 VDD.n2992 3.4105
R4638 VDD.n2916 VDD.n2860 3.4105
R4639 VDD.n4267 VDD.n2857 3.4105
R4640 VDD.n2942 VDD.n2941 3.4105
R4641 VDD.n4260 VDD.n4259 3.4105
R4642 VDD.n2959 VDD.n2935 3.4105
R4643 VDD.n4246 VDD.n2932 3.4105
R4644 VDD.n2983 VDD.n2982 3.4105
R4645 VDD.n4239 VDD.n4238 3.4105
R4646 VDD.n2995 VDD.n2987 3.4105
R4647 VDD.n4225 VDD.n4224 3.4105
R4648 VDD.n2899 VDD.n2898 3.4105
R4649 VDD.n2894 VDD.n2893 3.4105
R4650 VDD.n2796 VDD.n2795 3.4105
R4651 VDD.n2802 VDD.n2778 3.4105
R4652 VDD.n2783 VDD.n2780 3.4105
R4653 VDD.n2807 VDD.n2782 3.4105
R4654 VDD.n4300 VDD.n4299 3.4105
R4655 VDD.n2871 VDD.n2812 3.4105
R4656 VDD.n2881 VDD.n2866 3.4105
R4657 VDD.n2886 VDD.n2842 3.4105
R4658 VDD.n4324 VDD.n2750 3.4105
R4659 VDD.n2764 VDD.n2746 3.4105
R4660 VDD.n2737 VDD.n2736 3.4105
R4661 VDD.n4942 VDD.n4941 3.4105
R4662 VDD.n4948 VDD.n4947 3.4105
R4663 VDD.n4940 VDD.n1233 3.4105
R4664 VDD.n4950 VDD.n4949 3.4105
R4665 VDD.n4978 VDD.n1231 3.4105
R4666 VDD.n4978 VDD.n4977 3.4105
R4667 VDD.n4945 VDD.n1230 3.4105
R4668 VDD.n1223 VDD.n1222 3.4105
R4669 VDD.n1228 VDD.n1227 3.4105
R4670 VDD.n5908 VDD.n686 3.4105
R4671 VDD.n5910 VDD.n5909 3.4105
R4672 VDD.n5900 VDD.n687 3.4105
R4673 VDD.n5899 VDD.n5898 3.4105
R4674 VDD.n5868 VDD.n5866 3.4105
R4675 VDD.n5870 VDD.n5869 3.4105
R4676 VDD.n5864 VDD.n5863 3.4105
R4677 VDD.n5861 VDD.n703 3.4105
R4678 VDD.n5838 VDD.n719 3.4105
R4679 VDD.n5837 VDD.n5836 3.4105
R4680 VDD.n5817 VDD.n727 3.4105
R4681 VDD.n5816 VDD.n5815 3.4105
R4682 VDD.n5797 VDD.n749 3.4105
R4683 VDD.n5796 VDD.n5795 3.4105
R4684 VDD.n5774 VDD.n763 3.4105
R4685 VDD.n5773 VDD.n5772 3.4105
R4686 VDD.n5740 VDD.n5738 3.4105
R4687 VDD.n5742 VDD.n5741 3.4105
R4688 VDD.n5736 VDD.n777 3.4105
R4689 VDD.n5735 VDD.n5734 3.4105
R4690 VDD.n5715 VDD.n789 3.4105
R4691 VDD.n5714 VDD.n5713 3.4105
R4692 VDD.n5691 VDD.n803 3.4105
R4693 VDD.n5693 VDD.n5692 3.4105
R4694 VDD.n5683 VDD.n804 3.4105
R4695 VDD.n5682 VDD.n5681 3.4105
R4696 VDD.n5653 VDD.n819 3.4105
R4697 VDD.n5655 VDD.n5654 3.4105
R4698 VDD.n821 VDD.n820 3.4105
R4699 VDD.n5633 VDD.n5632 3.4105
R4700 VDD.n5627 VDD.n838 3.4105
R4701 VDD.n5626 VDD.n5625 3.4105
R4702 VDD.n5595 VDD.n5593 3.4105
R4703 VDD.n5597 VDD.n5596 3.4105
R4704 VDD.n5591 VDD.n5590 3.4105
R4705 VDD.n5588 VDD.n854 3.4105
R4706 VDD.n5569 VDD.n884 3.4105
R4707 VDD.n5568 VDD.n5567 3.4105
R4708 VDD.n5546 VDD.n898 3.4105
R4709 VDD.n5545 VDD.n5544 3.4105
R4710 VDD.n5512 VDD.n5510 3.4105
R4711 VDD.n5514 VDD.n5513 3.4105
R4712 VDD.n5508 VDD.n912 3.4105
R4713 VDD.n5507 VDD.n5506 3.4105
R4714 VDD.n5487 VDD.n924 3.4105
R4715 VDD.n5486 VDD.n5485 3.4105
R4716 VDD.n5463 VDD.n938 3.4105
R4717 VDD.n5465 VDD.n5464 3.4105
R4718 VDD.n5455 VDD.n939 3.4105
R4719 VDD.n5454 VDD.n5453 3.4105
R4720 VDD.n5425 VDD.n954 3.4105
R4721 VDD.n5427 VDD.n5426 3.4105
R4722 VDD.n956 VDD.n955 3.4105
R4723 VDD.n5405 VDD.n5404 3.4105
R4724 VDD.n5399 VDD.n973 3.4105
R4725 VDD.n5398 VDD.n5397 3.4105
R4726 VDD.n5367 VDD.n5365 3.4105
R4727 VDD.n5369 VDD.n5368 3.4105
R4728 VDD.n5363 VDD.n5362 3.4105
R4729 VDD.n5360 VDD.n989 3.4105
R4730 VDD.n5341 VDD.n1019 3.4105
R4731 VDD.n5340 VDD.n5339 3.4105
R4732 VDD.n5318 VDD.n1033 3.4105
R4733 VDD.n5317 VDD.n5316 3.4105
R4734 VDD.n5284 VDD.n5282 3.4105
R4735 VDD.n5286 VDD.n5285 3.4105
R4736 VDD.n5280 VDD.n1047 3.4105
R4737 VDD.n5279 VDD.n5278 3.4105
R4738 VDD.n5259 VDD.n1059 3.4105
R4739 VDD.n5258 VDD.n5257 3.4105
R4740 VDD.n5235 VDD.n1073 3.4105
R4741 VDD.n5237 VDD.n5236 3.4105
R4742 VDD.n5227 VDD.n1074 3.4105
R4743 VDD.n5226 VDD.n5225 3.4105
R4744 VDD.n5197 VDD.n1089 3.4105
R4745 VDD.n5199 VDD.n5198 3.4105
R4746 VDD.n1091 VDD.n1090 3.4105
R4747 VDD.n5177 VDD.n5176 3.4105
R4748 VDD.n5171 VDD.n1108 3.4105
R4749 VDD.n5170 VDD.n5169 3.4105
R4750 VDD.n5139 VDD.n5137 3.4105
R4751 VDD.n5141 VDD.n5140 3.4105
R4752 VDD.n5135 VDD.n5134 3.4105
R4753 VDD.n5132 VDD.n1124 3.4105
R4754 VDD.n5113 VDD.n1154 3.4105
R4755 VDD.n5112 VDD.n5111 3.4105
R4756 VDD.n5090 VDD.n1168 3.4105
R4757 VDD.n5089 VDD.n5088 3.4105
R4758 VDD.n5056 VDD.n5054 3.4105
R4759 VDD.n5058 VDD.n5057 3.4105
R4760 VDD.n5052 VDD.n1182 3.4105
R4761 VDD.n5051 VDD.n5050 3.4105
R4762 VDD.n5031 VDD.n1194 3.4105
R4763 VDD.n5030 VDD.n5029 3.4105
R4764 VDD.n669 VDD.n668 3.4105
R4765 VDD.n5904 VDD.n685 3.4105
R4766 VDD.n5897 VDD.n5896 3.4105
R4767 VDD.n5872 VDD.n5871 3.4105
R4768 VDD.n5839 VDD.n704 3.4105
R4769 VDD.n721 VDD.n720 3.4105
R4770 VDD.n5799 VDD.n5798 3.4105
R4771 VDD.n5776 VDD.n5775 3.4105
R4772 VDD.n5769 VDD.n766 3.4105
R4773 VDD.n5747 VDD.n5737 3.4105
R4774 VDD.n5717 VDD.n5716 3.4105
R4775 VDD.n5690 VDD.n5689 3.4105
R4776 VDD.n5687 VDD.n802 3.4105
R4777 VDD.n5680 VDD.n5679 3.4105
R4778 VDD.n5652 VDD.n817 3.4105
R4779 VDD.n5631 VDD.n837 3.4105
R4780 VDD.n5624 VDD.n5623 3.4105
R4781 VDD.n5599 VDD.n5598 3.4105
R4782 VDD.n5572 VDD.n5571 3.4105
R4783 VDD.n5548 VDD.n5547 3.4105
R4784 VDD.n5541 VDD.n901 3.4105
R4785 VDD.n5519 VDD.n5509 3.4105
R4786 VDD.n5489 VDD.n5488 3.4105
R4787 VDD.n5462 VDD.n5461 3.4105
R4788 VDD.n5459 VDD.n937 3.4105
R4789 VDD.n5452 VDD.n5451 3.4105
R4790 VDD.n5424 VDD.n952 3.4105
R4791 VDD.n5403 VDD.n972 3.4105
R4792 VDD.n5396 VDD.n5395 3.4105
R4793 VDD.n5371 VDD.n5370 3.4105
R4794 VDD.n5344 VDD.n5343 3.4105
R4795 VDD.n5320 VDD.n5319 3.4105
R4796 VDD.n5313 VDD.n1036 3.4105
R4797 VDD.n5291 VDD.n5281 3.4105
R4798 VDD.n5261 VDD.n5260 3.4105
R4799 VDD.n5234 VDD.n5233 3.4105
R4800 VDD.n5231 VDD.n1072 3.4105
R4801 VDD.n5224 VDD.n5223 3.4105
R4802 VDD.n5196 VDD.n1087 3.4105
R4803 VDD.n5175 VDD.n1107 3.4105
R4804 VDD.n5168 VDD.n5167 3.4105
R4805 VDD.n5143 VDD.n5142 3.4105
R4806 VDD.n5116 VDD.n5115 3.4105
R4807 VDD.n5092 VDD.n5091 3.4105
R4808 VDD.n5085 VDD.n1171 3.4105
R4809 VDD.n5063 VDD.n5053 3.4105
R4810 VDD.n5033 VDD.n5032 3.4105
R4811 VDD.n5028 VDD.n5027 3.4105
R4812 VDD.n5860 VDD.n5859 3.4105
R4813 VDD.n5844 VDD.n5842 3.4105
R4814 VDD.n702 VDD.n698 3.4105
R4815 VDD.n5862 VDD.n700 3.4105
R4816 VDD.n692 VDD.n688 3.4105
R4817 VDD.n5867 VDD.n691 3.4105
R4818 VDD.n5912 VDD.n5911 3.4105
R4819 VDD.n5901 VDD.n678 3.4105
R4820 VDD.n5905 VDD.n672 3.4105
R4821 VDD.n5835 VDD.n5834 3.4105
R4822 VDD.n5822 VDD.n5820 3.4105
R4823 VDD.n5719 VDD.n5718 3.4105
R4824 VDD.n5733 VDD.n5732 3.4105
R4825 VDD.n5749 VDD.n5748 3.4105
R4826 VDD.n5745 VDD.n5743 3.4105
R4827 VDD.n5766 VDD.n765 3.4105
R4828 VDD.n5771 VDD.n759 3.4105
R4829 VDD.n5778 VDD.n5777 3.4105
R4830 VDD.n5794 VDD.n5793 3.4105
R4831 VDD.n5801 VDD.n5800 3.4105
R4832 VDD.n5814 VDD.n5813 3.4105
R4833 VDD.n5688 VDD.n801 3.4105
R4834 VDD.n5712 VDD.n5711 3.4105
R4835 VDD.n843 VDD.n839 3.4105
R4836 VDD.n5594 VDD.n842 3.4105
R4837 VDD.n5635 VDD.n5634 3.4105
R4838 VDD.n5628 VDD.n831 3.4105
R4839 VDD.n5657 VDD.n5656 3.4105
R4840 VDD.n5649 VDD.n5648 3.4105
R4841 VDD.n809 VDD.n805 3.4105
R4842 VDD.n818 VDD.n808 3.4105
R4843 VDD.n5695 VDD.n5694 3.4105
R4844 VDD.n5684 VDD.n798 3.4105
R4845 VDD.n853 VDD.n849 3.4105
R4846 VDD.n5589 VDD.n851 3.4105
R4847 VDD.n5491 VDD.n5490 3.4105
R4848 VDD.n5505 VDD.n5504 3.4105
R4849 VDD.n5521 VDD.n5520 3.4105
R4850 VDD.n5517 VDD.n5515 3.4105
R4851 VDD.n5538 VDD.n900 3.4105
R4852 VDD.n5543 VDD.n894 3.4105
R4853 VDD.n5550 VDD.n5549 3.4105
R4854 VDD.n5566 VDD.n5565 3.4105
R4855 VDD.n5574 VDD.n5573 3.4105
R4856 VDD.n5587 VDD.n5586 3.4105
R4857 VDD.n5460 VDD.n936 3.4105
R4858 VDD.n5484 VDD.n5483 3.4105
R4859 VDD.n978 VDD.n974 3.4105
R4860 VDD.n5366 VDD.n977 3.4105
R4861 VDD.n5407 VDD.n5406 3.4105
R4862 VDD.n5400 VDD.n966 3.4105
R4863 VDD.n5429 VDD.n5428 3.4105
R4864 VDD.n5421 VDD.n5420 3.4105
R4865 VDD.n944 VDD.n940 3.4105
R4866 VDD.n953 VDD.n943 3.4105
R4867 VDD.n5467 VDD.n5466 3.4105
R4868 VDD.n5456 VDD.n933 3.4105
R4869 VDD.n988 VDD.n984 3.4105
R4870 VDD.n5361 VDD.n986 3.4105
R4871 VDD.n5263 VDD.n5262 3.4105
R4872 VDD.n5277 VDD.n5276 3.4105
R4873 VDD.n5293 VDD.n5292 3.4105
R4874 VDD.n5289 VDD.n5287 3.4105
R4875 VDD.n5310 VDD.n1035 3.4105
R4876 VDD.n5315 VDD.n1029 3.4105
R4877 VDD.n5322 VDD.n5321 3.4105
R4878 VDD.n5338 VDD.n5337 3.4105
R4879 VDD.n5346 VDD.n5345 3.4105
R4880 VDD.n5359 VDD.n5358 3.4105
R4881 VDD.n5232 VDD.n1071 3.4105
R4882 VDD.n5256 VDD.n5255 3.4105
R4883 VDD.n1113 VDD.n1109 3.4105
R4884 VDD.n5138 VDD.n1112 3.4105
R4885 VDD.n5179 VDD.n5178 3.4105
R4886 VDD.n5172 VDD.n1101 3.4105
R4887 VDD.n5201 VDD.n5200 3.4105
R4888 VDD.n5193 VDD.n5192 3.4105
R4889 VDD.n1079 VDD.n1075 3.4105
R4890 VDD.n1088 VDD.n1078 3.4105
R4891 VDD.n5239 VDD.n5238 3.4105
R4892 VDD.n5228 VDD.n1068 3.4105
R4893 VDD.n1123 VDD.n1119 3.4105
R4894 VDD.n5133 VDD.n1121 3.4105
R4895 VDD.n5065 VDD.n5064 3.4105
R4896 VDD.n5061 VDD.n5059 3.4105
R4897 VDD.n5082 VDD.n1170 3.4105
R4898 VDD.n5087 VDD.n1164 3.4105
R4899 VDD.n5094 VDD.n5093 3.4105
R4900 VDD.n5110 VDD.n5109 3.4105
R4901 VDD.n5118 VDD.n5117 3.4105
R4902 VDD.n5131 VDD.n5130 3.4105
R4903 VDD.n5049 VDD.n5048 3.4105
R4904 VDD.n5035 VDD.n5034 3.4105
R4905 VDD.n5022 VDD.n5021 3.4105
R4906 VDD.n6982 VDD.n6979 3.38568
R4907 VDD.n7015 VDD.n58 3.38568
R4908 VDD.n6756 VDD.n6753 3.38568
R4909 VDD.n6789 VDD.n192 3.38568
R4910 VDD.n6846 VDD.n6840 3.38568
R4911 VDD.n6530 VDD.n6527 3.38568
R4912 VDD.n6563 VDD.n326 3.38568
R4913 VDD.n6620 VDD.n6614 3.38568
R4914 VDD.n6304 VDD.n6301 3.38568
R4915 VDD.n6337 VDD.n460 3.38568
R4916 VDD.n6394 VDD.n6388 3.38568
R4917 VDD.n5729 VDD.n5728 3.38568
R4918 VDD.n5786 VDD.n5785 3.38568
R4919 VDD.n5501 VDD.n5500 3.38568
R4920 VDD.n5558 VDD.n5557 3.38568
R4921 VDD.n5273 VDD.n5272 3.38568
R4922 VDD.n5330 VDD.n5329 3.38568
R4923 VDD.n5045 VDD.n5044 3.38568
R4924 VDD.n5102 VDD.n5101 3.38568
R4925 VDD.n5885 VDD.n675 3.38568
R4926 VDD.n5852 VDD.n5851 3.38568
R4927 VDD.n5666 VDD.n5665 3.38568
R4928 VDD.n5612 VDD.n828 3.38568
R4929 VDD.n5438 VDD.n5437 3.38568
R4930 VDD.n5384 VDD.n963 3.38568
R4931 VDD.n5210 VDD.n5209 3.38568
R4932 VDD.n5156 VDD.n1098 3.38568
R4933 VDD.n6025 VDD.n646 3.38568
R4934 VDD.n7175 VDD.n17 3.38568
R4935 VDD.n6942 VDD.n115 3.38568
R4936 VDD.n6716 VDD.n249 3.38568
R4937 VDD.n6490 VDD.n383 3.38568
R4938 VDD.n6264 VDD.n517 3.38568
R4939 VDD.n6070 VDD.n6069 3.10353
R4940 VDD.n654 VDD.n653 3.10353
R4941 VDD.n5958 VDD.n656 3.10353
R4942 VDD.n5963 VDD.n5959 3.10353
R4943 VDD.n5968 VDD.n5967 3.10353
R4944 VDD.n6047 VDD.n5969 3.10353
R4945 VDD.n6044 VDD.n6042 3.10353
R4946 VDD.n6041 VDD.n5970 3.10353
R4947 VDD.n6016 VDD.n6013 3.10353
R4948 VDD.n6024 VDD.n6023 3.10353
R4949 VDD.n6196 VDD.n564 3.10353
R4950 VDD.n6195 VDD.n555 3.10353
R4951 VDD.n6217 VDD.n553 3.10353
R4952 VDD.n6216 VDD.n540 3.10353
R4953 VDD.n544 VDD.n541 3.10353
R4954 VDD.n6244 VDD.n538 3.10353
R4955 VDD.n6259 VDD.n529 3.10353
R4956 VDD.n6260 VDD.n527 3.10353
R4957 VDD.n6279 VDD.n518 3.10353
R4958 VDD.n6280 VDD.n507 3.10353
R4959 VDD.n516 VDD.n515 3.10353
R4960 VDD.n508 VDD.n496 3.10353
R4961 VDD.n495 VDD.n492 3.10353
R4962 VDD.n6307 VDD.n6306 3.10353
R4963 VDD.n494 VDD.n493 3.10353
R4964 VDD.n6332 VDD.n479 3.10353
R4965 VDD.n6339 VDD.n477 3.10353
R4966 VDD.n6340 VDD.n461 3.10353
R4967 VDD.n6365 VDD.n459 3.10353
R4968 VDD.n464 VDD.n458 3.10353
R4969 VDD.n6386 VDD.n449 3.10353
R4970 VDD.n6385 VDD.n446 3.10353
R4971 VDD.n6391 VDD.n447 3.10353
R4972 VDD.n6390 VDD.n432 3.10353
R4973 VDD.n6422 VDD.n430 3.10353
R4974 VDD.n6421 VDD.n421 3.10353
R4975 VDD.n6443 VDD.n419 3.10353
R4976 VDD.n6442 VDD.n406 3.10353
R4977 VDD.n410 VDD.n407 3.10353
R4978 VDD.n6470 VDD.n404 3.10353
R4979 VDD.n6485 VDD.n395 3.10353
R4980 VDD.n6486 VDD.n393 3.10353
R4981 VDD.n6505 VDD.n384 3.10353
R4982 VDD.n6506 VDD.n373 3.10353
R4983 VDD.n382 VDD.n381 3.10353
R4984 VDD.n374 VDD.n362 3.10353
R4985 VDD.n361 VDD.n358 3.10353
R4986 VDD.n6533 VDD.n6532 3.10353
R4987 VDD.n360 VDD.n359 3.10353
R4988 VDD.n6558 VDD.n345 3.10353
R4989 VDD.n6565 VDD.n343 3.10353
R4990 VDD.n6566 VDD.n327 3.10353
R4991 VDD.n6591 VDD.n325 3.10353
R4992 VDD.n330 VDD.n324 3.10353
R4993 VDD.n6612 VDD.n315 3.10353
R4994 VDD.n6611 VDD.n312 3.10353
R4995 VDD.n6617 VDD.n313 3.10353
R4996 VDD.n6616 VDD.n298 3.10353
R4997 VDD.n6648 VDD.n296 3.10353
R4998 VDD.n6647 VDD.n287 3.10353
R4999 VDD.n6669 VDD.n285 3.10353
R5000 VDD.n6668 VDD.n272 3.10353
R5001 VDD.n276 VDD.n273 3.10353
R5002 VDD.n6696 VDD.n270 3.10353
R5003 VDD.n6711 VDD.n261 3.10353
R5004 VDD.n6712 VDD.n259 3.10353
R5005 VDD.n6731 VDD.n250 3.10353
R5006 VDD.n6732 VDD.n239 3.10353
R5007 VDD.n248 VDD.n247 3.10353
R5008 VDD.n240 VDD.n228 3.10353
R5009 VDD.n227 VDD.n224 3.10353
R5010 VDD.n6759 VDD.n6758 3.10353
R5011 VDD.n226 VDD.n225 3.10353
R5012 VDD.n6784 VDD.n211 3.10353
R5013 VDD.n6791 VDD.n209 3.10353
R5014 VDD.n6792 VDD.n193 3.10353
R5015 VDD.n6817 VDD.n191 3.10353
R5016 VDD.n196 VDD.n190 3.10353
R5017 VDD.n6838 VDD.n181 3.10353
R5018 VDD.n6837 VDD.n178 3.10353
R5019 VDD.n6843 VDD.n179 3.10353
R5020 VDD.n6842 VDD.n164 3.10353
R5021 VDD.n6874 VDD.n162 3.10353
R5022 VDD.n6873 VDD.n153 3.10353
R5023 VDD.n6895 VDD.n151 3.10353
R5024 VDD.n6894 VDD.n138 3.10353
R5025 VDD.n142 VDD.n139 3.10353
R5026 VDD.n6922 VDD.n136 3.10353
R5027 VDD.n6937 VDD.n127 3.10353
R5028 VDD.n6938 VDD.n125 3.10353
R5029 VDD.n6957 VDD.n116 3.10353
R5030 VDD.n6958 VDD.n105 3.10353
R5031 VDD.n114 VDD.n113 3.10353
R5032 VDD.n106 VDD.n94 3.10353
R5033 VDD.n93 VDD.n90 3.10353
R5034 VDD.n6985 VDD.n6984 3.10353
R5035 VDD.n92 VDD.n91 3.10353
R5036 VDD.n7010 VDD.n77 3.10353
R5037 VDD.n7017 VDD.n75 3.10353
R5038 VDD.n7018 VDD.n59 3.10353
R5039 VDD.n7043 VDD.n57 3.10353
R5040 VDD.n62 VDD.n56 3.10353
R5041 VDD.n7069 VDD.n46 3.10353
R5042 VDD.n7068 VDD.n44 3.10353
R5043 VDD.n7220 VDD.n7219 3.10353
R5044 VDD.n25 VDD.n24 3.10353
R5045 VDD.n7108 VDD.n27 3.10353
R5046 VDD.n7113 VDD.n7109 3.10353
R5047 VDD.n7118 VDD.n7117 3.10353
R5048 VDD.n7197 VDD.n7119 3.10353
R5049 VDD.n7194 VDD.n7192 3.10353
R5050 VDD.n7191 VDD.n7120 3.10353
R5051 VDD.n7166 VDD.n7163 3.10353
R5052 VDD.n7174 VDD.n7173 3.10353
R5053 VDD.n2637 VDD.n2451 3.10353
R5054 VDD.n2638 VDD.n2445 3.10353
R5055 VDD.n2663 VDD.n2446 3.10353
R5056 VDD.n4369 VDD.n2644 3.10353
R5057 VDD.n2694 VDD.n2645 3.10353
R5058 VDD.n2700 VDD.n2695 3.10353
R5059 VDD.n2706 VDD.n2702 3.10353
R5060 VDD.n2707 VDD.n2688 3.10353
R5061 VDD.n2726 VDD.n2689 3.10353
R5062 VDD.n4342 VDD.n2713 3.10353
R5063 VDD.n1415 VDD.n1380 3.10353
R5064 VDD.n4867 VDD.n1397 3.10353
R5065 VDD.n1446 VDD.n1398 3.10353
R5066 VDD.n1452 VDD.n1447 3.10353
R5067 VDD.n1458 VDD.n1454 3.10353
R5068 VDD.n1459 VDD.n1440 3.10353
R5069 VDD.n1484 VDD.n1441 3.10353
R5070 VDD.n4840 VDD.n1465 3.10353
R5071 VDD.n1513 VDD.n1466 3.10353
R5072 VDD.n1517 VDD.n1516 3.10353
R5073 VDD.n1528 VDD.n1518 3.10353
R5074 VDD.n1521 VDD.n1508 3.10353
R5075 VDD.n4815 VDD.n1509 3.10353
R5076 VDD.n4814 VDD.n1535 3.10353
R5077 VDD.n1571 VDD.n1570 3.10353
R5078 VDD.n1569 VDD.n1558 3.10353
R5079 VDD.n4793 VDD.n1559 3.10353
R5080 VDD.n4792 VDD.n1577 3.10353
R5081 VDD.n1613 VDD.n1612 3.10353
R5082 VDD.n1611 VDD.n1600 3.10353
R5083 VDD.n4771 VDD.n1601 3.10353
R5084 VDD.n4770 VDD.n1619 3.10353
R5085 VDD.n1658 VDD.n1653 3.10353
R5086 VDD.n1659 VDD.n1648 3.10353
R5087 VDD.n1679 VDD.n1649 3.10353
R5088 VDD.n4746 VDD.n1665 3.10353
R5089 VDD.n1710 VDD.n1666 3.10353
R5090 VDD.n1716 VDD.n1711 3.10353
R5091 VDD.n1722 VDD.n1718 3.10353
R5092 VDD.n1723 VDD.n1704 3.10353
R5093 VDD.n1748 VDD.n1705 3.10353
R5094 VDD.n4719 VDD.n1729 3.10353
R5095 VDD.n1777 VDD.n1730 3.10353
R5096 VDD.n1781 VDD.n1780 3.10353
R5097 VDD.n1792 VDD.n1782 3.10353
R5098 VDD.n1785 VDD.n1772 3.10353
R5099 VDD.n4694 VDD.n1773 3.10353
R5100 VDD.n4693 VDD.n1799 3.10353
R5101 VDD.n1835 VDD.n1834 3.10353
R5102 VDD.n1833 VDD.n1822 3.10353
R5103 VDD.n4672 VDD.n1823 3.10353
R5104 VDD.n4671 VDD.n1841 3.10353
R5105 VDD.n1877 VDD.n1876 3.10353
R5106 VDD.n1875 VDD.n1864 3.10353
R5107 VDD.n4650 VDD.n1865 3.10353
R5108 VDD.n4649 VDD.n1883 3.10353
R5109 VDD.n1922 VDD.n1917 3.10353
R5110 VDD.n1923 VDD.n1912 3.10353
R5111 VDD.n1943 VDD.n1913 3.10353
R5112 VDD.n4625 VDD.n1929 3.10353
R5113 VDD.n1974 VDD.n1930 3.10353
R5114 VDD.n1980 VDD.n1975 3.10353
R5115 VDD.n1986 VDD.n1982 3.10353
R5116 VDD.n1987 VDD.n1968 3.10353
R5117 VDD.n2012 VDD.n1969 3.10353
R5118 VDD.n4598 VDD.n1993 3.10353
R5119 VDD.n2041 VDD.n1994 3.10353
R5120 VDD.n2045 VDD.n2044 3.10353
R5121 VDD.n2056 VDD.n2046 3.10353
R5122 VDD.n2049 VDD.n2036 3.10353
R5123 VDD.n4573 VDD.n2037 3.10353
R5124 VDD.n4572 VDD.n2063 3.10353
R5125 VDD.n2099 VDD.n2098 3.10353
R5126 VDD.n2097 VDD.n2086 3.10353
R5127 VDD.n4551 VDD.n2087 3.10353
R5128 VDD.n4550 VDD.n2105 3.10353
R5129 VDD.n2141 VDD.n2140 3.10353
R5130 VDD.n2139 VDD.n2128 3.10353
R5131 VDD.n4529 VDD.n2129 3.10353
R5132 VDD.n4528 VDD.n2147 3.10353
R5133 VDD.n2186 VDD.n2181 3.10353
R5134 VDD.n2187 VDD.n2176 3.10353
R5135 VDD.n2207 VDD.n2177 3.10353
R5136 VDD.n4504 VDD.n2193 3.10353
R5137 VDD.n2238 VDD.n2194 3.10353
R5138 VDD.n2244 VDD.n2239 3.10353
R5139 VDD.n2250 VDD.n2246 3.10353
R5140 VDD.n2251 VDD.n2232 3.10353
R5141 VDD.n2276 VDD.n2233 3.10353
R5142 VDD.n4477 VDD.n2257 3.10353
R5143 VDD.n2305 VDD.n2258 3.10353
R5144 VDD.n2309 VDD.n2308 3.10353
R5145 VDD.n2320 VDD.n2310 3.10353
R5146 VDD.n2313 VDD.n2300 3.10353
R5147 VDD.n4452 VDD.n2301 3.10353
R5148 VDD.n4451 VDD.n2327 3.10353
R5149 VDD.n2363 VDD.n2362 3.10353
R5150 VDD.n2361 VDD.n2350 3.10353
R5151 VDD.n4430 VDD.n2351 3.10353
R5152 VDD.n4429 VDD.n2369 3.10353
R5153 VDD.n2405 VDD.n2404 3.10353
R5154 VDD.n2403 VDD.n2392 3.10353
R5155 VDD.n4408 VDD.n2393 3.10353
R5156 VDD.n4407 VDD.n2411 3.10353
R5157 VDD.n1288 VDD.n1244 3.10353
R5158 VDD.n4919 VDD.n1249 3.10353
R5159 VDD.n1319 VDD.n1250 3.10353
R5160 VDD.n1325 VDD.n1320 3.10353
R5161 VDD.n1331 VDD.n1327 3.10353
R5162 VDD.n1332 VDD.n1313 3.10353
R5163 VDD.n1357 VDD.n1314 3.10353
R5164 VDD.n4892 VDD.n1338 3.10353
R5165 VDD.n1385 VDD.n1339 3.10353
R5166 VDD.n1389 VDD.n1388 3.10353
R5167 VDD.n2768 VDD.n2763 3.10353
R5168 VDD.n2769 VDD.n2753 3.10353
R5169 VDD.n2789 VDD.n2754 3.10353
R5170 VDD.n4316 VDD.n2775 3.10353
R5171 VDD.n2820 VDD.n2776 3.10353
R5172 VDD.n2826 VDD.n2821 3.10353
R5173 VDD.n2832 VDD.n2828 3.10353
R5174 VDD.n2833 VDD.n2814 3.10353
R5175 VDD.n2877 VDD.n2815 3.10353
R5176 VDD.n4289 VDD.n2839 3.10353
R5177 VDD.n2846 VDD.n2840 3.10353
R5178 VDD.n4280 VDD.n4279 3.10353
R5179 VDD.n4272 VDD.n2847 3.10353
R5180 VDD.n4271 VDD.n2853 3.10353
R5181 VDD.n2922 VDD.n2921 3.10353
R5182 VDD.n2920 VDD.n2910 3.10353
R5183 VDD.n4251 VDD.n2911 3.10353
R5184 VDD.n4250 VDD.n2928 3.10353
R5185 VDD.n2965 VDD.n2964 3.10353
R5186 VDD.n2963 VDD.n2953 3.10353
R5187 VDD.n4230 VDD.n2954 3.10353
R5188 VDD.n4229 VDD.n2971 3.10353
R5189 VDD.n3010 VDD.n3005 3.10353
R5190 VDD.n3011 VDD.n3000 3.10353
R5191 VDD.n3031 VDD.n3001 3.10353
R5192 VDD.n4205 VDD.n3017 3.10353
R5193 VDD.n3062 VDD.n3018 3.10353
R5194 VDD.n3068 VDD.n3063 3.10353
R5195 VDD.n3074 VDD.n3070 3.10353
R5196 VDD.n3075 VDD.n3056 3.10353
R5197 VDD.n3100 VDD.n3057 3.10353
R5198 VDD.n4178 VDD.n3081 3.10353
R5199 VDD.n3129 VDD.n3082 3.10353
R5200 VDD.n3133 VDD.n3132 3.10353
R5201 VDD.n3144 VDD.n3134 3.10353
R5202 VDD.n3137 VDD.n3124 3.10353
R5203 VDD.n4153 VDD.n3125 3.10353
R5204 VDD.n4152 VDD.n3151 3.10353
R5205 VDD.n3188 VDD.n3187 3.10353
R5206 VDD.n3186 VDD.n3176 3.10353
R5207 VDD.n4132 VDD.n3177 3.10353
R5208 VDD.n4131 VDD.n3194 3.10353
R5209 VDD.n3231 VDD.n3230 3.10353
R5210 VDD.n3229 VDD.n3219 3.10353
R5211 VDD.n4111 VDD.n3220 3.10353
R5212 VDD.n4110 VDD.n3237 3.10353
R5213 VDD.n3276 VDD.n3271 3.10353
R5214 VDD.n3277 VDD.n3266 3.10353
R5215 VDD.n3297 VDD.n3267 3.10353
R5216 VDD.n4086 VDD.n3283 3.10353
R5217 VDD.n3328 VDD.n3284 3.10353
R5218 VDD.n3334 VDD.n3329 3.10353
R5219 VDD.n3340 VDD.n3336 3.10353
R5220 VDD.n3341 VDD.n3322 3.10353
R5221 VDD.n3366 VDD.n3323 3.10353
R5222 VDD.n4059 VDD.n3347 3.10353
R5223 VDD.n3395 VDD.n3348 3.10353
R5224 VDD.n3399 VDD.n3398 3.10353
R5225 VDD.n3410 VDD.n3400 3.10353
R5226 VDD.n3403 VDD.n3390 3.10353
R5227 VDD.n4034 VDD.n3391 3.10353
R5228 VDD.n4033 VDD.n3417 3.10353
R5229 VDD.n3454 VDD.n3453 3.10353
R5230 VDD.n3452 VDD.n3442 3.10353
R5231 VDD.n4013 VDD.n3443 3.10353
R5232 VDD.n4012 VDD.n3460 3.10353
R5233 VDD.n3497 VDD.n3496 3.10353
R5234 VDD.n3495 VDD.n3485 3.10353
R5235 VDD.n3992 VDD.n3486 3.10353
R5236 VDD.n3991 VDD.n3503 3.10353
R5237 VDD.n3542 VDD.n3537 3.10353
R5238 VDD.n3543 VDD.n3532 3.10353
R5239 VDD.n3563 VDD.n3533 3.10353
R5240 VDD.n3967 VDD.n3549 3.10353
R5241 VDD.n3594 VDD.n3550 3.10353
R5242 VDD.n3600 VDD.n3595 3.10353
R5243 VDD.n3606 VDD.n3602 3.10353
R5244 VDD.n3607 VDD.n3588 3.10353
R5245 VDD.n3632 VDD.n3589 3.10353
R5246 VDD.n3940 VDD.n3613 3.10353
R5247 VDD.n3661 VDD.n3614 3.10353
R5248 VDD.n3665 VDD.n3664 3.10353
R5249 VDD.n3676 VDD.n3666 3.10353
R5250 VDD.n3669 VDD.n3656 3.10353
R5251 VDD.n3915 VDD.n3657 3.10353
R5252 VDD.n3914 VDD.n3683 3.10353
R5253 VDD.n3720 VDD.n3719 3.10353
R5254 VDD.n3718 VDD.n3708 3.10353
R5255 VDD.n3894 VDD.n3709 3.10353
R5256 VDD.n3893 VDD.n3726 3.10353
R5257 VDD.n3763 VDD.n3762 3.10353
R5258 VDD.n3761 VDD.n3751 3.10353
R5259 VDD.n3873 VDD.n3752 3.10353
R5260 VDD.n3872 VDD.n3769 3.10353
R5261 VDD.n5039 VDD.n1190 3.10353
R5262 VDD.n5040 VDD.n1188 3.10353
R5263 VDD.n5069 VDD.n1177 3.10353
R5264 VDD.n5071 VDD.n5070 3.10353
R5265 VDD.n5078 VDD.n1174 3.10353
R5266 VDD.n5077 VDD.n1161 3.10353
R5267 VDD.n1165 VDD.n1162 3.10353
R5268 VDD.n5106 VDD.n1159 3.10353
R5269 VDD.n5122 VDD.n1150 3.10353
R5270 VDD.n5123 VDD.n1130 3.10353
R5271 VDD.n1148 VDD.n1147 3.10353
R5272 VDD.n1140 VDD.n1131 3.10353
R5273 VDD.n1135 VDD.n1134 3.10353
R5274 VDD.n5151 VDD.n1117 3.10353
R5275 VDD.n5158 VDD.n1115 3.10353
R5276 VDD.n5159 VDD.n1099 3.10353
R5277 VDD.n5184 VDD.n1097 3.10353
R5278 VDD.n1102 VDD.n1096 3.10353
R5279 VDD.n5207 VDD.n1083 3.10353
R5280 VDD.n5206 VDD.n1084 3.10353
R5281 VDD.n5214 VDD.n5213 3.10353
R5282 VDD.n5215 VDD.n1066 3.10353
R5283 VDD.n5248 VDD.n1064 3.10353
R5284 VDD.n5252 VDD.n5249 3.10353
R5285 VDD.n5267 VDD.n1055 3.10353
R5286 VDD.n5268 VDD.n1053 3.10353
R5287 VDD.n5297 VDD.n1042 3.10353
R5288 VDD.n5299 VDD.n5298 3.10353
R5289 VDD.n5306 VDD.n1039 3.10353
R5290 VDD.n5305 VDD.n1026 3.10353
R5291 VDD.n1030 VDD.n1027 3.10353
R5292 VDD.n5334 VDD.n1024 3.10353
R5293 VDD.n5350 VDD.n1015 3.10353
R5294 VDD.n5351 VDD.n995 3.10353
R5295 VDD.n1013 VDD.n1012 3.10353
R5296 VDD.n1005 VDD.n996 3.10353
R5297 VDD.n1000 VDD.n999 3.10353
R5298 VDD.n5379 VDD.n982 3.10353
R5299 VDD.n5386 VDD.n980 3.10353
R5300 VDD.n5387 VDD.n964 3.10353
R5301 VDD.n5412 VDD.n962 3.10353
R5302 VDD.n967 VDD.n961 3.10353
R5303 VDD.n5435 VDD.n948 3.10353
R5304 VDD.n5434 VDD.n949 3.10353
R5305 VDD.n5442 VDD.n5441 3.10353
R5306 VDD.n5443 VDD.n931 3.10353
R5307 VDD.n5476 VDD.n929 3.10353
R5308 VDD.n5480 VDD.n5477 3.10353
R5309 VDD.n5495 VDD.n920 3.10353
R5310 VDD.n5496 VDD.n918 3.10353
R5311 VDD.n5525 VDD.n907 3.10353
R5312 VDD.n5527 VDD.n5526 3.10353
R5313 VDD.n5534 VDD.n904 3.10353
R5314 VDD.n5533 VDD.n891 3.10353
R5315 VDD.n895 VDD.n892 3.10353
R5316 VDD.n5562 VDD.n889 3.10353
R5317 VDD.n5578 VDD.n880 3.10353
R5318 VDD.n5579 VDD.n860 3.10353
R5319 VDD.n878 VDD.n877 3.10353
R5320 VDD.n870 VDD.n861 3.10353
R5321 VDD.n865 VDD.n864 3.10353
R5322 VDD.n5607 VDD.n847 3.10353
R5323 VDD.n5614 VDD.n845 3.10353
R5324 VDD.n5615 VDD.n829 3.10353
R5325 VDD.n5640 VDD.n827 3.10353
R5326 VDD.n832 VDD.n826 3.10353
R5327 VDD.n5663 VDD.n813 3.10353
R5328 VDD.n5662 VDD.n814 3.10353
R5329 VDD.n5670 VDD.n5669 3.10353
R5330 VDD.n5671 VDD.n796 3.10353
R5331 VDD.n5704 VDD.n794 3.10353
R5332 VDD.n5708 VDD.n5705 3.10353
R5333 VDD.n5723 VDD.n785 3.10353
R5334 VDD.n5724 VDD.n783 3.10353
R5335 VDD.n5753 VDD.n772 3.10353
R5336 VDD.n5755 VDD.n5754 3.10353
R5337 VDD.n5762 VDD.n769 3.10353
R5338 VDD.n5761 VDD.n756 3.10353
R5339 VDD.n760 VDD.n757 3.10353
R5340 VDD.n5790 VDD.n754 3.10353
R5341 VDD.n5805 VDD.n745 3.10353
R5342 VDD.n5806 VDD.n734 3.10353
R5343 VDD.n743 VDD.n742 3.10353
R5344 VDD.n735 VDD.n724 3.10353
R5345 VDD.n5829 VDD.n5828 3.10353
R5346 VDD.n5830 VDD.n716 3.10353
R5347 VDD.n714 VDD.n709 3.10353
R5348 VDD.n5855 VDD.n5854 3.10353
R5349 VDD.n711 VDD.n710 3.10353
R5350 VDD.n5880 VDD.n696 3.10353
R5351 VDD.n5887 VDD.n694 3.10353
R5352 VDD.n5888 VDD.n676 3.10353
R5353 VDD.n5917 VDD.n674 3.10353
R5354 VDD.n679 VDD.n673 3.10353
R5355 VDD.n608 VDD.n607 3.03311
R5356 VDD.n2481 VDD.n2474 3.03311
R5357 VDD.n4963 VDD.n4933 3.03311
R5358 VDD.n7277 VDD.n7276 3.03311
R5359 VDD.n1203 VDD 2.90898
R5360 VDD.n573 VDD 2.90898
R5361 VDD.n3823 VDD.t3 2.83209
R5362 VDD.n2540 VDD.t34 2.83209
R5363 VDD.n6123 VDD.n6122 2.64177
R5364 VDD.n2476 VDD.n2474 2.64177
R5365 VDD.n4954 VDD.n4933 2.64177
R5366 VDD.n7268 VDD.n7267 2.64177
R5367 VDD.n6071 VDD.n652 2.54483
R5368 VDD.n7221 VDD.n23 2.54336
R5369 VDD.n4341 VDD.n4340 2.54336
R5370 VDD.n1390 VDD.n1344 2.54336
R5371 VDD.n6137 VDD 2.54117
R5372 VDD.n631 VDD.n607 2.4386
R5373 VDD.n2600 VDD.n2484 2.4386
R5374 VDD.n4971 VDD.n1237 2.4386
R5375 VDD.n7276 VDD.n7266 2.4386
R5376 VDD.n6075 VDD.n639 2.28608
R5377 VDD.n7225 VDD.n10 2.28608
R5378 VDD.n2630 VDD.n2453 2.28608
R5379 VDD.n4927 VDD.n4926 2.28608
R5380 VDD.n6107 VDD.n6106 2.24869
R5381 VDD.n623 VDD.n622 2.24869
R5382 VDD.n6099 VDD.n6098 2.24869
R5383 VDD.n6154 VDD.n6148 2.24869
R5384 VDD.n6163 VDD.n6162 2.24869
R5385 VDD.n6145 VDD.n6141 2.24869
R5386 VDD.n587 VDD.n581 2.24869
R5387 VDD.n6171 VDD.n6170 2.24869
R5388 VDD.n5010 VDD.n5009 2.24869
R5389 VDD.n4997 VDD.n4991 2.24869
R5390 VDD.n5002 VDD.n5001 2.24869
R5391 VDD.n4988 VDD.n4984 2.24869
R5392 VDD.n1217 VDD.n1211 2.24869
R5393 VDD.n3827 VDD.n3826 2.24858
R5394 VDD.n3814 VDD.n3813 2.24858
R5395 VDD.n3817 VDD.n3816 2.24858
R5396 VDD.n3811 VDD.n3810 2.24858
R5397 VDD.n3807 VDD.n3806 2.24858
R5398 VDD.n2580 VDD.n2565 2.24858
R5399 VDD.n2574 VDD.n2566 2.24858
R5400 VDD.n2593 VDD.n2592 2.24858
R5401 VDD.n2543 VDD.n2542 2.24858
R5402 VDD.n2503 VDD.n2502 2.24858
R5403 VDD.n2496 VDD.n2488 2.24858
R5404 VDD.n2560 VDD.n2559 2.24858
R5405 VDD.n2551 VDD.n2550 2.24858
R5406 VDD.n6076 VDD.n6075 2.15377
R5407 VDD.n7226 VDD.n7225 2.15377
R5408 VDD.n2625 VDD.n2453 2.03414
R5409 VDD.n4927 VDD.n1241 2.03414
R5410 VDD.n1218 VDD.n638 1.99051
R5411 VDD.n588 VDD.n9 1.99051
R5412 VDD.n5927 VDD 1.98118
R5413 VDD.n5928 VDD 1.9603
R5414 VDD.n6079 VDD.n6078 1.94045
R5415 VDD.n6133 VDD.n6132 1.94045
R5416 VDD.n6088 VDD.n6087 1.94045
R5417 VDD.n7229 VDD.n7228 1.94045
R5418 VDD.n2623 VDD.n2429 1.94045
R5419 VDD.n1274 VDD.n1273 1.94045
R5420 VDD.n2604 VDD.n2603 1.94045
R5421 VDD.n2617 VDD.n2616 1.94045
R5422 VDD.n4975 VDD.n4974 1.94045
R5423 VDD.n4953 VDD.n4952 1.94045
R5424 VDD.n7257 VDD.n7256 1.94045
R5425 VDD.n7283 VDD.n7282 1.94045
R5426 VDD.n6082 VDD 1.7865
R5427 VDD.n6982 VDD.n6981 1.76521
R5428 VDD.n7044 VDD.n58 1.76521
R5429 VDD.n6870 VDD.n163 1.76521
R5430 VDD.n6891 VDD.n152 1.76521
R5431 VDD.n6918 VDD.n137 1.76521
R5432 VDD.n6921 VDD.n126 1.76521
R5433 VDD.n6942 VDD.n6941 1.76521
R5434 VDD.n6756 VDD.n6755 1.76521
R5435 VDD.n6818 VDD.n192 1.76521
R5436 VDD.n6846 VDD.n6845 1.76521
R5437 VDD.n6644 VDD.n297 1.76521
R5438 VDD.n6665 VDD.n286 1.76521
R5439 VDD.n6692 VDD.n271 1.76521
R5440 VDD.n6695 VDD.n260 1.76521
R5441 VDD.n6716 VDD.n6715 1.76521
R5442 VDD.n6530 VDD.n6529 1.76521
R5443 VDD.n6592 VDD.n326 1.76521
R5444 VDD.n6620 VDD.n6619 1.76521
R5445 VDD.n6418 VDD.n431 1.76521
R5446 VDD.n6439 VDD.n420 1.76521
R5447 VDD.n6466 VDD.n405 1.76521
R5448 VDD.n6469 VDD.n394 1.76521
R5449 VDD.n6490 VDD.n6489 1.76521
R5450 VDD.n6304 VDD.n6303 1.76521
R5451 VDD.n6366 VDD.n460 1.76521
R5452 VDD.n6394 VDD.n6393 1.76521
R5453 VDD.n6240 VDD.n539 1.76521
R5454 VDD.n6243 VDD.n528 1.76521
R5455 VDD.n6264 VDD.n6263 1.76521
R5456 VDD.n7222 VDD.n22 1.76521
R5457 VDD.n7175 VDD.n11 1.76521
R5458 VDD.n6072 VDD.n651 1.76521
R5459 VDD.n6025 VDD.n640 1.76521
R5460 VDD.n5827 VDD.n5825 1.76521
R5461 VDD.n5852 VDD.n713 1.76521
R5462 VDD.n5918 VDD.n675 1.76521
R5463 VDD.n5707 VDD.n784 1.76521
R5464 VDD.n5729 VDD.n5727 1.76521
R5465 VDD.n5785 VDD.n755 1.76521
R5466 VDD.n5810 VDD.n5809 1.76521
R5467 VDD.n868 VDD.n867 1.76521
R5468 VDD.n5641 VDD.n828 1.76521
R5469 VDD.n5668 VDD.n5666 1.76521
R5470 VDD.n5479 VDD.n919 1.76521
R5471 VDD.n5501 VDD.n5499 1.76521
R5472 VDD.n5557 VDD.n890 1.76521
R5473 VDD.n5583 VDD.n5582 1.76521
R5474 VDD.n1003 VDD.n1002 1.76521
R5475 VDD.n5413 VDD.n963 1.76521
R5476 VDD.n5440 VDD.n5438 1.76521
R5477 VDD.n5251 VDD.n1054 1.76521
R5478 VDD.n5273 VDD.n5271 1.76521
R5479 VDD.n5329 VDD.n1025 1.76521
R5480 VDD.n5355 VDD.n5354 1.76521
R5481 VDD.n1138 VDD.n1137 1.76521
R5482 VDD.n5185 VDD.n1098 1.76521
R5483 VDD.n5212 VDD.n5210 1.76521
R5484 VDD.n5045 VDD.n5043 1.76521
R5485 VDD.n5101 VDD.n1160 1.76521
R5486 VDD.n5127 VDD.n5126 1.76521
R5487 VDD.n4924 VDD.n1243 1.76521
R5488 VDD.n4920 VDD.n1248 1.76521
R5489 VDD.n1324 VDD.n1318 1.76521
R5490 VDD.n4897 VDD.n1315 1.76521
R5491 VDD.n4893 VDD.n1337 1.76521
R5492 VDD.n1391 VDD.n1384 1.76521
R5493 VDD.n4457 VDD.n2302 1.76521
R5494 VDD.n2364 VDD.n2326 1.76521
R5495 VDD.n4435 VDD.n2353 1.76521
R5496 VDD.n2406 VDD.n2368 1.76521
R5497 VDD.n4413 VDD.n2395 1.76521
R5498 VDD.n2536 VDD.n2410 1.76521
R5499 VDD.n4509 VDD.n2178 1.76521
R5500 VDD.n4505 VDD.n2192 1.76521
R5501 VDD.n2243 VDD.n2237 1.76521
R5502 VDD.n4482 VDD.n2234 1.76521
R5503 VDD.n4478 VDD.n2256 1.76521
R5504 VDD.n2322 VDD.n2304 1.76521
R5505 VDD.n4578 VDD.n2038 1.76521
R5506 VDD.n2100 VDD.n2062 1.76521
R5507 VDD.n4556 VDD.n2089 1.76521
R5508 VDD.n2142 VDD.n2104 1.76521
R5509 VDD.n4534 VDD.n2131 1.76521
R5510 VDD.n2182 VDD.n2146 1.76521
R5511 VDD.n4630 VDD.n1914 1.76521
R5512 VDD.n4626 VDD.n1928 1.76521
R5513 VDD.n1979 VDD.n1973 1.76521
R5514 VDD.n4603 VDD.n1970 1.76521
R5515 VDD.n4599 VDD.n1992 1.76521
R5516 VDD.n2058 VDD.n2040 1.76521
R5517 VDD.n4699 VDD.n1774 1.76521
R5518 VDD.n1836 VDD.n1798 1.76521
R5519 VDD.n4677 VDD.n1825 1.76521
R5520 VDD.n1878 VDD.n1840 1.76521
R5521 VDD.n4655 VDD.n1867 1.76521
R5522 VDD.n1918 VDD.n1882 1.76521
R5523 VDD.n4751 VDD.n1650 1.76521
R5524 VDD.n4747 VDD.n1664 1.76521
R5525 VDD.n1715 VDD.n1709 1.76521
R5526 VDD.n4724 VDD.n1706 1.76521
R5527 VDD.n4720 VDD.n1728 1.76521
R5528 VDD.n1794 VDD.n1776 1.76521
R5529 VDD.n4820 VDD.n1510 1.76521
R5530 VDD.n1572 VDD.n1534 1.76521
R5531 VDD.n4798 VDD.n1561 1.76521
R5532 VDD.n1614 VDD.n1576 1.76521
R5533 VDD.n4776 VDD.n1603 1.76521
R5534 VDD.n1654 VDD.n1618 1.76521
R5535 VDD.n4872 VDD.n1381 1.76521
R5536 VDD.n4868 VDD.n1396 1.76521
R5537 VDD.n1451 VDD.n1445 1.76521
R5538 VDD.n4845 VDD.n1442 1.76521
R5539 VDD.n4841 VDD.n1464 1.76521
R5540 VDD.n1530 VDD.n1512 1.76521
R5541 VDD.n2629 VDD.n2450 1.76521
R5542 VDD.n4374 VDD.n2447 1.76521
R5543 VDD.n4370 VDD.n2643 1.76521
R5544 VDD.n2699 VDD.n2693 1.76521
R5545 VDD.n4347 VDD.n2690 1.76521
R5546 VDD.n4343 VDD.n2712 1.76521
R5547 VDD.n3920 VDD.n3658 1.76521
R5548 VDD.n3721 VDD.n3682 1.76521
R5549 VDD.n3899 VDD.n3711 1.76521
R5550 VDD.n3764 VDD.n3725 1.76521
R5551 VDD.n3878 VDD.n3754 1.76521
R5552 VDD.n3819 VDD.n3768 1.76521
R5553 VDD.n3972 VDD.n3534 1.76521
R5554 VDD.n3968 VDD.n3548 1.76521
R5555 VDD.n3599 VDD.n3593 1.76521
R5556 VDD.n3945 VDD.n3590 1.76521
R5557 VDD.n3941 VDD.n3612 1.76521
R5558 VDD.n3678 VDD.n3660 1.76521
R5559 VDD.n4039 VDD.n3392 1.76521
R5560 VDD.n3455 VDD.n3416 1.76521
R5561 VDD.n4018 VDD.n3445 1.76521
R5562 VDD.n3498 VDD.n3459 1.76521
R5563 VDD.n3997 VDD.n3488 1.76521
R5564 VDD.n3538 VDD.n3502 1.76521
R5565 VDD.n4091 VDD.n3268 1.76521
R5566 VDD.n4087 VDD.n3282 1.76521
R5567 VDD.n3333 VDD.n3327 1.76521
R5568 VDD.n4064 VDD.n3324 1.76521
R5569 VDD.n4060 VDD.n3346 1.76521
R5570 VDD.n3412 VDD.n3394 1.76521
R5571 VDD.n4158 VDD.n3126 1.76521
R5572 VDD.n3189 VDD.n3150 1.76521
R5573 VDD.n4137 VDD.n3179 1.76521
R5574 VDD.n3232 VDD.n3193 1.76521
R5575 VDD.n4116 VDD.n3222 1.76521
R5576 VDD.n3272 VDD.n3236 1.76521
R5577 VDD.n4210 VDD.n3002 1.76521
R5578 VDD.n4206 VDD.n3016 1.76521
R5579 VDD.n3067 VDD.n3061 1.76521
R5580 VDD.n4183 VDD.n3058 1.76521
R5581 VDD.n4179 VDD.n3080 1.76521
R5582 VDD.n3146 VDD.n3128 1.76521
R5583 VDD.n4277 VDD.n2849 1.76521
R5584 VDD.n2923 VDD.n2852 1.76521
R5585 VDD.n4256 VDD.n2913 1.76521
R5586 VDD.n2966 VDD.n2927 1.76521
R5587 VDD.n4235 VDD.n2956 1.76521
R5588 VDD.n3006 VDD.n2970 1.76521
R5589 VDD.n2762 VDD.n2761 1.76521
R5590 VDD.n4321 VDD.n2755 1.76521
R5591 VDD.n4317 VDD.n2774 1.76521
R5592 VDD.n2825 VDD.n2819 1.76521
R5593 VDD.n4294 VDD.n2816 1.76521
R5594 VDD.n4290 VDD.n2838 1.76521
R5595 VDD.n6083 VDD 1.76349
R5596 VDD.n1203 VDD.t11 1.68435
R5597 VDD.n573 VDD.t60 1.68435
R5598 VDD.n26 VDD.n20 1.66612
R5599 VDD.n7116 VDD.n14 1.66612
R5600 VDD.n7193 VDD.n18 1.66612
R5601 VDD.n7164 VDD.n16 1.66612
R5602 VDD.n655 VDD.n649 1.66612
R5603 VDD.n5966 VDD.n643 1.66612
R5604 VDD.n6043 VDD.n647 1.66612
R5605 VDD.n6014 VDD.n645 1.66612
R5606 VDD.n5757 VDD.n5756 1.66612
R5607 VDD.n5789 VDD.n5788 1.66612
R5608 VDD.n5529 VDD.n5528 1.66612
R5609 VDD.n5561 VDD.n5560 1.66612
R5610 VDD.n5301 VDD.n5300 1.66612
R5611 VDD.n5333 VDD.n5332 1.66612
R5612 VDD.n5073 VDD.n5072 1.66612
R5613 VDD.n5105 VDD.n5104 1.66612
R5614 VDD.n5155 VDD.n5154 1.66612
R5615 VDD.n5188 VDD.n1082 1.66612
R5616 VDD.n5383 VDD.n5382 1.66612
R5617 VDD.n5416 VDD.n947 1.66612
R5618 VDD.n5611 VDD.n5610 1.66612
R5619 VDD.n5644 VDD.n812 1.66612
R5620 VDD.n5849 VDD.n5848 1.66612
R5621 VDD.n5884 VDD.n5883 1.66612
R5622 VDD.n5702 VDD.n5701 1.66612
R5623 VDD.n5474 VDD.n5473 1.66612
R5624 VDD.n5246 VDD.n5245 1.66612
R5625 VDD.n6299 VDD.n6298 1.66612
R5626 VDD.n6336 VDD.n6335 1.66612
R5627 VDD.n6369 VDD.n448 1.66612
R5628 VDD.n6525 VDD.n6524 1.66612
R5629 VDD.n6562 VDD.n6561 1.66612
R5630 VDD.n6595 VDD.n314 1.66612
R5631 VDD.n6751 VDD.n6750 1.66612
R5632 VDD.n6788 VDD.n6787 1.66612
R5633 VDD.n6821 VDD.n180 1.66612
R5634 VDD.n6977 VDD.n6976 1.66612
R5635 VDD.n7014 VDD.n7013 1.66612
R5636 VDD.n7047 VDD.n45 1.66612
R5637 VDD.n6961 VDD.n6960 1.66612
R5638 VDD.n6735 VDD.n6734 1.66612
R5639 VDD.n6509 VDD.n6508 1.66612
R5640 VDD.n6283 VDD.n6282 1.66612
R5641 VDD.n6193 VDD.n554 1.66612
R5642 VDD.n2475 VDD.n2464 1.35607
R5643 VDD.n3910 VDD.n3685 1.35607
R5644 VDD.n3902 VDD.n3901 1.35607
R5645 VDD.n3889 VDD.n3728 1.35607
R5646 VDD.n3881 VDD.n3880 1.35607
R5647 VDD.n3923 VDD.n3922 1.35607
R5648 VDD.n3965 VDD.n3552 1.35607
R5649 VDD.n3556 VDD.n3555 1.35607
R5650 VDD.n3947 VDD.n3586 1.35607
R5651 VDD.n3938 VDD.n3616 1.35607
R5652 VDD.n3975 VDD.n3974 1.35607
R5653 VDD.n4029 VDD.n3419 1.35607
R5654 VDD.n4021 VDD.n4020 1.35607
R5655 VDD.n4008 VDD.n3462 1.35607
R5656 VDD.n4000 VDD.n3999 1.35607
R5657 VDD.n4042 VDD.n4041 1.35607
R5658 VDD.n4084 VDD.n3286 1.35607
R5659 VDD.n3290 VDD.n3289 1.35607
R5660 VDD.n4066 VDD.n3320 1.35607
R5661 VDD.n4057 VDD.n3350 1.35607
R5662 VDD.n4094 VDD.n4093 1.35607
R5663 VDD.n4148 VDD.n3153 1.35607
R5664 VDD.n4140 VDD.n4139 1.35607
R5665 VDD.n4127 VDD.n3196 1.35607
R5666 VDD.n4119 VDD.n4118 1.35607
R5667 VDD.n4161 VDD.n4160 1.35607
R5668 VDD.n4203 VDD.n3020 1.35607
R5669 VDD.n3024 VDD.n3023 1.35607
R5670 VDD.n4185 VDD.n3054 1.35607
R5671 VDD.n4176 VDD.n3084 1.35607
R5672 VDD.n4213 VDD.n4212 1.35607
R5673 VDD.n4267 VDD.n2855 1.35607
R5674 VDD.n4259 VDD.n4258 1.35607
R5675 VDD.n4246 VDD.n2930 1.35607
R5676 VDD.n4238 VDD.n4237 1.35607
R5677 VDD.n2894 VDD.n2848 1.35607
R5678 VDD.n4314 VDD.n2778 1.35607
R5679 VDD.n2782 VDD.n2781 1.35607
R5680 VDD.n4296 VDD.n2812 1.35607
R5681 VDD.n4936 VDD.n4934 1.35607
R5682 VDD.n5845 VDD.n5844 1.35607
R5683 VDD.n700 VDD.n699 1.35607
R5684 VDD.n693 VDD.n691 1.35607
R5685 VDD.n5915 VDD.n678 1.35607
R5686 VDD.n5823 VDD.n5822 1.35607
R5687 VDD.n5732 VDD.n5731 1.35607
R5688 VDD.n5745 VDD.n5744 1.35607
R5689 VDD.n5783 VDD.n759 1.35607
R5690 VDD.n5793 VDD.n5792 1.35607
R5691 VDD.n5711 VDD.n5710 1.35607
R5692 VDD.n844 VDD.n842 1.35607
R5693 VDD.n5638 VDD.n831 1.35607
R5694 VDD.n5648 VDD.n5647 1.35607
R5695 VDD.n810 VDD.n808 1.35607
R5696 VDD.n851 VDD.n850 1.35607
R5697 VDD.n5504 VDD.n5503 1.35607
R5698 VDD.n5517 VDD.n5516 1.35607
R5699 VDD.n5555 VDD.n894 1.35607
R5700 VDD.n5565 VDD.n5564 1.35607
R5701 VDD.n5483 VDD.n5482 1.35607
R5702 VDD.n979 VDD.n977 1.35607
R5703 VDD.n5410 VDD.n966 1.35607
R5704 VDD.n5420 VDD.n5419 1.35607
R5705 VDD.n945 VDD.n943 1.35607
R5706 VDD.n986 VDD.n985 1.35607
R5707 VDD.n5276 VDD.n5275 1.35607
R5708 VDD.n5289 VDD.n5288 1.35607
R5709 VDD.n5327 VDD.n1029 1.35607
R5710 VDD.n5337 VDD.n5336 1.35607
R5711 VDD.n5255 VDD.n5254 1.35607
R5712 VDD.n1114 VDD.n1112 1.35607
R5713 VDD.n5182 VDD.n1101 1.35607
R5714 VDD.n5192 VDD.n5191 1.35607
R5715 VDD.n1080 VDD.n1078 1.35607
R5716 VDD.n1121 VDD.n1120 1.35607
R5717 VDD.n5061 VDD.n5060 1.35607
R5718 VDD.n5099 VDD.n1164 1.35607
R5719 VDD.n5109 VDD.n5108 1.35607
R5720 VDD.n5954 VDD.n5952 1.35607
R5721 VDD.n5957 VDD.n5956 1.35607
R5722 VDD.n6037 VDD.n5972 1.35607
R5723 VDD.n6028 VDD.n6027 1.35607
R5724 VDD.n6065 VDD.n658 1.35607
R5725 VDD.n6119 VDD.n6118 1.35607
R5726 VDD.n6211 VDD.n6210 1.35607
R5727 VDD.n6296 VDD.n6295 1.35607
R5728 VDD.n483 VDD.n482 1.35607
R5729 VDD.n476 VDD.n474 1.35607
R5730 VDD.n6363 VDD.n463 1.35607
R5731 VDD.n6373 VDD.n6372 1.35607
R5732 VDD.n6397 VDD.n6396 1.35607
R5733 VDD.n6522 VDD.n6521 1.35607
R5734 VDD.n349 VDD.n348 1.35607
R5735 VDD.n342 VDD.n340 1.35607
R5736 VDD.n6589 VDD.n329 1.35607
R5737 VDD.n6599 VDD.n6598 1.35607
R5738 VDD.n6623 VDD.n6622 1.35607
R5739 VDD.n6748 VDD.n6747 1.35607
R5740 VDD.n215 VDD.n214 1.35607
R5741 VDD.n208 VDD.n206 1.35607
R5742 VDD.n6815 VDD.n195 1.35607
R5743 VDD.n6825 VDD.n6824 1.35607
R5744 VDD.n6849 VDD.n6848 1.35607
R5745 VDD.n6974 VDD.n6973 1.35607
R5746 VDD.n81 VDD.n80 1.35607
R5747 VDD.n74 VDD.n72 1.35607
R5748 VDD.n7041 VDD.n61 1.35607
R5749 VDD.n7051 VDD.n7050 1.35607
R5750 VDD.n7073 VDD.n43 1.35607
R5751 VDD.n6945 VDD.n6944 1.35607
R5752 VDD.n6925 VDD.n6924 1.35607
R5753 VDD.n6916 VDD.n141 1.35607
R5754 VDD.n6889 VDD.n6888 1.35607
R5755 VDD.n6964 VDD.n6963 1.35607
R5756 VDD.n6868 VDD.n6867 1.35607
R5757 VDD.n6719 VDD.n6718 1.35607
R5758 VDD.n6699 VDD.n6698 1.35607
R5759 VDD.n6690 VDD.n275 1.35607
R5760 VDD.n6663 VDD.n6662 1.35607
R5761 VDD.n6738 VDD.n6737 1.35607
R5762 VDD.n6642 VDD.n6641 1.35607
R5763 VDD.n6493 VDD.n6492 1.35607
R5764 VDD.n6473 VDD.n6472 1.35607
R5765 VDD.n6464 VDD.n409 1.35607
R5766 VDD.n6437 VDD.n6436 1.35607
R5767 VDD.n6512 VDD.n6511 1.35607
R5768 VDD.n6416 VDD.n6415 1.35607
R5769 VDD.n6267 VDD.n6266 1.35607
R5770 VDD.n6247 VDD.n6246 1.35607
R5771 VDD.n6238 VDD.n543 1.35607
R5772 VDD.n6286 VDD.n6285 1.35607
R5773 VDD.n6190 VDD.n6189 1.35607
R5774 VDD.n7187 VDD.n7122 1.35607
R5775 VDD.n7107 VDD.n7106 1.35607
R5776 VDD.n7104 VDD.n7102 1.35607
R5777 VDD.n7215 VDD.n29 1.35607
R5778 VDD.n7178 VDD.n7177 1.35607
R5779 VDD.n2633 VDD.n2632 1.35607
R5780 VDD.n4376 VDD.n2443 1.35607
R5781 VDD.n4367 VDD.n2647 1.35607
R5782 VDD.n2651 VDD.n2650 1.35607
R5783 VDD.n4349 VDD.n2686 1.35607
R5784 VDD.n4874 VDD.n1377 1.35607
R5785 VDD.n4447 VDD.n2329 1.35607
R5786 VDD.n4438 VDD.n4437 1.35607
R5787 VDD.n4425 VDD.n2371 1.35607
R5788 VDD.n4416 VDD.n4415 1.35607
R5789 VDD.n4403 VDD.n2413 1.35607
R5790 VDD.n4460 VDD.n4459 1.35607
R5791 VDD.n4502 VDD.n2196 1.35607
R5792 VDD.n2200 VDD.n2199 1.35607
R5793 VDD.n4484 VDD.n2230 1.35607
R5794 VDD.n4475 VDD.n2260 1.35607
R5795 VDD.n2264 VDD.n2263 1.35607
R5796 VDD.n4512 VDD.n4511 1.35607
R5797 VDD.n4568 VDD.n2065 1.35607
R5798 VDD.n4559 VDD.n4558 1.35607
R5799 VDD.n4546 VDD.n2107 1.35607
R5800 VDD.n4537 VDD.n4536 1.35607
R5801 VDD.n4524 VDD.n2149 1.35607
R5802 VDD.n4581 VDD.n4580 1.35607
R5803 VDD.n4623 VDD.n1932 1.35607
R5804 VDD.n1936 VDD.n1935 1.35607
R5805 VDD.n4605 VDD.n1966 1.35607
R5806 VDD.n4596 VDD.n1996 1.35607
R5807 VDD.n2000 VDD.n1999 1.35607
R5808 VDD.n4633 VDD.n4632 1.35607
R5809 VDD.n4689 VDD.n1801 1.35607
R5810 VDD.n4680 VDD.n4679 1.35607
R5811 VDD.n4667 VDD.n1843 1.35607
R5812 VDD.n4658 VDD.n4657 1.35607
R5813 VDD.n4645 VDD.n1885 1.35607
R5814 VDD.n4702 VDD.n4701 1.35607
R5815 VDD.n4744 VDD.n1668 1.35607
R5816 VDD.n1672 VDD.n1671 1.35607
R5817 VDD.n4726 VDD.n1702 1.35607
R5818 VDD.n4717 VDD.n1732 1.35607
R5819 VDD.n1736 VDD.n1735 1.35607
R5820 VDD.n4754 VDD.n4753 1.35607
R5821 VDD.n4810 VDD.n1537 1.35607
R5822 VDD.n4801 VDD.n4800 1.35607
R5823 VDD.n4788 VDD.n1579 1.35607
R5824 VDD.n4779 VDD.n4778 1.35607
R5825 VDD.n4766 VDD.n1621 1.35607
R5826 VDD.n4823 VDD.n4822 1.35607
R5827 VDD.n1404 VDD.n1403 1.35607
R5828 VDD.n4847 VDD.n1438 1.35607
R5829 VDD.n4838 VDD.n1468 1.35607
R5830 VDD.n1472 VDD.n1471 1.35607
R5831 VDD.n4865 VDD.n1400 1.35607
R5832 VDD.n1285 VDD.n1245 1.35607
R5833 VDD.n4917 VDD.n1252 1.35607
R5834 VDD.n1256 VDD.n1255 1.35607
R5835 VDD.n4899 VDD.n1311 1.35607
R5836 VDD.n4890 VDD.n1341 1.35607
R5837 VDD.n4333 VDD.n4332 1.35607
R5838 VDD.n3868 VDD.n3771 1.35607
R5839 VDD.n3620 VDD.n3619 1.35607
R5840 VDD.n3987 VDD.n3505 1.35607
R5841 VDD.n3354 VDD.n3353 1.35607
R5842 VDD.n4106 VDD.n3239 1.35607
R5843 VDD.n3088 VDD.n3087 1.35607
R5844 VDD.n4225 VDD.n2973 1.35607
R5845 VDD.n4287 VDD.n2842 1.35607
R5846 VDD.n4324 VDD.n4323 1.35607
R5847 VDD.n5027 VDD.n5026 1.35607
R5848 VDD.n5923 VDD.n672 1.35607
R5849 VDD.n5813 VDD.n5812 1.35607
R5850 VDD.n5698 VDD.n798 1.35607
R5851 VDD.n5586 VDD.n5585 1.35607
R5852 VDD.n5470 VDD.n933 1.35607
R5853 VDD.n5358 VDD.n5357 1.35607
R5854 VDD.n5242 VDD.n1068 1.35607
R5855 VDD.n5130 VDD.n5129 1.35607
R5856 VDD.n5048 VDD.n5047 1.35607
R5857 VDD.n7264 VDD.n7263 1.35607
R5858 VDD.n3830 VDD.n3829 1.13981
R5859 VDD.n2506 VDD.n2505 1.13981
R5860 VDD.n6117 VDD.n6112 1.13717
R5861 VDD.n7151 VDD.n7146 1.13717
R5862 VDD.n7126 VDD.n7124 1.13717
R5863 VDD.n7136 VDD.n7135 1.13717
R5864 VDD.n7205 VDD.n7204 1.13717
R5865 VDD.n33 VDD.n31 1.13717
R5866 VDD.n7090 VDD.n7089 1.13717
R5867 VDD.n38 VDD.n37 1.13717
R5868 VDD.n7097 VDD.n7096 1.13717
R5869 VDD.n7207 VDD.n7206 1.13717
R5870 VDD.n7134 VDD.n7133 1.13717
R5871 VDD.n7185 VDD.n7184 1.13717
R5872 VDD.n7159 VDD.n7158 1.13717
R5873 VDD.n7058 VDD.n7057 1.13717
R5874 VDD.n6183 VDD.n566 1.13717
R5875 VDD.n41 VDD.n40 1.13717
R5876 VDD.n7054 VDD.n7053 1.13717
R5877 VDD.n54 VDD.n49 1.13717
R5878 VDD.n7033 VDD.n7032 1.13717
R5879 VDD.n67 VDD.n65 1.13717
R5880 VDD.n71 VDD.n70 1.13717
R5881 VDD.n7026 VDD.n7025 1.13717
R5882 VDD.n6995 VDD.n82 1.13717
R5883 VDD.n7003 VDD.n7002 1.13717
R5884 VDD.n6971 VDD.n6970 1.13717
R5885 VDD.n97 VDD.n85 1.13717
R5886 VDD.n6883 VDD.n156 1.13717
R5887 VDD.n6881 VDD.n155 1.13717
R5888 VDD.n6903 VDD.n146 1.13717
R5889 VDD.n6902 VDD.n6901 1.13717
R5890 VDD.n133 VDD.n132 1.13717
R5891 VDD.n6909 VDD.n134 1.13717
R5892 VDD.n122 VDD.n121 1.13717
R5893 VDD.n6931 VDD.n123 1.13717
R5894 VDD.n100 VDD.n99 1.13717
R5895 VDD.n6951 VDD.n101 1.13717
R5896 VDD.n6863 VDD.n167 1.13717
R5897 VDD.n6861 VDD.n166 1.13717
R5898 VDD.n6852 VDD.n6851 1.13717
R5899 VDD.n175 VDD.n171 1.13717
R5900 VDD.n6828 VDD.n6827 1.13717
R5901 VDD.n188 VDD.n184 1.13717
R5902 VDD.n6807 VDD.n6806 1.13717
R5903 VDD.n201 VDD.n199 1.13717
R5904 VDD.n205 VDD.n204 1.13717
R5905 VDD.n6800 VDD.n6799 1.13717
R5906 VDD.n6769 VDD.n216 1.13717
R5907 VDD.n6777 VDD.n6776 1.13717
R5908 VDD.n6745 VDD.n6744 1.13717
R5909 VDD.n231 VDD.n219 1.13717
R5910 VDD.n6657 VDD.n290 1.13717
R5911 VDD.n6655 VDD.n289 1.13717
R5912 VDD.n6677 VDD.n280 1.13717
R5913 VDD.n6676 VDD.n6675 1.13717
R5914 VDD.n267 VDD.n266 1.13717
R5915 VDD.n6683 VDD.n268 1.13717
R5916 VDD.n256 VDD.n255 1.13717
R5917 VDD.n6705 VDD.n257 1.13717
R5918 VDD.n234 VDD.n233 1.13717
R5919 VDD.n6725 VDD.n235 1.13717
R5920 VDD.n6637 VDD.n301 1.13717
R5921 VDD.n6635 VDD.n300 1.13717
R5922 VDD.n6626 VDD.n6625 1.13717
R5923 VDD.n309 VDD.n305 1.13717
R5924 VDD.n6602 VDD.n6601 1.13717
R5925 VDD.n322 VDD.n318 1.13717
R5926 VDD.n6581 VDD.n6580 1.13717
R5927 VDD.n335 VDD.n333 1.13717
R5928 VDD.n339 VDD.n338 1.13717
R5929 VDD.n6574 VDD.n6573 1.13717
R5930 VDD.n6543 VDD.n350 1.13717
R5931 VDD.n6551 VDD.n6550 1.13717
R5932 VDD.n6519 VDD.n6518 1.13717
R5933 VDD.n365 VDD.n353 1.13717
R5934 VDD.n6431 VDD.n424 1.13717
R5935 VDD.n6429 VDD.n423 1.13717
R5936 VDD.n6451 VDD.n414 1.13717
R5937 VDD.n6450 VDD.n6449 1.13717
R5938 VDD.n401 VDD.n400 1.13717
R5939 VDD.n6457 VDD.n402 1.13717
R5940 VDD.n390 VDD.n389 1.13717
R5941 VDD.n6479 VDD.n391 1.13717
R5942 VDD.n368 VDD.n367 1.13717
R5943 VDD.n6499 VDD.n369 1.13717
R5944 VDD.n6411 VDD.n435 1.13717
R5945 VDD.n6409 VDD.n434 1.13717
R5946 VDD.n6400 VDD.n6399 1.13717
R5947 VDD.n443 VDD.n439 1.13717
R5948 VDD.n6376 VDD.n6375 1.13717
R5949 VDD.n456 VDD.n452 1.13717
R5950 VDD.n6355 VDD.n6354 1.13717
R5951 VDD.n469 VDD.n467 1.13717
R5952 VDD.n473 VDD.n472 1.13717
R5953 VDD.n6348 VDD.n6347 1.13717
R5954 VDD.n6317 VDD.n484 1.13717
R5955 VDD.n6325 VDD.n6324 1.13717
R5956 VDD.n6293 VDD.n6292 1.13717
R5957 VDD.n499 VDD.n487 1.13717
R5958 VDD.n6225 VDD.n548 1.13717
R5959 VDD.n6224 VDD.n6223 1.13717
R5960 VDD.n535 VDD.n534 1.13717
R5961 VDD.n6231 VDD.n536 1.13717
R5962 VDD.n524 VDD.n523 1.13717
R5963 VDD.n6253 VDD.n525 1.13717
R5964 VDD.n502 VDD.n501 1.13717
R5965 VDD.n6273 VDD.n503 1.13717
R5966 VDD.n6203 VDD.n557 1.13717
R5967 VDD.n6205 VDD.n558 1.13717
R5968 VDD.n6185 VDD.n567 1.13717
R5969 VDD.n6009 VDD.n6008 1.13717
R5970 VDD.n5976 VDD.n5974 1.13717
R5971 VDD.n5986 VDD.n5985 1.13717
R5972 VDD.n6055 VDD.n6054 1.13717
R5973 VDD.n662 VDD.n660 1.13717
R5974 VDD.n5940 VDD.n5939 1.13717
R5975 VDD.n667 VDD.n666 1.13717
R5976 VDD.n5947 VDD.n5946 1.13717
R5977 VDD.n6057 VDD.n6056 1.13717
R5978 VDD.n5984 VDD.n5983 1.13717
R5979 VDD.n6035 VDD.n6034 1.13717
R5980 VDD.n6001 VDD.n5996 1.13717
R5981 VDD.n4386 VDD.n2434 1.13717
R5982 VDD.n1264 VDD.n1263 1.13717
R5983 VDD.n4883 VDD.n4882 1.13717
R5984 VDD.n1361 VDD.n1349 1.13717
R5985 VDD.n1309 VDD.n1307 1.13717
R5986 VDD.n4910 VDD.n4909 1.13717
R5987 VDD.n1292 VDD.n1260 1.13717
R5988 VDD.n1283 VDD.n1282 1.13717
R5989 VDD.n1300 VDD.n1299 1.13717
R5990 VDD.n4907 VDD.n1258 1.13717
R5991 VDD.n1353 VDD.n1352 1.13717
R5992 VDD.n1369 VDD.n1368 1.13717
R5993 VDD.n4880 VDD.n1347 1.13717
R5994 VDD.n2417 VDD.n2415 1.13717
R5995 VDD.n2420 VDD.n2389 1.13717
R5996 VDD.n2375 VDD.n2373 1.13717
R5997 VDD.n2378 VDD.n2347 1.13717
R5998 VDD.n2333 VDD.n2331 1.13717
R5999 VDD.n2336 VDD.n2297 1.13717
R6000 VDD.n4468 VDD.n4467 1.13717
R6001 VDD.n2280 VDD.n2268 1.13717
R6002 VDD.n2228 VDD.n2226 1.13717
R6003 VDD.n4495 VDD.n4494 1.13717
R6004 VDD.n2211 VDD.n2204 1.13717
R6005 VDD.n4514 VDD.n4513 1.13717
R6006 VDD.n2153 VDD.n2151 1.13717
R6007 VDD.n2156 VDD.n2125 1.13717
R6008 VDD.n2111 VDD.n2109 1.13717
R6009 VDD.n2114 VDD.n2083 1.13717
R6010 VDD.n2069 VDD.n2067 1.13717
R6011 VDD.n2072 VDD.n2033 1.13717
R6012 VDD.n4589 VDD.n4588 1.13717
R6013 VDD.n2016 VDD.n2004 1.13717
R6014 VDD.n1964 VDD.n1962 1.13717
R6015 VDD.n4616 VDD.n4615 1.13717
R6016 VDD.n1947 VDD.n1940 1.13717
R6017 VDD.n4635 VDD.n4634 1.13717
R6018 VDD.n1889 VDD.n1887 1.13717
R6019 VDD.n1892 VDD.n1861 1.13717
R6020 VDD.n1847 VDD.n1845 1.13717
R6021 VDD.n1850 VDD.n1819 1.13717
R6022 VDD.n1805 VDD.n1803 1.13717
R6023 VDD.n1808 VDD.n1769 1.13717
R6024 VDD.n4710 VDD.n4709 1.13717
R6025 VDD.n1752 VDD.n1740 1.13717
R6026 VDD.n1700 VDD.n1698 1.13717
R6027 VDD.n4737 VDD.n4736 1.13717
R6028 VDD.n1683 VDD.n1676 1.13717
R6029 VDD.n4756 VDD.n4755 1.13717
R6030 VDD.n1625 VDD.n1623 1.13717
R6031 VDD.n1628 VDD.n1597 1.13717
R6032 VDD.n1583 VDD.n1581 1.13717
R6033 VDD.n1586 VDD.n1555 1.13717
R6034 VDD.n1541 VDD.n1539 1.13717
R6035 VDD.n1544 VDD.n1505 1.13717
R6036 VDD.n4831 VDD.n4830 1.13717
R6037 VDD.n1488 VDD.n1476 1.13717
R6038 VDD.n1436 VDD.n1434 1.13717
R6039 VDD.n4858 VDD.n4857 1.13717
R6040 VDD.n1419 VDD.n1408 1.13717
R6041 VDD.n1376 VDD.n1375 1.13717
R6042 VDD.n1411 VDD.n1410 1.13717
R6043 VDD.n1427 VDD.n1426 1.13717
R6044 VDD.n4855 VDD.n1406 1.13717
R6045 VDD.n1480 VDD.n1479 1.13717
R6046 VDD.n1496 VDD.n1495 1.13717
R6047 VDD.n4828 VDD.n1474 1.13717
R6048 VDD.n1542 VDD.n1503 1.13717
R6049 VDD.n4808 VDD.n4807 1.13717
R6050 VDD.n1584 VDD.n1553 1.13717
R6051 VDD.n4786 VDD.n4785 1.13717
R6052 VDD.n1626 VDD.n1595 1.13717
R6053 VDD.n4764 VDD.n4763 1.13717
R6054 VDD.n1638 VDD.n1637 1.13717
R6055 VDD.n1691 VDD.n1690 1.13717
R6056 VDD.n4734 VDD.n1674 1.13717
R6057 VDD.n1744 VDD.n1743 1.13717
R6058 VDD.n1760 VDD.n1759 1.13717
R6059 VDD.n4707 VDD.n1738 1.13717
R6060 VDD.n1806 VDD.n1767 1.13717
R6061 VDD.n4687 VDD.n4686 1.13717
R6062 VDD.n1848 VDD.n1817 1.13717
R6063 VDD.n4665 VDD.n4664 1.13717
R6064 VDD.n1890 VDD.n1859 1.13717
R6065 VDD.n4643 VDD.n4642 1.13717
R6066 VDD.n1902 VDD.n1901 1.13717
R6067 VDD.n1955 VDD.n1954 1.13717
R6068 VDD.n4613 VDD.n1938 1.13717
R6069 VDD.n2008 VDD.n2007 1.13717
R6070 VDD.n2024 VDD.n2023 1.13717
R6071 VDD.n4586 VDD.n2002 1.13717
R6072 VDD.n2070 VDD.n2031 1.13717
R6073 VDD.n4566 VDD.n4565 1.13717
R6074 VDD.n2112 VDD.n2081 1.13717
R6075 VDD.n4544 VDD.n4543 1.13717
R6076 VDD.n2154 VDD.n2123 1.13717
R6077 VDD.n4522 VDD.n4521 1.13717
R6078 VDD.n2166 VDD.n2165 1.13717
R6079 VDD.n2219 VDD.n2218 1.13717
R6080 VDD.n4492 VDD.n2202 1.13717
R6081 VDD.n2272 VDD.n2271 1.13717
R6082 VDD.n2288 VDD.n2287 1.13717
R6083 VDD.n4465 VDD.n2266 1.13717
R6084 VDD.n2334 VDD.n2295 1.13717
R6085 VDD.n4445 VDD.n4444 1.13717
R6086 VDD.n2376 VDD.n2345 1.13717
R6087 VDD.n4423 VDD.n4422 1.13717
R6088 VDD.n2418 VDD.n2387 1.13717
R6089 VDD.n4401 VDD.n4400 1.13717
R6090 VDD.n2610 VDD.n2609 1.13717
R6091 VDD.n2733 VDD.n2715 1.13717
R6092 VDD.n2684 VDD.n2682 1.13717
R6093 VDD.n4360 VDD.n4359 1.13717
R6094 VDD.n2667 VDD.n2655 1.13717
R6095 VDD.n2441 VDD.n2439 1.13717
R6096 VDD.n4384 VDD.n2433 1.13717
R6097 VDD.n2659 VDD.n2658 1.13717
R6098 VDD.n2675 VDD.n2674 1.13717
R6099 VDD.n4357 VDD.n2653 1.13717
R6100 VDD.n2721 VDD.n2720 1.13717
R6101 VDD.n2735 VDD.n2716 1.13717
R6102 VDD.n2744 VDD.n2742 1.13717
R6103 VDD.n2747 VDD.n2745 1.13717
R6104 VDD.n2801 VDD.n2800 1.13717
R6105 VDD.n4304 VDD.n2784 1.13717
R6106 VDD.n2870 VDD.n2869 1.13717
R6107 VDD.n2885 VDD.n2865 1.13717
R6108 VDD.n2892 VDD.n2891 1.13717
R6109 VDD.n2903 VDD.n2859 1.13717
R6110 VDD.n2937 VDD.n2905 1.13717
R6111 VDD.n2946 VDD.n2934 1.13717
R6112 VDD.n2978 VDD.n2948 1.13717
R6113 VDD.n4223 VDD.n4222 1.13717
R6114 VDD.n2990 VDD.n2989 1.13717
R6115 VDD.n3043 VDD.n3042 1.13717
R6116 VDD.n4193 VDD.n3026 1.13717
R6117 VDD.n3096 VDD.n3095 1.13717
R6118 VDD.n3112 VDD.n3111 1.13717
R6119 VDD.n4166 VDD.n3090 1.13717
R6120 VDD.n3160 VDD.n3119 1.13717
R6121 VDD.n3169 VDD.n3157 1.13717
R6122 VDD.n3203 VDD.n3171 1.13717
R6123 VDD.n3212 VDD.n3200 1.13717
R6124 VDD.n3244 VDD.n3214 1.13717
R6125 VDD.n4104 VDD.n4103 1.13717
R6126 VDD.n3256 VDD.n3255 1.13717
R6127 VDD.n3309 VDD.n3308 1.13717
R6128 VDD.n4074 VDD.n3292 1.13717
R6129 VDD.n3362 VDD.n3361 1.13717
R6130 VDD.n3378 VDD.n3377 1.13717
R6131 VDD.n4047 VDD.n3356 1.13717
R6132 VDD.n3426 VDD.n3385 1.13717
R6133 VDD.n3435 VDD.n3423 1.13717
R6134 VDD.n3469 VDD.n3437 1.13717
R6135 VDD.n3478 VDD.n3466 1.13717
R6136 VDD.n3510 VDD.n3480 1.13717
R6137 VDD.n3985 VDD.n3984 1.13717
R6138 VDD.n3522 VDD.n3521 1.13717
R6139 VDD.n3575 VDD.n3574 1.13717
R6140 VDD.n3955 VDD.n3558 1.13717
R6141 VDD.n3628 VDD.n3627 1.13717
R6142 VDD.n3644 VDD.n3643 1.13717
R6143 VDD.n3928 VDD.n3622 1.13717
R6144 VDD.n3692 VDD.n3651 1.13717
R6145 VDD.n3701 VDD.n3689 1.13717
R6146 VDD.n3735 VDD.n3703 1.13717
R6147 VDD.n3744 VDD.n3732 1.13717
R6148 VDD.n3776 VDD.n3746 1.13717
R6149 VDD.n3866 VDD.n3865 1.13717
R6150 VDD.n3909 VDD.n3908 1.13717
R6151 VDD.n3737 VDD.n3705 1.13717
R6152 VDD.n3888 VDD.n3887 1.13717
R6153 VDD.n3778 VDD.n3748 1.13717
R6154 VDD.n3775 VDD.n3773 1.13717
R6155 VDD.n3694 VDD.n3653 1.13717
R6156 VDD.n3567 VDD.n3560 1.13717
R6157 VDD.n3958 VDD.n3957 1.13717
R6158 VDD.n3584 VDD.n3582 1.13717
R6159 VDD.n3636 VDD.n3624 1.13717
R6160 VDD.n3931 VDD.n3930 1.13717
R6161 VDD.n3977 VDD.n3976 1.13717
R6162 VDD.n4028 VDD.n4027 1.13717
R6163 VDD.n3471 VDD.n3439 1.13717
R6164 VDD.n4007 VDD.n4006 1.13717
R6165 VDD.n3512 VDD.n3482 1.13717
R6166 VDD.n3509 VDD.n3507 1.13717
R6167 VDD.n3428 VDD.n3387 1.13717
R6168 VDD.n3301 VDD.n3294 1.13717
R6169 VDD.n4077 VDD.n4076 1.13717
R6170 VDD.n3318 VDD.n3316 1.13717
R6171 VDD.n3370 VDD.n3358 1.13717
R6172 VDD.n4050 VDD.n4049 1.13717
R6173 VDD.n4096 VDD.n4095 1.13717
R6174 VDD.n4147 VDD.n4146 1.13717
R6175 VDD.n3205 VDD.n3173 1.13717
R6176 VDD.n4126 VDD.n4125 1.13717
R6177 VDD.n3246 VDD.n3216 1.13717
R6178 VDD.n3243 VDD.n3241 1.13717
R6179 VDD.n3162 VDD.n3121 1.13717
R6180 VDD.n3035 VDD.n3028 1.13717
R6181 VDD.n4196 VDD.n4195 1.13717
R6182 VDD.n3052 VDD.n3050 1.13717
R6183 VDD.n3104 VDD.n3092 1.13717
R6184 VDD.n4169 VDD.n4168 1.13717
R6185 VDD.n4215 VDD.n4214 1.13717
R6186 VDD.n4266 VDD.n4265 1.13717
R6187 VDD.n2939 VDD.n2907 1.13717
R6188 VDD.n4245 VDD.n4244 1.13717
R6189 VDD.n2980 VDD.n2950 1.13717
R6190 VDD.n2977 VDD.n2975 1.13717
R6191 VDD.n2895 VDD.n2862 1.13717
R6192 VDD.n2793 VDD.n2786 1.13717
R6193 VDD.n4307 VDD.n4306 1.13717
R6194 VDD.n2810 VDD.n2808 1.13717
R6195 VDD.n2884 VDD.n2883 1.13717
R6196 VDD.n4326 VDD.n4325 1.13717
R6197 VDD.n2738 VDD.n2737 1.13717
R6198 VDD.n4946 VDD.n4945 1.13717
R6199 VDD.n1196 VDD.n1195 1.13717
R6200 VDD.n1185 VDD.n1184 1.13717
R6201 VDD.n5055 VDD.n1183 1.13717
R6202 VDD.n5086 VDD.n1169 1.13717
R6203 VDD.n1156 VDD.n1155 1.13717
R6204 VDD.n5114 VDD.n1125 1.13717
R6205 VDD.n5136 VDD.n1122 1.13717
R6206 VDD.n1111 VDD.n1110 1.13717
R6207 VDD.n5174 VDD.n5173 1.13717
R6208 VDD.n5195 VDD.n5194 1.13717
R6209 VDD.n1077 VDD.n1076 1.13717
R6210 VDD.n5230 VDD.n5229 1.13717
R6211 VDD.n1061 VDD.n1060 1.13717
R6212 VDD.n1050 VDD.n1049 1.13717
R6213 VDD.n5283 VDD.n1048 1.13717
R6214 VDD.n5314 VDD.n1034 1.13717
R6215 VDD.n1021 VDD.n1020 1.13717
R6216 VDD.n5342 VDD.n990 1.13717
R6217 VDD.n5364 VDD.n987 1.13717
R6218 VDD.n976 VDD.n975 1.13717
R6219 VDD.n5402 VDD.n5401 1.13717
R6220 VDD.n5423 VDD.n5422 1.13717
R6221 VDD.n942 VDD.n941 1.13717
R6222 VDD.n5458 VDD.n5457 1.13717
R6223 VDD.n926 VDD.n925 1.13717
R6224 VDD.n915 VDD.n914 1.13717
R6225 VDD.n5511 VDD.n913 1.13717
R6226 VDD.n5542 VDD.n899 1.13717
R6227 VDD.n886 VDD.n885 1.13717
R6228 VDD.n5570 VDD.n855 1.13717
R6229 VDD.n5592 VDD.n852 1.13717
R6230 VDD.n841 VDD.n840 1.13717
R6231 VDD.n5630 VDD.n5629 1.13717
R6232 VDD.n5651 VDD.n5650 1.13717
R6233 VDD.n807 VDD.n806 1.13717
R6234 VDD.n5686 VDD.n5685 1.13717
R6235 VDD.n791 VDD.n790 1.13717
R6236 VDD.n780 VDD.n779 1.13717
R6237 VDD.n5739 VDD.n778 1.13717
R6238 VDD.n5770 VDD.n764 1.13717
R6239 VDD.n751 VDD.n750 1.13717
R6240 VDD.n729 VDD.n728 1.13717
R6241 VDD.n5819 VDD.n5818 1.13717
R6242 VDD.n5841 VDD.n5840 1.13717
R6243 VDD.n5865 VDD.n701 1.13717
R6244 VDD.n690 VDD.n689 1.13717
R6245 VDD.n5903 VDD.n5902 1.13717
R6246 VDD.n5907 VDD.n5906 1.13717
R6247 VDD.n5843 VDD.n704 1.13717
R6248 VDD.n5873 VDD.n5872 1.13717
R6249 VDD.n5896 VDD.n5895 1.13717
R6250 VDD.n685 VDD.n682 1.13717
R6251 VDD.n670 VDD.n669 1.13717
R6252 VDD.n5821 VDD.n721 1.13717
R6253 VDD.n5717 VDD.n781 1.13717
R6254 VDD.n5747 VDD.n5746 1.13717
R6255 VDD.n5769 VDD.n5768 1.13717
R6256 VDD.n5776 VDD.n752 1.13717
R6257 VDD.n5799 VDD.n730 1.13717
R6258 VDD.n5689 VDD.n792 1.13717
R6259 VDD.n5623 VDD.n5622 1.13717
R6260 VDD.n837 VDD.n835 1.13717
R6261 VDD.n823 VDD.n817 1.13717
R6262 VDD.n5679 VDD.n5678 1.13717
R6263 VDD.n802 VDD.n799 1.13717
R6264 VDD.n5600 VDD.n5599 1.13717
R6265 VDD.n5489 VDD.n916 1.13717
R6266 VDD.n5519 VDD.n5518 1.13717
R6267 VDD.n5541 VDD.n5540 1.13717
R6268 VDD.n5548 VDD.n887 1.13717
R6269 VDD.n5572 VDD.n856 1.13717
R6270 VDD.n5461 VDD.n927 1.13717
R6271 VDD.n5395 VDD.n5394 1.13717
R6272 VDD.n972 VDD.n970 1.13717
R6273 VDD.n958 VDD.n952 1.13717
R6274 VDD.n5451 VDD.n5450 1.13717
R6275 VDD.n937 VDD.n934 1.13717
R6276 VDD.n5372 VDD.n5371 1.13717
R6277 VDD.n5261 VDD.n1051 1.13717
R6278 VDD.n5291 VDD.n5290 1.13717
R6279 VDD.n5313 VDD.n5312 1.13717
R6280 VDD.n5320 VDD.n1022 1.13717
R6281 VDD.n5344 VDD.n991 1.13717
R6282 VDD.n5233 VDD.n1062 1.13717
R6283 VDD.n5167 VDD.n5166 1.13717
R6284 VDD.n1107 VDD.n1105 1.13717
R6285 VDD.n1093 VDD.n1087 1.13717
R6286 VDD.n5223 VDD.n5222 1.13717
R6287 VDD.n1072 VDD.n1069 1.13717
R6288 VDD.n5144 VDD.n5143 1.13717
R6289 VDD.n5063 VDD.n5062 1.13717
R6290 VDD.n5085 VDD.n5084 1.13717
R6291 VDD.n5092 VDD.n1157 1.13717
R6292 VDD.n5116 VDD.n1126 1.13717
R6293 VDD.n5033 VDD.n1186 1.13717
R6294 VDD.n5022 VDD.n1197 1.13717
R6295 VDD.n3786 VDD.n3785 1.13462
R6296 VDD.n3790 VDD.n3789 1.13462
R6297 VDD.n3794 VDD.n3793 1.13462
R6298 VDD.n3798 VDD.n3797 1.13462
R6299 VDD.n3802 VDD.n3801 1.13462
R6300 VDD.n2530 VDD.n2529 1.13462
R6301 VDD.n2557 VDD.n2556 1.13462
R6302 VDD.n2493 VDD.n2492 1.13462
R6303 VDD.n2499 VDD.n2498 1.13462
R6304 VDD.n2532 VDD.n2531 1.13462
R6305 VDD.n2590 VDD.n2589 1.13462
R6306 VDD.n2571 VDD.n2570 1.13462
R6307 VDD.n2577 VDD.n2576 1.13462
R6308 VDD.n597 VDD.n596 1.13005
R6309 VDD.n3841 VDD.n3840 1.13005
R6310 VDD.n2517 VDD.n2516 1.13005
R6311 VDD.n1227 VDD.n1226 1.13005
R6312 VDD.n3826 VDD.n3804 1.04044
R6313 VDD.n3814 VDD.n3812 1.04044
R6314 VDD.n3817 VDD.n3815 1.04044
R6315 VDD.n3811 VDD.n3809 1.04044
R6316 VDD.n3807 VDD.n3805 1.04044
R6317 VDD.n2578 VDD.n2565 1.04044
R6318 VDD.n2572 VDD.n2566 1.04044
R6319 VDD.n2593 VDD.n2567 1.04044
R6320 VDD.n2542 VDD.n2534 1.04044
R6321 VDD.n2502 VDD.n2501 1.04044
R6322 VDD.n2494 VDD.n2488 1.04044
R6323 VDD.n2560 VDD.n2489 1.04044
R6324 VDD.n2550 VDD.n2549 1.04044
R6325 VDD.n6108 VDD.n6107 1.04017
R6326 VDD.n624 VDD.n623 1.04017
R6327 VDD.n6100 VDD.n6099 1.04017
R6328 VDD.n6154 VDD.n6153 1.04017
R6329 VDD.n6164 VDD.n6163 1.04017
R6330 VDD.n6145 VDD.n6144 1.04017
R6331 VDD.n587 VDD.n586 1.04017
R6332 VDD.n6172 VDD.n6171 1.04017
R6333 VDD.n5011 VDD.n5010 1.04017
R6334 VDD.n4997 VDD.n4996 1.04017
R6335 VDD.n5003 VDD.n5002 1.04017
R6336 VDD.n4988 VDD.n4987 1.04017
R6337 VDD.n1217 VDD.n1216 1.04017
R6338 VDD.n6121 VDD.n607 1.01637
R6339 VDD.n2484 VDD.n2483 1.01637
R6340 VDD.n4965 VDD.n1237 1.01637
R6341 VDD.n7276 VDD.n7275 1.01637
R6342 VDD.n4980 VDD.n4979 0.936863
R6343 VDD.t11 VDD 0.918966
R6344 VDD.t60 VDD 0.918966
R6345 VDD.n632 VDD.n613 0.870766
R6346 VDD.n7238 VDD.n7237 0.870766
R6347 VDD.n6134 VDD.n601 0.870578
R6348 VDD.n2468 VDD.n2466 0.870578
R6349 VDD.n2615 VDD.n2614 0.870578
R6350 VDD.n4940 VDD.n1232 0.870578
R6351 VDD.n4951 VDD.n4950 0.870578
R6352 VDD.n7247 VDD.n7246 0.870578
R6353 VDD.n590 VDD.n589 0.853291
R6354 VDD.n1220 VDD.n1219 0.853291
R6355 VDD.n6118 VDD.n6117 0.853
R6356 VDD.n6 VDD.n5 0.853
R6357 VDD.n572 VDD.n571 0.853
R6358 VDD.n579 VDD.n571 0.853
R6359 VDD.n585 VDD.n584 0.853
R6360 VDD.n584 VDD.n575 0.853
R6361 VDD.n6143 VDD.n576 0.853
R6362 VDD.n6167 VDD.n576 0.853
R6363 VDD.n6166 VDD.n578 0.853
R6364 VDD.n6167 VDD.n6166 0.853
R6365 VDD.n6152 VDD.n6151 0.853
R6366 VDD.n6151 VDD.n575 0.853
R6367 VDD.n569 VDD.n568 0.853
R6368 VDD.n6102 VDD.n629 0.853
R6369 VDD.n6103 VDD.n6102 0.853
R6370 VDD.n626 VDD.n625 0.853
R6371 VDD.n627 VDD.n626 0.853
R6372 VDD.n618 VDD.n617 0.853
R6373 VDD.n627 VDD.n617 0.853
R6374 VDD.n635 VDD.n634 0.853
R6375 VDD.n3859 VDD.n3787 0.853
R6376 VDD.n3856 VDD.n3791 0.853
R6377 VDD.n3853 VDD.n3795 0.853
R6378 VDD.n3850 VDD.n3799 0.853
R6379 VDD.n3847 VDD.n3803 0.853
R6380 VDD.n1271 VDD.n1270 0.853
R6381 VDD.n2553 VDD.n2548 0.853
R6382 VDD.n2491 VDD.n2490 0.853
R6383 VDD.n2526 VDD.n2495 0.853
R6384 VDD.n2523 VDD.n2500 0.853
R6385 VDD.n2545 VDD.n2533 0.853
R6386 VDD.n2609 VDD.n2464 0.853
R6387 VDD.n2569 VDD.n2568 0.853
R6388 VDD.n2585 VDD.n2573 0.853
R6389 VDD.n2582 VDD.n2579 0.853
R6390 VDD.n4391 VDD.n2428 0.853
R6391 VDD.n4945 VDD.n4936 0.853
R6392 VDD.n1215 VDD.n1214 0.853
R6393 VDD.n1214 VDD.n1205 0.853
R6394 VDD.n4986 VDD.n1206 0.853
R6395 VDD.n5006 VDD.n1206 0.853
R6396 VDD.n5005 VDD.n1208 0.853
R6397 VDD.n5006 VDD.n5005 0.853
R6398 VDD.n4995 VDD.n4994 0.853
R6399 VDD.n4994 VDD.n1205 0.853
R6400 VDD.n1199 VDD.n1198 0.853
R6401 VDD.n1202 VDD.n1201 0.853
R6402 VDD.n1209 VDD.n1201 0.853
R6403 VDD.n7263 VDD.n7262 0.853
R6404 VDD.n3842 VDD.n3841 0.851407
R6405 VDD.n2518 VDD.n2517 0.851407
R6406 VDD.n7081 VDD.n23 0.84923
R6407 VDD.n4340 VDD.n4339 0.84923
R6408 VDD.n1345 VDD.n1344 0.84923
R6409 VDD.n5931 VDD.n652 0.849012
R6410 VDD.n6094 VDD.n630 0.813198
R6411 VDD.n6123 VDD.n6121 0.813198
R6412 VDD.n2483 VDD.n2474 0.813198
R6413 VDD.n2620 VDD.n2619 0.813198
R6414 VDD.n4965 VDD.n4933 0.813198
R6415 VDD.n4957 VDD.n4956 0.813198
R6416 VDD.n6156 VDD.n0 0.813198
R6417 VDD.n7275 VDD.n7268 0.813198
R6418 VDD.n2628 VDD.n2449 0.734658
R6419 VDD.n4373 VDD.n2641 0.734658
R6420 VDD.n4371 VDD.n2642 0.734658
R6421 VDD.n2698 VDD.n2692 0.734658
R6422 VDD.n4346 VDD.n2710 0.734658
R6423 VDD.n4344 VDD.n2711 0.734658
R6424 VDD.n2760 VDD.n2757 0.734658
R6425 VDD.n4320 VDD.n2772 0.734658
R6426 VDD.n4318 VDD.n2773 0.734658
R6427 VDD.n2824 VDD.n2818 0.734658
R6428 VDD.n4293 VDD.n2836 0.734658
R6429 VDD.n4291 VDD.n2837 0.734658
R6430 VDD.n4276 VDD.n4275 0.734658
R6431 VDD.n2924 VDD.n2851 0.734658
R6432 VDD.n4255 VDD.n4254 0.734658
R6433 VDD.n2967 VDD.n2926 0.734658
R6434 VDD.n4234 VDD.n4233 0.734658
R6435 VDD.n3007 VDD.n2969 0.734658
R6436 VDD.n4209 VDD.n3014 0.734658
R6437 VDD.n4207 VDD.n3015 0.734658
R6438 VDD.n3066 VDD.n3060 0.734658
R6439 VDD.n4182 VDD.n3078 0.734658
R6440 VDD.n4180 VDD.n3079 0.734658
R6441 VDD.n3147 VDD.n3127 0.734658
R6442 VDD.n4157 VDD.n4156 0.734658
R6443 VDD.n3190 VDD.n3149 0.734658
R6444 VDD.n4136 VDD.n4135 0.734658
R6445 VDD.n3233 VDD.n3192 0.734658
R6446 VDD.n4115 VDD.n4114 0.734658
R6447 VDD.n3273 VDD.n3235 0.734658
R6448 VDD.n4090 VDD.n3280 0.734658
R6449 VDD.n4088 VDD.n3281 0.734658
R6450 VDD.n3332 VDD.n3326 0.734658
R6451 VDD.n4063 VDD.n3344 0.734658
R6452 VDD.n4061 VDD.n3345 0.734658
R6453 VDD.n3413 VDD.n3393 0.734658
R6454 VDD.n4038 VDD.n4037 0.734658
R6455 VDD.n3456 VDD.n3415 0.734658
R6456 VDD.n4017 VDD.n4016 0.734658
R6457 VDD.n3499 VDD.n3458 0.734658
R6458 VDD.n3996 VDD.n3995 0.734658
R6459 VDD.n3539 VDD.n3501 0.734658
R6460 VDD.n3971 VDD.n3546 0.734658
R6461 VDD.n3969 VDD.n3547 0.734658
R6462 VDD.n3598 VDD.n3592 0.734658
R6463 VDD.n3944 VDD.n3610 0.734658
R6464 VDD.n3942 VDD.n3611 0.734658
R6465 VDD.n3679 VDD.n3659 0.734658
R6466 VDD.n3919 VDD.n3918 0.734658
R6467 VDD.n3722 VDD.n3681 0.734658
R6468 VDD.n3898 VDD.n3897 0.734658
R6469 VDD.n3765 VDD.n3724 0.734658
R6470 VDD.n3877 VDD.n3876 0.734658
R6471 VDD.n3818 VDD.n3767 0.734658
R6472 VDD.n3825 VDD.n3824 0.734658
R6473 VDD.n4923 VDD.n1242 0.734658
R6474 VDD.n4921 VDD.n1247 0.734658
R6475 VDD.n1323 VDD.n1317 0.734658
R6476 VDD.n4896 VDD.n1335 0.734658
R6477 VDD.n4894 VDD.n1336 0.734658
R6478 VDD.n1392 VDD.n1383 0.734658
R6479 VDD.n4871 VDD.n1394 0.734658
R6480 VDD.n4869 VDD.n1395 0.734658
R6481 VDD.n1450 VDD.n1444 0.734658
R6482 VDD.n4844 VDD.n1462 0.734658
R6483 VDD.n4842 VDD.n1463 0.734658
R6484 VDD.n1531 VDD.n1511 0.734658
R6485 VDD.n4819 VDD.n4818 0.734658
R6486 VDD.n1573 VDD.n1533 0.734658
R6487 VDD.n4797 VDD.n4796 0.734658
R6488 VDD.n1615 VDD.n1575 0.734658
R6489 VDD.n4775 VDD.n4774 0.734658
R6490 VDD.n1655 VDD.n1617 0.734658
R6491 VDD.n4750 VDD.n1662 0.734658
R6492 VDD.n4748 VDD.n1663 0.734658
R6493 VDD.n1714 VDD.n1708 0.734658
R6494 VDD.n4723 VDD.n1726 0.734658
R6495 VDD.n4721 VDD.n1727 0.734658
R6496 VDD.n1795 VDD.n1775 0.734658
R6497 VDD.n4698 VDD.n4697 0.734658
R6498 VDD.n1837 VDD.n1797 0.734658
R6499 VDD.n4676 VDD.n4675 0.734658
R6500 VDD.n1879 VDD.n1839 0.734658
R6501 VDD.n4654 VDD.n4653 0.734658
R6502 VDD.n1919 VDD.n1881 0.734658
R6503 VDD.n4629 VDD.n1926 0.734658
R6504 VDD.n4627 VDD.n1927 0.734658
R6505 VDD.n1978 VDD.n1972 0.734658
R6506 VDD.n4602 VDD.n1990 0.734658
R6507 VDD.n4600 VDD.n1991 0.734658
R6508 VDD.n2059 VDD.n2039 0.734658
R6509 VDD.n4577 VDD.n4576 0.734658
R6510 VDD.n2101 VDD.n2061 0.734658
R6511 VDD.n4555 VDD.n4554 0.734658
R6512 VDD.n2143 VDD.n2103 0.734658
R6513 VDD.n4533 VDD.n4532 0.734658
R6514 VDD.n2183 VDD.n2145 0.734658
R6515 VDD.n4508 VDD.n2190 0.734658
R6516 VDD.n4506 VDD.n2191 0.734658
R6517 VDD.n2242 VDD.n2236 0.734658
R6518 VDD.n4481 VDD.n2254 0.734658
R6519 VDD.n4479 VDD.n2255 0.734658
R6520 VDD.n2323 VDD.n2303 0.734658
R6521 VDD.n4456 VDD.n4455 0.734658
R6522 VDD.n2365 VDD.n2325 0.734658
R6523 VDD.n4434 VDD.n4433 0.734658
R6524 VDD.n2407 VDD.n2367 0.734658
R6525 VDD.n4412 VDD.n4411 0.734658
R6526 VDD.n2535 VDD.n2409 0.734658
R6527 VDD.n2561 VDD.n2487 0.734658
R6528 VDD.n3831 VDD.n3830 0.684595
R6529 VDD.n2507 VDD.n2506 0.684595
R6530 VDD.n7258 VDD.n7257 0.682713
R6531 VDD.n6133 VDD.n600 0.682713
R6532 VDD.n6087 VDD.n6086 0.682713
R6533 VDD.n2616 VDD.n2458 0.682713
R6534 VDD.n2605 VDD.n2604 0.682713
R6535 VDD.n4952 VDD.n4938 0.682713
R6536 VDD.n4976 VDD.n4975 0.682713
R6537 VDD.n7230 VDD.n7229 0.682707
R6538 VDD.n6177 VDD.n6176 0.682697
R6539 VDD.n5016 VDD.n5015 0.682697
R6540 VDD.n6080 VDD.n6079 0.682447
R6541 VDD.n4392 VDD.n2429 0.682447
R6542 VDD.n1273 VDD.n1272 0.682447
R6543 VDD.t8 VDD.n638 0.612811
R6544 VDD.t1 VDD.n9 0.612811
R6545 VDD.n5019 VDD 0.547714
R6546 VDD.n2850 VDD 0.534441
R6547 VDD.n3148 VDD 0.534441
R6548 VDD.n3414 VDD 0.534441
R6549 VDD.n3680 VDD 0.534441
R6550 VDD.n1532 VDD 0.534441
R6551 VDD.n1796 VDD 0.534441
R6552 VDD.n2060 VDD 0.534441
R6553 VDD.n2324 VDD 0.534441
R6554 VDD.n6073 VDD.n641 0.459733
R6555 VDD.n7223 VDD.n12 0.459733
R6556 VDD.t26 VDD.n4998 0.454532
R6557 VDD.t10 VDD.n6155 0.454532
R6558 VDD.n4998 VDD.t22 0.45205
R6559 VDD.n6155 VDD.t7 0.45205
R6560 VDD.n6130 VDD.n6129 0.406849
R6561 VDD.n2473 VDD.n2472 0.406849
R6562 VDD.n1236 VDD.n1235 0.406849
R6563 VDD.n7254 VDD.n7253 0.406849
R6564 VDD.n3843 VDD.n3842 0.370457
R6565 VDD.n2519 VDD.n2518 0.370457
R6566 VDD.n6138 VDD.n598 0.35535
R6567 VDD.n4981 VDD.n1228 0.35535
R6568 VDD.n7077 VDD 0.321584
R6569 VDD.n7078 VDD 0.317995
R6570 VDD.n5241 VDD.n1063 0.314894
R6571 VDD.n5469 VDD.n928 0.314894
R6572 VDD.n5697 VDD.n793 0.314894
R6573 VDD.n445 VDD.n433 0.314894
R6574 VDD.n311 VDD.n299 0.314894
R6575 VDD.n177 VDD.n165 0.314894
R6576 VDD.n2998 VDD.n2997 0.314894
R6577 VDD.n3264 VDD.n3263 0.314894
R6578 VDD.n3530 VDD.n3529 0.314894
R6579 VDD.n1646 VDD.n1645 0.314894
R6580 VDD.n1910 VDD.n1909 0.314894
R6581 VDD.n2174 VDD.n2173 0.314894
R6582 VDD.n1145 VDD.n1132 0.30353
R6583 VDD.n1010 VDD.n997 0.30353
R6584 VDD.n875 VDD.n862 0.30353
R6585 VDD.n740 VDD.n737 0.30353
R6586 VDD.n513 VDD.n510 0.30353
R6587 VDD.n379 VDD.n376 0.30353
R6588 VDD.n245 VDD.n242 0.30353
R6589 VDD.n111 VDD.n108 0.30353
R6590 VDD.n512 VDD.n511 0.30353
R6591 VDD.n378 VDD.n377 0.30353
R6592 VDD.n244 VDD.n243 0.30353
R6593 VDD.n110 VDD.n109 0.30353
R6594 VDD.n4283 VDD.n4282 0.30353
R6595 VDD.n3140 VDD.n3139 0.30353
R6596 VDD.n3406 VDD.n3405 0.30353
R6597 VDD.n3672 VDD.n3671 0.30353
R6598 VDD.n1524 VDD.n1523 0.30353
R6599 VDD.n1788 VDD.n1787 0.30353
R6600 VDD.n2052 VDD.n2051 0.30353
R6601 VDD.n2316 VDD.n2315 0.30353
R6602 VDD.n1525 VDD.n1520 0.30353
R6603 VDD.n1789 VDD.n1784 0.30353
R6604 VDD.n2053 VDD.n2048 0.30353
R6605 VDD.n2317 VDD.n2312 0.30353
R6606 VDD.n4284 VDD.n2844 0.30353
R6607 VDD.n3141 VDD.n3136 0.30353
R6608 VDD.n3407 VDD.n3402 0.30353
R6609 VDD.n3673 VDD.n3668 0.30353
R6610 VDD.n1144 VDD.n1143 0.30353
R6611 VDD.n1009 VDD.n1008 0.30353
R6612 VDD.n874 VDD.n873 0.30353
R6613 VDD.n739 VDD.n738 0.30353
R6614 VDD.n6407 VDD.n6405 0.288379
R6615 VDD.n6633 VDD.n6631 0.288379
R6616 VDD.n6859 VDD.n6857 0.288379
R6617 VDD.n1643 VDD.n1642 0.288379
R6618 VDD.n1907 VDD.n1906 0.288379
R6619 VDD.n2171 VDD.n2170 0.288379
R6620 VDD.n2995 VDD.n2994 0.288379
R6621 VDD.n3261 VDD.n3260 0.288379
R6622 VDD.n3527 VDD.n3526 0.288379
R6623 VDD.n5239 VDD.n1071 0.288379
R6624 VDD.n5467 VDD.n936 0.288379
R6625 VDD.n5695 VDD.n801 0.288379
R6626 VDD.n6180 VDD 0.266176
R6627 VDD.n6071 VDD.n6070 0.194439
R6628 VDD.n6066 VDD.n654 0.194439
R6629 VDD.n6066 VDD.n656 0.194439
R6630 VDD.n5965 VDD.n5963 0.194439
R6631 VDD.n5967 VDD.n5965 0.194439
R6632 VDD.n6047 VDD.n6046 0.194439
R6633 VDD.n6046 VDD.n6044 0.194439
R6634 VDD.n6012 VDD.n5970 0.194439
R6635 VDD.n6013 VDD.n6012 0.194439
R6636 VDD.n6026 VDD.n6024 0.194439
R6637 VDD.n6026 VDD.n639 0.194439
R6638 VDD.n6191 VDD.n564 0.194439
R6639 VDD.n6212 VDD.n555 0.194439
R6640 VDD.n6212 VDD.n553 0.194439
R6641 VDD.n6239 VDD.n540 0.194439
R6642 VDD.n6239 VDD.n541 0.194439
R6643 VDD.n6245 VDD.n6244 0.194439
R6644 VDD.n6245 VDD.n529 0.194439
R6645 VDD.n6265 VDD.n527 0.194439
R6646 VDD.n6265 VDD.n518 0.194439
R6647 VDD.n6284 VDD.n507 0.194439
R6648 VDD.n6284 VDD.n516 0.194439
R6649 VDD.n6297 VDD.n496 0.194439
R6650 VDD.n6297 VDD.n495 0.194439
R6651 VDD.n6306 VDD.n6305 0.194439
R6652 VDD.n6305 VDD.n494 0.194439
R6653 VDD.n6333 VDD.n6332 0.194439
R6654 VDD.n6333 VDD.n477 0.194439
R6655 VDD.n6364 VDD.n461 0.194439
R6656 VDD.n6365 VDD.n6364 0.194439
R6657 VDD.n6371 VDD.n458 0.194439
R6658 VDD.n6371 VDD.n449 0.194439
R6659 VDD.n6395 VDD.n446 0.194439
R6660 VDD.n6395 VDD.n447 0.194439
R6661 VDD.n6417 VDD.n432 0.194439
R6662 VDD.n6417 VDD.n430 0.194439
R6663 VDD.n6438 VDD.n421 0.194439
R6664 VDD.n6438 VDD.n419 0.194439
R6665 VDD.n6465 VDD.n406 0.194439
R6666 VDD.n6465 VDD.n407 0.194439
R6667 VDD.n6471 VDD.n6470 0.194439
R6668 VDD.n6471 VDD.n395 0.194439
R6669 VDD.n6491 VDD.n393 0.194439
R6670 VDD.n6491 VDD.n384 0.194439
R6671 VDD.n6510 VDD.n373 0.194439
R6672 VDD.n6510 VDD.n382 0.194439
R6673 VDD.n6523 VDD.n362 0.194439
R6674 VDD.n6523 VDD.n361 0.194439
R6675 VDD.n6532 VDD.n6531 0.194439
R6676 VDD.n6531 VDD.n360 0.194439
R6677 VDD.n6559 VDD.n6558 0.194439
R6678 VDD.n6559 VDD.n343 0.194439
R6679 VDD.n6590 VDD.n327 0.194439
R6680 VDD.n6591 VDD.n6590 0.194439
R6681 VDD.n6597 VDD.n324 0.194439
R6682 VDD.n6597 VDD.n315 0.194439
R6683 VDD.n6621 VDD.n312 0.194439
R6684 VDD.n6621 VDD.n313 0.194439
R6685 VDD.n6643 VDD.n298 0.194439
R6686 VDD.n6643 VDD.n296 0.194439
R6687 VDD.n6664 VDD.n287 0.194439
R6688 VDD.n6664 VDD.n285 0.194439
R6689 VDD.n6691 VDD.n272 0.194439
R6690 VDD.n6691 VDD.n273 0.194439
R6691 VDD.n6697 VDD.n6696 0.194439
R6692 VDD.n6697 VDD.n261 0.194439
R6693 VDD.n6717 VDD.n259 0.194439
R6694 VDD.n6717 VDD.n250 0.194439
R6695 VDD.n6736 VDD.n239 0.194439
R6696 VDD.n6736 VDD.n248 0.194439
R6697 VDD.n6749 VDD.n228 0.194439
R6698 VDD.n6749 VDD.n227 0.194439
R6699 VDD.n6758 VDD.n6757 0.194439
R6700 VDD.n6757 VDD.n226 0.194439
R6701 VDD.n6785 VDD.n6784 0.194439
R6702 VDD.n6785 VDD.n209 0.194439
R6703 VDD.n6816 VDD.n193 0.194439
R6704 VDD.n6817 VDD.n6816 0.194439
R6705 VDD.n6823 VDD.n190 0.194439
R6706 VDD.n6823 VDD.n181 0.194439
R6707 VDD.n6847 VDD.n178 0.194439
R6708 VDD.n6847 VDD.n179 0.194439
R6709 VDD.n6869 VDD.n164 0.194439
R6710 VDD.n6869 VDD.n162 0.194439
R6711 VDD.n6890 VDD.n153 0.194439
R6712 VDD.n6890 VDD.n151 0.194439
R6713 VDD.n6917 VDD.n138 0.194439
R6714 VDD.n6917 VDD.n139 0.194439
R6715 VDD.n6923 VDD.n6922 0.194439
R6716 VDD.n6923 VDD.n127 0.194439
R6717 VDD.n6943 VDD.n125 0.194439
R6718 VDD.n6943 VDD.n116 0.194439
R6719 VDD.n6962 VDD.n105 0.194439
R6720 VDD.n6962 VDD.n114 0.194439
R6721 VDD.n6975 VDD.n94 0.194439
R6722 VDD.n6975 VDD.n93 0.194439
R6723 VDD.n6984 VDD.n6983 0.194439
R6724 VDD.n6983 VDD.n92 0.194439
R6725 VDD.n7011 VDD.n7010 0.194439
R6726 VDD.n7011 VDD.n75 0.194439
R6727 VDD.n7042 VDD.n59 0.194439
R6728 VDD.n7043 VDD.n7042 0.194439
R6729 VDD.n7049 VDD.n56 0.194439
R6730 VDD.n7049 VDD.n46 0.194439
R6731 VDD.n7072 VDD.n44 0.194439
R6732 VDD.n7221 VDD.n7220 0.194439
R6733 VDD.n7216 VDD.n25 0.194439
R6734 VDD.n7216 VDD.n27 0.194439
R6735 VDD.n7115 VDD.n7113 0.194439
R6736 VDD.n7117 VDD.n7115 0.194439
R6737 VDD.n7197 VDD.n7196 0.194439
R6738 VDD.n7196 VDD.n7194 0.194439
R6739 VDD.n7162 VDD.n7120 0.194439
R6740 VDD.n7163 VDD.n7162 0.194439
R6741 VDD.n7176 VDD.n7174 0.194439
R6742 VDD.n7176 VDD.n10 0.194439
R6743 VDD.n2631 VDD.n2630 0.194439
R6744 VDD.n2631 VDD.n2451 0.194439
R6745 VDD.n4375 VDD.n2445 0.194439
R6746 VDD.n4375 VDD.n2446 0.194439
R6747 VDD.n4369 VDD.n4368 0.194439
R6748 VDD.n4368 VDD.n2645 0.194439
R6749 VDD.n2701 VDD.n2700 0.194439
R6750 VDD.n2702 VDD.n2701 0.194439
R6751 VDD.n4348 VDD.n2688 0.194439
R6752 VDD.n4348 VDD.n2689 0.194439
R6753 VDD.n4342 VDD.n4341 0.194439
R6754 VDD.n4873 VDD.n1380 0.194439
R6755 VDD.n4867 VDD.n4866 0.194439
R6756 VDD.n4866 VDD.n1398 0.194439
R6757 VDD.n1453 VDD.n1452 0.194439
R6758 VDD.n1454 VDD.n1453 0.194439
R6759 VDD.n4846 VDD.n1440 0.194439
R6760 VDD.n4846 VDD.n1441 0.194439
R6761 VDD.n4840 VDD.n4839 0.194439
R6762 VDD.n4839 VDD.n1466 0.194439
R6763 VDD.n1529 VDD.n1517 0.194439
R6764 VDD.n1529 VDD.n1528 0.194439
R6765 VDD.n4821 VDD.n1508 0.194439
R6766 VDD.n4821 VDD.n1509 0.194439
R6767 VDD.n1562 VDD.n1535 0.194439
R6768 VDD.n1571 VDD.n1562 0.194439
R6769 VDD.n4799 VDD.n1558 0.194439
R6770 VDD.n4799 VDD.n1559 0.194439
R6771 VDD.n1604 VDD.n1577 0.194439
R6772 VDD.n1613 VDD.n1604 0.194439
R6773 VDD.n4777 VDD.n1600 0.194439
R6774 VDD.n4777 VDD.n1601 0.194439
R6775 VDD.n1652 VDD.n1619 0.194439
R6776 VDD.n1653 VDD.n1652 0.194439
R6777 VDD.n4752 VDD.n1648 0.194439
R6778 VDD.n4752 VDD.n1649 0.194439
R6779 VDD.n4746 VDD.n4745 0.194439
R6780 VDD.n4745 VDD.n1666 0.194439
R6781 VDD.n1717 VDD.n1716 0.194439
R6782 VDD.n1718 VDD.n1717 0.194439
R6783 VDD.n4725 VDD.n1704 0.194439
R6784 VDD.n4725 VDD.n1705 0.194439
R6785 VDD.n4719 VDD.n4718 0.194439
R6786 VDD.n4718 VDD.n1730 0.194439
R6787 VDD.n1793 VDD.n1781 0.194439
R6788 VDD.n1793 VDD.n1792 0.194439
R6789 VDD.n4700 VDD.n1772 0.194439
R6790 VDD.n4700 VDD.n1773 0.194439
R6791 VDD.n1826 VDD.n1799 0.194439
R6792 VDD.n1835 VDD.n1826 0.194439
R6793 VDD.n4678 VDD.n1822 0.194439
R6794 VDD.n4678 VDD.n1823 0.194439
R6795 VDD.n1868 VDD.n1841 0.194439
R6796 VDD.n1877 VDD.n1868 0.194439
R6797 VDD.n4656 VDD.n1864 0.194439
R6798 VDD.n4656 VDD.n1865 0.194439
R6799 VDD.n1916 VDD.n1883 0.194439
R6800 VDD.n1917 VDD.n1916 0.194439
R6801 VDD.n4631 VDD.n1912 0.194439
R6802 VDD.n4631 VDD.n1913 0.194439
R6803 VDD.n4625 VDD.n4624 0.194439
R6804 VDD.n4624 VDD.n1930 0.194439
R6805 VDD.n1981 VDD.n1980 0.194439
R6806 VDD.n1982 VDD.n1981 0.194439
R6807 VDD.n4604 VDD.n1968 0.194439
R6808 VDD.n4604 VDD.n1969 0.194439
R6809 VDD.n4598 VDD.n4597 0.194439
R6810 VDD.n4597 VDD.n1994 0.194439
R6811 VDD.n2057 VDD.n2045 0.194439
R6812 VDD.n2057 VDD.n2056 0.194439
R6813 VDD.n4579 VDD.n2036 0.194439
R6814 VDD.n4579 VDD.n2037 0.194439
R6815 VDD.n2090 VDD.n2063 0.194439
R6816 VDD.n2099 VDD.n2090 0.194439
R6817 VDD.n4557 VDD.n2086 0.194439
R6818 VDD.n4557 VDD.n2087 0.194439
R6819 VDD.n2132 VDD.n2105 0.194439
R6820 VDD.n2141 VDD.n2132 0.194439
R6821 VDD.n4535 VDD.n2128 0.194439
R6822 VDD.n4535 VDD.n2129 0.194439
R6823 VDD.n2180 VDD.n2147 0.194439
R6824 VDD.n2181 VDD.n2180 0.194439
R6825 VDD.n4510 VDD.n2176 0.194439
R6826 VDD.n4510 VDD.n2177 0.194439
R6827 VDD.n4504 VDD.n4503 0.194439
R6828 VDD.n4503 VDD.n2194 0.194439
R6829 VDD.n2245 VDD.n2244 0.194439
R6830 VDD.n2246 VDD.n2245 0.194439
R6831 VDD.n4483 VDD.n2232 0.194439
R6832 VDD.n4483 VDD.n2233 0.194439
R6833 VDD.n4477 VDD.n4476 0.194439
R6834 VDD.n4476 VDD.n2258 0.194439
R6835 VDD.n2321 VDD.n2309 0.194439
R6836 VDD.n2321 VDD.n2320 0.194439
R6837 VDD.n4458 VDD.n2300 0.194439
R6838 VDD.n4458 VDD.n2301 0.194439
R6839 VDD.n2354 VDD.n2327 0.194439
R6840 VDD.n2363 VDD.n2354 0.194439
R6841 VDD.n4436 VDD.n2350 0.194439
R6842 VDD.n4436 VDD.n2351 0.194439
R6843 VDD.n2396 VDD.n2369 0.194439
R6844 VDD.n2405 VDD.n2396 0.194439
R6845 VDD.n4414 VDD.n2392 0.194439
R6846 VDD.n4414 VDD.n2393 0.194439
R6847 VDD.n2537 VDD.n2411 0.194439
R6848 VDD.n4926 VDD.n4925 0.194439
R6849 VDD.n4925 VDD.n1244 0.194439
R6850 VDD.n4919 VDD.n4918 0.194439
R6851 VDD.n4918 VDD.n1250 0.194439
R6852 VDD.n1326 VDD.n1325 0.194439
R6853 VDD.n1327 VDD.n1326 0.194439
R6854 VDD.n4898 VDD.n1313 0.194439
R6855 VDD.n4898 VDD.n1314 0.194439
R6856 VDD.n4892 VDD.n4891 0.194439
R6857 VDD.n4891 VDD.n1339 0.194439
R6858 VDD.n1390 VDD.n1389 0.194439
R6859 VDD.n2763 VDD.n2739 0.194439
R6860 VDD.n4322 VDD.n2753 0.194439
R6861 VDD.n4322 VDD.n2754 0.194439
R6862 VDD.n4316 VDD.n4315 0.194439
R6863 VDD.n4315 VDD.n2776 0.194439
R6864 VDD.n2827 VDD.n2826 0.194439
R6865 VDD.n2828 VDD.n2827 0.194439
R6866 VDD.n4295 VDD.n2814 0.194439
R6867 VDD.n4295 VDD.n2815 0.194439
R6868 VDD.n4289 VDD.n4288 0.194439
R6869 VDD.n4288 VDD.n2840 0.194439
R6870 VDD.n4279 VDD.n4278 0.194439
R6871 VDD.n4278 VDD.n2847 0.194439
R6872 VDD.n2914 VDD.n2853 0.194439
R6873 VDD.n2922 VDD.n2914 0.194439
R6874 VDD.n4257 VDD.n2910 0.194439
R6875 VDD.n4257 VDD.n2911 0.194439
R6876 VDD.n2957 VDD.n2928 0.194439
R6877 VDD.n2965 VDD.n2957 0.194439
R6878 VDD.n4236 VDD.n2953 0.194439
R6879 VDD.n4236 VDD.n2954 0.194439
R6880 VDD.n3004 VDD.n2971 0.194439
R6881 VDD.n3005 VDD.n3004 0.194439
R6882 VDD.n4211 VDD.n3000 0.194439
R6883 VDD.n4211 VDD.n3001 0.194439
R6884 VDD.n4205 VDD.n4204 0.194439
R6885 VDD.n4204 VDD.n3018 0.194439
R6886 VDD.n3069 VDD.n3068 0.194439
R6887 VDD.n3070 VDD.n3069 0.194439
R6888 VDD.n4184 VDD.n3056 0.194439
R6889 VDD.n4184 VDD.n3057 0.194439
R6890 VDD.n4178 VDD.n4177 0.194439
R6891 VDD.n4177 VDD.n3082 0.194439
R6892 VDD.n3145 VDD.n3133 0.194439
R6893 VDD.n3145 VDD.n3144 0.194439
R6894 VDD.n4159 VDD.n3124 0.194439
R6895 VDD.n4159 VDD.n3125 0.194439
R6896 VDD.n3180 VDD.n3151 0.194439
R6897 VDD.n3188 VDD.n3180 0.194439
R6898 VDD.n4138 VDD.n3176 0.194439
R6899 VDD.n4138 VDD.n3177 0.194439
R6900 VDD.n3223 VDD.n3194 0.194439
R6901 VDD.n3231 VDD.n3223 0.194439
R6902 VDD.n4117 VDD.n3219 0.194439
R6903 VDD.n4117 VDD.n3220 0.194439
R6904 VDD.n3270 VDD.n3237 0.194439
R6905 VDD.n3271 VDD.n3270 0.194439
R6906 VDD.n4092 VDD.n3266 0.194439
R6907 VDD.n4092 VDD.n3267 0.194439
R6908 VDD.n4086 VDD.n4085 0.194439
R6909 VDD.n4085 VDD.n3284 0.194439
R6910 VDD.n3335 VDD.n3334 0.194439
R6911 VDD.n3336 VDD.n3335 0.194439
R6912 VDD.n4065 VDD.n3322 0.194439
R6913 VDD.n4065 VDD.n3323 0.194439
R6914 VDD.n4059 VDD.n4058 0.194439
R6915 VDD.n4058 VDD.n3348 0.194439
R6916 VDD.n3411 VDD.n3399 0.194439
R6917 VDD.n3411 VDD.n3410 0.194439
R6918 VDD.n4040 VDD.n3390 0.194439
R6919 VDD.n4040 VDD.n3391 0.194439
R6920 VDD.n3446 VDD.n3417 0.194439
R6921 VDD.n3454 VDD.n3446 0.194439
R6922 VDD.n4019 VDD.n3442 0.194439
R6923 VDD.n4019 VDD.n3443 0.194439
R6924 VDD.n3489 VDD.n3460 0.194439
R6925 VDD.n3497 VDD.n3489 0.194439
R6926 VDD.n3998 VDD.n3485 0.194439
R6927 VDD.n3998 VDD.n3486 0.194439
R6928 VDD.n3536 VDD.n3503 0.194439
R6929 VDD.n3537 VDD.n3536 0.194439
R6930 VDD.n3973 VDD.n3532 0.194439
R6931 VDD.n3973 VDD.n3533 0.194439
R6932 VDD.n3967 VDD.n3966 0.194439
R6933 VDD.n3966 VDD.n3550 0.194439
R6934 VDD.n3601 VDD.n3600 0.194439
R6935 VDD.n3602 VDD.n3601 0.194439
R6936 VDD.n3946 VDD.n3588 0.194439
R6937 VDD.n3946 VDD.n3589 0.194439
R6938 VDD.n3940 VDD.n3939 0.194439
R6939 VDD.n3939 VDD.n3614 0.194439
R6940 VDD.n3677 VDD.n3665 0.194439
R6941 VDD.n3677 VDD.n3676 0.194439
R6942 VDD.n3921 VDD.n3656 0.194439
R6943 VDD.n3921 VDD.n3657 0.194439
R6944 VDD.n3712 VDD.n3683 0.194439
R6945 VDD.n3720 VDD.n3712 0.194439
R6946 VDD.n3900 VDD.n3708 0.194439
R6947 VDD.n3900 VDD.n3709 0.194439
R6948 VDD.n3755 VDD.n3726 0.194439
R6949 VDD.n3763 VDD.n3755 0.194439
R6950 VDD.n3879 VDD.n3751 0.194439
R6951 VDD.n3879 VDD.n3752 0.194439
R6952 VDD.n3820 VDD.n3769 0.194439
R6953 VDD.n5025 VDD.n1190 0.194439
R6954 VDD.n5046 VDD.n1188 0.194439
R6955 VDD.n5046 VDD.n1177 0.194439
R6956 VDD.n5071 VDD.n1175 0.194439
R6957 VDD.n1175 VDD.n1174 0.194439
R6958 VDD.n5100 VDD.n1161 0.194439
R6959 VDD.n5100 VDD.n1162 0.194439
R6960 VDD.n5107 VDD.n5106 0.194439
R6961 VDD.n5107 VDD.n1150 0.194439
R6962 VDD.n5128 VDD.n1130 0.194439
R6963 VDD.n5128 VDD.n1148 0.194439
R6964 VDD.n1140 VDD.n1139 0.194439
R6965 VDD.n1139 VDD.n1135 0.194439
R6966 VDD.n5152 VDD.n5151 0.194439
R6967 VDD.n5152 VDD.n1115 0.194439
R6968 VDD.n5183 VDD.n1099 0.194439
R6969 VDD.n5184 VDD.n5183 0.194439
R6970 VDD.n5190 VDD.n1096 0.194439
R6971 VDD.n5190 VDD.n1083 0.194439
R6972 VDD.n1084 VDD.n1081 0.194439
R6973 VDD.n5213 VDD.n1081 0.194439
R6974 VDD.n5243 VDD.n1066 0.194439
R6975 VDD.n5243 VDD.n1064 0.194439
R6976 VDD.n5253 VDD.n5252 0.194439
R6977 VDD.n5253 VDD.n1055 0.194439
R6978 VDD.n5274 VDD.n1053 0.194439
R6979 VDD.n5274 VDD.n1042 0.194439
R6980 VDD.n5299 VDD.n1040 0.194439
R6981 VDD.n1040 VDD.n1039 0.194439
R6982 VDD.n5328 VDD.n1026 0.194439
R6983 VDD.n5328 VDD.n1027 0.194439
R6984 VDD.n5335 VDD.n5334 0.194439
R6985 VDD.n5335 VDD.n1015 0.194439
R6986 VDD.n5356 VDD.n995 0.194439
R6987 VDD.n5356 VDD.n1013 0.194439
R6988 VDD.n1005 VDD.n1004 0.194439
R6989 VDD.n1004 VDD.n1000 0.194439
R6990 VDD.n5380 VDD.n5379 0.194439
R6991 VDD.n5380 VDD.n980 0.194439
R6992 VDD.n5411 VDD.n964 0.194439
R6993 VDD.n5412 VDD.n5411 0.194439
R6994 VDD.n5418 VDD.n961 0.194439
R6995 VDD.n5418 VDD.n948 0.194439
R6996 VDD.n949 VDD.n946 0.194439
R6997 VDD.n5441 VDD.n946 0.194439
R6998 VDD.n5471 VDD.n931 0.194439
R6999 VDD.n5471 VDD.n929 0.194439
R7000 VDD.n5481 VDD.n5480 0.194439
R7001 VDD.n5481 VDD.n920 0.194439
R7002 VDD.n5502 VDD.n918 0.194439
R7003 VDD.n5502 VDD.n907 0.194439
R7004 VDD.n5527 VDD.n905 0.194439
R7005 VDD.n905 VDD.n904 0.194439
R7006 VDD.n5556 VDD.n891 0.194439
R7007 VDD.n5556 VDD.n892 0.194439
R7008 VDD.n5563 VDD.n5562 0.194439
R7009 VDD.n5563 VDD.n880 0.194439
R7010 VDD.n5584 VDD.n860 0.194439
R7011 VDD.n5584 VDD.n878 0.194439
R7012 VDD.n870 VDD.n869 0.194439
R7013 VDD.n869 VDD.n865 0.194439
R7014 VDD.n5608 VDD.n5607 0.194439
R7015 VDD.n5608 VDD.n845 0.194439
R7016 VDD.n5639 VDD.n829 0.194439
R7017 VDD.n5640 VDD.n5639 0.194439
R7018 VDD.n5646 VDD.n826 0.194439
R7019 VDD.n5646 VDD.n813 0.194439
R7020 VDD.n814 VDD.n811 0.194439
R7021 VDD.n5669 VDD.n811 0.194439
R7022 VDD.n5699 VDD.n796 0.194439
R7023 VDD.n5699 VDD.n794 0.194439
R7024 VDD.n5709 VDD.n5708 0.194439
R7025 VDD.n5709 VDD.n785 0.194439
R7026 VDD.n5730 VDD.n783 0.194439
R7027 VDD.n5730 VDD.n772 0.194439
R7028 VDD.n5755 VDD.n770 0.194439
R7029 VDD.n770 VDD.n769 0.194439
R7030 VDD.n5784 VDD.n756 0.194439
R7031 VDD.n5784 VDD.n757 0.194439
R7032 VDD.n5791 VDD.n5790 0.194439
R7033 VDD.n5791 VDD.n745 0.194439
R7034 VDD.n5811 VDD.n734 0.194439
R7035 VDD.n5811 VDD.n743 0.194439
R7036 VDD.n5824 VDD.n724 0.194439
R7037 VDD.n5828 VDD.n5824 0.194439
R7038 VDD.n5846 VDD.n716 0.194439
R7039 VDD.n5846 VDD.n714 0.194439
R7040 VDD.n5854 VDD.n5853 0.194439
R7041 VDD.n5853 VDD.n711 0.194439
R7042 VDD.n5881 VDD.n5880 0.194439
R7043 VDD.n5881 VDD.n694 0.194439
R7044 VDD.n5916 VDD.n676 0.194439
R7045 VDD.n5917 VDD.n5916 0.194439
R7046 VDD.n5922 VDD.n673 0.194439
R7047 VDD.n7232 VDD 0.152702
R7048 VDD.n6078 VDD.n6077 0.132407
R7049 VDD.n7228 VDD.n7227 0.132407
R7050 VDD.n2624 VDD.n2623 0.13107
R7051 VDD.n1274 VDD.n1267 0.13107
R7052 VDD.n6078 VDD.n637 0.127283
R7053 VDD.n7228 VDD.n8 0.127283
R7054 VDD.n2623 VDD.n2452 0.127283
R7055 VDD.n1275 VDD.n1274 0.127283
R7056 VDD.n7233 VDD 0.1039
R7057 VDD.n5134 VDD.n5132 0.102103
R7058 VDD.n5362 VDD.n5360 0.102103
R7059 VDD.n5590 VDD.n5588 0.102103
R7060 VDD.n5815 VDD.n727 0.102103
R7061 VDD.n6288 VDD.n500 0.102103
R7062 VDD.n6514 VDD.n366 0.102103
R7063 VDD.n6740 VDD.n232 0.102103
R7064 VDD.n6966 VDD.n98 0.102103
R7065 VDD.n2887 VDD.n2864 0.102103
R7066 VDD.n4164 VDD.n4163 0.102103
R7067 VDD.n4045 VDD.n4044 0.102103
R7068 VDD.n3926 VDD.n3925 0.102103
R7069 VDD.n4826 VDD.n4825 0.102103
R7070 VDD.n4705 VDD.n4704 0.102103
R7071 VDD.n4584 VDD.n4583 0.102103
R7072 VDD.n4463 VDD.n4462 0.102103
R7073 VDD.n5237 VDD.n1073 0.100721
R7074 VDD.n5465 VDD.n938 0.100721
R7075 VDD.n5693 VDD.n803 0.100721
R7076 VDD.n6403 VDD.n437 0.100721
R7077 VDD.n6629 VDD.n303 0.100721
R7078 VDD.n6855 VDD.n169 0.100721
R7079 VDD.n4219 VDD.n4218 0.100721
R7080 VDD.n4100 VDD.n4099 0.100721
R7081 VDD.n3981 VDD.n3980 0.100721
R7082 VDD.n4760 VDD.n4759 0.100721
R7083 VDD.n4639 VDD.n4638 0.100721
R7084 VDD.n4518 VDD.n4517 0.100721
R7085 VDD.n6092 VDD.n6091 0.0981562
R7086 VDD.n7281 VDD.n7279 0.0981562
R7087 VDD.n2602 VDD.n2471 0.0877396
R7088 VDD.n4973 VDD.n1234 0.0877396
R7089 VDD.n7013 VDD.n7012 0.0847059
R7090 VDD.n7048 VDD.n7047 0.0847059
R7091 VDD.n6787 VDD.n6786 0.0847059
R7092 VDD.n6822 VDD.n6821 0.0847059
R7093 VDD.n6561 VDD.n6560 0.0847059
R7094 VDD.n6596 VDD.n6595 0.0847059
R7095 VDD.n6335 VDD.n6334 0.0847059
R7096 VDD.n6370 VDD.n6369 0.0847059
R7097 VDD.n6213 VDD.n554 0.0847059
R7098 VDD.n5848 VDD.n5847 0.0847059
R7099 VDD.n5883 VDD.n5882 0.0847059
R7100 VDD.n5610 VDD.n5609 0.0847059
R7101 VDD.n5645 VDD.n5644 0.0847059
R7102 VDD.n5701 VDD.n5700 0.0847059
R7103 VDD.n5382 VDD.n5381 0.0847059
R7104 VDD.n5417 VDD.n5416 0.0847059
R7105 VDD.n5473 VDD.n5472 0.0847059
R7106 VDD.n5154 VDD.n5153 0.0847059
R7107 VDD.n5189 VDD.n5188 0.0847059
R7108 VDD.n5245 VDD.n5244 0.0847059
R7109 VDD.n5788 VDD.n744 0.0847059
R7110 VDD.n5758 VDD.n5757 0.0847059
R7111 VDD.n5560 VDD.n879 0.0847059
R7112 VDD.n5530 VDD.n5529 0.0847059
R7113 VDD.n5332 VDD.n1014 0.0847059
R7114 VDD.n5302 VDD.n5301 0.0847059
R7115 VDD.n5104 VDD.n1149 0.0847059
R7116 VDD.n5074 VDD.n5073 0.0847059
R7117 VDD.n6011 VDD.n645 0.0847059
R7118 VDD.n6045 VDD.n647 0.0847059
R7119 VDD.n6067 VDD.n649 0.0847059
R7120 VDD.n5964 VDD.n643 0.0847059
R7121 VDD.n7217 VDD.n20 0.0847059
R7122 VDD.n7114 VDD.n14 0.0847059
R7123 VDD.n7195 VDD.n18 0.0847059
R7124 VDD.n7161 VDD.n16 0.0847059
R7125 VDD.n5999 VDD.n636 0.0796667
R7126 VDD.n7149 VDD.n7 0.0796667
R7127 VDD.n4389 VDD.n4388 0.0796667
R7128 VDD.n1277 VDD.n1266 0.0796667
R7129 VDD.n2562 VDD.t37 0.074533
R7130 VDD.n5037 VDD.n1187 0.0705758
R7131 VDD.n5067 VDD.n1179 0.0705758
R7132 VDD.n5080 VDD.n1163 0.0705758
R7133 VDD.n5095 VDD.n1158 0.0705758
R7134 VDD.n5120 VDD.n1128 0.0705758
R7135 VDD.n5147 VDD.n5146 0.0705758
R7136 VDD.n5164 VDD.n5163 0.0705758
R7137 VDD.n5181 VDD.n1104 0.0705758
R7138 VDD.n1095 VDD.n1085 0.0705758
R7139 VDD.n5220 VDD.n5219 0.0705758
R7140 VDD.n5265 VDD.n1052 0.0705758
R7141 VDD.n5295 VDD.n1044 0.0705758
R7142 VDD.n5308 VDD.n1028 0.0705758
R7143 VDD.n5323 VDD.n1023 0.0705758
R7144 VDD.n5348 VDD.n993 0.0705758
R7145 VDD.n5375 VDD.n5374 0.0705758
R7146 VDD.n5392 VDD.n5391 0.0705758
R7147 VDD.n5409 VDD.n969 0.0705758
R7148 VDD.n960 VDD.n950 0.0705758
R7149 VDD.n5448 VDD.n5447 0.0705758
R7150 VDD.n5493 VDD.n917 0.0705758
R7151 VDD.n5523 VDD.n909 0.0705758
R7152 VDD.n5536 VDD.n893 0.0705758
R7153 VDD.n5551 VDD.n888 0.0705758
R7154 VDD.n5576 VDD.n858 0.0705758
R7155 VDD.n5603 VDD.n5602 0.0705758
R7156 VDD.n5620 VDD.n5619 0.0705758
R7157 VDD.n5637 VDD.n834 0.0705758
R7158 VDD.n825 VDD.n815 0.0705758
R7159 VDD.n5676 VDD.n5675 0.0705758
R7160 VDD.n5721 VDD.n782 0.0705758
R7161 VDD.n5751 VDD.n774 0.0705758
R7162 VDD.n5764 VDD.n758 0.0705758
R7163 VDD.n5779 VDD.n753 0.0705758
R7164 VDD.n5803 VDD.n732 0.0705758
R7165 VDD.n5832 VDD.n723 0.0705758
R7166 VDD.n5857 VDD.n707 0.0705758
R7167 VDD.n5876 VDD.n5875 0.0705758
R7168 VDD.n5893 VDD.n5892 0.0705758
R7169 VDD.n5914 VDD.n681 0.0705758
R7170 VDD.n5937 VDD.n5936 0.0705758
R7171 VDD.n6064 VDD.n659 0.0705758
R7172 VDD.n6052 VDD.n6051 0.0705758
R7173 VDD.n5987 VDD.n5971 0.0705758
R7174 VDD.n6021 VDD.n6017 0.0705758
R7175 VDD.n6198 VDD.n556 0.0705758
R7176 VDD.n6219 VDD.n542 0.0705758
R7177 VDD.n6234 VDD.n537 0.0705758
R7178 VDD.n6257 VDD.n526 0.0705758
R7179 VDD.n6277 VDD.n505 0.0705758
R7180 VDD.n6309 VDD.n490 0.0705758
R7181 VDD.n6328 VDD.n6327 0.0705758
R7182 VDD.n6345 VDD.n6344 0.0705758
R7183 VDD.n6362 VDD.n466 0.0705758
R7184 VDD.n6383 VDD.n450 0.0705758
R7185 VDD.n6424 VDD.n422 0.0705758
R7186 VDD.n6445 VDD.n408 0.0705758
R7187 VDD.n6460 VDD.n403 0.0705758
R7188 VDD.n6483 VDD.n392 0.0705758
R7189 VDD.n6503 VDD.n371 0.0705758
R7190 VDD.n6535 VDD.n356 0.0705758
R7191 VDD.n6554 VDD.n6553 0.0705758
R7192 VDD.n6571 VDD.n6570 0.0705758
R7193 VDD.n6588 VDD.n332 0.0705758
R7194 VDD.n6609 VDD.n316 0.0705758
R7195 VDD.n6650 VDD.n288 0.0705758
R7196 VDD.n6671 VDD.n274 0.0705758
R7197 VDD.n6686 VDD.n269 0.0705758
R7198 VDD.n6709 VDD.n258 0.0705758
R7199 VDD.n6729 VDD.n237 0.0705758
R7200 VDD.n6761 VDD.n222 0.0705758
R7201 VDD.n6780 VDD.n6779 0.0705758
R7202 VDD.n6797 VDD.n6796 0.0705758
R7203 VDD.n6814 VDD.n198 0.0705758
R7204 VDD.n6835 VDD.n182 0.0705758
R7205 VDD.n6876 VDD.n154 0.0705758
R7206 VDD.n6897 VDD.n140 0.0705758
R7207 VDD.n6912 VDD.n135 0.0705758
R7208 VDD.n6935 VDD.n124 0.0705758
R7209 VDD.n6955 VDD.n103 0.0705758
R7210 VDD.n6987 VDD.n88 0.0705758
R7211 VDD.n7006 VDD.n7005 0.0705758
R7212 VDD.n7023 VDD.n7022 0.0705758
R7213 VDD.n7040 VDD.n64 0.0705758
R7214 VDD.n7066 VDD.n47 0.0705758
R7215 VDD.n7087 VDD.n7086 0.0705758
R7216 VDD.n7214 VDD.n30 0.0705758
R7217 VDD.n7202 VDD.n7201 0.0705758
R7218 VDD.n7137 VDD.n7121 0.0705758
R7219 VDD.n7171 VDD.n7167 0.0705758
R7220 VDD.n2766 VDD.n2751 0.0705758
R7221 VDD.n2791 VDD.n2777 0.0705758
R7222 VDD.n4310 VDD.n4309 0.0705758
R7223 VDD.n4297 VDD.n2811 0.0705758
R7224 VDD.n2879 VDD.n2841 0.0705758
R7225 VDD.n2896 VDD.n2854 0.0705758
R7226 VDD.n2918 VDD.n2915 0.0705758
R7227 VDD.n2929 VDD.n2909 0.0705758
R7228 VDD.n2961 VDD.n2958 0.0705758
R7229 VDD.n2972 VDD.n2952 0.0705758
R7230 VDD.n3033 VDD.n3019 0.0705758
R7231 VDD.n4199 VDD.n4198 0.0705758
R7232 VDD.n4186 VDD.n3053 0.0705758
R7233 VDD.n3102 VDD.n3083 0.0705758
R7234 VDD.n4172 VDD.n4171 0.0705758
R7235 VDD.n3152 VDD.n3123 0.0705758
R7236 VDD.n3184 VDD.n3181 0.0705758
R7237 VDD.n3195 VDD.n3175 0.0705758
R7238 VDD.n3227 VDD.n3224 0.0705758
R7239 VDD.n3238 VDD.n3218 0.0705758
R7240 VDD.n3299 VDD.n3285 0.0705758
R7241 VDD.n4080 VDD.n4079 0.0705758
R7242 VDD.n4067 VDD.n3319 0.0705758
R7243 VDD.n3368 VDD.n3349 0.0705758
R7244 VDD.n4053 VDD.n4052 0.0705758
R7245 VDD.n3418 VDD.n3389 0.0705758
R7246 VDD.n3450 VDD.n3447 0.0705758
R7247 VDD.n3461 VDD.n3441 0.0705758
R7248 VDD.n3493 VDD.n3490 0.0705758
R7249 VDD.n3504 VDD.n3484 0.0705758
R7250 VDD.n3565 VDD.n3551 0.0705758
R7251 VDD.n3961 VDD.n3960 0.0705758
R7252 VDD.n3948 VDD.n3585 0.0705758
R7253 VDD.n3634 VDD.n3615 0.0705758
R7254 VDD.n3934 VDD.n3933 0.0705758
R7255 VDD.n3684 VDD.n3655 0.0705758
R7256 VDD.n3716 VDD.n3713 0.0705758
R7257 VDD.n3727 VDD.n3707 0.0705758
R7258 VDD.n3759 VDD.n3756 0.0705758
R7259 VDD.n3770 VDD.n3750 0.0705758
R7260 VDD.n4377 VDD.n2442 0.0705758
R7261 VDD.n2665 VDD.n2646 0.0705758
R7262 VDD.n4363 VDD.n4362 0.0705758
R7263 VDD.n4350 VDD.n2685 0.0705758
R7264 VDD.n2728 VDD.n2714 0.0705758
R7265 VDD.n1417 VDD.n1399 0.0705758
R7266 VDD.n4861 VDD.n4860 0.0705758
R7267 VDD.n4848 VDD.n1437 0.0705758
R7268 VDD.n1486 VDD.n1467 0.0705758
R7269 VDD.n4834 VDD.n4833 0.0705758
R7270 VDD.n1536 VDD.n1507 0.0705758
R7271 VDD.n1567 VDD.n1563 0.0705758
R7272 VDD.n1578 VDD.n1557 0.0705758
R7273 VDD.n1609 VDD.n1605 0.0705758
R7274 VDD.n1620 VDD.n1599 0.0705758
R7275 VDD.n1681 VDD.n1667 0.0705758
R7276 VDD.n4740 VDD.n4739 0.0705758
R7277 VDD.n4727 VDD.n1701 0.0705758
R7278 VDD.n1750 VDD.n1731 0.0705758
R7279 VDD.n4713 VDD.n4712 0.0705758
R7280 VDD.n1800 VDD.n1771 0.0705758
R7281 VDD.n1831 VDD.n1827 0.0705758
R7282 VDD.n1842 VDD.n1821 0.0705758
R7283 VDD.n1873 VDD.n1869 0.0705758
R7284 VDD.n1884 VDD.n1863 0.0705758
R7285 VDD.n1945 VDD.n1931 0.0705758
R7286 VDD.n4619 VDD.n4618 0.0705758
R7287 VDD.n4606 VDD.n1965 0.0705758
R7288 VDD.n2014 VDD.n1995 0.0705758
R7289 VDD.n4592 VDD.n4591 0.0705758
R7290 VDD.n2064 VDD.n2035 0.0705758
R7291 VDD.n2095 VDD.n2091 0.0705758
R7292 VDD.n2106 VDD.n2085 0.0705758
R7293 VDD.n2137 VDD.n2133 0.0705758
R7294 VDD.n2148 VDD.n2127 0.0705758
R7295 VDD.n2209 VDD.n2195 0.0705758
R7296 VDD.n4498 VDD.n4497 0.0705758
R7297 VDD.n4485 VDD.n2229 0.0705758
R7298 VDD.n2278 VDD.n2259 0.0705758
R7299 VDD.n4471 VDD.n4470 0.0705758
R7300 VDD.n2328 VDD.n2299 0.0705758
R7301 VDD.n2359 VDD.n2355 0.0705758
R7302 VDD.n2370 VDD.n2349 0.0705758
R7303 VDD.n2401 VDD.n2397 0.0705758
R7304 VDD.n2412 VDD.n2391 0.0705758
R7305 VDD.n1290 VDD.n1251 0.0705758
R7306 VDD.n4913 VDD.n4912 0.0705758
R7307 VDD.n4900 VDD.n1310 0.0705758
R7308 VDD.n1359 VDD.n1340 0.0705758
R7309 VDD.n4886 VDD.n4885 0.0705758
R7310 VDD VDD.n4978 0.0693134
R7311 VDD.n7234 VDD 0.0680765
R7312 VDD.n4879 VDD 0.066192
R7313 VDD.n4337 VDD 0.066192
R7314 VDD.n2618 VDD.n2617 0.063
R7315 VDD.n4955 VDD.n4953 0.063
R7316 VDD.n6132 VDD.n602 0.0616979
R7317 VDD.n2603 VDD.n2602 0.0616979
R7318 VDD.n4974 VDD.n4973 0.0616979
R7319 VDD.n7256 VDD.n7250 0.0616979
R7320 VDD VDD.n602 0.0603958
R7321 VDD VDD.n2457 0.0603958
R7322 VDD VDD.n4959 0.0603958
R7323 VDD.n7250 VDD 0.0603958
R7324 VDD.n6132 VDD.n6131 0.0590938
R7325 VDD.n7256 VDD.n7255 0.0590938
R7326 VDD.n6092 VDD.n6088 0.0577917
R7327 VDD.n2617 VDD.n2457 0.0577917
R7328 VDD.n4959 VDD.n4953 0.0577917
R7329 VDD.n7283 VDD.n7281 0.0577917
R7330 VDD.n5935 VDD.n5932 0.0573182
R7331 VDD.n6062 VDD.n661 0.0573182
R7332 VDD.n6050 VDD.n5953 0.0573182
R7333 VDD.n5989 VDD.n5973 0.0573182
R7334 VDD.n6020 VDD.n6019 0.0573182
R7335 VDD.n6201 VDD.n6199 0.0573182
R7336 VDD.n6221 VDD.n6220 0.0573182
R7337 VDD.n6235 VDD.n6233 0.0573182
R7338 VDD.n6256 VDD.n6255 0.0573182
R7339 VDD.n6276 VDD.n6275 0.0573182
R7340 VDD.n6311 VDD.n6310 0.0573182
R7341 VDD.n6329 VDD.n481 0.0573182
R7342 VDD.n6343 VDD.n475 0.0573182
R7343 VDD.n6360 VDD.n468 0.0573182
R7344 VDD.n6382 VDD.n6381 0.0573182
R7345 VDD.n6427 VDD.n6425 0.0573182
R7346 VDD.n6447 VDD.n6446 0.0573182
R7347 VDD.n6461 VDD.n6459 0.0573182
R7348 VDD.n6482 VDD.n6481 0.0573182
R7349 VDD.n6502 VDD.n6501 0.0573182
R7350 VDD.n6537 VDD.n6536 0.0573182
R7351 VDD.n6555 VDD.n347 0.0573182
R7352 VDD.n6569 VDD.n341 0.0573182
R7353 VDD.n6586 VDD.n334 0.0573182
R7354 VDD.n6608 VDD.n6607 0.0573182
R7355 VDD.n6653 VDD.n6651 0.0573182
R7356 VDD.n6673 VDD.n6672 0.0573182
R7357 VDD.n6687 VDD.n6685 0.0573182
R7358 VDD.n6708 VDD.n6707 0.0573182
R7359 VDD.n6728 VDD.n6727 0.0573182
R7360 VDD.n6763 VDD.n6762 0.0573182
R7361 VDD.n6781 VDD.n213 0.0573182
R7362 VDD.n6795 VDD.n207 0.0573182
R7363 VDD.n6812 VDD.n200 0.0573182
R7364 VDD.n6834 VDD.n6833 0.0573182
R7365 VDD.n6879 VDD.n6877 0.0573182
R7366 VDD.n6899 VDD.n6898 0.0573182
R7367 VDD.n6913 VDD.n6911 0.0573182
R7368 VDD.n6934 VDD.n6933 0.0573182
R7369 VDD.n6954 VDD.n6953 0.0573182
R7370 VDD.n6989 VDD.n6988 0.0573182
R7371 VDD.n7007 VDD.n79 0.0573182
R7372 VDD.n7021 VDD.n73 0.0573182
R7373 VDD.n7038 VDD.n66 0.0573182
R7374 VDD.n7065 VDD.n7063 0.0573182
R7375 VDD.n7085 VDD.n7082 0.0573182
R7376 VDD.n7212 VDD.n32 0.0573182
R7377 VDD.n7200 VDD.n7103 0.0573182
R7378 VDD.n7139 VDD.n7123 0.0573182
R7379 VDD.n7170 VDD.n7169 0.0573182
R7380 VDD.n4379 VDD.n2440 0.0573182
R7381 VDD.n2669 VDD.n2666 0.0573182
R7382 VDD.n4364 VDD.n2649 0.0573182
R7383 VDD.n4352 VDD.n2683 0.0573182
R7384 VDD.n2731 VDD.n2729 0.0573182
R7385 VDD.n1421 VDD.n1418 0.0573182
R7386 VDD.n4862 VDD.n1402 0.0573182
R7387 VDD.n4850 VDD.n1435 0.0573182
R7388 VDD.n1490 VDD.n1487 0.0573182
R7389 VDD.n4835 VDD.n1470 0.0573182
R7390 VDD.n1546 VDD.n1538 0.0573182
R7391 VDD.n1566 VDD.n1565 0.0573182
R7392 VDD.n1588 VDD.n1580 0.0573182
R7393 VDD.n1608 VDD.n1607 0.0573182
R7394 VDD.n1630 VDD.n1622 0.0573182
R7395 VDD.n1685 VDD.n1682 0.0573182
R7396 VDD.n4741 VDD.n1670 0.0573182
R7397 VDD.n4729 VDD.n1699 0.0573182
R7398 VDD.n1754 VDD.n1751 0.0573182
R7399 VDD.n4714 VDD.n1734 0.0573182
R7400 VDD.n1810 VDD.n1802 0.0573182
R7401 VDD.n1830 VDD.n1829 0.0573182
R7402 VDD.n1852 VDD.n1844 0.0573182
R7403 VDD.n1872 VDD.n1871 0.0573182
R7404 VDD.n1894 VDD.n1886 0.0573182
R7405 VDD.n1949 VDD.n1946 0.0573182
R7406 VDD.n4620 VDD.n1934 0.0573182
R7407 VDD.n4608 VDD.n1963 0.0573182
R7408 VDD.n2018 VDD.n2015 0.0573182
R7409 VDD.n4593 VDD.n1998 0.0573182
R7410 VDD.n2074 VDD.n2066 0.0573182
R7411 VDD.n2094 VDD.n2093 0.0573182
R7412 VDD.n2116 VDD.n2108 0.0573182
R7413 VDD.n2136 VDD.n2135 0.0573182
R7414 VDD.n2158 VDD.n2150 0.0573182
R7415 VDD.n2213 VDD.n2210 0.0573182
R7416 VDD.n4499 VDD.n2198 0.0573182
R7417 VDD.n4487 VDD.n2227 0.0573182
R7418 VDD.n2282 VDD.n2279 0.0573182
R7419 VDD.n4472 VDD.n2262 0.0573182
R7420 VDD.n2338 VDD.n2330 0.0573182
R7421 VDD.n2358 VDD.n2357 0.0573182
R7422 VDD.n2380 VDD.n2372 0.0573182
R7423 VDD.n2400 VDD.n2399 0.0573182
R7424 VDD.n2422 VDD.n2414 0.0573182
R7425 VDD.n1294 VDD.n1291 0.0573182
R7426 VDD.n4914 VDD.n1254 0.0573182
R7427 VDD.n4902 VDD.n1308 0.0573182
R7428 VDD.n1363 VDD.n1360 0.0573182
R7429 VDD.n4887 VDD.n1343 0.0573182
R7430 VDD.n2765 VDD.n2764 0.0573182
R7431 VDD.n2795 VDD.n2792 0.0573182
R7432 VDD.n4311 VDD.n2780 0.0573182
R7433 VDD.n4299 VDD.n2809 0.0573182
R7434 VDD.n2881 VDD.n2880 0.0573182
R7435 VDD.n2898 VDD.n2856 0.0573182
R7436 VDD.n2917 VDD.n2916 0.0573182
R7437 VDD.n2941 VDD.n2931 0.0573182
R7438 VDD.n2960 VDD.n2959 0.0573182
R7439 VDD.n2982 VDD.n2974 0.0573182
R7440 VDD.n3037 VDD.n3034 0.0573182
R7441 VDD.n4200 VDD.n3022 0.0573182
R7442 VDD.n4188 VDD.n3051 0.0573182
R7443 VDD.n3106 VDD.n3103 0.0573182
R7444 VDD.n4173 VDD.n3086 0.0573182
R7445 VDD.n3164 VDD.n3154 0.0573182
R7446 VDD.n3183 VDD.n3182 0.0573182
R7447 VDD.n3207 VDD.n3197 0.0573182
R7448 VDD.n3226 VDD.n3225 0.0573182
R7449 VDD.n3248 VDD.n3240 0.0573182
R7450 VDD.n3303 VDD.n3300 0.0573182
R7451 VDD.n4081 VDD.n3288 0.0573182
R7452 VDD.n4069 VDD.n3317 0.0573182
R7453 VDD.n3372 VDD.n3369 0.0573182
R7454 VDD.n4054 VDD.n3352 0.0573182
R7455 VDD.n3430 VDD.n3420 0.0573182
R7456 VDD.n3449 VDD.n3448 0.0573182
R7457 VDD.n3473 VDD.n3463 0.0573182
R7458 VDD.n3492 VDD.n3491 0.0573182
R7459 VDD.n3514 VDD.n3506 0.0573182
R7460 VDD.n3569 VDD.n3566 0.0573182
R7461 VDD.n3962 VDD.n3554 0.0573182
R7462 VDD.n3950 VDD.n3583 0.0573182
R7463 VDD.n3638 VDD.n3635 0.0573182
R7464 VDD.n3935 VDD.n3618 0.0573182
R7465 VDD.n3696 VDD.n3686 0.0573182
R7466 VDD.n3715 VDD.n3714 0.0573182
R7467 VDD.n3739 VDD.n3729 0.0573182
R7468 VDD.n3758 VDD.n3757 0.0573182
R7469 VDD.n3780 VDD.n3772 0.0573182
R7470 VDD.n5036 VDD.n5035 0.0573182
R7471 VDD.n5066 VDD.n5065 0.0573182
R7472 VDD.n5082 VDD.n5081 0.0573182
R7473 VDD.n5096 VDD.n5094 0.0573182
R7474 VDD.n5119 VDD.n5118 0.0573182
R7475 VDD.n5148 VDD.n1119 0.0573182
R7476 VDD.n5162 VDD.n1113 0.0573182
R7477 VDD.n5179 VDD.n1106 0.0573182
R7478 VDD.n5202 VDD.n5201 0.0573182
R7479 VDD.n5218 VDD.n1079 0.0573182
R7480 VDD.n5264 VDD.n5263 0.0573182
R7481 VDD.n5294 VDD.n5293 0.0573182
R7482 VDD.n5310 VDD.n5309 0.0573182
R7483 VDD.n5324 VDD.n5322 0.0573182
R7484 VDD.n5347 VDD.n5346 0.0573182
R7485 VDD.n5376 VDD.n984 0.0573182
R7486 VDD.n5390 VDD.n978 0.0573182
R7487 VDD.n5407 VDD.n971 0.0573182
R7488 VDD.n5430 VDD.n5429 0.0573182
R7489 VDD.n5446 VDD.n944 0.0573182
R7490 VDD.n5492 VDD.n5491 0.0573182
R7491 VDD.n5522 VDD.n5521 0.0573182
R7492 VDD.n5538 VDD.n5537 0.0573182
R7493 VDD.n5552 VDD.n5550 0.0573182
R7494 VDD.n5575 VDD.n5574 0.0573182
R7495 VDD.n5604 VDD.n849 0.0573182
R7496 VDD.n5618 VDD.n843 0.0573182
R7497 VDD.n5635 VDD.n836 0.0573182
R7498 VDD.n5658 VDD.n5657 0.0573182
R7499 VDD.n5674 VDD.n809 0.0573182
R7500 VDD.n5720 VDD.n5719 0.0573182
R7501 VDD.n5750 VDD.n5749 0.0573182
R7502 VDD.n5766 VDD.n5765 0.0573182
R7503 VDD.n5780 VDD.n5778 0.0573182
R7504 VDD.n5802 VDD.n5801 0.0573182
R7505 VDD.n5834 VDD.n5833 0.0573182
R7506 VDD.n5859 VDD.n5858 0.0573182
R7507 VDD.n5877 VDD.n698 0.0573182
R7508 VDD.n5891 VDD.n692 0.0573182
R7509 VDD.n5912 VDD.n684 0.0573182
R7510 VDD.n4979 VDD.n1229 0.0533411
R7511 VDD.n4394 VDD.n4393 0.0533411
R7512 VDD.n6111 VDD.n613 0.0517727
R7513 VDD.n7237 VDD.n7236 0.0517727
R7514 VDD.n7233 VDD.n7232 0.0517053
R7515 VDD.n6083 VDD.n6082 0.0517053
R7516 VDD.n2614 VDD.n2460 0.0511623
R7517 VDD.n4950 VDD.n4939 0.0511623
R7518 VDD.n6079 VDD.n636 0.0455
R7519 VDD.n7229 VDD.n7 0.0455
R7520 VDD.n4389 VDD.n2429 0.0455
R7521 VDD.n1273 VDD.n1266 0.0455
R7522 VDD.n6114 VDD.n601 0.0438377
R7523 VDD.n2468 VDD.n2462 0.0438377
R7524 VDD.n4941 VDD.n4940 0.0438377
R7525 VDD.n7246 VDD.n7245 0.0438377
R7526 VDD.n5937 VDD.n652 0.0434423
R7527 VDD.n4340 VDD.n2714 0.0429349
R7528 VDD.n4885 VDD.n1344 0.0429349
R7529 VDD.n7087 VDD.n23 0.0429349
R7530 VDD.n633 VDD.n614 0.041625
R7531 VDD.n2613 VDD.n2612 0.041625
R7532 VDD.n4949 VDD.n4948 0.041625
R7533 VDD.n7242 VDD.n7241 0.041625
R7534 VDD VDD.n6180 0.0410684
R7535 VDD VDD.n5019 0.0410684
R7536 VDD.n6088 VDD 0.0408646
R7537 VDD VDD.n7283 0.0408646
R7538 VDD.n5047 VDD.n1187 0.0402727
R7539 VDD.n5060 VDD.n1179 0.0402727
R7540 VDD.n5099 VDD.n1163 0.0402727
R7541 VDD.n5108 VDD.n1158 0.0402727
R7542 VDD.n5129 VDD.n1128 0.0402727
R7543 VDD.n5146 VDD.n1120 0.0402727
R7544 VDD.n5164 VDD.n1114 0.0402727
R7545 VDD.n5182 VDD.n5181 0.0402727
R7546 VDD.n5191 VDD.n1095 0.0402727
R7547 VDD.n5220 VDD.n1080 0.0402727
R7548 VDD.n5242 VDD.n5241 0.0402727
R7549 VDD.n5254 VDD.n1063 0.0402727
R7550 VDD.n5275 VDD.n1052 0.0402727
R7551 VDD.n5288 VDD.n1044 0.0402727
R7552 VDD.n5327 VDD.n1028 0.0402727
R7553 VDD.n5336 VDD.n1023 0.0402727
R7554 VDD.n5357 VDD.n993 0.0402727
R7555 VDD.n5374 VDD.n985 0.0402727
R7556 VDD.n5392 VDD.n979 0.0402727
R7557 VDD.n5410 VDD.n5409 0.0402727
R7558 VDD.n5419 VDD.n960 0.0402727
R7559 VDD.n5448 VDD.n945 0.0402727
R7560 VDD.n5470 VDD.n5469 0.0402727
R7561 VDD.n5482 VDD.n928 0.0402727
R7562 VDD.n5503 VDD.n917 0.0402727
R7563 VDD.n5516 VDD.n909 0.0402727
R7564 VDD.n5555 VDD.n893 0.0402727
R7565 VDD.n5564 VDD.n888 0.0402727
R7566 VDD.n5585 VDD.n858 0.0402727
R7567 VDD.n5602 VDD.n850 0.0402727
R7568 VDD.n5620 VDD.n844 0.0402727
R7569 VDD.n5638 VDD.n5637 0.0402727
R7570 VDD.n5647 VDD.n825 0.0402727
R7571 VDD.n5676 VDD.n810 0.0402727
R7572 VDD.n5698 VDD.n5697 0.0402727
R7573 VDD.n5710 VDD.n793 0.0402727
R7574 VDD.n5731 VDD.n782 0.0402727
R7575 VDD.n5744 VDD.n774 0.0402727
R7576 VDD.n5783 VDD.n758 0.0402727
R7577 VDD.n5792 VDD.n753 0.0402727
R7578 VDD.n5812 VDD.n732 0.0402727
R7579 VDD.n5823 VDD.n723 0.0402727
R7580 VDD.n5845 VDD.n707 0.0402727
R7581 VDD.n5875 VDD.n699 0.0402727
R7582 VDD.n5893 VDD.n693 0.0402727
R7583 VDD.n5915 VDD.n5914 0.0402727
R7584 VDD.n6065 VDD.n6064 0.0402727
R7585 VDD.n6052 VDD.n5954 0.0402727
R7586 VDD.n5987 VDD.n5957 0.0402727
R7587 VDD.n6017 VDD.n5972 0.0402727
R7588 VDD.n6027 VDD.n637 0.0402727
R7589 VDD.n5935 VDD.n5934 0.0402727
R7590 VDD.n5961 VDD.n661 0.0402727
R7591 VDD.n6050 VDD.n6049 0.0402727
R7592 VDD.n6038 VDD.n5973 0.0402727
R7593 VDD.n6020 VDD.n5997 0.0402727
R7594 VDD.n6211 VDD.n556 0.0402727
R7595 VDD.n6238 VDD.n542 0.0402727
R7596 VDD.n6246 VDD.n537 0.0402727
R7597 VDD.n6266 VDD.n526 0.0402727
R7598 VDD.n6285 VDD.n505 0.0402727
R7599 VDD.n6296 VDD.n490 0.0402727
R7600 VDD.n6327 VDD.n482 0.0402727
R7601 VDD.n6345 VDD.n476 0.0402727
R7602 VDD.n6363 VDD.n6362 0.0402727
R7603 VDD.n6372 VDD.n450 0.0402727
R7604 VDD.n6396 VDD.n445 0.0402727
R7605 VDD.n6416 VDD.n433 0.0402727
R7606 VDD.n6437 VDD.n422 0.0402727
R7607 VDD.n6464 VDD.n408 0.0402727
R7608 VDD.n6472 VDD.n403 0.0402727
R7609 VDD.n6492 VDD.n392 0.0402727
R7610 VDD.n6511 VDD.n371 0.0402727
R7611 VDD.n6522 VDD.n356 0.0402727
R7612 VDD.n6553 VDD.n348 0.0402727
R7613 VDD.n6571 VDD.n342 0.0402727
R7614 VDD.n6589 VDD.n6588 0.0402727
R7615 VDD.n6598 VDD.n316 0.0402727
R7616 VDD.n6622 VDD.n311 0.0402727
R7617 VDD.n6642 VDD.n299 0.0402727
R7618 VDD.n6663 VDD.n288 0.0402727
R7619 VDD.n6690 VDD.n274 0.0402727
R7620 VDD.n6698 VDD.n269 0.0402727
R7621 VDD.n6718 VDD.n258 0.0402727
R7622 VDD.n6737 VDD.n237 0.0402727
R7623 VDD.n6748 VDD.n222 0.0402727
R7624 VDD.n6779 VDD.n214 0.0402727
R7625 VDD.n6797 VDD.n208 0.0402727
R7626 VDD.n6815 VDD.n6814 0.0402727
R7627 VDD.n6824 VDD.n182 0.0402727
R7628 VDD.n6848 VDD.n177 0.0402727
R7629 VDD.n6868 VDD.n165 0.0402727
R7630 VDD.n6889 VDD.n154 0.0402727
R7631 VDD.n6916 VDD.n140 0.0402727
R7632 VDD.n6924 VDD.n135 0.0402727
R7633 VDD.n6944 VDD.n124 0.0402727
R7634 VDD.n6963 VDD.n103 0.0402727
R7635 VDD.n6974 VDD.n88 0.0402727
R7636 VDD.n7005 VDD.n80 0.0402727
R7637 VDD.n7023 VDD.n74 0.0402727
R7638 VDD.n7041 VDD.n7040 0.0402727
R7639 VDD.n7050 VDD.n47 0.0402727
R7640 VDD.n6199 VDD.n562 0.0402727
R7641 VDD.n6220 VDD.n551 0.0402727
R7642 VDD.n6236 VDD.n6235 0.0402727
R7643 VDD.n6256 VDD.n531 0.0402727
R7644 VDD.n6276 VDD.n520 0.0402727
R7645 VDD.n512 VDD.n504 0.0402727
R7646 VDD.n511 VDD.n498 0.0402727
R7647 VDD.n6310 VDD.n489 0.0402727
R7648 VDD.n6330 VDD.n6329 0.0402727
R7649 VDD.n6343 VDD.n6342 0.0402727
R7650 VDD.n468 VDD.n455 0.0402727
R7651 VDD.n6382 VDD.n442 0.0402727
R7652 VDD.n6425 VDD.n428 0.0402727
R7653 VDD.n6446 VDD.n417 0.0402727
R7654 VDD.n6462 VDD.n6461 0.0402727
R7655 VDD.n6482 VDD.n397 0.0402727
R7656 VDD.n6502 VDD.n386 0.0402727
R7657 VDD.n378 VDD.n370 0.0402727
R7658 VDD.n377 VDD.n364 0.0402727
R7659 VDD.n6536 VDD.n355 0.0402727
R7660 VDD.n6556 VDD.n6555 0.0402727
R7661 VDD.n6569 VDD.n6568 0.0402727
R7662 VDD.n334 VDD.n321 0.0402727
R7663 VDD.n6608 VDD.n308 0.0402727
R7664 VDD.n6651 VDD.n294 0.0402727
R7665 VDD.n6672 VDD.n283 0.0402727
R7666 VDD.n6688 VDD.n6687 0.0402727
R7667 VDD.n6708 VDD.n263 0.0402727
R7668 VDD.n6728 VDD.n252 0.0402727
R7669 VDD.n244 VDD.n236 0.0402727
R7670 VDD.n243 VDD.n230 0.0402727
R7671 VDD.n6762 VDD.n221 0.0402727
R7672 VDD.n6782 VDD.n6781 0.0402727
R7673 VDD.n6795 VDD.n6794 0.0402727
R7674 VDD.n200 VDD.n187 0.0402727
R7675 VDD.n6834 VDD.n174 0.0402727
R7676 VDD.n6877 VDD.n160 0.0402727
R7677 VDD.n6898 VDD.n149 0.0402727
R7678 VDD.n6914 VDD.n6913 0.0402727
R7679 VDD.n6934 VDD.n129 0.0402727
R7680 VDD.n6954 VDD.n118 0.0402727
R7681 VDD.n110 VDD.n102 0.0402727
R7682 VDD.n109 VDD.n96 0.0402727
R7683 VDD.n6988 VDD.n87 0.0402727
R7684 VDD.n7008 VDD.n7007 0.0402727
R7685 VDD.n7021 VDD.n7020 0.0402727
R7686 VDD.n66 VDD.n53 0.0402727
R7687 VDD.n7065 VDD.n7064 0.0402727
R7688 VDD.n7215 VDD.n7214 0.0402727
R7689 VDD.n7202 VDD.n7104 0.0402727
R7690 VDD.n7137 VDD.n7107 0.0402727
R7691 VDD.n7167 VDD.n7122 0.0402727
R7692 VDD.n7177 VDD.n8 0.0402727
R7693 VDD.n7085 VDD.n7084 0.0402727
R7694 VDD.n7111 VDD.n32 0.0402727
R7695 VDD.n7200 VDD.n7199 0.0402727
R7696 VDD.n7188 VDD.n7123 0.0402727
R7697 VDD.n7170 VDD.n7147 0.0402727
R7698 VDD.n4323 VDD.n2751 0.0402727
R7699 VDD.n4314 VDD.n2777 0.0402727
R7700 VDD.n4309 VDD.n2781 0.0402727
R7701 VDD.n4297 VDD.n4296 0.0402727
R7702 VDD.n4287 VDD.n2841 0.0402727
R7703 VDD.n2896 VDD.n2848 0.0402727
R7704 VDD.n2915 VDD.n2855 0.0402727
R7705 VDD.n4258 VDD.n2909 0.0402727
R7706 VDD.n2958 VDD.n2930 0.0402727
R7707 VDD.n4237 VDD.n2952 0.0402727
R7708 VDD.n2997 VDD.n2973 0.0402727
R7709 VDD.n4212 VDD.n2998 0.0402727
R7710 VDD.n4203 VDD.n3019 0.0402727
R7711 VDD.n4198 VDD.n3023 0.0402727
R7712 VDD.n4186 VDD.n4185 0.0402727
R7713 VDD.n4176 VDD.n3083 0.0402727
R7714 VDD.n4171 VDD.n3087 0.0402727
R7715 VDD.n4160 VDD.n3123 0.0402727
R7716 VDD.n3181 VDD.n3153 0.0402727
R7717 VDD.n4139 VDD.n3175 0.0402727
R7718 VDD.n3224 VDD.n3196 0.0402727
R7719 VDD.n4118 VDD.n3218 0.0402727
R7720 VDD.n3263 VDD.n3239 0.0402727
R7721 VDD.n4093 VDD.n3264 0.0402727
R7722 VDD.n4084 VDD.n3285 0.0402727
R7723 VDD.n4079 VDD.n3289 0.0402727
R7724 VDD.n4067 VDD.n4066 0.0402727
R7725 VDD.n4057 VDD.n3349 0.0402727
R7726 VDD.n4052 VDD.n3353 0.0402727
R7727 VDD.n4041 VDD.n3389 0.0402727
R7728 VDD.n3447 VDD.n3419 0.0402727
R7729 VDD.n4020 VDD.n3441 0.0402727
R7730 VDD.n3490 VDD.n3462 0.0402727
R7731 VDD.n3999 VDD.n3484 0.0402727
R7732 VDD.n3529 VDD.n3505 0.0402727
R7733 VDD.n3974 VDD.n3530 0.0402727
R7734 VDD.n3965 VDD.n3551 0.0402727
R7735 VDD.n3960 VDD.n3555 0.0402727
R7736 VDD.n3948 VDD.n3947 0.0402727
R7737 VDD.n3938 VDD.n3615 0.0402727
R7738 VDD.n3933 VDD.n3619 0.0402727
R7739 VDD.n3922 VDD.n3655 0.0402727
R7740 VDD.n3713 VDD.n3685 0.0402727
R7741 VDD.n3901 VDD.n3707 0.0402727
R7742 VDD.n3756 VDD.n3728 0.0402727
R7743 VDD.n3880 VDD.n3750 0.0402727
R7744 VDD.n2632 VDD.n2452 0.0402727
R7745 VDD.n4377 VDD.n4376 0.0402727
R7746 VDD.n4367 VDD.n2646 0.0402727
R7747 VDD.n4362 VDD.n2650 0.0402727
R7748 VDD.n4350 VDD.n4349 0.0402727
R7749 VDD.n2634 VDD.n2440 0.0402727
R7750 VDD.n2666 VDD.n2662 0.0402727
R7751 VDD.n4365 VDD.n4364 0.0402727
R7752 VDD.n2703 VDD.n2683 0.0402727
R7753 VDD.n2729 VDD.n2725 0.0402727
R7754 VDD.n4865 VDD.n1399 0.0402727
R7755 VDD.n4860 VDD.n1403 0.0402727
R7756 VDD.n4848 VDD.n4847 0.0402727
R7757 VDD.n4838 VDD.n1467 0.0402727
R7758 VDD.n4833 VDD.n1471 0.0402727
R7759 VDD.n4822 VDD.n1507 0.0402727
R7760 VDD.n1563 VDD.n1537 0.0402727
R7761 VDD.n4800 VDD.n1557 0.0402727
R7762 VDD.n1605 VDD.n1579 0.0402727
R7763 VDD.n4778 VDD.n1599 0.0402727
R7764 VDD.n1645 VDD.n1621 0.0402727
R7765 VDD.n4753 VDD.n1646 0.0402727
R7766 VDD.n4744 VDD.n1667 0.0402727
R7767 VDD.n4739 VDD.n1671 0.0402727
R7768 VDD.n4727 VDD.n4726 0.0402727
R7769 VDD.n4717 VDD.n1731 0.0402727
R7770 VDD.n4712 VDD.n1735 0.0402727
R7771 VDD.n4701 VDD.n1771 0.0402727
R7772 VDD.n1827 VDD.n1801 0.0402727
R7773 VDD.n4679 VDD.n1821 0.0402727
R7774 VDD.n1869 VDD.n1843 0.0402727
R7775 VDD.n4657 VDD.n1863 0.0402727
R7776 VDD.n1909 VDD.n1885 0.0402727
R7777 VDD.n4632 VDD.n1910 0.0402727
R7778 VDD.n4623 VDD.n1931 0.0402727
R7779 VDD.n4618 VDD.n1935 0.0402727
R7780 VDD.n4606 VDD.n4605 0.0402727
R7781 VDD.n4596 VDD.n1995 0.0402727
R7782 VDD.n4591 VDD.n1999 0.0402727
R7783 VDD.n4580 VDD.n2035 0.0402727
R7784 VDD.n2091 VDD.n2065 0.0402727
R7785 VDD.n4558 VDD.n2085 0.0402727
R7786 VDD.n2133 VDD.n2107 0.0402727
R7787 VDD.n4536 VDD.n2127 0.0402727
R7788 VDD.n2173 VDD.n2149 0.0402727
R7789 VDD.n4511 VDD.n2174 0.0402727
R7790 VDD.n4502 VDD.n2195 0.0402727
R7791 VDD.n4497 VDD.n2199 0.0402727
R7792 VDD.n4485 VDD.n4484 0.0402727
R7793 VDD.n4475 VDD.n2259 0.0402727
R7794 VDD.n4470 VDD.n2263 0.0402727
R7795 VDD.n4459 VDD.n2299 0.0402727
R7796 VDD.n2355 VDD.n2329 0.0402727
R7797 VDD.n4437 VDD.n2349 0.0402727
R7798 VDD.n2397 VDD.n2371 0.0402727
R7799 VDD.n4415 VDD.n2391 0.0402727
R7800 VDD.n1418 VDD.n1414 0.0402727
R7801 VDD.n4863 VDD.n4862 0.0402727
R7802 VDD.n1455 VDD.n1435 0.0402727
R7803 VDD.n1487 VDD.n1483 0.0402727
R7804 VDD.n4836 VDD.n4835 0.0402727
R7805 VDD.n1526 VDD.n1525 0.0402727
R7806 VDD.n1520 VDD.n1504 0.0402727
R7807 VDD.n4811 VDD.n1538 0.0402727
R7808 VDD.n1566 VDD.n1554 0.0402727
R7809 VDD.n4789 VDD.n1580 0.0402727
R7810 VDD.n1608 VDD.n1596 0.0402727
R7811 VDD.n4767 VDD.n1622 0.0402727
R7812 VDD.n1682 VDD.n1640 0.0402727
R7813 VDD.n4742 VDD.n4741 0.0402727
R7814 VDD.n1719 VDD.n1699 0.0402727
R7815 VDD.n1751 VDD.n1747 0.0402727
R7816 VDD.n4715 VDD.n4714 0.0402727
R7817 VDD.n1790 VDD.n1789 0.0402727
R7818 VDD.n1784 VDD.n1768 0.0402727
R7819 VDD.n4690 VDD.n1802 0.0402727
R7820 VDD.n1830 VDD.n1818 0.0402727
R7821 VDD.n4668 VDD.n1844 0.0402727
R7822 VDD.n1872 VDD.n1860 0.0402727
R7823 VDD.n4646 VDD.n1886 0.0402727
R7824 VDD.n1946 VDD.n1904 0.0402727
R7825 VDD.n4621 VDD.n4620 0.0402727
R7826 VDD.n1983 VDD.n1963 0.0402727
R7827 VDD.n2015 VDD.n2011 0.0402727
R7828 VDD.n4594 VDD.n4593 0.0402727
R7829 VDD.n2054 VDD.n2053 0.0402727
R7830 VDD.n2048 VDD.n2032 0.0402727
R7831 VDD.n4569 VDD.n2066 0.0402727
R7832 VDD.n2094 VDD.n2082 0.0402727
R7833 VDD.n4547 VDD.n2108 0.0402727
R7834 VDD.n2136 VDD.n2124 0.0402727
R7835 VDD.n4525 VDD.n2150 0.0402727
R7836 VDD.n2210 VDD.n2168 0.0402727
R7837 VDD.n4500 VDD.n4499 0.0402727
R7838 VDD.n2247 VDD.n2227 0.0402727
R7839 VDD.n2279 VDD.n2275 0.0402727
R7840 VDD.n4473 VDD.n4472 0.0402727
R7841 VDD.n2318 VDD.n2317 0.0402727
R7842 VDD.n2312 VDD.n2296 0.0402727
R7843 VDD.n4448 VDD.n2330 0.0402727
R7844 VDD.n2358 VDD.n2346 0.0402727
R7845 VDD.n4426 VDD.n2372 0.0402727
R7846 VDD.n2400 VDD.n2388 0.0402727
R7847 VDD.n4404 VDD.n2414 0.0402727
R7848 VDD.n1275 VDD.n1245 0.0402727
R7849 VDD.n4917 VDD.n1251 0.0402727
R7850 VDD.n4912 VDD.n1255 0.0402727
R7851 VDD.n4900 VDD.n4899 0.0402727
R7852 VDD.n4890 VDD.n1340 0.0402727
R7853 VDD.n1291 VDD.n1286 0.0402727
R7854 VDD.n4915 VDD.n4914 0.0402727
R7855 VDD.n1328 VDD.n1308 0.0402727
R7856 VDD.n1360 VDD.n1356 0.0402727
R7857 VDD.n4888 VDD.n4887 0.0402727
R7858 VDD.n2765 VDD.n2741 0.0402727
R7859 VDD.n2792 VDD.n2749 0.0402727
R7860 VDD.n4312 VDD.n4311 0.0402727
R7861 VDD.n2829 VDD.n2809 0.0402727
R7862 VDD.n2880 VDD.n2876 0.0402727
R7863 VDD.n4285 VDD.n4284 0.0402727
R7864 VDD.n2863 VDD.n2844 0.0402727
R7865 VDD.n4268 VDD.n2856 0.0402727
R7866 VDD.n2917 VDD.n2906 0.0402727
R7867 VDD.n4247 VDD.n2931 0.0402727
R7868 VDD.n2960 VDD.n2949 0.0402727
R7869 VDD.n4226 VDD.n2974 0.0402727
R7870 VDD.n3034 VDD.n2993 0.0402727
R7871 VDD.n4201 VDD.n4200 0.0402727
R7872 VDD.n3071 VDD.n3051 0.0402727
R7873 VDD.n3103 VDD.n3099 0.0402727
R7874 VDD.n4174 VDD.n4173 0.0402727
R7875 VDD.n3142 VDD.n3141 0.0402727
R7876 VDD.n3136 VDD.n3120 0.0402727
R7877 VDD.n4149 VDD.n3154 0.0402727
R7878 VDD.n3183 VDD.n3172 0.0402727
R7879 VDD.n4128 VDD.n3197 0.0402727
R7880 VDD.n3226 VDD.n3215 0.0402727
R7881 VDD.n4107 VDD.n3240 0.0402727
R7882 VDD.n3300 VDD.n3259 0.0402727
R7883 VDD.n4082 VDD.n4081 0.0402727
R7884 VDD.n3337 VDD.n3317 0.0402727
R7885 VDD.n3369 VDD.n3365 0.0402727
R7886 VDD.n4055 VDD.n4054 0.0402727
R7887 VDD.n3408 VDD.n3407 0.0402727
R7888 VDD.n3402 VDD.n3386 0.0402727
R7889 VDD.n4030 VDD.n3420 0.0402727
R7890 VDD.n3449 VDD.n3438 0.0402727
R7891 VDD.n4009 VDD.n3463 0.0402727
R7892 VDD.n3492 VDD.n3481 0.0402727
R7893 VDD.n3988 VDD.n3506 0.0402727
R7894 VDD.n3566 VDD.n3525 0.0402727
R7895 VDD.n3963 VDD.n3962 0.0402727
R7896 VDD.n3603 VDD.n3583 0.0402727
R7897 VDD.n3635 VDD.n3631 0.0402727
R7898 VDD.n3936 VDD.n3935 0.0402727
R7899 VDD.n3674 VDD.n3673 0.0402727
R7900 VDD.n3668 VDD.n3652 0.0402727
R7901 VDD.n3911 VDD.n3686 0.0402727
R7902 VDD.n3715 VDD.n3704 0.0402727
R7903 VDD.n3890 VDD.n3729 0.0402727
R7904 VDD.n3758 VDD.n3747 0.0402727
R7905 VDD.n3869 VDD.n3772 0.0402727
R7906 VDD.n5036 VDD.n1192 0.0402727
R7907 VDD.n5066 VDD.n1180 0.0402727
R7908 VDD.n5081 VDD.n1172 0.0402727
R7909 VDD.n5097 VDD.n5096 0.0402727
R7910 VDD.n5119 VDD.n1152 0.0402727
R7911 VDD.n1144 VDD.n1127 0.0402727
R7912 VDD.n1143 VDD.n1142 0.0402727
R7913 VDD.n5149 VDD.n5148 0.0402727
R7914 VDD.n5162 VDD.n5161 0.0402727
R7915 VDD.n1106 VDD.n1092 0.0402727
R7916 VDD.n5203 VDD.n5202 0.0402727
R7917 VDD.n5218 VDD.n5217 0.0402727
R7918 VDD.n5264 VDD.n1057 0.0402727
R7919 VDD.n5294 VDD.n1045 0.0402727
R7920 VDD.n5309 VDD.n1037 0.0402727
R7921 VDD.n5325 VDD.n5324 0.0402727
R7922 VDD.n5347 VDD.n1017 0.0402727
R7923 VDD.n1009 VDD.n992 0.0402727
R7924 VDD.n1008 VDD.n1007 0.0402727
R7925 VDD.n5377 VDD.n5376 0.0402727
R7926 VDD.n5390 VDD.n5389 0.0402727
R7927 VDD.n971 VDD.n957 0.0402727
R7928 VDD.n5431 VDD.n5430 0.0402727
R7929 VDD.n5446 VDD.n5445 0.0402727
R7930 VDD.n5492 VDD.n922 0.0402727
R7931 VDD.n5522 VDD.n910 0.0402727
R7932 VDD.n5537 VDD.n902 0.0402727
R7933 VDD.n5553 VDD.n5552 0.0402727
R7934 VDD.n5575 VDD.n882 0.0402727
R7935 VDD.n874 VDD.n857 0.0402727
R7936 VDD.n873 VDD.n872 0.0402727
R7937 VDD.n5605 VDD.n5604 0.0402727
R7938 VDD.n5618 VDD.n5617 0.0402727
R7939 VDD.n836 VDD.n822 0.0402727
R7940 VDD.n5659 VDD.n5658 0.0402727
R7941 VDD.n5674 VDD.n5673 0.0402727
R7942 VDD.n5720 VDD.n787 0.0402727
R7943 VDD.n5750 VDD.n775 0.0402727
R7944 VDD.n5765 VDD.n767 0.0402727
R7945 VDD.n5781 VDD.n5780 0.0402727
R7946 VDD.n5802 VDD.n747 0.0402727
R7947 VDD.n739 VDD.n731 0.0402727
R7948 VDD.n738 VDD.n726 0.0402727
R7949 VDD.n5833 VDD.n718 0.0402727
R7950 VDD.n5858 VDD.n706 0.0402727
R7951 VDD.n5878 VDD.n5877 0.0402727
R7952 VDD.n5891 VDD.n5890 0.0402727
R7953 VDD.n684 VDD.n683 0.0402727
R7954 VDD.n2603 VDD 0.0369583
R7955 VDD.n2478 VDD 0.0369583
R7956 VDD.n4974 VDD 0.0369583
R7957 VDD.n4960 VDD 0.0369583
R7958 VDD.n6290 VDD.n6289 0.0368632
R7959 VDD.n6516 VDD.n6515 0.0368632
R7960 VDD.n6742 VDD.n6741 0.0368632
R7961 VDD.n6968 VDD.n6967 0.0368632
R7962 VDD.n5135 VDD.n1124 0.0368632
R7963 VDD.n5363 VDD.n989 0.0368632
R7964 VDD.n5591 VDD.n854 0.0368632
R7965 VDD.n5817 VDD.n5816 0.0368632
R7966 VDD.n5939 VDD.n5938 0.0364848
R7967 VDD.n6063 VDD.n660 0.0364848
R7968 VDD.n6054 VDD.n6053 0.0364848
R7969 VDD.n5988 VDD.n5986 0.0364848
R7970 VDD.n6018 VDD.n5974 0.0364848
R7971 VDD.n6009 VDD.n5998 0.0364848
R7972 VDD.n566 VDD.n565 0.0364848
R7973 VDD.n6200 VDD.n557 0.0364848
R7974 VDD.n6223 VDD.n6222 0.0364848
R7975 VDD.n546 VDD.n536 0.0364848
R7976 VDD.n532 VDD.n525 0.0364848
R7977 VDD.n521 VDD.n503 0.0364848
R7978 VDD.n499 VDD.n488 0.0364848
R7979 VDD.n6326 VDD.n6325 0.0364848
R7980 VDD.n6347 VDD.n6346 0.0364848
R7981 VDD.n6361 VDD.n467 0.0364848
R7982 VDD.n456 VDD.n451 0.0364848
R7983 VDD.n443 VDD.n438 0.0364848
R7984 VDD.n6406 VDD.n434 0.0364848
R7985 VDD.n6426 VDD.n423 0.0364848
R7986 VDD.n6449 VDD.n6448 0.0364848
R7987 VDD.n412 VDD.n402 0.0364848
R7988 VDD.n398 VDD.n391 0.0364848
R7989 VDD.n387 VDD.n369 0.0364848
R7990 VDD.n365 VDD.n354 0.0364848
R7991 VDD.n6552 VDD.n6551 0.0364848
R7992 VDD.n6573 VDD.n6572 0.0364848
R7993 VDD.n6587 VDD.n333 0.0364848
R7994 VDD.n322 VDD.n317 0.0364848
R7995 VDD.n309 VDD.n304 0.0364848
R7996 VDD.n6632 VDD.n300 0.0364848
R7997 VDD.n6652 VDD.n289 0.0364848
R7998 VDD.n6675 VDD.n6674 0.0364848
R7999 VDD.n278 VDD.n268 0.0364848
R8000 VDD.n264 VDD.n257 0.0364848
R8001 VDD.n253 VDD.n235 0.0364848
R8002 VDD.n231 VDD.n220 0.0364848
R8003 VDD.n6778 VDD.n6777 0.0364848
R8004 VDD.n6799 VDD.n6798 0.0364848
R8005 VDD.n6813 VDD.n199 0.0364848
R8006 VDD.n188 VDD.n183 0.0364848
R8007 VDD.n175 VDD.n170 0.0364848
R8008 VDD.n6858 VDD.n166 0.0364848
R8009 VDD.n6878 VDD.n155 0.0364848
R8010 VDD.n6901 VDD.n6900 0.0364848
R8011 VDD.n144 VDD.n134 0.0364848
R8012 VDD.n130 VDD.n123 0.0364848
R8013 VDD.n119 VDD.n101 0.0364848
R8014 VDD.n97 VDD.n86 0.0364848
R8015 VDD.n7004 VDD.n7003 0.0364848
R8016 VDD.n7025 VDD.n7024 0.0364848
R8017 VDD.n7039 VDD.n65 0.0364848
R8018 VDD.n54 VDD.n48 0.0364848
R8019 VDD.n7074 VDD.n41 0.0364848
R8020 VDD.n7089 VDD.n7088 0.0364848
R8021 VDD.n7213 VDD.n31 0.0364848
R8022 VDD.n7204 VDD.n7203 0.0364848
R8023 VDD.n7138 VDD.n7136 0.0364848
R8024 VDD.n7168 VDD.n7124 0.0364848
R8025 VDD.n7159 VDD.n7148 0.0364848
R8026 VDD.n2434 VDD.n2431 0.0364848
R8027 VDD.n4378 VDD.n2441 0.0364848
R8028 VDD.n2668 VDD.n2667 0.0364848
R8029 VDD.n4361 VDD.n4360 0.0364848
R8030 VDD.n4351 VDD.n2684 0.0364848
R8031 VDD.n2730 VDD.n2715 0.0364848
R8032 VDD.n4875 VDD.n1376 0.0364848
R8033 VDD.n1420 VDD.n1419 0.0364848
R8034 VDD.n4859 VDD.n4858 0.0364848
R8035 VDD.n4849 VDD.n1436 0.0364848
R8036 VDD.n1489 VDD.n1488 0.0364848
R8037 VDD.n4832 VDD.n4831 0.0364848
R8038 VDD.n1545 VDD.n1505 0.0364848
R8039 VDD.n1564 VDD.n1539 0.0364848
R8040 VDD.n1587 VDD.n1555 0.0364848
R8041 VDD.n1606 VDD.n1581 0.0364848
R8042 VDD.n1629 VDD.n1597 0.0364848
R8043 VDD.n1644 VDD.n1623 0.0364848
R8044 VDD.n4755 VDD.n1639 0.0364848
R8045 VDD.n1684 VDD.n1683 0.0364848
R8046 VDD.n4738 VDD.n4737 0.0364848
R8047 VDD.n4728 VDD.n1700 0.0364848
R8048 VDD.n1753 VDD.n1752 0.0364848
R8049 VDD.n4711 VDD.n4710 0.0364848
R8050 VDD.n1809 VDD.n1769 0.0364848
R8051 VDD.n1828 VDD.n1803 0.0364848
R8052 VDD.n1851 VDD.n1819 0.0364848
R8053 VDD.n1870 VDD.n1845 0.0364848
R8054 VDD.n1893 VDD.n1861 0.0364848
R8055 VDD.n1908 VDD.n1887 0.0364848
R8056 VDD.n4634 VDD.n1903 0.0364848
R8057 VDD.n1948 VDD.n1947 0.0364848
R8058 VDD.n4617 VDD.n4616 0.0364848
R8059 VDD.n4607 VDD.n1964 0.0364848
R8060 VDD.n2017 VDD.n2016 0.0364848
R8061 VDD.n4590 VDD.n4589 0.0364848
R8062 VDD.n2073 VDD.n2033 0.0364848
R8063 VDD.n2092 VDD.n2067 0.0364848
R8064 VDD.n2115 VDD.n2083 0.0364848
R8065 VDD.n2134 VDD.n2109 0.0364848
R8066 VDD.n2157 VDD.n2125 0.0364848
R8067 VDD.n2172 VDD.n2151 0.0364848
R8068 VDD.n4513 VDD.n2167 0.0364848
R8069 VDD.n2212 VDD.n2211 0.0364848
R8070 VDD.n4496 VDD.n4495 0.0364848
R8071 VDD.n4486 VDD.n2228 0.0364848
R8072 VDD.n2281 VDD.n2280 0.0364848
R8073 VDD.n4469 VDD.n4468 0.0364848
R8074 VDD.n2337 VDD.n2297 0.0364848
R8075 VDD.n2356 VDD.n2331 0.0364848
R8076 VDD.n2379 VDD.n2347 0.0364848
R8077 VDD.n2398 VDD.n2373 0.0364848
R8078 VDD.n2421 VDD.n2389 0.0364848
R8079 VDD.n4396 VDD.n2415 0.0364848
R8080 VDD.n1276 VDD.n1263 0.0364848
R8081 VDD.n1293 VDD.n1292 0.0364848
R8082 VDD.n4911 VDD.n4910 0.0364848
R8083 VDD.n4901 VDD.n1309 0.0364848
R8084 VDD.n1362 VDD.n1361 0.0364848
R8085 VDD.n4884 VDD.n4883 0.0364848
R8086 VDD.n4334 VDD.n2738 0.0364848
R8087 VDD.n4325 VDD.n2748 0.0364848
R8088 VDD.n2794 VDD.n2793 0.0364848
R8089 VDD.n4308 VDD.n4307 0.0364848
R8090 VDD.n4298 VDD.n2810 0.0364848
R8091 VDD.n2883 VDD.n2882 0.0364848
R8092 VDD.n2897 VDD.n2895 0.0364848
R8093 VDD.n4266 VDD.n2858 0.0364848
R8094 VDD.n2940 VDD.n2907 0.0364848
R8095 VDD.n4245 VDD.n2933 0.0364848
R8096 VDD.n2981 VDD.n2950 0.0364848
R8097 VDD.n2996 VDD.n2975 0.0364848
R8098 VDD.n4214 VDD.n2991 0.0364848
R8099 VDD.n3036 VDD.n3035 0.0364848
R8100 VDD.n4197 VDD.n4196 0.0364848
R8101 VDD.n4187 VDD.n3052 0.0364848
R8102 VDD.n3105 VDD.n3104 0.0364848
R8103 VDD.n4170 VDD.n4169 0.0364848
R8104 VDD.n3163 VDD.n3121 0.0364848
R8105 VDD.n4147 VDD.n3156 0.0364848
R8106 VDD.n3206 VDD.n3173 0.0364848
R8107 VDD.n4126 VDD.n3199 0.0364848
R8108 VDD.n3247 VDD.n3216 0.0364848
R8109 VDD.n3262 VDD.n3241 0.0364848
R8110 VDD.n4095 VDD.n3257 0.0364848
R8111 VDD.n3302 VDD.n3301 0.0364848
R8112 VDD.n4078 VDD.n4077 0.0364848
R8113 VDD.n4068 VDD.n3318 0.0364848
R8114 VDD.n3371 VDD.n3370 0.0364848
R8115 VDD.n4051 VDD.n4050 0.0364848
R8116 VDD.n3429 VDD.n3387 0.0364848
R8117 VDD.n4028 VDD.n3422 0.0364848
R8118 VDD.n3472 VDD.n3439 0.0364848
R8119 VDD.n4007 VDD.n3465 0.0364848
R8120 VDD.n3513 VDD.n3482 0.0364848
R8121 VDD.n3528 VDD.n3507 0.0364848
R8122 VDD.n3976 VDD.n3523 0.0364848
R8123 VDD.n3568 VDD.n3567 0.0364848
R8124 VDD.n3959 VDD.n3958 0.0364848
R8125 VDD.n3949 VDD.n3584 0.0364848
R8126 VDD.n3637 VDD.n3636 0.0364848
R8127 VDD.n3932 VDD.n3931 0.0364848
R8128 VDD.n3695 VDD.n3653 0.0364848
R8129 VDD.n3909 VDD.n3688 0.0364848
R8130 VDD.n3738 VDD.n3705 0.0364848
R8131 VDD.n3888 VDD.n3731 0.0364848
R8132 VDD.n3779 VDD.n3748 0.0364848
R8133 VDD.n3861 VDD.n3773 0.0364848
R8134 VDD.n5024 VDD.n1197 0.0364848
R8135 VDD.n1193 VDD.n1186 0.0364848
R8136 VDD.n5062 VDD.n1181 0.0364848
R8137 VDD.n5084 VDD.n5083 0.0364848
R8138 VDD.n1167 VDD.n1157 0.0364848
R8139 VDD.n1153 VDD.n1126 0.0364848
R8140 VDD.n5145 VDD.n5144 0.0364848
R8141 VDD.n5166 VDD.n5165 0.0364848
R8142 VDD.n5180 VDD.n1105 0.0364848
R8143 VDD.n1093 VDD.n1086 0.0364848
R8144 VDD.n5222 VDD.n5221 0.0364848
R8145 VDD.n5240 VDD.n1069 0.0364848
R8146 VDD.n1070 VDD.n1062 0.0364848
R8147 VDD.n1058 VDD.n1051 0.0364848
R8148 VDD.n5290 VDD.n1046 0.0364848
R8149 VDD.n5312 VDD.n5311 0.0364848
R8150 VDD.n1032 VDD.n1022 0.0364848
R8151 VDD.n1018 VDD.n991 0.0364848
R8152 VDD.n5373 VDD.n5372 0.0364848
R8153 VDD.n5394 VDD.n5393 0.0364848
R8154 VDD.n5408 VDD.n970 0.0364848
R8155 VDD.n958 VDD.n951 0.0364848
R8156 VDD.n5450 VDD.n5449 0.0364848
R8157 VDD.n5468 VDD.n934 0.0364848
R8158 VDD.n935 VDD.n927 0.0364848
R8159 VDD.n923 VDD.n916 0.0364848
R8160 VDD.n5518 VDD.n911 0.0364848
R8161 VDD.n5540 VDD.n5539 0.0364848
R8162 VDD.n897 VDD.n887 0.0364848
R8163 VDD.n883 VDD.n856 0.0364848
R8164 VDD.n5601 VDD.n5600 0.0364848
R8165 VDD.n5622 VDD.n5621 0.0364848
R8166 VDD.n5636 VDD.n835 0.0364848
R8167 VDD.n823 VDD.n816 0.0364848
R8168 VDD.n5678 VDD.n5677 0.0364848
R8169 VDD.n5696 VDD.n799 0.0364848
R8170 VDD.n800 VDD.n792 0.0364848
R8171 VDD.n788 VDD.n781 0.0364848
R8172 VDD.n5746 VDD.n776 0.0364848
R8173 VDD.n5768 VDD.n5767 0.0364848
R8174 VDD.n762 VDD.n752 0.0364848
R8175 VDD.n748 VDD.n730 0.0364848
R8176 VDD.n5821 VDD.n722 0.0364848
R8177 VDD.n5843 VDD.n705 0.0364848
R8178 VDD.n5874 VDD.n5873 0.0364848
R8179 VDD.n5895 VDD.n5894 0.0364848
R8180 VDD.n5913 VDD.n682 0.0364848
R8181 VDD.n5924 VDD.n670 0.0364848
R8182 VDD.n4827 VDD.n1501 0.0364844
R8183 VDD.n4706 VDD.n1765 0.0364844
R8184 VDD.n4585 VDD.n2029 0.0364844
R8185 VDD.n4464 VDD.n2293 0.0364844
R8186 VDD.n2889 VDD.n2888 0.0364844
R8187 VDD.n4165 VDD.n3117 0.0364844
R8188 VDD.n4046 VDD.n3383 0.0364844
R8189 VDD.n3927 VDD.n3649 0.0364844
R8190 VDD.n6115 VDD.n6113 0.0351948
R8191 VDD.n2469 VDD.n2467 0.0351948
R8192 VDD.n4942 VDD.n1233 0.0351948
R8193 VDD.n7260 VDD.n7259 0.0351948
R8194 VDD.n7263 VDD.n4 0.0309054
R8195 VDD.n6118 VDD.n611 0.0309054
R8196 VDD.n2480 VDD.n2479 0.0309054
R8197 VDD.n4962 VDD.n4961 0.0309054
R8198 VDD.n5038 VDD.n1191 0.030803
R8199 VDD.n5068 VDD.n1178 0.030803
R8200 VDD.n5079 VDD.n1173 0.030803
R8201 VDD.n5098 VDD.n1166 0.030803
R8202 VDD.n5121 VDD.n1151 0.030803
R8203 VDD.n1146 VDD.n1129 0.030803
R8204 VDD.n1141 VDD.n1133 0.030803
R8205 VDD.n5150 VDD.n1118 0.030803
R8206 VDD.n5160 VDD.n1100 0.030803
R8207 VDD.n1103 VDD.n1094 0.030803
R8208 VDD.n5205 VDD.n5204 0.030803
R8209 VDD.n5216 VDD.n1067 0.030803
R8210 VDD.n5266 VDD.n1056 0.030803
R8211 VDD.n5296 VDD.n1043 0.030803
R8212 VDD.n5307 VDD.n1038 0.030803
R8213 VDD.n5326 VDD.n1031 0.030803
R8214 VDD.n5349 VDD.n1016 0.030803
R8215 VDD.n1011 VDD.n994 0.030803
R8216 VDD.n1006 VDD.n998 0.030803
R8217 VDD.n5378 VDD.n983 0.030803
R8218 VDD.n5388 VDD.n965 0.030803
R8219 VDD.n968 VDD.n959 0.030803
R8220 VDD.n5433 VDD.n5432 0.030803
R8221 VDD.n5444 VDD.n932 0.030803
R8222 VDD.n5494 VDD.n921 0.030803
R8223 VDD.n5524 VDD.n908 0.030803
R8224 VDD.n5535 VDD.n903 0.030803
R8225 VDD.n5554 VDD.n896 0.030803
R8226 VDD.n5577 VDD.n881 0.030803
R8227 VDD.n876 VDD.n859 0.030803
R8228 VDD.n871 VDD.n863 0.030803
R8229 VDD.n5606 VDD.n848 0.030803
R8230 VDD.n5616 VDD.n830 0.030803
R8231 VDD.n833 VDD.n824 0.030803
R8232 VDD.n5661 VDD.n5660 0.030803
R8233 VDD.n5672 VDD.n797 0.030803
R8234 VDD.n5722 VDD.n786 0.030803
R8235 VDD.n5752 VDD.n773 0.030803
R8236 VDD.n5763 VDD.n768 0.030803
R8237 VDD.n5782 VDD.n761 0.030803
R8238 VDD.n5804 VDD.n746 0.030803
R8239 VDD.n741 VDD.n733 0.030803
R8240 VDD.n736 VDD.n725 0.030803
R8241 VDD.n5831 VDD.n717 0.030803
R8242 VDD.n5856 VDD.n708 0.030803
R8243 VDD.n5879 VDD.n697 0.030803
R8244 VDD.n5889 VDD.n677 0.030803
R8245 VDD.n680 VDD.n671 0.030803
R8246 VDD.n5933 VDD.n657 0.030803
R8247 VDD.n5962 VDD.n5960 0.030803
R8248 VDD.n6048 VDD.n5955 0.030803
R8249 VDD.n6040 VDD.n6039 0.030803
R8250 VDD.n6022 VDD.n6010 0.030803
R8251 VDD.n6197 VDD.n563 0.030803
R8252 VDD.n6218 VDD.n552 0.030803
R8253 VDD.n6237 VDD.n545 0.030803
R8254 VDD.n6258 VDD.n530 0.030803
R8255 VDD.n6278 VDD.n519 0.030803
R8256 VDD.n514 VDD.n506 0.030803
R8257 VDD.n509 VDD.n497 0.030803
R8258 VDD.n6308 VDD.n491 0.030803
R8259 VDD.n6331 VDD.n480 0.030803
R8260 VDD.n6341 VDD.n462 0.030803
R8261 VDD.n465 VDD.n457 0.030803
R8262 VDD.n6384 VDD.n444 0.030803
R8263 VDD.n6423 VDD.n429 0.030803
R8264 VDD.n6444 VDD.n418 0.030803
R8265 VDD.n6463 VDD.n411 0.030803
R8266 VDD.n6484 VDD.n396 0.030803
R8267 VDD.n6504 VDD.n385 0.030803
R8268 VDD.n380 VDD.n372 0.030803
R8269 VDD.n375 VDD.n363 0.030803
R8270 VDD.n6534 VDD.n357 0.030803
R8271 VDD.n6557 VDD.n346 0.030803
R8272 VDD.n6567 VDD.n328 0.030803
R8273 VDD.n331 VDD.n323 0.030803
R8274 VDD.n6610 VDD.n310 0.030803
R8275 VDD.n6649 VDD.n295 0.030803
R8276 VDD.n6670 VDD.n284 0.030803
R8277 VDD.n6689 VDD.n277 0.030803
R8278 VDD.n6710 VDD.n262 0.030803
R8279 VDD.n6730 VDD.n251 0.030803
R8280 VDD.n246 VDD.n238 0.030803
R8281 VDD.n241 VDD.n229 0.030803
R8282 VDD.n6760 VDD.n223 0.030803
R8283 VDD.n6783 VDD.n212 0.030803
R8284 VDD.n6793 VDD.n194 0.030803
R8285 VDD.n197 VDD.n189 0.030803
R8286 VDD.n6836 VDD.n176 0.030803
R8287 VDD.n6875 VDD.n161 0.030803
R8288 VDD.n6896 VDD.n150 0.030803
R8289 VDD.n6915 VDD.n143 0.030803
R8290 VDD.n6936 VDD.n128 0.030803
R8291 VDD.n6956 VDD.n117 0.030803
R8292 VDD.n112 VDD.n104 0.030803
R8293 VDD.n107 VDD.n95 0.030803
R8294 VDD.n6986 VDD.n89 0.030803
R8295 VDD.n7009 VDD.n78 0.030803
R8296 VDD.n7019 VDD.n60 0.030803
R8297 VDD.n63 VDD.n55 0.030803
R8298 VDD.n7067 VDD.n42 0.030803
R8299 VDD.n7083 VDD.n28 0.030803
R8300 VDD.n7112 VDD.n7110 0.030803
R8301 VDD.n7198 VDD.n7105 0.030803
R8302 VDD.n7190 VDD.n7189 0.030803
R8303 VDD.n7172 VDD.n7160 0.030803
R8304 VDD.n2767 VDD.n2740 0.030803
R8305 VDD.n2790 VDD.n2752 0.030803
R8306 VDD.n4313 VDD.n2779 0.030803
R8307 VDD.n2831 VDD.n2830 0.030803
R8308 VDD.n2878 VDD.n2813 0.030803
R8309 VDD.n4286 VDD.n2843 0.030803
R8310 VDD.n4281 VDD.n2845 0.030803
R8311 VDD.n4270 VDD.n4269 0.030803
R8312 VDD.n2919 VDD.n2908 0.030803
R8313 VDD.n4249 VDD.n4248 0.030803
R8314 VDD.n2962 VDD.n2951 0.030803
R8315 VDD.n4228 VDD.n4227 0.030803
R8316 VDD.n3032 VDD.n2999 0.030803
R8317 VDD.n4202 VDD.n3021 0.030803
R8318 VDD.n3073 VDD.n3072 0.030803
R8319 VDD.n3101 VDD.n3055 0.030803
R8320 VDD.n4175 VDD.n3085 0.030803
R8321 VDD.n3143 VDD.n3135 0.030803
R8322 VDD.n3138 VDD.n3122 0.030803
R8323 VDD.n4151 VDD.n4150 0.030803
R8324 VDD.n3185 VDD.n3174 0.030803
R8325 VDD.n4130 VDD.n4129 0.030803
R8326 VDD.n3228 VDD.n3217 0.030803
R8327 VDD.n4109 VDD.n4108 0.030803
R8328 VDD.n3298 VDD.n3265 0.030803
R8329 VDD.n4083 VDD.n3287 0.030803
R8330 VDD.n3339 VDD.n3338 0.030803
R8331 VDD.n3367 VDD.n3321 0.030803
R8332 VDD.n4056 VDD.n3351 0.030803
R8333 VDD.n3409 VDD.n3401 0.030803
R8334 VDD.n3404 VDD.n3388 0.030803
R8335 VDD.n4032 VDD.n4031 0.030803
R8336 VDD.n3451 VDD.n3440 0.030803
R8337 VDD.n4011 VDD.n4010 0.030803
R8338 VDD.n3494 VDD.n3483 0.030803
R8339 VDD.n3990 VDD.n3989 0.030803
R8340 VDD.n3564 VDD.n3531 0.030803
R8341 VDD.n3964 VDD.n3553 0.030803
R8342 VDD.n3605 VDD.n3604 0.030803
R8343 VDD.n3633 VDD.n3587 0.030803
R8344 VDD.n3937 VDD.n3617 0.030803
R8345 VDD.n3675 VDD.n3667 0.030803
R8346 VDD.n3670 VDD.n3654 0.030803
R8347 VDD.n3913 VDD.n3912 0.030803
R8348 VDD.n3717 VDD.n3706 0.030803
R8349 VDD.n3892 VDD.n3891 0.030803
R8350 VDD.n3760 VDD.n3749 0.030803
R8351 VDD.n3871 VDD.n3870 0.030803
R8352 VDD.n2636 VDD.n2635 0.030803
R8353 VDD.n2664 VDD.n2444 0.030803
R8354 VDD.n4366 VDD.n2648 0.030803
R8355 VDD.n2705 VDD.n2704 0.030803
R8356 VDD.n2727 VDD.n2687 0.030803
R8357 VDD.n1416 VDD.n1378 0.030803
R8358 VDD.n4864 VDD.n1401 0.030803
R8359 VDD.n1457 VDD.n1456 0.030803
R8360 VDD.n1485 VDD.n1439 0.030803
R8361 VDD.n4837 VDD.n1469 0.030803
R8362 VDD.n1527 VDD.n1519 0.030803
R8363 VDD.n1522 VDD.n1506 0.030803
R8364 VDD.n4813 VDD.n4812 0.030803
R8365 VDD.n1568 VDD.n1556 0.030803
R8366 VDD.n4791 VDD.n4790 0.030803
R8367 VDD.n1610 VDD.n1598 0.030803
R8368 VDD.n4769 VDD.n4768 0.030803
R8369 VDD.n1680 VDD.n1647 0.030803
R8370 VDD.n4743 VDD.n1669 0.030803
R8371 VDD.n1721 VDD.n1720 0.030803
R8372 VDD.n1749 VDD.n1703 0.030803
R8373 VDD.n4716 VDD.n1733 0.030803
R8374 VDD.n1791 VDD.n1783 0.030803
R8375 VDD.n1786 VDD.n1770 0.030803
R8376 VDD.n4692 VDD.n4691 0.030803
R8377 VDD.n1832 VDD.n1820 0.030803
R8378 VDD.n4670 VDD.n4669 0.030803
R8379 VDD.n1874 VDD.n1862 0.030803
R8380 VDD.n4648 VDD.n4647 0.030803
R8381 VDD.n1944 VDD.n1911 0.030803
R8382 VDD.n4622 VDD.n1933 0.030803
R8383 VDD.n1985 VDD.n1984 0.030803
R8384 VDD.n2013 VDD.n1967 0.030803
R8385 VDD.n4595 VDD.n1997 0.030803
R8386 VDD.n2055 VDD.n2047 0.030803
R8387 VDD.n2050 VDD.n2034 0.030803
R8388 VDD.n4571 VDD.n4570 0.030803
R8389 VDD.n2096 VDD.n2084 0.030803
R8390 VDD.n4549 VDD.n4548 0.030803
R8391 VDD.n2138 VDD.n2126 0.030803
R8392 VDD.n4527 VDD.n4526 0.030803
R8393 VDD.n2208 VDD.n2175 0.030803
R8394 VDD.n4501 VDD.n2197 0.030803
R8395 VDD.n2249 VDD.n2248 0.030803
R8396 VDD.n2277 VDD.n2231 0.030803
R8397 VDD.n4474 VDD.n2261 0.030803
R8398 VDD.n2319 VDD.n2311 0.030803
R8399 VDD.n2314 VDD.n2298 0.030803
R8400 VDD.n4450 VDD.n4449 0.030803
R8401 VDD.n2360 VDD.n2348 0.030803
R8402 VDD.n4428 VDD.n4427 0.030803
R8403 VDD.n2402 VDD.n2390 0.030803
R8404 VDD.n4406 VDD.n4405 0.030803
R8405 VDD.n1289 VDD.n1287 0.030803
R8406 VDD.n4916 VDD.n1253 0.030803
R8407 VDD.n1330 VDD.n1329 0.030803
R8408 VDD.n1358 VDD.n1312 0.030803
R8409 VDD.n4889 VDD.n1342 0.030803
R8410 VDD.n3 VDD.n2 0.0292162
R8411 VDD.n6090 VDD.n610 0.0292162
R8412 VDD.n2470 VDD.n2464 0.0292162
R8413 VDD.n4943 VDD.n4936 0.0292162
R8414 VDD VDD.n3860 0.0287804
R8415 VDD.n3846 VDD.n3845 0.0273994
R8416 VDD.n2522 VDD.n2521 0.0273994
R8417 VDD.n7079 VDD.n7078 0.026557
R8418 VDD.n5929 VDD.n5928 0.026557
R8419 VDD.n609 VDD 0.0265417
R8420 VDD VDD.n1 0.0265417
R8421 VDD.n4395 VDD.n4394 0.0263291
R8422 VDD.n6402 VDD 0.0257316
R8423 VDD.n6628 VDD 0.0257316
R8424 VDD.n6854 VDD 0.0257316
R8425 VDD VDD.n7076 0.0257316
R8426 VDD.n5236 VDD 0.0257316
R8427 VDD.n5464 VDD 0.0257316
R8428 VDD.n5692 VDD 0.0257316
R8429 VDD VDD.n5926 0.0257316
R8430 VDD.n4761 VDD 0.0254688
R8431 VDD.n4640 VDD 0.0254688
R8432 VDD.n4519 VDD 0.0254688
R8433 VDD.n4398 VDD 0.0254688
R8434 VDD.n4220 VDD 0.0254688
R8435 VDD.n4101 VDD 0.0254688
R8436 VDD.n3982 VDD 0.0254688
R8437 VDD.n3863 VDD 0.0254688
R8438 VDD.n3827 VDD.n3803 0.0252507
R8439 VDD.n3813 VDD.n3799 0.0252507
R8440 VDD.n3816 VDD.n3795 0.0252507
R8441 VDD.n3810 VDD.n3791 0.0252507
R8442 VDD.n3806 VDD.n3787 0.0252507
R8443 VDD.n2580 VDD.n2579 0.0252507
R8444 VDD.n2574 VDD.n2573 0.0252507
R8445 VDD.n2592 VDD.n2568 0.0252507
R8446 VDD.n2543 VDD.n2533 0.0252507
R8447 VDD.n2503 VDD.n2500 0.0252507
R8448 VDD.n2496 VDD.n2495 0.0252507
R8449 VDD.n2559 VDD.n2490 0.0252507
R8450 VDD.n2551 VDD.n2548 0.0252507
R8451 VDD.n6106 VDD.n618 0.0242893
R8452 VDD.n625 VDD.n622 0.0242893
R8453 VDD.n6098 VDD.n629 0.0242893
R8454 VDD.n6152 VDD.n6148 0.0242893
R8455 VDD.n6162 VDD.n578 0.0242893
R8456 VDD.n6143 VDD.n6141 0.0242893
R8457 VDD.n585 VDD.n581 0.0242893
R8458 VDD.n6170 VDD.n572 0.0242893
R8459 VDD.n5009 VDD.n1202 0.0242893
R8460 VDD.n4995 VDD.n4991 0.0242893
R8461 VDD.n5001 VDD.n1208 0.0242893
R8462 VDD.n4986 VDD.n4984 0.0242893
R8463 VDD.n1215 VDD.n1211 0.0242893
R8464 VDD.n6119 VDD.n609 0.0239375
R8465 VDD.n7264 VDD.n1 0.0239375
R8466 VDD.n595 VDD.n594 0.0234759
R8467 VDD.n3839 VDD.n3838 0.0234759
R8468 VDD.n2515 VDD.n2514 0.0234759
R8469 VDD.n1225 VDD.n1224 0.0234759
R8470 VDD.n6137 VDD 0.0234268
R8471 VDD.n6131 VDD 0.0226354
R8472 VDD.n2475 VDD.n2471 0.0226354
R8473 VDD.n2618 VDD 0.0226354
R8474 VDD.n4934 VDD.n1234 0.0226354
R8475 VDD.n4955 VDD 0.0226354
R8476 VDD.n7255 VDD 0.0226354
R8477 VDD.n2432 VDD.n2430 0.0212996
R8478 VDD.n1279 VDD.n1265 0.0212996
R8479 VDD.n6005 VDD.n6004 0.0206084
R8480 VDD.n7155 VDD.n7154 0.0206084
R8481 VDD.n5029 VDD.n5028 0.0205441
R8482 VDD.n5050 VDD.n5049 0.0205441
R8483 VDD.n5059 VDD.n5058 0.0205441
R8484 VDD.n5088 VDD.n5087 0.0205441
R8485 VDD.n5111 VDD.n5110 0.0205441
R8486 VDD.n5132 VDD.n5131 0.0205441
R8487 VDD.n5257 VDD.n5256 0.0205441
R8488 VDD.n5278 VDD.n5277 0.0205441
R8489 VDD.n5287 VDD.n5286 0.0205441
R8490 VDD.n5316 VDD.n5315 0.0205441
R8491 VDD.n5339 VDD.n5338 0.0205441
R8492 VDD.n5360 VDD.n5359 0.0205441
R8493 VDD.n5485 VDD.n5484 0.0205441
R8494 VDD.n5506 VDD.n5505 0.0205441
R8495 VDD.n5515 VDD.n5514 0.0205441
R8496 VDD.n5544 VDD.n5543 0.0205441
R8497 VDD.n5567 VDD.n5566 0.0205441
R8498 VDD.n5588 VDD.n5587 0.0205441
R8499 VDD.n5713 VDD.n5712 0.0205441
R8500 VDD.n5734 VDD.n5733 0.0205441
R8501 VDD.n5743 VDD.n5742 0.0205441
R8502 VDD.n5772 VDD.n5771 0.0205441
R8503 VDD.n5795 VDD.n5794 0.0205441
R8504 VDD.n5815 VDD.n5814 0.0205441
R8505 VDD.n6188 VDD.n6187 0.0205441
R8506 VDD.n6209 VDD.n6208 0.0205441
R8507 VDD.n6227 VDD.n6226 0.0205441
R8508 VDD.n6249 VDD.n6248 0.0205441
R8509 VDD.n6269 VDD.n6268 0.0205441
R8510 VDD.n6288 VDD.n6287 0.0205441
R8511 VDD.n6414 VDD.n6413 0.0205441
R8512 VDD.n6435 VDD.n6434 0.0205441
R8513 VDD.n6453 VDD.n6452 0.0205441
R8514 VDD.n6475 VDD.n6474 0.0205441
R8515 VDD.n6495 VDD.n6494 0.0205441
R8516 VDD.n6514 VDD.n6513 0.0205441
R8517 VDD.n6640 VDD.n6639 0.0205441
R8518 VDD.n6661 VDD.n6660 0.0205441
R8519 VDD.n6679 VDD.n6678 0.0205441
R8520 VDD.n6701 VDD.n6700 0.0205441
R8521 VDD.n6721 VDD.n6720 0.0205441
R8522 VDD.n6740 VDD.n6739 0.0205441
R8523 VDD.n6866 VDD.n6865 0.0205441
R8524 VDD.n6887 VDD.n6886 0.0205441
R8525 VDD.n6905 VDD.n6904 0.0205441
R8526 VDD.n6927 VDD.n6926 0.0205441
R8527 VDD.n6947 VDD.n6946 0.0205441
R8528 VDD.n6966 VDD.n6965 0.0205441
R8529 VDD.n4331 VDD.n4330 0.0205441
R8530 VDD.n2788 VDD.n2750 0.0205441
R8531 VDD.n2803 VDD.n2802 0.0205441
R8532 VDD.n4302 VDD.n2807 0.0205441
R8533 VDD.n2872 VDD.n2871 0.0205441
R8534 VDD.n2887 VDD.n2886 0.0205441
R8535 VDD.n3030 VDD.n2992 0.0205441
R8536 VDD.n3045 VDD.n3044 0.0205441
R8537 VDD.n4191 VDD.n3049 0.0205441
R8538 VDD.n3098 VDD.n3097 0.0205441
R8539 VDD.n3114 VDD.n3113 0.0205441
R8540 VDD.n4164 VDD.n3118 0.0205441
R8541 VDD.n3296 VDD.n3258 0.0205441
R8542 VDD.n3311 VDD.n3310 0.0205441
R8543 VDD.n4072 VDD.n3315 0.0205441
R8544 VDD.n3364 VDD.n3363 0.0205441
R8545 VDD.n3380 VDD.n3379 0.0205441
R8546 VDD.n4045 VDD.n3384 0.0205441
R8547 VDD.n3562 VDD.n3524 0.0205441
R8548 VDD.n3577 VDD.n3576 0.0205441
R8549 VDD.n3953 VDD.n3581 0.0205441
R8550 VDD.n3630 VDD.n3629 0.0205441
R8551 VDD.n3646 VDD.n3645 0.0205441
R8552 VDD.n3926 VDD.n3650 0.0205441
R8553 VDD.n4382 VDD.n2438 0.0205441
R8554 VDD.n2661 VDD.n2660 0.0205441
R8555 VDD.n2677 VDD.n2676 0.0205441
R8556 VDD.n4355 VDD.n2681 0.0205441
R8557 VDD.n2723 VDD.n2718 0.0205441
R8558 VDD.n1413 VDD.n1412 0.0205441
R8559 VDD.n1429 VDD.n1428 0.0205441
R8560 VDD.n4853 VDD.n1433 0.0205441
R8561 VDD.n1482 VDD.n1481 0.0205441
R8562 VDD.n1498 VDD.n1497 0.0205441
R8563 VDD.n4826 VDD.n1502 0.0205441
R8564 VDD.n1678 VDD.n1641 0.0205441
R8565 VDD.n1693 VDD.n1692 0.0205441
R8566 VDD.n4732 VDD.n1697 0.0205441
R8567 VDD.n1746 VDD.n1745 0.0205441
R8568 VDD.n1762 VDD.n1761 0.0205441
R8569 VDD.n4705 VDD.n1766 0.0205441
R8570 VDD.n1942 VDD.n1905 0.0205441
R8571 VDD.n1957 VDD.n1956 0.0205441
R8572 VDD.n4611 VDD.n1961 0.0205441
R8573 VDD.n2010 VDD.n2009 0.0205441
R8574 VDD.n2026 VDD.n2025 0.0205441
R8575 VDD.n4584 VDD.n2030 0.0205441
R8576 VDD.n2206 VDD.n2169 0.0205441
R8577 VDD.n2221 VDD.n2220 0.0205441
R8578 VDD.n4490 VDD.n2225 0.0205441
R8579 VDD.n2274 VDD.n2273 0.0205441
R8580 VDD.n2290 VDD.n2289 0.0205441
R8581 VDD.n4463 VDD.n2294 0.0205441
R8582 VDD.n1284 VDD.n1262 0.0205441
R8583 VDD.n1302 VDD.n1301 0.0205441
R8584 VDD.n4905 VDD.n1306 0.0205441
R8585 VDD.n1355 VDD.n1354 0.0205441
R8586 VDD.n1371 VDD.n1370 0.0205441
R8587 VDD.n5134 VDD.n5133 0.0198529
R8588 VDD.n5139 VDD.n5138 0.0198529
R8589 VDD.n5172 VDD.n5171 0.0198529
R8590 VDD.n5193 VDD.n1091 0.0198529
R8591 VDD.n1089 VDD.n1088 0.0198529
R8592 VDD.n5228 VDD.n5227 0.0198529
R8593 VDD.n5362 VDD.n5361 0.0198529
R8594 VDD.n5367 VDD.n5366 0.0198529
R8595 VDD.n5400 VDD.n5399 0.0198529
R8596 VDD.n5421 VDD.n956 0.0198529
R8597 VDD.n954 VDD.n953 0.0198529
R8598 VDD.n5456 VDD.n5455 0.0198529
R8599 VDD.n5590 VDD.n5589 0.0198529
R8600 VDD.n5595 VDD.n5594 0.0198529
R8601 VDD.n5628 VDD.n5627 0.0198529
R8602 VDD.n5649 VDD.n821 0.0198529
R8603 VDD.n819 VDD.n818 0.0198529
R8604 VDD.n5684 VDD.n5683 0.0198529
R8605 VDD.n5820 VDD.n727 0.0198529
R8606 VDD.n5842 VDD.n719 0.0198529
R8607 VDD.n5863 VDD.n5862 0.0198529
R8608 VDD.n5868 VDD.n5867 0.0198529
R8609 VDD.n5901 VDD.n5900 0.0198529
R8610 VDD.n5905 VDD.n686 0.0198529
R8611 VDD.n5945 VDD.n5944 0.0198529
R8612 VDD.n5950 VDD.n663 0.0198529
R8613 VDD.n5981 VDD.n5978 0.0198529
R8614 VDD.n6036 VDD.n5975 0.0198529
R8615 VDD.n6030 VDD.n6029 0.0198529
R8616 VDD.n6294 VDD.n500 0.0198529
R8617 VDD.n6315 VDD.n6314 0.0198529
R8618 VDD.n6320 VDD.n6319 0.0198529
R8619 VDD.n6353 VDD.n6352 0.0198529
R8620 VDD.n6374 VDD.n454 0.0198529
R8621 VDD.n6398 VDD.n441 0.0198529
R8622 VDD.n6520 VDD.n366 0.0198529
R8623 VDD.n6541 VDD.n6540 0.0198529
R8624 VDD.n6546 VDD.n6545 0.0198529
R8625 VDD.n6579 VDD.n6578 0.0198529
R8626 VDD.n6600 VDD.n320 0.0198529
R8627 VDD.n6624 VDD.n307 0.0198529
R8628 VDD.n6746 VDD.n232 0.0198529
R8629 VDD.n6767 VDD.n6766 0.0198529
R8630 VDD.n6772 VDD.n6771 0.0198529
R8631 VDD.n6805 VDD.n6804 0.0198529
R8632 VDD.n6826 VDD.n186 0.0198529
R8633 VDD.n6850 VDD.n173 0.0198529
R8634 VDD.n6972 VDD.n98 0.0198529
R8635 VDD.n6993 VDD.n6992 0.0198529
R8636 VDD.n6998 VDD.n6997 0.0198529
R8637 VDD.n7031 VDD.n7030 0.0198529
R8638 VDD.n7052 VDD.n52 0.0198529
R8639 VDD.n7056 VDD.n50 0.0198529
R8640 VDD.n7095 VDD.n7094 0.0198529
R8641 VDD.n7100 VDD.n34 0.0198529
R8642 VDD.n7131 VDD.n7128 0.0198529
R8643 VDD.n7186 VDD.n7125 0.0198529
R8644 VDD.n7180 VDD.n7179 0.0198529
R8645 VDD.n2893 VDD.n2864 0.0198529
R8646 VDD.n2901 VDD.n2857 0.0198529
R8647 VDD.n4261 VDD.n4260 0.0198529
R8648 VDD.n2944 VDD.n2932 0.0198529
R8649 VDD.n4240 VDD.n4239 0.0198529
R8650 VDD.n4224 VDD.n2976 0.0198529
R8651 VDD.n4163 VDD.n4162 0.0198529
R8652 VDD.n3167 VDD.n3155 0.0198529
R8653 VDD.n4142 VDD.n4141 0.0198529
R8654 VDD.n3210 VDD.n3198 0.0198529
R8655 VDD.n4121 VDD.n4120 0.0198529
R8656 VDD.n4105 VDD.n3242 0.0198529
R8657 VDD.n4044 VDD.n4043 0.0198529
R8658 VDD.n3433 VDD.n3421 0.0198529
R8659 VDD.n4023 VDD.n4022 0.0198529
R8660 VDD.n3476 VDD.n3464 0.0198529
R8661 VDD.n4002 VDD.n4001 0.0198529
R8662 VDD.n3986 VDD.n3508 0.0198529
R8663 VDD.n3925 VDD.n3924 0.0198529
R8664 VDD.n3699 VDD.n3687 0.0198529
R8665 VDD.n3904 VDD.n3903 0.0198529
R8666 VDD.n3742 VDD.n3730 0.0198529
R8667 VDD.n3883 VDD.n3882 0.0198529
R8668 VDD.n3867 VDD.n3774 0.0198529
R8669 VDD.n4825 VDD.n4824 0.0198529
R8670 VDD.n4809 VDD.n1540 0.0198529
R8671 VDD.n4803 VDD.n4802 0.0198529
R8672 VDD.n4787 VDD.n1582 0.0198529
R8673 VDD.n4781 VDD.n4780 0.0198529
R8674 VDD.n4765 VDD.n1624 0.0198529
R8675 VDD.n4704 VDD.n4703 0.0198529
R8676 VDD.n4688 VDD.n1804 0.0198529
R8677 VDD.n4682 VDD.n4681 0.0198529
R8678 VDD.n4666 VDD.n1846 0.0198529
R8679 VDD.n4660 VDD.n4659 0.0198529
R8680 VDD.n4644 VDD.n1888 0.0198529
R8681 VDD.n4583 VDD.n4582 0.0198529
R8682 VDD.n4567 VDD.n2068 0.0198529
R8683 VDD.n4561 VDD.n4560 0.0198529
R8684 VDD.n4545 VDD.n2110 0.0198529
R8685 VDD.n4539 VDD.n4538 0.0198529
R8686 VDD.n4523 VDD.n2152 0.0198529
R8687 VDD.n4462 VDD.n4461 0.0198529
R8688 VDD.n4446 VDD.n2332 0.0198529
R8689 VDD.n4440 VDD.n4439 0.0198529
R8690 VDD.n4424 VDD.n2374 0.0198529
R8691 VDD.n4418 VDD.n4417 0.0198529
R8692 VDD.n4402 VDD.n2416 0.0198529
R8693 VDD.n6112 VDD.n6111 0.0188117
R8694 VDD.n6114 VDD.n6112 0.0188117
R8695 VDD.n2610 VDD.n2462 0.0188117
R8696 VDD.n2611 VDD.n2610 0.0188117
R8697 VDD.n4946 VDD.n4941 0.0188117
R8698 VDD.n4947 VDD.n4946 0.0188117
R8699 VDD.n7245 VDD.n7244 0.0188117
R8700 VDD.n5023 VDD.n5022 0.0184706
R8701 VDD.n5034 VDD.n5033 0.0184706
R8702 VDD.n5064 VDD.n5063 0.0184706
R8703 VDD.n5085 VDD.n1170 0.0184706
R8704 VDD.n5093 VDD.n5092 0.0184706
R8705 VDD.n5117 VDD.n5116 0.0184706
R8706 VDD.n5143 VDD.n1123 0.0184706
R8707 VDD.n5167 VDD.n1109 0.0184706
R8708 VDD.n5178 VDD.n1107 0.0184706
R8709 VDD.n5200 VDD.n1087 0.0184706
R8710 VDD.n5223 VDD.n1075 0.0184706
R8711 VDD.n5238 VDD.n1072 0.0184706
R8712 VDD.n5233 VDD.n5232 0.0184706
R8713 VDD.n5262 VDD.n5261 0.0184706
R8714 VDD.n5292 VDD.n5291 0.0184706
R8715 VDD.n5313 VDD.n1035 0.0184706
R8716 VDD.n5321 VDD.n5320 0.0184706
R8717 VDD.n5345 VDD.n5344 0.0184706
R8718 VDD.n5371 VDD.n988 0.0184706
R8719 VDD.n5395 VDD.n974 0.0184706
R8720 VDD.n5406 VDD.n972 0.0184706
R8721 VDD.n5428 VDD.n952 0.0184706
R8722 VDD.n5451 VDD.n940 0.0184706
R8723 VDD.n5466 VDD.n937 0.0184706
R8724 VDD.n5461 VDD.n5460 0.0184706
R8725 VDD.n5490 VDD.n5489 0.0184706
R8726 VDD.n5520 VDD.n5519 0.0184706
R8727 VDD.n5541 VDD.n900 0.0184706
R8728 VDD.n5549 VDD.n5548 0.0184706
R8729 VDD.n5573 VDD.n5572 0.0184706
R8730 VDD.n5599 VDD.n853 0.0184706
R8731 VDD.n5623 VDD.n839 0.0184706
R8732 VDD.n5634 VDD.n837 0.0184706
R8733 VDD.n5656 VDD.n817 0.0184706
R8734 VDD.n5679 VDD.n805 0.0184706
R8735 VDD.n5694 VDD.n802 0.0184706
R8736 VDD.n5689 VDD.n5688 0.0184706
R8737 VDD.n5718 VDD.n5717 0.0184706
R8738 VDD.n5748 VDD.n5747 0.0184706
R8739 VDD.n5769 VDD.n765 0.0184706
R8740 VDD.n5777 VDD.n5776 0.0184706
R8741 VDD.n5800 VDD.n5799 0.0184706
R8742 VDD.n5835 VDD.n721 0.0184706
R8743 VDD.n5860 VDD.n704 0.0184706
R8744 VDD.n5872 VDD.n702 0.0184706
R8745 VDD.n5896 VDD.n688 0.0184706
R8746 VDD.n5911 VDD.n685 0.0184706
R8747 VDD.n5925 VDD.n669 0.0184706
R8748 VDD.n5940 VDD.n665 0.0184706
R8749 VDD.n6061 VDD.n662 0.0184706
R8750 VDD.n6055 VDD.n5951 0.0184706
R8751 VDD.n5990 VDD.n5985 0.0184706
R8752 VDD.n5995 VDD.n5976 0.0184706
R8753 VDD.n6008 VDD.n6000 0.0184706
R8754 VDD.n6183 VDD.n6182 0.0184706
R8755 VDD.n6203 VDD.n6202 0.0184706
R8756 VDD.n6224 VDD.n549 0.0184706
R8757 VDD.n6232 VDD.n6231 0.0184706
R8758 VDD.n6254 VDD.n6253 0.0184706
R8759 VDD.n6274 VDD.n6273 0.0184706
R8760 VDD.n6312 VDD.n487 0.0184706
R8761 VDD.n6324 VDD.n485 0.0184706
R8762 VDD.n6348 VDD.n471 0.0184706
R8763 VDD.n6359 VDD.n469 0.0184706
R8764 VDD.n6380 VDD.n452 0.0184706
R8765 VDD.n6404 VDD.n439 0.0184706
R8766 VDD.n6409 VDD.n6408 0.0184706
R8767 VDD.n6429 VDD.n6428 0.0184706
R8768 VDD.n6450 VDD.n415 0.0184706
R8769 VDD.n6458 VDD.n6457 0.0184706
R8770 VDD.n6480 VDD.n6479 0.0184706
R8771 VDD.n6500 VDD.n6499 0.0184706
R8772 VDD.n6538 VDD.n353 0.0184706
R8773 VDD.n6550 VDD.n351 0.0184706
R8774 VDD.n6574 VDD.n337 0.0184706
R8775 VDD.n6585 VDD.n335 0.0184706
R8776 VDD.n6606 VDD.n318 0.0184706
R8777 VDD.n6630 VDD.n305 0.0184706
R8778 VDD.n6635 VDD.n6634 0.0184706
R8779 VDD.n6655 VDD.n6654 0.0184706
R8780 VDD.n6676 VDD.n281 0.0184706
R8781 VDD.n6684 VDD.n6683 0.0184706
R8782 VDD.n6706 VDD.n6705 0.0184706
R8783 VDD.n6726 VDD.n6725 0.0184706
R8784 VDD.n6764 VDD.n219 0.0184706
R8785 VDD.n6776 VDD.n217 0.0184706
R8786 VDD.n6800 VDD.n203 0.0184706
R8787 VDD.n6811 VDD.n201 0.0184706
R8788 VDD.n6832 VDD.n184 0.0184706
R8789 VDD.n6856 VDD.n171 0.0184706
R8790 VDD.n6861 VDD.n6860 0.0184706
R8791 VDD.n6881 VDD.n6880 0.0184706
R8792 VDD.n6902 VDD.n147 0.0184706
R8793 VDD.n6910 VDD.n6909 0.0184706
R8794 VDD.n6932 VDD.n6931 0.0184706
R8795 VDD.n6952 VDD.n6951 0.0184706
R8796 VDD.n6990 VDD.n85 0.0184706
R8797 VDD.n7002 VDD.n83 0.0184706
R8798 VDD.n7026 VDD.n69 0.0184706
R8799 VDD.n7037 VDD.n67 0.0184706
R8800 VDD.n7062 VDD.n49 0.0184706
R8801 VDD.n7075 VDD.n40 0.0184706
R8802 VDD.n7090 VDD.n36 0.0184706
R8803 VDD.n7211 VDD.n33 0.0184706
R8804 VDD.n7205 VDD.n7101 0.0184706
R8805 VDD.n7140 VDD.n7135 0.0184706
R8806 VDD.n7145 VDD.n7126 0.0184706
R8807 VDD.n7158 VDD.n7150 0.0184706
R8808 VDD.n4335 VDD.n2737 0.0184706
R8809 VDD.n4326 VDD.n2746 0.0184706
R8810 VDD.n2796 VDD.n2786 0.0184706
R8811 VDD.n4306 VDD.n2783 0.0184706
R8812 VDD.n4300 VDD.n2808 0.0184706
R8813 VDD.n2884 VDD.n2866 0.0184706
R8814 VDD.n2899 VDD.n2862 0.0184706
R8815 VDD.n4265 VDD.n2860 0.0184706
R8816 VDD.n2942 VDD.n2939 0.0184706
R8817 VDD.n4244 VDD.n2935 0.0184706
R8818 VDD.n2983 VDD.n2980 0.0184706
R8819 VDD.n2987 VDD.n2977 0.0184706
R8820 VDD.n4215 VDD.n2988 0.0184706
R8821 VDD.n3038 VDD.n3028 0.0184706
R8822 VDD.n4195 VDD.n3025 0.0184706
R8823 VDD.n4189 VDD.n3050 0.0184706
R8824 VDD.n3107 VDD.n3092 0.0184706
R8825 VDD.n4168 VDD.n3089 0.0184706
R8826 VDD.n3165 VDD.n3162 0.0184706
R8827 VDD.n4146 VDD.n3158 0.0184706
R8828 VDD.n3208 VDD.n3205 0.0184706
R8829 VDD.n4125 VDD.n3201 0.0184706
R8830 VDD.n3249 VDD.n3246 0.0184706
R8831 VDD.n3253 VDD.n3243 0.0184706
R8832 VDD.n4096 VDD.n3254 0.0184706
R8833 VDD.n3304 VDD.n3294 0.0184706
R8834 VDD.n4076 VDD.n3291 0.0184706
R8835 VDD.n4070 VDD.n3316 0.0184706
R8836 VDD.n3373 VDD.n3358 0.0184706
R8837 VDD.n4049 VDD.n3355 0.0184706
R8838 VDD.n3431 VDD.n3428 0.0184706
R8839 VDD.n4027 VDD.n3424 0.0184706
R8840 VDD.n3474 VDD.n3471 0.0184706
R8841 VDD.n4006 VDD.n3467 0.0184706
R8842 VDD.n3515 VDD.n3512 0.0184706
R8843 VDD.n3519 VDD.n3509 0.0184706
R8844 VDD.n3977 VDD.n3520 0.0184706
R8845 VDD.n3570 VDD.n3560 0.0184706
R8846 VDD.n3957 VDD.n3557 0.0184706
R8847 VDD.n3951 VDD.n3582 0.0184706
R8848 VDD.n3639 VDD.n3624 0.0184706
R8849 VDD.n3930 VDD.n3621 0.0184706
R8850 VDD.n3697 VDD.n3694 0.0184706
R8851 VDD.n3908 VDD.n3690 0.0184706
R8852 VDD.n3740 VDD.n3737 0.0184706
R8853 VDD.n3887 VDD.n3733 0.0184706
R8854 VDD.n3781 VDD.n3778 0.0184706
R8855 VDD.n3862 VDD.n3775 0.0184706
R8856 VDD.n4387 VDD.n4386 0.0184706
R8857 VDD.n4380 VDD.n2439 0.0184706
R8858 VDD.n2670 VDD.n2655 0.0184706
R8859 VDD.n4359 VDD.n2652 0.0184706
R8860 VDD.n4353 VDD.n2682 0.0184706
R8861 VDD.n2733 VDD.n2732 0.0184706
R8862 VDD.n4876 VDD.n1375 0.0184706
R8863 VDD.n1422 VDD.n1408 0.0184706
R8864 VDD.n4857 VDD.n1405 0.0184706
R8865 VDD.n4851 VDD.n1434 0.0184706
R8866 VDD.n1491 VDD.n1476 0.0184706
R8867 VDD.n4830 VDD.n1473 0.0184706
R8868 VDD.n1547 VDD.n1544 0.0184706
R8869 VDD.n1552 VDD.n1541 0.0184706
R8870 VDD.n1589 VDD.n1586 0.0184706
R8871 VDD.n1594 VDD.n1583 0.0184706
R8872 VDD.n1631 VDD.n1628 0.0184706
R8873 VDD.n1635 VDD.n1625 0.0184706
R8874 VDD.n4756 VDD.n1636 0.0184706
R8875 VDD.n1686 VDD.n1676 0.0184706
R8876 VDD.n4736 VDD.n1673 0.0184706
R8877 VDD.n4730 VDD.n1698 0.0184706
R8878 VDD.n1755 VDD.n1740 0.0184706
R8879 VDD.n4709 VDD.n1737 0.0184706
R8880 VDD.n1811 VDD.n1808 0.0184706
R8881 VDD.n1816 VDD.n1805 0.0184706
R8882 VDD.n1853 VDD.n1850 0.0184706
R8883 VDD.n1858 VDD.n1847 0.0184706
R8884 VDD.n1895 VDD.n1892 0.0184706
R8885 VDD.n1899 VDD.n1889 0.0184706
R8886 VDD.n4635 VDD.n1900 0.0184706
R8887 VDD.n1950 VDD.n1940 0.0184706
R8888 VDD.n4615 VDD.n1937 0.0184706
R8889 VDD.n4609 VDD.n1962 0.0184706
R8890 VDD.n2019 VDD.n2004 0.0184706
R8891 VDD.n4588 VDD.n2001 0.0184706
R8892 VDD.n2075 VDD.n2072 0.0184706
R8893 VDD.n2080 VDD.n2069 0.0184706
R8894 VDD.n2117 VDD.n2114 0.0184706
R8895 VDD.n2122 VDD.n2111 0.0184706
R8896 VDD.n2159 VDD.n2156 0.0184706
R8897 VDD.n2163 VDD.n2153 0.0184706
R8898 VDD.n4514 VDD.n2164 0.0184706
R8899 VDD.n2214 VDD.n2204 0.0184706
R8900 VDD.n4494 VDD.n2201 0.0184706
R8901 VDD.n4488 VDD.n2226 0.0184706
R8902 VDD.n2283 VDD.n2268 0.0184706
R8903 VDD.n4467 VDD.n2265 0.0184706
R8904 VDD.n2339 VDD.n2336 0.0184706
R8905 VDD.n2344 VDD.n2333 0.0184706
R8906 VDD.n2381 VDD.n2378 0.0184706
R8907 VDD.n2386 VDD.n2375 0.0184706
R8908 VDD.n2423 VDD.n2420 0.0184706
R8909 VDD.n4397 VDD.n2417 0.0184706
R8910 VDD.n1278 VDD.n1264 0.0184706
R8911 VDD.n1295 VDD.n1260 0.0184706
R8912 VDD.n4909 VDD.n1257 0.0184706
R8913 VDD.n4903 VDD.n1307 0.0184706
R8914 VDD.n1364 VDD.n1349 0.0184706
R8915 VDD.n4882 VDD.n1346 0.0184706
R8916 VDD.n2481 VDD.n2477 0.0174271
R8917 VDD.n4963 VDD.n4935 0.0174271
R8918 VDD.n598 VDD.n589 0.0172857
R8919 VDD.n1228 VDD.n1219 0.0172857
R8920 VDD.n3852 VDD.n3851 0.0167579
R8921 VDD.n2528 VDD.n2527 0.0167579
R8922 VDD.n6089 VDD.n608 0.016125
R8923 VDD.n7278 VDD.n7277 0.016125
R8924 VDD VDD.n4395 0.0159219
R8925 VDD.n7077 VDD 0.0158368
R8926 VDD.n5927 VDD 0.0158368
R8927 VDD.n2584 VDD.n2583 0.0157919
R8928 VDD.n6105 VDD.n617 0.0156071
R8929 VDD.n6109 VDD.n617 0.0156071
R8930 VDD.n626 VDD.n621 0.0156071
R8931 VDD.n626 VDD.n616 0.0156071
R8932 VDD.n6102 VDD.n628 0.0156071
R8933 VDD.n6102 VDD.n6101 0.0156071
R8934 VDD.n6178 VDD.n569 0.0156071
R8935 VDD.n6151 VDD.n6150 0.0156071
R8936 VDD.n6151 VDD.n6149 0.0156071
R8937 VDD.n6166 VDD.n577 0.0156071
R8938 VDD.n6166 VDD.n6165 0.0156071
R8939 VDD.n6140 VDD.n576 0.0156071
R8940 VDD.n6142 VDD.n576 0.0156071
R8941 VDD.n584 VDD.n583 0.0156071
R8942 VDD.n584 VDD.n582 0.0156071
R8943 VDD.n6169 VDD.n571 0.0156071
R8944 VDD.n6173 VDD.n571 0.0156071
R8945 VDD.n5008 VDD.n1201 0.0156071
R8946 VDD.n5012 VDD.n1201 0.0156071
R8947 VDD.n5017 VDD.n1199 0.0156071
R8948 VDD.n4994 VDD.n4993 0.0156071
R8949 VDD.n4994 VDD.n4992 0.0156071
R8950 VDD.n5005 VDD.n1207 0.0156071
R8951 VDD.n5005 VDD.n5004 0.0156071
R8952 VDD.n4983 VDD.n1206 0.0156071
R8953 VDD.n4985 VDD.n1206 0.0156071
R8954 VDD.n1214 VDD.n1213 0.0156071
R8955 VDD.n1214 VDD.n1212 0.0156071
R8956 VDD.n3844 VDD.n3832 0.0156071
R8957 VDD.n3847 VDD.n3828 0.0156071
R8958 VDD.n3850 VDD.n3800 0.0156071
R8959 VDD.n3853 VDD.n3796 0.0156071
R8960 VDD.n3856 VDD.n3792 0.0156071
R8961 VDD.n3859 VDD.n3788 0.0156071
R8962 VDD.n2582 VDD.n2581 0.0156071
R8963 VDD.n2585 VDD.n2575 0.0156071
R8964 VDD.n2591 VDD.n2569 0.0156071
R8965 VDD.n2545 VDD.n2544 0.0156071
R8966 VDD.n2520 VDD.n2508 0.0156071
R8967 VDD.n2523 VDD.n2504 0.0156071
R8968 VDD.n2526 VDD.n2497 0.0156071
R8969 VDD.n2558 VDD.n2491 0.0156071
R8970 VDD.n2553 VDD.n2552 0.0156071
R8971 VDD.n6003 VDD.n635 0.0152558
R8972 VDD.n7153 VDD.n6 0.0152558
R8973 VDD.n4391 VDD.n4390 0.0152558
R8974 VDD.n1271 VDD.n1268 0.0152558
R8975 VDD.n596 VDD.n593 0.0148621
R8976 VDD.n3840 VDD.n3837 0.0148621
R8977 VDD.n2516 VDD.n2513 0.0148621
R8978 VDD.n1226 VDD.n1223 0.0148621
R8979 VDD.n3849 VDD.n3848 0.0148365
R8980 VDD.n2525 VDD.n2524 0.0148365
R8981 VDD.n5029 VDD.n1194 0.0143235
R8982 VDD.n5050 VDD.n1182 0.0143235
R8983 VDD.n5058 VDD.n5054 0.0143235
R8984 VDD.n5088 VDD.n1168 0.0143235
R8985 VDD.n5111 VDD.n1154 0.0143235
R8986 VDD.n5140 VDD.n5139 0.0143235
R8987 VDD.n5171 VDD.n5170 0.0143235
R8988 VDD.n5177 VDD.n1091 0.0143235
R8989 VDD.n5199 VDD.n1089 0.0143235
R8990 VDD.n5227 VDD.n5226 0.0143235
R8991 VDD.n5257 VDD.n1059 0.0143235
R8992 VDD.n5278 VDD.n1047 0.0143235
R8993 VDD.n5286 VDD.n5282 0.0143235
R8994 VDD.n5316 VDD.n1033 0.0143235
R8995 VDD.n5339 VDD.n1019 0.0143235
R8996 VDD.n5368 VDD.n5367 0.0143235
R8997 VDD.n5399 VDD.n5398 0.0143235
R8998 VDD.n5405 VDD.n956 0.0143235
R8999 VDD.n5427 VDD.n954 0.0143235
R9000 VDD.n5455 VDD.n5454 0.0143235
R9001 VDD.n5485 VDD.n924 0.0143235
R9002 VDD.n5506 VDD.n912 0.0143235
R9003 VDD.n5514 VDD.n5510 0.0143235
R9004 VDD.n5544 VDD.n898 0.0143235
R9005 VDD.n5567 VDD.n884 0.0143235
R9006 VDD.n5596 VDD.n5595 0.0143235
R9007 VDD.n5627 VDD.n5626 0.0143235
R9008 VDD.n5633 VDD.n821 0.0143235
R9009 VDD.n5655 VDD.n819 0.0143235
R9010 VDD.n5683 VDD.n5682 0.0143235
R9011 VDD.n5713 VDD.n789 0.0143235
R9012 VDD.n5734 VDD.n777 0.0143235
R9013 VDD.n5742 VDD.n5738 0.0143235
R9014 VDD.n5772 VDD.n763 0.0143235
R9015 VDD.n5795 VDD.n749 0.0143235
R9016 VDD.n5836 VDD.n719 0.0143235
R9017 VDD.n5863 VDD.n5861 0.0143235
R9018 VDD.n5869 VDD.n5868 0.0143235
R9019 VDD.n5900 VDD.n5899 0.0143235
R9020 VDD.n5910 VDD.n686 0.0143235
R9021 VDD.n5944 VDD.n5943 0.0143235
R9022 VDD.n6060 VDD.n663 0.0143235
R9023 VDD.n5981 VDD.n5980 0.0143235
R9024 VDD.n5991 VDD.n5975 0.0143235
R9025 VDD.n6031 VDD.n6030 0.0143235
R9026 VDD.n6187 VDD.n561 0.0143235
R9027 VDD.n6208 VDD.n559 0.0143235
R9028 VDD.n6227 VDD.n547 0.0143235
R9029 VDD.n6249 VDD.n533 0.0143235
R9030 VDD.n6269 VDD.n522 0.0143235
R9031 VDD.n6315 VDD.n6313 0.0143235
R9032 VDD.n6321 VDD.n6320 0.0143235
R9033 VDD.n6352 VDD.n6351 0.0143235
R9034 VDD.n6358 VDD.n454 0.0143235
R9035 VDD.n6379 VDD.n441 0.0143235
R9036 VDD.n6413 VDD.n427 0.0143235
R9037 VDD.n6434 VDD.n425 0.0143235
R9038 VDD.n6453 VDD.n413 0.0143235
R9039 VDD.n6475 VDD.n399 0.0143235
R9040 VDD.n6495 VDD.n388 0.0143235
R9041 VDD.n6541 VDD.n6539 0.0143235
R9042 VDD.n6547 VDD.n6546 0.0143235
R9043 VDD.n6578 VDD.n6577 0.0143235
R9044 VDD.n6584 VDD.n320 0.0143235
R9045 VDD.n6605 VDD.n307 0.0143235
R9046 VDD.n6639 VDD.n293 0.0143235
R9047 VDD.n6660 VDD.n291 0.0143235
R9048 VDD.n6679 VDD.n279 0.0143235
R9049 VDD.n6701 VDD.n265 0.0143235
R9050 VDD.n6721 VDD.n254 0.0143235
R9051 VDD.n6767 VDD.n6765 0.0143235
R9052 VDD.n6773 VDD.n6772 0.0143235
R9053 VDD.n6804 VDD.n6803 0.0143235
R9054 VDD.n6810 VDD.n186 0.0143235
R9055 VDD.n6831 VDD.n173 0.0143235
R9056 VDD.n6865 VDD.n159 0.0143235
R9057 VDD.n6886 VDD.n157 0.0143235
R9058 VDD.n6905 VDD.n145 0.0143235
R9059 VDD.n6927 VDD.n131 0.0143235
R9060 VDD.n6947 VDD.n120 0.0143235
R9061 VDD.n6993 VDD.n6991 0.0143235
R9062 VDD.n6999 VDD.n6998 0.0143235
R9063 VDD.n7030 VDD.n7029 0.0143235
R9064 VDD.n7036 VDD.n52 0.0143235
R9065 VDD.n7061 VDD.n50 0.0143235
R9066 VDD.n7094 VDD.n7093 0.0143235
R9067 VDD.n7210 VDD.n34 0.0143235
R9068 VDD.n7131 VDD.n7130 0.0143235
R9069 VDD.n7141 VDD.n7125 0.0143235
R9070 VDD.n7181 VDD.n7180 0.0143235
R9071 VDD.n4330 VDD.n2743 0.0143235
R9072 VDD.n2797 VDD.n2788 0.0143235
R9073 VDD.n2804 VDD.n2803 0.0143235
R9074 VDD.n4302 VDD.n4301 0.0143235
R9075 VDD.n2873 VDD.n2872 0.0143235
R9076 VDD.n2901 VDD.n2900 0.0143235
R9077 VDD.n4262 VDD.n4261 0.0143235
R9078 VDD.n2944 VDD.n2943 0.0143235
R9079 VDD.n4241 VDD.n4240 0.0143235
R9080 VDD.n2984 VDD.n2976 0.0143235
R9081 VDD.n3039 VDD.n3030 0.0143235
R9082 VDD.n3046 VDD.n3045 0.0143235
R9083 VDD.n4191 VDD.n4190 0.0143235
R9084 VDD.n3108 VDD.n3098 0.0143235
R9085 VDD.n3115 VDD.n3114 0.0143235
R9086 VDD.n3167 VDD.n3166 0.0143235
R9087 VDD.n4143 VDD.n4142 0.0143235
R9088 VDD.n3210 VDD.n3209 0.0143235
R9089 VDD.n4122 VDD.n4121 0.0143235
R9090 VDD.n3250 VDD.n3242 0.0143235
R9091 VDD.n3305 VDD.n3296 0.0143235
R9092 VDD.n3312 VDD.n3311 0.0143235
R9093 VDD.n4072 VDD.n4071 0.0143235
R9094 VDD.n3374 VDD.n3364 0.0143235
R9095 VDD.n3381 VDD.n3380 0.0143235
R9096 VDD.n3433 VDD.n3432 0.0143235
R9097 VDD.n4024 VDD.n4023 0.0143235
R9098 VDD.n3476 VDD.n3475 0.0143235
R9099 VDD.n4003 VDD.n4002 0.0143235
R9100 VDD.n3516 VDD.n3508 0.0143235
R9101 VDD.n3571 VDD.n3562 0.0143235
R9102 VDD.n3578 VDD.n3577 0.0143235
R9103 VDD.n3953 VDD.n3952 0.0143235
R9104 VDD.n3640 VDD.n3630 0.0143235
R9105 VDD.n3647 VDD.n3646 0.0143235
R9106 VDD.n3699 VDD.n3698 0.0143235
R9107 VDD.n3905 VDD.n3904 0.0143235
R9108 VDD.n3742 VDD.n3741 0.0143235
R9109 VDD.n3884 VDD.n3883 0.0143235
R9110 VDD.n3782 VDD.n3774 0.0143235
R9111 VDD.n4382 VDD.n4381 0.0143235
R9112 VDD.n2671 VDD.n2661 0.0143235
R9113 VDD.n2678 VDD.n2677 0.0143235
R9114 VDD.n4355 VDD.n4354 0.0143235
R9115 VDD.n2724 VDD.n2723 0.0143235
R9116 VDD.n1423 VDD.n1413 0.0143235
R9117 VDD.n1430 VDD.n1429 0.0143235
R9118 VDD.n4853 VDD.n4852 0.0143235
R9119 VDD.n1492 VDD.n1482 0.0143235
R9120 VDD.n1499 VDD.n1498 0.0143235
R9121 VDD.n1548 VDD.n1540 0.0143235
R9122 VDD.n4804 VDD.n4803 0.0143235
R9123 VDD.n1590 VDD.n1582 0.0143235
R9124 VDD.n4782 VDD.n4781 0.0143235
R9125 VDD.n1632 VDD.n1624 0.0143235
R9126 VDD.n1687 VDD.n1678 0.0143235
R9127 VDD.n1694 VDD.n1693 0.0143235
R9128 VDD.n4732 VDD.n4731 0.0143235
R9129 VDD.n1756 VDD.n1746 0.0143235
R9130 VDD.n1763 VDD.n1762 0.0143235
R9131 VDD.n1812 VDD.n1804 0.0143235
R9132 VDD.n4683 VDD.n4682 0.0143235
R9133 VDD.n1854 VDD.n1846 0.0143235
R9134 VDD.n4661 VDD.n4660 0.0143235
R9135 VDD.n1896 VDD.n1888 0.0143235
R9136 VDD.n1951 VDD.n1942 0.0143235
R9137 VDD.n1958 VDD.n1957 0.0143235
R9138 VDD.n4611 VDD.n4610 0.0143235
R9139 VDD.n2020 VDD.n2010 0.0143235
R9140 VDD.n2027 VDD.n2026 0.0143235
R9141 VDD.n2076 VDD.n2068 0.0143235
R9142 VDD.n4562 VDD.n4561 0.0143235
R9143 VDD.n2118 VDD.n2110 0.0143235
R9144 VDD.n4540 VDD.n4539 0.0143235
R9145 VDD.n2160 VDD.n2152 0.0143235
R9146 VDD.n2215 VDD.n2206 0.0143235
R9147 VDD.n2222 VDD.n2221 0.0143235
R9148 VDD.n4490 VDD.n4489 0.0143235
R9149 VDD.n2284 VDD.n2274 0.0143235
R9150 VDD.n2291 VDD.n2290 0.0143235
R9151 VDD.n2340 VDD.n2332 0.0143235
R9152 VDD.n4441 VDD.n4440 0.0143235
R9153 VDD.n2382 VDD.n2374 0.0143235
R9154 VDD.n4419 VDD.n4418 0.0143235
R9155 VDD.n2424 VDD.n2416 0.0143235
R9156 VDD.n1296 VDD.n1262 0.0143235
R9157 VDD.n1303 VDD.n1302 0.0143235
R9158 VDD.n4905 VDD.n4904 0.0143235
R9159 VDD.n1365 VDD.n1355 0.0143235
R9160 VDD.n1372 VDD.n1371 0.0143235
R9161 VDD.n3855 VDD.n3854 0.0140975
R9162 VDD.n2555 VDD.n2554 0.0140975
R9163 VDD.n7263 VDD.n3 0.0140135
R9164 VDD.n6118 VDD.n610 0.0140135
R9165 VDD.n2480 VDD.n2464 0.0140135
R9166 VDD.n4962 VDD.n4936 0.0140135
R9167 VDD.n5938 VDD.n5932 0.0137576
R9168 VDD.n6063 VDD.n6062 0.0137576
R9169 VDD.n6053 VDD.n5953 0.0137576
R9170 VDD.n5989 VDD.n5988 0.0137576
R9171 VDD.n6019 VDD.n6018 0.0137576
R9172 VDD.n5999 VDD.n5998 0.0137576
R9173 VDD.n6201 VDD.n6200 0.0137576
R9174 VDD.n6222 VDD.n6221 0.0137576
R9175 VDD.n6233 VDD.n546 0.0137576
R9176 VDD.n6255 VDD.n532 0.0137576
R9177 VDD.n6275 VDD.n521 0.0137576
R9178 VDD.n6311 VDD.n488 0.0137576
R9179 VDD.n6326 VDD.n481 0.0137576
R9180 VDD.n6346 VDD.n475 0.0137576
R9181 VDD.n6361 VDD.n6360 0.0137576
R9182 VDD.n6381 VDD.n451 0.0137576
R9183 VDD.n6405 VDD.n438 0.0137576
R9184 VDD.n6407 VDD.n6406 0.0137576
R9185 VDD.n6427 VDD.n6426 0.0137576
R9186 VDD.n6448 VDD.n6447 0.0137576
R9187 VDD.n6459 VDD.n412 0.0137576
R9188 VDD.n6481 VDD.n398 0.0137576
R9189 VDD.n6501 VDD.n387 0.0137576
R9190 VDD.n6537 VDD.n354 0.0137576
R9191 VDD.n6552 VDD.n347 0.0137576
R9192 VDD.n6572 VDD.n341 0.0137576
R9193 VDD.n6587 VDD.n6586 0.0137576
R9194 VDD.n6607 VDD.n317 0.0137576
R9195 VDD.n6631 VDD.n304 0.0137576
R9196 VDD.n6633 VDD.n6632 0.0137576
R9197 VDD.n6653 VDD.n6652 0.0137576
R9198 VDD.n6674 VDD.n6673 0.0137576
R9199 VDD.n6685 VDD.n278 0.0137576
R9200 VDD.n6707 VDD.n264 0.0137576
R9201 VDD.n6727 VDD.n253 0.0137576
R9202 VDD.n6763 VDD.n220 0.0137576
R9203 VDD.n6778 VDD.n213 0.0137576
R9204 VDD.n6798 VDD.n207 0.0137576
R9205 VDD.n6813 VDD.n6812 0.0137576
R9206 VDD.n6833 VDD.n183 0.0137576
R9207 VDD.n6857 VDD.n170 0.0137576
R9208 VDD.n6859 VDD.n6858 0.0137576
R9209 VDD.n6879 VDD.n6878 0.0137576
R9210 VDD.n6900 VDD.n6899 0.0137576
R9211 VDD.n6911 VDD.n144 0.0137576
R9212 VDD.n6933 VDD.n130 0.0137576
R9213 VDD.n6953 VDD.n119 0.0137576
R9214 VDD.n6989 VDD.n86 0.0137576
R9215 VDD.n7004 VDD.n79 0.0137576
R9216 VDD.n7024 VDD.n73 0.0137576
R9217 VDD.n7039 VDD.n7038 0.0137576
R9218 VDD.n7063 VDD.n48 0.0137576
R9219 VDD.n7088 VDD.n7082 0.0137576
R9220 VDD.n7213 VDD.n7212 0.0137576
R9221 VDD.n7203 VDD.n7103 0.0137576
R9222 VDD.n7139 VDD.n7138 0.0137576
R9223 VDD.n7169 VDD.n7168 0.0137576
R9224 VDD.n7149 VDD.n7148 0.0137576
R9225 VDD.n4388 VDD.n2431 0.0137576
R9226 VDD.n4379 VDD.n4378 0.0137576
R9227 VDD.n2669 VDD.n2668 0.0137576
R9228 VDD.n4361 VDD.n2649 0.0137576
R9229 VDD.n4352 VDD.n4351 0.0137576
R9230 VDD.n2731 VDD.n2730 0.0137576
R9231 VDD.n1421 VDD.n1420 0.0137576
R9232 VDD.n4859 VDD.n1402 0.0137576
R9233 VDD.n4850 VDD.n4849 0.0137576
R9234 VDD.n1490 VDD.n1489 0.0137576
R9235 VDD.n4832 VDD.n1470 0.0137576
R9236 VDD.n1546 VDD.n1545 0.0137576
R9237 VDD.n1565 VDD.n1564 0.0137576
R9238 VDD.n1588 VDD.n1587 0.0137576
R9239 VDD.n1607 VDD.n1606 0.0137576
R9240 VDD.n1630 VDD.n1629 0.0137576
R9241 VDD.n1644 VDD.n1643 0.0137576
R9242 VDD.n1642 VDD.n1639 0.0137576
R9243 VDD.n1685 VDD.n1684 0.0137576
R9244 VDD.n4738 VDD.n1670 0.0137576
R9245 VDD.n4729 VDD.n4728 0.0137576
R9246 VDD.n1754 VDD.n1753 0.0137576
R9247 VDD.n4711 VDD.n1734 0.0137576
R9248 VDD.n1810 VDD.n1809 0.0137576
R9249 VDD.n1829 VDD.n1828 0.0137576
R9250 VDD.n1852 VDD.n1851 0.0137576
R9251 VDD.n1871 VDD.n1870 0.0137576
R9252 VDD.n1894 VDD.n1893 0.0137576
R9253 VDD.n1908 VDD.n1907 0.0137576
R9254 VDD.n1906 VDD.n1903 0.0137576
R9255 VDD.n1949 VDD.n1948 0.0137576
R9256 VDD.n4617 VDD.n1934 0.0137576
R9257 VDD.n4608 VDD.n4607 0.0137576
R9258 VDD.n2018 VDD.n2017 0.0137576
R9259 VDD.n4590 VDD.n1998 0.0137576
R9260 VDD.n2074 VDD.n2073 0.0137576
R9261 VDD.n2093 VDD.n2092 0.0137576
R9262 VDD.n2116 VDD.n2115 0.0137576
R9263 VDD.n2135 VDD.n2134 0.0137576
R9264 VDD.n2158 VDD.n2157 0.0137576
R9265 VDD.n2172 VDD.n2171 0.0137576
R9266 VDD.n2170 VDD.n2167 0.0137576
R9267 VDD.n2213 VDD.n2212 0.0137576
R9268 VDD.n4496 VDD.n2198 0.0137576
R9269 VDD.n4487 VDD.n4486 0.0137576
R9270 VDD.n2282 VDD.n2281 0.0137576
R9271 VDD.n4469 VDD.n2262 0.0137576
R9272 VDD.n2338 VDD.n2337 0.0137576
R9273 VDD.n2357 VDD.n2356 0.0137576
R9274 VDD.n2380 VDD.n2379 0.0137576
R9275 VDD.n2399 VDD.n2398 0.0137576
R9276 VDD.n2422 VDD.n2421 0.0137576
R9277 VDD.n1277 VDD.n1276 0.0137576
R9278 VDD.n1294 VDD.n1293 0.0137576
R9279 VDD.n4911 VDD.n1254 0.0137576
R9280 VDD.n4902 VDD.n4901 0.0137576
R9281 VDD.n1363 VDD.n1362 0.0137576
R9282 VDD.n4884 VDD.n1343 0.0137576
R9283 VDD.n2764 VDD.n2748 0.0137576
R9284 VDD.n2795 VDD.n2794 0.0137576
R9285 VDD.n4308 VDD.n2780 0.0137576
R9286 VDD.n4299 VDD.n4298 0.0137576
R9287 VDD.n2882 VDD.n2881 0.0137576
R9288 VDD.n2898 VDD.n2897 0.0137576
R9289 VDD.n2916 VDD.n2858 0.0137576
R9290 VDD.n2941 VDD.n2940 0.0137576
R9291 VDD.n2959 VDD.n2933 0.0137576
R9292 VDD.n2982 VDD.n2981 0.0137576
R9293 VDD.n2996 VDD.n2995 0.0137576
R9294 VDD.n2994 VDD.n2991 0.0137576
R9295 VDD.n3037 VDD.n3036 0.0137576
R9296 VDD.n4197 VDD.n3022 0.0137576
R9297 VDD.n4188 VDD.n4187 0.0137576
R9298 VDD.n3106 VDD.n3105 0.0137576
R9299 VDD.n4170 VDD.n3086 0.0137576
R9300 VDD.n3164 VDD.n3163 0.0137576
R9301 VDD.n3182 VDD.n3156 0.0137576
R9302 VDD.n3207 VDD.n3206 0.0137576
R9303 VDD.n3225 VDD.n3199 0.0137576
R9304 VDD.n3248 VDD.n3247 0.0137576
R9305 VDD.n3262 VDD.n3261 0.0137576
R9306 VDD.n3260 VDD.n3257 0.0137576
R9307 VDD.n3303 VDD.n3302 0.0137576
R9308 VDD.n4078 VDD.n3288 0.0137576
R9309 VDD.n4069 VDD.n4068 0.0137576
R9310 VDD.n3372 VDD.n3371 0.0137576
R9311 VDD.n4051 VDD.n3352 0.0137576
R9312 VDD.n3430 VDD.n3429 0.0137576
R9313 VDD.n3448 VDD.n3422 0.0137576
R9314 VDD.n3473 VDD.n3472 0.0137576
R9315 VDD.n3491 VDD.n3465 0.0137576
R9316 VDD.n3514 VDD.n3513 0.0137576
R9317 VDD.n3528 VDD.n3527 0.0137576
R9318 VDD.n3526 VDD.n3523 0.0137576
R9319 VDD.n3569 VDD.n3568 0.0137576
R9320 VDD.n3959 VDD.n3554 0.0137576
R9321 VDD.n3950 VDD.n3949 0.0137576
R9322 VDD.n3638 VDD.n3637 0.0137576
R9323 VDD.n3932 VDD.n3618 0.0137576
R9324 VDD.n3696 VDD.n3695 0.0137576
R9325 VDD.n3714 VDD.n3688 0.0137576
R9326 VDD.n3739 VDD.n3738 0.0137576
R9327 VDD.n3757 VDD.n3731 0.0137576
R9328 VDD.n3780 VDD.n3779 0.0137576
R9329 VDD.n5035 VDD.n1193 0.0137576
R9330 VDD.n5065 VDD.n1181 0.0137576
R9331 VDD.n5083 VDD.n5082 0.0137576
R9332 VDD.n5094 VDD.n1167 0.0137576
R9333 VDD.n5118 VDD.n1153 0.0137576
R9334 VDD.n5145 VDD.n1119 0.0137576
R9335 VDD.n5165 VDD.n1113 0.0137576
R9336 VDD.n5180 VDD.n5179 0.0137576
R9337 VDD.n5201 VDD.n1086 0.0137576
R9338 VDD.n5221 VDD.n1079 0.0137576
R9339 VDD.n5240 VDD.n5239 0.0137576
R9340 VDD.n1071 VDD.n1070 0.0137576
R9341 VDD.n5263 VDD.n1058 0.0137576
R9342 VDD.n5293 VDD.n1046 0.0137576
R9343 VDD.n5311 VDD.n5310 0.0137576
R9344 VDD.n5322 VDD.n1032 0.0137576
R9345 VDD.n5346 VDD.n1018 0.0137576
R9346 VDD.n5373 VDD.n984 0.0137576
R9347 VDD.n5393 VDD.n978 0.0137576
R9348 VDD.n5408 VDD.n5407 0.0137576
R9349 VDD.n5429 VDD.n951 0.0137576
R9350 VDD.n5449 VDD.n944 0.0137576
R9351 VDD.n5468 VDD.n5467 0.0137576
R9352 VDD.n936 VDD.n935 0.0137576
R9353 VDD.n5491 VDD.n923 0.0137576
R9354 VDD.n5521 VDD.n911 0.0137576
R9355 VDD.n5539 VDD.n5538 0.0137576
R9356 VDD.n5550 VDD.n897 0.0137576
R9357 VDD.n5574 VDD.n883 0.0137576
R9358 VDD.n5601 VDD.n849 0.0137576
R9359 VDD.n5621 VDD.n843 0.0137576
R9360 VDD.n5636 VDD.n5635 0.0137576
R9361 VDD.n5657 VDD.n816 0.0137576
R9362 VDD.n5677 VDD.n809 0.0137576
R9363 VDD.n5696 VDD.n5695 0.0137576
R9364 VDD.n801 VDD.n800 0.0137576
R9365 VDD.n5719 VDD.n788 0.0137576
R9366 VDD.n5749 VDD.n776 0.0137576
R9367 VDD.n5767 VDD.n5766 0.0137576
R9368 VDD.n5778 VDD.n762 0.0137576
R9369 VDD.n5801 VDD.n748 0.0137576
R9370 VDD.n5834 VDD.n722 0.0137576
R9371 VDD.n5859 VDD.n705 0.0137576
R9372 VDD.n5874 VDD.n698 0.0137576
R9373 VDD.n5894 VDD.n692 0.0137576
R9374 VDD.n5913 VDD.n5912 0.0137576
R9375 VDD.n595 VDD.n591 0.0137243
R9376 VDD.n3839 VDD.n3835 0.0137243
R9377 VDD.n2515 VDD.n2511 0.0137243
R9378 VDD.n1225 VDD.n1221 0.0137243
R9379 VDD.n6117 VDD.n612 0.0137188
R9380 VDD.n6117 VDD.n6116 0.0137188
R9381 VDD.n2609 VDD.n2463 0.0137188
R9382 VDD.n2609 VDD.n2461 0.0137188
R9383 VDD.n4945 VDD.n4944 0.0137188
R9384 VDD.n4945 VDD.n4937 0.0137188
R9385 VDD.n7262 VDD.n7243 0.0137188
R9386 VDD.n7262 VDD.n7261 0.0137188
R9387 VDD.n2587 VDD.n2586 0.0134306
R9388 VDD.n4395 VDD.n2427 0.0133585
R9389 VDD.n6086 VDD.n633 0.0130393
R9390 VDD.n6113 VDD.n600 0.0130393
R9391 VDD.n2613 VDD.n2458 0.0130393
R9392 VDD.n2605 VDD.n2469 0.0130393
R9393 VDD.n4949 VDD.n4938 0.0130393
R9394 VDD.n4976 VDD.n1233 0.0130393
R9395 VDD.n7241 VDD.n7240 0.0130393
R9396 VDD.n7259 VDD.n7258 0.0130393
R9397 VDD.n3858 VDD.n3857 0.0129151
R9398 VDD.n2547 VDD.n2546 0.0129151
R9399 VDD.n2588 VDD 0.0108445
R9400 VDD.n597 VDD.n592 0.0105714
R9401 VDD.n3841 VDD.n3834 0.0105714
R9402 VDD.n3841 VDD.n3836 0.0105714
R9403 VDD.n2517 VDD.n2510 0.0105714
R9404 VDD.n2517 VDD.n2512 0.0105714
R9405 VDD.n1227 VDD.n1222 0.0105714
R9406 VDD.n2607 VDD.n2465 0.0105072
R9407 VDD.n6108 VDD.n618 0.0103794
R9408 VDD.n625 VDD.n624 0.0103794
R9409 VDD.n6100 VDD.n629 0.0103794
R9410 VDD.n6153 VDD.n6152 0.0103794
R9411 VDD.n6164 VDD.n578 0.0103794
R9412 VDD.n6144 VDD.n6143 0.0103794
R9413 VDD.n586 VDD.n585 0.0103794
R9414 VDD.n6172 VDD.n572 0.0103794
R9415 VDD.n5011 VDD.n1202 0.0103794
R9416 VDD.n4996 VDD.n4995 0.0103794
R9417 VDD.n5003 VDD.n1208 0.0103794
R9418 VDD.n4987 VDD.n4986 0.0103794
R9419 VDD.n1216 VDD.n1215 0.0103794
R9420 VDD.n5038 VDD.n5037 0.0099697
R9421 VDD.n5068 VDD.n5067 0.0099697
R9422 VDD.n5080 VDD.n5079 0.0099697
R9423 VDD.n5095 VDD.n1166 0.0099697
R9424 VDD.n5121 VDD.n5120 0.0099697
R9425 VDD.n1146 VDD.n1145 0.0099697
R9426 VDD.n1133 VDD.n1132 0.0099697
R9427 VDD.n5147 VDD.n1118 0.0099697
R9428 VDD.n5163 VDD.n5160 0.0099697
R9429 VDD.n1104 VDD.n1103 0.0099697
R9430 VDD.n5205 VDD.n1085 0.0099697
R9431 VDD.n5219 VDD.n5216 0.0099697
R9432 VDD.n5266 VDD.n5265 0.0099697
R9433 VDD.n5296 VDD.n5295 0.0099697
R9434 VDD.n5308 VDD.n5307 0.0099697
R9435 VDD.n5323 VDD.n1031 0.0099697
R9436 VDD.n5349 VDD.n5348 0.0099697
R9437 VDD.n1011 VDD.n1010 0.0099697
R9438 VDD.n998 VDD.n997 0.0099697
R9439 VDD.n5375 VDD.n983 0.0099697
R9440 VDD.n5391 VDD.n5388 0.0099697
R9441 VDD.n969 VDD.n968 0.0099697
R9442 VDD.n5433 VDD.n950 0.0099697
R9443 VDD.n5447 VDD.n5444 0.0099697
R9444 VDD.n5494 VDD.n5493 0.0099697
R9445 VDD.n5524 VDD.n5523 0.0099697
R9446 VDD.n5536 VDD.n5535 0.0099697
R9447 VDD.n5551 VDD.n896 0.0099697
R9448 VDD.n5577 VDD.n5576 0.0099697
R9449 VDD.n876 VDD.n875 0.0099697
R9450 VDD.n863 VDD.n862 0.0099697
R9451 VDD.n5603 VDD.n848 0.0099697
R9452 VDD.n5619 VDD.n5616 0.0099697
R9453 VDD.n834 VDD.n833 0.0099697
R9454 VDD.n5661 VDD.n815 0.0099697
R9455 VDD.n5675 VDD.n5672 0.0099697
R9456 VDD.n5722 VDD.n5721 0.0099697
R9457 VDD.n5752 VDD.n5751 0.0099697
R9458 VDD.n5764 VDD.n5763 0.0099697
R9459 VDD.n5779 VDD.n761 0.0099697
R9460 VDD.n5804 VDD.n5803 0.0099697
R9461 VDD.n741 VDD.n740 0.0099697
R9462 VDD.n737 VDD.n736 0.0099697
R9463 VDD.n5832 VDD.n5831 0.0099697
R9464 VDD.n5857 VDD.n5856 0.0099697
R9465 VDD.n5876 VDD.n697 0.0099697
R9466 VDD.n5892 VDD.n5889 0.0099697
R9467 VDD.n681 VDD.n680 0.0099697
R9468 VDD.n5936 VDD.n5933 0.0099697
R9469 VDD.n5960 VDD.n659 0.0099697
R9470 VDD.n6051 VDD.n5955 0.0099697
R9471 VDD.n6040 VDD.n5971 0.0099697
R9472 VDD.n6022 VDD.n6021 0.0099697
R9473 VDD.n6198 VDD.n6197 0.0099697
R9474 VDD.n6219 VDD.n6218 0.0099697
R9475 VDD.n6234 VDD.n545 0.0099697
R9476 VDD.n6258 VDD.n6257 0.0099697
R9477 VDD.n6278 VDD.n6277 0.0099697
R9478 VDD.n514 VDD.n513 0.0099697
R9479 VDD.n510 VDD.n509 0.0099697
R9480 VDD.n6309 VDD.n6308 0.0099697
R9481 VDD.n6328 VDD.n480 0.0099697
R9482 VDD.n6344 VDD.n6341 0.0099697
R9483 VDD.n466 VDD.n465 0.0099697
R9484 VDD.n6384 VDD.n6383 0.0099697
R9485 VDD.n6424 VDD.n6423 0.0099697
R9486 VDD.n6445 VDD.n6444 0.0099697
R9487 VDD.n6460 VDD.n411 0.0099697
R9488 VDD.n6484 VDD.n6483 0.0099697
R9489 VDD.n6504 VDD.n6503 0.0099697
R9490 VDD.n380 VDD.n379 0.0099697
R9491 VDD.n376 VDD.n375 0.0099697
R9492 VDD.n6535 VDD.n6534 0.0099697
R9493 VDD.n6554 VDD.n346 0.0099697
R9494 VDD.n6570 VDD.n6567 0.0099697
R9495 VDD.n332 VDD.n331 0.0099697
R9496 VDD.n6610 VDD.n6609 0.0099697
R9497 VDD.n6650 VDD.n6649 0.0099697
R9498 VDD.n6671 VDD.n6670 0.0099697
R9499 VDD.n6686 VDD.n277 0.0099697
R9500 VDD.n6710 VDD.n6709 0.0099697
R9501 VDD.n6730 VDD.n6729 0.0099697
R9502 VDD.n246 VDD.n245 0.0099697
R9503 VDD.n242 VDD.n241 0.0099697
R9504 VDD.n6761 VDD.n6760 0.0099697
R9505 VDD.n6780 VDD.n212 0.0099697
R9506 VDD.n6796 VDD.n6793 0.0099697
R9507 VDD.n198 VDD.n197 0.0099697
R9508 VDD.n6836 VDD.n6835 0.0099697
R9509 VDD.n6876 VDD.n6875 0.0099697
R9510 VDD.n6897 VDD.n6896 0.0099697
R9511 VDD.n6912 VDD.n143 0.0099697
R9512 VDD.n6936 VDD.n6935 0.0099697
R9513 VDD.n6956 VDD.n6955 0.0099697
R9514 VDD.n112 VDD.n111 0.0099697
R9515 VDD.n108 VDD.n107 0.0099697
R9516 VDD.n6987 VDD.n6986 0.0099697
R9517 VDD.n7006 VDD.n78 0.0099697
R9518 VDD.n7022 VDD.n7019 0.0099697
R9519 VDD.n64 VDD.n63 0.0099697
R9520 VDD.n7067 VDD.n7066 0.0099697
R9521 VDD.n7086 VDD.n7083 0.0099697
R9522 VDD.n7110 VDD.n30 0.0099697
R9523 VDD.n7201 VDD.n7105 0.0099697
R9524 VDD.n7190 VDD.n7121 0.0099697
R9525 VDD.n7172 VDD.n7171 0.0099697
R9526 VDD.n2767 VDD.n2766 0.0099697
R9527 VDD.n2791 VDD.n2790 0.0099697
R9528 VDD.n4310 VDD.n2779 0.0099697
R9529 VDD.n2831 VDD.n2811 0.0099697
R9530 VDD.n2879 VDD.n2878 0.0099697
R9531 VDD.n4283 VDD.n2843 0.0099697
R9532 VDD.n4282 VDD.n4281 0.0099697
R9533 VDD.n4270 VDD.n2854 0.0099697
R9534 VDD.n2919 VDD.n2918 0.0099697
R9535 VDD.n4249 VDD.n2929 0.0099697
R9536 VDD.n2962 VDD.n2961 0.0099697
R9537 VDD.n4228 VDD.n2972 0.0099697
R9538 VDD.n3033 VDD.n3032 0.0099697
R9539 VDD.n4199 VDD.n3021 0.0099697
R9540 VDD.n3073 VDD.n3053 0.0099697
R9541 VDD.n3102 VDD.n3101 0.0099697
R9542 VDD.n4172 VDD.n3085 0.0099697
R9543 VDD.n3140 VDD.n3135 0.0099697
R9544 VDD.n3139 VDD.n3138 0.0099697
R9545 VDD.n4151 VDD.n3152 0.0099697
R9546 VDD.n3185 VDD.n3184 0.0099697
R9547 VDD.n4130 VDD.n3195 0.0099697
R9548 VDD.n3228 VDD.n3227 0.0099697
R9549 VDD.n4109 VDD.n3238 0.0099697
R9550 VDD.n3299 VDD.n3298 0.0099697
R9551 VDD.n4080 VDD.n3287 0.0099697
R9552 VDD.n3339 VDD.n3319 0.0099697
R9553 VDD.n3368 VDD.n3367 0.0099697
R9554 VDD.n4053 VDD.n3351 0.0099697
R9555 VDD.n3406 VDD.n3401 0.0099697
R9556 VDD.n3405 VDD.n3404 0.0099697
R9557 VDD.n4032 VDD.n3418 0.0099697
R9558 VDD.n3451 VDD.n3450 0.0099697
R9559 VDD.n4011 VDD.n3461 0.0099697
R9560 VDD.n3494 VDD.n3493 0.0099697
R9561 VDD.n3990 VDD.n3504 0.0099697
R9562 VDD.n3565 VDD.n3564 0.0099697
R9563 VDD.n3961 VDD.n3553 0.0099697
R9564 VDD.n3605 VDD.n3585 0.0099697
R9565 VDD.n3634 VDD.n3633 0.0099697
R9566 VDD.n3934 VDD.n3617 0.0099697
R9567 VDD.n3672 VDD.n3667 0.0099697
R9568 VDD.n3671 VDD.n3670 0.0099697
R9569 VDD.n3913 VDD.n3684 0.0099697
R9570 VDD.n3717 VDD.n3716 0.0099697
R9571 VDD.n3892 VDD.n3727 0.0099697
R9572 VDD.n3760 VDD.n3759 0.0099697
R9573 VDD.n3871 VDD.n3770 0.0099697
R9574 VDD.n2636 VDD.n2442 0.0099697
R9575 VDD.n2665 VDD.n2664 0.0099697
R9576 VDD.n4363 VDD.n2648 0.0099697
R9577 VDD.n2705 VDD.n2685 0.0099697
R9578 VDD.n2728 VDD.n2727 0.0099697
R9579 VDD.n1417 VDD.n1416 0.0099697
R9580 VDD.n4861 VDD.n1401 0.0099697
R9581 VDD.n1457 VDD.n1437 0.0099697
R9582 VDD.n1486 VDD.n1485 0.0099697
R9583 VDD.n4834 VDD.n1469 0.0099697
R9584 VDD.n1524 VDD.n1519 0.0099697
R9585 VDD.n1523 VDD.n1522 0.0099697
R9586 VDD.n4813 VDD.n1536 0.0099697
R9587 VDD.n1568 VDD.n1567 0.0099697
R9588 VDD.n4791 VDD.n1578 0.0099697
R9589 VDD.n1610 VDD.n1609 0.0099697
R9590 VDD.n4769 VDD.n1620 0.0099697
R9591 VDD.n1681 VDD.n1680 0.0099697
R9592 VDD.n4740 VDD.n1669 0.0099697
R9593 VDD.n1721 VDD.n1701 0.0099697
R9594 VDD.n1750 VDD.n1749 0.0099697
R9595 VDD.n4713 VDD.n1733 0.0099697
R9596 VDD.n1788 VDD.n1783 0.0099697
R9597 VDD.n1787 VDD.n1786 0.0099697
R9598 VDD.n4692 VDD.n1800 0.0099697
R9599 VDD.n1832 VDD.n1831 0.0099697
R9600 VDD.n4670 VDD.n1842 0.0099697
R9601 VDD.n1874 VDD.n1873 0.0099697
R9602 VDD.n4648 VDD.n1884 0.0099697
R9603 VDD.n1945 VDD.n1944 0.0099697
R9604 VDD.n4619 VDD.n1933 0.0099697
R9605 VDD.n1985 VDD.n1965 0.0099697
R9606 VDD.n2014 VDD.n2013 0.0099697
R9607 VDD.n4592 VDD.n1997 0.0099697
R9608 VDD.n2052 VDD.n2047 0.0099697
R9609 VDD.n2051 VDD.n2050 0.0099697
R9610 VDD.n4571 VDD.n2064 0.0099697
R9611 VDD.n2096 VDD.n2095 0.0099697
R9612 VDD.n4549 VDD.n2106 0.0099697
R9613 VDD.n2138 VDD.n2137 0.0099697
R9614 VDD.n4527 VDD.n2148 0.0099697
R9615 VDD.n2209 VDD.n2208 0.0099697
R9616 VDD.n4498 VDD.n2197 0.0099697
R9617 VDD.n2249 VDD.n2229 0.0099697
R9618 VDD.n2278 VDD.n2277 0.0099697
R9619 VDD.n4471 VDD.n2261 0.0099697
R9620 VDD.n2316 VDD.n2311 0.0099697
R9621 VDD.n2315 VDD.n2314 0.0099697
R9622 VDD.n4450 VDD.n2328 0.0099697
R9623 VDD.n2360 VDD.n2359 0.0099697
R9624 VDD.n4428 VDD.n2370 0.0099697
R9625 VDD.n2402 VDD.n2401 0.0099697
R9626 VDD.n4406 VDD.n2412 0.0099697
R9627 VDD.n1290 VDD.n1289 0.0099697
R9628 VDD.n4913 VDD.n1253 0.0099697
R9629 VDD.n1330 VDD.n1310 0.0099697
R9630 VDD.n1359 VDD.n1358 0.0099697
R9631 VDD.n4886 VDD.n1342 0.0099697
R9632 VDD.n3804 VDD.n3803 0.00993793
R9633 VDD.n3812 VDD.n3799 0.00993793
R9634 VDD.n3815 VDD.n3795 0.00993793
R9635 VDD.n3809 VDD.n3791 0.00993793
R9636 VDD.n3805 VDD.n3787 0.00993793
R9637 VDD.n2579 VDD.n2578 0.00993793
R9638 VDD.n2573 VDD.n2572 0.00993793
R9639 VDD.n2568 VDD.n2567 0.00993793
R9640 VDD.n2534 VDD.n2533 0.00993793
R9641 VDD.n2501 VDD.n2500 0.00993793
R9642 VDD.n2495 VDD.n2494 0.00993793
R9643 VDD.n2490 VDD.n2489 0.00993793
R9644 VDD.n2549 VDD.n2548 0.00993793
R9645 VDD.n7156 VDD.n7152 0.00926684
R9646 VDD.n6006 VDD.n6002 0.00926684
R9647 VDD.n6136 VDD.n599 0.00895742
R9648 VDD.n1269 VDD 0.0089359
R9649 VDD VDD.n2435 0.0089359
R9650 VDD.n6186 VDD.n6185 0.00792105
R9651 VDD.n6250 VDD.n534 0.00792105
R9652 VDD.n6412 VDD.n6411 0.00792105
R9653 VDD.n6476 VDD.n400 0.00792105
R9654 VDD.n6638 VDD.n6637 0.00792105
R9655 VDD.n6702 VDD.n266 0.00792105
R9656 VDD.n6864 VDD.n6863 0.00792105
R9657 VDD.n6928 VDD.n132 0.00792105
R9658 VDD.n5030 VDD.n1195 0.00792105
R9659 VDD.n5089 VDD.n1169 0.00792105
R9660 VDD.n5258 VDD.n1060 0.00792105
R9661 VDD.n5317 VDD.n1034 0.00792105
R9662 VDD.n5486 VDD.n925 0.00792105
R9663 VDD.n5545 VDD.n899 0.00792105
R9664 VDD.n5714 VDD.n790 0.00792105
R9665 VDD.n5773 VDD.n764 0.00792105
R9666 VDD.n6207 VDD.n6205 0.00792105
R9667 VDD.n6228 VDD.n548 0.00792105
R9668 VDD.n6270 VDD.n523 0.00792105
R9669 VDD.n6289 VDD.n501 0.00792105
R9670 VDD.n6291 VDD.n486 0.00792105
R9671 VDD.n6323 VDD.n6322 0.00792105
R9672 VDD.n6350 VDD.n6349 0.00792105
R9673 VDD.n6357 VDD.n6356 0.00792105
R9674 VDD.n6378 VDD.n6377 0.00792105
R9675 VDD.n6402 VDD.n6401 0.00792105
R9676 VDD.n6433 VDD.n6431 0.00792105
R9677 VDD.n6454 VDD.n414 0.00792105
R9678 VDD.n6496 VDD.n389 0.00792105
R9679 VDD.n6515 VDD.n367 0.00792105
R9680 VDD.n6517 VDD.n352 0.00792105
R9681 VDD.n6549 VDD.n6548 0.00792105
R9682 VDD.n6576 VDD.n6575 0.00792105
R9683 VDD.n6583 VDD.n6582 0.00792105
R9684 VDD.n6604 VDD.n6603 0.00792105
R9685 VDD.n6628 VDD.n6627 0.00792105
R9686 VDD.n6659 VDD.n6657 0.00792105
R9687 VDD.n6680 VDD.n280 0.00792105
R9688 VDD.n6722 VDD.n255 0.00792105
R9689 VDD.n6741 VDD.n233 0.00792105
R9690 VDD.n6743 VDD.n218 0.00792105
R9691 VDD.n6775 VDD.n6774 0.00792105
R9692 VDD.n6802 VDD.n6801 0.00792105
R9693 VDD.n6809 VDD.n6808 0.00792105
R9694 VDD.n6830 VDD.n6829 0.00792105
R9695 VDD.n6854 VDD.n6853 0.00792105
R9696 VDD.n6885 VDD.n6883 0.00792105
R9697 VDD.n6906 VDD.n146 0.00792105
R9698 VDD.n6948 VDD.n121 0.00792105
R9699 VDD.n6967 VDD.n99 0.00792105
R9700 VDD.n6969 VDD.n84 0.00792105
R9701 VDD.n7001 VDD.n7000 0.00792105
R9702 VDD.n7028 VDD.n7027 0.00792105
R9703 VDD.n7035 VDD.n7034 0.00792105
R9704 VDD.n7060 VDD.n7055 0.00792105
R9705 VDD.n7076 VDD.n39 0.00792105
R9706 VDD.n5051 VDD.n1184 0.00792105
R9707 VDD.n5057 VDD.n5055 0.00792105
R9708 VDD.n5112 VDD.n1155 0.00792105
R9709 VDD.n5114 VDD.n1124 0.00792105
R9710 VDD.n5142 VDD.n5141 0.00792105
R9711 VDD.n5169 VDD.n5168 0.00792105
R9712 VDD.n5176 VDD.n5175 0.00792105
R9713 VDD.n5198 VDD.n5196 0.00792105
R9714 VDD.n5225 VDD.n5224 0.00792105
R9715 VDD.n5236 VDD.n5231 0.00792105
R9716 VDD.n5279 VDD.n1049 0.00792105
R9717 VDD.n5285 VDD.n5283 0.00792105
R9718 VDD.n5340 VDD.n1020 0.00792105
R9719 VDD.n5342 VDD.n989 0.00792105
R9720 VDD.n5370 VDD.n5369 0.00792105
R9721 VDD.n5397 VDD.n5396 0.00792105
R9722 VDD.n5404 VDD.n5403 0.00792105
R9723 VDD.n5426 VDD.n5424 0.00792105
R9724 VDD.n5453 VDD.n5452 0.00792105
R9725 VDD.n5464 VDD.n5459 0.00792105
R9726 VDD.n5507 VDD.n914 0.00792105
R9727 VDD.n5513 VDD.n5511 0.00792105
R9728 VDD.n5568 VDD.n885 0.00792105
R9729 VDD.n5570 VDD.n854 0.00792105
R9730 VDD.n5598 VDD.n5597 0.00792105
R9731 VDD.n5625 VDD.n5624 0.00792105
R9732 VDD.n5632 VDD.n5631 0.00792105
R9733 VDD.n5654 VDD.n5652 0.00792105
R9734 VDD.n5681 VDD.n5680 0.00792105
R9735 VDD.n5692 VDD.n5687 0.00792105
R9736 VDD.n5735 VDD.n779 0.00792105
R9737 VDD.n5741 VDD.n5739 0.00792105
R9738 VDD.n5796 VDD.n750 0.00792105
R9739 VDD.n5816 VDD.n728 0.00792105
R9740 VDD.n5837 VDD.n720 0.00792105
R9741 VDD.n5839 VDD.n703 0.00792105
R9742 VDD.n5871 VDD.n5870 0.00792105
R9743 VDD.n5898 VDD.n5897 0.00792105
R9744 VDD.n5909 VDD.n5904 0.00792105
R9745 VDD.n5926 VDD.n668 0.00792105
R9746 VDD.n1410 VDD.n1409 0.00784375
R9747 VDD.n1426 VDD.n1407 0.00784375
R9748 VDD.n4855 VDD.n4854 0.00784375
R9749 VDD.n1479 VDD.n1477 0.00784375
R9750 VDD.n1495 VDD.n1475 0.00784375
R9751 VDD.n4828 VDD.n4827 0.00784375
R9752 VDD.n1549 VDD.n1543 0.00784375
R9753 VDD.n4806 VDD.n4805 0.00784375
R9754 VDD.n1591 VDD.n1585 0.00784375
R9755 VDD.n4784 VDD.n4783 0.00784375
R9756 VDD.n1633 VDD.n1627 0.00784375
R9757 VDD.n4762 VDD.n4761 0.00784375
R9758 VDD.n1677 VDD.n1637 0.00784375
R9759 VDD.n1690 VDD.n1675 0.00784375
R9760 VDD.n4734 VDD.n4733 0.00784375
R9761 VDD.n1743 VDD.n1741 0.00784375
R9762 VDD.n1759 VDD.n1739 0.00784375
R9763 VDD.n4707 VDD.n4706 0.00784375
R9764 VDD.n1813 VDD.n1807 0.00784375
R9765 VDD.n4685 VDD.n4684 0.00784375
R9766 VDD.n1855 VDD.n1849 0.00784375
R9767 VDD.n4663 VDD.n4662 0.00784375
R9768 VDD.n1897 VDD.n1891 0.00784375
R9769 VDD.n4641 VDD.n4640 0.00784375
R9770 VDD.n1941 VDD.n1901 0.00784375
R9771 VDD.n1954 VDD.n1939 0.00784375
R9772 VDD.n4613 VDD.n4612 0.00784375
R9773 VDD.n2007 VDD.n2005 0.00784375
R9774 VDD.n2023 VDD.n2003 0.00784375
R9775 VDD.n4586 VDD.n4585 0.00784375
R9776 VDD.n2077 VDD.n2071 0.00784375
R9777 VDD.n4564 VDD.n4563 0.00784375
R9778 VDD.n2119 VDD.n2113 0.00784375
R9779 VDD.n4542 VDD.n4541 0.00784375
R9780 VDD.n2161 VDD.n2155 0.00784375
R9781 VDD.n4520 VDD.n4519 0.00784375
R9782 VDD.n2205 VDD.n2165 0.00784375
R9783 VDD.n2218 VDD.n2203 0.00784375
R9784 VDD.n4492 VDD.n4491 0.00784375
R9785 VDD.n2271 VDD.n2269 0.00784375
R9786 VDD.n2287 VDD.n2267 0.00784375
R9787 VDD.n4465 VDD.n4464 0.00784375
R9788 VDD.n2341 VDD.n2335 0.00784375
R9789 VDD.n4443 VDD.n4442 0.00784375
R9790 VDD.n2383 VDD.n2377 0.00784375
R9791 VDD.n4421 VDD.n4420 0.00784375
R9792 VDD.n2425 VDD.n2419 0.00784375
R9793 VDD.n4399 VDD.n4398 0.00784375
R9794 VDD.n4329 VDD.n2744 0.00784375
R9795 VDD.n2787 VDD.n2745 0.00784375
R9796 VDD.n2800 VDD.n2785 0.00784375
R9797 VDD.n4304 VDD.n4303 0.00784375
R9798 VDD.n2869 VDD.n2867 0.00784375
R9799 VDD.n2888 VDD.n2865 0.00784375
R9800 VDD.n2890 VDD.n2861 0.00784375
R9801 VDD.n4264 VDD.n4263 0.00784375
R9802 VDD.n2938 VDD.n2936 0.00784375
R9803 VDD.n4243 VDD.n4242 0.00784375
R9804 VDD.n2985 VDD.n2979 0.00784375
R9805 VDD.n4221 VDD.n4220 0.00784375
R9806 VDD.n3029 VDD.n2989 0.00784375
R9807 VDD.n3042 VDD.n3027 0.00784375
R9808 VDD.n4193 VDD.n4192 0.00784375
R9809 VDD.n3095 VDD.n3093 0.00784375
R9810 VDD.n3111 VDD.n3091 0.00784375
R9811 VDD.n4166 VDD.n4165 0.00784375
R9812 VDD.n3161 VDD.n3159 0.00784375
R9813 VDD.n4145 VDD.n4144 0.00784375
R9814 VDD.n3204 VDD.n3202 0.00784375
R9815 VDD.n4124 VDD.n4123 0.00784375
R9816 VDD.n3251 VDD.n3245 0.00784375
R9817 VDD.n4102 VDD.n4101 0.00784375
R9818 VDD.n3295 VDD.n3255 0.00784375
R9819 VDD.n3308 VDD.n3293 0.00784375
R9820 VDD.n4074 VDD.n4073 0.00784375
R9821 VDD.n3361 VDD.n3359 0.00784375
R9822 VDD.n3377 VDD.n3357 0.00784375
R9823 VDD.n4047 VDD.n4046 0.00784375
R9824 VDD.n3427 VDD.n3425 0.00784375
R9825 VDD.n4026 VDD.n4025 0.00784375
R9826 VDD.n3470 VDD.n3468 0.00784375
R9827 VDD.n4005 VDD.n4004 0.00784375
R9828 VDD.n3517 VDD.n3511 0.00784375
R9829 VDD.n3983 VDD.n3982 0.00784375
R9830 VDD.n3561 VDD.n3521 0.00784375
R9831 VDD.n3574 VDD.n3559 0.00784375
R9832 VDD.n3955 VDD.n3954 0.00784375
R9833 VDD.n3627 VDD.n3625 0.00784375
R9834 VDD.n3643 VDD.n3623 0.00784375
R9835 VDD.n3928 VDD.n3927 0.00784375
R9836 VDD.n3693 VDD.n3691 0.00784375
R9837 VDD.n3907 VDD.n3906 0.00784375
R9838 VDD.n3736 VDD.n3734 0.00784375
R9839 VDD.n3886 VDD.n3885 0.00784375
R9840 VDD.n3783 VDD.n3777 0.00784375
R9841 VDD.n3864 VDD.n3863 0.00784375
R9842 VDD.n7092 VDD.n7091 0.0078057
R9843 VDD.n7209 VDD.n7098 0.0078057
R9844 VDD.n7129 VDD.n7099 0.0078057
R9845 VDD.n7142 VDD.n7127 0.0078057
R9846 VDD.n7183 VDD.n7182 0.0078057
R9847 VDD.n7157 VDD.n7156 0.0078057
R9848 VDD.n7152 VDD.n5 0.0078057
R9849 VDD.n7231 VDD.n5 0.0078057
R9850 VDD.n5942 VDD.n5941 0.0078057
R9851 VDD.n6059 VDD.n5948 0.0078057
R9852 VDD.n5979 VDD.n5949 0.0078057
R9853 VDD.n5992 VDD.n5977 0.0078057
R9854 VDD.n6033 VDD.n6032 0.0078057
R9855 VDD.n6007 VDD.n6006 0.0078057
R9856 VDD.n6002 VDD.n634 0.0078057
R9857 VDD.n6081 VDD.n634 0.0078057
R9858 VDD.n1270 VDD.n1229 0.00773077
R9859 VDD.n1270 VDD.n1269 0.00773077
R9860 VDD.n1282 VDD.n1261 0.00773077
R9861 VDD.n1299 VDD.n1259 0.00773077
R9862 VDD.n4907 VDD.n4906 0.00773077
R9863 VDD.n1352 VDD.n1350 0.00773077
R9864 VDD.n1368 VDD.n1348 0.00773077
R9865 VDD.n4880 VDD.n4879 0.00773077
R9866 VDD.n4393 VDD.n2428 0.00773077
R9867 VDD.n2435 VDD.n2428 0.00773077
R9868 VDD.n4384 VDD.n4383 0.00773077
R9869 VDD.n2658 VDD.n2656 0.00773077
R9870 VDD.n2674 VDD.n2654 0.00773077
R9871 VDD.n4357 VDD.n4356 0.00773077
R9872 VDD.n2722 VDD.n2721 0.00773077
R9873 VDD.n4337 VDD.n2735 0.00773077
R9874 VDD.n6184 VDD.n6181 0.00767368
R9875 VDD.n6204 VDD.n560 0.00767368
R9876 VDD.n6206 VDD.n550 0.00767368
R9877 VDD.n6230 VDD.n6229 0.00767368
R9878 VDD.n6252 VDD.n6251 0.00767368
R9879 VDD.n6272 VDD.n6271 0.00767368
R9880 VDD.n6292 VDD.n6290 0.00767368
R9881 VDD.n6317 VDD.n6316 0.00767368
R9882 VDD.n6318 VDD.n472 0.00767368
R9883 VDD.n6355 VDD.n470 0.00767368
R9884 VDD.n6376 VDD.n453 0.00767368
R9885 VDD.n6400 VDD.n440 0.00767368
R9886 VDD.n6410 VDD.n436 0.00767368
R9887 VDD.n6430 VDD.n426 0.00767368
R9888 VDD.n6432 VDD.n416 0.00767368
R9889 VDD.n6456 VDD.n6455 0.00767368
R9890 VDD.n6478 VDD.n6477 0.00767368
R9891 VDD.n6498 VDD.n6497 0.00767368
R9892 VDD.n6518 VDD.n6516 0.00767368
R9893 VDD.n6543 VDD.n6542 0.00767368
R9894 VDD.n6544 VDD.n338 0.00767368
R9895 VDD.n6581 VDD.n336 0.00767368
R9896 VDD.n6602 VDD.n319 0.00767368
R9897 VDD.n6626 VDD.n306 0.00767368
R9898 VDD.n6636 VDD.n302 0.00767368
R9899 VDD.n6656 VDD.n292 0.00767368
R9900 VDD.n6658 VDD.n282 0.00767368
R9901 VDD.n6682 VDD.n6681 0.00767368
R9902 VDD.n6704 VDD.n6703 0.00767368
R9903 VDD.n6724 VDD.n6723 0.00767368
R9904 VDD.n6744 VDD.n6742 0.00767368
R9905 VDD.n6769 VDD.n6768 0.00767368
R9906 VDD.n6770 VDD.n204 0.00767368
R9907 VDD.n6807 VDD.n202 0.00767368
R9908 VDD.n6828 VDD.n185 0.00767368
R9909 VDD.n6852 VDD.n172 0.00767368
R9910 VDD.n6862 VDD.n168 0.00767368
R9911 VDD.n6882 VDD.n158 0.00767368
R9912 VDD.n6884 VDD.n148 0.00767368
R9913 VDD.n6908 VDD.n6907 0.00767368
R9914 VDD.n6930 VDD.n6929 0.00767368
R9915 VDD.n6950 VDD.n6949 0.00767368
R9916 VDD.n6970 VDD.n6968 0.00767368
R9917 VDD.n6995 VDD.n6994 0.00767368
R9918 VDD.n6996 VDD.n70 0.00767368
R9919 VDD.n7033 VDD.n68 0.00767368
R9920 VDD.n7054 VDD.n51 0.00767368
R9921 VDD.n7059 VDD.n7058 0.00767368
R9922 VDD.n5021 VDD.n5020 0.00767368
R9923 VDD.n5032 VDD.n5031 0.00767368
R9924 VDD.n5053 VDD.n5052 0.00767368
R9925 VDD.n5056 VDD.n1171 0.00767368
R9926 VDD.n5091 VDD.n5090 0.00767368
R9927 VDD.n5115 VDD.n5113 0.00767368
R9928 VDD.n5136 VDD.n5135 0.00767368
R9929 VDD.n5137 VDD.n1110 0.00767368
R9930 VDD.n5174 VDD.n1108 0.00767368
R9931 VDD.n5195 VDD.n1090 0.00767368
R9932 VDD.n5197 VDD.n1076 0.00767368
R9933 VDD.n5230 VDD.n1074 0.00767368
R9934 VDD.n5235 VDD.n5234 0.00767368
R9935 VDD.n5260 VDD.n5259 0.00767368
R9936 VDD.n5281 VDD.n5280 0.00767368
R9937 VDD.n5284 VDD.n1036 0.00767368
R9938 VDD.n5319 VDD.n5318 0.00767368
R9939 VDD.n5343 VDD.n5341 0.00767368
R9940 VDD.n5364 VDD.n5363 0.00767368
R9941 VDD.n5365 VDD.n975 0.00767368
R9942 VDD.n5402 VDD.n973 0.00767368
R9943 VDD.n5423 VDD.n955 0.00767368
R9944 VDD.n5425 VDD.n941 0.00767368
R9945 VDD.n5458 VDD.n939 0.00767368
R9946 VDD.n5463 VDD.n5462 0.00767368
R9947 VDD.n5488 VDD.n5487 0.00767368
R9948 VDD.n5509 VDD.n5508 0.00767368
R9949 VDD.n5512 VDD.n901 0.00767368
R9950 VDD.n5547 VDD.n5546 0.00767368
R9951 VDD.n5571 VDD.n5569 0.00767368
R9952 VDD.n5592 VDD.n5591 0.00767368
R9953 VDD.n5593 VDD.n840 0.00767368
R9954 VDD.n5630 VDD.n838 0.00767368
R9955 VDD.n5651 VDD.n820 0.00767368
R9956 VDD.n5653 VDD.n806 0.00767368
R9957 VDD.n5686 VDD.n804 0.00767368
R9958 VDD.n5691 VDD.n5690 0.00767368
R9959 VDD.n5716 VDD.n5715 0.00767368
R9960 VDD.n5737 VDD.n5736 0.00767368
R9961 VDD.n5740 VDD.n766 0.00767368
R9962 VDD.n5775 VDD.n5774 0.00767368
R9963 VDD.n5798 VDD.n5797 0.00767368
R9964 VDD.n5818 VDD.n5817 0.00767368
R9965 VDD.n5840 VDD.n5838 0.00767368
R9966 VDD.n5865 VDD.n5864 0.00767368
R9967 VDD.n5866 VDD.n689 0.00767368
R9968 VDD.n5903 VDD.n687 0.00767368
R9969 VDD.n5908 VDD.n5907 0.00767368
R9970 VDD.n4877 VDD.n1374 0.00759896
R9971 VDD.n1425 VDD.n1424 0.00759896
R9972 VDD.n4856 VDD.n1431 0.00759896
R9973 VDD.n1478 VDD.n1432 0.00759896
R9974 VDD.n1494 VDD.n1493 0.00759896
R9975 VDD.n4829 VDD.n1500 0.00759896
R9976 VDD.n1542 VDD.n1501 0.00759896
R9977 VDD.n4807 VDD.n1550 0.00759896
R9978 VDD.n1584 VDD.n1551 0.00759896
R9979 VDD.n4785 VDD.n1592 0.00759896
R9980 VDD.n1626 VDD.n1593 0.00759896
R9981 VDD.n4763 VDD.n1634 0.00759896
R9982 VDD.n4758 VDD.n4757 0.00759896
R9983 VDD.n1689 VDD.n1688 0.00759896
R9984 VDD.n4735 VDD.n1695 0.00759896
R9985 VDD.n1742 VDD.n1696 0.00759896
R9986 VDD.n1758 VDD.n1757 0.00759896
R9987 VDD.n4708 VDD.n1764 0.00759896
R9988 VDD.n1806 VDD.n1765 0.00759896
R9989 VDD.n4686 VDD.n1814 0.00759896
R9990 VDD.n1848 VDD.n1815 0.00759896
R9991 VDD.n4664 VDD.n1856 0.00759896
R9992 VDD.n1890 VDD.n1857 0.00759896
R9993 VDD.n4642 VDD.n1898 0.00759896
R9994 VDD.n4637 VDD.n4636 0.00759896
R9995 VDD.n1953 VDD.n1952 0.00759896
R9996 VDD.n4614 VDD.n1959 0.00759896
R9997 VDD.n2006 VDD.n1960 0.00759896
R9998 VDD.n2022 VDD.n2021 0.00759896
R9999 VDD.n4587 VDD.n2028 0.00759896
R10000 VDD.n2070 VDD.n2029 0.00759896
R10001 VDD.n4565 VDD.n2078 0.00759896
R10002 VDD.n2112 VDD.n2079 0.00759896
R10003 VDD.n4543 VDD.n2120 0.00759896
R10004 VDD.n2154 VDD.n2121 0.00759896
R10005 VDD.n4521 VDD.n2162 0.00759896
R10006 VDD.n4516 VDD.n4515 0.00759896
R10007 VDD.n2217 VDD.n2216 0.00759896
R10008 VDD.n4493 VDD.n2223 0.00759896
R10009 VDD.n2270 VDD.n2224 0.00759896
R10010 VDD.n2286 VDD.n2285 0.00759896
R10011 VDD.n4466 VDD.n2292 0.00759896
R10012 VDD.n2334 VDD.n2293 0.00759896
R10013 VDD.n4444 VDD.n2342 0.00759896
R10014 VDD.n2376 VDD.n2343 0.00759896
R10015 VDD.n4422 VDD.n2384 0.00759896
R10016 VDD.n2418 VDD.n2385 0.00759896
R10017 VDD.n4400 VDD.n2426 0.00759896
R10018 VDD.n4336 VDD.n2736 0.00759896
R10019 VDD.n4328 VDD.n4327 0.00759896
R10020 VDD.n2799 VDD.n2798 0.00759896
R10021 VDD.n4305 VDD.n2805 0.00759896
R10022 VDD.n2868 VDD.n2806 0.00759896
R10023 VDD.n2875 VDD.n2874 0.00759896
R10024 VDD.n2891 VDD.n2889 0.00759896
R10025 VDD.n2903 VDD.n2902 0.00759896
R10026 VDD.n2937 VDD.n2904 0.00759896
R10027 VDD.n2946 VDD.n2945 0.00759896
R10028 VDD.n2978 VDD.n2947 0.00759896
R10029 VDD.n4222 VDD.n2986 0.00759896
R10030 VDD.n4217 VDD.n4216 0.00759896
R10031 VDD.n3041 VDD.n3040 0.00759896
R10032 VDD.n4194 VDD.n3047 0.00759896
R10033 VDD.n3094 VDD.n3048 0.00759896
R10034 VDD.n3110 VDD.n3109 0.00759896
R10035 VDD.n4167 VDD.n3116 0.00759896
R10036 VDD.n3160 VDD.n3117 0.00759896
R10037 VDD.n3169 VDD.n3168 0.00759896
R10038 VDD.n3203 VDD.n3170 0.00759896
R10039 VDD.n3212 VDD.n3211 0.00759896
R10040 VDD.n3244 VDD.n3213 0.00759896
R10041 VDD.n4103 VDD.n3252 0.00759896
R10042 VDD.n4098 VDD.n4097 0.00759896
R10043 VDD.n3307 VDD.n3306 0.00759896
R10044 VDD.n4075 VDD.n3313 0.00759896
R10045 VDD.n3360 VDD.n3314 0.00759896
R10046 VDD.n3376 VDD.n3375 0.00759896
R10047 VDD.n4048 VDD.n3382 0.00759896
R10048 VDD.n3426 VDD.n3383 0.00759896
R10049 VDD.n3435 VDD.n3434 0.00759896
R10050 VDD.n3469 VDD.n3436 0.00759896
R10051 VDD.n3478 VDD.n3477 0.00759896
R10052 VDD.n3510 VDD.n3479 0.00759896
R10053 VDD.n3984 VDD.n3518 0.00759896
R10054 VDD.n3979 VDD.n3978 0.00759896
R10055 VDD.n3573 VDD.n3572 0.00759896
R10056 VDD.n3956 VDD.n3579 0.00759896
R10057 VDD.n3626 VDD.n3580 0.00759896
R10058 VDD.n3642 VDD.n3641 0.00759896
R10059 VDD.n3929 VDD.n3648 0.00759896
R10060 VDD.n3692 VDD.n3649 0.00759896
R10061 VDD.n3701 VDD.n3700 0.00759896
R10062 VDD.n3735 VDD.n3702 0.00759896
R10063 VDD.n3744 VDD.n3743 0.00759896
R10064 VDD.n3776 VDD.n3745 0.00759896
R10065 VDD.n3865 VDD.n3784 0.00759896
R10066 VDD.n7079 VDD.n37 0.00756218
R10067 VDD.n7097 VDD.n35 0.00756218
R10068 VDD.n7133 VDD.n7132 0.00756218
R10069 VDD.n7184 VDD.n7143 0.00756218
R10070 VDD.n5929 VDD.n666 0.00756218
R10071 VDD.n5947 VDD.n664 0.00756218
R10072 VDD.n5983 VDD.n5982 0.00756218
R10073 VDD.n6034 VDD.n5993 0.00756218
R10074 VDD.n7208 VDD.n7207 0.00756218
R10075 VDD.n7151 VDD.n7144 0.00756218
R10076 VDD.n6058 VDD.n6057 0.00756218
R10077 VDD.n6001 VDD.n5994 0.00756218
R10078 VDD.n1281 VDD.n1280 0.00748974
R10079 VDD.n1298 VDD.n1297 0.00748974
R10080 VDD.n4908 VDD.n1304 0.00748974
R10081 VDD.n1351 VDD.n1305 0.00748974
R10082 VDD.n1367 VDD.n1366 0.00748974
R10083 VDD.n4881 VDD.n1373 0.00748974
R10084 VDD.n4385 VDD.n2436 0.00748974
R10085 VDD.n2657 VDD.n2437 0.00748974
R10086 VDD.n2673 VDD.n2672 0.00748974
R10087 VDD.n4358 VDD.n2679 0.00748974
R10088 VDD.n2719 VDD.n2680 0.00748974
R10089 VDD.n2734 VDD.n2717 0.00748974
R10090 VDD.n6091 VDD.n6089 0.00701042
R10091 VDD.n6120 VDD.n608 0.00701042
R10092 VDD.n2478 VDD.n2477 0.00701042
R10093 VDD.n4960 VDD.n4935 0.00701042
R10094 VDD.n7279 VDD.n7278 0.00701042
R10095 VDD.n7277 VDD.n7265 0.00701042
R10096 VDD.n6084 VDD.n6083 0.0066978
R10097 VDD.n3847 VDD.n3802 0.00635126
R10098 VDD.n3850 VDD.n3798 0.00635126
R10099 VDD.n3853 VDD.n3794 0.00635126
R10100 VDD.n3856 VDD.n3790 0.00635126
R10101 VDD.n3859 VDD.n3786 0.00635126
R10102 VDD.n2582 VDD.n2577 0.00635126
R10103 VDD.n2585 VDD.n2571 0.00635126
R10104 VDD.n2589 VDD.n2569 0.00635126
R10105 VDD.n2545 VDD.n2532 0.00635126
R10106 VDD.n2523 VDD.n2499 0.00635126
R10107 VDD.n2526 VDD.n2493 0.00635126
R10108 VDD.n2556 VDD.n2491 0.00635126
R10109 VDD.n2553 VDD.n2530 0.00635126
R10110 VDD.n2482 VDD.n2475 0.00570833
R10111 VDD.n2482 VDD.n2481 0.00570833
R10112 VDD.n4964 VDD.n4934 0.00570833
R10113 VDD.n4964 VDD.n4963 0.00570833
R10114 VDD.n6186 VDD.n560 0.00544737
R10115 VDD.n6207 VDD.n6206 0.00544737
R10116 VDD.n6229 VDD.n6228 0.00544737
R10117 VDD.n6251 VDD.n6250 0.00544737
R10118 VDD.n6271 VDD.n6270 0.00544737
R10119 VDD.n6316 VDD.n486 0.00544737
R10120 VDD.n6322 VDD.n6318 0.00544737
R10121 VDD.n6350 VDD.n470 0.00544737
R10122 VDD.n6357 VDD.n453 0.00544737
R10123 VDD.n6378 VDD.n440 0.00544737
R10124 VDD.n6412 VDD.n426 0.00544737
R10125 VDD.n6433 VDD.n6432 0.00544737
R10126 VDD.n6455 VDD.n6454 0.00544737
R10127 VDD.n6477 VDD.n6476 0.00544737
R10128 VDD.n6497 VDD.n6496 0.00544737
R10129 VDD.n6542 VDD.n352 0.00544737
R10130 VDD.n6548 VDD.n6544 0.00544737
R10131 VDD.n6576 VDD.n336 0.00544737
R10132 VDD.n6583 VDD.n319 0.00544737
R10133 VDD.n6604 VDD.n306 0.00544737
R10134 VDD.n6638 VDD.n292 0.00544737
R10135 VDD.n6659 VDD.n6658 0.00544737
R10136 VDD.n6681 VDD.n6680 0.00544737
R10137 VDD.n6703 VDD.n6702 0.00544737
R10138 VDD.n6723 VDD.n6722 0.00544737
R10139 VDD.n6768 VDD.n218 0.00544737
R10140 VDD.n6774 VDD.n6770 0.00544737
R10141 VDD.n6802 VDD.n202 0.00544737
R10142 VDD.n6809 VDD.n185 0.00544737
R10143 VDD.n6830 VDD.n172 0.00544737
R10144 VDD.n6864 VDD.n158 0.00544737
R10145 VDD.n6885 VDD.n6884 0.00544737
R10146 VDD.n6907 VDD.n6906 0.00544737
R10147 VDD.n6929 VDD.n6928 0.00544737
R10148 VDD.n6949 VDD.n6948 0.00544737
R10149 VDD.n6994 VDD.n84 0.00544737
R10150 VDD.n7000 VDD.n6996 0.00544737
R10151 VDD.n7028 VDD.n68 0.00544737
R10152 VDD.n7035 VDD.n51 0.00544737
R10153 VDD.n7060 VDD.n7059 0.00544737
R10154 VDD.n5031 VDD.n5030 0.00544737
R10155 VDD.n5052 VDD.n5051 0.00544737
R10156 VDD.n5057 VDD.n5056 0.00544737
R10157 VDD.n5090 VDD.n5089 0.00544737
R10158 VDD.n5113 VDD.n5112 0.00544737
R10159 VDD.n5141 VDD.n5137 0.00544737
R10160 VDD.n5169 VDD.n1108 0.00544737
R10161 VDD.n5176 VDD.n1090 0.00544737
R10162 VDD.n5198 VDD.n5197 0.00544737
R10163 VDD.n5225 VDD.n1074 0.00544737
R10164 VDD.n5259 VDD.n5258 0.00544737
R10165 VDD.n5280 VDD.n5279 0.00544737
R10166 VDD.n5285 VDD.n5284 0.00544737
R10167 VDD.n5318 VDD.n5317 0.00544737
R10168 VDD.n5341 VDD.n5340 0.00544737
R10169 VDD.n5369 VDD.n5365 0.00544737
R10170 VDD.n5397 VDD.n973 0.00544737
R10171 VDD.n5404 VDD.n955 0.00544737
R10172 VDD.n5426 VDD.n5425 0.00544737
R10173 VDD.n5453 VDD.n939 0.00544737
R10174 VDD.n5487 VDD.n5486 0.00544737
R10175 VDD.n5508 VDD.n5507 0.00544737
R10176 VDD.n5513 VDD.n5512 0.00544737
R10177 VDD.n5546 VDD.n5545 0.00544737
R10178 VDD.n5569 VDD.n5568 0.00544737
R10179 VDD.n5597 VDD.n5593 0.00544737
R10180 VDD.n5625 VDD.n838 0.00544737
R10181 VDD.n5632 VDD.n820 0.00544737
R10182 VDD.n5654 VDD.n5653 0.00544737
R10183 VDD.n5681 VDD.n804 0.00544737
R10184 VDD.n5715 VDD.n5714 0.00544737
R10185 VDD.n5736 VDD.n5735 0.00544737
R10186 VDD.n5741 VDD.n5740 0.00544737
R10187 VDD.n5774 VDD.n5773 0.00544737
R10188 VDD.n5797 VDD.n5796 0.00544737
R10189 VDD.n5838 VDD.n5837 0.00544737
R10190 VDD.n5864 VDD.n703 0.00544737
R10191 VDD.n5870 VDD.n5866 0.00544737
R10192 VDD.n5898 VDD.n687 0.00544737
R10193 VDD.n5909 VDD.n5908 0.00544737
R10194 VDD.n1424 VDD.n1409 0.00539583
R10195 VDD.n1431 VDD.n1407 0.00539583
R10196 VDD.n4854 VDD.n1432 0.00539583
R10197 VDD.n1493 VDD.n1477 0.00539583
R10198 VDD.n1500 VDD.n1475 0.00539583
R10199 VDD.n1550 VDD.n1549 0.00539583
R10200 VDD.n4805 VDD.n1551 0.00539583
R10201 VDD.n1592 VDD.n1591 0.00539583
R10202 VDD.n4783 VDD.n1593 0.00539583
R10203 VDD.n1634 VDD.n1633 0.00539583
R10204 VDD.n1688 VDD.n1677 0.00539583
R10205 VDD.n1695 VDD.n1675 0.00539583
R10206 VDD.n4733 VDD.n1696 0.00539583
R10207 VDD.n1757 VDD.n1741 0.00539583
R10208 VDD.n1764 VDD.n1739 0.00539583
R10209 VDD.n1814 VDD.n1813 0.00539583
R10210 VDD.n4684 VDD.n1815 0.00539583
R10211 VDD.n1856 VDD.n1855 0.00539583
R10212 VDD.n4662 VDD.n1857 0.00539583
R10213 VDD.n1898 VDD.n1897 0.00539583
R10214 VDD.n1952 VDD.n1941 0.00539583
R10215 VDD.n1959 VDD.n1939 0.00539583
R10216 VDD.n4612 VDD.n1960 0.00539583
R10217 VDD.n2021 VDD.n2005 0.00539583
R10218 VDD.n2028 VDD.n2003 0.00539583
R10219 VDD.n2078 VDD.n2077 0.00539583
R10220 VDD.n4563 VDD.n2079 0.00539583
R10221 VDD.n2120 VDD.n2119 0.00539583
R10222 VDD.n4541 VDD.n2121 0.00539583
R10223 VDD.n2162 VDD.n2161 0.00539583
R10224 VDD.n2216 VDD.n2205 0.00539583
R10225 VDD.n2223 VDD.n2203 0.00539583
R10226 VDD.n4491 VDD.n2224 0.00539583
R10227 VDD.n2285 VDD.n2269 0.00539583
R10228 VDD.n2292 VDD.n2267 0.00539583
R10229 VDD.n2342 VDD.n2341 0.00539583
R10230 VDD.n4442 VDD.n2343 0.00539583
R10231 VDD.n2384 VDD.n2383 0.00539583
R10232 VDD.n4420 VDD.n2385 0.00539583
R10233 VDD.n2426 VDD.n2425 0.00539583
R10234 VDD.n4329 VDD.n4328 0.00539583
R10235 VDD.n2798 VDD.n2787 0.00539583
R10236 VDD.n2805 VDD.n2785 0.00539583
R10237 VDD.n4303 VDD.n2806 0.00539583
R10238 VDD.n2874 VDD.n2867 0.00539583
R10239 VDD.n2902 VDD.n2861 0.00539583
R10240 VDD.n4263 VDD.n2904 0.00539583
R10241 VDD.n2945 VDD.n2936 0.00539583
R10242 VDD.n4242 VDD.n2947 0.00539583
R10243 VDD.n2986 VDD.n2985 0.00539583
R10244 VDD.n3040 VDD.n3029 0.00539583
R10245 VDD.n3047 VDD.n3027 0.00539583
R10246 VDD.n4192 VDD.n3048 0.00539583
R10247 VDD.n3109 VDD.n3093 0.00539583
R10248 VDD.n3116 VDD.n3091 0.00539583
R10249 VDD.n3168 VDD.n3159 0.00539583
R10250 VDD.n4144 VDD.n3170 0.00539583
R10251 VDD.n3211 VDD.n3202 0.00539583
R10252 VDD.n4123 VDD.n3213 0.00539583
R10253 VDD.n3252 VDD.n3251 0.00539583
R10254 VDD.n3306 VDD.n3295 0.00539583
R10255 VDD.n3313 VDD.n3293 0.00539583
R10256 VDD.n4073 VDD.n3314 0.00539583
R10257 VDD.n3375 VDD.n3359 0.00539583
R10258 VDD.n3382 VDD.n3357 0.00539583
R10259 VDD.n3434 VDD.n3425 0.00539583
R10260 VDD.n4025 VDD.n3436 0.00539583
R10261 VDD.n3477 VDD.n3468 0.00539583
R10262 VDD.n4004 VDD.n3479 0.00539583
R10263 VDD.n3518 VDD.n3517 0.00539583
R10264 VDD.n3572 VDD.n3561 0.00539583
R10265 VDD.n3579 VDD.n3559 0.00539583
R10266 VDD.n3954 VDD.n3580 0.00539583
R10267 VDD.n3641 VDD.n3625 0.00539583
R10268 VDD.n3648 VDD.n3623 0.00539583
R10269 VDD.n3700 VDD.n3691 0.00539583
R10270 VDD.n3906 VDD.n3702 0.00539583
R10271 VDD.n3743 VDD.n3734 0.00539583
R10272 VDD.n3885 VDD.n3745 0.00539583
R10273 VDD.n3784 VDD.n3783 0.00539583
R10274 VDD.n7092 VDD.n35 0.00537047
R10275 VDD.n7209 VDD.n7208 0.00537047
R10276 VDD.n7132 VDD.n7129 0.00537047
R10277 VDD.n7143 VDD.n7142 0.00537047
R10278 VDD.n7182 VDD.n7144 0.00537047
R10279 VDD.n5942 VDD.n664 0.00537047
R10280 VDD.n6059 VDD.n6058 0.00537047
R10281 VDD.n5982 VDD.n5979 0.00537047
R10282 VDD.n5993 VDD.n5992 0.00537047
R10283 VDD.n6032 VDD.n5994 0.00537047
R10284 VDD.n1297 VDD.n1261 0.00532051
R10285 VDD.n1304 VDD.n1259 0.00532051
R10286 VDD.n4906 VDD.n1305 0.00532051
R10287 VDD.n1366 VDD.n1350 0.00532051
R10288 VDD.n1373 VDD.n1348 0.00532051
R10289 VDD.n4383 VDD.n2437 0.00532051
R10290 VDD.n2672 VDD.n2656 0.00532051
R10291 VDD.n2679 VDD.n2654 0.00532051
R10292 VDD.n4356 VDD.n2680 0.00532051
R10293 VDD.n2722 VDD.n2717 0.00532051
R10294 VDD.n3842 VDD.n3833 0.00518613
R10295 VDD.n2518 VDD.n2509 0.00518613
R10296 VDD.n6139 VDD.n6138 0.00511607
R10297 VDD.n4982 VDD.n4981 0.00511607
R10298 VDD.n3843 VDD.n3829 0.00493396
R10299 VDD.n3845 VDD.n3829 0.00493396
R10300 VDD.n3846 VDD.n3801 0.00493396
R10301 VDD.n3848 VDD.n3801 0.00493396
R10302 VDD.n3849 VDD.n3797 0.00493396
R10303 VDD.n3851 VDD.n3797 0.00493396
R10304 VDD.n3852 VDD.n3793 0.00493396
R10305 VDD.n3854 VDD.n3793 0.00493396
R10306 VDD.n3855 VDD.n3789 0.00493396
R10307 VDD.n3857 VDD.n3789 0.00493396
R10308 VDD.n3858 VDD.n3785 0.00493396
R10309 VDD.n3860 VDD.n3785 0.00493396
R10310 VDD.n2519 VDD.n2505 0.00493396
R10311 VDD.n2521 VDD.n2505 0.00493396
R10312 VDD.n2522 VDD.n2498 0.00493396
R10313 VDD.n2524 VDD.n2498 0.00493396
R10314 VDD.n2525 VDD.n2492 0.00493396
R10315 VDD.n2527 VDD.n2492 0.00493396
R10316 VDD.n2557 VDD.n2528 0.00493396
R10317 VDD.n2557 VDD.n2555 0.00493396
R10318 VDD.n2554 VDD.n2529 0.00493396
R10319 VDD.n2547 VDD.n2529 0.00493396
R10320 VDD.n2546 VDD.n2531 0.00493396
R10321 VDD.n2531 VDD.n2427 0.00493396
R10322 VDD.n6085 VDD.n632 0.00490305
R10323 VDD.n7239 VDD.n7238 0.00490305
R10324 VDD.n7230 VDD.n6 0.00480499
R10325 VDD.n6120 VDD.n6119 0.00440625
R10326 VDD.n7265 VDD.n7264 0.00440625
R10327 VDD.n4998 VDD.t21 0.00429204
R10328 VDD.n6155 VDD.t0 0.00429204
R10329 VDD.n5939 VDD.n5931 0.00428788
R10330 VDD.n660 VDD.n658 0.00428788
R10331 VDD.n6054 VDD.n5952 0.00428788
R10332 VDD.n5986 VDD.n5956 0.00428788
R10333 VDD.n6037 VDD.n5974 0.00428788
R10334 VDD.n6028 VDD.n6009 0.00428788
R10335 VDD.n6189 VDD.n566 0.00428788
R10336 VDD.n6210 VDD.n557 0.00428788
R10337 VDD.n6223 VDD.n543 0.00428788
R10338 VDD.n6247 VDD.n536 0.00428788
R10339 VDD.n6267 VDD.n525 0.00428788
R10340 VDD.n6286 VDD.n503 0.00428788
R10341 VDD.n6295 VDD.n499 0.00428788
R10342 VDD.n6325 VDD.n483 0.00428788
R10343 VDD.n6347 VDD.n474 0.00428788
R10344 VDD.n467 VDD.n463 0.00428788
R10345 VDD.n6373 VDD.n456 0.00428788
R10346 VDD.n6397 VDD.n443 0.00428788
R10347 VDD.n6415 VDD.n434 0.00428788
R10348 VDD.n6436 VDD.n423 0.00428788
R10349 VDD.n6449 VDD.n409 0.00428788
R10350 VDD.n6473 VDD.n402 0.00428788
R10351 VDD.n6493 VDD.n391 0.00428788
R10352 VDD.n6512 VDD.n369 0.00428788
R10353 VDD.n6521 VDD.n365 0.00428788
R10354 VDD.n6551 VDD.n349 0.00428788
R10355 VDD.n6573 VDD.n340 0.00428788
R10356 VDD.n333 VDD.n329 0.00428788
R10357 VDD.n6599 VDD.n322 0.00428788
R10358 VDD.n6623 VDD.n309 0.00428788
R10359 VDD.n6641 VDD.n300 0.00428788
R10360 VDD.n6662 VDD.n289 0.00428788
R10361 VDD.n6675 VDD.n275 0.00428788
R10362 VDD.n6699 VDD.n268 0.00428788
R10363 VDD.n6719 VDD.n257 0.00428788
R10364 VDD.n6738 VDD.n235 0.00428788
R10365 VDD.n6747 VDD.n231 0.00428788
R10366 VDD.n6777 VDD.n215 0.00428788
R10367 VDD.n6799 VDD.n206 0.00428788
R10368 VDD.n199 VDD.n195 0.00428788
R10369 VDD.n6825 VDD.n188 0.00428788
R10370 VDD.n6849 VDD.n175 0.00428788
R10371 VDD.n6867 VDD.n166 0.00428788
R10372 VDD.n6888 VDD.n155 0.00428788
R10373 VDD.n6901 VDD.n141 0.00428788
R10374 VDD.n6925 VDD.n134 0.00428788
R10375 VDD.n6945 VDD.n123 0.00428788
R10376 VDD.n6964 VDD.n101 0.00428788
R10377 VDD.n6973 VDD.n97 0.00428788
R10378 VDD.n7003 VDD.n81 0.00428788
R10379 VDD.n7025 VDD.n72 0.00428788
R10380 VDD.n65 VDD.n61 0.00428788
R10381 VDD.n7051 VDD.n54 0.00428788
R10382 VDD.n43 VDD.n41 0.00428788
R10383 VDD.n7089 VDD.n7081 0.00428788
R10384 VDD.n31 VDD.n29 0.00428788
R10385 VDD.n7204 VDD.n7102 0.00428788
R10386 VDD.n7136 VDD.n7106 0.00428788
R10387 VDD.n7187 VDD.n7124 0.00428788
R10388 VDD.n7178 VDD.n7159 0.00428788
R10389 VDD.n2633 VDD.n2434 0.00428788
R10390 VDD.n2443 VDD.n2441 0.00428788
R10391 VDD.n2667 VDD.n2647 0.00428788
R10392 VDD.n4360 VDD.n2651 0.00428788
R10393 VDD.n2686 VDD.n2684 0.00428788
R10394 VDD.n4339 VDD.n2715 0.00428788
R10395 VDD.n1377 VDD.n1376 0.00428788
R10396 VDD.n1419 VDD.n1400 0.00428788
R10397 VDD.n4858 VDD.n1404 0.00428788
R10398 VDD.n1438 VDD.n1436 0.00428788
R10399 VDD.n1488 VDD.n1468 0.00428788
R10400 VDD.n4831 VDD.n1472 0.00428788
R10401 VDD.n4823 VDD.n1505 0.00428788
R10402 VDD.n4810 VDD.n1539 0.00428788
R10403 VDD.n4801 VDD.n1555 0.00428788
R10404 VDD.n4788 VDD.n1581 0.00428788
R10405 VDD.n4779 VDD.n1597 0.00428788
R10406 VDD.n4766 VDD.n1623 0.00428788
R10407 VDD.n4755 VDD.n4754 0.00428788
R10408 VDD.n1683 VDD.n1668 0.00428788
R10409 VDD.n4737 VDD.n1672 0.00428788
R10410 VDD.n1702 VDD.n1700 0.00428788
R10411 VDD.n1752 VDD.n1732 0.00428788
R10412 VDD.n4710 VDD.n1736 0.00428788
R10413 VDD.n4702 VDD.n1769 0.00428788
R10414 VDD.n4689 VDD.n1803 0.00428788
R10415 VDD.n4680 VDD.n1819 0.00428788
R10416 VDD.n4667 VDD.n1845 0.00428788
R10417 VDD.n4658 VDD.n1861 0.00428788
R10418 VDD.n4645 VDD.n1887 0.00428788
R10419 VDD.n4634 VDD.n4633 0.00428788
R10420 VDD.n1947 VDD.n1932 0.00428788
R10421 VDD.n4616 VDD.n1936 0.00428788
R10422 VDD.n1966 VDD.n1964 0.00428788
R10423 VDD.n2016 VDD.n1996 0.00428788
R10424 VDD.n4589 VDD.n2000 0.00428788
R10425 VDD.n4581 VDD.n2033 0.00428788
R10426 VDD.n4568 VDD.n2067 0.00428788
R10427 VDD.n4559 VDD.n2083 0.00428788
R10428 VDD.n4546 VDD.n2109 0.00428788
R10429 VDD.n4537 VDD.n2125 0.00428788
R10430 VDD.n4524 VDD.n2151 0.00428788
R10431 VDD.n4513 VDD.n4512 0.00428788
R10432 VDD.n2211 VDD.n2196 0.00428788
R10433 VDD.n4495 VDD.n2200 0.00428788
R10434 VDD.n2230 VDD.n2228 0.00428788
R10435 VDD.n2280 VDD.n2260 0.00428788
R10436 VDD.n4468 VDD.n2264 0.00428788
R10437 VDD.n4460 VDD.n2297 0.00428788
R10438 VDD.n4447 VDD.n2331 0.00428788
R10439 VDD.n4438 VDD.n2347 0.00428788
R10440 VDD.n4425 VDD.n2373 0.00428788
R10441 VDD.n4416 VDD.n2389 0.00428788
R10442 VDD.n4403 VDD.n2415 0.00428788
R10443 VDD.n1285 VDD.n1263 0.00428788
R10444 VDD.n1292 VDD.n1252 0.00428788
R10445 VDD.n4910 VDD.n1256 0.00428788
R10446 VDD.n1311 VDD.n1309 0.00428788
R10447 VDD.n1361 VDD.n1341 0.00428788
R10448 VDD.n4883 VDD.n1345 0.00428788
R10449 VDD.n4332 VDD.n2738 0.00428788
R10450 VDD.n4325 VDD.n4324 0.00428788
R10451 VDD.n2793 VDD.n2778 0.00428788
R10452 VDD.n4307 VDD.n2782 0.00428788
R10453 VDD.n2812 VDD.n2810 0.00428788
R10454 VDD.n2883 VDD.n2842 0.00428788
R10455 VDD.n2895 VDD.n2894 0.00428788
R10456 VDD.n4267 VDD.n4266 0.00428788
R10457 VDD.n4259 VDD.n2907 0.00428788
R10458 VDD.n4246 VDD.n4245 0.00428788
R10459 VDD.n4238 VDD.n2950 0.00428788
R10460 VDD.n4225 VDD.n2975 0.00428788
R10461 VDD.n4214 VDD.n4213 0.00428788
R10462 VDD.n3035 VDD.n3020 0.00428788
R10463 VDD.n4196 VDD.n3024 0.00428788
R10464 VDD.n3054 VDD.n3052 0.00428788
R10465 VDD.n3104 VDD.n3084 0.00428788
R10466 VDD.n4169 VDD.n3088 0.00428788
R10467 VDD.n4161 VDD.n3121 0.00428788
R10468 VDD.n4148 VDD.n4147 0.00428788
R10469 VDD.n4140 VDD.n3173 0.00428788
R10470 VDD.n4127 VDD.n4126 0.00428788
R10471 VDD.n4119 VDD.n3216 0.00428788
R10472 VDD.n4106 VDD.n3241 0.00428788
R10473 VDD.n4095 VDD.n4094 0.00428788
R10474 VDD.n3301 VDD.n3286 0.00428788
R10475 VDD.n4077 VDD.n3290 0.00428788
R10476 VDD.n3320 VDD.n3318 0.00428788
R10477 VDD.n3370 VDD.n3350 0.00428788
R10478 VDD.n4050 VDD.n3354 0.00428788
R10479 VDD.n4042 VDD.n3387 0.00428788
R10480 VDD.n4029 VDD.n4028 0.00428788
R10481 VDD.n4021 VDD.n3439 0.00428788
R10482 VDD.n4008 VDD.n4007 0.00428788
R10483 VDD.n4000 VDD.n3482 0.00428788
R10484 VDD.n3987 VDD.n3507 0.00428788
R10485 VDD.n3976 VDD.n3975 0.00428788
R10486 VDD.n3567 VDD.n3552 0.00428788
R10487 VDD.n3958 VDD.n3556 0.00428788
R10488 VDD.n3586 VDD.n3584 0.00428788
R10489 VDD.n3636 VDD.n3616 0.00428788
R10490 VDD.n3931 VDD.n3620 0.00428788
R10491 VDD.n3923 VDD.n3653 0.00428788
R10492 VDD.n3910 VDD.n3909 0.00428788
R10493 VDD.n3902 VDD.n3705 0.00428788
R10494 VDD.n3889 VDD.n3888 0.00428788
R10495 VDD.n3881 VDD.n3748 0.00428788
R10496 VDD.n3868 VDD.n3773 0.00428788
R10497 VDD.n5027 VDD.n1197 0.00428788
R10498 VDD.n5048 VDD.n1186 0.00428788
R10499 VDD.n5062 VDD.n5061 0.00428788
R10500 VDD.n5084 VDD.n1164 0.00428788
R10501 VDD.n5109 VDD.n1157 0.00428788
R10502 VDD.n5130 VDD.n1126 0.00428788
R10503 VDD.n5144 VDD.n1121 0.00428788
R10504 VDD.n5166 VDD.n1112 0.00428788
R10505 VDD.n1105 VDD.n1101 0.00428788
R10506 VDD.n5192 VDD.n1093 0.00428788
R10507 VDD.n5222 VDD.n1078 0.00428788
R10508 VDD.n1069 VDD.n1068 0.00428788
R10509 VDD.n5255 VDD.n1062 0.00428788
R10510 VDD.n5276 VDD.n1051 0.00428788
R10511 VDD.n5290 VDD.n5289 0.00428788
R10512 VDD.n5312 VDD.n1029 0.00428788
R10513 VDD.n5337 VDD.n1022 0.00428788
R10514 VDD.n5358 VDD.n991 0.00428788
R10515 VDD.n5372 VDD.n986 0.00428788
R10516 VDD.n5394 VDD.n977 0.00428788
R10517 VDD.n970 VDD.n966 0.00428788
R10518 VDD.n5420 VDD.n958 0.00428788
R10519 VDD.n5450 VDD.n943 0.00428788
R10520 VDD.n934 VDD.n933 0.00428788
R10521 VDD.n5483 VDD.n927 0.00428788
R10522 VDD.n5504 VDD.n916 0.00428788
R10523 VDD.n5518 VDD.n5517 0.00428788
R10524 VDD.n5540 VDD.n894 0.00428788
R10525 VDD.n5565 VDD.n887 0.00428788
R10526 VDD.n5586 VDD.n856 0.00428788
R10527 VDD.n5600 VDD.n851 0.00428788
R10528 VDD.n5622 VDD.n842 0.00428788
R10529 VDD.n835 VDD.n831 0.00428788
R10530 VDD.n5648 VDD.n823 0.00428788
R10531 VDD.n5678 VDD.n808 0.00428788
R10532 VDD.n799 VDD.n798 0.00428788
R10533 VDD.n5711 VDD.n792 0.00428788
R10534 VDD.n5732 VDD.n781 0.00428788
R10535 VDD.n5746 VDD.n5745 0.00428788
R10536 VDD.n5768 VDD.n759 0.00428788
R10537 VDD.n5793 VDD.n752 0.00428788
R10538 VDD.n5813 VDD.n730 0.00428788
R10539 VDD.n5822 VDD.n5821 0.00428788
R10540 VDD.n5844 VDD.n5843 0.00428788
R10541 VDD.n5873 VDD.n700 0.00428788
R10542 VDD.n5895 VDD.n691 0.00428788
R10543 VDD.n682 VDD.n678 0.00428788
R10544 VDD.n672 VDD.n670 0.00428788
R10545 VDD.n6135 VDD.n6134 0.00428087
R10546 VDD.n2606 VDD.n2466 0.00428087
R10547 VDD.n2615 VDD.n2459 0.00428087
R10548 VDD.n4977 VDD.n1232 0.00428087
R10549 VDD.n4951 VDD.n1231 0.00428087
R10550 VDD.n7248 VDD.n7247 0.00428087
R10551 VDD.n6176 VDD.n569 0.00397409
R10552 VDD.n5015 VDD.n1199 0.00397409
R10553 VDD.n6080 VDD.n635 0.00391036
R10554 VDD.n4392 VDD.n4391 0.00391036
R10555 VDD.n1272 VDD.n1271 0.00391036
R10556 VDD.n2576 VDD.n2465 0.00387321
R10557 VDD.n2583 VDD.n2576 0.00387321
R10558 VDD.n2584 VDD.n2570 0.00387321
R10559 VDD.n2586 VDD.n2570 0.00387321
R10560 VDD.n2590 VDD.n2587 0.00387321
R10561 VDD.n2590 VDD.n2588 0.00387321
R10562 VDD.n6084 VDD.n620 0.00379258
R10563 VDD VDD.n7233 0.00364833
R10564 VDD.n6086 VDD.n6085 0.00360776
R10565 VDD.n6135 VDD.n600 0.00360776
R10566 VDD.n2606 VDD.n2605 0.00360776
R10567 VDD.n2459 VDD.n2458 0.00360776
R10568 VDD.n4977 VDD.n4976 0.00360776
R10569 VDD.n4938 VDD.n1231 0.00360776
R10570 VDD.n7240 VDD.n7239 0.00360776
R10571 VDD.n7258 VDD.n7248 0.00360776
R10572 VDD VDD.n6136 0.00353434
R10573 VDD.n597 VDD.n590 0.00351641
R10574 VDD.n1227 VDD.n1220 0.00351641
R10575 VDD.n5140 VDD.n1123 0.00326471
R10576 VDD.n5170 VDD.n1109 0.00326471
R10577 VDD.n5178 VDD.n5177 0.00326471
R10578 VDD.n5200 VDD.n5199 0.00326471
R10579 VDD.n5226 VDD.n1075 0.00326471
R10580 VDD.n5238 VDD.n5237 0.00326471
R10581 VDD.n5368 VDD.n988 0.00326471
R10582 VDD.n5398 VDD.n974 0.00326471
R10583 VDD.n5406 VDD.n5405 0.00326471
R10584 VDD.n5428 VDD.n5427 0.00326471
R10585 VDD.n5454 VDD.n940 0.00326471
R10586 VDD.n5466 VDD.n5465 0.00326471
R10587 VDD.n5596 VDD.n853 0.00326471
R10588 VDD.n5626 VDD.n839 0.00326471
R10589 VDD.n5634 VDD.n5633 0.00326471
R10590 VDD.n5656 VDD.n5655 0.00326471
R10591 VDD.n5682 VDD.n805 0.00326471
R10592 VDD.n5694 VDD.n5693 0.00326471
R10593 VDD.n5836 VDD.n5835 0.00326471
R10594 VDD.n5861 VDD.n5860 0.00326471
R10595 VDD.n5869 VDD.n702 0.00326471
R10596 VDD.n5899 VDD.n688 0.00326471
R10597 VDD.n5911 VDD.n5910 0.00326471
R10598 VDD.n5943 VDD.n665 0.00326471
R10599 VDD.n6061 VDD.n6060 0.00326471
R10600 VDD.n5980 VDD.n5951 0.00326471
R10601 VDD.n5991 VDD.n5990 0.00326471
R10602 VDD.n6031 VDD.n5995 0.00326471
R10603 VDD.n6005 VDD.n6000 0.00326471
R10604 VDD.n6313 VDD.n6312 0.00326471
R10605 VDD.n6321 VDD.n485 0.00326471
R10606 VDD.n6351 VDD.n471 0.00326471
R10607 VDD.n6359 VDD.n6358 0.00326471
R10608 VDD.n6380 VDD.n6379 0.00326471
R10609 VDD.n6404 VDD.n6403 0.00326471
R10610 VDD.n6539 VDD.n6538 0.00326471
R10611 VDD.n6547 VDD.n351 0.00326471
R10612 VDD.n6577 VDD.n337 0.00326471
R10613 VDD.n6585 VDD.n6584 0.00326471
R10614 VDD.n6606 VDD.n6605 0.00326471
R10615 VDD.n6630 VDD.n6629 0.00326471
R10616 VDD.n6765 VDD.n6764 0.00326471
R10617 VDD.n6773 VDD.n217 0.00326471
R10618 VDD.n6803 VDD.n203 0.00326471
R10619 VDD.n6811 VDD.n6810 0.00326471
R10620 VDD.n6832 VDD.n6831 0.00326471
R10621 VDD.n6856 VDD.n6855 0.00326471
R10622 VDD.n6991 VDD.n6990 0.00326471
R10623 VDD.n6999 VDD.n83 0.00326471
R10624 VDD.n7029 VDD.n69 0.00326471
R10625 VDD.n7037 VDD.n7036 0.00326471
R10626 VDD.n7062 VDD.n7061 0.00326471
R10627 VDD.n7093 VDD.n36 0.00326471
R10628 VDD.n7211 VDD.n7210 0.00326471
R10629 VDD.n7130 VDD.n7101 0.00326471
R10630 VDD.n7141 VDD.n7140 0.00326471
R10631 VDD.n7181 VDD.n7145 0.00326471
R10632 VDD.n7155 VDD.n7150 0.00326471
R10633 VDD.n2900 VDD.n2899 0.00326471
R10634 VDD.n4262 VDD.n2860 0.00326471
R10635 VDD.n2943 VDD.n2942 0.00326471
R10636 VDD.n4241 VDD.n2935 0.00326471
R10637 VDD.n2984 VDD.n2983 0.00326471
R10638 VDD.n4219 VDD.n2987 0.00326471
R10639 VDD.n3166 VDD.n3165 0.00326471
R10640 VDD.n4143 VDD.n3158 0.00326471
R10641 VDD.n3209 VDD.n3208 0.00326471
R10642 VDD.n4122 VDD.n3201 0.00326471
R10643 VDD.n3250 VDD.n3249 0.00326471
R10644 VDD.n4100 VDD.n3253 0.00326471
R10645 VDD.n3432 VDD.n3431 0.00326471
R10646 VDD.n4024 VDD.n3424 0.00326471
R10647 VDD.n3475 VDD.n3474 0.00326471
R10648 VDD.n4003 VDD.n3467 0.00326471
R10649 VDD.n3516 VDD.n3515 0.00326471
R10650 VDD.n3981 VDD.n3519 0.00326471
R10651 VDD.n3698 VDD.n3697 0.00326471
R10652 VDD.n3905 VDD.n3690 0.00326471
R10653 VDD.n3741 VDD.n3740 0.00326471
R10654 VDD.n3884 VDD.n3733 0.00326471
R10655 VDD.n3782 VDD.n3781 0.00326471
R10656 VDD.n1548 VDD.n1547 0.00326471
R10657 VDD.n4804 VDD.n1552 0.00326471
R10658 VDD.n1590 VDD.n1589 0.00326471
R10659 VDD.n4782 VDD.n1594 0.00326471
R10660 VDD.n1632 VDD.n1631 0.00326471
R10661 VDD.n4760 VDD.n1635 0.00326471
R10662 VDD.n1812 VDD.n1811 0.00326471
R10663 VDD.n4683 VDD.n1816 0.00326471
R10664 VDD.n1854 VDD.n1853 0.00326471
R10665 VDD.n4661 VDD.n1858 0.00326471
R10666 VDD.n1896 VDD.n1895 0.00326471
R10667 VDD.n4639 VDD.n1899 0.00326471
R10668 VDD.n2076 VDD.n2075 0.00326471
R10669 VDD.n4562 VDD.n2080 0.00326471
R10670 VDD.n2118 VDD.n2117 0.00326471
R10671 VDD.n4540 VDD.n2122 0.00326471
R10672 VDD.n2160 VDD.n2159 0.00326471
R10673 VDD.n4518 VDD.n2163 0.00326471
R10674 VDD.n2340 VDD.n2339 0.00326471
R10675 VDD.n4441 VDD.n2344 0.00326471
R10676 VDD.n2382 VDD.n2381 0.00326471
R10677 VDD.n4419 VDD.n2386 0.00326471
R10678 VDD.n2424 VDD.n2423 0.00326471
R10679 VDD.n5034 VDD.n1194 0.00257353
R10680 VDD.n5064 VDD.n1182 0.00257353
R10681 VDD.n5054 VDD.n1170 0.00257353
R10682 VDD.n5093 VDD.n1168 0.00257353
R10683 VDD.n5117 VDD.n1154 0.00257353
R10684 VDD.n5232 VDD.n1073 0.00257353
R10685 VDD.n5262 VDD.n1059 0.00257353
R10686 VDD.n5292 VDD.n1047 0.00257353
R10687 VDD.n5282 VDD.n1035 0.00257353
R10688 VDD.n5321 VDD.n1033 0.00257353
R10689 VDD.n5345 VDD.n1019 0.00257353
R10690 VDD.n5460 VDD.n938 0.00257353
R10691 VDD.n5490 VDD.n924 0.00257353
R10692 VDD.n5520 VDD.n912 0.00257353
R10693 VDD.n5510 VDD.n900 0.00257353
R10694 VDD.n5549 VDD.n898 0.00257353
R10695 VDD.n5573 VDD.n884 0.00257353
R10696 VDD.n5688 VDD.n803 0.00257353
R10697 VDD.n5718 VDD.n789 0.00257353
R10698 VDD.n5748 VDD.n777 0.00257353
R10699 VDD.n5738 VDD.n765 0.00257353
R10700 VDD.n5777 VDD.n763 0.00257353
R10701 VDD.n5800 VDD.n749 0.00257353
R10702 VDD.n6202 VDD.n561 0.00257353
R10703 VDD.n559 VDD.n549 0.00257353
R10704 VDD.n6232 VDD.n547 0.00257353
R10705 VDD.n6254 VDD.n533 0.00257353
R10706 VDD.n6274 VDD.n522 0.00257353
R10707 VDD.n6408 VDD.n437 0.00257353
R10708 VDD.n6428 VDD.n427 0.00257353
R10709 VDD.n425 VDD.n415 0.00257353
R10710 VDD.n6458 VDD.n413 0.00257353
R10711 VDD.n6480 VDD.n399 0.00257353
R10712 VDD.n6500 VDD.n388 0.00257353
R10713 VDD.n6634 VDD.n303 0.00257353
R10714 VDD.n6654 VDD.n293 0.00257353
R10715 VDD.n291 VDD.n281 0.00257353
R10716 VDD.n6684 VDD.n279 0.00257353
R10717 VDD.n6706 VDD.n265 0.00257353
R10718 VDD.n6726 VDD.n254 0.00257353
R10719 VDD.n6860 VDD.n169 0.00257353
R10720 VDD.n6880 VDD.n159 0.00257353
R10721 VDD.n157 VDD.n147 0.00257353
R10722 VDD.n6910 VDD.n145 0.00257353
R10723 VDD.n6932 VDD.n131 0.00257353
R10724 VDD.n6952 VDD.n120 0.00257353
R10725 VDD.n2746 VDD.n2743 0.00257353
R10726 VDD.n2797 VDD.n2796 0.00257353
R10727 VDD.n2804 VDD.n2783 0.00257353
R10728 VDD.n4301 VDD.n4300 0.00257353
R10729 VDD.n2873 VDD.n2866 0.00257353
R10730 VDD.n4218 VDD.n2988 0.00257353
R10731 VDD.n3039 VDD.n3038 0.00257353
R10732 VDD.n3046 VDD.n3025 0.00257353
R10733 VDD.n4190 VDD.n4189 0.00257353
R10734 VDD.n3108 VDD.n3107 0.00257353
R10735 VDD.n3115 VDD.n3089 0.00257353
R10736 VDD.n4099 VDD.n3254 0.00257353
R10737 VDD.n3305 VDD.n3304 0.00257353
R10738 VDD.n3312 VDD.n3291 0.00257353
R10739 VDD.n4071 VDD.n4070 0.00257353
R10740 VDD.n3374 VDD.n3373 0.00257353
R10741 VDD.n3381 VDD.n3355 0.00257353
R10742 VDD.n3980 VDD.n3520 0.00257353
R10743 VDD.n3571 VDD.n3570 0.00257353
R10744 VDD.n3578 VDD.n3557 0.00257353
R10745 VDD.n3952 VDD.n3951 0.00257353
R10746 VDD.n3640 VDD.n3639 0.00257353
R10747 VDD.n3647 VDD.n3621 0.00257353
R10748 VDD.n4387 VDD.n2432 0.00257353
R10749 VDD.n4381 VDD.n4380 0.00257353
R10750 VDD.n2671 VDD.n2670 0.00257353
R10751 VDD.n2678 VDD.n2652 0.00257353
R10752 VDD.n4354 VDD.n4353 0.00257353
R10753 VDD.n2732 VDD.n2724 0.00257353
R10754 VDD.n1423 VDD.n1422 0.00257353
R10755 VDD.n1430 VDD.n1405 0.00257353
R10756 VDD.n4852 VDD.n4851 0.00257353
R10757 VDD.n1492 VDD.n1491 0.00257353
R10758 VDD.n1499 VDD.n1473 0.00257353
R10759 VDD.n4759 VDD.n1636 0.00257353
R10760 VDD.n1687 VDD.n1686 0.00257353
R10761 VDD.n1694 VDD.n1673 0.00257353
R10762 VDD.n4731 VDD.n4730 0.00257353
R10763 VDD.n1756 VDD.n1755 0.00257353
R10764 VDD.n1763 VDD.n1737 0.00257353
R10765 VDD.n4638 VDD.n1900 0.00257353
R10766 VDD.n1951 VDD.n1950 0.00257353
R10767 VDD.n1958 VDD.n1937 0.00257353
R10768 VDD.n4610 VDD.n4609 0.00257353
R10769 VDD.n2020 VDD.n2019 0.00257353
R10770 VDD.n2027 VDD.n2001 0.00257353
R10771 VDD.n4517 VDD.n2164 0.00257353
R10772 VDD.n2215 VDD.n2214 0.00257353
R10773 VDD.n2222 VDD.n2201 0.00257353
R10774 VDD.n4489 VDD.n4488 0.00257353
R10775 VDD.n2284 VDD.n2283 0.00257353
R10776 VDD.n2291 VDD.n2265 0.00257353
R10777 VDD.n1279 VDD.n1278 0.00257353
R10778 VDD.n1296 VDD.n1295 0.00257353
R10779 VDD.n1303 VDD.n1257 0.00257353
R10780 VDD.n4904 VDD.n4903 0.00257353
R10781 VDD.n1365 VDD.n1364 0.00257353
R10782 VDD.n1372 VDD.n1346 0.00257353
R10783 VDD.n4394 VDD 0.00252392
R10784 VDD.n4979 VDD 0.00252392
R10785 VDD.n5026 VDD.n1191 0.00239394
R10786 VDD.n5047 VDD.n1178 0.00239394
R10787 VDD.n5060 VDD.n1173 0.00239394
R10788 VDD.n5099 VDD.n5098 0.00239394
R10789 VDD.n5108 VDD.n1151 0.00239394
R10790 VDD.n5129 VDD.n1129 0.00239394
R10791 VDD.n1141 VDD.n1120 0.00239394
R10792 VDD.n5150 VDD.n1114 0.00239394
R10793 VDD.n5182 VDD.n1100 0.00239394
R10794 VDD.n5191 VDD.n1094 0.00239394
R10795 VDD.n5204 VDD.n1080 0.00239394
R10796 VDD.n5242 VDD.n1067 0.00239394
R10797 VDD.n5254 VDD.n1056 0.00239394
R10798 VDD.n5275 VDD.n1043 0.00239394
R10799 VDD.n5288 VDD.n1038 0.00239394
R10800 VDD.n5327 VDD.n5326 0.00239394
R10801 VDD.n5336 VDD.n1016 0.00239394
R10802 VDD.n5357 VDD.n994 0.00239394
R10803 VDD.n1006 VDD.n985 0.00239394
R10804 VDD.n5378 VDD.n979 0.00239394
R10805 VDD.n5410 VDD.n965 0.00239394
R10806 VDD.n5419 VDD.n959 0.00239394
R10807 VDD.n5432 VDD.n945 0.00239394
R10808 VDD.n5470 VDD.n932 0.00239394
R10809 VDD.n5482 VDD.n921 0.00239394
R10810 VDD.n5503 VDD.n908 0.00239394
R10811 VDD.n5516 VDD.n903 0.00239394
R10812 VDD.n5555 VDD.n5554 0.00239394
R10813 VDD.n5564 VDD.n881 0.00239394
R10814 VDD.n5585 VDD.n859 0.00239394
R10815 VDD.n871 VDD.n850 0.00239394
R10816 VDD.n5606 VDD.n844 0.00239394
R10817 VDD.n5638 VDD.n830 0.00239394
R10818 VDD.n5647 VDD.n824 0.00239394
R10819 VDD.n5660 VDD.n810 0.00239394
R10820 VDD.n5698 VDD.n797 0.00239394
R10821 VDD.n5710 VDD.n786 0.00239394
R10822 VDD.n5731 VDD.n773 0.00239394
R10823 VDD.n5744 VDD.n768 0.00239394
R10824 VDD.n5783 VDD.n5782 0.00239394
R10825 VDD.n5792 VDD.n746 0.00239394
R10826 VDD.n5812 VDD.n733 0.00239394
R10827 VDD.n5823 VDD.n725 0.00239394
R10828 VDD.n5845 VDD.n717 0.00239394
R10829 VDD.n708 VDD.n699 0.00239394
R10830 VDD.n5879 VDD.n693 0.00239394
R10831 VDD.n5915 VDD.n677 0.00239394
R10832 VDD.n5923 VDD.n671 0.00239394
R10833 VDD.n6065 VDD.n657 0.00239394
R10834 VDD.n5962 VDD.n5954 0.00239394
R10835 VDD.n6048 VDD.n5957 0.00239394
R10836 VDD.n6039 VDD.n5972 0.00239394
R10837 VDD.n6027 VDD.n6010 0.00239394
R10838 VDD.n5934 VDD.n658 0.00239394
R10839 VDD.n5961 VDD.n5952 0.00239394
R10840 VDD.n6049 VDD.n5956 0.00239394
R10841 VDD.n6038 VDD.n6037 0.00239394
R10842 VDD.n6028 VDD.n5997 0.00239394
R10843 VDD.n6190 VDD.n563 0.00239394
R10844 VDD.n6211 VDD.n552 0.00239394
R10845 VDD.n6238 VDD.n6237 0.00239394
R10846 VDD.n6246 VDD.n530 0.00239394
R10847 VDD.n6266 VDD.n519 0.00239394
R10848 VDD.n6285 VDD.n506 0.00239394
R10849 VDD.n6296 VDD.n497 0.00239394
R10850 VDD.n491 VDD.n482 0.00239394
R10851 VDD.n6331 VDD.n476 0.00239394
R10852 VDD.n6363 VDD.n462 0.00239394
R10853 VDD.n6372 VDD.n457 0.00239394
R10854 VDD.n6396 VDD.n444 0.00239394
R10855 VDD.n6416 VDD.n429 0.00239394
R10856 VDD.n6437 VDD.n418 0.00239394
R10857 VDD.n6464 VDD.n6463 0.00239394
R10858 VDD.n6472 VDD.n396 0.00239394
R10859 VDD.n6492 VDD.n385 0.00239394
R10860 VDD.n6511 VDD.n372 0.00239394
R10861 VDD.n6522 VDD.n363 0.00239394
R10862 VDD.n357 VDD.n348 0.00239394
R10863 VDD.n6557 VDD.n342 0.00239394
R10864 VDD.n6589 VDD.n328 0.00239394
R10865 VDD.n6598 VDD.n323 0.00239394
R10866 VDD.n6622 VDD.n310 0.00239394
R10867 VDD.n6642 VDD.n295 0.00239394
R10868 VDD.n6663 VDD.n284 0.00239394
R10869 VDD.n6690 VDD.n6689 0.00239394
R10870 VDD.n6698 VDD.n262 0.00239394
R10871 VDD.n6718 VDD.n251 0.00239394
R10872 VDD.n6737 VDD.n238 0.00239394
R10873 VDD.n6748 VDD.n229 0.00239394
R10874 VDD.n223 VDD.n214 0.00239394
R10875 VDD.n6783 VDD.n208 0.00239394
R10876 VDD.n6815 VDD.n194 0.00239394
R10877 VDD.n6824 VDD.n189 0.00239394
R10878 VDD.n6848 VDD.n176 0.00239394
R10879 VDD.n6868 VDD.n161 0.00239394
R10880 VDD.n6889 VDD.n150 0.00239394
R10881 VDD.n6916 VDD.n6915 0.00239394
R10882 VDD.n6924 VDD.n128 0.00239394
R10883 VDD.n6944 VDD.n117 0.00239394
R10884 VDD.n6963 VDD.n104 0.00239394
R10885 VDD.n6974 VDD.n95 0.00239394
R10886 VDD.n89 VDD.n80 0.00239394
R10887 VDD.n7009 VDD.n74 0.00239394
R10888 VDD.n7041 VDD.n60 0.00239394
R10889 VDD.n7050 VDD.n55 0.00239394
R10890 VDD.n7073 VDD.n42 0.00239394
R10891 VDD.n6189 VDD.n562 0.00239394
R10892 VDD.n6210 VDD.n551 0.00239394
R10893 VDD.n6236 VDD.n543 0.00239394
R10894 VDD.n6247 VDD.n531 0.00239394
R10895 VDD.n6267 VDD.n520 0.00239394
R10896 VDD.n6286 VDD.n504 0.00239394
R10897 VDD.n6295 VDD.n498 0.00239394
R10898 VDD.n489 VDD.n483 0.00239394
R10899 VDD.n6330 VDD.n474 0.00239394
R10900 VDD.n6342 VDD.n463 0.00239394
R10901 VDD.n6373 VDD.n455 0.00239394
R10902 VDD.n6397 VDD.n442 0.00239394
R10903 VDD.n6415 VDD.n428 0.00239394
R10904 VDD.n6436 VDD.n417 0.00239394
R10905 VDD.n6462 VDD.n409 0.00239394
R10906 VDD.n6473 VDD.n397 0.00239394
R10907 VDD.n6493 VDD.n386 0.00239394
R10908 VDD.n6512 VDD.n370 0.00239394
R10909 VDD.n6521 VDD.n364 0.00239394
R10910 VDD.n355 VDD.n349 0.00239394
R10911 VDD.n6556 VDD.n340 0.00239394
R10912 VDD.n6568 VDD.n329 0.00239394
R10913 VDD.n6599 VDD.n321 0.00239394
R10914 VDD.n6623 VDD.n308 0.00239394
R10915 VDD.n6641 VDD.n294 0.00239394
R10916 VDD.n6662 VDD.n283 0.00239394
R10917 VDD.n6688 VDD.n275 0.00239394
R10918 VDD.n6699 VDD.n263 0.00239394
R10919 VDD.n6719 VDD.n252 0.00239394
R10920 VDD.n6738 VDD.n236 0.00239394
R10921 VDD.n6747 VDD.n230 0.00239394
R10922 VDD.n221 VDD.n215 0.00239394
R10923 VDD.n6782 VDD.n206 0.00239394
R10924 VDD.n6794 VDD.n195 0.00239394
R10925 VDD.n6825 VDD.n187 0.00239394
R10926 VDD.n6849 VDD.n174 0.00239394
R10927 VDD.n6867 VDD.n160 0.00239394
R10928 VDD.n6888 VDD.n149 0.00239394
R10929 VDD.n6914 VDD.n141 0.00239394
R10930 VDD.n6925 VDD.n129 0.00239394
R10931 VDD.n6945 VDD.n118 0.00239394
R10932 VDD.n6964 VDD.n102 0.00239394
R10933 VDD.n6973 VDD.n96 0.00239394
R10934 VDD.n87 VDD.n81 0.00239394
R10935 VDD.n7008 VDD.n72 0.00239394
R10936 VDD.n7020 VDD.n61 0.00239394
R10937 VDD.n7051 VDD.n53 0.00239394
R10938 VDD.n7064 VDD.n43 0.00239394
R10939 VDD.n7215 VDD.n28 0.00239394
R10940 VDD.n7112 VDD.n7104 0.00239394
R10941 VDD.n7198 VDD.n7107 0.00239394
R10942 VDD.n7189 VDD.n7122 0.00239394
R10943 VDD.n7177 VDD.n7160 0.00239394
R10944 VDD.n7084 VDD.n29 0.00239394
R10945 VDD.n7111 VDD.n7102 0.00239394
R10946 VDD.n7199 VDD.n7106 0.00239394
R10947 VDD.n7188 VDD.n7187 0.00239394
R10948 VDD.n7178 VDD.n7147 0.00239394
R10949 VDD.n4333 VDD.n2740 0.00239394
R10950 VDD.n4323 VDD.n2752 0.00239394
R10951 VDD.n4314 VDD.n4313 0.00239394
R10952 VDD.n2830 VDD.n2781 0.00239394
R10953 VDD.n4296 VDD.n2813 0.00239394
R10954 VDD.n4287 VDD.n4286 0.00239394
R10955 VDD.n2848 VDD.n2845 0.00239394
R10956 VDD.n4269 VDD.n2855 0.00239394
R10957 VDD.n4258 VDD.n2908 0.00239394
R10958 VDD.n4248 VDD.n2930 0.00239394
R10959 VDD.n4237 VDD.n2951 0.00239394
R10960 VDD.n4227 VDD.n2973 0.00239394
R10961 VDD.n4212 VDD.n2999 0.00239394
R10962 VDD.n4203 VDD.n4202 0.00239394
R10963 VDD.n3072 VDD.n3023 0.00239394
R10964 VDD.n4185 VDD.n3055 0.00239394
R10965 VDD.n4176 VDD.n4175 0.00239394
R10966 VDD.n3143 VDD.n3087 0.00239394
R10967 VDD.n4160 VDD.n3122 0.00239394
R10968 VDD.n4150 VDD.n3153 0.00239394
R10969 VDD.n4139 VDD.n3174 0.00239394
R10970 VDD.n4129 VDD.n3196 0.00239394
R10971 VDD.n4118 VDD.n3217 0.00239394
R10972 VDD.n4108 VDD.n3239 0.00239394
R10973 VDD.n4093 VDD.n3265 0.00239394
R10974 VDD.n4084 VDD.n4083 0.00239394
R10975 VDD.n3338 VDD.n3289 0.00239394
R10976 VDD.n4066 VDD.n3321 0.00239394
R10977 VDD.n4057 VDD.n4056 0.00239394
R10978 VDD.n3409 VDD.n3353 0.00239394
R10979 VDD.n4041 VDD.n3388 0.00239394
R10980 VDD.n4031 VDD.n3419 0.00239394
R10981 VDD.n4020 VDD.n3440 0.00239394
R10982 VDD.n4010 VDD.n3462 0.00239394
R10983 VDD.n3999 VDD.n3483 0.00239394
R10984 VDD.n3989 VDD.n3505 0.00239394
R10985 VDD.n3974 VDD.n3531 0.00239394
R10986 VDD.n3965 VDD.n3964 0.00239394
R10987 VDD.n3604 VDD.n3555 0.00239394
R10988 VDD.n3947 VDD.n3587 0.00239394
R10989 VDD.n3938 VDD.n3937 0.00239394
R10990 VDD.n3675 VDD.n3619 0.00239394
R10991 VDD.n3922 VDD.n3654 0.00239394
R10992 VDD.n3912 VDD.n3685 0.00239394
R10993 VDD.n3901 VDD.n3706 0.00239394
R10994 VDD.n3891 VDD.n3728 0.00239394
R10995 VDD.n3880 VDD.n3749 0.00239394
R10996 VDD.n3870 VDD.n3771 0.00239394
R10997 VDD.n2635 VDD.n2632 0.00239394
R10998 VDD.n4376 VDD.n2444 0.00239394
R10999 VDD.n4367 VDD.n4366 0.00239394
R11000 VDD.n2704 VDD.n2650 0.00239394
R11001 VDD.n4349 VDD.n2687 0.00239394
R11002 VDD.n2634 VDD.n2633 0.00239394
R11003 VDD.n2662 VDD.n2443 0.00239394
R11004 VDD.n4365 VDD.n2647 0.00239394
R11005 VDD.n2703 VDD.n2651 0.00239394
R11006 VDD.n2725 VDD.n2686 0.00239394
R11007 VDD.n4874 VDD.n1378 0.00239394
R11008 VDD.n4865 VDD.n4864 0.00239394
R11009 VDD.n1456 VDD.n1403 0.00239394
R11010 VDD.n4847 VDD.n1439 0.00239394
R11011 VDD.n4838 VDD.n4837 0.00239394
R11012 VDD.n1527 VDD.n1471 0.00239394
R11013 VDD.n4822 VDD.n1506 0.00239394
R11014 VDD.n4812 VDD.n1537 0.00239394
R11015 VDD.n4800 VDD.n1556 0.00239394
R11016 VDD.n4790 VDD.n1579 0.00239394
R11017 VDD.n4778 VDD.n1598 0.00239394
R11018 VDD.n4768 VDD.n1621 0.00239394
R11019 VDD.n4753 VDD.n1647 0.00239394
R11020 VDD.n4744 VDD.n4743 0.00239394
R11021 VDD.n1720 VDD.n1671 0.00239394
R11022 VDD.n4726 VDD.n1703 0.00239394
R11023 VDD.n4717 VDD.n4716 0.00239394
R11024 VDD.n1791 VDD.n1735 0.00239394
R11025 VDD.n4701 VDD.n1770 0.00239394
R11026 VDD.n4691 VDD.n1801 0.00239394
R11027 VDD.n4679 VDD.n1820 0.00239394
R11028 VDD.n4669 VDD.n1843 0.00239394
R11029 VDD.n4657 VDD.n1862 0.00239394
R11030 VDD.n4647 VDD.n1885 0.00239394
R11031 VDD.n4632 VDD.n1911 0.00239394
R11032 VDD.n4623 VDD.n4622 0.00239394
R11033 VDD.n1984 VDD.n1935 0.00239394
R11034 VDD.n4605 VDD.n1967 0.00239394
R11035 VDD.n4596 VDD.n4595 0.00239394
R11036 VDD.n2055 VDD.n1999 0.00239394
R11037 VDD.n4580 VDD.n2034 0.00239394
R11038 VDD.n4570 VDD.n2065 0.00239394
R11039 VDD.n4558 VDD.n2084 0.00239394
R11040 VDD.n4548 VDD.n2107 0.00239394
R11041 VDD.n4536 VDD.n2126 0.00239394
R11042 VDD.n4526 VDD.n2149 0.00239394
R11043 VDD.n4511 VDD.n2175 0.00239394
R11044 VDD.n4502 VDD.n4501 0.00239394
R11045 VDD.n2248 VDD.n2199 0.00239394
R11046 VDD.n4484 VDD.n2231 0.00239394
R11047 VDD.n4475 VDD.n4474 0.00239394
R11048 VDD.n2319 VDD.n2263 0.00239394
R11049 VDD.n4459 VDD.n2298 0.00239394
R11050 VDD.n4449 VDD.n2329 0.00239394
R11051 VDD.n4437 VDD.n2348 0.00239394
R11052 VDD.n4427 VDD.n2371 0.00239394
R11053 VDD.n4415 VDD.n2390 0.00239394
R11054 VDD.n4405 VDD.n2413 0.00239394
R11055 VDD.n1414 VDD.n1377 0.00239394
R11056 VDD.n4863 VDD.n1400 0.00239394
R11057 VDD.n1455 VDD.n1404 0.00239394
R11058 VDD.n1483 VDD.n1438 0.00239394
R11059 VDD.n4836 VDD.n1468 0.00239394
R11060 VDD.n1526 VDD.n1472 0.00239394
R11061 VDD.n4823 VDD.n1504 0.00239394
R11062 VDD.n4811 VDD.n4810 0.00239394
R11063 VDD.n4801 VDD.n1554 0.00239394
R11064 VDD.n4789 VDD.n4788 0.00239394
R11065 VDD.n4779 VDD.n1596 0.00239394
R11066 VDD.n4767 VDD.n4766 0.00239394
R11067 VDD.n4754 VDD.n1640 0.00239394
R11068 VDD.n4742 VDD.n1668 0.00239394
R11069 VDD.n1719 VDD.n1672 0.00239394
R11070 VDD.n1747 VDD.n1702 0.00239394
R11071 VDD.n4715 VDD.n1732 0.00239394
R11072 VDD.n1790 VDD.n1736 0.00239394
R11073 VDD.n4702 VDD.n1768 0.00239394
R11074 VDD.n4690 VDD.n4689 0.00239394
R11075 VDD.n4680 VDD.n1818 0.00239394
R11076 VDD.n4668 VDD.n4667 0.00239394
R11077 VDD.n4658 VDD.n1860 0.00239394
R11078 VDD.n4646 VDD.n4645 0.00239394
R11079 VDD.n4633 VDD.n1904 0.00239394
R11080 VDD.n4621 VDD.n1932 0.00239394
R11081 VDD.n1983 VDD.n1936 0.00239394
R11082 VDD.n2011 VDD.n1966 0.00239394
R11083 VDD.n4594 VDD.n1996 0.00239394
R11084 VDD.n2054 VDD.n2000 0.00239394
R11085 VDD.n4581 VDD.n2032 0.00239394
R11086 VDD.n4569 VDD.n4568 0.00239394
R11087 VDD.n4559 VDD.n2082 0.00239394
R11088 VDD.n4547 VDD.n4546 0.00239394
R11089 VDD.n4537 VDD.n2124 0.00239394
R11090 VDD.n4525 VDD.n4524 0.00239394
R11091 VDD.n4512 VDD.n2168 0.00239394
R11092 VDD.n4500 VDD.n2196 0.00239394
R11093 VDD.n2247 VDD.n2200 0.00239394
R11094 VDD.n2275 VDD.n2230 0.00239394
R11095 VDD.n4473 VDD.n2260 0.00239394
R11096 VDD.n2318 VDD.n2264 0.00239394
R11097 VDD.n4460 VDD.n2296 0.00239394
R11098 VDD.n4448 VDD.n4447 0.00239394
R11099 VDD.n4438 VDD.n2346 0.00239394
R11100 VDD.n4426 VDD.n4425 0.00239394
R11101 VDD.n4416 VDD.n2388 0.00239394
R11102 VDD.n4404 VDD.n4403 0.00239394
R11103 VDD.n1287 VDD.n1245 0.00239394
R11104 VDD.n4917 VDD.n4916 0.00239394
R11105 VDD.n1329 VDD.n1255 0.00239394
R11106 VDD.n4899 VDD.n1312 0.00239394
R11107 VDD.n4890 VDD.n4889 0.00239394
R11108 VDD.n1286 VDD.n1285 0.00239394
R11109 VDD.n4915 VDD.n1252 0.00239394
R11110 VDD.n1328 VDD.n1256 0.00239394
R11111 VDD.n1356 VDD.n1311 0.00239394
R11112 VDD.n4888 VDD.n1341 0.00239394
R11113 VDD.n4332 VDD.n2741 0.00239394
R11114 VDD.n4324 VDD.n2749 0.00239394
R11115 VDD.n4312 VDD.n2778 0.00239394
R11116 VDD.n2829 VDD.n2782 0.00239394
R11117 VDD.n2876 VDD.n2812 0.00239394
R11118 VDD.n4285 VDD.n2842 0.00239394
R11119 VDD.n2894 VDD.n2863 0.00239394
R11120 VDD.n4268 VDD.n4267 0.00239394
R11121 VDD.n4259 VDD.n2906 0.00239394
R11122 VDD.n4247 VDD.n4246 0.00239394
R11123 VDD.n4238 VDD.n2949 0.00239394
R11124 VDD.n4226 VDD.n4225 0.00239394
R11125 VDD.n4213 VDD.n2993 0.00239394
R11126 VDD.n4201 VDD.n3020 0.00239394
R11127 VDD.n3071 VDD.n3024 0.00239394
R11128 VDD.n3099 VDD.n3054 0.00239394
R11129 VDD.n4174 VDD.n3084 0.00239394
R11130 VDD.n3142 VDD.n3088 0.00239394
R11131 VDD.n4161 VDD.n3120 0.00239394
R11132 VDD.n4149 VDD.n4148 0.00239394
R11133 VDD.n4140 VDD.n3172 0.00239394
R11134 VDD.n4128 VDD.n4127 0.00239394
R11135 VDD.n4119 VDD.n3215 0.00239394
R11136 VDD.n4107 VDD.n4106 0.00239394
R11137 VDD.n4094 VDD.n3259 0.00239394
R11138 VDD.n4082 VDD.n3286 0.00239394
R11139 VDD.n3337 VDD.n3290 0.00239394
R11140 VDD.n3365 VDD.n3320 0.00239394
R11141 VDD.n4055 VDD.n3350 0.00239394
R11142 VDD.n3408 VDD.n3354 0.00239394
R11143 VDD.n4042 VDD.n3386 0.00239394
R11144 VDD.n4030 VDD.n4029 0.00239394
R11145 VDD.n4021 VDD.n3438 0.00239394
R11146 VDD.n4009 VDD.n4008 0.00239394
R11147 VDD.n4000 VDD.n3481 0.00239394
R11148 VDD.n3988 VDD.n3987 0.00239394
R11149 VDD.n3975 VDD.n3525 0.00239394
R11150 VDD.n3963 VDD.n3552 0.00239394
R11151 VDD.n3603 VDD.n3556 0.00239394
R11152 VDD.n3631 VDD.n3586 0.00239394
R11153 VDD.n3936 VDD.n3616 0.00239394
R11154 VDD.n3674 VDD.n3620 0.00239394
R11155 VDD.n3923 VDD.n3652 0.00239394
R11156 VDD.n3911 VDD.n3910 0.00239394
R11157 VDD.n3902 VDD.n3704 0.00239394
R11158 VDD.n3890 VDD.n3889 0.00239394
R11159 VDD.n3881 VDD.n3747 0.00239394
R11160 VDD.n3869 VDD.n3868 0.00239394
R11161 VDD.n5027 VDD.n1192 0.00239394
R11162 VDD.n5048 VDD.n1180 0.00239394
R11163 VDD.n5061 VDD.n1172 0.00239394
R11164 VDD.n5097 VDD.n1164 0.00239394
R11165 VDD.n5109 VDD.n1152 0.00239394
R11166 VDD.n5130 VDD.n1127 0.00239394
R11167 VDD.n1142 VDD.n1121 0.00239394
R11168 VDD.n5149 VDD.n1112 0.00239394
R11169 VDD.n5161 VDD.n1101 0.00239394
R11170 VDD.n5192 VDD.n1092 0.00239394
R11171 VDD.n5203 VDD.n1078 0.00239394
R11172 VDD.n5217 VDD.n1068 0.00239394
R11173 VDD.n5255 VDD.n1057 0.00239394
R11174 VDD.n5276 VDD.n1045 0.00239394
R11175 VDD.n5289 VDD.n1037 0.00239394
R11176 VDD.n5325 VDD.n1029 0.00239394
R11177 VDD.n5337 VDD.n1017 0.00239394
R11178 VDD.n5358 VDD.n992 0.00239394
R11179 VDD.n1007 VDD.n986 0.00239394
R11180 VDD.n5377 VDD.n977 0.00239394
R11181 VDD.n5389 VDD.n966 0.00239394
R11182 VDD.n5420 VDD.n957 0.00239394
R11183 VDD.n5431 VDD.n943 0.00239394
R11184 VDD.n5445 VDD.n933 0.00239394
R11185 VDD.n5483 VDD.n922 0.00239394
R11186 VDD.n5504 VDD.n910 0.00239394
R11187 VDD.n5517 VDD.n902 0.00239394
R11188 VDD.n5553 VDD.n894 0.00239394
R11189 VDD.n5565 VDD.n882 0.00239394
R11190 VDD.n5586 VDD.n857 0.00239394
R11191 VDD.n872 VDD.n851 0.00239394
R11192 VDD.n5605 VDD.n842 0.00239394
R11193 VDD.n5617 VDD.n831 0.00239394
R11194 VDD.n5648 VDD.n822 0.00239394
R11195 VDD.n5659 VDD.n808 0.00239394
R11196 VDD.n5673 VDD.n798 0.00239394
R11197 VDD.n5711 VDD.n787 0.00239394
R11198 VDD.n5732 VDD.n775 0.00239394
R11199 VDD.n5745 VDD.n767 0.00239394
R11200 VDD.n5781 VDD.n759 0.00239394
R11201 VDD.n5793 VDD.n747 0.00239394
R11202 VDD.n5813 VDD.n731 0.00239394
R11203 VDD.n5822 VDD.n726 0.00239394
R11204 VDD.n5844 VDD.n718 0.00239394
R11205 VDD.n706 VDD.n700 0.00239394
R11206 VDD.n5878 VDD.n691 0.00239394
R11207 VDD.n5890 VDD.n678 0.00239394
R11208 VDD.n683 VDD.n672 0.00239394
R11209 VDD.n3844 VDD.n3830 0.0021514
R11210 VDD.n2520 VDD.n2506 0.0021514
R11211 VDD.n6004 VDD.n6003 0.00213953
R11212 VDD.n7154 VDD.n7153 0.00213953
R11213 VDD.n4390 VDD.n2430 0.00213953
R11214 VDD.n1268 VDD.n1265 0.00213953
R11215 VDD.n614 VDD.n612 0.00196875
R11216 VDD.n6116 VDD.n6115 0.00196875
R11217 VDD.n6180 VDD.n6179 0.00196875
R11218 VDD.n2467 VDD.n2463 0.00196875
R11219 VDD.n2612 VDD.n2461 0.00196875
R11220 VDD.n4944 VDD.n4942 0.00196875
R11221 VDD.n4948 VDD.n4937 0.00196875
R11222 VDD.n5019 VDD.n5018 0.00196875
R11223 VDD.n7243 VDD.n7242 0.00196875
R11224 VDD.n7261 VDD.n7260 0.00196875
R11225 VDD VDD.n7231 0.00196114
R11226 VDD VDD.n6081 0.00196114
R11227 VDD.n6110 VDD.n599 0.00192033
R11228 VDD.n6138 VDD.n6137 0.00175893
R11229 VDD.n6175 VDD.n568 0.00175893
R11230 VDD.n6179 VDD.n568 0.00175893
R11231 VDD.n4981 VDD.n4980 0.00175893
R11232 VDD.n5014 VDD.n1198 0.00175893
R11233 VDD.n5018 VDD.n1198 0.00175893
R11234 VDD.n6104 VDD.n6103 0.00172665
R11235 VDD.n627 VDD.n615 0.00172665
R11236 VDD.n6168 VDD.n6167 0.00150714
R11237 VDD.n580 VDD.n579 0.00150714
R11238 VDD.n5007 VDD.n5006 0.00150714
R11239 VDD.n1210 VDD.n1209 0.00150714
R11240 VDD.n7232 VDD 0.00123057
R11241 VDD.n6082 VDD 0.00123057
R11242 VDD.n6175 VDD.n6174 0.00121339
R11243 VDD.n5014 VDD.n5013 0.00121339
R11244 VDD.n6104 VDD.n620 0.00121017
R11245 VDD.n6103 VDD.n627 0.00121017
R11246 VDD.n5022 VDD.n1196 0.00119118
R11247 VDD.n5028 VDD.n1196 0.00119118
R11248 VDD.n5033 VDD.n1185 0.00119118
R11249 VDD.n5049 VDD.n1185 0.00119118
R11250 VDD.n5063 VDD.n1183 0.00119118
R11251 VDD.n5059 VDD.n1183 0.00119118
R11252 VDD.n5086 VDD.n5085 0.00119118
R11253 VDD.n5087 VDD.n5086 0.00119118
R11254 VDD.n5092 VDD.n1156 0.00119118
R11255 VDD.n5110 VDD.n1156 0.00119118
R11256 VDD.n5116 VDD.n1125 0.00119118
R11257 VDD.n5131 VDD.n1125 0.00119118
R11258 VDD.n5133 VDD.n1122 0.00119118
R11259 VDD.n5143 VDD.n1122 0.00119118
R11260 VDD.n5138 VDD.n1111 0.00119118
R11261 VDD.n5167 VDD.n1111 0.00119118
R11262 VDD.n5173 VDD.n5172 0.00119118
R11263 VDD.n5173 VDD.n1107 0.00119118
R11264 VDD.n5194 VDD.n5193 0.00119118
R11265 VDD.n5194 VDD.n1087 0.00119118
R11266 VDD.n1088 VDD.n1077 0.00119118
R11267 VDD.n5223 VDD.n1077 0.00119118
R11268 VDD.n5229 VDD.n5228 0.00119118
R11269 VDD.n5229 VDD.n1072 0.00119118
R11270 VDD.n5233 VDD.n1061 0.00119118
R11271 VDD.n5256 VDD.n1061 0.00119118
R11272 VDD.n5261 VDD.n1050 0.00119118
R11273 VDD.n5277 VDD.n1050 0.00119118
R11274 VDD.n5291 VDD.n1048 0.00119118
R11275 VDD.n5287 VDD.n1048 0.00119118
R11276 VDD.n5314 VDD.n5313 0.00119118
R11277 VDD.n5315 VDD.n5314 0.00119118
R11278 VDD.n5320 VDD.n1021 0.00119118
R11279 VDD.n5338 VDD.n1021 0.00119118
R11280 VDD.n5344 VDD.n990 0.00119118
R11281 VDD.n5359 VDD.n990 0.00119118
R11282 VDD.n5361 VDD.n987 0.00119118
R11283 VDD.n5371 VDD.n987 0.00119118
R11284 VDD.n5366 VDD.n976 0.00119118
R11285 VDD.n5395 VDD.n976 0.00119118
R11286 VDD.n5401 VDD.n5400 0.00119118
R11287 VDD.n5401 VDD.n972 0.00119118
R11288 VDD.n5422 VDD.n5421 0.00119118
R11289 VDD.n5422 VDD.n952 0.00119118
R11290 VDD.n953 VDD.n942 0.00119118
R11291 VDD.n5451 VDD.n942 0.00119118
R11292 VDD.n5457 VDD.n5456 0.00119118
R11293 VDD.n5457 VDD.n937 0.00119118
R11294 VDD.n5461 VDD.n926 0.00119118
R11295 VDD.n5484 VDD.n926 0.00119118
R11296 VDD.n5489 VDD.n915 0.00119118
R11297 VDD.n5505 VDD.n915 0.00119118
R11298 VDD.n5519 VDD.n913 0.00119118
R11299 VDD.n5515 VDD.n913 0.00119118
R11300 VDD.n5542 VDD.n5541 0.00119118
R11301 VDD.n5543 VDD.n5542 0.00119118
R11302 VDD.n5548 VDD.n886 0.00119118
R11303 VDD.n5566 VDD.n886 0.00119118
R11304 VDD.n5572 VDD.n855 0.00119118
R11305 VDD.n5587 VDD.n855 0.00119118
R11306 VDD.n5589 VDD.n852 0.00119118
R11307 VDD.n5599 VDD.n852 0.00119118
R11308 VDD.n5594 VDD.n841 0.00119118
R11309 VDD.n5623 VDD.n841 0.00119118
R11310 VDD.n5629 VDD.n5628 0.00119118
R11311 VDD.n5629 VDD.n837 0.00119118
R11312 VDD.n5650 VDD.n5649 0.00119118
R11313 VDD.n5650 VDD.n817 0.00119118
R11314 VDD.n818 VDD.n807 0.00119118
R11315 VDD.n5679 VDD.n807 0.00119118
R11316 VDD.n5685 VDD.n5684 0.00119118
R11317 VDD.n5685 VDD.n802 0.00119118
R11318 VDD.n5689 VDD.n791 0.00119118
R11319 VDD.n5712 VDD.n791 0.00119118
R11320 VDD.n5717 VDD.n780 0.00119118
R11321 VDD.n5733 VDD.n780 0.00119118
R11322 VDD.n5747 VDD.n778 0.00119118
R11323 VDD.n5743 VDD.n778 0.00119118
R11324 VDD.n5770 VDD.n5769 0.00119118
R11325 VDD.n5771 VDD.n5770 0.00119118
R11326 VDD.n5776 VDD.n751 0.00119118
R11327 VDD.n5794 VDD.n751 0.00119118
R11328 VDD.n5799 VDD.n729 0.00119118
R11329 VDD.n5814 VDD.n729 0.00119118
R11330 VDD.n5820 VDD.n5819 0.00119118
R11331 VDD.n5819 VDD.n721 0.00119118
R11332 VDD.n5842 VDD.n5841 0.00119118
R11333 VDD.n5841 VDD.n704 0.00119118
R11334 VDD.n5862 VDD.n701 0.00119118
R11335 VDD.n5872 VDD.n701 0.00119118
R11336 VDD.n5867 VDD.n690 0.00119118
R11337 VDD.n5896 VDD.n690 0.00119118
R11338 VDD.n5902 VDD.n5901 0.00119118
R11339 VDD.n5902 VDD.n685 0.00119118
R11340 VDD.n5906 VDD.n5905 0.00119118
R11341 VDD.n5906 VDD.n669 0.00119118
R11342 VDD.n5930 VDD.n667 0.00119118
R11343 VDD.n5940 VDD.n667 0.00119118
R11344 VDD.n5946 VDD.n5945 0.00119118
R11345 VDD.n5946 VDD.n662 0.00119118
R11346 VDD.n6056 VDD.n5950 0.00119118
R11347 VDD.n6056 VDD.n6055 0.00119118
R11348 VDD.n5984 VDD.n5978 0.00119118
R11349 VDD.n5985 VDD.n5984 0.00119118
R11350 VDD.n6036 VDD.n6035 0.00119118
R11351 VDD.n6035 VDD.n5976 0.00119118
R11352 VDD.n6029 VDD.n5996 0.00119118
R11353 VDD.n6008 VDD.n5996 0.00119118
R11354 VDD.n6183 VDD.n567 0.00119118
R11355 VDD.n6188 VDD.n567 0.00119118
R11356 VDD.n6203 VDD.n558 0.00119118
R11357 VDD.n6209 VDD.n558 0.00119118
R11358 VDD.n6225 VDD.n6224 0.00119118
R11359 VDD.n6226 VDD.n6225 0.00119118
R11360 VDD.n6231 VDD.n535 0.00119118
R11361 VDD.n6248 VDD.n535 0.00119118
R11362 VDD.n6253 VDD.n524 0.00119118
R11363 VDD.n6268 VDD.n524 0.00119118
R11364 VDD.n6273 VDD.n502 0.00119118
R11365 VDD.n6287 VDD.n502 0.00119118
R11366 VDD.n6294 VDD.n6293 0.00119118
R11367 VDD.n6293 VDD.n487 0.00119118
R11368 VDD.n6314 VDD.n484 0.00119118
R11369 VDD.n6324 VDD.n484 0.00119118
R11370 VDD.n6319 VDD.n473 0.00119118
R11371 VDD.n6348 VDD.n473 0.00119118
R11372 VDD.n6354 VDD.n6353 0.00119118
R11373 VDD.n6354 VDD.n469 0.00119118
R11374 VDD.n6375 VDD.n6374 0.00119118
R11375 VDD.n6375 VDD.n452 0.00119118
R11376 VDD.n6399 VDD.n6398 0.00119118
R11377 VDD.n6399 VDD.n439 0.00119118
R11378 VDD.n6409 VDD.n435 0.00119118
R11379 VDD.n6414 VDD.n435 0.00119118
R11380 VDD.n6429 VDD.n424 0.00119118
R11381 VDD.n6435 VDD.n424 0.00119118
R11382 VDD.n6451 VDD.n6450 0.00119118
R11383 VDD.n6452 VDD.n6451 0.00119118
R11384 VDD.n6457 VDD.n401 0.00119118
R11385 VDD.n6474 VDD.n401 0.00119118
R11386 VDD.n6479 VDD.n390 0.00119118
R11387 VDD.n6494 VDD.n390 0.00119118
R11388 VDD.n6499 VDD.n368 0.00119118
R11389 VDD.n6513 VDD.n368 0.00119118
R11390 VDD.n6520 VDD.n6519 0.00119118
R11391 VDD.n6519 VDD.n353 0.00119118
R11392 VDD.n6540 VDD.n350 0.00119118
R11393 VDD.n6550 VDD.n350 0.00119118
R11394 VDD.n6545 VDD.n339 0.00119118
R11395 VDD.n6574 VDD.n339 0.00119118
R11396 VDD.n6580 VDD.n6579 0.00119118
R11397 VDD.n6580 VDD.n335 0.00119118
R11398 VDD.n6601 VDD.n6600 0.00119118
R11399 VDD.n6601 VDD.n318 0.00119118
R11400 VDD.n6625 VDD.n6624 0.00119118
R11401 VDD.n6625 VDD.n305 0.00119118
R11402 VDD.n6635 VDD.n301 0.00119118
R11403 VDD.n6640 VDD.n301 0.00119118
R11404 VDD.n6655 VDD.n290 0.00119118
R11405 VDD.n6661 VDD.n290 0.00119118
R11406 VDD.n6677 VDD.n6676 0.00119118
R11407 VDD.n6678 VDD.n6677 0.00119118
R11408 VDD.n6683 VDD.n267 0.00119118
R11409 VDD.n6700 VDD.n267 0.00119118
R11410 VDD.n6705 VDD.n256 0.00119118
R11411 VDD.n6720 VDD.n256 0.00119118
R11412 VDD.n6725 VDD.n234 0.00119118
R11413 VDD.n6739 VDD.n234 0.00119118
R11414 VDD.n6746 VDD.n6745 0.00119118
R11415 VDD.n6745 VDD.n219 0.00119118
R11416 VDD.n6766 VDD.n216 0.00119118
R11417 VDD.n6776 VDD.n216 0.00119118
R11418 VDD.n6771 VDD.n205 0.00119118
R11419 VDD.n6800 VDD.n205 0.00119118
R11420 VDD.n6806 VDD.n6805 0.00119118
R11421 VDD.n6806 VDD.n201 0.00119118
R11422 VDD.n6827 VDD.n6826 0.00119118
R11423 VDD.n6827 VDD.n184 0.00119118
R11424 VDD.n6851 VDD.n6850 0.00119118
R11425 VDD.n6851 VDD.n171 0.00119118
R11426 VDD.n6861 VDD.n167 0.00119118
R11427 VDD.n6866 VDD.n167 0.00119118
R11428 VDD.n6881 VDD.n156 0.00119118
R11429 VDD.n6887 VDD.n156 0.00119118
R11430 VDD.n6903 VDD.n6902 0.00119118
R11431 VDD.n6904 VDD.n6903 0.00119118
R11432 VDD.n6909 VDD.n133 0.00119118
R11433 VDD.n6926 VDD.n133 0.00119118
R11434 VDD.n6931 VDD.n122 0.00119118
R11435 VDD.n6946 VDD.n122 0.00119118
R11436 VDD.n6951 VDD.n100 0.00119118
R11437 VDD.n6965 VDD.n100 0.00119118
R11438 VDD.n6972 VDD.n6971 0.00119118
R11439 VDD.n6971 VDD.n85 0.00119118
R11440 VDD.n6992 VDD.n82 0.00119118
R11441 VDD.n7002 VDD.n82 0.00119118
R11442 VDD.n6997 VDD.n71 0.00119118
R11443 VDD.n7026 VDD.n71 0.00119118
R11444 VDD.n7032 VDD.n7031 0.00119118
R11445 VDD.n7032 VDD.n67 0.00119118
R11446 VDD.n7053 VDD.n7052 0.00119118
R11447 VDD.n7053 VDD.n49 0.00119118
R11448 VDD.n7057 VDD.n7056 0.00119118
R11449 VDD.n7057 VDD.n40 0.00119118
R11450 VDD.n7080 VDD.n38 0.00119118
R11451 VDD.n7090 VDD.n38 0.00119118
R11452 VDD.n7096 VDD.n7095 0.00119118
R11453 VDD.n7096 VDD.n33 0.00119118
R11454 VDD.n7206 VDD.n7100 0.00119118
R11455 VDD.n7206 VDD.n7205 0.00119118
R11456 VDD.n7134 VDD.n7128 0.00119118
R11457 VDD.n7135 VDD.n7134 0.00119118
R11458 VDD.n7186 VDD.n7185 0.00119118
R11459 VDD.n7185 VDD.n7126 0.00119118
R11460 VDD.n7179 VDD.n7146 0.00119118
R11461 VDD.n7158 VDD.n7146 0.00119118
R11462 VDD.n2742 VDD.n2737 0.00119118
R11463 VDD.n4331 VDD.n2742 0.00119118
R11464 VDD.n4326 VDD.n2747 0.00119118
R11465 VDD.n2750 VDD.n2747 0.00119118
R11466 VDD.n2801 VDD.n2786 0.00119118
R11467 VDD.n2802 VDD.n2801 0.00119118
R11468 VDD.n4306 VDD.n2784 0.00119118
R11469 VDD.n2807 VDD.n2784 0.00119118
R11470 VDD.n2870 VDD.n2808 0.00119118
R11471 VDD.n2871 VDD.n2870 0.00119118
R11472 VDD.n2885 VDD.n2884 0.00119118
R11473 VDD.n2886 VDD.n2885 0.00119118
R11474 VDD.n2893 VDD.n2892 0.00119118
R11475 VDD.n2892 VDD.n2862 0.00119118
R11476 VDD.n2859 VDD.n2857 0.00119118
R11477 VDD.n4265 VDD.n2859 0.00119118
R11478 VDD.n4260 VDD.n2905 0.00119118
R11479 VDD.n2939 VDD.n2905 0.00119118
R11480 VDD.n2934 VDD.n2932 0.00119118
R11481 VDD.n4244 VDD.n2934 0.00119118
R11482 VDD.n4239 VDD.n2948 0.00119118
R11483 VDD.n2980 VDD.n2948 0.00119118
R11484 VDD.n4224 VDD.n4223 0.00119118
R11485 VDD.n4223 VDD.n2977 0.00119118
R11486 VDD.n4215 VDD.n2990 0.00119118
R11487 VDD.n2992 VDD.n2990 0.00119118
R11488 VDD.n3043 VDD.n3028 0.00119118
R11489 VDD.n3044 VDD.n3043 0.00119118
R11490 VDD.n4195 VDD.n3026 0.00119118
R11491 VDD.n3049 VDD.n3026 0.00119118
R11492 VDD.n3096 VDD.n3050 0.00119118
R11493 VDD.n3097 VDD.n3096 0.00119118
R11494 VDD.n3112 VDD.n3092 0.00119118
R11495 VDD.n3113 VDD.n3112 0.00119118
R11496 VDD.n4168 VDD.n3090 0.00119118
R11497 VDD.n3118 VDD.n3090 0.00119118
R11498 VDD.n4162 VDD.n3119 0.00119118
R11499 VDD.n3162 VDD.n3119 0.00119118
R11500 VDD.n3157 VDD.n3155 0.00119118
R11501 VDD.n4146 VDD.n3157 0.00119118
R11502 VDD.n4141 VDD.n3171 0.00119118
R11503 VDD.n3205 VDD.n3171 0.00119118
R11504 VDD.n3200 VDD.n3198 0.00119118
R11505 VDD.n4125 VDD.n3200 0.00119118
R11506 VDD.n4120 VDD.n3214 0.00119118
R11507 VDD.n3246 VDD.n3214 0.00119118
R11508 VDD.n4105 VDD.n4104 0.00119118
R11509 VDD.n4104 VDD.n3243 0.00119118
R11510 VDD.n4096 VDD.n3256 0.00119118
R11511 VDD.n3258 VDD.n3256 0.00119118
R11512 VDD.n3309 VDD.n3294 0.00119118
R11513 VDD.n3310 VDD.n3309 0.00119118
R11514 VDD.n4076 VDD.n3292 0.00119118
R11515 VDD.n3315 VDD.n3292 0.00119118
R11516 VDD.n3362 VDD.n3316 0.00119118
R11517 VDD.n3363 VDD.n3362 0.00119118
R11518 VDD.n3378 VDD.n3358 0.00119118
R11519 VDD.n3379 VDD.n3378 0.00119118
R11520 VDD.n4049 VDD.n3356 0.00119118
R11521 VDD.n3384 VDD.n3356 0.00119118
R11522 VDD.n4043 VDD.n3385 0.00119118
R11523 VDD.n3428 VDD.n3385 0.00119118
R11524 VDD.n3423 VDD.n3421 0.00119118
R11525 VDD.n4027 VDD.n3423 0.00119118
R11526 VDD.n4022 VDD.n3437 0.00119118
R11527 VDD.n3471 VDD.n3437 0.00119118
R11528 VDD.n3466 VDD.n3464 0.00119118
R11529 VDD.n4006 VDD.n3466 0.00119118
R11530 VDD.n4001 VDD.n3480 0.00119118
R11531 VDD.n3512 VDD.n3480 0.00119118
R11532 VDD.n3986 VDD.n3985 0.00119118
R11533 VDD.n3985 VDD.n3509 0.00119118
R11534 VDD.n3977 VDD.n3522 0.00119118
R11535 VDD.n3524 VDD.n3522 0.00119118
R11536 VDD.n3575 VDD.n3560 0.00119118
R11537 VDD.n3576 VDD.n3575 0.00119118
R11538 VDD.n3957 VDD.n3558 0.00119118
R11539 VDD.n3581 VDD.n3558 0.00119118
R11540 VDD.n3628 VDD.n3582 0.00119118
R11541 VDD.n3629 VDD.n3628 0.00119118
R11542 VDD.n3644 VDD.n3624 0.00119118
R11543 VDD.n3645 VDD.n3644 0.00119118
R11544 VDD.n3930 VDD.n3622 0.00119118
R11545 VDD.n3650 VDD.n3622 0.00119118
R11546 VDD.n3924 VDD.n3651 0.00119118
R11547 VDD.n3694 VDD.n3651 0.00119118
R11548 VDD.n3689 VDD.n3687 0.00119118
R11549 VDD.n3908 VDD.n3689 0.00119118
R11550 VDD.n3903 VDD.n3703 0.00119118
R11551 VDD.n3737 VDD.n3703 0.00119118
R11552 VDD.n3732 VDD.n3730 0.00119118
R11553 VDD.n3887 VDD.n3732 0.00119118
R11554 VDD.n3882 VDD.n3746 0.00119118
R11555 VDD.n3778 VDD.n3746 0.00119118
R11556 VDD.n3867 VDD.n3866 0.00119118
R11557 VDD.n3866 VDD.n3775 0.00119118
R11558 VDD.n4386 VDD.n2433 0.00119118
R11559 VDD.n2438 VDD.n2433 0.00119118
R11560 VDD.n2659 VDD.n2439 0.00119118
R11561 VDD.n2660 VDD.n2659 0.00119118
R11562 VDD.n2675 VDD.n2655 0.00119118
R11563 VDD.n2676 VDD.n2675 0.00119118
R11564 VDD.n4359 VDD.n2653 0.00119118
R11565 VDD.n2681 VDD.n2653 0.00119118
R11566 VDD.n2720 VDD.n2682 0.00119118
R11567 VDD.n2720 VDD.n2718 0.00119118
R11568 VDD.n2733 VDD.n2716 0.00119118
R11569 VDD.n4338 VDD.n2716 0.00119118
R11570 VDD.n1411 VDD.n1375 0.00119118
R11571 VDD.n1412 VDD.n1411 0.00119118
R11572 VDD.n1427 VDD.n1408 0.00119118
R11573 VDD.n1428 VDD.n1427 0.00119118
R11574 VDD.n4857 VDD.n1406 0.00119118
R11575 VDD.n1433 VDD.n1406 0.00119118
R11576 VDD.n1480 VDD.n1434 0.00119118
R11577 VDD.n1481 VDD.n1480 0.00119118
R11578 VDD.n1496 VDD.n1476 0.00119118
R11579 VDD.n1497 VDD.n1496 0.00119118
R11580 VDD.n4830 VDD.n1474 0.00119118
R11581 VDD.n1502 VDD.n1474 0.00119118
R11582 VDD.n4824 VDD.n1503 0.00119118
R11583 VDD.n1544 VDD.n1503 0.00119118
R11584 VDD.n4809 VDD.n4808 0.00119118
R11585 VDD.n4808 VDD.n1541 0.00119118
R11586 VDD.n4802 VDD.n1553 0.00119118
R11587 VDD.n1586 VDD.n1553 0.00119118
R11588 VDD.n4787 VDD.n4786 0.00119118
R11589 VDD.n4786 VDD.n1583 0.00119118
R11590 VDD.n4780 VDD.n1595 0.00119118
R11591 VDD.n1628 VDD.n1595 0.00119118
R11592 VDD.n4765 VDD.n4764 0.00119118
R11593 VDD.n4764 VDD.n1625 0.00119118
R11594 VDD.n4756 VDD.n1638 0.00119118
R11595 VDD.n1641 VDD.n1638 0.00119118
R11596 VDD.n1691 VDD.n1676 0.00119118
R11597 VDD.n1692 VDD.n1691 0.00119118
R11598 VDD.n4736 VDD.n1674 0.00119118
R11599 VDD.n1697 VDD.n1674 0.00119118
R11600 VDD.n1744 VDD.n1698 0.00119118
R11601 VDD.n1745 VDD.n1744 0.00119118
R11602 VDD.n1760 VDD.n1740 0.00119118
R11603 VDD.n1761 VDD.n1760 0.00119118
R11604 VDD.n4709 VDD.n1738 0.00119118
R11605 VDD.n1766 VDD.n1738 0.00119118
R11606 VDD.n4703 VDD.n1767 0.00119118
R11607 VDD.n1808 VDD.n1767 0.00119118
R11608 VDD.n4688 VDD.n4687 0.00119118
R11609 VDD.n4687 VDD.n1805 0.00119118
R11610 VDD.n4681 VDD.n1817 0.00119118
R11611 VDD.n1850 VDD.n1817 0.00119118
R11612 VDD.n4666 VDD.n4665 0.00119118
R11613 VDD.n4665 VDD.n1847 0.00119118
R11614 VDD.n4659 VDD.n1859 0.00119118
R11615 VDD.n1892 VDD.n1859 0.00119118
R11616 VDD.n4644 VDD.n4643 0.00119118
R11617 VDD.n4643 VDD.n1889 0.00119118
R11618 VDD.n4635 VDD.n1902 0.00119118
R11619 VDD.n1905 VDD.n1902 0.00119118
R11620 VDD.n1955 VDD.n1940 0.00119118
R11621 VDD.n1956 VDD.n1955 0.00119118
R11622 VDD.n4615 VDD.n1938 0.00119118
R11623 VDD.n1961 VDD.n1938 0.00119118
R11624 VDD.n2008 VDD.n1962 0.00119118
R11625 VDD.n2009 VDD.n2008 0.00119118
R11626 VDD.n2024 VDD.n2004 0.00119118
R11627 VDD.n2025 VDD.n2024 0.00119118
R11628 VDD.n4588 VDD.n2002 0.00119118
R11629 VDD.n2030 VDD.n2002 0.00119118
R11630 VDD.n4582 VDD.n2031 0.00119118
R11631 VDD.n2072 VDD.n2031 0.00119118
R11632 VDD.n4567 VDD.n4566 0.00119118
R11633 VDD.n4566 VDD.n2069 0.00119118
R11634 VDD.n4560 VDD.n2081 0.00119118
R11635 VDD.n2114 VDD.n2081 0.00119118
R11636 VDD.n4545 VDD.n4544 0.00119118
R11637 VDD.n4544 VDD.n2111 0.00119118
R11638 VDD.n4538 VDD.n2123 0.00119118
R11639 VDD.n2156 VDD.n2123 0.00119118
R11640 VDD.n4523 VDD.n4522 0.00119118
R11641 VDD.n4522 VDD.n2153 0.00119118
R11642 VDD.n4514 VDD.n2166 0.00119118
R11643 VDD.n2169 VDD.n2166 0.00119118
R11644 VDD.n2219 VDD.n2204 0.00119118
R11645 VDD.n2220 VDD.n2219 0.00119118
R11646 VDD.n4494 VDD.n2202 0.00119118
R11647 VDD.n2225 VDD.n2202 0.00119118
R11648 VDD.n2272 VDD.n2226 0.00119118
R11649 VDD.n2273 VDD.n2272 0.00119118
R11650 VDD.n2288 VDD.n2268 0.00119118
R11651 VDD.n2289 VDD.n2288 0.00119118
R11652 VDD.n4467 VDD.n2266 0.00119118
R11653 VDD.n2294 VDD.n2266 0.00119118
R11654 VDD.n4461 VDD.n2295 0.00119118
R11655 VDD.n2336 VDD.n2295 0.00119118
R11656 VDD.n4446 VDD.n4445 0.00119118
R11657 VDD.n4445 VDD.n2333 0.00119118
R11658 VDD.n4439 VDD.n2345 0.00119118
R11659 VDD.n2378 VDD.n2345 0.00119118
R11660 VDD.n4424 VDD.n4423 0.00119118
R11661 VDD.n4423 VDD.n2375 0.00119118
R11662 VDD.n4417 VDD.n2387 0.00119118
R11663 VDD.n2420 VDD.n2387 0.00119118
R11664 VDD.n4402 VDD.n4401 0.00119118
R11665 VDD.n4401 VDD.n2417 0.00119118
R11666 VDD.n1283 VDD.n1264 0.00119118
R11667 VDD.n1284 VDD.n1283 0.00119118
R11668 VDD.n1300 VDD.n1260 0.00119118
R11669 VDD.n1301 VDD.n1300 0.00119118
R11670 VDD.n4909 VDD.n1258 0.00119118
R11671 VDD.n1306 VDD.n1258 0.00119118
R11672 VDD.n1353 VDD.n1307 0.00119118
R11673 VDD.n1354 VDD.n1353 0.00119118
R11674 VDD.n1369 VDD.n1349 0.00119118
R11675 VDD.n1370 VDD.n1369 0.00119118
R11676 VDD.n4882 VDD.n1347 0.00119118
R11677 VDD.n4878 VDD.n1347 0.00119118
R11678 VDD.n593 VDD.n591 0.0011215
R11679 VDD.n3837 VDD.n3835 0.0011215
R11680 VDD.n2513 VDD.n2511 0.0011215
R11681 VDD.n1223 VDD.n1221 0.0011215
R11682 VDD.n2611 VDD.n2460 0.00111039
R11683 VDD.n4947 VDD.n4939 0.00111039
R11684 VDD.n6111 VDD.n6110 0.00101648
R11685 VDD.n6181 VDD 0.000994737
R11686 VDD VDD.n436 0.000994737
R11687 VDD VDD.n302 0.000994737
R11688 VDD VDD.n168 0.000994737
R11689 VDD.n5020 VDD 0.000994737
R11690 VDD VDD.n5235 0.000994737
R11691 VDD VDD.n5463 0.000994737
R11692 VDD VDD.n5691 0.000994737
R11693 VDD VDD.n4877 0.000989583
R11694 VDD.n4758 VDD 0.000989583
R11695 VDD.n4637 VDD 0.000989583
R11696 VDD.n4516 VDD 0.000989583
R11697 VDD VDD.n4336 0.000989583
R11698 VDD.n4217 VDD 0.000989583
R11699 VDD.n4098 VDD 0.000989583
R11700 VDD.n3979 VDD 0.000989583
R11701 VDD.n1280 VDD 0.000982051
R11702 VDD.n2436 VDD 0.000982051
R11703 VDD.n2608 VDD.n2460 0.000837321
R11704 VDD.n4939 VDD.n1230 0.000837321
R11705 VDD.n7236 VDD.n7235 0.000837321
R11706 VDD.n6185 VDD.n6184 0.000747368
R11707 VDD.n6205 VDD.n6204 0.000747368
R11708 VDD.n550 VDD.n548 0.000747368
R11709 VDD.n6230 VDD.n534 0.000747368
R11710 VDD.n6252 VDD.n523 0.000747368
R11711 VDD.n6272 VDD.n501 0.000747368
R11712 VDD.n6292 VDD.n6291 0.000747368
R11713 VDD.n6323 VDD.n6317 0.000747368
R11714 VDD.n6349 VDD.n472 0.000747368
R11715 VDD.n6356 VDD.n6355 0.000747368
R11716 VDD.n6377 VDD.n6376 0.000747368
R11717 VDD.n6401 VDD.n6400 0.000747368
R11718 VDD.n6411 VDD.n6410 0.000747368
R11719 VDD.n6431 VDD.n6430 0.000747368
R11720 VDD.n416 VDD.n414 0.000747368
R11721 VDD.n6456 VDD.n400 0.000747368
R11722 VDD.n6478 VDD.n389 0.000747368
R11723 VDD.n6498 VDD.n367 0.000747368
R11724 VDD.n6518 VDD.n6517 0.000747368
R11725 VDD.n6549 VDD.n6543 0.000747368
R11726 VDD.n6575 VDD.n338 0.000747368
R11727 VDD.n6582 VDD.n6581 0.000747368
R11728 VDD.n6603 VDD.n6602 0.000747368
R11729 VDD.n6627 VDD.n6626 0.000747368
R11730 VDD.n6637 VDD.n6636 0.000747368
R11731 VDD.n6657 VDD.n6656 0.000747368
R11732 VDD.n282 VDD.n280 0.000747368
R11733 VDD.n6682 VDD.n266 0.000747368
R11734 VDD.n6704 VDD.n255 0.000747368
R11735 VDD.n6724 VDD.n233 0.000747368
R11736 VDD.n6744 VDD.n6743 0.000747368
R11737 VDD.n6775 VDD.n6769 0.000747368
R11738 VDD.n6801 VDD.n204 0.000747368
R11739 VDD.n6808 VDD.n6807 0.000747368
R11740 VDD.n6829 VDD.n6828 0.000747368
R11741 VDD.n6853 VDD.n6852 0.000747368
R11742 VDD.n6863 VDD.n6862 0.000747368
R11743 VDD.n6883 VDD.n6882 0.000747368
R11744 VDD.n148 VDD.n146 0.000747368
R11745 VDD.n6908 VDD.n132 0.000747368
R11746 VDD.n6930 VDD.n121 0.000747368
R11747 VDD.n6950 VDD.n99 0.000747368
R11748 VDD.n6970 VDD.n6969 0.000747368
R11749 VDD.n7001 VDD.n6995 0.000747368
R11750 VDD.n7027 VDD.n70 0.000747368
R11751 VDD.n7034 VDD.n7033 0.000747368
R11752 VDD.n7055 VDD.n7054 0.000747368
R11753 VDD.n7058 VDD.n39 0.000747368
R11754 VDD.n5021 VDD.n1195 0.000747368
R11755 VDD.n5032 VDD.n1184 0.000747368
R11756 VDD.n5055 VDD.n5053 0.000747368
R11757 VDD.n1171 VDD.n1169 0.000747368
R11758 VDD.n5091 VDD.n1155 0.000747368
R11759 VDD.n5115 VDD.n5114 0.000747368
R11760 VDD.n5142 VDD.n5136 0.000747368
R11761 VDD.n5168 VDD.n1110 0.000747368
R11762 VDD.n5175 VDD.n5174 0.000747368
R11763 VDD.n5196 VDD.n5195 0.000747368
R11764 VDD.n5224 VDD.n1076 0.000747368
R11765 VDD.n5231 VDD.n5230 0.000747368
R11766 VDD.n5234 VDD.n1060 0.000747368
R11767 VDD.n5260 VDD.n1049 0.000747368
R11768 VDD.n5283 VDD.n5281 0.000747368
R11769 VDD.n1036 VDD.n1034 0.000747368
R11770 VDD.n5319 VDD.n1020 0.000747368
R11771 VDD.n5343 VDD.n5342 0.000747368
R11772 VDD.n5370 VDD.n5364 0.000747368
R11773 VDD.n5396 VDD.n975 0.000747368
R11774 VDD.n5403 VDD.n5402 0.000747368
R11775 VDD.n5424 VDD.n5423 0.000747368
R11776 VDD.n5452 VDD.n941 0.000747368
R11777 VDD.n5459 VDD.n5458 0.000747368
R11778 VDD.n5462 VDD.n925 0.000747368
R11779 VDD.n5488 VDD.n914 0.000747368
R11780 VDD.n5511 VDD.n5509 0.000747368
R11781 VDD.n901 VDD.n899 0.000747368
R11782 VDD.n5547 VDD.n885 0.000747368
R11783 VDD.n5571 VDD.n5570 0.000747368
R11784 VDD.n5598 VDD.n5592 0.000747368
R11785 VDD.n5624 VDD.n840 0.000747368
R11786 VDD.n5631 VDD.n5630 0.000747368
R11787 VDD.n5652 VDD.n5651 0.000747368
R11788 VDD.n5680 VDD.n806 0.000747368
R11789 VDD.n5687 VDD.n5686 0.000747368
R11790 VDD.n5690 VDD.n790 0.000747368
R11791 VDD.n5716 VDD.n779 0.000747368
R11792 VDD.n5739 VDD.n5737 0.000747368
R11793 VDD.n766 VDD.n764 0.000747368
R11794 VDD.n5775 VDD.n750 0.000747368
R11795 VDD.n5798 VDD.n728 0.000747368
R11796 VDD.n5818 VDD.n720 0.000747368
R11797 VDD.n5840 VDD.n5839 0.000747368
R11798 VDD.n5871 VDD.n5865 0.000747368
R11799 VDD.n5897 VDD.n689 0.000747368
R11800 VDD.n5904 VDD.n5903 0.000747368
R11801 VDD.n5907 VDD.n668 0.000747368
R11802 VDD.n7078 VDD.n7077 0.000744792
R11803 VDD.n5928 VDD.n5927 0.000744792
R11804 VDD.n1410 VDD.n1374 0.000744792
R11805 VDD.n1426 VDD.n1425 0.000744792
R11806 VDD.n4856 VDD.n4855 0.000744792
R11807 VDD.n1479 VDD.n1478 0.000744792
R11808 VDD.n1495 VDD.n1494 0.000744792
R11809 VDD.n4829 VDD.n4828 0.000744792
R11810 VDD.n1543 VDD.n1542 0.000744792
R11811 VDD.n4807 VDD.n4806 0.000744792
R11812 VDD.n1585 VDD.n1584 0.000744792
R11813 VDD.n4785 VDD.n4784 0.000744792
R11814 VDD.n1627 VDD.n1626 0.000744792
R11815 VDD.n4763 VDD.n4762 0.000744792
R11816 VDD.n4757 VDD.n1637 0.000744792
R11817 VDD.n1690 VDD.n1689 0.000744792
R11818 VDD.n4735 VDD.n4734 0.000744792
R11819 VDD.n1743 VDD.n1742 0.000744792
R11820 VDD.n1759 VDD.n1758 0.000744792
R11821 VDD.n4708 VDD.n4707 0.000744792
R11822 VDD.n1807 VDD.n1806 0.000744792
R11823 VDD.n4686 VDD.n4685 0.000744792
R11824 VDD.n1849 VDD.n1848 0.000744792
R11825 VDD.n4664 VDD.n4663 0.000744792
R11826 VDD.n1891 VDD.n1890 0.000744792
R11827 VDD.n4642 VDD.n4641 0.000744792
R11828 VDD.n4636 VDD.n1901 0.000744792
R11829 VDD.n1954 VDD.n1953 0.000744792
R11830 VDD.n4614 VDD.n4613 0.000744792
R11831 VDD.n2007 VDD.n2006 0.000744792
R11832 VDD.n2023 VDD.n2022 0.000744792
R11833 VDD.n4587 VDD.n4586 0.000744792
R11834 VDD.n2071 VDD.n2070 0.000744792
R11835 VDD.n4565 VDD.n4564 0.000744792
R11836 VDD.n2113 VDD.n2112 0.000744792
R11837 VDD.n4543 VDD.n4542 0.000744792
R11838 VDD.n2155 VDD.n2154 0.000744792
R11839 VDD.n4521 VDD.n4520 0.000744792
R11840 VDD.n4515 VDD.n2165 0.000744792
R11841 VDD.n2218 VDD.n2217 0.000744792
R11842 VDD.n4493 VDD.n4492 0.000744792
R11843 VDD.n2271 VDD.n2270 0.000744792
R11844 VDD.n2287 VDD.n2286 0.000744792
R11845 VDD.n4466 VDD.n4465 0.000744792
R11846 VDD.n2335 VDD.n2334 0.000744792
R11847 VDD.n4444 VDD.n4443 0.000744792
R11848 VDD.n2377 VDD.n2376 0.000744792
R11849 VDD.n4422 VDD.n4421 0.000744792
R11850 VDD.n2419 VDD.n2418 0.000744792
R11851 VDD.n4400 VDD.n4399 0.000744792
R11852 VDD.n2744 VDD.n2736 0.000744792
R11853 VDD.n4327 VDD.n2745 0.000744792
R11854 VDD.n2800 VDD.n2799 0.000744792
R11855 VDD.n4305 VDD.n4304 0.000744792
R11856 VDD.n2869 VDD.n2868 0.000744792
R11857 VDD.n2875 VDD.n2865 0.000744792
R11858 VDD.n2891 VDD.n2890 0.000744792
R11859 VDD.n4264 VDD.n2903 0.000744792
R11860 VDD.n2938 VDD.n2937 0.000744792
R11861 VDD.n4243 VDD.n2946 0.000744792
R11862 VDD.n2979 VDD.n2978 0.000744792
R11863 VDD.n4222 VDD.n4221 0.000744792
R11864 VDD.n4216 VDD.n2989 0.000744792
R11865 VDD.n3042 VDD.n3041 0.000744792
R11866 VDD.n4194 VDD.n4193 0.000744792
R11867 VDD.n3095 VDD.n3094 0.000744792
R11868 VDD.n3111 VDD.n3110 0.000744792
R11869 VDD.n4167 VDD.n4166 0.000744792
R11870 VDD.n3161 VDD.n3160 0.000744792
R11871 VDD.n4145 VDD.n3169 0.000744792
R11872 VDD.n3204 VDD.n3203 0.000744792
R11873 VDD.n4124 VDD.n3212 0.000744792
R11874 VDD.n3245 VDD.n3244 0.000744792
R11875 VDD.n4103 VDD.n4102 0.000744792
R11876 VDD.n4097 VDD.n3255 0.000744792
R11877 VDD.n3308 VDD.n3307 0.000744792
R11878 VDD.n4075 VDD.n4074 0.000744792
R11879 VDD.n3361 VDD.n3360 0.000744792
R11880 VDD.n3377 VDD.n3376 0.000744792
R11881 VDD.n4048 VDD.n4047 0.000744792
R11882 VDD.n3427 VDD.n3426 0.000744792
R11883 VDD.n4026 VDD.n3435 0.000744792
R11884 VDD.n3470 VDD.n3469 0.000744792
R11885 VDD.n4005 VDD.n3478 0.000744792
R11886 VDD.n3511 VDD.n3510 0.000744792
R11887 VDD.n3984 VDD.n3983 0.000744792
R11888 VDD.n3978 VDD.n3521 0.000744792
R11889 VDD.n3574 VDD.n3573 0.000744792
R11890 VDD.n3956 VDD.n3955 0.000744792
R11891 VDD.n3627 VDD.n3626 0.000744792
R11892 VDD.n3643 VDD.n3642 0.000744792
R11893 VDD.n3929 VDD.n3928 0.000744792
R11894 VDD.n3693 VDD.n3692 0.000744792
R11895 VDD.n3907 VDD.n3701 0.000744792
R11896 VDD.n3736 VDD.n3735 0.000744792
R11897 VDD.n3886 VDD.n3744 0.000744792
R11898 VDD.n3777 VDD.n3776 0.000744792
R11899 VDD.n3865 VDD.n3864 0.000744792
R11900 VDD.n7091 VDD.n37 0.000743523
R11901 VDD.n7098 VDD.n7097 0.000743523
R11902 VDD.n7207 VDD.n7099 0.000743523
R11903 VDD.n7133 VDD.n7127 0.000743523
R11904 VDD.n7184 VDD.n7183 0.000743523
R11905 VDD.n7157 VDD.n7151 0.000743523
R11906 VDD.n5941 VDD.n666 0.000743523
R11907 VDD.n5948 VDD.n5947 0.000743523
R11908 VDD.n6057 VDD.n5949 0.000743523
R11909 VDD.n5983 VDD.n5977 0.000743523
R11910 VDD.n6034 VDD.n6033 0.000743523
R11911 VDD.n6007 VDD.n6001 0.000743523
R11912 VDD.n1282 VDD.n1281 0.000741026
R11913 VDD.n1299 VDD.n1298 0.000741026
R11914 VDD.n4908 VDD.n4907 0.000741026
R11915 VDD.n1352 VDD.n1351 0.000741026
R11916 VDD.n1368 VDD.n1367 0.000741026
R11917 VDD.n4881 VDD.n4880 0.000741026
R11918 VDD.n4385 VDD.n4384 0.000741026
R11919 VDD.n2658 VDD.n2657 0.000741026
R11920 VDD.n2674 VDD.n2673 0.000741026
R11921 VDD.n4358 VDD.n4357 0.000741026
R11922 VDD.n2721 VDD.n2719 0.000741026
R11923 VDD.n2735 VDD.n2734 0.000741026
R11924 VDD.n6168 VDD.n574 0.000709821
R11925 VDD.n579 VDD.n575 0.000709821
R11926 VDD.n6174 VDD.n570 0.000709821
R11927 VDD.n5007 VDD.n1204 0.000709821
R11928 VDD.n1209 VDD.n1205 0.000709821
R11929 VDD.n5013 VDD.n1200 0.000709821
R11930 VDD.n6111 VDD.n615 0.000693681
R11931 VDD.n2608 VDD.n2607 0.00061244
R11932 VDD.n4978 VDD.n1230 0.00061244
R11933 VDD.n7235 VDD.n7234 0.00061244
R11934 VDD.n6139 VDD.n574 0.000541964
R11935 VDD.n6167 VDD.n575 0.000541964
R11936 VDD.n580 VDD.n570 0.000541964
R11937 VDD.n4982 VDD.n1204 0.000541964
R11938 VDD.n5006 VDD.n1205 0.000541964
R11939 VDD.n1210 VDD.n1200 0.000541964
R11940 VSS VSS.n1325 2.45983e+06
R11941 VSS.n2362 VSS.n2361 553784
R11942 VSS.n2432 VSS.n2431 553379
R11943 VSS.n1324 VSS 22710.2
R11944 VSS.n259 VSS.n258 15644.4
R11945 VSS.n2167 VSS.n2166 15155.6
R11946 VSS.t55 VSS.n1258 1270.52
R11947 VSS.n2361 VSS.t53 1150.15
R11948 VSS.n2432 VSS.t58 1136.78
R11949 VSS.n1326 VSS 1043.16
R11950 VSS.n2341 VSS 1043.16
R11951 VSS.t39 VSS.n1316 1043.16
R11952 VSS.n1313 VSS.n1261 782.529
R11953 VSS.n2442 VSS 775.684
R11954 VSS.n1260 VSS 775.684
R11955 VSS.n700 VSS.t62 641.946
R11956 VSS.n1260 VSS.t55 641.946
R11957 VSS.n2505 VSS.n2504 626.532
R11958 VSS.n1377 VSS.n1376 626.532
R11959 VSS.n2234 VSS 601.824
R11960 VSS VSS.n1323 601.824
R11961 VSS.n1288 VSS.n1257 585
R11962 VSS.n1316 VSS.n1257 585
R11963 VSS.n1322 VSS.n1321 585
R11964 VSS.n1323 VSS.n1322 585
R11965 VSS.n1318 VSS.n1257 481.557
R11966 VSS.t33 VSS.n672 424.519
R11967 VSS.t82 VSS.n1228 424.519
R11968 VSS.n533 VSS.t12 360.841
R11969 VSS.t34 VSS.n2290 360.534
R11970 VSS.t21 VSS.n2430 360.534
R11971 VSS.n700 VSS 320.974
R11972 VSS.n2299 VSS 320.974
R11973 VSS.n1320 VSS.n1253 294.606
R11974 VSS.n259 VSS.t31 294.416
R11975 VSS.n702 VSS.n701 292.5
R11976 VSS.n701 VSS.n700 292.5
R11977 VSS.n2444 VSS.n2443 292.5
R11978 VSS.n2443 VSS.n2442 292.5
R11979 VSS.n2301 VSS.n2300 292.5
R11980 VSS.n2300 VSS.n2299 292.5
R11981 VSS.n1314 VSS.n1259 292.5
R11982 VSS.n1315 VSS.n1314 292.5
R11983 VSS.n1305 VSS.n1261 292.5
R11984 VSS.n1261 VSS.n1260 292.5
R11985 VSS.n1253 VSS.n1252 292.5
R11986 VSS.n1324 VSS.n1251 292.168
R11987 VSS.t20 VSS.t44 234.535
R11988 VSS.n688 VSS.n687 227.357
R11989 VSS.n2360 VSS.n2291 227.357
R11990 VSS.n2270 VSS.n2269 213.982
R11991 VSS.n1316 VSS.n1315 213.982
R11992 VSS.n2236 VSS.n2235 187.234
R11993 VSS.n1317 VSS.n1252 187.234
R11994 VSS.n1328 VSS.n1327 173.861
R11995 VSS.n2343 VSS.n2342 173.861
R11996 VSS.n1613 VSS.t79 153.446
R11997 VSS.n2086 VSS.t77 153.446
R11998 VSS.n397 VSS.t70 153.446
R11999 VSS.n1703 VSS.t36 153.446
R12000 VSS.n2007 VSS.t10 153.446
R12001 VSS.n1789 VSS.t2 153.446
R12002 VSS.n1760 VSS.t1 153.446
R12003 VSS.n465 VSS.t71 153.446
R12004 VSS.n2773 VSS.t32 153.446
R12005 VSS.n2737 VSS.t83 153.446
R12006 VSS.n75 VSS.t78 153.446
R12007 VSS.n999 VSS.t80 153.446
R12008 VSS.n187 VSS.t49 153.446
R12009 VSS.n871 VSS.t72 153.446
R12010 VSS.n903 VSS.t7 153.446
R12011 VSS.n2641 VSS.t81 153.446
R12012 VSS.n1328 VSS.t64 147.113
R12013 VSS.n2343 VSS.t5 147.113
R12014 VSS.n2236 VSS.t75 133.739
R12015 VSS.n2433 VSS.n2432 133.739
R12016 VSS.n2361 VSS.n2360 133.739
R12017 VSS.n1317 VSS.t39 133.739
R12018 VSS.t12 VSS.t66 114.87
R12019 VSS.t29 VSS.t73 114.87
R12020 VSS.n1569 VSS.t52 114.772
R12021 VSS.n629 VSS.t61 114.772
R12022 VSS.t46 VSS.t34 114.772
R12023 VSS.t19 VSS.t21 114.772
R12024 VSS.n2801 VSS.t57 114.772
R12025 VSS.n2577 VSS.t60 114.772
R12026 VSS.n423 VSS.t50 112.278
R12027 VSS.n1876 VSS.t51 112.278
R12028 VSS.n121 VSS.t37 112.278
R12029 VSS.n1008 VSS.t67 112.278
R12030 VSS.n2301 VSS.t54 107.195
R12031 VSS.n702 VSS.t63 107.195
R12032 VSS.n1305 VSS.t56 107.195
R12033 VSS.n2336 VSS.t6 107.195
R12034 VSS.n2444 VSS.t59 107.195
R12035 VSS.n2229 VSS.t76 107.195
R12036 VSS.n723 VSS.t65 107.195
R12037 VSS.n1254 VSS.t40 107.195
R12038 VSS.n2431 VSS.t20 103.544
R12039 VSS.t44 VSS.n2362 102.297
R12040 VSS.n689 VSS.n686 93.0283
R12041 VSS.n2359 VSS.n2292 93.0283
R12042 VSS.n2268 VSS.n2267 87.5561
R12043 VSS.n1314 VSS.n1257 87.5561
R12044 VSS.n1378 VSS.n1377 87.4012
R12045 VSS.n1230 VSS.n1229 87.4012
R12046 VSS.n2506 VSS.n2505 87.3268
R12047 VSS.n2375 VSS.n2374 87.3268
R12048 VSS.n1325 VSS.t23 82.4069
R12049 VSS.n766 VSS.t28 77.3934
R12050 VSS.n766 VSS.t27 77.3934
R12051 VSS.n512 VSS.t8 77.3934
R12052 VSS.n512 VSS.t11 77.3934
R12053 VSS.n335 VSS.t18 77.3934
R12054 VSS.n335 VSS.t17 77.3934
R12055 VSS.n2473 VSS.t45 77.3934
R12056 VSS.n2473 VSS.t47 77.3934
R12057 VSS.n2237 VSS.n2233 76.6116
R12058 VSS.n1318 VSS.n1253 76.6116
R12059 VSS.n1329 VSS.n727 71.1394
R12060 VSS.n2344 VSS.n2340 71.1394
R12061 VSS.t73 VSS.n1324 68.6725
R12062 VSS.n1377 VSS.t33 66.1753
R12063 VSS.n1229 VSS.t82 66.1753
R12064 VSS.n2505 VSS.t31 66.119
R12065 VSS.n2374 VSS.t69 66.119
R12066 VSS.t66 VSS.n532 58.6838
R12067 VSS.t38 VSS.n1568 57.3864
R12068 VSS.n2430 VSS.t41 57.3864
R12069 VSS.t30 VSS.n2800 57.3864
R12070 VSS.t68 VSS.n552 56.1389
R12071 VSS.t9 VSS.n2576 56.1389
R12072 VSS.n1327 VSS.n1326 53.4959
R12073 VSS.n2342 VSS.n2341 53.4959
R12074 VSS.n2169 VSS.n2168 51.1488
R12075 VSS.n261 VSS.n260 51.1488
R12076 VSS.n540 VSS.t0 47.4466
R12077 VSS.n728 VSS.t24 47.4466
R12078 VSS.n2280 VSS.t15 47.4062
R12079 VSS.n2389 VSS.t42 47.4062
R12080 VSS.n777 VSS.t74 43.7547
R12081 VSS.n2483 VSS.t35 43.7547
R12082 VSS.n522 VSS.t13 43.7547
R12083 VSS.n346 VSS.t22 43.7547
R12084 VSS.n540 VSS.t4 42.4523
R12085 VSS.n728 VSS.t25 42.4523
R12086 VSS.n2280 VSS.t14 42.4162
R12087 VSS.n1 VSS.t26 41.4448
R12088 VSS.n2504 VSS.t16 41.4448
R12089 VSS.n2458 VSS.t43 41.4448
R12090 VSS.n1376 VSS.t3 41.4448
R12091 VSS.n2235 VSS.n2234 40.1221
R12092 VSS.n1323 VSS.n1252 40.1221
R12093 VSS.n658 VSS.n657 38.7065
R12094 VSS.t52 VSS.t38 38.6736
R12095 VSS.t61 VSS.t68 38.6736
R12096 VSS.n629 VSS.n628 38.6736
R12097 VSS.n648 VSS.n647 38.6736
R12098 VSS.t57 VSS.t30 38.6736
R12099 VSS.t60 VSS.t9 38.6736
R12100 VSS.n1325 VSS.t29 37.4579
R12101 VSS.n669 VSS.n668 32.4636
R12102 VSS.n1306 VSS.n1262 23.9034
R12103 VSS.n1289 VSS.n1288 22.6545
R12104 VSS.n727 VSS.n726 21.8894
R12105 VSS.n2340 VSS.n2339 21.8894
R12106 VSS.n1355 VSS.t48 21.2264
R12107 VSS VSS.n1254 20.1079
R12108 VSS.n2229 VSS 20.1079
R12109 VSS.n1508 VSS.n1507 17.6406
R12110 VSS.n355 VSS.n354 17.6397
R12111 VSS.n2362 VSS.t46 17.4658
R12112 VSS.n2233 VSS.n2232 16.4172
R12113 VSS.n1322 VSS.n1253 16.4172
R12114 VSS.n2122 VSS.n2121 16.2182
R12115 VSS.n2111 VSS.n2110 16.2182
R12116 VSS.n2097 VSS.n2096 16.2182
R12117 VSS.n2431 VSS.t19 16.2182
R12118 VSS.n1126 VSS.n1125 16.2182
R12119 VSS.n2762 VSS.n2761 16.2182
R12120 VSS.n2748 VSS.n2747 16.2182
R12121 VSS.n2408 VSS 14.0497
R12122 VSS.n2433 VSS.n2270 13.3744
R12123 VSS.n1315 VSS.n1258 13.3744
R12124 VSS.n703 VSS.n702 13.1351
R12125 VSS.n2302 VSS.n2301 13.1351
R12126 VSS.n1306 VSS.n1305 13.1351
R12127 VSS.n1422 VSS.n1421 13.0195
R12128 VSS.n781 VSS 12.4783
R12129 VSS.n720 VSS.n719 9.3005
R12130 VSS.n718 VSS.n717 9.3005
R12131 VSS.n1330 VSS.n1329 9.3005
R12132 VSS.n1329 VSS.n1328 9.3005
R12133 VSS.n2246 VSS.n2245 9.3005
R12134 VSS.n2244 VSS.n2243 9.3005
R12135 VSS.n2436 VSS.n2434 9.3005
R12136 VSS.n2434 VSS.n2433 9.3005
R12137 VSS.n2238 VSS.n2237 9.3005
R12138 VSS.n2237 VSS.n2236 9.3005
R12139 VSS.n2345 VSS.n2344 9.3005
R12140 VSS.n2344 VSS.n2343 9.3005
R12141 VSS.n2352 VSS.n2351 9.3005
R12142 VSS.n2350 VSS.n2349 9.3005
R12143 VSS.n1290 VSS.n1289 9.3005
R12144 VSS.n1264 VSS.n1262 9.3005
R12145 VSS.n1313 VSS.n1312 9.3005
R12146 VSS.n1313 VSS.n1258 9.3005
R12147 VSS.n1319 VSS.n1256 9.3005
R12148 VSS.n1319 VSS.n1318 9.3005
R12149 VSS.n1318 VSS.n1317 9.3005
R12150 VSS.n1287 VSS.n1272 9.3005
R12151 VSS.n1286 VSS.n1285 9.3005
R12152 VSS.n1530 VSS.n1529 9.15497
R12153 VSS.n2211 VSS.n2210 9.15497
R12154 VSS.n656 VSS.n655 9.15497
R12155 VSS.n657 VSS.n656 9.15497
R12156 VSS.n671 VSS.n670 9.15497
R12157 VSS.n672 VSS.n671 9.15497
R12158 VSS.n530 VSS.n529 9.15497
R12159 VSS.n529 VSS.n528 9.15497
R12160 VSS.n542 VSS.n541 9.15497
R12161 VSS.n541 VSS.n540 9.15497
R12162 VSS.n535 VSS.n534 9.15497
R12163 VSS.n534 VSS.n533 9.15497
R12164 VSS.n1380 VSS.n1379 9.15497
R12165 VSS.n1379 VSS.n1378 9.15497
R12166 VSS.n627 VSS.n626 9.15497
R12167 VSS.n628 VSS.n627 9.15497
R12168 VSS.n646 VSS.n645 9.15497
R12169 VSS.n647 VSS.n646 9.15497
R12170 VSS.n1741 VSS.n1740 9.15497
R12171 VSS.n1740 VSS.n1739 9.15497
R12172 VSS.n1751 VSS.n1750 9.15497
R12173 VSS.n1750 VSS.n1749 9.15497
R12174 VSS.n1744 VSS.n1743 9.15497
R12175 VSS.n1743 VSS.n1742 9.15497
R12176 VSS.n1762 VSS.n1761 9.15497
R12177 VSS.n1761 VSS.n1760 9.15497
R12178 VSS.n1814 VSS.n1813 9.15497
R12179 VSS.n1813 VSS.n1812 9.15497
R12180 VSS.n1784 VSS.n1783 9.15497
R12181 VSS.n1783 VSS.n1782 9.15497
R12182 VSS.n1791 VSS.n1790 9.15497
R12183 VSS.n1790 VSS.n1789 9.15497
R12184 VSS.n1830 VSS.n1829 9.15497
R12185 VSS.n1829 VSS.n1828 9.15497
R12186 VSS.n1875 VSS.n1874 9.15497
R12187 VSS.n1874 VSS.n1873 9.15497
R12188 VSS.n1885 VSS.n1884 9.15497
R12189 VSS.n1884 VSS.n1883 9.15497
R12190 VSS.n1878 VSS.n1877 9.15497
R12191 VSS.n1877 VSS.n1876 9.15497
R12192 VSS.n1896 VSS.n1895 9.15497
R12193 VSS.n1895 VSS.n1894 9.15497
R12194 VSS.n1698 VSS.n1697 9.15497
R12195 VSS.n1697 VSS.n1696 9.15497
R12196 VSS.n1705 VSS.n1704 9.15497
R12197 VSS.n1704 VSS.n1703 9.15497
R12198 VSS.n1643 VSS.n1642 9.15497
R12199 VSS.n1642 VSS.n1641 9.15497
R12200 VSS.n1665 VSS.n1664 9.15497
R12201 VSS.n1664 VSS.n1663 9.15497
R12202 VSS.n2120 VSS.n2119 9.15497
R12203 VSS.n2121 VSS.n2120 9.15497
R12204 VSS.n2113 VSS.n2112 9.15497
R12205 VSS.n2112 VSS.n2111 9.15497
R12206 VSS.n2099 VSS.n2098 9.15497
R12207 VSS.n2098 VSS.n2097 9.15497
R12208 VSS.n1615 VSS.n1614 9.15497
R12209 VSS.n1614 VSS.n1613 9.15497
R12210 VSS.n1563 VSS.n1562 9.15497
R12211 VSS.n1562 VSS.n1561 9.15497
R12212 VSS.n1571 VSS.n1570 9.15497
R12213 VSS.n1570 VSS.n1569 9.15497
R12214 VSS.n2171 VSS.n2170 9.15497
R12215 VSS.n2170 VSS.n2169 9.15497
R12216 VSS.n2178 VSS.n2177 9.15497
R12217 VSS.n2177 VSS.n2176 9.15497
R12218 VSS.n1988 VSS.n1987 9.15497
R12219 VSS.n1987 VSS.n1986 9.15497
R12220 VSS.n1998 VSS.n1997 9.15497
R12221 VSS.n1997 VSS.n1996 9.15497
R12222 VSS.n1991 VSS.n1990 9.15497
R12223 VSS.n1990 VSS.n1989 9.15497
R12224 VSS.n2009 VSS.n2008 9.15497
R12225 VSS.n2008 VSS.n2007 9.15497
R12226 VSS.n1941 VSS.n1940 9.15497
R12227 VSS.n1940 VSS.n1939 9.15497
R12228 VSS.n1970 VSS.n1969 9.15497
R12229 VSS.n1969 VSS.n1968 9.15497
R12230 VSS.n1977 VSS.n1976 9.15497
R12231 VSS.n1976 VSS.n1975 9.15497
R12232 VSS.n425 VSS.n424 9.15497
R12233 VSS.n424 VSS.n423 9.15497
R12234 VSS.n378 VSS.n377 9.15497
R12235 VSS.n377 VSS.n376 9.15497
R12236 VSS.n388 VSS.n387 9.15497
R12237 VSS.n387 VSS.n386 9.15497
R12238 VSS.n381 VSS.n380 9.15497
R12239 VSS.n380 VSS.n379 9.15497
R12240 VSS.n399 VSS.n398 9.15497
R12241 VSS.n398 VSS.n397 9.15497
R12242 VSS.n2109 VSS.n2108 9.15497
R12243 VSS.n2110 VSS.n2109 9.15497
R12244 VSS.n2095 VSS.n2094 9.15497
R12245 VSS.n2096 VSS.n2095 9.15497
R12246 VSS.n2088 VSS.n2087 9.15497
R12247 VSS.n2087 VSS.n2086 9.15497
R12248 VSS.n2124 VSS.n2123 9.15497
R12249 VSS.n2123 VSS.n2122 9.15497
R12250 VSS.n1465 VSS.n1464 9.15497
R12251 VSS.n1464 VSS.n1463 9.15497
R12252 VSS.n460 VSS.n459 9.15497
R12253 VSS.n459 VSS.n458 9.15497
R12254 VSS.n467 VSS.n466 9.15497
R12255 VSS.n466 VSS.n465 9.15497
R12256 VSS.n442 VSS.n441 9.15497
R12257 VSS.n441 VSS.n440 9.15497
R12258 VSS.n650 VSS.n649 9.15497
R12259 VSS.n649 VSS.n648 9.15497
R12260 VSS.n660 VSS.n659 9.15497
R12261 VSS.n659 VSS.n658 9.15497
R12262 VSS.n667 VSS.n666 9.15497
R12263 VSS.n668 VSS.n667 9.15497
R12264 VSS.n631 VSS.n630 9.15497
R12265 VSS.n630 VSS.n629 9.15497
R12266 VSS.n2384 VSS.n2383 9.15497
R12267 VSS.n2383 VSS.n2382 9.15497
R12268 VSS.n2377 VSS.n2376 9.15497
R12269 VSS.n2376 VSS.n2375 9.15497
R12270 VSS.n2429 VSS.n2428 9.15497
R12271 VSS.n2430 VSS.n2429 9.15497
R12272 VSS.n2391 VSS.n2390 9.15497
R12273 VSS.n2390 VSS.n2389 9.15497
R12274 VSS.n2275 VSS.n2274 9.15497
R12275 VSS.n2274 VSS.n2273 9.15497
R12276 VSS.n2282 VSS.n2281 9.15497
R12277 VSS.n2281 VSS.n2280 9.15497
R12278 VSS.n2289 VSS.n2288 9.15497
R12279 VSS.n2290 VSS.n2289 9.15497
R12280 VSS.n2508 VSS.n2507 9.15497
R12281 VSS.n2507 VSS.n2506 9.15497
R12282 VSS.n2611 VSS.n2610 9.15497
R12283 VSS.n306 VSS.n305 9.15497
R12284 VSS.n1171 VSS.n1170 9.15497
R12285 VSS.n1170 VSS.n1169 9.15497
R12286 VSS.n1178 VSS.n1177 9.15497
R12287 VSS.n1177 VSS.n1176 9.15497
R12288 VSS.n168 VSS.n167 9.15497
R12289 VSS.n167 VSS.n166 9.15497
R12290 VSS.n178 VSS.n177 9.15497
R12291 VSS.n177 VSS.n176 9.15497
R12292 VSS.n171 VSS.n170 9.15497
R12293 VSS.n170 VSS.n169 9.15497
R12294 VSS.n189 VSS.n188 9.15497
R12295 VSS.n188 VSS.n187 9.15497
R12296 VSS.n136 VSS.n135 9.15497
R12297 VSS.n135 VSS.n134 9.15497
R12298 VSS.n155 VSS.n154 9.15497
R12299 VSS.n154 VSS.n153 9.15497
R12300 VSS.n162 VSS.n161 9.15497
R12301 VSS.n161 VSS.n160 9.15497
R12302 VSS.n123 VSS.n122 9.15497
R12303 VSS.n122 VSS.n121 9.15497
R12304 VSS.n56 VSS.n55 9.15497
R12305 VSS.n55 VSS.n54 9.15497
R12306 VSS.n66 VSS.n65 9.15497
R12307 VSS.n65 VSS.n64 9.15497
R12308 VSS.n59 VSS.n58 9.15497
R12309 VSS.n58 VSS.n57 9.15497
R12310 VSS.n77 VSS.n76 9.15497
R12311 VSS.n76 VSS.n75 9.15497
R12312 VSS.n2760 VSS.n2759 9.15497
R12313 VSS.n2761 VSS.n2760 9.15497
R12314 VSS.n2746 VSS.n2745 9.15497
R12315 VSS.n2747 VSS.n2746 9.15497
R12316 VSS.n2739 VSS.n2738 9.15497
R12317 VSS.n2738 VSS.n2737 9.15497
R12318 VSS.n1128 VSS.n1127 9.15497
R12319 VSS.n1127 VSS.n1126 9.15497
R12320 VSS.n2571 VSS.n2570 9.15497
R12321 VSS.n2570 VSS.n2569 9.15497
R12322 VSS.n2579 VSS.n2578 9.15497
R12323 VSS.n2578 VSS.n2577 9.15497
R12324 VSS.n2629 VSS.n2628 9.15497
R12325 VSS.n2628 VSS.n2627 9.15497
R12326 VSS.n2636 VSS.n2635 9.15497
R12327 VSS.n2635 VSS.n2634 9.15497
R12328 VSS.n2643 VSS.n2642 9.15497
R12329 VSS.n2642 VSS.n2641 9.15497
R12330 VSS.n235 VSS.n234 9.15497
R12331 VSS.n234 VSS.n233 9.15497
R12332 VSS.n1124 VSS.n45 9.15497
R12333 VSS.n1125 VSS.n1124 9.15497
R12334 VSS.n2764 VSS.n2763 9.15497
R12335 VSS.n2763 VSS.n2762 9.15497
R12336 VSS.n2750 VSS.n2749 9.15497
R12337 VSS.n2749 VSS.n2748 9.15497
R12338 VSS.n2775 VSS.n2774 9.15497
R12339 VSS.n2774 VSS.n2773 9.15497
R12340 VSS.n2795 VSS.n2794 9.15497
R12341 VSS.n2794 VSS.n2793 9.15497
R12342 VSS.n2803 VSS.n2802 9.15497
R12343 VSS.n2802 VSS.n2801 9.15497
R12344 VSS.n884 VSS.n883 9.15497
R12345 VSS.n883 VSS.n882 9.15497
R12346 VSS.n894 VSS.n893 9.15497
R12347 VSS.n893 VSS.n892 9.15497
R12348 VSS.n887 VSS.n886 9.15497
R12349 VSS.n886 VSS.n885 9.15497
R12350 VSS.n905 VSS.n904 9.15497
R12351 VSS.n904 VSS.n903 9.15497
R12352 VSS.n837 VSS.n836 9.15497
R12353 VSS.n836 VSS.n835 9.15497
R12354 VSS.n866 VSS.n865 9.15497
R12355 VSS.n865 VSS.n864 9.15497
R12356 VSS.n873 VSS.n872 9.15497
R12357 VSS.n872 VSS.n871 9.15497
R12358 VSS.n807 VSS.n806 9.15497
R12359 VSS.n806 VSS.n805 9.15497
R12360 VSS.n1007 VSS.n1006 9.15497
R12361 VSS.n1006 VSS.n1005 9.15497
R12362 VSS.n1017 VSS.n1016 9.15497
R12363 VSS.n1016 VSS.n1015 9.15497
R12364 VSS.n1010 VSS.n1009 9.15497
R12365 VSS.n1009 VSS.n1008 9.15497
R12366 VSS.n1028 VSS.n1027 9.15497
R12367 VSS.n1027 VSS.n1026 9.15497
R12368 VSS.n1092 VSS.n1091 9.15497
R12369 VSS.n1091 VSS.n1090 9.15497
R12370 VSS.n994 VSS.n993 9.15497
R12371 VSS.n993 VSS.n992 9.15497
R12372 VSS.n1001 VSS.n1000 9.15497
R12373 VSS.n1000 VSS.n999 9.15497
R12374 VSS.n1108 VSS.n1107 9.15497
R12375 VSS.n1107 VSS.n1106 9.15497
R12376 VSS.n263 VSS.n262 9.15497
R12377 VSS.n262 VSS.n261 9.15497
R12378 VSS.n271 VSS.n270 9.15497
R12379 VSS.n270 VSS.n269 9.15497
R12380 VSS.n1209 VSS.n1208 9.15497
R12381 VSS.n1208 VSS.n1207 9.15497
R12382 VSS.n1227 VSS.n1226 9.15497
R12383 VSS.n1228 VSS.n1227 9.15497
R12384 VSS.n730 VSS.n729 9.15497
R12385 VSS.n729 VSS.n728 9.15497
R12386 VSS.n1239 VSS.n1238 9.15497
R12387 VSS.n1238 VSS.n1237 9.15497
R12388 VSS.n1232 VSS.n1231 9.15497
R12389 VSS.n1231 VSS.n1230 9.15497
R12390 VSS.n1250 VSS.n1249 9.15497
R12391 VSS.n1251 VSS.n1250 9.15497
R12392 VSS.n2835 VSS.n2834 9.15497
R12393 VSS.n2834 VSS.n2833 9.15497
R12394 VSS.n2849 VSS.n2848 9.15497
R12395 VSS.n2848 VSS.n2847 9.15497
R12396 VSS.n690 VSS.n689 9.01392
R12397 VSS.n2359 VSS.n2358 9.01392
R12398 VSS.n2360 VSS.n2359 9.01392
R12399 VSS.n689 VSS.n688 9.01392
R12400 VSS.n2610 VSS.n2609 8.48574
R12401 VSS.n305 VSS.n304 8.48574
R12402 VSS.n2445 VSS.n2444 8.11658
R12403 VSS.n1305 VSS.n1304 8.11658
R12404 VSS.n702 VSS 7.93155
R12405 VSS.n2301 VSS 7.93155
R12406 VSS.n2230 VSS.n2229 7.90638
R12407 VSS.n1321 VSS.n1254 7.90638
R12408 VSS.n724 VSS.n723 7.52991
R12409 VSS.n2337 VSS.n2336 7.52991
R12410 VSS.n1228 VSS.n789 7.49199
R12411 VSS.n672 VSS.n669 6.24341
R12412 VSS.n260 VSS.n259 6.2381
R12413 VSS.n2434 VSS.n2268 5.47272
R12414 VSS.n1314 VSS.n1313 5.47272
R12415 VSS.n1296 VSS.n1269 5.18083
R12416 VSS.n2168 VSS.n2167 4.99058
R12417 VSS.n1274 VSS 4.7265
R12418 VSS.n704 VSS.n703 4.6505
R12419 VSS.n2441 VSS.n2440 4.6505
R12420 VSS.n2303 VSS.n2302 4.6505
R12421 VSS.n1307 VSS.n1306 4.6505
R12422 VSS VSS.n698 4.5005
R12423 VSS.n1332 VSS.n1331 4.5005
R12424 VSS.n2241 VSS.n2240 4.5005
R12425 VSS.n2347 VSS.n2346 4.5005
R12426 VSS VSS.n2298 4.5005
R12427 VSS.n1277 VSS.n1276 4.5005
R12428 VSS.n1284 VSS.n1283 4.5005
R12429 VSS.n1284 VSS.n1255 4.5005
R12430 VSS.n1303 VSS.n1302 4.5005
R12431 VSS.n1292 VSS.n1291 4.5005
R12432 VSS.n1311 VSS.n1310 4.5005
R12433 VSS.n1309 VSS.n1308 4.5005
R12434 VSS.n2240 VSS.n2239 3.76521
R12435 VSS.n1331 VSS.n722 3.76521
R12436 VSS.n2346 VSS.n2335 3.76521
R12437 VSS.n1286 VSS.n1255 3.76521
R12438 VSS.n533 VSS.n531 3.74624
R12439 VSS.n1278 VSS.n1277 3.45606
R12440 VSS.n2436 VSS.n2435 3.45447
R12441 VSS.n690 VSS.n685 3.45447
R12442 VSS.n2358 VSS.n2357 3.45447
R12443 VSS.n1312 VSS.n1262 3.45447
R12444 VSS.n1283 VSS.n1282 3.42401
R12445 VSS.n1302 VSS.n1301 3.42259
R12446 VSS.n937 VSS 3.42087
R12447 VSS.n1293 VSS.n1292 3.42064
R12448 VSS.n1309 VSS.n1266 3.41895
R12449 VSS.n1281 VSS.n1280 3.4105
R12450 VSS.n1297 VSS.n1296 3.4105
R12451 VSS.n1300 VSS.n1299 3.4105
R12452 VSS.n1279 VSS.n1271 3.4105
R12453 VSS.n1295 VSS.n1294 3.4105
R12454 VSS.n2864 VSS.n2863 3.4105
R12455 VSS.n2238 VSS.n2231 3.38874
R12456 VSS.n725 VSS.n724 3.38874
R12457 VSS.n2338 VSS.n2337 3.38874
R12458 VSS.n1320 VSS.n1319 3.38874
R12459 VSS.n2266 VSS.n2265 3.25129
R12460 VSS.n691 VSS.n684 3.25129
R12461 VSS.n2356 VSS.n2293 3.25129
R12462 VSS.n1288 VSS.n1259 3.25129
R12463 VSS.n1244 VSS.n730 3.03311
R12464 VSS.n265 VSS.n263 3.03311
R12465 VSS.n2630 VSS.n2629 3.03311
R12466 VSS.n1093 VSS.n1092 3.03311
R12467 VSS.n1022 VSS.n1007 3.03311
R12468 VSS.n838 VSS.n837 3.03311
R12469 VSS.n899 VSS.n884 3.03311
R12470 VSS.n2836 VSS.n2835 3.03311
R12471 VSS.n2769 VSS.n45 3.03311
R12472 VSS.n1210 VSS.n1209 3.03311
R12473 VSS.n2759 VSS.n2758 3.03311
R12474 VSS.n71 VSS.n56 3.03311
R12475 VSS.n137 VSS.n136 3.03311
R12476 VSS.n183 VSS.n168 3.03311
R12477 VSS.n2276 VSS.n2275 3.03311
R12478 VSS.n2428 VSS.n2427 3.03311
R12479 VSS.n1466 VSS.n1465 3.03311
R12480 VSS.n2108 VSS.n2107 3.03311
R12481 VSS.n393 VSS.n378 3.03311
R12482 VSS.n1942 VSS.n1941 3.03311
R12483 VSS.n2003 VSS.n1988 3.03311
R12484 VSS.n1644 VSS.n1643 3.03311
R12485 VSS.n1890 VSS.n1875 3.03311
R12486 VSS.n1815 VSS.n1814 3.03311
R12487 VSS.n1756 VSS.n1741 3.03311
R12488 VSS.n2212 VSS.n2211 3.03311
R12489 VSS.n2119 VSS.n2118 3.03311
R12490 VSS.n1509 VSS.n1508 3.03311
R12491 VSS.n1531 VSS.n1530 3.03311
R12492 VSS.n356 VSS.n355 3.03311
R12493 VSS.n547 VSS.n530 3.03311
R12494 VSS.n692 VSS.n691 3.03311
R12495 VSS.n543 VSS.n542 3.03311
R12496 VSS.n536 VSS.n535 3.03311
R12497 VSS.n1381 VSS.n1380 3.03311
R12498 VSS.n626 VSS.n625 3.03311
R12499 VSS.n645 VSS.n644 3.03311
R12500 VSS.n1752 VSS.n1751 3.03311
R12501 VSS.n1745 VSS.n1744 3.03311
R12502 VSS.n1763 VSS.n1762 3.03311
R12503 VSS.n1785 VSS.n1784 3.03311
R12504 VSS.n1792 VSS.n1791 3.03311
R12505 VSS.n1831 VSS.n1830 3.03311
R12506 VSS.n1886 VSS.n1885 3.03311
R12507 VSS.n1879 VSS.n1878 3.03311
R12508 VSS.n1897 VSS.n1896 3.03311
R12509 VSS.n1699 VSS.n1698 3.03311
R12510 VSS.n1706 VSS.n1705 3.03311
R12511 VSS.n1666 VSS.n1665 3.03311
R12512 VSS.n2114 VSS.n2113 3.03311
R12513 VSS.n2100 VSS.n2099 3.03311
R12514 VSS.n1616 VSS.n1615 3.03311
R12515 VSS.n1564 VSS.n1563 3.03311
R12516 VSS.n1572 VSS.n1571 3.03311
R12517 VSS.n2172 VSS.n2171 3.03311
R12518 VSS.n2179 VSS.n2178 3.03311
R12519 VSS.n1999 VSS.n1998 3.03311
R12520 VSS.n1992 VSS.n1991 3.03311
R12521 VSS.n2010 VSS.n2009 3.03311
R12522 VSS.n1971 VSS.n1970 3.03311
R12523 VSS.n1978 VSS.n1977 3.03311
R12524 VSS.n426 VSS.n425 3.03311
R12525 VSS.n389 VSS.n388 3.03311
R12526 VSS.n382 VSS.n381 3.03311
R12527 VSS.n400 VSS.n399 3.03311
R12528 VSS.n2094 VSS.n2093 3.03311
R12529 VSS.n2089 VSS.n2088 3.03311
R12530 VSS.n2125 VSS.n2124 3.03311
R12531 VSS.n461 VSS.n460 3.03311
R12532 VSS.n468 VSS.n467 3.03311
R12533 VSS.n443 VSS.n442 3.03311
R12534 VSS.n651 VSS.n650 3.03311
R12535 VSS.n661 VSS.n660 3.03311
R12536 VSS.n666 VSS.n665 3.03311
R12537 VSS.n632 VSS.n631 3.03311
R12538 VSS.n2385 VSS.n2384 3.03311
R12539 VSS.n2378 VSS.n2377 3.03311
R12540 VSS.n2392 VSS.n2391 3.03311
R12541 VSS.n2283 VSS.n2282 3.03311
R12542 VSS.n2288 VSS.n2287 3.03311
R12543 VSS.n2509 VSS.n2508 3.03311
R12544 VSS.n2356 VSS.n2355 3.03311
R12545 VSS.n2613 VSS.n2611 3.03311
R12546 VSS.n2559 VSS.n2558 3.03311
R12547 VSS.n307 VSS.n306 3.03311
R12548 VSS.n325 VSS.n324 3.03311
R12549 VSS.n1172 VSS.n1171 3.03311
R12550 VSS.n1179 VSS.n1178 3.03311
R12551 VSS.n179 VSS.n178 3.03311
R12552 VSS.n172 VSS.n171 3.03311
R12553 VSS.n190 VSS.n189 3.03311
R12554 VSS.n156 VSS.n155 3.03311
R12555 VSS.n163 VSS.n162 3.03311
R12556 VSS.n124 VSS.n123 3.03311
R12557 VSS.n67 VSS.n66 3.03311
R12558 VSS.n60 VSS.n59 3.03311
R12559 VSS.n78 VSS.n77 3.03311
R12560 VSS.n2745 VSS.n2744 3.03311
R12561 VSS.n2740 VSS.n2739 3.03311
R12562 VSS.n1129 VSS.n1128 3.03311
R12563 VSS.n2572 VSS.n2571 3.03311
R12564 VSS.n2580 VSS.n2579 3.03311
R12565 VSS.n2637 VSS.n2636 3.03311
R12566 VSS.n2644 VSS.n2643 3.03311
R12567 VSS.n236 VSS.n235 3.03311
R12568 VSS.n2765 VSS.n2764 3.03311
R12569 VSS.n2751 VSS.n2750 3.03311
R12570 VSS.n2776 VSS.n2775 3.03311
R12571 VSS.n2796 VSS.n2795 3.03311
R12572 VSS.n2804 VSS.n2803 3.03311
R12573 VSS.n895 VSS.n894 3.03311
R12574 VSS.n888 VSS.n887 3.03311
R12575 VSS.n906 VSS.n905 3.03311
R12576 VSS.n867 VSS.n866 3.03311
R12577 VSS.n874 VSS.n873 3.03311
R12578 VSS.n808 VSS.n807 3.03311
R12579 VSS.n1018 VSS.n1017 3.03311
R12580 VSS.n1011 VSS.n1010 3.03311
R12581 VSS.n1029 VSS.n1028 3.03311
R12582 VSS.n995 VSS.n994 3.03311
R12583 VSS.n1002 VSS.n1001 3.03311
R12584 VSS.n1109 VSS.n1108 3.03311
R12585 VSS.n272 VSS.n271 3.03311
R12586 VSS.n1226 VSS.n1225 3.03311
R12587 VSS.n1240 VSS.n1239 3.03311
R12588 VSS.n1233 VSS.n1232 3.03311
R12589 VSS.n1249 VSS.n1248 3.03311
R12590 VSS.n2850 VSS.n2849 3.03311
R12591 VSS.n2231 VSS.n2230 3.01226
R12592 VSS.n1330 VSS.n725 3.01226
R12593 VSS.n2345 VSS.n2338 3.01226
R12594 VSS.n1321 VSS.n1320 3.01226
R12595 VSS.n2437 VSS.n2436 2.28739
R12596 VSS.n1312 VSS.n1311 2.28739
R12597 VSS.n2502 VSS.n252 2.24031
R12598 VSS.n1374 VSS.n673 2.24031
R12599 VSS VSS.n2501 1.94963
R12600 VSS VSS.n1373 1.94963
R12601 VSS.n1331 VSS.n1330 1.50638
R12602 VSS.n2346 VSS.n2345 1.50638
R12603 VSS.n1287 VSS.n1286 1.50638
R12604 VSS.n1535 VSS.n1532 1.35607
R12605 VSS.n1337 VSS.n1336 1.35607
R12606 VSS.n715 VSS.n714 1.35607
R12607 VSS.n2227 VSS.n2226 1.35607
R12608 VSS.n2333 VSS.n2332 1.35607
R12609 VSS.n2354 VSS.n2309 1.35607
R12610 VSS.n2615 VSS.n2614 1.35607
R12611 VSS.n312 VSS.n308 1.35607
R12612 VSS.n328 VSS.n326 1.35607
R12613 VSS.n241 VSS.n238 1.35607
R12614 VSS.n814 VSS.n810 1.35607
R12615 VSS.n844 VSS.n840 1.35607
R12616 VSS.n1114 VSS.n1111 1.35607
R12617 VSS.n1097 VSS.n1094 1.35607
R12618 VSS.n2855 VSS.n2852 1.35607
R12619 VSS.n2838 VSS.n2837 1.35607
R12620 VSS.n1224 VSS.n1223 1.35607
R12621 VSS.n1214 VSS.n1211 1.35607
R12622 VSS.n130 VSS.n126 1.35607
R12623 VSS.n143 VSS.n139 1.35607
R12624 VSS.n1143 VSS.n1132 1.35607
R12625 VSS.n2426 VSS.n2425 1.35607
R12626 VSS.n432 VSS.n428 1.35607
R12627 VSS.n1948 VSS.n1944 1.35607
R12628 VSS.n2139 VSS.n2128 1.35607
R12629 VSS.n1837 VSS.n1833 1.35607
R12630 VSS.n1821 VSS.n1817 1.35607
R12631 VSS.n1670 VSS.n1667 1.35607
R12632 VSS.n1647 VSS.n1646 1.35607
R12633 VSS.n361 VSS.n358 1.35607
R12634 VSS.n2214 VSS.n2213 1.35607
R12635 VSS.n1514 VSS.n1511 1.35607
R12636 VSS.n707 VSS.n706 1.35607
R12637 VSS.n448 VSS.n445 1.35607
R12638 VSS.n1470 VSS.n1467 1.35607
R12639 VSS.n2264 VSS.n2263 1.35607
R12640 VSS.n2297 VSS.n2295 1.35607
R12641 VSS.n2561 VSS.n2560 1.35607
R12642 VSS.n1275 VSS.n1273 1.35607
R12643 VSS.n1265 VSS.n1263 1.35607
R12644 VSS.n779 VSS.n778 1.13981
R12645 VSS.n524 VSS.n523 1.13981
R12646 VSS.n348 VSS.n347 1.13981
R12647 VSS.n2485 VSS.n2484 1.13981
R12648 VSS.n1795 VSS.n1778 1.13845
R12649 VSS.n1294 VSS.n1270 1.13717
R12650 VSS.n2783 VSS.n16 1.13708
R12651 VSS.n294 VSS.n293 1.13696
R12652 VSS.n1370 VSS.n1369 1.13462
R12653 VSS.n2466 VSS.n2465 1.13462
R12654 VSS.n2866 VSS.n2865 1.13462
R12655 VSS.n785 VSS.n784 1.13388
R12656 VSS.n1157 VSS.n1156 1.13388
R12657 VSS.n1418 VSS.n1417 1.13388
R12658 VSS.n2412 VSS.n2411 1.13388
R12659 VSS.n2240 VSS.n2238 1.12991
R12660 VSS.n1319 VSS.n1255 1.12991
R12661 VSS.n1289 VSS.n1287 1.12991
R12662 VSS.n2449 VSS.n2447 1.04225
R12663 VSS.n1268 VSS.n1267 1.04225
R12664 VSS.n6 VSS.n5 1.04173
R12665 VSS.n2461 VSS.n2460 1.04145
R12666 VSS.n1233 VSS.n788 1.04008
R12667 VSS.n2645 VSS.n2644 1.04008
R12668 VSS.n1003 VSS.n1002 1.04008
R12669 VSS.n875 VSS.n874 1.04008
R12670 VSS.n1180 VSS.n1179 1.04008
R12671 VSS.n2740 VSS.n2736 1.04008
R12672 VSS.n164 VSS.n163 1.04008
R12673 VSS.n2378 VSS.n2373 1.04008
R12674 VSS.n469 VSS.n468 1.04008
R12675 VSS.n2089 VSS.n2085 1.04008
R12676 VSS.n1979 VSS.n1978 1.04008
R12677 VSS.n1707 VSS.n1706 1.04008
R12678 VSS.n1793 VSS.n1792 1.04008
R12679 VSS.n2180 VSS.n2179 1.03997
R12680 VSS.n2805 VSS.n2804 1.03985
R12681 VSS.n2581 VSS.n2580 1.03985
R12682 VSS.n273 VSS.n272 1.03985
R12683 VSS.n1030 VSS.n1029 1.03985
R12684 VSS.n907 VSS.n906 1.03985
R12685 VSS.n2777 VSS.n2776 1.03985
R12686 VSS.n79 VSS.n78 1.03985
R12687 VSS.n191 VSS.n190 1.03985
R12688 VSS.n2510 VSS.n2509 1.03985
R12689 VSS.n2011 VSS.n2010 1.03985
R12690 VSS.n401 VSS.n400 1.03985
R12691 VSS.n1764 VSS.n1763 1.03985
R12692 VSS.n1898 VSS.n1897 1.03985
R12693 VSS.n1617 VSS.n1616 1.03985
R12694 VSS.n1573 VSS.n1572 1.03985
R12695 VSS.n1382 VSS.n1381 1.03985
R12696 VSS.n625 VSS.n621 1.03985
R12697 VSS.n632 VSS.n551 1.03985
R12698 VSS.n2487 VSS.n2470 1.03084
R12699 VSS.n697 VSS.n696 0.878546
R12700 VSS.n1340 VSS.n1339 0.878359
R12701 VSS.n1280 VSS.n1278 0.871022
R12702 VSS.n1301 VSS.n1300 0.870834
R12703 VSS.n771 VSS.n769 0.853
R12704 VSS.n2864 VSS.n8 0.853
R12705 VSS.n277 VSS.n276 0.853
R12706 VSS.n242 VSS.n241 0.853
R12707 VSS.n967 VSS.n814 0.853
R12708 VSS.n967 VSS.n966 0.853
R12709 VSS.n938 VSS.n927 0.853
R12710 VSS.n943 VSS.n924 0.853
R12711 VSS.n948 VSS.n918 0.853
R12712 VSS.n953 VSS.n912 0.853
R12713 VSS.n877 VSS.n876 0.853
R12714 VSS.n856 VSS.n855 0.853
R12715 VSS.n845 VSS.n844 0.853
R12716 VSS.n954 VSS.n953 0.853
R12717 VSS.n2859 VSS.n2858 0.853
R12718 VSS.n2783 VSS.n2782 0.853
R12719 VSS.n2807 VSS.n2806 0.853
R12720 VSS.n2821 VSS.n2818 0.853
R12721 VSS.n2841 VSS.n2838 0.853
R12722 VSS.n2858 VSS.n2855 0.853
R12723 VSS.n2842 VSS.n2841 0.853
R12724 VSS.n2822 VSS.n2821 0.853
R12725 VSS.n2808 VSS.n2807 0.853
R12726 VSS.n1223 VSS.n1222 0.853
R12727 VSS.n1222 VSS.n1221 0.853
R12728 VSS.n1183 VSS.n1181 0.853
R12729 VSS.n1197 VSS.n1194 0.853
R12730 VSS.n1217 VSS.n1214 0.853
R12731 VSS.n1218 VSS.n1217 0.853
R12732 VSS.n1198 VSS.n1197 0.853
R12733 VSS.n1184 VSS.n1183 0.853
R12734 VSS.n2729 VSS.n84 0.853
R12735 VSS.n2729 VSS.n2728 0.853
R12736 VSS.n2710 VSS.n143 0.853
R12737 VSS.n2715 VSS.n130 0.853
R12738 VSS.n115 VSS.n114 0.853
R12739 VSS.n107 VSS.n106 0.853
R12740 VSS.n96 VSS.n95 0.853
R12741 VSS.n2716 VSS.n2715 0.853
R12742 VSS.n2735 VSS.n2734 0.853
R12743 VSS.n1155 VSS.n1143 0.853
R12744 VSS.n33 VSS.n31 0.853
R12745 VSS.n37 VSS.n28 0.853
R12746 VSS.n41 VSS.n22 0.853
R12747 VSS.n972 VSS.n802 0.853
R12748 VSS.n1051 VSS.n1046 0.853
R12749 VSS.n1056 VSS.n1041 0.853
R12750 VSS.n1061 VSS.n1035 0.853
R12751 VSS.n1066 VSS.n1004 0.853
R12752 VSS.n1080 VSS.n1077 0.853
R12753 VSS.n1100 VSS.n1097 0.853
R12754 VSS.n1117 VSS.n1114 0.853
R12755 VSS.n1118 VSS.n1117 0.853
R12756 VSS.n1101 VSS.n1100 0.853
R12757 VSS.n1081 VSS.n1080 0.853
R12758 VSS.n1067 VSS.n1066 0.853
R12759 VSS.n973 VSS.n972 0.853
R12760 VSS.n2695 VSS.n196 0.853
R12761 VSS.n2700 VSS.n165 0.853
R12762 VSS.n2705 VSS.n149 0.853
R12763 VSS.n2695 VSS.n2694 0.853
R12764 VSS.n213 VSS.n211 0.853
R12765 VSS.n218 VSS.n208 0.853
R12766 VSS.n223 VSS.n202 0.853
R12767 VSS.n2681 VSS.n242 0.853
R12768 VSS.n2649 VSS.n2646 0.853
R12769 VSS.n2663 VSS.n2660 0.853
R12770 VSS.n2677 VSS.n2674 0.853
R12771 VSS.n2678 VSS.n2677 0.853
R12772 VSS.n2664 VSS.n2663 0.853
R12773 VSS.n2650 VSS.n2649 0.853
R12774 VSS.n294 VSS.n286 0.853
R12775 VSS.n330 VSS.n328 0.853
R12776 VSS.n315 VSS.n312 0.853
R12777 VSS.n316 VSS.n315 0.853
R12778 VSS.n331 VSS.n330 0.853
R12779 VSS.n2500 VSS.n2499 0.853
R12780 VSS.n2501 VSS.n2500 0.853
R12781 VSS.n2372 VSS.n2371 0.853
R12782 VSS.n2219 VSS.n364 0.853
R12783 VSS.n2183 VSS.n2182 0.853
R12784 VSS.n2197 VSS.n2196 0.853
R12785 VSS.n2216 VSS.n2215 0.853
R12786 VSS.n364 VSS.n361 0.853
R12787 VSS.n2196 VSS.n2195 0.853
R12788 VSS.n2182 VSS.n2181 0.853
R12789 VSS.n2215 VSS.n2214 0.853
R12790 VSS.n1536 VSS.n1535 0.853
R12791 VSS.n1373 VSS.n1372 0.853
R12792 VSS.n714 VSS.n713 0.853
R12793 VSS.n1338 VSS.n1337 0.853
R12794 VSS.n708 VSS.n707 0.853
R12795 VSS.n449 VSS.n448 0.853
R12796 VSS.n1477 VSS.n449 0.853
R12797 VSS.n492 VSS.n490 0.853
R12798 VSS.n497 VSS.n487 0.853
R12799 VSS.n502 VSS.n481 0.853
R12800 VSS.n1434 VSS.n475 0.853
R12801 VSS.n1439 VSS.n470 0.853
R12802 VSS.n1453 VSS.n1450 0.853
R12803 VSS.n1473 VSS.n1470 0.853
R12804 VSS.n1474 VSS.n1473 0.853
R12805 VSS.n1454 VSS.n1453 0.853
R12806 VSS.n1440 VSS.n1439 0.853
R12807 VSS.n1434 VSS.n1433 0.853
R12808 VSS.n516 VSS.n515 0.853
R12809 VSS.n1416 VSS.n1402 0.853
R12810 VSS.n620 VSS.n619 0.853
R12811 VSS.n619 VSS.n618 0.853
R12812 VSS.n1723 VSS.n1722 0.853
R12813 VSS.n605 VSS.n604 0.853
R12814 VSS.n604 VSS.n603 0.853
R12815 VSS.n1734 VSS.n1733 0.853
R12816 VSS.n1770 VSS.n1769 0.853
R12817 VSS.n1805 VSS.n1804 0.853
R12818 VSS.n1795 VSS.n1794 0.853
R12819 VSS.n2033 VSS.n2031 0.853
R12820 VSS.n2037 VSS.n2028 0.853
R12821 VSS.n2042 VSS.n2022 0.853
R12822 VSS.n2047 VSS.n2016 0.853
R12823 VSS.n1981 VSS.n1980 0.853
R12824 VSS.n1960 VSS.n1959 0.853
R12825 VSS.n1949 VSS.n1948 0.853
R12826 VSS.n2061 VSS.n432 0.853
R12827 VSS.n2066 VSS.n421 0.853
R12828 VSS.n2061 VSS.n2060 0.853
R12829 VSS.n2048 VSS.n2047 0.853
R12830 VSS.n2084 VSS.n2083 0.853
R12831 VSS.n2154 VSS.n2139 0.853
R12832 VSS.n2155 VSS.n2154 0.853
R12833 VSS.n2070 VSS.n418 0.853
R12834 VSS.n2074 VSS.n412 0.853
R12835 VSS.n2078 VSS.n406 0.853
R12836 VSS.n1650 VSS.n1647 0.853
R12837 VSS.n1822 VSS.n1821 0.853
R12838 VSS.n1838 VSS.n1837 0.853
R12839 VSS.n1857 VSS.n1856 0.853
R12840 VSS.n1846 VSS.n1845 0.853
R12841 VSS.n1868 VSS.n1867 0.853
R12842 VSS.n1905 VSS.n1904 0.853
R12843 VSS.n1904 VSS.n1903 0.853
R12844 VSS.n1686 VSS.n1685 0.853
R12845 VSS.n1685 VSS.n1684 0.853
R12846 VSS.n1709 VSS.n1690 0.853
R12847 VSS.n1709 VSS.n1708 0.853
R12848 VSS.n1671 VSS.n1670 0.853
R12849 VSS.n1672 VSS.n1671 0.853
R12850 VSS.n1651 VSS.n1650 0.853
R12851 VSS.n1537 VSS.n1536 0.853
R12852 VSS.n1517 VSS.n1514 0.853
R12853 VSS.n1595 VSS.n1594 0.853
R12854 VSS.n1584 VSS.n1583 0.853
R12855 VSS.n1606 VSS.n1605 0.853
R12856 VSS.n1624 VSS.n1623 0.853
R12857 VSS.n1623 VSS.n1622 0.853
R12858 VSS.n1551 VSS.n1550 0.853
R12859 VSS.n1550 VSS.n1549 0.853
R12860 VSS.n1575 VSS.n1555 0.853
R12861 VSS.n1575 VSS.n1574 0.853
R12862 VSS.n1518 VSS.n1517 0.853
R12863 VSS.n340 VSS.n338 0.853
R12864 VSS.n2425 VSS.n2424 0.853
R12865 VSS.n2464 VSS.n2462 0.853
R12866 VSS.n2263 VSS.n2262 0.853
R12867 VSS.n2320 VSS.n2309 0.853
R12868 VSS.n2332 VSS.n2330 0.853
R12869 VSS.n2477 VSS.n2476 0.853
R12870 VSS.n2547 VSS.n2530 0.853
R12871 VSS.n2548 VSS.n2547 0.853
R12872 VSS.n2563 VSS.n2562 0.853
R12873 VSS.n2617 VSS.n2616 0.853
R12874 VSS.n2616 VSS.n2615 0.853
R12875 VSS.n2562 VSS.n2561 0.853
R12876 VSS.n2595 VSS.n2594 0.853
R12877 VSS.n2585 VSS.n2584 0.853
R12878 VSS.n1274 VSS.n1273 0.853
R12879 VSS.n1294 VSS.n1265 0.853
R12880 VSS.n787 VSS.n786 0.853
R12881 VSS.n2254 VSS.n2253 0.699777
R12882 VSS.n2329 VSS.n2328 0.699777
R12883 VSS.n2452 VSS.n2451 0.699516
R12884 VSS.n2314 VSS.n2313 0.699516
R12885 VSS.n773 VSS.n772 0.698382
R12886 VSS.n518 VSS.n517 0.698382
R12887 VSS.n342 VSS.n341 0.698382
R12888 VSS.n2479 VSS.n2478 0.698382
R12889 VSS.n778 VSS.n777 0.684595
R12890 VSS.n2484 VSS.n2483 0.684595
R12891 VSS.n523 VSS.n522 0.684595
R12892 VSS.n347 VSS.n346 0.684595
R12893 VSS.n1298 VSS.n1268 0.682713
R12894 VSS.n2450 VSS.n2449 0.682713
R12895 VSS.n1295 VSS 0.5645
R12896 VSS.n1296 VSS.n1295 0.4705
R12897 VSS.n343 VSS.n342 0.354051
R12898 VSS.n2480 VSS.n2479 0.354051
R12899 VSS.n519 VSS.n518 0.352782
R12900 VSS.n774 VSS.n773 0.352759
R12901 VSS.n2609 VSS.n2608 0.33661
R12902 VSS.n1507 VSS.n1506 0.336142
R12903 VSS.n1358 VSS.n1354 0.261125
R12904 VSS.n2470 VSS.n350 0.253125
R12905 VSS.n2470 VSS.n2469 0.249386
R12906 VSS.n1064 VSS.n1063 0.212
R12907 VSS.n970 VSS.n969 0.212
R12908 VSS.n880 VSS.n879 0.212
R12909 VSS.n2786 VSS.n2785 0.212
R12910 VSS.n2732 VSS.n2731 0.212
R12911 VSS.n118 VSS.n117 0.212
R12912 VSS.n2698 VSS.n2697 0.212
R12913 VSS.n2081 VSS.n2080 0.212
R12914 VSS.n2064 VSS.n2063 0.212
R12915 VSS.n1984 VSS.n1983 0.212
R12916 VSS.n1712 VSS.n1711 0.212
R12917 VSS.n1841 VSS.n1840 0.212
R12918 VSS.n1773 VSS.n1772 0.212
R12919 VSS.n1578 VSS.n1577 0.212
R12920 VSS.n1437 VSS.n1436 0.212
R12921 VSS.n2436 VSS.n2266 0.203675
R12922 VSS.n691 VSS.n690 0.203675
R12923 VSS.n2358 VSS.n2356 0.203675
R12924 VSS.n1312 VSS.n1259 0.203675
R12925 VSS.n2487 VSS.n2486 0.183261
R12926 VSS.n2325 VSS 0.180125
R12927 VSS.n2453 VSS 0.170375
R12928 VSS.n781 VSS.n780 0.127459
R12929 VSS.n2868 VSS 0.125741
R12930 VSS.n2408 VSS.n350 0.119277
R12931 VSS.n2497 VSS 0.112761
R12932 VSS.n2503 VSS 0.104812
R12933 VSS.n1375 VSS 0.104812
R12934 VSS.n1635 VSS 0.103332
R12935 VSS.n350 VSS.n349 0.101141
R12936 VSS.n1120 VSS 0.0994474
R12937 VSS.n2304 VSS.n2303 0.0929479
R12938 VSS.n1160 VSS 0.0903012
R12939 VSS.n1120 VSS 0.0897843
R12940 VSS.n2247 VSS.n2246 0.0825312
R12941 VSS.n1291 VSS.n1290 0.0825312
R12942 VSS.n1422 VSS 0.0801269
R12943 VSS.n2453 VSS 0.0763587
R12944 VSS.n827 VSS 0.0753227
R12945 VSS.n1335 VSS.n1334 0.0734167
R12946 VSS.n2311 VSS.n2310 0.0734167
R12947 VSS.n435 VSS 0.0724848
R12948 VSS.n696 VSS.n675 0.0714273
R12949 VSS VSS.n2868 0.0707673
R12950 VSS.n1421 VSS.n526 0.0702516
R12951 VSS.n1345 VSS.n1344 0.0698595
R12952 VSS.n1246 VSS.n1245 0.0685147
R12953 VSS.n1242 VSS.n1241 0.0685147
R12954 VSS.n1235 VSS.n1234 0.0685147
R12955 VSS.n2575 VSS.n2574 0.0685147
R12956 VSS.n268 VSS.n267 0.0685147
R12957 VSS.n2633 VSS.n2632 0.0685147
R12958 VSS.n2640 VSS.n2639 0.0685147
R12959 VSS.n991 VSS.n990 0.0685147
R12960 VSS.n998 VSS.n997 0.0685147
R12961 VSS.n1025 VSS.n1024 0.0685147
R12962 VSS.n1021 VSS.n1020 0.0685147
R12963 VSS.n1014 VSS.n1013 0.0685147
R12964 VSS.n870 VSS.n869 0.0685147
R12965 VSS.n902 VSS.n901 0.0685147
R12966 VSS.n898 VSS.n897 0.0685147
R12967 VSS.n891 VSS.n890 0.0685147
R12968 VSS.n2792 VSS.n2791 0.0685147
R12969 VSS.n2799 VSS.n2798 0.0685147
R12970 VSS.n2772 VSS.n2771 0.0685147
R12971 VSS.n2768 VSS.n2767 0.0685147
R12972 VSS.n2754 VSS.n2753 0.0685147
R12973 VSS.n1168 VSS.n1167 0.0685147
R12974 VSS.n1175 VSS.n1174 0.0685147
R12975 VSS.n1131 VSS.n1130 0.0685147
R12976 VSS.n2756 VSS.n2755 0.0685147
R12977 VSS.n2742 VSS.n2741 0.0685147
R12978 VSS.n74 VSS.n73 0.0685147
R12979 VSS.n70 VSS.n69 0.0685147
R12980 VSS.n63 VSS.n62 0.0685147
R12981 VSS.n159 VSS.n158 0.0685147
R12982 VSS.n186 VSS.n185 0.0685147
R12983 VSS.n182 VSS.n181 0.0685147
R12984 VSS.n175 VSS.n174 0.0685147
R12985 VSS.n2271 VSS.n251 0.0685147
R12986 VSS.n2278 VSS.n2277 0.0685147
R12987 VSS.n2285 VSS.n2284 0.0685147
R12988 VSS.n2394 VSS.n2393 0.0685147
R12989 VSS.n2387 VSS.n2386 0.0685147
R12990 VSS.n2380 VSS.n2379 0.0685147
R12991 VSS.n457 VSS.n456 0.0685147
R12992 VSS.n464 VSS.n463 0.0685147
R12993 VSS.n2006 VSS.n2005 0.0685147
R12994 VSS.n2002 VSS.n2001 0.0685147
R12995 VSS.n1995 VSS.n1994 0.0685147
R12996 VSS.n2127 VSS.n2126 0.0685147
R12997 VSS.n2105 VSS.n2104 0.0685147
R12998 VSS.n2091 VSS.n2090 0.0685147
R12999 VSS.n396 VSS.n395 0.0685147
R13000 VSS.n392 VSS.n391 0.0685147
R13001 VSS.n385 VSS.n384 0.0685147
R13002 VSS.n1974 VSS.n1973 0.0685147
R13003 VSS.n1759 VSS.n1758 0.0685147
R13004 VSS.n1755 VSS.n1754 0.0685147
R13005 VSS.n1748 VSS.n1747 0.0685147
R13006 VSS.n1695 VSS.n1694 0.0685147
R13007 VSS.n1702 VSS.n1701 0.0685147
R13008 VSS.n1893 VSS.n1892 0.0685147
R13009 VSS.n1889 VSS.n1888 0.0685147
R13010 VSS.n1882 VSS.n1881 0.0685147
R13011 VSS.n1788 VSS.n1787 0.0685147
R13012 VSS.n2165 VSS.n2164 0.0685147
R13013 VSS.n2175 VSS.n2174 0.0685147
R13014 VSS.n1612 VSS.n1611 0.0685147
R13015 VSS.n2117 VSS.n2116 0.0685147
R13016 VSS.n2103 VSS.n2102 0.0685147
R13017 VSS.n1560 VSS.n1559 0.0685147
R13018 VSS.n1567 VSS.n1566 0.0685147
R13019 VSS.n550 VSS.n549 0.0685147
R13020 VSS.n546 VSS.n545 0.0685147
R13021 VSS.n539 VSS.n538 0.0685147
R13022 VSS.n624 VSS.n623 0.0685147
R13023 VSS.n643 VSS.n642 0.0685147
R13024 VSS.n639 VSS.n638 0.0685147
R13025 VSS.n634 VSS.n633 0.0685147
R13026 VSS.n653 VSS.n652 0.0685147
R13027 VSS.n663 VSS.n662 0.0685147
R13028 VSS.n2447 VSS.n2441 0.0656042
R13029 VSS.n1307 VSS.n1267 0.0656042
R13030 VSS.n1652 VSS.n1499 0.06489
R13031 VSS.n705 VSS.n704 0.0643021
R13032 VSS.n2303 VSS.n2294 0.0643021
R13033 VSS.n1346 VSS.n1345 0.0637236
R13034 VSS.n1479 VSS.n1478 0.0635421
R13035 VSS.n2618 VSS.n243 0.0620273
R13036 VSS.n1160 VSS.n1120 0.061334
R13037 VSS.n2441 VSS 0.0603958
R13038 VSS VSS.n1307 0.0603958
R13039 VSS.n526 VSS.n525 0.0593248
R13040 VSS.n1344 VSS.n1343 0.0572917
R13041 VSS.n1921 VSS 0.0560168
R13042 VSS.n2 VSS 0.0548478
R13043 VSS.n2456 VSS 0.0548478
R13044 VSS.n1922 VSS.n1921 0.0524782
R13045 VSS.n1300 VSS.n1296 0.0518289
R13046 VSS.n1341 VSS.n1340 0.0517727
R13047 VSS.n718 VSS 0.0512812
R13048 VSS VSS.n2228 0.0512812
R13049 VSS VSS.n2352 0.0512812
R13050 VSS.n1276 VSS 0.0512812
R13051 VSS VSS.n351 0.0506333
R13052 VSS.n1927 VSS.n1922 0.0505748
R13053 VSS.n1479 VSS.n435 0.0496761
R13054 VSS VSS.n2452 0.0492848
R13055 VSS.n2862 VSS.n9 0.0491931
R13056 VSS.n735 VSS.n734 0.0482941
R13057 VSS.n741 VSS.n740 0.0482941
R13058 VSS.n747 VSS.n746 0.0482941
R13059 VSS.n282 VSS.n281 0.0482941
R13060 VSS.n300 VSS.n299 0.0482941
R13061 VSS.n1032 VSS.n1031 0.0482941
R13062 VSS.n1038 VSS.n1037 0.0482941
R13063 VSS.n812 VSS.n811 0.0482941
R13064 VSS.n842 VSS.n841 0.0482941
R13065 VSS.n853 VSS.n852 0.0482941
R13066 VSS.n909 VSS.n908 0.0482941
R13067 VSS.n915 VSS.n914 0.0482941
R13068 VSS.n921 VSS.n920 0.0482941
R13069 VSS.n2779 VSS.n2778 0.0482941
R13070 VSS.n19 VSS.n18 0.0482941
R13071 VSS.n25 VSS.n24 0.0482941
R13072 VSS.n1141 VSS.n1140 0.0482941
R13073 VSS.n1135 VSS.n1134 0.0482941
R13074 VSS.n50 VSS.n49 0.0482941
R13075 VSS.n81 VSS.n80 0.0482941
R13076 VSS.n92 VSS.n91 0.0482941
R13077 VSS.n103 VSS.n102 0.0482941
R13078 VSS.n128 VSS.n127 0.0482941
R13079 VSS.n141 VSS.n140 0.0482941
R13080 VSS.n147 VSS.n146 0.0482941
R13081 VSS.n193 VSS.n192 0.0482941
R13082 VSS.n199 VSS.n198 0.0482941
R13083 VSS.n205 VSS.n204 0.0482941
R13084 VSS.n2527 VSS.n2526 0.0482941
R13085 VSS.n2521 VSS.n2520 0.0482941
R13086 VSS.n2515 VSS.n2514 0.0482941
R13087 VSS.n2404 VSS.n2403 0.0482941
R13088 VSS.n2398 VSS.n2397 0.0482941
R13089 VSS.n2367 VSS.n2366 0.0482941
R13090 VSS.n2137 VSS.n2136 0.0482941
R13091 VSS.n2131 VSS.n2130 0.0482941
R13092 VSS.n373 VSS.n372 0.0482941
R13093 VSS.n403 VSS.n402 0.0482941
R13094 VSS.n409 VSS.n408 0.0482941
R13095 VSS.n415 VSS.n414 0.0482941
R13096 VSS.n430 VSS.n429 0.0482941
R13097 VSS.n1946 VSS.n1945 0.0482941
R13098 VSS.n1957 VSS.n1956 0.0482941
R13099 VSS.n2013 VSS.n2012 0.0482941
R13100 VSS.n2019 VSS.n2018 0.0482941
R13101 VSS.n2025 VSS.n2024 0.0482941
R13102 VSS.n1900 VSS.n1899 0.0482941
R13103 VSS.n1864 VSS.n1863 0.0482941
R13104 VSS.n1853 VSS.n1852 0.0482941
R13105 VSS.n1835 VSS.n1834 0.0482941
R13106 VSS.n1819 VSS.n1818 0.0482941
R13107 VSS.n1802 VSS.n1801 0.0482941
R13108 VSS.n1766 VSS.n1765 0.0482941
R13109 VSS.n1730 VSS.n1729 0.0482941
R13110 VSS.n1619 VSS.n1618 0.0482941
R13111 VSS.n1602 VSS.n1601 0.0482941
R13112 VSS.n1591 VSS.n1590 0.0482941
R13113 VSS.n1399 VSS.n1398 0.0482941
R13114 VSS.n1393 VSS.n1392 0.0482941
R13115 VSS.n1387 VSS.n1386 0.0482941
R13116 VSS.n569 VSS.n568 0.0482941
R13117 VSS.n563 VSS.n562 0.0482941
R13118 VSS.n557 VSS.n556 0.0482941
R13119 VSS.n472 VSS.n471 0.0482941
R13120 VSS.n478 VSS.n477 0.0482941
R13121 VSS.n484 VSS.n483 0.0482941
R13122 VSS.n2590 VSS.n2589 0.0482941
R13123 VSS.n2602 VSS.n2601 0.0482941
R13124 VSS.n817 VSS 0.0479063
R13125 VSS.n1365 VSS.n1364 0.0476858
R13126 VSS.n333 VSS 0.0471846
R13127 VSS.n1927 VSS 0.0466376
R13128 VSS.n1302 VSS.n1268 0.0444189
R13129 VSS.n2449 VSS.n2448 0.0444189
R13130 VSS.n8 VSS.n7 0.0434688
R13131 VSS.n2462 VSS.n2455 0.0434688
R13132 VSS.n707 VSS.n698 0.0427297
R13133 VSS.n2298 VSS.n2297 0.0427297
R13134 VSS.n2468 VSS.n2220 0.0425162
R13135 VSS.n936 VSS.n243 0.0424314
R13136 VSS.n769 VSS.n765 0.0415156
R13137 VSS.n2501 VSS.n253 0.0415156
R13138 VSS.n1373 VSS.n674 0.0415156
R13139 VSS.n515 VSS.n511 0.0415156
R13140 VSS.n338 VSS.n334 0.0415156
R13141 VSS.n2476 VSS.n2472 0.0415156
R13142 VSS.n711 VSS.n710 0.0411354
R13143 VSS.n2260 VSS.n2222 0.0411354
R13144 VSS.n2318 VSS.n2317 0.0411354
R13145 VSS.n1299 VSS.n1297 0.0411354
R13146 VSS.n1503 VSS.n351 0.039647
R13147 VSS.n2861 VSS.n2860 0.039516
R13148 VSS.n607 VSS 0.0393305
R13149 VSS.n1120 VSS.n1119 0.0392005
R13150 VSS.n1247 VSS.n1246 0.0391029
R13151 VSS.n1245 VSS.n1244 0.0391029
R13152 VSS.n1243 VSS.n1242 0.0391029
R13153 VSS.n1241 VSS.n1240 0.0391029
R13154 VSS.n1236 VSS.n1235 0.0391029
R13155 VSS.n1234 VSS.n1233 0.0391029
R13156 VSS.n733 VSS.n732 0.0391029
R13157 VSS.n737 VSS.n736 0.0391029
R13158 VSS.n739 VSS.n738 0.0391029
R13159 VSS.n743 VSS.n742 0.0391029
R13160 VSS.n745 VSS.n744 0.0391029
R13161 VSS.n749 VSS.n748 0.0391029
R13162 VSS.n2580 VSS.n2575 0.0391029
R13163 VSS.n2574 VSS.n2573 0.0391029
R13164 VSS.n2572 VSS.n2568 0.0391029
R13165 VSS.n2614 VSS.n2607 0.0391029
R13166 VSS.n2613 VSS.n2612 0.0391029
R13167 VSS.n2560 VSS.n2557 0.0391029
R13168 VSS.n272 VSS.n268 0.0391029
R13169 VSS.n267 VSS.n266 0.0391029
R13170 VSS.n265 VSS.n264 0.0391029
R13171 VSS.n308 VSS.n302 0.0391029
R13172 VSS.n307 VSS.n303 0.0391029
R13173 VSS.n326 VSS.n323 0.0391029
R13174 VSS.n275 VSS.n274 0.0391029
R13175 VSS.n286 VSS.n283 0.0391029
R13176 VSS.n285 VSS.n284 0.0391029
R13177 VSS.n312 VSS.n301 0.0391029
R13178 VSS.n311 VSS.n310 0.0391029
R13179 VSS.n328 VSS.n322 0.0391029
R13180 VSS.n238 VSS.n237 0.0391029
R13181 VSS.n2630 VSS.n2626 0.0391029
R13182 VSS.n2632 VSS.n2631 0.0391029
R13183 VSS.n2637 VSS.n2633 0.0391029
R13184 VSS.n2639 VSS.n2638 0.0391029
R13185 VSS.n2644 VSS.n2640 0.0391029
R13186 VSS.n241 VSS.n240 0.0391029
R13187 VSS.n2671 VSS.n2670 0.0391029
R13188 VSS.n2674 VSS.n2673 0.0391029
R13189 VSS.n2657 VSS.n2656 0.0391029
R13190 VSS.n2660 VSS.n2659 0.0391029
R13191 VSS.n2625 VSS.n2624 0.0391029
R13192 VSS.n1111 VSS.n1110 0.0391029
R13193 VSS.n1093 VSS.n1089 0.0391029
R13194 VSS.n995 VSS.n991 0.0391029
R13195 VSS.n997 VSS.n996 0.0391029
R13196 VSS.n1002 VSS.n998 0.0391029
R13197 VSS.n1114 VSS.n1113 0.0391029
R13198 VSS.n1088 VSS.n1087 0.0391029
R13199 VSS.n1097 VSS.n1096 0.0391029
R13200 VSS.n1074 VSS.n1073 0.0391029
R13201 VSS.n1077 VSS.n1076 0.0391029
R13202 VSS.n989 VSS.n988 0.0391029
R13203 VSS.n1029 VSS.n1025 0.0391029
R13204 VSS.n1024 VSS.n1023 0.0391029
R13205 VSS.n1022 VSS.n1021 0.0391029
R13206 VSS.n1020 VSS.n1019 0.0391029
R13207 VSS.n1018 VSS.n1014 0.0391029
R13208 VSS.n1013 VSS.n1012 0.0391029
R13209 VSS.n1034 VSS.n1033 0.0391029
R13210 VSS.n1041 VSS.n1036 0.0391029
R13211 VSS.n1040 VSS.n1039 0.0391029
R13212 VSS.n1046 VSS.n1042 0.0391029
R13213 VSS.n1045 VSS.n1044 0.0391029
R13214 VSS.n802 VSS.n800 0.0391029
R13215 VSS.n810 VSS.n809 0.0391029
R13216 VSS.n838 VSS.n834 0.0391029
R13217 VSS.n840 VSS.n839 0.0391029
R13218 VSS.n867 VSS.n863 0.0391029
R13219 VSS.n869 VSS.n868 0.0391029
R13220 VSS.n874 VSS.n870 0.0391029
R13221 VSS.n814 VSS.n813 0.0391029
R13222 VSS.n833 VSS.n832 0.0391029
R13223 VSS.n844 VSS.n843 0.0391029
R13224 VSS.n851 VSS.n850 0.0391029
R13225 VSS.n855 VSS.n854 0.0391029
R13226 VSS.n862 VSS.n861 0.0391029
R13227 VSS.n906 VSS.n902 0.0391029
R13228 VSS.n901 VSS.n900 0.0391029
R13229 VSS.n899 VSS.n898 0.0391029
R13230 VSS.n897 VSS.n896 0.0391029
R13231 VSS.n895 VSS.n891 0.0391029
R13232 VSS.n890 VSS.n889 0.0391029
R13233 VSS.n911 VSS.n910 0.0391029
R13234 VSS.n918 VSS.n913 0.0391029
R13235 VSS.n917 VSS.n916 0.0391029
R13236 VSS.n924 VSS.n919 0.0391029
R13237 VSS.n923 VSS.n922 0.0391029
R13238 VSS.n927 VSS.n925 0.0391029
R13239 VSS.n2852 VSS.n2851 0.0391029
R13240 VSS.n2836 VSS.n2832 0.0391029
R13241 VSS.n2796 VSS.n2792 0.0391029
R13242 VSS.n2798 VSS.n2797 0.0391029
R13243 VSS.n2804 VSS.n2799 0.0391029
R13244 VSS.n2855 VSS.n2854 0.0391029
R13245 VSS.n2829 VSS.n2828 0.0391029
R13246 VSS.n2838 VSS.n2831 0.0391029
R13247 VSS.n2815 VSS.n2814 0.0391029
R13248 VSS.n2818 VSS.n2817 0.0391029
R13249 VSS.n2790 VSS.n2789 0.0391029
R13250 VSS.n2776 VSS.n2772 0.0391029
R13251 VSS.n2771 VSS.n2770 0.0391029
R13252 VSS.n2769 VSS.n2768 0.0391029
R13253 VSS.n2767 VSS.n2766 0.0391029
R13254 VSS.n2765 VSS.n2754 0.0391029
R13255 VSS.n2753 VSS.n2752 0.0391029
R13256 VSS.n2781 VSS.n2780 0.0391029
R13257 VSS.n22 VSS.n17 0.0391029
R13258 VSS.n21 VSS.n20 0.0391029
R13259 VSS.n28 VSS.n23 0.0391029
R13260 VSS.n27 VSS.n26 0.0391029
R13261 VSS.n31 VSS.n29 0.0391029
R13262 VSS.n1224 VSS.n790 0.0391029
R13263 VSS.n1210 VSS.n1206 0.0391029
R13264 VSS.n1172 VSS.n1168 0.0391029
R13265 VSS.n1174 VSS.n1173 0.0391029
R13266 VSS.n1179 VSS.n1175 0.0391029
R13267 VSS.n1223 VSS.n793 0.0391029
R13268 VSS.n1205 VSS.n1204 0.0391029
R13269 VSS.n1214 VSS.n1213 0.0391029
R13270 VSS.n1191 VSS.n1190 0.0391029
R13271 VSS.n1194 VSS.n1193 0.0391029
R13272 VSS.n1166 VSS.n1165 0.0391029
R13273 VSS.n1132 VSS.n1131 0.0391029
R13274 VSS.n2757 VSS.n2756 0.0391029
R13275 VSS.n2743 VSS.n2742 0.0391029
R13276 VSS.n2741 VSS.n2740 0.0391029
R13277 VSS.n1143 VSS.n1142 0.0391029
R13278 VSS.n1139 VSS.n1138 0.0391029
R13279 VSS.n1137 VSS.n1136 0.0391029
R13280 VSS.n48 VSS.n47 0.0391029
R13281 VSS.n52 VSS.n51 0.0391029
R13282 VSS.n78 VSS.n74 0.0391029
R13283 VSS.n73 VSS.n72 0.0391029
R13284 VSS.n71 VSS.n70 0.0391029
R13285 VSS.n69 VSS.n68 0.0391029
R13286 VSS.n67 VSS.n63 0.0391029
R13287 VSS.n62 VSS.n61 0.0391029
R13288 VSS.n83 VSS.n82 0.0391029
R13289 VSS.n95 VSS.n90 0.0391029
R13290 VSS.n94 VSS.n93 0.0391029
R13291 VSS.n106 VSS.n101 0.0391029
R13292 VSS.n105 VSS.n104 0.0391029
R13293 VSS.n114 VSS.n112 0.0391029
R13294 VSS.n126 VSS.n125 0.0391029
R13295 VSS.n137 VSS.n133 0.0391029
R13296 VSS.n139 VSS.n138 0.0391029
R13297 VSS.n156 VSS.n152 0.0391029
R13298 VSS.n158 VSS.n157 0.0391029
R13299 VSS.n163 VSS.n159 0.0391029
R13300 VSS.n130 VSS.n129 0.0391029
R13301 VSS.n132 VSS.n131 0.0391029
R13302 VSS.n143 VSS.n142 0.0391029
R13303 VSS.n145 VSS.n144 0.0391029
R13304 VSS.n149 VSS.n148 0.0391029
R13305 VSS.n151 VSS.n150 0.0391029
R13306 VSS.n190 VSS.n186 0.0391029
R13307 VSS.n185 VSS.n184 0.0391029
R13308 VSS.n183 VSS.n182 0.0391029
R13309 VSS.n181 VSS.n180 0.0391029
R13310 VSS.n179 VSS.n175 0.0391029
R13311 VSS.n174 VSS.n173 0.0391029
R13312 VSS.n195 VSS.n194 0.0391029
R13313 VSS.n202 VSS.n197 0.0391029
R13314 VSS.n201 VSS.n200 0.0391029
R13315 VSS.n208 VSS.n203 0.0391029
R13316 VSS.n207 VSS.n206 0.0391029
R13317 VSS.n211 VSS.n209 0.0391029
R13318 VSS.n2509 VSS.n251 0.0391029
R13319 VSS.n2272 VSS.n2271 0.0391029
R13320 VSS.n2277 VSS.n2276 0.0391029
R13321 VSS.n2279 VSS.n2278 0.0391029
R13322 VSS.n2284 VSS.n2283 0.0391029
R13323 VSS.n2286 VSS.n2285 0.0391029
R13324 VSS.n2529 VSS.n2528 0.0391029
R13325 VSS.n2525 VSS.n2524 0.0391029
R13326 VSS.n2523 VSS.n2522 0.0391029
R13327 VSS.n2519 VSS.n2518 0.0391029
R13328 VSS.n2517 VSS.n2516 0.0391029
R13329 VSS.n2513 VSS.n2512 0.0391029
R13330 VSS.n2426 VSS.n2394 0.0391029
R13331 VSS.n2393 VSS.n2392 0.0391029
R13332 VSS.n2388 VSS.n2387 0.0391029
R13333 VSS.n2386 VSS.n2385 0.0391029
R13334 VSS.n2381 VSS.n2380 0.0391029
R13335 VSS.n2379 VSS.n2378 0.0391029
R13336 VSS.n2425 VSS.n2405 0.0391029
R13337 VSS.n2402 VSS.n2401 0.0391029
R13338 VSS.n2400 VSS.n2399 0.0391029
R13339 VSS.n2365 VSS.n2364 0.0391029
R13340 VSS.n2369 VSS.n2368 0.0391029
R13341 VSS.n445 VSS.n444 0.0391029
R13342 VSS.n1466 VSS.n1462 0.0391029
R13343 VSS.n461 VSS.n457 0.0391029
R13344 VSS.n463 VSS.n462 0.0391029
R13345 VSS.n468 VSS.n464 0.0391029
R13346 VSS.n448 VSS.n447 0.0391029
R13347 VSS.n1461 VSS.n1460 0.0391029
R13348 VSS.n1470 VSS.n1469 0.0391029
R13349 VSS.n1447 VSS.n1446 0.0391029
R13350 VSS.n1450 VSS.n1449 0.0391029
R13351 VSS.n455 VSS.n454 0.0391029
R13352 VSS.n2010 VSS.n2006 0.0391029
R13353 VSS.n2005 VSS.n2004 0.0391029
R13354 VSS.n2003 VSS.n2002 0.0391029
R13355 VSS.n2001 VSS.n2000 0.0391029
R13356 VSS.n1999 VSS.n1995 0.0391029
R13357 VSS.n1994 VSS.n1993 0.0391029
R13358 VSS.n2128 VSS.n2127 0.0391029
R13359 VSS.n2106 VSS.n2105 0.0391029
R13360 VSS.n2092 VSS.n2091 0.0391029
R13361 VSS.n2090 VSS.n2089 0.0391029
R13362 VSS.n2139 VSS.n2138 0.0391029
R13363 VSS.n2135 VSS.n2134 0.0391029
R13364 VSS.n2133 VSS.n2132 0.0391029
R13365 VSS.n371 VSS.n370 0.0391029
R13366 VSS.n375 VSS.n374 0.0391029
R13367 VSS.n400 VSS.n396 0.0391029
R13368 VSS.n395 VSS.n394 0.0391029
R13369 VSS.n393 VSS.n392 0.0391029
R13370 VSS.n391 VSS.n390 0.0391029
R13371 VSS.n389 VSS.n385 0.0391029
R13372 VSS.n384 VSS.n383 0.0391029
R13373 VSS.n405 VSS.n404 0.0391029
R13374 VSS.n412 VSS.n407 0.0391029
R13375 VSS.n411 VSS.n410 0.0391029
R13376 VSS.n418 VSS.n413 0.0391029
R13377 VSS.n417 VSS.n416 0.0391029
R13378 VSS.n421 VSS.n419 0.0391029
R13379 VSS.n428 VSS.n427 0.0391029
R13380 VSS.n1942 VSS.n1938 0.0391029
R13381 VSS.n1944 VSS.n1943 0.0391029
R13382 VSS.n1971 VSS.n1967 0.0391029
R13383 VSS.n1973 VSS.n1972 0.0391029
R13384 VSS.n1978 VSS.n1974 0.0391029
R13385 VSS.n432 VSS.n431 0.0391029
R13386 VSS.n1937 VSS.n1936 0.0391029
R13387 VSS.n1948 VSS.n1947 0.0391029
R13388 VSS.n1955 VSS.n1954 0.0391029
R13389 VSS.n1959 VSS.n1958 0.0391029
R13390 VSS.n1966 VSS.n1965 0.0391029
R13391 VSS.n2015 VSS.n2014 0.0391029
R13392 VSS.n2022 VSS.n2017 0.0391029
R13393 VSS.n2021 VSS.n2020 0.0391029
R13394 VSS.n2028 VSS.n2023 0.0391029
R13395 VSS.n2027 VSS.n2026 0.0391029
R13396 VSS.n2031 VSS.n2029 0.0391029
R13397 VSS.n1763 VSS.n1759 0.0391029
R13398 VSS.n1758 VSS.n1757 0.0391029
R13399 VSS.n1756 VSS.n1755 0.0391029
R13400 VSS.n1754 VSS.n1753 0.0391029
R13401 VSS.n1752 VSS.n1748 0.0391029
R13402 VSS.n1747 VSS.n1746 0.0391029
R13403 VSS.n1646 VSS.n1645 0.0391029
R13404 VSS.n1666 VSS.n1662 0.0391029
R13405 VSS.n1699 VSS.n1695 0.0391029
R13406 VSS.n1701 VSS.n1700 0.0391029
R13407 VSS.n1706 VSS.n1702 0.0391029
R13408 VSS.n1647 VSS.n1640 0.0391029
R13409 VSS.n1661 VSS.n1660 0.0391029
R13410 VSS.n1670 VSS.n1669 0.0391029
R13411 VSS.n1681 VSS.n1680 0.0391029
R13412 VSS.n1684 VSS.n1683 0.0391029
R13413 VSS.n1693 VSS.n1692 0.0391029
R13414 VSS.n1897 VSS.n1893 0.0391029
R13415 VSS.n1892 VSS.n1891 0.0391029
R13416 VSS.n1890 VSS.n1889 0.0391029
R13417 VSS.n1888 VSS.n1887 0.0391029
R13418 VSS.n1886 VSS.n1882 0.0391029
R13419 VSS.n1881 VSS.n1880 0.0391029
R13420 VSS.n1902 VSS.n1901 0.0391029
R13421 VSS.n1867 VSS.n1862 0.0391029
R13422 VSS.n1866 VSS.n1865 0.0391029
R13423 VSS.n1856 VSS.n1851 0.0391029
R13424 VSS.n1855 VSS.n1854 0.0391029
R13425 VSS.n1845 VSS.n1843 0.0391029
R13426 VSS.n1833 VSS.n1832 0.0391029
R13427 VSS.n1815 VSS.n1811 0.0391029
R13428 VSS.n1817 VSS.n1816 0.0391029
R13429 VSS.n1785 VSS.n1781 0.0391029
R13430 VSS.n1787 VSS.n1786 0.0391029
R13431 VSS.n1792 VSS.n1788 0.0391029
R13432 VSS.n1837 VSS.n1836 0.0391029
R13433 VSS.n1810 VSS.n1809 0.0391029
R13434 VSS.n1821 VSS.n1820 0.0391029
R13435 VSS.n1800 VSS.n1799 0.0391029
R13436 VSS.n1804 VSS.n1803 0.0391029
R13437 VSS.n1780 VSS.n1779 0.0391029
R13438 VSS.n1768 VSS.n1767 0.0391029
R13439 VSS.n1733 VSS.n1728 0.0391029
R13440 VSS.n1732 VSS.n1731 0.0391029
R13441 VSS.n1722 VSS.n1718 0.0391029
R13442 VSS.n1721 VSS.n1720 0.0391029
R13443 VSS.n603 VSS.n601 0.0391029
R13444 VSS.n358 VSS.n357 0.0391029
R13445 VSS.n2212 VSS.n2209 0.0391029
R13446 VSS.n2172 VSS.n2165 0.0391029
R13447 VSS.n2174 VSS.n2173 0.0391029
R13448 VSS.n2179 VSS.n2175 0.0391029
R13449 VSS.n361 VSS.n360 0.0391029
R13450 VSS.n2206 VSS.n2205 0.0391029
R13451 VSS.n2214 VSS.n2208 0.0391029
R13452 VSS.n2192 VSS.n2191 0.0391029
R13453 VSS.n2195 VSS.n2194 0.0391029
R13454 VSS.n2163 VSS.n2162 0.0391029
R13455 VSS.n1514 VSS.n1513 0.0391029
R13456 VSS.n1527 VSS.n1526 0.0391029
R13457 VSS.n1535 VSS.n1534 0.0391029
R13458 VSS.n1546 VSS.n1545 0.0391029
R13459 VSS.n1549 VSS.n1548 0.0391029
R13460 VSS.n1558 VSS.n1557 0.0391029
R13461 VSS.n1616 VSS.n1612 0.0391029
R13462 VSS.n1611 VSS.n368 0.0391029
R13463 VSS.n2118 VSS.n2117 0.0391029
R13464 VSS.n2116 VSS.n2115 0.0391029
R13465 VSS.n2114 VSS.n2103 0.0391029
R13466 VSS.n2102 VSS.n2101 0.0391029
R13467 VSS.n1621 VSS.n1620 0.0391029
R13468 VSS.n1605 VSS.n1600 0.0391029
R13469 VSS.n1604 VSS.n1603 0.0391029
R13470 VSS.n1594 VSS.n1589 0.0391029
R13471 VSS.n1593 VSS.n1592 0.0391029
R13472 VSS.n1583 VSS.n1581 0.0391029
R13473 VSS.n1511 VSS.n1510 0.0391029
R13474 VSS.n1531 VSS.n1528 0.0391029
R13475 VSS.n1564 VSS.n1560 0.0391029
R13476 VSS.n1566 VSS.n1565 0.0391029
R13477 VSS.n1572 VSS.n1567 0.0391029
R13478 VSS.n1381 VSS.n550 0.0391029
R13479 VSS.n549 VSS.n548 0.0391029
R13480 VSS.n547 VSS.n546 0.0391029
R13481 VSS.n545 VSS.n544 0.0391029
R13482 VSS.n543 VSS.n539 0.0391029
R13483 VSS.n538 VSS.n537 0.0391029
R13484 VSS.n1401 VSS.n1400 0.0391029
R13485 VSS.n1397 VSS.n1396 0.0391029
R13486 VSS.n1395 VSS.n1394 0.0391029
R13487 VSS.n1391 VSS.n1390 0.0391029
R13488 VSS.n1389 VSS.n1388 0.0391029
R13489 VSS.n1385 VSS.n1384 0.0391029
R13490 VSS.n625 VSS.n624 0.0391029
R13491 VSS.n623 VSS.n622 0.0391029
R13492 VSS.n644 VSS.n643 0.0391029
R13493 VSS.n642 VSS.n641 0.0391029
R13494 VSS.n640 VSS.n639 0.0391029
R13495 VSS.n638 VSS.n637 0.0391029
R13496 VSS.n571 VSS.n570 0.0391029
R13497 VSS.n567 VSS.n566 0.0391029
R13498 VSS.n565 VSS.n564 0.0391029
R13499 VSS.n561 VSS.n560 0.0391029
R13500 VSS.n559 VSS.n558 0.0391029
R13501 VSS.n555 VSS.n554 0.0391029
R13502 VSS.n633 VSS.n632 0.0391029
R13503 VSS.n635 VSS.n634 0.0391029
R13504 VSS.n652 VSS.n651 0.0391029
R13505 VSS.n654 VSS.n653 0.0391029
R13506 VSS.n662 VSS.n661 0.0391029
R13507 VSS.n664 VSS.n663 0.0391029
R13508 VSS.n474 VSS.n473 0.0391029
R13509 VSS.n481 VSS.n476 0.0391029
R13510 VSS.n480 VSS.n479 0.0391029
R13511 VSS.n487 VSS.n482 0.0391029
R13512 VSS.n486 VSS.n485 0.0391029
R13513 VSS.n490 VSS.n488 0.0391029
R13514 VSS.n2583 VSS.n2582 0.0391029
R13515 VSS.n2594 VSS.n2591 0.0391029
R13516 VSS.n2593 VSS.n2592 0.0391029
R13517 VSS.n2615 VSS.n2603 0.0391029
R13518 VSS.n2606 VSS.n2605 0.0391029
R13519 VSS.n2561 VSS.n2555 0.0391029
R13520 VSS.n2445 VSS 0.0378217
R13521 VSS.n1304 VSS 0.0378217
R13522 VSS.n1280 VSS.n1279 0.0376053
R13523 VSS.n1362 VSS.n1351 0.0375879
R13524 VSS.n2253 VSS.n2252 0.0361962
R13525 VSS.n2328 VSS.n2327 0.0361962
R13526 VSS.n2307 VSS.n2306 0.035973
R13527 VSS.n2309 VSS.n2308 0.035973
R13528 VSS.n694 VSS.n693 0.035973
R13529 VSS.n714 VSS.n695 0.035973
R13530 VSS.n2263 VSS.n2248 0.035973
R13531 VSS.n2250 VSS.n2249 0.035973
R13532 VSS.n1292 VSS.n1265 0.035973
R13533 VSS.n1310 VSS.n1309 0.035973
R13534 VSS.n2862 VSS.n2861 0.035918
R13535 VSS VSS.n2156 0.0358842
R13536 VSS.n1422 VSS.n509 0.0356615
R13537 VSS.n2498 VSS.n2497 0.0345671
R13538 VSS.n2447 VSS.n2446 0.0343542
R13539 VSS.n1303 VSS.n1267 0.0343542
R13540 VSS VSS.n2549 0.034115
R13541 VSS VSS.n2682 0.0338434
R13542 VSS.n706 VSS 0.0330521
R13543 VSS VSS.n2439 0.0330521
R13544 VSS VSS.n2295 0.0330521
R13545 VSS.n1308 VSS 0.0330521
R13546 VSS.n1283 VSS.n1273 0.0325946
R13547 VSS.n2332 VSS.n2312 0.0325946
R13548 VSS.n2226 VSS.n2225 0.0325946
R13549 VSS.n1337 VSS.n680 0.0325946
R13550 VSS.n936 VSS 0.0325669
R13551 VSS VSS.n716 0.03175
R13552 VSS.n2353 VSS 0.03175
R13553 VSS.n2693 VSS 0.0299577
R13554 VSS.n678 VSS.n677 0.029875
R13555 VSS.n2258 VSS.n2257 0.029875
R13556 VSS.n2323 VSS.n2322 0.029875
R13557 VSS.n1281 VSS.n1271 0.029875
R13558 VSS.n608 VSS 0.0298356
R13559 VSS VSS.n606 0.0298356
R13560 VSS.n1689 VSS 0.0298356
R13561 VSS VSS.n1915 0.0298356
R13562 VSS.n1554 VSS 0.0298356
R13563 VSS VSS.n1634 0.0298356
R13564 VSS VSS.n332 0.0297375
R13565 VSS.n956 VSS 0.0297375
R13566 VSS VSS.n10 0.0297375
R13567 VSS.n984 VSS 0.0297375
R13568 VSS.n3 VSS 0.0285374
R13569 VSS.n2457 VSS 0.0285374
R13570 VSS.n716 VSS.n715 0.0278438
R13571 VSS.n2264 VSS.n2247 0.0278438
R13572 VSS.n2354 VSS.n2353 0.0278438
R13573 VSS.n1291 VSS.n1263 0.0278438
R13574 VSS.n2157 VSS 0.0272339
R13575 VSS VSS.n450 0.0272339
R13576 VSS.n2050 VSS 0.0272339
R13577 VSS.n1423 VSS 0.0272339
R13578 VSS.n1483 VSS 0.0272339
R13579 VSS.n2861 VSS 0.0269789
R13580 VSS.n1636 VSS.n1635 0.0266812
R13581 VSS VSS.n1422 0.0263989
R13582 VSS.n1342 VSS.n1341 0.0261364
R13583 VSS.n2503 VSS.n2502 0.0257686
R13584 VSS.n1375 VSS.n1374 0.0257686
R13585 VSS.n1161 VSS 0.0256931
R13586 VSS.n2718 VSS 0.0256931
R13587 VSS.n2683 VSS 0.0256931
R13588 VSS VSS.n2496 0.0256931
R13589 VSS.n2550 VSS 0.0256931
R13590 VSS.n1343 VSS.n1342 0.0252818
R13591 VSS.n1499 VSS.n1493 0.025078
R13592 VSS VSS.n2487 0.024393
R13593 VSS.n2460 VSS.n2459 0.0241592
R13594 VSS.n5 VSS.n4 0.0241592
R13595 VSS VSS.n509 0.0240791
R13596 VSS.n767 VSS.n766 0.024008
R13597 VSS.n513 VSS.n512 0.024008
R13598 VSS.n336 VSS.n335 0.024008
R13599 VSS.n2474 VSS.n2473 0.024008
R13600 VSS.n289 VSS.n243 0.0227182
R13601 VSS.n1334 VSS 0.0226354
R13602 VSS.n2438 VSS.n2437 0.0226354
R13603 VSS.n2310 VSS 0.0226354
R13604 VSS.n1311 VSS.n1264 0.0226354
R13605 VSS.n2501 VSS.n252 0.0223823
R13606 VSS.n1373 VSS.n673 0.0223823
R13607 VSS.n732 VSS.n731 0.0219755
R13608 VSS.n328 VSS.n327 0.0219755
R13609 VSS.n241 VSS.n232 0.0219755
R13610 VSS.n1114 VSS.n1105 0.0219755
R13611 VSS.n802 VSS.n801 0.0219755
R13612 VSS.n814 VSS.n804 0.0219755
R13613 VSS.n927 VSS.n926 0.0219755
R13614 VSS.n2855 VSS.n2846 0.0219755
R13615 VSS.n31 VSS.n30 0.0219755
R13616 VSS.n1223 VSS.n791 0.0219755
R13617 VSS.n1143 VSS.n1123 0.0219755
R13618 VSS.n114 VSS.n113 0.0219755
R13619 VSS.n130 VSS.n120 0.0219755
R13620 VSS.n211 VSS.n210 0.0219755
R13621 VSS.n2512 VSS.n2511 0.0219755
R13622 VSS.n2425 VSS.n2395 0.0219755
R13623 VSS.n448 VSS.n439 0.0219755
R13624 VSS.n2139 VSS.n367 0.0219755
R13625 VSS.n421 VSS.n420 0.0219755
R13626 VSS.n432 VSS.n422 0.0219755
R13627 VSS.n2031 VSS.n2030 0.0219755
R13628 VSS.n1647 VSS.n1638 0.0219755
R13629 VSS.n1845 VSS.n1844 0.0219755
R13630 VSS.n1837 VSS.n1827 0.0219755
R13631 VSS.n603 VSS.n602 0.0219755
R13632 VSS.n361 VSS.n353 0.0219755
R13633 VSS.n1514 VSS.n1505 0.0219755
R13634 VSS.n1583 VSS.n1582 0.0219755
R13635 VSS.n1384 VSS.n1383 0.0219755
R13636 VSS.n554 VSS.n553 0.0219755
R13637 VSS.n490 VSS.n489 0.0219755
R13638 VSS.n2561 VSS.n2556 0.0219755
R13639 VSS.n692 VSS.n683 0.0213333
R13640 VSS.n2227 VSS.n2223 0.0213333
R13641 VSS.n2355 VSS.n2305 0.0213333
R13642 VSS.n1275 VSS.n1256 0.0213333
R13643 VSS.n2469 VSS.n2468 0.0211532
R13644 VSS VSS.n825 0.0201488
R13645 VSS.n1336 VSS.n1333 0.0200312
R13646 VSS.n2334 VSS.n2333 0.0200312
R13647 VSS VSS.n1480 0.0194262
R13648 VSS.n1916 VSS 0.0194262
R13649 VSS VSS.n1500 0.0194262
R13650 VSS VSS.n955 0.0193629
R13651 VSS VSS.n983 0.0193629
R13652 VSS.n826 VSS 0.0193629
R13653 VSS.n752 VSS.n751 0.0191618
R13654 VSS.n755 VSS.n754 0.0191618
R13655 VSS.n756 VSS.n755 0.0191618
R13656 VSS.n759 VSS.n758 0.0191618
R13657 VSS.n760 VSS.n759 0.0191618
R13658 VSS.n786 VSS.n762 0.0191618
R13659 VSS.n277 VSS.n257 0.0191618
R13660 VSS.n278 VSS.n277 0.0191618
R13661 VSS.n294 VSS.n280 0.0191618
R13662 VSS.n295 VSS.n294 0.0191618
R13663 VSS.n315 VSS.n298 0.0191618
R13664 VSS.n315 VSS.n314 0.0191618
R13665 VSS.n330 VSS.n320 0.0191618
R13666 VSS.n330 VSS.n329 0.0191618
R13667 VSS.n242 VSS.n229 0.0191618
R13668 VSS.n242 VSS.n231 0.0191618
R13669 VSS.n2677 VSS.n2668 0.0191618
R13670 VSS.n2677 VSS.n2676 0.0191618
R13671 VSS.n2663 VSS.n2654 0.0191618
R13672 VSS.n2663 VSS.n2662 0.0191618
R13673 VSS.n2649 VSS.n2622 0.0191618
R13674 VSS.n2649 VSS.n2648 0.0191618
R13675 VSS.n2585 VSS.n2567 0.0191618
R13676 VSS.n2586 VSS.n2585 0.0191618
R13677 VSS.n2595 VSS.n2588 0.0191618
R13678 VSS.n2596 VSS.n2595 0.0191618
R13679 VSS.n2616 VSS.n2598 0.0191618
R13680 VSS.n2616 VSS.n2600 0.0191618
R13681 VSS.n2562 VSS.n2552 0.0191618
R13682 VSS.n2562 VSS.n2553 0.0191618
R13683 VSS.n1117 VSS.n1104 0.0191618
R13684 VSS.n1117 VSS.n1116 0.0191618
R13685 VSS.n1100 VSS.n1085 0.0191618
R13686 VSS.n1100 VSS.n1099 0.0191618
R13687 VSS.n1080 VSS.n1071 0.0191618
R13688 VSS.n1080 VSS.n1079 0.0191618
R13689 VSS.n1066 VSS.n986 0.0191618
R13690 VSS.n1066 VSS.n1065 0.0191618
R13691 VSS.n1062 VSS.n1061 0.0191618
R13692 VSS.n1061 VSS.n1060 0.0191618
R13693 VSS.n1057 VSS.n1056 0.0191618
R13694 VSS.n1056 VSS.n1055 0.0191618
R13695 VSS.n1052 VSS.n1051 0.0191618
R13696 VSS.n1051 VSS.n1050 0.0191618
R13697 VSS.n972 VSS.n971 0.0191618
R13698 VSS.n968 VSS.n967 0.0191618
R13699 VSS.n967 VSS.n803 0.0191618
R13700 VSS.n845 VSS.n831 0.0191618
R13701 VSS.n846 VSS.n845 0.0191618
R13702 VSS.n856 VSS.n849 0.0191618
R13703 VSS.n857 VSS.n856 0.0191618
R13704 VSS.n877 VSS.n860 0.0191618
R13705 VSS.n878 VSS.n877 0.0191618
R13706 VSS.n953 VSS.n881 0.0191618
R13707 VSS.n953 VSS.n952 0.0191618
R13708 VSS.n949 VSS.n948 0.0191618
R13709 VSS.n948 VSS.n947 0.0191618
R13710 VSS.n944 VSS.n943 0.0191618
R13711 VSS.n943 VSS.n942 0.0191618
R13712 VSS.n939 VSS.n938 0.0191618
R13713 VSS.n938 VSS.n937 0.0191618
R13714 VSS.n2858 VSS.n2845 0.0191618
R13715 VSS.n2858 VSS.n2857 0.0191618
R13716 VSS.n2841 VSS.n2826 0.0191618
R13717 VSS.n2841 VSS.n2840 0.0191618
R13718 VSS.n2821 VSS.n2812 0.0191618
R13719 VSS.n2821 VSS.n2820 0.0191618
R13720 VSS.n2807 VSS.n12 0.0191618
R13721 VSS.n2807 VSS.n2787 0.0191618
R13722 VSS.n2784 VSS.n2783 0.0191618
R13723 VSS.n2783 VSS.n44 0.0191618
R13724 VSS.n42 VSS.n41 0.0191618
R13725 VSS.n41 VSS.n40 0.0191618
R13726 VSS.n38 VSS.n37 0.0191618
R13727 VSS.n37 VSS.n36 0.0191618
R13728 VSS.n34 VSS.n33 0.0191618
R13729 VSS.n1222 VSS.n794 0.0191618
R13730 VSS.n1222 VSS.n796 0.0191618
R13731 VSS.n1217 VSS.n1202 0.0191618
R13732 VSS.n1217 VSS.n1216 0.0191618
R13733 VSS.n1197 VSS.n1188 0.0191618
R13734 VSS.n1197 VSS.n1196 0.0191618
R13735 VSS.n1183 VSS.n1163 0.0191618
R13736 VSS.n1183 VSS.n1182 0.0191618
R13737 VSS.n1155 VSS.n1154 0.0191618
R13738 VSS.n1152 VSS.n1151 0.0191618
R13739 VSS.n1151 VSS.n1150 0.0191618
R13740 VSS.n1148 VSS.n1147 0.0191618
R13741 VSS.n1147 VSS.n1146 0.0191618
R13742 VSS.n2734 VSS.n2733 0.0191618
R13743 VSS.n2730 VSS.n2729 0.0191618
R13744 VSS.n2729 VSS.n53 0.0191618
R13745 VSS.n96 VSS.n89 0.0191618
R13746 VSS.n97 VSS.n96 0.0191618
R13747 VSS.n107 VSS.n100 0.0191618
R13748 VSS.n108 VSS.n107 0.0191618
R13749 VSS.n115 VSS.n111 0.0191618
R13750 VSS.n116 VSS.n115 0.0191618
R13751 VSS.n2715 VSS.n119 0.0191618
R13752 VSS.n2715 VSS.n2714 0.0191618
R13753 VSS.n2711 VSS.n2710 0.0191618
R13754 VSS.n2710 VSS.n2709 0.0191618
R13755 VSS.n2706 VSS.n2705 0.0191618
R13756 VSS.n2705 VSS.n2704 0.0191618
R13757 VSS.n2701 VSS.n2700 0.0191618
R13758 VSS.n2700 VSS.n2699 0.0191618
R13759 VSS.n2696 VSS.n2695 0.0191618
R13760 VSS.n2695 VSS.n227 0.0191618
R13761 VSS.n224 VSS.n223 0.0191618
R13762 VSS.n223 VSS.n222 0.0191618
R13763 VSS.n219 VSS.n218 0.0191618
R13764 VSS.n218 VSS.n217 0.0191618
R13765 VSS.n214 VSS.n213 0.0191618
R13766 VSS.n213 VSS.n212 0.0191618
R13767 VSS.n2547 VSS.n250 0.0191618
R13768 VSS.n2547 VSS.n2546 0.0191618
R13769 VSS.n2543 VSS.n2542 0.0191618
R13770 VSS.n2542 VSS.n2541 0.0191618
R13771 VSS.n2538 VSS.n2537 0.0191618
R13772 VSS.n2537 VSS.n2536 0.0191618
R13773 VSS.n2533 VSS.n2532 0.0191618
R13774 VSS.n2532 VSS.n2531 0.0191618
R13775 VSS.n2424 VSS.n2423 0.0191618
R13776 VSS.n2421 VSS.n2420 0.0191618
R13777 VSS.n2420 VSS.n2419 0.0191618
R13778 VSS.n2417 VSS.n2416 0.0191618
R13779 VSS.n2416 VSS.n2415 0.0191618
R13780 VSS.n2371 VSS.n2370 0.0191618
R13781 VSS.n2154 VSS.n366 0.0191618
R13782 VSS.n2154 VSS.n2153 0.0191618
R13783 VSS.n2150 VSS.n2149 0.0191618
R13784 VSS.n2149 VSS.n2148 0.0191618
R13785 VSS.n2145 VSS.n2144 0.0191618
R13786 VSS.n2144 VSS.n2143 0.0191618
R13787 VSS.n2083 VSS.n2082 0.0191618
R13788 VSS.n2079 VSS.n2078 0.0191618
R13789 VSS.n2078 VSS.n2077 0.0191618
R13790 VSS.n2075 VSS.n2074 0.0191618
R13791 VSS.n2074 VSS.n2073 0.0191618
R13792 VSS.n2071 VSS.n2070 0.0191618
R13793 VSS.n2070 VSS.n2069 0.0191618
R13794 VSS.n2067 VSS.n2066 0.0191618
R13795 VSS.n2066 VSS.n2065 0.0191618
R13796 VSS.n2062 VSS.n2061 0.0191618
R13797 VSS.n2061 VSS.n433 0.0191618
R13798 VSS.n1949 VSS.n1935 0.0191618
R13799 VSS.n1950 VSS.n1949 0.0191618
R13800 VSS.n1960 VSS.n1953 0.0191618
R13801 VSS.n1961 VSS.n1960 0.0191618
R13802 VSS.n1981 VSS.n1964 0.0191618
R13803 VSS.n1982 VSS.n1981 0.0191618
R13804 VSS.n2047 VSS.n1985 0.0191618
R13805 VSS.n2047 VSS.n2046 0.0191618
R13806 VSS.n2043 VSS.n2042 0.0191618
R13807 VSS.n2042 VSS.n2041 0.0191618
R13808 VSS.n2038 VSS.n2037 0.0191618
R13809 VSS.n2037 VSS.n2036 0.0191618
R13810 VSS.n2034 VSS.n2033 0.0191618
R13811 VSS.n1650 VSS.n1637 0.0191618
R13812 VSS.n1650 VSS.n1649 0.0191618
R13813 VSS.n1671 VSS.n1656 0.0191618
R13814 VSS.n1671 VSS.n1658 0.0191618
R13815 VSS.n1685 VSS.n1676 0.0191618
R13816 VSS.n1685 VSS.n1678 0.0191618
R13817 VSS.n1709 VSS.n1482 0.0191618
R13818 VSS.n1710 VSS.n1709 0.0191618
R13819 VSS.n1904 VSS.n1713 0.0191618
R13820 VSS.n1904 VSS.n1872 0.0191618
R13821 VSS.n1869 VSS.n1868 0.0191618
R13822 VSS.n1868 VSS.n1861 0.0191618
R13823 VSS.n1858 VSS.n1857 0.0191618
R13824 VSS.n1857 VSS.n1850 0.0191618
R13825 VSS.n1847 VSS.n1846 0.0191618
R13826 VSS.n1846 VSS.n1842 0.0191618
R13827 VSS.n1839 VSS.n1838 0.0191618
R13828 VSS.n1838 VSS.n1826 0.0191618
R13829 VSS.n1823 VSS.n1822 0.0191618
R13830 VSS.n1822 VSS.n1808 0.0191618
R13831 VSS.n1806 VSS.n1805 0.0191618
R13832 VSS.n1805 VSS.n1798 0.0191618
R13833 VSS.n1796 VSS.n1795 0.0191618
R13834 VSS.n1795 VSS.n1774 0.0191618
R13835 VSS.n1771 VSS.n1770 0.0191618
R13836 VSS.n1770 VSS.n1738 0.0191618
R13837 VSS.n1735 VSS.n1734 0.0191618
R13838 VSS.n1734 VSS.n1727 0.0191618
R13839 VSS.n1724 VSS.n1723 0.0191618
R13840 VSS.n1723 VSS.n1717 0.0191618
R13841 VSS.n604 VSS.n599 0.0191618
R13842 VSS.n364 VSS.n352 0.0191618
R13843 VSS.n364 VSS.n363 0.0191618
R13844 VSS.n2215 VSS.n2201 0.0191618
R13845 VSS.n2215 VSS.n2203 0.0191618
R13846 VSS.n2196 VSS.n2187 0.0191618
R13847 VSS.n2196 VSS.n2189 0.0191618
R13848 VSS.n2182 VSS.n2159 0.0191618
R13849 VSS.n2182 VSS.n2160 0.0191618
R13850 VSS.n1517 VSS.n1504 0.0191618
R13851 VSS.n1517 VSS.n1516 0.0191618
R13852 VSS.n1536 VSS.n1522 0.0191618
R13853 VSS.n1536 VSS.n1524 0.0191618
R13854 VSS.n1550 VSS.n1541 0.0191618
R13855 VSS.n1550 VSS.n1543 0.0191618
R13856 VSS.n1575 VSS.n1502 0.0191618
R13857 VSS.n1576 VSS.n1575 0.0191618
R13858 VSS.n1623 VSS.n1579 0.0191618
R13859 VSS.n1623 VSS.n1610 0.0191618
R13860 VSS.n1607 VSS.n1606 0.0191618
R13861 VSS.n1606 VSS.n1599 0.0191618
R13862 VSS.n1596 VSS.n1595 0.0191618
R13863 VSS.n1595 VSS.n1588 0.0191618
R13864 VSS.n1585 VSS.n1584 0.0191618
R13865 VSS.n1584 VSS.n1580 0.0191618
R13866 VSS.n1416 VSS.n1415 0.0191618
R13867 VSS.n1413 VSS.n1412 0.0191618
R13868 VSS.n1412 VSS.n1411 0.0191618
R13869 VSS.n1409 VSS.n1408 0.0191618
R13870 VSS.n1408 VSS.n1407 0.0191618
R13871 VSS.n1405 VSS.n1404 0.0191618
R13872 VSS.n619 VSS.n572 0.0191618
R13873 VSS.n619 VSS.n588 0.0191618
R13874 VSS.n585 VSS.n584 0.0191618
R13875 VSS.n584 VSS.n583 0.0191618
R13876 VSS.n580 VSS.n579 0.0191618
R13877 VSS.n579 VSS.n578 0.0191618
R13878 VSS.n575 VSS.n574 0.0191618
R13879 VSS.n574 VSS.n573 0.0191618
R13880 VSS.n449 VSS.n436 0.0191618
R13881 VSS.n449 VSS.n438 0.0191618
R13882 VSS.n1473 VSS.n1458 0.0191618
R13883 VSS.n1473 VSS.n1472 0.0191618
R13884 VSS.n1453 VSS.n1444 0.0191618
R13885 VSS.n1453 VSS.n1452 0.0191618
R13886 VSS.n1439 VSS.n452 0.0191618
R13887 VSS.n1439 VSS.n1438 0.0191618
R13888 VSS.n1435 VSS.n1434 0.0191618
R13889 VSS.n1434 VSS.n506 0.0191618
R13890 VSS.n503 VSS.n502 0.0191618
R13891 VSS.n502 VSS.n501 0.0191618
R13892 VSS.n498 VSS.n497 0.0191618
R13893 VSS.n497 VSS.n496 0.0191618
R13894 VSS.n493 VSS.n492 0.0191618
R13895 VSS.n492 VSS.n491 0.0191618
R13896 VSS.n1279 VSS.n1270 0.0190526
R13897 VSS.n1296 VSS.n1270 0.0190526
R13898 VSS VSS.n936 0.0189314
R13899 VSS.n2469 VSS.n351 0.0186413
R13900 VSS.n1160 VSS 0.0185144
R13901 VSS.n2252 VSS.n2251 0.0183481
R13902 VSS.n2251 VSS.n2221 0.0183481
R13903 VSS.n2326 VSS.n2325 0.0183481
R13904 VSS.n2327 VSS.n2326 0.0183481
R13905 VSS.n507 VSS 0.0177477
R13906 VSS VSS.n434 0.0177477
R13907 VSS VSS.n2049 0.0177477
R13908 VSS.n2459 VSS.n2458 0.0173735
R13909 VSS.n4 VSS.n1 0.0173735
R13910 VSS VSS.n85 0.0167536
R13911 VSS VSS.n2717 0.0167536
R13912 VSS.n1347 VSS.n1346 0.0164444
R13913 VSS.n776 VSS.n775 0.0156071
R13914 VSS.n771 VSS.n770 0.0156071
R13915 VSS.n2864 VSS.n0 0.0156071
R13916 VSS.n2482 VSS.n2481 0.0156071
R13917 VSS.n2500 VSS.n254 0.0156071
R13918 VSS.n2500 VSS.n255 0.0156071
R13919 VSS.n2464 VSS.n2463 0.0156071
R13920 VSS.n1372 VSS.n1371 0.0156071
R13921 VSS.n521 VSS.n520 0.0156071
R13922 VSS.n516 VSS.n510 0.0156071
R13923 VSS.n345 VSS.n344 0.0156071
R13924 VSS.n340 VSS.n339 0.0156071
R13925 VSS.n2477 VSS.n2471 0.0156071
R13926 VSS.n1927 VSS.n1926 0.0149953
R13927 VSS.n297 VSS.n296 0.0143235
R13928 VSS.n1059 VSS.n1058 0.0143235
R13929 VSS.n1054 VSS.n1053 0.0143235
R13930 VSS.n1049 VSS.n1048 0.0143235
R13931 VSS.n830 VSS.n829 0.0143235
R13932 VSS.n848 VSS.n847 0.0143235
R13933 VSS.n859 VSS.n858 0.0143235
R13934 VSS.n951 VSS.n950 0.0143235
R13935 VSS.n946 VSS.n945 0.0143235
R13936 VSS.n941 VSS.n940 0.0143235
R13937 VSS.n88 VSS.n87 0.0143235
R13938 VSS.n99 VSS.n98 0.0143235
R13939 VSS.n110 VSS.n109 0.0143235
R13940 VSS.n2713 VSS.n2712 0.0143235
R13941 VSS.n2708 VSS.n2707 0.0143235
R13942 VSS.n2703 VSS.n2702 0.0143235
R13943 VSS.n226 VSS.n225 0.0143235
R13944 VSS.n221 VSS.n220 0.0143235
R13945 VSS.n216 VSS.n215 0.0143235
R13946 VSS.n2545 VSS.n2544 0.0143235
R13947 VSS.n2540 VSS.n2539 0.0143235
R13948 VSS.n2535 VSS.n2534 0.0143235
R13949 VSS.n2152 VSS.n2151 0.0143235
R13950 VSS.n2147 VSS.n2146 0.0143235
R13951 VSS.n2142 VSS.n2141 0.0143235
R13952 VSS.n1934 VSS.n1933 0.0143235
R13953 VSS.n1952 VSS.n1951 0.0143235
R13954 VSS.n1963 VSS.n1962 0.0143235
R13955 VSS.n2045 VSS.n2044 0.0143235
R13956 VSS.n2040 VSS.n2039 0.0143235
R13957 VSS.n1871 VSS.n1870 0.0143235
R13958 VSS.n1860 VSS.n1859 0.0143235
R13959 VSS.n1849 VSS.n1848 0.0143235
R13960 VSS.n1825 VSS.n1824 0.0143235
R13961 VSS.n1737 VSS.n1736 0.0143235
R13962 VSS.n1726 VSS.n1725 0.0143235
R13963 VSS.n1716 VSS.n1715 0.0143235
R13964 VSS.n1609 VSS.n1608 0.0143235
R13965 VSS.n1598 VSS.n1597 0.0143235
R13966 VSS.n1587 VSS.n1586 0.0143235
R13967 VSS.n587 VSS.n586 0.0143235
R13968 VSS.n582 VSS.n581 0.0143235
R13969 VSS.n577 VSS.n576 0.0143235
R13970 VSS.n505 VSS.n504 0.0143235
R13971 VSS.n500 VSS.n499 0.0143235
R13972 VSS.n495 VSS.n494 0.0143235
R13973 VSS.n2504 VSS.n2503 0.0142993
R13974 VSS.n1376 VSS.n1375 0.0142993
R13975 VSS.n2618 VSS.n248 0.0138065
R13976 VSS.n768 VSS.n767 0.0137243
R13977 VSS.n514 VSS.n513 0.0137243
R13978 VSS.n337 VSS.n336 0.0137243
R13979 VSS.n2475 VSS.n2474 0.0137243
R13980 VSS.n709 VSS.n708 0.0137188
R13981 VSS.n713 VSS.n712 0.0137188
R13982 VSS.n1338 VSS.n679 0.0137188
R13983 VSS.n2256 VSS.n2255 0.0137188
R13984 VSS.n2262 VSS.n2259 0.0137188
R13985 VSS.n2262 VSS.n2261 0.0137188
R13986 VSS.n2316 VSS.n2315 0.0137188
R13987 VSS.n2320 VSS.n2319 0.0137188
R13988 VSS.n2321 VSS.n2320 0.0137188
R13989 VSS.n2330 VSS.n2324 0.0137188
R13990 VSS.n1282 VSS.n1274 0.0137188
R13991 VSS.n1294 VSS.n1293 0.0137188
R13992 VSS.n1294 VSS.n1266 0.0137188
R13993 VSS.n1332 VSS.n721 0.0135208
R13994 VSS.n2242 VSS.n2241 0.0135208
R13995 VSS.n2348 VSS.n2347 0.0135208
R13996 VSS.n1285 VSS.n1284 0.0135208
R13997 VSS.n2618 VSS 0.0133674
R13998 VSS.n1635 VSS 0.0131493
R13999 VSS.n2450 VSS.n2222 0.0130393
R14000 VSS.n1299 VSS.n1298 0.0130393
R14001 VSS.n2619 VSS.n2618 0.0128256
R14002 VSS.n1277 VSS.n1273 0.0123243
R14003 VSS.n2332 VSS.n2331 0.0123243
R14004 VSS.n2226 VSS.n2224 0.0123243
R14005 VSS.n1337 VSS.n681 0.0123243
R14006 VSS.n2502 VSS 0.0121822
R14007 VSS.n1374 VSS 0.0121822
R14008 VSS.n1499 VSS.n1498 0.0121325
R14009 VSS.n1921 VSS 0.012067
R14010 VSS.n1349 VSS.n1348 0.0116721
R14011 VSS.n734 VSS.n733 0.0115294
R14012 VSS.n740 VSS.n739 0.0115294
R14013 VSS.n746 VSS.n745 0.0115294
R14014 VSS.n283 VSS.n282 0.0115294
R14015 VSS.n301 VSS.n300 0.0115294
R14016 VSS.n322 VSS.n321 0.0115294
R14017 VSS.n240 VSS.n239 0.0115294
R14018 VSS.n2673 VSS.n2672 0.0115294
R14019 VSS.n2659 VSS.n2658 0.0115294
R14020 VSS.n1113 VSS.n1112 0.0115294
R14021 VSS.n1096 VSS.n1095 0.0115294
R14022 VSS.n1076 VSS.n1075 0.0115294
R14023 VSS.n800 VSS.n799 0.0115294
R14024 VSS.n813 VSS.n812 0.0115294
R14025 VSS.n843 VSS.n842 0.0115294
R14026 VSS.n854 VSS.n853 0.0115294
R14027 VSS.n2854 VSS.n2853 0.0115294
R14028 VSS.n2831 VSS.n2830 0.0115294
R14029 VSS.n2817 VSS.n2816 0.0115294
R14030 VSS.n793 VSS.n792 0.0115294
R14031 VSS.n1213 VSS.n1212 0.0115294
R14032 VSS.n1193 VSS.n1192 0.0115294
R14033 VSS.n1142 VSS.n1141 0.0115294
R14034 VSS.n1136 VSS.n1135 0.0115294
R14035 VSS.n49 VSS.n48 0.0115294
R14036 VSS.n129 VSS.n128 0.0115294
R14037 VSS.n142 VSS.n141 0.0115294
R14038 VSS.n148 VSS.n147 0.0115294
R14039 VSS.n2526 VSS.n2525 0.0115294
R14040 VSS.n2520 VSS.n2519 0.0115294
R14041 VSS.n2514 VSS.n2513 0.0115294
R14042 VSS.n2405 VSS.n2404 0.0115294
R14043 VSS.n2399 VSS.n2398 0.0115294
R14044 VSS.n2366 VSS.n2365 0.0115294
R14045 VSS.n447 VSS.n446 0.0115294
R14046 VSS.n1469 VSS.n1468 0.0115294
R14047 VSS.n1449 VSS.n1448 0.0115294
R14048 VSS.n2138 VSS.n2137 0.0115294
R14049 VSS.n2132 VSS.n2131 0.0115294
R14050 VSS.n372 VSS.n371 0.0115294
R14051 VSS.n431 VSS.n430 0.0115294
R14052 VSS.n1947 VSS.n1946 0.0115294
R14053 VSS.n1958 VSS.n1957 0.0115294
R14054 VSS.n1640 VSS.n1639 0.0115294
R14055 VSS.n1669 VSS.n1668 0.0115294
R14056 VSS.n1683 VSS.n1682 0.0115294
R14057 VSS.n1836 VSS.n1835 0.0115294
R14058 VSS.n1820 VSS.n1819 0.0115294
R14059 VSS.n1803 VSS.n1802 0.0115294
R14060 VSS.n601 VSS.n600 0.0115294
R14061 VSS.n360 VSS.n359 0.0115294
R14062 VSS.n2208 VSS.n2207 0.0115294
R14063 VSS.n2194 VSS.n2193 0.0115294
R14064 VSS.n1513 VSS.n1512 0.0115294
R14065 VSS.n1534 VSS.n1533 0.0115294
R14066 VSS.n1548 VSS.n1547 0.0115294
R14067 VSS.n1398 VSS.n1397 0.0115294
R14068 VSS.n1392 VSS.n1391 0.0115294
R14069 VSS.n1386 VSS.n1385 0.0115294
R14070 VSS.n568 VSS.n567 0.0115294
R14071 VSS.n562 VSS.n561 0.0115294
R14072 VSS.n556 VSS.n555 0.0115294
R14073 VSS.n2591 VSS.n2590 0.0115294
R14074 VSS.n2603 VSS.n2602 0.0115294
R14075 VSS.n2555 VSS.n2554 0.0115294
R14076 VSS.n3 VSS.n2 0.0113696
R14077 VSS.n2457 VSS.n2456 0.0113696
R14078 VSS.n8 VSS.n6 0.010716
R14079 VSS.n2462 VSS.n2461 0.0107133
R14080 VSS.n788 VSS.n787 0.0104679
R14081 VSS.n2646 VSS.n2645 0.0104679
R14082 VSS.n1004 VSS.n1003 0.0104679
R14083 VSS.n876 VSS.n875 0.0104679
R14084 VSS.n1181 VSS.n1180 0.0104679
R14085 VSS.n2736 VSS.n2735 0.0104679
R14086 VSS.n165 VSS.n164 0.0104679
R14087 VSS.n2373 VSS.n2372 0.0104679
R14088 VSS.n470 VSS.n469 0.0104679
R14089 VSS.n2085 VSS.n2084 0.0104679
R14090 VSS.n1980 VSS.n1979 0.0104679
R14091 VSS.n1708 VSS.n1707 0.0104679
R14092 VSS.n1794 VSS.n1793 0.0104679
R14093 VSS.n2181 VSS.n2180 0.0103933
R14094 VSS VSS.n289 0.0102662
R14095 VSS.n1160 VSS.n1159 0.010166
R14096 VSS.n825 VSS.n798 0.0100886
R14097 VSS.n753 VSS.n752 0.00997131
R14098 VSS.n754 VSS.n753 0.00997131
R14099 VSS.n757 VSS.n756 0.00997131
R14100 VSS.n758 VSS.n757 0.00997131
R14101 VSS.n761 VSS.n760 0.00997131
R14102 VSS.n762 VSS.n761 0.00997131
R14103 VSS.n279 VSS.n278 0.00997131
R14104 VSS.n280 VSS.n279 0.00997131
R14105 VSS.n2587 VSS.n2586 0.00997131
R14106 VSS.n2588 VSS.n2587 0.00997131
R14107 VSS.n2597 VSS.n2596 0.00997131
R14108 VSS.n2598 VSS.n2597 0.00997131
R14109 VSS.n44 VSS.n43 0.00997131
R14110 VSS.n43 VSS.n42 0.00997131
R14111 VSS.n40 VSS.n39 0.00997131
R14112 VSS.n39 VSS.n38 0.00997131
R14113 VSS.n36 VSS.n35 0.00997131
R14114 VSS.n35 VSS.n34 0.00997131
R14115 VSS.n1154 VSS.n1153 0.00997131
R14116 VSS.n1153 VSS.n1152 0.00997131
R14117 VSS.n1150 VSS.n1149 0.00997131
R14118 VSS.n1149 VSS.n1148 0.00997131
R14119 VSS.n1146 VSS.n1145 0.00997131
R14120 VSS.n1145 VSS.n1144 0.00997131
R14121 VSS.n2423 VSS.n2422 0.00997131
R14122 VSS.n2422 VSS.n2421 0.00997131
R14123 VSS.n2419 VSS.n2418 0.00997131
R14124 VSS.n2418 VSS.n2417 0.00997131
R14125 VSS.n2415 VSS.n2414 0.00997131
R14126 VSS.n2414 VSS.n2413 0.00997131
R14127 VSS.n2077 VSS.n2076 0.00997131
R14128 VSS.n2076 VSS.n2075 0.00997131
R14129 VSS.n2073 VSS.n2072 0.00997131
R14130 VSS.n2072 VSS.n2071 0.00997131
R14131 VSS.n2069 VSS.n2068 0.00997131
R14132 VSS.n2068 VSS.n2067 0.00997131
R14133 VSS.n2036 VSS.n2035 0.00997131
R14134 VSS.n2035 VSS.n2034 0.00997131
R14135 VSS.n1808 VSS.n1807 0.00997131
R14136 VSS.n1807 VSS.n1806 0.00997131
R14137 VSS.n1798 VSS.n1797 0.00997131
R14138 VSS.n1797 VSS.n1796 0.00997131
R14139 VSS.n1415 VSS.n1414 0.00997131
R14140 VSS.n1414 VSS.n1413 0.00997131
R14141 VSS.n1411 VSS.n1410 0.00997131
R14142 VSS.n1410 VSS.n1409 0.00997131
R14143 VSS.n1407 VSS.n1406 0.00997131
R14144 VSS.n1406 VSS.n1405 0.00997131
R14145 VSS VSS.n1160 0.00986931
R14146 VSS.n2806 VSS.n2805 0.0098203
R14147 VSS.n276 VSS.n273 0.0098203
R14148 VSS.n912 VSS.n907 0.0098203
R14149 VSS.n1035 VSS.n1030 0.0098203
R14150 VSS.n2782 VSS.n2777 0.0098203
R14151 VSS.n196 VSS.n191 0.0098203
R14152 VSS.n84 VSS.n79 0.0098203
R14153 VSS.n2530 VSS.n2510 0.0098203
R14154 VSS.n406 VSS.n401 0.0098203
R14155 VSS.n2016 VSS.n2011 0.0098203
R14156 VSS.n1903 VSS.n1898 0.0098203
R14157 VSS.n1769 VSS.n1764 0.0098203
R14158 VSS.n1622 VSS.n1617 0.0098203
R14159 VSS.n1574 VSS.n1573 0.0098203
R14160 VSS.n1402 VSS.n1382 0.0098203
R14161 VSS.n621 VSS.n620 0.0098203
R14162 VSS.n551 VSS.n475 0.0098203
R14163 VSS.n2584 VSS.n2581 0.0098203
R14164 VSS.n1922 VSS.n1479 0.00977288
R14165 VSS.n736 VSS.n735 0.00969118
R14166 VSS.n742 VSS.n741 0.00969118
R14167 VSS.n748 VSS.n747 0.00969118
R14168 VSS.n310 VSS.n309 0.00969118
R14169 VSS.n2670 VSS.n2669 0.00969118
R14170 VSS.n2656 VSS.n2655 0.00969118
R14171 VSS.n2624 VSS.n2623 0.00969118
R14172 VSS.n1087 VSS.n1086 0.00969118
R14173 VSS.n1073 VSS.n1072 0.00969118
R14174 VSS.n988 VSS.n987 0.00969118
R14175 VSS.n1033 VSS.n1032 0.00969118
R14176 VSS.n1039 VSS.n1038 0.00969118
R14177 VSS.n1044 VSS.n1043 0.00969118
R14178 VSS.n910 VSS.n909 0.00969118
R14179 VSS.n916 VSS.n915 0.00969118
R14180 VSS.n922 VSS.n921 0.00969118
R14181 VSS.n2828 VSS.n2827 0.00969118
R14182 VSS.n2814 VSS.n2813 0.00969118
R14183 VSS.n2789 VSS.n2788 0.00969118
R14184 VSS.n2780 VSS.n2779 0.00969118
R14185 VSS.n20 VSS.n19 0.00969118
R14186 VSS.n26 VSS.n25 0.00969118
R14187 VSS.n1204 VSS.n1203 0.00969118
R14188 VSS.n1190 VSS.n1189 0.00969118
R14189 VSS.n1165 VSS.n1164 0.00969118
R14190 VSS.n1140 VSS.n1139 0.00969118
R14191 VSS.n1134 VSS.n1133 0.00969118
R14192 VSS.n51 VSS.n50 0.00969118
R14193 VSS.n82 VSS.n81 0.00969118
R14194 VSS.n93 VSS.n92 0.00969118
R14195 VSS.n104 VSS.n103 0.00969118
R14196 VSS.n194 VSS.n193 0.00969118
R14197 VSS.n200 VSS.n199 0.00969118
R14198 VSS.n206 VSS.n205 0.00969118
R14199 VSS.n2528 VSS.n2527 0.00969118
R14200 VSS.n2522 VSS.n2521 0.00969118
R14201 VSS.n2516 VSS.n2515 0.00969118
R14202 VSS.n2403 VSS.n2402 0.00969118
R14203 VSS.n2397 VSS.n2396 0.00969118
R14204 VSS.n2368 VSS.n2367 0.00969118
R14205 VSS.n1460 VSS.n1459 0.00969118
R14206 VSS.n1446 VSS.n1445 0.00969118
R14207 VSS.n454 VSS.n453 0.00969118
R14208 VSS.n2136 VSS.n2135 0.00969118
R14209 VSS.n2130 VSS.n2129 0.00969118
R14210 VSS.n374 VSS.n373 0.00969118
R14211 VSS.n404 VSS.n403 0.00969118
R14212 VSS.n410 VSS.n409 0.00969118
R14213 VSS.n416 VSS.n415 0.00969118
R14214 VSS.n2014 VSS.n2013 0.00969118
R14215 VSS.n2020 VSS.n2019 0.00969118
R14216 VSS.n2026 VSS.n2025 0.00969118
R14217 VSS.n1660 VSS.n1659 0.00969118
R14218 VSS.n1680 VSS.n1679 0.00969118
R14219 VSS.n1692 VSS.n1691 0.00969118
R14220 VSS.n1901 VSS.n1900 0.00969118
R14221 VSS.n1865 VSS.n1864 0.00969118
R14222 VSS.n1854 VSS.n1853 0.00969118
R14223 VSS.n1767 VSS.n1766 0.00969118
R14224 VSS.n1731 VSS.n1730 0.00969118
R14225 VSS.n1720 VSS.n1719 0.00969118
R14226 VSS.n2205 VSS.n2204 0.00969118
R14227 VSS.n2191 VSS.n2190 0.00969118
R14228 VSS.n2162 VSS.n2161 0.00969118
R14229 VSS.n1526 VSS.n1525 0.00969118
R14230 VSS.n1545 VSS.n1544 0.00969118
R14231 VSS.n1557 VSS.n1556 0.00969118
R14232 VSS.n1620 VSS.n1619 0.00969118
R14233 VSS.n1603 VSS.n1602 0.00969118
R14234 VSS.n1592 VSS.n1591 0.00969118
R14235 VSS.n1400 VSS.n1399 0.00969118
R14236 VSS.n1394 VSS.n1393 0.00969118
R14237 VSS.n1388 VSS.n1387 0.00969118
R14238 VSS.n570 VSS.n569 0.00969118
R14239 VSS.n564 VSS.n563 0.00969118
R14240 VSS.n558 VSS.n557 0.00969118
R14241 VSS.n473 VSS.n472 0.00969118
R14242 VSS.n479 VSS.n478 0.00969118
R14243 VSS.n485 VSS.n484 0.00969118
R14244 VSS.n2605 VSS.n2604 0.00969118
R14245 VSS.n1336 VSS.n1335 0.00961458
R14246 VSS.n2228 VSS.n2227 0.00961458
R14247 VSS.n2333 VSS.n2311 0.00961458
R14248 VSS.n1276 VSS.n1275 0.00961458
R14249 VSS.n2497 VSS 0.009375
R14250 VSS VSS.n228 0.00844366
R14251 VSS.n348 VSS.n343 0.00816304
R14252 VSS.n349 VSS.n348 0.00816304
R14253 VSS.n2486 VSS.n2485 0.00816304
R14254 VSS.n2485 VSS.n2480 0.00816304
R14255 VSS.n2446 VSS.n2445 0.00811225
R14256 VSS.n1304 VSS.n1303 0.00811225
R14257 VSS.n4 VSS.n3 0.00809436
R14258 VSS.n2459 VSS.n2457 0.00809436
R14259 VSS.n1365 VSS 0.00774506
R14260 VSS.n1120 VSS 0.00759434
R14261 VSS.n751 VSS.n750 0.0075272
R14262 VSS.n1156 VSS.n1155 0.0075272
R14263 VSS.n33 VSS.n32 0.0075272
R14264 VSS.n2424 VSS.n2412 0.0075272
R14265 VSS.n1417 VSS.n1416 0.0075272
R14266 VSS.n1404 VSS.n1403 0.0075272
R14267 VSS.n2033 VSS.n2032 0.0075272
R14268 VSS.n786 VSS.n785 0.0075272
R14269 VSS.n683 VSS.n682 0.00701042
R14270 VSS.n2305 VSS.n2304 0.00701042
R14271 VSS.n2451 VSS.n2450 0.00673148
R14272 VSS.n825 VSS 0.00672253
R14273 VSS.n825 VSS.n824 0.00659014
R14274 VSS.n1120 VSS 0.00647324
R14275 VSS.n2865 VSS.n2864 0.00635126
R14276 VSS.n2465 VSS.n2464 0.00635126
R14277 VSS.n1372 VSS.n1370 0.00635126
R14278 VSS.n2863 VSS.n2862 0.00603245
R14279 VSS.n2468 VSS.n2467 0.00591449
R14280 VSS.n720 VSS.n718 0.00570833
R14281 VSS.n1333 VSS.n1332 0.00570833
R14282 VSS.n2244 VSS.n2242 0.00570833
R14283 VSS.n2439 VSS.n2438 0.00570833
R14284 VSS.n2352 VSS.n2350 0.00570833
R14285 VSS.n2347 VSS.n2334 0.00570833
R14286 VSS.n1285 VSS.n1272 0.00570833
R14287 VSS.n1308 VSS.n1264 0.00570833
R14288 VSS.n1422 VSS.n508 0.0055592
R14289 VSS.n589 VSS.n435 0.00531433
R14290 VSS.n2499 VSS.n333 0.00523154
R14291 VSS.n2499 VSS.n2498 0.00523154
R14292 VSS.n618 VSS.n607 0.00523154
R14293 VSS.n618 VSS.n617 0.00523154
R14294 VSS.n616 VSS.n615 0.00523154
R14295 VSS.n615 VSS.n614 0.00523154
R14296 VSS.n613 VSS.n612 0.00523154
R14297 VSS.n612 VSS.n611 0.00523154
R14298 VSS.n610 VSS.n609 0.00523154
R14299 VSS.n609 VSS.n608 0.00523154
R14300 VSS.n590 VSS.n589 0.00523154
R14301 VSS.n591 VSS.n590 0.00523154
R14302 VSS.n593 VSS.n592 0.00523154
R14303 VSS.n594 VSS.n593 0.00523154
R14304 VSS.n596 VSS.n595 0.00523154
R14305 VSS.n597 VSS.n596 0.00523154
R14306 VSS.n605 VSS.n598 0.00523154
R14307 VSS.n606 VSS.n605 0.00523154
R14308 VSS.n1651 VSS.n1636 0.00523154
R14309 VSS.n1672 VSS.n1654 0.00523154
R14310 VSS.n1673 VSS.n1672 0.00523154
R14311 VSS.n1686 VSS.n1674 0.00523154
R14312 VSS.n1687 VSS.n1686 0.00523154
R14313 VSS.n1690 VSS.n1688 0.00523154
R14314 VSS.n1690 VSS.n1689 0.00523154
R14315 VSS.n1905 VSS.n1480 0.00523154
R14316 VSS.n1906 VSS.n1905 0.00523154
R14317 VSS.n1908 VSS.n1907 0.00523154
R14318 VSS.n1909 VSS.n1908 0.00523154
R14319 VSS.n1911 VSS.n1910 0.00523154
R14320 VSS.n1912 VSS.n1911 0.00523154
R14321 VSS.n1914 VSS.n1913 0.00523154
R14322 VSS.n1915 VSS.n1914 0.00523154
R14323 VSS.n1917 VSS.n1916 0.00523154
R14324 VSS.n1918 VSS.n1917 0.00523154
R14325 VSS.n1920 VSS.n1919 0.00523154
R14326 VSS.n1518 VSS.n1503 0.00523154
R14327 VSS.n1519 VSS.n1518 0.00523154
R14328 VSS.n1537 VSS.n1520 0.00523154
R14329 VSS.n1538 VSS.n1537 0.00523154
R14330 VSS.n1551 VSS.n1539 0.00523154
R14331 VSS.n1552 VSS.n1551 0.00523154
R14332 VSS.n1555 VSS.n1553 0.00523154
R14333 VSS.n1555 VSS.n1554 0.00523154
R14334 VSS.n1624 VSS.n1500 0.00523154
R14335 VSS.n1625 VSS.n1624 0.00523154
R14336 VSS.n1627 VSS.n1626 0.00523154
R14337 VSS.n1628 VSS.n1627 0.00523154
R14338 VSS.n1630 VSS.n1629 0.00523154
R14339 VSS.n1631 VSS.n1630 0.00523154
R14340 VSS.n1633 VSS.n1632 0.00523154
R14341 VSS.n1634 VSS.n1633 0.00523154
R14342 VSS.n966 VSS.n965 0.00521572
R14343 VSS.n964 VSS.n963 0.00521572
R14344 VSS.n963 VSS.n962 0.00521572
R14345 VSS.n961 VSS.n960 0.00521572
R14346 VSS.n960 VSS.n959 0.00521572
R14347 VSS.n958 VSS.n957 0.00521572
R14348 VSS.n957 VSS.n956 0.00521572
R14349 VSS.n955 VSS.n954 0.00521572
R14350 VSS.n954 VSS.n828 0.00521572
R14351 VSS.n929 VSS.n928 0.00521572
R14352 VSS.n930 VSS.n929 0.00521572
R14353 VSS.n932 VSS.n931 0.00521572
R14354 VSS.n933 VSS.n932 0.00521572
R14355 VSS.n935 VSS.n934 0.00521572
R14356 VSS.n2860 VSS.n2859 0.00521572
R14357 VSS.n2859 VSS.n2844 0.00521572
R14358 VSS.n2843 VSS.n2842 0.00521572
R14359 VSS.n2842 VSS.n2824 0.00521572
R14360 VSS.n2823 VSS.n2822 0.00521572
R14361 VSS.n2822 VSS.n2810 0.00521572
R14362 VSS.n2809 VSS.n2808 0.00521572
R14363 VSS.n2808 VSS.n10 0.00521572
R14364 VSS.n1119 VSS.n1118 0.00521572
R14365 VSS.n1118 VSS.n1103 0.00521572
R14366 VSS.n1102 VSS.n1101 0.00521572
R14367 VSS.n1101 VSS.n1083 0.00521572
R14368 VSS.n1082 VSS.n1081 0.00521572
R14369 VSS.n1081 VSS.n1069 0.00521572
R14370 VSS.n1068 VSS.n1067 0.00521572
R14371 VSS.n1067 VSS.n984 0.00521572
R14372 VSS.n983 VSS.n982 0.00521572
R14373 VSS.n982 VSS.n981 0.00521572
R14374 VSS.n980 VSS.n979 0.00521572
R14375 VSS.n979 VSS.n978 0.00521572
R14376 VSS.n977 VSS.n976 0.00521572
R14377 VSS.n976 VSS.n975 0.00521572
R14378 VSS.n974 VSS.n973 0.00521572
R14379 VSS.n973 VSS.n798 0.00521572
R14380 VSS.n316 VSS.n256 0.00521572
R14381 VSS.n317 VSS.n316 0.00521572
R14382 VSS.n331 VSS.n318 0.00521572
R14383 VSS.n332 VSS.n331 0.00521572
R14384 VSS.n525 VSS.n524 0.00499045
R14385 VSS.n524 VSS.n519 0.00499045
R14386 VSS VSS.n351 0.00496556
R14387 VSS.n779 VSS.n774 0.00493396
R14388 VSS.n780 VSS.n779 0.00493396
R14389 VSS.n1278 VSS.n1274 0.00490287
R14390 VSS.n708 VSS.n697 0.00489761
R14391 VSS.n772 VSS.n771 0.00489326
R14392 VSS.n517 VSS.n516 0.00489326
R14393 VSS.n341 VSS.n340 0.00489326
R14394 VSS.n2478 VSS.n2477 0.00489326
R14395 VSS.n1924 VSS.n1923 0.00489252
R14396 VSS.n2220 VSS.n2219 0.00481193
R14397 VSS.n2219 VSS.n2218 0.00481193
R14398 VSS.n2217 VSS.n2216 0.00481193
R14399 VSS.n2216 VSS.n2199 0.00481193
R14400 VSS.n2198 VSS.n2197 0.00481193
R14401 VSS.n2197 VSS.n2185 0.00481193
R14402 VSS.n2184 VSS.n2183 0.00481193
R14403 VSS.n2183 VSS.n2157 0.00481193
R14404 VSS.n1478 VSS.n1477 0.00481193
R14405 VSS.n1477 VSS.n1476 0.00481193
R14406 VSS.n1475 VSS.n1474 0.00481193
R14407 VSS.n1474 VSS.n1456 0.00481193
R14408 VSS.n1455 VSS.n1454 0.00481193
R14409 VSS.n1454 VSS.n1442 0.00481193
R14410 VSS.n1441 VSS.n1440 0.00481193
R14411 VSS.n1440 VSS.n450 0.00481193
R14412 VSS.n1433 VSS.n507 0.00481193
R14413 VSS.n1433 VSS.n1432 0.00481193
R14414 VSS.n1431 VSS.n1430 0.00481193
R14415 VSS.n1430 VSS.n1429 0.00481193
R14416 VSS.n1428 VSS.n1427 0.00481193
R14417 VSS.n1427 VSS.n1426 0.00481193
R14418 VSS.n1425 VSS.n1424 0.00481193
R14419 VSS.n1424 VSS.n1423 0.00481193
R14420 VSS.n1484 VSS.n1483 0.00481193
R14421 VSS.n2060 VSS.n434 0.00481193
R14422 VSS.n2060 VSS.n2059 0.00481193
R14423 VSS.n2058 VSS.n2057 0.00481193
R14424 VSS.n2057 VSS.n2056 0.00481193
R14425 VSS.n2055 VSS.n2054 0.00481193
R14426 VSS.n2054 VSS.n2053 0.00481193
R14427 VSS.n2052 VSS.n2051 0.00481193
R14428 VSS.n2051 VSS.n2050 0.00481193
R14429 VSS.n2049 VSS.n2048 0.00481193
R14430 VSS.n2048 VSS.n1932 0.00481193
R14431 VSS.n1931 VSS.n1930 0.00481193
R14432 VSS.n1930 VSS.n1929 0.00481193
R14433 VSS.n2156 VSS.n2155 0.00481193
R14434 VSS.n2155 VSS.n365 0.00481193
R14435 VSS.n1486 VSS.n1485 0.00481193
R14436 VSS.n1487 VSS.n1486 0.00481193
R14437 VSS.n1489 VSS.n1488 0.00481193
R14438 VSS.n1490 VSS.n1489 0.00481193
R14439 VSS.n1492 VSS.n1491 0.00481193
R14440 VSS.n1493 VSS.n1492 0.00481193
R14441 VSS.n2861 VSS 0.00463641
R14442 VSS.n1653 VSS.n1652 0.00460067
R14443 VSS.n1926 VSS.n1925 0.00459245
R14444 VSS.n1221 VSS.n9 0.0045634
R14445 VSS.n1221 VSS.n1220 0.0045634
R14446 VSS.n1219 VSS.n1218 0.0045634
R14447 VSS.n1218 VSS.n1200 0.0045634
R14448 VSS.n1199 VSS.n1198 0.0045634
R14449 VSS.n1198 VSS.n1186 0.0045634
R14450 VSS.n1185 VSS.n1184 0.0045634
R14451 VSS.n1184 VSS.n1161 0.0045634
R14452 VSS.n2728 VSS.n85 0.0045634
R14453 VSS.n2728 VSS.n2727 0.0045634
R14454 VSS.n2726 VSS.n2725 0.0045634
R14455 VSS.n2725 VSS.n2724 0.0045634
R14456 VSS.n2723 VSS.n2722 0.0045634
R14457 VSS.n2722 VSS.n2721 0.0045634
R14458 VSS.n2720 VSS.n2719 0.0045634
R14459 VSS.n2719 VSS.n2718 0.0045634
R14460 VSS.n2717 VSS.n2716 0.0045634
R14461 VSS.n2716 VSS.n86 0.0045634
R14462 VSS.n816 VSS.n815 0.0045634
R14463 VSS.n2691 VSS.n2690 0.0045634
R14464 VSS.n2690 VSS.n2689 0.0045634
R14465 VSS.n2688 VSS.n2687 0.0045634
R14466 VSS.n2687 VSS.n2686 0.0045634
R14467 VSS.n2685 VSS.n2684 0.0045634
R14468 VSS.n2684 VSS.n2683 0.0045634
R14469 VSS.n2682 VSS.n2681 0.0045634
R14470 VSS.n2681 VSS.n2680 0.0045634
R14471 VSS.n2679 VSS.n2678 0.0045634
R14472 VSS.n2678 VSS.n2666 0.0045634
R14473 VSS.n2665 VSS.n2664 0.0045634
R14474 VSS.n2664 VSS.n2652 0.0045634
R14475 VSS.n2651 VSS.n2650 0.0045634
R14476 VSS.n2549 VSS.n2548 0.0045634
R14477 VSS.n2548 VSS.n249 0.0045634
R14478 VSS.n2489 VSS.n2488 0.0045634
R14479 VSS.n2490 VSS.n2489 0.0045634
R14480 VSS.n2492 VSS.n2491 0.0045634
R14481 VSS.n2493 VSS.n2492 0.0045634
R14482 VSS.n2495 VSS.n2494 0.0045634
R14483 VSS.n2496 VSS.n2495 0.0045634
R14484 VSS.n2617 VSS.n2565 0.0045634
R14485 VSS.n2564 VSS.n2563 0.0045634
R14486 VSS.n2563 VSS.n2550 0.0045634
R14487 VSS.n2255 VSS.n2254 0.00451955
R14488 VSS.n2330 VSS.n2329 0.00451955
R14489 VSS.n721 VSS.n720 0.00440625
R14490 VSS.n2241 VSS.n2223 0.00440625
R14491 VSS.n2246 VSS.n2244 0.00440625
R14492 VSS.n2350 VSS.n2348 0.00440625
R14493 VSS.n1284 VSS.n1256 0.00440625
R14494 VSS.n1290 VSS.n1272 0.00440625
R14495 VSS.n1921 VSS.n1920 0.00428523
R14496 VSS.n1301 VSS.n1269 0.0042807
R14497 VSS.n1339 VSS.n1338 0.00427564
R14498 VSS.n248 VSS.n247 0.00410644
R14499 VSS.n245 VSS.n244 0.00410644
R14500 VSS.n293 VSS.n287 0.00410644
R14501 VSS VSS.n509 0.00409203
R14502 VSS.n817 VSS.n816 0.00402161
R14503 VSS.n1498 VSS.n1497 0.00401501
R14504 VSS.n617 VSS.n616 0.00365436
R14505 VSS.n614 VSS.n613 0.00365436
R14506 VSS.n611 VSS.n610 0.00365436
R14507 VSS.n592 VSS.n591 0.00365436
R14508 VSS.n595 VSS.n594 0.00365436
R14509 VSS.n598 VSS.n597 0.00365436
R14510 VSS.n1654 VSS.n1653 0.00365436
R14511 VSS.n1674 VSS.n1673 0.00365436
R14512 VSS.n1688 VSS.n1687 0.00365436
R14513 VSS.n1907 VSS.n1906 0.00365436
R14514 VSS.n1910 VSS.n1909 0.00365436
R14515 VSS.n1913 VSS.n1912 0.00365436
R14516 VSS.n1919 VSS.n1918 0.00365436
R14517 VSS.n1520 VSS.n1519 0.00365436
R14518 VSS.n1539 VSS.n1538 0.00365436
R14519 VSS.n1553 VSS.n1552 0.00365436
R14520 VSS.n1626 VSS.n1625 0.00365436
R14521 VSS.n1629 VSS.n1628 0.00365436
R14522 VSS.n1632 VSS.n1631 0.00365436
R14523 VSS.n966 VSS.n827 0.00364381
R14524 VSS.n965 VSS.n964 0.00364381
R14525 VSS.n962 VSS.n961 0.00364381
R14526 VSS.n959 VSS.n958 0.00364381
R14527 VSS.n928 VSS.n828 0.00364381
R14528 VSS.n931 VSS.n930 0.00364381
R14529 VSS.n934 VSS.n933 0.00364381
R14530 VSS.n2844 VSS.n2843 0.00364381
R14531 VSS.n2824 VSS.n2823 0.00364381
R14532 VSS.n2810 VSS.n2809 0.00364381
R14533 VSS.n1103 VSS.n1102 0.00364381
R14534 VSS.n1083 VSS.n1082 0.00364381
R14535 VSS.n1069 VSS.n1068 0.00364381
R14536 VSS.n981 VSS.n980 0.00364381
R14537 VSS.n978 VSS.n977 0.00364381
R14538 VSS.n975 VSS.n974 0.00364381
R14539 VSS.n288 VSS.n256 0.00364381
R14540 VSS.n318 VSS.n317 0.00364381
R14541 VSS.n2315 VSS.n2314 0.00362372
R14542 VSS.n1298 VSS.n1269 0.00360776
R14543 VSS.n291 VSS.n290 0.00343981
R14544 VSS.n14 VSS.n13 0.0034393
R14545 VSS.n1159 VSS.n1158 0.0034393
R14546 VSS.n2218 VSS.n2217 0.00337462
R14547 VSS.n2199 VSS.n2198 0.00337462
R14548 VSS.n2185 VSS.n2184 0.00337462
R14549 VSS.n1476 VSS.n1475 0.00337462
R14550 VSS.n1456 VSS.n1455 0.00337462
R14551 VSS.n1442 VSS.n1441 0.00337462
R14552 VSS.n1432 VSS.n1431 0.00337462
R14553 VSS.n1429 VSS.n1428 0.00337462
R14554 VSS.n1426 VSS.n1425 0.00337462
R14555 VSS.n2059 VSS.n2058 0.00337462
R14556 VSS.n2056 VSS.n2055 0.00337462
R14557 VSS.n2053 VSS.n2052 0.00337462
R14558 VSS.n1932 VSS.n1931 0.00337462
R14559 VSS.n1929 VSS.n1928 0.00337462
R14560 VSS.n1485 VSS.n365 0.00337462
R14561 VSS.n1488 VSS.n1487 0.00337462
R14562 VSS.n1491 VSS.n1490 0.00337462
R14563 VSS.n1495 VSS.n1494 0.00334838
R14564 VSS.n1362 VSS.n1361 0.00324725
R14565 VSS.n1220 VSS.n1219 0.00320893
R14566 VSS.n1200 VSS.n1199 0.00320893
R14567 VSS.n1186 VSS.n1185 0.00320893
R14568 VSS.n2727 VSS.n2726 0.00320893
R14569 VSS.n2724 VSS.n2723 0.00320893
R14570 VSS.n2721 VSS.n2720 0.00320893
R14571 VSS.n815 VSS.n86 0.00320893
R14572 VSS.n2692 VSS.n2691 0.00320893
R14573 VSS.n2689 VSS.n2688 0.00320893
R14574 VSS.n2686 VSS.n2685 0.00320893
R14575 VSS.n2680 VSS.n2679 0.00320893
R14576 VSS.n2666 VSS.n2665 0.00320893
R14577 VSS.n2652 VSS.n2651 0.00320893
R14578 VSS.n2488 VSS.n249 0.00320893
R14579 VSS.n2491 VSS.n2490 0.00320893
R14580 VSS.n2494 VSS.n2493 0.00320893
R14581 VSS.n2618 VSS.n2617 0.00320893
R14582 VSS.n2565 VSS.n2564 0.00320893
R14583 VSS.n1776 VSS.n1775 0.00319485
R14584 VSS.n1777 VSS.n1776 0.00319485
R14585 VSS.n2693 VSS.n2692 0.00307349
R14586 VSS.n2650 VSS.n2620 0.00307349
R14587 VSS.n1925 VSS.n1924 0.00279583
R14588 VSS.n797 VSS.n16 0.00277266
R14589 VSS.n1122 VSS.n1121 0.00277266
R14590 VSS.n783 VSS.n782 0.00270045
R14591 VSS.n1499 VSS 0.00265596
R14592 VSS.n296 VSS.n295 0.00257353
R14593 VSS.n298 VSS.n297 0.00257353
R14594 VSS.n314 VSS.n313 0.00257353
R14595 VSS.n320 VSS.n319 0.00257353
R14596 VSS.n231 VSS.n230 0.00257353
R14597 VSS.n2668 VSS.n2667 0.00257353
R14598 VSS.n2676 VSS.n2675 0.00257353
R14599 VSS.n2654 VSS.n2653 0.00257353
R14600 VSS.n2662 VSS.n2661 0.00257353
R14601 VSS.n2622 VSS.n2621 0.00257353
R14602 VSS.n2648 VSS.n2647 0.00257353
R14603 VSS.n2567 VSS.n2566 0.00257353
R14604 VSS.n2600 VSS.n2599 0.00257353
R14605 VSS.n2552 VSS.n2551 0.00257353
R14606 VSS.n1116 VSS.n1115 0.00257353
R14607 VSS.n1085 VSS.n1084 0.00257353
R14608 VSS.n1099 VSS.n1098 0.00257353
R14609 VSS.n1071 VSS.n1070 0.00257353
R14610 VSS.n1079 VSS.n1078 0.00257353
R14611 VSS.n986 VSS.n985 0.00257353
R14612 VSS.n1065 VSS.n1064 0.00257353
R14613 VSS.n1063 VSS.n1062 0.00257353
R14614 VSS.n1060 VSS.n1059 0.00257353
R14615 VSS.n1058 VSS.n1057 0.00257353
R14616 VSS.n1055 VSS.n1054 0.00257353
R14617 VSS.n1053 VSS.n1052 0.00257353
R14618 VSS.n1050 VSS.n1049 0.00257353
R14619 VSS.n1048 VSS.n1047 0.00257353
R14620 VSS.n971 VSS.n970 0.00257353
R14621 VSS.n969 VSS.n968 0.00257353
R14622 VSS.n829 VSS.n803 0.00257353
R14623 VSS.n831 VSS.n830 0.00257353
R14624 VSS.n847 VSS.n846 0.00257353
R14625 VSS.n849 VSS.n848 0.00257353
R14626 VSS.n858 VSS.n857 0.00257353
R14627 VSS.n860 VSS.n859 0.00257353
R14628 VSS.n879 VSS.n878 0.00257353
R14629 VSS.n881 VSS.n880 0.00257353
R14630 VSS.n952 VSS.n951 0.00257353
R14631 VSS.n950 VSS.n949 0.00257353
R14632 VSS.n947 VSS.n946 0.00257353
R14633 VSS.n945 VSS.n944 0.00257353
R14634 VSS.n942 VSS.n941 0.00257353
R14635 VSS.n940 VSS.n939 0.00257353
R14636 VSS.n2857 VSS.n2856 0.00257353
R14637 VSS.n2826 VSS.n2825 0.00257353
R14638 VSS.n2840 VSS.n2839 0.00257353
R14639 VSS.n2812 VSS.n2811 0.00257353
R14640 VSS.n2820 VSS.n2819 0.00257353
R14641 VSS.n12 VSS.n11 0.00257353
R14642 VSS.n2787 VSS.n2786 0.00257353
R14643 VSS.n2785 VSS.n2784 0.00257353
R14644 VSS.n796 VSS.n795 0.00257353
R14645 VSS.n1202 VSS.n1201 0.00257353
R14646 VSS.n1216 VSS.n1215 0.00257353
R14647 VSS.n1188 VSS.n1187 0.00257353
R14648 VSS.n1196 VSS.n1195 0.00257353
R14649 VSS.n1163 VSS.n1162 0.00257353
R14650 VSS.n2733 VSS.n2732 0.00257353
R14651 VSS.n2731 VSS.n2730 0.00257353
R14652 VSS.n87 VSS.n53 0.00257353
R14653 VSS.n89 VSS.n88 0.00257353
R14654 VSS.n98 VSS.n97 0.00257353
R14655 VSS.n100 VSS.n99 0.00257353
R14656 VSS.n109 VSS.n108 0.00257353
R14657 VSS.n111 VSS.n110 0.00257353
R14658 VSS.n117 VSS.n116 0.00257353
R14659 VSS.n119 VSS.n118 0.00257353
R14660 VSS.n2714 VSS.n2713 0.00257353
R14661 VSS.n2712 VSS.n2711 0.00257353
R14662 VSS.n2709 VSS.n2708 0.00257353
R14663 VSS.n2707 VSS.n2706 0.00257353
R14664 VSS.n2704 VSS.n2703 0.00257353
R14665 VSS.n2702 VSS.n2701 0.00257353
R14666 VSS.n2699 VSS.n2698 0.00257353
R14667 VSS.n2697 VSS.n2696 0.00257353
R14668 VSS.n227 VSS.n226 0.00257353
R14669 VSS.n225 VSS.n224 0.00257353
R14670 VSS.n222 VSS.n221 0.00257353
R14671 VSS.n220 VSS.n219 0.00257353
R14672 VSS.n217 VSS.n216 0.00257353
R14673 VSS.n215 VSS.n214 0.00257353
R14674 VSS.n2546 VSS.n2545 0.00257353
R14675 VSS.n2544 VSS.n2543 0.00257353
R14676 VSS.n2541 VSS.n2540 0.00257353
R14677 VSS.n2539 VSS.n2538 0.00257353
R14678 VSS.n2536 VSS.n2535 0.00257353
R14679 VSS.n2534 VSS.n2533 0.00257353
R14680 VSS.n2153 VSS.n2152 0.00257353
R14681 VSS.n2151 VSS.n2150 0.00257353
R14682 VSS.n2148 VSS.n2147 0.00257353
R14683 VSS.n2146 VSS.n2145 0.00257353
R14684 VSS.n2143 VSS.n2142 0.00257353
R14685 VSS.n2141 VSS.n2140 0.00257353
R14686 VSS.n2082 VSS.n2081 0.00257353
R14687 VSS.n2080 VSS.n2079 0.00257353
R14688 VSS.n2065 VSS.n2064 0.00257353
R14689 VSS.n2063 VSS.n2062 0.00257353
R14690 VSS.n1933 VSS.n433 0.00257353
R14691 VSS.n1935 VSS.n1934 0.00257353
R14692 VSS.n1951 VSS.n1950 0.00257353
R14693 VSS.n1953 VSS.n1952 0.00257353
R14694 VSS.n1962 VSS.n1961 0.00257353
R14695 VSS.n1964 VSS.n1963 0.00257353
R14696 VSS.n1983 VSS.n1982 0.00257353
R14697 VSS.n1985 VSS.n1984 0.00257353
R14698 VSS.n2046 VSS.n2045 0.00257353
R14699 VSS.n2044 VSS.n2043 0.00257353
R14700 VSS.n2041 VSS.n2040 0.00257353
R14701 VSS.n2039 VSS.n2038 0.00257353
R14702 VSS.n1649 VSS.n1648 0.00257353
R14703 VSS.n1656 VSS.n1655 0.00257353
R14704 VSS.n1658 VSS.n1657 0.00257353
R14705 VSS.n1676 VSS.n1675 0.00257353
R14706 VSS.n1678 VSS.n1677 0.00257353
R14707 VSS.n1482 VSS.n1481 0.00257353
R14708 VSS.n1711 VSS.n1710 0.00257353
R14709 VSS.n1713 VSS.n1712 0.00257353
R14710 VSS.n1872 VSS.n1871 0.00257353
R14711 VSS.n1870 VSS.n1869 0.00257353
R14712 VSS.n1861 VSS.n1860 0.00257353
R14713 VSS.n1859 VSS.n1858 0.00257353
R14714 VSS.n1850 VSS.n1849 0.00257353
R14715 VSS.n1848 VSS.n1847 0.00257353
R14716 VSS.n1842 VSS.n1841 0.00257353
R14717 VSS.n1840 VSS.n1839 0.00257353
R14718 VSS.n1826 VSS.n1825 0.00257353
R14719 VSS.n1824 VSS.n1823 0.00257353
R14720 VSS.n1774 VSS.n1773 0.00257353
R14721 VSS.n1772 VSS.n1771 0.00257353
R14722 VSS.n1738 VSS.n1737 0.00257353
R14723 VSS.n1736 VSS.n1735 0.00257353
R14724 VSS.n1727 VSS.n1726 0.00257353
R14725 VSS.n1725 VSS.n1724 0.00257353
R14726 VSS.n1717 VSS.n1716 0.00257353
R14727 VSS.n1715 VSS.n1714 0.00257353
R14728 VSS.n363 VSS.n362 0.00257353
R14729 VSS.n2201 VSS.n2200 0.00257353
R14730 VSS.n2203 VSS.n2202 0.00257353
R14731 VSS.n2187 VSS.n2186 0.00257353
R14732 VSS.n2189 VSS.n2188 0.00257353
R14733 VSS.n2159 VSS.n2158 0.00257353
R14734 VSS.n1516 VSS.n1515 0.00257353
R14735 VSS.n1522 VSS.n1521 0.00257353
R14736 VSS.n1524 VSS.n1523 0.00257353
R14737 VSS.n1541 VSS.n1540 0.00257353
R14738 VSS.n1543 VSS.n1542 0.00257353
R14739 VSS.n1502 VSS.n1501 0.00257353
R14740 VSS.n1577 VSS.n1576 0.00257353
R14741 VSS.n1579 VSS.n1578 0.00257353
R14742 VSS.n1610 VSS.n1609 0.00257353
R14743 VSS.n1608 VSS.n1607 0.00257353
R14744 VSS.n1599 VSS.n1598 0.00257353
R14745 VSS.n1597 VSS.n1596 0.00257353
R14746 VSS.n1588 VSS.n1587 0.00257353
R14747 VSS.n1586 VSS.n1585 0.00257353
R14748 VSS.n588 VSS.n587 0.00257353
R14749 VSS.n586 VSS.n585 0.00257353
R14750 VSS.n583 VSS.n582 0.00257353
R14751 VSS.n581 VSS.n580 0.00257353
R14752 VSS.n578 VSS.n577 0.00257353
R14753 VSS.n576 VSS.n575 0.00257353
R14754 VSS.n438 VSS.n437 0.00257353
R14755 VSS.n1458 VSS.n1457 0.00257353
R14756 VSS.n1472 VSS.n1471 0.00257353
R14757 VSS.n1444 VSS.n1443 0.00257353
R14758 VSS.n1452 VSS.n1451 0.00257353
R14759 VSS.n452 VSS.n451 0.00257353
R14760 VSS.n1438 VSS.n1437 0.00257353
R14761 VSS.n1436 VSS.n1435 0.00257353
R14762 VSS.n506 VSS.n505 0.00257353
R14763 VSS.n504 VSS.n503 0.00257353
R14764 VSS.n501 VSS.n500 0.00257353
R14765 VSS.n499 VSS.n498 0.00257353
R14766 VSS.n496 VSS.n495 0.00257353
R14767 VSS.n494 VSS.n493 0.00257353
R14768 VSS.n293 VSS.n292 0.00255288
R14769 VSS.n246 VSS.n245 0.00255288
R14770 VSS.n247 VSS.n246 0.00255288
R14771 VSS.n1497 VSS.n1496 0.00250717
R14772 VSS.n820 VSS.n819 0.00248592
R14773 VSS.n823 VSS.n822 0.00248592
R14774 VSS.n824 VSS.n823 0.00248592
R14775 VSS.n2694 VSS.n228 0.00248592
R14776 VSS.n821 VSS.n820 0.00248592
R14777 VSS.n1363 VSS.n1350 0.00244755
R14778 VSS.n936 VSS.n935 0.00238629
R14779 VSS.n1248 VSS.n1247 0.00233824
R14780 VSS.n1244 VSS.n1243 0.00233824
R14781 VSS.n1240 VSS.n1236 0.00233824
R14782 VSS.n738 VSS.n737 0.00233824
R14783 VSS.n744 VSS.n743 0.00233824
R14784 VSS.n787 VSS.n749 0.00233824
R14785 VSS.n2573 VSS.n2572 0.00233824
R14786 VSS.n2614 VSS.n2613 0.00233824
R14787 VSS.n2560 VSS.n2559 0.00233824
R14788 VSS.n266 VSS.n265 0.00233824
R14789 VSS.n308 VSS.n307 0.00233824
R14790 VSS.n326 VSS.n325 0.00233824
R14791 VSS.n276 VSS.n275 0.00233824
R14792 VSS.n286 VSS.n285 0.00233824
R14793 VSS.n312 VSS.n311 0.00233824
R14794 VSS.n238 VSS.n236 0.00233824
R14795 VSS.n2631 VSS.n2630 0.00233824
R14796 VSS.n2638 VSS.n2637 0.00233824
R14797 VSS.n2674 VSS.n2671 0.00233824
R14798 VSS.n2660 VSS.n2657 0.00233824
R14799 VSS.n2646 VSS.n2625 0.00233824
R14800 VSS.n1111 VSS.n1109 0.00233824
R14801 VSS.n1094 VSS.n1093 0.00233824
R14802 VSS.n996 VSS.n995 0.00233824
R14803 VSS.n1097 VSS.n1088 0.00233824
R14804 VSS.n1077 VSS.n1074 0.00233824
R14805 VSS.n1004 VSS.n989 0.00233824
R14806 VSS.n1023 VSS.n1022 0.00233824
R14807 VSS.n1019 VSS.n1018 0.00233824
R14808 VSS.n1012 VSS.n1011 0.00233824
R14809 VSS.n1035 VSS.n1034 0.00233824
R14810 VSS.n1041 VSS.n1040 0.00233824
R14811 VSS.n1046 VSS.n1045 0.00233824
R14812 VSS.n810 VSS.n808 0.00233824
R14813 VSS.n840 VSS.n838 0.00233824
R14814 VSS.n868 VSS.n867 0.00233824
R14815 VSS.n844 VSS.n833 0.00233824
R14816 VSS.n855 VSS.n851 0.00233824
R14817 VSS.n876 VSS.n862 0.00233824
R14818 VSS.n900 VSS.n899 0.00233824
R14819 VSS.n896 VSS.n895 0.00233824
R14820 VSS.n889 VSS.n888 0.00233824
R14821 VSS.n912 VSS.n911 0.00233824
R14822 VSS.n918 VSS.n917 0.00233824
R14823 VSS.n924 VSS.n923 0.00233824
R14824 VSS.n2852 VSS.n2850 0.00233824
R14825 VSS.n2837 VSS.n2836 0.00233824
R14826 VSS.n2797 VSS.n2796 0.00233824
R14827 VSS.n2838 VSS.n2829 0.00233824
R14828 VSS.n2818 VSS.n2815 0.00233824
R14829 VSS.n2806 VSS.n2790 0.00233824
R14830 VSS.n2770 VSS.n2769 0.00233824
R14831 VSS.n2766 VSS.n2765 0.00233824
R14832 VSS.n2752 VSS.n2751 0.00233824
R14833 VSS.n2782 VSS.n2781 0.00233824
R14834 VSS.n22 VSS.n21 0.00233824
R14835 VSS.n28 VSS.n27 0.00233824
R14836 VSS.n1225 VSS.n1224 0.00233824
R14837 VSS.n1211 VSS.n1210 0.00233824
R14838 VSS.n1173 VSS.n1172 0.00233824
R14839 VSS.n1214 VSS.n1205 0.00233824
R14840 VSS.n1194 VSS.n1191 0.00233824
R14841 VSS.n1181 VSS.n1166 0.00233824
R14842 VSS.n1132 VSS.n1129 0.00233824
R14843 VSS.n2758 VSS.n2757 0.00233824
R14844 VSS.n2744 VSS.n2743 0.00233824
R14845 VSS.n1138 VSS.n1137 0.00233824
R14846 VSS.n47 VSS.n46 0.00233824
R14847 VSS.n2735 VSS.n52 0.00233824
R14848 VSS.n72 VSS.n71 0.00233824
R14849 VSS.n68 VSS.n67 0.00233824
R14850 VSS.n61 VSS.n60 0.00233824
R14851 VSS.n84 VSS.n83 0.00233824
R14852 VSS.n95 VSS.n94 0.00233824
R14853 VSS.n106 VSS.n105 0.00233824
R14854 VSS.n126 VSS.n124 0.00233824
R14855 VSS.n139 VSS.n137 0.00233824
R14856 VSS.n157 VSS.n156 0.00233824
R14857 VSS.n143 VSS.n132 0.00233824
R14858 VSS.n149 VSS.n145 0.00233824
R14859 VSS.n165 VSS.n151 0.00233824
R14860 VSS.n184 VSS.n183 0.00233824
R14861 VSS.n180 VSS.n179 0.00233824
R14862 VSS.n173 VSS.n172 0.00233824
R14863 VSS.n196 VSS.n195 0.00233824
R14864 VSS.n202 VSS.n201 0.00233824
R14865 VSS.n208 VSS.n207 0.00233824
R14866 VSS.n2276 VSS.n2272 0.00233824
R14867 VSS.n2283 VSS.n2279 0.00233824
R14868 VSS.n2287 VSS.n2286 0.00233824
R14869 VSS.n2530 VSS.n2529 0.00233824
R14870 VSS.n2524 VSS.n2523 0.00233824
R14871 VSS.n2518 VSS.n2517 0.00233824
R14872 VSS.n2427 VSS.n2426 0.00233824
R14873 VSS.n2392 VSS.n2388 0.00233824
R14874 VSS.n2385 VSS.n2381 0.00233824
R14875 VSS.n2401 VSS.n2400 0.00233824
R14876 VSS.n2364 VSS.n2363 0.00233824
R14877 VSS.n2372 VSS.n2369 0.00233824
R14878 VSS.n445 VSS.n443 0.00233824
R14879 VSS.n1467 VSS.n1466 0.00233824
R14880 VSS.n462 VSS.n461 0.00233824
R14881 VSS.n1470 VSS.n1461 0.00233824
R14882 VSS.n1450 VSS.n1447 0.00233824
R14883 VSS.n470 VSS.n455 0.00233824
R14884 VSS.n2004 VSS.n2003 0.00233824
R14885 VSS.n2000 VSS.n1999 0.00233824
R14886 VSS.n1993 VSS.n1992 0.00233824
R14887 VSS.n2128 VSS.n2125 0.00233824
R14888 VSS.n2107 VSS.n2106 0.00233824
R14889 VSS.n2093 VSS.n2092 0.00233824
R14890 VSS.n2134 VSS.n2133 0.00233824
R14891 VSS.n370 VSS.n369 0.00233824
R14892 VSS.n2084 VSS.n375 0.00233824
R14893 VSS.n394 VSS.n393 0.00233824
R14894 VSS.n390 VSS.n389 0.00233824
R14895 VSS.n383 VSS.n382 0.00233824
R14896 VSS.n406 VSS.n405 0.00233824
R14897 VSS.n412 VSS.n411 0.00233824
R14898 VSS.n418 VSS.n417 0.00233824
R14899 VSS.n428 VSS.n426 0.00233824
R14900 VSS.n1944 VSS.n1942 0.00233824
R14901 VSS.n1972 VSS.n1971 0.00233824
R14902 VSS.n1948 VSS.n1937 0.00233824
R14903 VSS.n1959 VSS.n1955 0.00233824
R14904 VSS.n1980 VSS.n1966 0.00233824
R14905 VSS.n2016 VSS.n2015 0.00233824
R14906 VSS.n2022 VSS.n2021 0.00233824
R14907 VSS.n2028 VSS.n2027 0.00233824
R14908 VSS.n1757 VSS.n1756 0.00233824
R14909 VSS.n1753 VSS.n1752 0.00233824
R14910 VSS.n1746 VSS.n1745 0.00233824
R14911 VSS.n1646 VSS.n1644 0.00233824
R14912 VSS.n1667 VSS.n1666 0.00233824
R14913 VSS.n1700 VSS.n1699 0.00233824
R14914 VSS.n1670 VSS.n1661 0.00233824
R14915 VSS.n1684 VSS.n1681 0.00233824
R14916 VSS.n1708 VSS.n1693 0.00233824
R14917 VSS.n1891 VSS.n1890 0.00233824
R14918 VSS.n1887 VSS.n1886 0.00233824
R14919 VSS.n1880 VSS.n1879 0.00233824
R14920 VSS.n1903 VSS.n1902 0.00233824
R14921 VSS.n1867 VSS.n1866 0.00233824
R14922 VSS.n1856 VSS.n1855 0.00233824
R14923 VSS.n1833 VSS.n1831 0.00233824
R14924 VSS.n1817 VSS.n1815 0.00233824
R14925 VSS.n1786 VSS.n1785 0.00233824
R14926 VSS.n1821 VSS.n1810 0.00233824
R14927 VSS.n1804 VSS.n1800 0.00233824
R14928 VSS.n1794 VSS.n1780 0.00233824
R14929 VSS.n1769 VSS.n1768 0.00233824
R14930 VSS.n1733 VSS.n1732 0.00233824
R14931 VSS.n1722 VSS.n1721 0.00233824
R14932 VSS.n358 VSS.n356 0.00233824
R14933 VSS.n2213 VSS.n2212 0.00233824
R14934 VSS.n2173 VSS.n2172 0.00233824
R14935 VSS.n2214 VSS.n2206 0.00233824
R14936 VSS.n2195 VSS.n2192 0.00233824
R14937 VSS.n2181 VSS.n2163 0.00233824
R14938 VSS.n1535 VSS.n1527 0.00233824
R14939 VSS.n1549 VSS.n1546 0.00233824
R14940 VSS.n1574 VSS.n1558 0.00233824
R14941 VSS.n2118 VSS.n368 0.00233824
R14942 VSS.n2115 VSS.n2114 0.00233824
R14943 VSS.n2101 VSS.n2100 0.00233824
R14944 VSS.n1622 VSS.n1621 0.00233824
R14945 VSS.n1605 VSS.n1604 0.00233824
R14946 VSS.n1594 VSS.n1593 0.00233824
R14947 VSS.n1511 VSS.n1509 0.00233824
R14948 VSS.n1532 VSS.n1531 0.00233824
R14949 VSS.n1565 VSS.n1564 0.00233824
R14950 VSS.n548 VSS.n547 0.00233824
R14951 VSS.n544 VSS.n543 0.00233824
R14952 VSS.n537 VSS.n536 0.00233824
R14953 VSS.n1402 VSS.n1401 0.00233824
R14954 VSS.n1396 VSS.n1395 0.00233824
R14955 VSS.n1390 VSS.n1389 0.00233824
R14956 VSS.n641 VSS.n640 0.00233824
R14957 VSS.n637 VSS.n636 0.00233824
R14958 VSS.n620 VSS.n571 0.00233824
R14959 VSS.n566 VSS.n565 0.00233824
R14960 VSS.n560 VSS.n559 0.00233824
R14961 VSS.n651 VSS.n635 0.00233824
R14962 VSS.n661 VSS.n654 0.00233824
R14963 VSS.n665 VSS.n664 0.00233824
R14964 VSS.n475 VSS.n474 0.00233824
R14965 VSS.n481 VSS.n480 0.00233824
R14966 VSS.n487 VSS.n486 0.00233824
R14967 VSS.n2584 VSS.n2583 0.00233824
R14968 VSS.n2594 VSS.n2593 0.00233824
R14969 VSS.n2615 VSS.n2606 0.00233824
R14970 VSS.n292 VSS.n291 0.00221991
R14971 VSS.n15 VSS.n14 0.00221938
R14972 VSS.n1158 VSS.n1157 0.00221938
R14973 VSS.n1353 VSS.n1352 0.00219508
R14974 VSS.n2309 VSS.n2307 0.00218919
R14975 VSS.n707 VSS.n699 0.00218919
R14976 VSS.n714 VSS.n694 0.00218919
R14977 VSS.n2263 VSS.n2250 0.00218919
R14978 VSS.n2297 VSS.n2296 0.00218919
R14979 VSS.n1310 VSS.n1265 0.00218919
R14980 VSS.n2467 VSS.n2466 0.00217458
R14981 VSS.n2466 VSS.n2454 0.00217458
R14982 VSS.n1496 VSS.n1495 0.00217419
R14983 VSS.n778 VSS.n776 0.0021514
R14984 VSS.n523 VSS.n521 0.0021514
R14985 VSS.n347 VSS.n345 0.0021514
R14986 VSS.n2484 VSS.n2482 0.0021514
R14987 VSS.n1778 VSS.n1777 0.00214684
R14988 VSS.n2410 VSS.n2409 0.00211602
R14989 VSS.n2407 VSS.n2406 0.00211602
R14990 VSS.n827 VSS.n826 0.00207191
R14991 VSS.n2867 VSS.n2866 0.00205116
R14992 VSS.n764 VSS.n763 0.00203379
R14993 VSS.n1369 VSS.n1366 0.00201776
R14994 VSS.n1420 VSS.n1419 0.00201154
R14995 VSS.n2620 VSS.n2619 0.00198991
R14996 VSS.n710 VSS.n709 0.00196875
R14997 VSS.n712 VSS.n711 0.00196875
R14998 VSS.n677 VSS.n676 0.00196875
R14999 VSS.n679 VSS.n678 0.00196875
R15000 VSS.n2257 VSS.n2256 0.00196875
R15001 VSS.n2259 VSS.n2258 0.00196875
R15002 VSS.n2261 VSS.n2260 0.00196875
R15003 VSS.n2317 VSS.n2316 0.00196875
R15004 VSS.n2319 VSS.n2318 0.00196875
R15005 VSS.n2322 VSS.n2321 0.00196875
R15006 VSS.n2324 VSS.n2323 0.00196875
R15007 VSS.n1282 VSS.n1281 0.00196875
R15008 VSS.n1293 VSS.n1271 0.00196875
R15009 VSS.n1297 VSS.n1266 0.00196875
R15010 VSS.n1360 VSS.n1359 0.00188889
R15011 VSS.n1157 VSS.n1122 0.00188633
R15012 VSS.n16 VSS.n15 0.00188633
R15013 VSS.n784 VSS.n783 0.00185004
R15014 VSS.n819 VSS.n818 0.00182394
R15015 VSS.n822 VSS.n821 0.00182394
R15016 VSS.n706 VSS.n705 0.00180208
R15017 VSS.n715 VSS.n692 0.00180208
R15018 VSS.n2437 VSS.n2264 0.00180208
R15019 VSS.n2295 VSS.n2294 0.00180208
R15020 VSS.n2355 VSS.n2354 0.00180208
R15021 VSS.n1311 VSS.n1263 0.00180208
R15022 VSS.n2866 VSS 0.00174092
R15023 VSS.n1369 VSS.n1368 0.00166362
R15024 VSS.n2411 VSS.n2407 0.00155801
R15025 VSS.n2411 VSS.n2410 0.00155801
R15026 VSS.n784 VSS.n764 0.00151689
R15027 VSS.n1419 VSS.n1418 0.00150577
R15028 VSS.n1364 VSS.n1363 0.00146875
R15029 VSS.n1363 VSS.n1362 0.00146875
R15030 VSS.n1364 VSS.n1347 0.00143699
R15031 VSS.n1775 VSS 0.0013785
R15032 VSS.n1343 VSS.n675 0.00135454
R15033 VSS.n1418 VSS.n527 0.00130947
R15034 VSS.n290 VSS 0.00123247
R15035 VSS.n2694 VSS.n2693 0.00122817
R15036 VSS.n1499 VSS.n1484 0.00121865
R15037 VSS.n1928 VSS.n1927 0.00121865
R15038 VSS.n527 VSS.n508 0.00120829
R15039 VSS.n1354 VSS.n1353 0.00115602
R15040 VSS.n1652 VSS.n1651 0.00113087
R15041 VSS.n769 VSS.n768 0.0011215
R15042 VSS.n515 VSS.n514 0.0011215
R15043 VSS.n338 VSS.n337 0.0011215
R15044 VSS.n2476 VSS.n2475 0.0011215
R15045 VSS.n1367 VSS 0.0011071
R15046 VSS VSS.n2221 0.00109494
R15047 VSS.n1358 VSS.n1357 0.00104413
R15048 VSS VSS.n797 0.00103208
R15049 VSS.n1357 VSS.n1356 0.00100447
R15050 VSS.n1363 VSS.n1349 0.000885246
R15051 VSS.n1368 VSS.n1367 0.000854144
R15052 VSS.n2406 VSS 0.000834917
R15053 VSS.n2454 VSS.n2453 0.000834917
R15054 VSS.n763 VSS 0.000810231
R15055 VSS.n2863 VSS 0.000810231
R15056 VSS.n2868 VSS.n2867 0.000810231
R15057 VSS.n1366 VSS.n1365 0.000803552
R15058 VSS.n1923 VSS 0.000792835
R15059 VSS.n818 VSS.n817 0.000764789
R15060 VSS.n244 VSS 0.000744156
R15061 VSS.n1494 VSS 0.000735
R15062 VSS.n1361 VSS.n1360 0.000677523
R15063 VSS.n1121 VSS 0.000677358
R15064 VSS.n2409 VSS.n2408 0.000667458
R15065 VSS.n289 VSS.n288 0.000657191
R15066 VSS.n782 VSS.n781 0.000655116
R15067 VSS VSS.n1420 0.000601184
R15068 VSS.n1421 VSS 0.000550592
R15069 VSS.n1356 VSS.n1355 0.000548599
R15070 VSS.n1359 VSS.n1358 0.000518408
R15071 x2.x10.Y.n5 x2.x10.Y.n0 304.151
R15072 x2.x10.Y x2.x10.Y.t3 154.8
R15073 x2.x10.Y x2.x10.Y.t6 154.8
R15074 x2.x10.Y x2.x10.Y.t9 154.8
R15075 x2.x10.Y x2.x10.Y.t4 154.8
R15076 x2.x10.Y x2.x10.Y.t2 154.8
R15077 x2.x10.Y x2.x10.Y.t5 154.8
R15078 x2.x10.Y x2.x10.Y.t8 154.8
R15079 x2.x10.Y x2.x10.Y.t7 154.8
R15080 x2.x10.Y.n2 x2.x10.Y.n0 143.207
R15081 x2.x10.Y x2.x10.Y.n5 134.663
R15082 x2.x10.Y x2.x10.Y.t0 116.097
R15083 x2.x10.Y.n3 x2.x10.Y.t1 25.626
R15084 x2.x10.Y.n1 x2.x10.Y 11.6875
R15085 x2.x10.Y.n4 x2.x10.Y.n3 9.14446
R15086 x2.x10.Y.n2 x2.x10.Y 7.45722
R15087 x2.x10.Y.n4 x2.x10.Y.n2 7.43775
R15088 x2.x10.Y.n1 x2.x10.Y 7.23528
R15089 x2.x10.Y x2.x10.Y.n1 5.04292
R15090 x2.x10.Y.n3 x2.x10.Y.n0 0.969421
R15091 x2.x10.Y.n5 x2.x10.Y.n4 0.652645
R15092 x2.x5[7].floating.n6 x2.x5[7].floating.t2 68.0345
R15093 x2.x5[7].floating.n27 x2.x5[7].floating.t1 68.0345
R15094 x2.x5[7].floating.n45 x2.x5[7].floating.t4 68.0345
R15095 x2.x5[7].floating.n57 x2.x5[7].floating.t7 68.0345
R15096 x2.x5[7].floating.n75 x2.x5[7].floating.t5 68.0345
R15097 x2.x5[7].floating.n87 x2.x5[7].floating.t0 68.0345
R15098 x2.x5[7].floating.n105 x2.x5[7].floating.t3 68.0345
R15099 x2.x5[7].floating.n116 x2.x5[7].floating.t6 68.0345
R15100 x2.x5[7].floating.n135 x2.x5[7].floating.n97 0.660401
R15101 x2.x5[7].floating.n144 x2.x5[7].floating.n82 0.660401
R15102 x2.x5[7].floating.n153 x2.x5[7].floating.n67 0.660401
R15103 x2.x5[7].floating.n162 x2.x5[7].floating.n52 0.660401
R15104 x2.x5[7].floating.n171 x2.x5[7].floating.n37 0.660401
R15105 x2.x5[7].floating.n11 x2.x5[7].floating.n10 0.320345
R15106 x2.x5[7].floating.n122 x2.x5[7].floating.n121 0.308269
R15107 x2.x5[7].floating.n123 x2.x5[7].floating.n122 0.173084
R15108 x2.x5[7].floating.n12 x2.x5[7].floating.n11 0.162103
R15109 x2.x5[7].floating.n122 x2.x5[7].floating 0.100688
R15110 x2.x5[7].floating.n11 x2.x5[7].floating 0.0755007
R15111 x2.x5[7].floating.n97 x2.x5[7].floating.n96 0.0716912
R15112 x2.x5[7].floating.n98 x2.x5[7].floating.n97 0.0716912
R15113 x2.x5[7].floating.n67 x2.x5[7].floating.n66 0.0716912
R15114 x2.x5[7].floating.n68 x2.x5[7].floating.n67 0.0716912
R15115 x2.x5[7].floating.n37 x2.x5[7].floating.n36 0.0716912
R15116 x2.x5[7].floating.n38 x2.x5[7].floating.n37 0.0716912
R15117 x2.x5[7].floating.n171 x2.x5[7].floating.n170 0.0716912
R15118 x2.x5[7].floating.n153 x2.x5[7].floating.n152 0.0716912
R15119 x2.x5[7].floating.n135 x2.x5[7].floating.n134 0.0716912
R15120 x2.x5[7].floating.n93 x2.x5[7].floating.n92 0.0557941
R15121 x2.x5[7].floating.n94 x2.x5[7].floating.n93 0.0557941
R15122 x2.x5[7].floating.n95 x2.x5[7].floating.n94 0.0557941
R15123 x2.x5[7].floating.n96 x2.x5[7].floating.n95 0.0557941
R15124 x2.x5[7].floating.n99 x2.x5[7].floating.n98 0.0557941
R15125 x2.x5[7].floating.n100 x2.x5[7].floating.n99 0.0557941
R15126 x2.x5[7].floating.n101 x2.x5[7].floating.n100 0.0557941
R15127 x2.x5[7].floating.n102 x2.x5[7].floating.n101 0.0557941
R15128 x2.x5[7].floating.n63 x2.x5[7].floating.n62 0.0557941
R15129 x2.x5[7].floating.n64 x2.x5[7].floating.n63 0.0557941
R15130 x2.x5[7].floating.n65 x2.x5[7].floating.n64 0.0557941
R15131 x2.x5[7].floating.n66 x2.x5[7].floating.n65 0.0557941
R15132 x2.x5[7].floating.n69 x2.x5[7].floating.n68 0.0557941
R15133 x2.x5[7].floating.n70 x2.x5[7].floating.n69 0.0557941
R15134 x2.x5[7].floating.n71 x2.x5[7].floating.n70 0.0557941
R15135 x2.x5[7].floating.n72 x2.x5[7].floating.n71 0.0557941
R15136 x2.x5[7].floating.n33 x2.x5[7].floating.n32 0.0557941
R15137 x2.x5[7].floating.n34 x2.x5[7].floating.n33 0.0557941
R15138 x2.x5[7].floating.n35 x2.x5[7].floating.n34 0.0557941
R15139 x2.x5[7].floating.n36 x2.x5[7].floating.n35 0.0557941
R15140 x2.x5[7].floating.n39 x2.x5[7].floating.n38 0.0557941
R15141 x2.x5[7].floating.n40 x2.x5[7].floating.n39 0.0557941
R15142 x2.x5[7].floating.n41 x2.x5[7].floating.n40 0.0557941
R15143 x2.x5[7].floating.n42 x2.x5[7].floating.n41 0.0557941
R15144 x2.x5[7].floating.n20 x2.x5[7].floating.n19 0.0557941
R15145 x2.x5[7].floating.n21 x2.x5[7].floating.n20 0.0557941
R15146 x2.x5[7].floating.n22 x2.x5[7].floating.n21 0.0557941
R15147 x2.x5[7].floating.n23 x2.x5[7].floating.n22 0.0557941
R15148 x2.x5[7].floating.n169 x2.x5[7].floating.n168 0.0557941
R15149 x2.x5[7].floating.n168 x2.x5[7].floating.n167 0.0557941
R15150 x2.x5[7].floating.n167 x2.x5[7].floating.n166 0.0557941
R15151 x2.x5[7].floating.n158 x2.x5[7].floating.n157 0.0557941
R15152 x2.x5[7].floating.n157 x2.x5[7].floating.n156 0.0557941
R15153 x2.x5[7].floating.n156 x2.x5[7].floating.n155 0.0557941
R15154 x2.x5[7].floating.n155 x2.x5[7].floating.n154 0.0557941
R15155 x2.x5[7].floating.n151 x2.x5[7].floating.n150 0.0557941
R15156 x2.x5[7].floating.n150 x2.x5[7].floating.n149 0.0557941
R15157 x2.x5[7].floating.n149 x2.x5[7].floating.n148 0.0557941
R15158 x2.x5[7].floating.n140 x2.x5[7].floating.n139 0.0557941
R15159 x2.x5[7].floating.n139 x2.x5[7].floating.n138 0.0557941
R15160 x2.x5[7].floating.n138 x2.x5[7].floating.n137 0.0557941
R15161 x2.x5[7].floating.n137 x2.x5[7].floating.n136 0.0557941
R15162 x2.x5[7].floating.n133 x2.x5[7].floating.n132 0.0557941
R15163 x2.x5[7].floating.n132 x2.x5[7].floating.n131 0.0557941
R15164 x2.x5[7].floating.n131 x2.x5[7].floating.n130 0.0557941
R15165 x2.x5[7].floating.n16 x2.x5[7].floating.n15 0.0537206
R15166 x2.x5[7].floating.n162 x2.x5[7].floating.n161 0.0537206
R15167 x2.x5[7].floating.n144 x2.x5[7].floating.n143 0.0537206
R15168 x2.x5[7].floating.n126 x2.x5[7].floating.n125 0.0537206
R15169 x2.x5[7].floating.n15 x2.x5[7].floating.n14 0.0530294
R15170 x2.x5[7].floating.n163 x2.x5[7].floating.n162 0.0530294
R15171 x2.x5[7].floating.n145 x2.x5[7].floating.n144 0.0530294
R15172 x2.x5[7].floating.n127 x2.x5[7].floating.n126 0.0530294
R15173 x2.x5[7].floating.n83 x2.x5[7].floating.n82 0.0529559
R15174 x2.x5[7].floating.n53 x2.x5[7].floating.n52 0.0529559
R15175 x2.x5[7].floating.n1 x2.x5[7].floating.n0 0.0529559
R15176 x2.x5[7].floating.n113 x2.x5[7].floating.n112 0.0529559
R15177 x2.x5[7].floating.n112 x2.x5[7].floating.n111 0.0524559
R15178 x2.x5[7].floating.n82 x2.x5[7].floating.n81 0.0524559
R15179 x2.x5[7].floating.n52 x2.x5[7].floating.n51 0.0524559
R15180 x2.x5[7].floating.n2 x2.x5[7].floating.n1 0.0524559
R15181 x2.x5[7].floating.n166 x2.x5[7].floating.n165 0.0523382
R15182 x2.x5[7].floating.n148 x2.x5[7].floating.n147 0.0523382
R15183 x2.x5[7].floating.n130 x2.x5[7].floating.n129 0.0523382
R15184 x2.x5[7].floating.n19 x2.x5[7].floating.n18 0.0516471
R15185 x2.x5[7].floating.n159 x2.x5[7].floating.n158 0.0516471
R15186 x2.x5[7].floating.n141 x2.x5[7].floating.n140 0.0516471
R15187 x2.x5[7].floating x2.x5[7].floating.n171 0.0495735
R15188 x2.x5[7].floating x2.x5[7].floating.n153 0.0495735
R15189 x2.x5[7].floating x2.x5[7].floating.n135 0.0495735
R15190 x2.x5[7].floating.n8 x2.x5[7].floating.n5 0.0408846
R15191 x2.x5[7].floating.n47 x2.x5[7].floating.n44 0.0408846
R15192 x2.x5[7].floating.n77 x2.x5[7].floating.n74 0.0408846
R15193 x2.x5[7].floating.n107 x2.x5[7].floating.n104 0.0408846
R15194 x2.x5[7].floating x2.x5[7].floating.n169 0.0336765
R15195 x2.x5[7].floating x2.x5[7].floating.n151 0.0336765
R15196 x2.x5[7].floating x2.x5[7].floating.n133 0.0336765
R15197 x2.x5[7].floating.n103 x2.x5[7].floating.n102 0.0271618
R15198 x2.x5[7].floating.n73 x2.x5[7].floating.n72 0.0271618
R15199 x2.x5[7].floating.n43 x2.x5[7].floating.n42 0.0271618
R15200 x2.x5[7].floating.n92 x2.x5[7].floating.n91 0.0266618
R15201 x2.x5[7].floating.n62 x2.x5[7].floating.n61 0.0266618
R15202 x2.x5[7].floating.n32 x2.x5[7].floating.n31 0.0266618
R15203 x2.x5[7].floating x2.x5[7].floating.n23 0.0226176
R15204 x2.x5[7].floating.n170 x2.x5[7].floating 0.0226176
R15205 x2.x5[7].floating.n154 x2.x5[7].floating 0.0226176
R15206 x2.x5[7].floating.n152 x2.x5[7].floating 0.0226176
R15207 x2.x5[7].floating.n136 x2.x5[7].floating 0.0226176
R15208 x2.x5[7].floating.n134 x2.x5[7].floating 0.0226176
R15209 x2.x5[7].floating.n119 x2.x5[7].floating.n118 0.021208
R15210 x2.x5[7].floating.n14 x2.x5[7].floating.n13 0.0191618
R15211 x2.x5[7].floating.n164 x2.x5[7].floating.n163 0.0191618
R15212 x2.x5[7].floating.n146 x2.x5[7].floating.n145 0.0191618
R15213 x2.x5[7].floating.n128 x2.x5[7].floating.n127 0.0191618
R15214 x2.x5[7].floating.n17 x2.x5[7].floating.n16 0.0184706
R15215 x2.x5[7].floating.n161 x2.x5[7].floating.n160 0.0184706
R15216 x2.x5[7].floating.n143 x2.x5[7].floating.n142 0.0184706
R15217 x2.x5[7].floating.n125 x2.x5[7].floating.n124 0.0184706
R15218 x2.x5[7].floating.n111 x2.x5[7].floating.n110 0.014
R15219 x2.x5[7].floating.n91 x2.x5[7].floating.n90 0.014
R15220 x2.x5[7].floating.n81 x2.x5[7].floating.n80 0.014
R15221 x2.x5[7].floating.n61 x2.x5[7].floating.n60 0.014
R15222 x2.x5[7].floating.n51 x2.x5[7].floating.n50 0.014
R15223 x2.x5[7].floating.n31 x2.x5[7].floating.n30 0.014
R15224 x2.x5[7].floating.n3 x2.x5[7].floating.n2 0.014
R15225 x2.x5[7].floating.n121 x2.x5[7].floating.n120 0.014
R15226 x2.x5[7].floating.n108 x2.x5[7].floating.n103 0.0135
R15227 x2.x5[7].floating.n84 x2.x5[7].floating.n83 0.0135
R15228 x2.x5[7].floating.n78 x2.x5[7].floating.n73 0.0135
R15229 x2.x5[7].floating.n54 x2.x5[7].floating.n53 0.0135
R15230 x2.x5[7].floating.n48 x2.x5[7].floating.n43 0.0135
R15231 x2.x5[7].floating.n10 x2.x5[7].floating.n9 0.0135
R15232 x2.x5[7].floating.n114 x2.x5[7].floating.n113 0.0135
R15233 x2.x5[7].floating.n29 x2.x5[7].floating.n26 0.0101154
R15234 x2.x5[7].floating.n59 x2.x5[7].floating.n56 0.0101154
R15235 x2.x5[7].floating.n89 x2.x5[7].floating.n86 0.0101154
R15236 x2.x5[7].floating.n18 x2.x5[7].floating.n17 0.00464706
R15237 x2.x5[7].floating.n160 x2.x5[7].floating.n159 0.00464706
R15238 x2.x5[7].floating.n142 x2.x5[7].floating.n141 0.00464706
R15239 x2.x5[7].floating.n124 x2.x5[7].floating.n123 0.00464706
R15240 x2.x5[7].floating.n13 x2.x5[7].floating.n12 0.00395588
R15241 x2.x5[7].floating.n165 x2.x5[7].floating.n164 0.00395588
R15242 x2.x5[7].floating.n147 x2.x5[7].floating.n146 0.00395588
R15243 x2.x5[7].floating.n129 x2.x5[7].floating.n128 0.00395588
R15244 x2.x5[7].floating.n109 x2.x5[7].floating.n108 0.0035
R15245 x2.x5[7].floating.n85 x2.x5[7].floating.n84 0.0035
R15246 x2.x5[7].floating.n79 x2.x5[7].floating.n78 0.0035
R15247 x2.x5[7].floating.n55 x2.x5[7].floating.n54 0.0035
R15248 x2.x5[7].floating.n49 x2.x5[7].floating.n48 0.0035
R15249 x2.x5[7].floating.n25 x2.x5[7].floating.n24 0.0035
R15250 x2.x5[7].floating.n9 x2.x5[7].floating.n4 0.0035
R15251 x2.x5[7].floating.n115 x2.x5[7].floating.n114 0.0035
R15252 x2.x5[7].floating.n110 x2.x5[7].floating.n109 0.003
R15253 x2.x5[7].floating.n90 x2.x5[7].floating.n85 0.003
R15254 x2.x5[7].floating.n80 x2.x5[7].floating.n79 0.003
R15255 x2.x5[7].floating.n60 x2.x5[7].floating.n55 0.003
R15256 x2.x5[7].floating.n50 x2.x5[7].floating.n49 0.003
R15257 x2.x5[7].floating.n30 x2.x5[7].floating.n25 0.003
R15258 x2.x5[7].floating.n4 x2.x5[7].floating.n3 0.003
R15259 x2.x5[7].floating.n120 x2.x5[7].floating.n115 0.003
R15260 x2.x5[7].floating.n28 x2.x5[7].floating.n27 0.00260608
R15261 x2.x5[7].floating.n58 x2.x5[7].floating.n57 0.00260608
R15262 x2.x5[7].floating.n88 x2.x5[7].floating.n87 0.00260608
R15263 x2.x5[7].floating.n117 x2.x5[7].floating.n116 0.00234008
R15264 x2.x5[7].floating.n119 x2.x5[7].floating.n117 0.00200725
R15265 x2.x5[7].floating.n7 x2.x5[7].floating.n6 0.00177054
R15266 x2.x5[7].floating.n46 x2.x5[7].floating.n45 0.00177054
R15267 x2.x5[7].floating.n76 x2.x5[7].floating.n75 0.00177054
R15268 x2.x5[7].floating.n106 x2.x5[7].floating.n105 0.00177054
R15269 x2.x5[7].floating.n8 x2.x5[7].floating.n7 0.00174992
R15270 x2.x5[7].floating.n47 x2.x5[7].floating.n46 0.00174992
R15271 x2.x5[7].floating.n77 x2.x5[7].floating.n76 0.00174992
R15272 x2.x5[7].floating.n107 x2.x5[7].floating.n106 0.00174992
R15273 x2.x5[7].floating.n29 x2.x5[7].floating.n28 0.00101477
R15274 x2.x5[7].floating.n59 x2.x5[7].floating.n58 0.00101477
R15275 x2.x5[7].floating.n89 x2.x5[7].floating.n88 0.00101477
R15276 x2.x5[7].floating.n108 x2.x5[7].floating.n107 0.00053972
R15277 x2.x5[7].floating.n90 x2.x5[7].floating.n89 0.00053972
R15278 x2.x5[7].floating.n78 x2.x5[7].floating.n77 0.00053972
R15279 x2.x5[7].floating.n60 x2.x5[7].floating.n59 0.00053972
R15280 x2.x5[7].floating.n48 x2.x5[7].floating.n47 0.00053972
R15281 x2.x5[7].floating.n30 x2.x5[7].floating.n29 0.00053972
R15282 x2.x5[7].floating.n9 x2.x5[7].floating.n8 0.00053972
R15283 x2.x5[7].floating.n120 x2.x5[7].floating.n119 0.00053972
R15284 in.t9 in.t21 221.72
R15285 in.t14 in.t9 221.72
R15286 in.t2 in.t14 221.72
R15287 in.t12 in.t2 221.72
R15288 in.t16 in.t12 221.72
R15289 in.t17 in.t1 221.72
R15290 in.t6 in.t17 221.72
R15291 in.t18 in.t6 221.72
R15292 in.t13 in.t18 221.72
R15293 in.t3 in.t13 221.72
R15294 in.t20 in.t3 221.72
R15295 in.t10 in.t20 221.72
R15296 in.t4 in.t8 221.72
R15297 in.t15 in.t4 221.72
R15298 in.t5 in.t15 221.72
R15299 in.t0 in.t5 221.72
R15300 in.t11 in.t0 221.72
R15301 in.t7 in.t11 221.72
R15302 in.t19 in.t7 221.72
R15303 in.n5 in.t16 154.8
R15304 in.n0 in 89.9738
R15305 in.n1 in.t10 78.7272
R15306 in.n0 in.t19 74.6592
R15307 in.n2 in 40.1672
R15308 in.n3 in.n1 32.1338
R15309 in in.n1 21.4227
R15310 in.n4 in.n0 21.3547
R15311 in.n4 in.n3 17.8279
R15312 in.n5 in.n4 13.4163
R15313 in.n2 in 11.8854
R15314 in.n3 in.n2 3.96214
R15315 in.n6 in 1.64944
R15316 in.n6 in 0.10169
R15317 in in.n6 0.00215441
R15318 in.n6 in.n5 0.00197059
R15319 sample_code1[1] sample_code1[1].t1 140.387
R15320 sample_code1[1].n0 sample_code1[1].t0 140.34
R15321 sample_code1[1].n0 sample_code1[1] 0.204269
R15322 sample_code1[1] sample_code1[1].n0 0.00197059
R15323 sample_code2[3].n0 sample_code2[3].t0 229.964
R15324 sample_code2[3].n0 sample_code2[3].t1 158.363
R15325 sample_code2[3].n1 sample_code2[3].n0 8.13263
R15326 sample_code2[3].n1 sample_code2[3] 2.67916
R15327 sample_code2[3] sample_code2[3].n2 2.1255
R15328 sample_code2[3] sample_code2[3].n1 1.84241
R15329 sample_code2[3].n2 sample_code2[3] 0.271333
R15330 sample_code2[3].n2 sample_code2[3] 0.0169729
R15331 x4.x10.Y x4.x10.Y.t5 154.847
R15332 x4.x10.Y x4.x10.Y.t8 154.8
R15333 x4.x10.Y x4.x10.Y.t9 154.8
R15334 x4.x10.Y x4.x10.Y.t2 154.8
R15335 x4.x10.Y x4.x10.Y.t3 154.8
R15336 x4.x10.Y x4.x10.Y.t4 154.8
R15337 x4.x10.Y x4.x10.Y.t6 154.8
R15338 x4.x10.Y x4.x10.Y.t7 154.8
R15339 x4.x10.Y.n0 x4.x10.Y 134.239
R15340 x4.x10.Y x4.x10.Y.t0 106.635
R15341 x4.x10.Y.n2 x4.x10.Y.t1 24.6567
R15342 x4.x10.Y.n5 x4.x10.Y.n4 12.4089
R15343 x4.x10.Y.n3 x4.x10.Y.n2 9.12522
R15344 x4.x10.Y.n4 x4.x10.Y.n3 7.34048
R15345 x4.x10.Y.n5 x4.x10.Y 2.22659
R15346 x4.x10.Y.n2 x4.x10.Y.n1 1.93377
R15347 x4.x10.Y x4.x10.Y.n5 1.55202
R15348 x4.x10.Y.n3 x4.x10.Y.n0 0.69928
R15349 x4.x5[7].floating.n95 x4.x5[7].floating.t7 68.0345
R15350 x4.x5[7].floating.n24 x4.x5[7].floating.t0 68.0345
R15351 x4.x5[7].floating.n42 x4.x5[7].floating.t1 68.0345
R15352 x4.x5[7].floating.n54 x4.x5[7].floating.t4 68.0345
R15353 x4.x5[7].floating.n154 x4.x5[7].floating.t2 68.0345
R15354 x4.x5[7].floating.n142 x4.x5[7].floating.t3 68.0345
R15355 x4.x5[7].floating.n12 x4.x5[7].floating.t5 68.0345
R15356 x4.x5[7].floating.n109 x4.x5[7].floating.t6 68.0345
R15357 x4.x5[7].floating.n73 x4.x5[7].floating.n35 0.660401
R15358 x4.x5[7].floating.n91 x4.x5[7].floating.n90 0.660401
R15359 x4.x5[7].floating.n130 x4.x5[7].floating.n20 0.660401
R15360 x4.x5[7].floating.n139 x4.x5[7].floating.n5 0.660401
R15361 x4.x5[7].floating.n121 x4.x5[7].floating.n120 0.660401
R15362 x4.x5[7].floating.n60 x4.x5[7].floating.n59 0.320345
R15363 x4.x5[7].floating.n160 x4.x5[7].floating.n159 0.308269
R15364 x4.x5[7].floating.n161 x4.x5[7].floating.n160 0.173084
R15365 x4.x5[7].floating.n61 x4.x5[7].floating.n60 0.162103
R15366 x4.x5[7].floating.n160 x4.x5[7].floating 0.100688
R15367 x4.x5[7].floating.n60 x4.x5[7].floating 0.0755007
R15368 x4.x5[7].floating.n36 x4.x5[7].floating.n35 0.0716912
R15369 x4.x5[7].floating.n35 x4.x5[7].floating.n34 0.0716912
R15370 x4.x5[7].floating.n6 x4.x5[7].floating.n5 0.0716912
R15371 x4.x5[7].floating.n5 x4.x5[7].floating.n4 0.0716912
R15372 x4.x5[7].floating.n74 x4.x5[7].floating.n73 0.0716912
R15373 x4.x5[7].floating.n122 x4.x5[7].floating.n121 0.0716912
R15374 x4.x5[7].floating.n140 x4.x5[7].floating.n139 0.0716912
R15375 x4.x5[7].floating.n120 x4.x5[7].floating.n105 0.0716912
R15376 x4.x5[7].floating.n120 x4.x5[7].floating.n119 0.0716912
R15377 x4.x5[7].floating.n40 x4.x5[7].floating.n39 0.0557941
R15378 x4.x5[7].floating.n39 x4.x5[7].floating.n38 0.0557941
R15379 x4.x5[7].floating.n38 x4.x5[7].floating.n37 0.0557941
R15380 x4.x5[7].floating.n37 x4.x5[7].floating.n36 0.0557941
R15381 x4.x5[7].floating.n34 x4.x5[7].floating.n33 0.0557941
R15382 x4.x5[7].floating.n33 x4.x5[7].floating.n32 0.0557941
R15383 x4.x5[7].floating.n32 x4.x5[7].floating.n31 0.0557941
R15384 x4.x5[7].floating.n31 x4.x5[7].floating.n30 0.0557941
R15385 x4.x5[7].floating.n10 x4.x5[7].floating.n9 0.0557941
R15386 x4.x5[7].floating.n9 x4.x5[7].floating.n8 0.0557941
R15387 x4.x5[7].floating.n8 x4.x5[7].floating.n7 0.0557941
R15388 x4.x5[7].floating.n7 x4.x5[7].floating.n6 0.0557941
R15389 x4.x5[7].floating.n4 x4.x5[7].floating.n3 0.0557941
R15390 x4.x5[7].floating.n3 x4.x5[7].floating.n2 0.0557941
R15391 x4.x5[7].floating.n2 x4.x5[7].floating.n1 0.0557941
R15392 x4.x5[7].floating.n1 x4.x5[7].floating.n0 0.0557941
R15393 x4.x5[7].floating.n69 x4.x5[7].floating.n68 0.0557941
R15394 x4.x5[7].floating.n70 x4.x5[7].floating.n69 0.0557941
R15395 x4.x5[7].floating.n71 x4.x5[7].floating.n70 0.0557941
R15396 x4.x5[7].floating.n72 x4.x5[7].floating.n71 0.0557941
R15397 x4.x5[7].floating.n76 x4.x5[7].floating.n75 0.0557941
R15398 x4.x5[7].floating.n77 x4.x5[7].floating.n76 0.0557941
R15399 x4.x5[7].floating.n78 x4.x5[7].floating.n77 0.0557941
R15400 x4.x5[7].floating.n86 x4.x5[7].floating.n85 0.0557941
R15401 x4.x5[7].floating.n85 x4.x5[7].floating.n84 0.0557941
R15402 x4.x5[7].floating.n84 x4.x5[7].floating.n83 0.0557941
R15403 x4.x5[7].floating.n83 x4.x5[7].floating.n82 0.0557941
R15404 x4.x5[7].floating.n124 x4.x5[7].floating.n123 0.0557941
R15405 x4.x5[7].floating.n125 x4.x5[7].floating.n124 0.0557941
R15406 x4.x5[7].floating.n126 x4.x5[7].floating.n125 0.0557941
R15407 x4.x5[7].floating.n135 x4.x5[7].floating.n134 0.0557941
R15408 x4.x5[7].floating.n136 x4.x5[7].floating.n135 0.0557941
R15409 x4.x5[7].floating.n137 x4.x5[7].floating.n136 0.0557941
R15410 x4.x5[7].floating.n138 x4.x5[7].floating.n137 0.0557941
R15411 x4.x5[7].floating.n171 x4.x5[7].floating.n170 0.0557941
R15412 x4.x5[7].floating.n170 x4.x5[7].floating.n169 0.0557941
R15413 x4.x5[7].floating.n169 x4.x5[7].floating.n168 0.0557941
R15414 x4.x5[7].floating.n102 x4.x5[7].floating.n101 0.0557941
R15415 x4.x5[7].floating.n103 x4.x5[7].floating.n102 0.0557941
R15416 x4.x5[7].floating.n104 x4.x5[7].floating.n103 0.0557941
R15417 x4.x5[7].floating.n105 x4.x5[7].floating.n104 0.0557941
R15418 x4.x5[7].floating.n119 x4.x5[7].floating.n118 0.0557941
R15419 x4.x5[7].floating.n118 x4.x5[7].floating.n117 0.0557941
R15420 x4.x5[7].floating.n117 x4.x5[7].floating.n116 0.0557941
R15421 x4.x5[7].floating.n116 x4.x5[7].floating.n115 0.0557941
R15422 x4.x5[7].floating.n65 x4.x5[7].floating.n64 0.0537206
R15423 x4.x5[7].floating.n90 x4.x5[7].floating.n89 0.0537206
R15424 x4.x5[7].floating.n131 x4.x5[7].floating.n130 0.0537206
R15425 x4.x5[7].floating.n164 x4.x5[7].floating.n163 0.0537206
R15426 x4.x5[7].floating.n64 x4.x5[7].floating.n63 0.0530294
R15427 x4.x5[7].floating.n90 x4.x5[7].floating.n81 0.0530294
R15428 x4.x5[7].floating.n130 x4.x5[7].floating.n129 0.0530294
R15429 x4.x5[7].floating.n165 x4.x5[7].floating.n164 0.0530294
R15430 x4.x5[7].floating.n92 x4.x5[7].floating.n91 0.0529559
R15431 x4.x5[7].floating.n50 x4.x5[7].floating.n49 0.0529559
R15432 x4.x5[7].floating.n20 x4.x5[7].floating.n19 0.0529559
R15433 x4.x5[7].floating.n151 x4.x5[7].floating.n150 0.0529559
R15434 x4.x5[7].floating.n51 x4.x5[7].floating.n50 0.0524559
R15435 x4.x5[7].floating.n91 x4.x5[7].floating.n21 0.0524559
R15436 x4.x5[7].floating.n106 x4.x5[7].floating.n20 0.0524559
R15437 x4.x5[7].floating.n150 x4.x5[7].floating.n149 0.0524559
R15438 x4.x5[7].floating.n79 x4.x5[7].floating.n78 0.0523382
R15439 x4.x5[7].floating.n127 x4.x5[7].floating.n126 0.0523382
R15440 x4.x5[7].floating.n168 x4.x5[7].floating.n167 0.0523382
R15441 x4.x5[7].floating.n68 x4.x5[7].floating.n67 0.0516471
R15442 x4.x5[7].floating.n87 x4.x5[7].floating.n86 0.0516471
R15443 x4.x5[7].floating.n134 x4.x5[7].floating.n133 0.0516471
R15444 x4.x5[7].floating.n73 x4.x5[7].floating 0.0495735
R15445 x4.x5[7].floating.n121 x4.x5[7].floating 0.0495735
R15446 x4.x5[7].floating.n139 x4.x5[7].floating 0.0495735
R15447 x4.x5[7].floating.n98 x4.x5[7].floating.n97 0.0408846
R15448 x4.x5[7].floating.n45 x4.x5[7].floating.n44 0.0408846
R15449 x4.x5[7].floating.n157 x4.x5[7].floating.n156 0.0408846
R15450 x4.x5[7].floating.n15 x4.x5[7].floating.n14 0.0408846
R15451 x4.x5[7].floating.n75 x4.x5[7].floating 0.0336765
R15452 x4.x5[7].floating.n123 x4.x5[7].floating 0.0336765
R15453 x4.x5[7].floating x4.x5[7].floating.n171 0.0336765
R15454 x4.x5[7].floating.n30 x4.x5[7].floating.n29 0.0271618
R15455 x4.x5[7].floating.n115 x4.x5[7].floating.n114 0.0271618
R15456 x4.x5[7].floating.n101 x4.x5[7].floating.n100 0.0266618
R15457 x4.x5[7].floating.n41 x4.x5[7].floating.n40 0.0266618
R15458 x4.x5[7].floating.n11 x4.x5[7].floating.n10 0.0266618
R15459 x4.x5[7].floating x4.x5[7].floating.n72 0.0226176
R15460 x4.x5[7].floating x4.x5[7].floating.n74 0.0226176
R15461 x4.x5[7].floating.n82 x4.x5[7].floating 0.0226176
R15462 x4.x5[7].floating x4.x5[7].floating.n122 0.0226176
R15463 x4.x5[7].floating x4.x5[7].floating.n138 0.0226176
R15464 x4.x5[7].floating x4.x5[7].floating.n140 0.0226176
R15465 x4.x5[7].floating.n63 x4.x5[7].floating.n62 0.0191618
R15466 x4.x5[7].floating.n81 x4.x5[7].floating.n80 0.0191618
R15467 x4.x5[7].floating.n129 x4.x5[7].floating.n128 0.0191618
R15468 x4.x5[7].floating.n166 x4.x5[7].floating.n165 0.0191618
R15469 x4.x5[7].floating.n66 x4.x5[7].floating.n65 0.0184706
R15470 x4.x5[7].floating.n89 x4.x5[7].floating.n88 0.0184706
R15471 x4.x5[7].floating.n132 x4.x5[7].floating.n131 0.0184706
R15472 x4.x5[7].floating.n163 x4.x5[7].floating.n162 0.0184706
R15473 x4.x5[7].floating.n100 x4.x5[7].floating.n99 0.014
R15474 x4.x5[7].floating.n52 x4.x5[7].floating.n51 0.014
R15475 x4.x5[7].floating.n46 x4.x5[7].floating.n41 0.014
R15476 x4.x5[7].floating.n22 x4.x5[7].floating.n21 0.014
R15477 x4.x5[7].floating.n16 x4.x5[7].floating.n11 0.014
R15478 x4.x5[7].floating.n149 x4.x5[7].floating.n148 0.014
R15479 x4.x5[7].floating.n159 x4.x5[7].floating.n158 0.014
R15480 x4.x5[7].floating.n107 x4.x5[7].floating.n106 0.014
R15481 x4.x5[7].floating.n93 x4.x5[7].floating.n92 0.0135
R15482 x4.x5[7].floating.n59 x4.x5[7].floating.n58 0.0135
R15483 x4.x5[7].floating.n49 x4.x5[7].floating.n48 0.0135
R15484 x4.x5[7].floating.n29 x4.x5[7].floating.n28 0.0135
R15485 x4.x5[7].floating.n19 x4.x5[7].floating.n18 0.0135
R15486 x4.x5[7].floating.n146 x4.x5[7].floating.n141 0.0135
R15487 x4.x5[7].floating.n152 x4.x5[7].floating.n151 0.0135
R15488 x4.x5[7].floating.n114 x4.x5[7].floating.n113 0.0135
R15489 x4.x5[7].floating.n27 x4.x5[7].floating.n26 0.0120385
R15490 x4.x5[7].floating.n57 x4.x5[7].floating.n56 0.0120385
R15491 x4.x5[7].floating.n145 x4.x5[7].floating.n144 0.0120385
R15492 x4.x5[7].floating.n112 x4.x5[7].floating.n111 0.0120385
R15493 x4.x5[7].floating.n67 x4.x5[7].floating.n66 0.00464706
R15494 x4.x5[7].floating.n88 x4.x5[7].floating.n87 0.00464706
R15495 x4.x5[7].floating.n133 x4.x5[7].floating.n132 0.00464706
R15496 x4.x5[7].floating.n162 x4.x5[7].floating.n161 0.00464706
R15497 x4.x5[7].floating.n62 x4.x5[7].floating.n61 0.00395588
R15498 x4.x5[7].floating.n80 x4.x5[7].floating.n79 0.00395588
R15499 x4.x5[7].floating.n128 x4.x5[7].floating.n127 0.00395588
R15500 x4.x5[7].floating.n167 x4.x5[7].floating.n166 0.00395588
R15501 x4.x5[7].floating.n110 x4.x5[7].floating.n109 0.00359614
R15502 x4.x5[7].floating.n25 x4.x5[7].floating.n24 0.00359614
R15503 x4.x5[7].floating.n55 x4.x5[7].floating.n54 0.00359614
R15504 x4.x5[7].floating.n143 x4.x5[7].floating.n142 0.00359614
R15505 x4.x5[7].floating.n94 x4.x5[7].floating.n93 0.0035
R15506 x4.x5[7].floating.n58 x4.x5[7].floating.n53 0.0035
R15507 x4.x5[7].floating.n48 x4.x5[7].floating.n47 0.0035
R15508 x4.x5[7].floating.n28 x4.x5[7].floating.n23 0.0035
R15509 x4.x5[7].floating.n18 x4.x5[7].floating.n17 0.0035
R15510 x4.x5[7].floating.n147 x4.x5[7].floating.n146 0.0035
R15511 x4.x5[7].floating.n153 x4.x5[7].floating.n152 0.0035
R15512 x4.x5[7].floating.n113 x4.x5[7].floating.n108 0.0035
R15513 x4.x5[7].floating.n99 x4.x5[7].floating.n94 0.003
R15514 x4.x5[7].floating.n53 x4.x5[7].floating.n52 0.003
R15515 x4.x5[7].floating.n47 x4.x5[7].floating.n46 0.003
R15516 x4.x5[7].floating.n23 x4.x5[7].floating.n22 0.003
R15517 x4.x5[7].floating.n17 x4.x5[7].floating.n16 0.003
R15518 x4.x5[7].floating.n148 x4.x5[7].floating.n147 0.003
R15519 x4.x5[7].floating.n158 x4.x5[7].floating.n153 0.003
R15520 x4.x5[7].floating.n108 x4.x5[7].floating.n107 0.003
R15521 x4.x5[7].floating.n155 x4.x5[7].floating.n154 0.00277942
R15522 x4.x5[7].floating.n96 x4.x5[7].floating.n95 0.0023396
R15523 x4.x5[7].floating.n43 x4.x5[7].floating.n42 0.0023396
R15524 x4.x5[7].floating.n13 x4.x5[7].floating.n12 0.0023396
R15525 x4.x5[7].floating.n157 x4.x5[7].floating.n155 0.00233747
R15526 x4.x5[7].floating.n98 x4.x5[7].floating.n96 0.00200689
R15527 x4.x5[7].floating.n45 x4.x5[7].floating.n43 0.00200689
R15528 x4.x5[7].floating.n15 x4.x5[7].floating.n13 0.00200689
R15529 x4.x5[7].floating.n27 x4.x5[7].floating.n25 0.0010233
R15530 x4.x5[7].floating.n57 x4.x5[7].floating.n55 0.0010233
R15531 x4.x5[7].floating.n145 x4.x5[7].floating.n143 0.0010233
R15532 x4.x5[7].floating.n112 x4.x5[7].floating.n110 0.0010233
R15533 x4.x5[7].floating.n99 x4.x5[7].floating.n98 0.00053972
R15534 x4.x5[7].floating.n58 x4.x5[7].floating.n57 0.00053972
R15535 x4.x5[7].floating.n46 x4.x5[7].floating.n45 0.00053972
R15536 x4.x5[7].floating.n28 x4.x5[7].floating.n27 0.00053972
R15537 x4.x5[7].floating.n16 x4.x5[7].floating.n15 0.00053972
R15538 x4.x5[7].floating.n146 x4.x5[7].floating.n145 0.00053972
R15539 x4.x5[7].floating.n158 x4.x5[7].floating.n157 0.00053972
R15540 x4.x5[7].floating.n113 x4.x5[7].floating.n112 0.00053972
R15541 sample_code2[1] sample_code2[1].t0 140.343
R15542 sample_code2[1].n0 sample_code2[1].t1 140.34
R15543 sample_code2[1] sample_code2[1].n0 0.247783
R15544 sample_code2[1].n0 sample_code2[1] 0.0466957
R15545 sample_code3[2] sample_code3[2].t0 140.387
R15546 sample_code3[2].n2 sample_code3[2].t2 140.34
R15547 sample_code3[2].n0 sample_code3[2].t3 140.34
R15548 sample_code3[2].n1 sample_code3[2].t1 140.34
R15549 sample_code3[2] sample_code3[2].n1 2.87278
R15550 sample_code3[2] sample_code3[2].n0 0.285826
R15551 sample_code3[2].n2 sample_code3[2] 0.220255
R15552 sample_code3[2].n1 sample_code3[2] 0.0466957
R15553 sample_code3[2].n0 sample_code3[2] 0.0466957
R15554 sample_code3[2] sample_code3[2].n2 0.00210741
R15555 out.n2 out.t5 107.647
R15556 out.n1 out.t4 107.647
R15557 out.n2 out.t3 91.5805
R15558 out.n1 out.t2 91.5805
R15559 out.n0 out.t1 68.3658
R15560 out.n2 out.n1 58.5727
R15561 out.n0 out.t0 41.7552
R15562 out.n3 out.n2 13.4143
R15563 out.n3 out.n0 0.501718
R15564 out out.n3 0.416261
R15565 x1.x10.Y x1.x10.Y.t5 154.847
R15566 x1.x10.Y x1.x10.Y.t6 154.8
R15567 x1.x10.Y x1.x10.Y.t8 154.8
R15568 x1.x10.Y x1.x10.Y.t9 154.8
R15569 x1.x10.Y x1.x10.Y.t4 154.8
R15570 x1.x10.Y x1.x10.Y.t2 154.8
R15571 x1.x10.Y x1.x10.Y.t3 154.8
R15572 x1.x10.Y x1.x10.Y.t7 154.8
R15573 x1.x10.Y.n0 x1.x10.Y 134.239
R15574 x1.x10.Y x1.x10.Y.t0 106.635
R15575 x1.x10.Y.n2 x1.x10.Y.t1 24.6567
R15576 x1.x10.Y.n5 x1.x10.Y.n4 12.4089
R15577 x1.x10.Y.n3 x1.x10.Y.n2 9.12522
R15578 x1.x10.Y.n4 x1.x10.Y.n3 7.34048
R15579 x1.x10.Y.n5 x1.x10.Y 2.22659
R15580 x1.x10.Y.n2 x1.x10.Y.n1 1.93377
R15581 x1.x10.Y x1.x10.Y.n5 1.55202
R15582 x1.x10.Y.n3 x1.x10.Y.n0 0.69928
R15583 x1.x5[7].floating.n122 x1.x5[7].floating.t7 68.0345
R15584 x1.x5[7].floating.n3 x1.x5[7].floating.t5 68.0345
R15585 x1.x5[7].floating.n21 x1.x5[7].floating.t0 68.0345
R15586 x1.x5[7].floating.n33 x1.x5[7].floating.t1 68.0345
R15587 x1.x5[7].floating.n51 x1.x5[7].floating.t3 68.0345
R15588 x1.x5[7].floating.n63 x1.x5[7].floating.t4 68.0345
R15589 x1.x5[7].floating.n154 x1.x5[7].floating.t2 68.0345
R15590 x1.x5[7].floating.n142 x1.x5[7].floating.t6 68.0345
R15591 x1.x5[7].floating.n82 x1.x5[7].floating.n44 0.660401
R15592 x1.x5[7].floating.n91 x1.x5[7].floating.n29 0.660401
R15593 x1.x5[7].floating.n100 x1.x5[7].floating.n14 0.660401
R15594 x1.x5[7].floating.n118 x1.x5[7].floating.n117 0.660401
R15595 x1.x5[7].floating.n139 x1.x5[7].floating.n138 0.660401
R15596 x1.x5[7].floating.n69 x1.x5[7].floating.n68 0.320345
R15597 x1.x5[7].floating.n160 x1.x5[7].floating.n159 0.308269
R15598 x1.x5[7].floating.n161 x1.x5[7].floating.n160 0.173084
R15599 x1.x5[7].floating.n70 x1.x5[7].floating.n69 0.162103
R15600 x1.x5[7].floating.n160 x1.x5[7].floating 0.100688
R15601 x1.x5[7].floating.n69 x1.x5[7].floating 0.0755007
R15602 x1.x5[7].floating.n45 x1.x5[7].floating.n44 0.0716912
R15603 x1.x5[7].floating.n44 x1.x5[7].floating.n43 0.0716912
R15604 x1.x5[7].floating.n15 x1.x5[7].floating.n14 0.0716912
R15605 x1.x5[7].floating.n14 x1.x5[7].floating.n13 0.0716912
R15606 x1.x5[7].floating.n83 x1.x5[7].floating.n82 0.0716912
R15607 x1.x5[7].floating.n101 x1.x5[7].floating.n100 0.0716912
R15608 x1.x5[7].floating.n140 x1.x5[7].floating.n139 0.0716912
R15609 x1.x5[7].floating.n138 x1.x5[7].floating.n132 0.0716912
R15610 x1.x5[7].floating.n138 x1.x5[7].floating.n137 0.0716912
R15611 x1.x5[7].floating.n49 x1.x5[7].floating.n48 0.0557941
R15612 x1.x5[7].floating.n48 x1.x5[7].floating.n47 0.0557941
R15613 x1.x5[7].floating.n47 x1.x5[7].floating.n46 0.0557941
R15614 x1.x5[7].floating.n46 x1.x5[7].floating.n45 0.0557941
R15615 x1.x5[7].floating.n43 x1.x5[7].floating.n42 0.0557941
R15616 x1.x5[7].floating.n42 x1.x5[7].floating.n41 0.0557941
R15617 x1.x5[7].floating.n41 x1.x5[7].floating.n40 0.0557941
R15618 x1.x5[7].floating.n40 x1.x5[7].floating.n39 0.0557941
R15619 x1.x5[7].floating.n19 x1.x5[7].floating.n18 0.0557941
R15620 x1.x5[7].floating.n18 x1.x5[7].floating.n17 0.0557941
R15621 x1.x5[7].floating.n17 x1.x5[7].floating.n16 0.0557941
R15622 x1.x5[7].floating.n16 x1.x5[7].floating.n15 0.0557941
R15623 x1.x5[7].floating.n13 x1.x5[7].floating.n12 0.0557941
R15624 x1.x5[7].floating.n12 x1.x5[7].floating.n11 0.0557941
R15625 x1.x5[7].floating.n11 x1.x5[7].floating.n10 0.0557941
R15626 x1.x5[7].floating.n10 x1.x5[7].floating.n9 0.0557941
R15627 x1.x5[7].floating.n78 x1.x5[7].floating.n77 0.0557941
R15628 x1.x5[7].floating.n79 x1.x5[7].floating.n78 0.0557941
R15629 x1.x5[7].floating.n80 x1.x5[7].floating.n79 0.0557941
R15630 x1.x5[7].floating.n81 x1.x5[7].floating.n80 0.0557941
R15631 x1.x5[7].floating.n85 x1.x5[7].floating.n84 0.0557941
R15632 x1.x5[7].floating.n86 x1.x5[7].floating.n85 0.0557941
R15633 x1.x5[7].floating.n87 x1.x5[7].floating.n86 0.0557941
R15634 x1.x5[7].floating.n96 x1.x5[7].floating.n95 0.0557941
R15635 x1.x5[7].floating.n97 x1.x5[7].floating.n96 0.0557941
R15636 x1.x5[7].floating.n98 x1.x5[7].floating.n97 0.0557941
R15637 x1.x5[7].floating.n99 x1.x5[7].floating.n98 0.0557941
R15638 x1.x5[7].floating.n103 x1.x5[7].floating.n102 0.0557941
R15639 x1.x5[7].floating.n104 x1.x5[7].floating.n103 0.0557941
R15640 x1.x5[7].floating.n105 x1.x5[7].floating.n104 0.0557941
R15641 x1.x5[7].floating.n113 x1.x5[7].floating.n112 0.0557941
R15642 x1.x5[7].floating.n112 x1.x5[7].floating.n111 0.0557941
R15643 x1.x5[7].floating.n111 x1.x5[7].floating.n110 0.0557941
R15644 x1.x5[7].floating.n110 x1.x5[7].floating.n109 0.0557941
R15645 x1.x5[7].floating.n171 x1.x5[7].floating.n170 0.0557941
R15646 x1.x5[7].floating.n170 x1.x5[7].floating.n169 0.0557941
R15647 x1.x5[7].floating.n169 x1.x5[7].floating.n168 0.0557941
R15648 x1.x5[7].floating.n129 x1.x5[7].floating.n128 0.0557941
R15649 x1.x5[7].floating.n130 x1.x5[7].floating.n129 0.0557941
R15650 x1.x5[7].floating.n131 x1.x5[7].floating.n130 0.0557941
R15651 x1.x5[7].floating.n132 x1.x5[7].floating.n131 0.0557941
R15652 x1.x5[7].floating.n137 x1.x5[7].floating.n136 0.0557941
R15653 x1.x5[7].floating.n136 x1.x5[7].floating.n135 0.0557941
R15654 x1.x5[7].floating.n135 x1.x5[7].floating.n134 0.0557941
R15655 x1.x5[7].floating.n134 x1.x5[7].floating.n133 0.0557941
R15656 x1.x5[7].floating.n74 x1.x5[7].floating.n73 0.0537206
R15657 x1.x5[7].floating.n92 x1.x5[7].floating.n91 0.0537206
R15658 x1.x5[7].floating.n117 x1.x5[7].floating.n116 0.0537206
R15659 x1.x5[7].floating.n164 x1.x5[7].floating.n163 0.0537206
R15660 x1.x5[7].floating.n73 x1.x5[7].floating.n72 0.0530294
R15661 x1.x5[7].floating.n91 x1.x5[7].floating.n90 0.0530294
R15662 x1.x5[7].floating.n117 x1.x5[7].floating.n108 0.0530294
R15663 x1.x5[7].floating.n165 x1.x5[7].floating.n164 0.0530294
R15664 x1.x5[7].floating.n119 x1.x5[7].floating.n118 0.0529559
R15665 x1.x5[7].floating.n59 x1.x5[7].floating.n58 0.0529559
R15666 x1.x5[7].floating.n29 x1.x5[7].floating.n28 0.0529559
R15667 x1.x5[7].floating.n151 x1.x5[7].floating.n150 0.0529559
R15668 x1.x5[7].floating.n60 x1.x5[7].floating.n59 0.0524559
R15669 x1.x5[7].floating.n30 x1.x5[7].floating.n29 0.0524559
R15670 x1.x5[7].floating.n118 x1.x5[7].floating.n0 0.0524559
R15671 x1.x5[7].floating.n150 x1.x5[7].floating.n149 0.0524559
R15672 x1.x5[7].floating.n88 x1.x5[7].floating.n87 0.0523382
R15673 x1.x5[7].floating.n106 x1.x5[7].floating.n105 0.0523382
R15674 x1.x5[7].floating.n168 x1.x5[7].floating.n167 0.0523382
R15675 x1.x5[7].floating.n77 x1.x5[7].floating.n76 0.0516471
R15676 x1.x5[7].floating.n95 x1.x5[7].floating.n94 0.0516471
R15677 x1.x5[7].floating.n114 x1.x5[7].floating.n113 0.0516471
R15678 x1.x5[7].floating.n82 x1.x5[7].floating 0.0495735
R15679 x1.x5[7].floating.n100 x1.x5[7].floating 0.0495735
R15680 x1.x5[7].floating.n139 x1.x5[7].floating 0.0495735
R15681 x1.x5[7].floating.n125 x1.x5[7].floating.n124 0.0408846
R15682 x1.x5[7].floating.n24 x1.x5[7].floating.n23 0.0408846
R15683 x1.x5[7].floating.n54 x1.x5[7].floating.n53 0.0408846
R15684 x1.x5[7].floating.n157 x1.x5[7].floating.n156 0.0408846
R15685 x1.x5[7].floating.n84 x1.x5[7].floating 0.0336765
R15686 x1.x5[7].floating.n102 x1.x5[7].floating 0.0336765
R15687 x1.x5[7].floating x1.x5[7].floating.n171 0.0336765
R15688 x1.x5[7].floating.n39 x1.x5[7].floating.n38 0.0271618
R15689 x1.x5[7].floating.n9 x1.x5[7].floating.n8 0.0271618
R15690 x1.x5[7].floating.n128 x1.x5[7].floating.n127 0.0266618
R15691 x1.x5[7].floating.n50 x1.x5[7].floating.n49 0.0266618
R15692 x1.x5[7].floating.n20 x1.x5[7].floating.n19 0.0266618
R15693 x1.x5[7].floating x1.x5[7].floating.n81 0.0226176
R15694 x1.x5[7].floating x1.x5[7].floating.n83 0.0226176
R15695 x1.x5[7].floating x1.x5[7].floating.n99 0.0226176
R15696 x1.x5[7].floating x1.x5[7].floating.n101 0.0226176
R15697 x1.x5[7].floating.n109 x1.x5[7].floating 0.0226176
R15698 x1.x5[7].floating x1.x5[7].floating.n140 0.0226176
R15699 x1.x5[7].floating.n72 x1.x5[7].floating.n71 0.0191618
R15700 x1.x5[7].floating.n90 x1.x5[7].floating.n89 0.0191618
R15701 x1.x5[7].floating.n108 x1.x5[7].floating.n107 0.0191618
R15702 x1.x5[7].floating.n166 x1.x5[7].floating.n165 0.0191618
R15703 x1.x5[7].floating.n75 x1.x5[7].floating.n74 0.0184706
R15704 x1.x5[7].floating.n93 x1.x5[7].floating.n92 0.0184706
R15705 x1.x5[7].floating.n116 x1.x5[7].floating.n115 0.0184706
R15706 x1.x5[7].floating.n163 x1.x5[7].floating.n162 0.0184706
R15707 x1.x5[7].floating.n127 x1.x5[7].floating.n126 0.014
R15708 x1.x5[7].floating.n61 x1.x5[7].floating.n60 0.014
R15709 x1.x5[7].floating.n55 x1.x5[7].floating.n50 0.014
R15710 x1.x5[7].floating.n31 x1.x5[7].floating.n30 0.014
R15711 x1.x5[7].floating.n25 x1.x5[7].floating.n20 0.014
R15712 x1.x5[7].floating.n1 x1.x5[7].floating.n0 0.014
R15713 x1.x5[7].floating.n159 x1.x5[7].floating.n158 0.014
R15714 x1.x5[7].floating.n149 x1.x5[7].floating.n148 0.014
R15715 x1.x5[7].floating.n120 x1.x5[7].floating.n119 0.0135
R15716 x1.x5[7].floating.n68 x1.x5[7].floating.n67 0.0135
R15717 x1.x5[7].floating.n58 x1.x5[7].floating.n57 0.0135
R15718 x1.x5[7].floating.n38 x1.x5[7].floating.n37 0.0135
R15719 x1.x5[7].floating.n28 x1.x5[7].floating.n27 0.0135
R15720 x1.x5[7].floating.n8 x1.x5[7].floating.n7 0.0135
R15721 x1.x5[7].floating.n152 x1.x5[7].floating.n151 0.0135
R15722 x1.x5[7].floating.n146 x1.x5[7].floating.n141 0.0135
R15723 x1.x5[7].floating.n6 x1.x5[7].floating.n5 0.0120385
R15724 x1.x5[7].floating.n36 x1.x5[7].floating.n35 0.0120385
R15725 x1.x5[7].floating.n66 x1.x5[7].floating.n65 0.0120385
R15726 x1.x5[7].floating.n145 x1.x5[7].floating.n144 0.0120385
R15727 x1.x5[7].floating.n76 x1.x5[7].floating.n75 0.00464706
R15728 x1.x5[7].floating.n94 x1.x5[7].floating.n93 0.00464706
R15729 x1.x5[7].floating.n115 x1.x5[7].floating.n114 0.00464706
R15730 x1.x5[7].floating.n162 x1.x5[7].floating.n161 0.00464706
R15731 x1.x5[7].floating.n71 x1.x5[7].floating.n70 0.00395588
R15732 x1.x5[7].floating.n89 x1.x5[7].floating.n88 0.00395588
R15733 x1.x5[7].floating.n107 x1.x5[7].floating.n106 0.00395588
R15734 x1.x5[7].floating.n167 x1.x5[7].floating.n166 0.00395588
R15735 x1.x5[7].floating.n143 x1.x5[7].floating.n142 0.00359614
R15736 x1.x5[7].floating.n4 x1.x5[7].floating.n3 0.00359614
R15737 x1.x5[7].floating.n34 x1.x5[7].floating.n33 0.00359614
R15738 x1.x5[7].floating.n64 x1.x5[7].floating.n63 0.00359614
R15739 x1.x5[7].floating.n121 x1.x5[7].floating.n120 0.0035
R15740 x1.x5[7].floating.n67 x1.x5[7].floating.n62 0.0035
R15741 x1.x5[7].floating.n57 x1.x5[7].floating.n56 0.0035
R15742 x1.x5[7].floating.n37 x1.x5[7].floating.n32 0.0035
R15743 x1.x5[7].floating.n27 x1.x5[7].floating.n26 0.0035
R15744 x1.x5[7].floating.n7 x1.x5[7].floating.n2 0.0035
R15745 x1.x5[7].floating.n153 x1.x5[7].floating.n152 0.0035
R15746 x1.x5[7].floating.n147 x1.x5[7].floating.n146 0.0035
R15747 x1.x5[7].floating.n126 x1.x5[7].floating.n121 0.003
R15748 x1.x5[7].floating.n62 x1.x5[7].floating.n61 0.003
R15749 x1.x5[7].floating.n56 x1.x5[7].floating.n55 0.003
R15750 x1.x5[7].floating.n32 x1.x5[7].floating.n31 0.003
R15751 x1.x5[7].floating.n26 x1.x5[7].floating.n25 0.003
R15752 x1.x5[7].floating.n2 x1.x5[7].floating.n1 0.003
R15753 x1.x5[7].floating.n158 x1.x5[7].floating.n153 0.003
R15754 x1.x5[7].floating.n148 x1.x5[7].floating.n147 0.003
R15755 x1.x5[7].floating.n155 x1.x5[7].floating.n154 0.00277942
R15756 x1.x5[7].floating.n123 x1.x5[7].floating.n122 0.0023396
R15757 x1.x5[7].floating.n22 x1.x5[7].floating.n21 0.0023396
R15758 x1.x5[7].floating.n52 x1.x5[7].floating.n51 0.0023396
R15759 x1.x5[7].floating.n157 x1.x5[7].floating.n155 0.00233747
R15760 x1.x5[7].floating.n125 x1.x5[7].floating.n123 0.00200689
R15761 x1.x5[7].floating.n24 x1.x5[7].floating.n22 0.00200689
R15762 x1.x5[7].floating.n54 x1.x5[7].floating.n52 0.00200689
R15763 x1.x5[7].floating.n6 x1.x5[7].floating.n4 0.0010233
R15764 x1.x5[7].floating.n36 x1.x5[7].floating.n34 0.0010233
R15765 x1.x5[7].floating.n66 x1.x5[7].floating.n64 0.0010233
R15766 x1.x5[7].floating.n145 x1.x5[7].floating.n143 0.0010233
R15767 x1.x5[7].floating.n126 x1.x5[7].floating.n125 0.00053972
R15768 x1.x5[7].floating.n67 x1.x5[7].floating.n66 0.00053972
R15769 x1.x5[7].floating.n55 x1.x5[7].floating.n54 0.00053972
R15770 x1.x5[7].floating.n37 x1.x5[7].floating.n36 0.00053972
R15771 x1.x5[7].floating.n25 x1.x5[7].floating.n24 0.00053972
R15772 x1.x5[7].floating.n7 x1.x5[7].floating.n6 0.00053972
R15773 x1.x5[7].floating.n158 x1.x5[7].floating.n157 0.00053972
R15774 x1.x5[7].floating.n146 x1.x5[7].floating.n145 0.00053972
R15775 sample_code0[1] sample_code0[1].t0 140.387
R15776 sample_code0[1].n0 sample_code0[1].t1 140.34
R15777 sample_code0[1].n0 sample_code0[1] 0.204621
R15778 sample_code0[1] sample_code0[1].n0 0.00216406
R15779 x3.x10.Y.n5 x3.x10.Y.n0 304.151
R15780 x3.x10.Y x3.x10.Y.t2 154.8
R15781 x3.x10.Y x3.x10.Y.t6 154.8
R15782 x3.x10.Y x3.x10.Y.t9 154.8
R15783 x3.x10.Y x3.x10.Y.t5 154.8
R15784 x3.x10.Y x3.x10.Y.t8 154.8
R15785 x3.x10.Y x3.x10.Y.t3 154.8
R15786 x3.x10.Y x3.x10.Y.t7 154.8
R15787 x3.x10.Y x3.x10.Y.t4 154.8
R15788 x3.x10.Y.n2 x3.x10.Y.n0 143.207
R15789 x3.x10.Y x3.x10.Y.n5 134.663
R15790 x3.x10.Y x3.x10.Y.t1 116.097
R15791 x3.x10.Y.n3 x3.x10.Y.t0 25.626
R15792 x3.x10.Y.n1 x3.x10.Y 11.6875
R15793 x3.x10.Y.n4 x3.x10.Y.n3 9.14446
R15794 x3.x10.Y.n2 x3.x10.Y 7.45722
R15795 x3.x10.Y.n4 x3.x10.Y.n2 7.43775
R15796 x3.x10.Y.n1 x3.x10.Y 7.23528
R15797 x3.x10.Y x3.x10.Y.n1 5.04292
R15798 x3.x10.Y.n3 x3.x10.Y.n0 0.969421
R15799 x3.x10.Y.n5 x3.x10.Y.n4 0.652645
R15800 x3.x5[7].floating.n6 x3.x5[7].floating.t5 68.0345
R15801 x3.x5[7].floating.n27 x3.x5[7].floating.t2 68.0345
R15802 x3.x5[7].floating.n57 x3.x5[7].floating.t1 68.0345
R15803 x3.x5[7].floating.n75 x3.x5[7].floating.t4 68.0345
R15804 x3.x5[7].floating.n87 x3.x5[7].floating.t0 68.0345
R15805 x3.x5[7].floating.n105 x3.x5[7].floating.t3 68.0345
R15806 x3.x5[7].floating.n117 x3.x5[7].floating.t7 68.0345
R15807 x3.x5[7].floating.n45 x3.x5[7].floating.t6 68.0345
R15808 x3.x5[7].floating.n135 x3.x5[7].floating.n97 0.660401
R15809 x3.x5[7].floating.n144 x3.x5[7].floating.n82 0.660401
R15810 x3.x5[7].floating.n153 x3.x5[7].floating.n67 0.660401
R15811 x3.x5[7].floating.n162 x3.x5[7].floating.n52 0.660401
R15812 x3.x5[7].floating.n171 x3.x5[7].floating.n37 0.660401
R15813 x3.x5[7].floating.n11 x3.x5[7].floating.n10 0.320345
R15814 x3.x5[7].floating.n122 x3.x5[7].floating.n121 0.308269
R15815 x3.x5[7].floating.n123 x3.x5[7].floating.n122 0.173084
R15816 x3.x5[7].floating.n12 x3.x5[7].floating.n11 0.162103
R15817 x3.x5[7].floating.n122 x3.x5[7].floating 0.100688
R15818 x3.x5[7].floating.n11 x3.x5[7].floating 0.0755007
R15819 x3.x5[7].floating.n97 x3.x5[7].floating.n96 0.0716912
R15820 x3.x5[7].floating.n98 x3.x5[7].floating.n97 0.0716912
R15821 x3.x5[7].floating.n67 x3.x5[7].floating.n66 0.0716912
R15822 x3.x5[7].floating.n68 x3.x5[7].floating.n67 0.0716912
R15823 x3.x5[7].floating.n37 x3.x5[7].floating.n36 0.0716912
R15824 x3.x5[7].floating.n38 x3.x5[7].floating.n37 0.0716912
R15825 x3.x5[7].floating.n171 x3.x5[7].floating.n170 0.0716912
R15826 x3.x5[7].floating.n153 x3.x5[7].floating.n152 0.0716912
R15827 x3.x5[7].floating.n135 x3.x5[7].floating.n134 0.0716912
R15828 x3.x5[7].floating.n93 x3.x5[7].floating.n92 0.0557941
R15829 x3.x5[7].floating.n94 x3.x5[7].floating.n93 0.0557941
R15830 x3.x5[7].floating.n95 x3.x5[7].floating.n94 0.0557941
R15831 x3.x5[7].floating.n96 x3.x5[7].floating.n95 0.0557941
R15832 x3.x5[7].floating.n99 x3.x5[7].floating.n98 0.0557941
R15833 x3.x5[7].floating.n100 x3.x5[7].floating.n99 0.0557941
R15834 x3.x5[7].floating.n101 x3.x5[7].floating.n100 0.0557941
R15835 x3.x5[7].floating.n102 x3.x5[7].floating.n101 0.0557941
R15836 x3.x5[7].floating.n63 x3.x5[7].floating.n62 0.0557941
R15837 x3.x5[7].floating.n64 x3.x5[7].floating.n63 0.0557941
R15838 x3.x5[7].floating.n65 x3.x5[7].floating.n64 0.0557941
R15839 x3.x5[7].floating.n66 x3.x5[7].floating.n65 0.0557941
R15840 x3.x5[7].floating.n69 x3.x5[7].floating.n68 0.0557941
R15841 x3.x5[7].floating.n70 x3.x5[7].floating.n69 0.0557941
R15842 x3.x5[7].floating.n71 x3.x5[7].floating.n70 0.0557941
R15843 x3.x5[7].floating.n72 x3.x5[7].floating.n71 0.0557941
R15844 x3.x5[7].floating.n33 x3.x5[7].floating.n32 0.0557941
R15845 x3.x5[7].floating.n34 x3.x5[7].floating.n33 0.0557941
R15846 x3.x5[7].floating.n35 x3.x5[7].floating.n34 0.0557941
R15847 x3.x5[7].floating.n36 x3.x5[7].floating.n35 0.0557941
R15848 x3.x5[7].floating.n39 x3.x5[7].floating.n38 0.0557941
R15849 x3.x5[7].floating.n40 x3.x5[7].floating.n39 0.0557941
R15850 x3.x5[7].floating.n41 x3.x5[7].floating.n40 0.0557941
R15851 x3.x5[7].floating.n42 x3.x5[7].floating.n41 0.0557941
R15852 x3.x5[7].floating.n20 x3.x5[7].floating.n19 0.0557941
R15853 x3.x5[7].floating.n21 x3.x5[7].floating.n20 0.0557941
R15854 x3.x5[7].floating.n22 x3.x5[7].floating.n21 0.0557941
R15855 x3.x5[7].floating.n23 x3.x5[7].floating.n22 0.0557941
R15856 x3.x5[7].floating.n169 x3.x5[7].floating.n168 0.0557941
R15857 x3.x5[7].floating.n168 x3.x5[7].floating.n167 0.0557941
R15858 x3.x5[7].floating.n167 x3.x5[7].floating.n166 0.0557941
R15859 x3.x5[7].floating.n158 x3.x5[7].floating.n157 0.0557941
R15860 x3.x5[7].floating.n157 x3.x5[7].floating.n156 0.0557941
R15861 x3.x5[7].floating.n156 x3.x5[7].floating.n155 0.0557941
R15862 x3.x5[7].floating.n155 x3.x5[7].floating.n154 0.0557941
R15863 x3.x5[7].floating.n151 x3.x5[7].floating.n150 0.0557941
R15864 x3.x5[7].floating.n150 x3.x5[7].floating.n149 0.0557941
R15865 x3.x5[7].floating.n149 x3.x5[7].floating.n148 0.0557941
R15866 x3.x5[7].floating.n140 x3.x5[7].floating.n139 0.0557941
R15867 x3.x5[7].floating.n139 x3.x5[7].floating.n138 0.0557941
R15868 x3.x5[7].floating.n138 x3.x5[7].floating.n137 0.0557941
R15869 x3.x5[7].floating.n137 x3.x5[7].floating.n136 0.0557941
R15870 x3.x5[7].floating.n133 x3.x5[7].floating.n132 0.0557941
R15871 x3.x5[7].floating.n132 x3.x5[7].floating.n131 0.0557941
R15872 x3.x5[7].floating.n131 x3.x5[7].floating.n130 0.0557941
R15873 x3.x5[7].floating.n16 x3.x5[7].floating.n15 0.0537206
R15874 x3.x5[7].floating.n162 x3.x5[7].floating.n161 0.0537206
R15875 x3.x5[7].floating.n144 x3.x5[7].floating.n143 0.0537206
R15876 x3.x5[7].floating.n126 x3.x5[7].floating.n125 0.0537206
R15877 x3.x5[7].floating.n15 x3.x5[7].floating.n14 0.0530294
R15878 x3.x5[7].floating.n163 x3.x5[7].floating.n162 0.0530294
R15879 x3.x5[7].floating.n145 x3.x5[7].floating.n144 0.0530294
R15880 x3.x5[7].floating.n127 x3.x5[7].floating.n126 0.0530294
R15881 x3.x5[7].floating.n113 x3.x5[7].floating.n112 0.0529559
R15882 x3.x5[7].floating.n83 x3.x5[7].floating.n82 0.0529559
R15883 x3.x5[7].floating.n53 x3.x5[7].floating.n52 0.0529559
R15884 x3.x5[7].floating.n1 x3.x5[7].floating.n0 0.0529559
R15885 x3.x5[7].floating.n112 x3.x5[7].floating.n111 0.0524559
R15886 x3.x5[7].floating.n82 x3.x5[7].floating.n81 0.0524559
R15887 x3.x5[7].floating.n52 x3.x5[7].floating.n51 0.0524559
R15888 x3.x5[7].floating.n2 x3.x5[7].floating.n1 0.0524559
R15889 x3.x5[7].floating.n166 x3.x5[7].floating.n165 0.0523382
R15890 x3.x5[7].floating.n148 x3.x5[7].floating.n147 0.0523382
R15891 x3.x5[7].floating.n130 x3.x5[7].floating.n129 0.0523382
R15892 x3.x5[7].floating.n19 x3.x5[7].floating.n18 0.0516471
R15893 x3.x5[7].floating.n159 x3.x5[7].floating.n158 0.0516471
R15894 x3.x5[7].floating.n141 x3.x5[7].floating.n140 0.0516471
R15895 x3.x5[7].floating x3.x5[7].floating.n171 0.0495735
R15896 x3.x5[7].floating x3.x5[7].floating.n153 0.0495735
R15897 x3.x5[7].floating x3.x5[7].floating.n135 0.0495735
R15898 x3.x5[7].floating.n8 x3.x5[7].floating.n5 0.0408846
R15899 x3.x5[7].floating.n77 x3.x5[7].floating.n74 0.0408846
R15900 x3.x5[7].floating.n107 x3.x5[7].floating.n104 0.0408846
R15901 x3.x5[7].floating.n47 x3.x5[7].floating.n44 0.0408846
R15902 x3.x5[7].floating x3.x5[7].floating.n169 0.0336765
R15903 x3.x5[7].floating x3.x5[7].floating.n151 0.0336765
R15904 x3.x5[7].floating x3.x5[7].floating.n133 0.0336765
R15905 x3.x5[7].floating.n103 x3.x5[7].floating.n102 0.0271618
R15906 x3.x5[7].floating.n73 x3.x5[7].floating.n72 0.0271618
R15907 x3.x5[7].floating.n43 x3.x5[7].floating.n42 0.0271618
R15908 x3.x5[7].floating.n92 x3.x5[7].floating.n91 0.0266618
R15909 x3.x5[7].floating.n62 x3.x5[7].floating.n61 0.0266618
R15910 x3.x5[7].floating.n32 x3.x5[7].floating.n31 0.0266618
R15911 x3.x5[7].floating x3.x5[7].floating.n23 0.0226176
R15912 x3.x5[7].floating.n170 x3.x5[7].floating 0.0226176
R15913 x3.x5[7].floating.n154 x3.x5[7].floating 0.0226176
R15914 x3.x5[7].floating.n152 x3.x5[7].floating 0.0226176
R15915 x3.x5[7].floating.n136 x3.x5[7].floating 0.0226176
R15916 x3.x5[7].floating.n134 x3.x5[7].floating 0.0226176
R15917 x3.x5[7].floating.n14 x3.x5[7].floating.n13 0.0191618
R15918 x3.x5[7].floating.n164 x3.x5[7].floating.n163 0.0191618
R15919 x3.x5[7].floating.n146 x3.x5[7].floating.n145 0.0191618
R15920 x3.x5[7].floating.n128 x3.x5[7].floating.n127 0.0191618
R15921 x3.x5[7].floating.n17 x3.x5[7].floating.n16 0.0184706
R15922 x3.x5[7].floating.n161 x3.x5[7].floating.n160 0.0184706
R15923 x3.x5[7].floating.n143 x3.x5[7].floating.n142 0.0184706
R15924 x3.x5[7].floating.n125 x3.x5[7].floating.n124 0.0184706
R15925 x3.x5[7].floating.n121 x3.x5[7].floating.n120 0.014
R15926 x3.x5[7].floating.n111 x3.x5[7].floating.n110 0.014
R15927 x3.x5[7].floating.n91 x3.x5[7].floating.n90 0.014
R15928 x3.x5[7].floating.n81 x3.x5[7].floating.n80 0.014
R15929 x3.x5[7].floating.n61 x3.x5[7].floating.n60 0.014
R15930 x3.x5[7].floating.n51 x3.x5[7].floating.n50 0.014
R15931 x3.x5[7].floating.n31 x3.x5[7].floating.n30 0.014
R15932 x3.x5[7].floating.n3 x3.x5[7].floating.n2 0.014
R15933 x3.x5[7].floating.n114 x3.x5[7].floating.n113 0.0135
R15934 x3.x5[7].floating.n108 x3.x5[7].floating.n103 0.0135
R15935 x3.x5[7].floating.n84 x3.x5[7].floating.n83 0.0135
R15936 x3.x5[7].floating.n78 x3.x5[7].floating.n73 0.0135
R15937 x3.x5[7].floating.n54 x3.x5[7].floating.n53 0.0135
R15938 x3.x5[7].floating.n48 x3.x5[7].floating.n43 0.0135
R15939 x3.x5[7].floating.n10 x3.x5[7].floating.n9 0.0135
R15940 x3.x5[7].floating.n29 x3.x5[7].floating.n26 0.0101154
R15941 x3.x5[7].floating.n59 x3.x5[7].floating.n56 0.0101154
R15942 x3.x5[7].floating.n89 x3.x5[7].floating.n86 0.0101154
R15943 x3.x5[7].floating.n119 x3.x5[7].floating.n116 0.0101154
R15944 x3.x5[7].floating.n18 x3.x5[7].floating.n17 0.00464706
R15945 x3.x5[7].floating.n160 x3.x5[7].floating.n159 0.00464706
R15946 x3.x5[7].floating.n142 x3.x5[7].floating.n141 0.00464706
R15947 x3.x5[7].floating.n124 x3.x5[7].floating.n123 0.00464706
R15948 x3.x5[7].floating.n13 x3.x5[7].floating.n12 0.00395588
R15949 x3.x5[7].floating.n165 x3.x5[7].floating.n164 0.00395588
R15950 x3.x5[7].floating.n147 x3.x5[7].floating.n146 0.00395588
R15951 x3.x5[7].floating.n129 x3.x5[7].floating.n128 0.00395588
R15952 x3.x5[7].floating.n115 x3.x5[7].floating.n114 0.0035
R15953 x3.x5[7].floating.n109 x3.x5[7].floating.n108 0.0035
R15954 x3.x5[7].floating.n85 x3.x5[7].floating.n84 0.0035
R15955 x3.x5[7].floating.n79 x3.x5[7].floating.n78 0.0035
R15956 x3.x5[7].floating.n55 x3.x5[7].floating.n54 0.0035
R15957 x3.x5[7].floating.n49 x3.x5[7].floating.n48 0.0035
R15958 x3.x5[7].floating.n25 x3.x5[7].floating.n24 0.0035
R15959 x3.x5[7].floating.n9 x3.x5[7].floating.n4 0.0035
R15960 x3.x5[7].floating.n120 x3.x5[7].floating.n115 0.003
R15961 x3.x5[7].floating.n110 x3.x5[7].floating.n109 0.003
R15962 x3.x5[7].floating.n90 x3.x5[7].floating.n85 0.003
R15963 x3.x5[7].floating.n80 x3.x5[7].floating.n79 0.003
R15964 x3.x5[7].floating.n60 x3.x5[7].floating.n55 0.003
R15965 x3.x5[7].floating.n50 x3.x5[7].floating.n49 0.003
R15966 x3.x5[7].floating.n30 x3.x5[7].floating.n25 0.003
R15967 x3.x5[7].floating.n4 x3.x5[7].floating.n3 0.003
R15968 x3.x5[7].floating.n28 x3.x5[7].floating.n27 0.00260608
R15969 x3.x5[7].floating.n58 x3.x5[7].floating.n57 0.00260608
R15970 x3.x5[7].floating.n88 x3.x5[7].floating.n87 0.00260608
R15971 x3.x5[7].floating.n118 x3.x5[7].floating.n117 0.00260608
R15972 x3.x5[7].floating.n46 x3.x5[7].floating.n45 0.00177054
R15973 x3.x5[7].floating.n7 x3.x5[7].floating.n6 0.00177054
R15974 x3.x5[7].floating.n76 x3.x5[7].floating.n75 0.00177054
R15975 x3.x5[7].floating.n106 x3.x5[7].floating.n105 0.00177054
R15976 x3.x5[7].floating.n47 x3.x5[7].floating.n46 0.00174992
R15977 x3.x5[7].floating.n8 x3.x5[7].floating.n7 0.00174992
R15978 x3.x5[7].floating.n77 x3.x5[7].floating.n76 0.00174992
R15979 x3.x5[7].floating.n107 x3.x5[7].floating.n106 0.00174992
R15980 x3.x5[7].floating.n29 x3.x5[7].floating.n28 0.00101477
R15981 x3.x5[7].floating.n59 x3.x5[7].floating.n58 0.00101477
R15982 x3.x5[7].floating.n89 x3.x5[7].floating.n88 0.00101477
R15983 x3.x5[7].floating.n119 x3.x5[7].floating.n118 0.00101477
R15984 x3.x5[7].floating.n120 x3.x5[7].floating.n119 0.00053972
R15985 x3.x5[7].floating.n108 x3.x5[7].floating.n107 0.00053972
R15986 x3.x5[7].floating.n90 x3.x5[7].floating.n89 0.00053972
R15987 x3.x5[7].floating.n78 x3.x5[7].floating.n77 0.00053972
R15988 x3.x5[7].floating.n60 x3.x5[7].floating.n59 0.00053972
R15989 x3.x5[7].floating.n30 x3.x5[7].floating.n29 0.00053972
R15990 x3.x5[7].floating.n9 x3.x5[7].floating.n8 0.00053972
R15991 x3.x5[7].floating.n48 x3.x5[7].floating.n47 0.00053972
R15992 sample_code0[3].n0 sample_code0[3].t1 229.971
R15993 sample_code0[3].n0 sample_code0[3].t0 158.35
R15994 sample_code0[3].n1 sample_code0[3].n0 8.50845
R15995 sample_code0[3].n1 sample_code0[3] 3.95275
R15996 sample_code0[3].n2 sample_code0[3].n1 1.73287
R15997 sample_code0[3].n3 sample_code0[3] 0.474765
R15998 sample_code0[3] sample_code0[3].n3 0.366977
R15999 sample_code0[3].n2 sample_code0[3] 0.339042
R16000 sample_code0[3].n3 sample_code0[3].n2 0.00334091
R16001 sample_code1[3].n0 sample_code1[3].t0 229.971
R16002 sample_code1[3].n0 sample_code1[3].t1 158.35
R16003 sample_code1[3].n1 sample_code1[3].n0 8.50845
R16004 sample_code1[3].n1 sample_code1[3] 3.95275
R16005 sample_code1[3].n2 sample_code1[3].n1 1.73287
R16006 sample_code1[3].n3 sample_code1[3] 0.474765
R16007 sample_code1[3] sample_code1[3].n3 0.366977
R16008 sample_code1[3].n2 sample_code1[3] 0.339042
R16009 sample_code1[3].n3 sample_code1[3].n2 0.00334091
R16010 sample_code0[2] sample_code0[2].t1 140.387
R16011 sample_code0[2].n2 sample_code0[2].t3 140.34
R16012 sample_code0[2].n1 sample_code0[2].t2 140.34
R16013 sample_code0[2].n0 sample_code0[2].t0 140.34
R16014 sample_code0[2].n2 sample_code0[2] 2.82997
R16015 sample_code0[2].n1 sample_code0[2] 0.285826
R16016 sample_code0[2] sample_code0[2].n0 0.264087
R16017 sample_code0[2] sample_code0[2].n1 0.0466957
R16018 sample_code0[2].n0 sample_code0[2] 0.0466957
R16019 sample_code0[2] sample_code0[2].n2 0.00224038
R16020 sample_code3[3].n0 sample_code3[3].t1 229.964
R16021 sample_code3[3].n0 sample_code3[3].t0 158.363
R16022 sample_code3[3].n1 sample_code3[3].n0 8.13263
R16023 sample_code3[3].n1 sample_code3[3] 2.67916
R16024 sample_code3[3] sample_code3[3].n2 2.1255
R16025 sample_code3[3] sample_code3[3].n1 1.84241
R16026 sample_code3[3].n2 sample_code3[3] 0.271333
R16027 sample_code3[3].n2 sample_code3[3] 0.0169729
R16028 sample_code1[2] sample_code1[2].t1 140.387
R16029 sample_code1[2].n2 sample_code1[2].t2 140.34
R16030 sample_code1[2].n1 sample_code1[2].t3 140.34
R16031 sample_code1[2].n0 sample_code1[2].t0 140.34
R16032 sample_code1[2].n2 sample_code1[2] 2.82956
R16033 sample_code1[2].n1 sample_code1[2] 0.285826
R16034 sample_code1[2] sample_code1[2].n0 0.264087
R16035 sample_code1[2] sample_code1[2].n1 0.0466957
R16036 sample_code1[2].n0 sample_code1[2] 0.0466957
R16037 sample_code1[2] sample_code1[2].n2 0.00202988
R16038 sample_code2[2] sample_code2[2].t1 140.387
R16039 sample_code2[2].n2 sample_code2[2].t3 140.34
R16040 sample_code2[2].n0 sample_code2[2].t2 140.34
R16041 sample_code2[2].n1 sample_code2[2].t0 140.34
R16042 sample_code2[2] sample_code2[2].n1 2.87278
R16043 sample_code2[2] sample_code2[2].n0 0.285826
R16044 sample_code2[2].n2 sample_code2[2] 0.219989
R16045 sample_code2[2].n1 sample_code2[2] 0.0466957
R16046 sample_code2[2].n0 sample_code2[2] 0.0466957
R16047 sample_code2[2] sample_code2[2].n2 0.00192617
R16048 sample_code3[0].n0 sample_code3[0].t0 140.34
R16049 sample_code3[0] sample_code3[0].n0 2.45601
R16050 sample_code3[0].n0 sample_code3[0] 0.0365169
R16051 sample_code3[1] sample_code3[1].t0 140.343
R16052 sample_code3[1].n0 sample_code3[1].t1 140.34
R16053 sample_code3[1] sample_code3[1].n0 0.247783
R16054 sample_code3[1].n0 sample_code3[1] 0.0466957
R16055 sample_code2[0].n0 sample_code2[0].t0 140.34
R16056 sample_code2[0].n1 sample_code2[0] 32.8219
R16057 sample_code2[0] sample_code2[0].n1 4.5955
R16058 sample_code2[0].n1 sample_code2[0].n0 2.46566
R16059 sample_code2[0].n0 sample_code2[0] 0.0365169
R16060 sample_code1[0] sample_code1[0].t0 140.376
R16061 sample_code1[0].n0 sample_code1[0] 54.4514
R16062 sample_code1[0] sample_code1[0].n0 4.7207
R16063 sample_code1[0].n0 sample_code1[0] 0.0117229
R16064 sample_code0[0] sample_code0[0].t0 140.376
R16065 sample_code0[0].n0 sample_code0[0] 24.5005
R16066 sample_code0[0] sample_code0[0].n0 4.42631
R16067 sample_code0[0].n0 sample_code0[0] 0.0238871
C0 a_7276_1674# a_7364_1812# 0.00227f
C1 sample_delay_offset sample_code3[2] 0.00886f
C2 sample_code1[2] a_7364_1398# 3.33e-19
C3 x1.x10.Y a_6465_2476# 6.93e-19
C4 x1.IN a_7276_1122# 0.0127f
C5 x4.x2.floating sample_code1[1] 1.73e-20
C6 VDD a_7364_2088# 1.29e-19
C7 sample_code1[1] x2.x9.output_stack 2.48e-21
C8 sample_code0[1] a_6465_2135# 3.4e-20
C9 a_6130_n299# x2.x2.floating 0.00177f
C10 sample_delay_offset x2.x6.SW 0.19f
C11 a_7276_1398# a_7364_1536# 0.00227f
C12 sample_code0[2] sample_code0[1] 1.3f
C13 a_6130_n299# sample_code2[0] 0.00672f
C14 a_680_3339# x4.x10.Y 1.49e-19
C15 VDD x2.IN 0.707f
C16 sample_code1[1] x3.IN 5.1e-20
C17 sample_code0[2] a_567_1950# 7.47e-20
C18 a_592_3477# x4.x6.floating 0.00578f
C19 x2.IN a_12767_n851# 0.00196f
C20 x1.x5[7].floating sample_code1[0] 0.00119f
C21 x4.x5[7].floating x4.x7.floating 0.182f
C22 x1.IN a_7364_2088# 0.00196f
C23 x2.x5[7].floating a_12726_n2240# 0.00154f
C24 x4.x7.floating a_727_1812# 0.00959f
C25 a_12767_n299# x2.x7.floating 8.52e-19
C26 a_12679_n161# x2.x4[3].floating 7.47e-19
C27 x4.x9.output_stack x1.x10.Y 1.93e-19
C28 a_7276_1122# a_7364_1260# 0.00227f
C29 a_6058_n161# x3.x7.floating 8.52e-19
C30 x4.x9.output_stack a_7276_1950# 5.22e-20
C31 a_592_3477# x4.x6.SW 5.11e-20
C32 VDD a_6465_2476# 0.212f
C33 x3.x4[3].floating sample_code2[1] 7.03e-20
C34 a_727_1812# a_655_1812# 0.00227f
C35 x2.x9.output_stack x2.x7.floating 0.185f
C36 x2.IN x2.x10.Y 0.0967f
C37 a_7389_3063# x1.x5[7].floating 0.00169f
C38 sample_code0[2] a_567_1398# 2.81e-19
C39 sample_delay_offset a_6130_n299# 0.00294f
C40 sample_delay_offset x1.x10.Y 0.0402f
C41 a_7301_3201# x1.x10.Y 2.35e-19
C42 a_12679_n713# a_12839_n851# 0.0388f
C43 a_6058_n713# a_6130_n851# 0.00227f
C44 VDD a_6130_n851# 0.00115f
C45 x1.IN a_7364_1536# 3.4e-19
C46 a_6105_n2102# a_6017_n2240# 0.0704f
C47 sample_delay_offset a_7276_1950# 0.0189f
C48 a_12726_n1964# a_12726_n2240# 0.0316f
C49 x4.x7.floating a_727_1260# 0.00925f
C50 VDD x2.x2.floating 0.0334f
C51 VDD sample_code2[0] 0.00338f
C52 a_6058_n713# x2.x2.floating 1.6e-19
C53 a_6058_n713# sample_code2[0] 1.03e-19
C54 x1.IN a_6465_2476# 0.15f
C55 a_727_1536# a_655_1536# 0.00227f
C56 a_12839_n23# x2.x7.floating 0.00218f
C57 sample_delay_offset a_7276_1398# 0.00299f
C58 sample_code2[2] x2.x3[1].floating 0.00624f
C59 a_6130_n299# a_5970_n437# 0.0388f
C60 x1.IN sample_code2[0] 4.21e-20
C61 VDD x4.x9.output_stack 0.594f
C62 a_12767_n161# a_12839_n299# 0.00227f
C63 a_6130_n23# a_6130_n299# 0.0316f
C64 a_5970_n161# x3.x6.SW 7.9e-20
C65 x2.x2.floating x2.x10.Y 0.00202f
C66 a_727_1260# a_655_1260# 0.00227f
C67 a_12679_n161# x2.x9.output_stack 8.05e-20
C68 sample_code2[0] x2.x10.Y 0.0124f
C69 a_12839_n851# x2.x6.SW 0.00179f
C70 x2.IN a_12839_n299# 0.0299f
C71 VDD sample_delay_offset 0.914f
C72 sample_delay_offset a_6058_n713# 0.00154f
C73 VDD a_7301_3201# 0.0923f
C74 x4.x7.floating sample_code1[0] 1.61e-20
C75 x3.x10.Y x2.x5[7].floating 0.00422f
C76 VDD a_40_n1036# 0.235f
C77 sample_code0[0] x4.x4[3].floating 8.34e-20
C78 x1.x9.output_stack x1.x4[3].floating 0.636f
C79 x1.IN x4.x9.output_stack 0.127f
C80 sample_delay_offset a_12767_n851# 0.00167f
C81 x3.x7.floating sample_code2[2] 1.63e-20
C82 a_592_3201# a_680_3063# 0.0704f
C83 sample_code3[2] sample_code2[1] 6.4e-20
C84 sample_code3[1] sample_code2[2] 2.96e-20
C85 x3.IN a_6105_n2378# 0.00832f
C86 x4.x4[3].floating a_727_1536# 8.29e-19
C87 x3.x7.floating x3.x6.floating 0.202f
C88 sample_code1[2] a_567_1122# 1.29e-19
C89 x1.IN sample_delay_offset 0.258f
C90 a_40_n1036# a_40_n1239# 0.0121f
C91 x1.IN a_7301_3201# 0.00866f
C92 a_12839_n23# a_12679_n161# 0.0388f
C93 x3.x6.floating a_6105_n1826# 0.00996f
C94 x1.x6.floating a_7436_1812# 0.00278f
C95 sample_delay_offset x2.x10.Y 0.0403f
C96 sample_delay_offset a_7364_1812# 0.00138f
C97 a_13174_2476# x2.IN 0.145f
C98 a_12679_n437# a_12679_n713# 0.0316f
C99 x2.IN x2.x6.floating 0.0299f
C100 x2.x6.SW a_12814_n1826# 0.00707f
C101 sample_code1[1] a_13174_2135# 3.4e-20
C102 sample_code1[2] sample_code1[1] 5.08f
C103 x3.x5[7].floating x3.x6.floating 1.18f
C104 x4.x10.Y x1.x6.SW 1.5e-20
C105 x2.IN a_12767_n713# 0.0013f
C106 x3.IN a_6058_n575# 7.93e-19
C107 x1.x6.floating a_7436_1260# 0.00109f
C108 sample_delay_offset a_7364_1260# 9.69e-19
C109 a_592_3477# x4.x10.Y 1.02e-19
C110 x2.x5[7].floating a_12814_n2378# 2.14e-19
C111 x4.x10.Y x4.x4[3].floating 0.00668f
C112 VDD x4.x6.floating 5.72f
C113 a_12679_n437# x2.x6.SW 1.28e-19
C114 a_592_3201# x4.x5[7].floating 2.76e-19
C115 sample_delay_offset a_12839_n299# 0.00298f
C116 VDD a_12839_n851# 0.00163f
C117 x1.x5[7].floating sample_code1[2] 0.0056f
C118 a_12814_n2102# a_12726_n2240# 0.0704f
C119 sample_delay_offset a_655_1950# 0.00155f
C120 a_6105_n2102# a_6105_n2378# 0.0316f
C121 VDD x4.x6.SW 0.423f
C122 VDD a_6749_n1036# 0.235f
C123 a_12839_n851# a_12767_n851# 0.00227f
C124 sample_code0[2] a_655_2088# 1.06e-19
C125 x2.x2.floating x2.x3[1].floating 1.17f
C126 x1.x10.Y x1.x3[1].floating 0.00302f
C127 sample_code2[0] x2.x3[1].floating 0.0326f
C128 x3.x9.output_stack sample_code2[2] 2.46e-20
C129 sample_code0[0] a_7276_1950# 0.00181f
C130 x1.x9.output_stack a_7364_2088# 0.00227f
C131 sample_delay_offset a_655_1398# 0.00103f
C132 x1.x9.output_stack x2.IN 0.127f
C133 sample_code3[0] sample_code2[2] 1.48e-20
C134 a_12839_n851# x2.x10.Y 1.69e-19
C135 x3.x9.output_stack x3.x6.floating 0.229f
C136 VDD sample_code2[1] 0.0183f
C137 sample_code0[2] a_655_1536# 3.62e-19
C138 a_6130_n851# x3.x7.floating 0.00409f
C139 sample_delay_offset x2.x6.floating 0.0706f
C140 VDD a_12814_n1826# 0.104f
C141 x3.x7.floating x2.x2.floating 0.0475f
C142 sample_code2[0] x3.x7.floating 0.0075f
C143 sample_code0[0] a_7276_1398# 0.00654f
C144 sample_code3[1] sample_code2[0] 3.47e-20
C145 sample_code1[0] x1.x4[3].floating 6.66e-20
C146 sample_delay_offset a_12767_n713# 0.00155f
C147 x3.x6.floating a_6749_n1239# 0.0013f
C148 x3.IN a_6058_n161# 2.42e-19
C149 sample_code2[2] x2.x4[3].floating 0.53f
C150 sample_delay_offset x2.x3[1].floating 7.23e-20
C151 sample_code1[1] a_567_1122# 8.94e-20
C152 x1.IN sample_code2[1] 4.93e-20
C153 x1.x9.output_stack a_6465_2476# 1.18e-20
C154 x2.x6.SW x2.x5[7].floating 0.00138f
C155 VDD x1.x3[1].floating 0.0301f
C156 VDD sample_code0[0] 0.00321f
C157 sample_code2[1] x2.x10.Y 6.64e-19
C158 sample_code2[0] x3.x5[7].floating 1.4e-20
C159 x2.x10.Y a_12814_n1826# 0.039f
C160 x3.x6.floating a_6017_n1964# 0.0194f
C161 a_6465_2135# x1.x7.floating 7.29e-19
C162 x4.x7.floating sample_code1[2] 1.87e-20
C163 x4.x10.Y x1.x10.Y 1.79e-20
C164 a_5970_n161# x3.x4[3].floating 7.47e-19
C165 sample_code0[2] x4.x4[3].floating 0.532f
C166 a_680_3063# x4.x9.output_stack 0.032f
C167 sample_delay_offset x3.x7.floating 0.261f
C168 a_6130_n575# a_6058_n575# 0.00227f
C169 sample_delay_offset sample_code3[1] 4.51e-19
C170 x1.IN sample_code0[0] 8.71e-19
C171 a_6058_n299# x2.x2.floating 2.21e-19
C172 a_40_n1036# sample_code3[1] 3.4e-20
C173 sample_delay_offset a_6105_n1826# 0.00273f
C174 a_6058_n299# sample_code2[0] 2.39e-19
C175 a_7301_3477# x1.x5[7].floating 2.14e-19
C176 VDD a_6058_n851# 1.29e-19
C177 a_680_3063# sample_delay_offset 3.64e-19
C178 x4.x9.output_stack x4.x3[1].floating 0.341f
C179 x1.x7.floating a_7364_1674# 8.52e-19
C180 x4.x9.output_stack x1.x9.output_stack 2.93e-20
C181 sample_delay_offset x3.x5[7].floating 0.00308f
C182 a_6465_2476# x4.x5[7].floating 0.0132f
C183 x2.x9.output_stack sample_code2[2] 0.322f
C184 sample_delay_offset x4.x3[1].floating 6.03e-20
C185 a_12839_n575# x2.x7.floating 0.00409f
C186 a_5970_n437# x3.x7.floating 0.00959f
C187 a_6130_n23# x3.x7.floating 0.00218f
C188 x3.IN sample_code2[2] 1.46e-19
C189 x1.x5[7].floating sample_code1[1] 0.0022f
C190 sample_delay_offset x1.x9.output_stack 0.262f
C191 x1.IN a_7364_1122# 1.34e-19
C192 x2.x9.output_stack x3.x6.floating 4.17e-19
C193 sample_code1[0] a_7276_1122# 6.54e-20
C194 VDD x4.x10.Y 2.7f
C195 x2.IN x2.x4[3].floating 6.65e-19
C196 x4.x2.floating a_7276_1674# 0.00177f
C197 a_5970_n713# x3.x6.SW 2.44e-19
C198 sample_delay_offset a_6058_n299# 0.00111f
C199 x3.IN x3.x6.floating 0.03f
C200 a_12767_n713# a_12839_n851# 0.00227f
C201 a_6130_n851# x3.x9.output_stack 0.0388f
C202 x1.x6.SW a_7436_1812# 2.44e-19
C203 a_12814_n2102# a_12814_n2378# 0.0316f
C204 a_6017_n2240# a_6105_n2378# 0.0704f
C205 a_567_1950# a_655_2088# 0.00227f
C206 x3.x9.output_stack x2.x2.floating 2.95e-19
C207 x3.IN a_6058_115# 1.34e-19
C208 x3.x9.output_stack sample_code2[0] 0.0111f
C209 x1.IN x4.x10.Y 1.23e-19
C210 VDD x2.x5[7].floating 44f
C211 x4.x2.floating a_7276_1122# 9.24e-19
C212 a_6749_n1036# x2.x3[1].floating 3.09e-19
C213 sample_code3[0] sample_code2[0] 1.74e-20
C214 x4.x9.output_stack x4.x5[7].floating 1.19f
C215 x1.x7.floating a_7436_1812# 0.00959f
C216 x4.x7.floating a_567_1674# 0.00409f
C217 x1.x6.SW a_7436_1260# 7.9e-20
C218 x3.x10.Y x3.x6.SW 0.788f
C219 x2.IN sample_code1[0] 0.0555f
C220 x4.x9.output_stack a_727_1812# 0.032f
C221 a_567_1674# a_655_1812# 0.00227f
C222 a_12839_n299# a_12679_n437# 0.0388f
C223 a_5970_n437# a_6058_n299# 0.00227f
C224 x2.x6.floating a_12814_n1826# 0.00996f
C225 a_680_3063# x4.x6.floating 0.0194f
C226 sample_delay_offset x4.x5[7].floating 0.00542f
C227 a_7301_3201# x4.x5[7].floating 4.61e-19
C228 sample_delay_offset a_7301_2925# 0.00273f
C229 x1.x10.Y x1.x2.floating 0.00202f
C230 sample_delay_offset a_727_1812# 0.0155f
C231 a_7301_3201# a_7301_2925# 0.0316f
C232 x3.x3[1].floating x3.x10.Y 0.00302f
C233 sample_code2[1] x2.x3[1].floating 0.226f
C234 sample_code2[0] x2.x4[3].floating 2.28e-21
C235 VDD a_12726_n1964# 0.0737f
C236 x2.IN a_12767_n299# 3.4e-19
C237 x1.x7.floating a_7436_1260# 0.00925f
C238 x4.x7.floating a_567_1122# 0.00218f
C239 a_6749_n1036# x3.x7.floating 7.29e-19
C240 sample_delay_offset x3.x9.output_stack 0.261f
C241 x4.x2.floating a_7364_2088# 2.02e-19
C242 x2.x10.Y x2.x5[7].floating 1.01f
C243 a_6465_2135# a_7276_1950# 0.00348f
C244 x3.x9.output_stack a_40_n1036# 0.00892f
C245 x4.x9.output_stack a_727_1260# 8.05e-20
C246 x2.IN x2.x9.output_stack 0.371f
C247 a_567_1398# a_655_1536# 0.00227f
C248 sample_delay_offset sample_code3[0] 0.00152f
C249 a_12679_n161# x2.x7.floating 0.00925f
C250 a_40_n1036# sample_code3[0] 0.00169f
C251 x4.x7.floating sample_code1[1] 1.73e-20
C252 sample_delay_offset a_6749_n1239# 0.00117f
C253 sample_delay_offset a_727_1260# 0.0126f
C254 sample_code0[1] x4.x4[3].floating 0.0296f
C255 x3.x7.floating sample_code2[1] 1.76e-20
C256 a_12679_n437# x2.x6.floating 0.00167f
C257 sample_code3[1] sample_code2[1] 3.2e-20
C258 x4.x2.floating a_7364_1536# 2.21e-19
C259 x3.x6.floating a_6105_n2102# 0.00996f
C260 x2.x10.Y a_12726_n1964# 4.2e-19
C261 a_5970_n161# a_6130_n299# 0.0388f
C262 x4.x4[3].floating a_567_1950# 1.17e-19
C263 sample_code1[2] x1.x4[3].floating 0.527f
C264 a_567_1122# a_655_1260# 0.00227f
C265 sample_delay_offset x2.x4[3].floating 0.0137f
C266 a_5970_n437# x3.x9.output_stack 1.74e-19
C267 x2.IN a_12839_n23# 0.029f
C268 x1.x6.SW x1.x6.floating 0.13f
C269 VDD a_592_2925# 0.103f
C270 x2.x6.SW a_12814_n2102# 9.98e-20
C271 VDD a_6465_2135# 0.235f
C272 VDD x1.x2.floating 0.0486f
C273 sample_delay_offset a_6017_n1964# 3.64e-19
C274 a_6130_n851# x2.x9.output_stack 5.22e-20
C275 VDD sample_code0[2] 0.0374f
C276 x4.x9.output_stack sample_code1[0] 2.42e-20
C277 x3.IN a_6130_n851# 0.0217f
C278 x3.x3[1].floating x3.x4[3].floating 1.19f
C279 x1.x4[3].floating a_7436_1536# 8.29e-19
C280 x2.x9.output_stack x2.x2.floating 0.193f
C281 x4.x4[3].floating a_567_1398# 1.17e-19
C282 x2.x9.output_stack sample_code2[0] 0.028f
C283 x1.x6.floating x1.x7.floating 0.202f
C284 x3.IN x2.x2.floating 0.0257f
C285 x3.IN sample_code2[0] 0.018f
C286 x4.x6.floating x4.x5[7].floating 1.18f
C287 sample_delay_offset sample_code1[0] 6.98f
C288 x1.IN a_6465_2135# 0.158f
C289 x4.x6.floating a_727_1812# 0.00278f
C290 x4.x9.output_stack x4.x2.floating 0.193f
C291 a_7276_1950# a_7436_1812# 0.0388f
C292 a_6058_n851# x3.x7.floating 8.52e-19
C293 x4.x6.SW x4.x5[7].floating 0.00138f
C294 sample_code1[2] a_7276_1674# 9.19e-20
C295 sample_delay_offset a_12767_n299# 0.00111f
C296 a_7389_3339# x1.x6.floating 0.0191f
C297 sample_code0[0] x4.x3[1].floating 0.0424f
C298 x1.x9.output_stack x1.x3[1].floating 0.341f
C299 x4.x6.SW a_727_1812# 2.44e-19
C300 a_7389_3063# sample_delay_offset 3.64e-19
C301 x1.IN a_7364_1674# 5.05e-19
C302 a_7301_3201# a_7389_3063# 0.0704f
C303 a_12726_n2240# a_12814_n2378# 0.0704f
C304 sample_delay_offset x4.x2.floating 0.0039f
C305 sample_delay_offset x2.x9.output_stack 0.264f
C306 x2.x5[7].floating x2.x6.floating 1.18f
C307 x4.x6.floating a_727_1260# 0.00109f
C308 x3.x9.output_stack a_6749_n1036# 6.54e-19
C309 sample_delay_offset x3.IN 0.258f
C310 sample_code1[2] a_7276_1122# 0.00747f
C311 a_7276_1674# a_7436_1536# 0.0388f
C312 sample_code1[0] a_6130_n23# 2.97e-20
C313 x2.x3[1].floating x2.x5[7].floating 0.8f
C314 x4.x6.SW a_727_1260# 7.9e-20
C315 a_6749_n1036# a_6749_n1239# 0.0121f
C316 x3.x2.floating sample_code2[2] 1.63e-20
C317 a_592_3477# a_680_3339# 0.0704f
C318 sample_code3[2] x3.x3[1].floating 0.00838f
C319 x2.x6.floating a_12726_n1964# 0.0194f
C320 a_12839_n851# x2.x4[3].floating 1.17e-19
C321 x3.x9.output_stack sample_code2[1] 4.73e-20
C322 a_5970_n713# x3.x4[3].floating 8.29e-19
C323 a_7276_1398# a_7436_1260# 0.0388f
C324 sample_delay_offset a_12839_n23# 0.00232f
C325 a_680_3063# x4.x10.Y 4.2e-19
C326 VDD a_12814_n2102# 0.0343f
C327 out x3.x10.Y 1.13e-19
C328 sample_code3[0] sample_code2[1] 1.6e-20
C329 x3.IN a_5970_n437# 0.0135f
C330 sample_code1[2] a_7364_2088# 8.1e-20
C331 sample_code0[2] a_655_1950# 1.36e-19
C332 x3.IN a_6130_n23# 0.0127f
C333 x2.IN a_13174_2135# 0.244f
C334 x4.x5[7].floating sample_code0[0] 0.00131f
C335 x1.IN a_7436_1812# 0.0135f
C336 x4.x10.Y x4.x3[1].floating 0.00302f
C337 x4.x7.floating a_655_1812# 8.52e-19
C338 x2.x5[7].floating a_6105_n1826# 1.79e-19
C339 sample_code1[1] x1.x4[3].floating 0.0226f
C340 x3.x4[3].floating x3.x10.Y 0.00668f
C341 sample_code2[1] x2.x4[3].floating 0.00929f
C342 a_727_1812# a_727_1536# 0.0316f
C343 a_7436_1812# a_7364_1812# 0.00227f
C344 sample_code1[2] a_7364_1536# 2.32e-19
C345 x1.x10.Y x1.x6.floating 0.0881f
C346 sample_code0[2] a_655_1398# 5.52e-19
C347 x3.x6.floating a_6017_n2240# 0.0191f
C348 x2.x10.Y a_12814_n2102# 2.35e-19
C349 sample_code1[0] a_6749_n1036# 3.76e-21
C350 a_6130_n299# x3.x6.SW 4.74e-20
C351 VDD sample_code0[1] 0.0182f
C352 a_567_1122# sample_code2[2] 2.86e-20
C353 a_12839_n575# a_12767_n575# 0.00227f
C354 x1.IN a_7436_1260# 0.0135f
C355 a_6130_n575# a_6130_n851# 0.0316f
C356 sample_delay_offset a_7364_1950# 0.00155f
C357 x4.x7.floating a_655_1260# 8.52e-19
C358 VDD a_567_1950# 0.00115f
C359 sample_delay_offset a_6105_n2102# 6.38e-19
C360 a_6130_n575# x2.x2.floating 0.00177f
C361 a_6130_n575# sample_code2[0] 0.00663f
C362 a_12839_n851# x2.x9.output_stack 0.0388f
C363 x3.x9.output_stack a_6058_n851# 0.00227f
C364 a_7436_1536# a_7364_1536# 0.00227f
C365 a_727_1536# a_727_1260# 0.0316f
C366 x2.x9.output_stack a_6749_n1036# 0.00892f
C367 x1.IN sample_code0[1] 5.47e-22
C368 x1.x5[7].floating x1.x4[3].floating 1.55f
C369 sample_delay_offset a_7364_1398# 0.00103f
C370 x3.IN a_6749_n1036# 0.157f
C371 a_12767_n575# x2.x7.floating 8.52e-19
C372 x4.x10.Y x4.x5[7].floating 1.01f
C373 a_12679_n437# x2.x4[3].floating 8.29e-19
C374 a_6058_n437# x3.x7.floating 8.52e-19
C375 a_7436_1260# a_7364_1260# 0.00227f
C376 VDD x1.x6.floating 5.87f
C377 x4.x9.output_stack sample_code1[2] 0.00469f
C378 VDD x3.x6.SW 0.45f
C379 x2.x9.output_stack sample_code2[1] 0.0705f
C380 sample_code1[0] x1.x3[1].floating 0.0394f
C381 sample_delay_offset a_6130_n575# 0.00378f
C382 sample_code0[0] sample_code1[0] 1.46e-20
C383 a_6058_n23# x2.x2.floating 2.21e-19
C384 x3.IN sample_code2[1] 1.94e-19
C385 a_6058_n23# sample_code2[0] 5.2e-19
C386 sample_code2[2] x2.x7.floating 0.0056f
C387 x2.x9.output_stack a_12814_n1826# 0.0702f
C388 sample_code1[1] a_7276_1122# 8.94e-20
C389 a_680_3063# a_592_2925# 0.0704f
C390 sample_code3[2] x3.x10.Y 0.00203f
C391 sample_delay_offset sample_code1[2] 0.0966f
C392 VDD x3.x3[1].floating 0.0301f
C393 x1.IN x1.x6.floating 0.03f
C394 x3.x9.output_stack x2.x5[7].floating 1.33e-19
C395 sample_code2[0] x3.x2.floating 1.9e-20
C396 x3.x6.SW x2.x10.Y 1.5e-20
C397 x4.x3[1].floating a_6465_2135# 3.09e-19
C398 sample_code0[2] x4.x3[1].floating 0.00115f
C399 a_5970_n161# x3.x7.floating 0.00925f
C400 sample_code0[0] x4.x2.floating 0.164f
C401 x1.x6.SW x1.x7.floating 9.72e-19
C402 x1.x9.output_stack x1.x2.floating 0.193f
C403 sample_delay_offset a_7436_1536# 0.0133f
C404 x1.x9.output_stack a_6465_2135# 6.54e-19
C405 a_5970_n437# a_6130_n575# 0.0388f
C406 a_12679_n437# a_12767_n299# 0.00227f
C407 x2.x6.floating a_12814_n2102# 0.00996f
C408 a_6749_n1239# x2.x5[7].floating 0.0132f
C409 sample_delay_offset a_6058_n23# 9.64e-19
C410 a_12679_n437# x2.x9.output_stack 1.74e-19
C411 VDD a_12726_n2240# 0.129f
C412 x2.IN sample_code1[1] 5.47e-22
C413 x2.IN a_12839_n575# 0.03f
C414 sample_code1[2] a_6130_n23# 2.07e-20
C415 a_567_1950# a_655_1950# 0.00227f
C416 VDD a_680_3339# 0.128f
C417 x2.x4[3].floating x2.x5[7].floating 1.55f
C418 x3.IN a_6058_n851# 0.00196f
C419 sample_delay_offset x3.x2.floating 0.00186f
C420 sample_code3[2] x3.x4[3].floating 0.536f
C421 a_40_n1036# x3.x2.floating 0.0104f
C422 a_6130_n299# x3.x10.Y 4.07e-20
C423 a_12767_n161# x2.x7.floating 8.52e-19
C424 a_567_1122# sample_code2[0] 2e-20
C425 a_567_1674# a_655_1674# 0.00227f
C426 x2.x10.Y a_12726_n2240# 1.49e-19
C427 x3.x6.floating a_6105_n2378# 0.00578f
C428 x2.IN x2.x7.floating 0.0261f
C429 a_6130_n23# a_6058_n23# 0.00227f
C430 a_592_2925# x4.x5[7].floating 2.76e-19
C431 a_5970_n713# a_6058_n713# 0.00227f
C432 x4.x6.floating sample_code1[2] 3.95e-22
C433 x2.IN x1.x5[7].floating 0.0199f
C434 x4.x5[7].floating sample_code0[2] 0.00564f
C435 sample_delay_offset a_567_1674# 0.00384f
C436 x2.x6.SW a_12814_n2378# 5.11e-20
C437 x4.x10.Y x4.x2.floating 0.00202f
C438 sample_delay_offset a_6017_n2240# 1.9e-19
C439 a_567_1398# a_655_1398# 0.00227f
C440 a_7301_3477# sample_delay_offset 3.28e-19
C441 x4.x6.SW sample_code1[2] 3.93e-21
C442 a_7301_3477# a_7301_3201# 0.0316f
C443 x1.x9.output_stack a_7436_1812# 0.032f
C444 sample_delay_offset a_567_1122# 0.0025f
C445 x2.x9.output_stack x2.x5[7].floating 1.19f
C446 x4.x9.output_stack sample_code1[1] 4.64e-20
C447 VDD x3.x10.Y 2.73f
C448 a_12679_n161# a_12767_n161# 0.00227f
C449 a_12767_115# a_12839_n23# 0.0022f
C450 x3.IN x2.x5[7].floating 0.0216f
C451 a_567_1122# a_655_1122# 0.0022f
C452 a_6130_n299# x3.x4[3].floating 1.17e-19
C453 a_5970_n161# x3.x9.output_stack 8.05e-20
C454 sample_delay_offset sample_code1[1] 0.0596f
C455 a_12679_n713# x2.x6.SW 2.44e-19
C456 x2.IN a_12679_n161# 0.0166f
C457 VDD a_655_2088# 1.29e-19
C458 x1.x10.Y x1.x6.SW 0.788f
C459 x1.x9.output_stack a_7436_1260# 8.05e-20
C460 sample_delay_offset a_12839_n575# 0.00382f
C461 x3.x10.Y a_40_n1239# 0.00127f
C462 x1.x6.SW a_7276_1950# 0.00179f
C463 x2.x9.output_stack a_12726_n1964# 0.032f
C464 VDD out 0.244f
C465 x3.x10.Y x2.x10.Y 1.79e-20
C466 sample_code0[1] x4.x3[1].floating 0.227f
C467 x1.x10.Y x1.x7.floating 0.00345f
C468 x1.x7.floating a_7276_1950# 0.00409f
C469 x1.x3[1].floating a_13174_2135# 3.09e-19
C470 sample_code1[2] x1.x3[1].floating 0.00115f
C471 sample_code1[0] x1.x2.floating 0.163f
C472 x1.x6.SW a_7276_1398# 4.74e-20
C473 a_6465_2135# sample_code1[0] 8.82e-21
C474 sample_code0[2] sample_code1[0] 5.83e-20
C475 sample_code0[0] sample_code1[2] 3.13f
C476 x3.x7.floating x3.x6.SW 9.72e-19
C477 sample_delay_offset x2.x7.floating 0.264f
C478 sample_code1[1] a_6130_n23# 2.46e-20
C479 out a_40_n1239# 0.145f
C480 x2.x6.floating a_12726_n2240# 0.0191f
C481 x3.x6.SW a_6105_n1826# 0.00707f
C482 sample_delay_offset x1.x5[7].floating 0.00308f
C483 VDD x3.x4[3].floating 0.0565f
C484 a_7301_3201# x1.x5[7].floating 2.76e-19
C485 a_7389_3339# x1.x10.Y 1.49e-19
C486 VDD a_12814_n2378# 0.112f
C487 x4.x6.SW a_567_1674# 8.11e-20
C488 VDD x1.x6.SW 0.452f
C489 x3.x2.floating sample_code2[1] 1.76e-20
C490 x1.x7.floating a_7276_1398# 0.00409f
C491 sample_code3[1] x3.x3[1].floating 0.23f
C492 x3.IN a_6058_n437# 5.05e-19
C493 x3.x6.SW x3.x5[7].floating 0.00138f
C494 x4.x2.floating a_6465_2135# 0.0104f
C495 sample_code1[2] a_7364_1122# 7.9e-19
C496 x2.x5[7].floating a_6105_n2102# 1.94e-19
C497 x1.x9.output_stack x1.x6.floating 0.229f
C498 VDD a_592_3477# 0.109f
C499 VDD x1.x7.floating 0.0315f
C500 x1.IN x1.x6.SW 0.0933f
C501 x4.x6.SW a_567_1122# 3.1e-20
C502 VDD x4.x4[3].floating 0.0565f
C503 x3.x3[1].floating x3.x5[7].floating 0.8f
C504 x4.x5[7].floating sample_code0[1] 0.00228f
C505 x4.x2.floating a_7364_1674# 2.21e-19
C506 x2.x10.Y a_12814_n2378# 1.02e-19
C507 sample_delay_offset a_12679_n161# 0.0124f
C508 a_12839_n575# a_12839_n851# 0.0316f
C509 x4.x10.Y sample_code1[2] 2.74e-20
C510 x1.IN x1.x7.floating 0.0242f
C511 a_567_1950# a_727_1812# 0.0388f
C512 x3.IN a_5970_n161# 0.0135f
C513 VDD a_7389_3339# 0.138f
C514 a_6058_n575# x2.x2.floating 2.21e-19
C515 sample_delay_offset a_6105_n2378# 3.28e-19
C516 a_6058_n575# sample_code2[0] 1.32e-19
C517 a_567_1122# sample_code2[1] 2.37e-20
C518 a_680_3339# a_680_3063# 0.0316f
C519 x4.x9.output_stack x4.x7.floating 0.185f
C520 x1.x7.floating a_7364_1812# 8.52e-19
C521 x1.x4[3].floating a_7276_1674# 1.17e-19
C522 x4.x7.floating a_655_1674# 8.52e-19
C523 VDD sample_code3[2] 0.0374f
C524 x4.x5[7].floating x1.x6.floating 0.0269f
C525 a_567_1674# a_727_1536# 0.0388f
C526 x1.IN a_7389_3339# 0.00847f
C527 a_12839_n851# x2.x7.floating 0.00409f
C528 sample_delay_offset x4.x7.floating 0.259f
C529 a_7301_2925# x1.x6.floating 0.00996f
C530 a_5970_n713# x3.x7.floating 0.00959f
C531 x1.x10.Y a_7276_1950# 1.69e-19
C532 x1.x7.floating a_7364_1260# 8.52e-19
C533 VDD x2.x6.SW 0.43f
C534 x1.x4[3].floating a_7276_1122# 7.17e-20
C535 sample_delay_offset a_655_1812# 0.00138f
C536 sample_code0[0] a_567_1122# 1.99e-19
C537 x3.x9.output_stack x3.x6.SW 0.164f
C538 x4.x2.floating a_7436_1812# 6.24e-19
C539 sample_delay_offset a_6058_n575# 0.00138f
C540 a_567_1398# a_727_1260# 0.0388f
C541 sample_code1[1] x1.x3[1].floating 0.224f
C542 x3.x9.output_stack x3.x3[1].floating 0.341f
C543 x3.x6.SW a_6749_n1239# 0.00208f
C544 x1.x10.Y a_7276_1398# 4.07e-20
C545 sample_code0[1] sample_code1[0] 2.91e-20
C546 sample_code0[0] sample_code1[1] 1.58e-20
C547 sample_delay_offset a_655_1260# 9.69e-19
C548 x3.x7.floating x3.x10.Y 0.00345f
C549 sample_code3[1] x3.x10.Y 6.71e-19
C550 x4.x2.floating a_7436_1260# 6.88e-19
C551 sample_code3[0] x3.x3[1].floating 0.0326f
C552 x3.x10.Y a_6105_n1826# 0.039f
C553 x2.x10.Y x2.x6.SW 0.788f
C554 a_7276_1122# sample_code2[2] 2.86e-20
C555 x4.x10.Y a_567_1674# 6.65e-20
C556 a_6058_n437# a_6130_n575# 0.00227f
C557 a_12679_n437# a_12839_n575# 0.0388f
C558 x2.x6.floating a_12814_n2378# 0.00578f
C559 VDD x1.x10.Y 2.73f
C560 VDD a_7276_1950# 0.00115f
C561 a_680_3339# x4.x5[7].floating 0.00154f
C562 a_6058_n161# x2.x2.floating 2.21e-19
C563 x3.x10.Y x3.x5[7].floating 1.01f
C564 a_6058_n161# sample_code2[0] 3.43e-19
C565 sample_code0[1] x4.x2.floating 0.0027f
C566 x2.IN a_12767_n575# 7.93e-19
C567 out sample_code3[1] 5.47e-22
C568 x1.x2.floating a_13174_2135# 0.0104f
C569 a_6465_2135# sample_code1[2] 0.00525f
C570 x1.x5[7].floating x1.x3[1].floating 0.8f
C571 x4.x10.Y a_567_1122# 2.2e-20
C572 sample_code0[2] sample_code1[2] 6.83e-20
C573 x1.IN x1.x10.Y 0.0967f
C574 x4.x6.floating x4.x7.floating 0.202f
C575 x2.x5[7].floating a_6017_n2240# 8.4e-20
C576 x1.IN a_7276_1950# 0.0217f
C577 a_12679_n437# x2.x7.floating 0.00959f
C578 x3.x4[3].floating x3.x7.floating 1.18f
C579 out x3.x5[7].floating 0.0199f
C580 sample_code3[1] x3.x4[3].floating 0.00929f
C581 x4.x6.SW x4.x7.floating 9.72e-19
C582 a_12679_n713# x2.x6.floating 0.00278f
C583 a_7364_1950# a_7436_1812# 0.00227f
C584 sample_code1[2] a_7364_1674# 1.7e-19
C585 a_12839_n299# x2.x6.SW 4.74e-20
C586 a_7389_3063# x1.x6.floating 0.0194f
C587 sample_delay_offset a_6058_n161# 0.00102f
C588 a_5970_n713# x3.x9.output_stack 0.032f
C589 a_12679_n713# a_12767_n713# 0.00227f
C590 x1.IN a_7276_1398# 0.0136f
C591 x2.x9.output_stack x3.x6.SW 3.62e-19
C592 VDD a_12767_n851# 1.29e-19
C593 x3.IN x3.x6.SW 0.0933f
C594 x3.x4[3].floating x3.x5[7].floating 1.55f
C595 a_7364_1674# a_7436_1536# 0.00227f
C596 VDD a_40_n1239# 0.211f
C597 VDD x1.IN 0.613f
C598 sample_code2[2] x2.x2.floating 1.63e-20
C599 sample_code2[0] sample_code2[2] 1.48e-20
C600 VDD x2.x10.Y 2.71f
C601 sample_delay_offset x1.x4[3].floating 0.00732f
C602 a_12679_n161# a_12679_n437# 0.0316f
C603 a_5970_n161# a_6058_n23# 0.00227f
C604 x2.x6.SW x2.x6.floating 0.13f
C605 x3.x9.output_stack x3.x10.Y 1.01f
C606 x1.x6.SW x1.x9.output_stack 0.164f
C607 a_7364_1398# a_7436_1260# 0.00227f
C608 sample_code2[0] x3.x6.floating 1.3e-21
C609 sample_code3[0] x3.x10.Y 0.0124f
C610 x2.IN a_12767_n161# 2.42e-19
C611 sample_code0[2] a_567_1674# 1.33e-19
C612 sample_delay_offset a_12767_n575# 0.00138f
C613 x3.x10.Y a_6749_n1239# 6.93e-19
C614 x2.x7.floating x2.x5[7].floating 0.182f
C615 x4.x9.output_stack sample_code2[2] 4.06e-21
C616 x4.x4[3].floating x4.x3[1].floating 1.19f
C617 sample_code0[0] x4.x7.floating 2.03e-20
C618 x2.x9.output_stack a_12726_n2240# 1.5e-19
C619 x1.x9.output_stack x1.x7.floating 0.185f
C620 a_6058_115# sample_code2[0] 8.2e-19
C621 a_592_3201# sample_delay_offset 6.38e-19
C622 x1.IN a_7364_1812# 7.93e-19
C623 sample_code3[2] x3.x7.floating 0.0056f
C624 x4.x7.floating a_727_1536# 0.00959f
C625 sample_code3[1] sample_code3[2] 0.882f
C626 x3.x9.output_stack out 0.127f
C627 a_7276_1122# sample_code2[0] 2e-20
C628 sample_delay_offset sample_code2[2] 6.08f
C629 a_7436_1812# a_7436_1536# 0.0316f
C630 x1.x10.Y a_13174_2476# 0.00127f
C631 sample_code0[2] a_567_1122# 0.0177f
C632 sample_code3[0] out 1.07e-19
C633 x3.x10.Y a_6017_n1964# 4.2e-19
C634 a_7389_3339# x1.x9.output_stack 1.5e-19
C635 sample_delay_offset x3.x6.floating 0.0706f
C636 x1.IN a_7364_1260# 1.8e-19
C637 VDD a_12839_n299# 4.84e-19
C638 sample_delay_offset a_7276_1674# 0.00384f
C639 sample_code3[2] x3.x5[7].floating 0.00568f
C640 x1.x6.SW x4.x5[7].floating 0.00313f
C641 x3.x6.SW a_6105_n2102# 9.98e-20
C642 x3.x9.output_stack x3.x4[3].floating 0.636f
C643 sample_code1[1] x1.x2.floating 0.0027f
C644 a_6465_2135# sample_code1[1] 9.55e-21
C645 a_7301_2925# x1.x6.SW 0.00707f
C646 sample_delay_offset a_6058_115# 5.66e-19
C647 sample_code0[2] sample_code1[1] 6.3e-20
C648 sample_code0[1] sample_code1[2] 3.42e-20
C649 a_7436_1536# a_7436_1260# 0.0316f
C650 x3.IN a_5970_n713# 0.0135f
C651 sample_code3[0] x3.x4[3].floating 2.28e-21
C652 a_592_3477# x4.x5[7].floating 2.14e-19
C653 sample_delay_offset a_7276_1122# 0.0025f
C654 a_6130_n23# sample_code2[2] 6.93e-20
C655 x4.x5[7].floating x4.x4[3].floating 1.55f
C656 x2.x5[7].floating a_6105_n2378# 3.13e-19
C657 a_5970_n437# x3.x6.floating 0.00167f
C658 a_12839_n299# x2.x10.Y 4.07e-20
C659 x4.x10.Y x4.x7.floating 0.00345f
C660 x4.x4[3].floating a_727_1812# 8.29e-19
C661 a_6130_n299# x3.x7.floating 0.00409f
C662 VDD a_13174_2476# 0.217f
C663 VDD x2.x6.floating 5.78f
C664 x2.x9.output_stack x3.x10.Y 1.93e-19
C665 a_6058_115# a_6130_n23# 0.0022f
C666 a_6130_n575# x3.x6.SW 8.11e-20
C667 sample_delay_offset a_12767_n161# 0.00103f
C668 a_592_3201# x4.x6.floating 0.00996f
C669 a_7389_3339# x4.x5[7].floating 1.78e-19
C670 x1.x5[7].floating x1.x2.floating 0.441f
C671 x3.IN x3.x10.Y 0.0967f
C672 x1.x6.floating sample_code1[2] 3.95e-22
C673 sample_delay_offset a_7364_2088# 0.00167f
C674 x4.x4[3].floating a_727_1260# 7.47e-19
C675 VDD x2.x3[1].floating 0.0301f
C676 a_6130_n851# x2.x2.floating 8.75e-19
C677 sample_delay_offset x2.IN 0.27f
C678 a_6130_n851# sample_code2[0] 0.00186f
C679 a_592_3201# x4.x6.SW 9.98e-20
C680 sample_code2[0] x2.x2.floating 0.167f
C681 x1.x10.Y x1.x9.output_stack 1.01f
C682 x2.x10.Y x2.x6.floating 0.0881f
C683 x4.x9.output_stack a_6465_2476# 0.00887f
C684 x3.x9.output_stack sample_code3[2] 0.334f
C685 x1.x6.floating a_7436_1536# 0.00167f
C686 x1.x9.output_stack a_7276_1950# 0.0388f
C687 sample_delay_offset a_7364_1536# 0.00111f
C688 a_6749_n1036# sample_code2[2] 8.96e-21
C689 a_6130_n299# a_6058_n299# 0.00227f
C690 a_12679_n713# x2.x4[3].floating 8.29e-19
C691 sample_code3[0] sample_code3[2] 1.89e-20
C692 VDD x3.x7.floating 0.0315f
C693 a_6058_n713# x3.x7.floating 8.52e-19
C694 VDD sample_code3[1] 0.0182f
C695 sample_delay_offset a_6465_2476# 0.00117f
C696 x2.x3[1].floating x2.x10.Y 0.00302f
C697 VDD a_6105_n1826# 0.11f
C698 a_567_1950# a_567_1674# 0.0316f
C699 VDD a_680_3063# 0.0732f
C700 sample_delay_offset a_6130_n851# 0.0189f
C701 sample_code1[0] x1.x7.floating 1.61e-20
C702 x1.x4[3].floating x1.x3[1].floating 1.19f
C703 x4.x4[3].floating sample_code1[0] 6.43e-20
C704 sample_delay_offset x2.x2.floating 0.00558f
C705 x3.IN x3.x4[3].floating 6.65e-19
C706 sample_code2[1] sample_code2[2] 4.67f
C707 sample_delay_offset sample_code2[0] 0.0609f
C708 VDD x3.x5[7].floating 43.9f
C709 sample_code0[1] a_567_1122# 3.36e-19
C710 VDD x4.x3[1].floating 0.0301f
C711 a_567_1674# a_567_1398# 0.0316f
C712 x3.x2.floating x3.x3[1].floating 1.17f
C713 VDD x1.x9.output_stack 0.596f
C714 x1.x10.Y x4.x5[7].floating 0.00422f
C715 x3.x10.Y a_6105_n2102# 2.35e-19
C716 a_12839_n23# a_12767_n23# 0.00227f
C717 x4.x2.floating x1.x7.floating 0.0475f
C718 a_7301_2925# x1.x10.Y 0.039f
C719 a_40_n1239# x3.x5[7].floating 0.0132f
C720 sample_code0[1] sample_code1[1] 3.15e-20
C721 sample_code0[2] x4.x7.floating 0.0173f
C722 sample_delay_offset x4.x9.output_stack 0.263f
C723 sample_delay_offset a_655_1674# 0.00123f
C724 a_6130_n575# a_5970_n713# 0.0388f
C725 a_12767_n437# a_12839_n575# 0.00227f
C726 sample_code0[2] a_655_1812# 1.81e-19
C727 a_5970_n437# x2.x2.floating 6.88e-19
C728 a_7301_3477# x1.x6.floating 0.00578f
C729 a_6130_n23# x2.x2.floating 9.24e-19
C730 a_12679_n713# x2.x9.output_stack 0.032f
C731 a_6130_n23# sample_code2[0] 0.0131f
C732 x1.IN x1.x9.output_stack 0.371f
C733 a_567_1398# a_567_1122# 0.0316f
C734 a_7276_1122# sample_code2[1] 2.37e-20
C735 x2.IN a_12839_n851# 0.038f
C736 a_7389_3339# a_7389_3063# 0.0316f
C737 a_7301_3201# sample_delay_offset 6.38e-19
C738 sample_code0[0] a_7276_1674# 0.00654f
C739 sample_delay_offset a_655_1122# 5.69e-19
C740 sample_code0[2] a_655_1260# 8.73e-19
C741 a_6130_n575# x3.x10.Y 6.65e-20
C742 a_12767_n437# x2.x7.floating 8.52e-19
C743 VDD x4.x5[7].floating 44f
C744 VDD a_7301_2925# 0.11f
C745 sample_code0[0] a_7276_1122# 0.00533f
C746 sample_delay_offset a_5970_n437# 0.0128f
C747 sample_delay_offset a_6130_n23# 0.00246f
C748 VDD x3.x9.output_stack 0.595f
C749 a_592_3201# x4.x10.Y 2.35e-19
C750 x2.x9.output_stack x2.x6.SW 0.164f
C751 x2.IN a_12814_n1826# 0.0175f
C752 VDD sample_code3[0] 0.00326f
C753 a_6130_n851# a_6749_n1036# 0.00348f
C754 x1.IN x4.x5[7].floating 0.0218f
C755 x1.x10.Y sample_code1[0] 0.0124f
C756 x1.IN a_7301_2925# 0.0175f
C757 VDD a_6749_n1239# 0.212f
C758 x3.x9.output_stack a_40_n1239# 0.00887f
C759 a_6749_n1036# x2.x2.floating 0.0104f
C760 x4.x9.output_stack x4.x6.floating 0.229f
C761 a_6749_n1036# sample_code2[0] 0.00699f
C762 x1.x7.floating a_7364_1950# 8.52e-19
C763 a_7276_1122# a_7364_1122# 0.0022f
C764 x1.x6.floating x1.x5[7].floating 1.18f
C765 VDD x2.x4[3].floating 0.0565f
C766 a_12839_n23# x2.x6.SW 3.1e-20
C767 sample_delay_offset x4.x6.floating 0.0706f
C768 a_6130_n575# x3.x4[3].floating 1.17e-19
C769 a_7389_3063# x1.x10.Y 4.2e-19
C770 x4.x6.SW x4.x9.output_stack 0.164f
C771 sample_code2[2] x2.x5[7].floating 0.0056f
C772 VDD a_6017_n1964# 0.0801f
C773 x3.x2.floating x3.x10.Y 0.00202f
C774 sample_code2[1] x2.x2.floating 0.00516f
C775 x1.x7.floating a_7364_1398# 8.52e-19
C776 sample_code2[0] sample_code2[1] 4.25f
C777 x2.IN a_12679_n437# 0.0166f
C778 x3.x6.floating x2.x5[7].floating 0.0231f
C779 x2.x10.Y a_6749_n1239# 0.00127f
C780 x3.IN a_6130_n299# 0.0136f
C781 x4.x2.floating a_7276_1950# 8.75e-19
C782 sample_delay_offset a_12839_n851# 0.0189f
C783 sample_delay_offset x4.x6.SW 0.19f
C784 x1.x6.SW sample_code1[2] 3.93e-21
C785 sample_delay_offset a_6749_n1036# 0.00652f
C786 x1.x9.output_stack a_13174_2476# 0.00887f
C787 VDD sample_code1[0] 0.00346f
C788 x2.x4[3].floating x2.x10.Y 0.00668f
C789 sample_code0[1] x4.x7.floating 2.21e-20
C790 x4.x9.output_stack sample_code2[1] 9.58e-22
C791 x4.x2.floating a_7276_1398# 0.00177f
C792 out x3.x2.floating 0.0191f
C793 a_5970_n161# a_6058_n161# 0.00227f
C794 x3.x10.Y a_6017_n2240# 1.49e-19
C795 sample_code1[2] x1.x7.floating 0.0129f
C796 x4.x7.floating a_567_1950# 0.00409f
C797 x4.x4[3].floating sample_code1[2] 7.49e-20
C798 x1.x6.SW a_7436_1536# 1.28e-19
C799 sample_delay_offset sample_code2[1] 0.0313f
C800 x2.IN a_12767_115# 1.34e-19
C801 a_655_1950# a_727_1812# 0.00227f
C802 x1.IN sample_code1[0] 1.38e-19
C803 VDD a_7389_3063# 0.0797f
C804 x3.x6.SW a_6105_n2378# 5.11e-20
C805 VDD x2.x9.output_stack 0.595f
C806 sample_delay_offset a_12814_n1826# 0.00273f
C807 a_6130_n851# a_6058_n851# 0.00227f
C808 VDD x4.x2.floating 0.0334f
C809 x3.x7.floating x3.x5[7].floating 0.182f
C810 a_592_3201# a_592_2925# 0.0316f
C811 sample_code3[1] x3.x5[7].floating 0.00224f
C812 x1.x7.floating a_7436_1536# 0.00959f
C813 x4.x9.output_stack sample_code0[0] 0.0321f
C814 x3.IN a_6058_n713# 0.0013f
C815 VDD x3.IN 0.612f
C816 a_6058_n851# x2.x2.floating 2.02e-19
C817 x4.x7.floating a_567_1398# 0.00409f
C818 a_6058_n851# sample_code2[0] 8.23e-20
C819 x2.x9.output_stack a_12767_n851# 0.00227f
C820 x3.x5[7].floating a_6105_n1826# 2.76e-19
C821 x4.x9.output_stack a_727_1536# 1.74e-19
C822 a_655_1674# a_727_1536# 0.00227f
C823 x1.IN a_7389_3063# 0.00921f
C824 sample_delay_offset x1.x3[1].floating 3.48e-20
C825 x2.IN x2.x5[7].floating 0.00127f
C826 a_6465_2135# sample_code2[2] 3.71e-21
C827 sample_delay_offset sample_code0[0] 0.0311f
C828 x1.IN x4.x2.floating 0.0257f
C829 x4.x10.Y a_6465_2476# 0.00127f
C830 a_12839_n299# x2.x4[3].floating 1.17e-19
C831 a_6058_n299# x3.x7.floating 8.52e-19
C832 a_6130_n23# sample_code2[1] 9.56e-20
C833 sample_delay_offset a_727_1536# 0.0133f
C834 VDD a_12839_n23# 4.84e-19
C835 x2.x9.output_stack x2.x10.Y 1.01f
C836 a_7276_1950# a_7364_1950# 0.00227f
C837 x4.x6.SW x4.x6.floating 0.13f
C838 x4.x2.floating a_7364_1812# 2.21e-19
C839 x3.IN x2.x10.Y 1.23e-19
C840 sample_delay_offset a_12679_n437# 0.0132f
C841 a_655_1398# a_727_1260# 0.00227f
C842 x2.IN a_12726_n1964# 0.00921f
C843 sample_delay_offset a_6058_n851# 0.00166f
C844 sample_delay_offset a_7364_1122# 5.69e-19
C845 a_7301_3477# x1.x6.SW 5.11e-20
C846 a_7276_1674# a_7364_1674# 0.00227f
C847 x4.x2.floating a_7364_1260# 2.21e-19
C848 x1.x4[3].floating a_7436_1812# 8.29e-19
C849 a_5970_n161# x3.x6.floating 0.00109f
C850 a_12839_n23# x2.x10.Y 2.2e-20
C851 x4.x4[3].floating a_567_1674# 1.17e-19
C852 x2.x2.floating x2.x5[7].floating 0.441f
C853 x4.x10.Y x4.x9.output_stack 1.01f
C854 sample_code2[0] x2.x5[7].floating 0.00119f
C855 a_6130_n299# a_6130_n575# 0.0316f
C856 sample_code3[2] x3.x2.floating 2.06e-20
C857 a_12839_n299# a_12767_n299# 0.00227f
C858 x3.x9.output_stack x3.x7.floating 0.185f
C859 a_680_3063# x4.x5[7].floating 0.00169f
C860 x3.x9.output_stack sample_code3[1] 0.0715f
C861 sample_delay_offset a_12767_115# 5.68e-19
C862 sample_delay_offset x4.x10.Y 0.0403f
C863 x2.x3[1].floating x2.x4[3].floating 1.19f
C864 a_7276_1398# a_7364_1398# 0.00227f
C865 VDD a_6105_n2102# 0.0945f
C866 x1.x10.Y sample_code1[2] 0.00201f
C867 x3.x9.output_stack a_6105_n1826# 0.0702f
C868 x1.x4[3].floating a_7436_1260# 7.47e-19
C869 a_6749_n1036# sample_code2[1] 4.37e-20
C870 x4.x4[3].floating a_567_1122# 7.17e-20
C871 sample_code1[2] a_7276_1950# 5.6e-20
C872 sample_code3[0] sample_code3[1] 0.459f
C873 x2.IN x1.x2.floating 0.0392f
C874 x4.x5[7].floating x4.x3[1].floating 0.8f
C875 x4.x6.floating sample_code0[0] 1.18e-19
C876 a_7301_3477# a_7389_3339# 0.0704f
C877 x1.IN a_7364_1950# 0.0013f
C878 x1.x9.output_stack x4.x5[7].floating 1.33e-19
C879 x3.x9.output_stack x3.x5[7].floating 1.19f
C880 sample_code1[1] x1.x7.floating 1.73e-20
C881 a_12767_n23# x2.x7.floating 8.52e-19
C882 x4.x6.floating a_727_1536# 0.00167f
C883 a_7301_2925# x1.x9.output_stack 0.0702f
C884 x4.x4[3].floating sample_code1[1] 6.93e-20
C885 sample_delay_offset x2.x5[7].floating 0.00542f
C886 sample_code3[0] x3.x5[7].floating 0.00121f
C887 a_7436_1812# a_7276_1674# 0.0388f
C888 x4.x6.SW sample_code0[0] 4.21e-21
C889 sample_code1[2] a_7276_1398# 1.74e-19
C890 x3.x10.Y a_6105_n2378# 1.02e-19
C891 a_12839_n23# a_12839_n299# 0.0316f
C892 x4.x6.SW a_727_1536# 1.28e-19
C893 x1.IN a_7364_1398# 2.42e-19
C894 a_6465_2476# a_6465_2135# 0.0121f
C895 x2.x9.output_stack x2.x6.floating 0.229f
C896 a_567_1122# sample_code3[2] 1.71e-20
C897 a_12839_n575# a_12679_n713# 0.0388f
C898 a_5970_n713# a_6058_n575# 0.00227f
C899 a_6105_n1826# a_6017_n1964# 0.0704f
C900 x1.x6.SW x1.x5[7].floating 0.00138f
C901 VDD a_13174_2135# 0.237f
C902 a_6058_n437# x2.x2.floating 2.21e-19
C903 sample_delay_offset a_12726_n1964# 3.64e-19
C904 a_6058_n437# sample_code2[0] 1.74e-19
C905 VDD sample_code1[2] 0.0376f
C906 a_7436_1536# a_7276_1398# 0.0388f
C907 x2.x9.output_stack x2.x3[1].floating 0.341f
C908 x3.x5[7].floating a_6017_n1964# 0.00169f
C909 x1.x5[7].floating x1.x7.floating 0.182f
C910 a_12679_n161# a_12767_n23# 0.00227f
C911 a_7301_2925# x4.x5[7].floating 1.79e-19
C912 a_12679_n713# x2.x7.floating 0.00959f
C913 x4.x10.Y x4.x6.floating 0.0881f
C914 x1.IN sample_code1[2] 0.0169f
C915 x4.x7.floating a_655_2088# 8.52e-19
C916 a_7436_1260# a_7276_1122# 0.0388f
C917 a_592_2925# x4.x9.output_stack 0.0702f
C918 x4.x9.output_stack a_6465_2135# 0.00892f
C919 x4.x9.output_stack sample_code0[2] 0.334f
C920 sample_code1[2] a_7364_1812# 1.29e-19
C921 a_12839_n575# x2.x6.SW 8.11e-20
C922 x2.x9.output_stack x3.x7.floating 3.32e-19
C923 sample_code0[2] a_655_1674# 2.5e-19
C924 x4.x3[1].floating sample_code1[0] 3.21e-20
C925 sample_delay_offset a_6058_n437# 0.00122f
C926 a_7389_3339# x1.x5[7].floating 0.00154f
C927 a_5970_n161# x2.x2.floating 6.88e-19
C928 x4.x10.Y x4.x6.SW 0.788f
C929 a_7301_3477# x1.x10.Y 1.02e-19
C930 x3.IN x3.x7.floating 0.0242f
C931 x1.x9.output_stack sample_code1[0] 0.0244f
C932 a_592_2925# sample_delay_offset 0.00273f
C933 x1.IN a_7436_1536# 0.0135f
C934 sample_delay_offset x1.x2.floating 0.00286f
C935 x2.IN a_12814_n2102# 0.00866f
C936 sample_delay_offset a_6465_2135# 0.00651f
C937 x3.IN a_6105_n1826# 0.0175f
C938 x4.x7.floating a_655_1536# 8.52e-19
C939 sample_delay_offset sample_code0[2] 0.0694f
C940 VDD x3.x2.floating 0.0334f
C941 x3.x9.output_stack sample_code3[0] 0.0285f
C942 sample_code1[2] a_7364_1260# 5.02e-19
C943 x3.x9.output_stack a_6749_n1239# 1.18e-20
C944 sample_code0[2] a_655_1122# 0.0013f
C945 x2.x7.floating x2.x6.SW 9.72e-19
C946 x3.x6.SW x3.x6.floating 0.13f
C947 x3.IN x3.x5[7].floating 0.00127f
C948 x4.x3[1].floating x4.x2.floating 1.17f
C949 a_7389_3063# x1.x9.output_stack 0.032f
C950 sample_delay_offset a_7364_1674# 0.00123f
C951 x1.x10.Y sample_code1[1] 6.64e-19
C952 x3.x3[1].floating sample_code2[2] 3.26e-20
C953 x1.x9.output_stack x4.x2.floating 2.95e-19
C954 a_5970_n437# a_6058_n437# 0.00227f
C955 sample_delay_offset a_5970_n161# 0.0121f
C956 VDD a_6017_n2240# 0.138f
C957 x3.x9.output_stack a_6017_n1964# 0.032f
C958 x2.IN a_12767_n437# 5.05e-19
C959 VDD a_7301_3477# 0.179f
C960 x3.IN a_6058_n299# 3.4e-19
C961 sample_code2[1] x2.x5[7].floating 0.0022f
C962 x4.x7.floating x4.x4[3].floating 1.18f
C963 a_680_3339# a_592_3201# 0.0704f
C964 x2.x5[7].floating a_12814_n1826# 2.76e-19
C965 x4.x10.Y sample_code0[0] 0.0125f
C966 sample_code1[0] x3.x9.output_stack 4.11e-21
C967 x1.IN a_7301_3477# 0.00832f
C968 x1.x10.Y x1.x5[7].floating 1.01f
C969 a_5970_n161# a_5970_n437# 0.0316f
C970 a_12679_n161# x2.x6.SW 7.9e-20
C971 a_6130_n23# a_5970_n161# 0.0388f
C972 a_592_2925# x4.x6.floating 0.00996f
C973 a_7389_3063# x4.x5[7].floating 4.88e-20
C974 VDD sample_code1[1] 0.0183f
C975 a_13174_2476# a_13174_2135# 0.0121f
C976 VDD a_12839_n575# 4.84e-19
C977 a_7389_3063# a_7301_2925# 0.0704f
C978 x4.x5[7].floating x4.x2.floating 0.441f
C979 x4.x6.floating sample_code0[2] 1.36e-19
C980 sample_delay_offset a_7436_1812# 0.0155f
C981 a_6105_n1826# a_6105_n2102# 0.0316f
C982 a_12814_n1826# a_12726_n1964# 0.0704f
C983 sample_delay_offset a_12814_n2102# 6.38e-19
C984 x3.x9.output_stack x2.x9.output_stack 2.93e-20
C985 a_592_2925# x4.x6.SW 0.00707f
C986 x3.IN x3.x9.output_stack 0.371f
C987 x4.x6.SW sample_code0[2] 9.76e-21
C988 x3.x5[7].floating a_6105_n2102# 2.76e-19
C989 x1.IN sample_code1[1] 1.86e-19
C990 sample_delay_offset a_7436_1260# 0.0126f
C991 x2.x9.output_stack a_6749_n1239# 0.00887f
C992 a_6465_2476# x1.x6.floating 0.0013f
C993 x4.x9.output_stack sample_code0[1] 0.0744f
C994 VDD x2.x7.floating 0.0321f
C995 a_5970_n713# x3.x6.floating 0.00278f
C996 a_12839_n575# x2.x10.Y 6.65e-20
C997 x3.IN a_6749_n1239# 0.15f
C998 a_6130_n575# x3.x7.floating 0.00409f
C999 VDD x1.x5[7].floating 44f
C1000 x4.x9.output_stack a_567_1950# 0.0388f
C1001 a_12767_n851# x2.x7.floating 8.52e-19
C1002 a_6130_n851# x3.x6.SW 0.00179f
C1003 x2.x9.output_stack x2.x4[3].floating 0.636f
C1004 sample_delay_offset sample_code0[1] 0.0287f
C1005 sample_delay_offset a_12767_n437# 0.00123f
C1006 sample_code2[0] x3.x6.SW 3.98e-21
C1007 sample_delay_offset a_567_1950# 0.0189f
C1008 x2.IN a_12726_n2240# 0.00847f
C1009 x3.IN a_6017_n1964# 0.00921f
C1010 x1.IN x1.x5[7].floating 0.00127f
C1011 x2.x7.floating x2.x10.Y 0.00345f
C1012 x3.x10.Y x3.x6.floating 0.0881f
C1013 sample_code2[0] x3.x3[1].floating 3.8e-20
C1014 x1.x3[1].floating x1.x2.floating 1.17f
C1015 x4.x9.output_stack x1.x6.floating 4.17e-19
C1016 x4.x2.floating sample_code1[0] 1.61e-20
C1017 a_12839_n23# x2.x4[3].floating 7.17e-20
C1018 x4.x3[1].floating sample_code1[2] 3.74e-20
C1019 sample_code1[0] x2.x9.output_stack 4.11e-21
C1020 sample_code0[0] a_6465_2135# 0.00169f
C1021 a_6058_n23# x3.x7.floating 8.52e-19
C1022 x1.x9.output_stack a_13174_2135# 0.00892f
C1023 sample_code0[2] sample_code0[0] 7.44e-20
C1024 sample_delay_offset a_567_1398# 0.00299f
C1025 sample_code1[0] x3.IN 6.06e-20
C1026 x1.x9.output_stack sample_code1[2] 0.333f
C1027 a_12839_n299# a_12839_n575# 0.0316f
C1028 sample_delay_offset x1.x6.floating 0.0706f
C1029 a_7301_3201# x1.x6.floating 0.00996f
C1030 VDD a_6105_n2378# 0.171f
C1031 sample_delay_offset x3.x6.SW 0.19f
C1032 sample_code3[1] x3.x2.floating 0.00656f
C1033 x1.x7.floating x1.x4[3].floating 1.18f
C1034 x1.x9.output_stack a_7436_1536# 1.74e-19
C1035 x3.IN x2.x9.output_stack 0.127f
C1036 sample_delay_offset x3.x3[1].floating 4.68e-20
C1037 x3.x4[3].floating sample_code2[2] 6.52e-20
C1038 x2.x5[7].floating a_12726_n1964# 0.00169f
C1039 a_40_n1036# x3.x3[1].floating 3.09e-19
C1040 a_12839_n299# x2.x7.floating 0.00409f
C1041 VDD x4.x7.floating 0.0282f
C1042 x3.x2.floating x3.x5[7].floating 0.441f
C1043 x4.x6.floating sample_code0[1] 1.27e-19
C1044 a_592_3477# a_592_3201# 0.0316f
C1045 a_5970_n437# x3.x6.SW 1.28e-19
C1046 a_6130_n23# x3.x6.SW 3.1e-20
C1047 x1.x6.SW a_7276_1674# 8.11e-20
C1048 a_592_2925# x4.x10.Y 0.039f
C1049 a_5970_n713# a_6130_n851# 0.0388f
C1050 a_680_3339# x4.x9.output_stack 1.5e-19
C1051 a_12679_n713# a_12767_n575# 0.00227f
C1052 x4.x5[7].floating sample_code1[2] 3.3e-21
C1053 a_6017_n1964# a_6105_n2102# 0.0704f
C1054 a_12814_n1826# a_12814_n2102# 0.0316f
C1055 x4.x6.SW sample_code0[1] 5.52e-21
C1056 x4.x10.Y sample_code0[2] 0.00203f
C1057 sample_delay_offset a_12726_n2240# 1.9e-19
C1058 a_5970_n713# x2.x2.floating 6.24e-19
C1059 a_567_1122# sample_code3[1] 1.48e-20
C1060 x4.x6.SW a_567_1950# 0.00179f
C1061 a_680_3339# sample_delay_offset 1.9e-19
C1062 x1.x7.floating a_7276_1674# 0.00409f
C1063 x3.x5[7].floating a_6017_n2240# 0.00154f
C1064 x2.x7.floating x2.x6.floating 0.202f
C1065 x1.x6.SW a_7276_1122# 3.1e-20
C1066 a_13174_2476# x1.x5[7].floating 0.0132f
C1067 a_12679_n161# a_12839_n299# 0.0388f
C1068 a_6058_n161# a_6130_n299# 0.00227f
C1069 a_12767_n713# x2.x7.floating 8.52e-19
C1070 a_6130_n851# x3.x10.Y 1.69e-19
C1071 x4.x6.SW a_567_1398# 4.74e-20
C1072 sample_code2[0] x3.x10.Y 2.78e-20
C1073 x1.x7.floating a_7276_1122# 0.00218f
C1074 sample_code3[2] sample_code2[2] 5.92e-20
C1075 x2.IN a_12767_n23# 1.8e-19
C1076 x4.x2.floating a_7364_1950# 1.6e-19
C1077 sample_delay_offset a_5970_n713# 0.015f
C1078 x2.IN a_12814_n2378# 0.00832f
C1079 x3.IN a_6105_n2102# 0.00866f
C1080 x3.x9.output_stack x3.x2.floating 0.193f
C1081 x4.x3[1].floating sample_code1[1] 3.46e-20
C1082 sample_code0[1] sample_code0[0] 2.72f
C1083 x1.x10.Y x1.x4[3].floating 0.00668f
C1084 x1.x9.output_stack sample_code1[1] 0.0731f
C1085 x4.x2.floating a_7364_1398# 2.21e-19
C1086 x1.x4[3].floating a_7276_1950# 1.17e-19
C1087 a_12679_n161# x2.x6.floating 0.00109f
C1088 sample_code3[0] x3.x2.floating 0.17f
C1089 x1.x7.floating a_7364_2088# 8.52e-19
C1090 sample_code1[0] a_13174_2135# 0.00169f
C1091 x4.x7.floating a_655_1950# 8.52e-19
C1092 sample_code1[2] sample_code1[0] 5.83e-20
C1093 sample_delay_offset x3.x10.Y 0.0402f
C1094 x4.x9.output_stack a_655_2088# 0.00227f
C1095 a_5970_n437# a_5970_n713# 0.0316f
C1096 a_727_1812# a_567_1674# 0.0388f
C1097 a_12679_n437# a_12767_n437# 0.00227f
C1098 x1.x6.SW a_6465_2476# 0.00208f
C1099 a_6130_n851# x3.x4[3].floating 1.17e-19
C1100 a_680_3339# x4.x6.floating 0.0191f
C1101 a_7301_3477# x4.x5[7].floating 4.6e-19
C1102 x2.IN a_12679_n713# 0.0166f
C1103 x3.x9.output_stack a_6017_n2240# 1.5e-19
C1104 x1.x7.floating a_7364_1536# 8.52e-19
C1105 x3.x3[1].floating sample_code2[1] 3.52e-20
C1106 sample_code2[0] x3.x4[3].floating 0.00915f
C1107 sample_delay_offset a_655_2088# 0.00167f
C1108 x1.x4[3].floating a_7276_1398# 1.17e-19
C1109 x4.x7.floating a_655_1398# 8.52e-19
C1110 x3.IN a_6130_n575# 0.0136f
C1111 x4.x2.floating sample_code1[2] 0.00611f
C1112 a_727_1536# a_567_1398# 0.0388f
C1113 sample_code1[2] x3.IN 4.34e-20
C1114 x2.x5[7].floating a_12814_n2102# 2.76e-19
C1115 x1.x9.output_stack x1.x5[7].floating 1.19f
C1116 a_40_n1036# out 0.149f
C1117 VDD x1.x4[3].floating 0.0565f
C1118 a_6130_n23# x3.x10.Y 2.2e-20
C1119 x1.x10.Y a_7276_1674# 6.65e-20
C1120 sample_delay_offset a_655_1536# 0.00111f
C1121 a_567_1122# sample_code3[0] 1.29e-20
C1122 a_7276_1950# a_7276_1674# 0.0316f
C1123 x4.x2.floating a_7436_1536# 6.88e-19
C1124 x4.x10.Y sample_code0[1] 6.94e-19
C1125 sample_delay_offset a_12767_n23# 9.67e-19
C1126 x4.x9.output_stack x1.x6.SW 3.62e-19
C1127 a_727_1260# a_567_1122# 0.0388f
C1128 sample_code1[1] x3.x9.output_stack 2.48e-21
C1129 x4.x10.Y a_567_1950# 1.69e-19
C1130 sample_delay_offset x3.x4[3].floating 0.00736f
C1131 a_12726_n1964# a_12814_n2102# 0.0704f
C1132 a_6017_n1964# a_6017_n2240# 0.0316f
C1133 x1.IN x1.x4[3].floating 6.65e-19
C1134 x2.IN x2.x6.SW 0.0928f
C1135 sample_delay_offset a_12814_n2378# 3.28e-19
C1136 x3.IN a_6058_n23# 1.8e-19
C1137 VDD a_592_3201# 0.0313f
C1138 x1.x10.Y a_7276_1122# 2.2e-20
C1139 a_7301_3201# x1.x6.SW 9.98e-20
C1140 sample_delay_offset x1.x6.SW 0.19f
C1141 a_7276_1674# a_7276_1398# 0.0316f
C1142 x4.x9.output_stack x1.x7.floating 3.32e-19
C1143 x4.x9.output_stack x4.x4[3].floating 0.636f
C1144 x3.x5[7].floating a_6105_n2378# 2.14e-19
C1145 VDD sample_code2[2] 0.0375f
C1146 x4.x10.Y a_567_1398# 4.07e-20
C1147 a_592_3477# sample_delay_offset 3.28e-19
C1148 sample_code3[2] sample_code2[0] 2.25f
C1149 sample_delay_offset x1.x7.floating 0.259f
C1150 VDD x3.x6.floating 5.87f
C1151 sample_delay_offset x4.x4[3].floating 0.00732f
C1152 a_7301_2925# x1.x5[7].floating 2.76e-19
C1153 a_12839_n575# x2.x4[3].floating 1.17e-19
C1154 a_6058_n575# x3.x7.floating 8.52e-19
C1155 a_5970_n437# x3.x4[3].floating 8.29e-19
C1156 a_6130_n23# x3.x4[3].floating 7.17e-20
C1157 a_7276_1398# a_7276_1122# 0.0316f
C1158 x1.IN sample_code2[2] 5.86e-20
C1159 sample_code1[0] a_567_1122# 6.54e-20
C1160 x1.x10.Y x2.IN 1.13e-19
C1161 a_7276_1950# a_7364_2088# 0.00227f
C1162 sample_code1[2] a_7364_1950# 1.01e-19
C1163 sample_delay_offset a_12679_n713# 0.0153f
C1164 sample_code2[2] x2.x10.Y 0.00201f
C1165 a_7389_3339# a_7301_3201# 0.0704f
C1166 a_7389_3339# sample_delay_offset 1.9e-19
C1167 x1.IN a_7276_1674# 0.0136f
C1168 x3.IN a_6017_n2240# 0.00847f
C1169 sample_code1[1] sample_code1[0] 6.51f
C1170 x3.x6.SW x2.x5[7].floating 0.00313f
C1171 x2.x4[3].floating x2.x7.floating 1.18f
C1172 a_12814_n2378# VSS 0.0953f
C1173 a_6105_n2378# VSS 0.0334f
C1174 a_12726_n2240# VSS 0.032f
C1175 a_6017_n2240# VSS 0.0233f
C1176 a_12814_n2102# VSS 0.0815f
C1177 a_6105_n2102# VSS 0.018f
C1178 a_12726_n1964# VSS 0.0402f
C1179 a_6017_n1964# VSS 0.0348f
C1180 a_12814_n1826# VSS 0.0147f
C1181 a_6105_n1826# VSS 0.00895f
C1182 x2.x6.floating VSS 0.353f
C1183 x2.x5[7].floating VSS 0.107p
C1184 a_6749_n1239# VSS 0.334f
C1185 x2.x6.SW VSS 0.299f
C1186 x2.x10.Y VSS 2.77f
C1187 x3.x6.floating VSS 0.218f
C1188 x3.x5[7].floating VSS 0.107p
C1189 a_40_n1239# VSS 0.319f
C1190 x3.x6.SW VSS 0.282f
C1191 x3.x10.Y VSS 2.75f
C1192 x2.x7.floating VSS 5.89f
C1193 x2.x4[3].floating VSS 21.7f
C1194 x2.x3[1].floating VSS 10.9f
C1195 x2.x2.floating VSS 6.35f
C1196 sample_code2[2] VSS 11.3f
C1197 sample_code2[1] VSS 10.4f
C1198 x3.x7.floating VSS 5.82f
C1199 x3.x4[3].floating VSS 21.7f
C1200 x3.x3[1].floating VSS 10.9f
C1201 x3.x2.floating VSS 6.42f
C1202 sample_code2[0] VSS -12f
C1203 a_12767_n851# VSS 6.32e-19
C1204 sample_code3[2] VSS 3.99f
C1205 sample_code3[1] VSS 1.27f
C1206 out VSS 0.43f
C1207 sample_code3[0] VSS 1.07f
C1208 a_6749_n1036# VSS 0.275f
C1209 x2.x9.output_stack VSS 1.54f
C1210 a_6058_n851# VSS 6.56e-19
C1211 a_40_n1036# VSS 0.295f
C1212 x3.x9.output_stack VSS 1.52f
C1213 a_12839_n851# VSS 0.103f
C1214 a_12767_n713# VSS 6.69e-19
C1215 a_6130_n851# VSS 0.114f
C1216 a_6058_n713# VSS 7.81e-19
C1217 a_12767_n575# VSS 7.52e-19
C1218 a_12679_n713# VSS 0.108f
C1219 a_6058_n575# VSS 7.43e-19
C1220 a_5970_n713# VSS 0.112f
C1221 a_12839_n575# VSS 0.0982f
C1222 a_12767_n437# VSS 0.00106f
C1223 a_6130_n575# VSS 0.11f
C1224 a_6058_n437# VSS 9.98e-19
C1225 a_12767_n299# VSS 0.00116f
C1226 a_12679_n437# VSS 0.111f
C1227 a_6058_n299# VSS 0.00109f
C1228 a_5970_n437# VSS 0.114f
C1229 a_12839_n299# VSS 0.0991f
C1230 a_12767_n161# VSS 0.00129f
C1231 a_6130_n299# VSS 0.111f
C1232 a_6058_n161# VSS 0.00121f
C1233 a_12767_n23# VSS 0.00145f
C1234 a_12679_n161# VSS 0.161f
C1235 a_6058_n23# VSS 0.00134f
C1236 a_5970_n161# VSS 0.165f
C1237 a_12839_n23# VSS 0.164f
C1238 a_12767_115# VSS 0.0049f
C1239 a_6130_n23# VSS 0.17f
C1240 a_6058_115# VSS 0.005f
C1241 x3.IN VSS 1.77f
C1242 a_7364_1122# VSS 0.005f
C1243 a_655_1122# VSS 0.00476f
C1244 a_7364_1260# VSS 0.00134f
C1245 a_7276_1122# VSS 0.17f
C1246 a_655_1260# VSS 0.00134f
C1247 a_567_1122# VSS 0.172f
C1248 a_7436_1260# VSS 0.165f
C1249 a_7364_1398# VSS 0.00121f
C1250 a_727_1260# VSS 0.165f
C1251 a_655_1398# VSS 0.00121f
C1252 a_7364_1536# VSS 0.00109f
C1253 a_7276_1398# VSS 0.111f
C1254 a_655_1536# VSS 0.00114f
C1255 a_567_1398# VSS 0.117f
C1256 a_7436_1536# VSS 0.114f
C1257 a_7364_1674# VSS 9.98e-19
C1258 a_727_1536# VSS 0.115f
C1259 a_655_1674# VSS 0.00157f
C1260 a_7364_1812# VSS 7.43e-19
C1261 a_7276_1674# VSS 0.11f
C1262 a_655_1812# VSS 7.43e-19
C1263 a_567_1674# VSS 0.115f
C1264 a_7436_1812# VSS 0.112f
C1265 a_7364_1950# VSS 7.81e-19
C1266 a_727_1812# VSS 0.112f
C1267 a_655_1950# VSS 6.69e-19
C1268 a_7364_2088# VSS 6.56e-19
C1269 a_7276_1950# VSS 0.114f
C1270 a_655_2088# VSS 6.32e-19
C1271 a_567_1950# VSS 0.12f
C1272 a_13174_2135# VSS 0.256f
C1273 x1.x2.floating VSS 6.41f
C1274 x1.x3[1].floating VSS 10.9f
C1275 x1.x4[3].floating VSS 21.7f
C1276 x1.x7.floating VSS 5.82f
C1277 sample_code1[0] VSS -50.7f
C1278 sample_code1[1] VSS 12f
C1279 sample_code1[2] VSS 8.97f
C1280 a_6465_2135# VSS 0.276f
C1281 x4.x2.floating VSS 6.35f
C1282 x4.x3[1].floating VSS 10.9f
C1283 x4.x4[3].floating VSS 21.7f
C1284 x4.x7.floating VSS 5.89f
C1285 sample_code0[0] VSS -4.98f
C1286 sample_code0[1] VSS 3.9f
C1287 sample_code0[2] VSS 2.4f
C1288 x1.x5[7].floating VSS 0.107p
C1289 x1.x6.floating VSS 0.218f
C1290 x2.IN VSS 3.34f
C1291 x4.x5[7].floating VSS 0.107p
C1292 x4.x6.floating VSS 0.403f
C1293 a_13174_2476# VSS 0.319f
C1294 a_6465_2476# VSS 0.334f
C1295 x1.x9.output_stack VSS 1.53f
C1296 x1.x6.SW VSS 0.282f
C1297 x1.x10.Y VSS 2.75f
C1298 x4.x9.output_stack VSS 1.51f
C1299 x4.x6.SW VSS 0.299f
C1300 x4.x10.Y VSS 2.76f
C1301 a_7301_2925# VSS 0.00895f
C1302 sample_delay_offset VSS 10.6f
C1303 a_592_2925# VSS 0.0147f
C1304 a_7389_3063# VSS 0.0348f
C1305 a_680_3063# VSS 0.0402f
C1306 a_7301_3201# VSS 0.0226f
C1307 a_592_3201# VSS 0.0815f
C1308 a_7389_3339# VSS 0.0236f
C1309 a_680_3339# VSS 0.032f
C1310 a_7301_3477# VSS 0.0292f
C1311 x1.IN VSS 1.77f
C1312 a_592_3477# VSS 0.0953f
C1313 VDD VSS 80.8f
C1314 sample_code0[0].t0 VSS 0.0571f
C1315 sample_code0[0].n0 VSS 12.1f
C1316 sample_code1[0].t0 VSS 0.0731f
C1317 sample_code1[0].n0 VSS 66f
C1318 sample_code2[0].t0 VSS 0.0529f
C1319 sample_code2[0].n0 VSS 0.923f
C1320 sample_code2[0].n1 VSS 19.7f
C1321 sample_code2[2].t0 VSS 0.0532f
C1322 sample_code2[2].t2 VSS 0.0532f
C1323 sample_code2[2].n0 VSS 0.211f
C1324 sample_code2[2].n1 VSS 0.702f
C1325 sample_code2[2].t1 VSS 0.0533f
C1326 sample_code2[2].t3 VSS 0.0532f
C1327 sample_code2[2].n2 VSS 1.3f
C1328 sample_code1[2].t0 VSS 0.0455f
C1329 sample_code1[2].n0 VSS 0.177f
C1330 sample_code1[2].t1 VSS 0.0456f
C1331 sample_code1[2].t3 VSS 0.0455f
C1332 sample_code1[2].n1 VSS 0.181f
C1333 sample_code1[2].t2 VSS 0.0455f
C1334 sample_code1[2].n2 VSS 1.69f
C1335 x3.x5[7].floating.n0 VSS 2.8f
C1336 x3.x5[7].floating.n1 VSS 51.3f
C1337 x3.x5[7].floating.n2 VSS 2.78f
C1338 x3.x5[7].floating.n3 VSS 1.06f
C1339 x3.x5[7].floating.n4 VSS 0.366f
C1340 x3.x5[7].floating.n5 VSS 1.16f
C1341 x3.x5[7].floating.t5 VSS 0.857f
C1342 x3.x5[7].floating.n6 VSS 6.48f
C1343 x3.x5[7].floating.n7 VSS 1.35f
C1344 x3.x5[7].floating.n8 VSS 2.18f
C1345 x3.x5[7].floating.n9 VSS 1.06f
C1346 x3.x5[7].floating.n10 VSS -15.2f
C1347 x3.x5[7].floating.n11 VSS -15.1f
C1348 x3.x5[7].floating.n12 VSS -41.5f
C1349 x3.x5[7].floating.n13 VSS 0.765f
C1350 x3.x5[7].floating.n14 VSS 2.46f
C1351 x3.x5[7].floating.n15 VSS 51.4f
C1352 x3.x5[7].floating.n16 VSS 2.46f
C1353 x3.x5[7].floating.n17 VSS 0.765f
C1354 x3.x5[7].floating.n18 VSS -33.4f
C1355 x3.x5[7].floating.n19 VSS -4.55f
C1356 x3.x5[7].floating.n20 VSS 3.82f
C1357 x3.x5[7].floating.n21 VSS -28.8f
C1358 x3.x5[7].floating.n22 VSS -7.06f
C1359 x3.x5[7].floating.n23 VSS 2.68f
C1360 x3.x5[7].floating.n24 VSS 1.06f
C1361 x3.x5[7].floating.n25 VSS 0.363f
C1362 x3.x5[7].floating.n26 VSS 1.21f
C1363 x3.x5[7].floating.t2 VSS 0.857f
C1364 x3.x5[7].floating.n27 VSS 6.65f
C1365 x3.x5[7].floating.n28 VSS 1.15f
C1366 x3.x5[7].floating.n29 VSS 2.16f
C1367 x3.x5[7].floating.n30 VSS 1.06f
C1368 x3.x5[7].floating.n31 VSS 2.22f
C1369 x3.x5[7].floating.n32 VSS -8f
C1370 x3.x5[7].floating.n33 VSS -28.8f
C1371 x3.x5[7].floating.n34 VSS 3.82f
C1372 x3.x5[7].floating.n35 VSS -7.06f
C1373 x3.x5[7].floating.n36 VSS -28.3f
C1374 x3.x5[7].floating.n37 VSS 52.6f
C1375 x3.x5[7].floating.n38 VSS -28.3f
C1376 x3.x5[7].floating.n39 VSS -7.06f
C1377 x3.x5[7].floating.n40 VSS 3.82f
C1378 x3.x5[7].floating.n41 VSS -28.8f
C1379 x3.x5[7].floating.n42 VSS -7.97f
C1380 x3.x5[7].floating.n43 VSS 2.21f
C1381 x3.x5[7].floating.n44 VSS 1.16f
C1382 x3.x5[7].floating.t6 VSS 0.857f
C1383 x3.x5[7].floating.n45 VSS 6.48f
C1384 x3.x5[7].floating.n46 VSS 1.35f
C1385 x3.x5[7].floating.n47 VSS 2.18f
C1386 x3.x5[7].floating.n48 VSS 1.06f
C1387 x3.x5[7].floating.n49 VSS 0.366f
C1388 x3.x5[7].floating.n50 VSS 1.06f
C1389 x3.x5[7].floating.n51 VSS 2.78f
C1390 x3.x5[7].floating.n52 VSS 51.3f
C1391 x3.x5[7].floating.n53 VSS 2.8f
C1392 x3.x5[7].floating.n54 VSS 1.06f
C1393 x3.x5[7].floating.n55 VSS 0.363f
C1394 x3.x5[7].floating.n56 VSS 1.21f
C1395 x3.x5[7].floating.t1 VSS 0.857f
C1396 x3.x5[7].floating.n57 VSS 6.65f
C1397 x3.x5[7].floating.n58 VSS 1.15f
C1398 x3.x5[7].floating.n59 VSS 2.16f
C1399 x3.x5[7].floating.n60 VSS 1.06f
C1400 x3.x5[7].floating.n61 VSS 2.22f
C1401 x3.x5[7].floating.n62 VSS -8f
C1402 x3.x5[7].floating.n63 VSS -28.8f
C1403 x3.x5[7].floating.n64 VSS 3.82f
C1404 x3.x5[7].floating.n65 VSS -7.06f
C1405 x3.x5[7].floating.n66 VSS -28.3f
C1406 x3.x5[7].floating.n67 VSS 52.6f
C1407 x3.x5[7].floating.n68 VSS -28.3f
C1408 x3.x5[7].floating.n69 VSS -7.06f
C1409 x3.x5[7].floating.n70 VSS 3.82f
C1410 x3.x5[7].floating.n71 VSS -28.8f
C1411 x3.x5[7].floating.n72 VSS -7.97f
C1412 x3.x5[7].floating.n73 VSS 2.21f
C1413 x3.x5[7].floating.n74 VSS 1.16f
C1414 x3.x5[7].floating.t4 VSS 0.857f
C1415 x3.x5[7].floating.n75 VSS 6.48f
C1416 x3.x5[7].floating.n76 VSS 1.35f
C1417 x3.x5[7].floating.n77 VSS 2.18f
C1418 x3.x5[7].floating.n78 VSS 1.06f
C1419 x3.x5[7].floating.n79 VSS 0.366f
C1420 x3.x5[7].floating.n80 VSS 1.06f
C1421 x3.x5[7].floating.n81 VSS 2.78f
C1422 x3.x5[7].floating.n82 VSS 51.3f
C1423 x3.x5[7].floating.n83 VSS 2.8f
C1424 x3.x5[7].floating.n84 VSS 1.06f
C1425 x3.x5[7].floating.n85 VSS 0.363f
C1426 x3.x5[7].floating.n86 VSS 1.21f
C1427 x3.x5[7].floating.t0 VSS 0.857f
C1428 x3.x5[7].floating.n87 VSS 6.65f
C1429 x3.x5[7].floating.n88 VSS 1.15f
C1430 x3.x5[7].floating.n89 VSS 2.16f
C1431 x3.x5[7].floating.n90 VSS 1.06f
C1432 x3.x5[7].floating.n91 VSS 2.22f
C1433 x3.x5[7].floating.n92 VSS -8f
C1434 x3.x5[7].floating.n93 VSS -28.8f
C1435 x3.x5[7].floating.n94 VSS 3.82f
C1436 x3.x5[7].floating.n95 VSS -7.06f
C1437 x3.x5[7].floating.n96 VSS -28.3f
C1438 x3.x5[7].floating.n97 VSS 52.6f
C1439 x3.x5[7].floating.n98 VSS -28.3f
C1440 x3.x5[7].floating.n99 VSS -7.06f
C1441 x3.x5[7].floating.n100 VSS 3.82f
C1442 x3.x5[7].floating.n101 VSS -28.8f
C1443 x3.x5[7].floating.n102 VSS -7.97f
C1444 x3.x5[7].floating.n103 VSS 2.21f
C1445 x3.x5[7].floating.n104 VSS 1.16f
C1446 x3.x5[7].floating.t3 VSS 0.857f
C1447 x3.x5[7].floating.n105 VSS 6.48f
C1448 x3.x5[7].floating.n106 VSS 1.35f
C1449 x3.x5[7].floating.n107 VSS 2.18f
C1450 x3.x5[7].floating.n108 VSS 1.06f
C1451 x3.x5[7].floating.n109 VSS 0.366f
C1452 x3.x5[7].floating.n110 VSS 1.06f
C1453 x3.x5[7].floating.n111 VSS 2.78f
C1454 x3.x5[7].floating.n112 VSS 51.3f
C1455 x3.x5[7].floating.n113 VSS 2.8f
C1456 x3.x5[7].floating.n114 VSS 1.06f
C1457 x3.x5[7].floating.n115 VSS 0.363f
C1458 x3.x5[7].floating.n116 VSS 1.21f
C1459 x3.x5[7].floating.t7 VSS 0.857f
C1460 x3.x5[7].floating.n117 VSS 6.65f
C1461 x3.x5[7].floating.n118 VSS 1.15f
C1462 x3.x5[7].floating.n119 VSS 2.16f
C1463 x3.x5[7].floating.n120 VSS 1.06f
C1464 x3.x5[7].floating.n121 VSS -17.3f
C1465 x3.x5[7].floating.n122 VSS -17.2f
C1466 x3.x5[7].floating.n123 VSS -43.5f
C1467 x3.x5[7].floating.n124 VSS 0.765f
C1468 x3.x5[7].floating.n125 VSS 2.46f
C1469 x3.x5[7].floating.n126 VSS 51.4f
C1470 x3.x5[7].floating.n127 VSS 2.46f
C1471 x3.x5[7].floating.n128 VSS 0.765f
C1472 x3.x5[7].floating.n129 VSS -32.9f
C1473 x3.x5[7].floating.n130 VSS -5f
C1474 x3.x5[7].floating.n131 VSS 3.82f
C1475 x3.x5[7].floating.n132 VSS -28.8f
C1476 x3.x5[7].floating.n133 VSS -7.82f
C1477 x3.x5[7].floating.n134 VSS 3.23f
C1478 x3.x5[7].floating.n135 VSS 51.9f
C1479 x3.x5[7].floating.n136 VSS 2.68f
C1480 x3.x5[7].floating.n137 VSS -7.06f
C1481 x3.x5[7].floating.n138 VSS -28.8f
C1482 x3.x5[7].floating.n139 VSS 3.82f
C1483 x3.x5[7].floating.n140 VSS -4.55f
C1484 x3.x5[7].floating.n141 VSS -33.4f
C1485 x3.x5[7].floating.n142 VSS 0.765f
C1486 x3.x5[7].floating.n143 VSS 2.46f
C1487 x3.x5[7].floating.n144 VSS 51.4f
C1488 x3.x5[7].floating.n145 VSS 2.46f
C1489 x3.x5[7].floating.n146 VSS 0.765f
C1490 x3.x5[7].floating.n147 VSS -32.9f
C1491 x3.x5[7].floating.n148 VSS -5f
C1492 x3.x5[7].floating.n149 VSS 3.82f
C1493 x3.x5[7].floating.n150 VSS -28.8f
C1494 x3.x5[7].floating.n151 VSS -7.82f
C1495 x3.x5[7].floating.n152 VSS 3.23f
C1496 x3.x5[7].floating.n153 VSS 51.9f
C1497 x3.x5[7].floating.n154 VSS 2.68f
C1498 x3.x5[7].floating.n155 VSS -7.06f
C1499 x3.x5[7].floating.n156 VSS -28.8f
C1500 x3.x5[7].floating.n157 VSS 3.82f
C1501 x3.x5[7].floating.n158 VSS -4.55f
C1502 x3.x5[7].floating.n159 VSS -33.4f
C1503 x3.x5[7].floating.n160 VSS 0.765f
C1504 x3.x5[7].floating.n161 VSS 2.46f
C1505 x3.x5[7].floating.n162 VSS 51.4f
C1506 x3.x5[7].floating.n163 VSS 2.46f
C1507 x3.x5[7].floating.n164 VSS 0.765f
C1508 x3.x5[7].floating.n165 VSS -32.9f
C1509 x3.x5[7].floating.n166 VSS -5f
C1510 x3.x5[7].floating.n167 VSS 3.82f
C1511 x3.x5[7].floating.n168 VSS -28.8f
C1512 x3.x5[7].floating.n169 VSS -7.82f
C1513 x3.x5[7].floating.n170 VSS 3.23f
C1514 x3.x5[7].floating.n171 VSS 51.9f
C1515 x3.x10.Y.n0 VSS 0.0359f
C1516 x3.x10.Y.t1 VSS 0.0526f
C1517 x3.x10.Y.n1 VSS 0.0169f
C1518 x3.x10.Y.n2 VSS 0.00704f
C1519 x3.x10.Y.t0 VSS 0.0181f
C1520 x3.x10.Y.n3 VSS 0.0188f
C1521 x3.x10.Y.n4 VSS 0.019f
C1522 x3.x10.Y.n5 VSS 0.221f
C1523 x3.x10.Y.t4 VSS 0.0167f
C1524 x3.x10.Y.t7 VSS 0.0167f
C1525 x3.x10.Y.t3 VSS 0.0167f
C1526 x3.x10.Y.t8 VSS 0.0167f
C1527 x3.x10.Y.t5 VSS 0.0167f
C1528 x3.x10.Y.t9 VSS 0.0167f
C1529 x3.x10.Y.t6 VSS 0.0167f
C1530 x3.x10.Y.t2 VSS 0.0167f
C1531 sample_code0[1].t0 VSS 0.0282f
C1532 sample_code0[1].t1 VSS 0.0282f
C1533 sample_code0[1].n0 VSS 0.694f
C1534 x1.x5[7].floating.n0 VSS 2.79f
C1535 x1.x5[7].floating.n1 VSS 1.06f
C1536 x1.x5[7].floating.n2 VSS 0.364f
C1537 x1.x5[7].floating.t5 VSS 0.859f
C1538 x1.x5[7].floating.n3 VSS 6.48f
C1539 x1.x5[7].floating.n4 VSS 1.15f
C1540 x1.x5[7].floating.n5 VSS 1.36f
C1541 x1.x5[7].floating.n6 VSS 2.2f
C1542 x1.x5[7].floating.n7 VSS 1.06f
C1543 x1.x5[7].floating.n8 VSS 2.23f
C1544 x1.x5[7].floating.n9 VSS -7.99f
C1545 x1.x5[7].floating.n10 VSS -28.9f
C1546 x1.x5[7].floating.n11 VSS 3.83f
C1547 x1.x5[7].floating.n12 VSS -7.07f
C1548 x1.x5[7].floating.n13 VSS -28.3f
C1549 x1.x5[7].floating.n14 VSS 52.7f
C1550 x1.x5[7].floating.n15 VSS -28.3f
C1551 x1.x5[7].floating.n16 VSS -7.07f
C1552 x1.x5[7].floating.n17 VSS 3.83f
C1553 x1.x5[7].floating.n18 VSS -28.9f
C1554 x1.x5[7].floating.n19 VSS -8.01f
C1555 x1.x5[7].floating.n20 VSS 2.21f
C1556 x1.x5[7].floating.t0 VSS 0.859f
C1557 x1.x5[7].floating.n21 VSS 6.65f
C1558 x1.x5[7].floating.n22 VSS 1.21f
C1559 x1.x5[7].floating.n23 VSS 1.17f
C1560 x1.x5[7].floating.n24 VSS 2.18f
C1561 x1.x5[7].floating.n25 VSS 1.06f
C1562 x1.x5[7].floating.n26 VSS 0.366f
C1563 x1.x5[7].floating.n27 VSS 1.06f
C1564 x1.x5[7].floating.n28 VSS 2.8f
C1565 x1.x5[7].floating.n29 VSS 51.4f
C1566 x1.x5[7].floating.n30 VSS 2.79f
C1567 x1.x5[7].floating.n31 VSS 1.06f
C1568 x1.x5[7].floating.n32 VSS 0.364f
C1569 x1.x5[7].floating.t1 VSS 0.859f
C1570 x1.x5[7].floating.n33 VSS 6.48f
C1571 x1.x5[7].floating.n34 VSS 1.15f
C1572 x1.x5[7].floating.n35 VSS 1.36f
C1573 x1.x5[7].floating.n36 VSS 2.2f
C1574 x1.x5[7].floating.n37 VSS 1.06f
C1575 x1.x5[7].floating.n38 VSS 2.23f
C1576 x1.x5[7].floating.n39 VSS -7.99f
C1577 x1.x5[7].floating.n40 VSS -28.9f
C1578 x1.x5[7].floating.n41 VSS 3.83f
C1579 x1.x5[7].floating.n42 VSS -7.07f
C1580 x1.x5[7].floating.n43 VSS -28.3f
C1581 x1.x5[7].floating.n44 VSS 52.7f
C1582 x1.x5[7].floating.n45 VSS -28.3f
C1583 x1.x5[7].floating.n46 VSS -7.07f
C1584 x1.x5[7].floating.n47 VSS 3.83f
C1585 x1.x5[7].floating.n48 VSS -28.9f
C1586 x1.x5[7].floating.n49 VSS -8.01f
C1587 x1.x5[7].floating.n50 VSS 2.21f
C1588 x1.x5[7].floating.t3 VSS 0.859f
C1589 x1.x5[7].floating.n51 VSS 6.65f
C1590 x1.x5[7].floating.n52 VSS 1.21f
C1591 x1.x5[7].floating.n53 VSS 1.17f
C1592 x1.x5[7].floating.n54 VSS 2.18f
C1593 x1.x5[7].floating.n55 VSS 1.06f
C1594 x1.x5[7].floating.n56 VSS 0.366f
C1595 x1.x5[7].floating.n57 VSS 1.06f
C1596 x1.x5[7].floating.n58 VSS 2.8f
C1597 x1.x5[7].floating.n59 VSS 51.4f
C1598 x1.x5[7].floating.n60 VSS 2.79f
C1599 x1.x5[7].floating.n61 VSS 1.06f
C1600 x1.x5[7].floating.n62 VSS 0.364f
C1601 x1.x5[7].floating.t4 VSS 0.859f
C1602 x1.x5[7].floating.n63 VSS 6.48f
C1603 x1.x5[7].floating.n64 VSS 1.15f
C1604 x1.x5[7].floating.n65 VSS 1.36f
C1605 x1.x5[7].floating.n66 VSS 2.2f
C1606 x1.x5[7].floating.n67 VSS 1.06f
C1607 x1.x5[7].floating.n68 VSS -15.2f
C1608 x1.x5[7].floating.n69 VSS -15.2f
C1609 x1.x5[7].floating.n70 VSS -41.6f
C1610 x1.x5[7].floating.n71 VSS 0.766f
C1611 x1.x5[7].floating.n72 VSS 2.47f
C1612 x1.x5[7].floating.n73 VSS 51.5f
C1613 x1.x5[7].floating.n74 VSS 2.47f
C1614 x1.x5[7].floating.n75 VSS 0.766f
C1615 x1.x5[7].floating.n76 VSS -33.5f
C1616 x1.x5[7].floating.n77 VSS -4.56f
C1617 x1.x5[7].floating.n78 VSS 3.83f
C1618 x1.x5[7].floating.n79 VSS -28.9f
C1619 x1.x5[7].floating.n80 VSS -7.07f
C1620 x1.x5[7].floating.n81 VSS 2.68f
C1621 x1.x5[7].floating.n82 VSS 52f
C1622 x1.x5[7].floating.n83 VSS 3.23f
C1623 x1.x5[7].floating.n84 VSS -7.84f
C1624 x1.x5[7].floating.n85 VSS -28.9f
C1625 x1.x5[7].floating.n86 VSS 3.83f
C1626 x1.x5[7].floating.n87 VSS -5.01f
C1627 x1.x5[7].floating.n88 VSS -33f
C1628 x1.x5[7].floating.n89 VSS 0.766f
C1629 x1.x5[7].floating.n90 VSS 2.47f
C1630 x1.x5[7].floating.n91 VSS 51.5f
C1631 x1.x5[7].floating.n92 VSS 2.47f
C1632 x1.x5[7].floating.n93 VSS 0.766f
C1633 x1.x5[7].floating.n94 VSS -33.5f
C1634 x1.x5[7].floating.n95 VSS -4.56f
C1635 x1.x5[7].floating.n96 VSS 3.83f
C1636 x1.x5[7].floating.n97 VSS -28.9f
C1637 x1.x5[7].floating.n98 VSS -7.07f
C1638 x1.x5[7].floating.n99 VSS 2.68f
C1639 x1.x5[7].floating.n100 VSS 52f
C1640 x1.x5[7].floating.n101 VSS 3.23f
C1641 x1.x5[7].floating.n102 VSS -7.84f
C1642 x1.x5[7].floating.n103 VSS -28.9f
C1643 x1.x5[7].floating.n104 VSS 3.83f
C1644 x1.x5[7].floating.n105 VSS -5.01f
C1645 x1.x5[7].floating.n106 VSS -33f
C1646 x1.x5[7].floating.n107 VSS 0.766f
C1647 x1.x5[7].floating.n108 VSS 2.47f
C1648 x1.x5[7].floating.n109 VSS 2.68f
C1649 x1.x5[7].floating.n110 VSS -7.07f
C1650 x1.x5[7].floating.n111 VSS -28.9f
C1651 x1.x5[7].floating.n112 VSS 3.83f
C1652 x1.x5[7].floating.n113 VSS -4.56f
C1653 x1.x5[7].floating.n114 VSS -33.5f
C1654 x1.x5[7].floating.n115 VSS 0.766f
C1655 x1.x5[7].floating.n116 VSS 2.47f
C1656 x1.x5[7].floating.n117 VSS 51.5f
C1657 x1.x5[7].floating.n118 VSS 51.4f
C1658 x1.x5[7].floating.n119 VSS 2.8f
C1659 x1.x5[7].floating.n120 VSS 1.06f
C1660 x1.x5[7].floating.n121 VSS 0.366f
C1661 x1.x5[7].floating.t7 VSS 0.859f
C1662 x1.x5[7].floating.n122 VSS 6.65f
C1663 x1.x5[7].floating.n123 VSS 1.21f
C1664 x1.x5[7].floating.n124 VSS 1.17f
C1665 x1.x5[7].floating.n125 VSS 2.18f
C1666 x1.x5[7].floating.n126 VSS 1.06f
C1667 x1.x5[7].floating.n127 VSS 2.21f
C1668 x1.x5[7].floating.n128 VSS -8.01f
C1669 x1.x5[7].floating.n129 VSS -28.9f
C1670 x1.x5[7].floating.n130 VSS 3.83f
C1671 x1.x5[7].floating.n131 VSS -7.07f
C1672 x1.x5[7].floating.n132 VSS -28.3f
C1673 x1.x5[7].floating.n133 VSS -7.99f
C1674 x1.x5[7].floating.n134 VSS -28.9f
C1675 x1.x5[7].floating.n135 VSS 3.83f
C1676 x1.x5[7].floating.n136 VSS -7.07f
C1677 x1.x5[7].floating.n137 VSS -28.3f
C1678 x1.x5[7].floating.n138 VSS 52.7f
C1679 x1.x5[7].floating.n139 VSS 52f
C1680 x1.x5[7].floating.n140 VSS 3.23f
C1681 x1.x5[7].floating.n141 VSS 2.23f
C1682 x1.x5[7].floating.t6 VSS 0.859f
C1683 x1.x5[7].floating.n142 VSS 6.48f
C1684 x1.x5[7].floating.n143 VSS 1.15f
C1685 x1.x5[7].floating.n144 VSS 1.36f
C1686 x1.x5[7].floating.n145 VSS 2.2f
C1687 x1.x5[7].floating.n146 VSS 1.06f
C1688 x1.x5[7].floating.n147 VSS 0.364f
C1689 x1.x5[7].floating.n148 VSS 1.06f
C1690 x1.x5[7].floating.n149 VSS 2.79f
C1691 x1.x5[7].floating.n150 VSS 51.4f
C1692 x1.x5[7].floating.n151 VSS 2.8f
C1693 x1.x5[7].floating.n152 VSS 1.06f
C1694 x1.x5[7].floating.n153 VSS 0.366f
C1695 x1.x5[7].floating.t2 VSS 0.859f
C1696 x1.x5[7].floating.n154 VSS 7.16f
C1697 x1.x5[7].floating.n155 VSS 1.21f
C1698 x1.x5[7].floating.n156 VSS 1.17f
C1699 x1.x5[7].floating.n157 VSS 1.67f
C1700 x1.x5[7].floating.n158 VSS 1.06f
C1701 x1.x5[7].floating.n159 VSS -17.4f
C1702 x1.x5[7].floating.n160 VSS -17.2f
C1703 x1.x5[7].floating.n161 VSS -43.6f
C1704 x1.x5[7].floating.n162 VSS 0.766f
C1705 x1.x5[7].floating.n163 VSS 2.47f
C1706 x1.x5[7].floating.n164 VSS 51.5f
C1707 x1.x5[7].floating.n165 VSS 2.47f
C1708 x1.x5[7].floating.n166 VSS 0.766f
C1709 x1.x5[7].floating.n167 VSS -33f
C1710 x1.x5[7].floating.n168 VSS -5.01f
C1711 x1.x5[7].floating.n169 VSS 3.83f
C1712 x1.x5[7].floating.n170 VSS -28.9f
C1713 x1.x5[7].floating.n171 VSS -7.84f
C1714 x1.x10.Y.t0 VSS 0.0462f
C1715 x1.x10.Y.t5 VSS 0.0167f
C1716 x1.x10.Y.t6 VSS 0.0167f
C1717 x1.x10.Y.t8 VSS 0.0167f
C1718 x1.x10.Y.t9 VSS 0.0167f
C1719 x1.x10.Y.t4 VSS 0.0167f
C1720 x1.x10.Y.t2 VSS 0.0167f
C1721 x1.x10.Y.t3 VSS 0.0167f
C1722 x1.x10.Y.t7 VSS 0.0167f
C1723 x1.x10.Y.n0 VSS 0.222f
C1724 x1.x10.Y.n1 VSS 0.0366f
C1725 x1.x10.Y.t1 VSS 0.0174f
C1726 x1.x10.Y.n2 VSS 0.0188f
C1727 x1.x10.Y.n3 VSS 0.0186f
C1728 x1.x10.Y.n4 VSS 0.0151f
C1729 x1.x10.Y.n5 VSS 0.0211f
C1730 sample_code3[2].t1 VSS 0.0192f
C1731 sample_code3[2].t3 VSS 0.0192f
C1732 sample_code3[2].n0 VSS 0.0764f
C1733 sample_code3[2].n1 VSS 0.254f
C1734 sample_code3[2].t0 VSS 0.0192f
C1735 sample_code3[2].t2 VSS 0.0192f
C1736 sample_code3[2].n2 VSS 0.425f
C1737 sample_code2[1].t1 VSS 0.0635f
C1738 sample_code2[1].n0 VSS 0.244f
C1739 sample_code2[1].t0 VSS 0.0635f
C1740 x4.x5[7].floating.n0 VSS -7.99f
C1741 x4.x5[7].floating.n1 VSS -28.9f
C1742 x4.x5[7].floating.n2 VSS 3.83f
C1743 x4.x5[7].floating.n3 VSS -7.07f
C1744 x4.x5[7].floating.n4 VSS -28.3f
C1745 x4.x5[7].floating.n5 VSS 52.7f
C1746 x4.x5[7].floating.n6 VSS -28.3f
C1747 x4.x5[7].floating.n7 VSS -7.07f
C1748 x4.x5[7].floating.n8 VSS 3.83f
C1749 x4.x5[7].floating.n9 VSS -28.9f
C1750 x4.x5[7].floating.n10 VSS -8.01f
C1751 x4.x5[7].floating.n11 VSS 2.21f
C1752 x4.x5[7].floating.t5 VSS 0.859f
C1753 x4.x5[7].floating.n12 VSS 6.65f
C1754 x4.x5[7].floating.n13 VSS 1.21f
C1755 x4.x5[7].floating.n14 VSS 1.17f
C1756 x4.x5[7].floating.n15 VSS 2.18f
C1757 x4.x5[7].floating.n16 VSS 1.06f
C1758 x4.x5[7].floating.n17 VSS 0.366f
C1759 x4.x5[7].floating.n18 VSS 1.06f
C1760 x4.x5[7].floating.n19 VSS 2.8f
C1761 x4.x5[7].floating.n20 VSS 51.4f
C1762 x4.x5[7].floating.n21 VSS 2.79f
C1763 x4.x5[7].floating.n22 VSS 1.06f
C1764 x4.x5[7].floating.n23 VSS 0.364f
C1765 x4.x5[7].floating.t0 VSS 0.859f
C1766 x4.x5[7].floating.n24 VSS 6.48f
C1767 x4.x5[7].floating.n25 VSS 1.15f
C1768 x4.x5[7].floating.n26 VSS 1.36f
C1769 x4.x5[7].floating.n27 VSS 2.2f
C1770 x4.x5[7].floating.n28 VSS 1.06f
C1771 x4.x5[7].floating.n29 VSS 2.23f
C1772 x4.x5[7].floating.n30 VSS -7.99f
C1773 x4.x5[7].floating.n31 VSS -28.9f
C1774 x4.x5[7].floating.n32 VSS 3.83f
C1775 x4.x5[7].floating.n33 VSS -7.07f
C1776 x4.x5[7].floating.n34 VSS -28.3f
C1777 x4.x5[7].floating.n35 VSS 52.7f
C1778 x4.x5[7].floating.n36 VSS -28.3f
C1779 x4.x5[7].floating.n37 VSS -7.07f
C1780 x4.x5[7].floating.n38 VSS 3.83f
C1781 x4.x5[7].floating.n39 VSS -28.9f
C1782 x4.x5[7].floating.n40 VSS -8.01f
C1783 x4.x5[7].floating.n41 VSS 2.21f
C1784 x4.x5[7].floating.t1 VSS 0.859f
C1785 x4.x5[7].floating.n42 VSS 6.65f
C1786 x4.x5[7].floating.n43 VSS 1.21f
C1787 x4.x5[7].floating.n44 VSS 1.17f
C1788 x4.x5[7].floating.n45 VSS 2.18f
C1789 x4.x5[7].floating.n46 VSS 1.06f
C1790 x4.x5[7].floating.n47 VSS 0.366f
C1791 x4.x5[7].floating.n48 VSS 1.06f
C1792 x4.x5[7].floating.n49 VSS 2.8f
C1793 x4.x5[7].floating.n50 VSS 51.4f
C1794 x4.x5[7].floating.n51 VSS 2.79f
C1795 x4.x5[7].floating.n52 VSS 1.06f
C1796 x4.x5[7].floating.n53 VSS 0.364f
C1797 x4.x5[7].floating.t4 VSS 0.859f
C1798 x4.x5[7].floating.n54 VSS 6.48f
C1799 x4.x5[7].floating.n55 VSS 1.15f
C1800 x4.x5[7].floating.n56 VSS 1.36f
C1801 x4.x5[7].floating.n57 VSS 2.2f
C1802 x4.x5[7].floating.n58 VSS 1.06f
C1803 x4.x5[7].floating.n59 VSS -15.2f
C1804 x4.x5[7].floating.n60 VSS -15.2f
C1805 x4.x5[7].floating.n61 VSS -41.6f
C1806 x4.x5[7].floating.n62 VSS 0.766f
C1807 x4.x5[7].floating.n63 VSS 2.47f
C1808 x4.x5[7].floating.n64 VSS 51.5f
C1809 x4.x5[7].floating.n65 VSS 2.47f
C1810 x4.x5[7].floating.n66 VSS 0.766f
C1811 x4.x5[7].floating.n67 VSS -33.5f
C1812 x4.x5[7].floating.n68 VSS -4.56f
C1813 x4.x5[7].floating.n69 VSS 3.83f
C1814 x4.x5[7].floating.n70 VSS -28.9f
C1815 x4.x5[7].floating.n71 VSS -7.07f
C1816 x4.x5[7].floating.n72 VSS 2.68f
C1817 x4.x5[7].floating.n73 VSS 52f
C1818 x4.x5[7].floating.n74 VSS 3.23f
C1819 x4.x5[7].floating.n75 VSS -7.84f
C1820 x4.x5[7].floating.n76 VSS -28.9f
C1821 x4.x5[7].floating.n77 VSS 3.83f
C1822 x4.x5[7].floating.n78 VSS -5.01f
C1823 x4.x5[7].floating.n79 VSS -33f
C1824 x4.x5[7].floating.n80 VSS 0.766f
C1825 x4.x5[7].floating.n81 VSS 2.47f
C1826 x4.x5[7].floating.n82 VSS 2.68f
C1827 x4.x5[7].floating.n83 VSS -7.07f
C1828 x4.x5[7].floating.n84 VSS -28.9f
C1829 x4.x5[7].floating.n85 VSS 3.83f
C1830 x4.x5[7].floating.n86 VSS -4.56f
C1831 x4.x5[7].floating.n87 VSS -33.5f
C1832 x4.x5[7].floating.n88 VSS 0.766f
C1833 x4.x5[7].floating.n89 VSS 2.47f
C1834 x4.x5[7].floating.n90 VSS 51.5f
C1835 x4.x5[7].floating.n91 VSS 51.4f
C1836 x4.x5[7].floating.n92 VSS 2.8f
C1837 x4.x5[7].floating.n93 VSS 1.06f
C1838 x4.x5[7].floating.n94 VSS 0.366f
C1839 x4.x5[7].floating.t7 VSS 0.859f
C1840 x4.x5[7].floating.n95 VSS 6.65f
C1841 x4.x5[7].floating.n96 VSS 1.21f
C1842 x4.x5[7].floating.n97 VSS 1.17f
C1843 x4.x5[7].floating.n98 VSS 2.18f
C1844 x4.x5[7].floating.n99 VSS 1.06f
C1845 x4.x5[7].floating.n100 VSS 2.21f
C1846 x4.x5[7].floating.n101 VSS -8.01f
C1847 x4.x5[7].floating.n102 VSS -28.9f
C1848 x4.x5[7].floating.n103 VSS 3.83f
C1849 x4.x5[7].floating.n104 VSS -7.07f
C1850 x4.x5[7].floating.n105 VSS -28.3f
C1851 x4.x5[7].floating.n106 VSS 2.79f
C1852 x4.x5[7].floating.n107 VSS 1.06f
C1853 x4.x5[7].floating.n108 VSS 0.364f
C1854 x4.x5[7].floating.t6 VSS 0.859f
C1855 x4.x5[7].floating.n109 VSS 6.48f
C1856 x4.x5[7].floating.n110 VSS 1.15f
C1857 x4.x5[7].floating.n111 VSS 1.36f
C1858 x4.x5[7].floating.n112 VSS 2.2f
C1859 x4.x5[7].floating.n113 VSS 1.06f
C1860 x4.x5[7].floating.n114 VSS 2.23f
C1861 x4.x5[7].floating.n115 VSS -7.99f
C1862 x4.x5[7].floating.n116 VSS -28.9f
C1863 x4.x5[7].floating.n117 VSS 3.83f
C1864 x4.x5[7].floating.n118 VSS -7.07f
C1865 x4.x5[7].floating.n119 VSS -28.3f
C1866 x4.x5[7].floating.n120 VSS 52.7f
C1867 x4.x5[7].floating.n121 VSS 52f
C1868 x4.x5[7].floating.n122 VSS 3.23f
C1869 x4.x5[7].floating.n123 VSS -7.84f
C1870 x4.x5[7].floating.n124 VSS -28.9f
C1871 x4.x5[7].floating.n125 VSS 3.83f
C1872 x4.x5[7].floating.n126 VSS -5.01f
C1873 x4.x5[7].floating.n127 VSS -33f
C1874 x4.x5[7].floating.n128 VSS 0.766f
C1875 x4.x5[7].floating.n129 VSS 2.47f
C1876 x4.x5[7].floating.n130 VSS 51.5f
C1877 x4.x5[7].floating.n131 VSS 2.47f
C1878 x4.x5[7].floating.n132 VSS 0.766f
C1879 x4.x5[7].floating.n133 VSS -33.5f
C1880 x4.x5[7].floating.n134 VSS -4.56f
C1881 x4.x5[7].floating.n135 VSS 3.83f
C1882 x4.x5[7].floating.n136 VSS -28.9f
C1883 x4.x5[7].floating.n137 VSS -7.07f
C1884 x4.x5[7].floating.n138 VSS 2.68f
C1885 x4.x5[7].floating.n139 VSS 52f
C1886 x4.x5[7].floating.n140 VSS 3.23f
C1887 x4.x5[7].floating.n141 VSS 2.23f
C1888 x4.x5[7].floating.t3 VSS 0.859f
C1889 x4.x5[7].floating.n142 VSS 6.48f
C1890 x4.x5[7].floating.n143 VSS 1.15f
C1891 x4.x5[7].floating.n144 VSS 1.36f
C1892 x4.x5[7].floating.n145 VSS 2.2f
C1893 x4.x5[7].floating.n146 VSS 1.06f
C1894 x4.x5[7].floating.n147 VSS 0.364f
C1895 x4.x5[7].floating.n148 VSS 1.06f
C1896 x4.x5[7].floating.n149 VSS 2.79f
C1897 x4.x5[7].floating.n150 VSS 51.4f
C1898 x4.x5[7].floating.n151 VSS 2.8f
C1899 x4.x5[7].floating.n152 VSS 1.06f
C1900 x4.x5[7].floating.n153 VSS 0.366f
C1901 x4.x5[7].floating.t2 VSS 0.859f
C1902 x4.x5[7].floating.n154 VSS 7.16f
C1903 x4.x5[7].floating.n155 VSS 1.21f
C1904 x4.x5[7].floating.n156 VSS 1.17f
C1905 x4.x5[7].floating.n157 VSS 1.67f
C1906 x4.x5[7].floating.n158 VSS 1.06f
C1907 x4.x5[7].floating.n159 VSS -17.4f
C1908 x4.x5[7].floating.n160 VSS -17.2f
C1909 x4.x5[7].floating.n161 VSS -43.6f
C1910 x4.x5[7].floating.n162 VSS 0.766f
C1911 x4.x5[7].floating.n163 VSS 2.47f
C1912 x4.x5[7].floating.n164 VSS 51.5f
C1913 x4.x5[7].floating.n165 VSS 2.47f
C1914 x4.x5[7].floating.n166 VSS 0.766f
C1915 x4.x5[7].floating.n167 VSS -33f
C1916 x4.x5[7].floating.n168 VSS -5.01f
C1917 x4.x5[7].floating.n169 VSS 3.83f
C1918 x4.x5[7].floating.n170 VSS -28.9f
C1919 x4.x5[7].floating.n171 VSS -7.84f
C1920 x4.x10.Y.t0 VSS 0.0462f
C1921 x4.x10.Y.t5 VSS 0.0167f
C1922 x4.x10.Y.t8 VSS 0.0167f
C1923 x4.x10.Y.t9 VSS 0.0167f
C1924 x4.x10.Y.t2 VSS 0.0167f
C1925 x4.x10.Y.t3 VSS 0.0167f
C1926 x4.x10.Y.t4 VSS 0.0167f
C1927 x4.x10.Y.t6 VSS 0.0167f
C1928 x4.x10.Y.t7 VSS 0.0167f
C1929 x4.x10.Y.n0 VSS 0.222f
C1930 x4.x10.Y.n1 VSS 0.0366f
C1931 x4.x10.Y.t1 VSS 0.0174f
C1932 x4.x10.Y.n2 VSS 0.0188f
C1933 x4.x10.Y.n3 VSS 0.0186f
C1934 x4.x10.Y.n4 VSS 0.0151f
C1935 x4.x10.Y.n5 VSS 0.0211f
C1936 sample_code1[1].t1 VSS 0.0649f
C1937 sample_code1[1].t0 VSS 0.0648f
C1938 sample_code1[1].n0 VSS 1.78f
C1939 x2.x5[7].floating.n0 VSS 2.8f
C1940 x2.x5[7].floating.n1 VSS 51.4f
C1941 x2.x5[7].floating.n2 VSS 2.79f
C1942 x2.x5[7].floating.n3 VSS 1.06f
C1943 x2.x5[7].floating.n4 VSS 0.367f
C1944 x2.x5[7].floating.n5 VSS 1.17f
C1945 x2.x5[7].floating.t2 VSS 0.859f
C1946 x2.x5[7].floating.n6 VSS 6.5f
C1947 x2.x5[7].floating.n7 VSS 1.36f
C1948 x2.x5[7].floating.n8 VSS 2.19f
C1949 x2.x5[7].floating.n9 VSS 1.06f
C1950 x2.x5[7].floating.n10 VSS -15.2f
C1951 x2.x5[7].floating.n11 VSS -15.2f
C1952 x2.x5[7].floating.n12 VSS -41.6f
C1953 x2.x5[7].floating.n13 VSS 0.766f
C1954 x2.x5[7].floating.n14 VSS 2.47f
C1955 x2.x5[7].floating.n15 VSS 51.5f
C1956 x2.x5[7].floating.n16 VSS 2.47f
C1957 x2.x5[7].floating.n17 VSS 0.766f
C1958 x2.x5[7].floating.n18 VSS -33.5f
C1959 x2.x5[7].floating.n19 VSS -4.56f
C1960 x2.x5[7].floating.n20 VSS 3.83f
C1961 x2.x5[7].floating.n21 VSS -28.9f
C1962 x2.x5[7].floating.n22 VSS -7.07f
C1963 x2.x5[7].floating.n23 VSS 2.68f
C1964 x2.x5[7].floating.n24 VSS 1.06f
C1965 x2.x5[7].floating.n25 VSS 0.364f
C1966 x2.x5[7].floating.n26 VSS 1.21f
C1967 x2.x5[7].floating.t1 VSS 0.859f
C1968 x2.x5[7].floating.n27 VSS 6.67f
C1969 x2.x5[7].floating.n28 VSS 1.15f
C1970 x2.x5[7].floating.n29 VSS 2.17f
C1971 x2.x5[7].floating.n30 VSS 1.06f
C1972 x2.x5[7].floating.n31 VSS 2.22f
C1973 x2.x5[7].floating.n32 VSS -8.01f
C1974 x2.x5[7].floating.n33 VSS -28.9f
C1975 x2.x5[7].floating.n34 VSS 3.83f
C1976 x2.x5[7].floating.n35 VSS -7.07f
C1977 x2.x5[7].floating.n36 VSS -28.3f
C1978 x2.x5[7].floating.n37 VSS 52.7f
C1979 x2.x5[7].floating.n38 VSS -28.3f
C1980 x2.x5[7].floating.n39 VSS -7.07f
C1981 x2.x5[7].floating.n40 VSS 3.83f
C1982 x2.x5[7].floating.n41 VSS -28.9f
C1983 x2.x5[7].floating.n42 VSS -7.99f
C1984 x2.x5[7].floating.n43 VSS 2.22f
C1985 x2.x5[7].floating.n44 VSS 1.17f
C1986 x2.x5[7].floating.t4 VSS 0.859f
C1987 x2.x5[7].floating.n45 VSS 6.5f
C1988 x2.x5[7].floating.n46 VSS 1.36f
C1989 x2.x5[7].floating.n47 VSS 2.19f
C1990 x2.x5[7].floating.n48 VSS 1.06f
C1991 x2.x5[7].floating.n49 VSS 0.367f
C1992 x2.x5[7].floating.n50 VSS 1.06f
C1993 x2.x5[7].floating.n51 VSS 2.79f
C1994 x2.x5[7].floating.n52 VSS 51.4f
C1995 x2.x5[7].floating.n53 VSS 2.8f
C1996 x2.x5[7].floating.n54 VSS 1.06f
C1997 x2.x5[7].floating.n55 VSS 0.364f
C1998 x2.x5[7].floating.n56 VSS 1.21f
C1999 x2.x5[7].floating.t7 VSS 0.859f
C2000 x2.x5[7].floating.n57 VSS 6.67f
C2001 x2.x5[7].floating.n58 VSS 1.15f
C2002 x2.x5[7].floating.n59 VSS 2.17f
C2003 x2.x5[7].floating.n60 VSS 1.06f
C2004 x2.x5[7].floating.n61 VSS 2.22f
C2005 x2.x5[7].floating.n62 VSS -8.01f
C2006 x2.x5[7].floating.n63 VSS -28.9f
C2007 x2.x5[7].floating.n64 VSS 3.83f
C2008 x2.x5[7].floating.n65 VSS -7.07f
C2009 x2.x5[7].floating.n66 VSS -28.3f
C2010 x2.x5[7].floating.n67 VSS 52.7f
C2011 x2.x5[7].floating.n68 VSS -28.3f
C2012 x2.x5[7].floating.n69 VSS -7.07f
C2013 x2.x5[7].floating.n70 VSS 3.83f
C2014 x2.x5[7].floating.n71 VSS -28.9f
C2015 x2.x5[7].floating.n72 VSS -7.99f
C2016 x2.x5[7].floating.n73 VSS 2.22f
C2017 x2.x5[7].floating.n74 VSS 1.17f
C2018 x2.x5[7].floating.t5 VSS 0.859f
C2019 x2.x5[7].floating.n75 VSS 6.5f
C2020 x2.x5[7].floating.n76 VSS 1.36f
C2021 x2.x5[7].floating.n77 VSS 2.19f
C2022 x2.x5[7].floating.n78 VSS 1.06f
C2023 x2.x5[7].floating.n79 VSS 0.367f
C2024 x2.x5[7].floating.n80 VSS 1.06f
C2025 x2.x5[7].floating.n81 VSS 2.79f
C2026 x2.x5[7].floating.n82 VSS 51.4f
C2027 x2.x5[7].floating.n83 VSS 2.8f
C2028 x2.x5[7].floating.n84 VSS 1.06f
C2029 x2.x5[7].floating.n85 VSS 0.364f
C2030 x2.x5[7].floating.n86 VSS 1.21f
C2031 x2.x5[7].floating.t0 VSS 0.859f
C2032 x2.x5[7].floating.n87 VSS 6.67f
C2033 x2.x5[7].floating.n88 VSS 1.15f
C2034 x2.x5[7].floating.n89 VSS 2.17f
C2035 x2.x5[7].floating.n90 VSS 1.06f
C2036 x2.x5[7].floating.n91 VSS 2.22f
C2037 x2.x5[7].floating.n92 VSS -8.01f
C2038 x2.x5[7].floating.n93 VSS -28.9f
C2039 x2.x5[7].floating.n94 VSS 3.83f
C2040 x2.x5[7].floating.n95 VSS -7.07f
C2041 x2.x5[7].floating.n96 VSS -28.3f
C2042 x2.x5[7].floating.n97 VSS 52.7f
C2043 x2.x5[7].floating.n98 VSS -28.3f
C2044 x2.x5[7].floating.n99 VSS -7.07f
C2045 x2.x5[7].floating.n100 VSS 3.83f
C2046 x2.x5[7].floating.n101 VSS -28.9f
C2047 x2.x5[7].floating.n102 VSS -7.99f
C2048 x2.x5[7].floating.n103 VSS 2.22f
C2049 x2.x5[7].floating.n104 VSS 1.17f
C2050 x2.x5[7].floating.t3 VSS 0.859f
C2051 x2.x5[7].floating.n105 VSS 6.5f
C2052 x2.x5[7].floating.n106 VSS 1.36f
C2053 x2.x5[7].floating.n107 VSS 2.19f
C2054 x2.x5[7].floating.n108 VSS 1.06f
C2055 x2.x5[7].floating.n109 VSS 0.367f
C2056 x2.x5[7].floating.n110 VSS 1.06f
C2057 x2.x5[7].floating.n111 VSS 2.79f
C2058 x2.x5[7].floating.n112 VSS 51.4f
C2059 x2.x5[7].floating.n113 VSS 2.8f
C2060 x2.x5[7].floating.n114 VSS 1.06f
C2061 x2.x5[7].floating.n115 VSS 0.366f
C2062 x2.x5[7].floating.t6 VSS 0.859f
C2063 x2.x5[7].floating.n116 VSS 7.13f
C2064 x2.x5[7].floating.n117 VSS 1.21f
C2065 x2.x5[7].floating.n118 VSS 1.16f
C2066 x2.x5[7].floating.n119 VSS 1.7f
C2067 x2.x5[7].floating.n120 VSS 1.06f
C2068 x2.x5[7].floating.n121 VSS -17.4f
C2069 x2.x5[7].floating.n122 VSS -17.2f
C2070 x2.x5[7].floating.n123 VSS -43.6f
C2071 x2.x5[7].floating.n124 VSS 0.766f
C2072 x2.x5[7].floating.n125 VSS 2.47f
C2073 x2.x5[7].floating.n126 VSS 51.5f
C2074 x2.x5[7].floating.n127 VSS 2.47f
C2075 x2.x5[7].floating.n128 VSS 0.766f
C2076 x2.x5[7].floating.n129 VSS -33f
C2077 x2.x5[7].floating.n130 VSS -5.01f
C2078 x2.x5[7].floating.n131 VSS 3.83f
C2079 x2.x5[7].floating.n132 VSS -28.9f
C2080 x2.x5[7].floating.n133 VSS -7.84f
C2081 x2.x5[7].floating.n134 VSS 3.23f
C2082 x2.x5[7].floating.n135 VSS 52f
C2083 x2.x5[7].floating.n136 VSS 2.68f
C2084 x2.x5[7].floating.n137 VSS -7.07f
C2085 x2.x5[7].floating.n138 VSS -28.9f
C2086 x2.x5[7].floating.n139 VSS 3.83f
C2087 x2.x5[7].floating.n140 VSS -4.56f
C2088 x2.x5[7].floating.n141 VSS -33.5f
C2089 x2.x5[7].floating.n142 VSS 0.766f
C2090 x2.x5[7].floating.n143 VSS 2.47f
C2091 x2.x5[7].floating.n144 VSS 51.5f
C2092 x2.x5[7].floating.n145 VSS 2.47f
C2093 x2.x5[7].floating.n146 VSS 0.766f
C2094 x2.x5[7].floating.n147 VSS -33f
C2095 x2.x5[7].floating.n148 VSS -5.01f
C2096 x2.x5[7].floating.n149 VSS 3.83f
C2097 x2.x5[7].floating.n150 VSS -28.9f
C2098 x2.x5[7].floating.n151 VSS -7.84f
C2099 x2.x5[7].floating.n152 VSS 3.23f
C2100 x2.x5[7].floating.n153 VSS 52f
C2101 x2.x5[7].floating.n154 VSS 2.68f
C2102 x2.x5[7].floating.n155 VSS -7.07f
C2103 x2.x5[7].floating.n156 VSS -28.9f
C2104 x2.x5[7].floating.n157 VSS 3.83f
C2105 x2.x5[7].floating.n158 VSS -4.56f
C2106 x2.x5[7].floating.n159 VSS -33.5f
C2107 x2.x5[7].floating.n160 VSS 0.766f
C2108 x2.x5[7].floating.n161 VSS 2.47f
C2109 x2.x5[7].floating.n162 VSS 51.5f
C2110 x2.x5[7].floating.n163 VSS 2.47f
C2111 x2.x5[7].floating.n164 VSS 0.766f
C2112 x2.x5[7].floating.n165 VSS -33f
C2113 x2.x5[7].floating.n166 VSS -5.01f
C2114 x2.x5[7].floating.n167 VSS 3.83f
C2115 x2.x5[7].floating.n168 VSS -28.9f
C2116 x2.x5[7].floating.n169 VSS -7.84f
C2117 x2.x5[7].floating.n170 VSS 3.23f
C2118 x2.x5[7].floating.n171 VSS 52f
C2119 x2.x10.Y.n0 VSS 0.0359f
C2120 x2.x10.Y.t0 VSS 0.0526f
C2121 x2.x10.Y.n1 VSS 0.0169f
C2122 x2.x10.Y.n2 VSS 0.00704f
C2123 x2.x10.Y.t1 VSS 0.0181f
C2124 x2.x10.Y.n3 VSS 0.0188f
C2125 x2.x10.Y.n4 VSS 0.019f
C2126 x2.x10.Y.n5 VSS 0.221f
C2127 x2.x10.Y.t7 VSS 0.0167f
C2128 x2.x10.Y.t8 VSS 0.0167f
C2129 x2.x10.Y.t5 VSS 0.0167f
C2130 x2.x10.Y.t2 VSS 0.0167f
C2131 x2.x10.Y.t4 VSS 0.0167f
C2132 x2.x10.Y.t9 VSS 0.0167f
C2133 x2.x10.Y.t6 VSS 0.0167f
C2134 x2.x10.Y.t3 VSS 0.0167f
C2135 VDD.t43 VSS 0.0509f
C2136 VDD.n0 VSS 0.0561f
C2137 VDD.n1 VSS 0.00873f
C2138 VDD.n2 VSS 0.00407f
C2139 VDD.n3 VSS 0.00443f
C2140 VDD.n4 VSS 0.00672f
C2141 VDD.n5 VSS 0.0277f
C2142 VDD.n6 VSS 0.0111f
C2143 VDD.n7 VSS 0.0122f
C2144 VDD.n8 VSS 0.0158f
C2145 VDD.n9 VSS 0.307f
C2146 VDD.n10 VSS 0.00302f
C2147 VDD.n11 VSS 0.00277f
C2148 VDD.n12 VSS 2.54f
C2149 VDD.n13 VSS 0.0129f
C2150 VDD.n15 VSS 0.0129f
C2151 VDD.n19 VSS 0.0129f
C2152 VDD.n22 VSS 0.00277f
C2153 VDD.n23 VSS 0.0576f
C2154 VDD.n24 VSS 0.00979f
C2155 VDD.n25 VSS 0.00269f
C2156 VDD.n26 VSS 0.00277f
C2157 VDD.n27 VSS 0.00269f
C2158 VDD.n28 VSS 0.00269f
C2159 VDD.n29 VSS 4.74e-19
C2160 VDD.n30 VSS 0.00663f
C2161 VDD.n31 VSS 0.00332f
C2162 VDD.n32 VSS 0.00806f
C2163 VDD.n33 VSS 0.00439f
C2164 VDD.n34 VSS 0.00781f
C2165 VDD.n35 VSS 0.0226f
C2166 VDD.n36 VSS -0.211f
C2167 VDD.n37 VSS 0.0139f
C2168 VDD.n38 VSS 3.26e-19
C2169 VDD.n39 VSS 0.0141f
C2170 VDD.n40 VSS 0.00439f
C2171 VDD.n41 VSS 0.00332f
C2172 VDD.n42 VSS 0.00269f
C2173 VDD.n43 VSS 4.74e-19
C2174 VDD.n44 VSS 0.00269f
C2175 VDD.n45 VSS 0.00277f
C2176 VDD.n46 VSS 0.00269f
C2177 VDD.n47 VSS 0.00916f
C2178 VDD.n48 VSS 0.00411f
C2179 VDD.n49 VSS 0.00439f
C2180 VDD.n50 VSS 0.00781f
C2181 VDD.n51 VSS 0.0223f
C2182 VDD.n52 VSS 0.00781f
C2183 VDD.n53 VSS 0.00348f
C2184 VDD.n54 VSS 0.00332f
C2185 VDD.n55 VSS 0.00269f
C2186 VDD.n56 VSS 0.00269f
C2187 VDD.n57 VSS 0.00979f
C2188 VDD.n58 VSS 0.0104f
C2189 VDD.n59 VSS 0.00269f
C2190 VDD.n60 VSS 0.00269f
C2191 VDD.n61 VSS 4.74e-19
C2192 VDD.n62 VSS 0.00979f
C2193 VDD.n63 VSS 0.00332f
C2194 VDD.n64 VSS 0.00663f
C2195 VDD.n65 VSS 0.00332f
C2196 VDD.n66 VSS 0.00806f
C2197 VDD.n67 VSS -0.0753f
C2198 VDD.n68 VSS 0.0223f
C2199 VDD.n69 VSS 0.00488f
C2200 VDD.n70 VSS -0.0782f
C2201 VDD.n71 VSS 3.26e-19
C2202 VDD.n72 VSS 4.74e-19
C2203 VDD.n73 VSS 0.00585f
C2204 VDD.n74 VSS 0.00348f
C2205 VDD.n75 VSS 0.00269f
C2206 VDD.n76 VSS 0.0129f
C2207 VDD.n77 VSS 0.00979f
C2208 VDD.n78 VSS 0.00332f
C2209 VDD.n79 VSS 0.00585f
C2210 VDD.n80 VSS 0.00348f
C2211 VDD.n81 VSS 4.74e-19
C2212 VDD.n82 VSS 3.26e-19
C2213 VDD.n83 VSS 0.00488f
C2214 VDD.n84 VSS 0.0227f
C2215 VDD.n85 VSS -0.0753f
C2216 VDD.n86 VSS 0.00411f
C2217 VDD.n87 VSS 0.00348f
C2218 VDD.n88 VSS 0.00916f
C2219 VDD.n89 VSS 0.00269f
C2220 VDD.n90 VSS 0.00979f
C2221 VDD.n91 VSS 0.00979f
C2222 VDD.n92 VSS 0.00269f
C2223 VDD.n93 VSS 0.00269f
C2224 VDD.n94 VSS 0.00269f
C2225 VDD.n95 VSS 0.00269f
C2226 VDD.n96 VSS 0.00348f
C2227 VDD.n97 VSS 0.00332f
C2228 VDD.n98 VSS 0.0285f
C2229 VDD.n99 VSS 0.0141f
C2230 VDD.n100 VSS 3.26e-19
C2231 VDD.n101 VSS 0.00332f
C2232 VDD.n102 VSS 0.00348f
C2233 VDD.n103 VSS 0.00916f
C2234 VDD.n104 VSS 0.00269f
C2235 VDD.n105 VSS 0.00269f
C2236 VDD.n106 VSS 0.0294f
C2237 VDD.n107 VSS 0.00332f
C2238 VDD.n108 VSS 0.0261f
C2239 VDD.n109 VSS 0.0286f
C2240 VDD.n110 VSS 0.0286f
C2241 VDD.n111 VSS 0.0261f
C2242 VDD.n112 VSS 0.00332f
C2243 VDD.n113 VSS 0.0294f
C2244 VDD.n114 VSS 0.00269f
C2245 VDD.n116 VSS 0.00269f
C2246 VDD.n117 VSS 0.00269f
C2247 VDD.n118 VSS 0.00348f
C2248 VDD.n119 VSS 0.00411f
C2249 VDD.n120 VSS 0.00374f
C2250 VDD.n121 VSS 0.0141f
C2251 VDD.n122 VSS 3.26e-19
C2252 VDD.n123 VSS 0.00332f
C2253 VDD.n124 VSS 0.00916f
C2254 VDD.n125 VSS 0.00269f
C2255 VDD.n126 VSS 0.0104f
C2256 VDD.n127 VSS 0.00269f
C2257 VDD.n128 VSS 0.00269f
C2258 VDD.n129 VSS 0.00348f
C2259 VDD.n130 VSS 0.00411f
C2260 VDD.n131 VSS 0.00374f
C2261 VDD.n132 VSS -0.0845f
C2262 VDD.n133 VSS 3.26e-19
C2263 VDD.n134 VSS 0.00332f
C2264 VDD.n135 VSS 0.00916f
C2265 VDD.n136 VSS 0.00979f
C2266 VDD.n137 VSS 0.00277f
C2267 VDD.n138 VSS 0.00269f
C2268 VDD.n139 VSS 0.00269f
C2269 VDD.n140 VSS 0.00916f
C2270 VDD.n141 VSS 4.74e-19
C2271 VDD.n142 VSS 0.00979f
C2272 VDD.n143 VSS 0.00332f
C2273 VDD.n144 VSS 0.00411f
C2274 VDD.n145 VSS 0.00374f
C2275 VDD.n146 VSS 0.0141f
C2276 VDD.n147 VSS -0.211f
C2277 VDD.n148 VSS 0.0136f
C2278 VDD.n149 VSS 0.00348f
C2279 VDD.n150 VSS 0.00269f
C2280 VDD.n151 VSS 0.00269f
C2281 VDD.n152 VSS 0.00277f
C2282 VDD.n153 VSS 0.00269f
C2283 VDD.n154 VSS 0.00916f
C2284 VDD.n155 VSS 0.00332f
C2285 VDD.n156 VSS 3.26e-19
C2286 VDD.n157 VSS 0.00374f
C2287 VDD.n158 VSS 0.0223f
C2288 VDD.n159 VSS 0.00374f
C2289 VDD.n160 VSS 0.00348f
C2290 VDD.n161 VSS 0.00269f
C2291 VDD.n162 VSS 0.00269f
C2292 VDD.n163 VSS 0.00277f
C2293 VDD.n164 VSS 0.00269f
C2294 VDD.n165 VSS 0.0295f
C2295 VDD.n166 VSS 0.00332f
C2296 VDD.n167 VSS 3.26e-19
C2297 VDD.n168 VSS 0.0141f
C2298 VDD.n169 VSS 0.0241f
C2299 VDD.n170 VSS 0.00411f
C2300 VDD.n171 VSS 0.00439f
C2301 VDD.n172 VSS -0.182f
C2302 VDD.n173 VSS 0.00781f
C2303 VDD.n174 VSS 0.00348f
C2304 VDD.n175 VSS 0.00332f
C2305 VDD.n176 VSS 0.00269f
C2306 VDD.n177 VSS 0.0295f
C2307 VDD.n178 VSS 0.00269f
C2308 VDD.n179 VSS 0.00269f
C2309 VDD.n180 VSS 0.00277f
C2310 VDD.n181 VSS 0.00269f
C2311 VDD.n182 VSS 0.00916f
C2312 VDD.n183 VSS 0.00411f
C2313 VDD.n184 VSS 0.00439f
C2314 VDD.n185 VSS 0.0223f
C2315 VDD.n186 VSS 0.00781f
C2316 VDD.n187 VSS 0.00348f
C2317 VDD.n188 VSS 0.00332f
C2318 VDD.n189 VSS 0.00269f
C2319 VDD.n190 VSS 0.00269f
C2320 VDD.n191 VSS 0.00979f
C2321 VDD.n192 VSS 0.0104f
C2322 VDD.n193 VSS 0.00269f
C2323 VDD.n194 VSS 0.00269f
C2324 VDD.n195 VSS 4.74e-19
C2325 VDD.n196 VSS 0.00979f
C2326 VDD.n197 VSS 0.00332f
C2327 VDD.n198 VSS 0.00663f
C2328 VDD.n199 VSS 0.00332f
C2329 VDD.n200 VSS 0.00806f
C2330 VDD.n201 VSS -0.0753f
C2331 VDD.n202 VSS 0.0223f
C2332 VDD.n203 VSS 0.00488f
C2333 VDD.n204 VSS -0.0782f
C2334 VDD.n205 VSS 3.26e-19
C2335 VDD.n206 VSS 4.74e-19
C2336 VDD.n207 VSS 0.00585f
C2337 VDD.n208 VSS 0.00348f
C2338 VDD.n209 VSS 0.00269f
C2339 VDD.n210 VSS 0.0129f
C2340 VDD.n211 VSS 0.00979f
C2341 VDD.n212 VSS 0.00332f
C2342 VDD.n213 VSS 0.00585f
C2343 VDD.n214 VSS 0.00348f
C2344 VDD.n215 VSS 4.74e-19
C2345 VDD.n216 VSS 3.26e-19
C2346 VDD.n217 VSS 0.00488f
C2347 VDD.n218 VSS 0.0227f
C2348 VDD.n219 VSS -0.0753f
C2349 VDD.n220 VSS 0.00411f
C2350 VDD.n221 VSS 0.00348f
C2351 VDD.n222 VSS 0.00916f
C2352 VDD.n223 VSS 0.00269f
C2353 VDD.n224 VSS 0.00979f
C2354 VDD.n225 VSS 0.00979f
C2355 VDD.n226 VSS 0.00269f
C2356 VDD.n227 VSS 0.00269f
C2357 VDD.n228 VSS 0.00269f
C2358 VDD.n229 VSS 0.00269f
C2359 VDD.n230 VSS 0.00348f
C2360 VDD.n231 VSS 0.00332f
C2361 VDD.n232 VSS 0.0285f
C2362 VDD.n233 VSS 0.0141f
C2363 VDD.n234 VSS 3.26e-19
C2364 VDD.n235 VSS 0.00332f
C2365 VDD.n236 VSS 0.00348f
C2366 VDD.n237 VSS 0.00916f
C2367 VDD.n238 VSS 0.00269f
C2368 VDD.n239 VSS 0.00269f
C2369 VDD.n240 VSS 0.0294f
C2370 VDD.n241 VSS 0.00332f
C2371 VDD.n242 VSS 0.0261f
C2372 VDD.n243 VSS 0.0286f
C2373 VDD.n244 VSS 0.0286f
C2374 VDD.n245 VSS 0.0261f
C2375 VDD.n246 VSS 0.00332f
C2376 VDD.n247 VSS 0.0294f
C2377 VDD.n248 VSS 0.00269f
C2378 VDD.n250 VSS 0.00269f
C2379 VDD.n251 VSS 0.00269f
C2380 VDD.n252 VSS 0.00348f
C2381 VDD.n253 VSS 0.00411f
C2382 VDD.n254 VSS 0.00374f
C2383 VDD.n255 VSS 0.0141f
C2384 VDD.n256 VSS 3.26e-19
C2385 VDD.n257 VSS 0.00332f
C2386 VDD.n258 VSS 0.00916f
C2387 VDD.n259 VSS 0.00269f
C2388 VDD.n260 VSS 0.0104f
C2389 VDD.n261 VSS 0.00269f
C2390 VDD.n262 VSS 0.00269f
C2391 VDD.n263 VSS 0.00348f
C2392 VDD.n264 VSS 0.00411f
C2393 VDD.n265 VSS 0.00374f
C2394 VDD.n266 VSS -0.0845f
C2395 VDD.n267 VSS 3.26e-19
C2396 VDD.n268 VSS 0.00332f
C2397 VDD.n269 VSS 0.00916f
C2398 VDD.n270 VSS 0.00979f
C2399 VDD.n271 VSS 0.00277f
C2400 VDD.n272 VSS 0.00269f
C2401 VDD.n273 VSS 0.00269f
C2402 VDD.n274 VSS 0.00916f
C2403 VDD.n275 VSS 4.74e-19
C2404 VDD.n276 VSS 0.00979f
C2405 VDD.n277 VSS 0.00332f
C2406 VDD.n278 VSS 0.00411f
C2407 VDD.n279 VSS 0.00374f
C2408 VDD.n280 VSS 0.0141f
C2409 VDD.n281 VSS -0.211f
C2410 VDD.n282 VSS 0.0136f
C2411 VDD.n283 VSS 0.00348f
C2412 VDD.n284 VSS 0.00269f
C2413 VDD.n285 VSS 0.00269f
C2414 VDD.n286 VSS 0.00277f
C2415 VDD.n287 VSS 0.00269f
C2416 VDD.n288 VSS 0.00916f
C2417 VDD.n289 VSS 0.00332f
C2418 VDD.n290 VSS 3.26e-19
C2419 VDD.n291 VSS 0.00374f
C2420 VDD.n292 VSS 0.0223f
C2421 VDD.n293 VSS 0.00374f
C2422 VDD.n294 VSS 0.00348f
C2423 VDD.n295 VSS 0.00269f
C2424 VDD.n296 VSS 0.00269f
C2425 VDD.n297 VSS 0.00277f
C2426 VDD.n298 VSS 0.00269f
C2427 VDD.n299 VSS 0.0295f
C2428 VDD.n300 VSS 0.00332f
C2429 VDD.n301 VSS 3.26e-19
C2430 VDD.n302 VSS 0.0141f
C2431 VDD.n303 VSS 0.0241f
C2432 VDD.n304 VSS 0.00411f
C2433 VDD.n305 VSS 0.00439f
C2434 VDD.n306 VSS -0.182f
C2435 VDD.n307 VSS 0.00781f
C2436 VDD.n308 VSS 0.00348f
C2437 VDD.n309 VSS 0.00332f
C2438 VDD.n310 VSS 0.00269f
C2439 VDD.n311 VSS 0.0295f
C2440 VDD.n312 VSS 0.00269f
C2441 VDD.n313 VSS 0.00269f
C2442 VDD.n314 VSS 0.00277f
C2443 VDD.n315 VSS 0.00269f
C2444 VDD.n316 VSS 0.00916f
C2445 VDD.n317 VSS 0.00411f
C2446 VDD.n318 VSS 0.00439f
C2447 VDD.n319 VSS 0.0223f
C2448 VDD.n320 VSS 0.00781f
C2449 VDD.n321 VSS 0.00348f
C2450 VDD.n322 VSS 0.00332f
C2451 VDD.n323 VSS 0.00269f
C2452 VDD.n324 VSS 0.00269f
C2453 VDD.n325 VSS 0.00979f
C2454 VDD.n326 VSS 0.0104f
C2455 VDD.n327 VSS 0.00269f
C2456 VDD.n328 VSS 0.00269f
C2457 VDD.n329 VSS 4.74e-19
C2458 VDD.n330 VSS 0.00979f
C2459 VDD.n331 VSS 0.00332f
C2460 VDD.n332 VSS 0.00663f
C2461 VDD.n333 VSS 0.00332f
C2462 VDD.n334 VSS 0.00806f
C2463 VDD.n335 VSS -0.0753f
C2464 VDD.n336 VSS 0.0223f
C2465 VDD.n337 VSS 0.00488f
C2466 VDD.n338 VSS -0.0782f
C2467 VDD.n339 VSS 3.26e-19
C2468 VDD.n340 VSS 4.74e-19
C2469 VDD.n341 VSS 0.00585f
C2470 VDD.n342 VSS 0.00348f
C2471 VDD.n343 VSS 0.00269f
C2472 VDD.n344 VSS 0.0129f
C2473 VDD.n345 VSS 0.00979f
C2474 VDD.n346 VSS 0.00332f
C2475 VDD.n347 VSS 0.00585f
C2476 VDD.n348 VSS 0.00348f
C2477 VDD.n349 VSS 4.74e-19
C2478 VDD.n350 VSS 3.26e-19
C2479 VDD.n351 VSS 0.00488f
C2480 VDD.n352 VSS 0.0227f
C2481 VDD.n353 VSS -0.0753f
C2482 VDD.n354 VSS 0.00411f
C2483 VDD.n355 VSS 0.00348f
C2484 VDD.n356 VSS 0.00916f
C2485 VDD.n357 VSS 0.00269f
C2486 VDD.n358 VSS 0.00979f
C2487 VDD.n359 VSS 0.00979f
C2488 VDD.n360 VSS 0.00269f
C2489 VDD.n361 VSS 0.00269f
C2490 VDD.n362 VSS 0.00269f
C2491 VDD.n363 VSS 0.00269f
C2492 VDD.n364 VSS 0.00348f
C2493 VDD.n365 VSS 0.00332f
C2494 VDD.n366 VSS 0.0285f
C2495 VDD.n367 VSS 0.0141f
C2496 VDD.n368 VSS 3.26e-19
C2497 VDD.n369 VSS 0.00332f
C2498 VDD.n370 VSS 0.00348f
C2499 VDD.n371 VSS 0.00916f
C2500 VDD.n372 VSS 0.00269f
C2501 VDD.n373 VSS 0.00269f
C2502 VDD.n374 VSS 0.0294f
C2503 VDD.n375 VSS 0.00332f
C2504 VDD.n376 VSS 0.0261f
C2505 VDD.n377 VSS 0.0286f
C2506 VDD.n378 VSS 0.0286f
C2507 VDD.n379 VSS 0.0261f
C2508 VDD.n380 VSS 0.00332f
C2509 VDD.n381 VSS 0.0294f
C2510 VDD.n382 VSS 0.00269f
C2511 VDD.n384 VSS 0.00269f
C2512 VDD.n385 VSS 0.00269f
C2513 VDD.n386 VSS 0.00348f
C2514 VDD.n387 VSS 0.00411f
C2515 VDD.n388 VSS 0.00374f
C2516 VDD.n389 VSS 0.0141f
C2517 VDD.n390 VSS 3.26e-19
C2518 VDD.n391 VSS 0.00332f
C2519 VDD.n392 VSS 0.00916f
C2520 VDD.n393 VSS 0.00269f
C2521 VDD.n394 VSS 0.0104f
C2522 VDD.n395 VSS 0.00269f
C2523 VDD.n396 VSS 0.00269f
C2524 VDD.n397 VSS 0.00348f
C2525 VDD.n398 VSS 0.00411f
C2526 VDD.n399 VSS 0.00374f
C2527 VDD.n400 VSS -0.0845f
C2528 VDD.n401 VSS 3.26e-19
C2529 VDD.n402 VSS 0.00332f
C2530 VDD.n403 VSS 0.00916f
C2531 VDD.n404 VSS 0.00979f
C2532 VDD.n405 VSS 0.00277f
C2533 VDD.n406 VSS 0.00269f
C2534 VDD.n407 VSS 0.00269f
C2535 VDD.n408 VSS 0.00916f
C2536 VDD.n409 VSS 4.74e-19
C2537 VDD.n410 VSS 0.00979f
C2538 VDD.n411 VSS 0.00332f
C2539 VDD.n412 VSS 0.00411f
C2540 VDD.n413 VSS 0.00374f
C2541 VDD.n414 VSS 0.0141f
C2542 VDD.n415 VSS -0.211f
C2543 VDD.n416 VSS 0.0136f
C2544 VDD.n417 VSS 0.00348f
C2545 VDD.n418 VSS 0.00269f
C2546 VDD.n419 VSS 0.00269f
C2547 VDD.n420 VSS 0.00277f
C2548 VDD.n421 VSS 0.00269f
C2549 VDD.n422 VSS 0.00916f
C2550 VDD.n423 VSS 0.00332f
C2551 VDD.n424 VSS 3.26e-19
C2552 VDD.n425 VSS 0.00374f
C2553 VDD.n426 VSS 0.0223f
C2554 VDD.n427 VSS 0.00374f
C2555 VDD.n428 VSS 0.00348f
C2556 VDD.n429 VSS 0.00269f
C2557 VDD.n430 VSS 0.00269f
C2558 VDD.n431 VSS 0.00277f
C2559 VDD.n432 VSS 0.00269f
C2560 VDD.n433 VSS 0.0295f
C2561 VDD.n434 VSS 0.00332f
C2562 VDD.n435 VSS 3.26e-19
C2563 VDD.n436 VSS 0.0141f
C2564 VDD.n437 VSS 0.0241f
C2565 VDD.n438 VSS 0.00411f
C2566 VDD.n439 VSS 0.00439f
C2567 VDD.n440 VSS -0.182f
C2568 VDD.n441 VSS 0.00781f
C2569 VDD.n442 VSS 0.00348f
C2570 VDD.n443 VSS 0.00332f
C2571 VDD.n444 VSS 0.00269f
C2572 VDD.n445 VSS 0.0295f
C2573 VDD.n446 VSS 0.00269f
C2574 VDD.n447 VSS 0.00269f
C2575 VDD.n448 VSS 0.00277f
C2576 VDD.n449 VSS 0.00269f
C2577 VDD.n450 VSS 0.00916f
C2578 VDD.n451 VSS 0.00411f
C2579 VDD.n452 VSS 0.00439f
C2580 VDD.n453 VSS 0.0223f
C2581 VDD.n454 VSS 0.00781f
C2582 VDD.n455 VSS 0.00348f
C2583 VDD.n456 VSS 0.00332f
C2584 VDD.n457 VSS 0.00269f
C2585 VDD.n458 VSS 0.00269f
C2586 VDD.n459 VSS 0.00979f
C2587 VDD.n460 VSS 0.0104f
C2588 VDD.n461 VSS 0.00269f
C2589 VDD.n462 VSS 0.00269f
C2590 VDD.n463 VSS 4.74e-19
C2591 VDD.n464 VSS 0.00979f
C2592 VDD.n465 VSS 0.00332f
C2593 VDD.n466 VSS 0.00663f
C2594 VDD.n467 VSS 0.00332f
C2595 VDD.n468 VSS 0.00806f
C2596 VDD.n469 VSS -0.0753f
C2597 VDD.n470 VSS 0.0223f
C2598 VDD.n471 VSS 0.00488f
C2599 VDD.n472 VSS -0.0782f
C2600 VDD.n473 VSS 3.26e-19
C2601 VDD.n474 VSS 4.74e-19
C2602 VDD.n475 VSS 0.00585f
C2603 VDD.n476 VSS 0.00348f
C2604 VDD.n477 VSS 0.00269f
C2605 VDD.n478 VSS 0.0129f
C2606 VDD.n479 VSS 0.00979f
C2607 VDD.n480 VSS 0.00332f
C2608 VDD.n481 VSS 0.00585f
C2609 VDD.n482 VSS 0.00348f
C2610 VDD.n483 VSS 4.74e-19
C2611 VDD.n484 VSS 3.26e-19
C2612 VDD.n485 VSS 0.00488f
C2613 VDD.n486 VSS 0.0227f
C2614 VDD.n487 VSS -0.0753f
C2615 VDD.n488 VSS 0.00411f
C2616 VDD.n489 VSS 0.00348f
C2617 VDD.n490 VSS 0.00916f
C2618 VDD.n491 VSS 0.00269f
C2619 VDD.n492 VSS 0.00979f
C2620 VDD.n493 VSS 0.00979f
C2621 VDD.n494 VSS 0.00269f
C2622 VDD.n495 VSS 0.00269f
C2623 VDD.n496 VSS 0.00269f
C2624 VDD.n497 VSS 0.00269f
C2625 VDD.n498 VSS 0.00348f
C2626 VDD.n499 VSS 0.00332f
C2627 VDD.n500 VSS 0.0285f
C2628 VDD.n501 VSS 0.0141f
C2629 VDD.n502 VSS 3.26e-19
C2630 VDD.n503 VSS 0.00332f
C2631 VDD.n504 VSS 0.00348f
C2632 VDD.n505 VSS 0.00916f
C2633 VDD.n506 VSS 0.00269f
C2634 VDD.n507 VSS 0.00269f
C2635 VDD.n508 VSS 0.0294f
C2636 VDD.n509 VSS 0.00332f
C2637 VDD.n510 VSS 0.0261f
C2638 VDD.n511 VSS 0.0286f
C2639 VDD.n512 VSS 0.0286f
C2640 VDD.n513 VSS 0.0261f
C2641 VDD.n514 VSS 0.00332f
C2642 VDD.n515 VSS 0.0294f
C2643 VDD.n516 VSS 0.00269f
C2644 VDD.n518 VSS 0.00269f
C2645 VDD.n519 VSS 0.00269f
C2646 VDD.n520 VSS 0.00348f
C2647 VDD.n521 VSS 0.00411f
C2648 VDD.n522 VSS 0.00374f
C2649 VDD.n523 VSS 0.0141f
C2650 VDD.n524 VSS 3.26e-19
C2651 VDD.n525 VSS 0.00332f
C2652 VDD.n526 VSS 0.00916f
C2653 VDD.n527 VSS 0.00269f
C2654 VDD.n528 VSS 0.0104f
C2655 VDD.n529 VSS 0.00269f
C2656 VDD.n530 VSS 0.00269f
C2657 VDD.n531 VSS 0.00348f
C2658 VDD.n532 VSS 0.00411f
C2659 VDD.n533 VSS 0.00374f
C2660 VDD.n534 VSS -0.0845f
C2661 VDD.n535 VSS 3.26e-19
C2662 VDD.n536 VSS 0.00332f
C2663 VDD.n537 VSS 0.00916f
C2664 VDD.n538 VSS 0.00979f
C2665 VDD.n539 VSS 0.00277f
C2666 VDD.n540 VSS 0.00269f
C2667 VDD.n541 VSS 0.00269f
C2668 VDD.n542 VSS 0.00916f
C2669 VDD.n543 VSS 4.74e-19
C2670 VDD.n544 VSS 0.00979f
C2671 VDD.n545 VSS 0.00332f
C2672 VDD.n546 VSS 0.00411f
C2673 VDD.n547 VSS 0.00374f
C2674 VDD.n548 VSS 0.0141f
C2675 VDD.n549 VSS -0.211f
C2676 VDD.n550 VSS 0.0136f
C2677 VDD.n551 VSS 0.00348f
C2678 VDD.n552 VSS 0.00269f
C2679 VDD.n553 VSS 0.00269f
C2680 VDD.n555 VSS 0.00269f
C2681 VDD.n556 VSS 0.00916f
C2682 VDD.n557 VSS 0.00332f
C2683 VDD.n558 VSS 3.26e-19
C2684 VDD.n559 VSS 0.00374f
C2685 VDD.n560 VSS 0.0223f
C2686 VDD.n561 VSS 0.00374f
C2687 VDD.n562 VSS 0.00348f
C2688 VDD.n563 VSS 0.00269f
C2689 VDD.n564 VSS 0.00269f
C2690 VDD.n565 VSS 0.0389f
C2691 VDD.n566 VSS 0.00332f
C2692 VDD.n567 VSS 3.26e-19
C2693 VDD.n568 VSS 0.161f
C2694 VDD.n569 VSS 0.0109f
C2695 VDD.n570 VSS 0.0161f
C2696 VDD.n571 VSS 0.0109f
C2697 VDD.n572 VSS 0.00634f
C2698 VDD.t60 VSS 0.253f
C2699 VDD.t1 VSS 1.66f
C2700 VDD.n573 VSS 0.471f
C2701 VDD.n574 VSS 0.0161f
C2702 VDD.n575 VSS 0.0161f
C2703 VDD.n576 VSS 0.0109f
C2704 VDD.n577 VSS 0.02f
C2705 VDD.n578 VSS 0.00634f
C2706 VDD.n579 VSS 0.0777f
C2707 VDD.n580 VSS 0.067f
C2708 VDD.n581 VSS 0.00824f
C2709 VDD.n582 VSS 0.02f
C2710 VDD.n583 VSS 0.02f
C2711 VDD.n584 VSS 0.0109f
C2712 VDD.n585 VSS 0.00634f
C2713 VDD.n586 VSS 0.00818f
C2714 VDD.n587 VSS 0.0813f
C2715 VDD.n588 VSS 2.02f
C2716 VDD.t71 VSS 2.26f
C2717 VDD.n589 VSS 0.0193f
C2718 VDD.n590 VSS 0.0171f
C2719 VDD.n591 VSS 0.00786f
C2720 VDD.n592 VSS 0.0168f
C2721 VDD.n593 VSS 0.00663f
C2722 VDD.t15 VSS 0.00663f
C2723 VDD.t13 VSS 0.00663f
C2724 VDD.n594 VSS 0.0163f
C2725 VDD.n595 VSS 0.0482f
C2726 VDD.n596 VSS 0.00805f
C2727 VDD.n597 VSS 0.0164f
C2728 VDD.n598 VSS 0.1f
C2729 VDD.n599 VSS 0.267f
C2730 VDD.n600 VSS 8.15e-19
C2731 VDD.n601 VSS 0.0409f
C2732 VDD.n602 VSS 0.0214f
C2733 VDD.t51 VSS 0.0509f
C2734 VDD.n603 VSS 0.00989f
C2735 VDD.n604 VSS 0.0124f
C2736 VDD.n605 VSS 0.131f
C2737 VDD.n606 VSS 0.014f
C2738 VDD.n607 VSS 0.00256f
C2739 VDD.n608 VSS 0.00391f
C2740 VDD.n609 VSS 0.00873f
C2741 VDD.n610 VSS 0.00443f
C2742 VDD.n611 VSS 0.00672f
C2743 VDD.n612 VSS 0.00689f
C2744 VDD.n613 VSS 0.0606f
C2745 VDD.n614 VSS 0.02f
C2746 VDD.n615 VSS 0.0383f
C2747 VDD.n616 VSS 0.02f
C2748 VDD.n617 VSS 0.0109f
C2749 VDD.n618 VSS 0.00634f
C2750 VDD.n619 VSS 0.199f
C2751 VDD.n620 VSS 0.108f
C2752 VDD.n621 VSS 0.02f
C2753 VDD.n622 VSS 0.00824f
C2754 VDD.n623 VSS 0.0813f
C2755 VDD.n624 VSS 0.00818f
C2756 VDD.n625 VSS 0.00634f
C2757 VDD.n626 VSS 0.0109f
C2758 VDD.n627 VSS 0.0523f
C2759 VDD.n628 VSS 0.02f
C2760 VDD.n629 VSS 0.00634f
C2761 VDD.t47 VSS 0.0509f
C2762 VDD.n630 VSS 0.0561f
C2763 VDD.n631 VSS 0.0109f
C2764 VDD.n632 VSS 0.0274f
C2765 VDD.n633 VSS 0.0261f
C2766 VDD.n634 VSS 0.0277f
C2767 VDD.n635 VSS 0.0111f
C2768 VDD.n636 VSS 0.0122f
C2769 VDD.n637 VSS 0.0158f
C2770 VDD.n638 VSS 0.307f
C2771 VDD.n639 VSS 0.00302f
C2772 VDD.n640 VSS 0.00277f
C2773 VDD.n641 VSS 2.57f
C2774 VDD.n642 VSS 0.0129f
C2775 VDD.n644 VSS 0.0129f
C2776 VDD.n648 VSS 0.0129f
C2777 VDD.n651 VSS 0.00277f
C2778 VDD.n652 VSS 0.0576f
C2779 VDD.n653 VSS 0.00979f
C2780 VDD.n654 VSS 0.00269f
C2781 VDD.n655 VSS 0.00277f
C2782 VDD.n656 VSS 0.00269f
C2783 VDD.n657 VSS 0.00269f
C2784 VDD.n658 VSS 4.74e-19
C2785 VDD.n659 VSS 0.00663f
C2786 VDD.n660 VSS 0.00332f
C2787 VDD.n661 VSS 0.00806f
C2788 VDD.n662 VSS 0.00439f
C2789 VDD.n663 VSS 0.00781f
C2790 VDD.n664 VSS 0.0226f
C2791 VDD.n665 VSS -0.211f
C2792 VDD.n666 VSS 0.0139f
C2793 VDD.n667 VSS 3.26e-19
C2794 VDD.n668 VSS 0.0141f
C2795 VDD.n669 VSS 0.00439f
C2796 VDD.n670 VSS 0.00332f
C2797 VDD.n671 VSS 0.00269f
C2798 VDD.n672 VSS 4.74e-19
C2799 VDD.n673 VSS 0.00269f
C2800 VDD.n674 VSS 0.00979f
C2801 VDD.n675 VSS 0.0104f
C2802 VDD.n676 VSS 0.00269f
C2803 VDD.n677 VSS 0.00269f
C2804 VDD.n678 VSS 4.74e-19
C2805 VDD.n679 VSS 0.00979f
C2806 VDD.n680 VSS 0.00332f
C2807 VDD.n681 VSS 0.00663f
C2808 VDD.n682 VSS 0.00332f
C2809 VDD.n683 VSS 0.00348f
C2810 VDD.n684 VSS 0.00806f
C2811 VDD.n685 VSS 0.00439f
C2812 VDD.n686 VSS 0.00781f
C2813 VDD.n687 VSS 0.0223f
C2814 VDD.n688 VSS -0.211f
C2815 VDD.n689 VSS 0.0136f
C2816 VDD.n690 VSS 3.26e-19
C2817 VDD.n691 VSS 4.74e-19
C2818 VDD.n692 VSS 0.00585f
C2819 VDD.n693 VSS 0.00348f
C2820 VDD.n694 VSS 0.00269f
C2821 VDD.n695 VSS 0.0129f
C2822 VDD.n696 VSS 0.00979f
C2823 VDD.n697 VSS 0.00332f
C2824 VDD.n698 VSS 0.00585f
C2825 VDD.n699 VSS 0.00348f
C2826 VDD.n700 VSS 4.74e-19
C2827 VDD.n701 VSS 3.26e-19
C2828 VDD.n702 VSS 0.00488f
C2829 VDD.n703 VSS 0.0227f
C2830 VDD.n704 VSS 0.00439f
C2831 VDD.n705 VSS 0.00411f
C2832 VDD.n706 VSS 0.00348f
C2833 VDD.n707 VSS 0.00916f
C2834 VDD.n708 VSS 0.00269f
C2835 VDD.n709 VSS 0.00979f
C2836 VDD.n710 VSS 0.00979f
C2837 VDD.n711 VSS 0.00269f
C2838 VDD.n713 VSS 0.00277f
C2839 VDD.n714 VSS 0.00269f
C2840 VDD.n715 VSS 0.0129f
C2841 VDD.n716 VSS 0.00269f
C2842 VDD.n717 VSS 0.00269f
C2843 VDD.n718 VSS 0.00348f
C2844 VDD.n719 VSS 0.00781f
C2845 VDD.n720 VSS 0.0141f
C2846 VDD.n721 VSS -0.0753f
C2847 VDD.n722 VSS 0.00411f
C2848 VDD.n723 VSS 0.00916f
C2849 VDD.n724 VSS 0.00269f
C2850 VDD.n725 VSS 0.00269f
C2851 VDD.n726 VSS 0.00348f
C2852 VDD.n727 VSS 0.0285f
C2853 VDD.n728 VSS 0.0141f
C2854 VDD.n729 VSS 3.26e-19
C2855 VDD.n730 VSS 0.00332f
C2856 VDD.n731 VSS 0.00348f
C2857 VDD.n732 VSS 0.00916f
C2858 VDD.n733 VSS 0.00269f
C2859 VDD.n734 VSS 0.00269f
C2860 VDD.n735 VSS 0.0294f
C2861 VDD.n736 VSS 0.00332f
C2862 VDD.n737 VSS 0.0261f
C2863 VDD.n738 VSS 0.0286f
C2864 VDD.n739 VSS 0.0286f
C2865 VDD.n740 VSS 0.0261f
C2866 VDD.n741 VSS 0.00332f
C2867 VDD.n742 VSS 0.0294f
C2868 VDD.n743 VSS 0.00269f
C2869 VDD.n744 VSS 0.0104f
C2870 VDD.n745 VSS 0.00269f
C2871 VDD.n746 VSS 0.00269f
C2872 VDD.n747 VSS 0.00348f
C2873 VDD.n748 VSS 0.00411f
C2874 VDD.n749 VSS 0.00374f
C2875 VDD.n750 VSS 0.0141f
C2876 VDD.n751 VSS 3.26e-19
C2877 VDD.n752 VSS 0.00332f
C2878 VDD.n753 VSS 0.00916f
C2879 VDD.n754 VSS 0.00979f
C2880 VDD.n755 VSS 0.00277f
C2881 VDD.n756 VSS 0.00269f
C2882 VDD.n757 VSS 0.00269f
C2883 VDD.n758 VSS 0.00916f
C2884 VDD.n759 VSS 4.74e-19
C2885 VDD.n760 VSS 0.00979f
C2886 VDD.n761 VSS 0.00332f
C2887 VDD.n762 VSS 0.00411f
C2888 VDD.n763 VSS 0.00374f
C2889 VDD.n764 VSS -0.0845f
C2890 VDD.n765 VSS 0.00472f
C2891 VDD.n766 VSS 0.0136f
C2892 VDD.n767 VSS 0.00348f
C2893 VDD.n768 VSS 0.00269f
C2894 VDD.n769 VSS 0.00269f
C2895 VDD.n770 VSS 3.16e-19
C2896 VDD.n771 VSS 0.0129f
C2897 VDD.n772 VSS 0.00269f
C2898 VDD.n773 VSS 0.00269f
C2899 VDD.n774 VSS 0.00916f
C2900 VDD.n775 VSS 0.00348f
C2901 VDD.n776 VSS 0.00411f
C2902 VDD.n777 VSS 0.00374f
C2903 VDD.n778 VSS 3.26e-19
C2904 VDD.n779 VSS 0.0141f
C2905 VDD.n780 VSS 3.26e-19
C2906 VDD.n781 VSS 0.00332f
C2907 VDD.n782 VSS 0.00916f
C2908 VDD.n783 VSS 0.00269f
C2909 VDD.n784 VSS 0.0104f
C2910 VDD.n785 VSS 0.00269f
C2911 VDD.n786 VSS 0.00269f
C2912 VDD.n787 VSS 0.00348f
C2913 VDD.n788 VSS 0.00411f
C2914 VDD.n789 VSS 0.00374f
C2915 VDD.n790 VSS -0.0845f
C2916 VDD.n791 VSS 3.26e-19
C2917 VDD.n792 VSS 0.00332f
C2918 VDD.n793 VSS 0.0295f
C2919 VDD.n794 VSS 0.00269f
C2920 VDD.n795 VSS 0.0129f
C2921 VDD.n796 VSS 0.00269f
C2922 VDD.n797 VSS 0.00269f
C2923 VDD.n798 VSS 4.74e-19
C2924 VDD.n799 VSS 0.00332f
C2925 VDD.n800 VSS 0.00411f
C2926 VDD.n801 VSS 0.0251f
C2927 VDD.n802 VSS 0.00439f
C2928 VDD.n803 VSS 0.0241f
C2929 VDD.n804 VSS -0.182f
C2930 VDD.n805 VSS 0.00488f
C2931 VDD.n806 VSS 0.0136f
C2932 VDD.n807 VSS 3.26e-19
C2933 VDD.n808 VSS 4.74e-19
C2934 VDD.n809 VSS 0.00585f
C2935 VDD.n810 VSS 0.00348f
C2936 VDD.n811 VSS 3.16e-19
C2937 VDD.n812 VSS 0.00277f
C2938 VDD.n813 VSS 0.00269f
C2939 VDD.n814 VSS 0.00269f
C2940 VDD.n815 VSS 0.00663f
C2941 VDD.n816 VSS 0.00411f
C2942 VDD.n817 VSS -0.0753f
C2943 VDD.n818 VSS 0.00472f
C2944 VDD.n819 VSS 0.00781f
C2945 VDD.n820 VSS 0.0223f
C2946 VDD.n821 VSS 0.00781f
C2947 VDD.n822 VSS 0.00348f
C2948 VDD.n823 VSS 0.00332f
C2949 VDD.n824 VSS 0.00269f
C2950 VDD.n825 VSS 0.00916f
C2951 VDD.n826 VSS 0.00269f
C2952 VDD.n827 VSS 0.00979f
C2953 VDD.n828 VSS 0.0104f
C2954 VDD.n829 VSS 0.00269f
C2955 VDD.n830 VSS 0.00269f
C2956 VDD.n831 VSS 4.74e-19
C2957 VDD.n832 VSS 0.00979f
C2958 VDD.n833 VSS 0.00332f
C2959 VDD.n834 VSS 0.00663f
C2960 VDD.n835 VSS 0.00332f
C2961 VDD.n836 VSS 0.00806f
C2962 VDD.n837 VSS 0.00439f
C2963 VDD.n838 VSS -0.182f
C2964 VDD.n839 VSS 0.00488f
C2965 VDD.n840 VSS 0.0136f
C2966 VDD.n841 VSS 3.26e-19
C2967 VDD.n842 VSS 4.74e-19
C2968 VDD.n843 VSS 0.00585f
C2969 VDD.n844 VSS 0.00348f
C2970 VDD.n845 VSS 0.00269f
C2971 VDD.n846 VSS 0.0129f
C2972 VDD.n847 VSS 0.00979f
C2973 VDD.n848 VSS 0.00332f
C2974 VDD.n849 VSS 0.00585f
C2975 VDD.n850 VSS 0.00348f
C2976 VDD.n851 VSS 4.74e-19
C2977 VDD.n852 VSS 3.26e-19
C2978 VDD.n853 VSS -0.211f
C2979 VDD.n854 VSS 0.0805f
C2980 VDD.n855 VSS 3.26e-19
C2981 VDD.n856 VSS 0.00332f
C2982 VDD.n857 VSS 0.00348f
C2983 VDD.n858 VSS 0.00916f
C2984 VDD.n859 VSS 0.00269f
C2985 VDD.n860 VSS 0.00269f
C2986 VDD.n861 VSS 0.0294f
C2987 VDD.n862 VSS 0.0261f
C2988 VDD.n863 VSS 0.00332f
C2989 VDD.n864 VSS 0.00979f
C2990 VDD.n865 VSS 0.00269f
C2991 VDD.n867 VSS 0.00277f
C2992 VDD.n868 VSS 0.0236f
C2993 VDD.n869 VSS 3.16e-19
C2994 VDD.n870 VSS 0.00269f
C2995 VDD.n871 VSS 0.00269f
C2996 VDD.n872 VSS 0.00348f
C2997 VDD.n873 VSS 0.0286f
C2998 VDD.n874 VSS 0.0286f
C2999 VDD.n875 VSS 0.0261f
C3000 VDD.n876 VSS 0.00332f
C3001 VDD.n877 VSS 0.0294f
C3002 VDD.n878 VSS 0.00269f
C3003 VDD.n879 VSS 0.0104f
C3004 VDD.n880 VSS 0.00269f
C3005 VDD.n881 VSS 0.00269f
C3006 VDD.n882 VSS 0.00348f
C3007 VDD.n883 VSS 0.00411f
C3008 VDD.n884 VSS 0.00374f
C3009 VDD.n885 VSS 0.0141f
C3010 VDD.n886 VSS 3.26e-19
C3011 VDD.n887 VSS 0.00332f
C3012 VDD.n888 VSS 0.00916f
C3013 VDD.n889 VSS 0.00979f
C3014 VDD.n890 VSS 0.00277f
C3015 VDD.n891 VSS 0.00269f
C3016 VDD.n892 VSS 0.00269f
C3017 VDD.n893 VSS 0.00916f
C3018 VDD.n894 VSS 4.74e-19
C3019 VDD.n895 VSS 0.00979f
C3020 VDD.n896 VSS 0.00332f
C3021 VDD.n897 VSS 0.00411f
C3022 VDD.n898 VSS 0.00374f
C3023 VDD.n899 VSS -0.0845f
C3024 VDD.n900 VSS 0.00472f
C3025 VDD.n901 VSS 0.0136f
C3026 VDD.n902 VSS 0.00348f
C3027 VDD.n903 VSS 0.00269f
C3028 VDD.n904 VSS 0.00269f
C3029 VDD.n905 VSS 3.16e-19
C3030 VDD.n906 VSS 0.0129f
C3031 VDD.n907 VSS 0.00269f
C3032 VDD.n908 VSS 0.00269f
C3033 VDD.n909 VSS 0.00916f
C3034 VDD.n910 VSS 0.00348f
C3035 VDD.n911 VSS 0.00411f
C3036 VDD.n912 VSS 0.00374f
C3037 VDD.n913 VSS 3.26e-19
C3038 VDD.n914 VSS 0.0141f
C3039 VDD.n915 VSS 3.26e-19
C3040 VDD.n916 VSS 0.00332f
C3041 VDD.n917 VSS 0.00916f
C3042 VDD.n918 VSS 0.00269f
C3043 VDD.n919 VSS 0.0104f
C3044 VDD.n920 VSS 0.00269f
C3045 VDD.n921 VSS 0.00269f
C3046 VDD.n922 VSS 0.00348f
C3047 VDD.n923 VSS 0.00411f
C3048 VDD.n924 VSS 0.00374f
C3049 VDD.n925 VSS -0.0845f
C3050 VDD.n926 VSS 3.26e-19
C3051 VDD.n927 VSS 0.00332f
C3052 VDD.n928 VSS 0.0295f
C3053 VDD.n929 VSS 0.00269f
C3054 VDD.n930 VSS 0.0129f
C3055 VDD.n931 VSS 0.00269f
C3056 VDD.n932 VSS 0.00269f
C3057 VDD.n933 VSS 4.74e-19
C3058 VDD.n934 VSS 0.00332f
C3059 VDD.n935 VSS 0.00411f
C3060 VDD.n936 VSS 0.0251f
C3061 VDD.n937 VSS 0.00439f
C3062 VDD.n938 VSS 0.0241f
C3063 VDD.n939 VSS -0.182f
C3064 VDD.n940 VSS 0.00488f
C3065 VDD.n941 VSS 0.0136f
C3066 VDD.n942 VSS 3.26e-19
C3067 VDD.n943 VSS 4.74e-19
C3068 VDD.n944 VSS 0.00585f
C3069 VDD.n945 VSS 0.00348f
C3070 VDD.n946 VSS 3.16e-19
C3071 VDD.n947 VSS 0.00277f
C3072 VDD.n948 VSS 0.00269f
C3073 VDD.n949 VSS 0.00269f
C3074 VDD.n950 VSS 0.00663f
C3075 VDD.n951 VSS 0.00411f
C3076 VDD.n952 VSS -0.0753f
C3077 VDD.n953 VSS 0.00472f
C3078 VDD.n954 VSS 0.00781f
C3079 VDD.n955 VSS 0.0223f
C3080 VDD.n956 VSS 0.00781f
C3081 VDD.n957 VSS 0.00348f
C3082 VDD.n958 VSS 0.00332f
C3083 VDD.n959 VSS 0.00269f
C3084 VDD.n960 VSS 0.00916f
C3085 VDD.n961 VSS 0.00269f
C3086 VDD.n962 VSS 0.00979f
C3087 VDD.n963 VSS 0.0104f
C3088 VDD.n964 VSS 0.00269f
C3089 VDD.n965 VSS 0.00269f
C3090 VDD.n966 VSS 4.74e-19
C3091 VDD.n967 VSS 0.00979f
C3092 VDD.n968 VSS 0.00332f
C3093 VDD.n969 VSS 0.00663f
C3094 VDD.n970 VSS 0.00332f
C3095 VDD.n971 VSS 0.00806f
C3096 VDD.n972 VSS 0.00439f
C3097 VDD.n973 VSS -0.182f
C3098 VDD.n974 VSS 0.00488f
C3099 VDD.n975 VSS 0.0136f
C3100 VDD.n976 VSS 3.26e-19
C3101 VDD.n977 VSS 4.74e-19
C3102 VDD.n978 VSS 0.00585f
C3103 VDD.n979 VSS 0.00348f
C3104 VDD.n980 VSS 0.00269f
C3105 VDD.n981 VSS 0.0129f
C3106 VDD.n982 VSS 0.00979f
C3107 VDD.n983 VSS 0.00332f
C3108 VDD.n984 VSS 0.00585f
C3109 VDD.n985 VSS 0.00348f
C3110 VDD.n986 VSS 4.74e-19
C3111 VDD.n987 VSS 3.26e-19
C3112 VDD.n988 VSS -0.211f
C3113 VDD.n989 VSS 0.0805f
C3114 VDD.n990 VSS 3.26e-19
C3115 VDD.n991 VSS 0.00332f
C3116 VDD.n992 VSS 0.00348f
C3117 VDD.n993 VSS 0.00916f
C3118 VDD.n994 VSS 0.00269f
C3119 VDD.n995 VSS 0.00269f
C3120 VDD.n996 VSS 0.0294f
C3121 VDD.n997 VSS 0.0261f
C3122 VDD.n998 VSS 0.00332f
C3123 VDD.n999 VSS 0.00979f
C3124 VDD.n1000 VSS 0.00269f
C3125 VDD.n1002 VSS 0.00277f
C3126 VDD.n1003 VSS 0.0236f
C3127 VDD.n1004 VSS 3.16e-19
C3128 VDD.n1005 VSS 0.00269f
C3129 VDD.n1006 VSS 0.00269f
C3130 VDD.n1007 VSS 0.00348f
C3131 VDD.n1008 VSS 0.0286f
C3132 VDD.n1009 VSS 0.0286f
C3133 VDD.n1010 VSS 0.0261f
C3134 VDD.n1011 VSS 0.00332f
C3135 VDD.n1012 VSS 0.0294f
C3136 VDD.n1013 VSS 0.00269f
C3137 VDD.n1014 VSS 0.0104f
C3138 VDD.n1015 VSS 0.00269f
C3139 VDD.n1016 VSS 0.00269f
C3140 VDD.n1017 VSS 0.00348f
C3141 VDD.n1018 VSS 0.00411f
C3142 VDD.n1019 VSS 0.00374f
C3143 VDD.n1020 VSS 0.0141f
C3144 VDD.n1021 VSS 3.26e-19
C3145 VDD.n1022 VSS 0.00332f
C3146 VDD.n1023 VSS 0.00916f
C3147 VDD.n1024 VSS 0.00979f
C3148 VDD.n1025 VSS 0.00277f
C3149 VDD.n1026 VSS 0.00269f
C3150 VDD.n1027 VSS 0.00269f
C3151 VDD.n1028 VSS 0.00916f
C3152 VDD.n1029 VSS 4.74e-19
C3153 VDD.n1030 VSS 0.00979f
C3154 VDD.n1031 VSS 0.00332f
C3155 VDD.n1032 VSS 0.00411f
C3156 VDD.n1033 VSS 0.00374f
C3157 VDD.n1034 VSS -0.0845f
C3158 VDD.n1035 VSS 0.00472f
C3159 VDD.n1036 VSS 0.0136f
C3160 VDD.n1037 VSS 0.00348f
C3161 VDD.n1038 VSS 0.00269f
C3162 VDD.n1039 VSS 0.00269f
C3163 VDD.n1040 VSS 3.16e-19
C3164 VDD.n1041 VSS 0.0129f
C3165 VDD.n1042 VSS 0.00269f
C3166 VDD.n1043 VSS 0.00269f
C3167 VDD.n1044 VSS 0.00916f
C3168 VDD.n1045 VSS 0.00348f
C3169 VDD.n1046 VSS 0.00411f
C3170 VDD.n1047 VSS 0.00374f
C3171 VDD.n1048 VSS 3.26e-19
C3172 VDD.n1049 VSS 0.0141f
C3173 VDD.n1050 VSS 3.26e-19
C3174 VDD.n1051 VSS 0.00332f
C3175 VDD.n1052 VSS 0.00916f
C3176 VDD.n1053 VSS 0.00269f
C3177 VDD.n1054 VSS 0.0104f
C3178 VDD.n1055 VSS 0.00269f
C3179 VDD.n1056 VSS 0.00269f
C3180 VDD.n1057 VSS 0.00348f
C3181 VDD.n1058 VSS 0.00411f
C3182 VDD.n1059 VSS 0.00374f
C3183 VDD.n1060 VSS -0.0845f
C3184 VDD.n1061 VSS 3.26e-19
C3185 VDD.n1062 VSS 0.00332f
C3186 VDD.n1063 VSS 0.0295f
C3187 VDD.n1064 VSS 0.00269f
C3188 VDD.n1065 VSS 0.0129f
C3189 VDD.n1066 VSS 0.00269f
C3190 VDD.n1067 VSS 0.00269f
C3191 VDD.n1068 VSS 4.74e-19
C3192 VDD.n1069 VSS 0.00332f
C3193 VDD.n1070 VSS 0.00411f
C3194 VDD.n1071 VSS 0.0251f
C3195 VDD.n1072 VSS 0.00439f
C3196 VDD.n1073 VSS 0.0241f
C3197 VDD.n1074 VSS -0.182f
C3198 VDD.n1075 VSS 0.00488f
C3199 VDD.n1076 VSS 0.0136f
C3200 VDD.n1077 VSS 3.26e-19
C3201 VDD.n1078 VSS 4.74e-19
C3202 VDD.n1079 VSS 0.00585f
C3203 VDD.n1080 VSS 0.00348f
C3204 VDD.n1081 VSS 3.16e-19
C3205 VDD.n1082 VSS 0.00277f
C3206 VDD.n1083 VSS 0.00269f
C3207 VDD.n1084 VSS 0.00269f
C3208 VDD.n1085 VSS 0.00663f
C3209 VDD.n1086 VSS 0.00411f
C3210 VDD.n1087 VSS -0.0753f
C3211 VDD.n1088 VSS 0.00472f
C3212 VDD.n1089 VSS 0.00781f
C3213 VDD.n1090 VSS 0.0223f
C3214 VDD.n1091 VSS 0.00781f
C3215 VDD.n1092 VSS 0.00348f
C3216 VDD.n1093 VSS 0.00332f
C3217 VDD.n1094 VSS 0.00269f
C3218 VDD.n1095 VSS 0.00916f
C3219 VDD.n1096 VSS 0.00269f
C3220 VDD.n1097 VSS 0.00979f
C3221 VDD.n1098 VSS 0.0104f
C3222 VDD.n1099 VSS 0.00269f
C3223 VDD.n1100 VSS 0.00269f
C3224 VDD.n1101 VSS 4.74e-19
C3225 VDD.n1102 VSS 0.00979f
C3226 VDD.n1103 VSS 0.00332f
C3227 VDD.n1104 VSS 0.00663f
C3228 VDD.n1105 VSS 0.00332f
C3229 VDD.n1106 VSS 0.00806f
C3230 VDD.n1107 VSS 0.00439f
C3231 VDD.n1108 VSS -0.182f
C3232 VDD.n1109 VSS 0.00488f
C3233 VDD.n1110 VSS 0.0136f
C3234 VDD.n1111 VSS 3.26e-19
C3235 VDD.n1112 VSS 4.74e-19
C3236 VDD.n1113 VSS 0.00585f
C3237 VDD.n1114 VSS 0.00348f
C3238 VDD.n1115 VSS 0.00269f
C3239 VDD.n1116 VSS 0.0129f
C3240 VDD.n1117 VSS 0.00979f
C3241 VDD.n1118 VSS 0.00332f
C3242 VDD.n1119 VSS 0.00585f
C3243 VDD.n1120 VSS 0.00348f
C3244 VDD.n1121 VSS 4.74e-19
C3245 VDD.n1122 VSS 3.26e-19
C3246 VDD.n1123 VSS -0.211f
C3247 VDD.n1124 VSS 0.0805f
C3248 VDD.n1125 VSS 3.26e-19
C3249 VDD.n1126 VSS 0.00332f
C3250 VDD.n1127 VSS 0.00348f
C3251 VDD.n1128 VSS 0.00916f
C3252 VDD.n1129 VSS 0.00269f
C3253 VDD.n1130 VSS 0.00269f
C3254 VDD.n1131 VSS 0.0294f
C3255 VDD.n1132 VSS 0.0261f
C3256 VDD.n1133 VSS 0.00332f
C3257 VDD.n1134 VSS 0.00979f
C3258 VDD.n1135 VSS 0.00269f
C3259 VDD.n1137 VSS 0.00277f
C3260 VDD.n1138 VSS 0.0236f
C3261 VDD.n1139 VSS 3.16e-19
C3262 VDD.n1140 VSS 0.00269f
C3263 VDD.n1141 VSS 0.00269f
C3264 VDD.n1142 VSS 0.00348f
C3265 VDD.n1143 VSS 0.0286f
C3266 VDD.n1144 VSS 0.0286f
C3267 VDD.n1145 VSS 0.0261f
C3268 VDD.n1146 VSS 0.00332f
C3269 VDD.n1147 VSS 0.0294f
C3270 VDD.n1148 VSS 0.00269f
C3271 VDD.n1149 VSS 0.0104f
C3272 VDD.n1150 VSS 0.00269f
C3273 VDD.n1151 VSS 0.00269f
C3274 VDD.n1152 VSS 0.00348f
C3275 VDD.n1153 VSS 0.00411f
C3276 VDD.n1154 VSS 0.00374f
C3277 VDD.n1155 VSS 0.0141f
C3278 VDD.n1156 VSS 3.26e-19
C3279 VDD.n1157 VSS 0.00332f
C3280 VDD.n1158 VSS 0.00916f
C3281 VDD.n1159 VSS 0.00979f
C3282 VDD.n1160 VSS 0.00277f
C3283 VDD.n1161 VSS 0.00269f
C3284 VDD.n1162 VSS 0.00269f
C3285 VDD.n1163 VSS 0.00916f
C3286 VDD.n1164 VSS 4.74e-19
C3287 VDD.n1165 VSS 0.00979f
C3288 VDD.n1166 VSS 0.00332f
C3289 VDD.n1167 VSS 0.00411f
C3290 VDD.n1168 VSS 0.00374f
C3291 VDD.n1169 VSS -0.0845f
C3292 VDD.n1170 VSS 0.00472f
C3293 VDD.n1171 VSS 0.0136f
C3294 VDD.n1172 VSS 0.00348f
C3295 VDD.n1173 VSS 0.00269f
C3296 VDD.n1174 VSS 0.00269f
C3297 VDD.n1175 VSS 3.16e-19
C3298 VDD.n1176 VSS 0.0129f
C3299 VDD.n1177 VSS 0.00269f
C3300 VDD.n1178 VSS 0.00269f
C3301 VDD.n1179 VSS 0.00916f
C3302 VDD.n1180 VSS 0.00348f
C3303 VDD.n1181 VSS 0.00411f
C3304 VDD.n1182 VSS 0.00374f
C3305 VDD.n1183 VSS 3.26e-19
C3306 VDD.n1184 VSS 0.0141f
C3307 VDD.n1185 VSS 3.26e-19
C3308 VDD.n1186 VSS 0.00332f
C3309 VDD.n1187 VSS 0.00916f
C3310 VDD.n1188 VSS 0.00269f
C3311 VDD.n1189 VSS 0.0276f
C3312 VDD.n1190 VSS 0.00269f
C3313 VDD.n1191 VSS 0.00269f
C3314 VDD.n1192 VSS 0.00348f
C3315 VDD.n1193 VSS 0.00411f
C3316 VDD.n1194 VSS 0.00374f
C3317 VDD.n1195 VSS -0.0845f
C3318 VDD.n1196 VSS 3.26e-19
C3319 VDD.n1197 VSS 0.00332f
C3320 VDD.n1198 VSS 0.161f
C3321 VDD.n1199 VSS 0.0109f
C3322 VDD.n1200 VSS 0.0161f
C3323 VDD.n1201 VSS 0.0109f
C3324 VDD.n1202 VSS 0.00634f
C3325 VDD.t11 VSS 0.253f
C3326 VDD.t8 VSS 1.66f
C3327 VDD.n1203 VSS 0.471f
C3328 VDD.n1204 VSS 0.0161f
C3329 VDD.n1205 VSS 0.0161f
C3330 VDD.n1206 VSS 0.0109f
C3331 VDD.n1207 VSS 0.02f
C3332 VDD.n1208 VSS 0.00634f
C3333 VDD.n1209 VSS 0.0777f
C3334 VDD.n1210 VSS 0.067f
C3335 VDD.n1211 VSS 0.00824f
C3336 VDD.n1212 VSS 0.02f
C3337 VDD.n1213 VSS 0.02f
C3338 VDD.n1214 VSS 0.0109f
C3339 VDD.n1215 VSS 0.00634f
C3340 VDD.n1216 VSS 0.00818f
C3341 VDD.n1217 VSS 0.0813f
C3342 VDD.n1218 VSS 2.02f
C3343 VDD.t16 VSS 2.26f
C3344 VDD.n1219 VSS 0.0193f
C3345 VDD.n1220 VSS 0.0171f
C3346 VDD.n1221 VSS 0.00786f
C3347 VDD.n1222 VSS 0.0168f
C3348 VDD.n1223 VSS 0.00663f
C3349 VDD.t24 VSS 0.00663f
C3350 VDD.t27 VSS 0.00663f
C3351 VDD.n1224 VSS 0.0163f
C3352 VDD.n1225 VSS 0.0482f
C3353 VDD.n1226 VSS 0.00805f
C3354 VDD.n1227 VSS 0.0164f
C3355 VDD.n1228 VSS 0.1f
C3356 VDD.n1229 VSS 0.113f
C3357 VDD.n1230 VSS 0.004f
C3358 VDD.n1231 VSS 0.0124f
C3359 VDD.n1232 VSS 0.016f
C3360 VDD.n1233 VSS 0.0232f
C3361 VDD.n1234 VSS 0.0193f
C3362 VDD.t76 VSS 0.0509f
C3363 VDD.n1235 VSS 0.0556f
C3364 VDD.n1236 VSS 0.00797f
C3365 VDD.n1237 VSS 0.00256f
C3366 VDD.n1238 VSS 0.0203f
C3367 VDD.n1239 VSS 0.00163f
C3368 VDD.n1240 VSS 0.0632f
C3369 VDD.t75 VSS 0.104f
C3370 VDD.t48 VSS 0.124f
C3371 VDD.n1241 VSS 0.0639f
C3372 VDD.n1242 VSS 0.0527f
C3373 VDD.n1243 VSS 0.00277f
C3374 VDD.n1244 VSS 0.00269f
C3375 VDD.n1245 VSS 0.00348f
C3376 VDD.n1246 VSS 0.0129f
C3377 VDD.n1247 VSS 0.198f
C3378 VDD.n1248 VSS 0.0104f
C3379 VDD.n1249 VSS 0.00979f
C3380 VDD.n1250 VSS 0.00269f
C3381 VDD.n1251 VSS 0.00916f
C3382 VDD.n1252 VSS 4.74e-19
C3383 VDD.n1253 VSS 0.00332f
C3384 VDD.n1254 VSS 0.00585f
C3385 VDD.n1255 VSS 0.00348f
C3386 VDD.n1256 VSS 4.74e-19
C3387 VDD.n1257 VSS -0.211f
C3388 VDD.n1258 VSS 3.26e-19
C3389 VDD.n1259 VSS 0.0233f
C3390 VDD.n1260 VSS 0.00439f
C3391 VDD.n1261 VSS -0.174f
C3392 VDD.n1262 VSS 0.00798f
C3393 VDD.n1263 VSS 0.00332f
C3394 VDD.n1264 VSS 0.00439f
C3395 VDD.n1265 VSS 0.0084f
C3396 VDD.n1266 VSS 0.0122f
C3397 VDD.t25 VSS 0.00583f
C3398 VDD.n1267 VSS 0.0574f
C3399 VDD.n1268 VSS 0.00618f
C3400 VDD.n1269 VSS 0.0303f
C3401 VDD.n1270 VSS 0.028f
C3402 VDD.n1271 VSS 0.0111f
C3403 VDD.n1272 VSS 0.00106f
C3404 VDD.n1273 VSS 0.0174f
C3405 VDD.n1274 VSS 0.0362f
C3406 VDD.n1275 VSS 0.0158f
C3407 VDD.n1276 VSS 0.00411f
C3408 VDD.n1277 VSS 0.00779f
C3409 VDD.n1278 VSS 0.00472f
C3410 VDD.n1279 VSS 0.00759f
C3411 VDD.n1280 VSS 0.0145f
C3412 VDD.n1281 VSS 0.014f
C3413 VDD.n1282 VSS -0.0841f
C3414 VDD.n1283 VSS 3.26e-19
C3415 VDD.n1284 VSS 0.00488f
C3416 VDD.n1285 VSS 4.74e-19
C3417 VDD.n1286 VSS 0.00348f
C3418 VDD.n1287 VSS 0.00269f
C3419 VDD.n1288 VSS 0.00979f
C3420 VDD.n1289 VSS 0.00332f
C3421 VDD.n1290 VSS 0.00663f
C3422 VDD.n1291 VSS 0.00806f
C3423 VDD.n1292 VSS 0.00332f
C3424 VDD.n1293 VSS 0.00411f
C3425 VDD.n1294 VSS 0.00585f
C3426 VDD.n1295 VSS 0.00472f
C3427 VDD.n1296 VSS 0.00374f
C3428 VDD.n1297 VSS 0.0229f
C3429 VDD.n1298 VSS 0.014f
C3430 VDD.n1299 VSS 0.0145f
C3431 VDD.n1300 VSS 3.26e-19
C3432 VDD.n1301 VSS 0.00488f
C3433 VDD.n1302 VSS 0.00798f
C3434 VDD.n1303 VSS 0.00374f
C3435 VDD.n1304 VSS 0.0229f
C3436 VDD.n1305 VSS 0.0229f
C3437 VDD.n1306 VSS 0.00488f
C3438 VDD.n1307 VSS 0.00439f
C3439 VDD.n1308 VSS 0.00806f
C3440 VDD.n1309 VSS 0.00332f
C3441 VDD.n1310 VSS 0.00663f
C3442 VDD.n1311 VSS 4.74e-19
C3443 VDD.n1312 VSS 0.00269f
C3444 VDD.n1313 VSS 0.00269f
C3445 VDD.n1314 VSS 0.00269f
C3446 VDD.n1315 VSS 0.00277f
C3447 VDD.n1316 VSS 0.0129f
C3448 VDD.n1317 VSS 0.198f
C3449 VDD.n1318 VSS 0.0104f
C3450 VDD.n1319 VSS 0.00979f
C3451 VDD.n1320 VSS 0.00979f
C3452 VDD.n1321 VSS 0.0129f
C3453 VDD.n1322 VSS 0.245f
C3454 VDD.n1323 VSS 0.0527f
C3455 VDD.n1324 VSS 0.00277f
C3456 VDD.n1325 VSS 0.00269f
C3457 VDD.n1326 VSS 3.16e-19
C3458 VDD.n1327 VSS 0.00269f
C3459 VDD.n1328 VSS 0.00348f
C3460 VDD.n1329 VSS 0.00269f
C3461 VDD.n1330 VSS 0.00332f
C3462 VDD.n1331 VSS 0.00979f
C3463 VDD.n1332 VSS 0.00979f
C3464 VDD.n1333 VSS 0.0129f
C3465 VDD.n1334 VSS 0.245f
C3466 VDD.n1335 VSS 0.0527f
C3467 VDD.n1336 VSS 0.198f
C3468 VDD.n1337 VSS 0.0104f
C3469 VDD.n1338 VSS 0.00979f
C3470 VDD.n1339 VSS 0.00269f
C3471 VDD.n1340 VSS 0.00916f
C3472 VDD.n1341 VSS 4.74e-19
C3473 VDD.n1342 VSS 0.00332f
C3474 VDD.n1343 VSS 0.00585f
C3475 VDD.n1344 VSS 0.0576f
C3476 VDD.n1345 VSS 0.0433f
C3477 VDD.n1346 VSS -0.211f
C3478 VDD.n1347 VSS 3.26e-19
C3479 VDD.n1348 VSS 0.0233f
C3480 VDD.n1349 VSS 0.00439f
C3481 VDD.n1350 VSS -0.174f
C3482 VDD.n1351 VSS 0.014f
C3483 VDD.n1352 VSS -0.0841f
C3484 VDD.n1353 VSS 3.26e-19
C3485 VDD.n1354 VSS 0.00488f
C3486 VDD.n1355 VSS 0.00798f
C3487 VDD.n1356 VSS 0.00348f
C3488 VDD.n1357 VSS 0.00979f
C3489 VDD.n1358 VSS 0.00332f
C3490 VDD.n1359 VSS 0.00663f
C3491 VDD.n1360 VSS 0.00806f
C3492 VDD.n1361 VSS 0.00332f
C3493 VDD.n1362 VSS 0.00411f
C3494 VDD.n1363 VSS 0.00585f
C3495 VDD.n1364 VSS 0.00472f
C3496 VDD.n1365 VSS 0.00374f
C3497 VDD.n1366 VSS 0.0229f
C3498 VDD.n1367 VSS 0.014f
C3499 VDD.n1368 VSS 0.0145f
C3500 VDD.n1369 VSS 3.26e-19
C3501 VDD.n1370 VSS 0.00488f
C3502 VDD.n1371 VSS 0.00798f
C3503 VDD.n1372 VSS 0.00374f
C3504 VDD.n1373 VSS 0.0229f
C3505 VDD.n1374 VSS 0.0138f
C3506 VDD.n1375 VSS 0.00439f
C3507 VDD.n1376 VSS 0.00332f
C3508 VDD.n1377 VSS 4.74e-19
C3509 VDD.n1378 VSS 0.00269f
C3510 VDD.n1379 VSS 0.018f
C3511 VDD.n1380 VSS 0.00269f
C3512 VDD.n1381 VSS 0.00277f
C3513 VDD.n1382 VSS 0.0129f
C3514 VDD.n1383 VSS 0.0527f
C3515 VDD.n1384 VSS 0.00277f
C3516 VDD.n1385 VSS 0.00979f
C3517 VDD.n1386 VSS 0.245f
C3518 VDD.n1387 VSS 0.0129f
C3519 VDD.n1388 VSS 0.00979f
C3520 VDD.n1389 VSS 0.00269f
C3521 VDD.n1390 VSS 0.0314f
C3522 VDD.n1391 VSS 0.0236f
C3523 VDD.n1392 VSS 0.124f
C3524 VDD.t31 VSS 0.49f
C3525 VDD.n1393 VSS 0.605f
C3526 VDD.n1394 VSS 0.0527f
C3527 VDD.n1395 VSS 0.198f
C3528 VDD.n1396 VSS 0.0104f
C3529 VDD.n1397 VSS 0.00979f
C3530 VDD.n1398 VSS 0.00269f
C3531 VDD.n1399 VSS 0.00916f
C3532 VDD.n1400 VSS 4.74e-19
C3533 VDD.n1401 VSS 0.00332f
C3534 VDD.n1402 VSS 0.00585f
C3535 VDD.n1403 VSS 0.00348f
C3536 VDD.n1404 VSS 4.74e-19
C3537 VDD.n1405 VSS -0.211f
C3538 VDD.n1406 VSS 3.26e-19
C3539 VDD.n1407 VSS 0.023f
C3540 VDD.n1408 VSS 0.00439f
C3541 VDD.n1409 VSS -0.174f
C3542 VDD.n1410 VSS -0.0844f
C3543 VDD.n1411 VSS 3.26e-19
C3544 VDD.n1412 VSS 0.00488f
C3545 VDD.n1413 VSS 0.00798f
C3546 VDD.n1414 VSS 0.00348f
C3547 VDD.n1415 VSS 0.00979f
C3548 VDD.n1416 VSS 0.00332f
C3549 VDD.n1417 VSS 0.00663f
C3550 VDD.n1418 VSS 0.00806f
C3551 VDD.n1419 VSS 0.00332f
C3552 VDD.n1420 VSS 0.00411f
C3553 VDD.n1421 VSS 0.00585f
C3554 VDD.n1422 VSS 0.00472f
C3555 VDD.n1423 VSS 0.00374f
C3556 VDD.n1424 VSS 0.0225f
C3557 VDD.n1425 VSS 0.0138f
C3558 VDD.n1426 VSS 0.0142f
C3559 VDD.n1427 VSS 3.26e-19
C3560 VDD.n1428 VSS 0.00488f
C3561 VDD.n1429 VSS 0.00798f
C3562 VDD.n1430 VSS 0.00374f
C3563 VDD.n1431 VSS 0.0225f
C3564 VDD.n1432 VSS 0.0225f
C3565 VDD.n1433 VSS 0.00488f
C3566 VDD.n1434 VSS 0.00439f
C3567 VDD.n1435 VSS 0.00806f
C3568 VDD.n1436 VSS 0.00332f
C3569 VDD.n1437 VSS 0.00663f
C3570 VDD.n1438 VSS 4.74e-19
C3571 VDD.n1439 VSS 0.00269f
C3572 VDD.n1440 VSS 0.00269f
C3573 VDD.n1441 VSS 0.00269f
C3574 VDD.n1442 VSS 0.00277f
C3575 VDD.n1443 VSS 0.0129f
C3576 VDD.n1444 VSS 0.198f
C3577 VDD.n1445 VSS 0.0104f
C3578 VDD.n1446 VSS 0.00979f
C3579 VDD.n1447 VSS 0.00979f
C3580 VDD.n1448 VSS 0.0129f
C3581 VDD.n1449 VSS 0.245f
C3582 VDD.n1450 VSS 0.0527f
C3583 VDD.n1451 VSS 0.00277f
C3584 VDD.n1452 VSS 0.00269f
C3585 VDD.n1453 VSS 3.16e-19
C3586 VDD.n1454 VSS 0.00269f
C3587 VDD.n1455 VSS 0.00348f
C3588 VDD.n1456 VSS 0.00269f
C3589 VDD.n1457 VSS 0.00332f
C3590 VDD.n1458 VSS 0.00979f
C3591 VDD.n1459 VSS 0.00979f
C3592 VDD.n1460 VSS 0.0129f
C3593 VDD.n1461 VSS 0.245f
C3594 VDD.n1462 VSS 0.0527f
C3595 VDD.n1463 VSS 0.198f
C3596 VDD.n1464 VSS 0.0104f
C3597 VDD.n1465 VSS 0.00979f
C3598 VDD.n1466 VSS 0.00269f
C3599 VDD.n1467 VSS 0.00916f
C3600 VDD.n1468 VSS 4.74e-19
C3601 VDD.n1469 VSS 0.00332f
C3602 VDD.n1470 VSS 0.00585f
C3603 VDD.n1471 VSS 0.00348f
C3604 VDD.n1472 VSS 4.74e-19
C3605 VDD.n1473 VSS -0.211f
C3606 VDD.n1474 VSS 3.26e-19
C3607 VDD.n1475 VSS 0.023f
C3608 VDD.n1476 VSS 0.00439f
C3609 VDD.n1477 VSS -0.174f
C3610 VDD.n1478 VSS 0.0138f
C3611 VDD.n1479 VSS -0.0844f
C3612 VDD.n1480 VSS 3.26e-19
C3613 VDD.n1481 VSS 0.00488f
C3614 VDD.n1482 VSS 0.00798f
C3615 VDD.n1483 VSS 0.00348f
C3616 VDD.n1484 VSS 0.00979f
C3617 VDD.n1485 VSS 0.00332f
C3618 VDD.n1486 VSS 0.00663f
C3619 VDD.n1487 VSS 0.00806f
C3620 VDD.n1488 VSS 0.00332f
C3621 VDD.n1489 VSS 0.00411f
C3622 VDD.n1490 VSS 0.00585f
C3623 VDD.n1491 VSS 0.00472f
C3624 VDD.n1492 VSS 0.00374f
C3625 VDD.n1493 VSS 0.0225f
C3626 VDD.n1494 VSS 0.0138f
C3627 VDD.n1495 VSS 0.0142f
C3628 VDD.n1496 VSS 3.26e-19
C3629 VDD.n1497 VSS 0.00488f
C3630 VDD.n1498 VSS 0.00798f
C3631 VDD.n1499 VSS 0.00374f
C3632 VDD.n1500 VSS 0.0225f
C3633 VDD.n1501 VSS 0.0809f
C3634 VDD.n1502 VSS 0.00488f
C3635 VDD.n1503 VSS 3.26e-19
C3636 VDD.n1504 VSS 0.00348f
C3637 VDD.n1505 VSS 0.00332f
C3638 VDD.n1506 VSS 0.00269f
C3639 VDD.n1507 VSS 0.00916f
C3640 VDD.n1508 VSS 0.00269f
C3641 VDD.n1509 VSS 0.00269f
C3642 VDD.n1510 VSS 0.00277f
C3643 VDD.n1511 VSS 0.0527f
C3644 VDD.n1512 VSS 0.00277f
C3645 VDD.n1513 VSS 0.00979f
C3646 VDD.n1514 VSS 0.245f
C3647 VDD.n1515 VSS 0.0129f
C3648 VDD.n1516 VSS 0.00979f
C3649 VDD.n1517 VSS 0.00269f
C3650 VDD.n1518 VSS 0.0294f
C3651 VDD.n1519 VSS 0.00332f
C3652 VDD.n1520 VSS 0.0286f
C3653 VDD.n1521 VSS 0.0294f
C3654 VDD.n1522 VSS 0.00332f
C3655 VDD.n1523 VSS 0.0261f
C3656 VDD.n1524 VSS 0.0261f
C3657 VDD.n1525 VSS 0.0286f
C3658 VDD.n1526 VSS 0.00348f
C3659 VDD.n1527 VSS 0.00269f
C3660 VDD.n1528 VSS 0.00269f
C3661 VDD.n1529 VSS 3.16e-19
C3662 VDD.n1530 VSS 0.0236f
C3663 VDD.n1531 VSS 0.124f
C3664 VDD.t66 VSS 0.47f
C3665 VDD.n1532 VSS 0.207f
C3666 VDD.t67 VSS 0.253f
C3667 VDD.n1533 VSS 0.198f
C3668 VDD.n1534 VSS 0.0104f
C3669 VDD.n1535 VSS 0.00269f
C3670 VDD.n1536 VSS 0.00663f
C3671 VDD.n1537 VSS 0.00348f
C3672 VDD.n1538 VSS 0.00806f
C3673 VDD.n1539 VSS 0.00332f
C3674 VDD.n1540 VSS 0.00781f
C3675 VDD.n1541 VSS 0.00439f
C3676 VDD.n1542 VSS 0.0138f
C3677 VDD.n1543 VSS 0.0142f
C3678 VDD.n1544 VSS -0.0753f
C3679 VDD.n1545 VSS 0.00411f
C3680 VDD.n1546 VSS 0.00585f
C3681 VDD.n1547 VSS -0.211f
C3682 VDD.n1548 VSS 0.00391f
C3683 VDD.n1549 VSS 0.023f
C3684 VDD.n1550 VSS 0.0225f
C3685 VDD.n1551 VSS -0.182f
C3686 VDD.n1552 VSS 0.00488f
C3687 VDD.n1553 VSS 3.26e-19
C3688 VDD.n1554 VSS 0.00348f
C3689 VDD.n1555 VSS 0.00332f
C3690 VDD.n1556 VSS 0.00269f
C3691 VDD.n1557 VSS 0.00916f
C3692 VDD.n1558 VSS 0.00269f
C3693 VDD.n1559 VSS 0.00269f
C3694 VDD.n1560 VSS 0.0129f
C3695 VDD.n1561 VSS 0.00277f
C3696 VDD.n1562 VSS 3.16e-19
C3697 VDD.n1563 VSS 0.00916f
C3698 VDD.n1564 VSS 0.00411f
C3699 VDD.n1565 VSS 0.00585f
C3700 VDD.n1566 VSS 0.00806f
C3701 VDD.n1567 VSS 0.00663f
C3702 VDD.n1568 VSS 0.00332f
C3703 VDD.n1569 VSS 0.00979f
C3704 VDD.n1570 VSS 0.00979f
C3705 VDD.n1571 VSS 0.00269f
C3706 VDD.n1572 VSS 0.00277f
C3707 VDD.n1573 VSS 0.0527f
C3708 VDD.n1574 VSS 0.245f
C3709 VDD.n1575 VSS 0.198f
C3710 VDD.n1576 VSS 0.0104f
C3711 VDD.n1577 VSS 0.00269f
C3712 VDD.n1578 VSS 0.00663f
C3713 VDD.n1579 VSS 0.00348f
C3714 VDD.n1580 VSS 0.00806f
C3715 VDD.n1581 VSS 0.00332f
C3716 VDD.n1582 VSS 0.00781f
C3717 VDD.n1583 VSS -0.0753f
C3718 VDD.n1584 VSS -0.078f
C3719 VDD.n1585 VSS 0.0142f
C3720 VDD.n1586 VSS 0.00439f
C3721 VDD.n1587 VSS 0.00411f
C3722 VDD.n1588 VSS 0.00585f
C3723 VDD.n1589 VSS 0.00488f
C3724 VDD.n1590 VSS 0.00391f
C3725 VDD.n1591 VSS 0.023f
C3726 VDD.n1592 VSS 0.0225f
C3727 VDD.n1593 VSS 0.0225f
C3728 VDD.n1594 VSS -0.211f
C3729 VDD.n1595 VSS 3.26e-19
C3730 VDD.n1596 VSS 0.00348f
C3731 VDD.n1597 VSS 0.00332f
C3732 VDD.n1598 VSS 0.00269f
C3733 VDD.n1599 VSS 0.00916f
C3734 VDD.n1600 VSS 0.00269f
C3735 VDD.n1601 VSS 0.00269f
C3736 VDD.n1602 VSS 0.0129f
C3737 VDD.n1603 VSS 0.00277f
C3738 VDD.n1604 VSS 3.16e-19
C3739 VDD.n1605 VSS 0.00916f
C3740 VDD.n1606 VSS 0.00411f
C3741 VDD.n1607 VSS 0.00585f
C3742 VDD.n1608 VSS 0.00806f
C3743 VDD.n1609 VSS 0.00663f
C3744 VDD.n1610 VSS 0.00332f
C3745 VDD.n1611 VSS 0.00979f
C3746 VDD.n1612 VSS 0.00979f
C3747 VDD.n1613 VSS 0.00269f
C3748 VDD.n1614 VSS 0.00277f
C3749 VDD.n1615 VSS 0.0527f
C3750 VDD.n1616 VSS 0.245f
C3751 VDD.n1617 VSS 0.198f
C3752 VDD.n1618 VSS 0.0104f
C3753 VDD.n1619 VSS 0.00269f
C3754 VDD.n1620 VSS 0.00663f
C3755 VDD.n1621 VSS 0.00348f
C3756 VDD.n1622 VSS 0.00806f
C3757 VDD.n1623 VSS 0.00332f
C3758 VDD.n1624 VSS 0.00781f
C3759 VDD.n1625 VSS 0.00439f
C3760 VDD.n1626 VSS 0.0138f
C3761 VDD.n1627 VSS 0.0142f
C3762 VDD.n1628 VSS 0.00439f
C3763 VDD.n1629 VSS 0.00411f
C3764 VDD.n1630 VSS 0.00585f
C3765 VDD.n1631 VSS 0.00488f
C3766 VDD.n1632 VSS 0.00391f
C3767 VDD.n1633 VSS 0.023f
C3768 VDD.n1634 VSS -0.182f
C3769 VDD.n1635 VSS 0.00488f
C3770 VDD.n1636 VSS 0.00472f
C3771 VDD.n1637 VSS -0.0844f
C3772 VDD.n1638 VSS 3.26e-19
C3773 VDD.n1639 VSS 0.00411f
C3774 VDD.n1640 VSS 0.00348f
C3775 VDD.n1641 VSS 0.00488f
C3776 VDD.n1642 VSS 0.0251f
C3777 VDD.n1643 VSS 0.0251f
C3778 VDD.n1644 VSS 0.00411f
C3779 VDD.n1645 VSS 0.0295f
C3780 VDD.n1646 VSS 0.0295f
C3781 VDD.n1647 VSS 0.00269f
C3782 VDD.n1648 VSS 0.00269f
C3783 VDD.n1649 VSS 0.00269f
C3784 VDD.n1650 VSS 0.00277f
C3785 VDD.n1651 VSS 0.0129f
C3786 VDD.n1652 VSS 3.16e-19
C3787 VDD.n1653 VSS 0.00269f
C3788 VDD.n1654 VSS 0.00277f
C3789 VDD.n1655 VSS 0.0527f
C3790 VDD.n1656 VSS 0.412f
C3791 VDD.n1657 VSS 0.0186f
C3792 VDD.n1658 VSS 0.03f
C3793 VDD.n1659 VSS 0.03f
C3794 VDD.n1660 VSS 0.0186f
C3795 VDD.n1661 VSS 0.226f
C3796 VDD.n1662 VSS 0.0527f
C3797 VDD.n1663 VSS 0.198f
C3798 VDD.n1664 VSS 0.0104f
C3799 VDD.n1665 VSS 0.00979f
C3800 VDD.n1666 VSS 0.00269f
C3801 VDD.n1667 VSS 0.00916f
C3802 VDD.n1668 VSS 4.74e-19
C3803 VDD.n1669 VSS 0.00332f
C3804 VDD.n1670 VSS 0.00585f
C3805 VDD.n1671 VSS 0.00348f
C3806 VDD.n1672 VSS 4.74e-19
C3807 VDD.n1673 VSS -0.211f
C3808 VDD.n1674 VSS 3.26e-19
C3809 VDD.n1675 VSS 0.023f
C3810 VDD.n1676 VSS 0.00439f
C3811 VDD.n1677 VSS -0.174f
C3812 VDD.n1678 VSS 0.00798f
C3813 VDD.n1679 VSS 0.00979f
C3814 VDD.n1680 VSS 0.00332f
C3815 VDD.n1681 VSS 0.00663f
C3816 VDD.n1682 VSS 0.00806f
C3817 VDD.n1683 VSS 0.00332f
C3818 VDD.n1684 VSS 0.00411f
C3819 VDD.n1685 VSS 0.00585f
C3820 VDD.n1686 VSS 0.00472f
C3821 VDD.n1687 VSS 0.00374f
C3822 VDD.n1688 VSS 0.0225f
C3823 VDD.n1689 VSS 0.0138f
C3824 VDD.n1690 VSS 0.0142f
C3825 VDD.n1691 VSS 3.26e-19
C3826 VDD.n1692 VSS 0.00488f
C3827 VDD.n1693 VSS 0.00798f
C3828 VDD.n1694 VSS 0.00374f
C3829 VDD.n1695 VSS 0.0225f
C3830 VDD.n1696 VSS 0.0225f
C3831 VDD.n1697 VSS 0.00488f
C3832 VDD.n1698 VSS 0.00439f
C3833 VDD.n1699 VSS 0.00806f
C3834 VDD.n1700 VSS 0.00332f
C3835 VDD.n1701 VSS 0.00663f
C3836 VDD.n1702 VSS 4.74e-19
C3837 VDD.n1703 VSS 0.00269f
C3838 VDD.n1704 VSS 0.00269f
C3839 VDD.n1705 VSS 0.00269f
C3840 VDD.n1706 VSS 0.00277f
C3841 VDD.n1707 VSS 0.0129f
C3842 VDD.n1708 VSS 0.198f
C3843 VDD.n1709 VSS 0.0104f
C3844 VDD.n1710 VSS 0.00979f
C3845 VDD.n1711 VSS 0.00979f
C3846 VDD.n1712 VSS 0.0129f
C3847 VDD.n1713 VSS 0.245f
C3848 VDD.n1714 VSS 0.0527f
C3849 VDD.n1715 VSS 0.00277f
C3850 VDD.n1716 VSS 0.00269f
C3851 VDD.n1717 VSS 3.16e-19
C3852 VDD.n1718 VSS 0.00269f
C3853 VDD.n1719 VSS 0.00348f
C3854 VDD.n1720 VSS 0.00269f
C3855 VDD.n1721 VSS 0.00332f
C3856 VDD.n1722 VSS 0.00979f
C3857 VDD.n1723 VSS 0.00979f
C3858 VDD.n1724 VSS 0.0129f
C3859 VDD.n1725 VSS 0.245f
C3860 VDD.n1726 VSS 0.0527f
C3861 VDD.n1727 VSS 0.198f
C3862 VDD.n1728 VSS 0.0104f
C3863 VDD.n1729 VSS 0.00979f
C3864 VDD.n1730 VSS 0.00269f
C3865 VDD.n1731 VSS 0.00916f
C3866 VDD.n1732 VSS 4.74e-19
C3867 VDD.n1733 VSS 0.00332f
C3868 VDD.n1734 VSS 0.00585f
C3869 VDD.n1735 VSS 0.00348f
C3870 VDD.n1736 VSS 4.74e-19
C3871 VDD.n1737 VSS -0.211f
C3872 VDD.n1738 VSS 3.26e-19
C3873 VDD.n1739 VSS 0.023f
C3874 VDD.n1740 VSS 0.00439f
C3875 VDD.n1741 VSS -0.174f
C3876 VDD.n1742 VSS 0.0138f
C3877 VDD.n1743 VSS -0.0844f
C3878 VDD.n1744 VSS 3.26e-19
C3879 VDD.n1745 VSS 0.00488f
C3880 VDD.n1746 VSS 0.00798f
C3881 VDD.n1747 VSS 0.00348f
C3882 VDD.n1748 VSS 0.00979f
C3883 VDD.n1749 VSS 0.00332f
C3884 VDD.n1750 VSS 0.00663f
C3885 VDD.n1751 VSS 0.00806f
C3886 VDD.n1752 VSS 0.00332f
C3887 VDD.n1753 VSS 0.00411f
C3888 VDD.n1754 VSS 0.00585f
C3889 VDD.n1755 VSS 0.00472f
C3890 VDD.n1756 VSS 0.00374f
C3891 VDD.n1757 VSS 0.0225f
C3892 VDD.n1758 VSS 0.0138f
C3893 VDD.n1759 VSS 0.0142f
C3894 VDD.n1760 VSS 3.26e-19
C3895 VDD.n1761 VSS 0.00488f
C3896 VDD.n1762 VSS 0.00798f
C3897 VDD.n1763 VSS 0.00374f
C3898 VDD.n1764 VSS 0.0225f
C3899 VDD.n1765 VSS 0.0809f
C3900 VDD.n1766 VSS 0.00488f
C3901 VDD.n1767 VSS 3.26e-19
C3902 VDD.n1768 VSS 0.00348f
C3903 VDD.n1769 VSS 0.00332f
C3904 VDD.n1770 VSS 0.00269f
C3905 VDD.n1771 VSS 0.00916f
C3906 VDD.n1772 VSS 0.00269f
C3907 VDD.n1773 VSS 0.00269f
C3908 VDD.n1774 VSS 0.00277f
C3909 VDD.n1775 VSS 0.0527f
C3910 VDD.n1776 VSS 0.00277f
C3911 VDD.n1777 VSS 0.00979f
C3912 VDD.n1778 VSS 0.245f
C3913 VDD.n1779 VSS 0.0129f
C3914 VDD.n1780 VSS 0.00979f
C3915 VDD.n1781 VSS 0.00269f
C3916 VDD.n1782 VSS 0.0294f
C3917 VDD.n1783 VSS 0.00332f
C3918 VDD.n1784 VSS 0.0286f
C3919 VDD.n1785 VSS 0.0294f
C3920 VDD.n1786 VSS 0.00332f
C3921 VDD.n1787 VSS 0.0261f
C3922 VDD.n1788 VSS 0.0261f
C3923 VDD.n1789 VSS 0.0286f
C3924 VDD.n1790 VSS 0.00348f
C3925 VDD.n1791 VSS 0.00269f
C3926 VDD.n1792 VSS 0.00269f
C3927 VDD.n1793 VSS 3.16e-19
C3928 VDD.n1794 VSS 0.0236f
C3929 VDD.n1795 VSS 0.124f
C3930 VDD.t20 VSS 0.47f
C3931 VDD.n1796 VSS 0.207f
C3932 VDD.t53 VSS 0.253f
C3933 VDD.n1797 VSS 0.198f
C3934 VDD.n1798 VSS 0.0104f
C3935 VDD.n1799 VSS 0.00269f
C3936 VDD.n1800 VSS 0.00663f
C3937 VDD.n1801 VSS 0.00348f
C3938 VDD.n1802 VSS 0.00806f
C3939 VDD.n1803 VSS 0.00332f
C3940 VDD.n1804 VSS 0.00781f
C3941 VDD.n1805 VSS 0.00439f
C3942 VDD.n1806 VSS 0.0138f
C3943 VDD.n1807 VSS 0.0142f
C3944 VDD.n1808 VSS -0.0753f
C3945 VDD.n1809 VSS 0.00411f
C3946 VDD.n1810 VSS 0.00585f
C3947 VDD.n1811 VSS -0.211f
C3948 VDD.n1812 VSS 0.00391f
C3949 VDD.n1813 VSS 0.023f
C3950 VDD.n1814 VSS 0.0225f
C3951 VDD.n1815 VSS -0.182f
C3952 VDD.n1816 VSS 0.00488f
C3953 VDD.n1817 VSS 3.26e-19
C3954 VDD.n1818 VSS 0.00348f
C3955 VDD.n1819 VSS 0.00332f
C3956 VDD.n1820 VSS 0.00269f
C3957 VDD.n1821 VSS 0.00916f
C3958 VDD.n1822 VSS 0.00269f
C3959 VDD.n1823 VSS 0.00269f
C3960 VDD.n1824 VSS 0.0129f
C3961 VDD.n1825 VSS 0.00277f
C3962 VDD.n1826 VSS 3.16e-19
C3963 VDD.n1827 VSS 0.00916f
C3964 VDD.n1828 VSS 0.00411f
C3965 VDD.n1829 VSS 0.00585f
C3966 VDD.n1830 VSS 0.00806f
C3967 VDD.n1831 VSS 0.00663f
C3968 VDD.n1832 VSS 0.00332f
C3969 VDD.n1833 VSS 0.00979f
C3970 VDD.n1834 VSS 0.00979f
C3971 VDD.n1835 VSS 0.00269f
C3972 VDD.n1836 VSS 0.00277f
C3973 VDD.n1837 VSS 0.0527f
C3974 VDD.n1838 VSS 0.245f
C3975 VDD.n1839 VSS 0.198f
C3976 VDD.n1840 VSS 0.0104f
C3977 VDD.n1841 VSS 0.00269f
C3978 VDD.n1842 VSS 0.00663f
C3979 VDD.n1843 VSS 0.00348f
C3980 VDD.n1844 VSS 0.00806f
C3981 VDD.n1845 VSS 0.00332f
C3982 VDD.n1846 VSS 0.00781f
C3983 VDD.n1847 VSS -0.0753f
C3984 VDD.n1848 VSS -0.078f
C3985 VDD.n1849 VSS 0.0142f
C3986 VDD.n1850 VSS 0.00439f
C3987 VDD.n1851 VSS 0.00411f
C3988 VDD.n1852 VSS 0.00585f
C3989 VDD.n1853 VSS 0.00488f
C3990 VDD.n1854 VSS 0.00391f
C3991 VDD.n1855 VSS 0.023f
C3992 VDD.n1856 VSS 0.0225f
C3993 VDD.n1857 VSS 0.0225f
C3994 VDD.n1858 VSS -0.211f
C3995 VDD.n1859 VSS 3.26e-19
C3996 VDD.n1860 VSS 0.00348f
C3997 VDD.n1861 VSS 0.00332f
C3998 VDD.n1862 VSS 0.00269f
C3999 VDD.n1863 VSS 0.00916f
C4000 VDD.n1864 VSS 0.00269f
C4001 VDD.n1865 VSS 0.00269f
C4002 VDD.n1866 VSS 0.0129f
C4003 VDD.n1867 VSS 0.00277f
C4004 VDD.n1868 VSS 3.16e-19
C4005 VDD.n1869 VSS 0.00916f
C4006 VDD.n1870 VSS 0.00411f
C4007 VDD.n1871 VSS 0.00585f
C4008 VDD.n1872 VSS 0.00806f
C4009 VDD.n1873 VSS 0.00663f
C4010 VDD.n1874 VSS 0.00332f
C4011 VDD.n1875 VSS 0.00979f
C4012 VDD.n1876 VSS 0.00979f
C4013 VDD.n1877 VSS 0.00269f
C4014 VDD.n1878 VSS 0.00277f
C4015 VDD.n1879 VSS 0.0527f
C4016 VDD.n1880 VSS 0.245f
C4017 VDD.n1881 VSS 0.198f
C4018 VDD.n1882 VSS 0.0104f
C4019 VDD.n1883 VSS 0.00269f
C4020 VDD.n1884 VSS 0.00663f
C4021 VDD.n1885 VSS 0.00348f
C4022 VDD.n1886 VSS 0.00806f
C4023 VDD.n1887 VSS 0.00332f
C4024 VDD.n1888 VSS 0.00781f
C4025 VDD.n1889 VSS 0.00439f
C4026 VDD.n1890 VSS 0.0138f
C4027 VDD.n1891 VSS 0.0142f
C4028 VDD.n1892 VSS 0.00439f
C4029 VDD.n1893 VSS 0.00411f
C4030 VDD.n1894 VSS 0.00585f
C4031 VDD.n1895 VSS 0.00488f
C4032 VDD.n1896 VSS 0.00391f
C4033 VDD.n1897 VSS 0.023f
C4034 VDD.n1898 VSS -0.182f
C4035 VDD.n1899 VSS 0.00488f
C4036 VDD.n1900 VSS 0.00472f
C4037 VDD.n1901 VSS -0.0844f
C4038 VDD.n1902 VSS 3.26e-19
C4039 VDD.n1903 VSS 0.00411f
C4040 VDD.n1904 VSS 0.00348f
C4041 VDD.n1905 VSS 0.00488f
C4042 VDD.n1906 VSS 0.0251f
C4043 VDD.n1907 VSS 0.0251f
C4044 VDD.n1908 VSS 0.00411f
C4045 VDD.n1909 VSS 0.0295f
C4046 VDD.n1910 VSS 0.0295f
C4047 VDD.n1911 VSS 0.00269f
C4048 VDD.n1912 VSS 0.00269f
C4049 VDD.n1913 VSS 0.00269f
C4050 VDD.n1914 VSS 0.00277f
C4051 VDD.n1915 VSS 0.0129f
C4052 VDD.n1916 VSS 3.16e-19
C4053 VDD.n1917 VSS 0.00269f
C4054 VDD.n1918 VSS 0.00277f
C4055 VDD.n1919 VSS 0.0527f
C4056 VDD.n1920 VSS 0.412f
C4057 VDD.n1921 VSS 0.0186f
C4058 VDD.n1922 VSS 0.03f
C4059 VDD.n1923 VSS 0.03f
C4060 VDD.n1924 VSS 0.0186f
C4061 VDD.n1925 VSS 0.226f
C4062 VDD.n1926 VSS 0.0527f
C4063 VDD.n1927 VSS 0.198f
C4064 VDD.n1928 VSS 0.0104f
C4065 VDD.n1929 VSS 0.00979f
C4066 VDD.n1930 VSS 0.00269f
C4067 VDD.n1931 VSS 0.00916f
C4068 VDD.n1932 VSS 4.74e-19
C4069 VDD.n1933 VSS 0.00332f
C4070 VDD.n1934 VSS 0.00585f
C4071 VDD.n1935 VSS 0.00348f
C4072 VDD.n1936 VSS 4.74e-19
C4073 VDD.n1937 VSS -0.211f
C4074 VDD.n1938 VSS 3.26e-19
C4075 VDD.n1939 VSS 0.023f
C4076 VDD.n1940 VSS 0.00439f
C4077 VDD.n1941 VSS -0.174f
C4078 VDD.n1942 VSS 0.00798f
C4079 VDD.n1943 VSS 0.00979f
C4080 VDD.n1944 VSS 0.00332f
C4081 VDD.n1945 VSS 0.00663f
C4082 VDD.n1946 VSS 0.00806f
C4083 VDD.n1947 VSS 0.00332f
C4084 VDD.n1948 VSS 0.00411f
C4085 VDD.n1949 VSS 0.00585f
C4086 VDD.n1950 VSS 0.00472f
C4087 VDD.n1951 VSS 0.00374f
C4088 VDD.n1952 VSS 0.0225f
C4089 VDD.n1953 VSS 0.0138f
C4090 VDD.n1954 VSS 0.0142f
C4091 VDD.n1955 VSS 3.26e-19
C4092 VDD.n1956 VSS 0.00488f
C4093 VDD.n1957 VSS 0.00798f
C4094 VDD.n1958 VSS 0.00374f
C4095 VDD.n1959 VSS 0.0225f
C4096 VDD.n1960 VSS 0.0225f
C4097 VDD.n1961 VSS 0.00488f
C4098 VDD.n1962 VSS 0.00439f
C4099 VDD.n1963 VSS 0.00806f
C4100 VDD.n1964 VSS 0.00332f
C4101 VDD.n1965 VSS 0.00663f
C4102 VDD.n1966 VSS 4.74e-19
C4103 VDD.n1967 VSS 0.00269f
C4104 VDD.n1968 VSS 0.00269f
C4105 VDD.n1969 VSS 0.00269f
C4106 VDD.n1970 VSS 0.00277f
C4107 VDD.n1971 VSS 0.0129f
C4108 VDD.n1972 VSS 0.198f
C4109 VDD.n1973 VSS 0.0104f
C4110 VDD.n1974 VSS 0.00979f
C4111 VDD.n1975 VSS 0.00979f
C4112 VDD.n1976 VSS 0.0129f
C4113 VDD.n1977 VSS 0.245f
C4114 VDD.n1978 VSS 0.0527f
C4115 VDD.n1979 VSS 0.00277f
C4116 VDD.n1980 VSS 0.00269f
C4117 VDD.n1981 VSS 3.16e-19
C4118 VDD.n1982 VSS 0.00269f
C4119 VDD.n1983 VSS 0.00348f
C4120 VDD.n1984 VSS 0.00269f
C4121 VDD.n1985 VSS 0.00332f
C4122 VDD.n1986 VSS 0.00979f
C4123 VDD.n1987 VSS 0.00979f
C4124 VDD.n1988 VSS 0.0129f
C4125 VDD.n1989 VSS 0.245f
C4126 VDD.n1990 VSS 0.0527f
C4127 VDD.n1991 VSS 0.198f
C4128 VDD.n1992 VSS 0.0104f
C4129 VDD.n1993 VSS 0.00979f
C4130 VDD.n1994 VSS 0.00269f
C4131 VDD.n1995 VSS 0.00916f
C4132 VDD.n1996 VSS 4.74e-19
C4133 VDD.n1997 VSS 0.00332f
C4134 VDD.n1998 VSS 0.00585f
C4135 VDD.n1999 VSS 0.00348f
C4136 VDD.n2000 VSS 4.74e-19
C4137 VDD.n2001 VSS -0.211f
C4138 VDD.n2002 VSS 3.26e-19
C4139 VDD.n2003 VSS 0.023f
C4140 VDD.n2004 VSS 0.00439f
C4141 VDD.n2005 VSS -0.174f
C4142 VDD.n2006 VSS 0.0138f
C4143 VDD.n2007 VSS -0.0844f
C4144 VDD.n2008 VSS 3.26e-19
C4145 VDD.n2009 VSS 0.00488f
C4146 VDD.n2010 VSS 0.00798f
C4147 VDD.n2011 VSS 0.00348f
C4148 VDD.n2012 VSS 0.00979f
C4149 VDD.n2013 VSS 0.00332f
C4150 VDD.n2014 VSS 0.00663f
C4151 VDD.n2015 VSS 0.00806f
C4152 VDD.n2016 VSS 0.00332f
C4153 VDD.n2017 VSS 0.00411f
C4154 VDD.n2018 VSS 0.00585f
C4155 VDD.n2019 VSS 0.00472f
C4156 VDD.n2020 VSS 0.00374f
C4157 VDD.n2021 VSS 0.0225f
C4158 VDD.n2022 VSS 0.0138f
C4159 VDD.n2023 VSS 0.0142f
C4160 VDD.n2024 VSS 3.26e-19
C4161 VDD.n2025 VSS 0.00488f
C4162 VDD.n2026 VSS 0.00798f
C4163 VDD.n2027 VSS 0.00374f
C4164 VDD.n2028 VSS 0.0225f
C4165 VDD.n2029 VSS 0.0809f
C4166 VDD.n2030 VSS 0.00488f
C4167 VDD.n2031 VSS 3.26e-19
C4168 VDD.n2032 VSS 0.00348f
C4169 VDD.n2033 VSS 0.00332f
C4170 VDD.n2034 VSS 0.00269f
C4171 VDD.n2035 VSS 0.00916f
C4172 VDD.n2036 VSS 0.00269f
C4173 VDD.n2037 VSS 0.00269f
C4174 VDD.n2038 VSS 0.00277f
C4175 VDD.n2039 VSS 0.0527f
C4176 VDD.n2040 VSS 0.00277f
C4177 VDD.n2041 VSS 0.00979f
C4178 VDD.n2042 VSS 0.245f
C4179 VDD.n2043 VSS 0.0129f
C4180 VDD.n2044 VSS 0.00979f
C4181 VDD.n2045 VSS 0.00269f
C4182 VDD.n2046 VSS 0.0294f
C4183 VDD.n2047 VSS 0.00332f
C4184 VDD.n2048 VSS 0.0286f
C4185 VDD.n2049 VSS 0.0294f
C4186 VDD.n2050 VSS 0.00332f
C4187 VDD.n2051 VSS 0.0261f
C4188 VDD.n2052 VSS 0.0261f
C4189 VDD.n2053 VSS 0.0286f
C4190 VDD.n2054 VSS 0.00348f
C4191 VDD.n2055 VSS 0.00269f
C4192 VDD.n2056 VSS 0.00269f
C4193 VDD.n2057 VSS 3.16e-19
C4194 VDD.n2058 VSS 0.0236f
C4195 VDD.n2059 VSS 0.124f
C4196 VDD.t72 VSS 0.47f
C4197 VDD.n2060 VSS 0.207f
C4198 VDD.t38 VSS 0.253f
C4199 VDD.n2061 VSS 0.198f
C4200 VDD.n2062 VSS 0.0104f
C4201 VDD.n2063 VSS 0.00269f
C4202 VDD.n2064 VSS 0.00663f
C4203 VDD.n2065 VSS 0.00348f
C4204 VDD.n2066 VSS 0.00806f
C4205 VDD.n2067 VSS 0.00332f
C4206 VDD.n2068 VSS 0.00781f
C4207 VDD.n2069 VSS 0.00439f
C4208 VDD.n2070 VSS 0.0138f
C4209 VDD.n2071 VSS 0.0142f
C4210 VDD.n2072 VSS -0.0753f
C4211 VDD.n2073 VSS 0.00411f
C4212 VDD.n2074 VSS 0.00585f
C4213 VDD.n2075 VSS -0.211f
C4214 VDD.n2076 VSS 0.00391f
C4215 VDD.n2077 VSS 0.023f
C4216 VDD.n2078 VSS 0.0225f
C4217 VDD.n2079 VSS -0.182f
C4218 VDD.n2080 VSS 0.00488f
C4219 VDD.n2081 VSS 3.26e-19
C4220 VDD.n2082 VSS 0.00348f
C4221 VDD.n2083 VSS 0.00332f
C4222 VDD.n2084 VSS 0.00269f
C4223 VDD.n2085 VSS 0.00916f
C4224 VDD.n2086 VSS 0.00269f
C4225 VDD.n2087 VSS 0.00269f
C4226 VDD.n2088 VSS 0.0129f
C4227 VDD.n2089 VSS 0.00277f
C4228 VDD.n2090 VSS 3.16e-19
C4229 VDD.n2091 VSS 0.00916f
C4230 VDD.n2092 VSS 0.00411f
C4231 VDD.n2093 VSS 0.00585f
C4232 VDD.n2094 VSS 0.00806f
C4233 VDD.n2095 VSS 0.00663f
C4234 VDD.n2096 VSS 0.00332f
C4235 VDD.n2097 VSS 0.00979f
C4236 VDD.n2098 VSS 0.00979f
C4237 VDD.n2099 VSS 0.00269f
C4238 VDD.n2100 VSS 0.00277f
C4239 VDD.n2101 VSS 0.0527f
C4240 VDD.n2102 VSS 0.245f
C4241 VDD.n2103 VSS 0.198f
C4242 VDD.n2104 VSS 0.0104f
C4243 VDD.n2105 VSS 0.00269f
C4244 VDD.n2106 VSS 0.00663f
C4245 VDD.n2107 VSS 0.00348f
C4246 VDD.n2108 VSS 0.00806f
C4247 VDD.n2109 VSS 0.00332f
C4248 VDD.n2110 VSS 0.00781f
C4249 VDD.n2111 VSS -0.0753f
C4250 VDD.n2112 VSS -0.078f
C4251 VDD.n2113 VSS 0.0142f
C4252 VDD.n2114 VSS 0.00439f
C4253 VDD.n2115 VSS 0.00411f
C4254 VDD.n2116 VSS 0.00585f
C4255 VDD.n2117 VSS 0.00488f
C4256 VDD.n2118 VSS 0.00391f
C4257 VDD.n2119 VSS 0.023f
C4258 VDD.n2120 VSS 0.0225f
C4259 VDD.n2121 VSS 0.0225f
C4260 VDD.n2122 VSS -0.211f
C4261 VDD.n2123 VSS 3.26e-19
C4262 VDD.n2124 VSS 0.00348f
C4263 VDD.n2125 VSS 0.00332f
C4264 VDD.n2126 VSS 0.00269f
C4265 VDD.n2127 VSS 0.00916f
C4266 VDD.n2128 VSS 0.00269f
C4267 VDD.n2129 VSS 0.00269f
C4268 VDD.n2130 VSS 0.0129f
C4269 VDD.n2131 VSS 0.00277f
C4270 VDD.n2132 VSS 3.16e-19
C4271 VDD.n2133 VSS 0.00916f
C4272 VDD.n2134 VSS 0.00411f
C4273 VDD.n2135 VSS 0.00585f
C4274 VDD.n2136 VSS 0.00806f
C4275 VDD.n2137 VSS 0.00663f
C4276 VDD.n2138 VSS 0.00332f
C4277 VDD.n2139 VSS 0.00979f
C4278 VDD.n2140 VSS 0.00979f
C4279 VDD.n2141 VSS 0.00269f
C4280 VDD.n2142 VSS 0.00277f
C4281 VDD.n2143 VSS 0.0527f
C4282 VDD.n2144 VSS 0.245f
C4283 VDD.n2145 VSS 0.198f
C4284 VDD.n2146 VSS 0.0104f
C4285 VDD.n2147 VSS 0.00269f
C4286 VDD.n2148 VSS 0.00663f
C4287 VDD.n2149 VSS 0.00348f
C4288 VDD.n2150 VSS 0.00806f
C4289 VDD.n2151 VSS 0.00332f
C4290 VDD.n2152 VSS 0.00781f
C4291 VDD.n2153 VSS 0.00439f
C4292 VDD.n2154 VSS 0.0138f
C4293 VDD.n2155 VSS 0.0142f
C4294 VDD.n2156 VSS 0.00439f
C4295 VDD.n2157 VSS 0.00411f
C4296 VDD.n2158 VSS 0.00585f
C4297 VDD.n2159 VSS 0.00488f
C4298 VDD.n2160 VSS 0.00391f
C4299 VDD.n2161 VSS 0.023f
C4300 VDD.n2162 VSS -0.182f
C4301 VDD.n2163 VSS 0.00488f
C4302 VDD.n2164 VSS 0.00472f
C4303 VDD.n2165 VSS -0.0844f
C4304 VDD.n2166 VSS 3.26e-19
C4305 VDD.n2167 VSS 0.00411f
C4306 VDD.n2168 VSS 0.00348f
C4307 VDD.n2169 VSS 0.00488f
C4308 VDD.n2170 VSS 0.0251f
C4309 VDD.n2171 VSS 0.0251f
C4310 VDD.n2172 VSS 0.00411f
C4311 VDD.n2173 VSS 0.0295f
C4312 VDD.n2174 VSS 0.0295f
C4313 VDD.n2175 VSS 0.00269f
C4314 VDD.n2176 VSS 0.00269f
C4315 VDD.n2177 VSS 0.00269f
C4316 VDD.n2178 VSS 0.00277f
C4317 VDD.n2179 VSS 0.0129f
C4318 VDD.n2180 VSS 3.16e-19
C4319 VDD.n2181 VSS 0.00269f
C4320 VDD.n2182 VSS 0.00277f
C4321 VDD.n2183 VSS 0.0527f
C4322 VDD.n2184 VSS 0.412f
C4323 VDD.n2185 VSS 0.0186f
C4324 VDD.n2186 VSS 0.03f
C4325 VDD.n2187 VSS 0.03f
C4326 VDD.n2188 VSS 0.0186f
C4327 VDD.n2189 VSS 0.226f
C4328 VDD.n2190 VSS 0.0527f
C4329 VDD.n2191 VSS 0.198f
C4330 VDD.n2192 VSS 0.0104f
C4331 VDD.n2193 VSS 0.00979f
C4332 VDD.n2194 VSS 0.00269f
C4333 VDD.n2195 VSS 0.00916f
C4334 VDD.n2196 VSS 4.74e-19
C4335 VDD.n2197 VSS 0.00332f
C4336 VDD.n2198 VSS 0.00585f
C4337 VDD.n2199 VSS 0.00348f
C4338 VDD.n2200 VSS 4.74e-19
C4339 VDD.n2201 VSS -0.211f
C4340 VDD.n2202 VSS 3.26e-19
C4341 VDD.n2203 VSS 0.023f
C4342 VDD.n2204 VSS 0.00439f
C4343 VDD.n2205 VSS -0.174f
C4344 VDD.n2206 VSS 0.00798f
C4345 VDD.n2207 VSS 0.00979f
C4346 VDD.n2208 VSS 0.00332f
C4347 VDD.n2209 VSS 0.00663f
C4348 VDD.n2210 VSS 0.00806f
C4349 VDD.n2211 VSS 0.00332f
C4350 VDD.n2212 VSS 0.00411f
C4351 VDD.n2213 VSS 0.00585f
C4352 VDD.n2214 VSS 0.00472f
C4353 VDD.n2215 VSS 0.00374f
C4354 VDD.n2216 VSS 0.0225f
C4355 VDD.n2217 VSS 0.0138f
C4356 VDD.n2218 VSS 0.0142f
C4357 VDD.n2219 VSS 3.26e-19
C4358 VDD.n2220 VSS 0.00488f
C4359 VDD.n2221 VSS 0.00798f
C4360 VDD.n2222 VSS 0.00374f
C4361 VDD.n2223 VSS 0.0225f
C4362 VDD.n2224 VSS 0.0225f
C4363 VDD.n2225 VSS 0.00488f
C4364 VDD.n2226 VSS 0.00439f
C4365 VDD.n2227 VSS 0.00806f
C4366 VDD.n2228 VSS 0.00332f
C4367 VDD.n2229 VSS 0.00663f
C4368 VDD.n2230 VSS 4.74e-19
C4369 VDD.n2231 VSS 0.00269f
C4370 VDD.n2232 VSS 0.00269f
C4371 VDD.n2233 VSS 0.00269f
C4372 VDD.n2234 VSS 0.00277f
C4373 VDD.n2235 VSS 0.0129f
C4374 VDD.n2236 VSS 0.198f
C4375 VDD.n2237 VSS 0.0104f
C4376 VDD.n2238 VSS 0.00979f
C4377 VDD.n2239 VSS 0.00979f
C4378 VDD.n2240 VSS 0.0129f
C4379 VDD.n2241 VSS 0.245f
C4380 VDD.n2242 VSS 0.0527f
C4381 VDD.n2243 VSS 0.00277f
C4382 VDD.n2244 VSS 0.00269f
C4383 VDD.n2245 VSS 3.16e-19
C4384 VDD.n2246 VSS 0.00269f
C4385 VDD.n2247 VSS 0.00348f
C4386 VDD.n2248 VSS 0.00269f
C4387 VDD.n2249 VSS 0.00332f
C4388 VDD.n2250 VSS 0.00979f
C4389 VDD.n2251 VSS 0.00979f
C4390 VDD.n2252 VSS 0.0129f
C4391 VDD.n2253 VSS 0.245f
C4392 VDD.n2254 VSS 0.0527f
C4393 VDD.n2255 VSS 0.198f
C4394 VDD.n2256 VSS 0.0104f
C4395 VDD.n2257 VSS 0.00979f
C4396 VDD.n2258 VSS 0.00269f
C4397 VDD.n2259 VSS 0.00916f
C4398 VDD.n2260 VSS 4.74e-19
C4399 VDD.n2261 VSS 0.00332f
C4400 VDD.n2262 VSS 0.00585f
C4401 VDD.n2263 VSS 0.00348f
C4402 VDD.n2264 VSS 4.74e-19
C4403 VDD.n2265 VSS -0.211f
C4404 VDD.n2266 VSS 3.26e-19
C4405 VDD.n2267 VSS 0.023f
C4406 VDD.n2268 VSS 0.00439f
C4407 VDD.n2269 VSS -0.174f
C4408 VDD.n2270 VSS 0.0138f
C4409 VDD.n2271 VSS -0.0844f
C4410 VDD.n2272 VSS 3.26e-19
C4411 VDD.n2273 VSS 0.00488f
C4412 VDD.n2274 VSS 0.00798f
C4413 VDD.n2275 VSS 0.00348f
C4414 VDD.n2276 VSS 0.00979f
C4415 VDD.n2277 VSS 0.00332f
C4416 VDD.n2278 VSS 0.00663f
C4417 VDD.n2279 VSS 0.00806f
C4418 VDD.n2280 VSS 0.00332f
C4419 VDD.n2281 VSS 0.00411f
C4420 VDD.n2282 VSS 0.00585f
C4421 VDD.n2283 VSS 0.00472f
C4422 VDD.n2284 VSS 0.00374f
C4423 VDD.n2285 VSS 0.0225f
C4424 VDD.n2286 VSS 0.0138f
C4425 VDD.n2287 VSS 0.0142f
C4426 VDD.n2288 VSS 3.26e-19
C4427 VDD.n2289 VSS 0.00488f
C4428 VDD.n2290 VSS 0.00798f
C4429 VDD.n2291 VSS 0.00374f
C4430 VDD.n2292 VSS 0.0225f
C4431 VDD.n2293 VSS 0.0809f
C4432 VDD.n2294 VSS 0.00488f
C4433 VDD.n2295 VSS 3.26e-19
C4434 VDD.n2296 VSS 0.00348f
C4435 VDD.n2297 VSS 0.00332f
C4436 VDD.n2298 VSS 0.00269f
C4437 VDD.n2299 VSS 0.00916f
C4438 VDD.n2300 VSS 0.00269f
C4439 VDD.n2301 VSS 0.00269f
C4440 VDD.n2302 VSS 0.00277f
C4441 VDD.n2303 VSS 0.0527f
C4442 VDD.n2304 VSS 0.00277f
C4443 VDD.n2305 VSS 0.00979f
C4444 VDD.n2306 VSS 0.245f
C4445 VDD.n2307 VSS 0.0129f
C4446 VDD.n2308 VSS 0.00979f
C4447 VDD.n2309 VSS 0.00269f
C4448 VDD.n2310 VSS 0.0294f
C4449 VDD.n2311 VSS 0.00332f
C4450 VDD.n2312 VSS 0.0286f
C4451 VDD.n2313 VSS 0.0294f
C4452 VDD.n2314 VSS 0.00332f
C4453 VDD.n2315 VSS 0.0261f
C4454 VDD.n2316 VSS 0.0261f
C4455 VDD.n2317 VSS 0.0286f
C4456 VDD.n2318 VSS 0.00348f
C4457 VDD.n2319 VSS 0.00269f
C4458 VDD.n2320 VSS 0.00269f
C4459 VDD.n2321 VSS 3.16e-19
C4460 VDD.n2322 VSS 0.0236f
C4461 VDD.n2323 VSS 0.124f
C4462 VDD.t28 VSS 0.47f
C4463 VDD.n2324 VSS 0.207f
C4464 VDD.t65 VSS 0.253f
C4465 VDD.n2325 VSS 0.198f
C4466 VDD.n2326 VSS 0.0104f
C4467 VDD.n2327 VSS 0.00269f
C4468 VDD.n2328 VSS 0.00663f
C4469 VDD.n2329 VSS 0.00348f
C4470 VDD.n2330 VSS 0.00806f
C4471 VDD.n2331 VSS 0.00332f
C4472 VDD.n2332 VSS 0.00781f
C4473 VDD.n2333 VSS 0.00439f
C4474 VDD.n2334 VSS 0.0138f
C4475 VDD.n2335 VSS 0.0142f
C4476 VDD.n2336 VSS -0.0753f
C4477 VDD.n2337 VSS 0.00411f
C4478 VDD.n2338 VSS 0.00585f
C4479 VDD.n2339 VSS -0.211f
C4480 VDD.n2340 VSS 0.00391f
C4481 VDD.n2341 VSS 0.023f
C4482 VDD.n2342 VSS 0.0225f
C4483 VDD.n2343 VSS -0.182f
C4484 VDD.n2344 VSS 0.00488f
C4485 VDD.n2345 VSS 3.26e-19
C4486 VDD.n2346 VSS 0.00348f
C4487 VDD.n2347 VSS 0.00332f
C4488 VDD.n2348 VSS 0.00269f
C4489 VDD.n2349 VSS 0.00916f
C4490 VDD.n2350 VSS 0.00269f
C4491 VDD.n2351 VSS 0.00269f
C4492 VDD.n2352 VSS 0.0129f
C4493 VDD.n2353 VSS 0.00277f
C4494 VDD.n2354 VSS 3.16e-19
C4495 VDD.n2355 VSS 0.00916f
C4496 VDD.n2356 VSS 0.00411f
C4497 VDD.n2357 VSS 0.00585f
C4498 VDD.n2358 VSS 0.00806f
C4499 VDD.n2359 VSS 0.00663f
C4500 VDD.n2360 VSS 0.00332f
C4501 VDD.n2361 VSS 0.00979f
C4502 VDD.n2362 VSS 0.00979f
C4503 VDD.n2363 VSS 0.00269f
C4504 VDD.n2364 VSS 0.00277f
C4505 VDD.n2365 VSS 0.0527f
C4506 VDD.n2366 VSS 0.245f
C4507 VDD.n2367 VSS 0.198f
C4508 VDD.n2368 VSS 0.0104f
C4509 VDD.n2369 VSS 0.00269f
C4510 VDD.n2370 VSS 0.00663f
C4511 VDD.n2371 VSS 0.00348f
C4512 VDD.n2372 VSS 0.00806f
C4513 VDD.n2373 VSS 0.00332f
C4514 VDD.n2374 VSS 0.00781f
C4515 VDD.n2375 VSS -0.0753f
C4516 VDD.n2376 VSS -0.078f
C4517 VDD.n2377 VSS 0.0142f
C4518 VDD.n2378 VSS 0.00439f
C4519 VDD.n2379 VSS 0.00411f
C4520 VDD.n2380 VSS 0.00585f
C4521 VDD.n2381 VSS 0.00488f
C4522 VDD.n2382 VSS 0.00391f
C4523 VDD.n2383 VSS 0.023f
C4524 VDD.n2384 VSS 0.0225f
C4525 VDD.n2385 VSS 0.0225f
C4526 VDD.n2386 VSS -0.211f
C4527 VDD.n2387 VSS 3.26e-19
C4528 VDD.n2388 VSS 0.00348f
C4529 VDD.n2389 VSS 0.00332f
C4530 VDD.n2390 VSS 0.00269f
C4531 VDD.n2391 VSS 0.00916f
C4532 VDD.n2392 VSS 0.00269f
C4533 VDD.n2393 VSS 0.00269f
C4534 VDD.n2394 VSS 0.0129f
C4535 VDD.n2395 VSS 0.00277f
C4536 VDD.n2396 VSS 3.16e-19
C4537 VDD.n2397 VSS 0.00916f
C4538 VDD.n2398 VSS 0.00411f
C4539 VDD.n2399 VSS 0.00585f
C4540 VDD.n2400 VSS 0.00806f
C4541 VDD.n2401 VSS 0.00663f
C4542 VDD.n2402 VSS 0.00332f
C4543 VDD.n2403 VSS 0.00979f
C4544 VDD.n2404 VSS 0.00979f
C4545 VDD.n2405 VSS 0.00269f
C4546 VDD.n2406 VSS 0.00277f
C4547 VDD.n2407 VSS 0.0527f
C4548 VDD.n2408 VSS 0.245f
C4549 VDD.n2409 VSS 0.198f
C4550 VDD.n2410 VSS 0.0104f
C4551 VDD.n2411 VSS 0.00269f
C4552 VDD.n2412 VSS 0.00663f
C4553 VDD.n2413 VSS 0.0422f
C4554 VDD.n2414 VSS 0.00806f
C4555 VDD.n2415 VSS 0.00332f
C4556 VDD.n2416 VSS 0.00781f
C4557 VDD.n2417 VSS 0.00439f
C4558 VDD.n2418 VSS 0.0138f
C4559 VDD.n2419 VSS 0.0142f
C4560 VDD.n2420 VSS 0.00439f
C4561 VDD.n2421 VSS 0.00411f
C4562 VDD.n2422 VSS 0.00585f
C4563 VDD.n2423 VSS 0.00488f
C4564 VDD.n2424 VSS 0.00391f
C4565 VDD.n2425 VSS 0.023f
C4566 VDD.n2426 VSS -0.182f
C4567 VDD.n2427 VSS 0.0891f
C4568 VDD.n2428 VSS 0.028f
C4569 VDD.n2429 VSS 0.0174f
C4570 VDD.n2430 VSS 0.0084f
C4571 VDD.n2431 VSS 0.00411f
C4572 VDD.n2432 VSS 0.00759f
C4573 VDD.n2433 VSS 3.26e-19
C4574 VDD.n2434 VSS 0.00332f
C4575 VDD.n2435 VSS 0.0303f
C4576 VDD.n2436 VSS 0.0145f
C4577 VDD.n2437 VSS 0.0229f
C4578 VDD.n2438 VSS 0.00488f
C4579 VDD.n2439 VSS 0.00439f
C4580 VDD.n2440 VSS 0.00806f
C4581 VDD.n2441 VSS 0.00332f
C4582 VDD.n2442 VSS 0.00663f
C4583 VDD.n2443 VSS 4.74e-19
C4584 VDD.n2444 VSS 0.00269f
C4585 VDD.n2445 VSS 0.00269f
C4586 VDD.n2446 VSS 0.00269f
C4587 VDD.n2447 VSS 0.00277f
C4588 VDD.n2448 VSS 0.0129f
C4589 VDD.n2449 VSS 0.198f
C4590 VDD.n2450 VSS 0.0104f
C4591 VDD.n2451 VSS 0.00269f
C4592 VDD.n2452 VSS 0.0158f
C4593 VDD.n2453 VSS 0.0087f
C4594 VDD.n2454 VSS 0.0186f
C4595 VDD.t44 VSS 0.299f
C4596 VDD.n2455 VSS 0.014f
C4597 VDD.n2456 VSS 0.0106f
C4598 VDD.t45 VSS 0.0509f
C4599 VDD.n2457 VSS 0.0207f
C4600 VDD.n2458 VSS 8.15e-19
C4601 VDD.n2459 VSS 0.0124f
C4602 VDD.n2460 VSS 0.0185f
C4603 VDD.n2461 VSS 0.00689f
C4604 VDD.n2462 VSS 0.0186f
C4605 VDD.n2463 VSS 0.0069f
C4606 VDD.n2464 VSS 0.00443f
C4607 VDD.n2465 VSS 0.119f
C4608 VDD.n2466 VSS 0.016f
C4609 VDD.n2467 VSS 0.017f
C4610 VDD.n2468 VSS 0.0409f
C4611 VDD.n2469 VSS 0.0232f
C4612 VDD.n2470 VSS 0.0069f
C4613 VDD.n2471 VSS 0.0193f
C4614 VDD.t59 VSS 0.0509f
C4615 VDD.n2472 VSS 0.0556f
C4616 VDD.n2473 VSS 0.00797f
C4617 VDD.n2474 VSS 0.00256f
C4618 VDD.n2475 VSS 0.00483f
C4619 VDD.n2476 VSS 0.0108f
C4620 VDD.n2477 VSS 0.00414f
C4621 VDD.n2478 VSS 0.00758f
C4622 VDD.n2479 VSS 0.0039f
C4623 VDD.n2480 VSS 0.00461f
C4624 VDD.n2481 VSS 0.00391f
C4625 VDD.n2482 VSS 0.00184f
C4626 VDD.n2483 VSS 0.00135f
C4627 VDD.n2484 VSS 0.00256f
C4628 VDD.n2485 VSS 0.0203f
C4629 VDD.n2486 VSS 0.00163f
C4630 VDD.t58 VSS 0.274f
C4631 VDD.t37 VSS 0.479f
C4632 VDD.n2487 VSS 0.0695f
C4633 VDD.n2488 VSS 0.0813f
C4634 VDD.n2489 VSS 0.00839f
C4635 VDD.n2490 VSS 0.00634f
C4636 VDD.n2491 VSS 0.0109f
C4637 VDD.n2492 VSS 0.0457f
C4638 VDD.n2493 VSS 0.0199f
C4639 VDD.n2494 VSS 0.00839f
C4640 VDD.n2495 VSS 0.00634f
C4641 VDD.n2496 VSS 0.0081f
C4642 VDD.n2497 VSS 0.02f
C4643 VDD.n2498 VSS 0.0457f
C4644 VDD.n2499 VSS 0.0199f
C4645 VDD.n2500 VSS 0.00634f
C4646 VDD.n2501 VSS 0.00839f
C4647 VDD.n2502 VSS 0.0813f
C4648 VDD.n2503 VSS 0.0081f
C4649 VDD.n2504 VSS 0.02f
C4650 VDD.n2505 VSS 0.0458f
C4651 VDD.n2506 VSS 0.0199f
C4652 VDD.t30 VSS 0.00943f
C4653 VDD.n2507 VSS 0.136f
C4654 VDD.n2508 VSS 0.02f
C4655 VDD.n2509 VSS 0.0193f
C4656 VDD.n2510 VSS 0.0168f
C4657 VDD.n2511 VSS 0.00786f
C4658 VDD.n2512 VSS 0.0172f
C4659 VDD.n2513 VSS 0.00659f
C4660 VDD.t36 VSS 0.00663f
C4661 VDD.t33 VSS 0.00663f
C4662 VDD.n2514 VSS 0.0163f
C4663 VDD.n2515 VSS 0.0482f
C4664 VDD.n2516 VSS 0.00805f
C4665 VDD.n2517 VSS 0.0164f
C4666 VDD.n2518 VSS 0.097f
C4667 VDD.n2519 VSS 0.116f
C4668 VDD.n2520 VSS 0.0109f
C4669 VDD.n2521 VSS 0.161f
C4670 VDD.n2522 VSS 0.161f
C4671 VDD.n2523 VSS 0.0109f
C4672 VDD.n2524 VSS 0.0967f
C4673 VDD.n2525 VSS 0.0967f
C4674 VDD.n2526 VSS 0.0109f
C4675 VDD.n2527 VSS 0.107f
C4676 VDD.n2528 VSS 0.107f
C4677 VDD.n2529 VSS 0.0457f
C4678 VDD.n2530 VSS 0.0199f
C4679 VDD.n2531 VSS 0.0457f
C4680 VDD.n2532 VSS 0.0199f
C4681 VDD.n2533 VSS 0.00634f
C4682 VDD.n2534 VSS 0.00839f
C4683 VDD.n2535 VSS 0.0527f
C4684 VDD.n2536 VSS 0.00277f
C4685 VDD.n2537 VSS 0.0418f
C4686 VDD.n2538 VSS 0.018f
C4687 VDD.n2539 VSS 0.413f
C4688 VDD.t29 VSS 0.555f
C4689 VDD.t34 VSS 0.308f
C4690 VDD.n2540 VSS 0.132f
C4691 VDD.n2541 VSS 0.149f
C4692 VDD.n2542 VSS 0.0813f
C4693 VDD.n2543 VSS 0.0081f
C4694 VDD.n2544 VSS 0.02f
C4695 VDD.n2545 VSS 0.0109f
C4696 VDD.n2546 VSS 0.0868f
C4697 VDD.n2547 VSS 0.0868f
C4698 VDD.n2548 VSS 0.00634f
C4699 VDD.n2549 VSS 0.00839f
C4700 VDD.n2550 VSS 0.0813f
C4701 VDD.n2551 VSS 0.0081f
C4702 VDD.n2552 VSS 0.02f
C4703 VDD.n2553 VSS 0.0109f
C4704 VDD.n2554 VSS 0.0929f
C4705 VDD.n2555 VSS 0.0929f
C4706 VDD.n2556 VSS 0.0199f
C4707 VDD.n2557 VSS 0.0457f
C4708 VDD.n2558 VSS 0.02f
C4709 VDD.n2559 VSS 0.0081f
C4710 VDD.n2560 VSS 0.0813f
C4711 VDD.n2561 VSS 0.215f
C4712 VDD.n2562 VSS 0.0941f
C4713 VDD.n2563 VSS 0.167f
C4714 VDD.n2564 VSS 0.553f
C4715 VDD.n2565 VSS 0.0813f
C4716 VDD.n2566 VSS 0.0813f
C4717 VDD.n2567 VSS 0.00839f
C4718 VDD.n2568 VSS 0.00634f
C4719 VDD.n2569 VSS 0.0109f
C4720 VDD.n2570 VSS 0.06f
C4721 VDD.n2571 VSS 0.0199f
C4722 VDD.n2572 VSS 0.00839f
C4723 VDD.n2573 VSS 0.00634f
C4724 VDD.n2574 VSS 0.0081f
C4725 VDD.n2575 VSS 0.02f
C4726 VDD.n2576 VSS 0.06f
C4727 VDD.n2577 VSS 0.0199f
C4728 VDD.n2578 VSS 0.00839f
C4729 VDD.n2579 VSS 0.00634f
C4730 VDD.n2580 VSS 0.0081f
C4731 VDD.n2581 VSS 0.02f
C4732 VDD.n2582 VSS 0.0109f
C4733 VDD.n2583 VSS 0.166f
C4734 VDD.n2584 VSS 0.166f
C4735 VDD.n2585 VSS 0.0109f
C4736 VDD.n2586 VSS 0.145f
C4737 VDD.n2587 VSS 0.145f
C4738 VDD.n2588 VSS 0.122f
C4739 VDD.n2589 VSS 0.0199f
C4740 VDD.n2590 VSS 0.06f
C4741 VDD.n2591 VSS 0.02f
C4742 VDD.n2592 VSS 0.0081f
C4743 VDD.n2593 VSS 0.0813f
C4744 VDD.n2594 VSS 0.297f
C4745 VDD.n2595 VSS 0.033f
C4746 VDD.n2596 VSS 0.0209f
C4747 VDD.n2597 VSS 0.0394f
C4748 VDD.n2598 VSS 0.199f
C4749 VDD.n2599 VSS 0.0124f
C4750 VDD.n2600 VSS 0.0109f
C4751 VDD.n2601 VSS 0.00997f
C4752 VDD.n2602 VSS 0.0262f
C4753 VDD.n2603 VSS 0.0172f
C4754 VDD.n2604 VSS 0.0197f
C4755 VDD.n2605 VSS 8.15e-19
C4756 VDD.n2606 VSS 0.0124f
C4757 VDD.n2607 VSS 0.09f
C4758 VDD.n2608 VSS 0.004f
C4759 VDD.n2609 VSS 0.0124f
C4760 VDD.n2610 VSS 0.0111f
C4761 VDD.n2611 VSS 0.00571f
C4762 VDD.n2612 VSS 0.02f
C4763 VDD.n2613 VSS 0.0261f
C4764 VDD.n2614 VSS 0.0604f
C4765 VDD.n2615 VSS 0.0274f
C4766 VDD.n2616 VSS 0.0198f
C4767 VDD.n2617 VSS 0.0211f
C4768 VDD.n2618 VSS 0.0233f
C4769 VDD.n2619 VSS 0.056f
C4770 VDD.n2620 VSS 0.00797f
C4771 VDD.n2621 VSS 0.0313f
C4772 VDD.n2622 VSS 0.246f
C4773 VDD.t32 VSS 0.739f
C4774 VDD.t35 VSS 0.00583f
C4775 VDD.n2623 VSS 0.0362f
C4776 VDD.n2624 VSS 0.0574f
C4777 VDD.n2625 VSS 0.0639f
C4778 VDD.n2626 VSS 0.442f
C4779 VDD.n2627 VSS 0.102f
C4780 VDD.n2628 VSS 0.0527f
C4781 VDD.n2629 VSS 0.00277f
C4782 VDD.n2630 VSS 0.00302f
C4783 VDD.n2631 VSS 3.16e-19
C4784 VDD.n2632 VSS 0.00348f
C4785 VDD.n2633 VSS 4.74e-19
C4786 VDD.n2634 VSS 0.00348f
C4787 VDD.n2635 VSS 0.00269f
C4788 VDD.n2636 VSS 0.00332f
C4789 VDD.n2637 VSS 0.00979f
C4790 VDD.n2638 VSS 0.00979f
C4791 VDD.n2639 VSS 0.0129f
C4792 VDD.n2640 VSS 0.245f
C4793 VDD.n2641 VSS 0.0527f
C4794 VDD.n2642 VSS 0.198f
C4795 VDD.n2643 VSS 0.0104f
C4796 VDD.n2644 VSS 0.00979f
C4797 VDD.n2645 VSS 0.00269f
C4798 VDD.n2646 VSS 0.00916f
C4799 VDD.n2647 VSS 4.74e-19
C4800 VDD.n2648 VSS 0.00332f
C4801 VDD.n2649 VSS 0.00585f
C4802 VDD.n2650 VSS 0.00348f
C4803 VDD.n2651 VSS 4.74e-19
C4804 VDD.n2652 VSS 0.00472f
C4805 VDD.n2653 VSS 3.26e-19
C4806 VDD.n2654 VSS 0.0233f
C4807 VDD.n2655 VSS -0.0753f
C4808 VDD.n2656 VSS 0.0233f
C4809 VDD.n2657 VSS 0.014f
C4810 VDD.n2658 VSS 0.0145f
C4811 VDD.n2659 VSS 3.26e-19
C4812 VDD.n2660 VSS 0.00488f
C4813 VDD.n2661 VSS 0.00798f
C4814 VDD.n2662 VSS 0.00348f
C4815 VDD.n2663 VSS 0.00979f
C4816 VDD.n2664 VSS 0.00332f
C4817 VDD.n2665 VSS 0.00663f
C4818 VDD.n2666 VSS 0.00806f
C4819 VDD.n2667 VSS 0.00332f
C4820 VDD.n2668 VSS 0.00411f
C4821 VDD.n2669 VSS 0.00585f
C4822 VDD.n2670 VSS -0.211f
C4823 VDD.n2671 VSS 0.00374f
C4824 VDD.n2672 VSS 0.0229f
C4825 VDD.n2673 VSS 0.014f
C4826 VDD.n2674 VSS 0.0145f
C4827 VDD.n2675 VSS 3.26e-19
C4828 VDD.n2676 VSS 0.00488f
C4829 VDD.n2677 VSS 0.00798f
C4830 VDD.n2678 VSS 0.00374f
C4831 VDD.n2679 VSS 0.0229f
C4832 VDD.n2680 VSS 0.0229f
C4833 VDD.n2681 VSS 0.00488f
C4834 VDD.n2682 VSS 0.00439f
C4835 VDD.n2683 VSS 0.00806f
C4836 VDD.n2684 VSS 0.00332f
C4837 VDD.n2685 VSS 0.00663f
C4838 VDD.n2686 VSS 4.74e-19
C4839 VDD.n2687 VSS 0.00269f
C4840 VDD.n2688 VSS 0.00269f
C4841 VDD.n2689 VSS 0.00269f
C4842 VDD.n2690 VSS 0.00277f
C4843 VDD.n2691 VSS 0.0129f
C4844 VDD.n2692 VSS 0.198f
C4845 VDD.n2693 VSS 0.0104f
C4846 VDD.n2694 VSS 0.00979f
C4847 VDD.n2695 VSS 0.00979f
C4848 VDD.n2696 VSS 0.0129f
C4849 VDD.n2697 VSS 0.245f
C4850 VDD.n2698 VSS 0.0527f
C4851 VDD.n2699 VSS 0.00277f
C4852 VDD.n2700 VSS 0.00269f
C4853 VDD.n2701 VSS 3.16e-19
C4854 VDD.n2702 VSS 0.00269f
C4855 VDD.n2703 VSS 0.00348f
C4856 VDD.n2704 VSS 0.00269f
C4857 VDD.n2705 VSS 0.00332f
C4858 VDD.n2706 VSS 0.00979f
C4859 VDD.n2707 VSS 0.00979f
C4860 VDD.n2708 VSS 0.0129f
C4861 VDD.n2709 VSS 0.245f
C4862 VDD.n2710 VSS 0.0527f
C4863 VDD.n2711 VSS 0.124f
C4864 VDD.n2712 VSS 0.0236f
C4865 VDD.n2713 VSS 0.00979f
C4866 VDD.n2714 VSS 0.0095f
C4867 VDD.n2715 VSS 0.00332f
C4868 VDD.n2716 VSS 3.26e-19
C4869 VDD.n2717 VSS 0.0229f
C4870 VDD.n2718 VSS 0.00488f
C4871 VDD.n2719 VSS 0.014f
C4872 VDD.n2720 VSS 3.26e-19
C4873 VDD.n2721 VSS 0.0145f
C4874 VDD.n2722 VSS 0.0233f
C4875 VDD.n2723 VSS 0.00798f
C4876 VDD.n2724 VSS 0.00374f
C4877 VDD.n2725 VSS 0.00348f
C4878 VDD.n2726 VSS 0.00979f
C4879 VDD.n2727 VSS 0.00332f
C4880 VDD.n2728 VSS 0.00663f
C4881 VDD.n2729 VSS 0.00806f
C4882 VDD.n2730 VSS 0.00411f
C4883 VDD.n2731 VSS 0.00585f
C4884 VDD.n2732 VSS -0.211f
C4885 VDD.n2733 VSS -0.0753f
C4886 VDD.n2734 VSS 0.014f
C4887 VDD.n2735 VSS 0.0145f
C4888 VDD.n2736 VSS 0.0138f
C4889 VDD.n2737 VSS 0.00439f
C4890 VDD.n2738 VSS 0.00332f
C4891 VDD.n2739 VSS 0.0418f
C4892 VDD.n2740 VSS 0.00269f
C4893 VDD.n2741 VSS 0.00348f
C4894 VDD.n2742 VSS 3.26e-19
C4895 VDD.n2743 VSS 0.00374f
C4896 VDD.n2744 VSS -0.0844f
C4897 VDD.n2745 VSS 0.0142f
C4898 VDD.n2746 VSS 0.00472f
C4899 VDD.n2747 VSS 3.26e-19
C4900 VDD.n2748 VSS 0.00411f
C4901 VDD.n2749 VSS 0.00348f
C4902 VDD.n2750 VSS 0.00488f
C4903 VDD.n2751 VSS 0.00916f
C4904 VDD.n2752 VSS 0.00269f
C4905 VDD.n2753 VSS 0.00269f
C4906 VDD.n2754 VSS 0.00269f
C4907 VDD.n2755 VSS 0.00277f
C4908 VDD.n2756 VSS 0.0129f
C4909 VDD.n2757 VSS 0.198f
C4910 VDD.n2758 VSS 0.018f
C4911 VDD.t56 VSS 0.49f
C4912 VDD.n2759 VSS 0.605f
C4913 VDD.n2760 VSS 0.0527f
C4914 VDD.n2761 VSS 0.00277f
C4915 VDD.n2762 VSS 0.0104f
C4916 VDD.n2763 VSS 0.00269f
C4917 VDD.n2764 VSS 0.00585f
C4918 VDD.n2765 VSS 0.00806f
C4919 VDD.n2766 VSS 0.00663f
C4920 VDD.n2767 VSS 0.00332f
C4921 VDD.n2768 VSS 0.00979f
C4922 VDD.n2769 VSS 0.00979f
C4923 VDD.n2770 VSS 0.0129f
C4924 VDD.n2771 VSS 0.245f
C4925 VDD.n2772 VSS 0.0527f
C4926 VDD.n2773 VSS 0.198f
C4927 VDD.n2774 VSS 0.0104f
C4928 VDD.n2775 VSS 0.00979f
C4929 VDD.n2776 VSS 0.00269f
C4930 VDD.n2777 VSS 0.00916f
C4931 VDD.n2778 VSS 4.74e-19
C4932 VDD.n2779 VSS 0.00332f
C4933 VDD.n2780 VSS 0.00585f
C4934 VDD.n2781 VSS 0.00348f
C4935 VDD.n2782 VSS 4.74e-19
C4936 VDD.n2783 VSS 0.00472f
C4937 VDD.n2784 VSS 3.26e-19
C4938 VDD.n2785 VSS 0.023f
C4939 VDD.n2786 VSS -0.0753f
C4940 VDD.n2787 VSS 0.023f
C4941 VDD.n2788 VSS 0.00798f
C4942 VDD.n2789 VSS 0.00979f
C4943 VDD.n2790 VSS 0.00332f
C4944 VDD.n2791 VSS 0.00663f
C4945 VDD.n2792 VSS 0.00806f
C4946 VDD.n2793 VSS 0.00332f
C4947 VDD.n2794 VSS 0.00411f
C4948 VDD.n2795 VSS 0.00585f
C4949 VDD.n2796 VSS -0.211f
C4950 VDD.n2797 VSS 0.00374f
C4951 VDD.n2798 VSS 0.0225f
C4952 VDD.n2799 VSS 0.0138f
C4953 VDD.n2800 VSS 0.0142f
C4954 VDD.n2801 VSS 3.26e-19
C4955 VDD.n2802 VSS 0.00488f
C4956 VDD.n2803 VSS 0.00798f
C4957 VDD.n2804 VSS 0.00374f
C4958 VDD.n2805 VSS 0.0225f
C4959 VDD.n2806 VSS 0.0225f
C4960 VDD.n2807 VSS 0.00488f
C4961 VDD.n2808 VSS 0.00439f
C4962 VDD.n2809 VSS 0.00806f
C4963 VDD.n2810 VSS 0.00332f
C4964 VDD.n2811 VSS 0.00663f
C4965 VDD.n2812 VSS 4.74e-19
C4966 VDD.n2813 VSS 0.00269f
C4967 VDD.n2814 VSS 0.00269f
C4968 VDD.n2815 VSS 0.00269f
C4969 VDD.n2816 VSS 0.00277f
C4970 VDD.n2817 VSS 0.0129f
C4971 VDD.n2818 VSS 0.198f
C4972 VDD.n2819 VSS 0.0104f
C4973 VDD.n2820 VSS 0.00979f
C4974 VDD.n2821 VSS 0.00979f
C4975 VDD.n2822 VSS 0.0129f
C4976 VDD.n2823 VSS 0.245f
C4977 VDD.n2824 VSS 0.0527f
C4978 VDD.n2825 VSS 0.00277f
C4979 VDD.n2826 VSS 0.00269f
C4980 VDD.n2827 VSS 3.16e-19
C4981 VDD.n2828 VSS 0.00269f
C4982 VDD.n2829 VSS 0.00348f
C4983 VDD.n2830 VSS 0.00269f
C4984 VDD.n2831 VSS 0.00332f
C4985 VDD.n2832 VSS 0.00979f
C4986 VDD.n2833 VSS 0.00979f
C4987 VDD.n2834 VSS 0.0129f
C4988 VDD.n2835 VSS 0.245f
C4989 VDD.n2836 VSS 0.0527f
C4990 VDD.n2837 VSS 0.124f
C4991 VDD.n2838 VSS 0.0236f
C4992 VDD.n2839 VSS 0.00979f
C4993 VDD.n2840 VSS 0.00269f
C4994 VDD.n2841 VSS 0.00916f
C4995 VDD.n2842 VSS 4.74e-19
C4996 VDD.n2843 VSS 0.00332f
C4997 VDD.n2844 VSS 0.0286f
C4998 VDD.n2845 VSS 0.00269f
C4999 VDD.n2846 VSS 0.0294f
C5000 VDD.n2847 VSS 0.00269f
C5001 VDD.n2848 VSS 0.00348f
C5002 VDD.n2849 VSS 0.00277f
C5003 VDD.t41 VSS 0.47f
C5004 VDD.n2850 VSS 0.207f
C5005 VDD.t68 VSS 0.253f
C5006 VDD.n2851 VSS 0.198f
C5007 VDD.n2852 VSS 0.0104f
C5008 VDD.n2853 VSS 0.00269f
C5009 VDD.n2854 VSS 0.00663f
C5010 VDD.n2855 VSS 0.00348f
C5011 VDD.n2856 VSS 0.00806f
C5012 VDD.n2857 VSS 0.00472f
C5013 VDD.n2858 VSS 0.00411f
C5014 VDD.n2859 VSS 3.26e-19
C5015 VDD.n2860 VSS 0.00488f
C5016 VDD.n2861 VSS 0.023f
C5017 VDD.n2862 VSS -0.0753f
C5018 VDD.n2863 VSS 0.00348f
C5019 VDD.n2864 VSS 0.0285f
C5020 VDD.n2865 VSS 0.0142f
C5021 VDD.n2866 VSS -0.211f
C5022 VDD.n2867 VSS 0.023f
C5023 VDD.n2868 VSS 0.0138f
C5024 VDD.n2869 VSS 0.0142f
C5025 VDD.n2870 VSS 3.26e-19
C5026 VDD.n2871 VSS 0.00488f
C5027 VDD.n2872 VSS 0.00798f
C5028 VDD.n2873 VSS 0.00374f
C5029 VDD.n2874 VSS 0.0225f
C5030 VDD.n2875 VSS 0.0138f
C5031 VDD.n2876 VSS 0.00348f
C5032 VDD.n2877 VSS 0.00979f
C5033 VDD.n2878 VSS 0.00332f
C5034 VDD.n2879 VSS 0.00663f
C5035 VDD.n2880 VSS 0.00806f
C5036 VDD.n2881 VSS 0.00585f
C5037 VDD.n2882 VSS 0.00411f
C5038 VDD.n2883 VSS 0.00332f
C5039 VDD.n2884 VSS -0.0753f
C5040 VDD.n2885 VSS 3.26e-19
C5041 VDD.n2886 VSS 0.00488f
C5042 VDD.n2887 VSS 0.0286f
C5043 VDD.n2888 VSS 0.0813f
C5044 VDD.n2889 VSS 0.0809f
C5045 VDD.n2890 VSS 0.0142f
C5046 VDD.n2891 VSS 0.0138f
C5047 VDD.n2892 VSS 3.26e-19
C5048 VDD.n2893 VSS 0.00472f
C5049 VDD.n2894 VSS 4.74e-19
C5050 VDD.n2895 VSS 0.00332f
C5051 VDD.n2896 VSS 0.00916f
C5052 VDD.n2897 VSS 0.00411f
C5053 VDD.n2898 VSS 0.00585f
C5054 VDD.n2899 VSS -0.211f
C5055 VDD.n2900 VSS 0.00391f
C5056 VDD.n2901 VSS 0.00781f
C5057 VDD.n2902 VSS 0.0225f
C5058 VDD.n2903 VSS 0.0138f
C5059 VDD.n2904 VSS -0.182f
C5060 VDD.n2905 VSS 3.26e-19
C5061 VDD.n2906 VSS 0.00348f
C5062 VDD.n2907 VSS 0.00332f
C5063 VDD.n2908 VSS 0.00269f
C5064 VDD.n2909 VSS 0.00916f
C5065 VDD.n2910 VSS 0.00269f
C5066 VDD.n2911 VSS 0.00269f
C5067 VDD.n2912 VSS 0.0129f
C5068 VDD.n2913 VSS 0.00277f
C5069 VDD.n2914 VSS 3.16e-19
C5070 VDD.n2915 VSS 0.00916f
C5071 VDD.n2916 VSS 0.00585f
C5072 VDD.n2917 VSS 0.00806f
C5073 VDD.n2918 VSS 0.00663f
C5074 VDD.n2919 VSS 0.00332f
C5075 VDD.n2920 VSS 0.00979f
C5076 VDD.n2921 VSS 0.00979f
C5077 VDD.n2922 VSS 0.00269f
C5078 VDD.n2923 VSS 0.00277f
C5079 VDD.n2924 VSS 0.0527f
C5080 VDD.n2925 VSS 0.245f
C5081 VDD.n2926 VSS 0.198f
C5082 VDD.n2927 VSS 0.0104f
C5083 VDD.n2928 VSS 0.00269f
C5084 VDD.n2929 VSS 0.00663f
C5085 VDD.n2930 VSS 0.00348f
C5086 VDD.n2931 VSS 0.00806f
C5087 VDD.n2932 VSS 0.00472f
C5088 VDD.n2933 VSS 0.00411f
C5089 VDD.n2934 VSS 3.26e-19
C5090 VDD.n2935 VSS -0.211f
C5091 VDD.n2936 VSS 0.023f
C5092 VDD.n2937 VSS -0.078f
C5093 VDD.n2938 VSS 0.0142f
C5094 VDD.n2939 VSS 0.00439f
C5095 VDD.n2940 VSS 0.00411f
C5096 VDD.n2941 VSS 0.00585f
C5097 VDD.n2942 VSS 0.00488f
C5098 VDD.n2943 VSS 0.00391f
C5099 VDD.n2944 VSS 0.00781f
C5100 VDD.n2945 VSS 0.0225f
C5101 VDD.n2946 VSS 0.0138f
C5102 VDD.n2947 VSS 0.0225f
C5103 VDD.n2948 VSS 3.26e-19
C5104 VDD.n2949 VSS 0.00348f
C5105 VDD.n2950 VSS 0.00332f
C5106 VDD.n2951 VSS 0.00269f
C5107 VDD.n2952 VSS 0.00916f
C5108 VDD.n2953 VSS 0.00269f
C5109 VDD.n2954 VSS 0.00269f
C5110 VDD.n2955 VSS 0.0129f
C5111 VDD.n2956 VSS 0.00277f
C5112 VDD.n2957 VSS 3.16e-19
C5113 VDD.n2958 VSS 0.00916f
C5114 VDD.n2959 VSS 0.00585f
C5115 VDD.n2960 VSS 0.00806f
C5116 VDD.n2961 VSS 0.00663f
C5117 VDD.n2962 VSS 0.00332f
C5118 VDD.n2963 VSS 0.00979f
C5119 VDD.n2964 VSS 0.00979f
C5120 VDD.n2965 VSS 0.00269f
C5121 VDD.n2966 VSS 0.00277f
C5122 VDD.n2967 VSS 0.0527f
C5123 VDD.n2968 VSS 0.245f
C5124 VDD.n2969 VSS 0.198f
C5125 VDD.n2970 VSS 0.0104f
C5126 VDD.n2971 VSS 0.00269f
C5127 VDD.n2972 VSS 0.00663f
C5128 VDD.n2973 VSS 0.00348f
C5129 VDD.n2974 VSS 0.00806f
C5130 VDD.n2975 VSS 0.00332f
C5131 VDD.n2976 VSS 0.00781f
C5132 VDD.n2977 VSS 0.00439f
C5133 VDD.n2978 VSS 0.0138f
C5134 VDD.n2979 VSS 0.0142f
C5135 VDD.n2980 VSS 0.00439f
C5136 VDD.n2981 VSS 0.00411f
C5137 VDD.n2982 VSS 0.00585f
C5138 VDD.n2983 VSS 0.00488f
C5139 VDD.n2984 VSS 0.00391f
C5140 VDD.n2985 VSS 0.023f
C5141 VDD.n2986 VSS -0.182f
C5142 VDD.n2987 VSS 0.00488f
C5143 VDD.n2988 VSS 0.00472f
C5144 VDD.n2989 VSS -0.0844f
C5145 VDD.n2990 VSS 3.26e-19
C5146 VDD.n2991 VSS 0.00411f
C5147 VDD.n2992 VSS 0.00488f
C5148 VDD.n2993 VSS 0.00348f
C5149 VDD.n2994 VSS 0.0251f
C5150 VDD.n2995 VSS 0.0251f
C5151 VDD.n2996 VSS 0.00411f
C5152 VDD.n2997 VSS 0.0295f
C5153 VDD.n2998 VSS 0.0295f
C5154 VDD.n2999 VSS 0.00269f
C5155 VDD.n3000 VSS 0.00269f
C5156 VDD.n3001 VSS 0.00269f
C5157 VDD.n3002 VSS 0.00277f
C5158 VDD.n3003 VSS 0.0129f
C5159 VDD.n3004 VSS 3.16e-19
C5160 VDD.n3005 VSS 0.00269f
C5161 VDD.n3006 VSS 0.00277f
C5162 VDD.n3007 VSS 0.0527f
C5163 VDD.n3008 VSS 0.412f
C5164 VDD.n3009 VSS 0.0186f
C5165 VDD.n3010 VSS 0.03f
C5166 VDD.n3011 VSS 0.03f
C5167 VDD.n3012 VSS 0.0186f
C5168 VDD.n3013 VSS 0.226f
C5169 VDD.n3014 VSS 0.0527f
C5170 VDD.n3015 VSS 0.198f
C5171 VDD.n3016 VSS 0.0104f
C5172 VDD.n3017 VSS 0.00979f
C5173 VDD.n3018 VSS 0.00269f
C5174 VDD.n3019 VSS 0.00916f
C5175 VDD.n3020 VSS 4.74e-19
C5176 VDD.n3021 VSS 0.00332f
C5177 VDD.n3022 VSS 0.00585f
C5178 VDD.n3023 VSS 0.00348f
C5179 VDD.n3024 VSS 4.74e-19
C5180 VDD.n3025 VSS -0.211f
C5181 VDD.n3026 VSS 3.26e-19
C5182 VDD.n3027 VSS 0.023f
C5183 VDD.n3028 VSS 0.00439f
C5184 VDD.n3029 VSS -0.174f
C5185 VDD.n3030 VSS 0.00798f
C5186 VDD.n3031 VSS 0.00979f
C5187 VDD.n3032 VSS 0.00332f
C5188 VDD.n3033 VSS 0.00663f
C5189 VDD.n3034 VSS 0.00806f
C5190 VDD.n3035 VSS 0.00332f
C5191 VDD.n3036 VSS 0.00411f
C5192 VDD.n3037 VSS 0.00585f
C5193 VDD.n3038 VSS 0.00472f
C5194 VDD.n3039 VSS 0.00374f
C5195 VDD.n3040 VSS 0.0225f
C5196 VDD.n3041 VSS 0.0138f
C5197 VDD.n3042 VSS 0.0142f
C5198 VDD.n3043 VSS 3.26e-19
C5199 VDD.n3044 VSS 0.00488f
C5200 VDD.n3045 VSS 0.00798f
C5201 VDD.n3046 VSS 0.00374f
C5202 VDD.n3047 VSS 0.0225f
C5203 VDD.n3048 VSS 0.0225f
C5204 VDD.n3049 VSS 0.00488f
C5205 VDD.n3050 VSS 0.00439f
C5206 VDD.n3051 VSS 0.00806f
C5207 VDD.n3052 VSS 0.00332f
C5208 VDD.n3053 VSS 0.00663f
C5209 VDD.n3054 VSS 4.74e-19
C5210 VDD.n3055 VSS 0.00269f
C5211 VDD.n3056 VSS 0.00269f
C5212 VDD.n3057 VSS 0.00269f
C5213 VDD.n3058 VSS 0.00277f
C5214 VDD.n3059 VSS 0.0129f
C5215 VDD.n3060 VSS 0.198f
C5216 VDD.n3061 VSS 0.0104f
C5217 VDD.n3062 VSS 0.00979f
C5218 VDD.n3063 VSS 0.00979f
C5219 VDD.n3064 VSS 0.0129f
C5220 VDD.n3065 VSS 0.245f
C5221 VDD.n3066 VSS 0.0527f
C5222 VDD.n3067 VSS 0.00277f
C5223 VDD.n3068 VSS 0.00269f
C5224 VDD.n3069 VSS 3.16e-19
C5225 VDD.n3070 VSS 0.00269f
C5226 VDD.n3071 VSS 0.00348f
C5227 VDD.n3072 VSS 0.00269f
C5228 VDD.n3073 VSS 0.00332f
C5229 VDD.n3074 VSS 0.00979f
C5230 VDD.n3075 VSS 0.00979f
C5231 VDD.n3076 VSS 0.0129f
C5232 VDD.n3077 VSS 0.245f
C5233 VDD.n3078 VSS 0.0527f
C5234 VDD.n3079 VSS 0.198f
C5235 VDD.n3080 VSS 0.0104f
C5236 VDD.n3081 VSS 0.00979f
C5237 VDD.n3082 VSS 0.00269f
C5238 VDD.n3083 VSS 0.00916f
C5239 VDD.n3084 VSS 4.74e-19
C5240 VDD.n3085 VSS 0.00332f
C5241 VDD.n3086 VSS 0.00585f
C5242 VDD.n3087 VSS 0.00348f
C5243 VDD.n3088 VSS 4.74e-19
C5244 VDD.n3089 VSS -0.211f
C5245 VDD.n3090 VSS 3.26e-19
C5246 VDD.n3091 VSS 0.023f
C5247 VDD.n3092 VSS 0.00439f
C5248 VDD.n3093 VSS -0.174f
C5249 VDD.n3094 VSS 0.0138f
C5250 VDD.n3095 VSS -0.0844f
C5251 VDD.n3096 VSS 3.26e-19
C5252 VDD.n3097 VSS 0.00488f
C5253 VDD.n3098 VSS 0.00798f
C5254 VDD.n3099 VSS 0.00348f
C5255 VDD.n3100 VSS 0.00979f
C5256 VDD.n3101 VSS 0.00332f
C5257 VDD.n3102 VSS 0.00663f
C5258 VDD.n3103 VSS 0.00806f
C5259 VDD.n3104 VSS 0.00332f
C5260 VDD.n3105 VSS 0.00411f
C5261 VDD.n3106 VSS 0.00585f
C5262 VDD.n3107 VSS 0.00472f
C5263 VDD.n3108 VSS 0.00374f
C5264 VDD.n3109 VSS 0.0225f
C5265 VDD.n3110 VSS 0.0138f
C5266 VDD.n3111 VSS 0.0142f
C5267 VDD.n3112 VSS 3.26e-19
C5268 VDD.n3113 VSS 0.00488f
C5269 VDD.n3114 VSS 0.00798f
C5270 VDD.n3115 VSS 0.00374f
C5271 VDD.n3116 VSS 0.0225f
C5272 VDD.n3117 VSS 0.0809f
C5273 VDD.n3118 VSS 0.00488f
C5274 VDD.n3119 VSS 3.26e-19
C5275 VDD.n3120 VSS 0.00348f
C5276 VDD.n3121 VSS 0.00332f
C5277 VDD.n3122 VSS 0.00269f
C5278 VDD.n3123 VSS 0.00916f
C5279 VDD.n3124 VSS 0.00269f
C5280 VDD.n3125 VSS 0.00269f
C5281 VDD.n3126 VSS 0.00277f
C5282 VDD.n3127 VSS 0.0527f
C5283 VDD.n3128 VSS 0.00277f
C5284 VDD.n3129 VSS 0.00979f
C5285 VDD.n3130 VSS 0.245f
C5286 VDD.n3131 VSS 0.0129f
C5287 VDD.n3132 VSS 0.00979f
C5288 VDD.n3133 VSS 0.00269f
C5289 VDD.n3134 VSS 0.0294f
C5290 VDD.n3135 VSS 0.00332f
C5291 VDD.n3136 VSS 0.0286f
C5292 VDD.n3137 VSS 0.0294f
C5293 VDD.n3138 VSS 0.00332f
C5294 VDD.n3139 VSS 0.0261f
C5295 VDD.n3140 VSS 0.0261f
C5296 VDD.n3141 VSS 0.0286f
C5297 VDD.n3142 VSS 0.00348f
C5298 VDD.n3143 VSS 0.00269f
C5299 VDD.n3144 VSS 0.00269f
C5300 VDD.n3145 VSS 3.16e-19
C5301 VDD.n3146 VSS 0.0236f
C5302 VDD.n3147 VSS 0.124f
C5303 VDD.t64 VSS 0.47f
C5304 VDD.n3148 VSS 0.207f
C5305 VDD.t74 VSS 0.253f
C5306 VDD.n3149 VSS 0.198f
C5307 VDD.n3150 VSS 0.0104f
C5308 VDD.n3151 VSS 0.00269f
C5309 VDD.n3152 VSS 0.00663f
C5310 VDD.n3153 VSS 0.00348f
C5311 VDD.n3154 VSS 0.00806f
C5312 VDD.n3155 VSS 0.00472f
C5313 VDD.n3156 VSS 0.00411f
C5314 VDD.n3157 VSS 3.26e-19
C5315 VDD.n3158 VSS 0.00488f
C5316 VDD.n3159 VSS 0.023f
C5317 VDD.n3160 VSS 0.0138f
C5318 VDD.n3161 VSS 0.0142f
C5319 VDD.n3162 VSS -0.0753f
C5320 VDD.n3163 VSS 0.00411f
C5321 VDD.n3164 VSS 0.00585f
C5322 VDD.n3165 VSS -0.211f
C5323 VDD.n3166 VSS 0.00391f
C5324 VDD.n3167 VSS 0.00781f
C5325 VDD.n3168 VSS 0.0225f
C5326 VDD.n3169 VSS 0.0138f
C5327 VDD.n3170 VSS -0.182f
C5328 VDD.n3171 VSS 3.26e-19
C5329 VDD.n3172 VSS 0.00348f
C5330 VDD.n3173 VSS 0.00332f
C5331 VDD.n3174 VSS 0.00269f
C5332 VDD.n3175 VSS 0.00916f
C5333 VDD.n3176 VSS 0.00269f
C5334 VDD.n3177 VSS 0.00269f
C5335 VDD.n3178 VSS 0.0129f
C5336 VDD.n3179 VSS 0.00277f
C5337 VDD.n3180 VSS 3.16e-19
C5338 VDD.n3181 VSS 0.00916f
C5339 VDD.n3182 VSS 0.00585f
C5340 VDD.n3183 VSS 0.00806f
C5341 VDD.n3184 VSS 0.00663f
C5342 VDD.n3185 VSS 0.00332f
C5343 VDD.n3186 VSS 0.00979f
C5344 VDD.n3187 VSS 0.00979f
C5345 VDD.n3188 VSS 0.00269f
C5346 VDD.n3189 VSS 0.00277f
C5347 VDD.n3190 VSS 0.0527f
C5348 VDD.n3191 VSS 0.245f
C5349 VDD.n3192 VSS 0.198f
C5350 VDD.n3193 VSS 0.0104f
C5351 VDD.n3194 VSS 0.00269f
C5352 VDD.n3195 VSS 0.00663f
C5353 VDD.n3196 VSS 0.00348f
C5354 VDD.n3197 VSS 0.00806f
C5355 VDD.n3198 VSS 0.00472f
C5356 VDD.n3199 VSS 0.00411f
C5357 VDD.n3200 VSS 3.26e-19
C5358 VDD.n3201 VSS -0.211f
C5359 VDD.n3202 VSS 0.023f
C5360 VDD.n3203 VSS -0.078f
C5361 VDD.n3204 VSS 0.0142f
C5362 VDD.n3205 VSS 0.00439f
C5363 VDD.n3206 VSS 0.00411f
C5364 VDD.n3207 VSS 0.00585f
C5365 VDD.n3208 VSS 0.00488f
C5366 VDD.n3209 VSS 0.00391f
C5367 VDD.n3210 VSS 0.00781f
C5368 VDD.n3211 VSS 0.0225f
C5369 VDD.n3212 VSS 0.0138f
C5370 VDD.n3213 VSS 0.0225f
C5371 VDD.n3214 VSS 3.26e-19
C5372 VDD.n3215 VSS 0.00348f
C5373 VDD.n3216 VSS 0.00332f
C5374 VDD.n3217 VSS 0.00269f
C5375 VDD.n3218 VSS 0.00916f
C5376 VDD.n3219 VSS 0.00269f
C5377 VDD.n3220 VSS 0.00269f
C5378 VDD.n3221 VSS 0.0129f
C5379 VDD.n3222 VSS 0.00277f
C5380 VDD.n3223 VSS 3.16e-19
C5381 VDD.n3224 VSS 0.00916f
C5382 VDD.n3225 VSS 0.00585f
C5383 VDD.n3226 VSS 0.00806f
C5384 VDD.n3227 VSS 0.00663f
C5385 VDD.n3228 VSS 0.00332f
C5386 VDD.n3229 VSS 0.00979f
C5387 VDD.n3230 VSS 0.00979f
C5388 VDD.n3231 VSS 0.00269f
C5389 VDD.n3232 VSS 0.00277f
C5390 VDD.n3233 VSS 0.0527f
C5391 VDD.n3234 VSS 0.245f
C5392 VDD.n3235 VSS 0.198f
C5393 VDD.n3236 VSS 0.0104f
C5394 VDD.n3237 VSS 0.00269f
C5395 VDD.n3238 VSS 0.00663f
C5396 VDD.n3239 VSS 0.00348f
C5397 VDD.n3240 VSS 0.00806f
C5398 VDD.n3241 VSS 0.00332f
C5399 VDD.n3242 VSS 0.00781f
C5400 VDD.n3243 VSS 0.00439f
C5401 VDD.n3244 VSS 0.0138f
C5402 VDD.n3245 VSS 0.0142f
C5403 VDD.n3246 VSS 0.00439f
C5404 VDD.n3247 VSS 0.00411f
C5405 VDD.n3248 VSS 0.00585f
C5406 VDD.n3249 VSS 0.00488f
C5407 VDD.n3250 VSS 0.00391f
C5408 VDD.n3251 VSS 0.023f
C5409 VDD.n3252 VSS -0.182f
C5410 VDD.n3253 VSS 0.00488f
C5411 VDD.n3254 VSS 0.00472f
C5412 VDD.n3255 VSS -0.0844f
C5413 VDD.n3256 VSS 3.26e-19
C5414 VDD.n3257 VSS 0.00411f
C5415 VDD.n3258 VSS 0.00488f
C5416 VDD.n3259 VSS 0.00348f
C5417 VDD.n3260 VSS 0.0251f
C5418 VDD.n3261 VSS 0.0251f
C5419 VDD.n3262 VSS 0.00411f
C5420 VDD.n3263 VSS 0.0295f
C5421 VDD.n3264 VSS 0.0295f
C5422 VDD.n3265 VSS 0.00269f
C5423 VDD.n3266 VSS 0.00269f
C5424 VDD.n3267 VSS 0.00269f
C5425 VDD.n3268 VSS 0.00277f
C5426 VDD.n3269 VSS 0.0129f
C5427 VDD.n3270 VSS 3.16e-19
C5428 VDD.n3271 VSS 0.00269f
C5429 VDD.n3272 VSS 0.00277f
C5430 VDD.n3273 VSS 0.0527f
C5431 VDD.n3274 VSS 0.412f
C5432 VDD.n3275 VSS 0.0186f
C5433 VDD.n3276 VSS 0.03f
C5434 VDD.n3277 VSS 0.03f
C5435 VDD.n3278 VSS 0.0186f
C5436 VDD.n3279 VSS 0.226f
C5437 VDD.n3280 VSS 0.0527f
C5438 VDD.n3281 VSS 0.198f
C5439 VDD.n3282 VSS 0.0104f
C5440 VDD.n3283 VSS 0.00979f
C5441 VDD.n3284 VSS 0.00269f
C5442 VDD.n3285 VSS 0.00916f
C5443 VDD.n3286 VSS 4.74e-19
C5444 VDD.n3287 VSS 0.00332f
C5445 VDD.n3288 VSS 0.00585f
C5446 VDD.n3289 VSS 0.00348f
C5447 VDD.n3290 VSS 4.74e-19
C5448 VDD.n3291 VSS -0.211f
C5449 VDD.n3292 VSS 3.26e-19
C5450 VDD.n3293 VSS 0.023f
C5451 VDD.n3294 VSS 0.00439f
C5452 VDD.n3295 VSS -0.174f
C5453 VDD.n3296 VSS 0.00798f
C5454 VDD.n3297 VSS 0.00979f
C5455 VDD.n3298 VSS 0.00332f
C5456 VDD.n3299 VSS 0.00663f
C5457 VDD.n3300 VSS 0.00806f
C5458 VDD.n3301 VSS 0.00332f
C5459 VDD.n3302 VSS 0.00411f
C5460 VDD.n3303 VSS 0.00585f
C5461 VDD.n3304 VSS 0.00472f
C5462 VDD.n3305 VSS 0.00374f
C5463 VDD.n3306 VSS 0.0225f
C5464 VDD.n3307 VSS 0.0138f
C5465 VDD.n3308 VSS 0.0142f
C5466 VDD.n3309 VSS 3.26e-19
C5467 VDD.n3310 VSS 0.00488f
C5468 VDD.n3311 VSS 0.00798f
C5469 VDD.n3312 VSS 0.00374f
C5470 VDD.n3313 VSS 0.0225f
C5471 VDD.n3314 VSS 0.0225f
C5472 VDD.n3315 VSS 0.00488f
C5473 VDD.n3316 VSS 0.00439f
C5474 VDD.n3317 VSS 0.00806f
C5475 VDD.n3318 VSS 0.00332f
C5476 VDD.n3319 VSS 0.00663f
C5477 VDD.n3320 VSS 4.74e-19
C5478 VDD.n3321 VSS 0.00269f
C5479 VDD.n3322 VSS 0.00269f
C5480 VDD.n3323 VSS 0.00269f
C5481 VDD.n3324 VSS 0.00277f
C5482 VDD.n3325 VSS 0.0129f
C5483 VDD.n3326 VSS 0.198f
C5484 VDD.n3327 VSS 0.0104f
C5485 VDD.n3328 VSS 0.00979f
C5486 VDD.n3329 VSS 0.00979f
C5487 VDD.n3330 VSS 0.0129f
C5488 VDD.n3331 VSS 0.245f
C5489 VDD.n3332 VSS 0.0527f
C5490 VDD.n3333 VSS 0.00277f
C5491 VDD.n3334 VSS 0.00269f
C5492 VDD.n3335 VSS 3.16e-19
C5493 VDD.n3336 VSS 0.00269f
C5494 VDD.n3337 VSS 0.00348f
C5495 VDD.n3338 VSS 0.00269f
C5496 VDD.n3339 VSS 0.00332f
C5497 VDD.n3340 VSS 0.00979f
C5498 VDD.n3341 VSS 0.00979f
C5499 VDD.n3342 VSS 0.0129f
C5500 VDD.n3343 VSS 0.245f
C5501 VDD.n3344 VSS 0.0527f
C5502 VDD.n3345 VSS 0.198f
C5503 VDD.n3346 VSS 0.0104f
C5504 VDD.n3347 VSS 0.00979f
C5505 VDD.n3348 VSS 0.00269f
C5506 VDD.n3349 VSS 0.00916f
C5507 VDD.n3350 VSS 4.74e-19
C5508 VDD.n3351 VSS 0.00332f
C5509 VDD.n3352 VSS 0.00585f
C5510 VDD.n3353 VSS 0.00348f
C5511 VDD.n3354 VSS 4.74e-19
C5512 VDD.n3355 VSS -0.211f
C5513 VDD.n3356 VSS 3.26e-19
C5514 VDD.n3357 VSS 0.023f
C5515 VDD.n3358 VSS 0.00439f
C5516 VDD.n3359 VSS -0.174f
C5517 VDD.n3360 VSS 0.0138f
C5518 VDD.n3361 VSS -0.0844f
C5519 VDD.n3362 VSS 3.26e-19
C5520 VDD.n3363 VSS 0.00488f
C5521 VDD.n3364 VSS 0.00798f
C5522 VDD.n3365 VSS 0.00348f
C5523 VDD.n3366 VSS 0.00979f
C5524 VDD.n3367 VSS 0.00332f
C5525 VDD.n3368 VSS 0.00663f
C5526 VDD.n3369 VSS 0.00806f
C5527 VDD.n3370 VSS 0.00332f
C5528 VDD.n3371 VSS 0.00411f
C5529 VDD.n3372 VSS 0.00585f
C5530 VDD.n3373 VSS 0.00472f
C5531 VDD.n3374 VSS 0.00374f
C5532 VDD.n3375 VSS 0.0225f
C5533 VDD.n3376 VSS 0.0138f
C5534 VDD.n3377 VSS 0.0142f
C5535 VDD.n3378 VSS 3.26e-19
C5536 VDD.n3379 VSS 0.00488f
C5537 VDD.n3380 VSS 0.00798f
C5538 VDD.n3381 VSS 0.00374f
C5539 VDD.n3382 VSS 0.0225f
C5540 VDD.n3383 VSS 0.0809f
C5541 VDD.n3384 VSS 0.00488f
C5542 VDD.n3385 VSS 3.26e-19
C5543 VDD.n3386 VSS 0.00348f
C5544 VDD.n3387 VSS 0.00332f
C5545 VDD.n3388 VSS 0.00269f
C5546 VDD.n3389 VSS 0.00916f
C5547 VDD.n3390 VSS 0.00269f
C5548 VDD.n3391 VSS 0.00269f
C5549 VDD.n3392 VSS 0.00277f
C5550 VDD.n3393 VSS 0.0527f
C5551 VDD.n3394 VSS 0.00277f
C5552 VDD.n3395 VSS 0.00979f
C5553 VDD.n3396 VSS 0.245f
C5554 VDD.n3397 VSS 0.0129f
C5555 VDD.n3398 VSS 0.00979f
C5556 VDD.n3399 VSS 0.00269f
C5557 VDD.n3400 VSS 0.0294f
C5558 VDD.n3401 VSS 0.00332f
C5559 VDD.n3402 VSS 0.0286f
C5560 VDD.n3403 VSS 0.0294f
C5561 VDD.n3404 VSS 0.00332f
C5562 VDD.n3405 VSS 0.0261f
C5563 VDD.n3406 VSS 0.0261f
C5564 VDD.n3407 VSS 0.0286f
C5565 VDD.n3408 VSS 0.00348f
C5566 VDD.n3409 VSS 0.00269f
C5567 VDD.n3410 VSS 0.00269f
C5568 VDD.n3411 VSS 3.16e-19
C5569 VDD.n3412 VSS 0.0236f
C5570 VDD.n3413 VSS 0.124f
C5571 VDD.t69 VSS 0.47f
C5572 VDD.n3414 VSS 0.207f
C5573 VDD.t70 VSS 0.253f
C5574 VDD.n3415 VSS 0.198f
C5575 VDD.n3416 VSS 0.0104f
C5576 VDD.n3417 VSS 0.00269f
C5577 VDD.n3418 VSS 0.00663f
C5578 VDD.n3419 VSS 0.00348f
C5579 VDD.n3420 VSS 0.00806f
C5580 VDD.n3421 VSS 0.00472f
C5581 VDD.n3422 VSS 0.00411f
C5582 VDD.n3423 VSS 3.26e-19
C5583 VDD.n3424 VSS 0.00488f
C5584 VDD.n3425 VSS 0.023f
C5585 VDD.n3426 VSS 0.0138f
C5586 VDD.n3427 VSS 0.0142f
C5587 VDD.n3428 VSS -0.0753f
C5588 VDD.n3429 VSS 0.00411f
C5589 VDD.n3430 VSS 0.00585f
C5590 VDD.n3431 VSS -0.211f
C5591 VDD.n3432 VSS 0.00391f
C5592 VDD.n3433 VSS 0.00781f
C5593 VDD.n3434 VSS 0.0225f
C5594 VDD.n3435 VSS 0.0138f
C5595 VDD.n3436 VSS -0.182f
C5596 VDD.n3437 VSS 3.26e-19
C5597 VDD.n3438 VSS 0.00348f
C5598 VDD.n3439 VSS 0.00332f
C5599 VDD.n3440 VSS 0.00269f
C5600 VDD.n3441 VSS 0.00916f
C5601 VDD.n3442 VSS 0.00269f
C5602 VDD.n3443 VSS 0.00269f
C5603 VDD.n3444 VSS 0.0129f
C5604 VDD.n3445 VSS 0.00277f
C5605 VDD.n3446 VSS 3.16e-19
C5606 VDD.n3447 VSS 0.00916f
C5607 VDD.n3448 VSS 0.00585f
C5608 VDD.n3449 VSS 0.00806f
C5609 VDD.n3450 VSS 0.00663f
C5610 VDD.n3451 VSS 0.00332f
C5611 VDD.n3452 VSS 0.00979f
C5612 VDD.n3453 VSS 0.00979f
C5613 VDD.n3454 VSS 0.00269f
C5614 VDD.n3455 VSS 0.00277f
C5615 VDD.n3456 VSS 0.0527f
C5616 VDD.n3457 VSS 0.245f
C5617 VDD.n3458 VSS 0.198f
C5618 VDD.n3459 VSS 0.0104f
C5619 VDD.n3460 VSS 0.00269f
C5620 VDD.n3461 VSS 0.00663f
C5621 VDD.n3462 VSS 0.00348f
C5622 VDD.n3463 VSS 0.00806f
C5623 VDD.n3464 VSS 0.00472f
C5624 VDD.n3465 VSS 0.00411f
C5625 VDD.n3466 VSS 3.26e-19
C5626 VDD.n3467 VSS -0.211f
C5627 VDD.n3468 VSS 0.023f
C5628 VDD.n3469 VSS -0.078f
C5629 VDD.n3470 VSS 0.0142f
C5630 VDD.n3471 VSS 0.00439f
C5631 VDD.n3472 VSS 0.00411f
C5632 VDD.n3473 VSS 0.00585f
C5633 VDD.n3474 VSS 0.00488f
C5634 VDD.n3475 VSS 0.00391f
C5635 VDD.n3476 VSS 0.00781f
C5636 VDD.n3477 VSS 0.0225f
C5637 VDD.n3478 VSS 0.0138f
C5638 VDD.n3479 VSS 0.0225f
C5639 VDD.n3480 VSS 3.26e-19
C5640 VDD.n3481 VSS 0.00348f
C5641 VDD.n3482 VSS 0.00332f
C5642 VDD.n3483 VSS 0.00269f
C5643 VDD.n3484 VSS 0.00916f
C5644 VDD.n3485 VSS 0.00269f
C5645 VDD.n3486 VSS 0.00269f
C5646 VDD.n3487 VSS 0.0129f
C5647 VDD.n3488 VSS 0.00277f
C5648 VDD.n3489 VSS 3.16e-19
C5649 VDD.n3490 VSS 0.00916f
C5650 VDD.n3491 VSS 0.00585f
C5651 VDD.n3492 VSS 0.00806f
C5652 VDD.n3493 VSS 0.00663f
C5653 VDD.n3494 VSS 0.00332f
C5654 VDD.n3495 VSS 0.00979f
C5655 VDD.n3496 VSS 0.00979f
C5656 VDD.n3497 VSS 0.00269f
C5657 VDD.n3498 VSS 0.00277f
C5658 VDD.n3499 VSS 0.0527f
C5659 VDD.n3500 VSS 0.245f
C5660 VDD.n3501 VSS 0.198f
C5661 VDD.n3502 VSS 0.0104f
C5662 VDD.n3503 VSS 0.00269f
C5663 VDD.n3504 VSS 0.00663f
C5664 VDD.n3505 VSS 0.00348f
C5665 VDD.n3506 VSS 0.00806f
C5666 VDD.n3507 VSS 0.00332f
C5667 VDD.n3508 VSS 0.00781f
C5668 VDD.n3509 VSS 0.00439f
C5669 VDD.n3510 VSS 0.0138f
C5670 VDD.n3511 VSS 0.0142f
C5671 VDD.n3512 VSS 0.00439f
C5672 VDD.n3513 VSS 0.00411f
C5673 VDD.n3514 VSS 0.00585f
C5674 VDD.n3515 VSS 0.00488f
C5675 VDD.n3516 VSS 0.00391f
C5676 VDD.n3517 VSS 0.023f
C5677 VDD.n3518 VSS -0.182f
C5678 VDD.n3519 VSS 0.00488f
C5679 VDD.n3520 VSS 0.00472f
C5680 VDD.n3521 VSS -0.0844f
C5681 VDD.n3522 VSS 3.26e-19
C5682 VDD.n3523 VSS 0.00411f
C5683 VDD.n3524 VSS 0.00488f
C5684 VDD.n3525 VSS 0.00348f
C5685 VDD.n3526 VSS 0.0251f
C5686 VDD.n3527 VSS 0.0251f
C5687 VDD.n3528 VSS 0.00411f
C5688 VDD.n3529 VSS 0.0295f
C5689 VDD.n3530 VSS 0.0295f
C5690 VDD.n3531 VSS 0.00269f
C5691 VDD.n3532 VSS 0.00269f
C5692 VDD.n3533 VSS 0.00269f
C5693 VDD.n3534 VSS 0.00277f
C5694 VDD.n3535 VSS 0.0129f
C5695 VDD.n3536 VSS 3.16e-19
C5696 VDD.n3537 VSS 0.00269f
C5697 VDD.n3538 VSS 0.00277f
C5698 VDD.n3539 VSS 0.0527f
C5699 VDD.n3540 VSS 0.412f
C5700 VDD.n3541 VSS 0.0186f
C5701 VDD.n3542 VSS 0.03f
C5702 VDD.n3543 VSS 0.03f
C5703 VDD.n3544 VSS 0.0186f
C5704 VDD.n3545 VSS 0.226f
C5705 VDD.n3546 VSS 0.0527f
C5706 VDD.n3547 VSS 0.198f
C5707 VDD.n3548 VSS 0.0104f
C5708 VDD.n3549 VSS 0.00979f
C5709 VDD.n3550 VSS 0.00269f
C5710 VDD.n3551 VSS 0.00916f
C5711 VDD.n3552 VSS 4.74e-19
C5712 VDD.n3553 VSS 0.00332f
C5713 VDD.n3554 VSS 0.00585f
C5714 VDD.n3555 VSS 0.00348f
C5715 VDD.n3556 VSS 4.74e-19
C5716 VDD.n3557 VSS -0.211f
C5717 VDD.n3558 VSS 3.26e-19
C5718 VDD.n3559 VSS 0.023f
C5719 VDD.n3560 VSS 0.00439f
C5720 VDD.n3561 VSS -0.174f
C5721 VDD.n3562 VSS 0.00798f
C5722 VDD.n3563 VSS 0.00979f
C5723 VDD.n3564 VSS 0.00332f
C5724 VDD.n3565 VSS 0.00663f
C5725 VDD.n3566 VSS 0.00806f
C5726 VDD.n3567 VSS 0.00332f
C5727 VDD.n3568 VSS 0.00411f
C5728 VDD.n3569 VSS 0.00585f
C5729 VDD.n3570 VSS 0.00472f
C5730 VDD.n3571 VSS 0.00374f
C5731 VDD.n3572 VSS 0.0225f
C5732 VDD.n3573 VSS 0.0138f
C5733 VDD.n3574 VSS 0.0142f
C5734 VDD.n3575 VSS 3.26e-19
C5735 VDD.n3576 VSS 0.00488f
C5736 VDD.n3577 VSS 0.00798f
C5737 VDD.n3578 VSS 0.00374f
C5738 VDD.n3579 VSS 0.0225f
C5739 VDD.n3580 VSS 0.0225f
C5740 VDD.n3581 VSS 0.00488f
C5741 VDD.n3582 VSS 0.00439f
C5742 VDD.n3583 VSS 0.00806f
C5743 VDD.n3584 VSS 0.00332f
C5744 VDD.n3585 VSS 0.00663f
C5745 VDD.n3586 VSS 4.74e-19
C5746 VDD.n3587 VSS 0.00269f
C5747 VDD.n3588 VSS 0.00269f
C5748 VDD.n3589 VSS 0.00269f
C5749 VDD.n3590 VSS 0.00277f
C5750 VDD.n3591 VSS 0.0129f
C5751 VDD.n3592 VSS 0.198f
C5752 VDD.n3593 VSS 0.0104f
C5753 VDD.n3594 VSS 0.00979f
C5754 VDD.n3595 VSS 0.00979f
C5755 VDD.n3596 VSS 0.0129f
C5756 VDD.n3597 VSS 0.245f
C5757 VDD.n3598 VSS 0.0527f
C5758 VDD.n3599 VSS 0.00277f
C5759 VDD.n3600 VSS 0.00269f
C5760 VDD.n3601 VSS 3.16e-19
C5761 VDD.n3602 VSS 0.00269f
C5762 VDD.n3603 VSS 0.00348f
C5763 VDD.n3604 VSS 0.00269f
C5764 VDD.n3605 VSS 0.00332f
C5765 VDD.n3606 VSS 0.00979f
C5766 VDD.n3607 VSS 0.00979f
C5767 VDD.n3608 VSS 0.0129f
C5768 VDD.n3609 VSS 0.245f
C5769 VDD.n3610 VSS 0.0527f
C5770 VDD.n3611 VSS 0.198f
C5771 VDD.n3612 VSS 0.0104f
C5772 VDD.n3613 VSS 0.00979f
C5773 VDD.n3614 VSS 0.00269f
C5774 VDD.n3615 VSS 0.00916f
C5775 VDD.n3616 VSS 4.74e-19
C5776 VDD.n3617 VSS 0.00332f
C5777 VDD.n3618 VSS 0.00585f
C5778 VDD.n3619 VSS 0.00348f
C5779 VDD.n3620 VSS 4.74e-19
C5780 VDD.n3621 VSS -0.211f
C5781 VDD.n3622 VSS 3.26e-19
C5782 VDD.n3623 VSS 0.023f
C5783 VDD.n3624 VSS 0.00439f
C5784 VDD.n3625 VSS -0.174f
C5785 VDD.n3626 VSS 0.0138f
C5786 VDD.n3627 VSS -0.0844f
C5787 VDD.n3628 VSS 3.26e-19
C5788 VDD.n3629 VSS 0.00488f
C5789 VDD.n3630 VSS 0.00798f
C5790 VDD.n3631 VSS 0.00348f
C5791 VDD.n3632 VSS 0.00979f
C5792 VDD.n3633 VSS 0.00332f
C5793 VDD.n3634 VSS 0.00663f
C5794 VDD.n3635 VSS 0.00806f
C5795 VDD.n3636 VSS 0.00332f
C5796 VDD.n3637 VSS 0.00411f
C5797 VDD.n3638 VSS 0.00585f
C5798 VDD.n3639 VSS 0.00472f
C5799 VDD.n3640 VSS 0.00374f
C5800 VDD.n3641 VSS 0.0225f
C5801 VDD.n3642 VSS 0.0138f
C5802 VDD.n3643 VSS 0.0142f
C5803 VDD.n3644 VSS 3.26e-19
C5804 VDD.n3645 VSS 0.00488f
C5805 VDD.n3646 VSS 0.00798f
C5806 VDD.n3647 VSS 0.00374f
C5807 VDD.n3648 VSS 0.0225f
C5808 VDD.n3649 VSS 0.0809f
C5809 VDD.n3650 VSS 0.00488f
C5810 VDD.n3651 VSS 3.26e-19
C5811 VDD.n3652 VSS 0.00348f
C5812 VDD.n3653 VSS 0.00332f
C5813 VDD.n3654 VSS 0.00269f
C5814 VDD.n3655 VSS 0.00916f
C5815 VDD.n3656 VSS 0.00269f
C5816 VDD.n3657 VSS 0.00269f
C5817 VDD.n3658 VSS 0.00277f
C5818 VDD.n3659 VSS 0.0527f
C5819 VDD.n3660 VSS 0.00277f
C5820 VDD.n3661 VSS 0.00979f
C5821 VDD.n3662 VSS 0.245f
C5822 VDD.n3663 VSS 0.0129f
C5823 VDD.n3664 VSS 0.00979f
C5824 VDD.n3665 VSS 0.00269f
C5825 VDD.n3666 VSS 0.0294f
C5826 VDD.n3667 VSS 0.00332f
C5827 VDD.n3668 VSS 0.0286f
C5828 VDD.n3669 VSS 0.0294f
C5829 VDD.n3670 VSS 0.00332f
C5830 VDD.n3671 VSS 0.0261f
C5831 VDD.n3672 VSS 0.0261f
C5832 VDD.n3673 VSS 0.0286f
C5833 VDD.n3674 VSS 0.00348f
C5834 VDD.n3675 VSS 0.00269f
C5835 VDD.n3676 VSS 0.00269f
C5836 VDD.n3677 VSS 3.16e-19
C5837 VDD.n3678 VSS 0.0236f
C5838 VDD.n3679 VSS 0.124f
C5839 VDD.t73 VSS 0.47f
C5840 VDD.n3680 VSS 0.207f
C5841 VDD.t2 VSS 0.253f
C5842 VDD.n3681 VSS 0.198f
C5843 VDD.n3682 VSS 0.0104f
C5844 VDD.n3683 VSS 0.00269f
C5845 VDD.n3684 VSS 0.00663f
C5846 VDD.n3685 VSS 0.00348f
C5847 VDD.n3686 VSS 0.00806f
C5848 VDD.n3687 VSS 0.00472f
C5849 VDD.n3688 VSS 0.00411f
C5850 VDD.n3689 VSS 3.26e-19
C5851 VDD.n3690 VSS 0.00488f
C5852 VDD.n3691 VSS 0.023f
C5853 VDD.n3692 VSS 0.0138f
C5854 VDD.n3693 VSS 0.0142f
C5855 VDD.n3694 VSS -0.0753f
C5856 VDD.n3695 VSS 0.00411f
C5857 VDD.n3696 VSS 0.00585f
C5858 VDD.n3697 VSS -0.211f
C5859 VDD.n3698 VSS 0.00391f
C5860 VDD.n3699 VSS 0.00781f
C5861 VDD.n3700 VSS 0.0225f
C5862 VDD.n3701 VSS 0.0138f
C5863 VDD.n3702 VSS -0.182f
C5864 VDD.n3703 VSS 3.26e-19
C5865 VDD.n3704 VSS 0.00348f
C5866 VDD.n3705 VSS 0.00332f
C5867 VDD.n3706 VSS 0.00269f
C5868 VDD.n3707 VSS 0.00916f
C5869 VDD.n3708 VSS 0.00269f
C5870 VDD.n3709 VSS 0.00269f
C5871 VDD.n3710 VSS 0.0129f
C5872 VDD.n3711 VSS 0.00277f
C5873 VDD.n3712 VSS 3.16e-19
C5874 VDD.n3713 VSS 0.00916f
C5875 VDD.n3714 VSS 0.00585f
C5876 VDD.n3715 VSS 0.00806f
C5877 VDD.n3716 VSS 0.00663f
C5878 VDD.n3717 VSS 0.00332f
C5879 VDD.n3718 VSS 0.00979f
C5880 VDD.n3719 VSS 0.00979f
C5881 VDD.n3720 VSS 0.00269f
C5882 VDD.n3721 VSS 0.00277f
C5883 VDD.n3722 VSS 0.0527f
C5884 VDD.n3723 VSS 0.245f
C5885 VDD.n3724 VSS 0.198f
C5886 VDD.n3725 VSS 0.0104f
C5887 VDD.n3726 VSS 0.00269f
C5888 VDD.n3727 VSS 0.00663f
C5889 VDD.n3728 VSS 0.00348f
C5890 VDD.n3729 VSS 0.00806f
C5891 VDD.n3730 VSS 0.00472f
C5892 VDD.n3731 VSS 0.00411f
C5893 VDD.n3732 VSS 3.26e-19
C5894 VDD.n3733 VSS -0.211f
C5895 VDD.n3734 VSS 0.023f
C5896 VDD.n3735 VSS -0.078f
C5897 VDD.n3736 VSS 0.0142f
C5898 VDD.n3737 VSS 0.00439f
C5899 VDD.n3738 VSS 0.00411f
C5900 VDD.n3739 VSS 0.00585f
C5901 VDD.n3740 VSS 0.00488f
C5902 VDD.n3741 VSS 0.00391f
C5903 VDD.n3742 VSS 0.00781f
C5904 VDD.n3743 VSS 0.0225f
C5905 VDD.n3744 VSS 0.0138f
C5906 VDD.n3745 VSS 0.0225f
C5907 VDD.n3746 VSS 3.26e-19
C5908 VDD.n3747 VSS 0.00348f
C5909 VDD.n3748 VSS 0.00332f
C5910 VDD.n3749 VSS 0.00269f
C5911 VDD.n3750 VSS 0.00916f
C5912 VDD.n3751 VSS 0.00269f
C5913 VDD.n3752 VSS 0.00269f
C5914 VDD.n3753 VSS 0.0129f
C5915 VDD.n3754 VSS 0.00277f
C5916 VDD.n3755 VSS 3.16e-19
C5917 VDD.n3756 VSS 0.00916f
C5918 VDD.n3757 VSS 0.00585f
C5919 VDD.n3758 VSS 0.00806f
C5920 VDD.n3759 VSS 0.00663f
C5921 VDD.n3760 VSS 0.00332f
C5922 VDD.n3761 VSS 0.00979f
C5923 VDD.n3762 VSS 0.00979f
C5924 VDD.n3763 VSS 0.00269f
C5925 VDD.n3764 VSS 0.00277f
C5926 VDD.n3765 VSS 0.0527f
C5927 VDD.n3766 VSS 0.245f
C5928 VDD.n3767 VSS 0.198f
C5929 VDD.n3768 VSS 0.0104f
C5930 VDD.n3769 VSS 0.00269f
C5931 VDD.n3770 VSS 0.00663f
C5932 VDD.n3771 VSS 0.0422f
C5933 VDD.n3772 VSS 0.00806f
C5934 VDD.n3773 VSS 0.00332f
C5935 VDD.n3774 VSS 0.00781f
C5936 VDD.n3775 VSS 0.00439f
C5937 VDD.n3776 VSS 0.0138f
C5938 VDD.n3777 VSS 0.0142f
C5939 VDD.n3778 VSS 0.00439f
C5940 VDD.n3779 VSS 0.00411f
C5941 VDD.n3780 VSS 0.00585f
C5942 VDD.n3781 VSS 0.00488f
C5943 VDD.n3782 VSS 0.00391f
C5944 VDD.n3783 VSS 0.023f
C5945 VDD.n3784 VSS -0.182f
C5946 VDD.n3785 VSS 0.0457f
C5947 VDD.n3786 VSS 0.0199f
C5948 VDD.n3787 VSS 0.00634f
C5949 VDD.n3788 VSS 0.02f
C5950 VDD.n3789 VSS 0.0457f
C5951 VDD.n3790 VSS 0.0199f
C5952 VDD.n3791 VSS 0.00634f
C5953 VDD.n3792 VSS 0.02f
C5954 VDD.n3793 VSS 0.0457f
C5955 VDD.n3794 VSS 0.0199f
C5956 VDD.n3795 VSS 0.00634f
C5957 VDD.n3796 VSS 0.02f
C5958 VDD.n3797 VSS 0.0457f
C5959 VDD.n3798 VSS 0.0199f
C5960 VDD.n3799 VSS 0.00634f
C5961 VDD.n3800 VSS 0.02f
C5962 VDD.n3801 VSS 0.0457f
C5963 VDD.n3802 VSS 0.0199f
C5964 VDD.n3803 VSS 0.00634f
C5965 VDD.n3804 VSS 0.00839f
C5966 VDD.n3805 VSS 0.00839f
C5967 VDD.n3806 VSS 0.0081f
C5968 VDD.n3807 VSS 0.0813f
C5969 VDD.n3808 VSS 0.149f
C5970 VDD.n3809 VSS 0.00839f
C5971 VDD.n3810 VSS 0.0081f
C5972 VDD.n3811 VSS 0.0813f
C5973 VDD.n3812 VSS 0.00839f
C5974 VDD.n3813 VSS 0.0081f
C5975 VDD.n3814 VSS 0.0813f
C5976 VDD.n3815 VSS 0.00839f
C5977 VDD.n3816 VSS 0.0081f
C5978 VDD.n3817 VSS 0.0813f
C5979 VDD.n3818 VSS 0.0527f
C5980 VDD.n3819 VSS 0.00277f
C5981 VDD.n3820 VSS 0.0418f
C5982 VDD.n3821 VSS 0.018f
C5983 VDD.n3822 VSS 0.413f
C5984 VDD.t5 VSS 0.555f
C5985 VDD.t3 VSS 0.308f
C5986 VDD.n3823 VSS 0.132f
C5987 VDD.t4 VSS 0.944f
C5988 VDD.n3824 VSS 0.212f
C5989 VDD.n3825 VSS 0.0695f
C5990 VDD.n3826 VSS 0.0813f
C5991 VDD.n3827 VSS 0.0081f
C5992 VDD.n3828 VSS 0.02f
C5993 VDD.n3829 VSS 0.0458f
C5994 VDD.n3830 VSS 0.0199f
C5995 VDD.t6 VSS 0.00943f
C5996 VDD.n3831 VSS 0.136f
C5997 VDD.n3832 VSS 0.02f
C5998 VDD.n3833 VSS 0.0193f
C5999 VDD.n3834 VSS 0.0168f
C6000 VDD.n3835 VSS 0.00786f
C6001 VDD.n3836 VSS 0.0172f
C6002 VDD.n3837 VSS 0.00659f
C6003 VDD.t52 VSS 0.00663f
C6004 VDD.t39 VSS 0.00663f
C6005 VDD.n3838 VSS 0.0163f
C6006 VDD.n3839 VSS 0.0482f
C6007 VDD.n3840 VSS 0.00805f
C6008 VDD.n3841 VSS 0.0164f
C6009 VDD.n3842 VSS 0.097f
C6010 VDD.n3843 VSS 0.116f
C6011 VDD.n3844 VSS 0.0109f
C6012 VDD.n3845 VSS 0.161f
C6013 VDD.n3846 VSS 0.161f
C6014 VDD.n3847 VSS 0.0109f
C6015 VDD.n3848 VSS 0.0967f
C6016 VDD.n3849 VSS 0.0967f
C6017 VDD.n3850 VSS 0.0109f
C6018 VDD.n3851 VSS 0.107f
C6019 VDD.n3852 VSS 0.107f
C6020 VDD.n3853 VSS 0.0109f
C6021 VDD.n3854 VSS 0.0929f
C6022 VDD.n3855 VSS 0.0929f
C6023 VDD.n3856 VSS 0.0109f
C6024 VDD.n3857 VSS 0.0868f
C6025 VDD.n3858 VSS 0.0868f
C6026 VDD.n3859 VSS 0.0109f
C6027 VDD.n3860 VSS 0.22f
C6028 VDD.n3861 VSS 0.0389f
C6029 VDD.n3862 VSS 0.0398f
C6030 VDD.n3863 VSS 0.0607f
C6031 VDD.n3864 VSS 0.0142f
C6032 VDD.n3865 VSS -0.078f
C6033 VDD.n3866 VSS 3.26e-19
C6034 VDD.n3867 VSS 0.00472f
C6035 VDD.n3868 VSS 4.74e-19
C6036 VDD.n3869 VSS 0.00348f
C6037 VDD.n3870 VSS 0.00269f
C6038 VDD.n3871 VSS 0.00332f
C6039 VDD.n3872 VSS 0.00979f
C6040 VDD.n3873 VSS 0.00979f
C6041 VDD.n3874 VSS 0.0129f
C6042 VDD.n3875 VSS 0.245f
C6043 VDD.n3876 VSS 0.0527f
C6044 VDD.n3877 VSS 0.198f
C6045 VDD.n3878 VSS 0.0104f
C6046 VDD.n3879 VSS 3.16e-19
C6047 VDD.n3880 VSS 0.00348f
C6048 VDD.n3881 VSS 4.74e-19
C6049 VDD.n3882 VSS 0.00472f
C6050 VDD.n3883 VSS 0.00781f
C6051 VDD.n3884 VSS 0.00391f
C6052 VDD.n3885 VSS 0.023f
C6053 VDD.n3886 VSS 0.0142f
C6054 VDD.n3887 VSS -0.0753f
C6055 VDD.n3888 VSS 0.00332f
C6056 VDD.n3889 VSS 4.74e-19
C6057 VDD.n3890 VSS 0.00348f
C6058 VDD.n3891 VSS 0.00269f
C6059 VDD.n3892 VSS 0.00332f
C6060 VDD.n3893 VSS 0.00979f
C6061 VDD.n3894 VSS 0.00979f
C6062 VDD.n3895 VSS 0.0129f
C6063 VDD.n3896 VSS 0.245f
C6064 VDD.n3897 VSS 0.0527f
C6065 VDD.n3898 VSS 0.198f
C6066 VDD.n3899 VSS 0.0104f
C6067 VDD.n3900 VSS 3.16e-19
C6068 VDD.n3901 VSS 0.00348f
C6069 VDD.n3902 VSS 4.74e-19
C6070 VDD.n3903 VSS 0.00472f
C6071 VDD.n3904 VSS 0.00781f
C6072 VDD.n3905 VSS 0.00391f
C6073 VDD.n3906 VSS 0.023f
C6074 VDD.n3907 VSS 0.0142f
C6075 VDD.n3908 VSS 0.00439f
C6076 VDD.n3909 VSS 0.00332f
C6077 VDD.n3910 VSS 4.74e-19
C6078 VDD.n3911 VSS 0.00348f
C6079 VDD.n3912 VSS 0.00269f
C6080 VDD.n3913 VSS 0.00332f
C6081 VDD.n3914 VSS 0.00979f
C6082 VDD.n3915 VSS 0.00979f
C6083 VDD.n3916 VSS 0.0129f
C6084 VDD.n3917 VSS 0.245f
C6085 VDD.n3918 VSS 0.0527f
C6086 VDD.n3919 VSS 0.124f
C6087 VDD.n3920 VSS 0.0236f
C6088 VDD.n3921 VSS 3.16e-19
C6089 VDD.n3922 VSS 0.00348f
C6090 VDD.n3923 VSS 4.74e-19
C6091 VDD.n3924 VSS 0.00472f
C6092 VDD.n3925 VSS 0.0285f
C6093 VDD.n3926 VSS 0.0286f
C6094 VDD.n3927 VSS 0.0813f
C6095 VDD.n3928 VSS 0.0142f
C6096 VDD.n3929 VSS 0.0138f
C6097 VDD.n3930 VSS -0.0753f
C6098 VDD.n3931 VSS 0.00332f
C6099 VDD.n3932 VSS 0.00411f
C6100 VDD.n3933 VSS 0.00916f
C6101 VDD.n3934 VSS 0.00663f
C6102 VDD.n3935 VSS 0.00806f
C6103 VDD.n3936 VSS 0.00348f
C6104 VDD.n3937 VSS 0.00269f
C6105 VDD.n3938 VSS 0.00348f
C6106 VDD.n3939 VSS 3.16e-19
C6107 VDD.n3940 VSS 0.00269f
C6108 VDD.n3941 VSS 0.00277f
C6109 VDD.n3942 VSS 0.0527f
C6110 VDD.n3943 VSS 0.245f
C6111 VDD.n3944 VSS 0.198f
C6112 VDD.n3945 VSS 0.0104f
C6113 VDD.n3946 VSS 3.16e-19
C6114 VDD.n3947 VSS 0.00348f
C6115 VDD.n3948 VSS 0.00916f
C6116 VDD.n3949 VSS 0.00411f
C6117 VDD.n3950 VSS 0.00585f
C6118 VDD.n3951 VSS 0.00472f
C6119 VDD.n3952 VSS 0.00374f
C6120 VDD.n3953 VSS 0.00798f
C6121 VDD.n3954 VSS 0.023f
C6122 VDD.n3955 VSS 0.0142f
C6123 VDD.n3956 VSS 0.0138f
C6124 VDD.n3957 VSS -0.0753f
C6125 VDD.n3958 VSS 0.00332f
C6126 VDD.n3959 VSS 0.00411f
C6127 VDD.n3960 VSS 0.00916f
C6128 VDD.n3961 VSS 0.00663f
C6129 VDD.n3962 VSS 0.00806f
C6130 VDD.n3963 VSS 0.00348f
C6131 VDD.n3964 VSS 0.00269f
C6132 VDD.n3965 VSS 0.00348f
C6133 VDD.n3966 VSS 3.16e-19
C6134 VDD.n3967 VSS 0.00269f
C6135 VDD.n3968 VSS 0.00277f
C6136 VDD.n3969 VSS 0.0527f
C6137 VDD.n3970 VSS 0.245f
C6138 VDD.n3971 VSS 0.198f
C6139 VDD.n3972 VSS 0.0104f
C6140 VDD.n3973 VSS 3.16e-19
C6141 VDD.n3974 VSS 0.00348f
C6142 VDD.n3975 VSS 4.74e-19
C6143 VDD.n3976 VSS 0.00332f
C6144 VDD.n3977 VSS 0.00439f
C6145 VDD.n3978 VSS 0.0138f
C6146 VDD.n3979 VSS 0.0142f
C6147 VDD.n3980 VSS 0.0241f
C6148 VDD.n3981 VSS 0.0243f
C6149 VDD.n3982 VSS 0.0607f
C6150 VDD.n3983 VSS 0.0142f
C6151 VDD.n3984 VSS -0.078f
C6152 VDD.n3985 VSS 3.26e-19
C6153 VDD.n3986 VSS 0.00472f
C6154 VDD.n3987 VSS 4.74e-19
C6155 VDD.n3988 VSS 0.00348f
C6156 VDD.n3989 VSS 0.00269f
C6157 VDD.n3990 VSS 0.00332f
C6158 VDD.n3991 VSS 0.00979f
C6159 VDD.n3992 VSS 0.00979f
C6160 VDD.n3993 VSS 0.0129f
C6161 VDD.n3994 VSS 0.245f
C6162 VDD.n3995 VSS 0.0527f
C6163 VDD.n3996 VSS 0.198f
C6164 VDD.n3997 VSS 0.0104f
C6165 VDD.n3998 VSS 3.16e-19
C6166 VDD.n3999 VSS 0.00348f
C6167 VDD.n4000 VSS 4.74e-19
C6168 VDD.n4001 VSS 0.00472f
C6169 VDD.n4002 VSS 0.00781f
C6170 VDD.n4003 VSS 0.00391f
C6171 VDD.n4004 VSS 0.023f
C6172 VDD.n4005 VSS 0.0142f
C6173 VDD.n4006 VSS -0.0753f
C6174 VDD.n4007 VSS 0.00332f
C6175 VDD.n4008 VSS 4.74e-19
C6176 VDD.n4009 VSS 0.00348f
C6177 VDD.n4010 VSS 0.00269f
C6178 VDD.n4011 VSS 0.00332f
C6179 VDD.n4012 VSS 0.00979f
C6180 VDD.n4013 VSS 0.00979f
C6181 VDD.n4014 VSS 0.0129f
C6182 VDD.n4015 VSS 0.245f
C6183 VDD.n4016 VSS 0.0527f
C6184 VDD.n4017 VSS 0.198f
C6185 VDD.n4018 VSS 0.0104f
C6186 VDD.n4019 VSS 3.16e-19
C6187 VDD.n4020 VSS 0.00348f
C6188 VDD.n4021 VSS 4.74e-19
C6189 VDD.n4022 VSS 0.00472f
C6190 VDD.n4023 VSS 0.00781f
C6191 VDD.n4024 VSS 0.00391f
C6192 VDD.n4025 VSS 0.023f
C6193 VDD.n4026 VSS 0.0142f
C6194 VDD.n4027 VSS 0.00439f
C6195 VDD.n4028 VSS 0.00332f
C6196 VDD.n4029 VSS 4.74e-19
C6197 VDD.n4030 VSS 0.00348f
C6198 VDD.n4031 VSS 0.00269f
C6199 VDD.n4032 VSS 0.00332f
C6200 VDD.n4033 VSS 0.00979f
C6201 VDD.n4034 VSS 0.00979f
C6202 VDD.n4035 VSS 0.0129f
C6203 VDD.n4036 VSS 0.245f
C6204 VDD.n4037 VSS 0.0527f
C6205 VDD.n4038 VSS 0.124f
C6206 VDD.n4039 VSS 0.0236f
C6207 VDD.n4040 VSS 3.16e-19
C6208 VDD.n4041 VSS 0.00348f
C6209 VDD.n4042 VSS 4.74e-19
C6210 VDD.n4043 VSS 0.00472f
C6211 VDD.n4044 VSS 0.0285f
C6212 VDD.n4045 VSS 0.0286f
C6213 VDD.n4046 VSS 0.0813f
C6214 VDD.n4047 VSS 0.0142f
C6215 VDD.n4048 VSS 0.0138f
C6216 VDD.n4049 VSS -0.0753f
C6217 VDD.n4050 VSS 0.00332f
C6218 VDD.n4051 VSS 0.00411f
C6219 VDD.n4052 VSS 0.00916f
C6220 VDD.n4053 VSS 0.00663f
C6221 VDD.n4054 VSS 0.00806f
C6222 VDD.n4055 VSS 0.00348f
C6223 VDD.n4056 VSS 0.00269f
C6224 VDD.n4057 VSS 0.00348f
C6225 VDD.n4058 VSS 3.16e-19
C6226 VDD.n4059 VSS 0.00269f
C6227 VDD.n4060 VSS 0.00277f
C6228 VDD.n4061 VSS 0.0527f
C6229 VDD.n4062 VSS 0.245f
C6230 VDD.n4063 VSS 0.198f
C6231 VDD.n4064 VSS 0.0104f
C6232 VDD.n4065 VSS 3.16e-19
C6233 VDD.n4066 VSS 0.00348f
C6234 VDD.n4067 VSS 0.00916f
C6235 VDD.n4068 VSS 0.00411f
C6236 VDD.n4069 VSS 0.00585f
C6237 VDD.n4070 VSS 0.00472f
C6238 VDD.n4071 VSS 0.00374f
C6239 VDD.n4072 VSS 0.00798f
C6240 VDD.n4073 VSS 0.023f
C6241 VDD.n4074 VSS 0.0142f
C6242 VDD.n4075 VSS 0.0138f
C6243 VDD.n4076 VSS -0.0753f
C6244 VDD.n4077 VSS 0.00332f
C6245 VDD.n4078 VSS 0.00411f
C6246 VDD.n4079 VSS 0.00916f
C6247 VDD.n4080 VSS 0.00663f
C6248 VDD.n4081 VSS 0.00806f
C6249 VDD.n4082 VSS 0.00348f
C6250 VDD.n4083 VSS 0.00269f
C6251 VDD.n4084 VSS 0.00348f
C6252 VDD.n4085 VSS 3.16e-19
C6253 VDD.n4086 VSS 0.00269f
C6254 VDD.n4087 VSS 0.00277f
C6255 VDD.n4088 VSS 0.0527f
C6256 VDD.n4089 VSS 0.245f
C6257 VDD.n4090 VSS 0.198f
C6258 VDD.n4091 VSS 0.0104f
C6259 VDD.n4092 VSS 3.16e-19
C6260 VDD.n4093 VSS 0.00348f
C6261 VDD.n4094 VSS 4.74e-19
C6262 VDD.n4095 VSS 0.00332f
C6263 VDD.n4096 VSS 0.00439f
C6264 VDD.n4097 VSS 0.0138f
C6265 VDD.n4098 VSS 0.0142f
C6266 VDD.n4099 VSS 0.0241f
C6267 VDD.n4100 VSS 0.0243f
C6268 VDD.n4101 VSS 0.0607f
C6269 VDD.n4102 VSS 0.0142f
C6270 VDD.n4103 VSS -0.078f
C6271 VDD.n4104 VSS 3.26e-19
C6272 VDD.n4105 VSS 0.00472f
C6273 VDD.n4106 VSS 4.74e-19
C6274 VDD.n4107 VSS 0.00348f
C6275 VDD.n4108 VSS 0.00269f
C6276 VDD.n4109 VSS 0.00332f
C6277 VDD.n4110 VSS 0.00979f
C6278 VDD.n4111 VSS 0.00979f
C6279 VDD.n4112 VSS 0.0129f
C6280 VDD.n4113 VSS 0.245f
C6281 VDD.n4114 VSS 0.0527f
C6282 VDD.n4115 VSS 0.198f
C6283 VDD.n4116 VSS 0.0104f
C6284 VDD.n4117 VSS 3.16e-19
C6285 VDD.n4118 VSS 0.00348f
C6286 VDD.n4119 VSS 4.74e-19
C6287 VDD.n4120 VSS 0.00472f
C6288 VDD.n4121 VSS 0.00781f
C6289 VDD.n4122 VSS 0.00391f
C6290 VDD.n4123 VSS 0.023f
C6291 VDD.n4124 VSS 0.0142f
C6292 VDD.n4125 VSS -0.0753f
C6293 VDD.n4126 VSS 0.00332f
C6294 VDD.n4127 VSS 4.74e-19
C6295 VDD.n4128 VSS 0.00348f
C6296 VDD.n4129 VSS 0.00269f
C6297 VDD.n4130 VSS 0.00332f
C6298 VDD.n4131 VSS 0.00979f
C6299 VDD.n4132 VSS 0.00979f
C6300 VDD.n4133 VSS 0.0129f
C6301 VDD.n4134 VSS 0.245f
C6302 VDD.n4135 VSS 0.0527f
C6303 VDD.n4136 VSS 0.198f
C6304 VDD.n4137 VSS 0.0104f
C6305 VDD.n4138 VSS 3.16e-19
C6306 VDD.n4139 VSS 0.00348f
C6307 VDD.n4140 VSS 4.74e-19
C6308 VDD.n4141 VSS 0.00472f
C6309 VDD.n4142 VSS 0.00781f
C6310 VDD.n4143 VSS 0.00391f
C6311 VDD.n4144 VSS 0.023f
C6312 VDD.n4145 VSS 0.0142f
C6313 VDD.n4146 VSS 0.00439f
C6314 VDD.n4147 VSS 0.00332f
C6315 VDD.n4148 VSS 4.74e-19
C6316 VDD.n4149 VSS 0.00348f
C6317 VDD.n4150 VSS 0.00269f
C6318 VDD.n4151 VSS 0.00332f
C6319 VDD.n4152 VSS 0.00979f
C6320 VDD.n4153 VSS 0.00979f
C6321 VDD.n4154 VSS 0.0129f
C6322 VDD.n4155 VSS 0.245f
C6323 VDD.n4156 VSS 0.0527f
C6324 VDD.n4157 VSS 0.124f
C6325 VDD.n4158 VSS 0.0236f
C6326 VDD.n4159 VSS 3.16e-19
C6327 VDD.n4160 VSS 0.00348f
C6328 VDD.n4161 VSS 4.74e-19
C6329 VDD.n4162 VSS 0.00472f
C6330 VDD.n4163 VSS 0.0285f
C6331 VDD.n4164 VSS 0.0286f
C6332 VDD.n4165 VSS 0.0813f
C6333 VDD.n4166 VSS 0.0142f
C6334 VDD.n4167 VSS 0.0138f
C6335 VDD.n4168 VSS -0.0753f
C6336 VDD.n4169 VSS 0.00332f
C6337 VDD.n4170 VSS 0.00411f
C6338 VDD.n4171 VSS 0.00916f
C6339 VDD.n4172 VSS 0.00663f
C6340 VDD.n4173 VSS 0.00806f
C6341 VDD.n4174 VSS 0.00348f
C6342 VDD.n4175 VSS 0.00269f
C6343 VDD.n4176 VSS 0.00348f
C6344 VDD.n4177 VSS 3.16e-19
C6345 VDD.n4178 VSS 0.00269f
C6346 VDD.n4179 VSS 0.00277f
C6347 VDD.n4180 VSS 0.0527f
C6348 VDD.n4181 VSS 0.245f
C6349 VDD.n4182 VSS 0.198f
C6350 VDD.n4183 VSS 0.0104f
C6351 VDD.n4184 VSS 3.16e-19
C6352 VDD.n4185 VSS 0.00348f
C6353 VDD.n4186 VSS 0.00916f
C6354 VDD.n4187 VSS 0.00411f
C6355 VDD.n4188 VSS 0.00585f
C6356 VDD.n4189 VSS 0.00472f
C6357 VDD.n4190 VSS 0.00374f
C6358 VDD.n4191 VSS 0.00798f
C6359 VDD.n4192 VSS 0.023f
C6360 VDD.n4193 VSS 0.0142f
C6361 VDD.n4194 VSS 0.0138f
C6362 VDD.n4195 VSS -0.0753f
C6363 VDD.n4196 VSS 0.00332f
C6364 VDD.n4197 VSS 0.00411f
C6365 VDD.n4198 VSS 0.00916f
C6366 VDD.n4199 VSS 0.00663f
C6367 VDD.n4200 VSS 0.00806f
C6368 VDD.n4201 VSS 0.00348f
C6369 VDD.n4202 VSS 0.00269f
C6370 VDD.n4203 VSS 0.00348f
C6371 VDD.n4204 VSS 3.16e-19
C6372 VDD.n4205 VSS 0.00269f
C6373 VDD.n4206 VSS 0.00277f
C6374 VDD.n4207 VSS 0.0527f
C6375 VDD.n4208 VSS 0.245f
C6376 VDD.n4209 VSS 0.198f
C6377 VDD.n4210 VSS 0.0104f
C6378 VDD.n4211 VSS 3.16e-19
C6379 VDD.n4212 VSS 0.00348f
C6380 VDD.n4213 VSS 4.74e-19
C6381 VDD.n4214 VSS 0.00332f
C6382 VDD.n4215 VSS 0.00439f
C6383 VDD.n4216 VSS 0.0138f
C6384 VDD.n4217 VSS 0.0142f
C6385 VDD.n4218 VSS 0.0241f
C6386 VDD.n4219 VSS 0.0243f
C6387 VDD.n4220 VSS 0.0607f
C6388 VDD.n4221 VSS 0.0142f
C6389 VDD.n4222 VSS -0.078f
C6390 VDD.n4223 VSS 3.26e-19
C6391 VDD.n4224 VSS 0.00472f
C6392 VDD.n4225 VSS 4.74e-19
C6393 VDD.n4226 VSS 0.00348f
C6394 VDD.n4227 VSS 0.00269f
C6395 VDD.n4228 VSS 0.00332f
C6396 VDD.n4229 VSS 0.00979f
C6397 VDD.n4230 VSS 0.00979f
C6398 VDD.n4231 VSS 0.0129f
C6399 VDD.n4232 VSS 0.245f
C6400 VDD.n4233 VSS 0.0527f
C6401 VDD.n4234 VSS 0.198f
C6402 VDD.n4235 VSS 0.0104f
C6403 VDD.n4236 VSS 3.16e-19
C6404 VDD.n4237 VSS 0.00348f
C6405 VDD.n4238 VSS 4.74e-19
C6406 VDD.n4239 VSS 0.00472f
C6407 VDD.n4240 VSS 0.00781f
C6408 VDD.n4241 VSS 0.00391f
C6409 VDD.n4242 VSS 0.023f
C6410 VDD.n4243 VSS 0.0142f
C6411 VDD.n4244 VSS -0.0753f
C6412 VDD.n4245 VSS 0.00332f
C6413 VDD.n4246 VSS 4.74e-19
C6414 VDD.n4247 VSS 0.00348f
C6415 VDD.n4248 VSS 0.00269f
C6416 VDD.n4249 VSS 0.00332f
C6417 VDD.n4250 VSS 0.00979f
C6418 VDD.n4251 VSS 0.00979f
C6419 VDD.n4252 VSS 0.0129f
C6420 VDD.n4253 VSS 0.245f
C6421 VDD.n4254 VSS 0.0527f
C6422 VDD.n4255 VSS 0.198f
C6423 VDD.n4256 VSS 0.0104f
C6424 VDD.n4257 VSS 3.16e-19
C6425 VDD.n4258 VSS 0.00348f
C6426 VDD.n4259 VSS 4.74e-19
C6427 VDD.n4260 VSS 0.00472f
C6428 VDD.n4261 VSS 0.00781f
C6429 VDD.n4262 VSS 0.00391f
C6430 VDD.n4263 VSS 0.023f
C6431 VDD.n4264 VSS 0.0142f
C6432 VDD.n4265 VSS 0.00439f
C6433 VDD.n4266 VSS 0.00332f
C6434 VDD.n4267 VSS 4.74e-19
C6435 VDD.n4268 VSS 0.00348f
C6436 VDD.n4269 VSS 0.00269f
C6437 VDD.n4270 VSS 0.00332f
C6438 VDD.n4271 VSS 0.00979f
C6439 VDD.n4272 VSS 0.00979f
C6440 VDD.n4273 VSS 0.0129f
C6441 VDD.n4274 VSS 0.245f
C6442 VDD.n4275 VSS 0.0527f
C6443 VDD.n4276 VSS 0.124f
C6444 VDD.n4277 VSS 0.0236f
C6445 VDD.n4278 VSS 3.16e-19
C6446 VDD.n4279 VSS 0.00269f
C6447 VDD.n4280 VSS 0.0294f
C6448 VDD.n4281 VSS 0.00332f
C6449 VDD.n4282 VSS 0.0261f
C6450 VDD.n4283 VSS 0.0261f
C6451 VDD.n4284 VSS 0.0286f
C6452 VDD.n4285 VSS 0.00348f
C6453 VDD.n4286 VSS 0.00269f
C6454 VDD.n4287 VSS 0.00348f
C6455 VDD.n4288 VSS 3.16e-19
C6456 VDD.n4289 VSS 0.00269f
C6457 VDD.n4290 VSS 0.00277f
C6458 VDD.n4291 VSS 0.0527f
C6459 VDD.n4292 VSS 0.245f
C6460 VDD.n4293 VSS 0.198f
C6461 VDD.n4294 VSS 0.0104f
C6462 VDD.n4295 VSS 3.16e-19
C6463 VDD.n4296 VSS 0.00348f
C6464 VDD.n4297 VSS 0.00916f
C6465 VDD.n4298 VSS 0.00411f
C6466 VDD.n4299 VSS 0.00585f
C6467 VDD.n4300 VSS 0.00472f
C6468 VDD.n4301 VSS 0.00374f
C6469 VDD.n4302 VSS 0.00798f
C6470 VDD.n4303 VSS -0.174f
C6471 VDD.n4304 VSS -0.0844f
C6472 VDD.n4305 VSS 0.0138f
C6473 VDD.n4306 VSS 0.00439f
C6474 VDD.n4307 VSS 0.00332f
C6475 VDD.n4308 VSS 0.00411f
C6476 VDD.n4309 VSS 0.00916f
C6477 VDD.n4310 VSS 0.00663f
C6478 VDD.n4311 VSS 0.00806f
C6479 VDD.n4312 VSS 0.00348f
C6480 VDD.n4313 VSS 0.00269f
C6481 VDD.n4314 VSS 0.00348f
C6482 VDD.n4315 VSS 3.16e-19
C6483 VDD.n4316 VSS 0.00269f
C6484 VDD.n4317 VSS 0.00277f
C6485 VDD.n4318 VSS 0.0527f
C6486 VDD.n4319 VSS 0.245f
C6487 VDD.n4320 VSS 0.198f
C6488 VDD.n4321 VSS 0.0104f
C6489 VDD.n4322 VSS 3.16e-19
C6490 VDD.n4323 VSS 0.00348f
C6491 VDD.n4324 VSS 4.74e-19
C6492 VDD.n4325 VSS 0.00332f
C6493 VDD.n4326 VSS 0.00439f
C6494 VDD.n4327 VSS 0.0138f
C6495 VDD.n4328 VSS 0.0225f
C6496 VDD.n4329 VSS -0.174f
C6497 VDD.n4330 VSS 0.00798f
C6498 VDD.n4331 VSS 0.00488f
C6499 VDD.n4332 VSS 4.74e-19
C6500 VDD.n4333 VSS 0.0422f
C6501 VDD.n4334 VSS 0.0389f
C6502 VDD.n4335 VSS 0.0398f
C6503 VDD.n4336 VSS 0.0143f
C6504 VDD.n4337 VSS 0.14f
C6505 VDD.n4338 VSS 0.0439f
C6506 VDD.n4339 VSS 0.0433f
C6507 VDD.n4340 VSS 0.0576f
C6508 VDD.n4341 VSS 0.0314f
C6509 VDD.n4342 VSS 0.00269f
C6510 VDD.n4343 VSS 0.00277f
C6511 VDD.n4344 VSS 0.0527f
C6512 VDD.n4345 VSS 0.245f
C6513 VDD.n4346 VSS 0.198f
C6514 VDD.n4347 VSS 0.0104f
C6515 VDD.n4348 VSS 3.16e-19
C6516 VDD.n4349 VSS 0.00348f
C6517 VDD.n4350 VSS 0.00916f
C6518 VDD.n4351 VSS 0.00411f
C6519 VDD.n4352 VSS 0.00585f
C6520 VDD.n4353 VSS 0.00472f
C6521 VDD.n4354 VSS 0.00374f
C6522 VDD.n4355 VSS 0.00798f
C6523 VDD.n4356 VSS -0.174f
C6524 VDD.n4357 VSS -0.0841f
C6525 VDD.n4358 VSS 0.014f
C6526 VDD.n4359 VSS 0.00439f
C6527 VDD.n4360 VSS 0.00332f
C6528 VDD.n4361 VSS 0.00411f
C6529 VDD.n4362 VSS 0.00916f
C6530 VDD.n4363 VSS 0.00663f
C6531 VDD.n4364 VSS 0.00806f
C6532 VDD.n4365 VSS 0.00348f
C6533 VDD.n4366 VSS 0.00269f
C6534 VDD.n4367 VSS 0.00348f
C6535 VDD.n4368 VSS 3.16e-19
C6536 VDD.n4369 VSS 0.00269f
C6537 VDD.n4370 VSS 0.00277f
C6538 VDD.n4371 VSS 0.0527f
C6539 VDD.n4372 VSS 0.245f
C6540 VDD.n4373 VSS 0.198f
C6541 VDD.n4374 VSS 0.0104f
C6542 VDD.n4375 VSS 3.16e-19
C6543 VDD.n4376 VSS 0.00348f
C6544 VDD.n4377 VSS 0.00916f
C6545 VDD.n4378 VSS 0.00411f
C6546 VDD.n4379 VSS 0.00585f
C6547 VDD.n4380 VSS 0.00472f
C6548 VDD.n4381 VSS 0.00374f
C6549 VDD.n4382 VSS 0.00798f
C6550 VDD.n4383 VSS -0.174f
C6551 VDD.n4384 VSS -0.0841f
C6552 VDD.n4385 VSS 0.014f
C6553 VDD.n4386 VSS 0.00439f
C6554 VDD.n4387 VSS 0.00472f
C6555 VDD.n4388 VSS 0.00779f
C6556 VDD.n4389 VSS 0.0122f
C6557 VDD.n4390 VSS 0.00618f
C6558 VDD.n4391 VSS 0.0111f
C6559 VDD.n4392 VSS 0.00106f
C6560 VDD.n4393 VSS 0.113f
C6561 VDD.n4394 VSS 0.331f
C6562 VDD.n4395 VSS 0.261f
C6563 VDD.n4396 VSS 0.0389f
C6564 VDD.n4397 VSS 0.0398f
C6565 VDD.n4398 VSS 0.0607f
C6566 VDD.n4399 VSS 0.0142f
C6567 VDD.n4400 VSS -0.078f
C6568 VDD.n4401 VSS 3.26e-19
C6569 VDD.n4402 VSS 0.00472f
C6570 VDD.n4403 VSS 4.74e-19
C6571 VDD.n4404 VSS 0.00348f
C6572 VDD.n4405 VSS 0.00269f
C6573 VDD.n4406 VSS 0.00332f
C6574 VDD.n4407 VSS 0.00979f
C6575 VDD.n4408 VSS 0.00979f
C6576 VDD.n4409 VSS 0.0129f
C6577 VDD.n4410 VSS 0.245f
C6578 VDD.n4411 VSS 0.0527f
C6579 VDD.n4412 VSS 0.198f
C6580 VDD.n4413 VSS 0.0104f
C6581 VDD.n4414 VSS 3.16e-19
C6582 VDD.n4415 VSS 0.00348f
C6583 VDD.n4416 VSS 4.74e-19
C6584 VDD.n4417 VSS 0.00472f
C6585 VDD.n4418 VSS 0.00781f
C6586 VDD.n4419 VSS 0.00391f
C6587 VDD.n4420 VSS 0.023f
C6588 VDD.n4421 VSS 0.0142f
C6589 VDD.n4422 VSS 0.0138f
C6590 VDD.n4423 VSS 3.26e-19
C6591 VDD.n4424 VSS 0.00472f
C6592 VDD.n4425 VSS 4.74e-19
C6593 VDD.n4426 VSS 0.00348f
C6594 VDD.n4427 VSS 0.00269f
C6595 VDD.n4428 VSS 0.00332f
C6596 VDD.n4429 VSS 0.00979f
C6597 VDD.n4430 VSS 0.00979f
C6598 VDD.n4431 VSS 0.0129f
C6599 VDD.n4432 VSS 0.245f
C6600 VDD.n4433 VSS 0.0527f
C6601 VDD.n4434 VSS 0.198f
C6602 VDD.n4435 VSS 0.0104f
C6603 VDD.n4436 VSS 3.16e-19
C6604 VDD.n4437 VSS 0.00348f
C6605 VDD.n4438 VSS 4.74e-19
C6606 VDD.n4439 VSS 0.00472f
C6607 VDD.n4440 VSS 0.00781f
C6608 VDD.n4441 VSS 0.00391f
C6609 VDD.n4442 VSS 0.023f
C6610 VDD.n4443 VSS 0.0142f
C6611 VDD.n4444 VSS 0.0138f
C6612 VDD.n4445 VSS 3.26e-19
C6613 VDD.n4446 VSS 0.00472f
C6614 VDD.n4447 VSS 4.74e-19
C6615 VDD.n4448 VSS 0.00348f
C6616 VDD.n4449 VSS 0.00269f
C6617 VDD.n4450 VSS 0.00332f
C6618 VDD.n4451 VSS 0.00979f
C6619 VDD.n4452 VSS 0.00979f
C6620 VDD.n4453 VSS 0.0129f
C6621 VDD.n4454 VSS 0.245f
C6622 VDD.n4455 VSS 0.0527f
C6623 VDD.n4456 VSS 0.124f
C6624 VDD.n4457 VSS 0.0236f
C6625 VDD.n4458 VSS 3.16e-19
C6626 VDD.n4459 VSS 0.00348f
C6627 VDD.n4460 VSS 4.74e-19
C6628 VDD.n4461 VSS 0.00472f
C6629 VDD.n4462 VSS 0.0285f
C6630 VDD.n4463 VSS 0.0286f
C6631 VDD.n4464 VSS 0.0813f
C6632 VDD.n4465 VSS 0.0142f
C6633 VDD.n4466 VSS 0.0138f
C6634 VDD.n4467 VSS -0.0753f
C6635 VDD.n4468 VSS 0.00332f
C6636 VDD.n4469 VSS 0.00411f
C6637 VDD.n4470 VSS 0.00916f
C6638 VDD.n4471 VSS 0.00663f
C6639 VDD.n4472 VSS 0.00806f
C6640 VDD.n4473 VSS 0.00348f
C6641 VDD.n4474 VSS 0.00269f
C6642 VDD.n4475 VSS 0.00348f
C6643 VDD.n4476 VSS 3.16e-19
C6644 VDD.n4477 VSS 0.00269f
C6645 VDD.n4478 VSS 0.00277f
C6646 VDD.n4479 VSS 0.0527f
C6647 VDD.n4480 VSS 0.245f
C6648 VDD.n4481 VSS 0.198f
C6649 VDD.n4482 VSS 0.0104f
C6650 VDD.n4483 VSS 3.16e-19
C6651 VDD.n4484 VSS 0.00348f
C6652 VDD.n4485 VSS 0.00916f
C6653 VDD.n4486 VSS 0.00411f
C6654 VDD.n4487 VSS 0.00585f
C6655 VDD.n4488 VSS 0.00472f
C6656 VDD.n4489 VSS 0.00374f
C6657 VDD.n4490 VSS 0.00798f
C6658 VDD.n4491 VSS 0.023f
C6659 VDD.n4492 VSS 0.0142f
C6660 VDD.n4493 VSS 0.0138f
C6661 VDD.n4494 VSS -0.0753f
C6662 VDD.n4495 VSS 0.00332f
C6663 VDD.n4496 VSS 0.00411f
C6664 VDD.n4497 VSS 0.00916f
C6665 VDD.n4498 VSS 0.00663f
C6666 VDD.n4499 VSS 0.00806f
C6667 VDD.n4500 VSS 0.00348f
C6668 VDD.n4501 VSS 0.00269f
C6669 VDD.n4502 VSS 0.00348f
C6670 VDD.n4503 VSS 3.16e-19
C6671 VDD.n4504 VSS 0.00269f
C6672 VDD.n4505 VSS 0.00277f
C6673 VDD.n4506 VSS 0.0527f
C6674 VDD.n4507 VSS 0.245f
C6675 VDD.n4508 VSS 0.198f
C6676 VDD.n4509 VSS 0.0104f
C6677 VDD.n4510 VSS 3.16e-19
C6678 VDD.n4511 VSS 0.00348f
C6679 VDD.n4512 VSS 4.74e-19
C6680 VDD.n4513 VSS 0.00332f
C6681 VDD.n4514 VSS 0.00439f
C6682 VDD.n4515 VSS 0.0138f
C6683 VDD.n4516 VSS 0.0142f
C6684 VDD.n4517 VSS 0.0241f
C6685 VDD.n4518 VSS 0.0243f
C6686 VDD.n4519 VSS 0.0607f
C6687 VDD.n4520 VSS 0.0142f
C6688 VDD.n4521 VSS -0.078f
C6689 VDD.n4522 VSS 3.26e-19
C6690 VDD.n4523 VSS 0.00472f
C6691 VDD.n4524 VSS 4.74e-19
C6692 VDD.n4525 VSS 0.00348f
C6693 VDD.n4526 VSS 0.00269f
C6694 VDD.n4527 VSS 0.00332f
C6695 VDD.n4528 VSS 0.00979f
C6696 VDD.n4529 VSS 0.00979f
C6697 VDD.n4530 VSS 0.0129f
C6698 VDD.n4531 VSS 0.245f
C6699 VDD.n4532 VSS 0.0527f
C6700 VDD.n4533 VSS 0.198f
C6701 VDD.n4534 VSS 0.0104f
C6702 VDD.n4535 VSS 3.16e-19
C6703 VDD.n4536 VSS 0.00348f
C6704 VDD.n4537 VSS 4.74e-19
C6705 VDD.n4538 VSS 0.00472f
C6706 VDD.n4539 VSS 0.00781f
C6707 VDD.n4540 VSS 0.00391f
C6708 VDD.n4541 VSS 0.023f
C6709 VDD.n4542 VSS 0.0142f
C6710 VDD.n4543 VSS 0.0138f
C6711 VDD.n4544 VSS 3.26e-19
C6712 VDD.n4545 VSS 0.00472f
C6713 VDD.n4546 VSS 4.74e-19
C6714 VDD.n4547 VSS 0.00348f
C6715 VDD.n4548 VSS 0.00269f
C6716 VDD.n4549 VSS 0.00332f
C6717 VDD.n4550 VSS 0.00979f
C6718 VDD.n4551 VSS 0.00979f
C6719 VDD.n4552 VSS 0.0129f
C6720 VDD.n4553 VSS 0.245f
C6721 VDD.n4554 VSS 0.0527f
C6722 VDD.n4555 VSS 0.198f
C6723 VDD.n4556 VSS 0.0104f
C6724 VDD.n4557 VSS 3.16e-19
C6725 VDD.n4558 VSS 0.00348f
C6726 VDD.n4559 VSS 4.74e-19
C6727 VDD.n4560 VSS 0.00472f
C6728 VDD.n4561 VSS 0.00781f
C6729 VDD.n4562 VSS 0.00391f
C6730 VDD.n4563 VSS 0.023f
C6731 VDD.n4564 VSS 0.0142f
C6732 VDD.n4565 VSS 0.0138f
C6733 VDD.n4566 VSS 3.26e-19
C6734 VDD.n4567 VSS 0.00472f
C6735 VDD.n4568 VSS 4.74e-19
C6736 VDD.n4569 VSS 0.00348f
C6737 VDD.n4570 VSS 0.00269f
C6738 VDD.n4571 VSS 0.00332f
C6739 VDD.n4572 VSS 0.00979f
C6740 VDD.n4573 VSS 0.00979f
C6741 VDD.n4574 VSS 0.0129f
C6742 VDD.n4575 VSS 0.245f
C6743 VDD.n4576 VSS 0.0527f
C6744 VDD.n4577 VSS 0.124f
C6745 VDD.n4578 VSS 0.0236f
C6746 VDD.n4579 VSS 3.16e-19
C6747 VDD.n4580 VSS 0.00348f
C6748 VDD.n4581 VSS 4.74e-19
C6749 VDD.n4582 VSS 0.00472f
C6750 VDD.n4583 VSS 0.0285f
C6751 VDD.n4584 VSS 0.0286f
C6752 VDD.n4585 VSS 0.0813f
C6753 VDD.n4586 VSS 0.0142f
C6754 VDD.n4587 VSS 0.0138f
C6755 VDD.n4588 VSS -0.0753f
C6756 VDD.n4589 VSS 0.00332f
C6757 VDD.n4590 VSS 0.00411f
C6758 VDD.n4591 VSS 0.00916f
C6759 VDD.n4592 VSS 0.00663f
C6760 VDD.n4593 VSS 0.00806f
C6761 VDD.n4594 VSS 0.00348f
C6762 VDD.n4595 VSS 0.00269f
C6763 VDD.n4596 VSS 0.00348f
C6764 VDD.n4597 VSS 3.16e-19
C6765 VDD.n4598 VSS 0.00269f
C6766 VDD.n4599 VSS 0.00277f
C6767 VDD.n4600 VSS 0.0527f
C6768 VDD.n4601 VSS 0.245f
C6769 VDD.n4602 VSS 0.198f
C6770 VDD.n4603 VSS 0.0104f
C6771 VDD.n4604 VSS 3.16e-19
C6772 VDD.n4605 VSS 0.00348f
C6773 VDD.n4606 VSS 0.00916f
C6774 VDD.n4607 VSS 0.00411f
C6775 VDD.n4608 VSS 0.00585f
C6776 VDD.n4609 VSS 0.00472f
C6777 VDD.n4610 VSS 0.00374f
C6778 VDD.n4611 VSS 0.00798f
C6779 VDD.n4612 VSS 0.023f
C6780 VDD.n4613 VSS 0.0142f
C6781 VDD.n4614 VSS 0.0138f
C6782 VDD.n4615 VSS -0.0753f
C6783 VDD.n4616 VSS 0.00332f
C6784 VDD.n4617 VSS 0.00411f
C6785 VDD.n4618 VSS 0.00916f
C6786 VDD.n4619 VSS 0.00663f
C6787 VDD.n4620 VSS 0.00806f
C6788 VDD.n4621 VSS 0.00348f
C6789 VDD.n4622 VSS 0.00269f
C6790 VDD.n4623 VSS 0.00348f
C6791 VDD.n4624 VSS 3.16e-19
C6792 VDD.n4625 VSS 0.00269f
C6793 VDD.n4626 VSS 0.00277f
C6794 VDD.n4627 VSS 0.0527f
C6795 VDD.n4628 VSS 0.245f
C6796 VDD.n4629 VSS 0.198f
C6797 VDD.n4630 VSS 0.0104f
C6798 VDD.n4631 VSS 3.16e-19
C6799 VDD.n4632 VSS 0.00348f
C6800 VDD.n4633 VSS 4.74e-19
C6801 VDD.n4634 VSS 0.00332f
C6802 VDD.n4635 VSS 0.00439f
C6803 VDD.n4636 VSS 0.0138f
C6804 VDD.n4637 VSS 0.0142f
C6805 VDD.n4638 VSS 0.0241f
C6806 VDD.n4639 VSS 0.0243f
C6807 VDD.n4640 VSS 0.0607f
C6808 VDD.n4641 VSS 0.0142f
C6809 VDD.n4642 VSS -0.078f
C6810 VDD.n4643 VSS 3.26e-19
C6811 VDD.n4644 VSS 0.00472f
C6812 VDD.n4645 VSS 4.74e-19
C6813 VDD.n4646 VSS 0.00348f
C6814 VDD.n4647 VSS 0.00269f
C6815 VDD.n4648 VSS 0.00332f
C6816 VDD.n4649 VSS 0.00979f
C6817 VDD.n4650 VSS 0.00979f
C6818 VDD.n4651 VSS 0.0129f
C6819 VDD.n4652 VSS 0.245f
C6820 VDD.n4653 VSS 0.0527f
C6821 VDD.n4654 VSS 0.198f
C6822 VDD.n4655 VSS 0.0104f
C6823 VDD.n4656 VSS 3.16e-19
C6824 VDD.n4657 VSS 0.00348f
C6825 VDD.n4658 VSS 4.74e-19
C6826 VDD.n4659 VSS 0.00472f
C6827 VDD.n4660 VSS 0.00781f
C6828 VDD.n4661 VSS 0.00391f
C6829 VDD.n4662 VSS 0.023f
C6830 VDD.n4663 VSS 0.0142f
C6831 VDD.n4664 VSS 0.0138f
C6832 VDD.n4665 VSS 3.26e-19
C6833 VDD.n4666 VSS 0.00472f
C6834 VDD.n4667 VSS 4.74e-19
C6835 VDD.n4668 VSS 0.00348f
C6836 VDD.n4669 VSS 0.00269f
C6837 VDD.n4670 VSS 0.00332f
C6838 VDD.n4671 VSS 0.00979f
C6839 VDD.n4672 VSS 0.00979f
C6840 VDD.n4673 VSS 0.0129f
C6841 VDD.n4674 VSS 0.245f
C6842 VDD.n4675 VSS 0.0527f
C6843 VDD.n4676 VSS 0.198f
C6844 VDD.n4677 VSS 0.0104f
C6845 VDD.n4678 VSS 3.16e-19
C6846 VDD.n4679 VSS 0.00348f
C6847 VDD.n4680 VSS 4.74e-19
C6848 VDD.n4681 VSS 0.00472f
C6849 VDD.n4682 VSS 0.00781f
C6850 VDD.n4683 VSS 0.00391f
C6851 VDD.n4684 VSS 0.023f
C6852 VDD.n4685 VSS 0.0142f
C6853 VDD.n4686 VSS 0.0138f
C6854 VDD.n4687 VSS 3.26e-19
C6855 VDD.n4688 VSS 0.00472f
C6856 VDD.n4689 VSS 4.74e-19
C6857 VDD.n4690 VSS 0.00348f
C6858 VDD.n4691 VSS 0.00269f
C6859 VDD.n4692 VSS 0.00332f
C6860 VDD.n4693 VSS 0.00979f
C6861 VDD.n4694 VSS 0.00979f
C6862 VDD.n4695 VSS 0.0129f
C6863 VDD.n4696 VSS 0.245f
C6864 VDD.n4697 VSS 0.0527f
C6865 VDD.n4698 VSS 0.124f
C6866 VDD.n4699 VSS 0.0236f
C6867 VDD.n4700 VSS 3.16e-19
C6868 VDD.n4701 VSS 0.00348f
C6869 VDD.n4702 VSS 4.74e-19
C6870 VDD.n4703 VSS 0.00472f
C6871 VDD.n4704 VSS 0.0285f
C6872 VDD.n4705 VSS 0.0286f
C6873 VDD.n4706 VSS 0.0813f
C6874 VDD.n4707 VSS 0.0142f
C6875 VDD.n4708 VSS 0.0138f
C6876 VDD.n4709 VSS -0.0753f
C6877 VDD.n4710 VSS 0.00332f
C6878 VDD.n4711 VSS 0.00411f
C6879 VDD.n4712 VSS 0.00916f
C6880 VDD.n4713 VSS 0.00663f
C6881 VDD.n4714 VSS 0.00806f
C6882 VDD.n4715 VSS 0.00348f
C6883 VDD.n4716 VSS 0.00269f
C6884 VDD.n4717 VSS 0.00348f
C6885 VDD.n4718 VSS 3.16e-19
C6886 VDD.n4719 VSS 0.00269f
C6887 VDD.n4720 VSS 0.00277f
C6888 VDD.n4721 VSS 0.0527f
C6889 VDD.n4722 VSS 0.245f
C6890 VDD.n4723 VSS 0.198f
C6891 VDD.n4724 VSS 0.0104f
C6892 VDD.n4725 VSS 3.16e-19
C6893 VDD.n4726 VSS 0.00348f
C6894 VDD.n4727 VSS 0.00916f
C6895 VDD.n4728 VSS 0.00411f
C6896 VDD.n4729 VSS 0.00585f
C6897 VDD.n4730 VSS 0.00472f
C6898 VDD.n4731 VSS 0.00374f
C6899 VDD.n4732 VSS 0.00798f
C6900 VDD.n4733 VSS 0.023f
C6901 VDD.n4734 VSS 0.0142f
C6902 VDD.n4735 VSS 0.0138f
C6903 VDD.n4736 VSS -0.0753f
C6904 VDD.n4737 VSS 0.00332f
C6905 VDD.n4738 VSS 0.00411f
C6906 VDD.n4739 VSS 0.00916f
C6907 VDD.n4740 VSS 0.00663f
C6908 VDD.n4741 VSS 0.00806f
C6909 VDD.n4742 VSS 0.00348f
C6910 VDD.n4743 VSS 0.00269f
C6911 VDD.n4744 VSS 0.00348f
C6912 VDD.n4745 VSS 3.16e-19
C6913 VDD.n4746 VSS 0.00269f
C6914 VDD.n4747 VSS 0.00277f
C6915 VDD.n4748 VSS 0.0527f
C6916 VDD.n4749 VSS 0.245f
C6917 VDD.n4750 VSS 0.198f
C6918 VDD.n4751 VSS 0.0104f
C6919 VDD.n4752 VSS 3.16e-19
C6920 VDD.n4753 VSS 0.00348f
C6921 VDD.n4754 VSS 4.74e-19
C6922 VDD.n4755 VSS 0.00332f
C6923 VDD.n4756 VSS 0.00439f
C6924 VDD.n4757 VSS 0.0138f
C6925 VDD.n4758 VSS 0.0142f
C6926 VDD.n4759 VSS 0.0241f
C6927 VDD.n4760 VSS 0.0243f
C6928 VDD.n4761 VSS 0.0607f
C6929 VDD.n4762 VSS 0.0142f
C6930 VDD.n4763 VSS -0.078f
C6931 VDD.n4764 VSS 3.26e-19
C6932 VDD.n4765 VSS 0.00472f
C6933 VDD.n4766 VSS 4.74e-19
C6934 VDD.n4767 VSS 0.00348f
C6935 VDD.n4768 VSS 0.00269f
C6936 VDD.n4769 VSS 0.00332f
C6937 VDD.n4770 VSS 0.00979f
C6938 VDD.n4771 VSS 0.00979f
C6939 VDD.n4772 VSS 0.0129f
C6940 VDD.n4773 VSS 0.245f
C6941 VDD.n4774 VSS 0.0527f
C6942 VDD.n4775 VSS 0.198f
C6943 VDD.n4776 VSS 0.0104f
C6944 VDD.n4777 VSS 3.16e-19
C6945 VDD.n4778 VSS 0.00348f
C6946 VDD.n4779 VSS 4.74e-19
C6947 VDD.n4780 VSS 0.00472f
C6948 VDD.n4781 VSS 0.00781f
C6949 VDD.n4782 VSS 0.00391f
C6950 VDD.n4783 VSS 0.023f
C6951 VDD.n4784 VSS 0.0142f
C6952 VDD.n4785 VSS 0.0138f
C6953 VDD.n4786 VSS 3.26e-19
C6954 VDD.n4787 VSS 0.00472f
C6955 VDD.n4788 VSS 4.74e-19
C6956 VDD.n4789 VSS 0.00348f
C6957 VDD.n4790 VSS 0.00269f
C6958 VDD.n4791 VSS 0.00332f
C6959 VDD.n4792 VSS 0.00979f
C6960 VDD.n4793 VSS 0.00979f
C6961 VDD.n4794 VSS 0.0129f
C6962 VDD.n4795 VSS 0.245f
C6963 VDD.n4796 VSS 0.0527f
C6964 VDD.n4797 VSS 0.198f
C6965 VDD.n4798 VSS 0.0104f
C6966 VDD.n4799 VSS 3.16e-19
C6967 VDD.n4800 VSS 0.00348f
C6968 VDD.n4801 VSS 4.74e-19
C6969 VDD.n4802 VSS 0.00472f
C6970 VDD.n4803 VSS 0.00781f
C6971 VDD.n4804 VSS 0.00391f
C6972 VDD.n4805 VSS 0.023f
C6973 VDD.n4806 VSS 0.0142f
C6974 VDD.n4807 VSS 0.0138f
C6975 VDD.n4808 VSS 3.26e-19
C6976 VDD.n4809 VSS 0.00472f
C6977 VDD.n4810 VSS 4.74e-19
C6978 VDD.n4811 VSS 0.00348f
C6979 VDD.n4812 VSS 0.00269f
C6980 VDD.n4813 VSS 0.00332f
C6981 VDD.n4814 VSS 0.00979f
C6982 VDD.n4815 VSS 0.00979f
C6983 VDD.n4816 VSS 0.0129f
C6984 VDD.n4817 VSS 0.245f
C6985 VDD.n4818 VSS 0.0527f
C6986 VDD.n4819 VSS 0.124f
C6987 VDD.n4820 VSS 0.0236f
C6988 VDD.n4821 VSS 3.16e-19
C6989 VDD.n4822 VSS 0.00348f
C6990 VDD.n4823 VSS 4.74e-19
C6991 VDD.n4824 VSS 0.00472f
C6992 VDD.n4825 VSS 0.0285f
C6993 VDD.n4826 VSS 0.0286f
C6994 VDD.n4827 VSS 0.0813f
C6995 VDD.n4828 VSS 0.0142f
C6996 VDD.n4829 VSS 0.0138f
C6997 VDD.n4830 VSS -0.0753f
C6998 VDD.n4831 VSS 0.00332f
C6999 VDD.n4832 VSS 0.00411f
C7000 VDD.n4833 VSS 0.00916f
C7001 VDD.n4834 VSS 0.00663f
C7002 VDD.n4835 VSS 0.00806f
C7003 VDD.n4836 VSS 0.00348f
C7004 VDD.n4837 VSS 0.00269f
C7005 VDD.n4838 VSS 0.00348f
C7006 VDD.n4839 VSS 3.16e-19
C7007 VDD.n4840 VSS 0.00269f
C7008 VDD.n4841 VSS 0.00277f
C7009 VDD.n4842 VSS 0.0527f
C7010 VDD.n4843 VSS 0.245f
C7011 VDD.n4844 VSS 0.198f
C7012 VDD.n4845 VSS 0.0104f
C7013 VDD.n4846 VSS 3.16e-19
C7014 VDD.n4847 VSS 0.00348f
C7015 VDD.n4848 VSS 0.00916f
C7016 VDD.n4849 VSS 0.00411f
C7017 VDD.n4850 VSS 0.00585f
C7018 VDD.n4851 VSS 0.00472f
C7019 VDD.n4852 VSS 0.00374f
C7020 VDD.n4853 VSS 0.00798f
C7021 VDD.n4854 VSS 0.023f
C7022 VDD.n4855 VSS 0.0142f
C7023 VDD.n4856 VSS 0.0138f
C7024 VDD.n4857 VSS -0.0753f
C7025 VDD.n4858 VSS 0.00332f
C7026 VDD.n4859 VSS 0.00411f
C7027 VDD.n4860 VSS 0.00916f
C7028 VDD.n4861 VSS 0.00663f
C7029 VDD.n4862 VSS 0.00806f
C7030 VDD.n4863 VSS 0.00348f
C7031 VDD.n4864 VSS 0.00269f
C7032 VDD.n4865 VSS 0.00348f
C7033 VDD.n4866 VSS 3.16e-19
C7034 VDD.n4867 VSS 0.00269f
C7035 VDD.n4868 VSS 0.00277f
C7036 VDD.n4869 VSS 0.0527f
C7037 VDD.n4870 VSS 0.245f
C7038 VDD.n4871 VSS 0.198f
C7039 VDD.n4872 VSS 0.0104f
C7040 VDD.n4873 VSS 0.0418f
C7041 VDD.n4874 VSS 0.0422f
C7042 VDD.n4875 VSS 0.0389f
C7043 VDD.n4876 VSS 0.0398f
C7044 VDD.n4877 VSS 0.0143f
C7045 VDD.n4878 VSS 0.0439f
C7046 VDD.n4879 VSS 0.14f
C7047 VDD.n4880 VSS 0.0145f
C7048 VDD.n4881 VSS 0.014f
C7049 VDD.n4882 VSS -0.0753f
C7050 VDD.n4883 VSS 0.00332f
C7051 VDD.n4884 VSS 0.00411f
C7052 VDD.n4885 VSS 0.0095f
C7053 VDD.n4886 VSS 0.00663f
C7054 VDD.n4887 VSS 0.00806f
C7055 VDD.n4888 VSS 0.00348f
C7056 VDD.n4889 VSS 0.00269f
C7057 VDD.n4890 VSS 0.00348f
C7058 VDD.n4891 VSS 3.16e-19
C7059 VDD.n4892 VSS 0.00269f
C7060 VDD.n4893 VSS 0.00277f
C7061 VDD.n4894 VSS 0.0527f
C7062 VDD.n4895 VSS 0.245f
C7063 VDD.n4896 VSS 0.198f
C7064 VDD.n4897 VSS 0.0104f
C7065 VDD.n4898 VSS 3.16e-19
C7066 VDD.n4899 VSS 0.00348f
C7067 VDD.n4900 VSS 0.00916f
C7068 VDD.n4901 VSS 0.00411f
C7069 VDD.n4902 VSS 0.00585f
C7070 VDD.n4903 VSS 0.00472f
C7071 VDD.n4904 VSS 0.00374f
C7072 VDD.n4905 VSS 0.00798f
C7073 VDD.n4906 VSS 0.0233f
C7074 VDD.n4907 VSS 0.0145f
C7075 VDD.n4908 VSS 0.014f
C7076 VDD.n4909 VSS -0.0753f
C7077 VDD.n4910 VSS 0.00332f
C7078 VDD.n4911 VSS 0.00411f
C7079 VDD.n4912 VSS 0.00916f
C7080 VDD.n4913 VSS 0.00663f
C7081 VDD.n4914 VSS 0.00806f
C7082 VDD.n4915 VSS 0.00348f
C7083 VDD.n4916 VSS 0.00269f
C7084 VDD.n4917 VSS 0.00348f
C7085 VDD.n4918 VSS 3.16e-19
C7086 VDD.n4919 VSS 0.00269f
C7087 VDD.n4920 VSS 0.00277f
C7088 VDD.n4921 VSS 0.0527f
C7089 VDD.n4922 VSS 0.245f
C7090 VDD.n4923 VSS 0.198f
C7091 VDD.n4924 VSS 0.0104f
C7092 VDD.n4925 VSS 3.16e-19
C7093 VDD.n4926 VSS 0.00302f
C7094 VDD.n4927 VSS 0.0087f
C7095 VDD.n4928 VSS 0.0186f
C7096 VDD.n4929 VSS 0.102f
C7097 VDD.n4930 VSS 0.442f
C7098 VDD.t23 VSS 0.797f
C7099 VDD.n4931 VSS 0.0931f
C7100 VDD.n4932 VSS 0.0313f
C7101 VDD.n4933 VSS 0.00256f
C7102 VDD.n4934 VSS 0.00483f
C7103 VDD.n4935 VSS 0.00414f
C7104 VDD.n4936 VSS 0.00443f
C7105 VDD.n4937 VSS 0.00689f
C7106 VDD.n4938 VSS 8.15e-19
C7107 VDD.n4939 VSS 0.0185f
C7108 VDD.n4940 VSS 0.0409f
C7109 VDD.n4941 VSS 0.0186f
C7110 VDD.n4942 VSS 0.017f
C7111 VDD.n4943 VSS 0.0069f
C7112 VDD.n4944 VSS 0.0069f
C7113 VDD.n4945 VSS 0.0124f
C7114 VDD.n4946 VSS 0.0111f
C7115 VDD.n4947 VSS 0.00571f
C7116 VDD.n4948 VSS 0.02f
C7117 VDD.n4949 VSS 0.0261f
C7118 VDD.n4950 VSS 0.0604f
C7119 VDD.n4951 VSS 0.0274f
C7120 VDD.n4952 VSS 0.0198f
C7121 VDD.n4953 VSS 0.0211f
C7122 VDD.n4954 VSS 0.0108f
C7123 VDD.t49 VSS 0.0509f
C7124 VDD.n4955 VSS 0.0233f
C7125 VDD.n4956 VSS 0.056f
C7126 VDD.n4957 VSS 0.00797f
C7127 VDD.n4958 VSS 0.0106f
C7128 VDD.n4959 VSS 0.0207f
C7129 VDD.n4960 VSS 0.00758f
C7130 VDD.n4961 VSS 0.0039f
C7131 VDD.n4962 VSS 0.00461f
C7132 VDD.n4963 VSS 0.00391f
C7133 VDD.n4964 VSS 0.00184f
C7134 VDD.n4965 VSS 0.00135f
C7135 VDD.n4966 VSS 0.014f
C7136 VDD.n4967 VSS 0.0914f
C7137 VDD.n4968 VSS 0.0149f
C7138 VDD.n4969 VSS 0.0755f
C7139 VDD.n4970 VSS 0.0124f
C7140 VDD.n4971 VSS 0.0109f
C7141 VDD.n4972 VSS 0.00997f
C7142 VDD.n4973 VSS 0.0262f
C7143 VDD.n4974 VSS 0.0172f
C7144 VDD.n4975 VSS 0.0197f
C7145 VDD.n4976 VSS 8.15e-19
C7146 VDD.n4977 VSS 0.0124f
C7147 VDD.n4978 VSS 0.613f
C7148 VDD.n4979 VSS 4.85f
C7149 VDD.n4980 VSS 8.83f
C7150 VDD.n4981 VSS 0.444f
C7151 VDD.n4982 VSS 0.298f
C7152 VDD.n4983 VSS 0.02f
C7153 VDD.n4984 VSS 0.00824f
C7154 VDD.n4985 VSS 0.02f
C7155 VDD.n4986 VSS 0.00634f
C7156 VDD.n4987 VSS 0.00818f
C7157 VDD.n4988 VSS 0.0813f
C7158 VDD.n4989 VSS 1.26f
C7159 VDD.n4990 VSS 1.83f
C7160 VDD.t9 VSS 1.75f
C7161 VDD.n4991 VSS 0.00824f
C7162 VDD.n4992 VSS 0.02f
C7163 VDD.n4993 VSS 0.02f
C7164 VDD.n4994 VSS 0.0109f
C7165 VDD.n4995 VSS 0.00634f
C7166 VDD.n4996 VSS 0.00818f
C7167 VDD.n4997 VSS 0.0813f
C7168 VDD.t21 VSS 0.428f
C7169 VDD.t22 VSS 0.896f
C7170 VDD.n4998 VSS 0.0156f
C7171 VDD.t26 VSS 2.21f
C7172 VDD.t62 VSS 6.67f
C7173 VDD.t14 VSS 5.45f
C7174 VDD.n4999 VSS 2.08f
C7175 VDD.t17 VSS 2.33f
C7176 VDD.n5000 VSS 2.08f
C7177 VDD.n5001 VSS 0.00824f
C7178 VDD.n5002 VSS 0.0813f
C7179 VDD.n5003 VSS 0.00818f
C7180 VDD.n5004 VSS 0.02f
C7181 VDD.n5005 VSS 0.0109f
C7182 VDD.n5006 VSS 0.067f
C7183 VDD.n5007 VSS 0.0777f
C7184 VDD.n5008 VSS 0.02f
C7185 VDD.n5009 VSS 0.00824f
C7186 VDD.n5010 VSS 0.0813f
C7187 VDD.n5011 VSS 0.00818f
C7188 VDD.n5012 VSS 0.02f
C7189 VDD.n5013 VSS 0.059f
C7190 VDD.n5014 VSS 0.126f
C7191 VDD.n5015 VSS 0.0199f
C7192 VDD.t63 VSS 0.00943f
C7193 VDD.n5016 VSS 0.136f
C7194 VDD.n5017 VSS 0.02f
C7195 VDD.n5018 VSS 0.174f
C7196 VDD.n5019 VSS 35.1f
C7197 VDD.n5020 VSS 0.0141f
C7198 VDD.n5021 VSS 0.0136f
C7199 VDD.n5022 VSS 0.00439f
C7200 VDD.n5023 VSS 0.0398f
C7201 VDD.n5024 VSS 0.0389f
C7202 VDD.n5025 VSS 0.0442f
C7203 VDD.n5026 VSS 0.0422f
C7204 VDD.n5027 VSS 4.74e-19
C7205 VDD.n5028 VSS 0.00488f
C7206 VDD.n5029 VSS 0.00798f
C7207 VDD.n5030 VSS -0.174f
C7208 VDD.n5031 VSS 0.0223f
C7209 VDD.n5032 VSS 0.0136f
C7210 VDD.n5033 VSS 0.00439f
C7211 VDD.n5034 VSS 0.00472f
C7212 VDD.n5035 VSS 0.00585f
C7213 VDD.n5036 VSS 0.00806f
C7214 VDD.n5037 VSS 0.00663f
C7215 VDD.n5038 VSS 0.00332f
C7216 VDD.n5039 VSS 0.00979f
C7217 VDD.n5040 VSS 0.00979f
C7218 VDD.n5041 VSS 0.0129f
C7219 VDD.n5043 VSS 0.00277f
C7220 VDD.n5045 VSS 0.0104f
C7221 VDD.n5046 VSS 3.16e-19
C7222 VDD.n5047 VSS 0.00348f
C7223 VDD.n5048 VSS 4.74e-19
C7224 VDD.n5049 VSS 0.00488f
C7225 VDD.n5050 VSS 0.00798f
C7226 VDD.n5051 VSS 0.0227f
C7227 VDD.n5052 VSS 0.0223f
C7228 VDD.n5053 VSS 0.0136f
C7229 VDD.n5054 VSS 0.00374f
C7230 VDD.n5055 VSS 0.0141f
C7231 VDD.n5056 VSS 0.0223f
C7232 VDD.n5057 VSS 0.0227f
C7233 VDD.n5058 VSS 0.00798f
C7234 VDD.n5059 VSS 0.00488f
C7235 VDD.n5060 VSS 0.00348f
C7236 VDD.n5061 VSS 4.74e-19
C7237 VDD.n5062 VSS 0.00332f
C7238 VDD.n5063 VSS -0.0753f
C7239 VDD.n5064 VSS -0.211f
C7240 VDD.n5065 VSS 0.00585f
C7241 VDD.n5066 VSS 0.00806f
C7242 VDD.n5067 VSS 0.00663f
C7243 VDD.n5068 VSS 0.00332f
C7244 VDD.n5069 VSS 0.00979f
C7245 VDD.n5070 VSS 0.00979f
C7246 VDD.n5071 VSS 0.00269f
C7247 VDD.n5072 VSS 0.00277f
C7248 VDD.n5074 VSS 0.0104f
C7249 VDD.n5076 VSS 0.0129f
C7250 VDD.n5077 VSS 0.00979f
C7251 VDD.n5078 VSS 0.00979f
C7252 VDD.n5079 VSS 0.00332f
C7253 VDD.n5080 VSS 0.00663f
C7254 VDD.n5081 VSS 0.00806f
C7255 VDD.n5082 VSS 0.00585f
C7256 VDD.n5083 VSS 0.00411f
C7257 VDD.n5084 VSS 0.00332f
C7258 VDD.n5085 VSS 0.00439f
C7259 VDD.n5086 VSS 3.26e-19
C7260 VDD.n5087 VSS 0.00488f
C7261 VDD.n5088 VSS 0.00798f
C7262 VDD.n5089 VSS -0.174f
C7263 VDD.n5090 VSS 0.0223f
C7264 VDD.n5091 VSS 0.0136f
C7265 VDD.n5092 VSS 0.00439f
C7266 VDD.n5093 VSS 0.00472f
C7267 VDD.n5094 VSS 0.00585f
C7268 VDD.n5095 VSS 0.00663f
C7269 VDD.n5096 VSS 0.00806f
C7270 VDD.n5097 VSS 0.00348f
C7271 VDD.n5098 VSS 0.00269f
C7272 VDD.n5099 VSS 0.00348f
C7273 VDD.n5100 VSS 3.16e-19
C7274 VDD.n5101 VSS 0.0104f
C7275 VDD.n5103 VSS 0.0129f
C7276 VDD.n5105 VSS 0.00277f
C7277 VDD.n5106 VSS 0.00269f
C7278 VDD.n5107 VSS 3.16e-19
C7279 VDD.n5108 VSS 0.00348f
C7280 VDD.n5109 VSS 4.74e-19
C7281 VDD.n5110 VSS 0.00488f
C7282 VDD.n5111 VSS 0.00798f
C7283 VDD.n5112 VSS 0.0227f
C7284 VDD.n5113 VSS 0.0223f
C7285 VDD.n5114 VSS 0.0141f
C7286 VDD.n5115 VSS 0.0136f
C7287 VDD.n5116 VSS -0.0753f
C7288 VDD.n5117 VSS -0.211f
C7289 VDD.n5118 VSS 0.00585f
C7290 VDD.n5119 VSS 0.00806f
C7291 VDD.n5120 VSS 0.00663f
C7292 VDD.n5121 VSS 0.00332f
C7293 VDD.n5122 VSS 0.00979f
C7294 VDD.n5123 VSS 0.00979f
C7295 VDD.n5124 VSS 0.0129f
C7296 VDD.n5126 VSS 0.00277f
C7297 VDD.n5127 VSS 0.0236f
C7298 VDD.n5128 VSS 3.16e-19
C7299 VDD.n5129 VSS 0.00348f
C7300 VDD.n5130 VSS 4.74e-19
C7301 VDD.n5131 VSS 0.00488f
C7302 VDD.n5132 VSS 0.0286f
C7303 VDD.n5133 VSS 0.00472f
C7304 VDD.n5134 VSS 0.0285f
C7305 VDD.n5135 VSS 0.08f
C7306 VDD.n5136 VSS 0.0136f
C7307 VDD.n5137 VSS 0.0223f
C7308 VDD.n5138 VSS 0.00472f
C7309 VDD.n5139 VSS 0.00781f
C7310 VDD.n5140 VSS 0.00391f
C7311 VDD.n5141 VSS 0.0227f
C7312 VDD.n5142 VSS 0.0141f
C7313 VDD.n5143 VSS -0.0753f
C7314 VDD.n5144 VSS 0.00332f
C7315 VDD.n5145 VSS 0.00411f
C7316 VDD.n5146 VSS 0.00916f
C7317 VDD.n5147 VSS 0.00663f
C7318 VDD.n5148 VSS 0.00806f
C7319 VDD.n5149 VSS 0.00348f
C7320 VDD.n5150 VSS 0.00269f
C7321 VDD.n5151 VSS 0.00269f
C7322 VDD.n5152 VSS 3.16e-19
C7323 VDD.n5153 VSS 0.0104f
C7324 VDD.n5155 VSS 0.00277f
C7325 VDD.n5157 VSS 0.0129f
C7326 VDD.n5158 VSS 0.00979f
C7327 VDD.n5159 VSS 0.00979f
C7328 VDD.n5160 VSS 0.00332f
C7329 VDD.n5161 VSS 0.00348f
C7330 VDD.n5162 VSS 0.00806f
C7331 VDD.n5163 VSS 0.00663f
C7332 VDD.n5164 VSS 0.00916f
C7333 VDD.n5165 VSS 0.00411f
C7334 VDD.n5166 VSS 0.00332f
C7335 VDD.n5167 VSS 0.00439f
C7336 VDD.n5168 VSS 0.0141f
C7337 VDD.n5169 VSS 0.0227f
C7338 VDD.n5170 VSS 0.00391f
C7339 VDD.n5171 VSS 0.00781f
C7340 VDD.n5172 VSS 0.00472f
C7341 VDD.n5173 VSS 3.26e-19
C7342 VDD.n5174 VSS -0.0782f
C7343 VDD.n5175 VSS 0.0141f
C7344 VDD.n5176 VSS 0.0227f
C7345 VDD.n5177 VSS 0.00391f
C7346 VDD.n5178 VSS 0.00488f
C7347 VDD.n5179 VSS 0.00585f
C7348 VDD.n5180 VSS 0.00411f
C7349 VDD.n5181 VSS 0.00916f
C7350 VDD.n5182 VSS 0.00348f
C7351 VDD.n5183 VSS 3.16e-19
C7352 VDD.n5184 VSS 0.00269f
C7353 VDD.n5185 VSS 0.00277f
C7354 VDD.n5187 VSS 0.0129f
C7355 VDD.n5189 VSS 0.0104f
C7356 VDD.n5190 VSS 3.16e-19
C7357 VDD.n5191 VSS 0.00348f
C7358 VDD.n5192 VSS 4.74e-19
C7359 VDD.n5193 VSS 0.00472f
C7360 VDD.n5194 VSS 3.26e-19
C7361 VDD.n5195 VSS 0.0136f
C7362 VDD.n5196 VSS 0.0141f
C7363 VDD.n5197 VSS 0.0223f
C7364 VDD.n5198 VSS 0.0227f
C7365 VDD.n5199 VSS 0.00391f
C7366 VDD.n5200 VSS -0.211f
C7367 VDD.n5201 VSS 0.00585f
C7368 VDD.n5202 VSS 0.00806f
C7369 VDD.n5203 VSS 0.00348f
C7370 VDD.n5204 VSS 0.00269f
C7371 VDD.n5205 VSS 0.00332f
C7372 VDD.n5206 VSS 0.00979f
C7373 VDD.n5207 VSS 0.00979f
C7374 VDD.n5208 VSS 0.0129f
C7375 VDD.n5210 VSS 0.0104f
C7376 VDD.n5212 VSS 0.00277f
C7377 VDD.n5213 VSS 0.00269f
C7378 VDD.n5214 VSS 0.00979f
C7379 VDD.n5215 VSS 0.00979f
C7380 VDD.n5216 VSS 0.00332f
C7381 VDD.n5217 VSS 0.00348f
C7382 VDD.n5218 VSS 0.00806f
C7383 VDD.n5219 VSS 0.00663f
C7384 VDD.n5220 VSS 0.00916f
C7385 VDD.n5221 VSS 0.00411f
C7386 VDD.n5222 VSS 0.00332f
C7387 VDD.n5223 VSS 0.00439f
C7388 VDD.n5224 VSS 0.0141f
C7389 VDD.n5225 VSS 0.0227f
C7390 VDD.n5226 VSS 0.00391f
C7391 VDD.n5227 VSS 0.00781f
C7392 VDD.n5228 VSS 0.00472f
C7393 VDD.n5229 VSS 3.26e-19
C7394 VDD.n5230 VSS -0.0782f
C7395 VDD.n5231 VSS 0.0141f
C7396 VDD.n5232 VSS 0.00472f
C7397 VDD.n5233 VSS 0.00439f
C7398 VDD.n5234 VSS 0.0136f
C7399 VDD.n5235 VSS 0.0141f
C7400 VDD.n5236 VSS 0.06f
C7401 VDD.n5237 VSS 0.0243f
C7402 VDD.n5238 VSS 0.00488f
C7403 VDD.n5239 VSS 0.0251f
C7404 VDD.n5240 VSS 0.00411f
C7405 VDD.n5241 VSS 0.0295f
C7406 VDD.n5242 VSS 0.00348f
C7407 VDD.n5243 VSS 3.16e-19
C7408 VDD.n5244 VSS 0.0104f
C7409 VDD.n5246 VSS 0.00277f
C7410 VDD.n5247 VSS 0.0186f
C7411 VDD.n5248 VSS 0.03f
C7412 VDD.n5249 VSS 0.0312f
C7413 VDD.n5250 VSS 0.0173f
C7414 VDD.n5251 VSS 0.00277f
C7415 VDD.n5252 VSS 0.00269f
C7416 VDD.n5253 VSS 3.16e-19
C7417 VDD.n5254 VSS 0.00348f
C7418 VDD.n5255 VSS 4.74e-19
C7419 VDD.n5256 VSS 0.00488f
C7420 VDD.n5257 VSS 0.00798f
C7421 VDD.n5258 VSS -0.174f
C7422 VDD.n5259 VSS 0.0223f
C7423 VDD.n5260 VSS 0.0136f
C7424 VDD.n5261 VSS 0.00439f
C7425 VDD.n5262 VSS 0.00472f
C7426 VDD.n5263 VSS 0.00585f
C7427 VDD.n5264 VSS 0.00806f
C7428 VDD.n5265 VSS 0.00663f
C7429 VDD.n5266 VSS 0.00332f
C7430 VDD.n5267 VSS 0.00979f
C7431 VDD.n5268 VSS 0.00979f
C7432 VDD.n5269 VSS 0.0129f
C7433 VDD.n5271 VSS 0.00277f
C7434 VDD.n5273 VSS 0.0104f
C7435 VDD.n5274 VSS 3.16e-19
C7436 VDD.n5275 VSS 0.00348f
C7437 VDD.n5276 VSS 4.74e-19
C7438 VDD.n5277 VSS 0.00488f
C7439 VDD.n5278 VSS 0.00798f
C7440 VDD.n5279 VSS 0.0227f
C7441 VDD.n5280 VSS 0.0223f
C7442 VDD.n5281 VSS 0.0136f
C7443 VDD.n5282 VSS 0.00374f
C7444 VDD.n5283 VSS 0.0141f
C7445 VDD.n5284 VSS 0.0223f
C7446 VDD.n5285 VSS 0.0227f
C7447 VDD.n5286 VSS 0.00798f
C7448 VDD.n5287 VSS 0.00488f
C7449 VDD.n5288 VSS 0.00348f
C7450 VDD.n5289 VSS 4.74e-19
C7451 VDD.n5290 VSS 0.00332f
C7452 VDD.n5291 VSS -0.0753f
C7453 VDD.n5292 VSS -0.211f
C7454 VDD.n5293 VSS 0.00585f
C7455 VDD.n5294 VSS 0.00806f
C7456 VDD.n5295 VSS 0.00663f
C7457 VDD.n5296 VSS 0.00332f
C7458 VDD.n5297 VSS 0.00979f
C7459 VDD.n5298 VSS 0.00979f
C7460 VDD.n5299 VSS 0.00269f
C7461 VDD.n5300 VSS 0.00277f
C7462 VDD.n5302 VSS 0.0104f
C7463 VDD.n5304 VSS 0.0129f
C7464 VDD.n5305 VSS 0.00979f
C7465 VDD.n5306 VSS 0.00979f
C7466 VDD.n5307 VSS 0.00332f
C7467 VDD.n5308 VSS 0.00663f
C7468 VDD.n5309 VSS 0.00806f
C7469 VDD.n5310 VSS 0.00585f
C7470 VDD.n5311 VSS 0.00411f
C7471 VDD.n5312 VSS 0.00332f
C7472 VDD.n5313 VSS 0.00439f
C7473 VDD.n5314 VSS 3.26e-19
C7474 VDD.n5315 VSS 0.00488f
C7475 VDD.n5316 VSS 0.00798f
C7476 VDD.n5317 VSS -0.174f
C7477 VDD.n5318 VSS 0.0223f
C7478 VDD.n5319 VSS 0.0136f
C7479 VDD.n5320 VSS 0.00439f
C7480 VDD.n5321 VSS 0.00472f
C7481 VDD.n5322 VSS 0.00585f
C7482 VDD.n5323 VSS 0.00663f
C7483 VDD.n5324 VSS 0.00806f
C7484 VDD.n5325 VSS 0.00348f
C7485 VDD.n5326 VSS 0.00269f
C7486 VDD.n5327 VSS 0.00348f
C7487 VDD.n5328 VSS 3.16e-19
C7488 VDD.n5329 VSS 0.0104f
C7489 VDD.n5331 VSS 0.0129f
C7490 VDD.n5333 VSS 0.00277f
C7491 VDD.n5334 VSS 0.00269f
C7492 VDD.n5335 VSS 3.16e-19
C7493 VDD.n5336 VSS 0.00348f
C7494 VDD.n5337 VSS 4.74e-19
C7495 VDD.n5338 VSS 0.00488f
C7496 VDD.n5339 VSS 0.00798f
C7497 VDD.n5340 VSS 0.0227f
C7498 VDD.n5341 VSS 0.0223f
C7499 VDD.n5342 VSS 0.0141f
C7500 VDD.n5343 VSS 0.0136f
C7501 VDD.n5344 VSS -0.0753f
C7502 VDD.n5345 VSS -0.211f
C7503 VDD.n5346 VSS 0.00585f
C7504 VDD.n5347 VSS 0.00806f
C7505 VDD.n5348 VSS 0.00663f
C7506 VDD.n5349 VSS 0.00332f
C7507 VDD.n5350 VSS 0.00979f
C7508 VDD.n5351 VSS 0.00979f
C7509 VDD.n5352 VSS 0.0129f
C7510 VDD.n5354 VSS 0.00277f
C7511 VDD.n5355 VSS 0.0236f
C7512 VDD.n5356 VSS 3.16e-19
C7513 VDD.n5357 VSS 0.00348f
C7514 VDD.n5358 VSS 4.74e-19
C7515 VDD.n5359 VSS 0.00488f
C7516 VDD.n5360 VSS 0.0286f
C7517 VDD.n5361 VSS 0.00472f
C7518 VDD.n5362 VSS 0.0285f
C7519 VDD.n5363 VSS 0.08f
C7520 VDD.n5364 VSS 0.0136f
C7521 VDD.n5365 VSS 0.0223f
C7522 VDD.n5366 VSS 0.00472f
C7523 VDD.n5367 VSS 0.00781f
C7524 VDD.n5368 VSS 0.00391f
C7525 VDD.n5369 VSS 0.0227f
C7526 VDD.n5370 VSS 0.0141f
C7527 VDD.n5371 VSS -0.0753f
C7528 VDD.n5372 VSS 0.00332f
C7529 VDD.n5373 VSS 0.00411f
C7530 VDD.n5374 VSS 0.00916f
C7531 VDD.n5375 VSS 0.00663f
C7532 VDD.n5376 VSS 0.00806f
C7533 VDD.n5377 VSS 0.00348f
C7534 VDD.n5378 VSS 0.00269f
C7535 VDD.n5379 VSS 0.00269f
C7536 VDD.n5380 VSS 3.16e-19
C7537 VDD.n5381 VSS 0.0104f
C7538 VDD.n5383 VSS 0.00277f
C7539 VDD.n5385 VSS 0.0129f
C7540 VDD.n5386 VSS 0.00979f
C7541 VDD.n5387 VSS 0.00979f
C7542 VDD.n5388 VSS 0.00332f
C7543 VDD.n5389 VSS 0.00348f
C7544 VDD.n5390 VSS 0.00806f
C7545 VDD.n5391 VSS 0.00663f
C7546 VDD.n5392 VSS 0.00916f
C7547 VDD.n5393 VSS 0.00411f
C7548 VDD.n5394 VSS 0.00332f
C7549 VDD.n5395 VSS 0.00439f
C7550 VDD.n5396 VSS 0.0141f
C7551 VDD.n5397 VSS 0.0227f
C7552 VDD.n5398 VSS 0.00391f
C7553 VDD.n5399 VSS 0.00781f
C7554 VDD.n5400 VSS 0.00472f
C7555 VDD.n5401 VSS 3.26e-19
C7556 VDD.n5402 VSS -0.0782f
C7557 VDD.n5403 VSS 0.0141f
C7558 VDD.n5404 VSS 0.0227f
C7559 VDD.n5405 VSS 0.00391f
C7560 VDD.n5406 VSS 0.00488f
C7561 VDD.n5407 VSS 0.00585f
C7562 VDD.n5408 VSS 0.00411f
C7563 VDD.n5409 VSS 0.00916f
C7564 VDD.n5410 VSS 0.00348f
C7565 VDD.n5411 VSS 3.16e-19
C7566 VDD.n5412 VSS 0.00269f
C7567 VDD.n5413 VSS 0.00277f
C7568 VDD.n5415 VSS 0.0129f
C7569 VDD.n5417 VSS 0.0104f
C7570 VDD.n5418 VSS 3.16e-19
C7571 VDD.n5419 VSS 0.00348f
C7572 VDD.n5420 VSS 4.74e-19
C7573 VDD.n5421 VSS 0.00472f
C7574 VDD.n5422 VSS 3.26e-19
C7575 VDD.n5423 VSS 0.0136f
C7576 VDD.n5424 VSS 0.0141f
C7577 VDD.n5425 VSS 0.0223f
C7578 VDD.n5426 VSS 0.0227f
C7579 VDD.n5427 VSS 0.00391f
C7580 VDD.n5428 VSS -0.211f
C7581 VDD.n5429 VSS 0.00585f
C7582 VDD.n5430 VSS 0.00806f
C7583 VDD.n5431 VSS 0.00348f
C7584 VDD.n5432 VSS 0.00269f
C7585 VDD.n5433 VSS 0.00332f
C7586 VDD.n5434 VSS 0.00979f
C7587 VDD.n5435 VSS 0.00979f
C7588 VDD.n5436 VSS 0.0129f
C7589 VDD.n5438 VSS 0.0104f
C7590 VDD.n5440 VSS 0.00277f
C7591 VDD.n5441 VSS 0.00269f
C7592 VDD.n5442 VSS 0.00979f
C7593 VDD.n5443 VSS 0.00979f
C7594 VDD.n5444 VSS 0.00332f
C7595 VDD.n5445 VSS 0.00348f
C7596 VDD.n5446 VSS 0.00806f
C7597 VDD.n5447 VSS 0.00663f
C7598 VDD.n5448 VSS 0.00916f
C7599 VDD.n5449 VSS 0.00411f
C7600 VDD.n5450 VSS 0.00332f
C7601 VDD.n5451 VSS 0.00439f
C7602 VDD.n5452 VSS 0.0141f
C7603 VDD.n5453 VSS 0.0227f
C7604 VDD.n5454 VSS 0.00391f
C7605 VDD.n5455 VSS 0.00781f
C7606 VDD.n5456 VSS 0.00472f
C7607 VDD.n5457 VSS 3.26e-19
C7608 VDD.n5458 VSS -0.0782f
C7609 VDD.n5459 VSS 0.0141f
C7610 VDD.n5460 VSS 0.00472f
C7611 VDD.n5461 VSS 0.00439f
C7612 VDD.n5462 VSS 0.0136f
C7613 VDD.n5463 VSS 0.0141f
C7614 VDD.n5464 VSS 0.06f
C7615 VDD.n5465 VSS 0.0243f
C7616 VDD.n5466 VSS 0.00488f
C7617 VDD.n5467 VSS 0.0251f
C7618 VDD.n5468 VSS 0.00411f
C7619 VDD.n5469 VSS 0.0295f
C7620 VDD.n5470 VSS 0.00348f
C7621 VDD.n5471 VSS 3.16e-19
C7622 VDD.n5472 VSS 0.0104f
C7623 VDD.n5474 VSS 0.00277f
C7624 VDD.n5475 VSS 0.0186f
C7625 VDD.n5476 VSS 0.03f
C7626 VDD.n5477 VSS 0.0312f
C7627 VDD.n5478 VSS 0.0173f
C7628 VDD.n5479 VSS 0.00277f
C7629 VDD.n5480 VSS 0.00269f
C7630 VDD.n5481 VSS 3.16e-19
C7631 VDD.n5482 VSS 0.00348f
C7632 VDD.n5483 VSS 4.74e-19
C7633 VDD.n5484 VSS 0.00488f
C7634 VDD.n5485 VSS 0.00798f
C7635 VDD.n5486 VSS -0.174f
C7636 VDD.n5487 VSS 0.0223f
C7637 VDD.n5488 VSS 0.0136f
C7638 VDD.n5489 VSS 0.00439f
C7639 VDD.n5490 VSS 0.00472f
C7640 VDD.n5491 VSS 0.00585f
C7641 VDD.n5492 VSS 0.00806f
C7642 VDD.n5493 VSS 0.00663f
C7643 VDD.n5494 VSS 0.00332f
C7644 VDD.n5495 VSS 0.00979f
C7645 VDD.n5496 VSS 0.00979f
C7646 VDD.n5497 VSS 0.0129f
C7647 VDD.n5499 VSS 0.00277f
C7648 VDD.n5501 VSS 0.0104f
C7649 VDD.n5502 VSS 3.16e-19
C7650 VDD.n5503 VSS 0.00348f
C7651 VDD.n5504 VSS 4.74e-19
C7652 VDD.n5505 VSS 0.00488f
C7653 VDD.n5506 VSS 0.00798f
C7654 VDD.n5507 VSS 0.0227f
C7655 VDD.n5508 VSS 0.0223f
C7656 VDD.n5509 VSS 0.0136f
C7657 VDD.n5510 VSS 0.00374f
C7658 VDD.n5511 VSS 0.0141f
C7659 VDD.n5512 VSS 0.0223f
C7660 VDD.n5513 VSS 0.0227f
C7661 VDD.n5514 VSS 0.00798f
C7662 VDD.n5515 VSS 0.00488f
C7663 VDD.n5516 VSS 0.00348f
C7664 VDD.n5517 VSS 4.74e-19
C7665 VDD.n5518 VSS 0.00332f
C7666 VDD.n5519 VSS -0.0753f
C7667 VDD.n5520 VSS -0.211f
C7668 VDD.n5521 VSS 0.00585f
C7669 VDD.n5522 VSS 0.00806f
C7670 VDD.n5523 VSS 0.00663f
C7671 VDD.n5524 VSS 0.00332f
C7672 VDD.n5525 VSS 0.00979f
C7673 VDD.n5526 VSS 0.00979f
C7674 VDD.n5527 VSS 0.00269f
C7675 VDD.n5528 VSS 0.00277f
C7676 VDD.n5530 VSS 0.0104f
C7677 VDD.n5532 VSS 0.0129f
C7678 VDD.n5533 VSS 0.00979f
C7679 VDD.n5534 VSS 0.00979f
C7680 VDD.n5535 VSS 0.00332f
C7681 VDD.n5536 VSS 0.00663f
C7682 VDD.n5537 VSS 0.00806f
C7683 VDD.n5538 VSS 0.00585f
C7684 VDD.n5539 VSS 0.00411f
C7685 VDD.n5540 VSS 0.00332f
C7686 VDD.n5541 VSS 0.00439f
C7687 VDD.n5542 VSS 3.26e-19
C7688 VDD.n5543 VSS 0.00488f
C7689 VDD.n5544 VSS 0.00798f
C7690 VDD.n5545 VSS -0.174f
C7691 VDD.n5546 VSS 0.0223f
C7692 VDD.n5547 VSS 0.0136f
C7693 VDD.n5548 VSS 0.00439f
C7694 VDD.n5549 VSS 0.00472f
C7695 VDD.n5550 VSS 0.00585f
C7696 VDD.n5551 VSS 0.00663f
C7697 VDD.n5552 VSS 0.00806f
C7698 VDD.n5553 VSS 0.00348f
C7699 VDD.n5554 VSS 0.00269f
C7700 VDD.n5555 VSS 0.00348f
C7701 VDD.n5556 VSS 3.16e-19
C7702 VDD.n5557 VSS 0.0104f
C7703 VDD.n5559 VSS 0.0129f
C7704 VDD.n5561 VSS 0.00277f
C7705 VDD.n5562 VSS 0.00269f
C7706 VDD.n5563 VSS 3.16e-19
C7707 VDD.n5564 VSS 0.00348f
C7708 VDD.n5565 VSS 4.74e-19
C7709 VDD.n5566 VSS 0.00488f
C7710 VDD.n5567 VSS 0.00798f
C7711 VDD.n5568 VSS 0.0227f
C7712 VDD.n5569 VSS 0.0223f
C7713 VDD.n5570 VSS 0.0141f
C7714 VDD.n5571 VSS 0.0136f
C7715 VDD.n5572 VSS -0.0753f
C7716 VDD.n5573 VSS -0.211f
C7717 VDD.n5574 VSS 0.00585f
C7718 VDD.n5575 VSS 0.00806f
C7719 VDD.n5576 VSS 0.00663f
C7720 VDD.n5577 VSS 0.00332f
C7721 VDD.n5578 VSS 0.00979f
C7722 VDD.n5579 VSS 0.00979f
C7723 VDD.n5580 VSS 0.0129f
C7724 VDD.n5582 VSS 0.00277f
C7725 VDD.n5583 VSS 0.0236f
C7726 VDD.n5584 VSS 3.16e-19
C7727 VDD.n5585 VSS 0.00348f
C7728 VDD.n5586 VSS 4.74e-19
C7729 VDD.n5587 VSS 0.00488f
C7730 VDD.n5588 VSS 0.0286f
C7731 VDD.n5589 VSS 0.00472f
C7732 VDD.n5590 VSS 0.0285f
C7733 VDD.n5591 VSS 0.08f
C7734 VDD.n5592 VSS 0.0136f
C7735 VDD.n5593 VSS 0.0223f
C7736 VDD.n5594 VSS 0.00472f
C7737 VDD.n5595 VSS 0.00781f
C7738 VDD.n5596 VSS 0.00391f
C7739 VDD.n5597 VSS 0.0227f
C7740 VDD.n5598 VSS 0.0141f
C7741 VDD.n5599 VSS -0.0753f
C7742 VDD.n5600 VSS 0.00332f
C7743 VDD.n5601 VSS 0.00411f
C7744 VDD.n5602 VSS 0.00916f
C7745 VDD.n5603 VSS 0.00663f
C7746 VDD.n5604 VSS 0.00806f
C7747 VDD.n5605 VSS 0.00348f
C7748 VDD.n5606 VSS 0.00269f
C7749 VDD.n5607 VSS 0.00269f
C7750 VDD.n5608 VSS 3.16e-19
C7751 VDD.n5609 VSS 0.0104f
C7752 VDD.n5611 VSS 0.00277f
C7753 VDD.n5613 VSS 0.0129f
C7754 VDD.n5614 VSS 0.00979f
C7755 VDD.n5615 VSS 0.00979f
C7756 VDD.n5616 VSS 0.00332f
C7757 VDD.n5617 VSS 0.00348f
C7758 VDD.n5618 VSS 0.00806f
C7759 VDD.n5619 VSS 0.00663f
C7760 VDD.n5620 VSS 0.00916f
C7761 VDD.n5621 VSS 0.00411f
C7762 VDD.n5622 VSS 0.00332f
C7763 VDD.n5623 VSS 0.00439f
C7764 VDD.n5624 VSS 0.0141f
C7765 VDD.n5625 VSS 0.0227f
C7766 VDD.n5626 VSS 0.00391f
C7767 VDD.n5627 VSS 0.00781f
C7768 VDD.n5628 VSS 0.00472f
C7769 VDD.n5629 VSS 3.26e-19
C7770 VDD.n5630 VSS -0.0782f
C7771 VDD.n5631 VSS 0.0141f
C7772 VDD.n5632 VSS 0.0227f
C7773 VDD.n5633 VSS 0.00391f
C7774 VDD.n5634 VSS 0.00488f
C7775 VDD.n5635 VSS 0.00585f
C7776 VDD.n5636 VSS 0.00411f
C7777 VDD.n5637 VSS 0.00916f
C7778 VDD.n5638 VSS 0.00348f
C7779 VDD.n5639 VSS 3.16e-19
C7780 VDD.n5640 VSS 0.00269f
C7781 VDD.n5641 VSS 0.00277f
C7782 VDD.n5643 VSS 0.0129f
C7783 VDD.n5645 VSS 0.0104f
C7784 VDD.n5646 VSS 3.16e-19
C7785 VDD.n5647 VSS 0.00348f
C7786 VDD.n5648 VSS 4.74e-19
C7787 VDD.n5649 VSS 0.00472f
C7788 VDD.n5650 VSS 3.26e-19
C7789 VDD.n5651 VSS 0.0136f
C7790 VDD.n5652 VSS 0.0141f
C7791 VDD.n5653 VSS 0.0223f
C7792 VDD.n5654 VSS 0.0227f
C7793 VDD.n5655 VSS 0.00391f
C7794 VDD.n5656 VSS -0.211f
C7795 VDD.n5657 VSS 0.00585f
C7796 VDD.n5658 VSS 0.00806f
C7797 VDD.n5659 VSS 0.00348f
C7798 VDD.n5660 VSS 0.00269f
C7799 VDD.n5661 VSS 0.00332f
C7800 VDD.n5662 VSS 0.00979f
C7801 VDD.n5663 VSS 0.00979f
C7802 VDD.n5664 VSS 0.0129f
C7803 VDD.n5666 VSS 0.0104f
C7804 VDD.n5668 VSS 0.00277f
C7805 VDD.n5669 VSS 0.00269f
C7806 VDD.n5670 VSS 0.00979f
C7807 VDD.n5671 VSS 0.00979f
C7808 VDD.n5672 VSS 0.00332f
C7809 VDD.n5673 VSS 0.00348f
C7810 VDD.n5674 VSS 0.00806f
C7811 VDD.n5675 VSS 0.00663f
C7812 VDD.n5676 VSS 0.00916f
C7813 VDD.n5677 VSS 0.00411f
C7814 VDD.n5678 VSS 0.00332f
C7815 VDD.n5679 VSS 0.00439f
C7816 VDD.n5680 VSS 0.0141f
C7817 VDD.n5681 VSS 0.0227f
C7818 VDD.n5682 VSS 0.00391f
C7819 VDD.n5683 VSS 0.00781f
C7820 VDD.n5684 VSS 0.00472f
C7821 VDD.n5685 VSS 3.26e-19
C7822 VDD.n5686 VSS -0.0782f
C7823 VDD.n5687 VSS 0.0141f
C7824 VDD.n5688 VSS 0.00472f
C7825 VDD.n5689 VSS 0.00439f
C7826 VDD.n5690 VSS 0.0136f
C7827 VDD.n5691 VSS 0.0141f
C7828 VDD.n5692 VSS 0.06f
C7829 VDD.n5693 VSS 0.0243f
C7830 VDD.n5694 VSS 0.00488f
C7831 VDD.n5695 VSS 0.0251f
C7832 VDD.n5696 VSS 0.00411f
C7833 VDD.n5697 VSS 0.0295f
C7834 VDD.n5698 VSS 0.00348f
C7835 VDD.n5699 VSS 3.16e-19
C7836 VDD.n5700 VSS 0.0104f
C7837 VDD.n5702 VSS 0.00277f
C7838 VDD.n5703 VSS 0.0186f
C7839 VDD.n5704 VSS 0.03f
C7840 VDD.n5705 VSS 0.0312f
C7841 VDD.n5706 VSS 0.0173f
C7842 VDD.n5707 VSS 0.00277f
C7843 VDD.n5708 VSS 0.00269f
C7844 VDD.n5709 VSS 3.16e-19
C7845 VDD.n5710 VSS 0.00348f
C7846 VDD.n5711 VSS 4.74e-19
C7847 VDD.n5712 VSS 0.00488f
C7848 VDD.n5713 VSS 0.00798f
C7849 VDD.n5714 VSS -0.174f
C7850 VDD.n5715 VSS 0.0223f
C7851 VDD.n5716 VSS 0.0136f
C7852 VDD.n5717 VSS 0.00439f
C7853 VDD.n5718 VSS 0.00472f
C7854 VDD.n5719 VSS 0.00585f
C7855 VDD.n5720 VSS 0.00806f
C7856 VDD.n5721 VSS 0.00663f
C7857 VDD.n5722 VSS 0.00332f
C7858 VDD.n5723 VSS 0.00979f
C7859 VDD.n5724 VSS 0.00979f
C7860 VDD.n5725 VSS 0.0129f
C7861 VDD.n5727 VSS 0.00277f
C7862 VDD.n5729 VSS 0.0104f
C7863 VDD.n5730 VSS 3.16e-19
C7864 VDD.n5731 VSS 0.00348f
C7865 VDD.n5732 VSS 4.74e-19
C7866 VDD.n5733 VSS 0.00488f
C7867 VDD.n5734 VSS 0.00798f
C7868 VDD.n5735 VSS 0.0227f
C7869 VDD.n5736 VSS 0.0223f
C7870 VDD.n5737 VSS 0.0136f
C7871 VDD.n5738 VSS 0.00374f
C7872 VDD.n5739 VSS 0.0141f
C7873 VDD.n5740 VSS 0.0223f
C7874 VDD.n5741 VSS 0.0227f
C7875 VDD.n5742 VSS 0.00798f
C7876 VDD.n5743 VSS 0.00488f
C7877 VDD.n5744 VSS 0.00348f
C7878 VDD.n5745 VSS 4.74e-19
C7879 VDD.n5746 VSS 0.00332f
C7880 VDD.n5747 VSS -0.0753f
C7881 VDD.n5748 VSS -0.211f
C7882 VDD.n5749 VSS 0.00585f
C7883 VDD.n5750 VSS 0.00806f
C7884 VDD.n5751 VSS 0.00663f
C7885 VDD.n5752 VSS 0.00332f
C7886 VDD.n5753 VSS 0.00979f
C7887 VDD.n5754 VSS 0.00979f
C7888 VDD.n5755 VSS 0.00269f
C7889 VDD.n5756 VSS 0.00277f
C7890 VDD.n5758 VSS 0.0104f
C7891 VDD.n5760 VSS 0.0129f
C7892 VDD.n5761 VSS 0.00979f
C7893 VDD.n5762 VSS 0.00979f
C7894 VDD.n5763 VSS 0.00332f
C7895 VDD.n5764 VSS 0.00663f
C7896 VDD.n5765 VSS 0.00806f
C7897 VDD.n5766 VSS 0.00585f
C7898 VDD.n5767 VSS 0.00411f
C7899 VDD.n5768 VSS 0.00332f
C7900 VDD.n5769 VSS 0.00439f
C7901 VDD.n5770 VSS 3.26e-19
C7902 VDD.n5771 VSS 0.00488f
C7903 VDD.n5772 VSS 0.00798f
C7904 VDD.n5773 VSS -0.174f
C7905 VDD.n5774 VSS 0.0223f
C7906 VDD.n5775 VSS 0.0136f
C7907 VDD.n5776 VSS 0.00439f
C7908 VDD.n5777 VSS 0.00472f
C7909 VDD.n5778 VSS 0.00585f
C7910 VDD.n5779 VSS 0.00663f
C7911 VDD.n5780 VSS 0.00806f
C7912 VDD.n5781 VSS 0.00348f
C7913 VDD.n5782 VSS 0.00269f
C7914 VDD.n5783 VSS 0.00348f
C7915 VDD.n5784 VSS 3.16e-19
C7916 VDD.n5785 VSS 0.0104f
C7917 VDD.n5787 VSS 0.0129f
C7918 VDD.n5789 VSS 0.00277f
C7919 VDD.n5790 VSS 0.00269f
C7920 VDD.n5791 VSS 3.16e-19
C7921 VDD.n5792 VSS 0.00348f
C7922 VDD.n5793 VSS 4.74e-19
C7923 VDD.n5794 VSS 0.00488f
C7924 VDD.n5795 VSS 0.00798f
C7925 VDD.n5796 VSS 0.0227f
C7926 VDD.n5797 VSS 0.0223f
C7927 VDD.n5798 VSS 0.0136f
C7928 VDD.n5799 VSS -0.0753f
C7929 VDD.n5800 VSS -0.211f
C7930 VDD.n5801 VSS 0.00585f
C7931 VDD.n5802 VSS 0.00806f
C7932 VDD.n5803 VSS 0.00663f
C7933 VDD.n5804 VSS 0.00332f
C7934 VDD.n5805 VSS 0.00979f
C7935 VDD.n5806 VSS 0.00979f
C7936 VDD.n5807 VSS 0.0129f
C7937 VDD.n5809 VSS 0.00277f
C7938 VDD.n5810 VSS 0.0236f
C7939 VDD.n5811 VSS 3.16e-19
C7940 VDD.n5812 VSS 0.00348f
C7941 VDD.n5813 VSS 4.74e-19
C7942 VDD.n5814 VSS 0.00488f
C7943 VDD.n5815 VSS 0.0286f
C7944 VDD.n5816 VSS 0.0805f
C7945 VDD.n5817 VSS 0.08f
C7946 VDD.n5818 VSS 0.0136f
C7947 VDD.n5819 VSS 3.26e-19
C7948 VDD.n5820 VSS 0.00472f
C7949 VDD.n5821 VSS 0.00332f
C7950 VDD.n5822 VSS 4.74e-19
C7951 VDD.n5823 VSS 0.00348f
C7952 VDD.n5824 VSS 3.16e-19
C7953 VDD.n5825 VSS 0.0236f
C7954 VDD.n5827 VSS 0.00277f
C7955 VDD.n5828 VSS 0.00269f
C7956 VDD.n5829 VSS 0.00979f
C7957 VDD.n5830 VSS 0.00979f
C7958 VDD.n5831 VSS 0.00332f
C7959 VDD.n5832 VSS 0.00663f
C7960 VDD.n5833 VSS 0.00806f
C7961 VDD.n5834 VSS 0.00585f
C7962 VDD.n5835 VSS -0.211f
C7963 VDD.n5836 VSS 0.00391f
C7964 VDD.n5837 VSS 0.0227f
C7965 VDD.n5838 VSS 0.0223f
C7966 VDD.n5839 VSS 0.0141f
C7967 VDD.n5840 VSS 0.0136f
C7968 VDD.n5841 VSS 3.26e-19
C7969 VDD.n5842 VSS 0.00472f
C7970 VDD.n5843 VSS 0.00332f
C7971 VDD.n5844 VSS 4.74e-19
C7972 VDD.n5845 VSS 0.00348f
C7973 VDD.n5846 VSS 3.16e-19
C7974 VDD.n5847 VSS 0.0104f
C7975 VDD.n5849 VSS 0.00277f
C7976 VDD.n5850 VSS 0.0129f
C7977 VDD.n5852 VSS 0.0104f
C7978 VDD.n5853 VSS 3.16e-19
C7979 VDD.n5854 VSS 0.00269f
C7980 VDD.n5855 VSS 0.00979f
C7981 VDD.n5856 VSS 0.00332f
C7982 VDD.n5857 VSS 0.00663f
C7983 VDD.n5858 VSS 0.00806f
C7984 VDD.n5859 VSS 0.00585f
C7985 VDD.n5860 VSS 0.00488f
C7986 VDD.n5861 VSS 0.00391f
C7987 VDD.n5862 VSS 0.00472f
C7988 VDD.n5863 VSS 0.00781f
C7989 VDD.n5864 VSS -0.182f
C7990 VDD.n5865 VSS -0.0782f
C7991 VDD.n5866 VSS 0.0223f
C7992 VDD.n5867 VSS 0.00472f
C7993 VDD.n5868 VSS 0.00781f
C7994 VDD.n5869 VSS 0.00391f
C7995 VDD.n5870 VSS 0.0227f
C7996 VDD.n5871 VSS 0.0141f
C7997 VDD.n5872 VSS 0.00439f
C7998 VDD.n5873 VSS 0.00332f
C7999 VDD.n5874 VSS 0.00411f
C8000 VDD.n5875 VSS 0.00916f
C8001 VDD.n5876 VSS 0.00663f
C8002 VDD.n5877 VSS 0.00806f
C8003 VDD.n5878 VSS 0.00348f
C8004 VDD.n5879 VSS 0.00269f
C8005 VDD.n5880 VSS 0.00269f
C8006 VDD.n5881 VSS 3.16e-19
C8007 VDD.n5882 VSS 0.0104f
C8008 VDD.n5884 VSS 0.00277f
C8009 VDD.n5886 VSS 0.0129f
C8010 VDD.n5887 VSS 0.00979f
C8011 VDD.n5888 VSS 0.00979f
C8012 VDD.n5889 VSS 0.00332f
C8013 VDD.n5890 VSS 0.00348f
C8014 VDD.n5891 VSS 0.00806f
C8015 VDD.n5892 VSS 0.00663f
C8016 VDD.n5893 VSS 0.00916f
C8017 VDD.n5894 VSS 0.00411f
C8018 VDD.n5895 VSS 0.00332f
C8019 VDD.n5896 VSS -0.0753f
C8020 VDD.n5897 VSS 0.0141f
C8021 VDD.n5898 VSS 0.0227f
C8022 VDD.n5899 VSS 0.00391f
C8023 VDD.n5900 VSS 0.00781f
C8024 VDD.n5901 VSS 0.00472f
C8025 VDD.n5902 VSS 3.26e-19
C8026 VDD.n5903 VSS 0.0136f
C8027 VDD.n5904 VSS 0.0141f
C8028 VDD.n5905 VSS 0.00472f
C8029 VDD.n5906 VSS 3.26e-19
C8030 VDD.n5907 VSS -0.0782f
C8031 VDD.n5908 VSS -0.182f
C8032 VDD.n5909 VSS 0.0227f
C8033 VDD.n5910 VSS 0.00391f
C8034 VDD.n5911 VSS 0.00488f
C8035 VDD.n5912 VSS 0.00585f
C8036 VDD.n5913 VSS 0.00411f
C8037 VDD.n5914 VSS 0.00916f
C8038 VDD.n5915 VSS 0.00348f
C8039 VDD.n5916 VSS 3.16e-19
C8040 VDD.n5917 VSS 0.00269f
C8041 VDD.n5918 VSS 0.00277f
C8042 VDD.n5920 VSS 0.0129f
C8043 VDD.n5921 VSS 0.0276f
C8044 VDD.n5922 VSS 0.0442f
C8045 VDD.n5923 VSS 0.0422f
C8046 VDD.n5924 VSS 0.0389f
C8047 VDD.n5925 VSS 0.0398f
C8048 VDD.n5926 VSS 0.0601f
C8049 VDD.n5927 VSS 3.67f
C8050 VDD.n5928 VSS 3.73f
C8051 VDD.n5929 VSS 0.063f
C8052 VDD.n5930 VSS 0.0439f
C8053 VDD.n5931 VSS 0.0433f
C8054 VDD.n5932 VSS 0.00585f
C8055 VDD.n5933 VSS 0.00332f
C8056 VDD.n5934 VSS 0.00348f
C8057 VDD.n5935 VSS 0.00806f
C8058 VDD.n5936 VSS 0.00663f
C8059 VDD.n5937 VSS 0.00956f
C8060 VDD.n5938 VSS 0.00411f
C8061 VDD.n5939 VSS 0.00332f
C8062 VDD.n5940 VSS -0.0753f
C8063 VDD.n5941 VSS 0.0143f
C8064 VDD.n5942 VSS 0.0231f
C8065 VDD.n5943 VSS 0.00391f
C8066 VDD.n5944 VSS 0.00781f
C8067 VDD.n5945 VSS 0.00472f
C8068 VDD.n5946 VSS 3.26e-19
C8069 VDD.n5947 VSS 0.0139f
C8070 VDD.n5948 VSS 0.0143f
C8071 VDD.n5949 VSS 0.0143f
C8072 VDD.n5950 VSS 0.00472f
C8073 VDD.n5951 VSS 0.00488f
C8074 VDD.n5952 VSS 4.74e-19
C8075 VDD.n5953 VSS 0.00585f
C8076 VDD.n5954 VSS 0.00348f
C8077 VDD.n5955 VSS 0.00332f
C8078 VDD.n5956 VSS 4.74e-19
C8079 VDD.n5957 VSS 0.00348f
C8080 VDD.n5958 VSS 0.00979f
C8081 VDD.n5959 VSS 0.00979f
C8082 VDD.n5960 VSS 0.00332f
C8083 VDD.n5961 VSS 0.00348f
C8084 VDD.n5962 VSS 0.00269f
C8085 VDD.n5963 VSS 0.00269f
C8086 VDD.n5964 VSS 0.0104f
C8087 VDD.n5965 VSS 3.16e-19
C8088 VDD.n5966 VSS 0.00277f
C8089 VDD.n5967 VSS 0.00269f
C8090 VDD.n5968 VSS 0.00979f
C8091 VDD.n5969 VSS 0.00979f
C8092 VDD.n5970 VSS 0.00269f
C8093 VDD.n5971 VSS 0.00663f
C8094 VDD.n5972 VSS 0.00348f
C8095 VDD.n5973 VSS 0.00806f
C8096 VDD.n5974 VSS 0.00332f
C8097 VDD.n5975 VSS 0.00781f
C8098 VDD.n5976 VSS 0.00439f
C8099 VDD.n5977 VSS 0.0143f
C8100 VDD.n5978 VSS 0.00472f
C8101 VDD.n5979 VSS 0.0231f
C8102 VDD.n5980 VSS 0.00391f
C8103 VDD.n5981 VSS 0.00781f
C8104 VDD.n5982 VSS 0.0226f
C8105 VDD.n5983 VSS 0.0139f
C8106 VDD.n5984 VSS 3.26e-19
C8107 VDD.n5985 VSS -0.0753f
C8108 VDD.n5986 VSS 0.00332f
C8109 VDD.n5987 VSS 0.00916f
C8110 VDD.n5988 VSS 0.00411f
C8111 VDD.n5989 VSS 0.00585f
C8112 VDD.n5990 VSS -0.211f
C8113 VDD.n5991 VSS 0.00391f
C8114 VDD.n5992 VSS 0.0231f
C8115 VDD.n5993 VSS 0.0226f
C8116 VDD.n5994 VSS -0.181f
C8117 VDD.n5995 VSS 0.00488f
C8118 VDD.n5996 VSS 3.26e-19
C8119 VDD.n5997 VSS 0.00348f
C8120 VDD.n5998 VSS 0.00411f
C8121 VDD.n5999 VSS 0.00779f
C8122 VDD.n6000 VSS 0.00488f
C8123 VDD.n6001 VSS -0.078f
C8124 VDD.n6002 VSS 0.0305f
C8125 VDD.n6003 VSS 0.00618f
C8126 VDD.n6004 VSS 0.00816f
C8127 VDD.n6005 VSS 0.00767f
C8128 VDD.n6006 VSS 0.0305f
C8129 VDD.n6007 VSS 0.0143f
C8130 VDD.n6008 VSS 0.00439f
C8131 VDD.n6009 VSS 0.00332f
C8132 VDD.n6010 VSS 0.00269f
C8133 VDD.n6011 VSS 0.0104f
C8134 VDD.n6012 VSS 3.16e-19
C8135 VDD.n6013 VSS 0.00269f
C8136 VDD.n6014 VSS 0.00277f
C8137 VDD.n6015 VSS 0.0129f
C8138 VDD.n6016 VSS 0.00979f
C8139 VDD.n6017 VSS 0.00916f
C8140 VDD.n6018 VSS 0.00411f
C8141 VDD.n6019 VSS 0.00585f
C8142 VDD.n6020 VSS 0.00806f
C8143 VDD.n6021 VSS 0.00663f
C8144 VDD.n6022 VSS 0.00332f
C8145 VDD.n6023 VSS 0.00979f
C8146 VDD.n6024 VSS 0.00269f
C8147 VDD.n6025 VSS 0.0104f
C8148 VDD.n6026 VSS 3.16e-19
C8149 VDD.n6027 VSS 0.00348f
C8150 VDD.n6028 VSS 4.74e-19
C8151 VDD.n6029 VSS 0.00472f
C8152 VDD.n6030 VSS 0.00781f
C8153 VDD.n6031 VSS 0.00391f
C8154 VDD.n6032 VSS 0.0231f
C8155 VDD.n6033 VSS 0.0143f
C8156 VDD.n6034 VSS 0.0139f
C8157 VDD.n6035 VSS 3.26e-19
C8158 VDD.n6036 VSS 0.00472f
C8159 VDD.n6037 VSS 4.74e-19
C8160 VDD.n6038 VSS 0.00348f
C8161 VDD.n6039 VSS 0.00269f
C8162 VDD.n6040 VSS 0.00332f
C8163 VDD.n6041 VSS 0.00979f
C8164 VDD.n6042 VSS 0.00979f
C8165 VDD.n6043 VSS 0.00277f
C8166 VDD.n6044 VSS 0.00269f
C8167 VDD.n6045 VSS 0.0104f
C8168 VDD.n6046 VSS 3.16e-19
C8169 VDD.n6047 VSS 0.00269f
C8170 VDD.n6048 VSS 0.00269f
C8171 VDD.n6049 VSS 0.00348f
C8172 VDD.n6050 VSS 0.00806f
C8173 VDD.n6051 VSS 0.00663f
C8174 VDD.n6052 VSS 0.00916f
C8175 VDD.n6053 VSS 0.00411f
C8176 VDD.n6054 VSS 0.00332f
C8177 VDD.n6055 VSS 0.00439f
C8178 VDD.n6056 VSS 3.26e-19
C8179 VDD.n6057 VSS -0.078f
C8180 VDD.n6058 VSS -0.181f
C8181 VDD.n6059 VSS 0.0231f
C8182 VDD.n6060 VSS 0.00391f
C8183 VDD.n6061 VSS 0.00488f
C8184 VDD.n6062 VSS 0.00585f
C8185 VDD.n6063 VSS 0.00411f
C8186 VDD.n6064 VSS 0.00916f
C8187 VDD.n6065 VSS 0.00348f
C8188 VDD.n6066 VSS 3.16e-19
C8189 VDD.n6067 VSS 0.0104f
C8190 VDD.n6068 VSS 0.0129f
C8191 VDD.n6069 VSS 0.00979f
C8192 VDD.n6070 VSS 0.00269f
C8193 VDD.n6071 VSS 0.0314f
C8194 VDD.n6072 VSS 0.0236f
C8195 VDD.n6073 VSS 0.46f
C8196 VDD.n6074 VSS 0.0173f
C8197 VDD.n6075 VSS 0.0102f
C8198 VDD.n6076 VSS 0.0633f
C8199 VDD.t12 VSS 0.00583f
C8200 VDD.n6077 VSS 0.0579f
C8201 VDD.n6078 VSS 0.0361f
C8202 VDD.n6079 VSS 0.0174f
C8203 VDD.n6080 VSS 0.00106f
C8204 VDD.n6081 VSS 0.0166f
C8205 VDD.n6082 VSS 3.48f
C8206 VDD.n6083 VSS 3.5f
C8207 VDD.n6084 VSS 0.256f
C8208 VDD.n6085 VSS 0.0124f
C8209 VDD.n6086 VSS 8.15e-19
C8210 VDD.n6087 VSS 0.0198f
C8211 VDD.n6088 VSS 0.0172f
C8212 VDD.n6089 VSS 0.00391f
C8213 VDD.n6090 VSS 0.00407f
C8214 VDD.n6091 VSS 0.0184f
C8215 VDD.n6092 VSS 0.0273f
C8216 VDD.n6093 VSS 0.0106f
C8217 VDD.n6094 VSS 0.00797f
C8218 VDD.n6095 VSS 0.0314f
C8219 VDD.n6096 VSS 0.172f
C8220 VDD.t46 VSS 0.191f
C8221 VDD.n6097 VSS 0.142f
C8222 VDD.n6098 VSS 0.00824f
C8223 VDD.n6099 VSS 0.0813f
C8224 VDD.n6100 VSS 0.00818f
C8225 VDD.n6101 VSS 0.02f
C8226 VDD.n6102 VSS 0.0109f
C8227 VDD.n6103 VSS 0.0523f
C8228 VDD.n6104 VSS 0.0523f
C8229 VDD.n6105 VSS 0.02f
C8230 VDD.n6106 VSS 0.00824f
C8231 VDD.n6107 VSS 0.0813f
C8232 VDD.n6108 VSS 0.00818f
C8233 VDD.n6109 VSS 0.02f
C8234 VDD.n6110 VSS 0.0523f
C8235 VDD.n6111 VSS 0.0402f
C8236 VDD.n6112 VSS 0.0111f
C8237 VDD.n6113 VSS 0.0232f
C8238 VDD.n6114 VSS 0.0186f
C8239 VDD.n6115 VSS 0.017f
C8240 VDD.n6116 VSS 0.0069f
C8241 VDD.n6117 VSS 0.0124f
C8242 VDD.n6118 VSS 0.00461f
C8243 VDD.n6119 VSS 0.00483f
C8244 VDD.n6120 VSS 0.00184f
C8245 VDD.n6121 VSS 0.00135f
C8246 VDD.n6122 VSS 0.0108f
C8247 VDD.n6123 VSS 0.00256f
C8248 VDD.n6124 VSS 0.00163f
C8249 VDD.n6125 VSS 0.0405f
C8250 VDD.n6126 VSS 0.205f
C8251 VDD.t50 VSS 0.279f
C8252 VDD.n6127 VSS 0.253f
C8253 VDD.n6128 VSS 0.0202f
C8254 VDD.n6129 VSS 0.00797f
C8255 VDD.n6130 VSS 0.0556f
C8256 VDD.n6131 VSS 0.0225f
C8257 VDD.n6132 VSS 0.0211f
C8258 VDD.n6133 VSS 0.0197f
C8259 VDD.n6134 VSS 0.016f
C8260 VDD.n6135 VSS 0.0124f
C8261 VDD.n6136 VSS 0.31f
C8262 VDD.n6137 VSS 2.06f
C8263 VDD.n6138 VSS 0.444f
C8264 VDD.n6139 VSS 0.298f
C8265 VDD.n6140 VSS 0.02f
C8266 VDD.n6141 VSS 0.00824f
C8267 VDD.n6142 VSS 0.02f
C8268 VDD.n6143 VSS 0.00634f
C8269 VDD.n6144 VSS 0.00818f
C8270 VDD.n6145 VSS 0.0813f
C8271 VDD.n6146 VSS 1.26f
C8272 VDD.n6147 VSS 1.7f
C8273 VDD.t57 VSS 1.75f
C8274 VDD.n6148 VSS 0.00824f
C8275 VDD.n6149 VSS 0.02f
C8276 VDD.n6150 VSS 0.02f
C8277 VDD.n6151 VSS 0.0109f
C8278 VDD.n6152 VSS 0.00634f
C8279 VDD.n6153 VSS 0.00818f
C8280 VDD.n6154 VSS 0.0813f
C8281 VDD.t0 VSS 0.428f
C8282 VDD.t7 VSS 0.896f
C8283 VDD.n6155 VSS 0.0156f
C8284 VDD.t10 VSS 2.21f
C8285 VDD.t18 VSS 6.67f
C8286 VDD.t77 VSS 5.11f
C8287 VDD.n6156 VSS 0.00797f
C8288 VDD.n6157 VSS 0.0314f
C8289 VDD.n6158 VSS 0.0632f
C8290 VDD.n6159 VSS 0.915f
C8291 VDD.n6160 VSS 1.59f
C8292 VDD.t40 VSS 2.33f
C8293 VDD.n6161 VSS 2.08f
C8294 VDD.n6162 VSS 0.00824f
C8295 VDD.n6163 VSS 0.0813f
C8296 VDD.n6164 VSS 0.00818f
C8297 VDD.n6165 VSS 0.02f
C8298 VDD.n6166 VSS 0.0109f
C8299 VDD.n6167 VSS 0.067f
C8300 VDD.n6168 VSS 0.0777f
C8301 VDD.n6169 VSS 0.02f
C8302 VDD.n6170 VSS 0.00824f
C8303 VDD.n6171 VSS 0.0813f
C8304 VDD.n6172 VSS 0.00818f
C8305 VDD.n6173 VSS 0.02f
C8306 VDD.n6174 VSS 0.059f
C8307 VDD.n6175 VSS 0.126f
C8308 VDD.n6176 VSS 0.0199f
C8309 VDD.t19 VSS 0.00943f
C8310 VDD.n6177 VSS 0.136f
C8311 VDD.n6178 VSS 0.02f
C8312 VDD.n6179 VSS 0.174f
C8313 VDD.n6180 VSS 17.1f
C8314 VDD.n6181 VSS 0.0141f
C8315 VDD.n6182 VSS 0.0398f
C8316 VDD.n6183 VSS 0.00439f
C8317 VDD.n6184 VSS 0.0136f
C8318 VDD.n6185 VSS -0.0845f
C8319 VDD.n6186 VSS -0.174f
C8320 VDD.n6187 VSS 0.00798f
C8321 VDD.n6188 VSS 0.00488f
C8322 VDD.n6189 VSS 4.74e-19
C8323 VDD.n6190 VSS 0.0422f
C8324 VDD.n6191 VSS 0.0515f
C8325 VDD.n6192 VSS 0.0202f
C8326 VDD.n6193 VSS 0.00277f
C8327 VDD.n6194 VSS 0.0129f
C8328 VDD.n6195 VSS 0.00979f
C8329 VDD.n6196 VSS 0.00979f
C8330 VDD.n6197 VSS 0.00332f
C8331 VDD.n6198 VSS 0.00663f
C8332 VDD.n6199 VSS 0.00806f
C8333 VDD.n6200 VSS 0.00411f
C8334 VDD.n6201 VSS 0.00585f
C8335 VDD.n6202 VSS 0.00472f
C8336 VDD.n6203 VSS 0.00439f
C8337 VDD.n6204 VSS 0.0136f
C8338 VDD.n6205 VSS 0.0141f
C8339 VDD.n6206 VSS 0.0223f
C8340 VDD.n6207 VSS 0.0227f
C8341 VDD.n6208 VSS 0.00798f
C8342 VDD.n6209 VSS 0.00488f
C8343 VDD.n6210 VSS 4.74e-19
C8344 VDD.n6211 VSS 0.00348f
C8345 VDD.n6212 VSS 3.16e-19
C8346 VDD.n6213 VSS 0.0104f
C8347 VDD.n6215 VSS 0.0129f
C8348 VDD.n6216 VSS 0.00979f
C8349 VDD.n6217 VSS 0.00979f
C8350 VDD.n6218 VSS 0.00332f
C8351 VDD.n6219 VSS 0.00663f
C8352 VDD.n6220 VSS 0.00806f
C8353 VDD.n6221 VSS 0.00585f
C8354 VDD.n6222 VSS 0.00411f
C8355 VDD.n6223 VSS 0.00332f
C8356 VDD.n6224 VSS -0.0753f
C8357 VDD.n6225 VSS 3.26e-19
C8358 VDD.n6226 VSS 0.00488f
C8359 VDD.n6227 VSS 0.00798f
C8360 VDD.n6228 VSS 0.0227f
C8361 VDD.n6229 VSS 0.0223f
C8362 VDD.n6230 VSS 0.0136f
C8363 VDD.n6231 VSS 0.00439f
C8364 VDD.n6232 VSS 0.00472f
C8365 VDD.n6233 VSS 0.00585f
C8366 VDD.n6234 VSS 0.00663f
C8367 VDD.n6235 VSS 0.00806f
C8368 VDD.n6236 VSS 0.00348f
C8369 VDD.n6237 VSS 0.00269f
C8370 VDD.n6238 VSS 0.00348f
C8371 VDD.n6239 VSS 3.16e-19
C8372 VDD.n6240 VSS 0.0104f
C8373 VDD.n6241 VSS 0.0129f
C8374 VDD.n6243 VSS 0.00277f
C8375 VDD.n6244 VSS 0.00269f
C8376 VDD.n6245 VSS 3.16e-19
C8377 VDD.n6246 VSS 0.00348f
C8378 VDD.n6247 VSS 4.74e-19
C8379 VDD.n6248 VSS 0.00488f
C8380 VDD.n6249 VSS 0.00798f
C8381 VDD.n6250 VSS -0.174f
C8382 VDD.n6251 VSS 0.0223f
C8383 VDD.n6252 VSS 0.0136f
C8384 VDD.n6253 VSS 0.00439f
C8385 VDD.n6254 VSS 0.00472f
C8386 VDD.n6255 VSS 0.00585f
C8387 VDD.n6256 VSS 0.00806f
C8388 VDD.n6257 VSS 0.00663f
C8389 VDD.n6258 VSS 0.00332f
C8390 VDD.n6259 VSS 0.00979f
C8391 VDD.n6260 VSS 0.00979f
C8392 VDD.n6261 VSS 0.0129f
C8393 VDD.n6263 VSS 0.00277f
C8394 VDD.n6264 VSS 0.0104f
C8395 VDD.n6265 VSS 3.16e-19
C8396 VDD.n6266 VSS 0.00348f
C8397 VDD.n6267 VSS 4.74e-19
C8398 VDD.n6268 VSS 0.00488f
C8399 VDD.n6269 VSS 0.00798f
C8400 VDD.n6270 VSS 0.0227f
C8401 VDD.n6271 VSS 0.0223f
C8402 VDD.n6272 VSS 0.0136f
C8403 VDD.n6273 VSS -0.0753f
C8404 VDD.n6274 VSS -0.211f
C8405 VDD.n6275 VSS 0.00585f
C8406 VDD.n6276 VSS 0.00806f
C8407 VDD.n6277 VSS 0.00663f
C8408 VDD.n6278 VSS 0.00332f
C8409 VDD.n6279 VSS 0.00979f
C8410 VDD.n6280 VSS 0.00979f
C8411 VDD.n6281 VSS 0.0129f
C8412 VDD.n6282 VSS 0.00277f
C8413 VDD.n6283 VSS 0.0234f
C8414 VDD.n6284 VSS 5.28e-19
C8415 VDD.n6285 VSS 0.00348f
C8416 VDD.n6286 VSS 4.74e-19
C8417 VDD.n6287 VSS 0.00488f
C8418 VDD.n6288 VSS 0.0286f
C8419 VDD.n6289 VSS 0.0805f
C8420 VDD.n6290 VSS 0.08f
C8421 VDD.n6291 VSS 0.0141f
C8422 VDD.n6292 VSS 0.0136f
C8423 VDD.n6293 VSS 3.26e-19
C8424 VDD.n6294 VSS 0.00472f
C8425 VDD.n6295 VSS 4.74e-19
C8426 VDD.n6296 VSS 0.00348f
C8427 VDD.n6297 VSS 5.28e-19
C8428 VDD.n6298 VSS 0.0234f
C8429 VDD.n6299 VSS 0.00277f
C8430 VDD.n6300 VSS 0.0129f
C8431 VDD.n6303 VSS 0.00277f
C8432 VDD.n6304 VSS 0.0104f
C8433 VDD.n6305 VSS 3.16e-19
C8434 VDD.n6306 VSS 0.00269f
C8435 VDD.n6307 VSS 0.00979f
C8436 VDD.n6308 VSS 0.00332f
C8437 VDD.n6309 VSS 0.00663f
C8438 VDD.n6310 VSS 0.00806f
C8439 VDD.n6311 VSS 0.00585f
C8440 VDD.n6312 VSS -0.211f
C8441 VDD.n6313 VSS 0.00391f
C8442 VDD.n6314 VSS 0.00472f
C8443 VDD.n6315 VSS 0.00781f
C8444 VDD.n6316 VSS 0.0223f
C8445 VDD.n6317 VSS 0.0136f
C8446 VDD.n6318 VSS -0.182f
C8447 VDD.n6319 VSS 0.00472f
C8448 VDD.n6320 VSS 0.00781f
C8449 VDD.n6321 VSS 0.00391f
C8450 VDD.n6322 VSS 0.0227f
C8451 VDD.n6323 VSS 0.0141f
C8452 VDD.n6324 VSS 0.00439f
C8453 VDD.n6325 VSS 0.00332f
C8454 VDD.n6326 VSS 0.00411f
C8455 VDD.n6327 VSS 0.00916f
C8456 VDD.n6328 VSS 0.00663f
C8457 VDD.n6329 VSS 0.00806f
C8458 VDD.n6330 VSS 0.00348f
C8459 VDD.n6331 VSS 0.00269f
C8460 VDD.n6332 VSS 0.00269f
C8461 VDD.n6333 VSS 3.16e-19
C8462 VDD.n6334 VSS 0.0104f
C8463 VDD.n6336 VSS 0.00277f
C8464 VDD.n6338 VSS 0.0129f
C8465 VDD.n6339 VSS 0.00979f
C8466 VDD.n6340 VSS 0.00979f
C8467 VDD.n6341 VSS 0.00332f
C8468 VDD.n6342 VSS 0.00348f
C8469 VDD.n6343 VSS 0.00806f
C8470 VDD.n6344 VSS 0.00663f
C8471 VDD.n6345 VSS 0.00916f
C8472 VDD.n6346 VSS 0.00411f
C8473 VDD.n6347 VSS 0.00332f
C8474 VDD.n6348 VSS 0.00439f
C8475 VDD.n6349 VSS 0.0141f
C8476 VDD.n6350 VSS 0.0227f
C8477 VDD.n6351 VSS 0.00391f
C8478 VDD.n6352 VSS 0.00781f
C8479 VDD.n6353 VSS 0.00472f
C8480 VDD.n6354 VSS 3.26e-19
C8481 VDD.n6355 VSS 0.0136f
C8482 VDD.n6356 VSS 0.0141f
C8483 VDD.n6357 VSS 0.0227f
C8484 VDD.n6358 VSS 0.00391f
C8485 VDD.n6359 VSS -0.211f
C8486 VDD.n6360 VSS 0.00585f
C8487 VDD.n6361 VSS 0.00411f
C8488 VDD.n6362 VSS 0.00916f
C8489 VDD.n6363 VSS 0.00348f
C8490 VDD.n6364 VSS 3.16e-19
C8491 VDD.n6365 VSS 0.00269f
C8492 VDD.n6366 VSS 0.00277f
C8493 VDD.n6368 VSS 0.0129f
C8494 VDD.n6370 VSS 0.0104f
C8495 VDD.n6371 VSS 3.16e-19
C8496 VDD.n6372 VSS 0.00348f
C8497 VDD.n6373 VSS 4.74e-19
C8498 VDD.n6374 VSS 0.00472f
C8499 VDD.n6375 VSS 3.26e-19
C8500 VDD.n6376 VSS 0.0136f
C8501 VDD.n6377 VSS 0.0141f
C8502 VDD.n6378 VSS 0.0227f
C8503 VDD.n6379 VSS 0.00391f
C8504 VDD.n6380 VSS 0.00488f
C8505 VDD.n6381 VSS 0.00585f
C8506 VDD.n6382 VSS 0.00806f
C8507 VDD.n6383 VSS 0.00663f
C8508 VDD.n6384 VSS 0.00332f
C8509 VDD.n6385 VSS 0.00979f
C8510 VDD.n6386 VSS 0.00979f
C8511 VDD.n6387 VSS 0.0129f
C8512 VDD.n6389 VSS 0.0173f
C8513 VDD.n6390 VSS 0.0312f
C8514 VDD.n6391 VSS 0.0312f
C8515 VDD.n6392 VSS 0.0173f
C8516 VDD.n6393 VSS 0.00277f
C8517 VDD.n6394 VSS 0.0104f
C8518 VDD.n6395 VSS 3.16e-19
C8519 VDD.n6396 VSS 0.00348f
C8520 VDD.n6397 VSS 4.74e-19
C8521 VDD.n6398 VSS 0.00472f
C8522 VDD.n6399 VSS 3.26e-19
C8523 VDD.n6400 VSS -0.0782f
C8524 VDD.n6401 VSS 0.0141f
C8525 VDD.n6402 VSS 0.06f
C8526 VDD.n6403 VSS 0.0243f
C8527 VDD.n6404 VSS 0.00488f
C8528 VDD.n6405 VSS 0.0251f
C8529 VDD.n6406 VSS 0.00411f
C8530 VDD.n6407 VSS 0.0251f
C8531 VDD.n6408 VSS 0.00472f
C8532 VDD.n6409 VSS 0.00439f
C8533 VDD.n6410 VSS 0.0136f
C8534 VDD.n6411 VSS -0.0845f
C8535 VDD.n6412 VSS -0.174f
C8536 VDD.n6413 VSS 0.00798f
C8537 VDD.n6414 VSS 0.00488f
C8538 VDD.n6415 VSS 4.74e-19
C8539 VDD.n6416 VSS 0.00348f
C8540 VDD.n6417 VSS 3.16e-19
C8541 VDD.n6418 VSS 0.0104f
C8542 VDD.n6420 VSS 0.0129f
C8543 VDD.n6421 VSS 0.00979f
C8544 VDD.n6422 VSS 0.00979f
C8545 VDD.n6423 VSS 0.00332f
C8546 VDD.n6424 VSS 0.00663f
C8547 VDD.n6425 VSS 0.00806f
C8548 VDD.n6426 VSS 0.00411f
C8549 VDD.n6427 VSS 0.00585f
C8550 VDD.n6428 VSS 0.00472f
C8551 VDD.n6429 VSS 0.00439f
C8552 VDD.n6430 VSS 0.0136f
C8553 VDD.n6431 VSS 0.0141f
C8554 VDD.n6432 VSS 0.0223f
C8555 VDD.n6433 VSS 0.0227f
C8556 VDD.n6434 VSS 0.00798f
C8557 VDD.n6435 VSS 0.00488f
C8558 VDD.n6436 VSS 4.74e-19
C8559 VDD.n6437 VSS 0.00348f
C8560 VDD.n6438 VSS 3.16e-19
C8561 VDD.n6439 VSS 0.0104f
C8562 VDD.n6441 VSS 0.0129f
C8563 VDD.n6442 VSS 0.00979f
C8564 VDD.n6443 VSS 0.00979f
C8565 VDD.n6444 VSS 0.00332f
C8566 VDD.n6445 VSS 0.00663f
C8567 VDD.n6446 VSS 0.00806f
C8568 VDD.n6447 VSS 0.00585f
C8569 VDD.n6448 VSS 0.00411f
C8570 VDD.n6449 VSS 0.00332f
C8571 VDD.n6450 VSS -0.0753f
C8572 VDD.n6451 VSS 3.26e-19
C8573 VDD.n6452 VSS 0.00488f
C8574 VDD.n6453 VSS 0.00798f
C8575 VDD.n6454 VSS 0.0227f
C8576 VDD.n6455 VSS 0.0223f
C8577 VDD.n6456 VSS 0.0136f
C8578 VDD.n6457 VSS 0.00439f
C8579 VDD.n6458 VSS 0.00472f
C8580 VDD.n6459 VSS 0.00585f
C8581 VDD.n6460 VSS 0.00663f
C8582 VDD.n6461 VSS 0.00806f
C8583 VDD.n6462 VSS 0.00348f
C8584 VDD.n6463 VSS 0.00269f
C8585 VDD.n6464 VSS 0.00348f
C8586 VDD.n6465 VSS 3.16e-19
C8587 VDD.n6466 VSS 0.0104f
C8588 VDD.n6467 VSS 0.0129f
C8589 VDD.n6469 VSS 0.00277f
C8590 VDD.n6470 VSS 0.00269f
C8591 VDD.n6471 VSS 3.16e-19
C8592 VDD.n6472 VSS 0.00348f
C8593 VDD.n6473 VSS 4.74e-19
C8594 VDD.n6474 VSS 0.00488f
C8595 VDD.n6475 VSS 0.00798f
C8596 VDD.n6476 VSS -0.174f
C8597 VDD.n6477 VSS 0.0223f
C8598 VDD.n6478 VSS 0.0136f
C8599 VDD.n6479 VSS 0.00439f
C8600 VDD.n6480 VSS 0.00472f
C8601 VDD.n6481 VSS 0.00585f
C8602 VDD.n6482 VSS 0.00806f
C8603 VDD.n6483 VSS 0.00663f
C8604 VDD.n6484 VSS 0.00332f
C8605 VDD.n6485 VSS 0.00979f
C8606 VDD.n6486 VSS 0.00979f
C8607 VDD.n6487 VSS 0.0129f
C8608 VDD.n6489 VSS 0.00277f
C8609 VDD.n6490 VSS 0.0104f
C8610 VDD.n6491 VSS 3.16e-19
C8611 VDD.n6492 VSS 0.00348f
C8612 VDD.n6493 VSS 4.74e-19
C8613 VDD.n6494 VSS 0.00488f
C8614 VDD.n6495 VSS 0.00798f
C8615 VDD.n6496 VSS 0.0227f
C8616 VDD.n6497 VSS 0.0223f
C8617 VDD.n6498 VSS 0.0136f
C8618 VDD.n6499 VSS -0.0753f
C8619 VDD.n6500 VSS -0.211f
C8620 VDD.n6501 VSS 0.00585f
C8621 VDD.n6502 VSS 0.00806f
C8622 VDD.n6503 VSS 0.00663f
C8623 VDD.n6504 VSS 0.00332f
C8624 VDD.n6505 VSS 0.00979f
C8625 VDD.n6506 VSS 0.00979f
C8626 VDD.n6507 VSS 0.0129f
C8627 VDD.n6508 VSS 0.00277f
C8628 VDD.n6509 VSS 0.0234f
C8629 VDD.n6510 VSS 5.28e-19
C8630 VDD.n6511 VSS 0.00348f
C8631 VDD.n6512 VSS 4.74e-19
C8632 VDD.n6513 VSS 0.00488f
C8633 VDD.n6514 VSS 0.0286f
C8634 VDD.n6515 VSS 0.0805f
C8635 VDD.n6516 VSS 0.08f
C8636 VDD.n6517 VSS 0.0141f
C8637 VDD.n6518 VSS 0.0136f
C8638 VDD.n6519 VSS 3.26e-19
C8639 VDD.n6520 VSS 0.00472f
C8640 VDD.n6521 VSS 4.74e-19
C8641 VDD.n6522 VSS 0.00348f
C8642 VDD.n6523 VSS 5.28e-19
C8643 VDD.n6524 VSS 0.0234f
C8644 VDD.n6525 VSS 0.00277f
C8645 VDD.n6526 VSS 0.0129f
C8646 VDD.n6529 VSS 0.00277f
C8647 VDD.n6530 VSS 0.0104f
C8648 VDD.n6531 VSS 3.16e-19
C8649 VDD.n6532 VSS 0.00269f
C8650 VDD.n6533 VSS 0.00979f
C8651 VDD.n6534 VSS 0.00332f
C8652 VDD.n6535 VSS 0.00663f
C8653 VDD.n6536 VSS 0.00806f
C8654 VDD.n6537 VSS 0.00585f
C8655 VDD.n6538 VSS -0.211f
C8656 VDD.n6539 VSS 0.00391f
C8657 VDD.n6540 VSS 0.00472f
C8658 VDD.n6541 VSS 0.00781f
C8659 VDD.n6542 VSS 0.0223f
C8660 VDD.n6543 VSS 0.0136f
C8661 VDD.n6544 VSS -0.182f
C8662 VDD.n6545 VSS 0.00472f
C8663 VDD.n6546 VSS 0.00781f
C8664 VDD.n6547 VSS 0.00391f
C8665 VDD.n6548 VSS 0.0227f
C8666 VDD.n6549 VSS 0.0141f
C8667 VDD.n6550 VSS 0.00439f
C8668 VDD.n6551 VSS 0.00332f
C8669 VDD.n6552 VSS 0.00411f
C8670 VDD.n6553 VSS 0.00916f
C8671 VDD.n6554 VSS 0.00663f
C8672 VDD.n6555 VSS 0.00806f
C8673 VDD.n6556 VSS 0.00348f
C8674 VDD.n6557 VSS 0.00269f
C8675 VDD.n6558 VSS 0.00269f
C8676 VDD.n6559 VSS 3.16e-19
C8677 VDD.n6560 VSS 0.0104f
C8678 VDD.n6562 VSS 0.00277f
C8679 VDD.n6564 VSS 0.0129f
C8680 VDD.n6565 VSS 0.00979f
C8681 VDD.n6566 VSS 0.00979f
C8682 VDD.n6567 VSS 0.00332f
C8683 VDD.n6568 VSS 0.00348f
C8684 VDD.n6569 VSS 0.00806f
C8685 VDD.n6570 VSS 0.00663f
C8686 VDD.n6571 VSS 0.00916f
C8687 VDD.n6572 VSS 0.00411f
C8688 VDD.n6573 VSS 0.00332f
C8689 VDD.n6574 VSS 0.00439f
C8690 VDD.n6575 VSS 0.0141f
C8691 VDD.n6576 VSS 0.0227f
C8692 VDD.n6577 VSS 0.00391f
C8693 VDD.n6578 VSS 0.00781f
C8694 VDD.n6579 VSS 0.00472f
C8695 VDD.n6580 VSS 3.26e-19
C8696 VDD.n6581 VSS 0.0136f
C8697 VDD.n6582 VSS 0.0141f
C8698 VDD.n6583 VSS 0.0227f
C8699 VDD.n6584 VSS 0.00391f
C8700 VDD.n6585 VSS -0.211f
C8701 VDD.n6586 VSS 0.00585f
C8702 VDD.n6587 VSS 0.00411f
C8703 VDD.n6588 VSS 0.00916f
C8704 VDD.n6589 VSS 0.00348f
C8705 VDD.n6590 VSS 3.16e-19
C8706 VDD.n6591 VSS 0.00269f
C8707 VDD.n6592 VSS 0.00277f
C8708 VDD.n6594 VSS 0.0129f
C8709 VDD.n6596 VSS 0.0104f
C8710 VDD.n6597 VSS 3.16e-19
C8711 VDD.n6598 VSS 0.00348f
C8712 VDD.n6599 VSS 4.74e-19
C8713 VDD.n6600 VSS 0.00472f
C8714 VDD.n6601 VSS 3.26e-19
C8715 VDD.n6602 VSS 0.0136f
C8716 VDD.n6603 VSS 0.0141f
C8717 VDD.n6604 VSS 0.0227f
C8718 VDD.n6605 VSS 0.00391f
C8719 VDD.n6606 VSS 0.00488f
C8720 VDD.n6607 VSS 0.00585f
C8721 VDD.n6608 VSS 0.00806f
C8722 VDD.n6609 VSS 0.00663f
C8723 VDD.n6610 VSS 0.00332f
C8724 VDD.n6611 VSS 0.00979f
C8725 VDD.n6612 VSS 0.00979f
C8726 VDD.n6613 VSS 0.0129f
C8727 VDD.n6615 VSS 0.0173f
C8728 VDD.n6616 VSS 0.0312f
C8729 VDD.n6617 VSS 0.0312f
C8730 VDD.n6618 VSS 0.0173f
C8731 VDD.n6619 VSS 0.00277f
C8732 VDD.n6620 VSS 0.0104f
C8733 VDD.n6621 VSS 3.16e-19
C8734 VDD.n6622 VSS 0.00348f
C8735 VDD.n6623 VSS 4.74e-19
C8736 VDD.n6624 VSS 0.00472f
C8737 VDD.n6625 VSS 3.26e-19
C8738 VDD.n6626 VSS -0.0782f
C8739 VDD.n6627 VSS 0.0141f
C8740 VDD.n6628 VSS 0.06f
C8741 VDD.n6629 VSS 0.0243f
C8742 VDD.n6630 VSS 0.00488f
C8743 VDD.n6631 VSS 0.0251f
C8744 VDD.n6632 VSS 0.00411f
C8745 VDD.n6633 VSS 0.0251f
C8746 VDD.n6634 VSS 0.00472f
C8747 VDD.n6635 VSS 0.00439f
C8748 VDD.n6636 VSS 0.0136f
C8749 VDD.n6637 VSS -0.0845f
C8750 VDD.n6638 VSS -0.174f
C8751 VDD.n6639 VSS 0.00798f
C8752 VDD.n6640 VSS 0.00488f
C8753 VDD.n6641 VSS 4.74e-19
C8754 VDD.n6642 VSS 0.00348f
C8755 VDD.n6643 VSS 3.16e-19
C8756 VDD.n6644 VSS 0.0104f
C8757 VDD.n6646 VSS 0.0129f
C8758 VDD.n6647 VSS 0.00979f
C8759 VDD.n6648 VSS 0.00979f
C8760 VDD.n6649 VSS 0.00332f
C8761 VDD.n6650 VSS 0.00663f
C8762 VDD.n6651 VSS 0.00806f
C8763 VDD.n6652 VSS 0.00411f
C8764 VDD.n6653 VSS 0.00585f
C8765 VDD.n6654 VSS 0.00472f
C8766 VDD.n6655 VSS 0.00439f
C8767 VDD.n6656 VSS 0.0136f
C8768 VDD.n6657 VSS 0.0141f
C8769 VDD.n6658 VSS 0.0223f
C8770 VDD.n6659 VSS 0.0227f
C8771 VDD.n6660 VSS 0.00798f
C8772 VDD.n6661 VSS 0.00488f
C8773 VDD.n6662 VSS 4.74e-19
C8774 VDD.n6663 VSS 0.00348f
C8775 VDD.n6664 VSS 3.16e-19
C8776 VDD.n6665 VSS 0.0104f
C8777 VDD.n6667 VSS 0.0129f
C8778 VDD.n6668 VSS 0.00979f
C8779 VDD.n6669 VSS 0.00979f
C8780 VDD.n6670 VSS 0.00332f
C8781 VDD.n6671 VSS 0.00663f
C8782 VDD.n6672 VSS 0.00806f
C8783 VDD.n6673 VSS 0.00585f
C8784 VDD.n6674 VSS 0.00411f
C8785 VDD.n6675 VSS 0.00332f
C8786 VDD.n6676 VSS -0.0753f
C8787 VDD.n6677 VSS 3.26e-19
C8788 VDD.n6678 VSS 0.00488f
C8789 VDD.n6679 VSS 0.00798f
C8790 VDD.n6680 VSS 0.0227f
C8791 VDD.n6681 VSS 0.0223f
C8792 VDD.n6682 VSS 0.0136f
C8793 VDD.n6683 VSS 0.00439f
C8794 VDD.n6684 VSS 0.00472f
C8795 VDD.n6685 VSS 0.00585f
C8796 VDD.n6686 VSS 0.00663f
C8797 VDD.n6687 VSS 0.00806f
C8798 VDD.n6688 VSS 0.00348f
C8799 VDD.n6689 VSS 0.00269f
C8800 VDD.n6690 VSS 0.00348f
C8801 VDD.n6691 VSS 3.16e-19
C8802 VDD.n6692 VSS 0.0104f
C8803 VDD.n6693 VSS 0.0129f
C8804 VDD.n6695 VSS 0.00277f
C8805 VDD.n6696 VSS 0.00269f
C8806 VDD.n6697 VSS 3.16e-19
C8807 VDD.n6698 VSS 0.00348f
C8808 VDD.n6699 VSS 4.74e-19
C8809 VDD.n6700 VSS 0.00488f
C8810 VDD.n6701 VSS 0.00798f
C8811 VDD.n6702 VSS -0.174f
C8812 VDD.n6703 VSS 0.0223f
C8813 VDD.n6704 VSS 0.0136f
C8814 VDD.n6705 VSS 0.00439f
C8815 VDD.n6706 VSS 0.00472f
C8816 VDD.n6707 VSS 0.00585f
C8817 VDD.n6708 VSS 0.00806f
C8818 VDD.n6709 VSS 0.00663f
C8819 VDD.n6710 VSS 0.00332f
C8820 VDD.n6711 VSS 0.00979f
C8821 VDD.n6712 VSS 0.00979f
C8822 VDD.n6713 VSS 0.0129f
C8823 VDD.n6715 VSS 0.00277f
C8824 VDD.n6716 VSS 0.0104f
C8825 VDD.n6717 VSS 3.16e-19
C8826 VDD.n6718 VSS 0.00348f
C8827 VDD.n6719 VSS 4.74e-19
C8828 VDD.n6720 VSS 0.00488f
C8829 VDD.n6721 VSS 0.00798f
C8830 VDD.n6722 VSS 0.0227f
C8831 VDD.n6723 VSS 0.0223f
C8832 VDD.n6724 VSS 0.0136f
C8833 VDD.n6725 VSS -0.0753f
C8834 VDD.n6726 VSS -0.211f
C8835 VDD.n6727 VSS 0.00585f
C8836 VDD.n6728 VSS 0.00806f
C8837 VDD.n6729 VSS 0.00663f
C8838 VDD.n6730 VSS 0.00332f
C8839 VDD.n6731 VSS 0.00979f
C8840 VDD.n6732 VSS 0.00979f
C8841 VDD.n6733 VSS 0.0129f
C8842 VDD.n6734 VSS 0.00277f
C8843 VDD.n6735 VSS 0.0234f
C8844 VDD.n6736 VSS 5.28e-19
C8845 VDD.n6737 VSS 0.00348f
C8846 VDD.n6738 VSS 4.74e-19
C8847 VDD.n6739 VSS 0.00488f
C8848 VDD.n6740 VSS 0.0286f
C8849 VDD.n6741 VSS 0.0805f
C8850 VDD.n6742 VSS 0.08f
C8851 VDD.n6743 VSS 0.0141f
C8852 VDD.n6744 VSS 0.0136f
C8853 VDD.n6745 VSS 3.26e-19
C8854 VDD.n6746 VSS 0.00472f
C8855 VDD.n6747 VSS 4.74e-19
C8856 VDD.n6748 VSS 0.00348f
C8857 VDD.n6749 VSS 5.28e-19
C8858 VDD.n6750 VSS 0.0234f
C8859 VDD.n6751 VSS 0.00277f
C8860 VDD.n6752 VSS 0.0129f
C8861 VDD.n6755 VSS 0.00277f
C8862 VDD.n6756 VSS 0.0104f
C8863 VDD.n6757 VSS 3.16e-19
C8864 VDD.n6758 VSS 0.00269f
C8865 VDD.n6759 VSS 0.00979f
C8866 VDD.n6760 VSS 0.00332f
C8867 VDD.n6761 VSS 0.00663f
C8868 VDD.n6762 VSS 0.00806f
C8869 VDD.n6763 VSS 0.00585f
C8870 VDD.n6764 VSS -0.211f
C8871 VDD.n6765 VSS 0.00391f
C8872 VDD.n6766 VSS 0.00472f
C8873 VDD.n6767 VSS 0.00781f
C8874 VDD.n6768 VSS 0.0223f
C8875 VDD.n6769 VSS 0.0136f
C8876 VDD.n6770 VSS -0.182f
C8877 VDD.n6771 VSS 0.00472f
C8878 VDD.n6772 VSS 0.00781f
C8879 VDD.n6773 VSS 0.00391f
C8880 VDD.n6774 VSS 0.0227f
C8881 VDD.n6775 VSS 0.0141f
C8882 VDD.n6776 VSS 0.00439f
C8883 VDD.n6777 VSS 0.00332f
C8884 VDD.n6778 VSS 0.00411f
C8885 VDD.n6779 VSS 0.00916f
C8886 VDD.n6780 VSS 0.00663f
C8887 VDD.n6781 VSS 0.00806f
C8888 VDD.n6782 VSS 0.00348f
C8889 VDD.n6783 VSS 0.00269f
C8890 VDD.n6784 VSS 0.00269f
C8891 VDD.n6785 VSS 3.16e-19
C8892 VDD.n6786 VSS 0.0104f
C8893 VDD.n6788 VSS 0.00277f
C8894 VDD.n6790 VSS 0.0129f
C8895 VDD.n6791 VSS 0.00979f
C8896 VDD.n6792 VSS 0.00979f
C8897 VDD.n6793 VSS 0.00332f
C8898 VDD.n6794 VSS 0.00348f
C8899 VDD.n6795 VSS 0.00806f
C8900 VDD.n6796 VSS 0.00663f
C8901 VDD.n6797 VSS 0.00916f
C8902 VDD.n6798 VSS 0.00411f
C8903 VDD.n6799 VSS 0.00332f
C8904 VDD.n6800 VSS 0.00439f
C8905 VDD.n6801 VSS 0.0141f
C8906 VDD.n6802 VSS 0.0227f
C8907 VDD.n6803 VSS 0.00391f
C8908 VDD.n6804 VSS 0.00781f
C8909 VDD.n6805 VSS 0.00472f
C8910 VDD.n6806 VSS 3.26e-19
C8911 VDD.n6807 VSS 0.0136f
C8912 VDD.n6808 VSS 0.0141f
C8913 VDD.n6809 VSS 0.0227f
C8914 VDD.n6810 VSS 0.00391f
C8915 VDD.n6811 VSS -0.211f
C8916 VDD.n6812 VSS 0.00585f
C8917 VDD.n6813 VSS 0.00411f
C8918 VDD.n6814 VSS 0.00916f
C8919 VDD.n6815 VSS 0.00348f
C8920 VDD.n6816 VSS 3.16e-19
C8921 VDD.n6817 VSS 0.00269f
C8922 VDD.n6818 VSS 0.00277f
C8923 VDD.n6820 VSS 0.0129f
C8924 VDD.n6822 VSS 0.0104f
C8925 VDD.n6823 VSS 3.16e-19
C8926 VDD.n6824 VSS 0.00348f
C8927 VDD.n6825 VSS 4.74e-19
C8928 VDD.n6826 VSS 0.00472f
C8929 VDD.n6827 VSS 3.26e-19
C8930 VDD.n6828 VSS 0.0136f
C8931 VDD.n6829 VSS 0.0141f
C8932 VDD.n6830 VSS 0.0227f
C8933 VDD.n6831 VSS 0.00391f
C8934 VDD.n6832 VSS 0.00488f
C8935 VDD.n6833 VSS 0.00585f
C8936 VDD.n6834 VSS 0.00806f
C8937 VDD.n6835 VSS 0.00663f
C8938 VDD.n6836 VSS 0.00332f
C8939 VDD.n6837 VSS 0.00979f
C8940 VDD.n6838 VSS 0.00979f
C8941 VDD.n6839 VSS 0.0129f
C8942 VDD.n6841 VSS 0.0173f
C8943 VDD.n6842 VSS 0.0312f
C8944 VDD.n6843 VSS 0.0312f
C8945 VDD.n6844 VSS 0.0173f
C8946 VDD.n6845 VSS 0.00277f
C8947 VDD.n6846 VSS 0.0104f
C8948 VDD.n6847 VSS 3.16e-19
C8949 VDD.n6848 VSS 0.00348f
C8950 VDD.n6849 VSS 4.74e-19
C8951 VDD.n6850 VSS 0.00472f
C8952 VDD.n6851 VSS 3.26e-19
C8953 VDD.n6852 VSS -0.0782f
C8954 VDD.n6853 VSS 0.0141f
C8955 VDD.n6854 VSS 0.06f
C8956 VDD.n6855 VSS 0.0243f
C8957 VDD.n6856 VSS 0.00488f
C8958 VDD.n6857 VSS 0.0251f
C8959 VDD.n6858 VSS 0.00411f
C8960 VDD.n6859 VSS 0.0251f
C8961 VDD.n6860 VSS 0.00472f
C8962 VDD.n6861 VSS 0.00439f
C8963 VDD.n6862 VSS 0.0136f
C8964 VDD.n6863 VSS -0.0845f
C8965 VDD.n6864 VSS -0.174f
C8966 VDD.n6865 VSS 0.00798f
C8967 VDD.n6866 VSS 0.00488f
C8968 VDD.n6867 VSS 4.74e-19
C8969 VDD.n6868 VSS 0.00348f
C8970 VDD.n6869 VSS 3.16e-19
C8971 VDD.n6870 VSS 0.0104f
C8972 VDD.n6872 VSS 0.0129f
C8973 VDD.n6873 VSS 0.00979f
C8974 VDD.n6874 VSS 0.00979f
C8975 VDD.n6875 VSS 0.00332f
C8976 VDD.n6876 VSS 0.00663f
C8977 VDD.n6877 VSS 0.00806f
C8978 VDD.n6878 VSS 0.00411f
C8979 VDD.n6879 VSS 0.00585f
C8980 VDD.n6880 VSS 0.00472f
C8981 VDD.n6881 VSS 0.00439f
C8982 VDD.n6882 VSS 0.0136f
C8983 VDD.n6883 VSS 0.0141f
C8984 VDD.n6884 VSS 0.0223f
C8985 VDD.n6885 VSS 0.0227f
C8986 VDD.n6886 VSS 0.00798f
C8987 VDD.n6887 VSS 0.00488f
C8988 VDD.n6888 VSS 4.74e-19
C8989 VDD.n6889 VSS 0.00348f
C8990 VDD.n6890 VSS 3.16e-19
C8991 VDD.n6891 VSS 0.0104f
C8992 VDD.n6893 VSS 0.0129f
C8993 VDD.n6894 VSS 0.00979f
C8994 VDD.n6895 VSS 0.00979f
C8995 VDD.n6896 VSS 0.00332f
C8996 VDD.n6897 VSS 0.00663f
C8997 VDD.n6898 VSS 0.00806f
C8998 VDD.n6899 VSS 0.00585f
C8999 VDD.n6900 VSS 0.00411f
C9000 VDD.n6901 VSS 0.00332f
C9001 VDD.n6902 VSS -0.0753f
C9002 VDD.n6903 VSS 3.26e-19
C9003 VDD.n6904 VSS 0.00488f
C9004 VDD.n6905 VSS 0.00798f
C9005 VDD.n6906 VSS 0.0227f
C9006 VDD.n6907 VSS 0.0223f
C9007 VDD.n6908 VSS 0.0136f
C9008 VDD.n6909 VSS 0.00439f
C9009 VDD.n6910 VSS 0.00472f
C9010 VDD.n6911 VSS 0.00585f
C9011 VDD.n6912 VSS 0.00663f
C9012 VDD.n6913 VSS 0.00806f
C9013 VDD.n6914 VSS 0.00348f
C9014 VDD.n6915 VSS 0.00269f
C9015 VDD.n6916 VSS 0.00348f
C9016 VDD.n6917 VSS 3.16e-19
C9017 VDD.n6918 VSS 0.0104f
C9018 VDD.n6919 VSS 0.0129f
C9019 VDD.n6921 VSS 0.00277f
C9020 VDD.n6922 VSS 0.00269f
C9021 VDD.n6923 VSS 3.16e-19
C9022 VDD.n6924 VSS 0.00348f
C9023 VDD.n6925 VSS 4.74e-19
C9024 VDD.n6926 VSS 0.00488f
C9025 VDD.n6927 VSS 0.00798f
C9026 VDD.n6928 VSS -0.174f
C9027 VDD.n6929 VSS 0.0223f
C9028 VDD.n6930 VSS 0.0136f
C9029 VDD.n6931 VSS 0.00439f
C9030 VDD.n6932 VSS 0.00472f
C9031 VDD.n6933 VSS 0.00585f
C9032 VDD.n6934 VSS 0.00806f
C9033 VDD.n6935 VSS 0.00663f
C9034 VDD.n6936 VSS 0.00332f
C9035 VDD.n6937 VSS 0.00979f
C9036 VDD.n6938 VSS 0.00979f
C9037 VDD.n6939 VSS 0.0129f
C9038 VDD.n6941 VSS 0.00277f
C9039 VDD.n6942 VSS 0.0104f
C9040 VDD.n6943 VSS 3.16e-19
C9041 VDD.n6944 VSS 0.00348f
C9042 VDD.n6945 VSS 4.74e-19
C9043 VDD.n6946 VSS 0.00488f
C9044 VDD.n6947 VSS 0.00798f
C9045 VDD.n6948 VSS 0.0227f
C9046 VDD.n6949 VSS 0.0223f
C9047 VDD.n6950 VSS 0.0136f
C9048 VDD.n6951 VSS -0.0753f
C9049 VDD.n6952 VSS -0.211f
C9050 VDD.n6953 VSS 0.00585f
C9051 VDD.n6954 VSS 0.00806f
C9052 VDD.n6955 VSS 0.00663f
C9053 VDD.n6956 VSS 0.00332f
C9054 VDD.n6957 VSS 0.00979f
C9055 VDD.n6958 VSS 0.00979f
C9056 VDD.n6959 VSS 0.0129f
C9057 VDD.n6960 VSS 0.00277f
C9058 VDD.n6961 VSS 0.0234f
C9059 VDD.n6962 VSS 5.28e-19
C9060 VDD.n6963 VSS 0.00348f
C9061 VDD.n6964 VSS 4.74e-19
C9062 VDD.n6965 VSS 0.00488f
C9063 VDD.n6966 VSS 0.0286f
C9064 VDD.n6967 VSS 0.0805f
C9065 VDD.n6968 VSS 0.08f
C9066 VDD.n6969 VSS 0.0141f
C9067 VDD.n6970 VSS 0.0136f
C9068 VDD.n6971 VSS 3.26e-19
C9069 VDD.n6972 VSS 0.00472f
C9070 VDD.n6973 VSS 4.74e-19
C9071 VDD.n6974 VSS 0.00348f
C9072 VDD.n6975 VSS 5.28e-19
C9073 VDD.n6976 VSS 0.0234f
C9074 VDD.n6977 VSS 0.00277f
C9075 VDD.n6978 VSS 0.0129f
C9076 VDD.n6981 VSS 0.00277f
C9077 VDD.n6982 VSS 0.0104f
C9078 VDD.n6983 VSS 3.16e-19
C9079 VDD.n6984 VSS 0.00269f
C9080 VDD.n6985 VSS 0.00979f
C9081 VDD.n6986 VSS 0.00332f
C9082 VDD.n6987 VSS 0.00663f
C9083 VDD.n6988 VSS 0.00806f
C9084 VDD.n6989 VSS 0.00585f
C9085 VDD.n6990 VSS -0.211f
C9086 VDD.n6991 VSS 0.00391f
C9087 VDD.n6992 VSS 0.00472f
C9088 VDD.n6993 VSS 0.00781f
C9089 VDD.n6994 VSS 0.0223f
C9090 VDD.n6995 VSS 0.0136f
C9091 VDD.n6996 VSS -0.182f
C9092 VDD.n6997 VSS 0.00472f
C9093 VDD.n6998 VSS 0.00781f
C9094 VDD.n6999 VSS 0.00391f
C9095 VDD.n7000 VSS 0.0227f
C9096 VDD.n7001 VSS 0.0141f
C9097 VDD.n7002 VSS 0.00439f
C9098 VDD.n7003 VSS 0.00332f
C9099 VDD.n7004 VSS 0.00411f
C9100 VDD.n7005 VSS 0.00916f
C9101 VDD.n7006 VSS 0.00663f
C9102 VDD.n7007 VSS 0.00806f
C9103 VDD.n7008 VSS 0.00348f
C9104 VDD.n7009 VSS 0.00269f
C9105 VDD.n7010 VSS 0.00269f
C9106 VDD.n7011 VSS 3.16e-19
C9107 VDD.n7012 VSS 0.0104f
C9108 VDD.n7014 VSS 0.00277f
C9109 VDD.n7016 VSS 0.0129f
C9110 VDD.n7017 VSS 0.00979f
C9111 VDD.n7018 VSS 0.00979f
C9112 VDD.n7019 VSS 0.00332f
C9113 VDD.n7020 VSS 0.00348f
C9114 VDD.n7021 VSS 0.00806f
C9115 VDD.n7022 VSS 0.00663f
C9116 VDD.n7023 VSS 0.00916f
C9117 VDD.n7024 VSS 0.00411f
C9118 VDD.n7025 VSS 0.00332f
C9119 VDD.n7026 VSS 0.00439f
C9120 VDD.n7027 VSS 0.0141f
C9121 VDD.n7028 VSS 0.0227f
C9122 VDD.n7029 VSS 0.00391f
C9123 VDD.n7030 VSS 0.00781f
C9124 VDD.n7031 VSS 0.00472f
C9125 VDD.n7032 VSS 3.26e-19
C9126 VDD.n7033 VSS 0.0136f
C9127 VDD.n7034 VSS 0.0141f
C9128 VDD.n7035 VSS 0.0227f
C9129 VDD.n7036 VSS 0.00391f
C9130 VDD.n7037 VSS -0.211f
C9131 VDD.n7038 VSS 0.00585f
C9132 VDD.n7039 VSS 0.00411f
C9133 VDD.n7040 VSS 0.00916f
C9134 VDD.n7041 VSS 0.00348f
C9135 VDD.n7042 VSS 3.16e-19
C9136 VDD.n7043 VSS 0.00269f
C9137 VDD.n7044 VSS 0.00277f
C9138 VDD.n7046 VSS 0.0129f
C9139 VDD.n7048 VSS 0.0104f
C9140 VDD.n7049 VSS 3.16e-19
C9141 VDD.n7050 VSS 0.00348f
C9142 VDD.n7051 VSS 4.74e-19
C9143 VDD.n7052 VSS 0.00472f
C9144 VDD.n7053 VSS 3.26e-19
C9145 VDD.n7054 VSS 0.0136f
C9146 VDD.n7055 VSS 0.0141f
C9147 VDD.n7056 VSS 0.00472f
C9148 VDD.n7057 VSS 3.26e-19
C9149 VDD.n7058 VSS -0.0782f
C9150 VDD.n7059 VSS -0.182f
C9151 VDD.n7060 VSS 0.0227f
C9152 VDD.n7061 VSS 0.00391f
C9153 VDD.n7062 VSS 0.00488f
C9154 VDD.n7063 VSS 0.00585f
C9155 VDD.n7064 VSS 0.00348f
C9156 VDD.n7065 VSS 0.00806f
C9157 VDD.n7066 VSS 0.00663f
C9158 VDD.n7067 VSS 0.00332f
C9159 VDD.n7068 VSS 0.00979f
C9160 VDD.n7069 VSS 0.00979f
C9161 VDD.n7070 VSS 0.0129f
C9162 VDD.n7071 VSS 0.0202f
C9163 VDD.n7072 VSS 0.0515f
C9164 VDD.n7073 VSS 0.0422f
C9165 VDD.n7074 VSS 0.0389f
C9166 VDD.n7075 VSS 0.0398f
C9167 VDD.n7076 VSS 0.0601f
C9168 VDD.n7077 VSS 0.619f
C9169 VDD.n7078 VSS 0.646f
C9170 VDD.n7079 VSS 0.063f
C9171 VDD.n7080 VSS 0.0439f
C9172 VDD.n7081 VSS 0.0433f
C9173 VDD.n7082 VSS 0.00585f
C9174 VDD.n7083 VSS 0.00332f
C9175 VDD.n7084 VSS 0.00348f
C9176 VDD.n7085 VSS 0.00806f
C9177 VDD.n7086 VSS 0.00663f
C9178 VDD.n7087 VSS 0.0095f
C9179 VDD.n7088 VSS 0.00411f
C9180 VDD.n7089 VSS 0.00332f
C9181 VDD.n7090 VSS -0.0753f
C9182 VDD.n7091 VSS 0.0143f
C9183 VDD.n7092 VSS 0.0231f
C9184 VDD.n7093 VSS 0.00391f
C9185 VDD.n7094 VSS 0.00781f
C9186 VDD.n7095 VSS 0.00472f
C9187 VDD.n7096 VSS 3.26e-19
C9188 VDD.n7097 VSS 0.0139f
C9189 VDD.n7098 VSS 0.0143f
C9190 VDD.n7099 VSS 0.0143f
C9191 VDD.n7100 VSS 0.00472f
C9192 VDD.n7101 VSS 0.00488f
C9193 VDD.n7102 VSS 4.74e-19
C9194 VDD.n7103 VSS 0.00585f
C9195 VDD.n7104 VSS 0.00348f
C9196 VDD.n7105 VSS 0.00332f
C9197 VDD.n7106 VSS 4.74e-19
C9198 VDD.n7107 VSS 0.00348f
C9199 VDD.n7108 VSS 0.00979f
C9200 VDD.n7109 VSS 0.00979f
C9201 VDD.n7110 VSS 0.00332f
C9202 VDD.n7111 VSS 0.00348f
C9203 VDD.n7112 VSS 0.00269f
C9204 VDD.n7113 VSS 0.00269f
C9205 VDD.n7114 VSS 0.0104f
C9206 VDD.n7115 VSS 3.16e-19
C9207 VDD.n7116 VSS 0.00277f
C9208 VDD.n7117 VSS 0.00269f
C9209 VDD.n7118 VSS 0.00979f
C9210 VDD.n7119 VSS 0.00979f
C9211 VDD.n7120 VSS 0.00269f
C9212 VDD.n7121 VSS 0.00663f
C9213 VDD.n7122 VSS 0.00348f
C9214 VDD.n7123 VSS 0.00806f
C9215 VDD.n7124 VSS 0.00332f
C9216 VDD.n7125 VSS 0.00781f
C9217 VDD.n7126 VSS 0.00439f
C9218 VDD.n7127 VSS 0.0143f
C9219 VDD.n7128 VSS 0.00472f
C9220 VDD.n7129 VSS 0.0231f
C9221 VDD.n7130 VSS 0.00391f
C9222 VDD.n7131 VSS 0.00781f
C9223 VDD.n7132 VSS 0.0226f
C9224 VDD.n7133 VSS 0.0139f
C9225 VDD.n7134 VSS 3.26e-19
C9226 VDD.n7135 VSS -0.0753f
C9227 VDD.n7136 VSS 0.00332f
C9228 VDD.n7137 VSS 0.00916f
C9229 VDD.n7138 VSS 0.00411f
C9230 VDD.n7139 VSS 0.00585f
C9231 VDD.n7140 VSS -0.211f
C9232 VDD.n7141 VSS 0.00391f
C9233 VDD.n7142 VSS 0.0231f
C9234 VDD.n7143 VSS 0.0226f
C9235 VDD.n7144 VSS -0.181f
C9236 VDD.n7145 VSS 0.00488f
C9237 VDD.n7146 VSS 3.26e-19
C9238 VDD.n7147 VSS 0.00348f
C9239 VDD.n7148 VSS 0.00411f
C9240 VDD.n7149 VSS 0.00779f
C9241 VDD.n7150 VSS 0.00488f
C9242 VDD.n7151 VSS -0.078f
C9243 VDD.n7152 VSS 0.0305f
C9244 VDD.n7153 VSS 0.00618f
C9245 VDD.n7154 VSS 0.00816f
C9246 VDD.n7155 VSS 0.00767f
C9247 VDD.n7156 VSS 0.0305f
C9248 VDD.n7157 VSS 0.0143f
C9249 VDD.n7158 VSS 0.00439f
C9250 VDD.n7159 VSS 0.00332f
C9251 VDD.n7160 VSS 0.00269f
C9252 VDD.n7161 VSS 0.0104f
C9253 VDD.n7162 VSS 3.16e-19
C9254 VDD.n7163 VSS 0.00269f
C9255 VDD.n7164 VSS 0.00277f
C9256 VDD.n7165 VSS 0.0129f
C9257 VDD.n7166 VSS 0.00979f
C9258 VDD.n7167 VSS 0.00916f
C9259 VDD.n7168 VSS 0.00411f
C9260 VDD.n7169 VSS 0.00585f
C9261 VDD.n7170 VSS 0.00806f
C9262 VDD.n7171 VSS 0.00663f
C9263 VDD.n7172 VSS 0.00332f
C9264 VDD.n7173 VSS 0.00979f
C9265 VDD.n7174 VSS 0.00269f
C9266 VDD.n7175 VSS 0.0104f
C9267 VDD.n7176 VSS 3.16e-19
C9268 VDD.n7177 VSS 0.00348f
C9269 VDD.n7178 VSS 4.74e-19
C9270 VDD.n7179 VSS 0.00472f
C9271 VDD.n7180 VSS 0.00781f
C9272 VDD.n7181 VSS 0.00391f
C9273 VDD.n7182 VSS 0.0231f
C9274 VDD.n7183 VSS 0.0143f
C9275 VDD.n7184 VSS 0.0139f
C9276 VDD.n7185 VSS 3.26e-19
C9277 VDD.n7186 VSS 0.00472f
C9278 VDD.n7187 VSS 4.74e-19
C9279 VDD.n7188 VSS 0.00348f
C9280 VDD.n7189 VSS 0.00269f
C9281 VDD.n7190 VSS 0.00332f
C9282 VDD.n7191 VSS 0.00979f
C9283 VDD.n7192 VSS 0.00979f
C9284 VDD.n7193 VSS 0.00277f
C9285 VDD.n7194 VSS 0.00269f
C9286 VDD.n7195 VSS 0.0104f
C9287 VDD.n7196 VSS 3.16e-19
C9288 VDD.n7197 VSS 0.00269f
C9289 VDD.n7198 VSS 0.00269f
C9290 VDD.n7199 VSS 0.00348f
C9291 VDD.n7200 VSS 0.00806f
C9292 VDD.n7201 VSS 0.00663f
C9293 VDD.n7202 VSS 0.00916f
C9294 VDD.n7203 VSS 0.00411f
C9295 VDD.n7204 VSS 0.00332f
C9296 VDD.n7205 VSS 0.00439f
C9297 VDD.n7206 VSS 3.26e-19
C9298 VDD.n7207 VSS -0.078f
C9299 VDD.n7208 VSS -0.181f
C9300 VDD.n7209 VSS 0.0231f
C9301 VDD.n7210 VSS 0.00391f
C9302 VDD.n7211 VSS 0.00488f
C9303 VDD.n7212 VSS 0.00585f
C9304 VDD.n7213 VSS 0.00411f
C9305 VDD.n7214 VSS 0.00916f
C9306 VDD.n7215 VSS 0.00348f
C9307 VDD.n7216 VSS 3.16e-19
C9308 VDD.n7217 VSS 0.0104f
C9309 VDD.n7218 VSS 0.0129f
C9310 VDD.n7219 VSS 0.00979f
C9311 VDD.n7220 VSS 0.00269f
C9312 VDD.n7221 VSS 0.0314f
C9313 VDD.n7222 VSS 0.0236f
C9314 VDD.n7223 VSS 0.46f
C9315 VDD.n7224 VSS 0.0173f
C9316 VDD.n7225 VSS 0.0102f
C9317 VDD.n7226 VSS 0.0633f
C9318 VDD.t61 VSS 0.00583f
C9319 VDD.n7227 VSS 0.0579f
C9320 VDD.n7228 VSS 0.0361f
C9321 VDD.n7229 VSS 0.0174f
C9322 VDD.n7230 VSS 0.00106f
C9323 VDD.n7231 VSS 0.0166f
C9324 VDD.n7232 VSS 0.384f
C9325 VDD.n7233 VSS 0.502f
C9326 VDD.n7234 VSS 0.602f
C9327 VDD.n7235 VSS 0.004f
C9328 VDD.n7236 VSS 0.024f
C9329 VDD.n7237 VSS 0.0606f
C9330 VDD.n7238 VSS 0.0274f
C9331 VDD.n7239 VSS 0.0124f
C9332 VDD.n7240 VSS 8.15e-19
C9333 VDD.n7241 VSS 0.0261f
C9334 VDD.n7242 VSS 0.02f
C9335 VDD.n7243 VSS 0.00689f
C9336 VDD.n7244 VSS 0.0111f
C9337 VDD.n7245 VSS 0.0186f
C9338 VDD.n7246 VSS 0.0409f
C9339 VDD.n7247 VSS 0.016f
C9340 VDD.n7248 VSS 0.0124f
C9341 VDD.n7249 VSS 0.00989f
C9342 VDD.n7250 VSS 0.0214f
C9343 VDD.t55 VSS 0.0509f
C9344 VDD.n7251 VSS 0.0931f
C9345 VDD.n7252 VSS 0.0202f
C9346 VDD.n7253 VSS 0.00797f
C9347 VDD.n7254 VSS 0.0556f
C9348 VDD.n7255 VSS 0.0225f
C9349 VDD.n7256 VSS 0.0211f
C9350 VDD.n7257 VSS 0.0197f
C9351 VDD.n7258 VSS 8.15e-19
C9352 VDD.n7259 VSS 0.0232f
C9353 VDD.n7260 VSS 0.017f
C9354 VDD.n7261 VSS 0.0069f
C9355 VDD.n7262 VSS 0.0124f
C9356 VDD.n7263 VSS 0.00461f
C9357 VDD.n7264 VSS 0.00483f
C9358 VDD.n7265 VSS 0.00184f
C9359 VDD.n7266 VSS 0.0109f
C9360 VDD.n7267 VSS 0.0108f
C9361 VDD.n7268 VSS 0.00256f
C9362 VDD.n7269 VSS 0.0124f
C9363 VDD.n7270 VSS 0.00163f
C9364 VDD.t42 VSS 0.125f
C9365 VDD.t54 VSS 0.103f
C9366 VDD.n7271 VSS 0.0755f
C9367 VDD.n7272 VSS 0.0149f
C9368 VDD.n7273 VSS 0.0914f
C9369 VDD.n7274 VSS 0.014f
C9370 VDD.n7275 VSS 0.00135f
C9371 VDD.n7276 VSS 0.00256f
C9372 VDD.n7277 VSS 0.00391f
C9373 VDD.n7278 VSS 0.00391f
C9374 VDD.n7279 VSS 0.0184f
C9375 VDD.n7280 VSS 0.0106f
C9376 VDD.n7281 VSS 0.0273f
C9377 VDD.n7282 VSS 0.0198f
C9378 VDD.n7283 VSS 0.0172f
C9379 sample_delay_offset.n0 VSS 0.00153f
C9380 sample_delay_offset.t5 VSS 0.0258f
C9381 sample_delay_offset.t9 VSS 0.0156f
C9382 sample_delay_offset.n1 VSS 0.0192f
C9383 sample_delay_offset.n2 VSS 0.0299f
C9384 sample_delay_offset.n3 VSS 0.0634f
C9385 sample_delay_offset.n4 VSS 0.0226f
C9386 sample_delay_offset.n5 VSS 0.234f
C9387 sample_delay_offset.t3 VSS 0.0137f
C9388 sample_delay_offset.n6 VSS 0.00687f
C9389 sample_delay_offset.t0 VSS 0.0258f
C9390 sample_delay_offset.t8 VSS 0.0162f
C9391 sample_delay_offset.n7 VSS 0.0487f
C9392 sample_delay_offset.n8 VSS 0.0097f
C9393 sample_delay_offset.n9 VSS 0.00293f
C9394 sample_delay_offset.n10 VSS 0.00236f
C9395 sample_delay_offset.n11 VSS 0.0027f
C9396 sample_delay_offset.n12 VSS 0.0114f
C9397 sample_delay_offset.n13 VSS 0.117f
C9398 sample_delay_offset.n14 VSS 0.259f
C9399 sample_delay_offset.t6 VSS 0.0137f
C9400 sample_delay_offset.n15 VSS 0.202f
C9401 sample_delay_offset.n16 VSS 1.44f
C9402 sample_delay_offset.n17 VSS 0.00687f
C9403 sample_delay_offset.t7 VSS 0.0258f
C9404 sample_delay_offset.t4 VSS 0.0162f
C9405 sample_delay_offset.n18 VSS 0.0487f
C9406 sample_delay_offset.n19 VSS 0.0097f
C9407 sample_delay_offset.n20 VSS 0.00293f
C9408 sample_delay_offset.n21 VSS 0.00236f
C9409 sample_delay_offset.n22 VSS 0.0027f
C9410 sample_delay_offset.n23 VSS 0.0114f
C9411 sample_delay_offset.n24 VSS 0.117f
C9412 sample_delay_offset.n25 VSS 0.259f
C9413 sample_delay_offset.t10 VSS 0.0137f
C9414 sample_delay_offset.n26 VSS 0.202f
C9415 sample_delay_offset.n27 VSS 0.331f
C9416 sample_delay_offset.n28 VSS 0.00153f
C9417 sample_delay_offset.t11 VSS 0.0258f
C9418 sample_delay_offset.t1 VSS 0.0156f
C9419 sample_delay_offset.n29 VSS 0.0192f
C9420 sample_delay_offset.n30 VSS 0.0299f
C9421 sample_delay_offset.n31 VSS 0.0634f
C9422 sample_delay_offset.n32 VSS 0.0226f
C9423 sample_delay_offset.n33 VSS 0.234f
C9424 sample_delay_offset.n34 VSS 0.106f
C9425 sample_delay_offset.t2 VSS 0.0137f
C9426 sample_delay_offset.n35 VSS 0.387f
C9427 sample_delay_offset.n36 VSS 1.95f
C9428 sample_delay_offset.n37 VSS 2.41f
C9429 sample_delay_offset.n38 VSS 3.16f
C9430 sample_delay_offset.n39 VSS 0.3f
C9431 sample_delay_offset.n40 VSS 0.106f
.ends

