magic
tech sky130A
timestamp 1698670603
<< pwell >>
rect 6617 -2967 6633 -2942
use hgu_cdac_cap_2  hgu_cdac_cap_2_0
timestamp 1698486325
transform 1 0 50 0 1 -3716
box -1470 13 -1134 1207
use hgu_cdac_cap_4  hgu_cdac_cap_4_0
timestamp 1698626624
transform 1 0 -1460 0 1 -5102
box 343 1399 982 2593
use hgu_cdac_cap_8  hgu_cdac_cap_8_0
timestamp 1698618791
transform 1 0 -854 0 1 -5102
box 343 1399 1588 2593
use hgu_cdac_cap_16  hgu_cdac_cap_16_0
timestamp 1698619766
transform 1 0 249 0 1 -7591
box 452 3888 2909 5082
use hgu_cdac_cap_32  hgu_cdac_cap_32_0
timestamp 1698622076
transform 1 0 -6419 0 1 -2445
box 9544 -1258 14425 -64
use hgu_cdac_cap_64  hgu_cdac_cap_64_0
timestamp 1698625969
transform 1 0 -8163 0 1 -5117
box 16136 1414 25865 2608
use hgu_cdac_unit  hgu_cdac_unit_0
timestamp 1698670284
transform 1 0 -2066 0 1 -3422
box 343 299 679 913
use hgu_cdac_unit  x1
timestamp 1698670284
transform 1 0 -2066 0 1 -4002
box 343 299 679 913
<< labels >>
flabel pwell 6617 -2967 6633 -2942 0 FreeSans 80 0 0 0 SUB
port 1 nsew
<< end >>
