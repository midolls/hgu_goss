* NGSPICE file created from test.ext - technology: sky130A

.subckt test vdd output input vss
X0 output input vdd vdd sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X1 output input vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
C0 input vdd 0.192f
C1 output vdd 0.166f
C2 input output 0.238f
.ends

