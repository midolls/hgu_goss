magic
tech sky130A
magscale 1 2
timestamp 1698061451
<< nwell >>
rect 991 5890 4184 6250
rect 992 5888 4176 5890
rect 984 5014 13040 5375
rect 544 4321 13040 4686
rect 3130 3771 13034 3821
rect 3132 3457 13034 3771
rect 996 2894 13031 2940
rect 996 2585 13028 2894
<< pwell >>
rect 993 5576 4167 5849
rect 1030 4706 12994 4978
rect 597 4016 12994 4282
rect 3210 3144 12993 3404
rect 1034 2271 12993 2555
<< psubdiff >>
rect 1035 5586 1064 5620
rect 1098 5586 1156 5620
rect 1190 5586 1248 5620
rect 1282 5586 1340 5620
rect 1374 5586 1432 5620
rect 1466 5586 1524 5620
rect 1558 5586 1616 5620
rect 1650 5586 1708 5620
rect 1742 5586 1800 5620
rect 1834 5586 1892 5620
rect 1926 5586 1984 5620
rect 2018 5586 2076 5620
rect 2110 5586 2168 5620
rect 2202 5586 2260 5620
rect 2294 5586 2352 5620
rect 2386 5586 2444 5620
rect 2478 5586 2536 5620
rect 2570 5586 2628 5620
rect 2662 5586 2720 5620
rect 2754 5586 2812 5620
rect 2846 5586 2904 5620
rect 2938 5586 2996 5620
rect 3030 5586 3088 5620
rect 3122 5586 3180 5620
rect 3214 5586 3272 5620
rect 3306 5586 3364 5620
rect 3398 5586 3456 5620
rect 3490 5586 3548 5620
rect 3582 5586 3640 5620
rect 3674 5586 3732 5620
rect 3766 5586 3824 5620
rect 3858 5586 3916 5620
rect 3950 5586 4008 5620
rect 4042 5586 4135 5620
rect 1034 4713 1063 4747
rect 1097 4713 1155 4747
rect 1189 4713 1247 4747
rect 1281 4713 1339 4747
rect 1373 4713 1431 4747
rect 1465 4713 1523 4747
rect 1557 4713 1615 4747
rect 1649 4713 1707 4747
rect 1741 4713 1799 4747
rect 1833 4713 1891 4747
rect 1925 4713 1983 4747
rect 2017 4713 2075 4747
rect 2109 4713 2167 4747
rect 2201 4713 2259 4747
rect 2293 4713 2351 4747
rect 2385 4713 2443 4747
rect 2477 4713 2535 4747
rect 2569 4713 2627 4747
rect 2661 4713 2719 4747
rect 2753 4713 2811 4747
rect 2845 4713 2903 4747
rect 2937 4713 2995 4747
rect 3029 4713 3087 4747
rect 3121 4713 3179 4747
rect 3213 4713 3271 4747
rect 3305 4713 3363 4747
rect 3397 4713 3455 4747
rect 3489 4713 3547 4747
rect 3581 4713 3639 4747
rect 3673 4713 3731 4747
rect 3765 4713 3823 4747
rect 3857 4713 3915 4747
rect 3949 4713 4007 4747
rect 4041 4713 4099 4747
rect 4133 4713 4191 4747
rect 4225 4713 4283 4747
rect 4317 4713 4375 4747
rect 4409 4713 4467 4747
rect 4501 4713 4559 4747
rect 4593 4713 4651 4747
rect 4685 4713 4743 4747
rect 4777 4713 4835 4747
rect 4869 4713 4927 4747
rect 4961 4713 5019 4747
rect 5053 4713 5111 4747
rect 5145 4713 5203 4747
rect 5237 4713 5295 4747
rect 5329 4713 5387 4747
rect 5421 4713 5479 4747
rect 5513 4713 5571 4747
rect 5605 4713 5663 4747
rect 5697 4713 5755 4747
rect 5789 4713 5847 4747
rect 5881 4713 5939 4747
rect 5973 4713 6031 4747
rect 6065 4713 6123 4747
rect 6157 4713 6215 4747
rect 6249 4713 6307 4747
rect 6341 4713 6399 4747
rect 6433 4713 6491 4747
rect 6525 4713 6583 4747
rect 6617 4713 6675 4747
rect 6709 4713 6767 4747
rect 6801 4713 6859 4747
rect 6893 4713 6951 4747
rect 6985 4713 7043 4747
rect 7077 4713 7135 4747
rect 7169 4713 7227 4747
rect 7261 4713 7319 4747
rect 7353 4713 7411 4747
rect 7445 4713 7503 4747
rect 7537 4713 7595 4747
rect 7629 4713 7687 4747
rect 7721 4713 7779 4747
rect 7813 4713 7871 4747
rect 7905 4713 7963 4747
rect 7997 4713 8055 4747
rect 8089 4713 8147 4747
rect 8181 4713 8239 4747
rect 8273 4713 8331 4747
rect 8365 4713 8423 4747
rect 8457 4713 8515 4747
rect 8549 4713 8607 4747
rect 8641 4713 8699 4747
rect 8733 4713 8791 4747
rect 8825 4713 8883 4747
rect 8917 4713 8975 4747
rect 9009 4713 9067 4747
rect 9101 4713 9159 4747
rect 9193 4713 9251 4747
rect 9285 4713 9343 4747
rect 9377 4713 9435 4747
rect 9469 4713 9527 4747
rect 9561 4713 9619 4747
rect 9653 4713 9711 4747
rect 9745 4713 9803 4747
rect 9837 4713 9895 4747
rect 9929 4713 9987 4747
rect 10021 4713 10079 4747
rect 10113 4713 10171 4747
rect 10205 4713 10263 4747
rect 10297 4713 10355 4747
rect 10389 4713 10447 4747
rect 10481 4713 10539 4747
rect 10573 4713 10631 4747
rect 10665 4713 10723 4747
rect 10757 4713 10815 4747
rect 10849 4713 10907 4747
rect 10941 4713 10999 4747
rect 11033 4713 11091 4747
rect 11125 4713 11183 4747
rect 11217 4713 11275 4747
rect 11309 4713 11367 4747
rect 11401 4713 11459 4747
rect 11493 4713 11551 4747
rect 11585 4713 11643 4747
rect 11677 4713 11735 4747
rect 11769 4713 11827 4747
rect 11861 4713 11919 4747
rect 11953 4713 12011 4747
rect 12045 4713 12103 4747
rect 12137 4713 12195 4747
rect 12229 4713 12287 4747
rect 12321 4713 12379 4747
rect 12413 4713 12471 4747
rect 12505 4713 12563 4747
rect 12597 4713 12655 4747
rect 12689 4713 12747 4747
rect 12781 4713 12839 4747
rect 12873 4713 12931 4747
rect 12965 4713 12994 4747
rect 594 4024 623 4058
rect 657 4024 715 4058
rect 749 4024 807 4058
rect 841 4024 899 4058
rect 933 4024 991 4058
rect 1025 4024 1083 4058
rect 1117 4024 1175 4058
rect 1209 4024 1267 4058
rect 1301 4024 1359 4058
rect 1393 4024 1451 4058
rect 1485 4024 1543 4058
rect 1577 4024 1635 4058
rect 1669 4024 1727 4058
rect 1761 4024 1819 4058
rect 1853 4024 1911 4058
rect 1945 4024 2003 4058
rect 2037 4024 2095 4058
rect 2129 4024 2187 4058
rect 2221 4024 2279 4058
rect 2313 4024 2371 4058
rect 2405 4024 2463 4058
rect 2497 4024 2555 4058
rect 2589 4024 2647 4058
rect 2681 4024 2739 4058
rect 2773 4024 2831 4058
rect 2865 4024 2923 4058
rect 2957 4024 3015 4058
rect 3049 4024 3107 4058
rect 3141 4024 3199 4058
rect 3233 4024 3291 4058
rect 3325 4024 3383 4058
rect 3417 4024 3475 4058
rect 3509 4024 3567 4058
rect 3601 4024 3659 4058
rect 3693 4024 3751 4058
rect 3785 4024 3843 4058
rect 3877 4024 3935 4058
rect 3969 4024 4027 4058
rect 4061 4024 4119 4058
rect 4153 4024 4211 4058
rect 4245 4024 4303 4058
rect 4337 4024 4395 4058
rect 4429 4024 4487 4058
rect 4521 4024 4579 4058
rect 4613 4024 4671 4058
rect 4705 4024 4763 4058
rect 4797 4024 4855 4058
rect 4889 4024 4947 4058
rect 4981 4024 5039 4058
rect 5073 4024 5131 4058
rect 5165 4024 5223 4058
rect 5257 4024 5315 4058
rect 5349 4024 5407 4058
rect 5441 4024 5499 4058
rect 5533 4024 5591 4058
rect 5625 4024 5683 4058
rect 5717 4024 5775 4058
rect 5809 4024 5867 4058
rect 5901 4024 5959 4058
rect 5993 4024 6051 4058
rect 6085 4024 6143 4058
rect 6177 4024 6235 4058
rect 6269 4024 6327 4058
rect 6361 4024 6419 4058
rect 6453 4024 6511 4058
rect 6545 4024 6603 4058
rect 6637 4024 6695 4058
rect 6729 4024 6787 4058
rect 6821 4024 6879 4058
rect 6913 4024 6971 4058
rect 7005 4024 7063 4058
rect 7097 4024 7155 4058
rect 7189 4024 7247 4058
rect 7281 4024 7339 4058
rect 7373 4024 7431 4058
rect 7465 4024 7523 4058
rect 7557 4024 7615 4058
rect 7649 4024 7707 4058
rect 7741 4024 7799 4058
rect 7833 4024 7891 4058
rect 7925 4024 7983 4058
rect 8017 4024 8075 4058
rect 8109 4024 8167 4058
rect 8201 4024 8259 4058
rect 8293 4024 8351 4058
rect 8385 4024 8443 4058
rect 8477 4024 8535 4058
rect 8569 4024 8627 4058
rect 8661 4024 8719 4058
rect 8753 4024 8811 4058
rect 8845 4024 8903 4058
rect 8937 4024 8995 4058
rect 9029 4024 9087 4058
rect 9121 4024 9179 4058
rect 9213 4024 9271 4058
rect 9305 4024 9363 4058
rect 9397 4024 9435 4058
rect 9469 4024 9527 4058
rect 9561 4024 9619 4058
rect 9653 4024 9711 4058
rect 9745 4024 9803 4058
rect 9837 4024 9895 4058
rect 9929 4024 9987 4058
rect 10021 4024 10079 4058
rect 10113 4024 10171 4058
rect 10205 4024 10263 4058
rect 10297 4024 10355 4058
rect 10389 4024 10447 4058
rect 10481 4024 10539 4058
rect 10573 4024 10631 4058
rect 10665 4024 10723 4058
rect 10757 4024 10815 4058
rect 10849 4024 10907 4058
rect 10941 4024 10999 4058
rect 11033 4024 11091 4058
rect 11125 4024 11183 4058
rect 11217 4024 11275 4058
rect 11309 4024 11367 4058
rect 11401 4024 11459 4058
rect 11493 4024 11551 4058
rect 11585 4024 11643 4058
rect 11677 4024 11735 4058
rect 11769 4024 11827 4058
rect 11861 4024 11919 4058
rect 11953 4024 12011 4058
rect 12045 4024 12103 4058
rect 12137 4024 12195 4058
rect 12229 4024 12287 4058
rect 12321 4024 12379 4058
rect 12413 4024 12471 4058
rect 12505 4024 12563 4058
rect 12597 4024 12655 4058
rect 12689 4024 12747 4058
rect 12781 4024 12839 4058
rect 12873 4024 12931 4058
rect 12965 4024 12994 4058
rect 3167 3151 3197 3185
rect 3231 3151 3289 3185
rect 3323 3151 3381 3185
rect 3415 3151 3473 3185
rect 3507 3151 3565 3185
rect 3599 3151 3657 3185
rect 3691 3151 3749 3185
rect 3783 3151 3841 3185
rect 3875 3151 3933 3185
rect 3967 3151 4025 3185
rect 4059 3151 4117 3185
rect 4151 3151 4209 3185
rect 4243 3151 4301 3185
rect 4335 3151 4393 3185
rect 4427 3151 4485 3185
rect 4519 3151 4577 3185
rect 4611 3151 4669 3185
rect 4703 3151 4761 3185
rect 4795 3151 4853 3185
rect 4887 3151 4945 3185
rect 4979 3151 5037 3185
rect 5071 3151 5129 3185
rect 5163 3151 5221 3185
rect 5255 3151 5313 3185
rect 5347 3151 5405 3185
rect 5439 3151 5497 3185
rect 5531 3151 5589 3185
rect 5623 3151 5681 3185
rect 5715 3151 5773 3185
rect 5807 3151 5865 3185
rect 5899 3151 5957 3185
rect 5991 3151 6049 3185
rect 6083 3151 6141 3185
rect 6175 3151 6233 3185
rect 6267 3151 6325 3185
rect 6359 3151 6417 3185
rect 6451 3151 6509 3185
rect 6543 3151 6601 3185
rect 6635 3151 6693 3185
rect 6727 3151 6785 3185
rect 6819 3151 6877 3185
rect 6911 3151 6969 3185
rect 7003 3151 7061 3185
rect 7095 3151 7153 3185
rect 7187 3151 7245 3185
rect 7279 3151 7337 3185
rect 7371 3151 7429 3185
rect 7463 3151 7521 3185
rect 7555 3151 7613 3185
rect 7647 3151 7705 3185
rect 7739 3151 7797 3185
rect 7831 3151 7889 3185
rect 7923 3151 7981 3185
rect 8015 3151 8073 3185
rect 8107 3151 8165 3185
rect 8199 3151 8257 3185
rect 8291 3151 8349 3185
rect 8383 3151 8441 3185
rect 8475 3151 8533 3185
rect 8567 3151 8625 3185
rect 8659 3151 8717 3185
rect 8751 3151 8809 3185
rect 8843 3151 8901 3185
rect 8935 3151 8993 3185
rect 9027 3151 9085 3185
rect 9119 3151 9177 3185
rect 9211 3151 9269 3185
rect 9303 3151 9361 3185
rect 9395 3151 9453 3185
rect 9487 3151 9545 3185
rect 9579 3151 9637 3185
rect 9671 3151 9729 3185
rect 9763 3151 9821 3185
rect 9855 3151 9894 3185
rect 9947 3151 9986 3185
rect 10039 3151 10078 3185
rect 10131 3151 10170 3185
rect 10223 3151 10262 3185
rect 10315 3151 10354 3185
rect 10407 3151 10446 3185
rect 10499 3151 10538 3185
rect 10591 3151 10630 3185
rect 10683 3151 10722 3185
rect 10775 3151 10814 3185
rect 10867 3151 10906 3185
rect 10959 3151 10998 3185
rect 11051 3151 11090 3185
rect 11143 3151 11182 3185
rect 11235 3151 11274 3185
rect 11327 3151 11366 3185
rect 11419 3151 11458 3185
rect 11511 3151 11550 3185
rect 11603 3151 11642 3185
rect 11695 3151 11734 3185
rect 11787 3151 11826 3185
rect 11879 3151 11918 3185
rect 11971 3151 12010 3185
rect 12044 3151 12102 3185
rect 12136 3151 12194 3185
rect 12228 3151 12286 3185
rect 12320 3151 12378 3185
rect 12412 3151 12470 3185
rect 12504 3151 12562 3185
rect 12596 3151 12654 3185
rect 12688 3151 12746 3185
rect 12780 3151 12838 3185
rect 12872 3151 12930 3185
rect 12964 3151 12992 3185
rect 1033 2278 1062 2312
rect 1096 2278 1154 2312
rect 1188 2278 1246 2312
rect 1280 2278 1338 2312
rect 1372 2278 1430 2312
rect 1464 2278 1522 2312
rect 1556 2278 1614 2312
rect 1648 2278 1706 2312
rect 1740 2278 1798 2312
rect 1832 2278 1890 2312
rect 1924 2278 1982 2312
rect 2016 2278 2074 2312
rect 2108 2278 2166 2312
rect 2200 2278 2258 2312
rect 2292 2278 2350 2312
rect 2384 2278 2442 2312
rect 2476 2278 2534 2312
rect 2568 2278 2626 2312
rect 2660 2278 2718 2312
rect 2752 2278 2810 2312
rect 2844 2278 2902 2312
rect 2936 2278 2994 2312
rect 3028 2278 3086 2312
rect 3120 2278 3178 2312
rect 3212 2278 3270 2312
rect 3304 2278 3362 2312
rect 3396 2278 3454 2312
rect 3488 2278 3546 2312
rect 3580 2278 3638 2312
rect 3672 2278 3730 2312
rect 3764 2278 3822 2312
rect 3856 2278 3914 2312
rect 3948 2278 4006 2312
rect 4040 2278 4098 2312
rect 4132 2278 4190 2312
rect 4224 2278 4282 2312
rect 4316 2278 4374 2312
rect 4408 2278 4466 2312
rect 4500 2278 4558 2312
rect 4592 2278 4650 2312
rect 4684 2278 4742 2312
rect 4776 2278 4834 2312
rect 4868 2278 4926 2312
rect 4960 2278 5018 2312
rect 5052 2278 5110 2312
rect 5144 2278 5202 2312
rect 5236 2278 5294 2312
rect 5328 2278 5386 2312
rect 5420 2278 5478 2312
rect 5512 2278 5570 2312
rect 5604 2278 5662 2312
rect 5696 2278 5754 2312
rect 5788 2278 5846 2312
rect 5880 2278 5938 2312
rect 5972 2278 6030 2312
rect 6064 2278 6122 2312
rect 6156 2278 6214 2312
rect 6248 2278 6306 2312
rect 6340 2278 6398 2312
rect 6432 2278 6490 2312
rect 6524 2278 6582 2312
rect 6616 2278 6674 2312
rect 6708 2278 6766 2312
rect 6800 2278 6858 2312
rect 6892 2278 6950 2312
rect 6984 2278 7042 2312
rect 7076 2278 7134 2312
rect 7168 2278 7226 2312
rect 7260 2278 7318 2312
rect 7352 2278 7410 2312
rect 7444 2278 7502 2312
rect 7536 2278 7594 2312
rect 7628 2278 7686 2312
rect 7720 2278 7778 2312
rect 7812 2278 7870 2312
rect 7904 2278 7962 2312
rect 7996 2278 8054 2312
rect 8088 2278 8146 2312
rect 8180 2278 8238 2312
rect 8272 2278 8330 2312
rect 8364 2278 8422 2312
rect 8456 2278 8514 2312
rect 8548 2278 8606 2312
rect 8640 2278 8698 2312
rect 8732 2278 8790 2312
rect 8824 2278 8882 2312
rect 8916 2278 8974 2312
rect 9008 2278 9066 2312
rect 9100 2278 9158 2312
rect 9192 2278 9250 2312
rect 9284 2278 9342 2312
rect 9376 2278 9434 2312
rect 9468 2278 9526 2312
rect 9560 2278 9618 2312
rect 9652 2278 9710 2312
rect 9744 2278 9802 2312
rect 9836 2278 9894 2312
rect 9928 2278 9986 2312
rect 10020 2278 10078 2312
rect 10112 2278 10170 2312
rect 10204 2278 10262 2312
rect 10296 2278 10354 2312
rect 10388 2278 10446 2312
rect 10480 2278 10538 2312
rect 10572 2278 10630 2312
rect 10664 2278 10722 2312
rect 10756 2278 10814 2312
rect 10848 2278 10906 2312
rect 10940 2278 10998 2312
rect 11032 2278 11090 2312
rect 11124 2278 11182 2312
rect 11216 2278 11274 2312
rect 11308 2278 11366 2312
rect 11400 2278 11458 2312
rect 11492 2278 11550 2312
rect 11584 2278 11642 2312
rect 11676 2278 11734 2312
rect 11768 2278 11826 2312
rect 11860 2278 11918 2312
rect 11952 2278 12010 2312
rect 12044 2278 12102 2312
rect 12136 2278 12194 2312
rect 12228 2278 12286 2312
rect 12320 2278 12378 2312
rect 12412 2278 12470 2312
rect 12504 2278 12562 2312
rect 12596 2278 12654 2312
rect 12688 2278 12746 2312
rect 12780 2278 12838 2312
rect 12872 2278 12930 2312
rect 12964 2278 12993 2312
<< nsubdiff >>
rect 1035 6178 1064 6212
rect 1098 6178 1156 6212
rect 1190 6178 1248 6212
rect 1282 6178 1340 6212
rect 1374 6178 1432 6212
rect 1466 6178 1524 6212
rect 1558 6178 1616 6212
rect 1650 6178 1679 6212
rect 2295 6178 2324 6212
rect 2358 6178 2416 6212
rect 2450 6178 2508 6212
rect 2542 6178 2600 6212
rect 2634 6178 2692 6212
rect 2726 6178 2784 6212
rect 2818 6178 2876 6212
rect 2910 6178 2968 6212
rect 3002 6178 3060 6212
rect 3094 6178 3152 6212
rect 3186 6178 3244 6212
rect 3278 6178 3336 6212
rect 3370 6178 3428 6212
rect 3462 6178 3520 6212
rect 3554 6178 3612 6212
rect 3646 6178 3704 6212
rect 3738 6178 3796 6212
rect 3830 6178 3888 6212
rect 3922 6178 3980 6212
rect 4014 6178 4072 6212
rect 4106 6178 4135 6212
rect 1034 5305 1063 5339
rect 1097 5305 1155 5339
rect 1189 5305 1247 5339
rect 1281 5305 1339 5339
rect 1373 5305 1431 5339
rect 1465 5305 1523 5339
rect 1557 5305 1615 5339
rect 1649 5305 1707 5339
rect 1741 5305 1799 5339
rect 1833 5305 1891 5339
rect 1925 5305 1983 5339
rect 2017 5305 2075 5339
rect 2109 5305 2167 5339
rect 2201 5305 2259 5339
rect 2293 5305 2351 5339
rect 2385 5305 2443 5339
rect 2477 5305 2535 5339
rect 2569 5305 2627 5339
rect 2661 5305 2719 5339
rect 2753 5305 2811 5339
rect 2845 5305 2895 5339
rect 3007 5305 3087 5339
rect 3121 5305 3179 5339
rect 3213 5305 3271 5339
rect 3305 5305 3363 5339
rect 3397 5305 3455 5339
rect 3489 5305 3547 5339
rect 3581 5305 3640 5339
rect 3674 5305 3731 5339
rect 3765 5305 3823 5339
rect 3857 5305 3915 5339
rect 3949 5305 4007 5339
rect 4041 5305 4139 5339
rect 4249 5305 4283 5339
rect 4317 5305 4375 5339
rect 4409 5305 4467 5339
rect 4501 5305 4559 5339
rect 4593 5305 4651 5339
rect 4685 5305 4743 5339
rect 4777 5305 4835 5339
rect 4869 5305 4927 5339
rect 4961 5305 5019 5339
rect 5053 5305 5111 5339
rect 5145 5305 5203 5339
rect 5237 5305 5295 5339
rect 5329 5305 5387 5339
rect 5421 5305 5479 5339
rect 5513 5305 5571 5339
rect 5605 5305 5663 5339
rect 5697 5305 5755 5339
rect 5789 5305 5847 5339
rect 5881 5305 5939 5339
rect 5973 5305 6031 5339
rect 6065 5305 6123 5339
rect 6157 5305 6215 5339
rect 6249 5305 6307 5339
rect 6341 5305 6399 5339
rect 6433 5305 6531 5339
rect 6641 5305 6675 5339
rect 6709 5305 6767 5339
rect 6801 5305 6859 5339
rect 6893 5305 6951 5339
rect 6985 5305 7043 5339
rect 7077 5305 7135 5339
rect 7169 5305 7227 5339
rect 7261 5305 7319 5339
rect 7353 5305 7411 5339
rect 7445 5305 7503 5339
rect 7537 5305 7595 5339
rect 7629 5305 7687 5339
rect 7721 5305 7779 5339
rect 7813 5305 7871 5339
rect 7905 5305 7963 5339
rect 7997 5305 8055 5339
rect 8089 5305 8147 5339
rect 8181 5305 8239 5339
rect 8273 5305 8331 5339
rect 8365 5305 8423 5339
rect 8457 5305 8515 5339
rect 8549 5305 8607 5339
rect 8641 5305 8699 5339
rect 8733 5305 8791 5339
rect 8825 5305 8923 5339
rect 9033 5305 9067 5339
rect 9101 5305 9159 5339
rect 9193 5305 9251 5339
rect 9285 5305 9343 5339
rect 9377 5305 9435 5339
rect 9469 5305 9527 5339
rect 9561 5305 9619 5339
rect 9653 5305 9711 5339
rect 9745 5305 9803 5339
rect 9837 5305 9895 5339
rect 9929 5305 9987 5339
rect 10021 5305 10079 5339
rect 10113 5305 10171 5339
rect 10205 5305 10263 5339
rect 10297 5305 10355 5339
rect 10389 5305 10447 5339
rect 10481 5305 10539 5339
rect 10573 5305 10631 5339
rect 10665 5305 10723 5339
rect 10757 5305 10815 5339
rect 10849 5305 10907 5339
rect 10941 5305 10999 5339
rect 11033 5305 11091 5339
rect 11125 5305 11183 5339
rect 11217 5305 11315 5339
rect 11425 5305 11459 5339
rect 11493 5305 11551 5339
rect 11585 5305 11643 5339
rect 11677 5305 11735 5339
rect 11769 5305 11827 5339
rect 11861 5305 11919 5339
rect 11953 5305 12011 5339
rect 12045 5305 12103 5339
rect 12137 5305 12195 5339
rect 12229 5305 12287 5339
rect 12321 5305 12379 5339
rect 12413 5305 12471 5339
rect 12505 5305 12563 5339
rect 12597 5305 12655 5339
rect 12689 5305 12747 5339
rect 12781 5305 12839 5339
rect 12873 5305 12931 5339
rect 12965 5305 12994 5339
rect 594 4616 623 4650
rect 657 4616 715 4650
rect 749 4616 807 4650
rect 841 4616 899 4650
rect 933 4616 991 4650
rect 1025 4616 1083 4650
rect 1117 4616 1175 4650
rect 1209 4616 1267 4650
rect 1301 4616 1359 4650
rect 1393 4616 1451 4650
rect 1485 4616 1543 4650
rect 1577 4616 1635 4650
rect 1669 4616 1727 4650
rect 1761 4616 1819 4650
rect 1853 4616 1911 4650
rect 1945 4616 2003 4650
rect 2037 4616 2095 4650
rect 2129 4616 2187 4650
rect 2221 4616 2279 4650
rect 2313 4616 2351 4650
rect 2405 4616 2443 4650
rect 2477 4616 2535 4650
rect 2569 4616 2627 4650
rect 2661 4616 2719 4650
rect 2753 4616 2811 4650
rect 2845 4616 2903 4650
rect 2937 4616 2995 4650
rect 3029 4616 3087 4650
rect 3121 4616 3179 4650
rect 3213 4616 3271 4650
rect 3305 4616 3363 4650
rect 3397 4616 3455 4650
rect 3489 4616 3547 4650
rect 3581 4616 3639 4650
rect 3673 4616 3731 4650
rect 3765 4616 3823 4650
rect 3857 4616 3915 4650
rect 3949 4616 4007 4650
rect 4041 4616 4099 4650
rect 4133 4616 4210 4650
rect 4320 4616 4375 4650
rect 4409 4616 4467 4650
rect 4501 4616 4559 4650
rect 4593 4616 4651 4650
rect 4685 4616 4743 4650
rect 4777 4616 4835 4650
rect 4869 4616 4927 4650
rect 4961 4616 5019 4650
rect 5053 4616 5111 4650
rect 5145 4616 5203 4650
rect 5237 4616 5295 4650
rect 5329 4616 5387 4650
rect 5421 4616 5479 4650
rect 5513 4616 5571 4650
rect 5605 4616 5663 4650
rect 5697 4616 5755 4650
rect 5789 4616 5847 4650
rect 5881 4616 5939 4650
rect 5973 4616 6031 4650
rect 6065 4616 6123 4650
rect 6157 4616 6215 4650
rect 6249 4616 6307 4650
rect 6341 4616 6399 4650
rect 6433 4616 6491 4650
rect 6525 4616 6602 4650
rect 6712 4616 6767 4650
rect 6801 4616 6859 4650
rect 6893 4616 6951 4650
rect 6985 4616 7043 4650
rect 7077 4616 7135 4650
rect 7169 4616 7227 4650
rect 7261 4616 7319 4650
rect 7353 4616 7411 4650
rect 7445 4616 7503 4650
rect 7537 4616 7595 4650
rect 7629 4616 7687 4650
rect 7721 4616 7779 4650
rect 7813 4616 7871 4650
rect 7905 4616 7963 4650
rect 7997 4616 8055 4650
rect 8089 4616 8147 4650
rect 8181 4616 8239 4650
rect 8273 4616 8331 4650
rect 8365 4616 8423 4650
rect 8457 4616 8515 4650
rect 8549 4616 8607 4650
rect 8641 4616 8699 4650
rect 8733 4616 8791 4650
rect 8825 4616 8883 4650
rect 8917 4616 8994 4650
rect 9104 4616 9159 4650
rect 9193 4616 9251 4650
rect 9285 4616 9343 4650
rect 9377 4616 9435 4650
rect 9469 4616 9527 4650
rect 9561 4616 9619 4650
rect 9653 4616 9711 4650
rect 9745 4616 9803 4650
rect 9837 4616 9895 4650
rect 9929 4616 9987 4650
rect 10021 4616 10079 4650
rect 10113 4616 10171 4650
rect 10205 4616 10263 4650
rect 10297 4616 10355 4650
rect 10389 4616 10447 4650
rect 10481 4616 10539 4650
rect 10573 4616 10631 4650
rect 10665 4616 10723 4650
rect 10757 4616 10815 4650
rect 10849 4616 10907 4650
rect 10941 4616 10999 4650
rect 11033 4616 11091 4650
rect 11125 4616 11183 4650
rect 11217 4616 11275 4650
rect 11309 4616 11386 4650
rect 11496 4616 11551 4650
rect 11585 4616 11643 4650
rect 11677 4616 11735 4650
rect 11769 4616 11827 4650
rect 11861 4616 11919 4650
rect 11953 4616 12011 4650
rect 12045 4616 12103 4650
rect 12137 4616 12195 4650
rect 12229 4616 12287 4650
rect 12321 4616 12379 4650
rect 12413 4616 12471 4650
rect 12505 4616 12563 4650
rect 12597 4616 12655 4650
rect 12689 4616 12747 4650
rect 12781 4616 12839 4650
rect 12873 4616 12931 4650
rect 12965 4616 12996 4650
rect 3168 3743 3197 3777
rect 3231 3743 3289 3777
rect 3323 3743 3381 3777
rect 3415 3743 3473 3777
rect 3507 3743 3565 3777
rect 3599 3743 3657 3777
rect 3691 3743 3749 3777
rect 3783 3743 3841 3777
rect 3875 3743 3933 3777
rect 3967 3743 4025 3777
rect 4059 3743 4117 3777
rect 4151 3743 4209 3777
rect 4243 3743 4301 3777
rect 4335 3743 4393 3777
rect 4427 3743 4485 3777
rect 4519 3743 4577 3777
rect 4611 3743 4669 3777
rect 4703 3743 4761 3777
rect 4795 3743 4853 3777
rect 4887 3743 4945 3777
rect 4979 3743 5018 3777
rect 5052 3743 5110 3777
rect 5144 3743 5202 3777
rect 5236 3743 5294 3777
rect 5328 3743 5386 3777
rect 5420 3743 5478 3777
rect 5512 3743 5570 3777
rect 5604 3743 5662 3777
rect 5696 3743 5754 3777
rect 5788 3743 5846 3777
rect 5880 3743 5938 3777
rect 5972 3743 6030 3777
rect 6064 3743 6122 3777
rect 6156 3743 6214 3777
rect 6248 3743 6306 3777
rect 6340 3743 6398 3777
rect 6432 3743 6490 3777
rect 6524 3743 6582 3777
rect 6616 3743 6674 3777
rect 6708 3743 6766 3777
rect 6800 3743 6858 3777
rect 6892 3743 6950 3777
rect 6984 3743 7042 3777
rect 7076 3743 7134 3777
rect 7168 3743 7226 3777
rect 7260 3743 7318 3777
rect 7352 3743 7410 3777
rect 7444 3743 7502 3777
rect 7536 3743 7594 3777
rect 7628 3743 7686 3777
rect 7720 3743 7778 3777
rect 7812 3743 7870 3777
rect 7904 3743 7962 3777
rect 7996 3743 8054 3777
rect 8088 3743 8146 3777
rect 8180 3743 8238 3777
rect 8272 3743 8330 3777
rect 8364 3743 8422 3777
rect 8456 3743 8514 3777
rect 8548 3743 8606 3777
rect 8640 3743 8698 3777
rect 8732 3743 8790 3777
rect 8824 3743 8882 3777
rect 8916 3743 8974 3777
rect 9008 3743 9066 3777
rect 9100 3743 9158 3777
rect 9192 3743 9250 3777
rect 9284 3743 9342 3777
rect 9376 3743 9434 3777
rect 9468 3743 9526 3777
rect 9560 3743 9618 3777
rect 9652 3743 9710 3777
rect 9744 3743 9802 3777
rect 9836 3743 9894 3777
rect 9928 3743 9986 3777
rect 10020 3743 10078 3777
rect 10112 3743 10170 3777
rect 10204 3743 10262 3777
rect 10296 3743 10354 3777
rect 10388 3743 10446 3777
rect 10480 3743 10538 3777
rect 10572 3743 10630 3777
rect 10664 3743 10722 3777
rect 10756 3743 10814 3777
rect 10848 3743 10906 3777
rect 10940 3743 10998 3777
rect 11032 3743 11090 3777
rect 11124 3743 11182 3777
rect 11216 3743 11274 3777
rect 11308 3743 11366 3777
rect 11400 3743 11458 3777
rect 11492 3743 11550 3777
rect 11584 3743 11642 3777
rect 11676 3743 11734 3777
rect 11768 3743 11826 3777
rect 11860 3743 11918 3777
rect 11952 3743 12010 3777
rect 12044 3743 12102 3777
rect 12136 3743 12194 3777
rect 12228 3743 12286 3777
rect 12320 3743 12378 3777
rect 12412 3743 12470 3777
rect 12504 3743 12562 3777
rect 12596 3743 12654 3777
rect 12688 3743 12746 3777
rect 12780 3743 12838 3777
rect 12872 3743 12930 3777
rect 12964 3743 12993 3777
rect 1033 2870 1062 2904
rect 1096 2870 1154 2904
rect 1188 2870 1246 2904
rect 1280 2870 1338 2904
rect 1372 2870 1430 2904
rect 1464 2870 1522 2904
rect 1556 2870 1614 2904
rect 1648 2870 1706 2904
rect 1740 2870 1798 2904
rect 1832 2870 1890 2904
rect 1924 2870 1982 2904
rect 2016 2870 2074 2904
rect 2108 2870 2166 2904
rect 2200 2870 2258 2904
rect 2292 2870 2350 2904
rect 2384 2870 2442 2904
rect 2476 2870 2534 2904
rect 2568 2870 2626 2904
rect 2660 2870 2718 2904
rect 2752 2870 2810 2904
rect 2844 2870 2902 2904
rect 2936 2870 2994 2904
rect 3028 2870 3086 2904
rect 3120 2870 3178 2904
rect 3212 2870 3270 2904
rect 3304 2870 3362 2904
rect 3396 2870 3454 2904
rect 3488 2870 3546 2904
rect 3580 2870 3638 2904
rect 3672 2870 3730 2904
rect 3764 2870 3822 2904
rect 3856 2870 3914 2904
rect 3948 2870 4006 2904
rect 4040 2870 4098 2904
rect 4132 2870 4190 2904
rect 4224 2870 4282 2904
rect 4316 2870 4374 2904
rect 4408 2870 4466 2904
rect 4500 2870 4558 2904
rect 4592 2870 4650 2904
rect 4684 2870 4742 2904
rect 4776 2870 4834 2904
rect 4868 2870 4926 2904
rect 4960 2870 5018 2904
rect 5052 2870 5110 2904
rect 5144 2870 5202 2904
rect 5236 2870 5294 2904
rect 5328 2870 5386 2904
rect 5420 2870 5478 2904
rect 5512 2870 5570 2904
rect 5604 2870 5662 2904
rect 5696 2870 5754 2904
rect 5788 2870 5846 2904
rect 5880 2870 5938 2904
rect 5972 2870 6030 2904
rect 6064 2870 6122 2904
rect 6156 2870 6214 2904
rect 6248 2870 6306 2904
rect 6340 2870 6398 2904
rect 6432 2870 6490 2904
rect 6524 2870 6582 2904
rect 6616 2870 6674 2904
rect 6708 2870 6766 2904
rect 6800 2870 6858 2904
rect 6892 2870 6950 2904
rect 6984 2870 7042 2904
rect 7076 2870 7134 2904
rect 7168 2870 7226 2904
rect 7260 2870 7318 2904
rect 7352 2870 7410 2904
rect 7444 2870 7502 2904
rect 7536 2870 7594 2904
rect 7628 2870 7686 2904
rect 7720 2870 7778 2904
rect 7812 2870 7870 2904
rect 7904 2870 7962 2904
rect 7996 2870 8054 2904
rect 8088 2870 8146 2904
rect 8180 2870 8238 2904
rect 8272 2870 8330 2904
rect 8364 2870 8422 2904
rect 8456 2870 8514 2904
rect 8548 2870 8606 2904
rect 8640 2870 8698 2904
rect 8732 2870 8790 2904
rect 8824 2870 8882 2904
rect 8916 2870 8974 2904
rect 9008 2870 9066 2904
rect 9100 2870 9158 2904
rect 9192 2870 9250 2904
rect 9284 2870 9342 2904
rect 9376 2870 9434 2904
rect 9468 2870 9526 2904
rect 9560 2870 9618 2904
rect 9652 2870 9710 2904
rect 9744 2870 9802 2904
rect 9836 2870 9894 2904
rect 9928 2870 9986 2904
rect 10020 2870 10078 2904
rect 10112 2870 10170 2904
rect 10204 2870 10262 2904
rect 10296 2870 10354 2904
rect 10388 2870 10446 2904
rect 10480 2870 10538 2904
rect 10572 2870 10630 2904
rect 10664 2870 10722 2904
rect 10756 2870 10814 2904
rect 10848 2870 10906 2904
rect 10940 2870 10998 2904
rect 11032 2870 11090 2904
rect 11124 2870 11182 2904
rect 11216 2870 11274 2904
rect 11308 2870 11366 2904
rect 11400 2870 11458 2904
rect 11492 2870 11550 2904
rect 11584 2870 11642 2904
rect 11676 2870 11734 2904
rect 11768 2870 11826 2904
rect 11860 2870 11918 2904
rect 11952 2870 12010 2904
rect 12044 2870 12102 2904
rect 12136 2870 12194 2904
rect 12228 2870 12286 2904
rect 12320 2870 12378 2904
rect 12412 2870 12470 2904
rect 12504 2870 12562 2904
rect 12596 2870 12654 2904
rect 12688 2870 12746 2904
rect 12780 2870 12838 2904
rect 12872 2870 12930 2904
rect 12964 2870 12993 2904
<< psubdiffcont >>
rect 1064 5586 1098 5620
rect 1156 5586 1190 5620
rect 1248 5586 1282 5620
rect 1340 5586 1374 5620
rect 1432 5586 1466 5620
rect 1524 5586 1558 5620
rect 1616 5586 1650 5620
rect 1708 5586 1742 5620
rect 1800 5586 1834 5620
rect 1892 5586 1926 5620
rect 1984 5586 2018 5620
rect 2076 5586 2110 5620
rect 2168 5586 2202 5620
rect 2260 5586 2294 5620
rect 2352 5586 2386 5620
rect 2444 5586 2478 5620
rect 2536 5586 2570 5620
rect 2628 5586 2662 5620
rect 2720 5586 2754 5620
rect 2812 5586 2846 5620
rect 2904 5586 2938 5620
rect 2996 5586 3030 5620
rect 3088 5586 3122 5620
rect 3180 5586 3214 5620
rect 3272 5586 3306 5620
rect 3364 5586 3398 5620
rect 3456 5586 3490 5620
rect 3548 5586 3582 5620
rect 3640 5586 3674 5620
rect 3732 5586 3766 5620
rect 3824 5586 3858 5620
rect 3916 5586 3950 5620
rect 4008 5586 4042 5620
rect 1063 4713 1097 4747
rect 1155 4713 1189 4747
rect 1247 4713 1281 4747
rect 1339 4713 1373 4747
rect 1431 4713 1465 4747
rect 1523 4713 1557 4747
rect 1615 4713 1649 4747
rect 1707 4713 1741 4747
rect 1799 4713 1833 4747
rect 1891 4713 1925 4747
rect 1983 4713 2017 4747
rect 2075 4713 2109 4747
rect 2167 4713 2201 4747
rect 2259 4713 2293 4747
rect 2351 4713 2385 4747
rect 2443 4713 2477 4747
rect 2535 4713 2569 4747
rect 2627 4713 2661 4747
rect 2719 4713 2753 4747
rect 2811 4713 2845 4747
rect 2903 4713 2937 4747
rect 2995 4713 3029 4747
rect 3087 4713 3121 4747
rect 3179 4713 3213 4747
rect 3271 4713 3305 4747
rect 3363 4713 3397 4747
rect 3455 4713 3489 4747
rect 3547 4713 3581 4747
rect 3639 4713 3673 4747
rect 3731 4713 3765 4747
rect 3823 4713 3857 4747
rect 3915 4713 3949 4747
rect 4007 4713 4041 4747
rect 4099 4713 4133 4747
rect 4191 4713 4225 4747
rect 4283 4713 4317 4747
rect 4375 4713 4409 4747
rect 4467 4713 4501 4747
rect 4559 4713 4593 4747
rect 4651 4713 4685 4747
rect 4743 4713 4777 4747
rect 4835 4713 4869 4747
rect 4927 4713 4961 4747
rect 5019 4713 5053 4747
rect 5111 4713 5145 4747
rect 5203 4713 5237 4747
rect 5295 4713 5329 4747
rect 5387 4713 5421 4747
rect 5479 4713 5513 4747
rect 5571 4713 5605 4747
rect 5663 4713 5697 4747
rect 5755 4713 5789 4747
rect 5847 4713 5881 4747
rect 5939 4713 5973 4747
rect 6031 4713 6065 4747
rect 6123 4713 6157 4747
rect 6215 4713 6249 4747
rect 6307 4713 6341 4747
rect 6399 4713 6433 4747
rect 6491 4713 6525 4747
rect 6583 4713 6617 4747
rect 6675 4713 6709 4747
rect 6767 4713 6801 4747
rect 6859 4713 6893 4747
rect 6951 4713 6985 4747
rect 7043 4713 7077 4747
rect 7135 4713 7169 4747
rect 7227 4713 7261 4747
rect 7319 4713 7353 4747
rect 7411 4713 7445 4747
rect 7503 4713 7537 4747
rect 7595 4713 7629 4747
rect 7687 4713 7721 4747
rect 7779 4713 7813 4747
rect 7871 4713 7905 4747
rect 7963 4713 7997 4747
rect 8055 4713 8089 4747
rect 8147 4713 8181 4747
rect 8239 4713 8273 4747
rect 8331 4713 8365 4747
rect 8423 4713 8457 4747
rect 8515 4713 8549 4747
rect 8607 4713 8641 4747
rect 8699 4713 8733 4747
rect 8791 4713 8825 4747
rect 8883 4713 8917 4747
rect 8975 4713 9009 4747
rect 9067 4713 9101 4747
rect 9159 4713 9193 4747
rect 9251 4713 9285 4747
rect 9343 4713 9377 4747
rect 9435 4713 9469 4747
rect 9527 4713 9561 4747
rect 9619 4713 9653 4747
rect 9711 4713 9745 4747
rect 9803 4713 9837 4747
rect 9895 4713 9929 4747
rect 9987 4713 10021 4747
rect 10079 4713 10113 4747
rect 10171 4713 10205 4747
rect 10263 4713 10297 4747
rect 10355 4713 10389 4747
rect 10447 4713 10481 4747
rect 10539 4713 10573 4747
rect 10631 4713 10665 4747
rect 10723 4713 10757 4747
rect 10815 4713 10849 4747
rect 10907 4713 10941 4747
rect 10999 4713 11033 4747
rect 11091 4713 11125 4747
rect 11183 4713 11217 4747
rect 11275 4713 11309 4747
rect 11367 4713 11401 4747
rect 11459 4713 11493 4747
rect 11551 4713 11585 4747
rect 11643 4713 11677 4747
rect 11735 4713 11769 4747
rect 11827 4713 11861 4747
rect 11919 4713 11953 4747
rect 12011 4713 12045 4747
rect 12103 4713 12137 4747
rect 12195 4713 12229 4747
rect 12287 4713 12321 4747
rect 12379 4713 12413 4747
rect 12471 4713 12505 4747
rect 12563 4713 12597 4747
rect 12655 4713 12689 4747
rect 12747 4713 12781 4747
rect 12839 4713 12873 4747
rect 12931 4713 12965 4747
rect 623 4024 657 4058
rect 715 4024 749 4058
rect 807 4024 841 4058
rect 899 4024 933 4058
rect 991 4024 1025 4058
rect 1083 4024 1117 4058
rect 1175 4024 1209 4058
rect 1267 4024 1301 4058
rect 1359 4024 1393 4058
rect 1451 4024 1485 4058
rect 1543 4024 1577 4058
rect 1635 4024 1669 4058
rect 1727 4024 1761 4058
rect 1819 4024 1853 4058
rect 1911 4024 1945 4058
rect 2003 4024 2037 4058
rect 2095 4024 2129 4058
rect 2187 4024 2221 4058
rect 2279 4024 2313 4058
rect 2371 4024 2405 4058
rect 2463 4024 2497 4058
rect 2555 4024 2589 4058
rect 2647 4024 2681 4058
rect 2739 4024 2773 4058
rect 2831 4024 2865 4058
rect 2923 4024 2957 4058
rect 3015 4024 3049 4058
rect 3107 4024 3141 4058
rect 3199 4024 3233 4058
rect 3291 4024 3325 4058
rect 3383 4024 3417 4058
rect 3475 4024 3509 4058
rect 3567 4024 3601 4058
rect 3659 4024 3693 4058
rect 3751 4024 3785 4058
rect 3843 4024 3877 4058
rect 3935 4024 3969 4058
rect 4027 4024 4061 4058
rect 4119 4024 4153 4058
rect 4211 4024 4245 4058
rect 4303 4024 4337 4058
rect 4395 4024 4429 4058
rect 4487 4024 4521 4058
rect 4579 4024 4613 4058
rect 4671 4024 4705 4058
rect 4763 4024 4797 4058
rect 4855 4024 4889 4058
rect 4947 4024 4981 4058
rect 5039 4024 5073 4058
rect 5131 4024 5165 4058
rect 5223 4024 5257 4058
rect 5315 4024 5349 4058
rect 5407 4024 5441 4058
rect 5499 4024 5533 4058
rect 5591 4024 5625 4058
rect 5683 4024 5717 4058
rect 5775 4024 5809 4058
rect 5867 4024 5901 4058
rect 5959 4024 5993 4058
rect 6051 4024 6085 4058
rect 6143 4024 6177 4058
rect 6235 4024 6269 4058
rect 6327 4024 6361 4058
rect 6419 4024 6453 4058
rect 6511 4024 6545 4058
rect 6603 4024 6637 4058
rect 6695 4024 6729 4058
rect 6787 4024 6821 4058
rect 6879 4024 6913 4058
rect 6971 4024 7005 4058
rect 7063 4024 7097 4058
rect 7155 4024 7189 4058
rect 7247 4024 7281 4058
rect 7339 4024 7373 4058
rect 7431 4024 7465 4058
rect 7523 4024 7557 4058
rect 7615 4024 7649 4058
rect 7707 4024 7741 4058
rect 7799 4024 7833 4058
rect 7891 4024 7925 4058
rect 7983 4024 8017 4058
rect 8075 4024 8109 4058
rect 8167 4024 8201 4058
rect 8259 4024 8293 4058
rect 8351 4024 8385 4058
rect 8443 4024 8477 4058
rect 8535 4024 8569 4058
rect 8627 4024 8661 4058
rect 8719 4024 8753 4058
rect 8811 4024 8845 4058
rect 8903 4024 8937 4058
rect 8995 4024 9029 4058
rect 9087 4024 9121 4058
rect 9179 4024 9213 4058
rect 9271 4024 9305 4058
rect 9363 4024 9397 4058
rect 9435 4024 9469 4058
rect 9527 4024 9561 4058
rect 9619 4024 9653 4058
rect 9711 4024 9745 4058
rect 9803 4024 9837 4058
rect 9895 4024 9929 4058
rect 9987 4024 10021 4058
rect 10079 4024 10113 4058
rect 10171 4024 10205 4058
rect 10263 4024 10297 4058
rect 10355 4024 10389 4058
rect 10447 4024 10481 4058
rect 10539 4024 10573 4058
rect 10631 4024 10665 4058
rect 10723 4024 10757 4058
rect 10815 4024 10849 4058
rect 10907 4024 10941 4058
rect 10999 4024 11033 4058
rect 11091 4024 11125 4058
rect 11183 4024 11217 4058
rect 11275 4024 11309 4058
rect 11367 4024 11401 4058
rect 11459 4024 11493 4058
rect 11551 4024 11585 4058
rect 11643 4024 11677 4058
rect 11735 4024 11769 4058
rect 11827 4024 11861 4058
rect 11919 4024 11953 4058
rect 12011 4024 12045 4058
rect 12103 4024 12137 4058
rect 12195 4024 12229 4058
rect 12287 4024 12321 4058
rect 12379 4024 12413 4058
rect 12471 4024 12505 4058
rect 12563 4024 12597 4058
rect 12655 4024 12689 4058
rect 12747 4024 12781 4058
rect 12839 4024 12873 4058
rect 12931 4024 12965 4058
rect 3197 3151 3231 3185
rect 3289 3151 3323 3185
rect 3381 3151 3415 3185
rect 3473 3151 3507 3185
rect 3565 3151 3599 3185
rect 3657 3151 3691 3185
rect 3749 3151 3783 3185
rect 3841 3151 3875 3185
rect 3933 3151 3967 3185
rect 4025 3151 4059 3185
rect 4117 3151 4151 3185
rect 4209 3151 4243 3185
rect 4301 3151 4335 3185
rect 4393 3151 4427 3185
rect 4485 3151 4519 3185
rect 4577 3151 4611 3185
rect 4669 3151 4703 3185
rect 4761 3151 4795 3185
rect 4853 3151 4887 3185
rect 4945 3151 4979 3185
rect 5037 3151 5071 3185
rect 5129 3151 5163 3185
rect 5221 3151 5255 3185
rect 5313 3151 5347 3185
rect 5405 3151 5439 3185
rect 5497 3151 5531 3185
rect 5589 3151 5623 3185
rect 5681 3151 5715 3185
rect 5773 3151 5807 3185
rect 5865 3151 5899 3185
rect 5957 3151 5991 3185
rect 6049 3151 6083 3185
rect 6141 3151 6175 3185
rect 6233 3151 6267 3185
rect 6325 3151 6359 3185
rect 6417 3151 6451 3185
rect 6509 3151 6543 3185
rect 6601 3151 6635 3185
rect 6693 3151 6727 3185
rect 6785 3151 6819 3185
rect 6877 3151 6911 3185
rect 6969 3151 7003 3185
rect 7061 3151 7095 3185
rect 7153 3151 7187 3185
rect 7245 3151 7279 3185
rect 7337 3151 7371 3185
rect 7429 3151 7463 3185
rect 7521 3151 7555 3185
rect 7613 3151 7647 3185
rect 7705 3151 7739 3185
rect 7797 3151 7831 3185
rect 7889 3151 7923 3185
rect 7981 3151 8015 3185
rect 8073 3151 8107 3185
rect 8165 3151 8199 3185
rect 8257 3151 8291 3185
rect 8349 3151 8383 3185
rect 8441 3151 8475 3185
rect 8533 3151 8567 3185
rect 8625 3151 8659 3185
rect 8717 3151 8751 3185
rect 8809 3151 8843 3185
rect 8901 3151 8935 3185
rect 8993 3151 9027 3185
rect 9085 3151 9119 3185
rect 9177 3151 9211 3185
rect 9269 3151 9303 3185
rect 9361 3151 9395 3185
rect 9453 3151 9487 3185
rect 9545 3151 9579 3185
rect 9637 3151 9671 3185
rect 9729 3151 9763 3185
rect 9821 3151 9855 3185
rect 9894 3151 9947 3185
rect 9986 3151 10039 3185
rect 10078 3151 10131 3185
rect 10170 3151 10223 3185
rect 10262 3151 10315 3185
rect 10354 3151 10407 3185
rect 10446 3151 10499 3185
rect 10538 3151 10591 3185
rect 10630 3151 10683 3185
rect 10722 3151 10775 3185
rect 10814 3151 10867 3185
rect 10906 3151 10959 3185
rect 10998 3151 11051 3185
rect 11090 3151 11143 3185
rect 11182 3151 11235 3185
rect 11274 3151 11327 3185
rect 11366 3151 11419 3185
rect 11458 3151 11511 3185
rect 11550 3151 11603 3185
rect 11642 3151 11695 3185
rect 11734 3151 11787 3185
rect 11826 3151 11879 3185
rect 11918 3151 11971 3185
rect 12010 3151 12044 3185
rect 12102 3151 12136 3185
rect 12194 3151 12228 3185
rect 12286 3151 12320 3185
rect 12378 3151 12412 3185
rect 12470 3151 12504 3185
rect 12562 3151 12596 3185
rect 12654 3151 12688 3185
rect 12746 3151 12780 3185
rect 12838 3151 12872 3185
rect 12930 3151 12964 3185
rect 1062 2278 1096 2312
rect 1154 2278 1188 2312
rect 1246 2278 1280 2312
rect 1338 2278 1372 2312
rect 1430 2278 1464 2312
rect 1522 2278 1556 2312
rect 1614 2278 1648 2312
rect 1706 2278 1740 2312
rect 1798 2278 1832 2312
rect 1890 2278 1924 2312
rect 1982 2278 2016 2312
rect 2074 2278 2108 2312
rect 2166 2278 2200 2312
rect 2258 2278 2292 2312
rect 2350 2278 2384 2312
rect 2442 2278 2476 2312
rect 2534 2278 2568 2312
rect 2626 2278 2660 2312
rect 2718 2278 2752 2312
rect 2810 2278 2844 2312
rect 2902 2278 2936 2312
rect 2994 2278 3028 2312
rect 3086 2278 3120 2312
rect 3178 2278 3212 2312
rect 3270 2278 3304 2312
rect 3362 2278 3396 2312
rect 3454 2278 3488 2312
rect 3546 2278 3580 2312
rect 3638 2278 3672 2312
rect 3730 2278 3764 2312
rect 3822 2278 3856 2312
rect 3914 2278 3948 2312
rect 4006 2278 4040 2312
rect 4098 2278 4132 2312
rect 4190 2278 4224 2312
rect 4282 2278 4316 2312
rect 4374 2278 4408 2312
rect 4466 2278 4500 2312
rect 4558 2278 4592 2312
rect 4650 2278 4684 2312
rect 4742 2278 4776 2312
rect 4834 2278 4868 2312
rect 4926 2278 4960 2312
rect 5018 2278 5052 2312
rect 5110 2278 5144 2312
rect 5202 2278 5236 2312
rect 5294 2278 5328 2312
rect 5386 2278 5420 2312
rect 5478 2278 5512 2312
rect 5570 2278 5604 2312
rect 5662 2278 5696 2312
rect 5754 2278 5788 2312
rect 5846 2278 5880 2312
rect 5938 2278 5972 2312
rect 6030 2278 6064 2312
rect 6122 2278 6156 2312
rect 6214 2278 6248 2312
rect 6306 2278 6340 2312
rect 6398 2278 6432 2312
rect 6490 2278 6524 2312
rect 6582 2278 6616 2312
rect 6674 2278 6708 2312
rect 6766 2278 6800 2312
rect 6858 2278 6892 2312
rect 6950 2278 6984 2312
rect 7042 2278 7076 2312
rect 7134 2278 7168 2312
rect 7226 2278 7260 2312
rect 7318 2278 7352 2312
rect 7410 2278 7444 2312
rect 7502 2278 7536 2312
rect 7594 2278 7628 2312
rect 7686 2278 7720 2312
rect 7778 2278 7812 2312
rect 7870 2278 7904 2312
rect 7962 2278 7996 2312
rect 8054 2278 8088 2312
rect 8146 2278 8180 2312
rect 8238 2278 8272 2312
rect 8330 2278 8364 2312
rect 8422 2278 8456 2312
rect 8514 2278 8548 2312
rect 8606 2278 8640 2312
rect 8698 2278 8732 2312
rect 8790 2278 8824 2312
rect 8882 2278 8916 2312
rect 8974 2278 9008 2312
rect 9066 2278 9100 2312
rect 9158 2278 9192 2312
rect 9250 2278 9284 2312
rect 9342 2278 9376 2312
rect 9434 2278 9468 2312
rect 9526 2278 9560 2312
rect 9618 2278 9652 2312
rect 9710 2278 9744 2312
rect 9802 2278 9836 2312
rect 9894 2278 9928 2312
rect 9986 2278 10020 2312
rect 10078 2278 10112 2312
rect 10170 2278 10204 2312
rect 10262 2278 10296 2312
rect 10354 2278 10388 2312
rect 10446 2278 10480 2312
rect 10538 2278 10572 2312
rect 10630 2278 10664 2312
rect 10722 2278 10756 2312
rect 10814 2278 10848 2312
rect 10906 2278 10940 2312
rect 10998 2278 11032 2312
rect 11090 2278 11124 2312
rect 11182 2278 11216 2312
rect 11274 2278 11308 2312
rect 11366 2278 11400 2312
rect 11458 2278 11492 2312
rect 11550 2278 11584 2312
rect 11642 2278 11676 2312
rect 11734 2278 11768 2312
rect 11826 2278 11860 2312
rect 11918 2278 11952 2312
rect 12010 2278 12044 2312
rect 12102 2278 12136 2312
rect 12194 2278 12228 2312
rect 12286 2278 12320 2312
rect 12378 2278 12412 2312
rect 12470 2278 12504 2312
rect 12562 2278 12596 2312
rect 12654 2278 12688 2312
rect 12746 2278 12780 2312
rect 12838 2278 12872 2312
rect 12930 2278 12964 2312
<< nsubdiffcont >>
rect 1064 6178 1098 6212
rect 1156 6178 1190 6212
rect 1248 6178 1282 6212
rect 1340 6178 1374 6212
rect 1432 6178 1466 6212
rect 1524 6178 1558 6212
rect 1616 6178 1650 6212
rect 2324 6178 2358 6212
rect 2416 6178 2450 6212
rect 2508 6178 2542 6212
rect 2600 6178 2634 6212
rect 2692 6178 2726 6212
rect 2784 6178 2818 6212
rect 2876 6178 2910 6212
rect 2968 6178 3002 6212
rect 3060 6178 3094 6212
rect 3152 6178 3186 6212
rect 3244 6178 3278 6212
rect 3336 6178 3370 6212
rect 3428 6178 3462 6212
rect 3520 6178 3554 6212
rect 3612 6178 3646 6212
rect 3704 6178 3738 6212
rect 3796 6178 3830 6212
rect 3888 6178 3922 6212
rect 3980 6178 4014 6212
rect 4072 6178 4106 6212
rect 1063 5305 1097 5339
rect 1155 5305 1189 5339
rect 1247 5305 1281 5339
rect 1339 5305 1373 5339
rect 1431 5305 1465 5339
rect 1523 5305 1557 5339
rect 1615 5305 1649 5339
rect 1707 5305 1741 5339
rect 1799 5305 1833 5339
rect 1891 5305 1925 5339
rect 1983 5305 2017 5339
rect 2075 5305 2109 5339
rect 2167 5305 2201 5339
rect 2259 5305 2293 5339
rect 2351 5305 2385 5339
rect 2443 5305 2477 5339
rect 2535 5305 2569 5339
rect 2627 5305 2661 5339
rect 2719 5305 2753 5339
rect 2811 5305 2845 5339
rect 3087 5305 3121 5339
rect 3179 5305 3213 5339
rect 3271 5305 3305 5339
rect 3363 5305 3397 5339
rect 3455 5305 3489 5339
rect 3547 5305 3581 5339
rect 3640 5305 3674 5339
rect 3731 5305 3765 5339
rect 3823 5305 3857 5339
rect 3915 5305 3949 5339
rect 4007 5305 4041 5339
rect 4283 5305 4317 5339
rect 4375 5305 4409 5339
rect 4467 5305 4501 5339
rect 4559 5305 4593 5339
rect 4651 5305 4685 5339
rect 4743 5305 4777 5339
rect 4835 5305 4869 5339
rect 4927 5305 4961 5339
rect 5019 5305 5053 5339
rect 5111 5305 5145 5339
rect 5203 5305 5237 5339
rect 5295 5305 5329 5339
rect 5387 5305 5421 5339
rect 5479 5305 5513 5339
rect 5571 5305 5605 5339
rect 5663 5305 5697 5339
rect 5755 5305 5789 5339
rect 5847 5305 5881 5339
rect 5939 5305 5973 5339
rect 6031 5305 6065 5339
rect 6123 5305 6157 5339
rect 6215 5305 6249 5339
rect 6307 5305 6341 5339
rect 6399 5305 6433 5339
rect 6675 5305 6709 5339
rect 6767 5305 6801 5339
rect 6859 5305 6893 5339
rect 6951 5305 6985 5339
rect 7043 5305 7077 5339
rect 7135 5305 7169 5339
rect 7227 5305 7261 5339
rect 7319 5305 7353 5339
rect 7411 5305 7445 5339
rect 7503 5305 7537 5339
rect 7595 5305 7629 5339
rect 7687 5305 7721 5339
rect 7779 5305 7813 5339
rect 7871 5305 7905 5339
rect 7963 5305 7997 5339
rect 8055 5305 8089 5339
rect 8147 5305 8181 5339
rect 8239 5305 8273 5339
rect 8331 5305 8365 5339
rect 8423 5305 8457 5339
rect 8515 5305 8549 5339
rect 8607 5305 8641 5339
rect 8699 5305 8733 5339
rect 8791 5305 8825 5339
rect 9067 5305 9101 5339
rect 9159 5305 9193 5339
rect 9251 5305 9285 5339
rect 9343 5305 9377 5339
rect 9435 5305 9469 5339
rect 9527 5305 9561 5339
rect 9619 5305 9653 5339
rect 9711 5305 9745 5339
rect 9803 5305 9837 5339
rect 9895 5305 9929 5339
rect 9987 5305 10021 5339
rect 10079 5305 10113 5339
rect 10171 5305 10205 5339
rect 10263 5305 10297 5339
rect 10355 5305 10389 5339
rect 10447 5305 10481 5339
rect 10539 5305 10573 5339
rect 10631 5305 10665 5339
rect 10723 5305 10757 5339
rect 10815 5305 10849 5339
rect 10907 5305 10941 5339
rect 10999 5305 11033 5339
rect 11091 5305 11125 5339
rect 11183 5305 11217 5339
rect 11459 5305 11493 5339
rect 11551 5305 11585 5339
rect 11643 5305 11677 5339
rect 11735 5305 11769 5339
rect 11827 5305 11861 5339
rect 11919 5305 11953 5339
rect 12011 5305 12045 5339
rect 12103 5305 12137 5339
rect 12195 5305 12229 5339
rect 12287 5305 12321 5339
rect 12379 5305 12413 5339
rect 12471 5305 12505 5339
rect 12563 5305 12597 5339
rect 12655 5305 12689 5339
rect 12747 5305 12781 5339
rect 12839 5305 12873 5339
rect 12931 5305 12965 5339
rect 623 4616 657 4650
rect 715 4616 749 4650
rect 807 4616 841 4650
rect 899 4616 933 4650
rect 991 4616 1025 4650
rect 1083 4616 1117 4650
rect 1175 4616 1209 4650
rect 1267 4616 1301 4650
rect 1359 4616 1393 4650
rect 1451 4616 1485 4650
rect 1543 4616 1577 4650
rect 1635 4616 1669 4650
rect 1727 4616 1761 4650
rect 1819 4616 1853 4650
rect 1911 4616 1945 4650
rect 2003 4616 2037 4650
rect 2095 4616 2129 4650
rect 2187 4616 2221 4650
rect 2279 4616 2313 4650
rect 2351 4616 2405 4650
rect 2443 4616 2477 4650
rect 2535 4616 2569 4650
rect 2627 4616 2661 4650
rect 2719 4616 2753 4650
rect 2811 4616 2845 4650
rect 2903 4616 2937 4650
rect 2995 4616 3029 4650
rect 3087 4616 3121 4650
rect 3179 4616 3213 4650
rect 3271 4616 3305 4650
rect 3363 4616 3397 4650
rect 3455 4616 3489 4650
rect 3547 4616 3581 4650
rect 3639 4616 3673 4650
rect 3731 4616 3765 4650
rect 3823 4616 3857 4650
rect 3915 4616 3949 4650
rect 4007 4616 4041 4650
rect 4099 4616 4133 4650
rect 4375 4616 4409 4650
rect 4467 4616 4501 4650
rect 4559 4616 4593 4650
rect 4651 4616 4685 4650
rect 4743 4616 4777 4650
rect 4835 4616 4869 4650
rect 4927 4616 4961 4650
rect 5019 4616 5053 4650
rect 5111 4616 5145 4650
rect 5203 4616 5237 4650
rect 5295 4616 5329 4650
rect 5387 4616 5421 4650
rect 5479 4616 5513 4650
rect 5571 4616 5605 4650
rect 5663 4616 5697 4650
rect 5755 4616 5789 4650
rect 5847 4616 5881 4650
rect 5939 4616 5973 4650
rect 6031 4616 6065 4650
rect 6123 4616 6157 4650
rect 6215 4616 6249 4650
rect 6307 4616 6341 4650
rect 6399 4616 6433 4650
rect 6491 4616 6525 4650
rect 6767 4616 6801 4650
rect 6859 4616 6893 4650
rect 6951 4616 6985 4650
rect 7043 4616 7077 4650
rect 7135 4616 7169 4650
rect 7227 4616 7261 4650
rect 7319 4616 7353 4650
rect 7411 4616 7445 4650
rect 7503 4616 7537 4650
rect 7595 4616 7629 4650
rect 7687 4616 7721 4650
rect 7779 4616 7813 4650
rect 7871 4616 7905 4650
rect 7963 4616 7997 4650
rect 8055 4616 8089 4650
rect 8147 4616 8181 4650
rect 8239 4616 8273 4650
rect 8331 4616 8365 4650
rect 8423 4616 8457 4650
rect 8515 4616 8549 4650
rect 8607 4616 8641 4650
rect 8699 4616 8733 4650
rect 8791 4616 8825 4650
rect 8883 4616 8917 4650
rect 9159 4616 9193 4650
rect 9251 4616 9285 4650
rect 9343 4616 9377 4650
rect 9435 4616 9469 4650
rect 9527 4616 9561 4650
rect 9619 4616 9653 4650
rect 9711 4616 9745 4650
rect 9803 4616 9837 4650
rect 9895 4616 9929 4650
rect 9987 4616 10021 4650
rect 10079 4616 10113 4650
rect 10171 4616 10205 4650
rect 10263 4616 10297 4650
rect 10355 4616 10389 4650
rect 10447 4616 10481 4650
rect 10539 4616 10573 4650
rect 10631 4616 10665 4650
rect 10723 4616 10757 4650
rect 10815 4616 10849 4650
rect 10907 4616 10941 4650
rect 10999 4616 11033 4650
rect 11091 4616 11125 4650
rect 11183 4616 11217 4650
rect 11275 4616 11309 4650
rect 11551 4616 11585 4650
rect 11643 4616 11677 4650
rect 11735 4616 11769 4650
rect 11827 4616 11861 4650
rect 11919 4616 11953 4650
rect 12011 4616 12045 4650
rect 12103 4616 12137 4650
rect 12195 4616 12229 4650
rect 12287 4616 12321 4650
rect 12379 4616 12413 4650
rect 12471 4616 12505 4650
rect 12563 4616 12597 4650
rect 12655 4616 12689 4650
rect 12747 4616 12781 4650
rect 12839 4616 12873 4650
rect 12931 4616 12965 4650
rect 3197 3743 3231 3777
rect 3289 3743 3323 3777
rect 3381 3743 3415 3777
rect 3473 3743 3507 3777
rect 3565 3743 3599 3777
rect 3657 3743 3691 3777
rect 3749 3743 3783 3777
rect 3841 3743 3875 3777
rect 3933 3743 3967 3777
rect 4025 3743 4059 3777
rect 4117 3743 4151 3777
rect 4209 3743 4243 3777
rect 4301 3743 4335 3777
rect 4393 3743 4427 3777
rect 4485 3743 4519 3777
rect 4577 3743 4611 3777
rect 4669 3743 4703 3777
rect 4761 3743 4795 3777
rect 4853 3743 4887 3777
rect 4945 3743 4979 3777
rect 5018 3743 5052 3777
rect 5110 3743 5144 3777
rect 5202 3743 5236 3777
rect 5294 3743 5328 3777
rect 5386 3743 5420 3777
rect 5478 3743 5512 3777
rect 5570 3743 5604 3777
rect 5662 3743 5696 3777
rect 5754 3743 5788 3777
rect 5846 3743 5880 3777
rect 5938 3743 5972 3777
rect 6030 3743 6064 3777
rect 6122 3743 6156 3777
rect 6214 3743 6248 3777
rect 6306 3743 6340 3777
rect 6398 3743 6432 3777
rect 6490 3743 6524 3777
rect 6582 3743 6616 3777
rect 6674 3743 6708 3777
rect 6766 3743 6800 3777
rect 6858 3743 6892 3777
rect 6950 3743 6984 3777
rect 7042 3743 7076 3777
rect 7134 3743 7168 3777
rect 7226 3743 7260 3777
rect 7318 3743 7352 3777
rect 7410 3743 7444 3777
rect 7502 3743 7536 3777
rect 7594 3743 7628 3777
rect 7686 3743 7720 3777
rect 7778 3743 7812 3777
rect 7870 3743 7904 3777
rect 7962 3743 7996 3777
rect 8054 3743 8088 3777
rect 8146 3743 8180 3777
rect 8238 3743 8272 3777
rect 8330 3743 8364 3777
rect 8422 3743 8456 3777
rect 8514 3743 8548 3777
rect 8606 3743 8640 3777
rect 8698 3743 8732 3777
rect 8790 3743 8824 3777
rect 8882 3743 8916 3777
rect 8974 3743 9008 3777
rect 9066 3743 9100 3777
rect 9158 3743 9192 3777
rect 9250 3743 9284 3777
rect 9342 3743 9376 3777
rect 9434 3743 9468 3777
rect 9526 3743 9560 3777
rect 9618 3743 9652 3777
rect 9710 3743 9744 3777
rect 9802 3743 9836 3777
rect 9894 3743 9928 3777
rect 9986 3743 10020 3777
rect 10078 3743 10112 3777
rect 10170 3743 10204 3777
rect 10262 3743 10296 3777
rect 10354 3743 10388 3777
rect 10446 3743 10480 3777
rect 10538 3743 10572 3777
rect 10630 3743 10664 3777
rect 10722 3743 10756 3777
rect 10814 3743 10848 3777
rect 10906 3743 10940 3777
rect 10998 3743 11032 3777
rect 11090 3743 11124 3777
rect 11182 3743 11216 3777
rect 11274 3743 11308 3777
rect 11366 3743 11400 3777
rect 11458 3743 11492 3777
rect 11550 3743 11584 3777
rect 11642 3743 11676 3777
rect 11734 3743 11768 3777
rect 11826 3743 11860 3777
rect 11918 3743 11952 3777
rect 12010 3743 12044 3777
rect 12102 3743 12136 3777
rect 12194 3743 12228 3777
rect 12286 3743 12320 3777
rect 12378 3743 12412 3777
rect 12470 3743 12504 3777
rect 12562 3743 12596 3777
rect 12654 3743 12688 3777
rect 12746 3743 12780 3777
rect 12838 3743 12872 3777
rect 12930 3743 12964 3777
rect 1062 2870 1096 2904
rect 1154 2870 1188 2904
rect 1246 2870 1280 2904
rect 1338 2870 1372 2904
rect 1430 2870 1464 2904
rect 1522 2870 1556 2904
rect 1614 2870 1648 2904
rect 1706 2870 1740 2904
rect 1798 2870 1832 2904
rect 1890 2870 1924 2904
rect 1982 2870 2016 2904
rect 2074 2870 2108 2904
rect 2166 2870 2200 2904
rect 2258 2870 2292 2904
rect 2350 2870 2384 2904
rect 2442 2870 2476 2904
rect 2534 2870 2568 2904
rect 2626 2870 2660 2904
rect 2718 2870 2752 2904
rect 2810 2870 2844 2904
rect 2902 2870 2936 2904
rect 2994 2870 3028 2904
rect 3086 2870 3120 2904
rect 3178 2870 3212 2904
rect 3270 2870 3304 2904
rect 3362 2870 3396 2904
rect 3454 2870 3488 2904
rect 3546 2870 3580 2904
rect 3638 2870 3672 2904
rect 3730 2870 3764 2904
rect 3822 2870 3856 2904
rect 3914 2870 3948 2904
rect 4006 2870 4040 2904
rect 4098 2870 4132 2904
rect 4190 2870 4224 2904
rect 4282 2870 4316 2904
rect 4374 2870 4408 2904
rect 4466 2870 4500 2904
rect 4558 2870 4592 2904
rect 4650 2870 4684 2904
rect 4742 2870 4776 2904
rect 4834 2870 4868 2904
rect 4926 2870 4960 2904
rect 5018 2870 5052 2904
rect 5110 2870 5144 2904
rect 5202 2870 5236 2904
rect 5294 2870 5328 2904
rect 5386 2870 5420 2904
rect 5478 2870 5512 2904
rect 5570 2870 5604 2904
rect 5662 2870 5696 2904
rect 5754 2870 5788 2904
rect 5846 2870 5880 2904
rect 5938 2870 5972 2904
rect 6030 2870 6064 2904
rect 6122 2870 6156 2904
rect 6214 2870 6248 2904
rect 6306 2870 6340 2904
rect 6398 2870 6432 2904
rect 6490 2870 6524 2904
rect 6582 2870 6616 2904
rect 6674 2870 6708 2904
rect 6766 2870 6800 2904
rect 6858 2870 6892 2904
rect 6950 2870 6984 2904
rect 7042 2870 7076 2904
rect 7134 2870 7168 2904
rect 7226 2870 7260 2904
rect 7318 2870 7352 2904
rect 7410 2870 7444 2904
rect 7502 2870 7536 2904
rect 7594 2870 7628 2904
rect 7686 2870 7720 2904
rect 7778 2870 7812 2904
rect 7870 2870 7904 2904
rect 7962 2870 7996 2904
rect 8054 2870 8088 2904
rect 8146 2870 8180 2904
rect 8238 2870 8272 2904
rect 8330 2870 8364 2904
rect 8422 2870 8456 2904
rect 8514 2870 8548 2904
rect 8606 2870 8640 2904
rect 8698 2870 8732 2904
rect 8790 2870 8824 2904
rect 8882 2870 8916 2904
rect 8974 2870 9008 2904
rect 9066 2870 9100 2904
rect 9158 2870 9192 2904
rect 9250 2870 9284 2904
rect 9342 2870 9376 2904
rect 9434 2870 9468 2904
rect 9526 2870 9560 2904
rect 9618 2870 9652 2904
rect 9710 2870 9744 2904
rect 9802 2870 9836 2904
rect 9894 2870 9928 2904
rect 9986 2870 10020 2904
rect 10078 2870 10112 2904
rect 10170 2870 10204 2904
rect 10262 2870 10296 2904
rect 10354 2870 10388 2904
rect 10446 2870 10480 2904
rect 10538 2870 10572 2904
rect 10630 2870 10664 2904
rect 10722 2870 10756 2904
rect 10814 2870 10848 2904
rect 10906 2870 10940 2904
rect 10998 2870 11032 2904
rect 11090 2870 11124 2904
rect 11182 2870 11216 2904
rect 11274 2870 11308 2904
rect 11366 2870 11400 2904
rect 11458 2870 11492 2904
rect 11550 2870 11584 2904
rect 11642 2870 11676 2904
rect 11734 2870 11768 2904
rect 11826 2870 11860 2904
rect 11918 2870 11952 2904
rect 12010 2870 12044 2904
rect 12102 2870 12136 2904
rect 12194 2870 12228 2904
rect 12286 2870 12320 2904
rect 12378 2870 12412 2904
rect 12470 2870 12504 2904
rect 12562 2870 12596 2904
rect 12654 2870 12688 2904
rect 12746 2870 12780 2904
rect 12838 2870 12872 2904
rect 12930 2870 12964 2904
<< poly >>
rect 2918 5330 2984 5340
rect 2918 5296 2934 5330
rect 2968 5296 2984 5330
rect 4161 5333 4227 5343
rect 2918 5286 2984 5296
rect 4161 5299 4177 5333
rect 4211 5299 4227 5333
rect 6553 5335 6619 5345
rect 4161 5289 4227 5299
rect 6553 5301 6569 5335
rect 6603 5301 6619 5335
rect 8945 5335 9011 5345
rect 6553 5291 6619 5301
rect 8945 5301 8961 5335
rect 8995 5301 9011 5335
rect 11337 5336 11403 5346
rect 8945 5291 9011 5301
rect 11337 5302 11353 5336
rect 11387 5302 11403 5336
rect 11337 5292 11403 5302
rect 2937 5209 2967 5286
rect 4180 5277 4210 5289
rect 6572 5276 6602 5291
rect 8964 5276 8994 5291
rect 11356 5277 11386 5292
rect 4232 4647 4298 4657
rect 4232 4613 4248 4647
rect 4282 4613 4298 4647
rect 6624 4647 6690 4657
rect 4232 4603 4298 4613
rect 6624 4613 6640 4647
rect 6674 4613 6690 4647
rect 9016 4647 9082 4657
rect 6624 4603 6690 4613
rect 9016 4613 9032 4647
rect 9066 4613 9082 4647
rect 11408 4647 11474 4657
rect 9016 4603 9082 4613
rect 11408 4613 11424 4647
rect 11458 4613 11474 4647
rect 11408 4603 11474 4613
rect 4251 4588 4281 4603
rect 6643 4588 6673 4603
rect 9035 4588 9065 4603
rect 11427 4588 11457 4603
<< polycont >>
rect 2934 5296 2968 5330
rect 4177 5299 4211 5333
rect 6569 5301 6603 5335
rect 8961 5301 8995 5335
rect 11353 5302 11387 5336
rect 4248 4613 4282 4647
rect 6640 4613 6674 4647
rect 9032 4613 9066 4647
rect 11424 4613 11458 4647
<< locali >>
rect 1035 6178 1064 6212
rect 1098 6178 1156 6212
rect 1190 6178 1248 6212
rect 1282 6178 1340 6212
rect 1374 6178 1432 6212
rect 1466 6178 1524 6212
rect 1558 6178 1616 6212
rect 1650 6178 1679 6212
rect 2295 6178 2324 6212
rect 2358 6178 2416 6212
rect 2450 6178 2508 6212
rect 2542 6178 2600 6212
rect 2634 6178 2692 6212
rect 2726 6178 2784 6212
rect 2818 6178 2876 6212
rect 2910 6178 2968 6212
rect 3002 6178 3060 6212
rect 3094 6178 3152 6212
rect 3186 6178 3244 6212
rect 3278 6178 3336 6212
rect 3370 6178 3428 6212
rect 3462 6178 3520 6212
rect 3554 6178 3612 6212
rect 3646 6178 3704 6212
rect 3738 6178 3796 6212
rect 3830 6178 3888 6212
rect 3922 6178 3980 6212
rect 4014 6178 4072 6212
rect 4106 6178 4135 6212
rect 1035 6154 1679 6178
rect 1271 5846 1361 5884
rect 1540 5849 1712 5883
rect 1746 5849 1756 5883
rect 4133 5625 4136 5644
rect 1035 5620 4136 5625
rect 1035 5586 1064 5620
rect 1098 5586 1156 5620
rect 1190 5586 1248 5620
rect 1282 5586 1340 5620
rect 1374 5586 1432 5620
rect 1466 5586 1524 5620
rect 1558 5586 1616 5620
rect 1650 5586 1708 5620
rect 1742 5586 1800 5620
rect 1834 5586 1892 5620
rect 1926 5586 1984 5620
rect 2018 5586 2076 5620
rect 2110 5586 2168 5620
rect 2202 5586 2260 5620
rect 2294 5586 2352 5620
rect 2386 5586 2444 5620
rect 2478 5586 2536 5620
rect 2570 5586 2628 5620
rect 2662 5586 2720 5620
rect 2754 5586 2812 5620
rect 2846 5586 2904 5620
rect 2938 5586 2996 5620
rect 3030 5586 3088 5620
rect 3122 5586 3180 5620
rect 3214 5586 3272 5620
rect 3306 5586 3364 5620
rect 3398 5586 3456 5620
rect 3490 5586 3548 5620
rect 3582 5586 3640 5620
rect 3674 5586 3732 5620
rect 3766 5586 3824 5620
rect 3858 5586 3916 5620
rect 3950 5586 4008 5620
rect 4042 5586 4136 5620
rect 1034 5305 1063 5339
rect 1097 5305 1155 5339
rect 1189 5305 1247 5339
rect 1281 5305 1339 5339
rect 1373 5305 1431 5339
rect 1465 5305 1523 5339
rect 1557 5305 1615 5339
rect 1649 5305 1707 5339
rect 1741 5305 1799 5339
rect 1833 5305 1891 5339
rect 1925 5305 1983 5339
rect 2017 5305 2075 5339
rect 2109 5305 2167 5339
rect 2201 5305 2259 5339
rect 2293 5305 2351 5339
rect 2385 5305 2443 5339
rect 2477 5305 2535 5339
rect 2569 5305 2627 5339
rect 2661 5305 2719 5339
rect 2753 5305 2811 5339
rect 2845 5330 3087 5339
rect 2845 5305 2934 5330
rect 2918 5296 2934 5305
rect 2968 5305 3087 5330
rect 3121 5305 3179 5339
rect 3213 5305 3271 5339
rect 3305 5305 3363 5339
rect 3397 5305 3455 5339
rect 3489 5305 3547 5339
rect 3581 5305 3640 5339
rect 3674 5305 3731 5339
rect 3765 5305 3823 5339
rect 3857 5305 3915 5339
rect 3949 5305 4007 5339
rect 4041 5333 4283 5339
rect 4041 5305 4177 5333
rect 2968 5296 2984 5305
rect 4161 5299 4177 5305
rect 4211 5305 4283 5333
rect 4317 5305 4375 5339
rect 4409 5305 4467 5339
rect 4501 5305 4559 5339
rect 4593 5305 4651 5339
rect 4685 5305 4743 5339
rect 4777 5305 4835 5339
rect 4869 5305 4927 5339
rect 4961 5305 5019 5339
rect 5053 5305 5111 5339
rect 5145 5305 5203 5339
rect 5237 5305 5295 5339
rect 5329 5305 5387 5339
rect 5421 5305 5479 5339
rect 5513 5305 5571 5339
rect 5605 5305 5663 5339
rect 5697 5305 5755 5339
rect 5789 5305 5847 5339
rect 5881 5305 5939 5339
rect 5973 5305 6031 5339
rect 6065 5305 6123 5339
rect 6157 5305 6215 5339
rect 6249 5305 6307 5339
rect 6341 5305 6399 5339
rect 6433 5335 6675 5339
rect 6433 5305 6569 5335
rect 4211 5299 4227 5305
rect 4161 5296 4227 5299
rect 6553 5301 6569 5305
rect 6603 5305 6675 5335
rect 6709 5305 6767 5339
rect 6801 5305 6859 5339
rect 6893 5305 6951 5339
rect 6985 5305 7043 5339
rect 7077 5305 7135 5339
rect 7169 5305 7227 5339
rect 7261 5305 7319 5339
rect 7353 5305 7411 5339
rect 7445 5305 7503 5339
rect 7537 5305 7595 5339
rect 7629 5305 7687 5339
rect 7721 5305 7779 5339
rect 7813 5305 7871 5339
rect 7905 5305 7963 5339
rect 7997 5305 8055 5339
rect 8089 5305 8147 5339
rect 8181 5305 8239 5339
rect 8273 5305 8331 5339
rect 8365 5305 8423 5339
rect 8457 5305 8515 5339
rect 8549 5305 8607 5339
rect 8641 5305 8699 5339
rect 8733 5305 8791 5339
rect 8825 5335 9067 5339
rect 8825 5305 8961 5335
rect 6603 5301 6619 5305
rect 2918 5286 2984 5296
rect 6553 5291 6619 5301
rect 8945 5301 8961 5305
rect 8995 5305 9067 5335
rect 9101 5305 9159 5339
rect 9193 5305 9251 5339
rect 9285 5305 9343 5339
rect 9377 5305 9435 5339
rect 9469 5305 9527 5339
rect 9561 5305 9619 5339
rect 9653 5305 9711 5339
rect 9745 5305 9803 5339
rect 9837 5305 9895 5339
rect 9929 5305 9987 5339
rect 10021 5305 10079 5339
rect 10113 5305 10171 5339
rect 10205 5305 10263 5339
rect 10297 5305 10355 5339
rect 10389 5305 10447 5339
rect 10481 5305 10539 5339
rect 10573 5305 10631 5339
rect 10665 5305 10723 5339
rect 10757 5305 10815 5339
rect 10849 5305 10907 5339
rect 10941 5305 10999 5339
rect 11033 5305 11091 5339
rect 11125 5305 11183 5339
rect 11217 5336 11459 5339
rect 11217 5305 11353 5336
rect 8995 5301 9011 5305
rect 8945 5291 9011 5301
rect 11337 5302 11353 5305
rect 11387 5305 11459 5336
rect 11493 5305 11551 5339
rect 11585 5305 11643 5339
rect 11677 5305 11735 5339
rect 11769 5305 11827 5339
rect 11861 5305 11919 5339
rect 11953 5305 12011 5339
rect 12045 5305 12103 5339
rect 12137 5305 12195 5339
rect 12229 5305 12287 5339
rect 12321 5305 12379 5339
rect 12413 5305 12471 5339
rect 12505 5305 12563 5339
rect 12597 5305 12655 5339
rect 12689 5305 12747 5339
rect 12781 5305 12839 5339
rect 12873 5305 12931 5339
rect 12965 5305 12994 5339
rect 11387 5302 11403 5305
rect 11337 5292 11403 5302
rect 1034 4713 1063 4747
rect 1097 4713 1155 4747
rect 1189 4713 1247 4747
rect 1281 4713 1339 4747
rect 1373 4713 1431 4747
rect 1465 4713 1523 4747
rect 1557 4713 1615 4747
rect 1649 4713 1707 4747
rect 1741 4713 1799 4747
rect 1833 4713 1891 4747
rect 1925 4713 1983 4747
rect 2017 4713 2075 4747
rect 2109 4713 2167 4747
rect 2201 4713 2259 4747
rect 2293 4713 2351 4747
rect 2385 4713 2443 4747
rect 2477 4713 2535 4747
rect 2569 4713 2627 4747
rect 2661 4713 2719 4747
rect 2753 4713 2811 4747
rect 2845 4713 2903 4747
rect 2937 4713 2995 4747
rect 3029 4713 3087 4747
rect 3121 4713 3179 4747
rect 3213 4713 3271 4747
rect 3305 4713 3363 4747
rect 3397 4713 3455 4747
rect 3489 4713 3547 4747
rect 3581 4713 3639 4747
rect 3673 4713 3731 4747
rect 3765 4713 3823 4747
rect 3857 4713 3915 4747
rect 3949 4713 4007 4747
rect 4041 4713 4099 4747
rect 4133 4713 4191 4747
rect 4225 4713 4283 4747
rect 4317 4713 4375 4747
rect 4409 4713 4467 4747
rect 4501 4713 4559 4747
rect 4593 4713 4651 4747
rect 4685 4713 4743 4747
rect 4777 4713 4835 4747
rect 4869 4713 4927 4747
rect 4961 4713 5019 4747
rect 5053 4713 5111 4747
rect 5145 4713 5203 4747
rect 5237 4713 5295 4747
rect 5329 4713 5387 4747
rect 5421 4713 5479 4747
rect 5513 4713 5571 4747
rect 5605 4713 5663 4747
rect 5697 4713 5755 4747
rect 5789 4713 5847 4747
rect 5881 4713 5939 4747
rect 5973 4713 6031 4747
rect 6065 4713 6123 4747
rect 6157 4713 6215 4747
rect 6249 4713 6307 4747
rect 6341 4713 6399 4747
rect 6433 4713 6491 4747
rect 6525 4713 6583 4747
rect 6617 4713 6675 4747
rect 6709 4713 6767 4747
rect 6801 4713 6859 4747
rect 6893 4713 6951 4747
rect 6985 4713 7043 4747
rect 7077 4713 7135 4747
rect 7169 4713 7227 4747
rect 7261 4713 7319 4747
rect 7353 4713 7411 4747
rect 7445 4713 7503 4747
rect 7537 4713 7595 4747
rect 7629 4713 7687 4747
rect 7721 4713 7779 4747
rect 7813 4713 7871 4747
rect 7905 4713 7963 4747
rect 7997 4713 8055 4747
rect 8089 4713 8147 4747
rect 8181 4713 8239 4747
rect 8273 4713 8331 4747
rect 8365 4713 8423 4747
rect 8457 4713 8515 4747
rect 8549 4713 8607 4747
rect 8641 4713 8699 4747
rect 8733 4713 8791 4747
rect 8825 4713 8883 4747
rect 8917 4713 8975 4747
rect 9009 4713 9067 4747
rect 9101 4713 9159 4747
rect 9193 4713 9251 4747
rect 9285 4713 9343 4747
rect 9377 4713 9435 4747
rect 9469 4713 9527 4747
rect 9561 4713 9619 4747
rect 9653 4713 9711 4747
rect 9745 4713 9803 4747
rect 9837 4713 9895 4747
rect 9929 4713 9987 4747
rect 10021 4713 10079 4747
rect 10113 4713 10171 4747
rect 10205 4713 10263 4747
rect 10297 4713 10355 4747
rect 10389 4713 10447 4747
rect 10481 4713 10539 4747
rect 10573 4713 10631 4747
rect 10665 4713 10723 4747
rect 10757 4713 10815 4747
rect 10849 4713 10907 4747
rect 10941 4713 10999 4747
rect 11033 4713 11091 4747
rect 11125 4713 11183 4747
rect 11217 4713 11275 4747
rect 11309 4713 11367 4747
rect 11401 4713 11459 4747
rect 11493 4713 11551 4747
rect 11585 4713 11643 4747
rect 11677 4713 11735 4747
rect 11769 4713 11827 4747
rect 11861 4713 11919 4747
rect 11953 4713 12011 4747
rect 12045 4713 12103 4747
rect 12137 4713 12195 4747
rect 12229 4713 12287 4747
rect 12321 4713 12379 4747
rect 12413 4713 12471 4747
rect 12505 4713 12563 4747
rect 12597 4713 12655 4747
rect 12689 4713 12747 4747
rect 12781 4713 12839 4747
rect 12873 4713 12931 4747
rect 12965 4713 12994 4747
rect 594 4616 623 4650
rect 657 4616 715 4650
rect 749 4616 807 4650
rect 841 4616 899 4650
rect 933 4616 991 4650
rect 1025 4616 1083 4650
rect 1117 4616 1175 4650
rect 1209 4616 1267 4650
rect 1301 4616 1359 4650
rect 1393 4616 1451 4650
rect 1485 4616 1543 4650
rect 1577 4616 1635 4650
rect 1669 4616 1727 4650
rect 1761 4616 1819 4650
rect 1853 4616 1911 4650
rect 1945 4616 2003 4650
rect 2037 4616 2095 4650
rect 2129 4616 2187 4650
rect 2221 4616 2279 4650
rect 2313 4616 2351 4650
rect 2405 4616 2443 4650
rect 2477 4616 2535 4650
rect 2569 4616 2627 4650
rect 2661 4616 2719 4650
rect 2753 4616 2811 4650
rect 2845 4616 2903 4650
rect 2937 4616 2995 4650
rect 3029 4616 3087 4650
rect 3121 4616 3179 4650
rect 3213 4616 3271 4650
rect 3305 4616 3363 4650
rect 3397 4616 3455 4650
rect 3489 4616 3547 4650
rect 3581 4616 3639 4650
rect 3673 4616 3731 4650
rect 3765 4616 3823 4650
rect 3857 4616 3915 4650
rect 3949 4616 4007 4650
rect 4041 4616 4099 4650
rect 4133 4647 4375 4650
rect 4133 4616 4248 4647
rect 4232 4613 4248 4616
rect 4282 4616 4375 4647
rect 4409 4616 4467 4650
rect 4501 4616 4559 4650
rect 4593 4616 4651 4650
rect 4685 4616 4743 4650
rect 4777 4616 4835 4650
rect 4869 4616 4927 4650
rect 4961 4616 5019 4650
rect 5053 4616 5111 4650
rect 5145 4616 5203 4650
rect 5237 4616 5295 4650
rect 5329 4616 5387 4650
rect 5421 4616 5479 4650
rect 5513 4616 5571 4650
rect 5605 4616 5663 4650
rect 5697 4616 5755 4650
rect 5789 4616 5847 4650
rect 5881 4616 5939 4650
rect 5973 4616 6031 4650
rect 6065 4616 6123 4650
rect 6157 4616 6215 4650
rect 6249 4616 6307 4650
rect 6341 4616 6399 4650
rect 6433 4616 6491 4650
rect 6525 4647 6767 4650
rect 6525 4616 6640 4647
rect 4282 4613 4298 4616
rect 4232 4603 4298 4613
rect 6624 4613 6640 4616
rect 6674 4616 6767 4647
rect 6801 4616 6859 4650
rect 6893 4616 6951 4650
rect 6985 4616 7043 4650
rect 7077 4616 7135 4650
rect 7169 4616 7227 4650
rect 7261 4616 7319 4650
rect 7353 4616 7411 4650
rect 7445 4616 7503 4650
rect 7537 4616 7595 4650
rect 7629 4616 7687 4650
rect 7721 4616 7779 4650
rect 7813 4616 7871 4650
rect 7905 4616 7963 4650
rect 7997 4616 8055 4650
rect 8089 4616 8147 4650
rect 8181 4616 8239 4650
rect 8273 4616 8331 4650
rect 8365 4616 8423 4650
rect 8457 4616 8515 4650
rect 8549 4616 8607 4650
rect 8641 4616 8699 4650
rect 8733 4616 8791 4650
rect 8825 4616 8883 4650
rect 8917 4647 9159 4650
rect 8917 4616 9032 4647
rect 6674 4613 6690 4616
rect 6624 4603 6690 4613
rect 9016 4613 9032 4616
rect 9066 4616 9159 4647
rect 9193 4616 9251 4650
rect 9285 4616 9343 4650
rect 9377 4616 9435 4650
rect 9469 4616 9527 4650
rect 9561 4616 9619 4650
rect 9653 4616 9711 4650
rect 9745 4616 9803 4650
rect 9837 4616 9895 4650
rect 9929 4616 9987 4650
rect 10021 4616 10079 4650
rect 10113 4616 10171 4650
rect 10205 4616 10263 4650
rect 10297 4616 10355 4650
rect 10389 4616 10447 4650
rect 10481 4616 10539 4650
rect 10573 4616 10631 4650
rect 10665 4616 10723 4650
rect 10757 4616 10815 4650
rect 10849 4616 10907 4650
rect 10941 4616 10999 4650
rect 11033 4616 11091 4650
rect 11125 4616 11183 4650
rect 11217 4616 11275 4650
rect 11309 4647 11551 4650
rect 11309 4616 11424 4647
rect 9066 4613 9082 4616
rect 9016 4603 9082 4613
rect 11408 4613 11424 4616
rect 11458 4616 11551 4647
rect 11585 4616 11643 4650
rect 11677 4616 11735 4650
rect 11769 4616 11827 4650
rect 11861 4616 11919 4650
rect 11953 4616 12011 4650
rect 12045 4616 12103 4650
rect 12137 4616 12195 4650
rect 12229 4616 12287 4650
rect 12321 4616 12379 4650
rect 12413 4616 12471 4650
rect 12505 4618 12563 4650
rect 12505 4616 12554 4618
rect 12597 4618 12655 4650
rect 12689 4618 12747 4650
rect 12781 4618 12839 4650
rect 12873 4618 12931 4650
rect 12965 4616 12994 4650
rect 11458 4613 11474 4616
rect 11408 4603 11474 4613
rect 831 4282 931 4327
rect 1267 4280 1464 4320
rect 594 4024 623 4058
rect 657 4024 715 4058
rect 749 4024 807 4058
rect 841 4024 899 4058
rect 933 4024 991 4058
rect 1025 4024 1083 4058
rect 1117 4024 1175 4058
rect 1209 4024 1267 4058
rect 1301 4024 1359 4058
rect 1393 4024 1451 4058
rect 1485 4024 1543 4058
rect 1577 4024 1635 4058
rect 1669 4024 1727 4058
rect 1761 4024 1819 4058
rect 1853 4024 1911 4058
rect 1945 4024 2003 4058
rect 2037 4024 2095 4058
rect 2129 4024 2187 4058
rect 2221 4024 2279 4058
rect 2313 4024 2371 4058
rect 2405 4024 2463 4058
rect 2497 4024 2555 4058
rect 2589 4024 2647 4058
rect 2681 4024 2739 4058
rect 2773 4024 2831 4058
rect 2865 4024 2923 4058
rect 2957 4024 3015 4058
rect 3049 4024 3107 4058
rect 3141 4024 3199 4058
rect 3233 4024 3291 4058
rect 3325 4024 3383 4058
rect 3417 4024 3475 4058
rect 3509 4024 3567 4058
rect 3601 4024 3659 4058
rect 3693 4024 3751 4058
rect 3785 4024 3843 4058
rect 3877 4024 3935 4058
rect 3969 4024 4027 4058
rect 4061 4024 4119 4058
rect 4153 4024 4211 4058
rect 4245 4024 4303 4058
rect 4337 4024 4395 4058
rect 4429 4024 4487 4058
rect 4521 4024 4579 4058
rect 4613 4024 4671 4058
rect 4705 4024 4763 4058
rect 4797 4024 4855 4058
rect 4889 4024 4947 4058
rect 4981 4024 5039 4058
rect 5073 4024 5131 4058
rect 5165 4024 5223 4058
rect 5257 4024 5315 4058
rect 5349 4024 5407 4058
rect 5441 4024 5499 4058
rect 5533 4024 5591 4058
rect 5625 4024 5683 4058
rect 5717 4024 5775 4058
rect 5809 4024 5867 4058
rect 5901 4024 5959 4058
rect 5993 4024 6051 4058
rect 6085 4024 6143 4058
rect 6177 4024 6235 4058
rect 6269 4024 6327 4058
rect 6361 4024 6419 4058
rect 6453 4024 6511 4058
rect 6545 4024 6603 4058
rect 6637 4024 6695 4058
rect 6729 4024 6787 4058
rect 6821 4024 6879 4058
rect 6913 4024 6971 4058
rect 7005 4024 7063 4058
rect 7097 4024 7155 4058
rect 7189 4024 7247 4058
rect 7281 4024 7339 4058
rect 7373 4024 7431 4058
rect 7465 4024 7523 4058
rect 7557 4024 7615 4058
rect 7649 4024 7707 4058
rect 7741 4024 7799 4058
rect 7833 4024 7891 4058
rect 7925 4024 7983 4058
rect 8017 4024 8075 4058
rect 8109 4024 8167 4058
rect 8201 4024 8259 4058
rect 8293 4024 8351 4058
rect 8385 4024 8443 4058
rect 8477 4024 8535 4058
rect 8569 4024 8627 4058
rect 8661 4024 8719 4058
rect 8753 4024 8811 4058
rect 8845 4024 8903 4058
rect 8937 4024 8995 4058
rect 9029 4024 9087 4058
rect 9121 4024 9179 4058
rect 9213 4024 9271 4058
rect 9305 4024 9363 4058
rect 9397 4024 9435 4058
rect 9469 4024 9527 4058
rect 9561 4024 9619 4058
rect 9653 4024 9711 4058
rect 9745 4024 9803 4058
rect 9837 4024 9895 4058
rect 9929 4024 9987 4058
rect 10021 4024 10079 4058
rect 10113 4024 10171 4058
rect 10205 4024 10263 4058
rect 10297 4024 10355 4058
rect 10389 4024 10447 4058
rect 10481 4024 10539 4058
rect 10573 4024 10631 4058
rect 10665 4024 10723 4058
rect 10757 4024 10815 4058
rect 10849 4024 10907 4058
rect 10941 4024 10999 4058
rect 11033 4024 11091 4058
rect 11125 4024 11183 4058
rect 11217 4024 11275 4058
rect 11309 4024 11367 4058
rect 11401 4024 11459 4058
rect 11493 4024 11551 4058
rect 11585 4024 11643 4058
rect 11677 4024 11735 4058
rect 11769 4024 11827 4058
rect 11861 4024 11919 4058
rect 11953 4024 12011 4058
rect 12045 4024 12103 4058
rect 12137 4024 12195 4058
rect 12229 4024 12287 4058
rect 12321 4024 12379 4058
rect 12413 4024 12471 4058
rect 12505 4024 12563 4058
rect 12597 4024 12655 4058
rect 12689 4024 12747 4058
rect 12781 4024 12839 4058
rect 12873 4024 12931 4058
rect 12965 4024 12994 4058
rect 3168 3743 3197 3777
rect 3231 3743 3289 3777
rect 3323 3743 3381 3777
rect 3415 3743 3473 3777
rect 3507 3743 3565 3777
rect 3599 3743 3657 3777
rect 3691 3743 3749 3777
rect 3783 3743 3841 3777
rect 3875 3743 3933 3777
rect 3967 3743 4025 3777
rect 4059 3743 4117 3777
rect 4151 3743 4209 3777
rect 4243 3743 4301 3777
rect 4335 3743 4393 3777
rect 4427 3743 4485 3777
rect 4519 3743 4577 3777
rect 4611 3743 4669 3777
rect 4703 3743 4761 3777
rect 4795 3743 4853 3777
rect 4887 3743 4945 3777
rect 4979 3743 5018 3777
rect 5052 3743 5110 3777
rect 5144 3743 5202 3777
rect 5236 3743 5294 3777
rect 5328 3743 5386 3777
rect 5420 3743 5478 3777
rect 5512 3743 5570 3777
rect 5604 3743 5662 3777
rect 5696 3743 5754 3777
rect 5788 3743 5846 3777
rect 5880 3743 5938 3777
rect 5972 3743 6030 3777
rect 6064 3743 6122 3777
rect 6156 3743 6214 3777
rect 6248 3743 6306 3777
rect 6340 3743 6398 3777
rect 6432 3743 6490 3777
rect 6524 3743 6582 3777
rect 6616 3743 6674 3777
rect 6708 3743 6766 3777
rect 6800 3743 6858 3777
rect 6892 3743 6950 3777
rect 6984 3743 7042 3777
rect 7076 3743 7134 3777
rect 7168 3743 7226 3777
rect 7260 3743 7318 3777
rect 7352 3743 7410 3777
rect 7444 3743 7502 3777
rect 7536 3743 7594 3777
rect 7628 3743 7686 3777
rect 7720 3743 7778 3777
rect 7812 3743 7870 3777
rect 7904 3743 7962 3777
rect 7996 3743 8054 3777
rect 8088 3743 8146 3777
rect 8180 3743 8238 3777
rect 8272 3743 8330 3777
rect 8364 3743 8422 3777
rect 8456 3743 8514 3777
rect 8548 3743 8606 3777
rect 8640 3743 8698 3777
rect 8732 3743 8790 3777
rect 8824 3743 8882 3777
rect 8916 3743 8974 3777
rect 9008 3743 9066 3777
rect 9100 3743 9158 3777
rect 9192 3743 9250 3777
rect 9284 3743 9342 3777
rect 9376 3743 9434 3777
rect 9468 3743 9526 3777
rect 9560 3743 9618 3777
rect 9652 3743 9710 3777
rect 9744 3743 9802 3777
rect 9836 3743 9894 3777
rect 9928 3743 9986 3777
rect 10020 3743 10078 3777
rect 10112 3743 10170 3777
rect 10204 3743 10262 3777
rect 10296 3743 10354 3777
rect 10388 3743 10446 3777
rect 10480 3743 10538 3777
rect 10572 3743 10630 3777
rect 10664 3743 10722 3777
rect 10756 3743 10814 3777
rect 10848 3743 10906 3777
rect 10940 3743 10998 3777
rect 11032 3743 11090 3777
rect 11124 3743 11182 3777
rect 11216 3743 11274 3777
rect 11308 3743 11366 3777
rect 11400 3743 11458 3777
rect 11492 3743 11550 3777
rect 11584 3743 11642 3777
rect 11676 3743 11734 3777
rect 11768 3743 11826 3777
rect 11860 3743 11918 3777
rect 11952 3743 12010 3777
rect 12044 3743 12102 3777
rect 12136 3743 12194 3777
rect 12228 3743 12286 3777
rect 12320 3743 12378 3777
rect 12412 3743 12470 3777
rect 12504 3743 12562 3777
rect 12596 3743 12654 3777
rect 12688 3743 12746 3777
rect 12780 3743 12838 3777
rect 12872 3743 12930 3777
rect 12964 3743 12993 3777
rect 3160 3446 3236 3455
rect 3160 3412 3162 3446
rect 3196 3412 3236 3446
rect 3160 3407 3236 3412
rect 5770 3423 5896 3471
rect 8169 3424 8295 3472
rect 10553 3415 10679 3463
rect 3167 3151 3197 3185
rect 3231 3151 3289 3185
rect 3323 3151 3381 3185
rect 3415 3151 3473 3185
rect 3507 3151 3565 3185
rect 3599 3151 3657 3185
rect 3691 3151 3749 3185
rect 3783 3151 3841 3185
rect 3875 3151 3933 3185
rect 3967 3151 4025 3185
rect 4059 3151 4117 3185
rect 4151 3151 4209 3185
rect 4243 3151 4301 3185
rect 4335 3151 4393 3185
rect 4427 3151 4485 3185
rect 4519 3151 4577 3185
rect 4611 3151 4669 3185
rect 4703 3151 4761 3185
rect 4795 3151 4853 3185
rect 4887 3151 4945 3185
rect 4979 3151 5037 3185
rect 5071 3151 5129 3185
rect 5163 3151 5221 3185
rect 5255 3151 5313 3185
rect 5347 3151 5405 3185
rect 5439 3151 5497 3185
rect 5531 3151 5589 3185
rect 5623 3151 5681 3185
rect 5715 3151 5773 3185
rect 5807 3151 5865 3185
rect 5899 3151 5957 3185
rect 5991 3151 6049 3185
rect 6083 3151 6141 3185
rect 6175 3151 6233 3185
rect 6267 3151 6325 3185
rect 6359 3151 6417 3185
rect 6451 3151 6509 3185
rect 6543 3151 6601 3185
rect 6635 3151 6693 3185
rect 6727 3151 6785 3185
rect 6819 3151 6877 3185
rect 6911 3151 6969 3185
rect 7003 3151 7061 3185
rect 7095 3151 7153 3185
rect 7187 3151 7245 3185
rect 7279 3151 7337 3185
rect 7371 3151 7429 3185
rect 7463 3151 7521 3185
rect 7555 3151 7613 3185
rect 7647 3151 7705 3185
rect 7739 3151 7797 3185
rect 7831 3151 7889 3185
rect 7923 3151 7981 3185
rect 8015 3151 8073 3185
rect 8107 3151 8165 3185
rect 8199 3151 8257 3185
rect 8291 3151 8349 3185
rect 8383 3151 8441 3185
rect 8475 3151 8533 3185
rect 8567 3151 8625 3185
rect 8659 3151 8717 3185
rect 8751 3151 8809 3185
rect 8843 3151 8901 3185
rect 8935 3151 8993 3185
rect 9027 3151 9085 3185
rect 9119 3151 9177 3185
rect 9211 3151 9269 3185
rect 9303 3151 9361 3185
rect 9395 3151 9453 3185
rect 9487 3151 9545 3185
rect 9579 3151 9637 3185
rect 9671 3151 9729 3185
rect 9763 3151 9821 3185
rect 9855 3151 9894 3185
rect 9947 3151 9986 3185
rect 10039 3151 10078 3185
rect 10131 3151 10170 3185
rect 10223 3151 10262 3185
rect 10315 3151 10354 3185
rect 10407 3151 10446 3185
rect 10499 3151 10538 3185
rect 10591 3151 10630 3185
rect 10683 3151 10722 3185
rect 10775 3151 10814 3185
rect 10867 3151 10906 3185
rect 10959 3151 10998 3185
rect 11051 3151 11090 3185
rect 11143 3151 11182 3185
rect 11235 3151 11274 3185
rect 11327 3151 11366 3185
rect 11419 3151 11458 3185
rect 11511 3151 11550 3185
rect 11603 3151 11642 3185
rect 11695 3151 11734 3185
rect 11787 3151 11826 3185
rect 11879 3151 11918 3185
rect 11971 3151 12010 3185
rect 12044 3151 12102 3185
rect 12136 3151 12194 3185
rect 12228 3151 12286 3185
rect 12320 3151 12378 3185
rect 12412 3151 12470 3185
rect 12504 3151 12562 3185
rect 12596 3151 12654 3185
rect 12688 3151 12746 3185
rect 12780 3151 12838 3185
rect 12872 3151 12930 3185
rect 12964 3151 12992 3185
rect 1033 2870 1062 2904
rect 1096 2870 1154 2904
rect 1188 2870 1246 2904
rect 1280 2870 1338 2904
rect 1372 2870 1430 2904
rect 1464 2870 1522 2904
rect 1556 2870 1614 2904
rect 1648 2870 1706 2904
rect 1740 2870 1798 2904
rect 1832 2870 1890 2904
rect 1924 2870 1982 2904
rect 2016 2870 2074 2904
rect 2108 2870 2166 2904
rect 2200 2870 2258 2904
rect 2292 2870 2350 2904
rect 2384 2870 2442 2904
rect 2476 2870 2534 2904
rect 2568 2870 2626 2904
rect 2660 2870 2718 2904
rect 2752 2870 2810 2904
rect 2844 2870 2902 2904
rect 2936 2870 2994 2904
rect 3028 2870 3086 2904
rect 3120 2870 3178 2904
rect 3212 2870 3270 2904
rect 3304 2870 3362 2904
rect 3396 2870 3454 2904
rect 3488 2870 3546 2904
rect 3580 2870 3638 2904
rect 3672 2870 3730 2904
rect 3764 2870 3822 2904
rect 3856 2870 3914 2904
rect 3948 2870 4006 2904
rect 4040 2870 4098 2904
rect 4132 2870 4190 2904
rect 4224 2870 4282 2904
rect 4316 2870 4374 2904
rect 4408 2870 4466 2904
rect 4500 2870 4558 2904
rect 4592 2870 4650 2904
rect 4684 2870 4742 2904
rect 4776 2870 4834 2904
rect 4868 2870 4926 2904
rect 4960 2870 5018 2904
rect 5052 2870 5110 2904
rect 5144 2870 5202 2904
rect 5236 2870 5294 2904
rect 5328 2870 5386 2904
rect 5420 2870 5478 2904
rect 5512 2870 5570 2904
rect 5604 2870 5662 2904
rect 5696 2870 5754 2904
rect 5788 2870 5846 2904
rect 5880 2870 5938 2904
rect 5972 2870 6030 2904
rect 6064 2870 6122 2904
rect 6156 2870 6214 2904
rect 6248 2870 6306 2904
rect 6340 2870 6398 2904
rect 6432 2870 6490 2904
rect 6524 2870 6582 2904
rect 6616 2870 6674 2904
rect 6708 2870 6766 2904
rect 6800 2870 6858 2904
rect 6892 2870 6950 2904
rect 6984 2870 7042 2904
rect 7076 2870 7134 2904
rect 7168 2870 7226 2904
rect 7260 2870 7318 2904
rect 7352 2870 7410 2904
rect 7444 2870 7502 2904
rect 7536 2870 7594 2904
rect 7628 2870 7686 2904
rect 7720 2870 7778 2904
rect 7812 2870 7870 2904
rect 7904 2870 7962 2904
rect 7996 2870 8054 2904
rect 8088 2870 8146 2904
rect 8180 2870 8238 2904
rect 8272 2870 8330 2904
rect 8364 2870 8422 2904
rect 8456 2870 8514 2904
rect 8548 2870 8606 2904
rect 8640 2870 8698 2904
rect 8732 2870 8790 2904
rect 8824 2870 8882 2904
rect 8916 2870 8974 2904
rect 9008 2870 9066 2904
rect 9100 2870 9158 2904
rect 9192 2870 9250 2904
rect 9284 2870 9342 2904
rect 9376 2870 9434 2904
rect 9468 2870 9526 2904
rect 9560 2870 9618 2904
rect 9652 2870 9710 2904
rect 9744 2870 9802 2904
rect 9836 2870 9894 2904
rect 9928 2870 9986 2904
rect 10020 2870 10078 2904
rect 10112 2870 10170 2904
rect 10204 2870 10262 2904
rect 10296 2870 10354 2904
rect 10388 2870 10446 2904
rect 10480 2870 10538 2904
rect 10572 2870 10630 2904
rect 10664 2870 10722 2904
rect 10756 2870 10814 2904
rect 10848 2870 10906 2904
rect 10940 2870 10998 2904
rect 11032 2870 11090 2904
rect 11124 2870 11182 2904
rect 11216 2870 11274 2904
rect 11308 2870 11366 2904
rect 11400 2870 11458 2904
rect 11492 2870 11550 2904
rect 11584 2870 11642 2904
rect 11676 2870 11734 2904
rect 11768 2870 11826 2904
rect 11860 2870 11918 2904
rect 11952 2870 12010 2904
rect 12044 2870 12102 2904
rect 12136 2870 12194 2904
rect 12228 2870 12286 2904
rect 12320 2870 12378 2904
rect 12412 2870 12470 2904
rect 12504 2870 12562 2904
rect 12596 2870 12654 2904
rect 12688 2870 12746 2904
rect 12780 2870 12838 2904
rect 12872 2870 12930 2904
rect 12964 2870 12993 2904
rect 3348 2534 3474 2582
rect 5737 2537 5863 2585
rect 8135 2538 8261 2586
rect 10516 2527 10642 2575
rect 1033 2278 1062 2312
rect 1096 2278 1154 2312
rect 1188 2278 1246 2312
rect 1280 2278 1338 2312
rect 1372 2278 1430 2312
rect 1464 2278 1522 2312
rect 1556 2278 1614 2312
rect 1648 2278 1706 2312
rect 1740 2278 1798 2312
rect 1832 2278 1890 2312
rect 1924 2278 1982 2312
rect 2016 2278 2074 2312
rect 2108 2278 2166 2312
rect 2200 2278 2258 2312
rect 2292 2278 2350 2312
rect 2384 2278 2442 2312
rect 2476 2278 2534 2312
rect 2568 2278 2626 2312
rect 2660 2278 2718 2312
rect 2752 2278 2810 2312
rect 2844 2278 2902 2312
rect 2936 2278 2994 2312
rect 3028 2278 3086 2312
rect 3120 2278 3178 2312
rect 3212 2278 3270 2312
rect 3304 2278 3362 2312
rect 3396 2278 3454 2312
rect 3488 2278 3546 2312
rect 3580 2278 3638 2312
rect 3672 2278 3730 2312
rect 3764 2278 3822 2312
rect 3856 2278 3914 2312
rect 3948 2278 4006 2312
rect 4040 2278 4098 2312
rect 4132 2278 4190 2312
rect 4224 2278 4282 2312
rect 4316 2278 4374 2312
rect 4408 2278 4466 2312
rect 4500 2278 4558 2312
rect 4592 2278 4650 2312
rect 4684 2278 4742 2312
rect 4776 2278 4834 2312
rect 4868 2278 4926 2312
rect 4960 2278 5018 2312
rect 5052 2278 5110 2312
rect 5144 2278 5202 2312
rect 5236 2278 5294 2312
rect 5328 2278 5386 2312
rect 5420 2278 5478 2312
rect 5512 2278 5570 2312
rect 5604 2278 5662 2312
rect 5696 2278 5754 2312
rect 5788 2278 5846 2312
rect 5880 2278 5938 2312
rect 5972 2278 6030 2312
rect 6064 2278 6122 2312
rect 6156 2278 6214 2312
rect 6248 2278 6306 2312
rect 6340 2278 6398 2312
rect 6432 2278 6490 2312
rect 6524 2278 6582 2312
rect 6616 2278 6674 2312
rect 6708 2278 6766 2312
rect 6800 2278 6858 2312
rect 6892 2278 6950 2312
rect 6984 2278 7042 2312
rect 7076 2278 7134 2312
rect 7168 2278 7226 2312
rect 7260 2278 7318 2312
rect 7352 2278 7410 2312
rect 7444 2278 7502 2312
rect 7536 2278 7594 2312
rect 7628 2278 7686 2312
rect 7720 2278 7778 2312
rect 7812 2278 7870 2312
rect 7904 2278 7962 2312
rect 7996 2278 8054 2312
rect 8088 2278 8146 2312
rect 8180 2278 8238 2312
rect 8272 2278 8330 2312
rect 8364 2278 8422 2312
rect 8456 2278 8514 2312
rect 8548 2278 8606 2312
rect 8640 2278 8698 2312
rect 8732 2278 8790 2312
rect 8824 2278 8882 2312
rect 8916 2278 8974 2312
rect 9008 2278 9066 2312
rect 9100 2278 9158 2312
rect 9192 2278 9250 2312
rect 9284 2278 9342 2312
rect 9376 2278 9434 2312
rect 9468 2278 9526 2312
rect 9560 2278 9618 2312
rect 9652 2278 9710 2312
rect 9744 2278 9802 2312
rect 9836 2278 9894 2312
rect 9928 2278 9986 2312
rect 10020 2278 10078 2312
rect 10112 2278 10170 2312
rect 10204 2278 10262 2312
rect 10296 2278 10354 2312
rect 10388 2278 10446 2312
rect 10480 2278 10538 2312
rect 10572 2278 10630 2312
rect 10664 2278 10722 2312
rect 10756 2278 10814 2312
rect 10848 2278 10906 2312
rect 10940 2278 10998 2312
rect 11032 2278 11090 2312
rect 11124 2278 11182 2312
rect 11216 2278 11274 2312
rect 11308 2278 11366 2312
rect 11400 2278 11458 2312
rect 11492 2278 11550 2312
rect 11584 2278 11642 2312
rect 11676 2278 11734 2312
rect 11768 2278 11826 2312
rect 11860 2278 11918 2312
rect 11952 2278 12010 2312
rect 12044 2278 12102 2312
rect 12136 2278 12194 2312
rect 12228 2278 12286 2312
rect 12320 2278 12378 2312
rect 12412 2278 12470 2312
rect 12504 2278 12562 2312
rect 12596 2278 12654 2312
rect 12688 2278 12746 2312
rect 12780 2278 12838 2312
rect 12872 2278 12930 2312
rect 12964 2278 12993 2312
<< viali >>
rect 1068 5849 1102 5883
rect 1712 5849 1746 5883
rect 2410 5846 2444 5880
rect 3138 5850 3172 5884
rect 3519 5779 3553 5813
rect 3613 5779 3647 5813
rect 2778 5709 2812 5743
rect 3891 5718 3925 5752
rect 12931 5167 12965 5201
rect 1428 5040 1462 5074
rect 3368 5047 3402 5081
rect 3779 5043 3813 5077
rect 5757 5046 5791 5080
rect 6168 5042 6202 5076
rect 8152 5044 8186 5078
rect 8563 5040 8597 5074
rect 10543 5043 10577 5077
rect 10954 5039 10988 5073
rect 1067 4960 1101 4994
rect 3457 4960 3491 4994
rect 5305 4977 5339 5011
rect 5850 4961 5884 4995
rect 7695 4978 7729 5012
rect 8242 4960 8276 4994
rect 10086 4980 10120 5014
rect 10637 4962 10671 4996
rect 12477 4978 12511 5012
rect 3087 4849 3121 4883
rect 5476 4860 5510 4894
rect 5748 4872 5782 4906
rect 7864 4863 7898 4897
rect 8144 4861 8178 4895
rect 10261 4846 10295 4880
rect 10544 4877 10578 4911
rect 12652 4847 12686 4881
rect 12939 4877 12973 4911
rect 3452 4490 3486 4524
rect 2538 4454 2572 4488
rect 5430 4352 5464 4386
rect 5841 4356 5875 4390
rect 7822 4352 7856 4386
rect 8233 4356 8267 4390
rect 10214 4353 10248 4387
rect 10625 4357 10659 4391
rect 12575 4349 12609 4383
rect 12930 4341 12964 4375
rect 625 4284 659 4318
rect 3898 4288 3932 4322
rect 5750 4267 5784 4301
rect 6292 4290 6326 4324
rect 8147 4268 8181 4302
rect 8682 4291 8716 4325
rect 10538 4268 10572 4302
rect 11076 4288 11110 4322
rect 5845 4188 5879 4222
rect 3366 4153 3400 4187
rect 6131 4149 6165 4183
rect 8245 4175 8279 4209
rect 10633 4183 10667 4217
rect 8519 4148 8553 4182
rect 10913 4154 10947 4188
rect 3347 3486 3381 3520
rect 3162 3412 3196 3446
rect 3455 3411 3489 3445
rect 3784 3419 3818 3453
rect 5303 3412 5337 3446
rect 6200 3415 6234 3449
rect 7693 3420 7727 3454
rect 8587 3415 8621 3449
rect 10084 3416 10118 3450
rect 10990 3414 11024 3448
rect 12476 3415 12510 3449
rect 8149 3313 8183 3347
rect 10541 3314 10575 3348
rect 12931 3317 12965 3351
rect 3015 2598 3049 2632
rect 5396 2595 5430 2629
rect 7787 2599 7821 2633
rect 10176 2600 10210 2634
rect 12570 2600 12604 2634
rect 1503 2538 1537 2572
rect 3896 2543 3930 2577
rect 6290 2543 6324 2577
rect 8682 2544 8716 2578
rect 11075 2545 11109 2579
rect 12927 2549 12961 2583
rect 1059 2413 1093 2447
rect 3450 2436 3484 2470
rect 5841 2435 5875 2469
rect 8236 2438 8270 2472
rect 10625 2436 10659 2470
<< metal1 >>
rect -773 6211 -392 6343
rect 95 6218 230 6219
rect 376 6218 12090 6219
rect 95 6211 12090 6218
rect -773 6128 12090 6211
rect -773 5345 -392 6128
rect 95 6123 12090 6128
rect 220 6122 418 6123
rect 83 5947 117 5952
rect 83 5919 2907 5947
rect 83 5918 117 5919
rect 8120 5903 8173 5910
rect 1056 5883 1122 5890
rect 86 5881 120 5882
rect 1056 5881 1068 5883
rect 86 5853 1068 5881
rect 86 5848 120 5853
rect 1056 5849 1068 5853
rect 1102 5849 1122 5883
rect 1056 5838 1122 5849
rect 1690 5839 1697 5891
rect 1749 5839 1758 5891
rect 2013 5890 2079 5891
rect 2013 5838 2020 5890
rect 2072 5876 2079 5890
rect 2397 5881 2455 5886
rect 3124 5884 3184 5890
rect 2397 5880 2457 5881
rect 2397 5876 2410 5880
rect 2072 5848 2410 5876
rect 2072 5838 2079 5848
rect 2397 5846 2410 5848
rect 2444 5846 2457 5880
rect 2397 5845 2457 5846
rect 3124 5850 3138 5884
rect 3172 5881 3184 5884
rect 3172 5853 8120 5881
rect 3172 5850 3184 5853
rect 2397 5840 2455 5845
rect 3124 5840 3184 5850
rect 8172 5851 8173 5903
rect 8120 5844 8173 5851
rect 10528 5827 10581 5834
rect 88 5810 122 5816
rect 3503 5813 3566 5820
rect 3503 5810 3519 5813
rect 87 5782 3519 5810
rect 3503 5779 3519 5782
rect 3553 5779 3566 5813
rect 3503 5772 3566 5779
rect 3596 5769 3602 5821
rect 3654 5769 3660 5821
rect 3727 5787 10528 5815
rect 2766 5743 2825 5750
rect 2766 5709 2778 5743
rect 2812 5731 2825 5743
rect 3727 5741 3756 5787
rect 10580 5775 10581 5827
rect 10528 5768 10581 5775
rect 3727 5731 3755 5741
rect 2812 5709 3755 5731
rect 2766 5703 3755 5709
rect 3875 5707 3882 5759
rect 3934 5734 3941 5759
rect 5724 5734 5731 5759
rect 3934 5707 5731 5734
rect 5783 5707 5790 5759
rect 3875 5706 5790 5707
rect 446 5675 576 5676
rect 44 5665 12039 5675
rect 13338 5672 13694 5936
rect 12278 5665 13694 5672
rect 44 5638 13694 5665
rect 40 5604 13694 5638
rect 44 5596 13694 5604
rect 44 5589 13238 5596
rect 44 5580 12039 5589
rect 44 5579 450 5580
rect 504 5579 12039 5580
rect 1053 5516 1119 5517
rect 1053 5505 1060 5516
rect 1039 5477 1060 5505
rect 1053 5464 1060 5477
rect 1112 5505 1119 5516
rect 1714 5516 1780 5517
rect 1714 5505 1721 5516
rect 1112 5477 1721 5505
rect 1112 5464 1119 5477
rect 1714 5464 1721 5477
rect 1773 5505 1780 5516
rect 3444 5516 3510 5517
rect 3444 5505 3451 5516
rect 1773 5477 3451 5505
rect 1773 5464 1780 5477
rect 3444 5464 3451 5477
rect 3503 5505 3510 5516
rect 5827 5516 5893 5517
rect 5827 5505 5834 5516
rect 3503 5477 5834 5505
rect 3503 5464 3510 5477
rect 5827 5464 5834 5477
rect 5886 5505 5893 5516
rect 8222 5516 8288 5517
rect 8222 5505 8229 5516
rect 5886 5477 8229 5505
rect 5886 5464 5893 5477
rect 8222 5464 8229 5477
rect 8281 5505 8288 5516
rect 10617 5516 10683 5517
rect 10617 5505 10624 5516
rect 8281 5477 10624 5505
rect 8281 5464 8288 5477
rect 10617 5464 10624 5477
rect 10676 5505 10683 5516
rect 12913 5516 12979 5517
rect 12913 5505 12920 5516
rect 10676 5477 12920 5505
rect 10676 5464 10683 5477
rect 12913 5464 12920 5477
rect 12972 5464 12979 5516
rect 13338 5402 13694 5596
rect 36 5374 13694 5402
rect 36 5345 13030 5346
rect -773 5293 13030 5345
rect -773 5262 13031 5293
rect -773 4650 -392 5262
rect 36 5250 13031 5262
rect 12557 5215 12589 5216
rect 12557 5211 12638 5215
rect 12557 5159 12563 5211
rect 12615 5201 12638 5211
rect 12918 5201 12977 5207
rect 12615 5167 12931 5201
rect 12965 5167 12977 5201
rect 12615 5166 12977 5167
rect 12615 5159 12638 5166
rect 12918 5160 12977 5166
rect 12557 5150 12638 5159
rect 12557 5149 12589 5150
rect 1411 5074 1474 5081
rect 2015 5074 2022 5086
rect 1411 5040 1428 5074
rect 1462 5046 2022 5074
rect 1462 5040 1474 5046
rect 1411 5034 1474 5040
rect 2015 5034 2022 5046
rect 2074 5034 2081 5086
rect 3356 5081 3415 5087
rect 3356 5047 3368 5081
rect 3402 5077 3415 5081
rect 3767 5077 3826 5083
rect 3402 5049 3779 5077
rect 3402 5047 3415 5049
rect 3356 5040 3415 5047
rect 3767 5043 3779 5049
rect 3813 5043 3826 5077
rect 3767 5036 3826 5043
rect 5745 5080 5804 5086
rect 5745 5046 5757 5080
rect 5791 5076 5804 5080
rect 6156 5076 6215 5082
rect 5791 5048 6168 5076
rect 5791 5046 5804 5048
rect 5745 5039 5804 5046
rect 6156 5042 6168 5048
rect 6202 5042 6215 5076
rect 6156 5035 6215 5042
rect 8140 5078 8199 5084
rect 8140 5044 8152 5078
rect 8186 5074 8199 5078
rect 8551 5074 8610 5080
rect 8186 5046 8563 5074
rect 8186 5044 8199 5046
rect 8140 5037 8199 5044
rect 8551 5040 8563 5046
rect 8597 5040 8610 5074
rect 8551 5033 8610 5040
rect 10531 5077 10590 5083
rect 10531 5043 10543 5077
rect 10577 5073 10590 5077
rect 10942 5073 11001 5079
rect 10577 5045 10954 5073
rect 10577 5043 10590 5045
rect 10531 5036 10590 5043
rect 10942 5039 10954 5045
rect 10988 5039 11001 5073
rect 10942 5032 11001 5039
rect 1052 5003 1118 5004
rect 1052 4951 1059 5003
rect 1111 4951 1118 5003
rect 3442 5003 3508 5004
rect 3442 4951 3449 5003
rect 3501 4951 3508 5003
rect 5286 4970 5293 5022
rect 5345 4970 5351 5022
rect 7686 5021 7739 5028
rect 5835 5004 5901 5005
rect 5835 4952 5842 5004
rect 5894 4952 5901 5004
rect 7738 4969 7739 5021
rect 10077 5023 10130 5030
rect 7686 4962 7739 4969
rect 8227 5003 8293 5004
rect 8227 4951 8234 5003
rect 8286 4951 8293 5003
rect 10129 4971 10130 5023
rect 12468 5021 12521 5028
rect 10077 4964 10130 4971
rect 10622 5005 10688 5006
rect 10622 4953 10629 5005
rect 10681 4953 10688 5005
rect 12520 4969 12521 5021
rect 12468 4962 12521 4969
rect 2520 4948 2586 4949
rect 2520 4896 2527 4948
rect 2579 4896 2586 4948
rect 5576 4915 5629 4922
rect 10372 4920 10425 4927
rect 12767 4920 12820 4927
rect 5460 4904 5524 4910
rect 3070 4890 3136 4891
rect 3070 4838 3077 4890
rect 3129 4838 3136 4890
rect 5460 4852 5467 4904
rect 5519 4852 5524 4904
rect 5576 4863 5577 4915
rect 5737 4911 5798 4915
rect 5736 4906 5798 4911
rect 5629 4872 5748 4906
rect 5782 4872 5798 4906
rect 5736 4867 5798 4872
rect 5737 4864 5798 4867
rect 5576 4856 5629 4863
rect 7850 4860 7856 4912
rect 7908 4860 7914 4912
rect 7850 4852 7914 4860
rect 7972 4904 8025 4911
rect 7972 4852 7973 4904
rect 8135 4900 8196 4905
rect 8132 4895 8196 4900
rect 8025 4861 8144 4895
rect 8178 4861 8196 4895
rect 8132 4856 8196 4861
rect 8135 4854 8196 4856
rect 10252 4889 10305 4896
rect 5460 4851 5524 4852
rect 5460 4846 5523 4851
rect 7972 4845 8025 4852
rect 10304 4837 10305 4889
rect 10372 4868 10373 4920
rect 10532 4911 10593 4920
rect 10425 4877 10544 4911
rect 10578 4877 10593 4911
rect 10532 4869 10593 4877
rect 12643 4890 12696 4897
rect 10372 4861 10425 4868
rect 10252 4830 10305 4837
rect 12695 4838 12696 4890
rect 12767 4868 12768 4920
rect 12926 4911 12987 4920
rect 12820 4877 12939 4911
rect 12973 4877 12987 4911
rect 12926 4869 12987 4877
rect 12767 4861 12820 4868
rect 12643 4831 12696 4838
rect 32 4795 13027 4802
rect 13338 4795 13694 5374
rect 32 4719 13694 4795
rect 32 4706 13027 4719
rect 32 4650 13027 4657
rect -773 4567 13027 4650
rect -773 3779 -392 4567
rect 32 4561 13027 4567
rect 2527 4498 2580 4505
rect 2527 4446 2528 4498
rect 3436 4480 3442 4532
rect 3494 4480 3500 4532
rect 5833 4514 5899 4515
rect 5833 4462 5840 4514
rect 5892 4499 5899 4514
rect 8224 4514 8290 4515
rect 5892 4462 5952 4499
rect 8224 4462 8231 4514
rect 8283 4499 8290 4514
rect 10618 4505 10671 4511
rect 8283 4462 8344 4499
rect 2527 4439 2580 4446
rect 5833 4397 5886 4404
rect 5833 4396 5834 4397
rect 5417 4386 5476 4392
rect 5828 4386 5834 4396
rect 5417 4352 5430 4386
rect 5464 4358 5834 4386
rect 5464 4352 5476 4358
rect 5417 4345 5476 4352
rect 5828 4349 5834 4358
rect 5833 4345 5834 4349
rect 5886 4349 5887 4396
rect 3888 4332 3941 4339
rect 5833 4338 5886 4345
rect 617 4328 682 4329
rect 414 4319 448 4322
rect 611 4319 682 4328
rect 412 4318 682 4319
rect 412 4291 625 4318
rect 414 4288 448 4291
rect 611 4284 625 4291
rect 659 4284 682 4318
rect 611 4278 682 4284
rect 617 4277 682 4278
rect 3940 4280 3941 4332
rect 3888 4273 3941 4280
rect 5736 4307 5786 4308
rect 5736 4305 5796 4307
rect 5915 4305 5952 4462
rect 8221 4396 8274 4402
rect 8220 4395 8279 4396
rect 7809 4386 7868 4392
rect 8220 4386 8222 4395
rect 7809 4352 7822 4386
rect 7856 4358 8222 4386
rect 7856 4352 7868 4358
rect 7809 4345 7868 4352
rect 8220 4349 8222 4358
rect 8221 4343 8222 4349
rect 8274 4349 8279 4395
rect 5736 4301 5952 4305
rect 5736 4267 5750 4301
rect 5784 4268 5952 4301
rect 6283 4333 6336 4340
rect 8221 4336 8274 4343
rect 6335 4281 6336 4333
rect 6283 4274 6336 4281
rect 8133 4305 8190 4308
rect 8307 4305 8344 4462
rect 10618 4453 10619 4505
rect 10671 4462 10736 4499
rect 10618 4445 10671 4453
rect 10613 4397 10666 4403
rect 10612 4396 10671 4397
rect 10201 4387 10260 4393
rect 10612 4387 10614 4396
rect 10201 4353 10214 4387
rect 10248 4359 10614 4387
rect 10248 4353 10260 4359
rect 10201 4346 10260 4353
rect 10612 4350 10614 4359
rect 10613 4344 10614 4350
rect 10666 4350 10671 4396
rect 8133 4302 8344 4305
rect 8133 4268 8147 4302
rect 8181 4268 8344 4302
rect 8673 4334 8726 4341
rect 10613 4337 10666 4344
rect 8725 4282 8726 4334
rect 8673 4275 8726 4282
rect 10525 4305 10579 4309
rect 10699 4305 10736 4462
rect 12558 4388 12629 4396
rect 10525 4302 10736 4305
rect 10525 4268 10538 4302
rect 10572 4268 10736 4302
rect 11067 4331 11120 4338
rect 12558 4336 12566 4388
rect 12618 4336 12629 4388
rect 11119 4279 11120 4331
rect 12914 4331 12920 4383
rect 12972 4331 12978 4383
rect 12914 4330 12978 4331
rect 11067 4272 11120 4279
rect 5784 4267 5796 4268
rect 5736 4260 5796 4267
rect 8133 4255 8190 4268
rect 10525 4257 10579 4268
rect 5976 4229 6029 4236
rect 5831 4222 5893 4228
rect 3349 4194 3415 4195
rect 3349 4142 3356 4194
rect 3408 4142 3415 4194
rect 5831 4188 5845 4222
rect 5879 4221 5893 4222
rect 5879 4188 5976 4221
rect 5831 4187 5976 4188
rect 5831 4182 5893 4187
rect 6028 4177 6029 4229
rect 8227 4209 8294 4219
rect 8398 4218 8451 4225
rect 5976 4170 6029 4177
rect 6118 4183 6171 4195
rect 6118 4149 6131 4183
rect 6165 4174 6171 4183
rect 6567 4193 6633 4194
rect 6567 4174 6574 4193
rect 6165 4149 6574 4174
rect 6118 4146 6574 4149
rect 6118 4143 6171 4146
rect 6567 4141 6574 4146
rect 6626 4174 6633 4193
rect 8227 4175 8245 4209
rect 8279 4175 8398 4209
rect 6626 4146 6832 4174
rect 8227 4165 8294 4175
rect 8450 4166 8451 4218
rect 10615 4217 10682 4227
rect 10786 4226 10839 4233
rect 8959 4194 9025 4195
rect 8398 4159 8451 4166
rect 8507 4182 8565 4189
rect 8507 4148 8519 4182
rect 8553 4173 8565 4182
rect 8959 4173 8966 4194
rect 8553 4148 8966 4173
rect 6626 4141 6633 4146
rect 8507 4145 8966 4148
rect 8507 4142 8565 4145
rect 8959 4142 8966 4145
rect 9018 4173 9025 4194
rect 10615 4183 10633 4217
rect 10667 4183 10786 4217
rect 10615 4173 10682 4183
rect 10838 4174 10839 4226
rect 11348 4195 11414 4196
rect 9018 4145 9225 4173
rect 10786 4167 10839 4174
rect 10898 4188 10959 4194
rect 10898 4154 10913 4188
rect 10947 4174 10959 4188
rect 11348 4174 11355 4195
rect 10947 4154 11355 4174
rect 10898 4146 11355 4154
rect 9018 4142 9025 4145
rect 10898 4142 10959 4146
rect 11348 4143 11355 4146
rect 11407 4174 11414 4195
rect 11407 4146 11617 4174
rect 11407 4143 11414 4146
rect 93 4104 13088 4113
rect 13338 4104 13694 4719
rect 93 4028 13694 4104
rect 93 4017 13088 4028
rect 3349 3952 3415 3953
rect 1489 3941 1496 3952
rect 1484 3912 1496 3941
rect 1489 3900 1496 3912
rect 1548 3941 1555 3952
rect 3349 3941 3356 3952
rect 1548 3912 3356 3941
rect 1548 3900 1555 3912
rect 3349 3900 3356 3912
rect 3408 3941 3415 3952
rect 3881 3952 3947 3953
rect 3881 3941 3888 3952
rect 3408 3912 3888 3941
rect 3408 3900 3415 3912
rect 3881 3900 3888 3912
rect 3940 3941 3947 3952
rect 5285 3952 5351 3953
rect 5285 3941 5292 3952
rect 3940 3913 5292 3941
rect 3940 3900 3947 3913
rect 5285 3900 5292 3913
rect 5344 3941 5351 3952
rect 6270 3952 6336 3953
rect 6270 3941 6277 3952
rect 5344 3913 6277 3941
rect 5344 3900 5351 3913
rect 6270 3900 6277 3913
rect 6329 3941 6336 3952
rect 7677 3952 7743 3953
rect 7677 3941 7684 3952
rect 6329 3913 7684 3941
rect 6329 3900 6336 3913
rect 7677 3900 7684 3913
rect 7736 3941 7743 3952
rect 8660 3952 8726 3953
rect 8660 3941 8667 3952
rect 7736 3913 8667 3941
rect 7736 3900 7743 3913
rect 8660 3900 8667 3913
rect 8719 3941 8726 3952
rect 10074 3952 10140 3953
rect 10074 3941 10081 3952
rect 8719 3913 10081 3941
rect 8719 3900 8726 3913
rect 10074 3900 10081 3913
rect 10133 3941 10140 3952
rect 11050 3952 11116 3953
rect 11050 3941 11057 3952
rect 10133 3913 11057 3941
rect 10133 3900 10140 3913
rect 11050 3900 11057 3913
rect 11109 3941 11116 3952
rect 12462 3952 12528 3953
rect 12462 3941 12469 3952
rect 11109 3913 12469 3941
rect 11109 3900 11116 3913
rect 12462 3900 12469 3913
rect 12521 3941 12528 3952
rect 12521 3913 12941 3941
rect 12521 3900 12528 3913
rect 13338 3840 13694 4028
rect 113 3812 13694 3840
rect 110 3779 13105 3784
rect -773 3696 13105 3779
rect -773 2907 -392 3696
rect 110 3688 13105 3696
rect 2614 3524 2681 3525
rect 2614 3472 2622 3524
rect 2674 3499 2681 3524
rect 3060 3523 3126 3524
rect 3060 3499 3067 3523
rect 2674 3472 3067 3499
rect 2622 3471 3067 3472
rect 3119 3471 3126 3523
rect 3333 3520 3394 3527
rect 3333 3486 3347 3520
rect 3381 3515 3394 3520
rect 4181 3515 4189 3524
rect 3381 3487 4189 3515
rect 3381 3486 3394 3487
rect 3333 3480 3394 3486
rect 4181 3472 4189 3487
rect 4241 3472 4248 3524
rect 7684 3463 7737 3470
rect 2012 3451 2078 3452
rect 412 3443 446 3448
rect 2012 3443 2019 3451
rect 412 3415 2019 3443
rect 412 3414 446 3415
rect 2012 3399 2019 3415
rect 2071 3443 2078 3451
rect 3156 3446 3202 3458
rect 3156 3443 3162 3446
rect 2071 3415 3162 3443
rect 2071 3399 2078 3415
rect 3156 3412 3162 3415
rect 3196 3412 3202 3446
rect 3156 3400 3202 3412
rect 3446 3445 3495 3458
rect 3446 3411 3455 3445
rect 3489 3411 3495 3445
rect 3446 3404 3495 3411
rect 3541 3453 3837 3459
rect 3541 3420 3784 3453
rect 3453 3240 3492 3404
rect 3541 3240 3580 3420
rect 3776 3419 3784 3420
rect 3818 3419 3837 3453
rect 3776 3407 3837 3419
rect 5293 3453 5346 3460
rect 5345 3401 5346 3453
rect 6184 3405 6191 3457
rect 6243 3405 6250 3457
rect 7736 3411 7737 3463
rect 10075 3459 10128 3466
rect 7684 3404 7737 3411
rect 8571 3405 8578 3457
rect 8630 3405 8637 3457
rect 10127 3407 10128 3459
rect 12467 3458 12520 3465
rect 5293 3394 5346 3401
rect 10075 3400 10128 3407
rect 10974 3404 10981 3456
rect 11033 3404 11040 3456
rect 12519 3406 12520 3458
rect 12467 3399 12520 3406
rect 4175 3387 4239 3388
rect 4175 3335 4181 3387
rect 4233 3335 4239 3387
rect 6568 3386 6634 3387
rect 11348 3386 11414 3387
rect 6568 3334 6575 3386
rect 6627 3334 6634 3386
rect 8962 3385 9028 3386
rect 8141 3355 8194 3362
rect 8193 3303 8194 3355
rect 8962 3333 8969 3385
rect 9021 3333 9028 3385
rect 10533 3356 10586 3363
rect 8141 3296 8194 3303
rect 10585 3304 10586 3356
rect 11348 3334 11355 3386
rect 11407 3334 11414 3386
rect 12923 3359 12976 3366
rect 10533 3297 10586 3304
rect 12975 3307 12976 3359
rect 12923 3300 12976 3307
rect 89 3231 13084 3240
rect 13338 3231 13694 3812
rect 89 3155 13694 3231
rect 89 3144 13084 3155
rect 414 3066 448 3071
rect 3000 3066 3007 3077
rect 412 3038 3007 3066
rect 414 3037 448 3038
rect 3000 3025 3007 3038
rect 3059 3066 3066 3077
rect 5380 3066 5387 3078
rect 3059 3038 5387 3066
rect 3059 3025 3066 3038
rect 5380 3026 5387 3038
rect 5439 3066 5446 3078
rect 6179 3066 6186 3077
rect 5439 3038 6186 3066
rect 5439 3026 5446 3038
rect 6179 3025 6186 3038
rect 6238 3066 6245 3077
rect 7773 3066 7780 3077
rect 6238 3038 7780 3066
rect 6238 3025 6245 3038
rect 7773 3025 7780 3038
rect 7832 3066 7839 3077
rect 8568 3066 8575 3078
rect 7832 3038 8575 3066
rect 7832 3025 7839 3038
rect 8568 3026 8575 3038
rect 8627 3066 8634 3078
rect 10160 3066 10167 3077
rect 8627 3038 10167 3066
rect 8627 3026 8634 3038
rect 10160 3025 10167 3038
rect 10219 3066 10226 3077
rect 10977 3066 10984 3078
rect 10219 3038 10984 3066
rect 10219 3025 10226 3038
rect 10977 3026 10984 3038
rect 11036 3066 11043 3078
rect 12555 3066 12562 3078
rect 11036 3038 12562 3066
rect 11036 3026 11043 3038
rect 12555 3026 12562 3038
rect 12614 3066 12621 3078
rect 12614 3038 12998 3066
rect 12614 3026 12621 3038
rect 13338 2968 13694 3155
rect 179 2940 13694 2968
rect 179 2939 13058 2940
rect 217 2907 13212 2911
rect -773 2824 13212 2907
rect -773 2464 -392 2824
rect 217 2815 13212 2824
rect 2999 2588 3006 2640
rect 3058 2588 3065 2640
rect 3887 2588 3940 2595
rect 1488 2530 1498 2582
rect 1550 2530 1562 2582
rect 1488 2528 1562 2530
rect 3887 2536 3888 2588
rect 5380 2585 5387 2637
rect 5439 2585 5446 2637
rect 6281 2586 6334 2593
rect 7771 2589 7778 2641
rect 7830 2589 7837 2641
rect 3887 2529 3940 2536
rect 6333 2534 6334 2586
rect 6281 2527 6334 2534
rect 8673 2587 8726 2594
rect 10160 2590 10167 2642
rect 10219 2590 10226 2642
rect 8725 2535 8726 2587
rect 8673 2528 8726 2535
rect 11066 2588 11119 2595
rect 12554 2590 12561 2642
rect 12613 2590 12620 2642
rect 12919 2595 12971 2597
rect 12916 2591 12973 2595
rect 11118 2536 11119 2588
rect 12916 2539 12919 2591
rect 12971 2539 12973 2591
rect 12916 2536 12973 2539
rect 11066 2529 11119 2536
rect 12919 2533 12971 2536
rect 2612 2514 2678 2515
rect 2612 2462 2619 2514
rect 2671 2462 2678 2514
rect 3442 2478 3495 2485
rect 1051 2455 1104 2462
rect 1103 2403 1104 2455
rect 3494 2426 3495 2478
rect 3442 2419 3495 2426
rect 5017 2438 5051 2506
rect 5833 2477 5886 2484
rect 5460 2438 5466 2447
rect 5017 2410 5466 2438
rect 1051 2396 1104 2403
rect 5460 2395 5466 2410
rect 5518 2395 5524 2447
rect 5885 2425 5886 2477
rect 5833 2418 5886 2425
rect 7409 2438 7443 2506
rect 8228 2480 8281 2487
rect 7852 2438 7858 2447
rect 7409 2410 7858 2438
rect 7852 2395 7858 2410
rect 7910 2395 7916 2447
rect 8280 2428 8281 2480
rect 8228 2421 8281 2428
rect 9801 2438 9835 2506
rect 10617 2478 10670 2485
rect 10244 2438 10250 2447
rect 9801 2410 10250 2438
rect 10244 2395 10250 2410
rect 10302 2395 10308 2447
rect 10669 2426 10670 2478
rect 10617 2419 10670 2426
rect 12193 2438 12227 2506
rect 12635 2438 12641 2447
rect 12193 2410 12641 2438
rect 12635 2395 12641 2410
rect 12693 2395 12699 2447
rect 244 2361 13239 2367
rect 13338 2361 13694 2940
rect 244 2285 13694 2361
rect 244 2271 13239 2285
rect 13338 2260 13694 2285
<< via1 >>
rect 1697 5883 1749 5891
rect 1697 5849 1712 5883
rect 1712 5849 1746 5883
rect 1746 5849 1749 5883
rect 1697 5839 1749 5849
rect 2020 5838 2072 5890
rect 8120 5851 8172 5903
rect 3602 5813 3654 5821
rect 3602 5779 3613 5813
rect 3613 5779 3647 5813
rect 3647 5779 3654 5813
rect 3602 5769 3654 5779
rect 10528 5775 10580 5827
rect 3882 5752 3934 5759
rect 3882 5718 3891 5752
rect 3891 5718 3925 5752
rect 3925 5718 3934 5752
rect 3882 5707 3934 5718
rect 5731 5707 5783 5759
rect 1060 5464 1112 5516
rect 1721 5464 1773 5516
rect 3451 5464 3503 5516
rect 5834 5464 5886 5516
rect 8229 5464 8281 5516
rect 10624 5464 10676 5516
rect 12920 5464 12972 5516
rect 12563 5159 12615 5211
rect 2022 5034 2074 5086
rect 1059 4994 1111 5003
rect 1059 4960 1067 4994
rect 1067 4960 1101 4994
rect 1101 4960 1111 4994
rect 1059 4951 1111 4960
rect 3449 4994 3501 5003
rect 3449 4960 3457 4994
rect 3457 4960 3491 4994
rect 3491 4960 3501 4994
rect 3449 4951 3501 4960
rect 5293 5011 5345 5022
rect 5293 4977 5305 5011
rect 5305 4977 5339 5011
rect 5339 4977 5345 5011
rect 5293 4970 5345 4977
rect 7686 5012 7738 5021
rect 5842 4995 5894 5004
rect 5842 4961 5850 4995
rect 5850 4961 5884 4995
rect 5884 4961 5894 4995
rect 5842 4952 5894 4961
rect 7686 4978 7695 5012
rect 7695 4978 7729 5012
rect 7729 4978 7738 5012
rect 7686 4969 7738 4978
rect 10077 5014 10129 5023
rect 8234 4994 8286 5003
rect 8234 4960 8242 4994
rect 8242 4960 8276 4994
rect 8276 4960 8286 4994
rect 8234 4951 8286 4960
rect 10077 4980 10086 5014
rect 10086 4980 10120 5014
rect 10120 4980 10129 5014
rect 10077 4971 10129 4980
rect 12468 5012 12520 5021
rect 10629 4996 10681 5005
rect 10629 4962 10637 4996
rect 10637 4962 10671 4996
rect 10671 4962 10681 4996
rect 10629 4953 10681 4962
rect 12468 4978 12477 5012
rect 12477 4978 12511 5012
rect 12511 4978 12520 5012
rect 12468 4969 12520 4978
rect 2527 4896 2579 4948
rect 3077 4883 3129 4890
rect 3077 4849 3087 4883
rect 3087 4849 3121 4883
rect 3121 4849 3129 4883
rect 3077 4838 3129 4849
rect 5467 4894 5519 4904
rect 5467 4860 5476 4894
rect 5476 4860 5510 4894
rect 5510 4860 5519 4894
rect 5467 4852 5519 4860
rect 5577 4863 5629 4915
rect 7856 4897 7908 4912
rect 7856 4863 7864 4897
rect 7864 4863 7898 4897
rect 7898 4863 7908 4897
rect 7856 4860 7908 4863
rect 7973 4852 8025 4904
rect 10252 4880 10304 4889
rect 10252 4846 10261 4880
rect 10261 4846 10295 4880
rect 10295 4846 10304 4880
rect 10252 4837 10304 4846
rect 10373 4868 10425 4920
rect 12643 4881 12695 4890
rect 12643 4847 12652 4881
rect 12652 4847 12686 4881
rect 12686 4847 12695 4881
rect 12643 4838 12695 4847
rect 12768 4868 12820 4920
rect 2528 4488 2580 4498
rect 2528 4454 2538 4488
rect 2538 4454 2572 4488
rect 2572 4454 2580 4488
rect 3442 4524 3494 4532
rect 3442 4490 3452 4524
rect 3452 4490 3486 4524
rect 3486 4490 3494 4524
rect 3442 4480 3494 4490
rect 5840 4462 5892 4514
rect 8231 4462 8283 4514
rect 2528 4446 2580 4454
rect 5834 4390 5886 4397
rect 5834 4356 5841 4390
rect 5841 4356 5875 4390
rect 5875 4356 5886 4390
rect 5834 4345 5886 4356
rect 3888 4322 3940 4332
rect 3888 4288 3898 4322
rect 3898 4288 3932 4322
rect 3932 4288 3940 4322
rect 3888 4280 3940 4288
rect 8222 4390 8274 4395
rect 8222 4356 8233 4390
rect 8233 4356 8267 4390
rect 8267 4356 8274 4390
rect 8222 4343 8274 4356
rect 6283 4324 6335 4333
rect 6283 4290 6292 4324
rect 6292 4290 6326 4324
rect 6326 4290 6335 4324
rect 6283 4281 6335 4290
rect 10619 4453 10671 4505
rect 10614 4391 10666 4396
rect 10614 4357 10625 4391
rect 10625 4357 10659 4391
rect 10659 4357 10666 4391
rect 10614 4344 10666 4357
rect 8673 4325 8725 4334
rect 8673 4291 8682 4325
rect 8682 4291 8716 4325
rect 8716 4291 8725 4325
rect 8673 4282 8725 4291
rect 12566 4383 12618 4388
rect 12566 4349 12575 4383
rect 12575 4349 12609 4383
rect 12609 4349 12618 4383
rect 12566 4336 12618 4349
rect 11067 4322 11119 4331
rect 11067 4288 11076 4322
rect 11076 4288 11110 4322
rect 11110 4288 11119 4322
rect 11067 4279 11119 4288
rect 12920 4375 12972 4383
rect 12920 4341 12930 4375
rect 12930 4341 12964 4375
rect 12964 4341 12972 4375
rect 12920 4331 12972 4341
rect 3356 4187 3408 4194
rect 3356 4153 3366 4187
rect 3366 4153 3400 4187
rect 3400 4153 3408 4187
rect 3356 4142 3408 4153
rect 5976 4177 6028 4229
rect 6574 4141 6626 4193
rect 8398 4166 8450 4218
rect 8966 4142 9018 4194
rect 10786 4174 10838 4226
rect 11355 4143 11407 4195
rect 1496 3900 1548 3952
rect 3356 3900 3408 3952
rect 3888 3900 3940 3952
rect 5292 3900 5344 3952
rect 6277 3900 6329 3952
rect 7684 3900 7736 3952
rect 8667 3900 8719 3952
rect 10081 3900 10133 3952
rect 11057 3900 11109 3952
rect 12469 3900 12521 3952
rect 2622 3472 2674 3524
rect 3067 3471 3119 3523
rect 4189 3472 4241 3524
rect 2019 3399 2071 3451
rect 5293 3446 5345 3453
rect 5293 3412 5303 3446
rect 5303 3412 5337 3446
rect 5337 3412 5345 3446
rect 5293 3401 5345 3412
rect 6191 3449 6243 3457
rect 6191 3415 6200 3449
rect 6200 3415 6234 3449
rect 6234 3415 6243 3449
rect 6191 3405 6243 3415
rect 7684 3454 7736 3463
rect 7684 3420 7693 3454
rect 7693 3420 7727 3454
rect 7727 3420 7736 3454
rect 7684 3411 7736 3420
rect 8578 3449 8630 3457
rect 8578 3415 8587 3449
rect 8587 3415 8621 3449
rect 8621 3415 8630 3449
rect 8578 3405 8630 3415
rect 10075 3450 10127 3459
rect 10075 3416 10084 3450
rect 10084 3416 10118 3450
rect 10118 3416 10127 3450
rect 10075 3407 10127 3416
rect 10981 3448 11033 3456
rect 10981 3414 10990 3448
rect 10990 3414 11024 3448
rect 11024 3414 11033 3448
rect 10981 3404 11033 3414
rect 12467 3449 12519 3458
rect 12467 3415 12476 3449
rect 12476 3415 12510 3449
rect 12510 3415 12519 3449
rect 12467 3406 12519 3415
rect 4181 3335 4233 3387
rect 6575 3334 6627 3386
rect 8141 3347 8193 3355
rect 8141 3313 8149 3347
rect 8149 3313 8183 3347
rect 8183 3313 8193 3347
rect 8141 3303 8193 3313
rect 8969 3333 9021 3385
rect 10533 3348 10585 3356
rect 10533 3314 10541 3348
rect 10541 3314 10575 3348
rect 10575 3314 10585 3348
rect 10533 3304 10585 3314
rect 11355 3334 11407 3386
rect 12923 3351 12975 3359
rect 12923 3317 12931 3351
rect 12931 3317 12965 3351
rect 12965 3317 12975 3351
rect 12923 3307 12975 3317
rect 3007 3025 3059 3077
rect 5387 3026 5439 3078
rect 6186 3025 6238 3077
rect 7780 3025 7832 3077
rect 8575 3026 8627 3078
rect 10167 3025 10219 3077
rect 10984 3026 11036 3078
rect 12562 3026 12614 3078
rect 3006 2632 3058 2640
rect 3006 2598 3015 2632
rect 3015 2598 3049 2632
rect 3049 2598 3058 2632
rect 3006 2588 3058 2598
rect 1498 2572 1550 2582
rect 1498 2538 1503 2572
rect 1503 2538 1537 2572
rect 1537 2538 1550 2572
rect 1498 2530 1550 2538
rect 3888 2577 3940 2588
rect 5387 2629 5439 2637
rect 5387 2595 5396 2629
rect 5396 2595 5430 2629
rect 5430 2595 5439 2629
rect 5387 2585 5439 2595
rect 7778 2633 7830 2641
rect 7778 2599 7787 2633
rect 7787 2599 7821 2633
rect 7821 2599 7830 2633
rect 7778 2589 7830 2599
rect 3888 2543 3896 2577
rect 3896 2543 3930 2577
rect 3930 2543 3940 2577
rect 3888 2536 3940 2543
rect 6281 2577 6333 2586
rect 6281 2543 6290 2577
rect 6290 2543 6324 2577
rect 6324 2543 6333 2577
rect 6281 2534 6333 2543
rect 10167 2634 10219 2642
rect 10167 2600 10176 2634
rect 10176 2600 10210 2634
rect 10210 2600 10219 2634
rect 10167 2590 10219 2600
rect 8673 2578 8725 2587
rect 8673 2544 8682 2578
rect 8682 2544 8716 2578
rect 8716 2544 8725 2578
rect 8673 2535 8725 2544
rect 12561 2634 12613 2642
rect 12561 2600 12570 2634
rect 12570 2600 12604 2634
rect 12604 2600 12613 2634
rect 12561 2590 12613 2600
rect 11066 2579 11118 2588
rect 11066 2545 11075 2579
rect 11075 2545 11109 2579
rect 11109 2545 11118 2579
rect 11066 2536 11118 2545
rect 12919 2583 12971 2591
rect 12919 2549 12927 2583
rect 12927 2549 12961 2583
rect 12961 2549 12971 2583
rect 12919 2539 12971 2549
rect 2619 2462 2671 2514
rect 3442 2470 3494 2478
rect 1051 2447 1103 2455
rect 1051 2413 1059 2447
rect 1059 2413 1093 2447
rect 1093 2413 1103 2447
rect 1051 2403 1103 2413
rect 3442 2436 3450 2470
rect 3450 2436 3484 2470
rect 3484 2436 3494 2470
rect 3442 2426 3494 2436
rect 5833 2469 5885 2477
rect 5466 2395 5518 2447
rect 5833 2435 5841 2469
rect 5841 2435 5875 2469
rect 5875 2435 5885 2469
rect 5833 2425 5885 2435
rect 8228 2472 8280 2480
rect 7858 2395 7910 2447
rect 8228 2438 8236 2472
rect 8236 2438 8270 2472
rect 8270 2438 8280 2472
rect 8228 2428 8280 2438
rect 10617 2470 10669 2478
rect 10250 2395 10302 2447
rect 10617 2436 10625 2470
rect 10625 2436 10659 2470
rect 10659 2436 10669 2470
rect 10617 2426 10669 2436
rect 12641 2395 12693 2447
<< metal2 >>
rect 8120 5903 8173 5910
rect 1690 5839 1697 5891
rect 1749 5839 1758 5891
rect 1730 5517 1758 5839
rect 2013 5890 2079 5891
rect 2013 5838 2020 5890
rect 2072 5838 2079 5890
rect 8172 5851 8173 5903
rect 8120 5844 8173 5851
rect 1053 5516 1119 5517
rect 1053 5464 1060 5516
rect 1112 5464 1119 5516
rect 1714 5516 1780 5517
rect 1714 5464 1721 5516
rect 1773 5464 1780 5516
rect 1071 5029 1099 5464
rect 2032 5086 2060 5838
rect 3596 5769 3602 5821
rect 3654 5769 3660 5821
rect 3444 5516 3510 5517
rect 3444 5464 3451 5516
rect 3503 5464 3510 5516
rect 2015 5034 2022 5086
rect 2074 5034 2081 5086
rect 1070 5004 1099 5029
rect 1052 5003 1118 5004
rect 1052 4951 1059 5003
rect 1111 4951 1118 5003
rect 1489 3900 1496 3952
rect 1548 3900 1555 3952
rect 1508 2582 1536 3900
rect 2032 3452 2060 5034
rect 3464 5004 3492 5464
rect 3442 5003 3508 5004
rect 3442 4951 3449 5003
rect 3501 4951 3508 5003
rect 2520 4948 2586 4949
rect 2520 4896 2527 4948
rect 2579 4896 2586 4948
rect 2535 4505 2568 4896
rect 3070 4890 3136 4891
rect 3070 4838 3077 4890
rect 3129 4838 3136 4890
rect 2527 4498 2580 4505
rect 2527 4446 2528 4498
rect 2527 4439 2580 4446
rect 2616 3525 2681 3526
rect 2615 3524 2681 3525
rect 3094 3524 3122 4838
rect 3436 4480 3442 4532
rect 3494 4525 3500 4532
rect 3608 4525 3641 5769
rect 3875 5707 3882 5759
rect 3934 5707 3941 5759
rect 5724 5707 5731 5759
rect 5783 5707 5790 5759
rect 3875 5706 3941 5707
rect 5286 4970 5293 5022
rect 5345 4970 5351 5022
rect 3494 4490 3641 4525
rect 3494 4480 3500 4490
rect 3888 4332 3941 4339
rect 3940 4280 3941 4332
rect 3888 4273 3941 4280
rect 3349 4194 3415 4195
rect 3349 4142 3356 4194
rect 3408 4142 3415 4194
rect 3369 3953 3397 4142
rect 3900 3953 3928 4273
rect 5305 3953 5333 4970
rect 5576 4915 5629 4922
rect 5460 4904 5524 4910
rect 5460 4852 5467 4904
rect 5519 4852 5524 4904
rect 5576 4863 5577 4915
rect 5576 4856 5629 4863
rect 5460 4851 5524 4852
rect 5460 4846 5523 4851
rect 3349 3952 3415 3953
rect 3349 3900 3356 3952
rect 3408 3900 3415 3952
rect 3881 3952 3947 3953
rect 3881 3900 3888 3952
rect 3940 3900 3947 3952
rect 5285 3952 5351 3953
rect 5285 3900 5292 3952
rect 5344 3900 5351 3952
rect 2615 3472 2622 3524
rect 2674 3472 2681 3524
rect 3060 3523 3126 3524
rect 2012 3451 2078 3452
rect 2012 3399 2019 3451
rect 2071 3399 2078 3451
rect 1488 2530 1498 2582
rect 1550 2530 1562 2582
rect 1488 2528 1562 2530
rect 2629 2515 2657 3472
rect 3060 3471 3067 3523
rect 3119 3471 3126 3523
rect 3000 3025 3007 3077
rect 3059 3025 3066 3077
rect 3020 2640 3048 3025
rect 2999 2588 3006 2640
rect 3058 2588 3065 2640
rect 3900 2595 3928 3900
rect 4181 3472 4189 3524
rect 4241 3472 4248 3524
rect 4194 3388 4222 3472
rect 5305 3460 5333 3900
rect 5293 3453 5346 3460
rect 5345 3401 5346 3453
rect 5293 3394 5346 3401
rect 4175 3387 4239 3388
rect 4175 3335 4181 3387
rect 4233 3335 4239 3387
rect 5380 3026 5387 3078
rect 5439 3026 5446 3078
rect 5400 2637 5428 3026
rect 3887 2588 3940 2595
rect 3887 2536 3888 2588
rect 5380 2585 5387 2637
rect 5439 2585 5446 2637
rect 3887 2529 3940 2536
rect 2612 2514 2678 2515
rect 2612 2462 2619 2514
rect 2671 2462 2678 2514
rect 3442 2478 3495 2485
rect 1051 2455 1104 2462
rect 1103 2403 1104 2455
rect 3494 2426 3495 2478
rect 5476 2447 5509 4846
rect 3442 2419 3495 2426
rect 1051 2396 1104 2403
rect 1063 1784 1091 2396
rect 3454 1784 3482 2419
rect 5460 2395 5466 2447
rect 5518 2395 5524 2447
rect 5476 2392 5509 2395
rect 1058 1750 1092 1784
rect 3450 1750 3484 1784
rect 5589 1782 5617 4856
rect 5739 4390 5772 5707
rect 5827 5516 5893 5517
rect 5827 5464 5834 5516
rect 5886 5464 5893 5516
rect 5847 5005 5875 5464
rect 7686 5021 7739 5028
rect 5835 5004 5901 5005
rect 5835 4952 5842 5004
rect 5894 4952 5901 5004
rect 7738 4969 7739 5021
rect 7686 4962 7739 4969
rect 5847 4515 5875 4952
rect 5833 4514 5899 4515
rect 5833 4462 5840 4514
rect 5892 4462 5899 4514
rect 5833 4397 5886 4404
rect 5833 4390 5834 4397
rect 5739 4356 5834 4390
rect 5833 4345 5834 4356
rect 5833 4338 5886 4345
rect 6283 4333 6336 4340
rect 6335 4281 6336 4333
rect 6283 4274 6336 4281
rect 5976 4229 6029 4236
rect 6028 4177 6029 4229
rect 5976 4170 6029 4177
rect 5833 2477 5886 2484
rect 5885 2425 5886 2477
rect 5833 2418 5886 2425
rect 5845 1782 5873 2418
rect 1063 1748 1091 1750
rect 3454 1748 3482 1750
rect 5586 1748 5620 1782
rect 5844 1748 5878 1782
rect 5988 1779 6016 4170
rect 6292 3953 6320 4274
rect 6567 4193 6633 4194
rect 6567 4141 6574 4193
rect 6626 4141 6633 4193
rect 6270 3952 6336 3953
rect 6270 3900 6277 3952
rect 6329 3900 6336 3952
rect 6184 3405 6191 3457
rect 6243 3405 6250 3457
rect 6197 3077 6225 3405
rect 6179 3025 6186 3077
rect 6238 3025 6245 3077
rect 6292 2593 6320 3900
rect 6584 3387 6612 4141
rect 7697 3953 7725 4962
rect 7850 4860 7856 4912
rect 7908 4860 7914 4912
rect 7850 4852 7914 4860
rect 7972 4904 8025 4911
rect 7972 4852 7973 4904
rect 7677 3952 7743 3953
rect 7677 3900 7684 3952
rect 7736 3900 7743 3952
rect 7697 3470 7725 3900
rect 7684 3463 7737 3470
rect 7736 3411 7737 3463
rect 7684 3404 7737 3411
rect 6568 3386 6634 3387
rect 6568 3334 6575 3386
rect 6627 3334 6634 3386
rect 7773 3025 7780 3077
rect 7832 3025 7839 3077
rect 7793 2641 7821 3025
rect 6281 2586 6334 2593
rect 7771 2589 7778 2641
rect 7830 2589 7837 2641
rect 6333 2534 6334 2586
rect 6281 2527 6334 2534
rect 7867 2447 7900 4852
rect 7972 4845 8025 4852
rect 7852 2395 7858 2447
rect 7910 2395 7916 2447
rect 7985 1784 8013 4845
rect 8129 4390 8162 5844
rect 10528 5827 10581 5834
rect 10580 5775 10581 5827
rect 10528 5768 10581 5775
rect 8222 5516 8288 5517
rect 8222 5464 8229 5516
rect 8281 5464 8288 5516
rect 8242 5004 8270 5464
rect 10077 5023 10130 5030
rect 8227 5003 8293 5004
rect 8227 4951 8234 5003
rect 8286 4951 8293 5003
rect 10129 4971 10130 5023
rect 10077 4964 10130 4971
rect 8242 4515 8270 4951
rect 8224 4514 8290 4515
rect 8224 4462 8231 4514
rect 8283 4462 8290 4514
rect 8221 4395 8274 4402
rect 8221 4390 8222 4395
rect 8129 4356 8222 4390
rect 8130 4355 8222 4356
rect 8221 4343 8222 4355
rect 8221 4336 8274 4343
rect 8673 4334 8726 4341
rect 8725 4282 8726 4334
rect 8673 4275 8726 4282
rect 8398 4218 8451 4225
rect 8450 4166 8451 4218
rect 8398 4159 8451 4166
rect 8141 3355 8194 3362
rect 8193 3303 8194 3355
rect 8141 3296 8194 3303
rect 8153 1898 8181 3296
rect 8228 2480 8281 2487
rect 8280 2428 8281 2480
rect 8228 2421 8281 2428
rect 8151 1864 8185 1898
rect 5986 1745 6020 1779
rect 7982 1750 8016 1784
rect 7985 1748 8013 1750
rect 8153 1748 8181 1864
rect 8240 1844 8268 2421
rect 8238 1810 8272 1844
rect 8240 1748 8268 1810
rect 8410 1779 8438 4159
rect 8684 3953 8712 4275
rect 8959 4194 9025 4195
rect 8959 4142 8966 4194
rect 9018 4142 9025 4194
rect 8660 3952 8726 3953
rect 8660 3900 8667 3952
rect 8719 3900 8726 3952
rect 8571 3405 8578 3457
rect 8630 3405 8637 3457
rect 8586 3078 8614 3405
rect 8568 3026 8575 3078
rect 8627 3026 8634 3078
rect 8684 2594 8712 3900
rect 8977 3386 9005 4142
rect 10089 3953 10117 4964
rect 10372 4920 10425 4927
rect 10252 4889 10305 4896
rect 10304 4837 10305 4889
rect 10372 4868 10373 4920
rect 10372 4861 10425 4868
rect 10252 4830 10305 4837
rect 10074 3952 10140 3953
rect 10074 3900 10081 3952
rect 10133 3900 10140 3952
rect 10089 3466 10117 3900
rect 10075 3459 10128 3466
rect 10127 3407 10128 3459
rect 10075 3400 10128 3407
rect 8962 3385 9028 3386
rect 8962 3333 8969 3385
rect 9021 3333 9028 3385
rect 10160 3025 10167 3077
rect 10219 3025 10226 3077
rect 10180 2642 10208 3025
rect 8673 2587 8726 2594
rect 10160 2590 10167 2642
rect 10219 2590 10226 2642
rect 8725 2535 8726 2587
rect 8673 2528 8726 2535
rect 10259 2447 10292 4830
rect 10244 2395 10250 2447
rect 10302 2395 10308 2447
rect 10385 1779 10413 4861
rect 10537 4391 10570 5768
rect 10617 5516 10683 5517
rect 10617 5464 10624 5516
rect 10676 5464 10683 5516
rect 12913 5516 12979 5517
rect 12913 5464 12920 5516
rect 12972 5464 12979 5516
rect 10637 5006 10665 5464
rect 12557 5211 12622 5216
rect 12557 5159 12563 5211
rect 12615 5159 12622 5211
rect 12557 5149 12622 5159
rect 12468 5021 12521 5028
rect 10622 5005 10688 5006
rect 10622 4953 10629 5005
rect 10681 4953 10688 5005
rect 12520 4969 12521 5021
rect 12468 4962 12521 4969
rect 10637 4511 10665 4953
rect 10618 4505 10671 4511
rect 10618 4453 10619 4505
rect 10618 4445 10671 4453
rect 10613 4396 10666 4403
rect 10613 4391 10614 4396
rect 10537 4357 10614 4391
rect 10613 4344 10614 4357
rect 10613 4337 10666 4344
rect 11067 4331 11120 4338
rect 11119 4279 11120 4331
rect 11067 4272 11120 4279
rect 10786 4226 10839 4233
rect 10838 4174 10839 4226
rect 10786 4167 10839 4174
rect 10533 3356 10586 3363
rect 10585 3304 10586 3356
rect 10533 3297 10586 3304
rect 10545 1870 10573 3297
rect 10617 2478 10670 2485
rect 10669 2426 10670 2478
rect 10617 2419 10670 2426
rect 10629 1870 10657 2419
rect 10544 1836 10578 1870
rect 10627 1836 10661 1870
rect 8406 1745 8440 1779
rect 10382 1745 10416 1779
rect 10545 1748 10573 1836
rect 10629 1748 10657 1836
rect 10798 1782 10826 4167
rect 11076 3953 11104 4272
rect 11348 4195 11414 4196
rect 11348 4143 11355 4195
rect 11407 4143 11414 4195
rect 11050 3952 11116 3953
rect 11050 3900 11057 3952
rect 11109 3900 11116 3952
rect 10974 3404 10981 3456
rect 11033 3404 11040 3456
rect 10995 3078 11023 3404
rect 10977 3026 10984 3078
rect 11036 3026 11043 3078
rect 11076 2595 11104 3900
rect 11369 3387 11397 4143
rect 12481 3953 12509 4962
rect 12575 4388 12608 5149
rect 12933 5148 12961 5464
rect 12767 4920 12820 4927
rect 12643 4890 12696 4897
rect 12695 4838 12696 4890
rect 12767 4868 12768 4920
rect 12767 4861 12820 4868
rect 12643 4831 12696 4838
rect 12560 4336 12566 4388
rect 12618 4336 12624 4388
rect 12462 3952 12528 3953
rect 12462 3900 12469 3952
rect 12521 3900 12528 3952
rect 12481 3465 12509 3900
rect 12467 3458 12520 3465
rect 12519 3406 12520 3458
rect 12467 3399 12520 3406
rect 11348 3386 11414 3387
rect 11348 3334 11355 3386
rect 11407 3334 11414 3386
rect 12555 3026 12562 3078
rect 12614 3026 12621 3078
rect 12575 2642 12603 3026
rect 11066 2588 11119 2595
rect 12554 2590 12561 2642
rect 12613 2590 12620 2642
rect 11118 2536 11119 2588
rect 11066 2529 11119 2536
rect 12652 2447 12685 4831
rect 12635 2395 12641 2447
rect 12693 2395 12699 2447
rect 10795 1748 10829 1782
rect 12780 1779 12808 4861
rect 12932 4383 12965 5148
rect 12914 4331 12920 4383
rect 12972 4331 12978 4383
rect 12914 4330 12978 4331
rect 12923 3359 12976 3366
rect 12975 3307 12976 3359
rect 12923 3300 12976 3307
rect 12935 2597 12963 3300
rect 12919 2591 12971 2597
rect 12919 2533 12971 2539
rect 12935 1854 12963 2533
rect 12932 1820 12966 1854
rect 12776 1745 12810 1779
rect 12935 1748 12963 1820
use sky130_fd_sc_hd__mux4_4  sky130_fd_sc_hd__mux4_4_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform -1 0 4135 0 1 5627
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_1  x1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1697295826
transform 1 0 594 0 1 4065
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  x2
timestamp 1697295826
transform 1 0 1035 0 1 5627
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  x3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1697295826
transform 1 0 870 0 1 4065
box -38 -48 590 592
use sky130_fd_sc_hd__buf_16  x4 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 1402 0 1 4065
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_2  x5 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 1311 0 1 5627
box -38 -48 406 592
use sky130_fd_sc_hd__dfbbp_1  x20 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1697358018
transform 1 0 1034 0 1 4754
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbp_1  x27
timestamp 1697358018
transform 1 0 3426 0 1 4754
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbp_1  x30
timestamp 1697358018
transform 1 0 5818 0 1 4754
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbp_1  x33
timestamp 1697358018
transform 1 0 8210 0 1 4754
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbp_1  x36
timestamp 1697358018
transform 1 0 10602 0 1 4754
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbp_1  x39
timestamp 1697358018
transform -1 0 12994 0 1 4065
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbp_1  x42
timestamp 1697358018
transform -1 0 10602 0 1 4065
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbp_1  x45
timestamp 1697358018
transform -1 0 8210 0 1 4065
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbp_1  x48
timestamp 1697358018
transform -1 0 5818 0 1 4065
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbp_1  x51
timestamp 1697358018
transform -1 0 3425 0 1 2319
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbp_1  x54
timestamp 1697358018
transform -1 0 5817 0 1 2319
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbp_1  x57
timestamp 1697358018
transform -1 0 8209 0 1 2319
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbp_1  x60
timestamp 1697358018
transform -1 0 10601 0 1 2319
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbp_1  x63
timestamp 1697358018
transform -1 0 12993 0 1 2319
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbp_1  x66
timestamp 1697358018
transform 1 0 10601 0 1 3192
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbp_1  x69
timestamp 1697358018
transform 1 0 8209 0 1 3192
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbp_1  x72
timestamp 1697358018
transform 1 0 5817 0 1 3192
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbp_1  x75
timestamp 1697358018
transform 1 0 3425 0 1 3192
box -38 -48 2430 592
use sky130_fd_sc_hd__inv_1  x77 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1697965495
transform 1 0 3168 0 1 3192
box -38 -48 314 592
<< labels >>
flabel metal1 86 5848 120 5882 0 FreeSans 480 0 0 0 clk_sar
port 45 nsew
flabel metal1 88 5782 122 5816 0 FreeSans 480 0 0 0 sel_bit[1]
port 5 nsew
flabel metal1 83 5918 117 5952 0 FreeSans 480 0 0 0 sel_bit[0]
port 4 nsew
flabel metal2 1058 1750 1092 1784 0 FreeSans 480 0 0 0 D[7]
port 9 nsew
flabel metal2 3450 1750 3484 1784 0 FreeSans 480 0 0 0 D[6]
port 10 nsew
flabel metal2 5844 1748 5878 1782 0 FreeSans 480 0 0 0 D[5]
port 12 nsew
flabel metal2 7982 1750 8016 1784 0 FreeSans 480 0 0 0 check[5]
port 14 nsew
flabel metal2 8406 1745 8440 1779 0 FreeSans 480 0 0 0 check[1]
port 15 nsew
flabel metal2 10382 1745 10416 1779 0 FreeSans 480 0 0 0 check[4]
port 16 nsew
flabel metal2 10795 1748 10829 1782 0 FreeSans 480 0 0 0 check[2]
port 17 nsew
flabel metal2 12776 1745 12810 1779 0 FreeSans 480 0 0 0 check[3]
port 18 nsew
flabel metal2 10627 1836 10661 1870 0 FreeSans 480 0 0 0 D[3]
port 20 nsew
flabel metal2 10544 1836 10578 1870 0 FreeSans 480 0 0 0 D[1]
port 21 nsew
flabel metal1 414 4288 448 4322 0 FreeSans 480 0 0 0 reset
port 6 nsew
flabel metal2 5586 1748 5620 1782 0 FreeSans 480 0 0 0 check[6]
port 11 nsew
flabel metal2 8238 1810 8272 1844 0 FreeSans 480 0 0 0 D[4]
port 22 nsew
flabel metal2 8151 1864 8185 1898 0 FreeSans 480 0 0 0 D[0]
port 24 nsew
flabel metal2 12932 1820 12966 1854 0 FreeSans 480 0 0 0 D[2]
port 19 nsew
flabel metal1 412 3414 446 3448 0 FreeSans 480 0 0 0 eob
port 7 nsew
flabel metal2 5986 1745 6020 1779 0 FreeSans 480 0 0 0 check[0]
port 13 nsew
flabel metal1 414 3037 448 3071 0 FreeSans 480 0 0 0 comparator_out
port 8 nsew
flabel metal1 100 6154 134 6188 0 FreeSans 480 0 0 0 VDD
port 47 nsew
flabel metal1 40 5604 74 5638 0 FreeSans 480 0 0 0 VSS
port 49 nsew
<< end >>
