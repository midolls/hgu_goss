magic
tech sky130A
magscale 1 2
timestamp 1700722492
<< nwell >>
rect -3292 7457 -3185 7829
rect -3397 6176 -3134 6839
<< metal1 >>
rect -8566 13488 -8560 13540
rect -8508 13538 -8502 13540
rect -8508 13491 -8447 13538
rect -8508 13488 -8502 13491
rect -6358 9031 -6352 9083
rect -6300 9031 -6294 9083
rect -950 8781 -944 8791
rect -6199 8751 -944 8781
rect -950 8739 -944 8751
rect -892 8781 -886 8791
rect -892 8751 -877 8781
rect -892 8739 -886 8751
rect -1043 8711 -1037 8721
rect -6199 8681 -1037 8711
rect -1043 8669 -1037 8681
rect -985 8711 -979 8721
rect -985 8681 -877 8711
rect -985 8669 -979 8681
rect -1505 8641 -1499 8653
rect -6199 8611 -1499 8641
rect -1505 8601 -1499 8611
rect -1447 8641 -1441 8653
rect -1447 8611 -877 8641
rect -1447 8601 -1441 8611
rect -1783 8572 -1777 8583
rect -2377 8571 -1777 8572
rect -6199 8541 -1777 8571
rect -1783 8531 -1777 8541
rect -1725 8572 -1719 8583
rect -1725 8571 -1087 8572
rect -1725 8541 -877 8571
rect -1725 8531 -1719 8541
rect -1633 8502 -1627 8513
rect -6199 8472 -1627 8502
rect -1633 8461 -1627 8472
rect -1575 8502 -1569 8513
rect -1575 8472 -877 8502
rect -1575 8461 -1569 8472
rect -2297 8432 -2291 8443
rect -6199 8402 -2291 8432
rect -2297 8391 -2291 8402
rect -2239 8432 -2233 8443
rect -2239 8402 -877 8432
rect -2239 8391 -2233 8402
rect -1225 8363 -1219 8373
rect -6199 8333 -1219 8363
rect -1225 8321 -1219 8333
rect -1167 8363 -1161 8373
rect -1167 8333 -877 8363
rect -1167 8321 -1161 8333
rect -3234 8293 -3228 8304
rect -6199 8263 -3228 8293
rect -3234 8252 -3228 8263
rect -3176 8293 -3170 8304
rect -3176 8263 -877 8293
rect -3176 8252 -3170 8263
rect -3321 8223 -3315 8233
rect -6199 8193 -3315 8223
rect -3321 8181 -3315 8193
rect -3263 8223 -3257 8233
rect -3263 8193 -877 8223
rect -3263 8181 -3257 8193
rect -3683 8153 -3677 8165
rect -6199 8123 -3677 8153
rect -3683 8113 -3677 8123
rect -3625 8153 -3619 8165
rect -3625 8123 -877 8153
rect -3625 8113 -3619 8123
rect -3961 8084 -3955 8095
rect -6199 8054 -3955 8084
rect -3961 8043 -3955 8054
rect -3903 8084 -3897 8095
rect -3903 8054 -877 8084
rect -3903 8043 -3897 8054
rect -3811 8014 -3805 8025
rect -6199 7984 -3805 8014
rect -3811 7973 -3805 7984
rect -3753 8014 -3747 8025
rect -3753 7984 -877 8014
rect -3753 7973 -3747 7984
rect -4475 7944 -4469 7955
rect -6199 7914 -4469 7944
rect -4475 7903 -4469 7914
rect -4417 7944 -4411 7955
rect -4417 7914 -877 7944
rect -4417 7903 -4411 7914
rect -3408 7875 -3402 7885
rect -6199 7845 -3402 7875
rect -3408 7833 -3402 7845
rect -3350 7875 -3344 7885
rect -3350 7845 -877 7875
rect -3350 7833 -3344 7845
rect -8565 7651 -8559 7703
rect -8507 7689 -8501 7703
rect -3334 7691 -3158 7787
rect -8507 7661 -5970 7689
rect -8507 7651 -8501 7661
rect -5998 5599 -5970 7661
rect -3447 7051 -3150 7243
rect -3443 6411 -3146 6603
rect -3421 5867 -3160 5963
rect -5397 5658 -5391 5674
rect -5422 5623 -5391 5658
rect -5397 5622 -5391 5623
rect -5339 5658 -5333 5674
rect -5339 5623 164 5658
rect -5339 5622 -5333 5623
rect -6011 5547 -6005 5599
rect -5953 5547 -5947 5599
rect -1314 5465 -1308 5517
rect -1256 5506 -1250 5517
rect -1128 5506 -1122 5516
rect -1256 5476 -1122 5506
rect -1256 5465 -1250 5476
rect -1128 5464 -1122 5476
rect -1070 5464 -1064 5516
rect -1589 5396 -1583 5448
rect -1531 5436 -1525 5448
rect -1214 5436 -1208 5446
rect -1531 5406 -1208 5436
rect -1531 5396 -1525 5406
rect -1214 5394 -1208 5406
rect -1156 5394 -1150 5446
rect -1864 5326 -1858 5378
rect -1806 5366 -1800 5378
rect -1301 5366 -1295 5377
rect -1806 5336 -1295 5366
rect -1806 5326 -1800 5336
rect -1301 5325 -1295 5336
rect -1243 5325 -1237 5377
rect -2406 5256 -2400 5308
rect -2348 5297 -2342 5308
rect -1387 5297 -1381 5307
rect -2348 5267 -1381 5297
rect -2348 5256 -2342 5267
rect -1387 5255 -1381 5267
rect -1329 5255 -1323 5307
rect -2971 5187 -2965 5239
rect -2913 5227 -2907 5239
rect -1474 5227 -1468 5238
rect -2913 5197 -1468 5227
rect -2913 5187 -2907 5197
rect -1474 5186 -1468 5197
rect -1416 5186 -1410 5238
rect -3235 5117 -3229 5169
rect -3177 5158 -3171 5169
rect -1560 5158 -1554 5168
rect -3177 5128 -1554 5158
rect -3177 5117 -3171 5128
rect -1560 5116 -1554 5128
rect -1502 5116 -1496 5168
rect -3323 5047 -3317 5099
rect -3265 5088 -3259 5099
rect -1646 5088 -1640 5098
rect -3265 5058 -1640 5088
rect -3265 5047 -3259 5058
rect -1646 5046 -1640 5058
rect -1588 5046 -1582 5098
rect -3497 4977 -3491 5029
rect -3439 5018 -3433 5029
rect -1732 5018 -1726 5028
rect -3439 4988 -1726 5018
rect -3439 4977 -3433 4988
rect -1732 4976 -1726 4988
rect -1674 4976 -1668 5028
rect -3770 4908 -3764 4960
rect -3712 4948 -3706 4960
rect -1819 4948 -1813 4959
rect -3712 4918 -1813 4948
rect -3712 4908 -3706 4918
rect -1819 4907 -1813 4918
rect -1761 4907 -1755 4959
rect -4049 4838 -4043 4890
rect -3991 4879 -3985 4890
rect -1905 4879 -1899 4889
rect -3991 4849 -1899 4879
rect -3991 4838 -3985 4849
rect -1905 4837 -1899 4849
rect -1847 4837 -1841 4889
rect -4596 4769 -4590 4821
rect -4538 4809 -4532 4821
rect -1991 4809 -1985 4819
rect -4538 4779 -1985 4809
rect -4538 4769 -4532 4779
rect -1991 4767 -1985 4779
rect -1933 4767 -1927 4819
rect -5147 4699 -5141 4751
rect -5089 4739 -5083 4751
rect -2078 4739 -2072 4750
rect -5089 4709 -2072 4739
rect -5089 4699 -5083 4709
rect -2078 4698 -2072 4709
rect -2020 4698 -2014 4750
rect -1352 -153 -1346 -101
rect -1294 -111 -1288 -101
rect -1294 -141 14484 -111
rect -1294 -153 -1288 -141
rect -804 -223 -798 -171
rect -746 -181 -740 -171
rect -746 -211 14484 -181
rect -746 -223 -740 -211
rect -537 -292 -531 -240
rect -479 -251 -473 -240
rect -479 -281 14484 -251
rect -479 -292 -473 -281
rect -251 -362 -245 -310
rect -193 -320 -187 -310
rect -193 -350 14484 -320
rect -193 -362 -187 -350
rect -24 -431 -18 -379
rect 34 -390 40 -379
rect 34 -420 14484 -390
rect 34 -431 40 -420
rect 112 -501 118 -449
rect 170 -459 176 -449
rect 170 -489 14484 -459
rect 170 -501 176 -489
rect 448 -571 454 -519
rect 506 -529 512 -519
rect 506 -559 14484 -529
rect 506 -571 512 -559
rect 994 -641 1000 -589
rect 1052 -599 1058 -589
rect 1052 -629 14484 -599
rect 1052 -641 1058 -629
rect 1541 -710 1547 -658
rect 1599 -669 1605 -658
rect 1599 -699 14484 -669
rect 1599 -710 1605 -699
rect 1827 -780 1833 -728
rect 1885 -738 1891 -728
rect 1885 -768 14484 -738
rect 1885 -780 1891 -768
rect 2093 -850 2099 -798
rect 2151 -808 2157 -798
rect 2151 -838 14484 -808
rect 2151 -850 2157 -838
rect 2338 -919 2344 -867
rect 2396 -878 2402 -867
rect 2396 -908 14484 -878
rect 2396 -919 2402 -908
rect 2476 -988 2482 -936
rect 2534 -947 2540 -936
rect 2534 -977 14484 -947
rect 2534 -988 2540 -977
rect -164 -3047 -158 -3035
rect -2409 -3077 -158 -3047
rect -164 -3087 -158 -3077
rect -106 -3047 -100 -3035
rect -106 -3077 2642 -3047
rect -106 -3087 -100 -3077
rect -1236 -3116 -1230 -3105
rect -2409 -3146 -1230 -3116
rect -1236 -3157 -1230 -3146
rect -1178 -3116 -1172 -3105
rect -1178 -3146 2642 -3116
rect -1178 -3157 -1172 -3146
rect -572 -3186 -566 -3175
rect -2409 -3216 -566 -3186
rect -572 -3227 -566 -3216
rect -514 -3186 -508 -3175
rect -514 -3216 2642 -3186
rect -514 -3227 -508 -3216
rect -722 -3256 -716 -3245
rect -2409 -3286 -716 -3256
rect -722 -3297 -716 -3286
rect -664 -3256 -658 -3245
rect -664 -3286 2642 -3256
rect -664 -3297 -658 -3286
rect -444 -3325 -438 -3315
rect -2409 -3355 -438 -3325
rect -444 -3367 -438 -3355
rect -386 -3325 -380 -3315
rect -386 -3355 2642 -3325
rect -386 -3367 -380 -3355
rect -22 -3395 -16 -3383
rect -2409 -3425 -16 -3395
rect -22 -3435 -16 -3425
rect 36 -3395 42 -3383
rect 36 -3425 2642 -3395
rect 36 -3435 42 -3425
rect 112 -3465 118 -3453
rect -2409 -3495 118 -3465
rect 112 -3505 118 -3495
rect 170 -3465 176 -3453
rect 170 -3495 2642 -3465
rect 170 -3505 176 -3495
rect 2190 -3535 2196 -3523
rect -2409 -3565 2196 -3535
rect 2190 -3575 2196 -3565
rect 2248 -3535 2254 -3523
rect 2248 -3565 2642 -3535
rect 2248 -3575 2254 -3565
rect 1118 -3604 1124 -3593
rect -2409 -3634 1124 -3604
rect 1118 -3645 1124 -3634
rect 1176 -3604 1182 -3593
rect 1176 -3634 2642 -3604
rect 1176 -3645 1182 -3634
rect 1782 -3674 1788 -3663
rect -2409 -3704 1788 -3674
rect 1782 -3715 1788 -3704
rect 1840 -3674 1846 -3663
rect 1840 -3704 2642 -3674
rect 1840 -3715 1846 -3704
rect 1632 -3743 1638 -3733
rect -2409 -3773 1638 -3743
rect 1038 -3774 1638 -3773
rect 1632 -3785 1638 -3774
rect 1690 -3743 1696 -3733
rect 1690 -3773 2642 -3743
rect 1690 -3774 2328 -3773
rect 1690 -3785 1696 -3774
rect 1910 -3813 1916 -3803
rect -2409 -3843 1916 -3813
rect 1910 -3855 1916 -3843
rect 1968 -3813 1974 -3803
rect 1968 -3843 2642 -3813
rect 1968 -3855 1974 -3843
rect 2337 -3883 2343 -3871
rect -2409 -3913 2343 -3883
rect 2337 -3923 2343 -3913
rect 2395 -3883 2401 -3871
rect 2395 -3913 2642 -3883
rect 2395 -3923 2401 -3913
rect 2481 -3953 2487 -3941
rect -2410 -3983 2487 -3953
rect 2481 -3993 2487 -3983
rect 2539 -3953 2545 -3941
rect 2539 -3983 2641 -3953
rect 2539 -3993 2545 -3983
<< via1 >>
rect -8560 13488 -8508 13540
rect -6352 9031 -6300 9083
rect -944 8739 -892 8791
rect -1037 8669 -985 8721
rect -1499 8601 -1447 8653
rect -1777 8531 -1725 8583
rect -1627 8461 -1575 8513
rect -2291 8391 -2239 8443
rect -1219 8321 -1167 8373
rect -3228 8252 -3176 8304
rect -3315 8181 -3263 8233
rect -3677 8113 -3625 8165
rect -3955 8043 -3903 8095
rect -3805 7973 -3753 8025
rect -4469 7903 -4417 7955
rect -3402 7833 -3350 7885
rect -8559 7651 -8507 7703
rect -5391 5622 -5339 5674
rect -6005 5547 -5953 5599
rect -1308 5465 -1256 5517
rect -1122 5464 -1070 5516
rect -1583 5396 -1531 5448
rect -1208 5394 -1156 5446
rect -1858 5326 -1806 5378
rect -1295 5325 -1243 5377
rect -2400 5256 -2348 5308
rect -1381 5255 -1329 5307
rect -2965 5187 -2913 5239
rect -1468 5186 -1416 5238
rect -3229 5117 -3177 5169
rect -1554 5116 -1502 5168
rect -3317 5047 -3265 5099
rect -1640 5046 -1588 5098
rect -3491 4977 -3439 5029
rect -1726 4976 -1674 5028
rect -3764 4908 -3712 4960
rect -1813 4907 -1761 4959
rect -4043 4838 -3991 4890
rect -1899 4837 -1847 4889
rect -4590 4769 -4538 4821
rect -1985 4767 -1933 4819
rect -5141 4699 -5089 4751
rect -2072 4698 -2020 4750
rect -1346 -153 -1294 -101
rect -798 -223 -746 -171
rect -531 -292 -479 -240
rect -245 -362 -193 -310
rect -18 -431 34 -379
rect 118 -501 170 -449
rect 454 -571 506 -519
rect 1000 -641 1052 -589
rect 1547 -710 1599 -658
rect 1833 -780 1885 -728
rect 2099 -850 2151 -798
rect 2344 -919 2396 -867
rect 2482 -988 2534 -936
rect -158 -3087 -106 -3035
rect -1230 -3157 -1178 -3105
rect -566 -3227 -514 -3175
rect -716 -3297 -664 -3245
rect -438 -3367 -386 -3315
rect -16 -3435 36 -3383
rect 118 -3505 170 -3453
rect 2196 -3575 2248 -3523
rect 1124 -3645 1176 -3593
rect 1788 -3715 1840 -3663
rect 1638 -3785 1690 -3733
rect 1916 -3855 1968 -3803
rect 2343 -3923 2395 -3871
rect 2487 -3993 2539 -3941
<< metal2 >>
rect -8566 13488 -8560 13540
rect -8508 13488 -8502 13540
rect -8552 7703 -8524 13488
rect -6358 9031 -6352 9083
rect -6300 9031 -6294 9083
rect -8565 7651 -8559 7703
rect -8507 7651 -8501 7703
rect -6338 7614 -6310 9031
rect -950 8739 -944 8791
rect -892 8739 -886 8791
rect -1043 8669 -1037 8721
rect -985 8669 -979 8721
rect -1505 8601 -1499 8653
rect -1447 8601 -1441 8653
rect -1783 8531 -1777 8583
rect -1725 8531 -1719 8583
rect -2297 8391 -2291 8443
rect -2239 8391 -2233 8443
rect -3234 8252 -3228 8304
rect -3176 8252 -3170 8304
rect -3321 8181 -3315 8233
rect -3263 8181 -3257 8233
rect -3683 8113 -3677 8165
rect -3625 8113 -3619 8165
rect -3961 8043 -3955 8095
rect -3903 8043 -3897 8095
rect -4475 7903 -4469 7955
rect -4417 7903 -4411 7955
rect -4464 7819 -4423 7903
rect -3945 7819 -3904 8043
rect -3811 7973 -3805 8025
rect -3753 7973 -3747 8025
rect -3801 7819 -3760 7973
rect -3669 7819 -3628 8113
rect -3408 7833 -3402 7885
rect -3350 7833 -3344 7885
rect -3391 7819 -3350 7833
rect -5397 5622 -5391 5674
rect -5339 5622 -5333 5674
rect -6011 5547 -6005 5599
rect -5953 5547 -5947 5599
rect -5135 4751 -5093 5833
rect -4586 4821 -4544 5828
rect -4038 4890 -3996 5830
rect -3758 4960 -3716 5831
rect -3486 5029 -3444 5827
rect -3312 5099 -3270 8181
rect -3223 5169 -3181 8252
rect -2286 7819 -2245 8391
rect -1767 7819 -1726 8531
rect -1633 8461 -1627 8513
rect -1575 8461 -1569 8513
rect -1623 7819 -1582 8461
rect -1491 7819 -1450 8601
rect -1225 8321 -1219 8373
rect -1167 8321 -1161 8373
rect -1213 7819 -1172 8321
rect -2959 5239 -2917 5824
rect -2395 5308 -2353 5829
rect -1852 5378 -1810 5832
rect -1578 5448 -1536 5832
rect -1303 5517 -1261 5840
rect -1314 5465 -1308 5517
rect -1256 5465 -1250 5517
rect -1128 5464 -1122 5516
rect -1070 5464 -1064 5516
rect -1589 5396 -1583 5448
rect -1531 5396 -1525 5448
rect -1214 5394 -1208 5446
rect -1156 5394 -1150 5446
rect -1864 5326 -1858 5378
rect -1806 5326 -1800 5378
rect -1301 5325 -1295 5377
rect -1243 5325 -1237 5377
rect -2406 5256 -2400 5308
rect -2348 5256 -2342 5308
rect -1387 5255 -1381 5307
rect -1329 5255 -1323 5307
rect -2971 5187 -2965 5239
rect -2913 5187 -2907 5239
rect -1474 5186 -1468 5238
rect -1416 5186 -1410 5238
rect -3235 5117 -3229 5169
rect -3177 5117 -3171 5169
rect -1560 5116 -1554 5168
rect -1502 5116 -1496 5168
rect -3323 5047 -3317 5099
rect -3265 5047 -3259 5099
rect -1646 5046 -1640 5098
rect -1588 5046 -1582 5098
rect -3497 4977 -3491 5029
rect -3439 4977 -3433 5029
rect -1732 4976 -1726 5028
rect -1674 4976 -1668 5028
rect -3770 4908 -3764 4960
rect -3712 4908 -3706 4960
rect -1819 4907 -1813 4959
rect -1761 4907 -1755 4959
rect -4049 4838 -4043 4890
rect -3991 4838 -3985 4890
rect -1905 4837 -1899 4889
rect -1847 4837 -1841 4889
rect -4596 4769 -4590 4821
rect -4538 4769 -4532 4821
rect -1991 4767 -1985 4819
rect -1933 4767 -1927 4819
rect -5147 4699 -5141 4751
rect -5089 4699 -5083 4751
rect -2078 4698 -2072 4750
rect -2020 4698 -2014 4750
rect -2062 4590 -2020 4698
rect -1980 4590 -1938 4767
rect -1896 4590 -1854 4837
rect -1808 4590 -1766 4907
rect -1721 4590 -1679 4976
rect -1635 4590 -1593 5046
rect -1549 4590 -1507 5116
rect -1462 4590 -1420 5186
rect -1376 4590 -1334 5255
rect -1290 4590 -1248 5325
rect -1203 4590 -1161 5394
rect -1118 4590 -1076 5464
rect -1031 4591 -989 8669
rect -944 4591 -902 8739
rect -1352 -153 -1346 -101
rect -1294 -153 -1288 -101
rect -1902 -987 -1860 -219
rect -1340 -1032 -1298 -153
rect -804 -223 -798 -171
rect -746 -223 -740 -171
rect -794 -1032 -752 -223
rect -537 -292 -531 -240
rect -479 -292 -473 -240
rect -526 -1032 -484 -292
rect -251 -362 -245 -310
rect -193 -362 -187 -310
rect -239 -1032 -197 -362
rect -24 -431 -18 -379
rect 34 -431 40 -379
rect -1225 -3105 -1184 -2843
rect -1236 -3157 -1230 -3105
rect -1178 -3157 -1172 -3105
rect -706 -3245 -665 -2963
rect -562 -3175 -521 -2916
rect -572 -3227 -566 -3175
rect -514 -3227 -508 -3175
rect -722 -3297 -716 -3245
rect -664 -3297 -658 -3245
rect -430 -3315 -389 -3028
rect -164 -3087 -158 -3035
rect -106 -3087 -100 -3035
rect -444 -3367 -438 -3315
rect -386 -3367 -380 -3315
rect -13 -3383 29 -431
rect 112 -501 118 -449
rect 170 -501 176 -449
rect -22 -3435 -16 -3383
rect 36 -3435 42 -3383
rect 123 -3453 165 -501
rect 448 -571 454 -519
rect 506 -571 512 -519
rect 460 -1032 502 -571
rect 994 -641 1000 -589
rect 1052 -641 1058 -589
rect 1006 -1032 1048 -641
rect 1541 -710 1547 -658
rect 1599 -710 1605 -658
rect 1552 -1032 1594 -710
rect 1827 -780 1833 -728
rect 1885 -780 1891 -728
rect 1839 -1032 1881 -780
rect 2093 -850 2099 -798
rect 2151 -850 2157 -798
rect 2104 -1032 2146 -850
rect 2338 -919 2344 -867
rect 2396 -919 2402 -867
rect 112 -3505 118 -3453
rect 170 -3505 176 -3453
rect 1129 -3593 1170 -2750
rect 1118 -3645 1124 -3593
rect 1176 -3645 1182 -3593
rect 1648 -3733 1689 -2891
rect 1792 -3663 1833 -2805
rect 1782 -3715 1788 -3663
rect 1840 -3715 1846 -3663
rect 1632 -3785 1638 -3733
rect 1690 -3785 1696 -3733
rect 1924 -3803 1965 -2945
rect 2202 -3523 2243 -3017
rect 2190 -3575 2196 -3523
rect 2248 -3575 2254 -3523
rect 1910 -3855 1916 -3803
rect 1968 -3855 1974 -3803
rect 2349 -3871 2391 -919
rect 2476 -988 2482 -936
rect 2534 -988 2540 -936
rect 2337 -3923 2343 -3871
rect 2395 -3923 2401 -3871
rect 2487 -3941 2529 -988
rect 2481 -3993 2487 -3941
rect 2539 -3993 2545 -3941
<< metal4 >>
rect -5346 9209 -4382 9215
rect -5756 9030 -4382 9209
rect -5756 8938 -5568 9030
rect -5378 9028 -4382 9030
rect -5378 8938 -5174 9028
rect -5756 8936 -5174 8938
rect -4984 9026 -4382 9028
rect -4984 8936 -4767 9026
rect -5756 8934 -4767 8936
rect -4577 8934 -4382 9026
rect -5756 7770 -4382 8934
rect -3171 9018 -2207 9177
rect -3171 8926 -3042 9018
rect -2852 9014 -2207 9018
rect -2852 8926 -2616 9014
rect -3171 8922 -2616 8926
rect -2426 8922 -2207 9014
rect -5756 7764 -4792 7770
rect -5756 5870 -5344 7764
rect -3171 7733 -2207 8922
rect -6144 4549 -5862 5189
rect -4300 4549 -3323 5974
rect -1171 5863 -699 7792
rect -6144 4255 -2585 4549
rect -6144 4251 -5862 4255
use hgu_cdac_half  hgu_cdac_half_0
timestamp 1700485439
transform 1 0 -49110 0 -1 6793
box -459 -645 39606 6456
use hgu_cdac_half  hgu_cdac_half_1
timestamp 1700485439
transform 1 0 -49110 0 1 8403
box -459 -645 39606 6456
use hgu_cdac_sw_buffer  hgu_cdac_sw_buffer_0
timestamp 1699539897
transform -1 0 -315 0 -1 -3772
box -270 -2798 1830 -714
use hgu_cdac_sw_buffer  hgu_cdac_sw_buffer_1
timestamp 1699539897
transform -1 0 2039 0 -1 -3768
box -270 -2798 1830 -714
use hgu_cdac_sw_buffer  hgu_cdac_sw_buffer_2
timestamp 1699539897
transform -1 0 -1376 0 1 8596
box -270 -2798 1830 -714
use hgu_cdac_sw_buffer  hgu_cdac_sw_buffer_3
timestamp 1699539897
transform -1 0 -3554 0 1 8595
box -270 -2798 1830 -714
use hgu_comp_flat  hgu_comp_flat_0
timestamp 1698719859
transform 1 0 -9082 0 1 7042
box 338 -1940 3788 618
use hgu_sarlogic_flat  hgu_sarlogic_flat_0
timestamp 1700302578
transform 1 0 -10778 0 1 1681
box 2064 -1908 31250 13749
use hgu_tah  hgu_tah_0
timestamp 1699832401
transform 1 0 -51671 0 1 3641
box 711 297 1858 5355
use hgu_vgen_vref  hgu_vgen_vref_0
timestamp 1700722492
transform -1 0 -50750 0 1 -30367
box 0 0 22370 76000
<< end >>
