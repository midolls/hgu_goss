magic
tech sky130A
magscale 1 2
timestamp 1699537245
<< nwell >>
rect 12283 10064 18880 10661
rect 12234 10063 18880 10064
rect 11754 9696 18880 10063
rect 12283 9634 18880 9696
rect 12283 9367 18878 9634
rect 12928 9301 13146 9367
rect 13660 9304 14004 9367
rect 14872 9304 15216 9367
rect 16084 9304 16428 9367
rect 17296 9304 17640 9367
rect 18070 9319 18878 9367
rect 18070 9318 18289 9319
rect 13332 6641 18192 7303
rect 13332 5361 18192 6023
<< pwell >>
rect 11834 9456 12020 9638
rect 12024 9456 12210 9638
rect 11834 9452 11855 9456
rect 11821 9418 11855 9452
rect 12189 9452 12210 9456
rect 12189 9418 12223 9452
rect 18570 9215 18839 9261
rect 18473 9079 18839 9215
rect 18501 9041 18535 9079
rect 13400 7543 13434 7581
rect 15792 7543 15826 7581
rect 13371 7407 15761 7543
rect 15763 7407 18153 7543
rect 14152 7363 14606 7407
rect 14927 7363 15761 7407
rect 16544 7363 16998 7407
rect 17319 7363 18153 7407
rect 15294 7361 15761 7363
rect 17686 7361 18153 7363
rect 15294 6581 15761 6583
rect 17686 6581 18153 6583
rect 14152 6537 14606 6581
rect 14927 6537 15761 6581
rect 16544 6537 16998 6581
rect 17319 6537 18153 6581
rect 13371 6401 15761 6537
rect 15763 6401 18153 6537
rect 13400 6363 13434 6401
rect 15792 6363 15826 6401
rect 13400 6263 13434 6301
rect 15792 6263 15826 6301
rect 13371 6127 15761 6263
rect 15763 6127 18153 6263
rect 14152 6083 14606 6127
rect 14927 6083 15761 6127
rect 16544 6083 16998 6127
rect 17319 6083 18153 6127
rect 15294 6081 15761 6083
rect 17686 6081 18153 6083
rect 15294 5301 15761 5303
rect 17686 5301 18153 5303
rect 14152 5257 14606 5301
rect 14927 5257 15761 5301
rect 16544 5257 16998 5301
rect 17319 5257 18153 5301
rect 13371 5121 15761 5257
rect 15763 5121 18153 5257
rect 13400 5083 13434 5121
rect 15792 5083 15826 5121
<< nmos >>
rect 13375 9152 13405 9236
rect 14107 9152 14137 9236
rect 14229 9152 14259 9236
rect 15319 9152 15349 9236
rect 15441 9152 15471 9236
rect 16657 9152 16687 9236
rect 16779 9152 16809 9236
rect 17513 9152 17543 9236
rect 18165 9153 18195 9237
rect 18257 9153 18287 9237
rect 18353 9153 18383 9237
rect 12355 8968 12385 9052
rect 12427 8968 12457 9052
rect 18165 9015 18195 9099
rect 12355 8830 12385 8914
rect 12427 8830 12457 8914
rect 12355 8692 12385 8776
rect 12427 8692 12457 8776
rect 12355 8554 12385 8638
rect 12427 8554 12457 8638
rect 12355 8416 12385 8500
rect 12427 8416 12457 8500
rect 12355 8278 12385 8362
rect 12427 8278 12457 8362
rect 12355 8140 12385 8224
rect 12427 8140 12457 8224
rect 12355 8002 12385 8086
rect 12427 8002 12457 8086
<< scnmos >>
rect 11912 9482 11942 9612
rect 12102 9482 12132 9612
rect 18551 9105 18581 9189
rect 18646 9105 18676 9235
rect 18730 9105 18760 9235
rect 13449 7433 13479 7517
rect 13533 7433 13563 7517
rect 13721 7433 13751 7517
rect 13816 7445 13846 7517
rect 13922 7445 13952 7517
rect 14018 7433 14048 7517
rect 14128 7433 14158 7517
rect 14228 7389 14258 7517
rect 14312 7389 14342 7517
rect 14500 7389 14530 7517
rect 14595 7445 14625 7517
rect 14704 7445 14734 7517
rect 14799 7433 14829 7517
rect 14885 7433 14915 7517
rect 15003 7389 15033 7517
rect 15087 7389 15117 7517
rect 15275 7433 15305 7517
rect 15370 7387 15400 7517
rect 15558 7433 15588 7517
rect 15653 7387 15683 7517
rect 15841 7433 15871 7517
rect 15925 7433 15955 7517
rect 16113 7433 16143 7517
rect 16208 7445 16238 7517
rect 16314 7445 16344 7517
rect 16410 7433 16440 7517
rect 16520 7433 16550 7517
rect 16620 7389 16650 7517
rect 16704 7389 16734 7517
rect 16892 7389 16922 7517
rect 16987 7445 17017 7517
rect 17096 7445 17126 7517
rect 17191 7433 17221 7517
rect 17277 7433 17307 7517
rect 17395 7389 17425 7517
rect 17479 7389 17509 7517
rect 17667 7433 17697 7517
rect 17762 7387 17792 7517
rect 17950 7433 17980 7517
rect 18045 7387 18075 7517
rect 13449 6427 13479 6511
rect 13533 6427 13563 6511
rect 13721 6427 13751 6511
rect 13816 6427 13846 6499
rect 13922 6427 13952 6499
rect 14018 6427 14048 6511
rect 14128 6427 14158 6511
rect 14228 6427 14258 6555
rect 14312 6427 14342 6555
rect 14500 6427 14530 6555
rect 14595 6427 14625 6499
rect 14704 6427 14734 6499
rect 14799 6427 14829 6511
rect 14885 6427 14915 6511
rect 15003 6427 15033 6555
rect 15087 6427 15117 6555
rect 15275 6427 15305 6511
rect 15370 6427 15400 6557
rect 15558 6427 15588 6511
rect 15653 6427 15683 6557
rect 15841 6427 15871 6511
rect 15925 6427 15955 6511
rect 16113 6427 16143 6511
rect 16208 6427 16238 6499
rect 16314 6427 16344 6499
rect 16410 6427 16440 6511
rect 16520 6427 16550 6511
rect 16620 6427 16650 6555
rect 16704 6427 16734 6555
rect 16892 6427 16922 6555
rect 16987 6427 17017 6499
rect 17096 6427 17126 6499
rect 17191 6427 17221 6511
rect 17277 6427 17307 6511
rect 17395 6427 17425 6555
rect 17479 6427 17509 6555
rect 17667 6427 17697 6511
rect 17762 6427 17792 6557
rect 17950 6427 17980 6511
rect 18045 6427 18075 6557
rect 13449 6153 13479 6237
rect 13533 6153 13563 6237
rect 13721 6153 13751 6237
rect 13816 6165 13846 6237
rect 13922 6165 13952 6237
rect 14018 6153 14048 6237
rect 14128 6153 14158 6237
rect 14228 6109 14258 6237
rect 14312 6109 14342 6237
rect 14500 6109 14530 6237
rect 14595 6165 14625 6237
rect 14704 6165 14734 6237
rect 14799 6153 14829 6237
rect 14885 6153 14915 6237
rect 15003 6109 15033 6237
rect 15087 6109 15117 6237
rect 15275 6153 15305 6237
rect 15370 6107 15400 6237
rect 15558 6153 15588 6237
rect 15653 6107 15683 6237
rect 15841 6153 15871 6237
rect 15925 6153 15955 6237
rect 16113 6153 16143 6237
rect 16208 6165 16238 6237
rect 16314 6165 16344 6237
rect 16410 6153 16440 6237
rect 16520 6153 16550 6237
rect 16620 6109 16650 6237
rect 16704 6109 16734 6237
rect 16892 6109 16922 6237
rect 16987 6165 17017 6237
rect 17096 6165 17126 6237
rect 17191 6153 17221 6237
rect 17277 6153 17307 6237
rect 17395 6109 17425 6237
rect 17479 6109 17509 6237
rect 17667 6153 17697 6237
rect 17762 6107 17792 6237
rect 17950 6153 17980 6237
rect 18045 6107 18075 6237
rect 13449 5147 13479 5231
rect 13533 5147 13563 5231
rect 13721 5147 13751 5231
rect 13816 5147 13846 5219
rect 13922 5147 13952 5219
rect 14018 5147 14048 5231
rect 14128 5147 14158 5231
rect 14228 5147 14258 5275
rect 14312 5147 14342 5275
rect 14500 5147 14530 5275
rect 14595 5147 14625 5219
rect 14704 5147 14734 5219
rect 14799 5147 14829 5231
rect 14885 5147 14915 5231
rect 15003 5147 15033 5275
rect 15087 5147 15117 5275
rect 15275 5147 15305 5231
rect 15370 5147 15400 5277
rect 15558 5147 15588 5231
rect 15653 5147 15683 5277
rect 15841 5147 15871 5231
rect 15925 5147 15955 5231
rect 16113 5147 16143 5231
rect 16208 5147 16238 5219
rect 16314 5147 16344 5219
rect 16410 5147 16440 5231
rect 16520 5147 16550 5231
rect 16620 5147 16650 5275
rect 16704 5147 16734 5275
rect 16892 5147 16922 5275
rect 16987 5147 17017 5219
rect 17096 5147 17126 5219
rect 17191 5147 17221 5231
rect 17277 5147 17307 5231
rect 17395 5147 17425 5275
rect 17479 5147 17509 5275
rect 17667 5147 17697 5231
rect 17762 5147 17792 5277
rect 17950 5147 17980 5231
rect 18045 5147 18075 5277
<< pmos >>
rect 13022 9350 13052 9434
rect 13754 9353 13784 9437
rect 13880 9353 13910 9437
rect 14966 9353 14996 9437
rect 15092 9353 15122 9437
rect 16178 9353 16208 9437
rect 16304 9353 16334 9437
rect 17390 9353 17420 9437
rect 17516 9353 17546 9437
<< scpmoshvt >>
rect 11912 9732 11942 9932
rect 12102 9732 12132 9932
rect 18551 9419 18581 9547
rect 18646 9355 18676 9555
rect 18730 9355 18760 9555
rect 13449 7073 13479 7201
rect 13533 7073 13563 7201
rect 13721 7067 13751 7151
rect 13814 7067 13844 7151
rect 13898 7067 13928 7151
rect 14018 7067 14048 7151
rect 14124 7067 14154 7151
rect 14232 7067 14262 7235
rect 14316 7067 14346 7235
rect 14453 7067 14483 7235
rect 14597 7067 14627 7151
rect 14681 7067 14711 7151
rect 14799 7067 14829 7151
rect 14907 7067 14937 7151
rect 15003 7067 15033 7235
rect 15075 7067 15105 7235
rect 15273 7135 15303 7263
rect 15370 7067 15400 7267
rect 15558 7083 15588 7211
rect 15653 7067 15683 7267
rect 15841 7073 15871 7201
rect 15925 7073 15955 7201
rect 16113 7067 16143 7151
rect 16206 7067 16236 7151
rect 16290 7067 16320 7151
rect 16410 7067 16440 7151
rect 16516 7067 16546 7151
rect 16624 7067 16654 7235
rect 16708 7067 16738 7235
rect 16845 7067 16875 7235
rect 16989 7067 17019 7151
rect 17073 7067 17103 7151
rect 17191 7067 17221 7151
rect 17299 7067 17329 7151
rect 17395 7067 17425 7235
rect 17467 7067 17497 7235
rect 17665 7135 17695 7263
rect 17762 7067 17792 7267
rect 17950 7083 17980 7211
rect 18045 7067 18075 7267
rect 13449 6743 13479 6871
rect 13533 6743 13563 6871
rect 13721 6793 13751 6877
rect 13814 6793 13844 6877
rect 13898 6793 13928 6877
rect 14018 6793 14048 6877
rect 14124 6793 14154 6877
rect 14232 6709 14262 6877
rect 14316 6709 14346 6877
rect 14453 6709 14483 6877
rect 14597 6793 14627 6877
rect 14681 6793 14711 6877
rect 14799 6793 14829 6877
rect 14907 6793 14937 6877
rect 15003 6709 15033 6877
rect 15075 6709 15105 6877
rect 15273 6681 15303 6809
rect 15370 6677 15400 6877
rect 15558 6733 15588 6861
rect 15653 6677 15683 6877
rect 15841 6743 15871 6871
rect 15925 6743 15955 6871
rect 16113 6793 16143 6877
rect 16206 6793 16236 6877
rect 16290 6793 16320 6877
rect 16410 6793 16440 6877
rect 16516 6793 16546 6877
rect 16624 6709 16654 6877
rect 16708 6709 16738 6877
rect 16845 6709 16875 6877
rect 16989 6793 17019 6877
rect 17073 6793 17103 6877
rect 17191 6793 17221 6877
rect 17299 6793 17329 6877
rect 17395 6709 17425 6877
rect 17467 6709 17497 6877
rect 17665 6681 17695 6809
rect 17762 6677 17792 6877
rect 17950 6733 17980 6861
rect 18045 6677 18075 6877
rect 13449 5793 13479 5921
rect 13533 5793 13563 5921
rect 13721 5787 13751 5871
rect 13814 5787 13844 5871
rect 13898 5787 13928 5871
rect 14018 5787 14048 5871
rect 14124 5787 14154 5871
rect 14232 5787 14262 5955
rect 14316 5787 14346 5955
rect 14453 5787 14483 5955
rect 14597 5787 14627 5871
rect 14681 5787 14711 5871
rect 14799 5787 14829 5871
rect 14907 5787 14937 5871
rect 15003 5787 15033 5955
rect 15075 5787 15105 5955
rect 15273 5855 15303 5983
rect 15370 5787 15400 5987
rect 15558 5803 15588 5931
rect 15653 5787 15683 5987
rect 15841 5793 15871 5921
rect 15925 5793 15955 5921
rect 16113 5787 16143 5871
rect 16206 5787 16236 5871
rect 16290 5787 16320 5871
rect 16410 5787 16440 5871
rect 16516 5787 16546 5871
rect 16624 5787 16654 5955
rect 16708 5787 16738 5955
rect 16845 5787 16875 5955
rect 16989 5787 17019 5871
rect 17073 5787 17103 5871
rect 17191 5787 17221 5871
rect 17299 5787 17329 5871
rect 17395 5787 17425 5955
rect 17467 5787 17497 5955
rect 17665 5855 17695 5983
rect 17762 5787 17792 5987
rect 17950 5803 17980 5931
rect 18045 5787 18075 5987
rect 13449 5463 13479 5591
rect 13533 5463 13563 5591
rect 13721 5513 13751 5597
rect 13814 5513 13844 5597
rect 13898 5513 13928 5597
rect 14018 5513 14048 5597
rect 14124 5513 14154 5597
rect 14232 5429 14262 5597
rect 14316 5429 14346 5597
rect 14453 5429 14483 5597
rect 14597 5513 14627 5597
rect 14681 5513 14711 5597
rect 14799 5513 14829 5597
rect 14907 5513 14937 5597
rect 15003 5429 15033 5597
rect 15075 5429 15105 5597
rect 15273 5401 15303 5529
rect 15370 5397 15400 5597
rect 15558 5453 15588 5581
rect 15653 5397 15683 5597
rect 15841 5463 15871 5591
rect 15925 5463 15955 5591
rect 16113 5513 16143 5597
rect 16206 5513 16236 5597
rect 16290 5513 16320 5597
rect 16410 5513 16440 5597
rect 16516 5513 16546 5597
rect 16624 5429 16654 5597
rect 16708 5429 16738 5597
rect 16845 5429 16875 5597
rect 16989 5513 17019 5597
rect 17073 5513 17103 5597
rect 17191 5513 17221 5597
rect 17299 5513 17329 5597
rect 17395 5429 17425 5597
rect 17467 5429 17497 5597
rect 17665 5401 17695 5529
rect 17762 5397 17792 5597
rect 17950 5453 17980 5581
rect 18045 5397 18075 5597
<< pmoshvt >>
rect 12380 10495 12410 10579
rect 12380 10357 12410 10441
rect 12380 10219 12410 10303
rect 12380 10081 12410 10165
rect 12380 9943 12410 10027
rect 12380 9805 12410 9889
rect 18165 9494 18195 9578
rect 18165 9356 18195 9440
rect 18257 9356 18287 9440
rect 18353 9356 18383 9440
<< ndiff >>
rect 11860 9600 11912 9612
rect 11860 9566 11868 9600
rect 11902 9566 11912 9600
rect 11860 9532 11912 9566
rect 11860 9498 11868 9532
rect 11902 9498 11912 9532
rect 11860 9482 11912 9498
rect 11942 9600 11994 9612
rect 11942 9566 11952 9600
rect 11986 9566 11994 9600
rect 11942 9532 11994 9566
rect 11942 9498 11952 9532
rect 11986 9498 11994 9532
rect 11942 9482 11994 9498
rect 12050 9600 12102 9612
rect 12050 9566 12058 9600
rect 12092 9566 12102 9600
rect 12050 9532 12102 9566
rect 12050 9498 12058 9532
rect 12092 9498 12102 9532
rect 12050 9482 12102 9498
rect 12132 9600 12184 9612
rect 12132 9566 12142 9600
rect 12176 9566 12184 9600
rect 12132 9532 12184 9566
rect 12132 9498 12142 9532
rect 12176 9498 12184 9532
rect 12132 9482 12184 9498
rect 13317 9224 13375 9236
rect 13317 9164 13329 9224
rect 13363 9164 13375 9224
rect 13317 9152 13375 9164
rect 13405 9224 13463 9236
rect 13405 9164 13419 9224
rect 13453 9164 13463 9224
rect 13405 9152 13463 9164
rect 14049 9224 14107 9236
rect 14049 9164 14061 9224
rect 14095 9164 14107 9224
rect 14049 9152 14107 9164
rect 14137 9224 14229 9236
rect 14137 9164 14168 9224
rect 14202 9164 14229 9224
rect 14137 9152 14229 9164
rect 14259 9224 14317 9236
rect 14259 9164 14271 9224
rect 14305 9164 14317 9224
rect 14259 9152 14317 9164
rect 15261 9224 15319 9236
rect 15261 9164 15273 9224
rect 15307 9164 15319 9224
rect 15261 9152 15319 9164
rect 15349 9224 15441 9236
rect 15349 9164 15379 9224
rect 15413 9164 15441 9224
rect 15349 9152 15441 9164
rect 15471 9224 15529 9236
rect 15471 9164 15483 9224
rect 15517 9164 15529 9224
rect 15471 9152 15529 9164
rect 16599 9224 16657 9236
rect 16599 9164 16611 9224
rect 16645 9164 16657 9224
rect 16599 9152 16657 9164
rect 16687 9224 16779 9236
rect 16687 9164 16719 9224
rect 16753 9164 16779 9224
rect 16687 9152 16779 9164
rect 16809 9224 16867 9236
rect 16809 9164 16821 9224
rect 16855 9164 16867 9224
rect 16809 9152 16867 9164
rect 17454 9224 17513 9236
rect 17454 9164 17466 9224
rect 17500 9164 17513 9224
rect 17454 9152 17513 9164
rect 17543 9224 17601 9236
rect 17543 9164 17555 9224
rect 17589 9164 17601 9224
rect 17543 9152 17601 9164
rect 18107 9225 18165 9237
rect 18107 9165 18119 9225
rect 18153 9165 18165 9225
rect 18107 9153 18165 9165
rect 18195 9225 18257 9237
rect 18195 9165 18207 9225
rect 18241 9165 18257 9225
rect 18195 9153 18257 9165
rect 18287 9225 18353 9237
rect 18287 9165 18303 9225
rect 18337 9165 18353 9225
rect 18287 9153 18353 9165
rect 18383 9225 18445 9237
rect 18383 9165 18399 9225
rect 18433 9165 18445 9225
rect 18596 9189 18646 9235
rect 18383 9153 18445 9165
rect 18499 9164 18551 9189
rect 18499 9130 18507 9164
rect 18541 9130 18551 9164
rect 18499 9105 18551 9130
rect 18581 9151 18646 9189
rect 18581 9117 18600 9151
rect 18634 9117 18646 9151
rect 18581 9105 18646 9117
rect 18676 9181 18730 9235
rect 18676 9147 18686 9181
rect 18720 9147 18730 9181
rect 18676 9105 18730 9147
rect 18760 9223 18813 9235
rect 18760 9189 18770 9223
rect 18804 9189 18813 9223
rect 18760 9155 18813 9189
rect 18760 9121 18770 9155
rect 18804 9121 18813 9155
rect 18760 9105 18813 9121
rect 18107 9087 18165 9099
rect 12297 9040 12355 9052
rect 12297 8980 12309 9040
rect 12343 8980 12355 9040
rect 12297 8968 12355 8980
rect 12385 8968 12427 9052
rect 12457 9040 12515 9052
rect 12457 8980 12469 9040
rect 12503 8980 12515 9040
rect 18107 9027 18119 9087
rect 18153 9027 18165 9087
rect 18107 9015 18165 9027
rect 18195 9087 18253 9099
rect 18195 9027 18207 9087
rect 18241 9027 18253 9087
rect 18195 9015 18253 9027
rect 12457 8968 12515 8980
rect 12297 8902 12355 8914
rect 12297 8842 12309 8902
rect 12343 8842 12355 8902
rect 12297 8830 12355 8842
rect 12385 8830 12427 8914
rect 12457 8902 12515 8914
rect 12457 8842 12469 8902
rect 12503 8842 12515 8902
rect 12457 8830 12515 8842
rect 12297 8764 12355 8776
rect 12297 8704 12309 8764
rect 12343 8704 12355 8764
rect 12297 8692 12355 8704
rect 12385 8692 12427 8776
rect 12457 8764 12515 8776
rect 12457 8704 12469 8764
rect 12503 8704 12515 8764
rect 12457 8692 12515 8704
rect 12297 8626 12355 8638
rect 12297 8566 12309 8626
rect 12343 8566 12355 8626
rect 12297 8554 12355 8566
rect 12385 8554 12427 8638
rect 12457 8626 12515 8638
rect 12457 8566 12469 8626
rect 12503 8566 12515 8626
rect 12457 8554 12515 8566
rect 12297 8488 12355 8500
rect 12297 8428 12309 8488
rect 12343 8428 12355 8488
rect 12297 8416 12355 8428
rect 12385 8416 12427 8500
rect 12457 8488 12515 8500
rect 12457 8428 12469 8488
rect 12503 8428 12515 8488
rect 12457 8416 12515 8428
rect 12297 8350 12355 8362
rect 12297 8290 12309 8350
rect 12343 8290 12355 8350
rect 12297 8278 12355 8290
rect 12385 8278 12427 8362
rect 12457 8350 12515 8362
rect 12457 8290 12469 8350
rect 12503 8290 12515 8350
rect 12457 8278 12515 8290
rect 12297 8212 12355 8224
rect 12297 8152 12309 8212
rect 12343 8152 12355 8212
rect 12297 8140 12355 8152
rect 12385 8140 12427 8224
rect 12457 8212 12515 8224
rect 12457 8152 12469 8212
rect 12503 8152 12515 8212
rect 12457 8140 12515 8152
rect 12297 8074 12355 8086
rect 12297 8014 12309 8074
rect 12343 8014 12355 8074
rect 12297 8002 12355 8014
rect 12385 8002 12427 8086
rect 12457 8074 12515 8086
rect 12457 8014 12469 8074
rect 12503 8014 12515 8074
rect 12457 8002 12515 8014
rect 13397 7479 13449 7517
rect 13397 7445 13405 7479
rect 13439 7445 13449 7479
rect 13397 7433 13449 7445
rect 13479 7505 13533 7517
rect 13479 7471 13489 7505
rect 13523 7471 13533 7505
rect 13479 7433 13533 7471
rect 13563 7479 13615 7517
rect 13563 7445 13573 7479
rect 13607 7445 13615 7479
rect 13563 7433 13615 7445
rect 13669 7505 13721 7517
rect 13669 7471 13677 7505
rect 13711 7471 13721 7505
rect 13669 7433 13721 7471
rect 13751 7487 13816 7517
rect 13751 7453 13761 7487
rect 13795 7453 13816 7487
rect 13751 7445 13816 7453
rect 13846 7505 13922 7517
rect 13846 7471 13867 7505
rect 13901 7471 13922 7505
rect 13846 7445 13922 7471
rect 13952 7445 14018 7517
rect 13751 7433 13801 7445
rect 13967 7433 14018 7445
rect 14048 7509 14128 7517
rect 14048 7475 14084 7509
rect 14118 7475 14128 7509
rect 14048 7433 14128 7475
rect 14158 7489 14228 7517
rect 14158 7455 14168 7489
rect 14202 7455 14228 7489
rect 14158 7433 14228 7455
rect 14178 7389 14228 7433
rect 14258 7445 14312 7517
rect 14258 7411 14268 7445
rect 14302 7411 14312 7445
rect 14258 7389 14312 7411
rect 14342 7471 14394 7517
rect 14342 7437 14352 7471
rect 14386 7437 14394 7471
rect 14342 7389 14394 7437
rect 14448 7505 14500 7517
rect 14448 7471 14456 7505
rect 14490 7471 14500 7505
rect 14448 7389 14500 7471
rect 14530 7445 14595 7517
rect 14625 7505 14704 7517
rect 14625 7471 14650 7505
rect 14684 7471 14704 7505
rect 14625 7445 14704 7471
rect 14734 7445 14799 7517
rect 14530 7389 14580 7445
rect 14749 7433 14799 7445
rect 14829 7509 14885 7517
rect 14829 7475 14841 7509
rect 14875 7475 14885 7509
rect 14829 7433 14885 7475
rect 14915 7489 15003 7517
rect 14915 7455 14943 7489
rect 14977 7455 15003 7489
rect 14915 7433 15003 7455
rect 14953 7389 15003 7433
rect 15033 7445 15087 7517
rect 15033 7411 15043 7445
rect 15077 7411 15087 7445
rect 15033 7389 15087 7411
rect 15117 7497 15169 7517
rect 15117 7463 15127 7497
rect 15161 7463 15169 7497
rect 15117 7389 15169 7463
rect 15223 7495 15275 7517
rect 15223 7461 15231 7495
rect 15265 7461 15275 7495
rect 15223 7433 15275 7461
rect 15305 7505 15370 7517
rect 15305 7471 15326 7505
rect 15360 7471 15370 7505
rect 15305 7433 15370 7471
rect 15320 7387 15370 7433
rect 15400 7471 15452 7517
rect 15400 7437 15410 7471
rect 15444 7437 15452 7471
rect 15400 7387 15452 7437
rect 15506 7479 15558 7517
rect 15506 7445 15514 7479
rect 15548 7445 15558 7479
rect 15506 7433 15558 7445
rect 15588 7505 15653 7517
rect 15588 7471 15609 7505
rect 15643 7471 15653 7505
rect 15588 7433 15653 7471
rect 15603 7387 15653 7433
rect 15683 7469 15735 7517
rect 15683 7435 15693 7469
rect 15727 7435 15735 7469
rect 15683 7387 15735 7435
rect 15789 7479 15841 7517
rect 15789 7445 15797 7479
rect 15831 7445 15841 7479
rect 15789 7433 15841 7445
rect 15871 7505 15925 7517
rect 15871 7471 15881 7505
rect 15915 7471 15925 7505
rect 15871 7433 15925 7471
rect 15955 7479 16007 7517
rect 15955 7445 15965 7479
rect 15999 7445 16007 7479
rect 15955 7433 16007 7445
rect 16061 7505 16113 7517
rect 16061 7471 16069 7505
rect 16103 7471 16113 7505
rect 16061 7433 16113 7471
rect 16143 7487 16208 7517
rect 16143 7453 16153 7487
rect 16187 7453 16208 7487
rect 16143 7445 16208 7453
rect 16238 7505 16314 7517
rect 16238 7471 16259 7505
rect 16293 7471 16314 7505
rect 16238 7445 16314 7471
rect 16344 7445 16410 7517
rect 16143 7433 16193 7445
rect 16359 7433 16410 7445
rect 16440 7509 16520 7517
rect 16440 7475 16476 7509
rect 16510 7475 16520 7509
rect 16440 7433 16520 7475
rect 16550 7489 16620 7517
rect 16550 7455 16560 7489
rect 16594 7455 16620 7489
rect 16550 7433 16620 7455
rect 16570 7389 16620 7433
rect 16650 7445 16704 7517
rect 16650 7411 16660 7445
rect 16694 7411 16704 7445
rect 16650 7389 16704 7411
rect 16734 7471 16786 7517
rect 16734 7437 16744 7471
rect 16778 7437 16786 7471
rect 16734 7389 16786 7437
rect 16840 7505 16892 7517
rect 16840 7471 16848 7505
rect 16882 7471 16892 7505
rect 16840 7389 16892 7471
rect 16922 7445 16987 7517
rect 17017 7505 17096 7517
rect 17017 7471 17042 7505
rect 17076 7471 17096 7505
rect 17017 7445 17096 7471
rect 17126 7445 17191 7517
rect 16922 7389 16972 7445
rect 17141 7433 17191 7445
rect 17221 7509 17277 7517
rect 17221 7475 17233 7509
rect 17267 7475 17277 7509
rect 17221 7433 17277 7475
rect 17307 7489 17395 7517
rect 17307 7455 17335 7489
rect 17369 7455 17395 7489
rect 17307 7433 17395 7455
rect 17345 7389 17395 7433
rect 17425 7445 17479 7517
rect 17425 7411 17435 7445
rect 17469 7411 17479 7445
rect 17425 7389 17479 7411
rect 17509 7497 17561 7517
rect 17509 7463 17519 7497
rect 17553 7463 17561 7497
rect 17509 7389 17561 7463
rect 17615 7495 17667 7517
rect 17615 7461 17623 7495
rect 17657 7461 17667 7495
rect 17615 7433 17667 7461
rect 17697 7505 17762 7517
rect 17697 7471 17718 7505
rect 17752 7471 17762 7505
rect 17697 7433 17762 7471
rect 17712 7387 17762 7433
rect 17792 7471 17844 7517
rect 17792 7437 17802 7471
rect 17836 7437 17844 7471
rect 17792 7387 17844 7437
rect 17898 7479 17950 7517
rect 17898 7445 17906 7479
rect 17940 7445 17950 7479
rect 17898 7433 17950 7445
rect 17980 7505 18045 7517
rect 17980 7471 18001 7505
rect 18035 7471 18045 7505
rect 17980 7433 18045 7471
rect 17995 7387 18045 7433
rect 18075 7469 18127 7517
rect 18075 7435 18085 7469
rect 18119 7435 18127 7469
rect 18075 7387 18127 7435
rect 13397 6499 13449 6511
rect 13397 6465 13405 6499
rect 13439 6465 13449 6499
rect 13397 6427 13449 6465
rect 13479 6473 13533 6511
rect 13479 6439 13489 6473
rect 13523 6439 13533 6473
rect 13479 6427 13533 6439
rect 13563 6499 13615 6511
rect 13563 6465 13573 6499
rect 13607 6465 13615 6499
rect 13563 6427 13615 6465
rect 13669 6473 13721 6511
rect 13669 6439 13677 6473
rect 13711 6439 13721 6473
rect 13669 6427 13721 6439
rect 13751 6499 13801 6511
rect 14178 6511 14228 6555
rect 13967 6499 14018 6511
rect 13751 6491 13816 6499
rect 13751 6457 13761 6491
rect 13795 6457 13816 6491
rect 13751 6427 13816 6457
rect 13846 6473 13922 6499
rect 13846 6439 13867 6473
rect 13901 6439 13922 6473
rect 13846 6427 13922 6439
rect 13952 6427 14018 6499
rect 14048 6469 14128 6511
rect 14048 6435 14084 6469
rect 14118 6435 14128 6469
rect 14048 6427 14128 6435
rect 14158 6489 14228 6511
rect 14158 6455 14168 6489
rect 14202 6455 14228 6489
rect 14158 6427 14228 6455
rect 14258 6533 14312 6555
rect 14258 6499 14268 6533
rect 14302 6499 14312 6533
rect 14258 6427 14312 6499
rect 14342 6507 14394 6555
rect 14342 6473 14352 6507
rect 14386 6473 14394 6507
rect 14342 6427 14394 6473
rect 14448 6473 14500 6555
rect 14448 6439 14456 6473
rect 14490 6439 14500 6473
rect 14448 6427 14500 6439
rect 14530 6499 14580 6555
rect 14953 6511 15003 6555
rect 14749 6499 14799 6511
rect 14530 6427 14595 6499
rect 14625 6473 14704 6499
rect 14625 6439 14650 6473
rect 14684 6439 14704 6473
rect 14625 6427 14704 6439
rect 14734 6427 14799 6499
rect 14829 6469 14885 6511
rect 14829 6435 14841 6469
rect 14875 6435 14885 6469
rect 14829 6427 14885 6435
rect 14915 6489 15003 6511
rect 14915 6455 14943 6489
rect 14977 6455 15003 6489
rect 14915 6427 15003 6455
rect 15033 6533 15087 6555
rect 15033 6499 15043 6533
rect 15077 6499 15087 6533
rect 15033 6427 15087 6499
rect 15117 6481 15169 6555
rect 15320 6511 15370 6557
rect 15117 6447 15127 6481
rect 15161 6447 15169 6481
rect 15117 6427 15169 6447
rect 15223 6483 15275 6511
rect 15223 6449 15231 6483
rect 15265 6449 15275 6483
rect 15223 6427 15275 6449
rect 15305 6473 15370 6511
rect 15305 6439 15326 6473
rect 15360 6439 15370 6473
rect 15305 6427 15370 6439
rect 15400 6507 15452 6557
rect 15603 6511 15653 6557
rect 15400 6473 15410 6507
rect 15444 6473 15452 6507
rect 15400 6427 15452 6473
rect 15506 6499 15558 6511
rect 15506 6465 15514 6499
rect 15548 6465 15558 6499
rect 15506 6427 15558 6465
rect 15588 6473 15653 6511
rect 15588 6439 15609 6473
rect 15643 6439 15653 6473
rect 15588 6427 15653 6439
rect 15683 6509 15735 6557
rect 15683 6475 15693 6509
rect 15727 6475 15735 6509
rect 15683 6427 15735 6475
rect 15789 6499 15841 6511
rect 15789 6465 15797 6499
rect 15831 6465 15841 6499
rect 15789 6427 15841 6465
rect 15871 6473 15925 6511
rect 15871 6439 15881 6473
rect 15915 6439 15925 6473
rect 15871 6427 15925 6439
rect 15955 6499 16007 6511
rect 15955 6465 15965 6499
rect 15999 6465 16007 6499
rect 15955 6427 16007 6465
rect 16061 6473 16113 6511
rect 16061 6439 16069 6473
rect 16103 6439 16113 6473
rect 16061 6427 16113 6439
rect 16143 6499 16193 6511
rect 16570 6511 16620 6555
rect 16359 6499 16410 6511
rect 16143 6491 16208 6499
rect 16143 6457 16153 6491
rect 16187 6457 16208 6491
rect 16143 6427 16208 6457
rect 16238 6473 16314 6499
rect 16238 6439 16259 6473
rect 16293 6439 16314 6473
rect 16238 6427 16314 6439
rect 16344 6427 16410 6499
rect 16440 6469 16520 6511
rect 16440 6435 16476 6469
rect 16510 6435 16520 6469
rect 16440 6427 16520 6435
rect 16550 6489 16620 6511
rect 16550 6455 16560 6489
rect 16594 6455 16620 6489
rect 16550 6427 16620 6455
rect 16650 6533 16704 6555
rect 16650 6499 16660 6533
rect 16694 6499 16704 6533
rect 16650 6427 16704 6499
rect 16734 6507 16786 6555
rect 16734 6473 16744 6507
rect 16778 6473 16786 6507
rect 16734 6427 16786 6473
rect 16840 6473 16892 6555
rect 16840 6439 16848 6473
rect 16882 6439 16892 6473
rect 16840 6427 16892 6439
rect 16922 6499 16972 6555
rect 17345 6511 17395 6555
rect 17141 6499 17191 6511
rect 16922 6427 16987 6499
rect 17017 6473 17096 6499
rect 17017 6439 17042 6473
rect 17076 6439 17096 6473
rect 17017 6427 17096 6439
rect 17126 6427 17191 6499
rect 17221 6469 17277 6511
rect 17221 6435 17233 6469
rect 17267 6435 17277 6469
rect 17221 6427 17277 6435
rect 17307 6489 17395 6511
rect 17307 6455 17335 6489
rect 17369 6455 17395 6489
rect 17307 6427 17395 6455
rect 17425 6533 17479 6555
rect 17425 6499 17435 6533
rect 17469 6499 17479 6533
rect 17425 6427 17479 6499
rect 17509 6481 17561 6555
rect 17712 6511 17762 6557
rect 17509 6447 17519 6481
rect 17553 6447 17561 6481
rect 17509 6427 17561 6447
rect 17615 6483 17667 6511
rect 17615 6449 17623 6483
rect 17657 6449 17667 6483
rect 17615 6427 17667 6449
rect 17697 6473 17762 6511
rect 17697 6439 17718 6473
rect 17752 6439 17762 6473
rect 17697 6427 17762 6439
rect 17792 6507 17844 6557
rect 17995 6511 18045 6557
rect 17792 6473 17802 6507
rect 17836 6473 17844 6507
rect 17792 6427 17844 6473
rect 17898 6499 17950 6511
rect 17898 6465 17906 6499
rect 17940 6465 17950 6499
rect 17898 6427 17950 6465
rect 17980 6473 18045 6511
rect 17980 6439 18001 6473
rect 18035 6439 18045 6473
rect 17980 6427 18045 6439
rect 18075 6509 18127 6557
rect 18075 6475 18085 6509
rect 18119 6475 18127 6509
rect 18075 6427 18127 6475
rect 13397 6199 13449 6237
rect 13397 6165 13405 6199
rect 13439 6165 13449 6199
rect 13397 6153 13449 6165
rect 13479 6225 13533 6237
rect 13479 6191 13489 6225
rect 13523 6191 13533 6225
rect 13479 6153 13533 6191
rect 13563 6199 13615 6237
rect 13563 6165 13573 6199
rect 13607 6165 13615 6199
rect 13563 6153 13615 6165
rect 13669 6225 13721 6237
rect 13669 6191 13677 6225
rect 13711 6191 13721 6225
rect 13669 6153 13721 6191
rect 13751 6207 13816 6237
rect 13751 6173 13761 6207
rect 13795 6173 13816 6207
rect 13751 6165 13816 6173
rect 13846 6225 13922 6237
rect 13846 6191 13867 6225
rect 13901 6191 13922 6225
rect 13846 6165 13922 6191
rect 13952 6165 14018 6237
rect 13751 6153 13801 6165
rect 13967 6153 14018 6165
rect 14048 6229 14128 6237
rect 14048 6195 14084 6229
rect 14118 6195 14128 6229
rect 14048 6153 14128 6195
rect 14158 6209 14228 6237
rect 14158 6175 14168 6209
rect 14202 6175 14228 6209
rect 14158 6153 14228 6175
rect 14178 6109 14228 6153
rect 14258 6165 14312 6237
rect 14258 6131 14268 6165
rect 14302 6131 14312 6165
rect 14258 6109 14312 6131
rect 14342 6191 14394 6237
rect 14342 6157 14352 6191
rect 14386 6157 14394 6191
rect 14342 6109 14394 6157
rect 14448 6225 14500 6237
rect 14448 6191 14456 6225
rect 14490 6191 14500 6225
rect 14448 6109 14500 6191
rect 14530 6165 14595 6237
rect 14625 6225 14704 6237
rect 14625 6191 14650 6225
rect 14684 6191 14704 6225
rect 14625 6165 14704 6191
rect 14734 6165 14799 6237
rect 14530 6109 14580 6165
rect 14749 6153 14799 6165
rect 14829 6229 14885 6237
rect 14829 6195 14841 6229
rect 14875 6195 14885 6229
rect 14829 6153 14885 6195
rect 14915 6209 15003 6237
rect 14915 6175 14943 6209
rect 14977 6175 15003 6209
rect 14915 6153 15003 6175
rect 14953 6109 15003 6153
rect 15033 6165 15087 6237
rect 15033 6131 15043 6165
rect 15077 6131 15087 6165
rect 15033 6109 15087 6131
rect 15117 6217 15169 6237
rect 15117 6183 15127 6217
rect 15161 6183 15169 6217
rect 15117 6109 15169 6183
rect 15223 6215 15275 6237
rect 15223 6181 15231 6215
rect 15265 6181 15275 6215
rect 15223 6153 15275 6181
rect 15305 6225 15370 6237
rect 15305 6191 15326 6225
rect 15360 6191 15370 6225
rect 15305 6153 15370 6191
rect 15320 6107 15370 6153
rect 15400 6191 15452 6237
rect 15400 6157 15410 6191
rect 15444 6157 15452 6191
rect 15400 6107 15452 6157
rect 15506 6199 15558 6237
rect 15506 6165 15514 6199
rect 15548 6165 15558 6199
rect 15506 6153 15558 6165
rect 15588 6225 15653 6237
rect 15588 6191 15609 6225
rect 15643 6191 15653 6225
rect 15588 6153 15653 6191
rect 15603 6107 15653 6153
rect 15683 6189 15735 6237
rect 15683 6155 15693 6189
rect 15727 6155 15735 6189
rect 15683 6107 15735 6155
rect 15789 6199 15841 6237
rect 15789 6165 15797 6199
rect 15831 6165 15841 6199
rect 15789 6153 15841 6165
rect 15871 6225 15925 6237
rect 15871 6191 15881 6225
rect 15915 6191 15925 6225
rect 15871 6153 15925 6191
rect 15955 6199 16007 6237
rect 15955 6165 15965 6199
rect 15999 6165 16007 6199
rect 15955 6153 16007 6165
rect 16061 6225 16113 6237
rect 16061 6191 16069 6225
rect 16103 6191 16113 6225
rect 16061 6153 16113 6191
rect 16143 6207 16208 6237
rect 16143 6173 16153 6207
rect 16187 6173 16208 6207
rect 16143 6165 16208 6173
rect 16238 6225 16314 6237
rect 16238 6191 16259 6225
rect 16293 6191 16314 6225
rect 16238 6165 16314 6191
rect 16344 6165 16410 6237
rect 16143 6153 16193 6165
rect 16359 6153 16410 6165
rect 16440 6229 16520 6237
rect 16440 6195 16476 6229
rect 16510 6195 16520 6229
rect 16440 6153 16520 6195
rect 16550 6209 16620 6237
rect 16550 6175 16560 6209
rect 16594 6175 16620 6209
rect 16550 6153 16620 6175
rect 16570 6109 16620 6153
rect 16650 6165 16704 6237
rect 16650 6131 16660 6165
rect 16694 6131 16704 6165
rect 16650 6109 16704 6131
rect 16734 6191 16786 6237
rect 16734 6157 16744 6191
rect 16778 6157 16786 6191
rect 16734 6109 16786 6157
rect 16840 6225 16892 6237
rect 16840 6191 16848 6225
rect 16882 6191 16892 6225
rect 16840 6109 16892 6191
rect 16922 6165 16987 6237
rect 17017 6225 17096 6237
rect 17017 6191 17042 6225
rect 17076 6191 17096 6225
rect 17017 6165 17096 6191
rect 17126 6165 17191 6237
rect 16922 6109 16972 6165
rect 17141 6153 17191 6165
rect 17221 6229 17277 6237
rect 17221 6195 17233 6229
rect 17267 6195 17277 6229
rect 17221 6153 17277 6195
rect 17307 6209 17395 6237
rect 17307 6175 17335 6209
rect 17369 6175 17395 6209
rect 17307 6153 17395 6175
rect 17345 6109 17395 6153
rect 17425 6165 17479 6237
rect 17425 6131 17435 6165
rect 17469 6131 17479 6165
rect 17425 6109 17479 6131
rect 17509 6217 17561 6237
rect 17509 6183 17519 6217
rect 17553 6183 17561 6217
rect 17509 6109 17561 6183
rect 17615 6215 17667 6237
rect 17615 6181 17623 6215
rect 17657 6181 17667 6215
rect 17615 6153 17667 6181
rect 17697 6225 17762 6237
rect 17697 6191 17718 6225
rect 17752 6191 17762 6225
rect 17697 6153 17762 6191
rect 17712 6107 17762 6153
rect 17792 6191 17844 6237
rect 17792 6157 17802 6191
rect 17836 6157 17844 6191
rect 17792 6107 17844 6157
rect 17898 6199 17950 6237
rect 17898 6165 17906 6199
rect 17940 6165 17950 6199
rect 17898 6153 17950 6165
rect 17980 6225 18045 6237
rect 17980 6191 18001 6225
rect 18035 6191 18045 6225
rect 17980 6153 18045 6191
rect 17995 6107 18045 6153
rect 18075 6189 18127 6237
rect 18075 6155 18085 6189
rect 18119 6155 18127 6189
rect 18075 6107 18127 6155
rect 13397 5219 13449 5231
rect 13397 5185 13405 5219
rect 13439 5185 13449 5219
rect 13397 5147 13449 5185
rect 13479 5193 13533 5231
rect 13479 5159 13489 5193
rect 13523 5159 13533 5193
rect 13479 5147 13533 5159
rect 13563 5219 13615 5231
rect 13563 5185 13573 5219
rect 13607 5185 13615 5219
rect 13563 5147 13615 5185
rect 13669 5193 13721 5231
rect 13669 5159 13677 5193
rect 13711 5159 13721 5193
rect 13669 5147 13721 5159
rect 13751 5219 13801 5231
rect 14178 5231 14228 5275
rect 13967 5219 14018 5231
rect 13751 5211 13816 5219
rect 13751 5177 13761 5211
rect 13795 5177 13816 5211
rect 13751 5147 13816 5177
rect 13846 5193 13922 5219
rect 13846 5159 13867 5193
rect 13901 5159 13922 5193
rect 13846 5147 13922 5159
rect 13952 5147 14018 5219
rect 14048 5189 14128 5231
rect 14048 5155 14084 5189
rect 14118 5155 14128 5189
rect 14048 5147 14128 5155
rect 14158 5209 14228 5231
rect 14158 5175 14168 5209
rect 14202 5175 14228 5209
rect 14158 5147 14228 5175
rect 14258 5253 14312 5275
rect 14258 5219 14268 5253
rect 14302 5219 14312 5253
rect 14258 5147 14312 5219
rect 14342 5227 14394 5275
rect 14342 5193 14352 5227
rect 14386 5193 14394 5227
rect 14342 5147 14394 5193
rect 14448 5193 14500 5275
rect 14448 5159 14456 5193
rect 14490 5159 14500 5193
rect 14448 5147 14500 5159
rect 14530 5219 14580 5275
rect 14953 5231 15003 5275
rect 14749 5219 14799 5231
rect 14530 5147 14595 5219
rect 14625 5193 14704 5219
rect 14625 5159 14650 5193
rect 14684 5159 14704 5193
rect 14625 5147 14704 5159
rect 14734 5147 14799 5219
rect 14829 5189 14885 5231
rect 14829 5155 14841 5189
rect 14875 5155 14885 5189
rect 14829 5147 14885 5155
rect 14915 5209 15003 5231
rect 14915 5175 14943 5209
rect 14977 5175 15003 5209
rect 14915 5147 15003 5175
rect 15033 5253 15087 5275
rect 15033 5219 15043 5253
rect 15077 5219 15087 5253
rect 15033 5147 15087 5219
rect 15117 5201 15169 5275
rect 15320 5231 15370 5277
rect 15117 5167 15127 5201
rect 15161 5167 15169 5201
rect 15117 5147 15169 5167
rect 15223 5203 15275 5231
rect 15223 5169 15231 5203
rect 15265 5169 15275 5203
rect 15223 5147 15275 5169
rect 15305 5193 15370 5231
rect 15305 5159 15326 5193
rect 15360 5159 15370 5193
rect 15305 5147 15370 5159
rect 15400 5227 15452 5277
rect 15603 5231 15653 5277
rect 15400 5193 15410 5227
rect 15444 5193 15452 5227
rect 15400 5147 15452 5193
rect 15506 5219 15558 5231
rect 15506 5185 15514 5219
rect 15548 5185 15558 5219
rect 15506 5147 15558 5185
rect 15588 5193 15653 5231
rect 15588 5159 15609 5193
rect 15643 5159 15653 5193
rect 15588 5147 15653 5159
rect 15683 5229 15735 5277
rect 15683 5195 15693 5229
rect 15727 5195 15735 5229
rect 15683 5147 15735 5195
rect 15789 5219 15841 5231
rect 15789 5185 15797 5219
rect 15831 5185 15841 5219
rect 15789 5147 15841 5185
rect 15871 5193 15925 5231
rect 15871 5159 15881 5193
rect 15915 5159 15925 5193
rect 15871 5147 15925 5159
rect 15955 5219 16007 5231
rect 15955 5185 15965 5219
rect 15999 5185 16007 5219
rect 15955 5147 16007 5185
rect 16061 5193 16113 5231
rect 16061 5159 16069 5193
rect 16103 5159 16113 5193
rect 16061 5147 16113 5159
rect 16143 5219 16193 5231
rect 16570 5231 16620 5275
rect 16359 5219 16410 5231
rect 16143 5211 16208 5219
rect 16143 5177 16153 5211
rect 16187 5177 16208 5211
rect 16143 5147 16208 5177
rect 16238 5193 16314 5219
rect 16238 5159 16259 5193
rect 16293 5159 16314 5193
rect 16238 5147 16314 5159
rect 16344 5147 16410 5219
rect 16440 5189 16520 5231
rect 16440 5155 16476 5189
rect 16510 5155 16520 5189
rect 16440 5147 16520 5155
rect 16550 5209 16620 5231
rect 16550 5175 16560 5209
rect 16594 5175 16620 5209
rect 16550 5147 16620 5175
rect 16650 5253 16704 5275
rect 16650 5219 16660 5253
rect 16694 5219 16704 5253
rect 16650 5147 16704 5219
rect 16734 5227 16786 5275
rect 16734 5193 16744 5227
rect 16778 5193 16786 5227
rect 16734 5147 16786 5193
rect 16840 5193 16892 5275
rect 16840 5159 16848 5193
rect 16882 5159 16892 5193
rect 16840 5147 16892 5159
rect 16922 5219 16972 5275
rect 17345 5231 17395 5275
rect 17141 5219 17191 5231
rect 16922 5147 16987 5219
rect 17017 5193 17096 5219
rect 17017 5159 17042 5193
rect 17076 5159 17096 5193
rect 17017 5147 17096 5159
rect 17126 5147 17191 5219
rect 17221 5189 17277 5231
rect 17221 5155 17233 5189
rect 17267 5155 17277 5189
rect 17221 5147 17277 5155
rect 17307 5209 17395 5231
rect 17307 5175 17335 5209
rect 17369 5175 17395 5209
rect 17307 5147 17395 5175
rect 17425 5253 17479 5275
rect 17425 5219 17435 5253
rect 17469 5219 17479 5253
rect 17425 5147 17479 5219
rect 17509 5201 17561 5275
rect 17712 5231 17762 5277
rect 17509 5167 17519 5201
rect 17553 5167 17561 5201
rect 17509 5147 17561 5167
rect 17615 5203 17667 5231
rect 17615 5169 17623 5203
rect 17657 5169 17667 5203
rect 17615 5147 17667 5169
rect 17697 5193 17762 5231
rect 17697 5159 17718 5193
rect 17752 5159 17762 5193
rect 17697 5147 17762 5159
rect 17792 5227 17844 5277
rect 17995 5231 18045 5277
rect 17792 5193 17802 5227
rect 17836 5193 17844 5227
rect 17792 5147 17844 5193
rect 17898 5219 17950 5231
rect 17898 5185 17906 5219
rect 17940 5185 17950 5219
rect 17898 5147 17950 5185
rect 17980 5193 18045 5231
rect 17980 5159 18001 5193
rect 18035 5159 18045 5193
rect 17980 5147 18045 5159
rect 18075 5229 18127 5277
rect 18075 5195 18085 5229
rect 18119 5195 18127 5229
rect 18075 5147 18127 5195
<< pdiff >>
rect 12322 10567 12380 10579
rect 12322 10507 12334 10567
rect 12368 10507 12380 10567
rect 12322 10495 12380 10507
rect 12410 10567 12468 10579
rect 12410 10507 12422 10567
rect 12456 10507 12468 10567
rect 12410 10495 12468 10507
rect 12322 10429 12380 10441
rect 12322 10369 12334 10429
rect 12368 10369 12380 10429
rect 12322 10357 12380 10369
rect 12410 10429 12468 10441
rect 12410 10369 12422 10429
rect 12456 10369 12468 10429
rect 12410 10357 12468 10369
rect 12322 10291 12380 10303
rect 12322 10231 12334 10291
rect 12368 10231 12380 10291
rect 12322 10219 12380 10231
rect 12410 10291 12468 10303
rect 12410 10231 12422 10291
rect 12456 10231 12468 10291
rect 12410 10219 12468 10231
rect 12322 10153 12380 10165
rect 12322 10093 12334 10153
rect 12368 10093 12380 10153
rect 12322 10081 12380 10093
rect 12410 10153 12468 10165
rect 12410 10093 12422 10153
rect 12456 10093 12468 10153
rect 12410 10081 12468 10093
rect 12322 10015 12380 10027
rect 12322 9955 12334 10015
rect 12368 9955 12380 10015
rect 12322 9943 12380 9955
rect 12410 10015 12468 10027
rect 12410 9955 12422 10015
rect 12456 9955 12468 10015
rect 12410 9943 12468 9955
rect 11860 9920 11912 9932
rect 11860 9886 11868 9920
rect 11902 9886 11912 9920
rect 11860 9852 11912 9886
rect 11860 9818 11868 9852
rect 11902 9818 11912 9852
rect 11860 9784 11912 9818
rect 11860 9750 11868 9784
rect 11902 9750 11912 9784
rect 11860 9732 11912 9750
rect 11942 9920 11994 9932
rect 11942 9886 11952 9920
rect 11986 9886 11994 9920
rect 11942 9852 11994 9886
rect 11942 9818 11952 9852
rect 11986 9818 11994 9852
rect 11942 9784 11994 9818
rect 11942 9750 11952 9784
rect 11986 9750 11994 9784
rect 11942 9732 11994 9750
rect 12050 9920 12102 9932
rect 12050 9886 12058 9920
rect 12092 9886 12102 9920
rect 12050 9852 12102 9886
rect 12050 9818 12058 9852
rect 12092 9818 12102 9852
rect 12050 9784 12102 9818
rect 12050 9750 12058 9784
rect 12092 9750 12102 9784
rect 12050 9732 12102 9750
rect 12132 9920 12184 9932
rect 12132 9886 12142 9920
rect 12176 9886 12184 9920
rect 12132 9852 12184 9886
rect 12132 9818 12142 9852
rect 12176 9818 12184 9852
rect 12132 9784 12184 9818
rect 12322 9877 12380 9889
rect 12322 9817 12334 9877
rect 12368 9817 12380 9877
rect 12322 9805 12380 9817
rect 12410 9877 12468 9889
rect 12410 9817 12422 9877
rect 12456 9817 12468 9877
rect 12410 9805 12468 9817
rect 12132 9750 12142 9784
rect 12176 9750 12184 9784
rect 12132 9732 12184 9750
rect 18107 9566 18165 9578
rect 18107 9506 18119 9566
rect 18153 9506 18165 9566
rect 18107 9494 18165 9506
rect 18195 9566 18253 9578
rect 18195 9506 18207 9566
rect 18241 9506 18253 9566
rect 18596 9547 18646 9555
rect 18195 9494 18253 9506
rect 18499 9535 18551 9547
rect 18499 9501 18507 9535
rect 18541 9501 18551 9535
rect 18499 9467 18551 9501
rect 12964 9422 13022 9434
rect 12964 9362 12976 9422
rect 13010 9362 13022 9422
rect 12964 9350 13022 9362
rect 13052 9425 13110 9434
rect 13052 9365 13064 9425
rect 13098 9365 13110 9425
rect 13052 9350 13110 9365
rect 13696 9425 13754 9437
rect 13696 9365 13708 9425
rect 13742 9365 13754 9425
rect 13696 9353 13754 9365
rect 13784 9425 13880 9437
rect 13784 9365 13813 9425
rect 13847 9365 13880 9425
rect 13784 9353 13880 9365
rect 13910 9425 13968 9437
rect 13910 9365 13922 9425
rect 13956 9365 13968 9425
rect 13910 9353 13968 9365
rect 14908 9425 14966 9437
rect 14908 9365 14920 9425
rect 14954 9365 14966 9425
rect 14908 9353 14966 9365
rect 14996 9425 15092 9437
rect 14996 9365 15024 9425
rect 15058 9365 15092 9425
rect 14996 9353 15092 9365
rect 15122 9425 15180 9437
rect 15122 9365 15134 9425
rect 15168 9365 15180 9425
rect 15122 9353 15180 9365
rect 16120 9425 16178 9437
rect 16120 9365 16132 9425
rect 16166 9365 16178 9425
rect 16120 9353 16178 9365
rect 16208 9425 16304 9437
rect 16208 9365 16237 9425
rect 16271 9365 16304 9425
rect 16208 9353 16304 9365
rect 16334 9425 16392 9437
rect 16334 9365 16346 9425
rect 16380 9365 16392 9425
rect 16334 9353 16392 9365
rect 17332 9425 17390 9437
rect 17332 9365 17344 9425
rect 17378 9365 17390 9425
rect 17332 9353 17390 9365
rect 17420 9425 17516 9437
rect 17420 9365 17451 9425
rect 17485 9365 17516 9425
rect 17420 9353 17516 9365
rect 17546 9425 17604 9437
rect 17546 9365 17558 9425
rect 17592 9365 17604 9425
rect 17546 9353 17604 9365
rect 18107 9428 18165 9440
rect 18107 9368 18119 9428
rect 18153 9368 18165 9428
rect 18107 9356 18165 9368
rect 18195 9428 18257 9440
rect 18195 9368 18207 9428
rect 18241 9368 18257 9428
rect 18195 9356 18257 9368
rect 18287 9428 18353 9440
rect 18287 9368 18303 9428
rect 18337 9368 18353 9428
rect 18287 9356 18353 9368
rect 18383 9428 18445 9440
rect 18383 9368 18399 9428
rect 18433 9368 18445 9428
rect 18499 9433 18507 9467
rect 18541 9433 18551 9467
rect 18499 9419 18551 9433
rect 18581 9535 18646 9547
rect 18581 9501 18600 9535
rect 18634 9501 18646 9535
rect 18581 9467 18646 9501
rect 18581 9433 18600 9467
rect 18634 9433 18646 9467
rect 18581 9419 18646 9433
rect 18383 9356 18445 9368
rect 18596 9355 18646 9419
rect 18676 9519 18730 9555
rect 18676 9485 18686 9519
rect 18720 9485 18730 9519
rect 18676 9438 18730 9485
rect 18676 9404 18686 9438
rect 18720 9404 18730 9438
rect 18676 9355 18730 9404
rect 18760 9543 18813 9555
rect 18760 9509 18770 9543
rect 18804 9509 18813 9543
rect 18760 9475 18813 9509
rect 18760 9441 18770 9475
rect 18804 9441 18813 9475
rect 18760 9407 18813 9441
rect 18760 9373 18770 9407
rect 18804 9373 18813 9407
rect 18760 9355 18813 9373
rect 13397 7189 13449 7201
rect 13397 7155 13405 7189
rect 13439 7155 13449 7189
rect 13397 7121 13449 7155
rect 13397 7087 13405 7121
rect 13439 7087 13449 7121
rect 13397 7073 13449 7087
rect 13479 7137 13533 7201
rect 13479 7103 13489 7137
rect 13523 7103 13533 7137
rect 13479 7073 13533 7103
rect 13563 7189 13615 7201
rect 13563 7155 13573 7189
rect 13607 7155 13615 7189
rect 13563 7121 13615 7155
rect 14170 7207 14232 7235
rect 14170 7173 14188 7207
rect 14222 7173 14232 7207
rect 14170 7151 14232 7173
rect 13563 7087 13573 7121
rect 13607 7087 13615 7121
rect 13563 7073 13615 7087
rect 13669 7137 13721 7151
rect 13669 7103 13677 7137
rect 13711 7103 13721 7137
rect 13669 7067 13721 7103
rect 13751 7121 13814 7151
rect 13751 7087 13761 7121
rect 13795 7087 13814 7121
rect 13751 7067 13814 7087
rect 13844 7114 13898 7151
rect 13844 7080 13854 7114
rect 13888 7080 13898 7114
rect 13844 7067 13898 7080
rect 13928 7067 14018 7151
rect 14048 7123 14124 7151
rect 14048 7089 14068 7123
rect 14102 7089 14124 7123
rect 14048 7067 14124 7089
rect 14154 7139 14232 7151
rect 14154 7105 14188 7139
rect 14222 7105 14232 7139
rect 14154 7067 14232 7105
rect 14262 7067 14316 7235
rect 14346 7181 14453 7235
rect 14346 7147 14362 7181
rect 14396 7147 14453 7181
rect 14346 7113 14453 7147
rect 14346 7079 14362 7113
rect 14396 7079 14453 7113
rect 14346 7067 14453 7079
rect 14483 7151 14535 7235
rect 15320 7263 15370 7267
rect 15221 7249 15273 7263
rect 14952 7151 15003 7235
rect 14483 7067 14597 7151
rect 14627 7114 14681 7151
rect 14627 7080 14637 7114
rect 14671 7080 14681 7114
rect 14627 7067 14681 7080
rect 14711 7067 14799 7151
rect 14829 7113 14907 7151
rect 14829 7079 14851 7113
rect 14885 7079 14907 7113
rect 14829 7067 14907 7079
rect 14937 7139 15003 7151
rect 14937 7105 14959 7139
rect 14993 7105 15003 7139
rect 14937 7067 15003 7105
rect 15033 7067 15075 7235
rect 15105 7113 15157 7235
rect 15221 7215 15229 7249
rect 15263 7215 15273 7249
rect 15221 7135 15273 7215
rect 15303 7135 15370 7263
rect 15105 7079 15115 7113
rect 15149 7079 15157 7113
rect 15318 7113 15370 7135
rect 15105 7067 15157 7079
rect 15318 7079 15326 7113
rect 15360 7079 15370 7113
rect 15318 7067 15370 7079
rect 15400 7218 15452 7267
rect 15400 7184 15410 7218
rect 15444 7184 15452 7218
rect 15603 7211 15653 7267
rect 15400 7150 15452 7184
rect 15400 7116 15410 7150
rect 15444 7116 15452 7150
rect 15400 7067 15452 7116
rect 15506 7199 15558 7211
rect 15506 7165 15514 7199
rect 15548 7165 15558 7199
rect 15506 7131 15558 7165
rect 15506 7097 15514 7131
rect 15548 7097 15558 7131
rect 15506 7083 15558 7097
rect 15588 7193 15653 7211
rect 15588 7159 15609 7193
rect 15643 7159 15653 7193
rect 15588 7125 15653 7159
rect 15588 7091 15609 7125
rect 15643 7091 15653 7125
rect 15588 7083 15653 7091
rect 15603 7067 15653 7083
rect 15683 7217 15735 7267
rect 15683 7183 15693 7217
rect 15727 7183 15735 7217
rect 15683 7149 15735 7183
rect 15683 7115 15693 7149
rect 15727 7115 15735 7149
rect 15683 7067 15735 7115
rect 15789 7189 15841 7201
rect 15789 7155 15797 7189
rect 15831 7155 15841 7189
rect 15789 7121 15841 7155
rect 15789 7087 15797 7121
rect 15831 7087 15841 7121
rect 15789 7073 15841 7087
rect 15871 7137 15925 7201
rect 15871 7103 15881 7137
rect 15915 7103 15925 7137
rect 15871 7073 15925 7103
rect 15955 7189 16007 7201
rect 15955 7155 15965 7189
rect 15999 7155 16007 7189
rect 15955 7121 16007 7155
rect 16562 7207 16624 7235
rect 16562 7173 16580 7207
rect 16614 7173 16624 7207
rect 16562 7151 16624 7173
rect 15955 7087 15965 7121
rect 15999 7087 16007 7121
rect 15955 7073 16007 7087
rect 16061 7137 16113 7151
rect 16061 7103 16069 7137
rect 16103 7103 16113 7137
rect 16061 7067 16113 7103
rect 16143 7121 16206 7151
rect 16143 7087 16153 7121
rect 16187 7087 16206 7121
rect 16143 7067 16206 7087
rect 16236 7114 16290 7151
rect 16236 7080 16246 7114
rect 16280 7080 16290 7114
rect 16236 7067 16290 7080
rect 16320 7067 16410 7151
rect 16440 7123 16516 7151
rect 16440 7089 16460 7123
rect 16494 7089 16516 7123
rect 16440 7067 16516 7089
rect 16546 7139 16624 7151
rect 16546 7105 16580 7139
rect 16614 7105 16624 7139
rect 16546 7067 16624 7105
rect 16654 7067 16708 7235
rect 16738 7181 16845 7235
rect 16738 7147 16754 7181
rect 16788 7147 16845 7181
rect 16738 7113 16845 7147
rect 16738 7079 16754 7113
rect 16788 7079 16845 7113
rect 16738 7067 16845 7079
rect 16875 7151 16927 7235
rect 17712 7263 17762 7267
rect 17613 7249 17665 7263
rect 17344 7151 17395 7235
rect 16875 7067 16989 7151
rect 17019 7114 17073 7151
rect 17019 7080 17029 7114
rect 17063 7080 17073 7114
rect 17019 7067 17073 7080
rect 17103 7067 17191 7151
rect 17221 7113 17299 7151
rect 17221 7079 17243 7113
rect 17277 7079 17299 7113
rect 17221 7067 17299 7079
rect 17329 7139 17395 7151
rect 17329 7105 17351 7139
rect 17385 7105 17395 7139
rect 17329 7067 17395 7105
rect 17425 7067 17467 7235
rect 17497 7113 17549 7235
rect 17613 7215 17621 7249
rect 17655 7215 17665 7249
rect 17613 7135 17665 7215
rect 17695 7135 17762 7263
rect 17497 7079 17507 7113
rect 17541 7079 17549 7113
rect 17710 7113 17762 7135
rect 17497 7067 17549 7079
rect 17710 7079 17718 7113
rect 17752 7079 17762 7113
rect 17710 7067 17762 7079
rect 17792 7218 17844 7267
rect 17792 7184 17802 7218
rect 17836 7184 17844 7218
rect 17995 7211 18045 7267
rect 17792 7150 17844 7184
rect 17792 7116 17802 7150
rect 17836 7116 17844 7150
rect 17792 7067 17844 7116
rect 17898 7199 17950 7211
rect 17898 7165 17906 7199
rect 17940 7165 17950 7199
rect 17898 7131 17950 7165
rect 17898 7097 17906 7131
rect 17940 7097 17950 7131
rect 17898 7083 17950 7097
rect 17980 7193 18045 7211
rect 17980 7159 18001 7193
rect 18035 7159 18045 7193
rect 17980 7125 18045 7159
rect 17980 7091 18001 7125
rect 18035 7091 18045 7125
rect 17980 7083 18045 7091
rect 17995 7067 18045 7083
rect 18075 7217 18127 7267
rect 18075 7183 18085 7217
rect 18119 7183 18127 7217
rect 18075 7149 18127 7183
rect 18075 7115 18085 7149
rect 18119 7115 18127 7149
rect 18075 7067 18127 7115
rect 13397 6857 13449 6871
rect 13397 6823 13405 6857
rect 13439 6823 13449 6857
rect 13397 6789 13449 6823
rect 13397 6755 13405 6789
rect 13439 6755 13449 6789
rect 13397 6743 13449 6755
rect 13479 6841 13533 6871
rect 13479 6807 13489 6841
rect 13523 6807 13533 6841
rect 13479 6743 13533 6807
rect 13563 6857 13615 6871
rect 13563 6823 13573 6857
rect 13607 6823 13615 6857
rect 13563 6789 13615 6823
rect 13669 6841 13721 6877
rect 13669 6807 13677 6841
rect 13711 6807 13721 6841
rect 13669 6793 13721 6807
rect 13751 6857 13814 6877
rect 13751 6823 13761 6857
rect 13795 6823 13814 6857
rect 13751 6793 13814 6823
rect 13844 6864 13898 6877
rect 13844 6830 13854 6864
rect 13888 6830 13898 6864
rect 13844 6793 13898 6830
rect 13928 6793 14018 6877
rect 14048 6855 14124 6877
rect 14048 6821 14068 6855
rect 14102 6821 14124 6855
rect 14048 6793 14124 6821
rect 14154 6839 14232 6877
rect 14154 6805 14188 6839
rect 14222 6805 14232 6839
rect 14154 6793 14232 6805
rect 13563 6755 13573 6789
rect 13607 6755 13615 6789
rect 13563 6743 13615 6755
rect 14170 6771 14232 6793
rect 14170 6737 14188 6771
rect 14222 6737 14232 6771
rect 14170 6709 14232 6737
rect 14262 6709 14316 6877
rect 14346 6865 14453 6877
rect 14346 6831 14362 6865
rect 14396 6831 14453 6865
rect 14346 6797 14453 6831
rect 14346 6763 14362 6797
rect 14396 6763 14453 6797
rect 14346 6709 14453 6763
rect 14483 6793 14597 6877
rect 14627 6864 14681 6877
rect 14627 6830 14637 6864
rect 14671 6830 14681 6864
rect 14627 6793 14681 6830
rect 14711 6793 14799 6877
rect 14829 6865 14907 6877
rect 14829 6831 14851 6865
rect 14885 6831 14907 6865
rect 14829 6793 14907 6831
rect 14937 6839 15003 6877
rect 14937 6805 14959 6839
rect 14993 6805 15003 6839
rect 14937 6793 15003 6805
rect 14483 6709 14535 6793
rect 14952 6709 15003 6793
rect 15033 6709 15075 6877
rect 15105 6865 15157 6877
rect 15105 6831 15115 6865
rect 15149 6831 15157 6865
rect 15318 6865 15370 6877
rect 15105 6709 15157 6831
rect 15318 6831 15326 6865
rect 15360 6831 15370 6865
rect 15318 6809 15370 6831
rect 15221 6729 15273 6809
rect 15221 6695 15229 6729
rect 15263 6695 15273 6729
rect 15221 6681 15273 6695
rect 15303 6681 15370 6809
rect 15320 6677 15370 6681
rect 15400 6828 15452 6877
rect 15603 6861 15653 6877
rect 15400 6794 15410 6828
rect 15444 6794 15452 6828
rect 15400 6760 15452 6794
rect 15400 6726 15410 6760
rect 15444 6726 15452 6760
rect 15506 6847 15558 6861
rect 15506 6813 15514 6847
rect 15548 6813 15558 6847
rect 15506 6779 15558 6813
rect 15506 6745 15514 6779
rect 15548 6745 15558 6779
rect 15506 6733 15558 6745
rect 15588 6853 15653 6861
rect 15588 6819 15609 6853
rect 15643 6819 15653 6853
rect 15588 6785 15653 6819
rect 15588 6751 15609 6785
rect 15643 6751 15653 6785
rect 15588 6733 15653 6751
rect 15400 6677 15452 6726
rect 15603 6677 15653 6733
rect 15683 6829 15735 6877
rect 15683 6795 15693 6829
rect 15727 6795 15735 6829
rect 15683 6761 15735 6795
rect 15683 6727 15693 6761
rect 15727 6727 15735 6761
rect 15789 6857 15841 6871
rect 15789 6823 15797 6857
rect 15831 6823 15841 6857
rect 15789 6789 15841 6823
rect 15789 6755 15797 6789
rect 15831 6755 15841 6789
rect 15789 6743 15841 6755
rect 15871 6841 15925 6871
rect 15871 6807 15881 6841
rect 15915 6807 15925 6841
rect 15871 6743 15925 6807
rect 15955 6857 16007 6871
rect 15955 6823 15965 6857
rect 15999 6823 16007 6857
rect 15955 6789 16007 6823
rect 16061 6841 16113 6877
rect 16061 6807 16069 6841
rect 16103 6807 16113 6841
rect 16061 6793 16113 6807
rect 16143 6857 16206 6877
rect 16143 6823 16153 6857
rect 16187 6823 16206 6857
rect 16143 6793 16206 6823
rect 16236 6864 16290 6877
rect 16236 6830 16246 6864
rect 16280 6830 16290 6864
rect 16236 6793 16290 6830
rect 16320 6793 16410 6877
rect 16440 6855 16516 6877
rect 16440 6821 16460 6855
rect 16494 6821 16516 6855
rect 16440 6793 16516 6821
rect 16546 6839 16624 6877
rect 16546 6805 16580 6839
rect 16614 6805 16624 6839
rect 16546 6793 16624 6805
rect 15955 6755 15965 6789
rect 15999 6755 16007 6789
rect 15955 6743 16007 6755
rect 15683 6677 15735 6727
rect 16562 6771 16624 6793
rect 16562 6737 16580 6771
rect 16614 6737 16624 6771
rect 16562 6709 16624 6737
rect 16654 6709 16708 6877
rect 16738 6865 16845 6877
rect 16738 6831 16754 6865
rect 16788 6831 16845 6865
rect 16738 6797 16845 6831
rect 16738 6763 16754 6797
rect 16788 6763 16845 6797
rect 16738 6709 16845 6763
rect 16875 6793 16989 6877
rect 17019 6864 17073 6877
rect 17019 6830 17029 6864
rect 17063 6830 17073 6864
rect 17019 6793 17073 6830
rect 17103 6793 17191 6877
rect 17221 6865 17299 6877
rect 17221 6831 17243 6865
rect 17277 6831 17299 6865
rect 17221 6793 17299 6831
rect 17329 6839 17395 6877
rect 17329 6805 17351 6839
rect 17385 6805 17395 6839
rect 17329 6793 17395 6805
rect 16875 6709 16927 6793
rect 17344 6709 17395 6793
rect 17425 6709 17467 6877
rect 17497 6865 17549 6877
rect 17497 6831 17507 6865
rect 17541 6831 17549 6865
rect 17710 6865 17762 6877
rect 17497 6709 17549 6831
rect 17710 6831 17718 6865
rect 17752 6831 17762 6865
rect 17710 6809 17762 6831
rect 17613 6729 17665 6809
rect 17613 6695 17621 6729
rect 17655 6695 17665 6729
rect 17613 6681 17665 6695
rect 17695 6681 17762 6809
rect 17712 6677 17762 6681
rect 17792 6828 17844 6877
rect 17995 6861 18045 6877
rect 17792 6794 17802 6828
rect 17836 6794 17844 6828
rect 17792 6760 17844 6794
rect 17792 6726 17802 6760
rect 17836 6726 17844 6760
rect 17898 6847 17950 6861
rect 17898 6813 17906 6847
rect 17940 6813 17950 6847
rect 17898 6779 17950 6813
rect 17898 6745 17906 6779
rect 17940 6745 17950 6779
rect 17898 6733 17950 6745
rect 17980 6853 18045 6861
rect 17980 6819 18001 6853
rect 18035 6819 18045 6853
rect 17980 6785 18045 6819
rect 17980 6751 18001 6785
rect 18035 6751 18045 6785
rect 17980 6733 18045 6751
rect 17792 6677 17844 6726
rect 17995 6677 18045 6733
rect 18075 6829 18127 6877
rect 18075 6795 18085 6829
rect 18119 6795 18127 6829
rect 18075 6761 18127 6795
rect 18075 6727 18085 6761
rect 18119 6727 18127 6761
rect 18075 6677 18127 6727
rect 13397 5909 13449 5921
rect 13397 5875 13405 5909
rect 13439 5875 13449 5909
rect 13397 5841 13449 5875
rect 13397 5807 13405 5841
rect 13439 5807 13449 5841
rect 13397 5793 13449 5807
rect 13479 5857 13533 5921
rect 13479 5823 13489 5857
rect 13523 5823 13533 5857
rect 13479 5793 13533 5823
rect 13563 5909 13615 5921
rect 13563 5875 13573 5909
rect 13607 5875 13615 5909
rect 13563 5841 13615 5875
rect 14170 5927 14232 5955
rect 14170 5893 14188 5927
rect 14222 5893 14232 5927
rect 14170 5871 14232 5893
rect 13563 5807 13573 5841
rect 13607 5807 13615 5841
rect 13563 5793 13615 5807
rect 13669 5857 13721 5871
rect 13669 5823 13677 5857
rect 13711 5823 13721 5857
rect 13669 5787 13721 5823
rect 13751 5841 13814 5871
rect 13751 5807 13761 5841
rect 13795 5807 13814 5841
rect 13751 5787 13814 5807
rect 13844 5834 13898 5871
rect 13844 5800 13854 5834
rect 13888 5800 13898 5834
rect 13844 5787 13898 5800
rect 13928 5787 14018 5871
rect 14048 5843 14124 5871
rect 14048 5809 14068 5843
rect 14102 5809 14124 5843
rect 14048 5787 14124 5809
rect 14154 5859 14232 5871
rect 14154 5825 14188 5859
rect 14222 5825 14232 5859
rect 14154 5787 14232 5825
rect 14262 5787 14316 5955
rect 14346 5901 14453 5955
rect 14346 5867 14362 5901
rect 14396 5867 14453 5901
rect 14346 5833 14453 5867
rect 14346 5799 14362 5833
rect 14396 5799 14453 5833
rect 14346 5787 14453 5799
rect 14483 5871 14535 5955
rect 15320 5983 15370 5987
rect 15221 5969 15273 5983
rect 14952 5871 15003 5955
rect 14483 5787 14597 5871
rect 14627 5834 14681 5871
rect 14627 5800 14637 5834
rect 14671 5800 14681 5834
rect 14627 5787 14681 5800
rect 14711 5787 14799 5871
rect 14829 5833 14907 5871
rect 14829 5799 14851 5833
rect 14885 5799 14907 5833
rect 14829 5787 14907 5799
rect 14937 5859 15003 5871
rect 14937 5825 14959 5859
rect 14993 5825 15003 5859
rect 14937 5787 15003 5825
rect 15033 5787 15075 5955
rect 15105 5833 15157 5955
rect 15221 5935 15229 5969
rect 15263 5935 15273 5969
rect 15221 5855 15273 5935
rect 15303 5855 15370 5983
rect 15105 5799 15115 5833
rect 15149 5799 15157 5833
rect 15318 5833 15370 5855
rect 15105 5787 15157 5799
rect 15318 5799 15326 5833
rect 15360 5799 15370 5833
rect 15318 5787 15370 5799
rect 15400 5938 15452 5987
rect 15400 5904 15410 5938
rect 15444 5904 15452 5938
rect 15603 5931 15653 5987
rect 15400 5870 15452 5904
rect 15400 5836 15410 5870
rect 15444 5836 15452 5870
rect 15400 5787 15452 5836
rect 15506 5919 15558 5931
rect 15506 5885 15514 5919
rect 15548 5885 15558 5919
rect 15506 5851 15558 5885
rect 15506 5817 15514 5851
rect 15548 5817 15558 5851
rect 15506 5803 15558 5817
rect 15588 5913 15653 5931
rect 15588 5879 15609 5913
rect 15643 5879 15653 5913
rect 15588 5845 15653 5879
rect 15588 5811 15609 5845
rect 15643 5811 15653 5845
rect 15588 5803 15653 5811
rect 15603 5787 15653 5803
rect 15683 5937 15735 5987
rect 15683 5903 15693 5937
rect 15727 5903 15735 5937
rect 15683 5869 15735 5903
rect 15683 5835 15693 5869
rect 15727 5835 15735 5869
rect 15683 5787 15735 5835
rect 15789 5909 15841 5921
rect 15789 5875 15797 5909
rect 15831 5875 15841 5909
rect 15789 5841 15841 5875
rect 15789 5807 15797 5841
rect 15831 5807 15841 5841
rect 15789 5793 15841 5807
rect 15871 5857 15925 5921
rect 15871 5823 15881 5857
rect 15915 5823 15925 5857
rect 15871 5793 15925 5823
rect 15955 5909 16007 5921
rect 15955 5875 15965 5909
rect 15999 5875 16007 5909
rect 15955 5841 16007 5875
rect 16562 5927 16624 5955
rect 16562 5893 16580 5927
rect 16614 5893 16624 5927
rect 16562 5871 16624 5893
rect 15955 5807 15965 5841
rect 15999 5807 16007 5841
rect 15955 5793 16007 5807
rect 16061 5857 16113 5871
rect 16061 5823 16069 5857
rect 16103 5823 16113 5857
rect 16061 5787 16113 5823
rect 16143 5841 16206 5871
rect 16143 5807 16153 5841
rect 16187 5807 16206 5841
rect 16143 5787 16206 5807
rect 16236 5834 16290 5871
rect 16236 5800 16246 5834
rect 16280 5800 16290 5834
rect 16236 5787 16290 5800
rect 16320 5787 16410 5871
rect 16440 5843 16516 5871
rect 16440 5809 16460 5843
rect 16494 5809 16516 5843
rect 16440 5787 16516 5809
rect 16546 5859 16624 5871
rect 16546 5825 16580 5859
rect 16614 5825 16624 5859
rect 16546 5787 16624 5825
rect 16654 5787 16708 5955
rect 16738 5901 16845 5955
rect 16738 5867 16754 5901
rect 16788 5867 16845 5901
rect 16738 5833 16845 5867
rect 16738 5799 16754 5833
rect 16788 5799 16845 5833
rect 16738 5787 16845 5799
rect 16875 5871 16927 5955
rect 17712 5983 17762 5987
rect 17613 5969 17665 5983
rect 17344 5871 17395 5955
rect 16875 5787 16989 5871
rect 17019 5834 17073 5871
rect 17019 5800 17029 5834
rect 17063 5800 17073 5834
rect 17019 5787 17073 5800
rect 17103 5787 17191 5871
rect 17221 5833 17299 5871
rect 17221 5799 17243 5833
rect 17277 5799 17299 5833
rect 17221 5787 17299 5799
rect 17329 5859 17395 5871
rect 17329 5825 17351 5859
rect 17385 5825 17395 5859
rect 17329 5787 17395 5825
rect 17425 5787 17467 5955
rect 17497 5833 17549 5955
rect 17613 5935 17621 5969
rect 17655 5935 17665 5969
rect 17613 5855 17665 5935
rect 17695 5855 17762 5983
rect 17497 5799 17507 5833
rect 17541 5799 17549 5833
rect 17710 5833 17762 5855
rect 17497 5787 17549 5799
rect 17710 5799 17718 5833
rect 17752 5799 17762 5833
rect 17710 5787 17762 5799
rect 17792 5938 17844 5987
rect 17792 5904 17802 5938
rect 17836 5904 17844 5938
rect 17995 5931 18045 5987
rect 17792 5870 17844 5904
rect 17792 5836 17802 5870
rect 17836 5836 17844 5870
rect 17792 5787 17844 5836
rect 17898 5919 17950 5931
rect 17898 5885 17906 5919
rect 17940 5885 17950 5919
rect 17898 5851 17950 5885
rect 17898 5817 17906 5851
rect 17940 5817 17950 5851
rect 17898 5803 17950 5817
rect 17980 5913 18045 5931
rect 17980 5879 18001 5913
rect 18035 5879 18045 5913
rect 17980 5845 18045 5879
rect 17980 5811 18001 5845
rect 18035 5811 18045 5845
rect 17980 5803 18045 5811
rect 17995 5787 18045 5803
rect 18075 5937 18127 5987
rect 18075 5903 18085 5937
rect 18119 5903 18127 5937
rect 18075 5869 18127 5903
rect 18075 5835 18085 5869
rect 18119 5835 18127 5869
rect 18075 5787 18127 5835
rect 13397 5577 13449 5591
rect 13397 5543 13405 5577
rect 13439 5543 13449 5577
rect 13397 5509 13449 5543
rect 13397 5475 13405 5509
rect 13439 5475 13449 5509
rect 13397 5463 13449 5475
rect 13479 5561 13533 5591
rect 13479 5527 13489 5561
rect 13523 5527 13533 5561
rect 13479 5463 13533 5527
rect 13563 5577 13615 5591
rect 13563 5543 13573 5577
rect 13607 5543 13615 5577
rect 13563 5509 13615 5543
rect 13669 5561 13721 5597
rect 13669 5527 13677 5561
rect 13711 5527 13721 5561
rect 13669 5513 13721 5527
rect 13751 5577 13814 5597
rect 13751 5543 13761 5577
rect 13795 5543 13814 5577
rect 13751 5513 13814 5543
rect 13844 5584 13898 5597
rect 13844 5550 13854 5584
rect 13888 5550 13898 5584
rect 13844 5513 13898 5550
rect 13928 5513 14018 5597
rect 14048 5575 14124 5597
rect 14048 5541 14068 5575
rect 14102 5541 14124 5575
rect 14048 5513 14124 5541
rect 14154 5559 14232 5597
rect 14154 5525 14188 5559
rect 14222 5525 14232 5559
rect 14154 5513 14232 5525
rect 13563 5475 13573 5509
rect 13607 5475 13615 5509
rect 13563 5463 13615 5475
rect 14170 5491 14232 5513
rect 14170 5457 14188 5491
rect 14222 5457 14232 5491
rect 14170 5429 14232 5457
rect 14262 5429 14316 5597
rect 14346 5585 14453 5597
rect 14346 5551 14362 5585
rect 14396 5551 14453 5585
rect 14346 5517 14453 5551
rect 14346 5483 14362 5517
rect 14396 5483 14453 5517
rect 14346 5429 14453 5483
rect 14483 5513 14597 5597
rect 14627 5584 14681 5597
rect 14627 5550 14637 5584
rect 14671 5550 14681 5584
rect 14627 5513 14681 5550
rect 14711 5513 14799 5597
rect 14829 5585 14907 5597
rect 14829 5551 14851 5585
rect 14885 5551 14907 5585
rect 14829 5513 14907 5551
rect 14937 5559 15003 5597
rect 14937 5525 14959 5559
rect 14993 5525 15003 5559
rect 14937 5513 15003 5525
rect 14483 5429 14535 5513
rect 14952 5429 15003 5513
rect 15033 5429 15075 5597
rect 15105 5585 15157 5597
rect 15105 5551 15115 5585
rect 15149 5551 15157 5585
rect 15318 5585 15370 5597
rect 15105 5429 15157 5551
rect 15318 5551 15326 5585
rect 15360 5551 15370 5585
rect 15318 5529 15370 5551
rect 15221 5449 15273 5529
rect 15221 5415 15229 5449
rect 15263 5415 15273 5449
rect 15221 5401 15273 5415
rect 15303 5401 15370 5529
rect 15320 5397 15370 5401
rect 15400 5548 15452 5597
rect 15603 5581 15653 5597
rect 15400 5514 15410 5548
rect 15444 5514 15452 5548
rect 15400 5480 15452 5514
rect 15400 5446 15410 5480
rect 15444 5446 15452 5480
rect 15506 5567 15558 5581
rect 15506 5533 15514 5567
rect 15548 5533 15558 5567
rect 15506 5499 15558 5533
rect 15506 5465 15514 5499
rect 15548 5465 15558 5499
rect 15506 5453 15558 5465
rect 15588 5573 15653 5581
rect 15588 5539 15609 5573
rect 15643 5539 15653 5573
rect 15588 5505 15653 5539
rect 15588 5471 15609 5505
rect 15643 5471 15653 5505
rect 15588 5453 15653 5471
rect 15400 5397 15452 5446
rect 15603 5397 15653 5453
rect 15683 5549 15735 5597
rect 15683 5515 15693 5549
rect 15727 5515 15735 5549
rect 15683 5481 15735 5515
rect 15683 5447 15693 5481
rect 15727 5447 15735 5481
rect 15789 5577 15841 5591
rect 15789 5543 15797 5577
rect 15831 5543 15841 5577
rect 15789 5509 15841 5543
rect 15789 5475 15797 5509
rect 15831 5475 15841 5509
rect 15789 5463 15841 5475
rect 15871 5561 15925 5591
rect 15871 5527 15881 5561
rect 15915 5527 15925 5561
rect 15871 5463 15925 5527
rect 15955 5577 16007 5591
rect 15955 5543 15965 5577
rect 15999 5543 16007 5577
rect 15955 5509 16007 5543
rect 16061 5561 16113 5597
rect 16061 5527 16069 5561
rect 16103 5527 16113 5561
rect 16061 5513 16113 5527
rect 16143 5577 16206 5597
rect 16143 5543 16153 5577
rect 16187 5543 16206 5577
rect 16143 5513 16206 5543
rect 16236 5584 16290 5597
rect 16236 5550 16246 5584
rect 16280 5550 16290 5584
rect 16236 5513 16290 5550
rect 16320 5513 16410 5597
rect 16440 5575 16516 5597
rect 16440 5541 16460 5575
rect 16494 5541 16516 5575
rect 16440 5513 16516 5541
rect 16546 5559 16624 5597
rect 16546 5525 16580 5559
rect 16614 5525 16624 5559
rect 16546 5513 16624 5525
rect 15955 5475 15965 5509
rect 15999 5475 16007 5509
rect 15955 5463 16007 5475
rect 15683 5397 15735 5447
rect 16562 5491 16624 5513
rect 16562 5457 16580 5491
rect 16614 5457 16624 5491
rect 16562 5429 16624 5457
rect 16654 5429 16708 5597
rect 16738 5585 16845 5597
rect 16738 5551 16754 5585
rect 16788 5551 16845 5585
rect 16738 5517 16845 5551
rect 16738 5483 16754 5517
rect 16788 5483 16845 5517
rect 16738 5429 16845 5483
rect 16875 5513 16989 5597
rect 17019 5584 17073 5597
rect 17019 5550 17029 5584
rect 17063 5550 17073 5584
rect 17019 5513 17073 5550
rect 17103 5513 17191 5597
rect 17221 5585 17299 5597
rect 17221 5551 17243 5585
rect 17277 5551 17299 5585
rect 17221 5513 17299 5551
rect 17329 5559 17395 5597
rect 17329 5525 17351 5559
rect 17385 5525 17395 5559
rect 17329 5513 17395 5525
rect 16875 5429 16927 5513
rect 17344 5429 17395 5513
rect 17425 5429 17467 5597
rect 17497 5585 17549 5597
rect 17497 5551 17507 5585
rect 17541 5551 17549 5585
rect 17710 5585 17762 5597
rect 17497 5429 17549 5551
rect 17710 5551 17718 5585
rect 17752 5551 17762 5585
rect 17710 5529 17762 5551
rect 17613 5449 17665 5529
rect 17613 5415 17621 5449
rect 17655 5415 17665 5449
rect 17613 5401 17665 5415
rect 17695 5401 17762 5529
rect 17712 5397 17762 5401
rect 17792 5548 17844 5597
rect 17995 5581 18045 5597
rect 17792 5514 17802 5548
rect 17836 5514 17844 5548
rect 17792 5480 17844 5514
rect 17792 5446 17802 5480
rect 17836 5446 17844 5480
rect 17898 5567 17950 5581
rect 17898 5533 17906 5567
rect 17940 5533 17950 5567
rect 17898 5499 17950 5533
rect 17898 5465 17906 5499
rect 17940 5465 17950 5499
rect 17898 5453 17950 5465
rect 17980 5573 18045 5581
rect 17980 5539 18001 5573
rect 18035 5539 18045 5573
rect 17980 5505 18045 5539
rect 17980 5471 18001 5505
rect 18035 5471 18045 5505
rect 17980 5453 18045 5471
rect 17792 5397 17844 5446
rect 17995 5397 18045 5453
rect 18075 5549 18127 5597
rect 18075 5515 18085 5549
rect 18119 5515 18127 5549
rect 18075 5481 18127 5515
rect 18075 5447 18085 5481
rect 18119 5447 18127 5481
rect 18075 5397 18127 5447
<< ndiffc >>
rect 11868 9566 11902 9600
rect 11868 9498 11902 9532
rect 11952 9566 11986 9600
rect 11952 9498 11986 9532
rect 12058 9566 12092 9600
rect 12058 9498 12092 9532
rect 12142 9566 12176 9600
rect 12142 9498 12176 9532
rect 13329 9164 13363 9224
rect 13419 9164 13453 9224
rect 14061 9164 14095 9224
rect 14168 9164 14202 9224
rect 14271 9164 14305 9224
rect 15273 9164 15307 9224
rect 15379 9164 15413 9224
rect 15483 9164 15517 9224
rect 16611 9164 16645 9224
rect 16719 9164 16753 9224
rect 16821 9164 16855 9224
rect 17466 9164 17500 9224
rect 17555 9164 17589 9224
rect 18119 9165 18153 9225
rect 18207 9165 18241 9225
rect 18303 9165 18337 9225
rect 18399 9165 18433 9225
rect 18507 9130 18541 9164
rect 18600 9117 18634 9151
rect 18686 9147 18720 9181
rect 18770 9189 18804 9223
rect 18770 9121 18804 9155
rect 12309 8980 12343 9040
rect 12469 8980 12503 9040
rect 18119 9027 18153 9087
rect 18207 9027 18241 9087
rect 12309 8842 12343 8902
rect 12469 8842 12503 8902
rect 12309 8704 12343 8764
rect 12469 8704 12503 8764
rect 12309 8566 12343 8626
rect 12469 8566 12503 8626
rect 12309 8428 12343 8488
rect 12469 8428 12503 8488
rect 12309 8290 12343 8350
rect 12469 8290 12503 8350
rect 12309 8152 12343 8212
rect 12469 8152 12503 8212
rect 12309 8014 12343 8074
rect 12469 8014 12503 8074
rect 13405 7445 13439 7479
rect 13489 7471 13523 7505
rect 13573 7445 13607 7479
rect 13677 7471 13711 7505
rect 13761 7453 13795 7487
rect 13867 7471 13901 7505
rect 14084 7475 14118 7509
rect 14168 7455 14202 7489
rect 14268 7411 14302 7445
rect 14352 7437 14386 7471
rect 14456 7471 14490 7505
rect 14650 7471 14684 7505
rect 14841 7475 14875 7509
rect 14943 7455 14977 7489
rect 15043 7411 15077 7445
rect 15127 7463 15161 7497
rect 15231 7461 15265 7495
rect 15326 7471 15360 7505
rect 15410 7437 15444 7471
rect 15514 7445 15548 7479
rect 15609 7471 15643 7505
rect 15693 7435 15727 7469
rect 15797 7445 15831 7479
rect 15881 7471 15915 7505
rect 15965 7445 15999 7479
rect 16069 7471 16103 7505
rect 16153 7453 16187 7487
rect 16259 7471 16293 7505
rect 16476 7475 16510 7509
rect 16560 7455 16594 7489
rect 16660 7411 16694 7445
rect 16744 7437 16778 7471
rect 16848 7471 16882 7505
rect 17042 7471 17076 7505
rect 17233 7475 17267 7509
rect 17335 7455 17369 7489
rect 17435 7411 17469 7445
rect 17519 7463 17553 7497
rect 17623 7461 17657 7495
rect 17718 7471 17752 7505
rect 17802 7437 17836 7471
rect 17906 7445 17940 7479
rect 18001 7471 18035 7505
rect 18085 7435 18119 7469
rect 13405 6465 13439 6499
rect 13489 6439 13523 6473
rect 13573 6465 13607 6499
rect 13677 6439 13711 6473
rect 13761 6457 13795 6491
rect 13867 6439 13901 6473
rect 14084 6435 14118 6469
rect 14168 6455 14202 6489
rect 14268 6499 14302 6533
rect 14352 6473 14386 6507
rect 14456 6439 14490 6473
rect 14650 6439 14684 6473
rect 14841 6435 14875 6469
rect 14943 6455 14977 6489
rect 15043 6499 15077 6533
rect 15127 6447 15161 6481
rect 15231 6449 15265 6483
rect 15326 6439 15360 6473
rect 15410 6473 15444 6507
rect 15514 6465 15548 6499
rect 15609 6439 15643 6473
rect 15693 6475 15727 6509
rect 15797 6465 15831 6499
rect 15881 6439 15915 6473
rect 15965 6465 15999 6499
rect 16069 6439 16103 6473
rect 16153 6457 16187 6491
rect 16259 6439 16293 6473
rect 16476 6435 16510 6469
rect 16560 6455 16594 6489
rect 16660 6499 16694 6533
rect 16744 6473 16778 6507
rect 16848 6439 16882 6473
rect 17042 6439 17076 6473
rect 17233 6435 17267 6469
rect 17335 6455 17369 6489
rect 17435 6499 17469 6533
rect 17519 6447 17553 6481
rect 17623 6449 17657 6483
rect 17718 6439 17752 6473
rect 17802 6473 17836 6507
rect 17906 6465 17940 6499
rect 18001 6439 18035 6473
rect 18085 6475 18119 6509
rect 13405 6165 13439 6199
rect 13489 6191 13523 6225
rect 13573 6165 13607 6199
rect 13677 6191 13711 6225
rect 13761 6173 13795 6207
rect 13867 6191 13901 6225
rect 14084 6195 14118 6229
rect 14168 6175 14202 6209
rect 14268 6131 14302 6165
rect 14352 6157 14386 6191
rect 14456 6191 14490 6225
rect 14650 6191 14684 6225
rect 14841 6195 14875 6229
rect 14943 6175 14977 6209
rect 15043 6131 15077 6165
rect 15127 6183 15161 6217
rect 15231 6181 15265 6215
rect 15326 6191 15360 6225
rect 15410 6157 15444 6191
rect 15514 6165 15548 6199
rect 15609 6191 15643 6225
rect 15693 6155 15727 6189
rect 15797 6165 15831 6199
rect 15881 6191 15915 6225
rect 15965 6165 15999 6199
rect 16069 6191 16103 6225
rect 16153 6173 16187 6207
rect 16259 6191 16293 6225
rect 16476 6195 16510 6229
rect 16560 6175 16594 6209
rect 16660 6131 16694 6165
rect 16744 6157 16778 6191
rect 16848 6191 16882 6225
rect 17042 6191 17076 6225
rect 17233 6195 17267 6229
rect 17335 6175 17369 6209
rect 17435 6131 17469 6165
rect 17519 6183 17553 6217
rect 17623 6181 17657 6215
rect 17718 6191 17752 6225
rect 17802 6157 17836 6191
rect 17906 6165 17940 6199
rect 18001 6191 18035 6225
rect 18085 6155 18119 6189
rect 13405 5185 13439 5219
rect 13489 5159 13523 5193
rect 13573 5185 13607 5219
rect 13677 5159 13711 5193
rect 13761 5177 13795 5211
rect 13867 5159 13901 5193
rect 14084 5155 14118 5189
rect 14168 5175 14202 5209
rect 14268 5219 14302 5253
rect 14352 5193 14386 5227
rect 14456 5159 14490 5193
rect 14650 5159 14684 5193
rect 14841 5155 14875 5189
rect 14943 5175 14977 5209
rect 15043 5219 15077 5253
rect 15127 5167 15161 5201
rect 15231 5169 15265 5203
rect 15326 5159 15360 5193
rect 15410 5193 15444 5227
rect 15514 5185 15548 5219
rect 15609 5159 15643 5193
rect 15693 5195 15727 5229
rect 15797 5185 15831 5219
rect 15881 5159 15915 5193
rect 15965 5185 15999 5219
rect 16069 5159 16103 5193
rect 16153 5177 16187 5211
rect 16259 5159 16293 5193
rect 16476 5155 16510 5189
rect 16560 5175 16594 5209
rect 16660 5219 16694 5253
rect 16744 5193 16778 5227
rect 16848 5159 16882 5193
rect 17042 5159 17076 5193
rect 17233 5155 17267 5189
rect 17335 5175 17369 5209
rect 17435 5219 17469 5253
rect 17519 5167 17553 5201
rect 17623 5169 17657 5203
rect 17718 5159 17752 5193
rect 17802 5193 17836 5227
rect 17906 5185 17940 5219
rect 18001 5159 18035 5193
rect 18085 5195 18119 5229
<< pdiffc >>
rect 12334 10507 12368 10567
rect 12422 10507 12456 10567
rect 12334 10369 12368 10429
rect 12422 10369 12456 10429
rect 12334 10231 12368 10291
rect 12422 10231 12456 10291
rect 12334 10093 12368 10153
rect 12422 10093 12456 10153
rect 12334 9955 12368 10015
rect 12422 9955 12456 10015
rect 11868 9886 11902 9920
rect 11868 9818 11902 9852
rect 11868 9750 11902 9784
rect 11952 9886 11986 9920
rect 11952 9818 11986 9852
rect 11952 9750 11986 9784
rect 12058 9886 12092 9920
rect 12058 9818 12092 9852
rect 12058 9750 12092 9784
rect 12142 9886 12176 9920
rect 12142 9818 12176 9852
rect 12334 9817 12368 9877
rect 12422 9817 12456 9877
rect 12142 9750 12176 9784
rect 18119 9506 18153 9566
rect 18207 9506 18241 9566
rect 18507 9501 18541 9535
rect 12976 9362 13010 9422
rect 13064 9365 13098 9425
rect 13708 9365 13742 9425
rect 13813 9365 13847 9425
rect 13922 9365 13956 9425
rect 14920 9365 14954 9425
rect 15024 9365 15058 9425
rect 15134 9365 15168 9425
rect 16132 9365 16166 9425
rect 16237 9365 16271 9425
rect 16346 9365 16380 9425
rect 17344 9365 17378 9425
rect 17451 9365 17485 9425
rect 17558 9365 17592 9425
rect 18119 9368 18153 9428
rect 18207 9368 18241 9428
rect 18303 9368 18337 9428
rect 18399 9368 18433 9428
rect 18507 9433 18541 9467
rect 18600 9501 18634 9535
rect 18600 9433 18634 9467
rect 18686 9485 18720 9519
rect 18686 9404 18720 9438
rect 18770 9509 18804 9543
rect 18770 9441 18804 9475
rect 18770 9373 18804 9407
rect 13405 7155 13439 7189
rect 13405 7087 13439 7121
rect 13489 7103 13523 7137
rect 13573 7155 13607 7189
rect 14188 7173 14222 7207
rect 13573 7087 13607 7121
rect 13677 7103 13711 7137
rect 13761 7087 13795 7121
rect 13854 7080 13888 7114
rect 14068 7089 14102 7123
rect 14188 7105 14222 7139
rect 14362 7147 14396 7181
rect 14362 7079 14396 7113
rect 14637 7080 14671 7114
rect 14851 7079 14885 7113
rect 14959 7105 14993 7139
rect 15229 7215 15263 7249
rect 15115 7079 15149 7113
rect 15326 7079 15360 7113
rect 15410 7184 15444 7218
rect 15410 7116 15444 7150
rect 15514 7165 15548 7199
rect 15514 7097 15548 7131
rect 15609 7159 15643 7193
rect 15609 7091 15643 7125
rect 15693 7183 15727 7217
rect 15693 7115 15727 7149
rect 15797 7155 15831 7189
rect 15797 7087 15831 7121
rect 15881 7103 15915 7137
rect 15965 7155 15999 7189
rect 16580 7173 16614 7207
rect 15965 7087 15999 7121
rect 16069 7103 16103 7137
rect 16153 7087 16187 7121
rect 16246 7080 16280 7114
rect 16460 7089 16494 7123
rect 16580 7105 16614 7139
rect 16754 7147 16788 7181
rect 16754 7079 16788 7113
rect 17029 7080 17063 7114
rect 17243 7079 17277 7113
rect 17351 7105 17385 7139
rect 17621 7215 17655 7249
rect 17507 7079 17541 7113
rect 17718 7079 17752 7113
rect 17802 7184 17836 7218
rect 17802 7116 17836 7150
rect 17906 7165 17940 7199
rect 17906 7097 17940 7131
rect 18001 7159 18035 7193
rect 18001 7091 18035 7125
rect 18085 7183 18119 7217
rect 18085 7115 18119 7149
rect 13405 6823 13439 6857
rect 13405 6755 13439 6789
rect 13489 6807 13523 6841
rect 13573 6823 13607 6857
rect 13677 6807 13711 6841
rect 13761 6823 13795 6857
rect 13854 6830 13888 6864
rect 14068 6821 14102 6855
rect 14188 6805 14222 6839
rect 13573 6755 13607 6789
rect 14188 6737 14222 6771
rect 14362 6831 14396 6865
rect 14362 6763 14396 6797
rect 14637 6830 14671 6864
rect 14851 6831 14885 6865
rect 14959 6805 14993 6839
rect 15115 6831 15149 6865
rect 15326 6831 15360 6865
rect 15229 6695 15263 6729
rect 15410 6794 15444 6828
rect 15410 6726 15444 6760
rect 15514 6813 15548 6847
rect 15514 6745 15548 6779
rect 15609 6819 15643 6853
rect 15609 6751 15643 6785
rect 15693 6795 15727 6829
rect 15693 6727 15727 6761
rect 15797 6823 15831 6857
rect 15797 6755 15831 6789
rect 15881 6807 15915 6841
rect 15965 6823 15999 6857
rect 16069 6807 16103 6841
rect 16153 6823 16187 6857
rect 16246 6830 16280 6864
rect 16460 6821 16494 6855
rect 16580 6805 16614 6839
rect 15965 6755 15999 6789
rect 16580 6737 16614 6771
rect 16754 6831 16788 6865
rect 16754 6763 16788 6797
rect 17029 6830 17063 6864
rect 17243 6831 17277 6865
rect 17351 6805 17385 6839
rect 17507 6831 17541 6865
rect 17718 6831 17752 6865
rect 17621 6695 17655 6729
rect 17802 6794 17836 6828
rect 17802 6726 17836 6760
rect 17906 6813 17940 6847
rect 17906 6745 17940 6779
rect 18001 6819 18035 6853
rect 18001 6751 18035 6785
rect 18085 6795 18119 6829
rect 18085 6727 18119 6761
rect 13405 5875 13439 5909
rect 13405 5807 13439 5841
rect 13489 5823 13523 5857
rect 13573 5875 13607 5909
rect 14188 5893 14222 5927
rect 13573 5807 13607 5841
rect 13677 5823 13711 5857
rect 13761 5807 13795 5841
rect 13854 5800 13888 5834
rect 14068 5809 14102 5843
rect 14188 5825 14222 5859
rect 14362 5867 14396 5901
rect 14362 5799 14396 5833
rect 14637 5800 14671 5834
rect 14851 5799 14885 5833
rect 14959 5825 14993 5859
rect 15229 5935 15263 5969
rect 15115 5799 15149 5833
rect 15326 5799 15360 5833
rect 15410 5904 15444 5938
rect 15410 5836 15444 5870
rect 15514 5885 15548 5919
rect 15514 5817 15548 5851
rect 15609 5879 15643 5913
rect 15609 5811 15643 5845
rect 15693 5903 15727 5937
rect 15693 5835 15727 5869
rect 15797 5875 15831 5909
rect 15797 5807 15831 5841
rect 15881 5823 15915 5857
rect 15965 5875 15999 5909
rect 16580 5893 16614 5927
rect 15965 5807 15999 5841
rect 16069 5823 16103 5857
rect 16153 5807 16187 5841
rect 16246 5800 16280 5834
rect 16460 5809 16494 5843
rect 16580 5825 16614 5859
rect 16754 5867 16788 5901
rect 16754 5799 16788 5833
rect 17029 5800 17063 5834
rect 17243 5799 17277 5833
rect 17351 5825 17385 5859
rect 17621 5935 17655 5969
rect 17507 5799 17541 5833
rect 17718 5799 17752 5833
rect 17802 5904 17836 5938
rect 17802 5836 17836 5870
rect 17906 5885 17940 5919
rect 17906 5817 17940 5851
rect 18001 5879 18035 5913
rect 18001 5811 18035 5845
rect 18085 5903 18119 5937
rect 18085 5835 18119 5869
rect 13405 5543 13439 5577
rect 13405 5475 13439 5509
rect 13489 5527 13523 5561
rect 13573 5543 13607 5577
rect 13677 5527 13711 5561
rect 13761 5543 13795 5577
rect 13854 5550 13888 5584
rect 14068 5541 14102 5575
rect 14188 5525 14222 5559
rect 13573 5475 13607 5509
rect 14188 5457 14222 5491
rect 14362 5551 14396 5585
rect 14362 5483 14396 5517
rect 14637 5550 14671 5584
rect 14851 5551 14885 5585
rect 14959 5525 14993 5559
rect 15115 5551 15149 5585
rect 15326 5551 15360 5585
rect 15229 5415 15263 5449
rect 15410 5514 15444 5548
rect 15410 5446 15444 5480
rect 15514 5533 15548 5567
rect 15514 5465 15548 5499
rect 15609 5539 15643 5573
rect 15609 5471 15643 5505
rect 15693 5515 15727 5549
rect 15693 5447 15727 5481
rect 15797 5543 15831 5577
rect 15797 5475 15831 5509
rect 15881 5527 15915 5561
rect 15965 5543 15999 5577
rect 16069 5527 16103 5561
rect 16153 5543 16187 5577
rect 16246 5550 16280 5584
rect 16460 5541 16494 5575
rect 16580 5525 16614 5559
rect 15965 5475 15999 5509
rect 16580 5457 16614 5491
rect 16754 5551 16788 5585
rect 16754 5483 16788 5517
rect 17029 5550 17063 5584
rect 17243 5551 17277 5585
rect 17351 5525 17385 5559
rect 17507 5551 17541 5585
rect 17718 5551 17752 5585
rect 17621 5415 17655 5449
rect 17802 5514 17836 5548
rect 17802 5446 17836 5480
rect 17906 5533 17940 5567
rect 17906 5465 17940 5499
rect 18001 5539 18035 5573
rect 18001 5471 18035 5505
rect 18085 5515 18119 5549
rect 18085 5447 18119 5481
<< psubdiff >>
rect 11862 9389 11886 9423
rect 11920 9389 12004 9423
rect 12038 9389 12148 9423
rect 12182 9389 12224 9423
rect 11862 9387 12224 9389
rect 18473 9040 18593 9041
rect 18473 9006 18501 9040
rect 18535 9007 18593 9040
rect 18627 9007 18685 9041
rect 18719 9007 18778 9041
rect 18812 9007 18842 9041
rect 18535 9006 18842 9007
rect 18473 9005 18842 9006
rect 12586 8198 12690 8233
rect 12586 8164 12617 8198
rect 12651 8164 12690 8198
rect 12586 8135 12690 8164
rect 12984 8027 13316 8043
rect 12984 7993 13010 8027
rect 13044 7993 13090 8027
rect 13124 7993 13170 8027
rect 13204 7993 13250 8027
rect 13284 7993 13316 8027
rect 12984 7975 13316 7993
rect 13716 8027 14048 8043
rect 13716 7993 13742 8027
rect 13776 7993 13822 8027
rect 13856 7993 13902 8027
rect 13936 7993 13982 8027
rect 14016 7993 14048 8027
rect 13716 7975 14048 7993
rect 14318 8027 14650 8043
rect 14318 7993 14350 8027
rect 14384 7993 14430 8027
rect 14464 7993 14510 8027
rect 14544 7993 14590 8027
rect 14624 7993 14650 8027
rect 14318 7975 14650 7993
rect 14928 8027 15260 8043
rect 14928 7993 14954 8027
rect 14988 7993 15034 8027
rect 15068 7993 15114 8027
rect 15148 7993 15194 8027
rect 15228 7993 15260 8027
rect 14928 7975 15260 7993
rect 15530 8027 15862 8043
rect 15530 7993 15562 8027
rect 15596 7993 15642 8027
rect 15676 7993 15722 8027
rect 15756 7993 15802 8027
rect 15836 7993 15862 8027
rect 15530 7975 15862 7993
rect 16266 8027 16598 8043
rect 16266 7993 16292 8027
rect 16326 7993 16372 8027
rect 16406 7993 16452 8027
rect 16486 7993 16532 8027
rect 16566 7993 16598 8027
rect 16266 7975 16598 7993
rect 16868 8027 17200 8043
rect 16868 7993 16900 8027
rect 16934 7993 16980 8027
rect 17014 7993 17060 8027
rect 17094 7993 17140 8027
rect 17174 7993 17200 8027
rect 16868 7975 17200 7993
rect 17602 8027 17934 8043
rect 17602 7993 17634 8027
rect 17668 7993 17714 8027
rect 17748 7993 17794 8027
rect 17828 7993 17874 8027
rect 17908 7993 17934 8027
rect 17602 7975 17934 7993
rect 13370 7581 13399 7615
rect 13433 7581 13491 7615
rect 13525 7581 13583 7615
rect 13617 7581 13675 7615
rect 13709 7581 13767 7615
rect 13801 7581 13859 7615
rect 13893 7581 13951 7615
rect 13985 7581 14043 7615
rect 14077 7581 14135 7615
rect 14169 7581 14226 7615
rect 14260 7581 14319 7615
rect 14353 7581 14411 7615
rect 14445 7581 14503 7615
rect 14537 7581 14595 7615
rect 14629 7581 14687 7615
rect 14721 7581 14779 7615
rect 14813 7581 14871 7615
rect 14905 7581 14963 7615
rect 14997 7581 15055 7615
rect 15089 7581 15147 7615
rect 15181 7581 15239 7615
rect 15273 7581 15331 7615
rect 15365 7581 15423 7615
rect 15457 7581 15515 7615
rect 15549 7581 15607 7615
rect 15641 7581 15699 7615
rect 15733 7581 15791 7615
rect 15825 7581 15883 7615
rect 15917 7581 15975 7615
rect 16009 7581 16067 7615
rect 16101 7581 16159 7615
rect 16193 7581 16251 7615
rect 16285 7581 16343 7615
rect 16377 7581 16435 7615
rect 16469 7581 16527 7615
rect 16561 7581 16619 7615
rect 16653 7581 16711 7615
rect 16745 7581 16803 7615
rect 16837 7581 16895 7615
rect 16929 7581 16987 7615
rect 17021 7581 17079 7615
rect 17113 7581 17171 7615
rect 17205 7581 17263 7615
rect 17297 7581 17355 7615
rect 17389 7581 17447 7615
rect 17481 7581 17539 7615
rect 17573 7581 17631 7615
rect 17665 7581 17723 7615
rect 17757 7581 17815 7615
rect 17849 7581 17907 7615
rect 17941 7581 17999 7615
rect 18033 7581 18091 7615
rect 18125 7581 18154 7615
rect 13370 6316 13399 6350
rect 13433 6316 13491 6350
rect 13525 6316 13583 6350
rect 13617 6316 13675 6350
rect 13709 6316 13767 6350
rect 13801 6316 13859 6350
rect 13893 6316 13951 6350
rect 13985 6316 14043 6350
rect 14077 6316 14135 6350
rect 14169 6316 14227 6350
rect 14261 6316 14319 6350
rect 14353 6316 14411 6350
rect 14445 6316 14503 6350
rect 14537 6316 14595 6350
rect 14629 6316 14687 6350
rect 14721 6316 14779 6350
rect 14813 6316 14871 6350
rect 14905 6316 14964 6350
rect 14998 6316 15055 6350
rect 15089 6316 15147 6350
rect 15181 6316 15239 6350
rect 15273 6316 15332 6350
rect 15366 6316 15423 6350
rect 15457 6316 15515 6350
rect 15549 6316 15607 6350
rect 15641 6316 15699 6350
rect 15733 6316 15791 6350
rect 15825 6316 15883 6350
rect 15917 6316 15975 6350
rect 16009 6316 16067 6350
rect 16101 6316 16159 6350
rect 16193 6316 16251 6350
rect 16285 6316 16343 6350
rect 16377 6316 16435 6350
rect 16469 6316 16526 6350
rect 16560 6316 16618 6350
rect 16652 6316 16711 6350
rect 16745 6316 16803 6350
rect 16837 6316 16895 6350
rect 16929 6316 16986 6350
rect 17020 6316 17079 6350
rect 17113 6316 17170 6350
rect 17204 6316 17263 6350
rect 17297 6316 17355 6350
rect 17389 6316 17447 6350
rect 17481 6316 17539 6350
rect 17573 6316 17631 6350
rect 17665 6316 17723 6350
rect 17757 6316 17815 6350
rect 17849 6316 17907 6350
rect 17941 6316 17999 6350
rect 18033 6316 18091 6350
rect 18125 6316 18154 6350
rect 13370 5049 13399 5083
rect 13433 5049 13491 5083
rect 13525 5049 13583 5083
rect 13617 5049 13675 5083
rect 13709 5049 13767 5083
rect 13801 5049 13859 5083
rect 13893 5049 13951 5083
rect 13985 5049 14043 5083
rect 14077 5049 14135 5083
rect 14169 5049 14227 5083
rect 14261 5049 14319 5083
rect 14353 5049 14411 5083
rect 14445 5049 14503 5083
rect 14537 5049 14595 5083
rect 14629 5049 14687 5083
rect 14721 5049 14779 5083
rect 14813 5049 14871 5083
rect 14905 5049 14963 5083
rect 14997 5049 15055 5083
rect 15089 5049 15147 5083
rect 15181 5049 15239 5083
rect 15273 5049 15331 5083
rect 15365 5049 15423 5083
rect 15457 5049 15515 5083
rect 15549 5049 15607 5083
rect 15641 5049 15699 5083
rect 15733 5049 15791 5083
rect 15825 5049 15883 5083
rect 15917 5049 15975 5083
rect 16009 5049 16067 5083
rect 16101 5049 16159 5083
rect 16193 5049 16251 5083
rect 16285 5049 16343 5083
rect 16377 5049 16435 5083
rect 16469 5049 16527 5083
rect 16561 5049 16619 5083
rect 16653 5049 16711 5083
rect 16745 5049 16803 5083
rect 16837 5049 16895 5083
rect 16929 5049 16987 5083
rect 17021 5049 17079 5083
rect 17113 5049 17171 5083
rect 17205 5049 17263 5083
rect 17297 5049 17355 5083
rect 17389 5049 17447 5083
rect 17481 5049 17539 5083
rect 17573 5049 17631 5083
rect 17665 5049 17723 5083
rect 17757 5049 17815 5083
rect 17849 5049 17907 5083
rect 17941 5049 17999 5083
rect 18033 5049 18091 5083
rect 18125 5049 18154 5083
<< nsubdiff >>
rect 12532 10591 13070 10611
rect 12532 10557 12580 10591
rect 12614 10557 12660 10591
rect 12694 10557 12740 10591
rect 12774 10557 12820 10591
rect 12854 10557 12900 10591
rect 12934 10557 12980 10591
rect 13014 10557 13070 10591
rect 12532 10543 13070 10557
rect 13264 10594 13802 10614
rect 13264 10560 13312 10594
rect 13346 10560 13392 10594
rect 13426 10560 13472 10594
rect 13506 10560 13552 10594
rect 13586 10560 13632 10594
rect 13666 10560 13712 10594
rect 13746 10560 13802 10594
rect 13264 10546 13802 10560
rect 13862 10594 14400 10614
rect 13862 10560 13918 10594
rect 13952 10560 13998 10594
rect 14032 10560 14078 10594
rect 14112 10560 14158 10594
rect 14192 10560 14238 10594
rect 14272 10560 14318 10594
rect 14352 10560 14400 10594
rect 13862 10546 14400 10560
rect 14476 10594 15014 10614
rect 14476 10560 14524 10594
rect 14558 10560 14604 10594
rect 14638 10560 14684 10594
rect 14718 10560 14764 10594
rect 14798 10560 14844 10594
rect 14878 10560 14924 10594
rect 14958 10560 15014 10594
rect 14476 10546 15014 10560
rect 15074 10594 15612 10614
rect 15074 10560 15130 10594
rect 15164 10560 15210 10594
rect 15244 10560 15290 10594
rect 15324 10560 15370 10594
rect 15404 10560 15450 10594
rect 15484 10560 15530 10594
rect 15564 10560 15612 10594
rect 15074 10546 15612 10560
rect 15688 10594 16226 10614
rect 15688 10560 15736 10594
rect 15770 10560 15816 10594
rect 15850 10560 15896 10594
rect 15930 10560 15976 10594
rect 16010 10560 16056 10594
rect 16090 10560 16136 10594
rect 16170 10560 16226 10594
rect 15688 10546 16226 10560
rect 16286 10594 16824 10614
rect 16286 10560 16342 10594
rect 16376 10560 16422 10594
rect 16456 10560 16502 10594
rect 16536 10560 16582 10594
rect 16616 10560 16662 10594
rect 16696 10560 16742 10594
rect 16776 10560 16824 10594
rect 16286 10546 16824 10560
rect 16900 10594 17438 10614
rect 16900 10560 16948 10594
rect 16982 10560 17028 10594
rect 17062 10560 17108 10594
rect 17142 10560 17188 10594
rect 17222 10560 17268 10594
rect 17302 10560 17348 10594
rect 17382 10560 17438 10594
rect 16900 10546 17438 10560
rect 17498 10594 18036 10614
rect 17498 10560 17554 10594
rect 17588 10560 17634 10594
rect 17668 10560 17714 10594
rect 17748 10560 17794 10594
rect 17828 10560 17874 10594
rect 17908 10560 17954 10594
rect 17988 10560 18036 10594
rect 17498 10546 18036 10560
rect 18268 10543 18354 10569
rect 18268 10509 18294 10543
rect 18328 10509 18354 10543
rect 18268 10483 18354 10509
rect 12522 10413 12605 10438
rect 12522 10378 12547 10413
rect 12581 10378 12605 10413
rect 12522 10354 12605 10378
rect 18273 10399 18359 10425
rect 18273 10365 18299 10399
rect 18333 10365 18359 10399
rect 18273 10339 18359 10365
rect 18274 10247 18360 10273
rect 18274 10213 18300 10247
rect 18334 10213 18360 10247
rect 18274 10187 18360 10213
rect 18274 10077 18360 10103
rect 18274 10043 18300 10077
rect 18334 10043 18360 10077
rect 11836 10025 12252 10027
rect 11836 9991 11866 10025
rect 11900 9991 11996 10025
rect 12030 9991 12142 10025
rect 12176 9991 12252 10025
rect 11836 9987 12252 9991
rect 18274 10017 18360 10043
rect 18273 9920 18359 9946
rect 18273 9886 18299 9920
rect 18333 9886 18359 9920
rect 18273 9860 18359 9886
rect 18472 9652 18841 9654
rect 18472 9618 18501 9652
rect 18535 9618 18684 9652
rect 18718 9618 18841 9652
rect 13370 6955 13400 6989
rect 13434 6955 13491 6989
rect 13525 6955 13584 6989
rect 13618 6955 13675 6989
rect 13709 6955 13766 6989
rect 13800 6955 13860 6989
rect 13894 6955 13951 6989
rect 13985 6955 14044 6989
rect 14078 6955 14135 6989
rect 14169 6955 14227 6989
rect 14261 6955 14318 6989
rect 14352 6955 14411 6989
rect 14445 6955 14504 6989
rect 14538 6955 14595 6989
rect 14629 6955 14687 6989
rect 14721 6955 14779 6989
rect 14813 6955 14871 6989
rect 14905 6955 14963 6989
rect 14997 6955 15055 6989
rect 15089 6955 15147 6989
rect 15181 6955 15240 6989
rect 15274 6955 15330 6989
rect 15364 6955 15423 6989
rect 15457 6955 15516 6989
rect 15550 6955 15608 6989
rect 15642 6955 15699 6989
rect 15733 6955 15792 6989
rect 15826 6955 15884 6989
rect 15918 6955 15976 6989
rect 16010 6955 16068 6989
rect 16102 6955 16160 6989
rect 16194 6955 16252 6989
rect 16286 6955 16343 6989
rect 16377 6955 16434 6989
rect 16468 6955 16527 6989
rect 16561 6955 16620 6989
rect 16654 6955 16712 6989
rect 16746 6955 16803 6989
rect 16837 6955 16897 6989
rect 16931 6955 16987 6989
rect 17021 6955 17078 6989
rect 17112 6955 17171 6989
rect 17205 6955 17264 6989
rect 17298 6955 17356 6989
rect 17390 6955 17447 6989
rect 17481 6955 17539 6989
rect 17573 6955 17631 6989
rect 17665 6955 17722 6989
rect 17756 6955 17814 6989
rect 17848 6955 17907 6989
rect 17941 6955 17999 6989
rect 18033 6955 18091 6989
rect 18125 6955 18154 6989
rect 13370 5674 13402 5708
rect 13436 5674 13492 5708
rect 13526 5674 13585 5708
rect 13619 5674 13675 5708
rect 13709 5674 13766 5708
rect 13800 5674 13860 5708
rect 13894 5674 13951 5708
rect 13985 5674 14043 5708
rect 14077 5674 14135 5708
rect 14169 5674 14228 5708
rect 14262 5674 14319 5708
rect 14353 5674 14411 5708
rect 14445 5674 14503 5708
rect 14537 5674 14595 5708
rect 14629 5674 14688 5708
rect 14722 5674 14779 5708
rect 14813 5674 14870 5708
rect 14904 5674 14963 5708
rect 14997 5674 15056 5708
rect 15090 5674 15147 5708
rect 15181 5674 15239 5708
rect 15273 5674 15331 5708
rect 15365 5674 15423 5708
rect 15457 5674 15516 5708
rect 15550 5674 15606 5708
rect 15640 5674 15699 5708
rect 15733 5674 15791 5708
rect 15825 5674 15884 5708
rect 15918 5674 15978 5708
rect 16012 5674 16067 5708
rect 16101 5674 16159 5708
rect 16193 5674 16251 5708
rect 16285 5674 16343 5708
rect 16377 5674 16435 5708
rect 16469 5674 16527 5708
rect 16561 5674 16619 5708
rect 16653 5674 16711 5708
rect 16745 5674 16803 5708
rect 16837 5674 16895 5708
rect 16929 5674 16987 5708
rect 17021 5674 17079 5708
rect 17113 5674 17171 5708
rect 17205 5674 17263 5708
rect 17297 5674 17355 5708
rect 17389 5674 17447 5708
rect 17481 5674 17539 5708
rect 17573 5674 17631 5708
rect 17665 5674 17723 5708
rect 17757 5674 17815 5708
rect 17849 5674 17907 5708
rect 17941 5674 18000 5708
rect 18034 5674 18091 5708
rect 18125 5674 18154 5708
<< psubdiffcont >>
rect 11886 9389 11920 9423
rect 12004 9389 12038 9423
rect 12148 9389 12182 9423
rect 18501 9006 18535 9040
rect 18593 9007 18627 9041
rect 18685 9007 18719 9041
rect 18778 9007 18812 9041
rect 12617 8164 12651 8198
rect 13010 7993 13044 8027
rect 13090 7993 13124 8027
rect 13170 7993 13204 8027
rect 13250 7993 13284 8027
rect 13742 7993 13776 8027
rect 13822 7993 13856 8027
rect 13902 7993 13936 8027
rect 13982 7993 14016 8027
rect 14350 7993 14384 8027
rect 14430 7993 14464 8027
rect 14510 7993 14544 8027
rect 14590 7993 14624 8027
rect 14954 7993 14988 8027
rect 15034 7993 15068 8027
rect 15114 7993 15148 8027
rect 15194 7993 15228 8027
rect 15562 7993 15596 8027
rect 15642 7993 15676 8027
rect 15722 7993 15756 8027
rect 15802 7993 15836 8027
rect 16292 7993 16326 8027
rect 16372 7993 16406 8027
rect 16452 7993 16486 8027
rect 16532 7993 16566 8027
rect 16900 7993 16934 8027
rect 16980 7993 17014 8027
rect 17060 7993 17094 8027
rect 17140 7993 17174 8027
rect 17634 7993 17668 8027
rect 17714 7993 17748 8027
rect 17794 7993 17828 8027
rect 17874 7993 17908 8027
rect 13399 7581 13433 7615
rect 13491 7581 13525 7615
rect 13583 7581 13617 7615
rect 13675 7581 13709 7615
rect 13767 7581 13801 7615
rect 13859 7581 13893 7615
rect 13951 7581 13985 7615
rect 14043 7581 14077 7615
rect 14135 7581 14169 7615
rect 14226 7581 14260 7615
rect 14319 7581 14353 7615
rect 14411 7581 14445 7615
rect 14503 7581 14537 7615
rect 14595 7581 14629 7615
rect 14687 7581 14721 7615
rect 14779 7581 14813 7615
rect 14871 7581 14905 7615
rect 14963 7581 14997 7615
rect 15055 7581 15089 7615
rect 15147 7581 15181 7615
rect 15239 7581 15273 7615
rect 15331 7581 15365 7615
rect 15423 7581 15457 7615
rect 15515 7581 15549 7615
rect 15607 7581 15641 7615
rect 15699 7581 15733 7615
rect 15791 7581 15825 7615
rect 15883 7581 15917 7615
rect 15975 7581 16009 7615
rect 16067 7581 16101 7615
rect 16159 7581 16193 7615
rect 16251 7581 16285 7615
rect 16343 7581 16377 7615
rect 16435 7581 16469 7615
rect 16527 7581 16561 7615
rect 16619 7581 16653 7615
rect 16711 7581 16745 7615
rect 16803 7581 16837 7615
rect 16895 7581 16929 7615
rect 16987 7581 17021 7615
rect 17079 7581 17113 7615
rect 17171 7581 17205 7615
rect 17263 7581 17297 7615
rect 17355 7581 17389 7615
rect 17447 7581 17481 7615
rect 17539 7581 17573 7615
rect 17631 7581 17665 7615
rect 17723 7581 17757 7615
rect 17815 7581 17849 7615
rect 17907 7581 17941 7615
rect 17999 7581 18033 7615
rect 18091 7581 18125 7615
rect 13399 6316 13433 6350
rect 13491 6316 13525 6350
rect 13583 6316 13617 6350
rect 13675 6316 13709 6350
rect 13767 6316 13801 6350
rect 13859 6316 13893 6350
rect 13951 6316 13985 6350
rect 14043 6316 14077 6350
rect 14135 6316 14169 6350
rect 14227 6316 14261 6350
rect 14319 6316 14353 6350
rect 14411 6316 14445 6350
rect 14503 6316 14537 6350
rect 14595 6316 14629 6350
rect 14687 6316 14721 6350
rect 14779 6316 14813 6350
rect 14871 6316 14905 6350
rect 14964 6316 14998 6350
rect 15055 6316 15089 6350
rect 15147 6316 15181 6350
rect 15239 6316 15273 6350
rect 15332 6316 15366 6350
rect 15423 6316 15457 6350
rect 15515 6316 15549 6350
rect 15607 6316 15641 6350
rect 15699 6316 15733 6350
rect 15791 6316 15825 6350
rect 15883 6316 15917 6350
rect 15975 6316 16009 6350
rect 16067 6316 16101 6350
rect 16159 6316 16193 6350
rect 16251 6316 16285 6350
rect 16343 6316 16377 6350
rect 16435 6316 16469 6350
rect 16526 6316 16560 6350
rect 16618 6316 16652 6350
rect 16711 6316 16745 6350
rect 16803 6316 16837 6350
rect 16895 6316 16929 6350
rect 16986 6316 17020 6350
rect 17079 6316 17113 6350
rect 17170 6316 17204 6350
rect 17263 6316 17297 6350
rect 17355 6316 17389 6350
rect 17447 6316 17481 6350
rect 17539 6316 17573 6350
rect 17631 6316 17665 6350
rect 17723 6316 17757 6350
rect 17815 6316 17849 6350
rect 17907 6316 17941 6350
rect 17999 6316 18033 6350
rect 18091 6316 18125 6350
rect 13399 5049 13433 5083
rect 13491 5049 13525 5083
rect 13583 5049 13617 5083
rect 13675 5049 13709 5083
rect 13767 5049 13801 5083
rect 13859 5049 13893 5083
rect 13951 5049 13985 5083
rect 14043 5049 14077 5083
rect 14135 5049 14169 5083
rect 14227 5049 14261 5083
rect 14319 5049 14353 5083
rect 14411 5049 14445 5083
rect 14503 5049 14537 5083
rect 14595 5049 14629 5083
rect 14687 5049 14721 5083
rect 14779 5049 14813 5083
rect 14871 5049 14905 5083
rect 14963 5049 14997 5083
rect 15055 5049 15089 5083
rect 15147 5049 15181 5083
rect 15239 5049 15273 5083
rect 15331 5049 15365 5083
rect 15423 5049 15457 5083
rect 15515 5049 15549 5083
rect 15607 5049 15641 5083
rect 15699 5049 15733 5083
rect 15791 5049 15825 5083
rect 15883 5049 15917 5083
rect 15975 5049 16009 5083
rect 16067 5049 16101 5083
rect 16159 5049 16193 5083
rect 16251 5049 16285 5083
rect 16343 5049 16377 5083
rect 16435 5049 16469 5083
rect 16527 5049 16561 5083
rect 16619 5049 16653 5083
rect 16711 5049 16745 5083
rect 16803 5049 16837 5083
rect 16895 5049 16929 5083
rect 16987 5049 17021 5083
rect 17079 5049 17113 5083
rect 17171 5049 17205 5083
rect 17263 5049 17297 5083
rect 17355 5049 17389 5083
rect 17447 5049 17481 5083
rect 17539 5049 17573 5083
rect 17631 5049 17665 5083
rect 17723 5049 17757 5083
rect 17815 5049 17849 5083
rect 17907 5049 17941 5083
rect 17999 5049 18033 5083
rect 18091 5049 18125 5083
<< nsubdiffcont >>
rect 12580 10557 12614 10591
rect 12660 10557 12694 10591
rect 12740 10557 12774 10591
rect 12820 10557 12854 10591
rect 12900 10557 12934 10591
rect 12980 10557 13014 10591
rect 13312 10560 13346 10594
rect 13392 10560 13426 10594
rect 13472 10560 13506 10594
rect 13552 10560 13586 10594
rect 13632 10560 13666 10594
rect 13712 10560 13746 10594
rect 13918 10560 13952 10594
rect 13998 10560 14032 10594
rect 14078 10560 14112 10594
rect 14158 10560 14192 10594
rect 14238 10560 14272 10594
rect 14318 10560 14352 10594
rect 14524 10560 14558 10594
rect 14604 10560 14638 10594
rect 14684 10560 14718 10594
rect 14764 10560 14798 10594
rect 14844 10560 14878 10594
rect 14924 10560 14958 10594
rect 15130 10560 15164 10594
rect 15210 10560 15244 10594
rect 15290 10560 15324 10594
rect 15370 10560 15404 10594
rect 15450 10560 15484 10594
rect 15530 10560 15564 10594
rect 15736 10560 15770 10594
rect 15816 10560 15850 10594
rect 15896 10560 15930 10594
rect 15976 10560 16010 10594
rect 16056 10560 16090 10594
rect 16136 10560 16170 10594
rect 16342 10560 16376 10594
rect 16422 10560 16456 10594
rect 16502 10560 16536 10594
rect 16582 10560 16616 10594
rect 16662 10560 16696 10594
rect 16742 10560 16776 10594
rect 16948 10560 16982 10594
rect 17028 10560 17062 10594
rect 17108 10560 17142 10594
rect 17188 10560 17222 10594
rect 17268 10560 17302 10594
rect 17348 10560 17382 10594
rect 17554 10560 17588 10594
rect 17634 10560 17668 10594
rect 17714 10560 17748 10594
rect 17794 10560 17828 10594
rect 17874 10560 17908 10594
rect 17954 10560 17988 10594
rect 18294 10509 18328 10543
rect 12547 10378 12581 10413
rect 18299 10365 18333 10399
rect 18300 10213 18334 10247
rect 18300 10043 18334 10077
rect 11866 9991 11900 10025
rect 11996 9991 12030 10025
rect 12142 9991 12176 10025
rect 18299 9886 18333 9920
rect 18501 9618 18535 9652
rect 18684 9618 18718 9652
rect 13400 6955 13434 6989
rect 13491 6955 13525 6989
rect 13584 6955 13618 6989
rect 13675 6955 13709 6989
rect 13766 6955 13800 6989
rect 13860 6955 13894 6989
rect 13951 6955 13985 6989
rect 14044 6955 14078 6989
rect 14135 6955 14169 6989
rect 14227 6955 14261 6989
rect 14318 6955 14352 6989
rect 14411 6955 14445 6989
rect 14504 6955 14538 6989
rect 14595 6955 14629 6989
rect 14687 6955 14721 6989
rect 14779 6955 14813 6989
rect 14871 6955 14905 6989
rect 14963 6955 14997 6989
rect 15055 6955 15089 6989
rect 15147 6955 15181 6989
rect 15240 6955 15274 6989
rect 15330 6955 15364 6989
rect 15423 6955 15457 6989
rect 15516 6955 15550 6989
rect 15608 6955 15642 6989
rect 15699 6955 15733 6989
rect 15792 6955 15826 6989
rect 15884 6955 15918 6989
rect 15976 6955 16010 6989
rect 16068 6955 16102 6989
rect 16160 6955 16194 6989
rect 16252 6955 16286 6989
rect 16343 6955 16377 6989
rect 16434 6955 16468 6989
rect 16527 6955 16561 6989
rect 16620 6955 16654 6989
rect 16712 6955 16746 6989
rect 16803 6955 16837 6989
rect 16897 6955 16931 6989
rect 16987 6955 17021 6989
rect 17078 6955 17112 6989
rect 17171 6955 17205 6989
rect 17264 6955 17298 6989
rect 17356 6955 17390 6989
rect 17447 6955 17481 6989
rect 17539 6955 17573 6989
rect 17631 6955 17665 6989
rect 17722 6955 17756 6989
rect 17814 6955 17848 6989
rect 17907 6955 17941 6989
rect 17999 6955 18033 6989
rect 18091 6955 18125 6989
rect 13402 5674 13436 5708
rect 13492 5674 13526 5708
rect 13585 5674 13619 5708
rect 13675 5674 13709 5708
rect 13766 5674 13800 5708
rect 13860 5674 13894 5708
rect 13951 5674 13985 5708
rect 14043 5674 14077 5708
rect 14135 5674 14169 5708
rect 14228 5674 14262 5708
rect 14319 5674 14353 5708
rect 14411 5674 14445 5708
rect 14503 5674 14537 5708
rect 14595 5674 14629 5708
rect 14688 5674 14722 5708
rect 14779 5674 14813 5708
rect 14870 5674 14904 5708
rect 14963 5674 14997 5708
rect 15056 5674 15090 5708
rect 15147 5674 15181 5708
rect 15239 5674 15273 5708
rect 15331 5674 15365 5708
rect 15423 5674 15457 5708
rect 15516 5674 15550 5708
rect 15606 5674 15640 5708
rect 15699 5674 15733 5708
rect 15791 5674 15825 5708
rect 15884 5674 15918 5708
rect 15978 5674 16012 5708
rect 16067 5674 16101 5708
rect 16159 5674 16193 5708
rect 16251 5674 16285 5708
rect 16343 5674 16377 5708
rect 16435 5674 16469 5708
rect 16527 5674 16561 5708
rect 16619 5674 16653 5708
rect 16711 5674 16745 5708
rect 16803 5674 16837 5708
rect 16895 5674 16929 5708
rect 16987 5674 17021 5708
rect 17079 5674 17113 5708
rect 17171 5674 17205 5708
rect 17263 5674 17297 5708
rect 17355 5674 17389 5708
rect 17447 5674 17481 5708
rect 17539 5674 17573 5708
rect 17631 5674 17665 5708
rect 17723 5674 17757 5708
rect 17815 5674 17849 5708
rect 17907 5674 17941 5708
rect 18000 5674 18034 5708
rect 18091 5674 18125 5708
<< poly >>
rect 12380 10579 12410 10609
rect 12380 10441 12410 10495
rect 12380 10303 12410 10357
rect 12380 10165 12410 10219
rect 12380 10027 12410 10081
rect 11912 9932 11942 9958
rect 12102 9932 12132 9958
rect 12380 9889 12410 9943
rect 12380 9774 12410 9805
rect 12362 9758 12428 9774
rect 11912 9700 11942 9732
rect 11856 9684 11942 9700
rect 11856 9650 11872 9684
rect 11906 9650 11942 9684
rect 11856 9634 11942 9650
rect 11912 9612 11942 9634
rect 12102 9700 12132 9732
rect 12362 9724 12378 9758
rect 12412 9724 12428 9758
rect 12362 9708 12428 9724
rect 12102 9684 12188 9700
rect 12102 9650 12138 9684
rect 12172 9650 12188 9684
rect 12102 9634 12188 9650
rect 12102 9612 12132 9634
rect 18165 9578 18195 9609
rect 13004 9515 13070 9531
rect 11912 9456 11942 9482
rect 12102 9456 12132 9482
rect 13004 9481 13020 9515
rect 13054 9481 13070 9515
rect 13004 9465 13070 9481
rect 13736 9518 13802 9534
rect 13736 9484 13752 9518
rect 13786 9484 13802 9518
rect 13736 9468 13802 9484
rect 13862 9518 13928 9534
rect 13862 9484 13878 9518
rect 13912 9484 13928 9518
rect 13862 9468 13928 9484
rect 14948 9518 15014 9534
rect 14948 9484 14964 9518
rect 14998 9484 15014 9518
rect 14948 9468 15014 9484
rect 15074 9518 15140 9534
rect 15074 9484 15090 9518
rect 15124 9484 15140 9518
rect 15074 9468 15140 9484
rect 16160 9518 16226 9534
rect 16160 9484 16176 9518
rect 16210 9484 16226 9518
rect 16160 9468 16226 9484
rect 16286 9518 16352 9534
rect 16286 9484 16302 9518
rect 16336 9484 16352 9518
rect 16286 9468 16352 9484
rect 17372 9518 17438 9534
rect 17372 9484 17388 9518
rect 17422 9484 17438 9518
rect 17372 9468 17438 9484
rect 17498 9518 17564 9534
rect 17498 9484 17514 9518
rect 17548 9484 17564 9518
rect 18551 9547 18581 9573
rect 18646 9555 18676 9581
rect 18730 9555 18760 9581
rect 17498 9468 17564 9484
rect 13022 9434 13052 9465
rect 13754 9437 13784 9468
rect 13880 9437 13910 9468
rect 14966 9437 14996 9468
rect 15092 9437 15122 9468
rect 16178 9437 16208 9468
rect 16304 9437 16334 9468
rect 17390 9437 17420 9468
rect 17516 9437 17546 9468
rect 18165 9440 18195 9494
rect 18257 9440 18287 9466
rect 18353 9440 18383 9471
rect 13022 9322 13052 9350
rect 13754 9325 13784 9353
rect 13880 9325 13910 9353
rect 14966 9325 14996 9353
rect 15092 9325 15122 9353
rect 16178 9325 16208 9353
rect 16304 9325 16334 9353
rect 17390 9325 17420 9353
rect 17516 9325 17546 9353
rect 18165 9331 18195 9356
rect 18036 9311 18195 9331
rect 18257 9331 18287 9356
rect 18353 9331 18383 9356
rect 18257 9325 18383 9331
rect 18036 9277 18048 9311
rect 18082 9277 18195 9311
rect 13375 9236 13405 9262
rect 14107 9236 14137 9262
rect 14229 9236 14259 9262
rect 15319 9236 15349 9262
rect 15441 9236 15471 9262
rect 16657 9236 16687 9262
rect 16779 9236 16809 9262
rect 17513 9236 17543 9262
rect 18036 9258 18195 9277
rect 18239 9309 18383 9325
rect 18551 9323 18581 9419
rect 18646 9323 18676 9355
rect 18730 9323 18760 9355
rect 18239 9275 18255 9309
rect 18289 9275 18383 9309
rect 18239 9259 18383 9275
rect 18165 9237 18195 9258
rect 18257 9252 18383 9259
rect 18499 9307 18581 9323
rect 18499 9273 18509 9307
rect 18543 9273 18581 9307
rect 18499 9257 18581 9273
rect 18623 9307 18760 9323
rect 18623 9273 18633 9307
rect 18667 9273 18760 9307
rect 18623 9257 18760 9273
rect 18257 9237 18287 9252
rect 18353 9237 18383 9252
rect 18551 9189 18581 9257
rect 18646 9235 18676 9257
rect 18730 9235 18760 9257
rect 12373 9124 12439 9140
rect 13375 9130 13405 9152
rect 14107 9130 14137 9152
rect 14229 9130 14259 9152
rect 15319 9130 15349 9152
rect 15441 9130 15471 9152
rect 16657 9130 16687 9152
rect 16779 9130 16809 9152
rect 17513 9130 17543 9152
rect 12373 9097 12389 9124
rect 12355 9090 12389 9097
rect 12423 9097 12439 9124
rect 13357 9114 13423 9130
rect 12423 9090 12457 9097
rect 12355 9067 12457 9090
rect 12355 9052 12385 9067
rect 12427 9052 12457 9067
rect 13357 9080 13373 9114
rect 13407 9080 13423 9114
rect 13357 9064 13423 9080
rect 14089 9114 14155 9130
rect 14089 9080 14105 9114
rect 14139 9080 14155 9114
rect 14089 9064 14155 9080
rect 14211 9114 14277 9130
rect 14211 9080 14227 9114
rect 14261 9080 14277 9114
rect 14211 9064 14277 9080
rect 15301 9114 15367 9130
rect 15301 9080 15317 9114
rect 15351 9080 15367 9114
rect 15301 9064 15367 9080
rect 15423 9114 15489 9130
rect 15423 9080 15439 9114
rect 15473 9080 15489 9114
rect 15423 9064 15489 9080
rect 16639 9114 16705 9130
rect 16639 9080 16655 9114
rect 16689 9080 16705 9114
rect 16639 9064 16705 9080
rect 16761 9114 16827 9130
rect 16761 9080 16777 9114
rect 16811 9080 16827 9114
rect 16761 9064 16827 9080
rect 17495 9114 17561 9130
rect 17495 9080 17511 9114
rect 17545 9080 17561 9114
rect 18165 9099 18195 9153
rect 18257 9127 18287 9153
rect 18353 9127 18383 9153
rect 17495 9064 17561 9080
rect 18551 9079 18581 9105
rect 18646 9079 18676 9105
rect 18730 9079 18760 9105
rect 18165 8988 18195 9015
rect 12355 8914 12385 8968
rect 12427 8914 12457 8968
rect 12355 8776 12385 8830
rect 12427 8776 12457 8830
rect 12355 8638 12385 8692
rect 12427 8638 12457 8692
rect 12355 8500 12385 8554
rect 12427 8500 12457 8554
rect 12355 8362 12385 8416
rect 12427 8362 12457 8416
rect 12355 8224 12385 8278
rect 12427 8224 12457 8278
rect 12355 8086 12385 8140
rect 12427 8086 12457 8140
rect 12355 7976 12385 8002
rect 12427 7976 12457 8002
rect 13449 7517 13479 7543
rect 13533 7517 13563 7543
rect 13721 7517 13751 7543
rect 13816 7517 13846 7543
rect 13922 7517 13952 7543
rect 14018 7517 14048 7543
rect 14128 7517 14158 7543
rect 14228 7517 14258 7543
rect 14312 7517 14342 7543
rect 14500 7517 14530 7543
rect 14595 7517 14625 7543
rect 14704 7517 14734 7543
rect 14799 7517 14829 7543
rect 14885 7517 14915 7543
rect 15003 7517 15033 7543
rect 15087 7517 15117 7543
rect 15275 7517 15305 7543
rect 15370 7517 15400 7543
rect 15558 7517 15588 7543
rect 15653 7517 15683 7543
rect 15841 7517 15871 7543
rect 15925 7517 15955 7543
rect 16113 7517 16143 7543
rect 16208 7517 16238 7543
rect 16314 7517 16344 7543
rect 16410 7517 16440 7543
rect 16520 7517 16550 7543
rect 16620 7517 16650 7543
rect 16704 7517 16734 7543
rect 16892 7517 16922 7543
rect 16987 7517 17017 7543
rect 17096 7517 17126 7543
rect 17191 7517 17221 7543
rect 17277 7517 17307 7543
rect 17395 7517 17425 7543
rect 17479 7517 17509 7543
rect 17667 7517 17697 7543
rect 17762 7517 17792 7543
rect 17950 7517 17980 7543
rect 18045 7517 18075 7543
rect 13449 7418 13479 7433
rect 13416 7388 13479 7418
rect 13416 7350 13446 7388
rect 13391 7334 13446 7350
rect 13533 7344 13563 7433
rect 13721 7363 13751 7433
rect 13816 7423 13846 7445
rect 13816 7407 13880 7423
rect 13816 7373 13836 7407
rect 13870 7373 13880 7407
rect 13391 7300 13402 7334
rect 13436 7300 13446 7334
rect 13391 7284 13446 7300
rect 13488 7334 13563 7344
rect 13488 7300 13504 7334
rect 13538 7300 13563 7334
rect 13488 7290 13563 7300
rect 13710 7347 13764 7363
rect 13816 7357 13880 7373
rect 13922 7411 13952 7445
rect 13922 7395 13976 7411
rect 13922 7361 13932 7395
rect 13966 7361 13976 7395
rect 13710 7313 13720 7347
rect 13754 7313 13764 7347
rect 13922 7345 13976 7361
rect 13922 7315 13952 7345
rect 13710 7297 13764 7313
rect 13416 7246 13446 7284
rect 13416 7216 13479 7246
rect 13449 7201 13479 7216
rect 13533 7201 13563 7290
rect 13721 7151 13751 7297
rect 13814 7285 13952 7315
rect 13814 7151 13844 7285
rect 14018 7249 14048 7433
rect 14128 7401 14158 7433
rect 14094 7385 14158 7401
rect 14595 7423 14625 7445
rect 14595 7407 14662 7423
rect 14094 7351 14104 7385
rect 14138 7371 14158 7385
rect 14138 7351 14154 7371
rect 14094 7335 14154 7351
rect 13886 7233 13952 7243
rect 13886 7199 13902 7233
rect 13936 7199 13952 7233
rect 13886 7189 13952 7199
rect 14018 7233 14082 7249
rect 14018 7199 14038 7233
rect 14072 7199 14082 7233
rect 13898 7151 13928 7189
rect 14018 7183 14082 7199
rect 14018 7151 14048 7183
rect 14124 7151 14154 7335
rect 14228 7333 14258 7389
rect 14312 7333 14342 7389
rect 14500 7367 14530 7389
rect 14476 7351 14530 7367
rect 14595 7373 14618 7407
rect 14652 7373 14662 7407
rect 14595 7357 14662 7373
rect 14196 7317 14262 7333
rect 14196 7283 14206 7317
rect 14240 7283 14262 7317
rect 14196 7267 14262 7283
rect 14312 7317 14402 7333
rect 14476 7331 14486 7351
rect 14312 7283 14358 7317
rect 14392 7283 14402 7317
rect 14312 7267 14402 7283
rect 14453 7317 14486 7331
rect 14520 7317 14530 7351
rect 14453 7301 14530 7317
rect 14704 7315 14734 7445
rect 14232 7235 14262 7267
rect 14316 7235 14346 7267
rect 14453 7235 14483 7301
rect 14597 7285 14734 7315
rect 14597 7249 14627 7285
rect 13449 7047 13479 7073
rect 13533 7047 13563 7073
rect 14573 7233 14627 7249
rect 14799 7249 14829 7433
rect 14885 7401 14915 7433
rect 14871 7385 14937 7401
rect 14871 7351 14881 7385
rect 14915 7351 14937 7385
rect 14871 7335 14937 7351
rect 15003 7349 15033 7389
rect 14573 7199 14583 7233
rect 14617 7199 14627 7233
rect 14573 7183 14627 7199
rect 14669 7233 14735 7243
rect 14669 7199 14685 7233
rect 14719 7199 14735 7233
rect 14669 7189 14735 7199
rect 14799 7233 14865 7249
rect 14799 7199 14821 7233
rect 14855 7199 14865 7233
rect 14597 7151 14627 7183
rect 14681 7151 14711 7189
rect 14799 7183 14865 7199
rect 14799 7151 14829 7183
rect 14907 7151 14937 7335
rect 14979 7333 15033 7349
rect 14979 7299 14989 7333
rect 15023 7299 15033 7333
rect 14979 7283 15033 7299
rect 15087 7333 15117 7389
rect 15275 7361 15305 7433
rect 15558 7418 15588 7433
rect 15532 7388 15588 7418
rect 15370 7365 15400 7387
rect 15242 7345 15306 7361
rect 15087 7317 15171 7333
rect 15087 7297 15127 7317
rect 15003 7235 15033 7283
rect 15075 7283 15127 7297
rect 15161 7283 15171 7317
rect 15242 7311 15258 7345
rect 15292 7311 15306 7345
rect 15242 7295 15306 7311
rect 15348 7359 15400 7365
rect 15532 7359 15562 7388
rect 15841 7418 15871 7433
rect 15808 7388 15871 7418
rect 15653 7365 15683 7387
rect 15348 7349 15562 7359
rect 15348 7315 15358 7349
rect 15392 7315 15562 7349
rect 15348 7305 15562 7315
rect 15348 7299 15400 7305
rect 15075 7267 15171 7283
rect 15075 7235 15105 7267
rect 15273 7263 15303 7295
rect 15370 7267 15400 7299
rect 15273 7109 15303 7135
rect 15532 7257 15562 7305
rect 15624 7349 15683 7365
rect 15808 7350 15838 7388
rect 15624 7315 15634 7349
rect 15668 7315 15683 7349
rect 15624 7299 15683 7315
rect 15653 7267 15683 7299
rect 15783 7334 15838 7350
rect 15925 7344 15955 7433
rect 16113 7363 16143 7433
rect 16208 7423 16238 7445
rect 16208 7407 16272 7423
rect 16208 7373 16228 7407
rect 16262 7373 16272 7407
rect 15783 7300 15794 7334
rect 15828 7300 15838 7334
rect 15783 7284 15838 7300
rect 15880 7334 15955 7344
rect 15880 7300 15896 7334
rect 15930 7300 15955 7334
rect 15880 7290 15955 7300
rect 16102 7347 16156 7363
rect 16208 7357 16272 7373
rect 16314 7411 16344 7445
rect 16314 7395 16368 7411
rect 16314 7361 16324 7395
rect 16358 7361 16368 7395
rect 16102 7313 16112 7347
rect 16146 7313 16156 7347
rect 16314 7345 16368 7361
rect 16314 7315 16344 7345
rect 16102 7297 16156 7313
rect 15532 7227 15588 7257
rect 15558 7211 15588 7227
rect 13721 7041 13751 7067
rect 13814 7041 13844 7067
rect 13898 7041 13928 7067
rect 14018 7041 14048 7067
rect 14124 7041 14154 7067
rect 14232 7041 14262 7067
rect 14316 7041 14346 7067
rect 14453 7041 14483 7067
rect 14597 7041 14627 7067
rect 14681 7041 14711 7067
rect 14799 7041 14829 7067
rect 14907 7041 14937 7067
rect 15003 7041 15033 7067
rect 15075 7041 15105 7067
rect 15370 7041 15400 7067
rect 15558 7057 15588 7083
rect 15808 7246 15838 7284
rect 15808 7216 15871 7246
rect 15841 7201 15871 7216
rect 15925 7201 15955 7290
rect 16113 7151 16143 7297
rect 16206 7285 16344 7315
rect 16206 7151 16236 7285
rect 16410 7249 16440 7433
rect 16520 7401 16550 7433
rect 16486 7385 16550 7401
rect 16987 7423 17017 7445
rect 16987 7407 17054 7423
rect 16486 7351 16496 7385
rect 16530 7371 16550 7385
rect 16530 7351 16546 7371
rect 16486 7335 16546 7351
rect 16278 7233 16344 7243
rect 16278 7199 16294 7233
rect 16328 7199 16344 7233
rect 16278 7189 16344 7199
rect 16410 7233 16474 7249
rect 16410 7199 16430 7233
rect 16464 7199 16474 7233
rect 16290 7151 16320 7189
rect 16410 7183 16474 7199
rect 16410 7151 16440 7183
rect 16516 7151 16546 7335
rect 16620 7333 16650 7389
rect 16704 7333 16734 7389
rect 16892 7367 16922 7389
rect 16868 7351 16922 7367
rect 16987 7373 17010 7407
rect 17044 7373 17054 7407
rect 16987 7357 17054 7373
rect 16588 7317 16654 7333
rect 16588 7283 16598 7317
rect 16632 7283 16654 7317
rect 16588 7267 16654 7283
rect 16704 7317 16794 7333
rect 16868 7331 16878 7351
rect 16704 7283 16750 7317
rect 16784 7283 16794 7317
rect 16704 7267 16794 7283
rect 16845 7317 16878 7331
rect 16912 7317 16922 7351
rect 16845 7301 16922 7317
rect 17096 7315 17126 7445
rect 16624 7235 16654 7267
rect 16708 7235 16738 7267
rect 16845 7235 16875 7301
rect 16989 7285 17126 7315
rect 16989 7249 17019 7285
rect 15653 7041 15683 7067
rect 15841 7047 15871 7073
rect 15925 7047 15955 7073
rect 16965 7233 17019 7249
rect 17191 7249 17221 7433
rect 17277 7401 17307 7433
rect 17263 7385 17329 7401
rect 17263 7351 17273 7385
rect 17307 7351 17329 7385
rect 17263 7335 17329 7351
rect 17395 7349 17425 7389
rect 16965 7199 16975 7233
rect 17009 7199 17019 7233
rect 16965 7183 17019 7199
rect 17061 7233 17127 7243
rect 17061 7199 17077 7233
rect 17111 7199 17127 7233
rect 17061 7189 17127 7199
rect 17191 7233 17257 7249
rect 17191 7199 17213 7233
rect 17247 7199 17257 7233
rect 16989 7151 17019 7183
rect 17073 7151 17103 7189
rect 17191 7183 17257 7199
rect 17191 7151 17221 7183
rect 17299 7151 17329 7335
rect 17371 7333 17425 7349
rect 17371 7299 17381 7333
rect 17415 7299 17425 7333
rect 17371 7283 17425 7299
rect 17479 7333 17509 7389
rect 17667 7361 17697 7433
rect 17950 7418 17980 7433
rect 17924 7388 17980 7418
rect 17762 7365 17792 7387
rect 17634 7345 17698 7361
rect 17479 7317 17563 7333
rect 17479 7297 17519 7317
rect 17395 7235 17425 7283
rect 17467 7283 17519 7297
rect 17553 7283 17563 7317
rect 17634 7311 17650 7345
rect 17684 7311 17698 7345
rect 17634 7295 17698 7311
rect 17740 7359 17792 7365
rect 17924 7359 17954 7388
rect 18045 7365 18075 7387
rect 17740 7349 17954 7359
rect 17740 7315 17750 7349
rect 17784 7315 17954 7349
rect 17740 7305 17954 7315
rect 17740 7299 17792 7305
rect 17467 7267 17563 7283
rect 17467 7235 17497 7267
rect 17665 7263 17695 7295
rect 17762 7267 17792 7299
rect 17665 7109 17695 7135
rect 17924 7257 17954 7305
rect 18016 7349 18075 7365
rect 18016 7315 18026 7349
rect 18060 7315 18075 7349
rect 18016 7299 18075 7315
rect 18045 7267 18075 7299
rect 17924 7227 17980 7257
rect 17950 7211 17980 7227
rect 16113 7041 16143 7067
rect 16206 7041 16236 7067
rect 16290 7041 16320 7067
rect 16410 7041 16440 7067
rect 16516 7041 16546 7067
rect 16624 7041 16654 7067
rect 16708 7041 16738 7067
rect 16845 7041 16875 7067
rect 16989 7041 17019 7067
rect 17073 7041 17103 7067
rect 17191 7041 17221 7067
rect 17299 7041 17329 7067
rect 17395 7041 17425 7067
rect 17467 7041 17497 7067
rect 17762 7041 17792 7067
rect 17950 7057 17980 7083
rect 18045 7041 18075 7067
rect 13449 6871 13479 6897
rect 13533 6871 13563 6897
rect 13721 6877 13751 6903
rect 13814 6877 13844 6903
rect 13898 6877 13928 6903
rect 14018 6877 14048 6903
rect 14124 6877 14154 6903
rect 14232 6877 14262 6903
rect 14316 6877 14346 6903
rect 14453 6877 14483 6903
rect 14597 6877 14627 6903
rect 14681 6877 14711 6903
rect 14799 6877 14829 6903
rect 14907 6877 14937 6903
rect 15003 6877 15033 6903
rect 15075 6877 15105 6903
rect 15370 6877 15400 6903
rect 13449 6728 13479 6743
rect 13416 6698 13479 6728
rect 13416 6660 13446 6698
rect 13391 6644 13446 6660
rect 13533 6654 13563 6743
rect 13391 6610 13402 6644
rect 13436 6610 13446 6644
rect 13391 6594 13446 6610
rect 13488 6644 13563 6654
rect 13721 6647 13751 6793
rect 13814 6659 13844 6793
rect 13898 6755 13928 6793
rect 14018 6761 14048 6793
rect 13886 6745 13952 6755
rect 13886 6711 13902 6745
rect 13936 6711 13952 6745
rect 13886 6701 13952 6711
rect 14018 6745 14082 6761
rect 14018 6711 14038 6745
rect 14072 6711 14082 6745
rect 14018 6695 14082 6711
rect 13488 6610 13504 6644
rect 13538 6610 13563 6644
rect 13488 6600 13563 6610
rect 13416 6556 13446 6594
rect 13416 6526 13479 6556
rect 13449 6511 13479 6526
rect 13533 6511 13563 6600
rect 13710 6631 13764 6647
rect 13710 6597 13720 6631
rect 13754 6597 13764 6631
rect 13814 6629 13952 6659
rect 13710 6581 13764 6597
rect 13922 6599 13952 6629
rect 13721 6511 13751 6581
rect 13816 6571 13880 6587
rect 13816 6537 13836 6571
rect 13870 6537 13880 6571
rect 13816 6521 13880 6537
rect 13922 6583 13976 6599
rect 13922 6549 13932 6583
rect 13966 6549 13976 6583
rect 13922 6533 13976 6549
rect 13816 6499 13846 6521
rect 13922 6499 13952 6533
rect 14018 6511 14048 6695
rect 14124 6609 14154 6793
rect 14597 6761 14627 6793
rect 14573 6745 14627 6761
rect 14681 6755 14711 6793
rect 14799 6761 14829 6793
rect 14573 6711 14583 6745
rect 14617 6711 14627 6745
rect 14232 6677 14262 6709
rect 14316 6677 14346 6709
rect 14196 6661 14262 6677
rect 14196 6627 14206 6661
rect 14240 6627 14262 6661
rect 14196 6611 14262 6627
rect 14312 6661 14402 6677
rect 14312 6627 14358 6661
rect 14392 6627 14402 6661
rect 14312 6611 14402 6627
rect 14453 6643 14483 6709
rect 14573 6695 14627 6711
rect 14669 6745 14735 6755
rect 14669 6711 14685 6745
rect 14719 6711 14735 6745
rect 14669 6701 14735 6711
rect 14799 6745 14865 6761
rect 14799 6711 14821 6745
rect 14855 6711 14865 6745
rect 14597 6659 14627 6695
rect 14799 6695 14865 6711
rect 14453 6627 14530 6643
rect 14597 6629 14734 6659
rect 14453 6613 14486 6627
rect 14094 6593 14154 6609
rect 14094 6559 14104 6593
rect 14138 6573 14154 6593
rect 14138 6559 14158 6573
rect 14094 6543 14158 6559
rect 14228 6555 14258 6611
rect 14312 6555 14342 6611
rect 14476 6593 14486 6613
rect 14520 6593 14530 6627
rect 14476 6577 14530 6593
rect 14500 6555 14530 6577
rect 14595 6571 14662 6587
rect 14128 6511 14158 6543
rect 14595 6537 14618 6571
rect 14652 6537 14662 6571
rect 14595 6521 14662 6537
rect 14595 6499 14625 6521
rect 14704 6499 14734 6629
rect 14799 6511 14829 6695
rect 14907 6609 14937 6793
rect 15273 6809 15303 6835
rect 15003 6661 15033 6709
rect 14871 6593 14937 6609
rect 14979 6645 15033 6661
rect 15075 6677 15105 6709
rect 15075 6661 15171 6677
rect 15075 6647 15127 6661
rect 14979 6611 14989 6645
rect 15023 6611 15033 6645
rect 14979 6595 15033 6611
rect 14871 6559 14881 6593
rect 14915 6559 14937 6593
rect 14871 6543 14937 6559
rect 15003 6555 15033 6595
rect 15087 6627 15127 6647
rect 15161 6627 15171 6661
rect 15273 6649 15303 6681
rect 15558 6861 15588 6887
rect 15653 6877 15683 6903
rect 15558 6717 15588 6733
rect 15532 6687 15588 6717
rect 15087 6611 15171 6627
rect 15242 6633 15306 6649
rect 15370 6645 15400 6677
rect 15087 6555 15117 6611
rect 15242 6599 15258 6633
rect 15292 6599 15306 6633
rect 15242 6583 15306 6599
rect 15348 6639 15400 6645
rect 15532 6639 15562 6687
rect 15841 6871 15871 6897
rect 15925 6871 15955 6897
rect 16113 6877 16143 6903
rect 16206 6877 16236 6903
rect 16290 6877 16320 6903
rect 16410 6877 16440 6903
rect 16516 6877 16546 6903
rect 16624 6877 16654 6903
rect 16708 6877 16738 6903
rect 16845 6877 16875 6903
rect 16989 6877 17019 6903
rect 17073 6877 17103 6903
rect 17191 6877 17221 6903
rect 17299 6877 17329 6903
rect 17395 6877 17425 6903
rect 17467 6877 17497 6903
rect 17762 6877 17792 6903
rect 15841 6728 15871 6743
rect 15808 6698 15871 6728
rect 15653 6645 15683 6677
rect 15808 6660 15838 6698
rect 15348 6629 15562 6639
rect 15348 6595 15358 6629
rect 15392 6595 15562 6629
rect 15348 6585 15562 6595
rect 14885 6511 14915 6543
rect 15275 6511 15305 6583
rect 15348 6579 15400 6585
rect 15370 6557 15400 6579
rect 15532 6556 15562 6585
rect 15624 6629 15683 6645
rect 15624 6595 15634 6629
rect 15668 6595 15683 6629
rect 15624 6579 15683 6595
rect 15783 6644 15838 6660
rect 15925 6654 15955 6743
rect 15783 6610 15794 6644
rect 15828 6610 15838 6644
rect 15783 6594 15838 6610
rect 15880 6644 15955 6654
rect 16113 6647 16143 6793
rect 16206 6659 16236 6793
rect 16290 6755 16320 6793
rect 16410 6761 16440 6793
rect 16278 6745 16344 6755
rect 16278 6711 16294 6745
rect 16328 6711 16344 6745
rect 16278 6701 16344 6711
rect 16410 6745 16474 6761
rect 16410 6711 16430 6745
rect 16464 6711 16474 6745
rect 16410 6695 16474 6711
rect 15880 6610 15896 6644
rect 15930 6610 15955 6644
rect 15880 6600 15955 6610
rect 15653 6557 15683 6579
rect 15532 6526 15588 6556
rect 15558 6511 15588 6526
rect 15808 6556 15838 6594
rect 15808 6526 15871 6556
rect 15841 6511 15871 6526
rect 15925 6511 15955 6600
rect 16102 6631 16156 6647
rect 16102 6597 16112 6631
rect 16146 6597 16156 6631
rect 16206 6629 16344 6659
rect 16102 6581 16156 6597
rect 16314 6599 16344 6629
rect 16113 6511 16143 6581
rect 16208 6571 16272 6587
rect 16208 6537 16228 6571
rect 16262 6537 16272 6571
rect 16208 6521 16272 6537
rect 16314 6583 16368 6599
rect 16314 6549 16324 6583
rect 16358 6549 16368 6583
rect 16314 6533 16368 6549
rect 16208 6499 16238 6521
rect 16314 6499 16344 6533
rect 16410 6511 16440 6695
rect 16516 6609 16546 6793
rect 16989 6761 17019 6793
rect 16965 6745 17019 6761
rect 17073 6755 17103 6793
rect 17191 6761 17221 6793
rect 16965 6711 16975 6745
rect 17009 6711 17019 6745
rect 16624 6677 16654 6709
rect 16708 6677 16738 6709
rect 16588 6661 16654 6677
rect 16588 6627 16598 6661
rect 16632 6627 16654 6661
rect 16588 6611 16654 6627
rect 16704 6661 16794 6677
rect 16704 6627 16750 6661
rect 16784 6627 16794 6661
rect 16704 6611 16794 6627
rect 16845 6643 16875 6709
rect 16965 6695 17019 6711
rect 17061 6745 17127 6755
rect 17061 6711 17077 6745
rect 17111 6711 17127 6745
rect 17061 6701 17127 6711
rect 17191 6745 17257 6761
rect 17191 6711 17213 6745
rect 17247 6711 17257 6745
rect 16989 6659 17019 6695
rect 17191 6695 17257 6711
rect 16845 6627 16922 6643
rect 16989 6629 17126 6659
rect 16845 6613 16878 6627
rect 16486 6593 16546 6609
rect 16486 6559 16496 6593
rect 16530 6573 16546 6593
rect 16530 6559 16550 6573
rect 16486 6543 16550 6559
rect 16620 6555 16650 6611
rect 16704 6555 16734 6611
rect 16868 6593 16878 6613
rect 16912 6593 16922 6627
rect 16868 6577 16922 6593
rect 16892 6555 16922 6577
rect 16987 6571 17054 6587
rect 16520 6511 16550 6543
rect 16987 6537 17010 6571
rect 17044 6537 17054 6571
rect 16987 6521 17054 6537
rect 16987 6499 17017 6521
rect 17096 6499 17126 6629
rect 17191 6511 17221 6695
rect 17299 6609 17329 6793
rect 17665 6809 17695 6835
rect 17395 6661 17425 6709
rect 17263 6593 17329 6609
rect 17371 6645 17425 6661
rect 17467 6677 17497 6709
rect 17467 6661 17563 6677
rect 17467 6647 17519 6661
rect 17371 6611 17381 6645
rect 17415 6611 17425 6645
rect 17371 6595 17425 6611
rect 17263 6559 17273 6593
rect 17307 6559 17329 6593
rect 17263 6543 17329 6559
rect 17395 6555 17425 6595
rect 17479 6627 17519 6647
rect 17553 6627 17563 6661
rect 17665 6649 17695 6681
rect 17950 6861 17980 6887
rect 18045 6877 18075 6903
rect 17950 6717 17980 6733
rect 17924 6687 17980 6717
rect 17479 6611 17563 6627
rect 17634 6633 17698 6649
rect 17762 6645 17792 6677
rect 17479 6555 17509 6611
rect 17634 6599 17650 6633
rect 17684 6599 17698 6633
rect 17634 6583 17698 6599
rect 17740 6639 17792 6645
rect 17924 6639 17954 6687
rect 18045 6645 18075 6677
rect 17740 6629 17954 6639
rect 17740 6595 17750 6629
rect 17784 6595 17954 6629
rect 17740 6585 17954 6595
rect 17277 6511 17307 6543
rect 17667 6511 17697 6583
rect 17740 6579 17792 6585
rect 17762 6557 17792 6579
rect 17924 6556 17954 6585
rect 18016 6629 18075 6645
rect 18016 6595 18026 6629
rect 18060 6595 18075 6629
rect 18016 6579 18075 6595
rect 18045 6557 18075 6579
rect 17924 6526 17980 6556
rect 17950 6511 17980 6526
rect 13449 6401 13479 6427
rect 13533 6401 13563 6427
rect 13721 6401 13751 6427
rect 13816 6401 13846 6427
rect 13922 6401 13952 6427
rect 14018 6401 14048 6427
rect 14128 6401 14158 6427
rect 14228 6401 14258 6427
rect 14312 6401 14342 6427
rect 14500 6401 14530 6427
rect 14595 6401 14625 6427
rect 14704 6401 14734 6427
rect 14799 6401 14829 6427
rect 14885 6401 14915 6427
rect 15003 6401 15033 6427
rect 15087 6401 15117 6427
rect 15275 6401 15305 6427
rect 15370 6401 15400 6427
rect 15558 6401 15588 6427
rect 15653 6401 15683 6427
rect 15841 6401 15871 6427
rect 15925 6401 15955 6427
rect 16113 6401 16143 6427
rect 16208 6401 16238 6427
rect 16314 6401 16344 6427
rect 16410 6401 16440 6427
rect 16520 6401 16550 6427
rect 16620 6401 16650 6427
rect 16704 6401 16734 6427
rect 16892 6401 16922 6427
rect 16987 6401 17017 6427
rect 17096 6401 17126 6427
rect 17191 6401 17221 6427
rect 17277 6401 17307 6427
rect 17395 6401 17425 6427
rect 17479 6401 17509 6427
rect 17667 6401 17697 6427
rect 17762 6401 17792 6427
rect 17950 6401 17980 6427
rect 18045 6401 18075 6427
rect 13449 6237 13479 6263
rect 13533 6237 13563 6263
rect 13721 6237 13751 6263
rect 13816 6237 13846 6263
rect 13922 6237 13952 6263
rect 14018 6237 14048 6263
rect 14128 6237 14158 6263
rect 14228 6237 14258 6263
rect 14312 6237 14342 6263
rect 14500 6237 14530 6263
rect 14595 6237 14625 6263
rect 14704 6237 14734 6263
rect 14799 6237 14829 6263
rect 14885 6237 14915 6263
rect 15003 6237 15033 6263
rect 15087 6237 15117 6263
rect 15275 6237 15305 6263
rect 15370 6237 15400 6263
rect 15558 6237 15588 6263
rect 15653 6237 15683 6263
rect 15841 6237 15871 6263
rect 15925 6237 15955 6263
rect 16113 6237 16143 6263
rect 16208 6237 16238 6263
rect 16314 6237 16344 6263
rect 16410 6237 16440 6263
rect 16520 6237 16550 6263
rect 16620 6237 16650 6263
rect 16704 6237 16734 6263
rect 16892 6237 16922 6263
rect 16987 6237 17017 6263
rect 17096 6237 17126 6263
rect 17191 6237 17221 6263
rect 17277 6237 17307 6263
rect 17395 6237 17425 6263
rect 17479 6237 17509 6263
rect 17667 6237 17697 6263
rect 17762 6237 17792 6263
rect 17950 6237 17980 6263
rect 18045 6237 18075 6263
rect 13449 6138 13479 6153
rect 13416 6108 13479 6138
rect 13416 6070 13446 6108
rect 13391 6054 13446 6070
rect 13533 6064 13563 6153
rect 13721 6083 13751 6153
rect 13816 6143 13846 6165
rect 13816 6127 13880 6143
rect 13816 6093 13836 6127
rect 13870 6093 13880 6127
rect 13391 6020 13402 6054
rect 13436 6020 13446 6054
rect 13391 6004 13446 6020
rect 13488 6054 13563 6064
rect 13488 6020 13504 6054
rect 13538 6020 13563 6054
rect 13488 6010 13563 6020
rect 13710 6067 13764 6083
rect 13816 6077 13880 6093
rect 13922 6131 13952 6165
rect 13922 6115 13976 6131
rect 13922 6081 13932 6115
rect 13966 6081 13976 6115
rect 13710 6033 13720 6067
rect 13754 6033 13764 6067
rect 13922 6065 13976 6081
rect 13922 6035 13952 6065
rect 13710 6017 13764 6033
rect 13416 5966 13446 6004
rect 13416 5936 13479 5966
rect 13449 5921 13479 5936
rect 13533 5921 13563 6010
rect 13721 5871 13751 6017
rect 13814 6005 13952 6035
rect 13814 5871 13844 6005
rect 14018 5969 14048 6153
rect 14128 6121 14158 6153
rect 14094 6105 14158 6121
rect 14595 6143 14625 6165
rect 14595 6127 14662 6143
rect 14094 6071 14104 6105
rect 14138 6091 14158 6105
rect 14138 6071 14154 6091
rect 14094 6055 14154 6071
rect 13886 5953 13952 5963
rect 13886 5919 13902 5953
rect 13936 5919 13952 5953
rect 13886 5909 13952 5919
rect 14018 5953 14082 5969
rect 14018 5919 14038 5953
rect 14072 5919 14082 5953
rect 13898 5871 13928 5909
rect 14018 5903 14082 5919
rect 14018 5871 14048 5903
rect 14124 5871 14154 6055
rect 14228 6053 14258 6109
rect 14312 6053 14342 6109
rect 14500 6087 14530 6109
rect 14476 6071 14530 6087
rect 14595 6093 14618 6127
rect 14652 6093 14662 6127
rect 14595 6077 14662 6093
rect 14196 6037 14262 6053
rect 14196 6003 14206 6037
rect 14240 6003 14262 6037
rect 14196 5987 14262 6003
rect 14312 6037 14402 6053
rect 14476 6051 14486 6071
rect 14312 6003 14358 6037
rect 14392 6003 14402 6037
rect 14312 5987 14402 6003
rect 14453 6037 14486 6051
rect 14520 6037 14530 6071
rect 14453 6021 14530 6037
rect 14704 6035 14734 6165
rect 14232 5955 14262 5987
rect 14316 5955 14346 5987
rect 14453 5955 14483 6021
rect 14597 6005 14734 6035
rect 14597 5969 14627 6005
rect 13449 5767 13479 5793
rect 13533 5767 13563 5793
rect 14573 5953 14627 5969
rect 14799 5969 14829 6153
rect 14885 6121 14915 6153
rect 14871 6105 14937 6121
rect 14871 6071 14881 6105
rect 14915 6071 14937 6105
rect 14871 6055 14937 6071
rect 15003 6069 15033 6109
rect 14573 5919 14583 5953
rect 14617 5919 14627 5953
rect 14573 5903 14627 5919
rect 14669 5953 14735 5963
rect 14669 5919 14685 5953
rect 14719 5919 14735 5953
rect 14669 5909 14735 5919
rect 14799 5953 14865 5969
rect 14799 5919 14821 5953
rect 14855 5919 14865 5953
rect 14597 5871 14627 5903
rect 14681 5871 14711 5909
rect 14799 5903 14865 5919
rect 14799 5871 14829 5903
rect 14907 5871 14937 6055
rect 14979 6053 15033 6069
rect 14979 6019 14989 6053
rect 15023 6019 15033 6053
rect 14979 6003 15033 6019
rect 15087 6053 15117 6109
rect 15275 6081 15305 6153
rect 15558 6138 15588 6153
rect 15532 6108 15588 6138
rect 15370 6085 15400 6107
rect 15242 6065 15306 6081
rect 15087 6037 15171 6053
rect 15087 6017 15127 6037
rect 15003 5955 15033 6003
rect 15075 6003 15127 6017
rect 15161 6003 15171 6037
rect 15242 6031 15258 6065
rect 15292 6031 15306 6065
rect 15242 6015 15306 6031
rect 15348 6079 15400 6085
rect 15532 6079 15562 6108
rect 15841 6138 15871 6153
rect 15808 6108 15871 6138
rect 15653 6085 15683 6107
rect 15348 6069 15562 6079
rect 15348 6035 15358 6069
rect 15392 6035 15562 6069
rect 15348 6025 15562 6035
rect 15348 6019 15400 6025
rect 15075 5987 15171 6003
rect 15075 5955 15105 5987
rect 15273 5983 15303 6015
rect 15370 5987 15400 6019
rect 15273 5829 15303 5855
rect 15532 5977 15562 6025
rect 15624 6069 15683 6085
rect 15808 6070 15838 6108
rect 15624 6035 15634 6069
rect 15668 6035 15683 6069
rect 15624 6019 15683 6035
rect 15653 5987 15683 6019
rect 15783 6054 15838 6070
rect 15925 6064 15955 6153
rect 16113 6083 16143 6153
rect 16208 6143 16238 6165
rect 16208 6127 16272 6143
rect 16208 6093 16228 6127
rect 16262 6093 16272 6127
rect 15783 6020 15794 6054
rect 15828 6020 15838 6054
rect 15783 6004 15838 6020
rect 15880 6054 15955 6064
rect 15880 6020 15896 6054
rect 15930 6020 15955 6054
rect 15880 6010 15955 6020
rect 16102 6067 16156 6083
rect 16208 6077 16272 6093
rect 16314 6131 16344 6165
rect 16314 6115 16368 6131
rect 16314 6081 16324 6115
rect 16358 6081 16368 6115
rect 16102 6033 16112 6067
rect 16146 6033 16156 6067
rect 16314 6065 16368 6081
rect 16314 6035 16344 6065
rect 16102 6017 16156 6033
rect 15532 5947 15588 5977
rect 15558 5931 15588 5947
rect 13721 5761 13751 5787
rect 13814 5761 13844 5787
rect 13898 5761 13928 5787
rect 14018 5761 14048 5787
rect 14124 5761 14154 5787
rect 14232 5761 14262 5787
rect 14316 5761 14346 5787
rect 14453 5761 14483 5787
rect 14597 5761 14627 5787
rect 14681 5761 14711 5787
rect 14799 5761 14829 5787
rect 14907 5761 14937 5787
rect 15003 5761 15033 5787
rect 15075 5761 15105 5787
rect 15370 5761 15400 5787
rect 15558 5777 15588 5803
rect 15808 5966 15838 6004
rect 15808 5936 15871 5966
rect 15841 5921 15871 5936
rect 15925 5921 15955 6010
rect 16113 5871 16143 6017
rect 16206 6005 16344 6035
rect 16206 5871 16236 6005
rect 16410 5969 16440 6153
rect 16520 6121 16550 6153
rect 16486 6105 16550 6121
rect 16987 6143 17017 6165
rect 16987 6127 17054 6143
rect 16486 6071 16496 6105
rect 16530 6091 16550 6105
rect 16530 6071 16546 6091
rect 16486 6055 16546 6071
rect 16278 5953 16344 5963
rect 16278 5919 16294 5953
rect 16328 5919 16344 5953
rect 16278 5909 16344 5919
rect 16410 5953 16474 5969
rect 16410 5919 16430 5953
rect 16464 5919 16474 5953
rect 16290 5871 16320 5909
rect 16410 5903 16474 5919
rect 16410 5871 16440 5903
rect 16516 5871 16546 6055
rect 16620 6053 16650 6109
rect 16704 6053 16734 6109
rect 16892 6087 16922 6109
rect 16868 6071 16922 6087
rect 16987 6093 17010 6127
rect 17044 6093 17054 6127
rect 16987 6077 17054 6093
rect 16588 6037 16654 6053
rect 16588 6003 16598 6037
rect 16632 6003 16654 6037
rect 16588 5987 16654 6003
rect 16704 6037 16794 6053
rect 16868 6051 16878 6071
rect 16704 6003 16750 6037
rect 16784 6003 16794 6037
rect 16704 5987 16794 6003
rect 16845 6037 16878 6051
rect 16912 6037 16922 6071
rect 16845 6021 16922 6037
rect 17096 6035 17126 6165
rect 16624 5955 16654 5987
rect 16708 5955 16738 5987
rect 16845 5955 16875 6021
rect 16989 6005 17126 6035
rect 16989 5969 17019 6005
rect 15653 5761 15683 5787
rect 15841 5767 15871 5793
rect 15925 5767 15955 5793
rect 16965 5953 17019 5969
rect 17191 5969 17221 6153
rect 17277 6121 17307 6153
rect 17263 6105 17329 6121
rect 17263 6071 17273 6105
rect 17307 6071 17329 6105
rect 17263 6055 17329 6071
rect 17395 6069 17425 6109
rect 16965 5919 16975 5953
rect 17009 5919 17019 5953
rect 16965 5903 17019 5919
rect 17061 5953 17127 5963
rect 17061 5919 17077 5953
rect 17111 5919 17127 5953
rect 17061 5909 17127 5919
rect 17191 5953 17257 5969
rect 17191 5919 17213 5953
rect 17247 5919 17257 5953
rect 16989 5871 17019 5903
rect 17073 5871 17103 5909
rect 17191 5903 17257 5919
rect 17191 5871 17221 5903
rect 17299 5871 17329 6055
rect 17371 6053 17425 6069
rect 17371 6019 17381 6053
rect 17415 6019 17425 6053
rect 17371 6003 17425 6019
rect 17479 6053 17509 6109
rect 17667 6081 17697 6153
rect 17950 6138 17980 6153
rect 17924 6108 17980 6138
rect 17762 6085 17792 6107
rect 17634 6065 17698 6081
rect 17479 6037 17563 6053
rect 17479 6017 17519 6037
rect 17395 5955 17425 6003
rect 17467 6003 17519 6017
rect 17553 6003 17563 6037
rect 17634 6031 17650 6065
rect 17684 6031 17698 6065
rect 17634 6015 17698 6031
rect 17740 6079 17792 6085
rect 17924 6079 17954 6108
rect 18045 6085 18075 6107
rect 17740 6069 17954 6079
rect 17740 6035 17750 6069
rect 17784 6035 17954 6069
rect 17740 6025 17954 6035
rect 17740 6019 17792 6025
rect 17467 5987 17563 6003
rect 17467 5955 17497 5987
rect 17665 5983 17695 6015
rect 17762 5987 17792 6019
rect 17665 5829 17695 5855
rect 17924 5977 17954 6025
rect 18016 6069 18075 6085
rect 18016 6035 18026 6069
rect 18060 6035 18075 6069
rect 18016 6019 18075 6035
rect 18045 5987 18075 6019
rect 17924 5947 17980 5977
rect 17950 5931 17980 5947
rect 16113 5761 16143 5787
rect 16206 5761 16236 5787
rect 16290 5761 16320 5787
rect 16410 5761 16440 5787
rect 16516 5761 16546 5787
rect 16624 5761 16654 5787
rect 16708 5761 16738 5787
rect 16845 5761 16875 5787
rect 16989 5761 17019 5787
rect 17073 5761 17103 5787
rect 17191 5761 17221 5787
rect 17299 5761 17329 5787
rect 17395 5761 17425 5787
rect 17467 5761 17497 5787
rect 17762 5761 17792 5787
rect 17950 5777 17980 5803
rect 18045 5761 18075 5787
rect 13449 5591 13479 5617
rect 13533 5591 13563 5617
rect 13721 5597 13751 5623
rect 13814 5597 13844 5623
rect 13898 5597 13928 5623
rect 14018 5597 14048 5623
rect 14124 5597 14154 5623
rect 14232 5597 14262 5623
rect 14316 5597 14346 5623
rect 14453 5597 14483 5623
rect 14597 5597 14627 5623
rect 14681 5597 14711 5623
rect 14799 5597 14829 5623
rect 14907 5597 14937 5623
rect 15003 5597 15033 5623
rect 15075 5597 15105 5623
rect 15370 5597 15400 5623
rect 13449 5448 13479 5463
rect 13416 5418 13479 5448
rect 13416 5380 13446 5418
rect 13391 5364 13446 5380
rect 13533 5374 13563 5463
rect 13391 5330 13402 5364
rect 13436 5330 13446 5364
rect 13391 5314 13446 5330
rect 13488 5364 13563 5374
rect 13721 5367 13751 5513
rect 13814 5379 13844 5513
rect 13898 5475 13928 5513
rect 14018 5481 14048 5513
rect 13886 5465 13952 5475
rect 13886 5431 13902 5465
rect 13936 5431 13952 5465
rect 13886 5421 13952 5431
rect 14018 5465 14082 5481
rect 14018 5431 14038 5465
rect 14072 5431 14082 5465
rect 14018 5415 14082 5431
rect 13488 5330 13504 5364
rect 13538 5330 13563 5364
rect 13488 5320 13563 5330
rect 13416 5276 13446 5314
rect 13416 5246 13479 5276
rect 13449 5231 13479 5246
rect 13533 5231 13563 5320
rect 13710 5351 13764 5367
rect 13710 5317 13720 5351
rect 13754 5317 13764 5351
rect 13814 5349 13952 5379
rect 13710 5301 13764 5317
rect 13922 5319 13952 5349
rect 13721 5231 13751 5301
rect 13816 5291 13880 5307
rect 13816 5257 13836 5291
rect 13870 5257 13880 5291
rect 13816 5241 13880 5257
rect 13922 5303 13976 5319
rect 13922 5269 13932 5303
rect 13966 5269 13976 5303
rect 13922 5253 13976 5269
rect 13816 5219 13846 5241
rect 13922 5219 13952 5253
rect 14018 5231 14048 5415
rect 14124 5329 14154 5513
rect 14597 5481 14627 5513
rect 14573 5465 14627 5481
rect 14681 5475 14711 5513
rect 14799 5481 14829 5513
rect 14573 5431 14583 5465
rect 14617 5431 14627 5465
rect 14232 5397 14262 5429
rect 14316 5397 14346 5429
rect 14196 5381 14262 5397
rect 14196 5347 14206 5381
rect 14240 5347 14262 5381
rect 14196 5331 14262 5347
rect 14312 5381 14402 5397
rect 14312 5347 14358 5381
rect 14392 5347 14402 5381
rect 14312 5331 14402 5347
rect 14453 5363 14483 5429
rect 14573 5415 14627 5431
rect 14669 5465 14735 5475
rect 14669 5431 14685 5465
rect 14719 5431 14735 5465
rect 14669 5421 14735 5431
rect 14799 5465 14865 5481
rect 14799 5431 14821 5465
rect 14855 5431 14865 5465
rect 14597 5379 14627 5415
rect 14799 5415 14865 5431
rect 14453 5347 14530 5363
rect 14597 5349 14734 5379
rect 14453 5333 14486 5347
rect 14094 5313 14154 5329
rect 14094 5279 14104 5313
rect 14138 5293 14154 5313
rect 14138 5279 14158 5293
rect 14094 5263 14158 5279
rect 14228 5275 14258 5331
rect 14312 5275 14342 5331
rect 14476 5313 14486 5333
rect 14520 5313 14530 5347
rect 14476 5297 14530 5313
rect 14500 5275 14530 5297
rect 14595 5291 14662 5307
rect 14128 5231 14158 5263
rect 14595 5257 14618 5291
rect 14652 5257 14662 5291
rect 14595 5241 14662 5257
rect 14595 5219 14625 5241
rect 14704 5219 14734 5349
rect 14799 5231 14829 5415
rect 14907 5329 14937 5513
rect 15273 5529 15303 5555
rect 15003 5381 15033 5429
rect 14871 5313 14937 5329
rect 14979 5365 15033 5381
rect 15075 5397 15105 5429
rect 15075 5381 15171 5397
rect 15075 5367 15127 5381
rect 14979 5331 14989 5365
rect 15023 5331 15033 5365
rect 14979 5315 15033 5331
rect 14871 5279 14881 5313
rect 14915 5279 14937 5313
rect 14871 5263 14937 5279
rect 15003 5275 15033 5315
rect 15087 5347 15127 5367
rect 15161 5347 15171 5381
rect 15273 5369 15303 5401
rect 15558 5581 15588 5607
rect 15653 5597 15683 5623
rect 15558 5437 15588 5453
rect 15532 5407 15588 5437
rect 15087 5331 15171 5347
rect 15242 5353 15306 5369
rect 15370 5365 15400 5397
rect 15087 5275 15117 5331
rect 15242 5319 15258 5353
rect 15292 5319 15306 5353
rect 15242 5303 15306 5319
rect 15348 5359 15400 5365
rect 15532 5359 15562 5407
rect 15841 5591 15871 5617
rect 15925 5591 15955 5617
rect 16113 5597 16143 5623
rect 16206 5597 16236 5623
rect 16290 5597 16320 5623
rect 16410 5597 16440 5623
rect 16516 5597 16546 5623
rect 16624 5597 16654 5623
rect 16708 5597 16738 5623
rect 16845 5597 16875 5623
rect 16989 5597 17019 5623
rect 17073 5597 17103 5623
rect 17191 5597 17221 5623
rect 17299 5597 17329 5623
rect 17395 5597 17425 5623
rect 17467 5597 17497 5623
rect 17762 5597 17792 5623
rect 15841 5448 15871 5463
rect 15808 5418 15871 5448
rect 15653 5365 15683 5397
rect 15808 5380 15838 5418
rect 15348 5349 15562 5359
rect 15348 5315 15358 5349
rect 15392 5315 15562 5349
rect 15348 5305 15562 5315
rect 14885 5231 14915 5263
rect 15275 5231 15305 5303
rect 15348 5299 15400 5305
rect 15370 5277 15400 5299
rect 15532 5276 15562 5305
rect 15624 5349 15683 5365
rect 15624 5315 15634 5349
rect 15668 5315 15683 5349
rect 15624 5299 15683 5315
rect 15783 5364 15838 5380
rect 15925 5374 15955 5463
rect 15783 5330 15794 5364
rect 15828 5330 15838 5364
rect 15783 5314 15838 5330
rect 15880 5364 15955 5374
rect 16113 5367 16143 5513
rect 16206 5379 16236 5513
rect 16290 5475 16320 5513
rect 16410 5481 16440 5513
rect 16278 5465 16344 5475
rect 16278 5431 16294 5465
rect 16328 5431 16344 5465
rect 16278 5421 16344 5431
rect 16410 5465 16474 5481
rect 16410 5431 16430 5465
rect 16464 5431 16474 5465
rect 16410 5415 16474 5431
rect 15880 5330 15896 5364
rect 15930 5330 15955 5364
rect 15880 5320 15955 5330
rect 15653 5277 15683 5299
rect 15532 5246 15588 5276
rect 15558 5231 15588 5246
rect 15808 5276 15838 5314
rect 15808 5246 15871 5276
rect 15841 5231 15871 5246
rect 15925 5231 15955 5320
rect 16102 5351 16156 5367
rect 16102 5317 16112 5351
rect 16146 5317 16156 5351
rect 16206 5349 16344 5379
rect 16102 5301 16156 5317
rect 16314 5319 16344 5349
rect 16113 5231 16143 5301
rect 16208 5291 16272 5307
rect 16208 5257 16228 5291
rect 16262 5257 16272 5291
rect 16208 5241 16272 5257
rect 16314 5303 16368 5319
rect 16314 5269 16324 5303
rect 16358 5269 16368 5303
rect 16314 5253 16368 5269
rect 16208 5219 16238 5241
rect 16314 5219 16344 5253
rect 16410 5231 16440 5415
rect 16516 5329 16546 5513
rect 16989 5481 17019 5513
rect 16965 5465 17019 5481
rect 17073 5475 17103 5513
rect 17191 5481 17221 5513
rect 16965 5431 16975 5465
rect 17009 5431 17019 5465
rect 16624 5397 16654 5429
rect 16708 5397 16738 5429
rect 16588 5381 16654 5397
rect 16588 5347 16598 5381
rect 16632 5347 16654 5381
rect 16588 5331 16654 5347
rect 16704 5381 16794 5397
rect 16704 5347 16750 5381
rect 16784 5347 16794 5381
rect 16704 5331 16794 5347
rect 16845 5363 16875 5429
rect 16965 5415 17019 5431
rect 17061 5465 17127 5475
rect 17061 5431 17077 5465
rect 17111 5431 17127 5465
rect 17061 5421 17127 5431
rect 17191 5465 17257 5481
rect 17191 5431 17213 5465
rect 17247 5431 17257 5465
rect 16989 5379 17019 5415
rect 17191 5415 17257 5431
rect 16845 5347 16922 5363
rect 16989 5349 17126 5379
rect 16845 5333 16878 5347
rect 16486 5313 16546 5329
rect 16486 5279 16496 5313
rect 16530 5293 16546 5313
rect 16530 5279 16550 5293
rect 16486 5263 16550 5279
rect 16620 5275 16650 5331
rect 16704 5275 16734 5331
rect 16868 5313 16878 5333
rect 16912 5313 16922 5347
rect 16868 5297 16922 5313
rect 16892 5275 16922 5297
rect 16987 5291 17054 5307
rect 16520 5231 16550 5263
rect 16987 5257 17010 5291
rect 17044 5257 17054 5291
rect 16987 5241 17054 5257
rect 16987 5219 17017 5241
rect 17096 5219 17126 5349
rect 17191 5231 17221 5415
rect 17299 5329 17329 5513
rect 17665 5529 17695 5555
rect 17395 5381 17425 5429
rect 17263 5313 17329 5329
rect 17371 5365 17425 5381
rect 17467 5397 17497 5429
rect 17467 5381 17563 5397
rect 17467 5367 17519 5381
rect 17371 5331 17381 5365
rect 17415 5331 17425 5365
rect 17371 5315 17425 5331
rect 17263 5279 17273 5313
rect 17307 5279 17329 5313
rect 17263 5263 17329 5279
rect 17395 5275 17425 5315
rect 17479 5347 17519 5367
rect 17553 5347 17563 5381
rect 17665 5369 17695 5401
rect 17950 5581 17980 5607
rect 18045 5597 18075 5623
rect 17950 5437 17980 5453
rect 17924 5407 17980 5437
rect 17479 5331 17563 5347
rect 17634 5353 17698 5369
rect 17762 5365 17792 5397
rect 17479 5275 17509 5331
rect 17634 5319 17650 5353
rect 17684 5319 17698 5353
rect 17634 5303 17698 5319
rect 17740 5359 17792 5365
rect 17924 5359 17954 5407
rect 18045 5365 18075 5397
rect 17740 5349 17954 5359
rect 17740 5315 17750 5349
rect 17784 5315 17954 5349
rect 17740 5305 17954 5315
rect 17277 5231 17307 5263
rect 17667 5231 17697 5303
rect 17740 5299 17792 5305
rect 17762 5277 17792 5299
rect 17924 5276 17954 5305
rect 18016 5349 18075 5365
rect 18016 5315 18026 5349
rect 18060 5315 18075 5349
rect 18016 5299 18075 5315
rect 18045 5277 18075 5299
rect 17924 5246 17980 5276
rect 17950 5231 17980 5246
rect 13449 5121 13479 5147
rect 13533 5121 13563 5147
rect 13721 5121 13751 5147
rect 13816 5121 13846 5147
rect 13922 5121 13952 5147
rect 14018 5121 14048 5147
rect 14128 5121 14158 5147
rect 14228 5121 14258 5147
rect 14312 5121 14342 5147
rect 14500 5121 14530 5147
rect 14595 5121 14625 5147
rect 14704 5121 14734 5147
rect 14799 5121 14829 5147
rect 14885 5121 14915 5147
rect 15003 5121 15033 5147
rect 15087 5121 15117 5147
rect 15275 5121 15305 5147
rect 15370 5121 15400 5147
rect 15558 5121 15588 5147
rect 15653 5121 15683 5147
rect 15841 5121 15871 5147
rect 15925 5121 15955 5147
rect 16113 5121 16143 5147
rect 16208 5121 16238 5147
rect 16314 5121 16344 5147
rect 16410 5121 16440 5147
rect 16520 5121 16550 5147
rect 16620 5121 16650 5147
rect 16704 5121 16734 5147
rect 16892 5121 16922 5147
rect 16987 5121 17017 5147
rect 17096 5121 17126 5147
rect 17191 5121 17221 5147
rect 17277 5121 17307 5147
rect 17395 5121 17425 5147
rect 17479 5121 17509 5147
rect 17667 5121 17697 5147
rect 17762 5121 17792 5147
rect 17950 5121 17980 5147
rect 18045 5121 18075 5147
<< polycont >>
rect 11872 9650 11906 9684
rect 12378 9724 12412 9758
rect 12138 9650 12172 9684
rect 13020 9481 13054 9515
rect 13752 9484 13786 9518
rect 13878 9484 13912 9518
rect 14964 9484 14998 9518
rect 15090 9484 15124 9518
rect 16176 9484 16210 9518
rect 16302 9484 16336 9518
rect 17388 9484 17422 9518
rect 17514 9484 17548 9518
rect 18048 9277 18082 9311
rect 18255 9275 18289 9309
rect 18509 9273 18543 9307
rect 18633 9273 18667 9307
rect 12389 9090 12423 9124
rect 13373 9080 13407 9114
rect 14105 9080 14139 9114
rect 14227 9080 14261 9114
rect 15317 9080 15351 9114
rect 15439 9080 15473 9114
rect 16655 9080 16689 9114
rect 16777 9080 16811 9114
rect 17511 9080 17545 9114
rect 13836 7373 13870 7407
rect 13402 7300 13436 7334
rect 13504 7300 13538 7334
rect 13932 7361 13966 7395
rect 13720 7313 13754 7347
rect 14104 7351 14138 7385
rect 13902 7199 13936 7233
rect 14038 7199 14072 7233
rect 14618 7373 14652 7407
rect 14206 7283 14240 7317
rect 14358 7283 14392 7317
rect 14486 7317 14520 7351
rect 14881 7351 14915 7385
rect 14583 7199 14617 7233
rect 14685 7199 14719 7233
rect 14821 7199 14855 7233
rect 14989 7299 15023 7333
rect 15127 7283 15161 7317
rect 15258 7311 15292 7345
rect 15358 7315 15392 7349
rect 15634 7315 15668 7349
rect 16228 7373 16262 7407
rect 15794 7300 15828 7334
rect 15896 7300 15930 7334
rect 16324 7361 16358 7395
rect 16112 7313 16146 7347
rect 16496 7351 16530 7385
rect 16294 7199 16328 7233
rect 16430 7199 16464 7233
rect 17010 7373 17044 7407
rect 16598 7283 16632 7317
rect 16750 7283 16784 7317
rect 16878 7317 16912 7351
rect 17273 7351 17307 7385
rect 16975 7199 17009 7233
rect 17077 7199 17111 7233
rect 17213 7199 17247 7233
rect 17381 7299 17415 7333
rect 17519 7283 17553 7317
rect 17650 7311 17684 7345
rect 17750 7315 17784 7349
rect 18026 7315 18060 7349
rect 13402 6610 13436 6644
rect 13902 6711 13936 6745
rect 14038 6711 14072 6745
rect 13504 6610 13538 6644
rect 13720 6597 13754 6631
rect 13836 6537 13870 6571
rect 13932 6549 13966 6583
rect 14583 6711 14617 6745
rect 14206 6627 14240 6661
rect 14358 6627 14392 6661
rect 14685 6711 14719 6745
rect 14821 6711 14855 6745
rect 14104 6559 14138 6593
rect 14486 6593 14520 6627
rect 14618 6537 14652 6571
rect 14989 6611 15023 6645
rect 14881 6559 14915 6593
rect 15127 6627 15161 6661
rect 15258 6599 15292 6633
rect 15358 6595 15392 6629
rect 15634 6595 15668 6629
rect 15794 6610 15828 6644
rect 16294 6711 16328 6745
rect 16430 6711 16464 6745
rect 15896 6610 15930 6644
rect 16112 6597 16146 6631
rect 16228 6537 16262 6571
rect 16324 6549 16358 6583
rect 16975 6711 17009 6745
rect 16598 6627 16632 6661
rect 16750 6627 16784 6661
rect 17077 6711 17111 6745
rect 17213 6711 17247 6745
rect 16496 6559 16530 6593
rect 16878 6593 16912 6627
rect 17010 6537 17044 6571
rect 17381 6611 17415 6645
rect 17273 6559 17307 6593
rect 17519 6627 17553 6661
rect 17650 6599 17684 6633
rect 17750 6595 17784 6629
rect 18026 6595 18060 6629
rect 13836 6093 13870 6127
rect 13402 6020 13436 6054
rect 13504 6020 13538 6054
rect 13932 6081 13966 6115
rect 13720 6033 13754 6067
rect 14104 6071 14138 6105
rect 13902 5919 13936 5953
rect 14038 5919 14072 5953
rect 14618 6093 14652 6127
rect 14206 6003 14240 6037
rect 14358 6003 14392 6037
rect 14486 6037 14520 6071
rect 14881 6071 14915 6105
rect 14583 5919 14617 5953
rect 14685 5919 14719 5953
rect 14821 5919 14855 5953
rect 14989 6019 15023 6053
rect 15127 6003 15161 6037
rect 15258 6031 15292 6065
rect 15358 6035 15392 6069
rect 15634 6035 15668 6069
rect 16228 6093 16262 6127
rect 15794 6020 15828 6054
rect 15896 6020 15930 6054
rect 16324 6081 16358 6115
rect 16112 6033 16146 6067
rect 16496 6071 16530 6105
rect 16294 5919 16328 5953
rect 16430 5919 16464 5953
rect 17010 6093 17044 6127
rect 16598 6003 16632 6037
rect 16750 6003 16784 6037
rect 16878 6037 16912 6071
rect 17273 6071 17307 6105
rect 16975 5919 17009 5953
rect 17077 5919 17111 5953
rect 17213 5919 17247 5953
rect 17381 6019 17415 6053
rect 17519 6003 17553 6037
rect 17650 6031 17684 6065
rect 17750 6035 17784 6069
rect 18026 6035 18060 6069
rect 13402 5330 13436 5364
rect 13902 5431 13936 5465
rect 14038 5431 14072 5465
rect 13504 5330 13538 5364
rect 13720 5317 13754 5351
rect 13836 5257 13870 5291
rect 13932 5269 13966 5303
rect 14583 5431 14617 5465
rect 14206 5347 14240 5381
rect 14358 5347 14392 5381
rect 14685 5431 14719 5465
rect 14821 5431 14855 5465
rect 14104 5279 14138 5313
rect 14486 5313 14520 5347
rect 14618 5257 14652 5291
rect 14989 5331 15023 5365
rect 14881 5279 14915 5313
rect 15127 5347 15161 5381
rect 15258 5319 15292 5353
rect 15358 5315 15392 5349
rect 15634 5315 15668 5349
rect 15794 5330 15828 5364
rect 16294 5431 16328 5465
rect 16430 5431 16464 5465
rect 15896 5330 15930 5364
rect 16112 5317 16146 5351
rect 16228 5257 16262 5291
rect 16324 5269 16358 5303
rect 16975 5431 17009 5465
rect 16598 5347 16632 5381
rect 16750 5347 16784 5381
rect 17077 5431 17111 5465
rect 17213 5431 17247 5465
rect 16496 5279 16530 5313
rect 16878 5313 16912 5347
rect 17010 5257 17044 5291
rect 17381 5331 17415 5365
rect 17273 5279 17307 5313
rect 17519 5347 17553 5381
rect 17650 5319 17684 5353
rect 17750 5315 17784 5349
rect 18026 5315 18060 5349
<< locali >>
rect 12464 10591 13134 10609
rect 12464 10583 12580 10591
rect 12334 10567 12368 10583
rect 12334 10491 12368 10507
rect 12422 10567 12580 10583
rect 12456 10557 12580 10567
rect 12616 10557 12660 10591
rect 12696 10557 12740 10591
rect 12776 10557 12820 10591
rect 12856 10557 12900 10591
rect 12936 10557 12980 10591
rect 13016 10557 13134 10591
rect 12456 10543 13134 10557
rect 13196 10594 18104 10612
rect 13196 10560 13312 10594
rect 13348 10560 13392 10594
rect 13428 10560 13472 10594
rect 13508 10560 13552 10594
rect 13588 10560 13632 10594
rect 13668 10560 13712 10594
rect 13748 10560 13916 10594
rect 13952 10560 13996 10594
rect 14032 10560 14076 10594
rect 14112 10560 14156 10594
rect 14192 10560 14236 10594
rect 14272 10560 14316 10594
rect 14352 10560 14524 10594
rect 14560 10560 14604 10594
rect 14640 10560 14684 10594
rect 14720 10560 14764 10594
rect 14800 10560 14844 10594
rect 14880 10560 14924 10594
rect 14960 10560 15128 10594
rect 15164 10560 15208 10594
rect 15244 10560 15288 10594
rect 15324 10560 15368 10594
rect 15404 10560 15448 10594
rect 15484 10560 15528 10594
rect 15564 10560 15736 10594
rect 15772 10560 15816 10594
rect 15852 10560 15896 10594
rect 15932 10560 15976 10594
rect 16012 10560 16056 10594
rect 16092 10560 16136 10594
rect 16172 10560 16340 10594
rect 16376 10560 16420 10594
rect 16456 10560 16500 10594
rect 16536 10560 16580 10594
rect 16616 10560 16660 10594
rect 16696 10560 16740 10594
rect 16776 10560 16948 10594
rect 16984 10560 17028 10594
rect 17064 10560 17108 10594
rect 17144 10560 17188 10594
rect 17224 10560 17268 10594
rect 17304 10560 17348 10594
rect 17384 10560 17552 10594
rect 17588 10560 17632 10594
rect 17668 10560 17712 10594
rect 17748 10560 17792 10594
rect 17828 10560 17872 10594
rect 17908 10560 17952 10594
rect 17988 10560 18104 10594
rect 13196 10546 18104 10560
rect 18268 10543 18354 10569
rect 12456 10507 12592 10543
rect 12422 10502 12592 10507
rect 12422 10491 12456 10502
rect 12334 10429 12368 10445
rect 12334 10353 12368 10369
rect 12422 10429 12456 10445
rect 12535 10438 12592 10502
rect 18268 10509 18294 10543
rect 18328 10509 18354 10543
rect 18268 10483 18354 10509
rect 12422 10353 12456 10369
rect 12522 10413 12605 10438
rect 12522 10378 12547 10413
rect 12581 10378 12605 10413
rect 12522 10354 12605 10378
rect 18273 10399 18359 10425
rect 18273 10365 18299 10399
rect 18333 10365 18359 10399
rect 18273 10339 18359 10365
rect 12334 10291 12368 10307
rect 12334 10215 12368 10231
rect 12422 10291 12456 10307
rect 12422 10215 12456 10231
rect 18274 10247 18360 10273
rect 18274 10213 18300 10247
rect 18334 10213 18360 10247
rect 18274 10187 18360 10213
rect 12334 10153 12368 10169
rect 12334 10077 12368 10093
rect 12422 10153 12456 10169
rect 12422 10077 12456 10093
rect 18274 10077 18360 10103
rect 18274 10043 18300 10077
rect 18334 10043 18360 10077
rect 11850 9996 11866 10025
rect 11792 9962 11821 9996
rect 11855 9991 11866 9996
rect 11900 9996 11916 10025
rect 11980 9996 11996 10025
rect 12030 9996 12050 10025
rect 12126 9996 12142 10025
rect 11900 9991 11913 9996
rect 11855 9962 11913 9991
rect 11947 9991 11996 9996
rect 11947 9962 12005 9991
rect 12039 9962 12097 9996
rect 12131 9991 12142 9996
rect 12176 9996 12196 10025
rect 12334 10015 12368 10031
rect 12176 9991 12189 9996
rect 12131 9962 12189 9991
rect 12223 9962 12252 9996
rect 11860 9920 11902 9962
rect 11860 9886 11868 9920
rect 11860 9852 11902 9886
rect 11860 9818 11868 9852
rect 11860 9784 11902 9818
rect 11860 9750 11868 9784
rect 11860 9734 11902 9750
rect 11936 9920 12002 9928
rect 11936 9886 11952 9920
rect 11986 9886 12002 9920
rect 11936 9853 12002 9886
rect 11936 9819 11949 9853
rect 11983 9852 12002 9853
rect 11936 9818 11952 9819
rect 11986 9818 12002 9852
rect 11936 9784 12002 9818
rect 11936 9750 11952 9784
rect 11986 9750 12002 9784
rect 11936 9732 12002 9750
rect 11856 9688 11922 9698
rect 11856 9654 11868 9688
rect 11902 9684 11922 9688
rect 11856 9650 11872 9654
rect 11906 9650 11922 9684
rect 11856 9600 11902 9616
rect 11956 9612 12002 9732
rect 11856 9566 11868 9600
rect 11856 9532 11902 9566
rect 11856 9498 11868 9532
rect 11856 9452 11902 9498
rect 11936 9600 12002 9612
rect 11936 9566 11952 9600
rect 11986 9566 12002 9600
rect 11936 9532 12002 9566
rect 11936 9498 11952 9532
rect 11986 9498 12002 9532
rect 11936 9486 12002 9498
rect 12042 9920 12108 9928
rect 12042 9886 12058 9920
rect 12092 9886 12108 9920
rect 12042 9852 12108 9886
rect 12042 9818 12058 9852
rect 12092 9818 12108 9852
rect 12042 9798 12108 9818
rect 12042 9750 12058 9798
rect 12092 9750 12108 9798
rect 12042 9732 12108 9750
rect 12142 9920 12184 9962
rect 12334 9939 12368 9955
rect 12422 10015 12456 10031
rect 18274 10017 18360 10043
rect 12422 9939 12456 9955
rect 12176 9886 12184 9920
rect 18273 9920 18359 9946
rect 12142 9852 12184 9886
rect 12176 9818 12184 9852
rect 12142 9784 12184 9818
rect 12334 9877 12368 9893
rect 12334 9801 12368 9817
rect 12422 9877 12456 9893
rect 18273 9886 18299 9920
rect 18333 9886 18359 9920
rect 18273 9860 18359 9886
rect 12422 9801 12456 9817
rect 12176 9750 12184 9784
rect 12142 9734 12184 9750
rect 12042 9612 12088 9732
rect 12362 9724 12378 9758
rect 12412 9724 12428 9758
rect 12122 9687 12188 9698
rect 12122 9684 12142 9687
rect 12122 9650 12138 9684
rect 12176 9653 12188 9687
rect 12172 9650 12188 9653
rect 12272 9688 12321 9700
rect 12272 9654 12281 9688
rect 12315 9683 12321 9688
rect 12315 9654 12604 9683
rect 12272 9648 12604 9654
rect 12272 9641 12321 9648
rect 12569 9625 12604 9648
rect 18472 9652 18841 9654
rect 12042 9600 12108 9612
rect 12042 9566 12058 9600
rect 12092 9566 12108 9600
rect 12042 9532 12108 9566
rect 12042 9498 12058 9532
rect 12092 9498 12108 9532
rect 12042 9486 12108 9498
rect 12142 9600 12188 9616
rect 12569 9613 12618 9625
rect 12176 9566 12188 9600
rect 12142 9532 12188 9566
rect 12310 9595 12359 9607
rect 12310 9561 12319 9595
rect 12353 9561 12520 9595
rect 12569 9579 12578 9613
rect 12612 9579 12618 9613
rect 18472 9585 18501 9652
rect 18535 9619 18684 9652
rect 18718 9619 18841 9652
rect 18535 9585 18593 9619
rect 18627 9618 18684 9619
rect 18627 9585 18685 9618
rect 18719 9585 18777 9619
rect 18811 9618 18841 9619
rect 18811 9585 18840 9618
rect 12569 9566 12618 9579
rect 18119 9566 18153 9582
rect 12310 9548 12359 9561
rect 12176 9498 12188 9532
rect 12142 9452 12188 9498
rect 12479 9519 12520 9561
rect 12570 9520 12619 9532
rect 12570 9519 12579 9520
rect 12479 9486 12579 9519
rect 12613 9486 12619 9520
rect 12479 9485 12619 9486
rect 12570 9473 12619 9485
rect 13004 9481 13020 9515
rect 13054 9481 13070 9515
rect 13736 9484 13752 9518
rect 13786 9484 13802 9518
rect 13862 9484 13878 9518
rect 13912 9484 13928 9518
rect 14948 9484 14964 9518
rect 14998 9484 15014 9518
rect 15074 9484 15090 9518
rect 15124 9484 15140 9518
rect 16160 9484 16176 9518
rect 16210 9484 16226 9518
rect 16286 9484 16302 9518
rect 16336 9484 16352 9518
rect 17372 9484 17388 9518
rect 17422 9484 17438 9518
rect 17498 9484 17514 9518
rect 17548 9484 17564 9518
rect 18119 9490 18153 9506
rect 18207 9566 18241 9582
rect 18207 9490 18241 9506
rect 18507 9535 18541 9551
rect 18507 9467 18541 9501
rect 11792 9418 11821 9452
rect 11855 9423 11913 9452
rect 11947 9423 12005 9452
rect 11855 9418 11886 9423
rect 11947 9418 12004 9423
rect 12039 9418 12097 9452
rect 12131 9423 12189 9452
rect 12131 9418 12148 9423
rect 11870 9389 11886 9418
rect 11920 9389 11946 9418
rect 11988 9389 12004 9418
rect 12038 9389 12064 9418
rect 12130 9389 12148 9418
rect 12182 9418 12189 9423
rect 12223 9418 12252 9452
rect 12976 9422 13010 9438
rect 12182 9389 12198 9418
rect 12976 9346 13010 9362
rect 13064 9425 13098 9441
rect 13064 9349 13098 9365
rect 13708 9425 13742 9441
rect 13708 9349 13742 9365
rect 13813 9425 13847 9441
rect 13813 9349 13847 9365
rect 13922 9425 13956 9441
rect 13922 9349 13956 9365
rect 14920 9425 14954 9441
rect 14920 9349 14954 9365
rect 15024 9425 15058 9441
rect 15024 9349 15058 9365
rect 15134 9425 15168 9441
rect 15134 9349 15168 9365
rect 16132 9425 16166 9441
rect 16132 9349 16166 9365
rect 16237 9425 16271 9441
rect 16237 9349 16271 9365
rect 16346 9425 16380 9441
rect 16346 9349 16380 9365
rect 17344 9425 17378 9441
rect 17344 9349 17378 9365
rect 17451 9425 17485 9441
rect 17451 9349 17485 9365
rect 17558 9425 17592 9441
rect 17558 9349 17592 9365
rect 18119 9428 18153 9444
rect 18119 9352 18153 9368
rect 18207 9428 18241 9444
rect 18207 9352 18241 9368
rect 18303 9428 18337 9444
rect 18303 9352 18337 9368
rect 18399 9428 18433 9444
rect 18399 9352 18433 9368
rect 18584 9535 18650 9585
rect 18584 9501 18600 9535
rect 18634 9501 18650 9535
rect 18584 9467 18650 9501
rect 18584 9433 18600 9467
rect 18634 9433 18650 9467
rect 18684 9519 18735 9551
rect 18684 9485 18686 9519
rect 18720 9485 18735 9519
rect 18684 9438 18735 9485
rect 18507 9399 18541 9433
rect 18684 9404 18686 9438
rect 18720 9404 18735 9438
rect 18507 9365 18650 9399
rect 18684 9370 18735 9404
rect 18032 9277 18048 9311
rect 18082 9277 18098 9311
rect 18489 9309 18560 9329
rect 18239 9275 18255 9309
rect 18289 9275 18305 9309
rect 18489 9275 18495 9309
rect 18529 9307 18560 9309
rect 18489 9273 18509 9275
rect 18543 9273 18560 9307
rect 18489 9255 18560 9273
rect 18616 9323 18650 9365
rect 18616 9307 18667 9323
rect 18616 9273 18633 9307
rect 18616 9257 18667 9273
rect 18701 9309 18735 9370
rect 18770 9543 18822 9585
rect 18804 9509 18822 9543
rect 18770 9475 18822 9509
rect 18804 9441 18822 9475
rect 18770 9407 18822 9441
rect 18804 9373 18822 9407
rect 18770 9355 18822 9373
rect 18701 9275 18702 9309
rect 13329 9224 13363 9240
rect 13329 9148 13363 9164
rect 13419 9224 13453 9240
rect 13419 9148 13453 9164
rect 14061 9224 14095 9240
rect 14061 9148 14095 9164
rect 14168 9224 14202 9240
rect 14168 9148 14202 9164
rect 14271 9224 14305 9240
rect 14271 9148 14305 9164
rect 15273 9224 15307 9240
rect 15273 9148 15307 9164
rect 15379 9224 15413 9240
rect 15379 9148 15413 9164
rect 15483 9224 15517 9240
rect 15483 9148 15517 9164
rect 16611 9224 16645 9240
rect 16611 9148 16645 9164
rect 16719 9224 16753 9240
rect 16719 9148 16753 9164
rect 16821 9224 16855 9240
rect 16821 9148 16855 9164
rect 17466 9224 17500 9240
rect 17466 9148 17500 9164
rect 17555 9224 17589 9240
rect 17555 9148 17589 9164
rect 18119 9225 18153 9241
rect 18119 9149 18153 9165
rect 18207 9225 18241 9241
rect 18207 9149 18241 9165
rect 18303 9225 18337 9241
rect 18303 9149 18337 9165
rect 18399 9225 18433 9241
rect 18616 9219 18650 9257
rect 18701 9224 18735 9275
rect 18399 9149 18433 9165
rect 18507 9185 18650 9219
rect 18507 9164 18541 9185
rect 18684 9181 18735 9224
rect 12373 9090 12389 9124
rect 12423 9090 12439 9124
rect 13357 9080 13373 9114
rect 13407 9080 13423 9114
rect 14089 9080 14105 9114
rect 14139 9080 14155 9114
rect 14211 9080 14227 9114
rect 14261 9080 14277 9114
rect 15301 9080 15317 9114
rect 15351 9080 15367 9114
rect 15423 9080 15439 9114
rect 15473 9080 15489 9114
rect 16639 9080 16655 9114
rect 16689 9080 16705 9114
rect 16761 9080 16777 9114
rect 16811 9080 16827 9114
rect 17495 9080 17511 9114
rect 17545 9080 17561 9114
rect 18507 9109 18541 9130
rect 18584 9117 18600 9151
rect 18634 9117 18650 9151
rect 18119 9087 18153 9103
rect 12309 9040 12343 9056
rect 12309 8964 12343 8980
rect 12469 9040 12503 9056
rect 18119 9011 18153 9027
rect 18207 9087 18241 9103
rect 18584 9075 18650 9117
rect 18684 9147 18686 9181
rect 18720 9147 18735 9181
rect 18684 9109 18735 9147
rect 18770 9223 18822 9243
rect 18804 9189 18822 9223
rect 18770 9155 18822 9189
rect 18804 9121 18822 9155
rect 18770 9075 18822 9121
rect 18472 9041 18501 9075
rect 18535 9041 18593 9075
rect 18207 9011 18241 9027
rect 18473 9040 18593 9041
rect 18473 9006 18501 9040
rect 18535 9007 18593 9040
rect 18627 9007 18685 9075
rect 18719 9041 18777 9075
rect 18811 9041 18840 9075
rect 18719 9007 18778 9041
rect 18812 9007 18842 9041
rect 18535 9006 18842 9007
rect 18473 9005 18842 9006
rect 12469 8964 12503 8980
rect 12309 8902 12343 8918
rect 12309 8826 12343 8842
rect 12469 8902 12503 8918
rect 12469 8826 12503 8842
rect 12309 8764 12343 8780
rect 12309 8688 12343 8704
rect 12469 8764 12503 8780
rect 12469 8688 12503 8704
rect 12309 8626 12343 8642
rect 12309 8550 12343 8566
rect 12469 8626 12503 8642
rect 12469 8550 12503 8566
rect 12309 8488 12343 8504
rect 12309 8412 12343 8428
rect 12469 8488 12503 8504
rect 12469 8412 12503 8428
rect 12309 8350 12343 8366
rect 12309 8274 12343 8290
rect 12469 8350 12503 8366
rect 12469 8274 12503 8290
rect 12309 8212 12343 8228
rect 12309 8136 12343 8152
rect 12469 8212 12503 8228
rect 12469 8136 12503 8152
rect 12585 8198 12690 8233
rect 12585 8164 12617 8198
rect 12651 8164 12690 8198
rect 12585 8135 12690 8164
rect 12309 8074 12343 8090
rect 12309 7998 12343 8014
rect 12469 8080 12503 8090
rect 12599 8080 12676 8135
rect 12469 8074 12676 8080
rect 12503 8014 12676 8074
rect 12469 8011 12676 8014
rect 12984 8027 13316 8043
rect 12469 7998 12503 8011
rect 12984 7993 13010 8027
rect 13044 7993 13090 8027
rect 13124 7993 13170 8027
rect 13204 7993 13250 8027
rect 13284 7993 13316 8027
rect 12984 7975 13316 7993
rect 13716 8027 14048 8043
rect 13716 7993 13742 8027
rect 13776 7993 13822 8027
rect 13856 7993 13902 8027
rect 13936 7993 13982 8027
rect 14016 7993 14048 8027
rect 13716 7975 14048 7993
rect 14318 8027 14650 8043
rect 14318 7993 14350 8027
rect 14384 7993 14430 8027
rect 14464 7993 14510 8027
rect 14544 7993 14590 8027
rect 14624 7993 14650 8027
rect 14318 7975 14650 7993
rect 14928 8027 15260 8043
rect 14928 7993 14954 8027
rect 14988 7993 15034 8027
rect 15068 7993 15114 8027
rect 15148 7993 15194 8027
rect 15228 7993 15260 8027
rect 14928 7975 15260 7993
rect 15530 8027 15862 8043
rect 15530 7993 15562 8027
rect 15596 7993 15642 8027
rect 15676 7993 15722 8027
rect 15756 7993 15802 8027
rect 15836 7993 15862 8027
rect 15530 7975 15862 7993
rect 16266 8027 16598 8043
rect 16266 7993 16292 8027
rect 16326 7993 16372 8027
rect 16406 7993 16452 8027
rect 16486 7993 16532 8027
rect 16566 7993 16598 8027
rect 16266 7975 16598 7993
rect 16868 8027 17200 8043
rect 16868 7993 16900 8027
rect 16934 7993 16980 8027
rect 17014 7993 17060 8027
rect 17094 7993 17140 8027
rect 17174 7993 17200 8027
rect 16868 7975 17200 7993
rect 17602 8027 17934 8043
rect 17602 7993 17634 8027
rect 17668 7993 17714 8027
rect 17748 7993 17794 8027
rect 17828 7993 17874 8027
rect 17908 7993 17934 8027
rect 17602 7975 17934 7993
rect 13370 7547 13399 7615
rect 13433 7547 13491 7615
rect 13525 7547 13583 7615
rect 13617 7547 13675 7615
rect 13709 7547 13767 7615
rect 13801 7547 13859 7615
rect 13893 7547 13951 7615
rect 13985 7547 14043 7615
rect 14077 7547 14135 7615
rect 14169 7581 14226 7615
rect 14260 7581 14319 7615
rect 14169 7547 14227 7581
rect 14261 7547 14319 7581
rect 14353 7547 14411 7615
rect 14445 7547 14503 7615
rect 14537 7547 14595 7615
rect 14629 7547 14687 7615
rect 14721 7547 14779 7615
rect 14813 7547 14871 7615
rect 14905 7547 14963 7615
rect 14997 7547 15055 7615
rect 15089 7547 15147 7615
rect 15181 7547 15239 7615
rect 15273 7547 15331 7615
rect 15365 7547 15423 7615
rect 15457 7547 15515 7615
rect 15549 7547 15607 7615
rect 15641 7547 15699 7615
rect 15733 7547 15791 7615
rect 15825 7547 15883 7615
rect 15917 7547 15975 7615
rect 16009 7547 16067 7615
rect 16101 7547 16159 7615
rect 16193 7547 16251 7615
rect 16285 7547 16343 7615
rect 16377 7547 16435 7615
rect 16469 7547 16527 7615
rect 16561 7547 16619 7615
rect 16653 7547 16711 7615
rect 16745 7547 16803 7615
rect 16837 7547 16895 7615
rect 16929 7547 16987 7615
rect 17021 7547 17079 7615
rect 17113 7547 17171 7615
rect 17205 7547 17263 7615
rect 17297 7547 17355 7615
rect 17389 7547 17447 7615
rect 17481 7547 17539 7615
rect 17573 7547 17631 7615
rect 17665 7547 17723 7615
rect 17757 7547 17815 7615
rect 17849 7547 17907 7615
rect 17941 7547 17999 7615
rect 18033 7547 18091 7615
rect 18125 7547 18154 7615
rect 13473 7505 13539 7547
rect 13387 7479 13439 7495
rect 13387 7445 13405 7479
rect 13473 7471 13489 7505
rect 13523 7471 13539 7505
rect 13657 7505 13727 7547
rect 13573 7479 13618 7495
rect 13387 7437 13439 7445
rect 13607 7445 13618 7479
rect 13657 7471 13677 7505
rect 13711 7471 13727 7505
rect 13851 7505 14050 7511
rect 13761 7487 13795 7503
rect 13387 7403 13538 7437
rect 13387 7355 13458 7369
rect 13387 7334 13416 7355
rect 13387 7300 13402 7334
rect 13450 7321 13458 7355
rect 13436 7300 13458 7321
rect 13387 7239 13458 7300
rect 13492 7334 13538 7403
rect 13492 7300 13504 7334
rect 13492 7207 13538 7300
rect 13387 7189 13492 7205
rect 13387 7155 13405 7189
rect 13439 7173 13492 7189
rect 13526 7173 13538 7207
rect 13439 7171 13538 7173
rect 13573 7411 13618 7445
rect 13851 7471 13867 7505
rect 13901 7471 14050 7505
rect 13761 7437 13795 7453
rect 13573 7377 13584 7411
rect 13573 7189 13618 7377
rect 13387 7121 13439 7155
rect 13607 7155 13618 7189
rect 13652 7399 13795 7437
rect 13836 7407 13880 7423
rect 13652 7205 13686 7399
rect 13870 7373 13880 7407
rect 13720 7347 13802 7363
rect 13754 7313 13802 7347
rect 13720 7281 13802 7313
rect 13720 7247 13736 7281
rect 13770 7247 13802 7281
rect 13720 7239 13802 7247
rect 13836 7249 13880 7373
rect 13916 7411 13982 7435
rect 13916 7395 13948 7411
rect 13916 7361 13932 7395
rect 13966 7361 13982 7377
rect 14016 7325 14050 7471
rect 14084 7509 14118 7547
rect 14084 7459 14118 7475
rect 14152 7489 14386 7513
rect 14152 7455 14168 7489
rect 14202 7479 14386 7489
rect 14202 7455 14218 7479
rect 14352 7471 14386 7479
rect 14440 7505 14506 7547
rect 14440 7471 14456 7505
rect 14490 7471 14506 7505
rect 14634 7505 14787 7511
rect 14634 7471 14650 7505
rect 14684 7471 14787 7505
rect 14088 7411 14170 7417
rect 14252 7411 14268 7445
rect 14302 7411 14318 7445
rect 14352 7421 14386 7437
rect 14088 7385 14136 7411
rect 14088 7351 14104 7385
rect 14138 7371 14170 7377
rect 14274 7385 14318 7411
rect 14595 7407 14652 7423
rect 14138 7351 14154 7371
rect 14274 7351 14536 7385
rect 13970 7317 14050 7325
rect 14196 7317 14240 7333
rect 13970 7283 14206 7317
rect 13836 7233 13936 7249
rect 13836 7207 13902 7233
rect 13652 7171 13795 7205
rect 13836 7173 13860 7207
rect 13894 7199 13902 7207
rect 13894 7173 13936 7199
rect 13387 7087 13405 7121
rect 13387 7071 13439 7087
rect 13473 7103 13489 7137
rect 13523 7103 13539 7137
rect 13473 7037 13539 7103
rect 13573 7121 13618 7155
rect 13607 7087 13618 7121
rect 13573 7071 13618 7087
rect 13657 7103 13677 7137
rect 13711 7103 13727 7137
rect 13657 7037 13727 7103
rect 13761 7121 13795 7171
rect 13970 7114 14004 7283
rect 14190 7267 14240 7283
rect 14038 7233 14088 7249
rect 14072 7207 14088 7233
rect 14274 7207 14308 7351
rect 14470 7317 14486 7351
rect 14520 7317 14536 7351
rect 14595 7373 14618 7407
rect 14595 7343 14652 7373
rect 14342 7283 14358 7317
rect 14392 7283 14408 7317
rect 14595 7309 14596 7343
rect 14630 7339 14652 7343
rect 14630 7309 14719 7339
rect 14595 7303 14719 7309
rect 14342 7281 14408 7283
rect 14342 7275 14543 7281
rect 14342 7241 14504 7275
rect 14538 7241 14543 7275
rect 14342 7233 14543 7241
rect 14583 7233 14630 7249
rect 14072 7199 14188 7207
rect 14038 7173 14188 7199
rect 14222 7173 14308 7207
rect 14617 7207 14630 7233
rect 14038 7157 14308 7173
rect 14188 7139 14222 7157
rect 13761 7071 13795 7087
rect 13838 7080 13854 7114
rect 13888 7080 14004 7114
rect 14052 7089 14068 7123
rect 14102 7089 14128 7123
rect 14188 7089 14222 7105
rect 14346 7147 14362 7181
rect 14396 7147 14412 7181
rect 14583 7173 14596 7199
rect 14678 7233 14719 7303
rect 14678 7199 14685 7233
rect 14678 7183 14719 7199
rect 14753 7317 14787 7471
rect 14823 7509 14875 7547
rect 14823 7475 14841 7509
rect 14823 7459 14875 7475
rect 14927 7497 15161 7513
rect 14927 7489 15127 7497
rect 14927 7455 14943 7489
rect 14977 7479 15127 7489
rect 14977 7455 14993 7479
rect 15127 7447 15161 7463
rect 15218 7495 15265 7511
rect 15218 7461 15231 7495
rect 14862 7411 14937 7417
rect 14862 7377 14872 7411
rect 14906 7385 14937 7411
rect 15027 7411 15043 7445
rect 15077 7411 15093 7445
rect 15218 7413 15265 7461
rect 15027 7408 15093 7411
rect 14862 7351 14881 7377
rect 14915 7351 14937 7385
rect 14979 7333 15023 7349
rect 14979 7317 14989 7333
rect 14753 7299 14989 7317
rect 14753 7283 15023 7299
rect 14583 7167 14630 7173
rect 14346 7113 14412 7147
rect 14753 7114 14787 7283
rect 14821 7233 14871 7249
rect 14855 7199 14871 7233
rect 14821 7181 14871 7199
rect 15057 7181 15093 7408
rect 15127 7379 15265 7413
rect 15310 7505 15376 7547
rect 15310 7471 15326 7505
rect 15360 7471 15376 7505
rect 15310 7403 15376 7471
rect 15410 7471 15467 7513
rect 15444 7437 15467 7471
rect 15410 7421 15467 7437
rect 15127 7317 15182 7379
rect 15342 7349 15392 7365
rect 15161 7283 15182 7317
rect 15233 7340 15258 7345
rect 15233 7306 15255 7340
rect 15292 7311 15308 7345
rect 15289 7306 15308 7311
rect 15233 7299 15308 7306
rect 15342 7315 15358 7349
rect 15342 7299 15392 7315
rect 15127 7275 15182 7283
rect 15127 7241 15148 7275
rect 15182 7241 15229 7249
rect 15127 7215 15229 7241
rect 15263 7215 15279 7249
rect 15342 7181 15376 7299
rect 15426 7238 15467 7421
rect 14821 7147 15376 7181
rect 15410 7218 15467 7238
rect 15444 7184 15467 7218
rect 15410 7150 15467 7184
rect 14052 7037 14128 7089
rect 14346 7079 14362 7113
rect 14396 7079 14412 7113
rect 14621 7080 14637 7114
rect 14671 7080 14787 7114
rect 14959 7139 14993 7147
rect 14346 7037 14412 7079
rect 14835 7079 14851 7113
rect 14885 7079 14911 7113
rect 15444 7116 15467 7150
rect 14959 7089 14993 7105
rect 14835 7037 14911 7079
rect 15099 7079 15115 7113
rect 15149 7079 15326 7113
rect 15360 7079 15376 7113
rect 15099 7037 15376 7079
rect 15410 7071 15467 7116
rect 15501 7479 15564 7513
rect 15501 7445 15514 7479
rect 15548 7445 15564 7479
rect 15600 7505 15659 7547
rect 15600 7471 15609 7505
rect 15643 7471 15659 7505
rect 15600 7455 15659 7471
rect 15693 7469 15745 7513
rect 15865 7505 15931 7547
rect 15501 7365 15564 7445
rect 15727 7435 15745 7469
rect 15693 7399 15745 7435
rect 15779 7479 15831 7495
rect 15779 7445 15797 7479
rect 15865 7471 15881 7505
rect 15915 7471 15931 7505
rect 16049 7505 16119 7547
rect 15965 7479 16010 7495
rect 15779 7437 15831 7445
rect 15999 7445 16010 7479
rect 16049 7471 16069 7505
rect 16103 7471 16119 7505
rect 16243 7505 16442 7511
rect 16153 7487 16187 7503
rect 15779 7403 15930 7437
rect 15501 7349 15668 7365
rect 15501 7315 15634 7349
rect 15501 7299 15668 7315
rect 15501 7199 15564 7299
rect 15702 7275 15745 7399
rect 15693 7217 15745 7275
rect 15779 7334 15850 7369
rect 15779 7300 15794 7334
rect 15828 7310 15850 7334
rect 15779 7276 15805 7300
rect 15839 7276 15850 7310
rect 15779 7239 15850 7276
rect 15884 7334 15930 7403
rect 15884 7300 15896 7334
rect 15501 7165 15514 7199
rect 15548 7165 15564 7199
rect 15501 7131 15564 7165
rect 15501 7097 15514 7131
rect 15548 7097 15564 7131
rect 15501 7081 15564 7097
rect 15600 7193 15659 7211
rect 15600 7159 15609 7193
rect 15643 7159 15659 7193
rect 15600 7125 15659 7159
rect 15600 7091 15609 7125
rect 15643 7091 15659 7125
rect 15600 7037 15659 7091
rect 15727 7183 15745 7217
rect 15884 7207 15930 7300
rect 15693 7149 15745 7183
rect 15727 7143 15745 7149
rect 15693 7109 15703 7115
rect 15737 7109 15745 7143
rect 15693 7071 15745 7109
rect 15779 7189 15884 7205
rect 15779 7155 15797 7189
rect 15831 7173 15884 7189
rect 15918 7173 15930 7207
rect 15831 7171 15930 7173
rect 15965 7411 16010 7445
rect 16243 7471 16259 7505
rect 16293 7471 16442 7505
rect 16153 7437 16187 7453
rect 15965 7377 15976 7411
rect 15965 7189 16010 7377
rect 15779 7121 15831 7155
rect 15999 7155 16010 7189
rect 16044 7399 16187 7437
rect 16228 7407 16272 7423
rect 16044 7205 16078 7399
rect 16262 7373 16272 7407
rect 16112 7347 16194 7363
rect 16146 7343 16194 7347
rect 16112 7309 16138 7313
rect 16172 7309 16194 7343
rect 16112 7239 16194 7309
rect 16228 7249 16272 7373
rect 16308 7411 16374 7435
rect 16308 7395 16340 7411
rect 16308 7361 16324 7395
rect 16358 7361 16374 7377
rect 16408 7325 16442 7471
rect 16476 7509 16510 7547
rect 16476 7459 16510 7475
rect 16544 7489 16778 7513
rect 16544 7455 16560 7489
rect 16594 7479 16778 7489
rect 16594 7455 16610 7479
rect 16744 7471 16778 7479
rect 16832 7505 16898 7547
rect 16832 7471 16848 7505
rect 16882 7471 16898 7505
rect 17026 7505 17179 7511
rect 17026 7471 17042 7505
rect 17076 7471 17179 7505
rect 16480 7411 16562 7417
rect 16644 7411 16660 7445
rect 16694 7411 16710 7445
rect 16744 7421 16778 7437
rect 16480 7385 16528 7411
rect 16480 7351 16496 7385
rect 16530 7371 16562 7377
rect 16666 7385 16710 7411
rect 16987 7407 17044 7423
rect 16530 7351 16546 7371
rect 16666 7351 16928 7385
rect 16362 7317 16442 7325
rect 16588 7317 16632 7333
rect 16362 7283 16598 7317
rect 16228 7233 16328 7249
rect 16228 7207 16294 7233
rect 16044 7171 16187 7205
rect 16228 7173 16252 7207
rect 16286 7199 16294 7207
rect 16286 7173 16328 7199
rect 15779 7087 15797 7121
rect 15779 7071 15831 7087
rect 15865 7103 15881 7137
rect 15915 7103 15931 7137
rect 15865 7037 15931 7103
rect 15965 7121 16010 7155
rect 15999 7087 16010 7121
rect 15965 7071 16010 7087
rect 16049 7103 16069 7137
rect 16103 7103 16119 7137
rect 16049 7037 16119 7103
rect 16153 7121 16187 7171
rect 16362 7114 16396 7283
rect 16582 7267 16632 7283
rect 16430 7233 16480 7249
rect 16464 7207 16480 7233
rect 16666 7207 16700 7351
rect 16862 7317 16878 7351
rect 16912 7317 16928 7351
rect 16987 7373 17010 7407
rect 16987 7343 17044 7373
rect 16734 7283 16750 7317
rect 16784 7283 16800 7317
rect 16987 7309 16988 7343
rect 17022 7339 17044 7343
rect 17022 7309 17111 7339
rect 16987 7303 17111 7309
rect 16734 7281 16800 7283
rect 16734 7275 16935 7281
rect 16734 7241 16896 7275
rect 16930 7241 16935 7275
rect 16734 7233 16935 7241
rect 16975 7233 17022 7249
rect 16464 7199 16580 7207
rect 16430 7173 16580 7199
rect 16614 7173 16700 7207
rect 17009 7207 17022 7233
rect 16430 7157 16700 7173
rect 16580 7139 16614 7157
rect 16153 7071 16187 7087
rect 16230 7080 16246 7114
rect 16280 7080 16396 7114
rect 16444 7089 16460 7123
rect 16494 7089 16520 7123
rect 16580 7089 16614 7105
rect 16738 7147 16754 7181
rect 16788 7147 16804 7181
rect 16975 7173 16988 7199
rect 17070 7233 17111 7303
rect 17070 7199 17077 7233
rect 17070 7183 17111 7199
rect 17145 7317 17179 7471
rect 17215 7509 17267 7547
rect 17215 7475 17233 7509
rect 17215 7459 17267 7475
rect 17319 7497 17553 7513
rect 17319 7489 17519 7497
rect 17319 7455 17335 7489
rect 17369 7479 17519 7489
rect 17369 7455 17385 7479
rect 17519 7447 17553 7463
rect 17610 7495 17657 7511
rect 17610 7461 17623 7495
rect 17254 7411 17329 7417
rect 17254 7377 17264 7411
rect 17298 7385 17329 7411
rect 17419 7411 17435 7445
rect 17469 7411 17485 7445
rect 17610 7413 17657 7461
rect 17419 7408 17485 7411
rect 17254 7351 17273 7377
rect 17307 7351 17329 7385
rect 17371 7333 17415 7349
rect 17371 7317 17381 7333
rect 17145 7299 17381 7317
rect 17145 7283 17415 7299
rect 16975 7167 17022 7173
rect 16738 7113 16804 7147
rect 17145 7114 17179 7283
rect 17213 7233 17263 7249
rect 17247 7199 17263 7233
rect 17213 7181 17263 7199
rect 17449 7181 17485 7408
rect 17519 7379 17657 7413
rect 17702 7505 17768 7547
rect 17702 7471 17718 7505
rect 17752 7471 17768 7505
rect 17702 7403 17768 7471
rect 17802 7471 17859 7513
rect 17836 7437 17859 7471
rect 17802 7421 17859 7437
rect 17519 7317 17574 7379
rect 17734 7349 17784 7365
rect 17553 7283 17574 7317
rect 17625 7311 17650 7345
rect 17684 7344 17700 7345
rect 17625 7310 17654 7311
rect 17688 7310 17700 7344
rect 17625 7299 17700 7310
rect 17734 7315 17750 7349
rect 17734 7299 17784 7315
rect 17519 7275 17574 7283
rect 17519 7241 17540 7275
rect 17574 7241 17621 7249
rect 17519 7215 17621 7241
rect 17655 7215 17671 7249
rect 17734 7181 17768 7299
rect 17818 7238 17859 7421
rect 17213 7147 17768 7181
rect 17802 7218 17859 7238
rect 17836 7184 17859 7218
rect 17802 7150 17859 7184
rect 16444 7037 16520 7089
rect 16738 7079 16754 7113
rect 16788 7079 16804 7113
rect 17013 7080 17029 7114
rect 17063 7080 17179 7114
rect 17351 7139 17385 7147
rect 16738 7037 16804 7079
rect 17227 7079 17243 7113
rect 17277 7079 17303 7113
rect 17836 7116 17859 7150
rect 17351 7089 17385 7105
rect 17227 7037 17303 7079
rect 17491 7079 17507 7113
rect 17541 7079 17718 7113
rect 17752 7079 17768 7113
rect 17491 7037 17768 7079
rect 17802 7071 17859 7116
rect 17893 7479 17956 7513
rect 17893 7445 17906 7479
rect 17940 7445 17956 7479
rect 17992 7505 18051 7547
rect 17992 7471 18001 7505
rect 18035 7471 18051 7505
rect 17992 7455 18051 7471
rect 18085 7469 18137 7513
rect 18119 7460 18137 7469
rect 17893 7365 17956 7445
rect 18085 7426 18091 7435
rect 18125 7426 18137 7460
rect 18085 7399 18137 7426
rect 17893 7349 18060 7365
rect 17893 7315 18026 7349
rect 17893 7299 18060 7315
rect 17893 7199 17956 7299
rect 18094 7275 18137 7399
rect 18085 7217 18137 7275
rect 17893 7165 17906 7199
rect 17940 7165 17956 7199
rect 17893 7131 17956 7165
rect 17893 7097 17906 7131
rect 17940 7097 17956 7131
rect 17893 7081 17956 7097
rect 17992 7193 18051 7211
rect 17992 7159 18001 7193
rect 18035 7159 18051 7193
rect 17992 7125 18051 7159
rect 17992 7091 18001 7125
rect 18035 7091 18051 7125
rect 17992 7037 18051 7091
rect 18119 7183 18137 7217
rect 18085 7149 18137 7183
rect 18119 7115 18137 7149
rect 18085 7071 18137 7115
rect 13370 7003 13399 7037
rect 13433 7003 13491 7037
rect 13525 7003 13583 7037
rect 13617 7003 13675 7037
rect 13709 7003 13767 7037
rect 13801 7003 13859 7037
rect 13893 7003 13951 7037
rect 13985 7003 14043 7037
rect 14077 7003 14135 7037
rect 14169 7003 14227 7037
rect 14261 7003 14319 7037
rect 14353 7003 14411 7037
rect 14445 7003 14503 7037
rect 14537 7003 14595 7037
rect 14629 7003 14687 7037
rect 14721 7003 14779 7037
rect 14813 7003 14871 7037
rect 14905 7003 14963 7037
rect 14997 7003 15055 7037
rect 15089 7003 15147 7037
rect 15181 7003 15239 7037
rect 15273 7003 15331 7037
rect 15365 7003 15423 7037
rect 15457 7003 15515 7037
rect 15549 7003 15607 7037
rect 15641 7003 15699 7037
rect 15733 7003 15791 7037
rect 15825 7003 15883 7037
rect 15917 7003 15975 7037
rect 16009 7003 16067 7037
rect 16101 7003 16159 7037
rect 16193 7003 16251 7037
rect 16285 7003 16343 7037
rect 16377 7003 16435 7037
rect 16469 7003 16527 7037
rect 16561 7003 16619 7037
rect 16653 7003 16711 7037
rect 16745 7003 16803 7037
rect 16837 7003 16895 7037
rect 16929 7003 16987 7037
rect 17021 7003 17079 7037
rect 17113 7003 17171 7037
rect 17205 7003 17263 7037
rect 17297 7003 17355 7037
rect 17389 7003 17447 7037
rect 17481 7003 17539 7037
rect 17573 7003 17631 7037
rect 17665 7003 17723 7037
rect 17757 7003 17815 7037
rect 17849 7003 17907 7037
rect 17941 7003 17999 7037
rect 18033 7003 18091 7037
rect 18125 7003 18154 7037
rect 13370 6989 18154 7003
rect 13370 6955 13400 6989
rect 13434 6955 13491 6989
rect 13525 6955 13584 6989
rect 13618 6955 13675 6989
rect 13709 6955 13766 6989
rect 13800 6955 13860 6989
rect 13894 6955 13951 6989
rect 13985 6955 14044 6989
rect 14078 6955 14135 6989
rect 14169 6955 14227 6989
rect 14261 6955 14318 6989
rect 14352 6955 14411 6989
rect 14445 6955 14504 6989
rect 14538 6955 14595 6989
rect 14629 6955 14687 6989
rect 14721 6955 14779 6989
rect 14813 6955 14871 6989
rect 14905 6955 14963 6989
rect 14997 6955 15055 6989
rect 15089 6955 15147 6989
rect 15181 6955 15240 6989
rect 15274 6955 15330 6989
rect 15364 6955 15423 6989
rect 15457 6955 15516 6989
rect 15550 6955 15608 6989
rect 15642 6955 15699 6989
rect 15733 6955 15792 6989
rect 15826 6955 15884 6989
rect 15918 6955 15976 6989
rect 16010 6955 16068 6989
rect 16102 6955 16160 6989
rect 16194 6955 16252 6989
rect 16286 6955 16343 6989
rect 16377 6955 16434 6989
rect 16468 6955 16527 6989
rect 16561 6955 16620 6989
rect 16654 6955 16712 6989
rect 16746 6955 16803 6989
rect 16837 6955 16897 6989
rect 16931 6955 16987 6989
rect 17021 6955 17078 6989
rect 17112 6955 17171 6989
rect 17205 6955 17264 6989
rect 17298 6955 17356 6989
rect 17390 6955 17447 6989
rect 17481 6955 17539 6989
rect 17573 6955 17631 6989
rect 17665 6955 17722 6989
rect 17756 6955 17814 6989
rect 17848 6955 17907 6989
rect 17941 6955 17999 6989
rect 18033 6955 18091 6989
rect 18125 6955 18154 6989
rect 13370 6941 18154 6955
rect 13370 6907 13399 6941
rect 13433 6907 13491 6941
rect 13525 6907 13583 6941
rect 13617 6907 13675 6941
rect 13709 6907 13767 6941
rect 13801 6907 13859 6941
rect 13893 6907 13951 6941
rect 13985 6907 14043 6941
rect 14077 6907 14135 6941
rect 14169 6907 14227 6941
rect 14261 6907 14319 6941
rect 14353 6907 14411 6941
rect 14445 6907 14503 6941
rect 14537 6907 14595 6941
rect 14629 6907 14687 6941
rect 14721 6907 14779 6941
rect 14813 6907 14871 6941
rect 14905 6907 14963 6941
rect 14997 6907 15055 6941
rect 15089 6907 15147 6941
rect 15181 6907 15239 6941
rect 15273 6907 15331 6941
rect 15365 6907 15423 6941
rect 15457 6907 15515 6941
rect 15549 6907 15607 6941
rect 15641 6907 15699 6941
rect 15733 6907 15791 6941
rect 15825 6907 15883 6941
rect 15917 6907 15975 6941
rect 16009 6907 16067 6941
rect 16101 6907 16159 6941
rect 16193 6907 16251 6941
rect 16285 6907 16343 6941
rect 16377 6907 16435 6941
rect 16469 6907 16527 6941
rect 16561 6907 16619 6941
rect 16653 6907 16711 6941
rect 16745 6907 16803 6941
rect 16837 6907 16895 6941
rect 16929 6907 16987 6941
rect 17021 6907 17079 6941
rect 17113 6907 17171 6941
rect 17205 6907 17263 6941
rect 17297 6907 17355 6941
rect 17389 6907 17447 6941
rect 17481 6907 17539 6941
rect 17573 6907 17631 6941
rect 17665 6907 17723 6941
rect 17757 6907 17815 6941
rect 17849 6907 17907 6941
rect 17941 6907 17999 6941
rect 18033 6907 18091 6941
rect 18125 6907 18154 6941
rect 13387 6857 13439 6873
rect 13387 6823 13405 6857
rect 13387 6789 13439 6823
rect 13473 6841 13539 6907
rect 13473 6807 13489 6841
rect 13523 6807 13539 6841
rect 13573 6857 13618 6873
rect 13607 6823 13618 6857
rect 13387 6755 13405 6789
rect 13573 6789 13618 6823
rect 13657 6841 13727 6907
rect 13657 6807 13677 6841
rect 13711 6807 13727 6841
rect 13761 6857 13795 6873
rect 13838 6830 13854 6864
rect 13888 6830 14004 6864
rect 13439 6771 13538 6773
rect 13439 6755 13492 6771
rect 13387 6739 13492 6755
rect 13526 6737 13538 6771
rect 13387 6671 13411 6705
rect 13445 6671 13458 6705
rect 13387 6644 13458 6671
rect 13387 6610 13402 6644
rect 13436 6610 13458 6644
rect 13387 6575 13458 6610
rect 13492 6644 13538 6737
rect 13492 6610 13504 6644
rect 13492 6541 13538 6610
rect 13387 6507 13538 6541
rect 13607 6755 13618 6789
rect 13761 6773 13795 6823
rect 13573 6567 13618 6755
rect 13573 6533 13584 6567
rect 13387 6499 13439 6507
rect 13387 6465 13405 6499
rect 13573 6499 13618 6533
rect 13652 6739 13795 6773
rect 13652 6545 13686 6739
rect 13836 6737 13860 6771
rect 13894 6745 13936 6771
rect 13894 6737 13902 6745
rect 13836 6711 13902 6737
rect 13720 6635 13802 6705
rect 13720 6631 13741 6635
rect 13775 6601 13802 6635
rect 13754 6597 13802 6601
rect 13720 6581 13802 6597
rect 13836 6695 13936 6711
rect 13836 6571 13880 6695
rect 13970 6661 14004 6830
rect 14052 6855 14128 6907
rect 14346 6865 14412 6907
rect 14052 6821 14068 6855
rect 14102 6821 14128 6855
rect 14188 6839 14222 6855
rect 14188 6787 14222 6805
rect 14346 6831 14362 6865
rect 14396 6831 14412 6865
rect 14835 6865 14911 6907
rect 14346 6797 14412 6831
rect 14621 6830 14637 6864
rect 14671 6830 14787 6864
rect 14835 6831 14851 6865
rect 14885 6831 14911 6865
rect 15099 6865 15376 6907
rect 14959 6839 14993 6855
rect 14038 6771 14308 6787
rect 14038 6745 14188 6771
rect 14072 6737 14188 6745
rect 14222 6737 14308 6771
rect 14346 6763 14362 6797
rect 14396 6763 14412 6797
rect 14583 6771 14630 6777
rect 14072 6711 14088 6737
rect 14038 6695 14088 6711
rect 14190 6661 14240 6677
rect 13970 6627 14206 6661
rect 13970 6619 14050 6627
rect 13652 6507 13795 6545
rect 13870 6537 13880 6571
rect 13836 6521 13880 6537
rect 13916 6549 13932 6583
rect 13966 6567 13982 6583
rect 13916 6533 13948 6549
rect 13916 6509 13982 6533
rect 13387 6449 13439 6465
rect 13473 6439 13489 6473
rect 13523 6439 13539 6473
rect 13607 6465 13618 6499
rect 13761 6491 13795 6507
rect 13573 6449 13618 6465
rect 13473 6397 13539 6439
rect 13657 6439 13677 6473
rect 13711 6439 13727 6473
rect 14016 6473 14050 6619
rect 14196 6611 14240 6627
rect 14274 6593 14308 6737
rect 14583 6745 14596 6771
rect 14617 6711 14630 6737
rect 14342 6703 14543 6711
rect 14342 6669 14504 6703
rect 14538 6669 14543 6703
rect 14583 6695 14630 6711
rect 14678 6745 14719 6761
rect 14678 6711 14685 6745
rect 14342 6663 14543 6669
rect 14342 6661 14408 6663
rect 14342 6627 14358 6661
rect 14392 6627 14408 6661
rect 14678 6641 14719 6711
rect 14595 6635 14719 6641
rect 14470 6593 14486 6627
rect 14520 6593 14536 6627
rect 14088 6559 14104 6593
rect 14138 6573 14154 6593
rect 14138 6567 14170 6573
rect 14088 6533 14136 6559
rect 14274 6559 14536 6593
rect 14595 6601 14596 6635
rect 14630 6605 14719 6635
rect 14753 6661 14787 6830
rect 15099 6831 15115 6865
rect 15149 6831 15326 6865
rect 15360 6831 15376 6865
rect 14959 6797 14993 6805
rect 15410 6828 15467 6873
rect 14821 6763 15376 6797
rect 14821 6745 14871 6763
rect 14855 6711 14871 6745
rect 14821 6695 14871 6711
rect 14753 6645 15023 6661
rect 14753 6627 14989 6645
rect 14630 6601 14652 6605
rect 14595 6571 14652 6601
rect 14274 6533 14318 6559
rect 14088 6527 14170 6533
rect 14252 6499 14268 6533
rect 14302 6499 14318 6533
rect 14595 6537 14618 6571
rect 14352 6507 14386 6523
rect 14595 6521 14652 6537
rect 13761 6441 13795 6457
rect 13657 6397 13727 6439
rect 13851 6439 13867 6473
rect 13901 6439 14050 6473
rect 13851 6433 14050 6439
rect 14084 6469 14118 6485
rect 14084 6397 14118 6435
rect 14152 6455 14168 6489
rect 14202 6465 14218 6489
rect 14753 6473 14787 6627
rect 14979 6611 14989 6627
rect 14979 6595 15023 6611
rect 14862 6567 14881 6593
rect 14862 6533 14872 6567
rect 14915 6559 14937 6593
rect 14906 6533 14937 6559
rect 15057 6536 15093 6763
rect 14862 6527 14937 6533
rect 15027 6533 15093 6536
rect 15027 6499 15043 6533
rect 15077 6499 15093 6533
rect 15127 6703 15229 6729
rect 15127 6669 15148 6703
rect 15182 6695 15229 6703
rect 15263 6695 15279 6729
rect 15127 6661 15182 6669
rect 15161 6627 15182 6661
rect 15342 6645 15376 6763
rect 15444 6794 15467 6828
rect 15410 6760 15467 6794
rect 15444 6726 15467 6760
rect 15410 6706 15467 6726
rect 15127 6565 15182 6627
rect 15233 6633 15308 6645
rect 15233 6599 15256 6633
rect 15292 6599 15308 6633
rect 15342 6629 15392 6645
rect 15342 6595 15358 6629
rect 15342 6579 15392 6595
rect 15127 6531 15265 6565
rect 14352 6465 14386 6473
rect 14202 6455 14386 6465
rect 14152 6431 14386 6455
rect 14440 6439 14456 6473
rect 14490 6439 14506 6473
rect 14440 6397 14506 6439
rect 14634 6439 14650 6473
rect 14684 6439 14787 6473
rect 14634 6433 14787 6439
rect 14823 6469 14875 6485
rect 14823 6435 14841 6469
rect 14823 6397 14875 6435
rect 14927 6455 14943 6489
rect 14977 6465 14993 6489
rect 15127 6481 15161 6497
rect 14977 6455 15127 6465
rect 14927 6447 15127 6455
rect 14927 6431 15161 6447
rect 15218 6483 15265 6531
rect 15218 6449 15231 6483
rect 15218 6433 15265 6449
rect 15310 6473 15376 6541
rect 15426 6523 15467 6706
rect 15310 6439 15326 6473
rect 15360 6439 15376 6473
rect 15310 6397 15376 6439
rect 15410 6507 15467 6523
rect 15444 6473 15467 6507
rect 15410 6431 15467 6473
rect 15501 6847 15564 6863
rect 15501 6813 15514 6847
rect 15548 6813 15564 6847
rect 15501 6779 15564 6813
rect 15501 6745 15514 6779
rect 15548 6745 15564 6779
rect 15501 6645 15564 6745
rect 15600 6853 15659 6907
rect 15600 6819 15609 6853
rect 15643 6819 15659 6853
rect 15600 6785 15659 6819
rect 15600 6751 15609 6785
rect 15643 6751 15659 6785
rect 15600 6733 15659 6751
rect 15693 6831 15745 6873
rect 15693 6829 15702 6831
rect 15736 6797 15745 6831
rect 15727 6795 15745 6797
rect 15693 6761 15745 6795
rect 15727 6727 15745 6761
rect 15779 6857 15831 6873
rect 15779 6823 15797 6857
rect 15779 6789 15831 6823
rect 15865 6841 15931 6907
rect 15865 6807 15881 6841
rect 15915 6807 15931 6841
rect 15965 6857 16010 6873
rect 15999 6823 16010 6857
rect 15779 6755 15797 6789
rect 15965 6789 16010 6823
rect 16049 6841 16119 6907
rect 16049 6807 16069 6841
rect 16103 6807 16119 6841
rect 16153 6857 16187 6873
rect 16230 6830 16246 6864
rect 16280 6830 16396 6864
rect 15831 6771 15930 6773
rect 15831 6755 15884 6771
rect 15779 6739 15884 6755
rect 15693 6669 15745 6727
rect 15918 6737 15930 6771
rect 15501 6629 15668 6645
rect 15501 6595 15634 6629
rect 15501 6579 15668 6595
rect 15501 6499 15564 6579
rect 15702 6545 15745 6669
rect 15779 6662 15850 6705
rect 15779 6644 15806 6662
rect 15779 6610 15794 6644
rect 15840 6628 15850 6662
rect 15828 6610 15850 6628
rect 15779 6575 15850 6610
rect 15884 6644 15930 6737
rect 15884 6610 15896 6644
rect 15501 6465 15514 6499
rect 15548 6465 15564 6499
rect 15693 6509 15745 6545
rect 15884 6541 15930 6610
rect 15501 6431 15564 6465
rect 15600 6473 15659 6489
rect 15600 6439 15609 6473
rect 15643 6439 15659 6473
rect 15600 6397 15659 6439
rect 15727 6475 15745 6509
rect 15693 6431 15745 6475
rect 15779 6507 15930 6541
rect 15999 6755 16010 6789
rect 16153 6773 16187 6823
rect 15965 6567 16010 6755
rect 15965 6533 15976 6567
rect 15779 6499 15831 6507
rect 15779 6465 15797 6499
rect 15965 6499 16010 6533
rect 16044 6739 16187 6773
rect 16044 6545 16078 6739
rect 16228 6737 16252 6771
rect 16286 6745 16328 6771
rect 16286 6737 16294 6745
rect 16228 6711 16294 6737
rect 16112 6634 16194 6705
rect 16112 6631 16139 6634
rect 16173 6600 16194 6634
rect 16146 6597 16194 6600
rect 16112 6581 16194 6597
rect 16228 6695 16328 6711
rect 16228 6571 16272 6695
rect 16362 6661 16396 6830
rect 16444 6855 16520 6907
rect 16738 6865 16804 6907
rect 16444 6821 16460 6855
rect 16494 6821 16520 6855
rect 16580 6839 16614 6855
rect 16580 6787 16614 6805
rect 16738 6831 16754 6865
rect 16788 6831 16804 6865
rect 17227 6865 17303 6907
rect 16738 6797 16804 6831
rect 17013 6830 17029 6864
rect 17063 6830 17179 6864
rect 17227 6831 17243 6865
rect 17277 6831 17303 6865
rect 17491 6865 17768 6907
rect 17351 6839 17385 6855
rect 16430 6771 16700 6787
rect 16430 6745 16580 6771
rect 16464 6737 16580 6745
rect 16614 6737 16700 6771
rect 16738 6763 16754 6797
rect 16788 6763 16804 6797
rect 16975 6771 17022 6777
rect 16464 6711 16480 6737
rect 16430 6695 16480 6711
rect 16582 6661 16632 6677
rect 16362 6627 16598 6661
rect 16362 6619 16442 6627
rect 16044 6507 16187 6545
rect 16262 6537 16272 6571
rect 16228 6521 16272 6537
rect 16308 6549 16324 6583
rect 16358 6567 16374 6583
rect 16308 6533 16340 6549
rect 16308 6509 16374 6533
rect 15779 6449 15831 6465
rect 15865 6439 15881 6473
rect 15915 6439 15931 6473
rect 15999 6465 16010 6499
rect 16153 6491 16187 6507
rect 15965 6449 16010 6465
rect 15865 6397 15931 6439
rect 16049 6439 16069 6473
rect 16103 6439 16119 6473
rect 16408 6473 16442 6619
rect 16588 6611 16632 6627
rect 16666 6593 16700 6737
rect 16975 6745 16988 6771
rect 17009 6711 17022 6737
rect 16734 6703 16935 6711
rect 16734 6669 16896 6703
rect 16930 6669 16935 6703
rect 16975 6695 17022 6711
rect 17070 6745 17111 6761
rect 17070 6711 17077 6745
rect 16734 6663 16935 6669
rect 16734 6661 16800 6663
rect 16734 6627 16750 6661
rect 16784 6627 16800 6661
rect 17070 6641 17111 6711
rect 16987 6635 17111 6641
rect 16862 6593 16878 6627
rect 16912 6593 16928 6627
rect 16480 6559 16496 6593
rect 16530 6573 16546 6593
rect 16530 6567 16562 6573
rect 16480 6533 16528 6559
rect 16666 6559 16928 6593
rect 16987 6601 16988 6635
rect 17022 6605 17111 6635
rect 17145 6661 17179 6830
rect 17491 6831 17507 6865
rect 17541 6831 17718 6865
rect 17752 6831 17768 6865
rect 17351 6797 17385 6805
rect 17802 6828 17859 6873
rect 17213 6763 17768 6797
rect 17213 6745 17263 6763
rect 17247 6711 17263 6745
rect 17213 6695 17263 6711
rect 17145 6645 17415 6661
rect 17145 6627 17381 6645
rect 17022 6601 17044 6605
rect 16987 6571 17044 6601
rect 16666 6533 16710 6559
rect 16480 6527 16562 6533
rect 16644 6499 16660 6533
rect 16694 6499 16710 6533
rect 16987 6537 17010 6571
rect 16744 6507 16778 6523
rect 16987 6521 17044 6537
rect 16153 6441 16187 6457
rect 16049 6397 16119 6439
rect 16243 6439 16259 6473
rect 16293 6439 16442 6473
rect 16243 6433 16442 6439
rect 16476 6469 16510 6485
rect 16476 6397 16510 6435
rect 16544 6455 16560 6489
rect 16594 6465 16610 6489
rect 17145 6473 17179 6627
rect 17371 6611 17381 6627
rect 17371 6595 17415 6611
rect 17254 6567 17273 6593
rect 17254 6533 17264 6567
rect 17307 6559 17329 6593
rect 17298 6533 17329 6559
rect 17449 6536 17485 6763
rect 17254 6527 17329 6533
rect 17419 6533 17485 6536
rect 17419 6499 17435 6533
rect 17469 6499 17485 6533
rect 17519 6703 17621 6729
rect 17519 6669 17540 6703
rect 17574 6695 17621 6703
rect 17655 6695 17671 6729
rect 17519 6661 17574 6669
rect 17553 6627 17574 6661
rect 17734 6645 17768 6763
rect 17836 6794 17859 6828
rect 17802 6760 17859 6794
rect 17836 6726 17859 6760
rect 17802 6706 17859 6726
rect 17519 6565 17574 6627
rect 17625 6634 17700 6645
rect 17625 6600 17649 6634
rect 17683 6633 17700 6634
rect 17625 6599 17650 6600
rect 17684 6599 17700 6633
rect 17734 6629 17784 6645
rect 17734 6595 17750 6629
rect 17734 6579 17784 6595
rect 17519 6531 17657 6565
rect 16744 6465 16778 6473
rect 16594 6455 16778 6465
rect 16544 6431 16778 6455
rect 16832 6439 16848 6473
rect 16882 6439 16898 6473
rect 16832 6397 16898 6439
rect 17026 6439 17042 6473
rect 17076 6439 17179 6473
rect 17026 6433 17179 6439
rect 17215 6469 17267 6485
rect 17215 6435 17233 6469
rect 17215 6397 17267 6435
rect 17319 6455 17335 6489
rect 17369 6465 17385 6489
rect 17519 6481 17553 6497
rect 17369 6455 17519 6465
rect 17319 6447 17519 6455
rect 17319 6431 17553 6447
rect 17610 6483 17657 6531
rect 17610 6449 17623 6483
rect 17610 6433 17657 6449
rect 17702 6473 17768 6541
rect 17818 6523 17859 6706
rect 17702 6439 17718 6473
rect 17752 6439 17768 6473
rect 17702 6397 17768 6439
rect 17802 6507 17859 6523
rect 17836 6473 17859 6507
rect 17802 6431 17859 6473
rect 17893 6847 17956 6863
rect 17893 6813 17906 6847
rect 17940 6813 17956 6847
rect 17893 6779 17956 6813
rect 17893 6745 17906 6779
rect 17940 6745 17956 6779
rect 17893 6645 17956 6745
rect 17992 6853 18051 6907
rect 17992 6819 18001 6853
rect 18035 6819 18051 6853
rect 17992 6785 18051 6819
rect 17992 6751 18001 6785
rect 18035 6751 18051 6785
rect 17992 6733 18051 6751
rect 18085 6829 18137 6873
rect 18119 6795 18137 6829
rect 18085 6761 18137 6795
rect 18119 6727 18137 6761
rect 18085 6669 18137 6727
rect 17893 6629 18060 6645
rect 17893 6595 18026 6629
rect 17893 6579 18060 6595
rect 17893 6499 17956 6579
rect 18094 6545 18137 6669
rect 17893 6465 17906 6499
rect 17940 6465 17956 6499
rect 18085 6509 18137 6545
rect 18119 6502 18137 6509
rect 17893 6431 17956 6465
rect 17992 6473 18051 6489
rect 17992 6439 18001 6473
rect 18035 6439 18051 6473
rect 17992 6397 18051 6439
rect 18085 6468 18092 6475
rect 18126 6468 18137 6502
rect 18085 6431 18137 6468
rect 13370 6363 13399 6397
rect 13433 6363 13491 6397
rect 13525 6363 13583 6397
rect 13617 6363 13675 6397
rect 13709 6363 13767 6397
rect 13801 6363 13859 6397
rect 13893 6363 13951 6397
rect 13985 6363 14043 6397
rect 14077 6363 14135 6397
rect 14169 6363 14227 6397
rect 14261 6363 14319 6397
rect 14353 6363 14411 6397
rect 14445 6363 14503 6397
rect 14537 6363 14595 6397
rect 14629 6363 14687 6397
rect 14721 6363 14779 6397
rect 14813 6363 14871 6397
rect 14905 6363 14963 6397
rect 14997 6363 15055 6397
rect 15089 6363 15147 6397
rect 15181 6363 15239 6397
rect 15273 6363 15331 6397
rect 15365 6363 15423 6397
rect 15457 6363 15515 6397
rect 15549 6363 15607 6397
rect 15641 6363 15699 6397
rect 15733 6363 15791 6397
rect 15825 6363 15883 6397
rect 15917 6363 15975 6397
rect 16009 6363 16067 6397
rect 16101 6363 16159 6397
rect 16193 6363 16251 6397
rect 16285 6363 16343 6397
rect 16377 6363 16435 6397
rect 16469 6363 16527 6397
rect 16561 6363 16619 6397
rect 16653 6363 16711 6397
rect 16745 6363 16803 6397
rect 16837 6363 16895 6397
rect 16929 6363 16987 6397
rect 17021 6363 17079 6397
rect 17113 6363 17171 6397
rect 17205 6363 17263 6397
rect 17297 6363 17355 6397
rect 17389 6363 17447 6397
rect 17481 6363 17539 6397
rect 17573 6363 17631 6397
rect 17665 6363 17723 6397
rect 17757 6363 17815 6397
rect 17849 6363 17907 6397
rect 17941 6363 17999 6397
rect 18033 6363 18091 6397
rect 18125 6363 18154 6397
rect 13370 6350 18154 6363
rect 13370 6316 13399 6350
rect 13433 6316 13491 6350
rect 13525 6316 13583 6350
rect 13617 6316 13675 6350
rect 13709 6316 13767 6350
rect 13801 6316 13859 6350
rect 13893 6316 13951 6350
rect 13985 6316 14043 6350
rect 14077 6316 14135 6350
rect 14169 6316 14227 6350
rect 14261 6316 14319 6350
rect 14353 6316 14411 6350
rect 14445 6316 14503 6350
rect 14537 6316 14595 6350
rect 14629 6316 14687 6350
rect 14721 6316 14779 6350
rect 14813 6316 14871 6350
rect 14905 6316 14964 6350
rect 14998 6316 15055 6350
rect 15089 6316 15147 6350
rect 15181 6316 15239 6350
rect 15273 6316 15332 6350
rect 15366 6316 15423 6350
rect 15457 6316 15515 6350
rect 15549 6316 15607 6350
rect 15641 6316 15699 6350
rect 15733 6316 15791 6350
rect 15825 6316 15883 6350
rect 15917 6316 15975 6350
rect 16009 6316 16067 6350
rect 16101 6316 16159 6350
rect 16193 6316 16251 6350
rect 16285 6316 16343 6350
rect 16377 6316 16435 6350
rect 16469 6316 16526 6350
rect 16560 6316 16618 6350
rect 16652 6316 16711 6350
rect 16745 6316 16803 6350
rect 16837 6316 16895 6350
rect 16929 6316 16986 6350
rect 17020 6316 17079 6350
rect 17113 6316 17170 6350
rect 17204 6316 17263 6350
rect 17297 6316 17355 6350
rect 17389 6316 17447 6350
rect 17481 6316 17539 6350
rect 17573 6316 17631 6350
rect 17665 6316 17723 6350
rect 17757 6316 17815 6350
rect 17849 6316 17907 6350
rect 17941 6316 17999 6350
rect 18033 6316 18091 6350
rect 18125 6316 18154 6350
rect 13370 6301 18154 6316
rect 13370 6267 13399 6301
rect 13433 6267 13491 6301
rect 13525 6267 13583 6301
rect 13617 6267 13675 6301
rect 13709 6267 13767 6301
rect 13801 6267 13859 6301
rect 13893 6267 13951 6301
rect 13985 6267 14043 6301
rect 14077 6267 14135 6301
rect 14169 6267 14227 6301
rect 14261 6267 14319 6301
rect 14353 6267 14411 6301
rect 14445 6267 14503 6301
rect 14537 6267 14595 6301
rect 14629 6267 14687 6301
rect 14721 6267 14779 6301
rect 14813 6267 14871 6301
rect 14905 6267 14963 6301
rect 14997 6267 15055 6301
rect 15089 6267 15147 6301
rect 15181 6267 15239 6301
rect 15273 6267 15331 6301
rect 15365 6267 15423 6301
rect 15457 6267 15515 6301
rect 15549 6267 15607 6301
rect 15641 6267 15699 6301
rect 15733 6267 15791 6301
rect 15825 6267 15883 6301
rect 15917 6267 15975 6301
rect 16009 6267 16067 6301
rect 16101 6267 16159 6301
rect 16193 6267 16251 6301
rect 16285 6267 16343 6301
rect 16377 6267 16435 6301
rect 16469 6267 16527 6301
rect 16561 6267 16619 6301
rect 16653 6267 16711 6301
rect 16745 6267 16803 6301
rect 16837 6267 16895 6301
rect 16929 6267 16987 6301
rect 17021 6267 17079 6301
rect 17113 6267 17171 6301
rect 17205 6267 17263 6301
rect 17297 6267 17355 6301
rect 17389 6267 17447 6301
rect 17481 6267 17539 6301
rect 17573 6267 17631 6301
rect 17665 6267 17723 6301
rect 17757 6267 17815 6301
rect 17849 6267 17907 6301
rect 17941 6267 17999 6301
rect 18033 6267 18091 6301
rect 18125 6267 18154 6301
rect 13473 6225 13539 6267
rect 13387 6199 13439 6215
rect 13387 6165 13405 6199
rect 13473 6191 13489 6225
rect 13523 6191 13539 6225
rect 13657 6225 13727 6267
rect 13573 6199 13618 6215
rect 13387 6157 13439 6165
rect 13607 6165 13618 6199
rect 13657 6191 13677 6225
rect 13711 6191 13727 6225
rect 13851 6225 14050 6231
rect 13761 6207 13795 6223
rect 13387 6123 13538 6157
rect 13387 6055 13419 6089
rect 13453 6055 13458 6089
rect 13387 6054 13458 6055
rect 13387 6020 13402 6054
rect 13436 6020 13458 6054
rect 13387 5959 13458 6020
rect 13492 6054 13538 6123
rect 13492 6020 13504 6054
rect 13492 5927 13538 6020
rect 13387 5909 13492 5925
rect 13387 5875 13405 5909
rect 13439 5893 13492 5909
rect 13526 5893 13538 5927
rect 13439 5891 13538 5893
rect 13573 6131 13618 6165
rect 13851 6191 13867 6225
rect 13901 6191 14050 6225
rect 13761 6157 13795 6173
rect 13573 6097 13584 6131
rect 13573 5909 13618 6097
rect 13387 5841 13439 5875
rect 13607 5875 13618 5909
rect 13652 6119 13795 6157
rect 13836 6127 13880 6143
rect 13652 5925 13686 6119
rect 13870 6093 13880 6127
rect 13720 6067 13802 6083
rect 13754 6033 13802 6067
rect 13720 6005 13802 6033
rect 13720 5971 13746 6005
rect 13780 5971 13802 6005
rect 13720 5959 13802 5971
rect 13836 5969 13880 6093
rect 13916 6131 13982 6155
rect 13916 6115 13948 6131
rect 13916 6081 13932 6115
rect 13966 6081 13982 6097
rect 14016 6045 14050 6191
rect 14084 6229 14118 6267
rect 14084 6179 14118 6195
rect 14152 6209 14386 6233
rect 14152 6175 14168 6209
rect 14202 6199 14386 6209
rect 14202 6175 14218 6199
rect 14352 6191 14386 6199
rect 14440 6225 14506 6267
rect 14440 6191 14456 6225
rect 14490 6191 14506 6225
rect 14634 6225 14787 6231
rect 14634 6191 14650 6225
rect 14684 6191 14787 6225
rect 14088 6131 14170 6137
rect 14252 6131 14268 6165
rect 14302 6131 14318 6165
rect 14352 6141 14386 6157
rect 14088 6105 14136 6131
rect 14088 6071 14104 6105
rect 14138 6091 14170 6097
rect 14274 6105 14318 6131
rect 14595 6127 14652 6143
rect 14138 6071 14154 6091
rect 14274 6071 14536 6105
rect 13970 6037 14050 6045
rect 14196 6037 14240 6053
rect 13970 6003 14206 6037
rect 13836 5953 13936 5969
rect 13836 5927 13902 5953
rect 13652 5891 13795 5925
rect 13836 5893 13860 5927
rect 13894 5919 13902 5927
rect 13894 5893 13936 5919
rect 13387 5807 13405 5841
rect 13387 5791 13439 5807
rect 13473 5823 13489 5857
rect 13523 5823 13539 5857
rect 13473 5757 13539 5823
rect 13573 5841 13618 5875
rect 13607 5807 13618 5841
rect 13573 5791 13618 5807
rect 13657 5823 13677 5857
rect 13711 5823 13727 5857
rect 13657 5757 13727 5823
rect 13761 5841 13795 5891
rect 13970 5834 14004 6003
rect 14190 5987 14240 6003
rect 14038 5953 14088 5969
rect 14072 5927 14088 5953
rect 14274 5927 14308 6071
rect 14470 6037 14486 6071
rect 14520 6037 14536 6071
rect 14595 6093 14618 6127
rect 14595 6063 14652 6093
rect 14342 6003 14358 6037
rect 14392 6003 14408 6037
rect 14595 6029 14596 6063
rect 14630 6059 14652 6063
rect 14630 6029 14719 6059
rect 14595 6023 14719 6029
rect 14342 6001 14408 6003
rect 14342 5995 14543 6001
rect 14342 5961 14504 5995
rect 14538 5961 14543 5995
rect 14342 5953 14543 5961
rect 14583 5953 14630 5969
rect 14072 5919 14188 5927
rect 14038 5893 14188 5919
rect 14222 5893 14308 5927
rect 14617 5927 14630 5953
rect 14038 5877 14308 5893
rect 14188 5859 14222 5877
rect 13761 5791 13795 5807
rect 13838 5800 13854 5834
rect 13888 5800 14004 5834
rect 14052 5809 14068 5843
rect 14102 5809 14128 5843
rect 14188 5809 14222 5825
rect 14346 5867 14362 5901
rect 14396 5867 14412 5901
rect 14583 5893 14596 5919
rect 14678 5953 14719 6023
rect 14678 5919 14685 5953
rect 14678 5903 14719 5919
rect 14753 6037 14787 6191
rect 14823 6229 14875 6267
rect 14823 6195 14841 6229
rect 14823 6179 14875 6195
rect 14927 6217 15161 6233
rect 14927 6209 15127 6217
rect 14927 6175 14943 6209
rect 14977 6199 15127 6209
rect 14977 6175 14993 6199
rect 15127 6167 15161 6183
rect 15218 6215 15265 6231
rect 15218 6181 15231 6215
rect 14862 6131 14937 6137
rect 14862 6097 14872 6131
rect 14906 6105 14937 6131
rect 15027 6131 15043 6165
rect 15077 6131 15093 6165
rect 15218 6133 15265 6181
rect 15027 6128 15093 6131
rect 14862 6071 14881 6097
rect 14915 6071 14937 6105
rect 14979 6053 15023 6069
rect 14979 6037 14989 6053
rect 14753 6019 14989 6037
rect 14753 6003 15023 6019
rect 14583 5887 14630 5893
rect 14346 5833 14412 5867
rect 14753 5834 14787 6003
rect 14821 5953 14871 5969
rect 14855 5919 14871 5953
rect 14821 5901 14871 5919
rect 15057 5901 15093 6128
rect 15127 6099 15265 6133
rect 15310 6225 15376 6267
rect 15310 6191 15326 6225
rect 15360 6191 15376 6225
rect 15310 6123 15376 6191
rect 15410 6191 15467 6233
rect 15444 6157 15467 6191
rect 15410 6141 15467 6157
rect 15127 6037 15182 6099
rect 15342 6069 15392 6085
rect 15161 6003 15182 6037
rect 15233 6031 15258 6065
rect 15292 6063 15308 6065
rect 15233 6029 15265 6031
rect 15299 6029 15308 6063
rect 15233 6019 15308 6029
rect 15342 6035 15358 6069
rect 15342 6019 15392 6035
rect 15127 5995 15182 6003
rect 15127 5961 15148 5995
rect 15182 5961 15229 5969
rect 15127 5935 15229 5961
rect 15263 5935 15279 5969
rect 15342 5901 15376 6019
rect 15426 5958 15467 6141
rect 14821 5867 15376 5901
rect 15410 5938 15467 5958
rect 15444 5904 15467 5938
rect 15410 5870 15467 5904
rect 14052 5757 14128 5809
rect 14346 5799 14362 5833
rect 14396 5799 14412 5833
rect 14621 5800 14637 5834
rect 14671 5800 14787 5834
rect 14959 5859 14993 5867
rect 14346 5757 14412 5799
rect 14835 5799 14851 5833
rect 14885 5799 14911 5833
rect 15444 5836 15467 5870
rect 14959 5809 14993 5825
rect 14835 5757 14911 5799
rect 15099 5799 15115 5833
rect 15149 5799 15326 5833
rect 15360 5799 15376 5833
rect 15099 5757 15376 5799
rect 15410 5791 15467 5836
rect 15501 6199 15564 6233
rect 15501 6165 15514 6199
rect 15548 6165 15564 6199
rect 15600 6225 15659 6267
rect 15600 6191 15609 6225
rect 15643 6191 15659 6225
rect 15600 6175 15659 6191
rect 15693 6189 15745 6233
rect 15865 6225 15931 6267
rect 15501 6085 15564 6165
rect 15727 6155 15745 6189
rect 15693 6119 15745 6155
rect 15779 6199 15831 6215
rect 15779 6165 15797 6199
rect 15865 6191 15881 6225
rect 15915 6191 15931 6225
rect 16049 6225 16119 6267
rect 15965 6199 16010 6215
rect 15779 6157 15831 6165
rect 15999 6165 16010 6199
rect 16049 6191 16069 6225
rect 16103 6191 16119 6225
rect 16243 6225 16442 6231
rect 16153 6207 16187 6223
rect 15779 6123 15930 6157
rect 15501 6069 15668 6085
rect 15501 6035 15634 6069
rect 15501 6019 15668 6035
rect 15501 5919 15564 6019
rect 15702 5995 15745 6119
rect 15693 5937 15745 5995
rect 15779 6054 15850 6089
rect 15779 6020 15794 6054
rect 15828 6045 15850 6054
rect 15779 6011 15803 6020
rect 15837 6011 15850 6045
rect 15779 5959 15850 6011
rect 15884 6054 15930 6123
rect 15884 6020 15896 6054
rect 15501 5885 15514 5919
rect 15548 5885 15564 5919
rect 15501 5851 15564 5885
rect 15501 5817 15514 5851
rect 15548 5817 15564 5851
rect 15501 5801 15564 5817
rect 15600 5913 15659 5931
rect 15600 5879 15609 5913
rect 15643 5879 15659 5913
rect 15600 5845 15659 5879
rect 15600 5811 15609 5845
rect 15643 5811 15659 5845
rect 15600 5757 15659 5811
rect 15727 5903 15745 5937
rect 15884 5927 15930 6020
rect 15693 5869 15745 5903
rect 15727 5868 15745 5869
rect 15693 5834 15699 5835
rect 15733 5834 15745 5868
rect 15693 5791 15745 5834
rect 15779 5909 15884 5925
rect 15779 5875 15797 5909
rect 15831 5893 15884 5909
rect 15918 5893 15930 5927
rect 15831 5891 15930 5893
rect 15965 6131 16010 6165
rect 16243 6191 16259 6225
rect 16293 6191 16442 6225
rect 16153 6157 16187 6173
rect 15965 6097 15976 6131
rect 15965 5909 16010 6097
rect 15779 5841 15831 5875
rect 15999 5875 16010 5909
rect 16044 6119 16187 6157
rect 16228 6127 16272 6143
rect 16044 5925 16078 6119
rect 16262 6093 16272 6127
rect 16112 6067 16194 6083
rect 16146 6062 16194 6067
rect 16112 6028 16140 6033
rect 16174 6028 16194 6062
rect 16112 5959 16194 6028
rect 16228 5969 16272 6093
rect 16308 6131 16374 6155
rect 16308 6115 16340 6131
rect 16308 6081 16324 6115
rect 16358 6081 16374 6097
rect 16408 6045 16442 6191
rect 16476 6229 16510 6267
rect 16476 6179 16510 6195
rect 16544 6209 16778 6233
rect 16544 6175 16560 6209
rect 16594 6199 16778 6209
rect 16594 6175 16610 6199
rect 16744 6191 16778 6199
rect 16832 6225 16898 6267
rect 16832 6191 16848 6225
rect 16882 6191 16898 6225
rect 17026 6225 17179 6231
rect 17026 6191 17042 6225
rect 17076 6191 17179 6225
rect 16480 6131 16562 6137
rect 16644 6131 16660 6165
rect 16694 6131 16710 6165
rect 16744 6141 16778 6157
rect 16480 6105 16528 6131
rect 16480 6071 16496 6105
rect 16530 6091 16562 6097
rect 16666 6105 16710 6131
rect 16987 6127 17044 6143
rect 16530 6071 16546 6091
rect 16666 6071 16928 6105
rect 16362 6037 16442 6045
rect 16588 6037 16632 6053
rect 16362 6003 16598 6037
rect 16228 5953 16328 5969
rect 16228 5927 16294 5953
rect 16044 5891 16187 5925
rect 16228 5893 16252 5927
rect 16286 5919 16294 5927
rect 16286 5893 16328 5919
rect 15779 5807 15797 5841
rect 15779 5791 15831 5807
rect 15865 5823 15881 5857
rect 15915 5823 15931 5857
rect 15865 5757 15931 5823
rect 15965 5841 16010 5875
rect 15999 5807 16010 5841
rect 15965 5791 16010 5807
rect 16049 5823 16069 5857
rect 16103 5823 16119 5857
rect 16049 5757 16119 5823
rect 16153 5841 16187 5891
rect 16362 5834 16396 6003
rect 16582 5987 16632 6003
rect 16430 5953 16480 5969
rect 16464 5927 16480 5953
rect 16666 5927 16700 6071
rect 16862 6037 16878 6071
rect 16912 6037 16928 6071
rect 16987 6093 17010 6127
rect 16987 6063 17044 6093
rect 16734 6003 16750 6037
rect 16784 6003 16800 6037
rect 16987 6029 16988 6063
rect 17022 6059 17044 6063
rect 17022 6029 17111 6059
rect 16987 6023 17111 6029
rect 16734 6001 16800 6003
rect 16734 5995 16935 6001
rect 16734 5961 16896 5995
rect 16930 5961 16935 5995
rect 16734 5953 16935 5961
rect 16975 5953 17022 5969
rect 16464 5919 16580 5927
rect 16430 5893 16580 5919
rect 16614 5893 16700 5927
rect 17009 5927 17022 5953
rect 16430 5877 16700 5893
rect 16580 5859 16614 5877
rect 16153 5791 16187 5807
rect 16230 5800 16246 5834
rect 16280 5800 16396 5834
rect 16444 5809 16460 5843
rect 16494 5809 16520 5843
rect 16580 5809 16614 5825
rect 16738 5867 16754 5901
rect 16788 5867 16804 5901
rect 16975 5893 16988 5919
rect 17070 5953 17111 6023
rect 17070 5919 17077 5953
rect 17070 5903 17111 5919
rect 17145 6037 17179 6191
rect 17215 6229 17267 6267
rect 17215 6195 17233 6229
rect 17215 6179 17267 6195
rect 17319 6217 17553 6233
rect 17319 6209 17519 6217
rect 17319 6175 17335 6209
rect 17369 6199 17519 6209
rect 17369 6175 17385 6199
rect 17519 6167 17553 6183
rect 17610 6215 17657 6231
rect 17610 6181 17623 6215
rect 17254 6131 17329 6137
rect 17254 6097 17264 6131
rect 17298 6105 17329 6131
rect 17419 6131 17435 6165
rect 17469 6131 17485 6165
rect 17610 6133 17657 6181
rect 17419 6128 17485 6131
rect 17254 6071 17273 6097
rect 17307 6071 17329 6105
rect 17371 6053 17415 6069
rect 17371 6037 17381 6053
rect 17145 6019 17381 6037
rect 17145 6003 17415 6019
rect 16975 5887 17022 5893
rect 16738 5833 16804 5867
rect 17145 5834 17179 6003
rect 17213 5953 17263 5969
rect 17247 5919 17263 5953
rect 17213 5901 17263 5919
rect 17449 5901 17485 6128
rect 17519 6099 17657 6133
rect 17702 6225 17768 6267
rect 17702 6191 17718 6225
rect 17752 6191 17768 6225
rect 17702 6123 17768 6191
rect 17802 6191 17859 6233
rect 17836 6157 17859 6191
rect 17802 6141 17859 6157
rect 17519 6037 17574 6099
rect 17734 6069 17784 6085
rect 17553 6003 17574 6037
rect 17625 6031 17649 6065
rect 17684 6031 17700 6065
rect 17625 6019 17700 6031
rect 17734 6035 17750 6069
rect 17734 6019 17784 6035
rect 17519 5995 17574 6003
rect 17519 5961 17540 5995
rect 17574 5961 17621 5969
rect 17519 5935 17621 5961
rect 17655 5935 17671 5969
rect 17734 5901 17768 6019
rect 17818 5958 17859 6141
rect 17213 5867 17768 5901
rect 17802 5938 17859 5958
rect 17836 5904 17859 5938
rect 17802 5870 17859 5904
rect 16444 5757 16520 5809
rect 16738 5799 16754 5833
rect 16788 5799 16804 5833
rect 17013 5800 17029 5834
rect 17063 5800 17179 5834
rect 17351 5859 17385 5867
rect 16738 5757 16804 5799
rect 17227 5799 17243 5833
rect 17277 5799 17303 5833
rect 17836 5836 17859 5870
rect 17351 5809 17385 5825
rect 17227 5757 17303 5799
rect 17491 5799 17507 5833
rect 17541 5799 17718 5833
rect 17752 5799 17768 5833
rect 17491 5757 17768 5799
rect 17802 5791 17859 5836
rect 17893 6199 17956 6233
rect 17893 6165 17906 6199
rect 17940 6165 17956 6199
rect 17992 6225 18051 6267
rect 17992 6191 18001 6225
rect 18035 6191 18051 6225
rect 17992 6175 18051 6191
rect 18085 6189 18137 6233
rect 18119 6179 18137 6189
rect 17893 6085 17956 6165
rect 18085 6145 18086 6155
rect 18120 6145 18137 6179
rect 18085 6119 18137 6145
rect 17893 6069 18060 6085
rect 17893 6035 18026 6069
rect 17893 6019 18060 6035
rect 17893 5919 17956 6019
rect 18094 5995 18137 6119
rect 18085 5937 18137 5995
rect 17893 5885 17906 5919
rect 17940 5885 17956 5919
rect 17893 5851 17956 5885
rect 17893 5817 17906 5851
rect 17940 5817 17956 5851
rect 17893 5801 17956 5817
rect 17992 5913 18051 5931
rect 17992 5879 18001 5913
rect 18035 5879 18051 5913
rect 17992 5845 18051 5879
rect 17992 5811 18001 5845
rect 18035 5811 18051 5845
rect 17992 5757 18051 5811
rect 18119 5903 18137 5937
rect 18085 5869 18137 5903
rect 18119 5835 18137 5869
rect 18085 5791 18137 5835
rect 13370 5723 13399 5757
rect 13433 5723 13491 5757
rect 13525 5723 13583 5757
rect 13617 5723 13675 5757
rect 13709 5723 13767 5757
rect 13801 5723 13859 5757
rect 13893 5723 13951 5757
rect 13985 5723 14043 5757
rect 14077 5723 14135 5757
rect 14169 5723 14227 5757
rect 14261 5723 14319 5757
rect 14353 5723 14411 5757
rect 14445 5723 14503 5757
rect 14537 5723 14595 5757
rect 14629 5723 14687 5757
rect 14721 5723 14779 5757
rect 14813 5723 14871 5757
rect 14905 5723 14963 5757
rect 14997 5723 15055 5757
rect 15089 5723 15147 5757
rect 15181 5723 15239 5757
rect 15273 5723 15331 5757
rect 15365 5723 15423 5757
rect 15457 5723 15515 5757
rect 15549 5723 15607 5757
rect 15641 5723 15699 5757
rect 15733 5723 15791 5757
rect 15825 5723 15883 5757
rect 15917 5723 15975 5757
rect 16009 5723 16067 5757
rect 16101 5723 16159 5757
rect 16193 5723 16251 5757
rect 16285 5723 16343 5757
rect 16377 5723 16435 5757
rect 16469 5723 16527 5757
rect 16561 5723 16619 5757
rect 16653 5723 16711 5757
rect 16745 5723 16803 5757
rect 16837 5723 16895 5757
rect 16929 5723 16987 5757
rect 17021 5723 17079 5757
rect 17113 5723 17171 5757
rect 17205 5723 17263 5757
rect 17297 5723 17355 5757
rect 17389 5723 17447 5757
rect 17481 5723 17539 5757
rect 17573 5723 17631 5757
rect 17665 5723 17723 5757
rect 17757 5723 17815 5757
rect 17849 5723 17907 5757
rect 17941 5723 17999 5757
rect 18033 5723 18091 5757
rect 18125 5723 18154 5757
rect 13370 5708 18154 5723
rect 13370 5674 13402 5708
rect 13436 5674 13492 5708
rect 13526 5674 13585 5708
rect 13619 5674 13675 5708
rect 13709 5674 13766 5708
rect 13800 5674 13860 5708
rect 13894 5674 13951 5708
rect 13985 5674 14043 5708
rect 14077 5674 14135 5708
rect 14169 5674 14228 5708
rect 14262 5674 14319 5708
rect 14353 5674 14411 5708
rect 14445 5674 14503 5708
rect 14537 5674 14595 5708
rect 14629 5674 14688 5708
rect 14722 5674 14779 5708
rect 14813 5674 14870 5708
rect 14904 5674 14963 5708
rect 14997 5674 15056 5708
rect 15090 5674 15147 5708
rect 15181 5674 15239 5708
rect 15273 5674 15331 5708
rect 15365 5674 15423 5708
rect 15457 5674 15516 5708
rect 15550 5674 15606 5708
rect 15640 5674 15699 5708
rect 15733 5674 15791 5708
rect 15825 5674 15884 5708
rect 15918 5674 15978 5708
rect 16012 5674 16067 5708
rect 16101 5674 16159 5708
rect 16193 5674 16251 5708
rect 16285 5674 16343 5708
rect 16377 5674 16435 5708
rect 16469 5674 16527 5708
rect 16561 5674 16619 5708
rect 16653 5674 16711 5708
rect 16745 5674 16803 5708
rect 16837 5674 16895 5708
rect 16929 5674 16987 5708
rect 17021 5674 17079 5708
rect 17113 5674 17171 5708
rect 17205 5674 17263 5708
rect 17297 5674 17355 5708
rect 17389 5674 17447 5708
rect 17481 5674 17539 5708
rect 17573 5674 17631 5708
rect 17665 5674 17723 5708
rect 17757 5674 17815 5708
rect 17849 5674 17907 5708
rect 17941 5674 18000 5708
rect 18034 5674 18091 5708
rect 18125 5674 18154 5708
rect 13370 5661 18154 5674
rect 13370 5627 13399 5661
rect 13433 5627 13491 5661
rect 13525 5627 13583 5661
rect 13617 5627 13675 5661
rect 13709 5627 13767 5661
rect 13801 5627 13859 5661
rect 13893 5627 13951 5661
rect 13985 5627 14043 5661
rect 14077 5627 14135 5661
rect 14169 5627 14227 5661
rect 14261 5627 14319 5661
rect 14353 5627 14411 5661
rect 14445 5627 14503 5661
rect 14537 5627 14595 5661
rect 14629 5627 14687 5661
rect 14721 5627 14779 5661
rect 14813 5627 14871 5661
rect 14905 5627 14963 5661
rect 14997 5627 15055 5661
rect 15089 5627 15147 5661
rect 15181 5627 15239 5661
rect 15273 5627 15331 5661
rect 15365 5627 15423 5661
rect 15457 5627 15515 5661
rect 15549 5627 15607 5661
rect 15641 5627 15699 5661
rect 15733 5627 15791 5661
rect 15825 5627 15883 5661
rect 15917 5627 15975 5661
rect 16009 5627 16067 5661
rect 16101 5627 16159 5661
rect 16193 5627 16251 5661
rect 16285 5627 16343 5661
rect 16377 5627 16435 5661
rect 16469 5627 16527 5661
rect 16561 5627 16619 5661
rect 16653 5627 16711 5661
rect 16745 5627 16803 5661
rect 16837 5627 16895 5661
rect 16929 5627 16987 5661
rect 17021 5627 17079 5661
rect 17113 5627 17171 5661
rect 17205 5627 17263 5661
rect 17297 5627 17355 5661
rect 17389 5627 17447 5661
rect 17481 5627 17539 5661
rect 17573 5627 17631 5661
rect 17665 5627 17723 5661
rect 17757 5627 17815 5661
rect 17849 5627 17907 5661
rect 17941 5627 17999 5661
rect 18033 5627 18091 5661
rect 18125 5627 18154 5661
rect 13387 5577 13439 5593
rect 13387 5543 13405 5577
rect 13387 5509 13439 5543
rect 13473 5561 13539 5627
rect 13473 5527 13489 5561
rect 13523 5527 13539 5561
rect 13573 5577 13618 5593
rect 13607 5543 13618 5577
rect 13387 5475 13405 5509
rect 13573 5509 13618 5543
rect 13657 5561 13727 5627
rect 13657 5527 13677 5561
rect 13711 5527 13727 5561
rect 13761 5577 13795 5593
rect 13838 5550 13854 5584
rect 13888 5550 14004 5584
rect 13439 5491 13538 5493
rect 13439 5475 13492 5491
rect 13387 5459 13492 5475
rect 13526 5457 13538 5491
rect 13387 5364 13458 5425
rect 13387 5330 13402 5364
rect 13436 5330 13458 5364
rect 13387 5329 13458 5330
rect 13387 5295 13415 5329
rect 13449 5295 13458 5329
rect 13492 5364 13538 5457
rect 13492 5330 13504 5364
rect 13492 5261 13538 5330
rect 13387 5227 13538 5261
rect 13607 5475 13618 5509
rect 13761 5493 13795 5543
rect 13573 5287 13618 5475
rect 13573 5253 13584 5287
rect 13387 5219 13439 5227
rect 13387 5185 13405 5219
rect 13573 5219 13618 5253
rect 13652 5459 13795 5493
rect 13652 5265 13686 5459
rect 13836 5457 13860 5491
rect 13894 5465 13936 5491
rect 13894 5457 13902 5465
rect 13836 5431 13902 5457
rect 13720 5413 13802 5425
rect 13720 5379 13743 5413
rect 13777 5379 13802 5413
rect 13720 5351 13802 5379
rect 13754 5317 13802 5351
rect 13720 5301 13802 5317
rect 13836 5415 13936 5431
rect 13836 5291 13880 5415
rect 13970 5381 14004 5550
rect 14052 5575 14128 5627
rect 14346 5585 14412 5627
rect 14052 5541 14068 5575
rect 14102 5541 14128 5575
rect 14188 5559 14222 5575
rect 14188 5507 14222 5525
rect 14346 5551 14362 5585
rect 14396 5551 14412 5585
rect 14835 5585 14911 5627
rect 14346 5517 14412 5551
rect 14621 5550 14637 5584
rect 14671 5550 14787 5584
rect 14835 5551 14851 5585
rect 14885 5551 14911 5585
rect 15099 5585 15376 5627
rect 14959 5559 14993 5575
rect 14038 5491 14308 5507
rect 14038 5465 14188 5491
rect 14072 5457 14188 5465
rect 14222 5457 14308 5491
rect 14346 5483 14362 5517
rect 14396 5483 14412 5517
rect 14583 5491 14630 5497
rect 14072 5431 14088 5457
rect 14038 5415 14088 5431
rect 14190 5381 14240 5397
rect 13970 5347 14206 5381
rect 13970 5339 14050 5347
rect 13652 5227 13795 5265
rect 13870 5257 13880 5291
rect 13836 5241 13880 5257
rect 13916 5269 13932 5303
rect 13966 5287 13982 5303
rect 13916 5253 13948 5269
rect 13916 5229 13982 5253
rect 13387 5169 13439 5185
rect 13473 5159 13489 5193
rect 13523 5159 13539 5193
rect 13607 5185 13618 5219
rect 13761 5211 13795 5227
rect 13573 5169 13618 5185
rect 13473 5117 13539 5159
rect 13657 5159 13677 5193
rect 13711 5159 13727 5193
rect 14016 5193 14050 5339
rect 14196 5331 14240 5347
rect 14274 5313 14308 5457
rect 14583 5465 14596 5491
rect 14617 5431 14630 5457
rect 14342 5423 14543 5431
rect 14342 5389 14504 5423
rect 14538 5389 14543 5423
rect 14583 5415 14630 5431
rect 14678 5465 14719 5481
rect 14678 5431 14685 5465
rect 14342 5383 14543 5389
rect 14342 5381 14408 5383
rect 14342 5347 14358 5381
rect 14392 5347 14408 5381
rect 14678 5361 14719 5431
rect 14595 5355 14719 5361
rect 14470 5313 14486 5347
rect 14520 5313 14536 5347
rect 14088 5279 14104 5313
rect 14138 5293 14154 5313
rect 14138 5287 14170 5293
rect 14088 5253 14136 5279
rect 14274 5279 14536 5313
rect 14595 5321 14596 5355
rect 14630 5325 14719 5355
rect 14753 5381 14787 5550
rect 15099 5551 15115 5585
rect 15149 5551 15326 5585
rect 15360 5551 15376 5585
rect 14959 5517 14993 5525
rect 15410 5548 15467 5593
rect 14821 5483 15376 5517
rect 14821 5465 14871 5483
rect 14855 5431 14871 5465
rect 14821 5415 14871 5431
rect 14753 5365 15023 5381
rect 14753 5347 14989 5365
rect 14630 5321 14652 5325
rect 14595 5291 14652 5321
rect 14274 5253 14318 5279
rect 14088 5247 14170 5253
rect 14252 5219 14268 5253
rect 14302 5219 14318 5253
rect 14595 5257 14618 5291
rect 14352 5227 14386 5243
rect 14595 5241 14652 5257
rect 13761 5161 13795 5177
rect 13657 5117 13727 5159
rect 13851 5159 13867 5193
rect 13901 5159 14050 5193
rect 13851 5153 14050 5159
rect 14084 5189 14118 5205
rect 14084 5117 14118 5155
rect 14152 5175 14168 5209
rect 14202 5185 14218 5209
rect 14753 5193 14787 5347
rect 14979 5331 14989 5347
rect 14979 5315 15023 5331
rect 14862 5287 14881 5313
rect 14862 5253 14872 5287
rect 14915 5279 14937 5313
rect 14906 5253 14937 5279
rect 15057 5256 15093 5483
rect 14862 5247 14937 5253
rect 15027 5253 15093 5256
rect 15027 5219 15043 5253
rect 15077 5219 15093 5253
rect 15127 5423 15229 5449
rect 15127 5389 15148 5423
rect 15182 5415 15229 5423
rect 15263 5415 15279 5449
rect 15127 5381 15182 5389
rect 15161 5347 15182 5381
rect 15342 5365 15376 5483
rect 15444 5514 15467 5548
rect 15410 5480 15467 5514
rect 15444 5446 15467 5480
rect 15410 5426 15467 5446
rect 15127 5285 15182 5347
rect 15233 5353 15308 5365
rect 15233 5319 15257 5353
rect 15292 5319 15308 5353
rect 15342 5349 15392 5365
rect 15342 5315 15358 5349
rect 15342 5299 15392 5315
rect 15127 5251 15265 5285
rect 14352 5185 14386 5193
rect 14202 5175 14386 5185
rect 14152 5151 14386 5175
rect 14440 5159 14456 5193
rect 14490 5159 14506 5193
rect 14440 5117 14506 5159
rect 14634 5159 14650 5193
rect 14684 5159 14787 5193
rect 14634 5153 14787 5159
rect 14823 5189 14875 5205
rect 14823 5155 14841 5189
rect 14823 5117 14875 5155
rect 14927 5175 14943 5209
rect 14977 5185 14993 5209
rect 15127 5201 15161 5217
rect 14977 5175 15127 5185
rect 14927 5167 15127 5175
rect 14927 5151 15161 5167
rect 15218 5203 15265 5251
rect 15218 5169 15231 5203
rect 15218 5153 15265 5169
rect 15310 5193 15376 5261
rect 15426 5243 15467 5426
rect 15310 5159 15326 5193
rect 15360 5159 15376 5193
rect 15310 5117 15376 5159
rect 15410 5227 15467 5243
rect 15444 5193 15467 5227
rect 15410 5151 15467 5193
rect 15501 5567 15564 5583
rect 15501 5533 15514 5567
rect 15548 5533 15564 5567
rect 15501 5499 15564 5533
rect 15501 5465 15514 5499
rect 15548 5465 15564 5499
rect 15501 5365 15564 5465
rect 15600 5573 15659 5627
rect 15600 5539 15609 5573
rect 15643 5539 15659 5573
rect 15600 5505 15659 5539
rect 15600 5471 15609 5505
rect 15643 5471 15659 5505
rect 15600 5453 15659 5471
rect 15693 5553 15745 5593
rect 15693 5549 15699 5553
rect 15733 5519 15745 5553
rect 15727 5515 15745 5519
rect 15693 5481 15745 5515
rect 15727 5447 15745 5481
rect 15779 5577 15831 5593
rect 15779 5543 15797 5577
rect 15779 5509 15831 5543
rect 15865 5561 15931 5627
rect 15865 5527 15881 5561
rect 15915 5527 15931 5561
rect 15965 5577 16010 5593
rect 15999 5543 16010 5577
rect 15779 5475 15797 5509
rect 15965 5509 16010 5543
rect 16049 5561 16119 5627
rect 16049 5527 16069 5561
rect 16103 5527 16119 5561
rect 16153 5577 16187 5593
rect 16230 5550 16246 5584
rect 16280 5550 16396 5584
rect 15831 5491 15930 5493
rect 15831 5475 15884 5491
rect 15779 5459 15884 5475
rect 15693 5389 15745 5447
rect 15918 5457 15930 5491
rect 15501 5349 15668 5365
rect 15501 5315 15634 5349
rect 15501 5299 15668 5315
rect 15501 5219 15564 5299
rect 15702 5265 15745 5389
rect 15779 5364 15850 5425
rect 15779 5330 15794 5364
rect 15828 5359 15850 5364
rect 15779 5325 15804 5330
rect 15838 5325 15850 5359
rect 15779 5295 15850 5325
rect 15884 5364 15930 5457
rect 15884 5330 15896 5364
rect 15501 5185 15514 5219
rect 15548 5185 15564 5219
rect 15693 5229 15745 5265
rect 15884 5261 15930 5330
rect 15501 5151 15564 5185
rect 15600 5193 15659 5209
rect 15600 5159 15609 5193
rect 15643 5159 15659 5193
rect 15600 5117 15659 5159
rect 15727 5195 15745 5229
rect 15693 5151 15745 5195
rect 15779 5227 15930 5261
rect 15999 5475 16010 5509
rect 16153 5493 16187 5543
rect 15965 5287 16010 5475
rect 15965 5253 15976 5287
rect 15779 5219 15831 5227
rect 15779 5185 15797 5219
rect 15965 5219 16010 5253
rect 16044 5459 16187 5493
rect 16044 5265 16078 5459
rect 16228 5457 16252 5491
rect 16286 5465 16328 5491
rect 16286 5457 16294 5465
rect 16228 5431 16294 5457
rect 16112 5354 16194 5425
rect 16112 5351 16141 5354
rect 16175 5320 16194 5354
rect 16146 5317 16194 5320
rect 16112 5301 16194 5317
rect 16228 5415 16328 5431
rect 16228 5291 16272 5415
rect 16362 5381 16396 5550
rect 16444 5575 16520 5627
rect 16738 5585 16804 5627
rect 16444 5541 16460 5575
rect 16494 5541 16520 5575
rect 16580 5559 16614 5575
rect 16580 5507 16614 5525
rect 16738 5551 16754 5585
rect 16788 5551 16804 5585
rect 17227 5585 17303 5627
rect 16738 5517 16804 5551
rect 17013 5550 17029 5584
rect 17063 5550 17179 5584
rect 17227 5551 17243 5585
rect 17277 5551 17303 5585
rect 17491 5585 17768 5627
rect 17351 5559 17385 5575
rect 16430 5491 16700 5507
rect 16430 5465 16580 5491
rect 16464 5457 16580 5465
rect 16614 5457 16700 5491
rect 16738 5483 16754 5517
rect 16788 5483 16804 5517
rect 16975 5491 17022 5497
rect 16464 5431 16480 5457
rect 16430 5415 16480 5431
rect 16582 5381 16632 5397
rect 16362 5347 16598 5381
rect 16362 5339 16442 5347
rect 16044 5227 16187 5265
rect 16262 5257 16272 5291
rect 16228 5241 16272 5257
rect 16308 5269 16324 5303
rect 16358 5287 16374 5303
rect 16308 5253 16340 5269
rect 16308 5229 16374 5253
rect 15779 5169 15831 5185
rect 15865 5159 15881 5193
rect 15915 5159 15931 5193
rect 15999 5185 16010 5219
rect 16153 5211 16187 5227
rect 15965 5169 16010 5185
rect 15865 5117 15931 5159
rect 16049 5159 16069 5193
rect 16103 5159 16119 5193
rect 16408 5193 16442 5339
rect 16588 5331 16632 5347
rect 16666 5313 16700 5457
rect 16975 5465 16988 5491
rect 17009 5431 17022 5457
rect 16734 5423 16935 5431
rect 16734 5389 16896 5423
rect 16930 5389 16935 5423
rect 16975 5415 17022 5431
rect 17070 5465 17111 5481
rect 17070 5431 17077 5465
rect 16734 5383 16935 5389
rect 16734 5381 16800 5383
rect 16734 5347 16750 5381
rect 16784 5347 16800 5381
rect 17070 5361 17111 5431
rect 16987 5355 17111 5361
rect 16862 5313 16878 5347
rect 16912 5313 16928 5347
rect 16480 5279 16496 5313
rect 16530 5293 16546 5313
rect 16530 5287 16562 5293
rect 16480 5253 16528 5279
rect 16666 5279 16928 5313
rect 16987 5321 16988 5355
rect 17022 5325 17111 5355
rect 17145 5381 17179 5550
rect 17491 5551 17507 5585
rect 17541 5551 17718 5585
rect 17752 5551 17768 5585
rect 17351 5517 17385 5525
rect 17802 5548 17859 5593
rect 17213 5483 17768 5517
rect 17213 5465 17263 5483
rect 17247 5431 17263 5465
rect 17213 5415 17263 5431
rect 17145 5365 17415 5381
rect 17145 5347 17381 5365
rect 17022 5321 17044 5325
rect 16987 5291 17044 5321
rect 16666 5253 16710 5279
rect 16480 5247 16562 5253
rect 16644 5219 16660 5253
rect 16694 5219 16710 5253
rect 16987 5257 17010 5291
rect 16744 5227 16778 5243
rect 16987 5241 17044 5257
rect 16153 5161 16187 5177
rect 16049 5117 16119 5159
rect 16243 5159 16259 5193
rect 16293 5159 16442 5193
rect 16243 5153 16442 5159
rect 16476 5189 16510 5205
rect 16476 5117 16510 5155
rect 16544 5175 16560 5209
rect 16594 5185 16610 5209
rect 17145 5193 17179 5347
rect 17371 5331 17381 5347
rect 17371 5315 17415 5331
rect 17254 5287 17273 5313
rect 17254 5253 17264 5287
rect 17307 5279 17329 5313
rect 17298 5253 17329 5279
rect 17449 5256 17485 5483
rect 17254 5247 17329 5253
rect 17419 5253 17485 5256
rect 17419 5219 17435 5253
rect 17469 5219 17485 5253
rect 17519 5423 17621 5449
rect 17519 5389 17540 5423
rect 17574 5415 17621 5423
rect 17655 5415 17671 5449
rect 17519 5381 17574 5389
rect 17553 5347 17574 5381
rect 17734 5365 17768 5483
rect 17836 5514 17859 5548
rect 17802 5480 17859 5514
rect 17836 5446 17859 5480
rect 17802 5426 17859 5446
rect 17519 5285 17574 5347
rect 17625 5354 17700 5365
rect 17625 5320 17649 5354
rect 17683 5353 17700 5354
rect 17625 5319 17650 5320
rect 17684 5319 17700 5353
rect 17734 5349 17784 5365
rect 17734 5315 17750 5349
rect 17734 5299 17784 5315
rect 17519 5251 17657 5285
rect 16744 5185 16778 5193
rect 16594 5175 16778 5185
rect 16544 5151 16778 5175
rect 16832 5159 16848 5193
rect 16882 5159 16898 5193
rect 16832 5117 16898 5159
rect 17026 5159 17042 5193
rect 17076 5159 17179 5193
rect 17026 5153 17179 5159
rect 17215 5189 17267 5205
rect 17215 5155 17233 5189
rect 17215 5117 17267 5155
rect 17319 5175 17335 5209
rect 17369 5185 17385 5209
rect 17519 5201 17553 5217
rect 17369 5175 17519 5185
rect 17319 5167 17519 5175
rect 17319 5151 17553 5167
rect 17610 5203 17657 5251
rect 17610 5169 17623 5203
rect 17610 5153 17657 5169
rect 17702 5193 17768 5261
rect 17818 5243 17859 5426
rect 17702 5159 17718 5193
rect 17752 5159 17768 5193
rect 17702 5117 17768 5159
rect 17802 5227 17859 5243
rect 17836 5193 17859 5227
rect 17802 5151 17859 5193
rect 17893 5567 17956 5583
rect 17893 5533 17906 5567
rect 17940 5533 17956 5567
rect 17893 5499 17956 5533
rect 17893 5465 17906 5499
rect 17940 5465 17956 5499
rect 17893 5365 17956 5465
rect 17992 5573 18051 5627
rect 17992 5539 18001 5573
rect 18035 5539 18051 5573
rect 17992 5505 18051 5539
rect 17992 5471 18001 5505
rect 18035 5471 18051 5505
rect 17992 5453 18051 5471
rect 18085 5549 18137 5593
rect 18119 5515 18137 5549
rect 18085 5481 18137 5515
rect 18119 5447 18137 5481
rect 18085 5389 18137 5447
rect 17893 5349 18060 5365
rect 17893 5315 18026 5349
rect 17893 5299 18060 5315
rect 17893 5219 17956 5299
rect 18094 5265 18137 5389
rect 17893 5185 17906 5219
rect 17940 5185 17956 5219
rect 18085 5229 18137 5265
rect 18119 5220 18137 5229
rect 17893 5151 17956 5185
rect 17992 5193 18051 5209
rect 17992 5159 18001 5193
rect 18035 5159 18051 5193
rect 17992 5117 18051 5159
rect 18085 5186 18087 5195
rect 18121 5186 18137 5220
rect 18085 5151 18137 5186
rect 13370 5049 13399 5117
rect 13433 5049 13491 5117
rect 13525 5049 13583 5117
rect 13617 5049 13675 5117
rect 13709 5049 13767 5117
rect 13801 5049 13859 5117
rect 13893 5049 13951 5117
rect 13985 5049 14043 5117
rect 14077 5049 14135 5117
rect 14169 5049 14227 5117
rect 14261 5049 14319 5117
rect 14353 5049 14411 5117
rect 14445 5049 14503 5117
rect 14537 5049 14595 5117
rect 14629 5049 14687 5117
rect 14721 5049 14779 5117
rect 14813 5049 14871 5117
rect 14905 5049 14963 5117
rect 14997 5049 15055 5117
rect 15089 5049 15147 5117
rect 15181 5049 15239 5117
rect 15273 5049 15331 5117
rect 15365 5049 15423 5117
rect 15457 5049 15515 5117
rect 15549 5049 15607 5117
rect 15641 5049 15699 5117
rect 15733 5049 15791 5117
rect 15825 5049 15883 5117
rect 15917 5049 15975 5117
rect 16009 5049 16067 5117
rect 16101 5049 16159 5117
rect 16193 5049 16251 5117
rect 16285 5049 16343 5117
rect 16377 5049 16435 5117
rect 16469 5049 16527 5117
rect 16561 5049 16619 5117
rect 16653 5049 16711 5117
rect 16745 5049 16803 5117
rect 16837 5049 16895 5117
rect 16929 5049 16987 5117
rect 17021 5049 17079 5117
rect 17113 5049 17171 5117
rect 17205 5049 17263 5117
rect 17297 5049 17355 5117
rect 17389 5049 17447 5117
rect 17481 5049 17539 5117
rect 17573 5049 17631 5117
rect 17665 5049 17723 5117
rect 17757 5049 17815 5117
rect 17849 5049 17907 5117
rect 17941 5049 17999 5117
rect 18033 5049 18091 5117
rect 18125 5049 18154 5117
<< viali >>
rect 12334 10507 12368 10567
rect 12422 10507 12456 10567
rect 12582 10557 12614 10591
rect 12614 10557 12616 10591
rect 12662 10557 12694 10591
rect 12694 10557 12696 10591
rect 12742 10557 12774 10591
rect 12774 10557 12776 10591
rect 12822 10557 12854 10591
rect 12854 10557 12856 10591
rect 12902 10557 12934 10591
rect 12934 10557 12936 10591
rect 12982 10557 13014 10591
rect 13014 10557 13016 10591
rect 13314 10560 13346 10594
rect 13346 10560 13348 10594
rect 13394 10560 13426 10594
rect 13426 10560 13428 10594
rect 13474 10560 13506 10594
rect 13506 10560 13508 10594
rect 13554 10560 13586 10594
rect 13586 10560 13588 10594
rect 13634 10560 13666 10594
rect 13666 10560 13668 10594
rect 13714 10560 13746 10594
rect 13746 10560 13748 10594
rect 13916 10560 13918 10594
rect 13918 10560 13950 10594
rect 13996 10560 13998 10594
rect 13998 10560 14030 10594
rect 14076 10560 14078 10594
rect 14078 10560 14110 10594
rect 14156 10560 14158 10594
rect 14158 10560 14190 10594
rect 14236 10560 14238 10594
rect 14238 10560 14270 10594
rect 14316 10560 14318 10594
rect 14318 10560 14350 10594
rect 14526 10560 14558 10594
rect 14558 10560 14560 10594
rect 14606 10560 14638 10594
rect 14638 10560 14640 10594
rect 14686 10560 14718 10594
rect 14718 10560 14720 10594
rect 14766 10560 14798 10594
rect 14798 10560 14800 10594
rect 14846 10560 14878 10594
rect 14878 10560 14880 10594
rect 14926 10560 14958 10594
rect 14958 10560 14960 10594
rect 15128 10560 15130 10594
rect 15130 10560 15162 10594
rect 15208 10560 15210 10594
rect 15210 10560 15242 10594
rect 15288 10560 15290 10594
rect 15290 10560 15322 10594
rect 15368 10560 15370 10594
rect 15370 10560 15402 10594
rect 15448 10560 15450 10594
rect 15450 10560 15482 10594
rect 15528 10560 15530 10594
rect 15530 10560 15562 10594
rect 15738 10560 15770 10594
rect 15770 10560 15772 10594
rect 15818 10560 15850 10594
rect 15850 10560 15852 10594
rect 15898 10560 15930 10594
rect 15930 10560 15932 10594
rect 15978 10560 16010 10594
rect 16010 10560 16012 10594
rect 16058 10560 16090 10594
rect 16090 10560 16092 10594
rect 16138 10560 16170 10594
rect 16170 10560 16172 10594
rect 16340 10560 16342 10594
rect 16342 10560 16374 10594
rect 16420 10560 16422 10594
rect 16422 10560 16454 10594
rect 16500 10560 16502 10594
rect 16502 10560 16534 10594
rect 16580 10560 16582 10594
rect 16582 10560 16614 10594
rect 16660 10560 16662 10594
rect 16662 10560 16694 10594
rect 16740 10560 16742 10594
rect 16742 10560 16774 10594
rect 16950 10560 16982 10594
rect 16982 10560 16984 10594
rect 17030 10560 17062 10594
rect 17062 10560 17064 10594
rect 17110 10560 17142 10594
rect 17142 10560 17144 10594
rect 17190 10560 17222 10594
rect 17222 10560 17224 10594
rect 17270 10560 17302 10594
rect 17302 10560 17304 10594
rect 17350 10560 17382 10594
rect 17382 10560 17384 10594
rect 17552 10560 17554 10594
rect 17554 10560 17586 10594
rect 17632 10560 17634 10594
rect 17634 10560 17666 10594
rect 17712 10560 17714 10594
rect 17714 10560 17746 10594
rect 17792 10560 17794 10594
rect 17794 10560 17826 10594
rect 17872 10560 17874 10594
rect 17874 10560 17906 10594
rect 17952 10560 17954 10594
rect 17954 10560 17986 10594
rect 12334 10369 12368 10429
rect 18294 10509 18328 10543
rect 12422 10369 12456 10429
rect 18299 10365 18333 10399
rect 12334 10231 12368 10291
rect 12422 10231 12456 10291
rect 18300 10213 18334 10247
rect 12334 10093 12368 10153
rect 12422 10093 12456 10153
rect 18300 10043 18334 10077
rect 11821 9962 11855 9996
rect 11913 9962 11947 9996
rect 12005 9991 12030 9996
rect 12030 9991 12039 9996
rect 12005 9962 12039 9991
rect 12097 9962 12131 9996
rect 12189 9962 12223 9996
rect 11949 9852 11983 9853
rect 11949 9819 11952 9852
rect 11952 9819 11983 9852
rect 11868 9684 11902 9688
rect 11868 9654 11872 9684
rect 11872 9654 11902 9684
rect 12058 9784 12092 9798
rect 12058 9764 12092 9784
rect 12334 9955 12368 10015
rect 12422 9955 12456 10015
rect 12334 9817 12368 9877
rect 12422 9817 12456 9877
rect 18299 9886 18333 9920
rect 12378 9724 12412 9758
rect 12142 9684 12176 9687
rect 12142 9653 12172 9684
rect 12172 9653 12176 9684
rect 12281 9654 12315 9688
rect 12319 9561 12353 9595
rect 12578 9579 12612 9613
rect 18501 9618 18535 9619
rect 18501 9585 18535 9618
rect 18593 9585 18627 9619
rect 18685 9618 18718 9619
rect 18718 9618 18719 9619
rect 18685 9585 18719 9618
rect 18777 9585 18811 9619
rect 12579 9486 12613 9520
rect 13020 9481 13054 9515
rect 13752 9484 13786 9518
rect 13878 9484 13912 9518
rect 14964 9484 14998 9518
rect 15090 9484 15124 9518
rect 16176 9484 16210 9518
rect 16302 9484 16336 9518
rect 17388 9484 17422 9518
rect 17514 9484 17548 9518
rect 18119 9506 18153 9566
rect 18207 9506 18241 9566
rect 11821 9418 11855 9452
rect 11913 9423 11947 9452
rect 12005 9423 12039 9452
rect 11913 9418 11920 9423
rect 11920 9418 11947 9423
rect 12005 9418 12038 9423
rect 12038 9418 12039 9423
rect 12097 9418 12131 9452
rect 12189 9418 12223 9452
rect 12976 9362 13010 9422
rect 13064 9365 13098 9425
rect 13708 9365 13742 9425
rect 13813 9365 13847 9425
rect 13922 9365 13956 9425
rect 14920 9365 14954 9425
rect 15024 9365 15058 9425
rect 15134 9365 15168 9425
rect 16132 9365 16166 9425
rect 16237 9365 16271 9425
rect 16346 9365 16380 9425
rect 17344 9365 17378 9425
rect 17451 9365 17485 9425
rect 17558 9365 17592 9425
rect 18119 9368 18153 9428
rect 18207 9368 18241 9428
rect 18303 9368 18337 9428
rect 18399 9368 18433 9428
rect 18048 9277 18082 9311
rect 18255 9275 18289 9309
rect 18495 9307 18529 9309
rect 18495 9275 18509 9307
rect 18509 9275 18529 9307
rect 18702 9275 18736 9309
rect 13329 9164 13363 9224
rect 13419 9164 13453 9224
rect 14061 9164 14095 9224
rect 14168 9164 14202 9224
rect 14271 9164 14305 9224
rect 15273 9164 15307 9224
rect 15379 9164 15413 9224
rect 15483 9164 15517 9224
rect 16611 9164 16645 9224
rect 16719 9164 16753 9224
rect 16821 9164 16855 9224
rect 17466 9164 17500 9224
rect 17555 9164 17589 9224
rect 18119 9165 18153 9225
rect 18207 9165 18241 9225
rect 18303 9165 18337 9225
rect 18399 9165 18433 9225
rect 12389 9090 12423 9124
rect 13373 9080 13407 9114
rect 14105 9080 14139 9114
rect 14227 9080 14261 9114
rect 15317 9080 15351 9114
rect 15439 9080 15473 9114
rect 16655 9080 16689 9114
rect 16777 9080 16811 9114
rect 17511 9080 17545 9114
rect 12309 8980 12343 9040
rect 12469 8980 12503 9040
rect 18119 9027 18153 9087
rect 18207 9027 18241 9087
rect 18501 9041 18535 9075
rect 18593 9041 18627 9075
rect 18685 9041 18719 9075
rect 18777 9041 18811 9075
rect 12309 8842 12343 8902
rect 12469 8842 12503 8902
rect 12309 8704 12343 8764
rect 12469 8704 12503 8764
rect 12309 8566 12343 8626
rect 12469 8566 12503 8626
rect 12309 8428 12343 8488
rect 12469 8428 12503 8488
rect 12309 8290 12343 8350
rect 12469 8290 12503 8350
rect 12309 8152 12343 8212
rect 12469 8152 12503 8212
rect 12309 8014 12343 8074
rect 12469 8014 12503 8074
rect 13010 7993 13044 8027
rect 13090 7993 13124 8027
rect 13170 7993 13204 8027
rect 13250 7993 13284 8027
rect 13742 7993 13776 8027
rect 13822 7993 13856 8027
rect 13902 7993 13936 8027
rect 13982 7993 14016 8027
rect 14350 7993 14384 8027
rect 14430 7993 14464 8027
rect 14510 7993 14544 8027
rect 14590 7993 14624 8027
rect 14954 7993 14988 8027
rect 15034 7993 15068 8027
rect 15114 7993 15148 8027
rect 15194 7993 15228 8027
rect 15562 7993 15596 8027
rect 15642 7993 15676 8027
rect 15722 7993 15756 8027
rect 15802 7993 15836 8027
rect 16292 7993 16326 8027
rect 16372 7993 16406 8027
rect 16452 7993 16486 8027
rect 16532 7993 16566 8027
rect 16900 7993 16934 8027
rect 16980 7993 17014 8027
rect 17060 7993 17094 8027
rect 17140 7993 17174 8027
rect 17634 7993 17668 8027
rect 17714 7993 17748 8027
rect 17794 7993 17828 8027
rect 17874 7993 17908 8027
rect 13399 7547 13433 7581
rect 13491 7547 13525 7581
rect 13583 7547 13617 7581
rect 13675 7547 13709 7581
rect 13767 7547 13801 7581
rect 13859 7547 13893 7581
rect 13951 7547 13985 7581
rect 14043 7547 14077 7581
rect 14135 7547 14169 7581
rect 14227 7547 14261 7581
rect 14319 7547 14353 7581
rect 14411 7547 14445 7581
rect 14503 7547 14537 7581
rect 14595 7547 14629 7581
rect 14687 7547 14721 7581
rect 14779 7547 14813 7581
rect 14871 7547 14905 7581
rect 14963 7547 14997 7581
rect 15055 7547 15089 7581
rect 15147 7547 15181 7581
rect 15239 7547 15273 7581
rect 15331 7547 15365 7581
rect 15423 7547 15457 7581
rect 15515 7547 15549 7581
rect 15607 7547 15641 7581
rect 15699 7547 15733 7581
rect 15791 7547 15825 7581
rect 15883 7547 15917 7581
rect 15975 7547 16009 7581
rect 16067 7547 16101 7581
rect 16159 7547 16193 7581
rect 16251 7547 16285 7581
rect 16343 7547 16377 7581
rect 16435 7547 16469 7581
rect 16527 7547 16561 7581
rect 16619 7547 16653 7581
rect 16711 7547 16745 7581
rect 16803 7547 16837 7581
rect 16895 7547 16929 7581
rect 16987 7547 17021 7581
rect 17079 7547 17113 7581
rect 17171 7547 17205 7581
rect 17263 7547 17297 7581
rect 17355 7547 17389 7581
rect 17447 7547 17481 7581
rect 17539 7547 17573 7581
rect 17631 7547 17665 7581
rect 17723 7547 17757 7581
rect 17815 7547 17849 7581
rect 17907 7547 17941 7581
rect 17999 7547 18033 7581
rect 18091 7547 18125 7581
rect 13416 7334 13450 7355
rect 13416 7321 13436 7334
rect 13436 7321 13450 7334
rect 13492 7173 13526 7207
rect 13584 7377 13618 7411
rect 13736 7247 13770 7281
rect 13948 7395 13982 7411
rect 13948 7377 13966 7395
rect 13966 7377 13982 7395
rect 14136 7385 14170 7411
rect 14136 7377 14138 7385
rect 14138 7377 14170 7385
rect 13860 7173 13894 7207
rect 14596 7309 14630 7343
rect 14504 7241 14538 7275
rect 14596 7199 14617 7207
rect 14617 7199 14630 7207
rect 14596 7173 14630 7199
rect 14872 7385 14906 7411
rect 14872 7377 14881 7385
rect 14881 7377 14906 7385
rect 15255 7311 15258 7340
rect 15258 7311 15289 7340
rect 15255 7306 15289 7311
rect 15148 7241 15182 7275
rect 15805 7300 15828 7310
rect 15828 7300 15839 7310
rect 15805 7276 15839 7300
rect 15703 7115 15727 7143
rect 15727 7115 15737 7143
rect 15703 7109 15737 7115
rect 15884 7173 15918 7207
rect 15976 7377 16010 7411
rect 16138 7313 16146 7343
rect 16146 7313 16172 7343
rect 16138 7309 16172 7313
rect 16340 7395 16374 7411
rect 16340 7377 16358 7395
rect 16358 7377 16374 7395
rect 16528 7385 16562 7411
rect 16528 7377 16530 7385
rect 16530 7377 16562 7385
rect 16252 7173 16286 7207
rect 16988 7309 17022 7343
rect 16896 7241 16930 7275
rect 16988 7199 17009 7207
rect 17009 7199 17022 7207
rect 16988 7173 17022 7199
rect 17264 7385 17298 7411
rect 17264 7377 17273 7385
rect 17273 7377 17298 7385
rect 17654 7311 17684 7344
rect 17684 7311 17688 7344
rect 17654 7310 17688 7311
rect 17540 7241 17574 7275
rect 18091 7435 18119 7460
rect 18119 7435 18125 7460
rect 18091 7426 18125 7435
rect 13399 7003 13433 7037
rect 13491 7003 13525 7037
rect 13583 7003 13617 7037
rect 13675 7003 13709 7037
rect 13767 7003 13801 7037
rect 13859 7003 13893 7037
rect 13951 7003 13985 7037
rect 14043 7003 14077 7037
rect 14135 7003 14169 7037
rect 14227 7003 14261 7037
rect 14319 7003 14353 7037
rect 14411 7003 14445 7037
rect 14503 7003 14537 7037
rect 14595 7003 14629 7037
rect 14687 7003 14721 7037
rect 14779 7003 14813 7037
rect 14871 7003 14905 7037
rect 14963 7003 14997 7037
rect 15055 7003 15089 7037
rect 15147 7003 15181 7037
rect 15239 7003 15273 7037
rect 15331 7003 15365 7037
rect 15423 7003 15457 7037
rect 15515 7003 15549 7037
rect 15607 7003 15641 7037
rect 15699 7003 15733 7037
rect 15791 7003 15825 7037
rect 15883 7003 15917 7037
rect 15975 7003 16009 7037
rect 16067 7003 16101 7037
rect 16159 7003 16193 7037
rect 16251 7003 16285 7037
rect 16343 7003 16377 7037
rect 16435 7003 16469 7037
rect 16527 7003 16561 7037
rect 16619 7003 16653 7037
rect 16711 7003 16745 7037
rect 16803 7003 16837 7037
rect 16895 7003 16929 7037
rect 16987 7003 17021 7037
rect 17079 7003 17113 7037
rect 17171 7003 17205 7037
rect 17263 7003 17297 7037
rect 17355 7003 17389 7037
rect 17447 7003 17481 7037
rect 17539 7003 17573 7037
rect 17631 7003 17665 7037
rect 17723 7003 17757 7037
rect 17815 7003 17849 7037
rect 17907 7003 17941 7037
rect 17999 7003 18033 7037
rect 18091 7003 18125 7037
rect 13399 6907 13433 6941
rect 13491 6907 13525 6941
rect 13583 6907 13617 6941
rect 13675 6907 13709 6941
rect 13767 6907 13801 6941
rect 13859 6907 13893 6941
rect 13951 6907 13985 6941
rect 14043 6907 14077 6941
rect 14135 6907 14169 6941
rect 14227 6907 14261 6941
rect 14319 6907 14353 6941
rect 14411 6907 14445 6941
rect 14503 6907 14537 6941
rect 14595 6907 14629 6941
rect 14687 6907 14721 6941
rect 14779 6907 14813 6941
rect 14871 6907 14905 6941
rect 14963 6907 14997 6941
rect 15055 6907 15089 6941
rect 15147 6907 15181 6941
rect 15239 6907 15273 6941
rect 15331 6907 15365 6941
rect 15423 6907 15457 6941
rect 15515 6907 15549 6941
rect 15607 6907 15641 6941
rect 15699 6907 15733 6941
rect 15791 6907 15825 6941
rect 15883 6907 15917 6941
rect 15975 6907 16009 6941
rect 16067 6907 16101 6941
rect 16159 6907 16193 6941
rect 16251 6907 16285 6941
rect 16343 6907 16377 6941
rect 16435 6907 16469 6941
rect 16527 6907 16561 6941
rect 16619 6907 16653 6941
rect 16711 6907 16745 6941
rect 16803 6907 16837 6941
rect 16895 6907 16929 6941
rect 16987 6907 17021 6941
rect 17079 6907 17113 6941
rect 17171 6907 17205 6941
rect 17263 6907 17297 6941
rect 17355 6907 17389 6941
rect 17447 6907 17481 6941
rect 17539 6907 17573 6941
rect 17631 6907 17665 6941
rect 17723 6907 17757 6941
rect 17815 6907 17849 6941
rect 17907 6907 17941 6941
rect 17999 6907 18033 6941
rect 18091 6907 18125 6941
rect 13492 6737 13526 6771
rect 13411 6671 13445 6705
rect 13584 6533 13618 6567
rect 13860 6737 13894 6771
rect 13741 6631 13775 6635
rect 13741 6601 13754 6631
rect 13754 6601 13775 6631
rect 13948 6549 13966 6567
rect 13966 6549 13982 6567
rect 13948 6533 13982 6549
rect 14596 6745 14630 6771
rect 14596 6737 14617 6745
rect 14617 6737 14630 6745
rect 14504 6669 14538 6703
rect 14136 6559 14138 6567
rect 14138 6559 14170 6567
rect 14136 6533 14170 6559
rect 14596 6601 14630 6635
rect 14872 6559 14881 6567
rect 14881 6559 14906 6567
rect 14872 6533 14906 6559
rect 15148 6669 15182 6703
rect 15256 6599 15258 6633
rect 15258 6599 15290 6633
rect 15702 6829 15736 6831
rect 15702 6797 15727 6829
rect 15727 6797 15736 6829
rect 15884 6737 15918 6771
rect 15806 6644 15840 6662
rect 15806 6628 15828 6644
rect 15828 6628 15840 6644
rect 15976 6533 16010 6567
rect 16252 6737 16286 6771
rect 16139 6631 16173 6634
rect 16139 6600 16146 6631
rect 16146 6600 16173 6631
rect 16340 6549 16358 6567
rect 16358 6549 16374 6567
rect 16340 6533 16374 6549
rect 16988 6745 17022 6771
rect 16988 6737 17009 6745
rect 17009 6737 17022 6745
rect 16896 6669 16930 6703
rect 16528 6559 16530 6567
rect 16530 6559 16562 6567
rect 16528 6533 16562 6559
rect 16988 6601 17022 6635
rect 17264 6559 17273 6567
rect 17273 6559 17298 6567
rect 17264 6533 17298 6559
rect 17540 6669 17574 6703
rect 17649 6633 17683 6634
rect 17649 6600 17650 6633
rect 17650 6600 17683 6633
rect 18092 6475 18119 6502
rect 18119 6475 18126 6502
rect 18092 6468 18126 6475
rect 13399 6363 13433 6397
rect 13491 6363 13525 6397
rect 13583 6363 13617 6397
rect 13675 6363 13709 6397
rect 13767 6363 13801 6397
rect 13859 6363 13893 6397
rect 13951 6363 13985 6397
rect 14043 6363 14077 6397
rect 14135 6363 14169 6397
rect 14227 6363 14261 6397
rect 14319 6363 14353 6397
rect 14411 6363 14445 6397
rect 14503 6363 14537 6397
rect 14595 6363 14629 6397
rect 14687 6363 14721 6397
rect 14779 6363 14813 6397
rect 14871 6363 14905 6397
rect 14963 6363 14997 6397
rect 15055 6363 15089 6397
rect 15147 6363 15181 6397
rect 15239 6363 15273 6397
rect 15331 6363 15365 6397
rect 15423 6363 15457 6397
rect 15515 6363 15549 6397
rect 15607 6363 15641 6397
rect 15699 6363 15733 6397
rect 15791 6363 15825 6397
rect 15883 6363 15917 6397
rect 15975 6363 16009 6397
rect 16067 6363 16101 6397
rect 16159 6363 16193 6397
rect 16251 6363 16285 6397
rect 16343 6363 16377 6397
rect 16435 6363 16469 6397
rect 16527 6363 16561 6397
rect 16619 6363 16653 6397
rect 16711 6363 16745 6397
rect 16803 6363 16837 6397
rect 16895 6363 16929 6397
rect 16987 6363 17021 6397
rect 17079 6363 17113 6397
rect 17171 6363 17205 6397
rect 17263 6363 17297 6397
rect 17355 6363 17389 6397
rect 17447 6363 17481 6397
rect 17539 6363 17573 6397
rect 17631 6363 17665 6397
rect 17723 6363 17757 6397
rect 17815 6363 17849 6397
rect 17907 6363 17941 6397
rect 17999 6363 18033 6397
rect 18091 6363 18125 6397
rect 13399 6267 13433 6301
rect 13491 6267 13525 6301
rect 13583 6267 13617 6301
rect 13675 6267 13709 6301
rect 13767 6267 13801 6301
rect 13859 6267 13893 6301
rect 13951 6267 13985 6301
rect 14043 6267 14077 6301
rect 14135 6267 14169 6301
rect 14227 6267 14261 6301
rect 14319 6267 14353 6301
rect 14411 6267 14445 6301
rect 14503 6267 14537 6301
rect 14595 6267 14629 6301
rect 14687 6267 14721 6301
rect 14779 6267 14813 6301
rect 14871 6267 14905 6301
rect 14963 6267 14997 6301
rect 15055 6267 15089 6301
rect 15147 6267 15181 6301
rect 15239 6267 15273 6301
rect 15331 6267 15365 6301
rect 15423 6267 15457 6301
rect 15515 6267 15549 6301
rect 15607 6267 15641 6301
rect 15699 6267 15733 6301
rect 15791 6267 15825 6301
rect 15883 6267 15917 6301
rect 15975 6267 16009 6301
rect 16067 6267 16101 6301
rect 16159 6267 16193 6301
rect 16251 6267 16285 6301
rect 16343 6267 16377 6301
rect 16435 6267 16469 6301
rect 16527 6267 16561 6301
rect 16619 6267 16653 6301
rect 16711 6267 16745 6301
rect 16803 6267 16837 6301
rect 16895 6267 16929 6301
rect 16987 6267 17021 6301
rect 17079 6267 17113 6301
rect 17171 6267 17205 6301
rect 17263 6267 17297 6301
rect 17355 6267 17389 6301
rect 17447 6267 17481 6301
rect 17539 6267 17573 6301
rect 17631 6267 17665 6301
rect 17723 6267 17757 6301
rect 17815 6267 17849 6301
rect 17907 6267 17941 6301
rect 17999 6267 18033 6301
rect 18091 6267 18125 6301
rect 13419 6055 13453 6089
rect 13492 5893 13526 5927
rect 13584 6097 13618 6131
rect 13746 5971 13780 6005
rect 13948 6115 13982 6131
rect 13948 6097 13966 6115
rect 13966 6097 13982 6115
rect 14136 6105 14170 6131
rect 14136 6097 14138 6105
rect 14138 6097 14170 6105
rect 13860 5893 13894 5927
rect 14596 6029 14630 6063
rect 14504 5961 14538 5995
rect 14596 5919 14617 5927
rect 14617 5919 14630 5927
rect 14596 5893 14630 5919
rect 14872 6105 14906 6131
rect 14872 6097 14881 6105
rect 14881 6097 14906 6105
rect 15265 6031 15292 6063
rect 15292 6031 15299 6063
rect 15265 6029 15299 6031
rect 15148 5961 15182 5995
rect 15803 6020 15828 6045
rect 15828 6020 15837 6045
rect 15803 6011 15837 6020
rect 15699 5835 15727 5868
rect 15727 5835 15733 5868
rect 15699 5834 15733 5835
rect 15884 5893 15918 5927
rect 15976 6097 16010 6131
rect 16140 6033 16146 6062
rect 16146 6033 16174 6062
rect 16140 6028 16174 6033
rect 16340 6115 16374 6131
rect 16340 6097 16358 6115
rect 16358 6097 16374 6115
rect 16528 6105 16562 6131
rect 16528 6097 16530 6105
rect 16530 6097 16562 6105
rect 16252 5893 16286 5927
rect 16988 6029 17022 6063
rect 16896 5961 16930 5995
rect 16988 5919 17009 5927
rect 17009 5919 17022 5927
rect 16988 5893 17022 5919
rect 17264 6105 17298 6131
rect 17264 6097 17273 6105
rect 17273 6097 17298 6105
rect 17649 6031 17650 6065
rect 17650 6031 17683 6065
rect 17540 5961 17574 5995
rect 18086 6155 18119 6179
rect 18119 6155 18120 6179
rect 18086 6145 18120 6155
rect 13399 5723 13433 5757
rect 13491 5723 13525 5757
rect 13583 5723 13617 5757
rect 13675 5723 13709 5757
rect 13767 5723 13801 5757
rect 13859 5723 13893 5757
rect 13951 5723 13985 5757
rect 14043 5723 14077 5757
rect 14135 5723 14169 5757
rect 14227 5723 14261 5757
rect 14319 5723 14353 5757
rect 14411 5723 14445 5757
rect 14503 5723 14537 5757
rect 14595 5723 14629 5757
rect 14687 5723 14721 5757
rect 14779 5723 14813 5757
rect 14871 5723 14905 5757
rect 14963 5723 14997 5757
rect 15055 5723 15089 5757
rect 15147 5723 15181 5757
rect 15239 5723 15273 5757
rect 15331 5723 15365 5757
rect 15423 5723 15457 5757
rect 15515 5723 15549 5757
rect 15607 5723 15641 5757
rect 15699 5723 15733 5757
rect 15791 5723 15825 5757
rect 15883 5723 15917 5757
rect 15975 5723 16009 5757
rect 16067 5723 16101 5757
rect 16159 5723 16193 5757
rect 16251 5723 16285 5757
rect 16343 5723 16377 5757
rect 16435 5723 16469 5757
rect 16527 5723 16561 5757
rect 16619 5723 16653 5757
rect 16711 5723 16745 5757
rect 16803 5723 16837 5757
rect 16895 5723 16929 5757
rect 16987 5723 17021 5757
rect 17079 5723 17113 5757
rect 17171 5723 17205 5757
rect 17263 5723 17297 5757
rect 17355 5723 17389 5757
rect 17447 5723 17481 5757
rect 17539 5723 17573 5757
rect 17631 5723 17665 5757
rect 17723 5723 17757 5757
rect 17815 5723 17849 5757
rect 17907 5723 17941 5757
rect 17999 5723 18033 5757
rect 18091 5723 18125 5757
rect 13399 5627 13433 5661
rect 13491 5627 13525 5661
rect 13583 5627 13617 5661
rect 13675 5627 13709 5661
rect 13767 5627 13801 5661
rect 13859 5627 13893 5661
rect 13951 5627 13985 5661
rect 14043 5627 14077 5661
rect 14135 5627 14169 5661
rect 14227 5627 14261 5661
rect 14319 5627 14353 5661
rect 14411 5627 14445 5661
rect 14503 5627 14537 5661
rect 14595 5627 14629 5661
rect 14687 5627 14721 5661
rect 14779 5627 14813 5661
rect 14871 5627 14905 5661
rect 14963 5627 14997 5661
rect 15055 5627 15089 5661
rect 15147 5627 15181 5661
rect 15239 5627 15273 5661
rect 15331 5627 15365 5661
rect 15423 5627 15457 5661
rect 15515 5627 15549 5661
rect 15607 5627 15641 5661
rect 15699 5627 15733 5661
rect 15791 5627 15825 5661
rect 15883 5627 15917 5661
rect 15975 5627 16009 5661
rect 16067 5627 16101 5661
rect 16159 5627 16193 5661
rect 16251 5627 16285 5661
rect 16343 5627 16377 5661
rect 16435 5627 16469 5661
rect 16527 5627 16561 5661
rect 16619 5627 16653 5661
rect 16711 5627 16745 5661
rect 16803 5627 16837 5661
rect 16895 5627 16929 5661
rect 16987 5627 17021 5661
rect 17079 5627 17113 5661
rect 17171 5627 17205 5661
rect 17263 5627 17297 5661
rect 17355 5627 17389 5661
rect 17447 5627 17481 5661
rect 17539 5627 17573 5661
rect 17631 5627 17665 5661
rect 17723 5627 17757 5661
rect 17815 5627 17849 5661
rect 17907 5627 17941 5661
rect 17999 5627 18033 5661
rect 18091 5627 18125 5661
rect 13492 5457 13526 5491
rect 13415 5295 13449 5329
rect 13584 5253 13618 5287
rect 13860 5457 13894 5491
rect 13743 5379 13777 5413
rect 13948 5269 13966 5287
rect 13966 5269 13982 5287
rect 13948 5253 13982 5269
rect 14596 5465 14630 5491
rect 14596 5457 14617 5465
rect 14617 5457 14630 5465
rect 14504 5389 14538 5423
rect 14136 5279 14138 5287
rect 14138 5279 14170 5287
rect 14136 5253 14170 5279
rect 14596 5321 14630 5355
rect 14872 5279 14881 5287
rect 14881 5279 14906 5287
rect 14872 5253 14906 5279
rect 15148 5389 15182 5423
rect 15257 5319 15258 5353
rect 15258 5319 15291 5353
rect 15699 5549 15733 5553
rect 15699 5519 15727 5549
rect 15727 5519 15733 5549
rect 15884 5457 15918 5491
rect 15804 5330 15828 5359
rect 15828 5330 15838 5359
rect 15804 5325 15838 5330
rect 15976 5253 16010 5287
rect 16252 5457 16286 5491
rect 16141 5351 16175 5354
rect 16141 5320 16146 5351
rect 16146 5320 16175 5351
rect 16340 5269 16358 5287
rect 16358 5269 16374 5287
rect 16340 5253 16374 5269
rect 16988 5465 17022 5491
rect 16988 5457 17009 5465
rect 17009 5457 17022 5465
rect 16896 5389 16930 5423
rect 16528 5279 16530 5287
rect 16530 5279 16562 5287
rect 16528 5253 16562 5279
rect 16988 5321 17022 5355
rect 17264 5279 17273 5287
rect 17273 5279 17298 5287
rect 17264 5253 17298 5279
rect 17540 5389 17574 5423
rect 17649 5353 17683 5354
rect 17649 5320 17650 5353
rect 17650 5320 17683 5353
rect 18087 5195 18119 5220
rect 18119 5195 18121 5220
rect 18087 5186 18121 5195
rect 13399 5083 13433 5117
rect 13491 5083 13525 5117
rect 13583 5083 13617 5117
rect 13675 5083 13709 5117
rect 13767 5083 13801 5117
rect 13859 5083 13893 5117
rect 13951 5083 13985 5117
rect 14043 5083 14077 5117
rect 14135 5083 14169 5117
rect 14227 5083 14261 5117
rect 14319 5083 14353 5117
rect 14411 5083 14445 5117
rect 14503 5083 14537 5117
rect 14595 5083 14629 5117
rect 14687 5083 14721 5117
rect 14779 5083 14813 5117
rect 14871 5083 14905 5117
rect 14963 5083 14997 5117
rect 15055 5083 15089 5117
rect 15147 5083 15181 5117
rect 15239 5083 15273 5117
rect 15331 5083 15365 5117
rect 15423 5083 15457 5117
rect 15515 5083 15549 5117
rect 15607 5083 15641 5117
rect 15699 5083 15733 5117
rect 15791 5083 15825 5117
rect 15883 5083 15917 5117
rect 15975 5083 16009 5117
rect 16067 5083 16101 5117
rect 16159 5083 16193 5117
rect 16251 5083 16285 5117
rect 16343 5083 16377 5117
rect 16435 5083 16469 5117
rect 16527 5083 16561 5117
rect 16619 5083 16653 5117
rect 16711 5083 16745 5117
rect 16803 5083 16837 5117
rect 16895 5083 16929 5117
rect 16987 5083 17021 5117
rect 17079 5083 17113 5117
rect 17171 5083 17205 5117
rect 17263 5083 17297 5117
rect 17355 5083 17389 5117
rect 17447 5083 17481 5117
rect 17539 5083 17573 5117
rect 17631 5083 17665 5117
rect 17723 5083 17757 5117
rect 17815 5083 17849 5117
rect 17907 5083 17941 5117
rect 17999 5083 18033 5117
rect 18091 5083 18125 5117
<< metal1 >>
rect 12455 10612 12545 10628
rect 12455 10601 12474 10612
rect 12437 10579 12474 10601
rect 12328 10567 12374 10579
rect 12328 10507 12334 10567
rect 12368 10507 12374 10567
rect 12328 10429 12374 10507
rect 12416 10567 12474 10579
rect 12416 10507 12422 10567
rect 12456 10560 12474 10567
rect 12526 10609 12545 10612
rect 12526 10603 13134 10609
rect 12526 10560 12572 10603
rect 12456 10551 12572 10560
rect 12624 10551 12652 10603
rect 12704 10551 12732 10603
rect 12784 10551 12812 10603
rect 12864 10551 12892 10603
rect 12944 10551 12972 10603
rect 13024 10551 13134 10603
rect 12456 10543 13134 10551
rect 13196 10606 18104 10612
rect 13196 10554 13304 10606
rect 13356 10554 13384 10606
rect 13436 10554 13464 10606
rect 13516 10554 13544 10606
rect 13596 10554 13624 10606
rect 13676 10554 13704 10606
rect 13756 10554 13908 10606
rect 13960 10554 13988 10606
rect 14040 10554 14068 10606
rect 14120 10554 14148 10606
rect 14200 10554 14228 10606
rect 14280 10554 14308 10606
rect 14360 10554 14516 10606
rect 14568 10554 14596 10606
rect 14648 10554 14676 10606
rect 14728 10554 14756 10606
rect 14808 10554 14836 10606
rect 14888 10554 14916 10606
rect 14968 10554 15120 10606
rect 15172 10554 15200 10606
rect 15252 10554 15280 10606
rect 15332 10554 15360 10606
rect 15412 10554 15440 10606
rect 15492 10554 15520 10606
rect 15572 10554 15728 10606
rect 15780 10554 15808 10606
rect 15860 10554 15888 10606
rect 15940 10554 15968 10606
rect 16020 10554 16048 10606
rect 16100 10554 16128 10606
rect 16180 10554 16332 10606
rect 16384 10554 16412 10606
rect 16464 10554 16492 10606
rect 16544 10554 16572 10606
rect 16624 10554 16652 10606
rect 16704 10554 16732 10606
rect 16784 10554 16940 10606
rect 16992 10554 17020 10606
rect 17072 10554 17100 10606
rect 17152 10554 17180 10606
rect 17232 10554 17260 10606
rect 17312 10554 17340 10606
rect 17392 10554 17544 10606
rect 17596 10554 17624 10606
rect 17676 10554 17704 10606
rect 17756 10554 17784 10606
rect 17836 10554 17864 10606
rect 17916 10554 17944 10606
rect 17996 10554 18104 10606
rect 13196 10546 18104 10554
rect 18264 10550 18354 10566
rect 12456 10513 12490 10543
rect 12456 10507 12462 10513
rect 12416 10495 12462 10507
rect 18264 10498 18283 10550
rect 18335 10498 18354 10550
rect 18264 10482 18354 10498
rect 12328 10369 12334 10429
rect 12368 10369 12374 10429
rect 12328 10357 12374 10369
rect 12416 10429 12462 10441
rect 12416 10369 12422 10429
rect 12456 10369 12462 10429
rect 12328 10291 12374 10303
rect 12328 10231 12334 10291
rect 12368 10231 12374 10291
rect 12328 10153 12374 10231
rect 12416 10291 12462 10369
rect 18269 10406 18359 10422
rect 18269 10354 18288 10406
rect 18340 10354 18359 10406
rect 18269 10338 18359 10354
rect 12416 10231 12422 10291
rect 12456 10231 12462 10291
rect 12416 10219 12462 10231
rect 18270 10254 18360 10270
rect 18270 10202 18289 10254
rect 18341 10202 18360 10254
rect 18270 10186 18360 10202
rect 12328 10093 12334 10153
rect 12368 10093 12374 10153
rect 12328 10081 12374 10093
rect 12416 10153 12462 10165
rect 12416 10093 12422 10153
rect 12456 10093 12462 10153
rect 11792 10007 12252 10027
rect 11792 9996 11857 10007
rect 11792 9962 11821 9996
rect 11855 9962 11857 9996
rect 11792 9955 11857 9962
rect 11909 10006 12132 10007
rect 11909 9996 11988 10006
rect 12040 9996 12132 10006
rect 11909 9962 11913 9996
rect 11947 9962 11988 9996
rect 12040 9962 12097 9996
rect 12131 9962 12132 9996
rect 11909 9955 11988 9962
rect 11792 9954 11988 9955
rect 12040 9955 12132 9962
rect 12184 9996 12252 10007
rect 12184 9962 12189 9996
rect 12223 9962 12252 9996
rect 12184 9955 12252 9962
rect 12040 9954 12252 9955
rect 11792 9931 12252 9954
rect 12328 10015 12374 10027
rect 12328 9955 12334 10015
rect 12368 9955 12374 10015
rect 12328 9877 12374 9955
rect 12416 10015 12462 10093
rect 18270 10084 18360 10100
rect 18270 10032 18289 10084
rect 18341 10032 18360 10084
rect 18270 10016 18360 10032
rect 12416 9955 12422 10015
rect 12456 9955 12462 10015
rect 12416 9943 12462 9955
rect 18269 9927 18359 9943
rect 11937 9853 12300 9860
rect 11937 9819 11949 9853
rect 11983 9832 12300 9853
rect 11983 9819 11995 9832
rect 11937 9812 11995 9819
rect 12042 9798 12109 9804
rect 12042 9764 12058 9798
rect 12092 9785 12109 9798
rect 12092 9764 12244 9785
rect 12042 9757 12244 9764
rect 12122 9696 12188 9698
rect 11860 9691 11914 9695
rect 11859 9688 11914 9691
rect 11730 9654 11868 9688
rect 11902 9654 11914 9688
rect 11859 9651 11914 9654
rect 11859 9647 11913 9651
rect 12122 9644 12130 9696
rect 12182 9644 12188 9696
rect 12122 9643 12188 9644
rect 12216 9613 12244 9757
rect 12272 9700 12300 9832
rect 12328 9817 12334 9877
rect 12368 9817 12374 9877
rect 12328 9805 12374 9817
rect 12416 9877 12519 9889
rect 12416 9817 12422 9877
rect 12456 9817 12519 9877
rect 18269 9875 18288 9927
rect 18340 9875 18359 9927
rect 18269 9859 18359 9875
rect 12416 9805 12519 9817
rect 12366 9758 12435 9764
rect 12366 9724 12378 9758
rect 12412 9724 12435 9758
rect 12366 9718 12435 9724
rect 12272 9688 12321 9700
rect 12272 9654 12281 9688
rect 12315 9654 12321 9688
rect 12272 9641 12321 9654
rect 12216 9595 12359 9613
rect 12216 9585 12319 9595
rect 12310 9561 12319 9585
rect 12353 9561 12359 9595
rect 12310 9548 12359 9561
rect 11792 9461 12252 9483
rect 11792 9452 11875 9461
rect 11927 9452 11995 9461
rect 12047 9452 12138 9461
rect 12190 9452 12252 9461
rect 11792 9418 11821 9452
rect 11855 9418 11875 9452
rect 11947 9418 11995 9452
rect 12047 9418 12097 9452
rect 12131 9418 12138 9452
rect 12223 9418 12252 9452
rect 11792 9409 11875 9418
rect 11927 9409 11995 9418
rect 12047 9409 12138 9418
rect 12190 9409 12252 9418
rect 11792 9387 12252 9409
rect 12387 9318 12435 9718
rect 11767 9271 12435 9318
rect 12387 9130 12435 9271
rect 12377 9124 12435 9130
rect 12136 9118 12201 9119
rect 12136 9117 12142 9118
rect 12030 9069 12142 9117
rect 12136 9066 12142 9069
rect 12194 9066 12201 9118
rect 12377 9090 12389 9124
rect 12423 9090 12435 9124
rect 12377 9084 12435 9090
rect 12473 9315 12519 9805
rect 18187 9685 18277 9701
rect 18187 9674 18206 9685
rect 18112 9633 18206 9674
rect 18258 9633 18277 9685
rect 18564 9693 18654 9709
rect 18564 9682 18583 9693
rect 18545 9650 18583 9682
rect 12569 9618 12618 9625
rect 12569 9613 13188 9618
rect 12569 9579 12578 9613
rect 12612 9579 13188 9613
rect 12569 9571 13188 9579
rect 12569 9566 12618 9571
rect 12570 9524 12619 9532
rect 13139 9524 13188 9571
rect 18112 9615 18277 9633
rect 18472 9641 18583 9650
rect 18635 9650 18654 9693
rect 18764 9693 18854 9709
rect 18764 9682 18783 9693
rect 18745 9650 18783 9682
rect 18635 9641 18783 9650
rect 18835 9641 18854 9693
rect 18472 9623 18854 9641
rect 18472 9619 18840 9623
rect 18112 9569 18159 9615
rect 18472 9585 18501 9619
rect 18535 9585 18593 9619
rect 18627 9585 18685 9619
rect 18719 9585 18777 9619
rect 18811 9585 18840 9619
rect 18113 9566 18159 9569
rect 12570 9520 13071 9524
rect 12570 9486 12579 9520
rect 12613 9515 13071 9520
rect 12613 9486 13020 9515
rect 12570 9481 13020 9486
rect 13054 9481 13071 9515
rect 12570 9478 13071 9481
rect 13139 9518 17560 9524
rect 13139 9484 13752 9518
rect 13786 9484 13878 9518
rect 13912 9484 14964 9518
rect 14998 9484 15090 9518
rect 15124 9484 16176 9518
rect 16210 9484 16302 9518
rect 16336 9484 17388 9518
rect 17422 9484 17514 9518
rect 17548 9484 17560 9518
rect 18113 9506 18119 9566
rect 18153 9506 18159 9566
rect 18113 9494 18159 9506
rect 18201 9566 18247 9578
rect 18201 9506 18207 9566
rect 18241 9506 18247 9566
rect 18472 9554 18840 9585
rect 18201 9497 18247 9506
rect 13139 9478 17560 9484
rect 12570 9477 13066 9478
rect 13139 9477 13585 9478
rect 12570 9473 12619 9477
rect 13008 9475 13066 9477
rect 18201 9468 18439 9497
rect 12970 9426 13016 9434
rect 12947 9425 13026 9426
rect 12947 9361 12954 9425
rect 13018 9361 13026 9425
rect 13058 9425 13104 9437
rect 13702 9429 13748 9437
rect 13058 9365 13064 9425
rect 13098 9365 13104 9425
rect 12970 9350 13016 9361
rect 13058 9315 13104 9365
rect 13679 9428 13758 9429
rect 13679 9364 13686 9428
rect 13750 9364 13758 9428
rect 13807 9425 13853 9437
rect 13916 9429 13962 9437
rect 14914 9429 14960 9437
rect 13807 9365 13813 9425
rect 13847 9365 13853 9425
rect 13702 9353 13748 9364
rect 13807 9315 13853 9365
rect 13906 9428 13985 9429
rect 13906 9364 13914 9428
rect 13978 9364 13985 9428
rect 14891 9428 14970 9429
rect 14891 9364 14898 9428
rect 14962 9364 14970 9428
rect 15018 9425 15064 9437
rect 15128 9429 15174 9437
rect 16126 9429 16172 9437
rect 15018 9365 15024 9425
rect 15058 9365 15064 9425
rect 13916 9353 13962 9364
rect 14914 9353 14960 9364
rect 15018 9315 15064 9365
rect 15118 9428 15197 9429
rect 15118 9364 15126 9428
rect 15190 9364 15197 9428
rect 16103 9428 16182 9429
rect 16103 9364 16110 9428
rect 16174 9364 16182 9428
rect 16231 9425 16277 9437
rect 16340 9429 16386 9437
rect 17338 9429 17384 9437
rect 16231 9365 16237 9425
rect 16271 9365 16277 9425
rect 15128 9353 15174 9364
rect 16126 9353 16172 9364
rect 16231 9315 16277 9365
rect 16330 9428 16409 9429
rect 16330 9364 16338 9428
rect 16402 9364 16409 9428
rect 17315 9428 17394 9429
rect 17315 9364 17322 9428
rect 17386 9364 17394 9428
rect 17445 9425 17491 9437
rect 17552 9429 17598 9437
rect 17445 9365 17451 9425
rect 17485 9365 17491 9425
rect 16340 9353 16386 9364
rect 17338 9353 17384 9364
rect 17445 9315 17491 9365
rect 17542 9428 17621 9429
rect 17542 9364 17550 9428
rect 17614 9364 17621 9428
rect 18113 9428 18159 9440
rect 18113 9368 18119 9428
rect 18153 9368 18159 9428
rect 17552 9353 17598 9364
rect 18113 9356 18159 9368
rect 18201 9428 18247 9468
rect 18201 9368 18207 9428
rect 18241 9368 18247 9428
rect 18201 9356 18247 9368
rect 18275 9428 18365 9440
rect 18275 9424 18303 9428
rect 18337 9424 18365 9428
rect 18275 9372 18294 9424
rect 18346 9372 18365 9424
rect 18275 9368 18303 9372
rect 18337 9368 18365 9372
rect 18275 9356 18365 9368
rect 18393 9428 18439 9468
rect 18393 9368 18399 9428
rect 18433 9368 18439 9428
rect 18393 9356 18439 9368
rect 18032 9315 18098 9317
rect 12473 9311 18098 9315
rect 12473 9277 18048 9311
rect 18082 9277 18098 9311
rect 12473 9273 18098 9277
rect 12473 9052 12519 9273
rect 13323 9226 13369 9236
rect 13301 9162 13310 9226
rect 13374 9162 13383 9226
rect 13301 9161 13383 9162
rect 13413 9224 13459 9273
rect 14055 9226 14101 9236
rect 13413 9164 13419 9224
rect 13453 9164 13459 9224
rect 13323 9152 13369 9161
rect 13413 9152 13459 9164
rect 14033 9162 14042 9226
rect 14106 9162 14115 9226
rect 14033 9161 14115 9162
rect 14162 9224 14208 9273
rect 14265 9226 14311 9236
rect 15267 9226 15313 9236
rect 14162 9164 14168 9224
rect 14202 9164 14208 9224
rect 14055 9152 14101 9161
rect 14162 9152 14208 9164
rect 14251 9162 14260 9226
rect 14324 9162 14333 9226
rect 14251 9161 14333 9162
rect 15245 9162 15254 9226
rect 15318 9162 15327 9226
rect 15245 9161 15327 9162
rect 15373 9224 15419 9273
rect 15477 9226 15523 9236
rect 16605 9226 16651 9236
rect 15373 9164 15379 9224
rect 15413 9164 15419 9224
rect 14265 9152 14311 9161
rect 15267 9152 15313 9161
rect 15373 9152 15419 9164
rect 15463 9162 15472 9226
rect 15536 9162 15545 9226
rect 15463 9161 15545 9162
rect 16583 9162 16592 9226
rect 16656 9162 16665 9226
rect 16583 9161 16665 9162
rect 16713 9224 16759 9273
rect 16815 9226 16861 9236
rect 16713 9164 16719 9224
rect 16753 9164 16759 9224
rect 15477 9152 15523 9161
rect 16605 9152 16651 9161
rect 16713 9152 16759 9164
rect 16801 9162 16810 9226
rect 16874 9162 16883 9226
rect 16801 9161 16883 9162
rect 17460 9224 17506 9273
rect 18036 9271 18098 9273
rect 18131 9308 18159 9356
rect 18243 9309 18542 9315
rect 18243 9308 18255 9309
rect 18131 9279 18255 9308
rect 18131 9237 18159 9279
rect 18243 9275 18255 9279
rect 18289 9275 18495 9309
rect 18529 9275 18542 9309
rect 18243 9269 18542 9275
rect 18690 9309 18748 9315
rect 18690 9275 18702 9309
rect 18736 9306 18748 9309
rect 18736 9278 18897 9306
rect 18736 9275 18748 9278
rect 18690 9269 18748 9275
rect 17549 9226 17595 9236
rect 17460 9164 17466 9224
rect 17500 9164 17506 9224
rect 16815 9152 16861 9161
rect 17460 9152 17506 9164
rect 17535 9162 17544 9226
rect 17608 9162 17617 9226
rect 17535 9161 17617 9162
rect 18113 9225 18159 9237
rect 18113 9165 18119 9225
rect 18153 9165 18159 9225
rect 17549 9152 17595 9161
rect 18113 9153 18159 9165
rect 18201 9225 18247 9237
rect 18201 9165 18207 9225
rect 18241 9165 18247 9225
rect 18201 9125 18247 9165
rect 18275 9225 18365 9237
rect 18275 9221 18303 9225
rect 18337 9221 18365 9225
rect 18275 9169 18294 9221
rect 18346 9169 18365 9221
rect 18275 9165 18303 9169
rect 18337 9165 18365 9169
rect 18275 9153 18365 9165
rect 18393 9225 18439 9237
rect 18393 9165 18399 9225
rect 18433 9165 18439 9225
rect 18393 9125 18439 9165
rect 17501 9120 17560 9123
rect 12623 9066 12630 9118
rect 12682 9116 12688 9118
rect 13361 9116 13419 9120
rect 12682 9114 13419 9116
rect 12682 9080 13373 9114
rect 13407 9099 13419 9114
rect 14093 9114 15489 9120
rect 13407 9080 13421 9099
rect 12682 9069 13421 9080
rect 14093 9080 14105 9114
rect 14139 9080 14227 9114
rect 14261 9080 15317 9114
rect 15351 9080 15439 9114
rect 15473 9080 15489 9114
rect 14093 9074 15489 9080
rect 16643 9114 16827 9120
rect 16643 9080 16655 9114
rect 16689 9080 16777 9114
rect 16811 9080 16827 9114
rect 16643 9074 16827 9080
rect 17499 9114 17560 9120
rect 17499 9080 17511 9114
rect 17545 9080 17560 9114
rect 17499 9074 17560 9080
rect 12682 9066 12688 9069
rect 12623 9065 12688 9066
rect 13363 9064 13421 9069
rect 12303 9040 12349 9052
rect 12303 8980 12309 9040
rect 12343 8980 12349 9040
rect 12303 8902 12349 8980
rect 12463 9040 12519 9052
rect 12463 8980 12469 9040
rect 12503 8980 12519 9040
rect 12463 8968 12519 8980
rect 12303 8842 12309 8902
rect 12343 8842 12349 8902
rect 12303 8830 12349 8842
rect 12463 8902 12509 8914
rect 12463 8842 12469 8902
rect 12503 8842 12509 8902
rect 12303 8764 12349 8776
rect 12303 8704 12309 8764
rect 12343 8704 12349 8764
rect 12303 8626 12349 8704
rect 12463 8764 12509 8842
rect 12463 8704 12469 8764
rect 12503 8704 12509 8764
rect 12463 8692 12509 8704
rect 12303 8566 12309 8626
rect 12343 8566 12349 8626
rect 12303 8554 12349 8566
rect 12463 8626 12509 8638
rect 12463 8566 12469 8626
rect 12503 8566 12509 8626
rect 12303 8488 12349 8500
rect 12303 8428 12309 8488
rect 12343 8428 12349 8488
rect 12303 8350 12349 8428
rect 12463 8488 12509 8566
rect 12463 8428 12469 8488
rect 12503 8428 12509 8488
rect 12463 8416 12509 8428
rect 12303 8290 12309 8350
rect 12343 8290 12349 8350
rect 12303 8278 12349 8290
rect 12463 8350 12509 8362
rect 12463 8290 12469 8350
rect 12503 8290 12509 8350
rect 12303 8212 12349 8224
rect 12303 8152 12309 8212
rect 12343 8152 12349 8212
rect 12303 8074 12349 8152
rect 12463 8212 12509 8290
rect 12463 8152 12469 8212
rect 12503 8152 12509 8212
rect 12463 8140 12509 8152
rect 12303 8014 12309 8074
rect 12343 8014 12349 8074
rect 12463 8074 12509 8086
rect 12463 8050 12469 8074
rect 12303 8002 12349 8014
rect 12424 8034 12469 8050
rect 12503 8050 12509 8074
rect 12503 8034 12531 8050
rect 12424 7982 12460 8034
rect 12512 7982 12531 8034
rect 12424 7966 12531 7982
rect 12984 8037 13316 8043
rect 12984 7985 13002 8037
rect 13054 7985 13082 8037
rect 13134 7985 13162 8037
rect 13214 7985 13242 8037
rect 13294 7985 13316 8037
rect 12984 7975 13316 7985
rect 13716 8037 14048 8043
rect 13716 7985 13734 8037
rect 13786 7985 13814 8037
rect 13866 7985 13894 8037
rect 13946 7985 13974 8037
rect 14026 7985 14048 8037
rect 13716 7975 14048 7985
rect 14219 7946 14277 9074
rect 14318 8037 14650 8043
rect 14318 7985 14340 8037
rect 14392 7985 14420 8037
rect 14472 7985 14500 8037
rect 14552 7985 14580 8037
rect 14632 7985 14650 8037
rect 14318 7975 14650 7985
rect 14928 8037 15260 8043
rect 14928 7985 14946 8037
rect 14998 7985 15026 8037
rect 15078 7985 15106 8037
rect 15158 7985 15186 8037
rect 15238 7985 15260 8037
rect 14928 7975 15260 7985
rect 15530 8037 15862 8043
rect 15530 7985 15552 8037
rect 15604 7985 15632 8037
rect 15684 7985 15712 8037
rect 15764 7985 15792 8037
rect 15844 7985 15862 8037
rect 15530 7975 15862 7985
rect 16266 8037 16598 8043
rect 16266 7985 16284 8037
rect 16336 7985 16364 8037
rect 16416 7985 16444 8037
rect 16496 7985 16524 8037
rect 16576 7985 16598 8037
rect 16266 7975 16598 7985
rect 13338 7918 14277 7946
rect 16645 7890 16703 9074
rect 16868 8037 17200 8043
rect 16868 7985 16890 8037
rect 16942 7985 16970 8037
rect 17022 7985 17050 8037
rect 17102 7985 17130 8037
rect 17182 7985 17200 8037
rect 16868 7975 17200 7985
rect 13338 7862 16703 7890
rect 17501 7834 17560 9074
rect 18113 9087 18159 9099
rect 18113 9027 18119 9087
rect 18153 9027 18159 9087
rect 18113 8975 18159 9027
rect 18201 9096 18439 9125
rect 18201 9087 18247 9096
rect 18201 9027 18207 9087
rect 18241 9027 18247 9087
rect 18472 9075 18840 9106
rect 18472 9067 18501 9075
rect 18201 9015 18247 9027
rect 18358 9051 18501 9067
rect 18358 8999 18394 9051
rect 18446 9041 18501 9051
rect 18535 9041 18593 9075
rect 18627 9041 18685 9075
rect 18719 9041 18777 9075
rect 18811 9067 18840 9075
rect 18811 9041 18841 9067
rect 18446 8999 18841 9041
rect 18358 8983 18841 8999
rect 18113 8959 18274 8975
rect 18113 8907 18203 8959
rect 18255 8907 18274 8959
rect 18113 8891 18274 8907
rect 13338 7806 17560 7834
rect 17602 8037 17934 8043
rect 17602 7985 17624 8037
rect 17676 7985 17704 8037
rect 17756 7985 17784 8037
rect 17836 7985 17864 8037
rect 17916 7985 17934 8037
rect 17602 7778 17934 7985
rect 13285 7750 17934 7778
rect 13285 7612 13339 7750
rect 13409 7655 13415 7707
rect 13467 7695 13473 7707
rect 15803 7695 15809 7707
rect 13467 7667 15809 7695
rect 13467 7655 13473 7667
rect 15803 7655 15809 7667
rect 15861 7695 15867 7707
rect 18869 7695 18897 9278
rect 15861 7667 18897 7695
rect 15861 7655 15867 7667
rect 13491 7612 13525 7615
rect 13583 7612 13617 7615
rect 13675 7612 13709 7615
rect 13767 7612 13801 7615
rect 13859 7612 13893 7615
rect 13951 7612 13985 7615
rect 14043 7612 14077 7615
rect 14135 7612 14169 7615
rect 14226 7612 14260 7615
rect 14319 7612 14353 7615
rect 14411 7612 14445 7615
rect 14503 7612 14537 7615
rect 14595 7612 14629 7615
rect 14687 7612 14721 7615
rect 14779 7612 14813 7615
rect 14871 7612 14905 7615
rect 14963 7612 14997 7615
rect 15055 7612 15089 7615
rect 15147 7612 15181 7615
rect 15239 7612 15273 7615
rect 15331 7612 15365 7615
rect 15423 7612 15457 7615
rect 15515 7612 15549 7615
rect 15607 7612 15641 7615
rect 15699 7612 15733 7615
rect 15791 7612 15825 7615
rect 15883 7612 15917 7615
rect 15975 7612 16009 7615
rect 16067 7612 16101 7615
rect 16159 7612 16193 7615
rect 16251 7612 16285 7615
rect 16343 7612 16377 7615
rect 16435 7612 16469 7615
rect 16527 7612 16561 7615
rect 16619 7612 16653 7615
rect 16711 7612 16745 7615
rect 16803 7612 16837 7615
rect 16895 7612 16929 7615
rect 16987 7612 17021 7615
rect 17079 7612 17113 7615
rect 17171 7612 17205 7615
rect 17263 7612 17297 7615
rect 17355 7612 17389 7615
rect 17447 7612 17481 7615
rect 17539 7612 17573 7615
rect 17631 7612 17665 7615
rect 17723 7612 17757 7615
rect 17815 7612 17849 7615
rect 17907 7612 17941 7615
rect 17999 7612 18033 7615
rect 18091 7612 18125 7615
rect 13285 7596 18154 7612
rect 13285 7595 16903 7596
rect 13285 7592 14539 7595
rect 13285 7590 14107 7592
rect 13285 7589 13906 7590
rect 13285 7581 13507 7589
rect 13559 7588 13906 7589
rect 13559 7581 13681 7588
rect 13733 7581 13906 7588
rect 13958 7581 14107 7590
rect 14159 7590 14539 7592
rect 14159 7581 14330 7590
rect 14382 7581 14539 7590
rect 13285 7547 13399 7581
rect 13433 7547 13491 7581
rect 13559 7547 13583 7581
rect 13617 7547 13675 7581
rect 13733 7547 13767 7581
rect 13801 7547 13859 7581
rect 13893 7547 13906 7581
rect 13985 7547 14043 7581
rect 14077 7547 14107 7581
rect 14169 7547 14227 7581
rect 14261 7547 14319 7581
rect 14382 7547 14411 7581
rect 14445 7547 14503 7581
rect 14537 7547 14539 7581
rect 13285 7537 13507 7547
rect 13559 7537 13681 7547
rect 13285 7536 13681 7537
rect 13733 7538 13906 7547
rect 13958 7540 14107 7547
rect 14159 7540 14330 7547
rect 13958 7538 14330 7540
rect 14382 7543 14539 7547
rect 14591 7592 15162 7595
rect 14591 7588 14957 7592
rect 14591 7581 14767 7588
rect 14819 7581 14957 7588
rect 15009 7581 15162 7592
rect 15214 7581 15361 7595
rect 15413 7590 15965 7595
rect 15413 7581 15577 7590
rect 15629 7581 15965 7590
rect 16017 7593 16903 7595
rect 16017 7592 16674 7593
rect 16017 7590 16442 7592
rect 16017 7581 16200 7590
rect 16252 7581 16442 7590
rect 16494 7581 16674 7592
rect 16726 7581 16903 7593
rect 16955 7595 18154 7596
rect 16955 7592 18036 7595
rect 16955 7588 17370 7592
rect 16955 7581 17152 7588
rect 17204 7581 17370 7588
rect 17422 7590 18036 7592
rect 17422 7588 17820 7590
rect 17422 7581 17599 7588
rect 17651 7581 17820 7588
rect 17872 7581 18036 7590
rect 14591 7547 14595 7581
rect 14629 7547 14687 7581
rect 14721 7547 14767 7581
rect 14819 7547 14871 7581
rect 14905 7547 14957 7581
rect 15009 7547 15055 7581
rect 15089 7547 15147 7581
rect 15214 7547 15239 7581
rect 15273 7547 15331 7581
rect 15413 7547 15423 7581
rect 15457 7547 15515 7581
rect 15549 7547 15577 7581
rect 15641 7547 15699 7581
rect 15733 7547 15791 7581
rect 15825 7547 15883 7581
rect 15917 7547 15965 7581
rect 16017 7547 16067 7581
rect 16101 7547 16159 7581
rect 16193 7547 16200 7581
rect 16285 7547 16343 7581
rect 16377 7547 16435 7581
rect 16494 7547 16527 7581
rect 16561 7547 16619 7581
rect 16653 7547 16674 7581
rect 16745 7547 16803 7581
rect 16837 7547 16895 7581
rect 16955 7547 16987 7581
rect 17021 7547 17079 7581
rect 17113 7547 17152 7581
rect 17205 7547 17263 7581
rect 17297 7547 17355 7581
rect 17422 7547 17447 7581
rect 17481 7547 17539 7581
rect 17573 7547 17599 7581
rect 17665 7547 17723 7581
rect 17757 7547 17815 7581
rect 17872 7547 17907 7581
rect 17941 7547 17999 7581
rect 18033 7547 18036 7581
rect 14591 7543 14767 7547
rect 14382 7538 14767 7543
rect 13733 7536 14767 7538
rect 14819 7540 14957 7547
rect 15009 7543 15162 7547
rect 15214 7543 15361 7547
rect 15413 7543 15577 7547
rect 15009 7540 15577 7543
rect 14819 7538 15577 7540
rect 15629 7543 15965 7547
rect 16017 7543 16200 7547
rect 15629 7538 16200 7543
rect 16252 7540 16442 7547
rect 16494 7541 16674 7547
rect 16726 7544 16903 7547
rect 16955 7544 17152 7547
rect 16726 7541 17152 7544
rect 16494 7540 17152 7541
rect 16252 7538 17152 7540
rect 14819 7536 17152 7538
rect 17204 7540 17370 7547
rect 17422 7540 17599 7547
rect 17204 7536 17599 7540
rect 17651 7538 17820 7547
rect 17872 7543 18036 7547
rect 18088 7581 18154 7595
rect 18088 7547 18091 7581
rect 18125 7547 18154 7581
rect 18088 7543 18154 7547
rect 17872 7538 18154 7543
rect 17651 7536 18154 7538
rect 13285 7516 18154 7536
rect 13289 7476 13334 7486
rect 13289 7448 15907 7476
rect 18207 7466 18252 7476
rect 18078 7460 18252 7466
rect 13289 7438 13334 7448
rect 13572 7411 13630 7417
rect 13572 7377 13584 7411
rect 13618 7408 13630 7411
rect 13936 7411 13994 7417
rect 13936 7408 13948 7411
rect 13618 7380 13948 7408
rect 13618 7377 13630 7380
rect 13572 7371 13630 7377
rect 13936 7377 13948 7380
rect 13982 7377 13994 7411
rect 13936 7371 13994 7377
rect 14124 7411 14182 7417
rect 14124 7377 14136 7411
rect 14170 7408 14182 7411
rect 14860 7411 14918 7417
rect 14860 7408 14872 7411
rect 14170 7402 14872 7408
rect 14906 7402 14918 7411
rect 14170 7380 14865 7402
rect 14170 7377 14182 7380
rect 14124 7371 14182 7377
rect 13406 7364 13458 7370
rect 13955 7340 13994 7371
rect 14858 7350 14865 7380
rect 14917 7350 14924 7402
rect 14584 7343 14642 7349
rect 14584 7340 14596 7343
rect 13955 7312 14596 7340
rect 13406 7306 13458 7312
rect 14584 7309 14596 7312
rect 14630 7309 14642 7343
rect 14584 7303 14642 7309
rect 15243 7299 15250 7351
rect 15302 7299 15309 7351
rect 15878 7342 15906 7448
rect 18078 7426 18091 7460
rect 18125 7437 18252 7460
rect 18125 7426 18137 7437
rect 18207 7428 18252 7437
rect 18078 7420 18137 7426
rect 15964 7411 16022 7417
rect 15964 7377 15976 7411
rect 16010 7408 16022 7411
rect 16328 7411 16386 7417
rect 16328 7408 16340 7411
rect 16010 7380 16340 7408
rect 16010 7377 16022 7380
rect 15964 7371 16022 7377
rect 16328 7377 16340 7380
rect 16374 7377 16386 7411
rect 16328 7371 16386 7377
rect 16516 7411 16574 7417
rect 16516 7377 16528 7411
rect 16562 7408 16574 7411
rect 17252 7411 17310 7417
rect 17252 7408 17264 7411
rect 16562 7401 17264 7408
rect 17298 7401 17310 7411
rect 16562 7380 17260 7401
rect 16562 7377 16574 7380
rect 16516 7371 16574 7377
rect 17252 7371 17260 7380
rect 16120 7343 16187 7352
rect 16120 7342 16138 7343
rect 15798 7322 15850 7328
rect 15878 7314 16138 7342
rect 13721 7281 13782 7287
rect 13297 7269 13342 7280
rect 13721 7269 13736 7281
rect 13297 7247 13736 7269
rect 13770 7247 13782 7281
rect 13297 7241 13782 7247
rect 14492 7275 14550 7281
rect 14492 7241 14504 7275
rect 14538 7272 14550 7275
rect 15136 7275 15194 7281
rect 15136 7272 15148 7275
rect 14538 7244 15148 7272
rect 14538 7241 14550 7244
rect 13297 7232 13342 7241
rect 14492 7235 14550 7241
rect 15136 7241 15148 7244
rect 15182 7241 15194 7275
rect 16120 7309 16138 7314
rect 16172 7309 16187 7343
rect 16347 7340 16386 7371
rect 17253 7349 17260 7371
rect 17312 7349 17319 7401
rect 16976 7343 17034 7349
rect 16976 7340 16988 7343
rect 16347 7312 16988 7340
rect 16120 7301 16187 7309
rect 16976 7309 16988 7312
rect 17022 7309 17034 7343
rect 16976 7303 17034 7309
rect 17638 7300 17645 7352
rect 17697 7300 17704 7352
rect 15798 7264 15850 7270
rect 16884 7275 16942 7281
rect 15136 7235 15194 7241
rect 16884 7241 16896 7275
rect 16930 7272 16942 7275
rect 17528 7275 17586 7281
rect 17528 7272 17540 7275
rect 16930 7244 17540 7272
rect 16930 7241 16942 7244
rect 16884 7235 16942 7241
rect 17528 7241 17540 7244
rect 17574 7241 17586 7275
rect 17528 7235 17586 7241
rect 13480 7207 13538 7213
rect 13480 7173 13492 7207
rect 13526 7204 13538 7207
rect 13848 7207 13906 7213
rect 13848 7204 13860 7207
rect 13526 7176 13860 7204
rect 13526 7173 13538 7176
rect 13480 7167 13538 7173
rect 13848 7173 13860 7176
rect 13894 7204 13906 7207
rect 14584 7207 14642 7213
rect 14584 7204 14596 7207
rect 13894 7176 14596 7204
rect 13894 7173 13906 7176
rect 13848 7167 13906 7173
rect 14584 7173 14596 7176
rect 14630 7173 14642 7207
rect 14584 7167 14642 7173
rect 15872 7207 15930 7213
rect 15872 7173 15884 7207
rect 15918 7204 15930 7207
rect 16240 7207 16298 7213
rect 16240 7204 16252 7207
rect 15918 7176 16252 7204
rect 15918 7173 15930 7176
rect 15872 7167 15930 7173
rect 16240 7173 16252 7176
rect 16286 7204 16298 7207
rect 16976 7207 17034 7213
rect 16976 7204 16988 7207
rect 16286 7176 16988 7204
rect 16286 7173 16298 7176
rect 16240 7167 16298 7173
rect 16976 7173 16988 7176
rect 17022 7173 17034 7207
rect 16976 7167 17034 7173
rect 15691 7143 15749 7150
rect 15691 7109 15703 7143
rect 15737 7136 15749 7143
rect 18207 7136 18252 7146
rect 15737 7109 18252 7136
rect 15691 7108 18252 7109
rect 15691 7102 15749 7108
rect 18207 7098 18252 7108
rect 13370 7037 18154 7068
rect 13370 7003 13399 7037
rect 13433 7003 13491 7037
rect 13525 7006 13583 7037
rect 13561 7003 13583 7006
rect 13617 7003 13675 7037
rect 13709 7004 13767 7037
rect 13736 7003 13767 7004
rect 13801 7003 13859 7037
rect 13893 7006 13951 7037
rect 13933 7003 13951 7006
rect 13985 7003 14043 7037
rect 14077 7009 14135 7037
rect 14077 7003 14100 7009
rect 14169 7003 14227 7037
rect 14261 7003 14319 7037
rect 14353 7005 14411 7037
rect 14384 7003 14411 7005
rect 14445 7003 14503 7037
rect 14537 7012 14595 7037
rect 14537 7003 14556 7012
rect 14629 7003 14687 7037
rect 14721 7003 14779 7037
rect 14813 7003 14871 7037
rect 14905 7003 14963 7037
rect 14997 7003 15055 7037
rect 15089 7003 15147 7037
rect 15181 7003 15239 7037
rect 15273 7003 15331 7037
rect 15365 7003 15423 7037
rect 15457 7003 15515 7037
rect 15549 7003 15607 7037
rect 15641 7003 15699 7037
rect 15733 7003 15791 7037
rect 15825 7003 15883 7037
rect 15917 7003 15975 7037
rect 16009 7003 16067 7037
rect 16101 7003 16159 7037
rect 16193 7003 16251 7037
rect 16285 7003 16343 7037
rect 16377 7003 16435 7037
rect 16469 7003 16527 7037
rect 16561 7003 16619 7037
rect 16653 7003 16711 7037
rect 16745 7003 16803 7037
rect 16837 7003 16895 7037
rect 16929 7003 16987 7037
rect 17021 7003 17079 7037
rect 17113 7003 17171 7037
rect 17205 7003 17263 7037
rect 17297 7003 17355 7037
rect 17389 7003 17447 7037
rect 17481 7003 17539 7037
rect 17573 7003 17631 7037
rect 17665 7003 17723 7037
rect 17757 7003 17815 7037
rect 17849 7003 17907 7037
rect 17941 7003 17999 7037
rect 18033 7003 18091 7037
rect 18125 7003 18154 7037
rect 13370 6954 13509 7003
rect 13561 6954 13684 7003
rect 13370 6952 13684 6954
rect 13736 6954 13881 7003
rect 13933 6957 14100 7003
rect 14152 6957 14332 7003
rect 13933 6954 14332 6957
rect 13736 6953 14332 6954
rect 14384 6960 14556 7003
rect 14608 7002 17985 7003
rect 14608 7000 17763 7002
rect 14608 6960 14768 7000
rect 14384 6953 14768 6960
rect 13736 6952 14768 6953
rect 13370 6948 14768 6952
rect 14820 6996 17763 7000
rect 14820 6948 14990 6996
rect 13370 6944 14990 6948
rect 15042 6995 17763 6996
rect 15042 6993 16727 6995
rect 15042 6944 15213 6993
rect 13370 6941 15213 6944
rect 15265 6941 15423 6993
rect 15475 6941 15636 6993
rect 15688 6991 16727 6993
rect 15688 6990 16535 6991
rect 15688 6989 16356 6990
rect 15688 6986 16155 6989
rect 15688 6941 15953 6986
rect 16005 6941 16155 6986
rect 16207 6941 16356 6989
rect 16408 6941 16535 6990
rect 16587 6943 16727 6991
rect 16779 6993 17555 6995
rect 16779 6992 17349 6993
rect 16779 6943 16912 6992
rect 16587 6941 16912 6943
rect 16964 6991 17349 6992
rect 16964 6941 17144 6991
rect 17196 6941 17349 6991
rect 17401 6943 17555 6993
rect 17607 6992 17763 6995
rect 17607 6943 17655 6992
rect 17401 6941 17655 6943
rect 17707 6950 17763 6992
rect 17815 6951 17985 7002
rect 18037 6951 18154 7003
rect 17815 6950 18154 6951
rect 17707 6941 18154 6950
rect 13370 6907 13399 6941
rect 13433 6907 13491 6941
rect 13525 6907 13583 6941
rect 13617 6907 13675 6941
rect 13709 6907 13767 6941
rect 13801 6907 13859 6941
rect 13893 6907 13951 6941
rect 13985 6907 14043 6941
rect 14077 6907 14135 6941
rect 14169 6907 14227 6941
rect 14261 6907 14319 6941
rect 14353 6907 14411 6941
rect 14445 6907 14503 6941
rect 14537 6907 14595 6941
rect 14629 6907 14687 6941
rect 14721 6907 14779 6941
rect 14813 6907 14871 6941
rect 14905 6907 14963 6941
rect 14997 6907 15055 6941
rect 15089 6907 15147 6941
rect 15181 6907 15239 6941
rect 15273 6907 15331 6941
rect 15365 6907 15423 6941
rect 15457 6907 15515 6941
rect 15549 6907 15607 6941
rect 15641 6907 15699 6941
rect 15733 6907 15791 6941
rect 15825 6907 15883 6941
rect 15917 6934 15953 6941
rect 15917 6907 15975 6934
rect 16009 6907 16067 6941
rect 16101 6937 16155 6941
rect 16207 6937 16251 6941
rect 16101 6907 16159 6937
rect 16193 6907 16251 6937
rect 16285 6907 16343 6941
rect 16408 6938 16435 6941
rect 16377 6907 16435 6938
rect 16469 6907 16527 6941
rect 16587 6939 16619 6941
rect 16561 6907 16619 6939
rect 16653 6907 16711 6941
rect 16745 6907 16803 6941
rect 16837 6907 16895 6941
rect 16964 6940 16987 6941
rect 16929 6907 16987 6940
rect 17021 6907 17079 6941
rect 17113 6939 17144 6941
rect 17113 6907 17171 6939
rect 17205 6907 17263 6941
rect 17297 6907 17355 6941
rect 17389 6907 17447 6941
rect 17481 6907 17539 6941
rect 17573 6907 17631 6941
rect 17707 6940 17723 6941
rect 17665 6907 17723 6940
rect 17757 6907 17815 6941
rect 17849 6907 17907 6941
rect 17941 6907 17999 6941
rect 18033 6907 18091 6941
rect 18125 6907 18154 6941
rect 13370 6876 18154 6907
rect 18207 6837 18252 6847
rect 15689 6831 18252 6837
rect 15689 6797 15702 6831
rect 15736 6809 18252 6831
rect 15736 6797 15750 6809
rect 18207 6799 18252 6809
rect 15689 6790 15750 6797
rect 13480 6771 13538 6777
rect 13480 6737 13492 6771
rect 13526 6768 13538 6771
rect 13848 6771 13906 6777
rect 13848 6768 13860 6771
rect 13526 6740 13860 6768
rect 13526 6737 13538 6740
rect 13480 6731 13538 6737
rect 13848 6737 13860 6740
rect 13894 6768 13906 6771
rect 14584 6771 14642 6777
rect 14584 6768 14596 6771
rect 13894 6740 14596 6768
rect 13894 6737 13906 6740
rect 13848 6731 13906 6737
rect 14584 6737 14596 6740
rect 14630 6737 14642 6771
rect 14584 6731 14642 6737
rect 15872 6771 15930 6777
rect 15872 6737 15884 6771
rect 15918 6768 15930 6771
rect 16240 6771 16298 6777
rect 16240 6768 16252 6771
rect 15918 6740 16252 6768
rect 15918 6737 15930 6740
rect 15872 6731 15930 6737
rect 16240 6737 16252 6740
rect 16286 6768 16298 6771
rect 16976 6771 17034 6777
rect 16976 6768 16988 6771
rect 16286 6740 16988 6768
rect 16286 6737 16298 6740
rect 16240 6731 16298 6737
rect 16976 6737 16988 6740
rect 17022 6737 17034 6771
rect 16976 6731 17034 6737
rect 13401 6715 13453 6721
rect 14492 6703 14550 6709
rect 14492 6669 14504 6703
rect 14538 6700 14550 6703
rect 15136 6703 15194 6709
rect 15136 6700 15148 6703
rect 14538 6672 15148 6700
rect 14538 6669 14550 6672
rect 14492 6663 14550 6669
rect 15136 6669 15148 6672
rect 15182 6669 15194 6703
rect 16884 6703 16942 6709
rect 15136 6663 15194 6669
rect 15797 6673 15849 6679
rect 13401 6657 13453 6663
rect 16884 6669 16896 6703
rect 16930 6700 16942 6703
rect 17528 6703 17586 6709
rect 17528 6700 17540 6703
rect 16930 6672 17540 6700
rect 16930 6669 16942 6672
rect 16884 6663 16942 6669
rect 17528 6669 17540 6672
rect 17574 6669 17586 6703
rect 17528 6663 17586 6669
rect 13307 6629 13352 6639
rect 13723 6635 13790 6644
rect 13723 6629 13741 6635
rect 13307 6601 13741 6629
rect 13775 6601 13790 6635
rect 14584 6635 14642 6641
rect 14584 6632 14596 6635
rect 13307 6591 13352 6601
rect 13723 6593 13790 6601
rect 13955 6604 14596 6632
rect 13955 6573 13994 6604
rect 14584 6601 14596 6604
rect 14630 6601 14642 6635
rect 14584 6595 14642 6601
rect 15242 6588 15248 6640
rect 15300 6588 15306 6640
rect 16121 6634 16188 6643
rect 16121 6629 16139 6634
rect 15797 6615 15849 6621
rect 15885 6601 16139 6629
rect 13572 6567 13630 6573
rect 13572 6533 13584 6567
rect 13618 6564 13630 6567
rect 13936 6567 13994 6573
rect 13936 6564 13948 6567
rect 13618 6536 13948 6564
rect 13618 6533 13630 6536
rect 13572 6527 13630 6533
rect 13936 6533 13948 6536
rect 13982 6533 13994 6567
rect 13936 6527 13994 6533
rect 14124 6567 14182 6573
rect 14124 6533 14136 6567
rect 14170 6564 14182 6567
rect 14484 6564 14490 6576
rect 14170 6536 14490 6564
rect 14170 6533 14182 6536
rect 14124 6527 14182 6533
rect 14484 6524 14490 6536
rect 14542 6564 14548 6576
rect 14860 6567 14918 6573
rect 14860 6564 14872 6567
rect 14542 6536 14872 6564
rect 14542 6524 14548 6536
rect 14860 6533 14872 6536
rect 14906 6533 14918 6567
rect 14860 6527 14918 6533
rect 14484 6523 14548 6524
rect 13310 6495 13355 6505
rect 15885 6495 15913 6601
rect 16121 6600 16139 6601
rect 16173 6600 16188 6634
rect 16976 6635 17034 6641
rect 16976 6632 16988 6635
rect 16121 6592 16188 6600
rect 16347 6604 16988 6632
rect 16347 6573 16386 6604
rect 16976 6601 16988 6604
rect 17022 6601 17034 6635
rect 16976 6595 17034 6601
rect 17635 6589 17641 6641
rect 17693 6589 17699 6641
rect 15964 6567 16022 6573
rect 15964 6533 15976 6567
rect 16010 6564 16022 6567
rect 16328 6567 16386 6573
rect 16328 6564 16340 6567
rect 16010 6536 16340 6564
rect 16010 6533 16022 6536
rect 15964 6527 16022 6533
rect 16328 6533 16340 6536
rect 16374 6533 16386 6567
rect 16328 6527 16386 6533
rect 16516 6567 16574 6573
rect 16516 6533 16528 6567
rect 16562 6564 16574 6567
rect 16879 6564 16885 6576
rect 16562 6536 16885 6564
rect 16562 6533 16574 6536
rect 16516 6527 16574 6533
rect 16879 6524 16885 6536
rect 16937 6564 16943 6576
rect 17252 6567 17310 6573
rect 17252 6564 17264 6567
rect 16937 6536 17264 6564
rect 16937 6524 16943 6536
rect 17252 6533 17264 6536
rect 17298 6533 17310 6567
rect 17252 6527 17310 6533
rect 18080 6502 18137 6514
rect 13310 6467 15914 6495
rect 18080 6468 18092 6502
rect 18126 6499 18137 6502
rect 18212 6499 18257 6505
rect 18126 6468 18257 6499
rect 13310 6457 13355 6467
rect 18080 6465 18257 6468
rect 18080 6462 18137 6465
rect 18212 6457 18257 6465
rect 13370 6397 18154 6428
rect 13370 6363 13399 6397
rect 13433 6363 13491 6397
rect 13525 6363 13583 6397
rect 13617 6363 13675 6397
rect 13709 6363 13767 6397
rect 13801 6363 13859 6397
rect 13893 6363 13951 6397
rect 13985 6363 14043 6397
rect 14077 6363 14135 6397
rect 14169 6363 14227 6397
rect 14261 6363 14319 6397
rect 14353 6363 14411 6397
rect 14445 6363 14503 6397
rect 14537 6363 14595 6397
rect 14629 6363 14687 6397
rect 14721 6363 14779 6397
rect 14813 6363 14871 6397
rect 14905 6363 14963 6397
rect 14997 6363 15055 6397
rect 15089 6363 15147 6397
rect 15181 6363 15239 6397
rect 15273 6363 15331 6397
rect 15365 6363 15423 6397
rect 15457 6363 15515 6397
rect 15549 6363 15607 6397
rect 15641 6363 15699 6397
rect 15733 6363 15791 6397
rect 15825 6363 15883 6397
rect 15917 6363 15975 6397
rect 16009 6363 16067 6397
rect 16101 6363 16159 6397
rect 16193 6363 16251 6397
rect 16285 6363 16343 6397
rect 16377 6363 16435 6397
rect 16469 6363 16527 6397
rect 16561 6363 16619 6397
rect 16653 6363 16711 6397
rect 16745 6363 16803 6397
rect 16837 6366 16895 6397
rect 16929 6366 16987 6397
rect 16837 6363 16879 6366
rect 16931 6363 16987 6366
rect 17021 6363 17079 6397
rect 17113 6363 17171 6397
rect 17205 6363 17263 6397
rect 17297 6363 17355 6397
rect 17389 6363 17447 6397
rect 17481 6363 17539 6397
rect 17573 6363 17631 6397
rect 17665 6363 17723 6397
rect 17757 6363 17815 6397
rect 17849 6363 17907 6397
rect 17941 6363 17999 6397
rect 18033 6363 18091 6397
rect 18125 6363 18154 6397
rect 13370 6362 13958 6363
rect 13370 6357 13752 6362
rect 13370 6305 13536 6357
rect 13588 6310 13752 6357
rect 13804 6311 13958 6362
rect 14010 6360 16656 6363
rect 14010 6359 16211 6360
rect 14010 6357 14581 6359
rect 14010 6355 14356 6357
rect 14010 6311 14160 6355
rect 13804 6310 14160 6311
rect 13588 6305 14160 6310
rect 13370 6303 14160 6305
rect 14212 6305 14356 6355
rect 14408 6307 14581 6357
rect 14633 6358 15679 6359
rect 14633 6355 15239 6358
rect 14633 6307 14796 6355
rect 14408 6305 14796 6307
rect 14212 6303 14796 6305
rect 14848 6303 15031 6355
rect 15083 6306 15239 6355
rect 15291 6306 15481 6358
rect 15533 6307 15679 6358
rect 15731 6307 15986 6359
rect 16038 6308 16211 6359
rect 16263 6359 16656 6360
rect 16263 6308 16440 6359
rect 16038 6307 16440 6308
rect 16492 6311 16656 6359
rect 16708 6314 16879 6363
rect 16931 6362 18154 6363
rect 16931 6314 17103 6362
rect 16708 6311 17103 6314
rect 16492 6310 17103 6311
rect 17155 6355 18154 6362
rect 17155 6354 17981 6355
rect 17155 6351 17754 6354
rect 17155 6310 17330 6351
rect 16492 6307 17330 6310
rect 15533 6306 17330 6307
rect 15083 6303 17330 6306
rect 13370 6301 17330 6303
rect 17382 6350 17754 6351
rect 17382 6301 17543 6350
rect 17595 6302 17754 6350
rect 17806 6303 17981 6354
rect 18033 6303 18154 6355
rect 17806 6302 18154 6303
rect 17595 6301 18154 6302
rect 13370 6267 13399 6301
rect 13433 6267 13491 6301
rect 13525 6267 13583 6301
rect 13617 6267 13675 6301
rect 13709 6267 13767 6301
rect 13801 6267 13859 6301
rect 13893 6267 13951 6301
rect 13985 6267 14043 6301
rect 14077 6267 14135 6301
rect 14169 6267 14227 6301
rect 14261 6267 14319 6301
rect 14353 6267 14411 6301
rect 14445 6267 14503 6301
rect 14537 6267 14595 6301
rect 14629 6267 14687 6301
rect 14721 6267 14779 6301
rect 14813 6267 14871 6301
rect 14905 6267 14963 6301
rect 14997 6267 15055 6301
rect 15089 6267 15147 6301
rect 15181 6267 15239 6301
rect 15273 6267 15331 6301
rect 15365 6267 15423 6301
rect 15457 6267 15515 6301
rect 15549 6267 15607 6301
rect 15641 6267 15699 6301
rect 15733 6267 15791 6301
rect 15825 6267 15883 6301
rect 15917 6267 15975 6301
rect 16009 6267 16067 6301
rect 16101 6267 16159 6301
rect 16193 6267 16251 6301
rect 16285 6267 16343 6301
rect 16377 6267 16435 6301
rect 16469 6267 16527 6301
rect 16561 6267 16619 6301
rect 16653 6267 16711 6301
rect 16745 6267 16803 6301
rect 16837 6267 16895 6301
rect 16929 6267 16987 6301
rect 17021 6267 17079 6301
rect 17113 6267 17171 6301
rect 17205 6267 17263 6301
rect 17297 6299 17330 6301
rect 17297 6267 17355 6299
rect 17389 6267 17447 6301
rect 17481 6267 17539 6301
rect 17595 6298 17631 6301
rect 17573 6267 17631 6298
rect 17665 6267 17723 6301
rect 17757 6267 17815 6301
rect 17849 6267 17907 6301
rect 17941 6267 17999 6301
rect 18033 6267 18091 6301
rect 18125 6267 18154 6301
rect 13370 6236 18154 6267
rect 13297 6196 13342 6205
rect 13297 6168 15928 6196
rect 18203 6189 18248 6195
rect 18070 6179 18248 6189
rect 13297 6157 13342 6168
rect 13572 6131 13630 6137
rect 13409 6100 13461 6106
rect 13572 6097 13584 6131
rect 13618 6128 13630 6131
rect 13936 6131 13994 6137
rect 13936 6128 13948 6131
rect 13618 6100 13948 6128
rect 13618 6097 13630 6100
rect 13572 6091 13630 6097
rect 13936 6097 13948 6100
rect 13982 6097 13994 6131
rect 13936 6091 13994 6097
rect 14124 6131 14182 6137
rect 14124 6097 14136 6131
rect 14170 6128 14182 6131
rect 14860 6131 14918 6137
rect 14860 6128 14872 6131
rect 14906 6128 14918 6131
rect 14170 6100 14870 6128
rect 14170 6097 14182 6100
rect 14124 6091 14182 6097
rect 14860 6091 14870 6100
rect 13409 6042 13461 6048
rect 13955 6060 13994 6091
rect 14863 6076 14870 6091
rect 14922 6076 14929 6128
rect 14584 6063 14642 6069
rect 14584 6060 14596 6063
rect 13955 6032 14596 6060
rect 14584 6029 14596 6032
rect 14630 6029 14642 6063
rect 14584 6023 14642 6029
rect 15246 6017 15253 6069
rect 15305 6017 15312 6069
rect 15796 6057 15848 6063
rect 13728 6005 13795 6014
rect 13298 5990 13343 6002
rect 13728 5990 13746 6005
rect 13298 5971 13746 5990
rect 13780 5971 13795 6005
rect 15899 6062 15927 6168
rect 18070 6145 18086 6179
rect 18120 6155 18248 6179
rect 18120 6145 18137 6155
rect 18203 6147 18248 6155
rect 15964 6131 16022 6137
rect 15964 6097 15976 6131
rect 16010 6128 16022 6131
rect 16328 6131 16386 6137
rect 16328 6128 16340 6131
rect 16010 6100 16340 6128
rect 16010 6097 16022 6100
rect 15964 6091 16022 6097
rect 16328 6097 16340 6100
rect 16374 6097 16386 6131
rect 16328 6091 16386 6097
rect 16516 6131 16574 6137
rect 16516 6097 16528 6131
rect 16562 6128 16574 6131
rect 17252 6131 17310 6137
rect 18070 6135 18137 6145
rect 17252 6130 17264 6131
rect 17298 6130 17310 6131
rect 17252 6128 17262 6130
rect 16562 6100 17262 6128
rect 16562 6097 16574 6100
rect 16516 6091 16574 6097
rect 17252 6091 17262 6100
rect 16122 6062 16189 6071
rect 15899 6034 16140 6062
rect 16122 6028 16140 6034
rect 16174 6028 16189 6062
rect 16347 6060 16386 6091
rect 17255 6078 17262 6091
rect 17314 6078 17321 6130
rect 16976 6063 17034 6069
rect 16976 6060 16988 6063
rect 16347 6032 16988 6060
rect 16122 6020 16189 6028
rect 16976 6029 16988 6032
rect 17022 6029 17034 6063
rect 16976 6023 17034 6029
rect 17632 6024 17639 6076
rect 17691 6024 17698 6076
rect 13298 5963 13795 5971
rect 14492 5995 14550 6001
rect 13298 5962 13744 5963
rect 13298 5954 13343 5962
rect 14492 5961 14504 5995
rect 14538 5992 14550 5995
rect 15136 5995 15194 6001
rect 15796 5999 15848 6005
rect 15136 5992 15148 5995
rect 14538 5964 15148 5992
rect 14538 5961 14550 5964
rect 14492 5955 14550 5961
rect 15136 5961 15148 5964
rect 15182 5961 15194 5995
rect 15136 5955 15194 5961
rect 16884 5995 16942 6001
rect 16884 5961 16896 5995
rect 16930 5992 16942 5995
rect 17528 5995 17586 6001
rect 17528 5992 17540 5995
rect 16930 5964 17540 5992
rect 16930 5961 16942 5964
rect 16884 5955 16942 5961
rect 17528 5961 17540 5964
rect 17574 5961 17586 5995
rect 17528 5955 17586 5961
rect 13480 5927 13538 5933
rect 13480 5893 13492 5927
rect 13526 5924 13538 5927
rect 13848 5927 13906 5933
rect 13848 5924 13860 5927
rect 13526 5896 13860 5924
rect 13526 5893 13538 5896
rect 13480 5887 13538 5893
rect 13848 5893 13860 5896
rect 13894 5924 13906 5927
rect 14584 5927 14642 5933
rect 14584 5924 14596 5927
rect 13894 5896 14596 5924
rect 13894 5893 13906 5896
rect 13848 5887 13906 5893
rect 14584 5893 14596 5896
rect 14630 5893 14642 5927
rect 14584 5887 14642 5893
rect 15872 5927 15930 5933
rect 15872 5893 15884 5927
rect 15918 5924 15930 5927
rect 16240 5927 16298 5933
rect 16240 5924 16252 5927
rect 15918 5896 16252 5924
rect 15918 5893 15930 5896
rect 15872 5887 15930 5893
rect 16240 5893 16252 5896
rect 16286 5924 16298 5927
rect 16976 5927 17034 5933
rect 16976 5924 16988 5927
rect 16286 5896 16988 5924
rect 16286 5893 16298 5896
rect 16240 5887 16298 5893
rect 16976 5893 16988 5896
rect 17022 5893 17034 5927
rect 16976 5887 17034 5893
rect 15684 5868 15747 5874
rect 15684 5834 15699 5868
rect 15733 5855 15747 5868
rect 18206 5855 18251 5864
rect 15733 5834 18251 5855
rect 15684 5827 18251 5834
rect 18206 5816 18251 5827
rect 13370 5757 18154 5788
rect 13370 5723 13399 5757
rect 13433 5723 13491 5757
rect 13525 5723 13583 5757
rect 13617 5723 13675 5757
rect 13709 5723 13767 5757
rect 13801 5723 13859 5757
rect 13893 5723 13951 5757
rect 13985 5723 14043 5757
rect 14077 5723 14135 5757
rect 14169 5723 14227 5757
rect 14261 5723 14319 5757
rect 14353 5723 14411 5757
rect 14445 5723 14503 5757
rect 14537 5723 14595 5757
rect 14629 5723 14687 5757
rect 14721 5723 14779 5757
rect 14813 5723 14871 5757
rect 14905 5723 14963 5757
rect 14997 5723 15055 5757
rect 15089 5723 15147 5757
rect 15181 5726 15239 5757
rect 15181 5723 15188 5726
rect 15273 5723 15331 5757
rect 15365 5723 15423 5757
rect 15457 5728 15515 5757
rect 15478 5723 15515 5728
rect 15549 5723 15607 5757
rect 15641 5730 15699 5757
rect 15691 5723 15699 5730
rect 15733 5723 15791 5757
rect 15825 5723 15883 5757
rect 15917 5723 15975 5757
rect 16009 5723 16067 5757
rect 16101 5723 16159 5757
rect 16193 5723 16251 5757
rect 16285 5723 16343 5757
rect 16377 5723 16435 5757
rect 16469 5723 16527 5757
rect 16561 5723 16619 5757
rect 16653 5723 16711 5757
rect 16745 5723 16803 5757
rect 16837 5723 16895 5757
rect 16929 5723 16987 5757
rect 17021 5723 17079 5757
rect 17113 5723 17171 5757
rect 17205 5723 17263 5757
rect 17297 5723 17355 5757
rect 17389 5723 17447 5757
rect 17481 5723 17539 5757
rect 17573 5723 17631 5757
rect 17665 5723 17723 5757
rect 17757 5723 17815 5757
rect 17849 5723 17907 5757
rect 17941 5723 17999 5757
rect 18033 5723 18091 5757
rect 18125 5723 18154 5757
rect 13370 5722 15188 5723
rect 13370 5721 14756 5722
rect 13370 5712 13787 5721
rect 13370 5661 13562 5712
rect 13614 5669 13787 5712
rect 13839 5718 14285 5721
rect 13839 5669 14064 5718
rect 13614 5666 14064 5669
rect 14116 5669 14285 5718
rect 14337 5718 14756 5721
rect 14337 5669 14530 5718
rect 14116 5666 14530 5669
rect 14582 5670 14756 5718
rect 14808 5720 15188 5722
rect 14808 5670 14968 5720
rect 14582 5668 14968 5670
rect 15020 5674 15188 5720
rect 15240 5676 15426 5723
rect 15478 5678 15639 5723
rect 15691 5721 18154 5723
rect 15691 5720 16373 5721
rect 15691 5678 16026 5720
rect 15478 5676 16026 5678
rect 15240 5674 16026 5676
rect 15020 5668 16026 5674
rect 16078 5669 16373 5720
rect 16425 5718 18154 5721
rect 16425 5716 17032 5718
rect 16425 5669 16609 5716
rect 16078 5668 16609 5669
rect 14582 5666 16609 5668
rect 13614 5664 16609 5666
rect 16661 5664 16793 5716
rect 16845 5666 17032 5716
rect 17084 5717 18154 5718
rect 17084 5714 17802 5717
rect 17084 5666 17235 5714
rect 16845 5664 17235 5666
rect 13614 5662 17235 5664
rect 17287 5713 17802 5714
rect 17287 5711 17611 5713
rect 17287 5662 17420 5711
rect 13614 5661 17420 5662
rect 17472 5661 17611 5711
rect 17663 5665 17802 5713
rect 17854 5713 18154 5717
rect 17854 5665 17988 5713
rect 17663 5661 17988 5665
rect 18040 5661 18154 5713
rect 13370 5627 13399 5661
rect 13433 5627 13491 5661
rect 13525 5660 13562 5661
rect 13525 5627 13583 5660
rect 13617 5627 13675 5661
rect 13709 5627 13767 5661
rect 13801 5627 13859 5661
rect 13893 5627 13951 5661
rect 13985 5627 14043 5661
rect 14077 5627 14135 5661
rect 14169 5627 14227 5661
rect 14261 5627 14319 5661
rect 14353 5627 14411 5661
rect 14445 5627 14503 5661
rect 14537 5627 14595 5661
rect 14629 5627 14687 5661
rect 14721 5627 14779 5661
rect 14813 5627 14871 5661
rect 14905 5627 14963 5661
rect 14997 5627 15055 5661
rect 15089 5627 15147 5661
rect 15181 5627 15239 5661
rect 15273 5627 15331 5661
rect 15365 5627 15423 5661
rect 15457 5627 15515 5661
rect 15549 5627 15607 5661
rect 15641 5627 15699 5661
rect 15733 5627 15791 5661
rect 15825 5627 15883 5661
rect 15917 5627 15975 5661
rect 16009 5627 16067 5661
rect 16101 5627 16159 5661
rect 16193 5627 16251 5661
rect 16285 5627 16343 5661
rect 16377 5627 16435 5661
rect 16469 5627 16527 5661
rect 16561 5627 16619 5661
rect 16653 5627 16711 5661
rect 16745 5627 16803 5661
rect 16837 5627 16895 5661
rect 16929 5627 16987 5661
rect 17021 5627 17079 5661
rect 17113 5627 17171 5661
rect 17205 5627 17263 5661
rect 17297 5627 17355 5661
rect 17389 5659 17420 5661
rect 17389 5627 17447 5659
rect 17481 5627 17539 5661
rect 17573 5627 17631 5661
rect 17665 5627 17723 5661
rect 17757 5627 17815 5661
rect 17849 5627 17907 5661
rect 17941 5627 17999 5661
rect 18033 5627 18091 5661
rect 18125 5627 18154 5661
rect 13370 5596 18154 5627
rect 18209 5560 18254 5568
rect 15687 5553 18254 5560
rect 15687 5519 15699 5553
rect 15733 5532 18254 5553
rect 15733 5519 15745 5532
rect 18209 5520 18254 5532
rect 15687 5512 15745 5519
rect 13480 5491 13538 5497
rect 13480 5457 13492 5491
rect 13526 5488 13538 5491
rect 13848 5491 13906 5497
rect 13848 5488 13860 5491
rect 13526 5460 13860 5488
rect 13526 5457 13538 5460
rect 13480 5451 13538 5457
rect 13848 5457 13860 5460
rect 13894 5488 13906 5491
rect 14584 5491 14642 5497
rect 14584 5488 14596 5491
rect 13894 5460 14596 5488
rect 13894 5457 13906 5460
rect 13848 5451 13906 5457
rect 14584 5457 14596 5460
rect 14630 5457 14642 5491
rect 14584 5451 14642 5457
rect 15872 5491 15930 5497
rect 15872 5457 15884 5491
rect 15918 5488 15930 5491
rect 16240 5491 16298 5497
rect 16240 5488 16252 5491
rect 15918 5460 16252 5488
rect 15918 5457 15930 5460
rect 15872 5451 15930 5457
rect 16240 5457 16252 5460
rect 16286 5488 16298 5491
rect 16976 5491 17034 5497
rect 16976 5488 16988 5491
rect 16286 5460 16988 5488
rect 16286 5457 16298 5460
rect 16240 5451 16298 5457
rect 16976 5457 16988 5460
rect 17022 5457 17034 5491
rect 16976 5451 17034 5457
rect 13285 5412 13330 5424
rect 14492 5423 14550 5429
rect 13725 5413 13792 5422
rect 13725 5412 13743 5413
rect 13285 5384 13743 5412
rect 13285 5376 13330 5384
rect 13725 5379 13743 5384
rect 13777 5379 13792 5413
rect 14492 5389 14504 5423
rect 14538 5420 14550 5423
rect 15136 5423 15194 5429
rect 15136 5420 15148 5423
rect 14538 5392 15148 5420
rect 14538 5389 14550 5392
rect 14492 5383 14550 5389
rect 15136 5389 15148 5392
rect 15182 5389 15194 5423
rect 15136 5383 15194 5389
rect 16884 5423 16942 5429
rect 16884 5389 16896 5423
rect 16930 5420 16942 5423
rect 17528 5423 17586 5429
rect 17528 5420 17540 5423
rect 16930 5392 17540 5420
rect 16930 5389 16942 5392
rect 16884 5383 16942 5389
rect 17528 5389 17540 5392
rect 17574 5389 17586 5423
rect 17528 5383 17586 5389
rect 13725 5371 13792 5379
rect 15797 5370 15849 5376
rect 15242 5361 15307 5362
rect 14584 5355 14642 5361
rect 14584 5352 14596 5355
rect 13404 5340 13456 5346
rect 13955 5324 14596 5352
rect 13955 5293 13994 5324
rect 14584 5321 14596 5324
rect 14630 5321 14642 5355
rect 14584 5315 14642 5321
rect 15242 5309 15248 5361
rect 15300 5309 15307 5361
rect 16123 5354 16190 5363
rect 17634 5362 17698 5363
rect 16123 5349 16141 5354
rect 15797 5312 15849 5318
rect 15886 5321 16141 5349
rect 13404 5282 13456 5288
rect 13572 5287 13630 5293
rect 13572 5253 13584 5287
rect 13618 5284 13630 5287
rect 13936 5287 13994 5293
rect 13936 5284 13948 5287
rect 13618 5256 13948 5284
rect 13618 5253 13630 5256
rect 13572 5247 13630 5253
rect 13936 5253 13948 5256
rect 13982 5253 13994 5287
rect 13936 5247 13994 5253
rect 14124 5287 14182 5293
rect 14124 5253 14136 5287
rect 14170 5284 14182 5287
rect 14491 5284 14499 5296
rect 14170 5256 14499 5284
rect 14170 5253 14182 5256
rect 14124 5247 14182 5253
rect 14491 5244 14499 5256
rect 14551 5284 14557 5296
rect 14860 5287 14918 5293
rect 14860 5284 14872 5287
rect 14551 5256 14872 5284
rect 14551 5244 14557 5256
rect 14860 5253 14872 5256
rect 14906 5253 14918 5287
rect 14860 5247 14918 5253
rect 13282 5215 13327 5225
rect 15886 5215 15914 5321
rect 16123 5320 16141 5321
rect 16175 5320 16190 5354
rect 16976 5355 17034 5361
rect 16976 5352 16988 5355
rect 16123 5312 16190 5320
rect 16347 5324 16988 5352
rect 16347 5293 16386 5324
rect 16976 5321 16988 5324
rect 17022 5321 17034 5355
rect 16976 5315 17034 5321
rect 17634 5310 17640 5362
rect 17692 5310 17698 5362
rect 15964 5287 16022 5293
rect 15964 5253 15976 5287
rect 16010 5284 16022 5287
rect 16328 5287 16386 5293
rect 16328 5284 16340 5287
rect 16010 5256 16340 5284
rect 16010 5253 16022 5256
rect 15964 5247 16022 5253
rect 16328 5253 16340 5256
rect 16374 5253 16386 5287
rect 16328 5247 16386 5253
rect 16516 5287 16574 5293
rect 16516 5253 16528 5287
rect 16562 5284 16574 5287
rect 16882 5284 16889 5296
rect 16562 5256 16889 5284
rect 16562 5253 16574 5256
rect 16516 5247 16574 5253
rect 16882 5244 16889 5256
rect 16942 5284 16949 5296
rect 17252 5287 17310 5293
rect 17252 5284 17264 5287
rect 16942 5256 17264 5284
rect 16942 5244 16949 5256
rect 17252 5253 17264 5256
rect 17298 5253 17310 5287
rect 17252 5247 17310 5253
rect 18075 5220 18133 5227
rect 13282 5187 15915 5215
rect 13282 5177 13327 5187
rect 18075 5186 18087 5220
rect 18121 5218 18133 5220
rect 18205 5218 18250 5224
rect 18121 5186 18250 5218
rect 18075 5184 18250 5186
rect 18075 5180 18133 5184
rect 18205 5176 18250 5184
rect 13370 5132 18154 5148
rect 13370 5131 16150 5132
rect 13370 5130 13826 5131
rect 13370 5117 13435 5130
rect 13370 5083 13399 5117
rect 13433 5083 13435 5117
rect 13370 5078 13435 5083
rect 13487 5126 13826 5130
rect 13487 5117 13640 5126
rect 13692 5117 13826 5126
rect 13878 5129 16150 5131
rect 13878 5124 14239 5129
rect 13878 5117 14020 5124
rect 14072 5117 14239 5124
rect 14291 5117 14449 5129
rect 13487 5083 13491 5117
rect 13525 5083 13583 5117
rect 13617 5083 13640 5117
rect 13709 5083 13767 5117
rect 13801 5083 13826 5117
rect 13893 5083 13951 5117
rect 13985 5083 14020 5117
rect 14077 5083 14135 5117
rect 14169 5083 14227 5117
rect 14291 5083 14319 5117
rect 14353 5083 14411 5117
rect 14445 5083 14449 5117
rect 13487 5078 13640 5083
rect 13370 5074 13640 5078
rect 13692 5079 13826 5083
rect 13878 5079 14020 5083
rect 13692 5074 14020 5079
rect 13370 5072 14020 5074
rect 14072 5077 14239 5083
rect 14291 5077 14449 5083
rect 14501 5126 15932 5129
rect 14501 5117 14678 5126
rect 14730 5117 14924 5126
rect 14976 5117 15198 5126
rect 15250 5117 15473 5126
rect 15525 5117 15709 5126
rect 15761 5117 15932 5126
rect 15984 5117 16150 5129
rect 16202 5130 18154 5132
rect 16202 5126 17595 5130
rect 16202 5125 17175 5126
rect 16202 5123 16567 5125
rect 16202 5117 16328 5123
rect 16380 5117 16567 5123
rect 14501 5083 14503 5117
rect 14537 5083 14595 5117
rect 14629 5083 14678 5117
rect 14730 5083 14779 5117
rect 14813 5083 14871 5117
rect 14905 5083 14924 5117
rect 14997 5083 15055 5117
rect 15089 5083 15147 5117
rect 15181 5083 15198 5117
rect 15273 5083 15331 5117
rect 15365 5083 15423 5117
rect 15457 5083 15473 5117
rect 15549 5083 15607 5117
rect 15641 5083 15699 5117
rect 15761 5083 15791 5117
rect 15825 5083 15883 5117
rect 15917 5083 15932 5117
rect 16009 5083 16067 5117
rect 16101 5083 16150 5117
rect 16202 5083 16251 5117
rect 16285 5083 16328 5117
rect 16380 5083 16435 5117
rect 16469 5083 16527 5117
rect 16561 5083 16567 5117
rect 14501 5077 14678 5083
rect 14072 5074 14678 5077
rect 14730 5074 14924 5083
rect 14976 5074 15198 5083
rect 15250 5074 15473 5083
rect 15525 5074 15709 5083
rect 15761 5077 15932 5083
rect 15984 5080 16150 5083
rect 16202 5080 16328 5083
rect 15984 5077 16328 5080
rect 15761 5074 16328 5077
rect 14072 5072 16328 5074
rect 13370 5071 16328 5072
rect 16380 5073 16567 5083
rect 16619 5117 16764 5125
rect 16816 5117 16962 5125
rect 17014 5117 17175 5125
rect 17227 5125 17595 5126
rect 17227 5117 17398 5125
rect 17450 5117 17595 5125
rect 17647 5128 18154 5130
rect 17647 5117 17811 5128
rect 17863 5117 18020 5128
rect 18072 5117 18154 5128
rect 16653 5083 16711 5117
rect 16745 5083 16764 5117
rect 16837 5083 16895 5117
rect 16929 5083 16962 5117
rect 17021 5083 17079 5117
rect 17113 5083 17171 5117
rect 17227 5083 17263 5117
rect 17297 5083 17355 5117
rect 17389 5083 17398 5117
rect 17481 5083 17539 5117
rect 17573 5083 17595 5117
rect 17665 5083 17723 5117
rect 17757 5083 17811 5117
rect 17863 5083 17907 5117
rect 17941 5083 17999 5117
rect 18072 5083 18091 5117
rect 18125 5083 18154 5117
rect 16619 5073 16764 5083
rect 16816 5073 16962 5083
rect 17014 5074 17175 5083
rect 17227 5074 17398 5083
rect 17014 5073 17398 5074
rect 17450 5078 17595 5083
rect 17647 5078 17811 5083
rect 17450 5076 17811 5078
rect 17863 5076 18020 5083
rect 18072 5076 18154 5083
rect 17450 5073 18154 5076
rect 16380 5071 18154 5073
rect 13370 5052 18154 5071
rect 13399 5049 13433 5052
rect 13491 5049 13525 5052
rect 13583 5049 13617 5052
rect 13675 5049 13709 5052
rect 13767 5049 13801 5052
rect 13859 5049 13893 5052
rect 13951 5049 13985 5052
rect 14043 5049 14077 5052
rect 14135 5049 14169 5052
rect 14227 5049 14261 5052
rect 14319 5049 14353 5052
rect 14411 5049 14445 5052
rect 14503 5049 14537 5052
rect 14595 5049 14629 5052
rect 14687 5049 14721 5052
rect 14779 5049 14813 5052
rect 14871 5049 14905 5052
rect 14963 5049 14997 5052
rect 15055 5049 15089 5052
rect 15147 5049 15181 5052
rect 15239 5049 15273 5052
rect 15331 5049 15365 5052
rect 15423 5049 15457 5052
rect 15515 5049 15549 5052
rect 15607 5049 15641 5052
rect 15699 5049 15733 5052
rect 15791 5049 15825 5052
rect 15883 5049 15917 5052
rect 15975 5049 16009 5052
rect 16067 5049 16101 5052
rect 16159 5049 16193 5052
rect 16251 5049 16285 5052
rect 16343 5049 16377 5052
rect 16435 5049 16469 5052
rect 16527 5049 16561 5052
rect 16619 5049 16653 5052
rect 16711 5049 16745 5052
rect 16803 5049 16837 5052
rect 16895 5049 16929 5052
rect 16987 5049 17021 5052
rect 17079 5049 17113 5052
rect 17171 5049 17205 5052
rect 17263 5049 17297 5052
rect 17355 5049 17389 5052
rect 17447 5049 17481 5052
rect 17539 5049 17573 5052
rect 17631 5049 17665 5052
rect 17723 5049 17757 5052
rect 17815 5049 17849 5052
rect 17907 5049 17941 5052
rect 17999 5049 18033 5052
rect 18091 5049 18125 5052
<< via1 >>
rect 12474 10560 12526 10612
rect 12572 10591 12624 10603
rect 12572 10557 12582 10591
rect 12582 10557 12616 10591
rect 12616 10557 12624 10591
rect 12572 10551 12624 10557
rect 12652 10591 12704 10603
rect 12652 10557 12662 10591
rect 12662 10557 12696 10591
rect 12696 10557 12704 10591
rect 12652 10551 12704 10557
rect 12732 10591 12784 10603
rect 12732 10557 12742 10591
rect 12742 10557 12776 10591
rect 12776 10557 12784 10591
rect 12732 10551 12784 10557
rect 12812 10591 12864 10603
rect 12812 10557 12822 10591
rect 12822 10557 12856 10591
rect 12856 10557 12864 10591
rect 12812 10551 12864 10557
rect 12892 10591 12944 10603
rect 12892 10557 12902 10591
rect 12902 10557 12936 10591
rect 12936 10557 12944 10591
rect 12892 10551 12944 10557
rect 12972 10591 13024 10603
rect 12972 10557 12982 10591
rect 12982 10557 13016 10591
rect 13016 10557 13024 10591
rect 12972 10551 13024 10557
rect 13304 10594 13356 10606
rect 13304 10560 13314 10594
rect 13314 10560 13348 10594
rect 13348 10560 13356 10594
rect 13304 10554 13356 10560
rect 13384 10594 13436 10606
rect 13384 10560 13394 10594
rect 13394 10560 13428 10594
rect 13428 10560 13436 10594
rect 13384 10554 13436 10560
rect 13464 10594 13516 10606
rect 13464 10560 13474 10594
rect 13474 10560 13508 10594
rect 13508 10560 13516 10594
rect 13464 10554 13516 10560
rect 13544 10594 13596 10606
rect 13544 10560 13554 10594
rect 13554 10560 13588 10594
rect 13588 10560 13596 10594
rect 13544 10554 13596 10560
rect 13624 10594 13676 10606
rect 13624 10560 13634 10594
rect 13634 10560 13668 10594
rect 13668 10560 13676 10594
rect 13624 10554 13676 10560
rect 13704 10594 13756 10606
rect 13704 10560 13714 10594
rect 13714 10560 13748 10594
rect 13748 10560 13756 10594
rect 13704 10554 13756 10560
rect 13908 10594 13960 10606
rect 13908 10560 13916 10594
rect 13916 10560 13950 10594
rect 13950 10560 13960 10594
rect 13908 10554 13960 10560
rect 13988 10594 14040 10606
rect 13988 10560 13996 10594
rect 13996 10560 14030 10594
rect 14030 10560 14040 10594
rect 13988 10554 14040 10560
rect 14068 10594 14120 10606
rect 14068 10560 14076 10594
rect 14076 10560 14110 10594
rect 14110 10560 14120 10594
rect 14068 10554 14120 10560
rect 14148 10594 14200 10606
rect 14148 10560 14156 10594
rect 14156 10560 14190 10594
rect 14190 10560 14200 10594
rect 14148 10554 14200 10560
rect 14228 10594 14280 10606
rect 14228 10560 14236 10594
rect 14236 10560 14270 10594
rect 14270 10560 14280 10594
rect 14228 10554 14280 10560
rect 14308 10594 14360 10606
rect 14308 10560 14316 10594
rect 14316 10560 14350 10594
rect 14350 10560 14360 10594
rect 14308 10554 14360 10560
rect 14516 10594 14568 10606
rect 14516 10560 14526 10594
rect 14526 10560 14560 10594
rect 14560 10560 14568 10594
rect 14516 10554 14568 10560
rect 14596 10594 14648 10606
rect 14596 10560 14606 10594
rect 14606 10560 14640 10594
rect 14640 10560 14648 10594
rect 14596 10554 14648 10560
rect 14676 10594 14728 10606
rect 14676 10560 14686 10594
rect 14686 10560 14720 10594
rect 14720 10560 14728 10594
rect 14676 10554 14728 10560
rect 14756 10594 14808 10606
rect 14756 10560 14766 10594
rect 14766 10560 14800 10594
rect 14800 10560 14808 10594
rect 14756 10554 14808 10560
rect 14836 10594 14888 10606
rect 14836 10560 14846 10594
rect 14846 10560 14880 10594
rect 14880 10560 14888 10594
rect 14836 10554 14888 10560
rect 14916 10594 14968 10606
rect 14916 10560 14926 10594
rect 14926 10560 14960 10594
rect 14960 10560 14968 10594
rect 14916 10554 14968 10560
rect 15120 10594 15172 10606
rect 15120 10560 15128 10594
rect 15128 10560 15162 10594
rect 15162 10560 15172 10594
rect 15120 10554 15172 10560
rect 15200 10594 15252 10606
rect 15200 10560 15208 10594
rect 15208 10560 15242 10594
rect 15242 10560 15252 10594
rect 15200 10554 15252 10560
rect 15280 10594 15332 10606
rect 15280 10560 15288 10594
rect 15288 10560 15322 10594
rect 15322 10560 15332 10594
rect 15280 10554 15332 10560
rect 15360 10594 15412 10606
rect 15360 10560 15368 10594
rect 15368 10560 15402 10594
rect 15402 10560 15412 10594
rect 15360 10554 15412 10560
rect 15440 10594 15492 10606
rect 15440 10560 15448 10594
rect 15448 10560 15482 10594
rect 15482 10560 15492 10594
rect 15440 10554 15492 10560
rect 15520 10594 15572 10606
rect 15520 10560 15528 10594
rect 15528 10560 15562 10594
rect 15562 10560 15572 10594
rect 15520 10554 15572 10560
rect 15728 10594 15780 10606
rect 15728 10560 15738 10594
rect 15738 10560 15772 10594
rect 15772 10560 15780 10594
rect 15728 10554 15780 10560
rect 15808 10594 15860 10606
rect 15808 10560 15818 10594
rect 15818 10560 15852 10594
rect 15852 10560 15860 10594
rect 15808 10554 15860 10560
rect 15888 10594 15940 10606
rect 15888 10560 15898 10594
rect 15898 10560 15932 10594
rect 15932 10560 15940 10594
rect 15888 10554 15940 10560
rect 15968 10594 16020 10606
rect 15968 10560 15978 10594
rect 15978 10560 16012 10594
rect 16012 10560 16020 10594
rect 15968 10554 16020 10560
rect 16048 10594 16100 10606
rect 16048 10560 16058 10594
rect 16058 10560 16092 10594
rect 16092 10560 16100 10594
rect 16048 10554 16100 10560
rect 16128 10594 16180 10606
rect 16128 10560 16138 10594
rect 16138 10560 16172 10594
rect 16172 10560 16180 10594
rect 16128 10554 16180 10560
rect 16332 10594 16384 10606
rect 16332 10560 16340 10594
rect 16340 10560 16374 10594
rect 16374 10560 16384 10594
rect 16332 10554 16384 10560
rect 16412 10594 16464 10606
rect 16412 10560 16420 10594
rect 16420 10560 16454 10594
rect 16454 10560 16464 10594
rect 16412 10554 16464 10560
rect 16492 10594 16544 10606
rect 16492 10560 16500 10594
rect 16500 10560 16534 10594
rect 16534 10560 16544 10594
rect 16492 10554 16544 10560
rect 16572 10594 16624 10606
rect 16572 10560 16580 10594
rect 16580 10560 16614 10594
rect 16614 10560 16624 10594
rect 16572 10554 16624 10560
rect 16652 10594 16704 10606
rect 16652 10560 16660 10594
rect 16660 10560 16694 10594
rect 16694 10560 16704 10594
rect 16652 10554 16704 10560
rect 16732 10594 16784 10606
rect 16732 10560 16740 10594
rect 16740 10560 16774 10594
rect 16774 10560 16784 10594
rect 16732 10554 16784 10560
rect 16940 10594 16992 10606
rect 16940 10560 16950 10594
rect 16950 10560 16984 10594
rect 16984 10560 16992 10594
rect 16940 10554 16992 10560
rect 17020 10594 17072 10606
rect 17020 10560 17030 10594
rect 17030 10560 17064 10594
rect 17064 10560 17072 10594
rect 17020 10554 17072 10560
rect 17100 10594 17152 10606
rect 17100 10560 17110 10594
rect 17110 10560 17144 10594
rect 17144 10560 17152 10594
rect 17100 10554 17152 10560
rect 17180 10594 17232 10606
rect 17180 10560 17190 10594
rect 17190 10560 17224 10594
rect 17224 10560 17232 10594
rect 17180 10554 17232 10560
rect 17260 10594 17312 10606
rect 17260 10560 17270 10594
rect 17270 10560 17304 10594
rect 17304 10560 17312 10594
rect 17260 10554 17312 10560
rect 17340 10594 17392 10606
rect 17340 10560 17350 10594
rect 17350 10560 17384 10594
rect 17384 10560 17392 10594
rect 17340 10554 17392 10560
rect 17544 10594 17596 10606
rect 17544 10560 17552 10594
rect 17552 10560 17586 10594
rect 17586 10560 17596 10594
rect 17544 10554 17596 10560
rect 17624 10594 17676 10606
rect 17624 10560 17632 10594
rect 17632 10560 17666 10594
rect 17666 10560 17676 10594
rect 17624 10554 17676 10560
rect 17704 10594 17756 10606
rect 17704 10560 17712 10594
rect 17712 10560 17746 10594
rect 17746 10560 17756 10594
rect 17704 10554 17756 10560
rect 17784 10594 17836 10606
rect 17784 10560 17792 10594
rect 17792 10560 17826 10594
rect 17826 10560 17836 10594
rect 17784 10554 17836 10560
rect 17864 10594 17916 10606
rect 17864 10560 17872 10594
rect 17872 10560 17906 10594
rect 17906 10560 17916 10594
rect 17864 10554 17916 10560
rect 17944 10594 17996 10606
rect 17944 10560 17952 10594
rect 17952 10560 17986 10594
rect 17986 10560 17996 10594
rect 17944 10554 17996 10560
rect 18283 10543 18335 10550
rect 18283 10509 18294 10543
rect 18294 10509 18328 10543
rect 18328 10509 18335 10543
rect 18283 10498 18335 10509
rect 18288 10399 18340 10406
rect 18288 10365 18299 10399
rect 18299 10365 18333 10399
rect 18333 10365 18340 10399
rect 18288 10354 18340 10365
rect 18289 10247 18341 10254
rect 18289 10213 18300 10247
rect 18300 10213 18334 10247
rect 18334 10213 18341 10247
rect 18289 10202 18341 10213
rect 11857 9955 11909 10007
rect 11988 9996 12040 10006
rect 11988 9962 12005 9996
rect 12005 9962 12039 9996
rect 12039 9962 12040 9996
rect 11988 9954 12040 9962
rect 12132 9955 12184 10007
rect 18289 10077 18341 10084
rect 18289 10043 18300 10077
rect 18300 10043 18334 10077
rect 18334 10043 18341 10077
rect 18289 10032 18341 10043
rect 12130 9687 12182 9696
rect 12130 9653 12142 9687
rect 12142 9653 12176 9687
rect 12176 9653 12182 9687
rect 12130 9644 12182 9653
rect 18288 9920 18340 9927
rect 18288 9886 18299 9920
rect 18299 9886 18333 9920
rect 18333 9886 18340 9920
rect 18288 9875 18340 9886
rect 11875 9452 11927 9461
rect 11995 9452 12047 9461
rect 12138 9452 12190 9461
rect 11875 9418 11913 9452
rect 11913 9418 11927 9452
rect 11995 9418 12005 9452
rect 12005 9418 12039 9452
rect 12039 9418 12047 9452
rect 12138 9418 12189 9452
rect 12189 9418 12190 9452
rect 11875 9409 11927 9418
rect 11995 9409 12047 9418
rect 12138 9409 12190 9418
rect 12142 9066 12194 9118
rect 18206 9633 18258 9685
rect 18583 9641 18635 9693
rect 18783 9641 18835 9693
rect 12954 9422 13018 9425
rect 12954 9362 12976 9422
rect 12976 9362 13010 9422
rect 13010 9362 13018 9422
rect 12954 9361 13018 9362
rect 13686 9425 13750 9428
rect 13686 9365 13708 9425
rect 13708 9365 13742 9425
rect 13742 9365 13750 9425
rect 13686 9364 13750 9365
rect 13914 9425 13978 9428
rect 13914 9365 13922 9425
rect 13922 9365 13956 9425
rect 13956 9365 13978 9425
rect 13914 9364 13978 9365
rect 14898 9425 14962 9428
rect 14898 9365 14920 9425
rect 14920 9365 14954 9425
rect 14954 9365 14962 9425
rect 14898 9364 14962 9365
rect 15126 9425 15190 9428
rect 15126 9365 15134 9425
rect 15134 9365 15168 9425
rect 15168 9365 15190 9425
rect 15126 9364 15190 9365
rect 16110 9425 16174 9428
rect 16110 9365 16132 9425
rect 16132 9365 16166 9425
rect 16166 9365 16174 9425
rect 16110 9364 16174 9365
rect 16338 9425 16402 9428
rect 16338 9365 16346 9425
rect 16346 9365 16380 9425
rect 16380 9365 16402 9425
rect 16338 9364 16402 9365
rect 17322 9425 17386 9428
rect 17322 9365 17344 9425
rect 17344 9365 17378 9425
rect 17378 9365 17386 9425
rect 17322 9364 17386 9365
rect 17550 9425 17614 9428
rect 17550 9365 17558 9425
rect 17558 9365 17592 9425
rect 17592 9365 17614 9425
rect 17550 9364 17614 9365
rect 18294 9372 18303 9424
rect 18303 9372 18337 9424
rect 18337 9372 18346 9424
rect 13310 9224 13374 9226
rect 13310 9164 13329 9224
rect 13329 9164 13363 9224
rect 13363 9164 13374 9224
rect 13310 9162 13374 9164
rect 14042 9224 14106 9226
rect 14042 9164 14061 9224
rect 14061 9164 14095 9224
rect 14095 9164 14106 9224
rect 14042 9162 14106 9164
rect 14260 9224 14324 9226
rect 14260 9164 14271 9224
rect 14271 9164 14305 9224
rect 14305 9164 14324 9224
rect 14260 9162 14324 9164
rect 15254 9224 15318 9226
rect 15254 9164 15273 9224
rect 15273 9164 15307 9224
rect 15307 9164 15318 9224
rect 15254 9162 15318 9164
rect 15472 9224 15536 9226
rect 15472 9164 15483 9224
rect 15483 9164 15517 9224
rect 15517 9164 15536 9224
rect 15472 9162 15536 9164
rect 16592 9224 16656 9226
rect 16592 9164 16611 9224
rect 16611 9164 16645 9224
rect 16645 9164 16656 9224
rect 16592 9162 16656 9164
rect 16810 9224 16874 9226
rect 16810 9164 16821 9224
rect 16821 9164 16855 9224
rect 16855 9164 16874 9224
rect 16810 9162 16874 9164
rect 17544 9224 17608 9226
rect 17544 9164 17555 9224
rect 17555 9164 17589 9224
rect 17589 9164 17608 9224
rect 17544 9162 17608 9164
rect 18294 9169 18303 9221
rect 18303 9169 18337 9221
rect 18337 9169 18346 9221
rect 12630 9066 12682 9118
rect 12460 8014 12469 8034
rect 12469 8014 12503 8034
rect 12503 8014 12512 8034
rect 12460 7982 12512 8014
rect 13002 8027 13054 8037
rect 13002 7993 13010 8027
rect 13010 7993 13044 8027
rect 13044 7993 13054 8027
rect 13002 7985 13054 7993
rect 13082 8027 13134 8037
rect 13082 7993 13090 8027
rect 13090 7993 13124 8027
rect 13124 7993 13134 8027
rect 13082 7985 13134 7993
rect 13162 8027 13214 8037
rect 13162 7993 13170 8027
rect 13170 7993 13204 8027
rect 13204 7993 13214 8027
rect 13162 7985 13214 7993
rect 13242 8027 13294 8037
rect 13242 7993 13250 8027
rect 13250 7993 13284 8027
rect 13284 7993 13294 8027
rect 13242 7985 13294 7993
rect 13734 8027 13786 8037
rect 13734 7993 13742 8027
rect 13742 7993 13776 8027
rect 13776 7993 13786 8027
rect 13734 7985 13786 7993
rect 13814 8027 13866 8037
rect 13814 7993 13822 8027
rect 13822 7993 13856 8027
rect 13856 7993 13866 8027
rect 13814 7985 13866 7993
rect 13894 8027 13946 8037
rect 13894 7993 13902 8027
rect 13902 7993 13936 8027
rect 13936 7993 13946 8027
rect 13894 7985 13946 7993
rect 13974 8027 14026 8037
rect 13974 7993 13982 8027
rect 13982 7993 14016 8027
rect 14016 7993 14026 8027
rect 13974 7985 14026 7993
rect 14340 8027 14392 8037
rect 14340 7993 14350 8027
rect 14350 7993 14384 8027
rect 14384 7993 14392 8027
rect 14340 7985 14392 7993
rect 14420 8027 14472 8037
rect 14420 7993 14430 8027
rect 14430 7993 14464 8027
rect 14464 7993 14472 8027
rect 14420 7985 14472 7993
rect 14500 8027 14552 8037
rect 14500 7993 14510 8027
rect 14510 7993 14544 8027
rect 14544 7993 14552 8027
rect 14500 7985 14552 7993
rect 14580 8027 14632 8037
rect 14580 7993 14590 8027
rect 14590 7993 14624 8027
rect 14624 7993 14632 8027
rect 14580 7985 14632 7993
rect 14946 8027 14998 8037
rect 14946 7993 14954 8027
rect 14954 7993 14988 8027
rect 14988 7993 14998 8027
rect 14946 7985 14998 7993
rect 15026 8027 15078 8037
rect 15026 7993 15034 8027
rect 15034 7993 15068 8027
rect 15068 7993 15078 8027
rect 15026 7985 15078 7993
rect 15106 8027 15158 8037
rect 15106 7993 15114 8027
rect 15114 7993 15148 8027
rect 15148 7993 15158 8027
rect 15106 7985 15158 7993
rect 15186 8027 15238 8037
rect 15186 7993 15194 8027
rect 15194 7993 15228 8027
rect 15228 7993 15238 8027
rect 15186 7985 15238 7993
rect 15552 8027 15604 8037
rect 15552 7993 15562 8027
rect 15562 7993 15596 8027
rect 15596 7993 15604 8027
rect 15552 7985 15604 7993
rect 15632 8027 15684 8037
rect 15632 7993 15642 8027
rect 15642 7993 15676 8027
rect 15676 7993 15684 8027
rect 15632 7985 15684 7993
rect 15712 8027 15764 8037
rect 15712 7993 15722 8027
rect 15722 7993 15756 8027
rect 15756 7993 15764 8027
rect 15712 7985 15764 7993
rect 15792 8027 15844 8037
rect 15792 7993 15802 8027
rect 15802 7993 15836 8027
rect 15836 7993 15844 8027
rect 15792 7985 15844 7993
rect 16284 8027 16336 8037
rect 16284 7993 16292 8027
rect 16292 7993 16326 8027
rect 16326 7993 16336 8027
rect 16284 7985 16336 7993
rect 16364 8027 16416 8037
rect 16364 7993 16372 8027
rect 16372 7993 16406 8027
rect 16406 7993 16416 8027
rect 16364 7985 16416 7993
rect 16444 8027 16496 8037
rect 16444 7993 16452 8027
rect 16452 7993 16486 8027
rect 16486 7993 16496 8027
rect 16444 7985 16496 7993
rect 16524 8027 16576 8037
rect 16524 7993 16532 8027
rect 16532 7993 16566 8027
rect 16566 7993 16576 8027
rect 16524 7985 16576 7993
rect 16890 8027 16942 8037
rect 16890 7993 16900 8027
rect 16900 7993 16934 8027
rect 16934 7993 16942 8027
rect 16890 7985 16942 7993
rect 16970 8027 17022 8037
rect 16970 7993 16980 8027
rect 16980 7993 17014 8027
rect 17014 7993 17022 8027
rect 16970 7985 17022 7993
rect 17050 8027 17102 8037
rect 17050 7993 17060 8027
rect 17060 7993 17094 8027
rect 17094 7993 17102 8027
rect 17050 7985 17102 7993
rect 17130 8027 17182 8037
rect 17130 7993 17140 8027
rect 17140 7993 17174 8027
rect 17174 7993 17182 8027
rect 17130 7985 17182 7993
rect 18394 8999 18446 9051
rect 18203 8907 18255 8959
rect 17624 8027 17676 8037
rect 17624 7993 17634 8027
rect 17634 7993 17668 8027
rect 17668 7993 17676 8027
rect 17624 7985 17676 7993
rect 17704 8027 17756 8037
rect 17704 7993 17714 8027
rect 17714 7993 17748 8027
rect 17748 7993 17756 8027
rect 17704 7985 17756 7993
rect 17784 8027 17836 8037
rect 17784 7993 17794 8027
rect 17794 7993 17828 8027
rect 17828 7993 17836 8027
rect 17784 7985 17836 7993
rect 17864 8027 17916 8037
rect 17864 7993 17874 8027
rect 17874 7993 17908 8027
rect 17908 7993 17916 8027
rect 17864 7985 17916 7993
rect 13415 7655 13467 7707
rect 15809 7655 15861 7707
rect 13507 7581 13559 7589
rect 13681 7581 13733 7588
rect 13906 7581 13958 7590
rect 14107 7581 14159 7592
rect 14330 7581 14382 7590
rect 13507 7547 13525 7581
rect 13525 7547 13559 7581
rect 13681 7547 13709 7581
rect 13709 7547 13733 7581
rect 13906 7547 13951 7581
rect 13951 7547 13958 7581
rect 14107 7547 14135 7581
rect 14135 7547 14159 7581
rect 14330 7547 14353 7581
rect 14353 7547 14382 7581
rect 13507 7537 13559 7547
rect 13681 7536 13733 7547
rect 13906 7538 13958 7547
rect 14107 7540 14159 7547
rect 14330 7538 14382 7547
rect 14539 7543 14591 7595
rect 14767 7581 14819 7588
rect 14957 7581 15009 7592
rect 15162 7581 15214 7595
rect 15361 7581 15413 7595
rect 15577 7581 15629 7590
rect 15965 7581 16017 7595
rect 16200 7581 16252 7590
rect 16442 7581 16494 7592
rect 16674 7581 16726 7593
rect 16903 7581 16955 7596
rect 17152 7581 17204 7588
rect 17370 7581 17422 7592
rect 17599 7581 17651 7588
rect 17820 7581 17872 7590
rect 14767 7547 14779 7581
rect 14779 7547 14813 7581
rect 14813 7547 14819 7581
rect 14957 7547 14963 7581
rect 14963 7547 14997 7581
rect 14997 7547 15009 7581
rect 15162 7547 15181 7581
rect 15181 7547 15214 7581
rect 15361 7547 15365 7581
rect 15365 7547 15413 7581
rect 15577 7547 15607 7581
rect 15607 7547 15629 7581
rect 15965 7547 15975 7581
rect 15975 7547 16009 7581
rect 16009 7547 16017 7581
rect 16200 7547 16251 7581
rect 16251 7547 16252 7581
rect 16442 7547 16469 7581
rect 16469 7547 16494 7581
rect 16674 7547 16711 7581
rect 16711 7547 16726 7581
rect 16903 7547 16929 7581
rect 16929 7547 16955 7581
rect 17152 7547 17171 7581
rect 17171 7547 17204 7581
rect 17370 7547 17389 7581
rect 17389 7547 17422 7581
rect 17599 7547 17631 7581
rect 17631 7547 17651 7581
rect 17820 7547 17849 7581
rect 17849 7547 17872 7581
rect 14767 7536 14819 7547
rect 14957 7540 15009 7547
rect 15162 7543 15214 7547
rect 15361 7543 15413 7547
rect 15577 7538 15629 7547
rect 15965 7543 16017 7547
rect 16200 7538 16252 7547
rect 16442 7540 16494 7547
rect 16674 7541 16726 7547
rect 16903 7544 16955 7547
rect 17152 7536 17204 7547
rect 17370 7540 17422 7547
rect 17599 7536 17651 7547
rect 17820 7538 17872 7547
rect 18036 7543 18088 7595
rect 13406 7355 13458 7364
rect 13406 7321 13416 7355
rect 13416 7321 13450 7355
rect 13450 7321 13458 7355
rect 13406 7312 13458 7321
rect 14865 7377 14872 7402
rect 14872 7377 14906 7402
rect 14906 7377 14917 7402
rect 14865 7350 14917 7377
rect 15250 7340 15302 7351
rect 15250 7306 15255 7340
rect 15255 7306 15289 7340
rect 15289 7306 15302 7340
rect 15250 7299 15302 7306
rect 17260 7377 17264 7401
rect 17264 7377 17298 7401
rect 17298 7377 17312 7401
rect 15798 7310 15850 7322
rect 15798 7276 15805 7310
rect 15805 7276 15839 7310
rect 15839 7276 15850 7310
rect 17260 7349 17312 7377
rect 17645 7344 17697 7352
rect 17645 7310 17654 7344
rect 17654 7310 17688 7344
rect 17688 7310 17697 7344
rect 17645 7300 17697 7310
rect 15798 7270 15850 7276
rect 13509 7003 13525 7006
rect 13525 7003 13561 7006
rect 13684 7003 13709 7004
rect 13709 7003 13736 7004
rect 13881 7003 13893 7006
rect 13893 7003 13933 7006
rect 14100 7003 14135 7009
rect 14135 7003 14152 7009
rect 14332 7003 14353 7005
rect 14353 7003 14384 7005
rect 14556 7003 14595 7012
rect 14595 7003 14608 7012
rect 13509 6954 13561 7003
rect 13684 6952 13736 7003
rect 13881 6954 13933 7003
rect 14100 6957 14152 7003
rect 14332 6953 14384 7003
rect 14556 6960 14608 7003
rect 14768 6948 14820 7000
rect 14990 6944 15042 6996
rect 15213 6941 15265 6993
rect 15423 6941 15475 6993
rect 15636 6941 15688 6993
rect 15953 6941 16005 6986
rect 16155 6941 16207 6989
rect 16356 6941 16408 6990
rect 16535 6941 16587 6991
rect 16727 6943 16779 6995
rect 16912 6941 16964 6992
rect 17144 6941 17196 6991
rect 17349 6941 17401 6993
rect 17555 6943 17607 6995
rect 17655 6941 17707 6992
rect 17763 6950 17815 7002
rect 17985 6951 18037 7003
rect 15953 6934 15975 6941
rect 15975 6934 16005 6941
rect 16155 6937 16159 6941
rect 16159 6937 16193 6941
rect 16193 6937 16207 6941
rect 16356 6938 16377 6941
rect 16377 6938 16408 6941
rect 16535 6939 16561 6941
rect 16561 6939 16587 6941
rect 16912 6940 16929 6941
rect 16929 6940 16964 6941
rect 17144 6939 17171 6941
rect 17171 6939 17196 6941
rect 17655 6940 17665 6941
rect 17665 6940 17707 6941
rect 13401 6705 13453 6715
rect 13401 6671 13411 6705
rect 13411 6671 13445 6705
rect 13445 6671 13453 6705
rect 13401 6663 13453 6671
rect 15797 6662 15849 6673
rect 15248 6633 15300 6640
rect 15248 6599 15256 6633
rect 15256 6599 15290 6633
rect 15290 6599 15300 6633
rect 15248 6588 15300 6599
rect 15797 6628 15806 6662
rect 15806 6628 15840 6662
rect 15840 6628 15849 6662
rect 15797 6621 15849 6628
rect 14490 6524 14542 6576
rect 17641 6634 17693 6641
rect 17641 6600 17649 6634
rect 17649 6600 17683 6634
rect 17683 6600 17693 6634
rect 17641 6589 17693 6600
rect 16885 6524 16937 6576
rect 16879 6363 16895 6366
rect 16895 6363 16929 6366
rect 16929 6363 16931 6366
rect 13536 6305 13588 6357
rect 13752 6310 13804 6362
rect 13958 6311 14010 6363
rect 14160 6303 14212 6355
rect 14356 6305 14408 6357
rect 14581 6307 14633 6359
rect 14796 6303 14848 6355
rect 15031 6303 15083 6355
rect 15239 6306 15291 6358
rect 15481 6306 15533 6358
rect 15679 6307 15731 6359
rect 15986 6307 16038 6359
rect 16211 6308 16263 6360
rect 16440 6307 16492 6359
rect 16656 6311 16708 6363
rect 16879 6314 16931 6363
rect 17103 6310 17155 6362
rect 17330 6301 17382 6351
rect 17543 6301 17595 6350
rect 17754 6302 17806 6354
rect 17981 6303 18033 6355
rect 17330 6299 17355 6301
rect 17355 6299 17382 6301
rect 17543 6298 17573 6301
rect 17573 6298 17595 6301
rect 13409 6089 13461 6100
rect 14870 6097 14872 6128
rect 14872 6097 14906 6128
rect 14906 6097 14922 6128
rect 13409 6055 13419 6089
rect 13419 6055 13453 6089
rect 13453 6055 13461 6089
rect 13409 6048 13461 6055
rect 14870 6076 14922 6097
rect 15253 6063 15305 6069
rect 15253 6029 15265 6063
rect 15265 6029 15299 6063
rect 15299 6029 15305 6063
rect 15253 6017 15305 6029
rect 15796 6045 15848 6057
rect 15796 6011 15803 6045
rect 15803 6011 15837 6045
rect 15837 6011 15848 6045
rect 17262 6097 17264 6130
rect 17264 6097 17298 6130
rect 17298 6097 17314 6130
rect 17262 6078 17314 6097
rect 17639 6065 17691 6076
rect 17639 6031 17649 6065
rect 17649 6031 17683 6065
rect 17683 6031 17691 6065
rect 17639 6024 17691 6031
rect 15796 6005 15848 6011
rect 15188 5723 15239 5726
rect 15239 5723 15240 5726
rect 15426 5723 15457 5728
rect 15457 5723 15478 5728
rect 15639 5723 15641 5730
rect 15641 5723 15691 5730
rect 13562 5661 13614 5712
rect 13787 5669 13839 5721
rect 14064 5666 14116 5718
rect 14285 5669 14337 5721
rect 14530 5666 14582 5718
rect 14756 5670 14808 5722
rect 14968 5668 15020 5720
rect 15188 5674 15240 5723
rect 15426 5676 15478 5723
rect 15639 5678 15691 5723
rect 16026 5668 16078 5720
rect 16373 5669 16425 5721
rect 16609 5664 16661 5716
rect 16793 5664 16845 5716
rect 17032 5666 17084 5718
rect 17235 5662 17287 5714
rect 17420 5661 17472 5711
rect 17611 5661 17663 5713
rect 17802 5665 17854 5717
rect 17988 5661 18040 5713
rect 13562 5660 13583 5661
rect 13583 5660 13614 5661
rect 17420 5659 17447 5661
rect 17447 5659 17472 5661
rect 13404 5329 13456 5340
rect 13404 5295 13415 5329
rect 13415 5295 13449 5329
rect 13449 5295 13456 5329
rect 13404 5288 13456 5295
rect 15248 5353 15300 5361
rect 15248 5319 15257 5353
rect 15257 5319 15291 5353
rect 15291 5319 15300 5353
rect 15248 5309 15300 5319
rect 15797 5359 15849 5370
rect 15797 5325 15804 5359
rect 15804 5325 15838 5359
rect 15838 5325 15849 5359
rect 15797 5318 15849 5325
rect 14499 5244 14551 5296
rect 17640 5354 17692 5362
rect 17640 5320 17649 5354
rect 17649 5320 17683 5354
rect 17683 5320 17692 5354
rect 17640 5310 17692 5320
rect 16889 5244 16942 5296
rect 13435 5078 13487 5130
rect 13640 5117 13692 5126
rect 13826 5117 13878 5131
rect 14020 5117 14072 5124
rect 14239 5117 14291 5129
rect 13640 5083 13675 5117
rect 13675 5083 13692 5117
rect 13826 5083 13859 5117
rect 13859 5083 13878 5117
rect 14020 5083 14043 5117
rect 14043 5083 14072 5117
rect 14239 5083 14261 5117
rect 14261 5083 14291 5117
rect 13640 5074 13692 5083
rect 13826 5079 13878 5083
rect 14020 5072 14072 5083
rect 14239 5077 14291 5083
rect 14449 5077 14501 5129
rect 14678 5117 14730 5126
rect 14924 5117 14976 5126
rect 15198 5117 15250 5126
rect 15473 5117 15525 5126
rect 15709 5117 15761 5126
rect 15932 5117 15984 5129
rect 16150 5117 16202 5132
rect 16328 5117 16380 5123
rect 14678 5083 14687 5117
rect 14687 5083 14721 5117
rect 14721 5083 14730 5117
rect 14924 5083 14963 5117
rect 14963 5083 14976 5117
rect 15198 5083 15239 5117
rect 15239 5083 15250 5117
rect 15473 5083 15515 5117
rect 15515 5083 15525 5117
rect 15709 5083 15733 5117
rect 15733 5083 15761 5117
rect 15932 5083 15975 5117
rect 15975 5083 15984 5117
rect 16150 5083 16159 5117
rect 16159 5083 16193 5117
rect 16193 5083 16202 5117
rect 16328 5083 16343 5117
rect 16343 5083 16377 5117
rect 16377 5083 16380 5117
rect 14678 5074 14730 5083
rect 14924 5074 14976 5083
rect 15198 5074 15250 5083
rect 15473 5074 15525 5083
rect 15709 5074 15761 5083
rect 15932 5077 15984 5083
rect 16150 5080 16202 5083
rect 16328 5071 16380 5083
rect 16567 5073 16619 5125
rect 16764 5117 16816 5125
rect 16962 5117 17014 5125
rect 17175 5117 17227 5126
rect 17398 5117 17450 5125
rect 17595 5117 17647 5130
rect 17811 5117 17863 5128
rect 18020 5117 18072 5128
rect 16764 5083 16803 5117
rect 16803 5083 16816 5117
rect 16962 5083 16987 5117
rect 16987 5083 17014 5117
rect 17175 5083 17205 5117
rect 17205 5083 17227 5117
rect 17398 5083 17447 5117
rect 17447 5083 17450 5117
rect 17595 5083 17631 5117
rect 17631 5083 17647 5117
rect 17811 5083 17815 5117
rect 17815 5083 17849 5117
rect 17849 5083 17863 5117
rect 18020 5083 18033 5117
rect 18033 5083 18072 5117
rect 16764 5073 16816 5083
rect 16962 5073 17014 5083
rect 17175 5074 17227 5083
rect 17398 5073 17450 5083
rect 17595 5078 17647 5083
rect 17811 5076 17863 5083
rect 18020 5076 18072 5083
<< metal2 >>
rect 12463 10614 12537 10618
rect 12463 10558 12472 10614
rect 12528 10609 12537 10614
rect 12528 10605 13134 10609
rect 12528 10558 12568 10605
rect 12463 10554 12568 10558
rect 12464 10549 12568 10554
rect 12624 10549 12648 10605
rect 12704 10549 12728 10605
rect 12784 10549 12808 10605
rect 12864 10549 12888 10605
rect 12944 10549 12968 10605
rect 13024 10549 13134 10605
rect 12464 10543 13134 10549
rect 13196 10608 18104 10612
rect 13196 10552 13300 10608
rect 13356 10552 13380 10608
rect 13436 10552 13460 10608
rect 13516 10552 13540 10608
rect 13596 10552 13620 10608
rect 13676 10552 13700 10608
rect 13756 10552 13908 10608
rect 13964 10552 13988 10608
rect 14044 10552 14068 10608
rect 14124 10552 14148 10608
rect 14204 10552 14228 10608
rect 14284 10552 14308 10608
rect 14364 10552 14512 10608
rect 14568 10552 14592 10608
rect 14648 10552 14672 10608
rect 14728 10552 14752 10608
rect 14808 10552 14832 10608
rect 14888 10552 14912 10608
rect 14968 10552 15120 10608
rect 15176 10552 15200 10608
rect 15256 10552 15280 10608
rect 15336 10552 15360 10608
rect 15416 10552 15440 10608
rect 15496 10552 15520 10608
rect 15576 10552 15724 10608
rect 15780 10552 15804 10608
rect 15860 10552 15884 10608
rect 15940 10552 15964 10608
rect 16020 10552 16044 10608
rect 16100 10552 16124 10608
rect 16180 10552 16332 10608
rect 16388 10552 16412 10608
rect 16468 10552 16492 10608
rect 16548 10552 16572 10608
rect 16628 10552 16652 10608
rect 16708 10552 16732 10608
rect 16788 10552 16936 10608
rect 16992 10552 17016 10608
rect 17072 10552 17096 10608
rect 17152 10552 17176 10608
rect 17232 10552 17256 10608
rect 17312 10552 17336 10608
rect 17392 10552 17544 10608
rect 17600 10552 17624 10608
rect 17680 10552 17704 10608
rect 17760 10552 17784 10608
rect 17840 10552 17864 10608
rect 17920 10552 17944 10608
rect 18000 10552 18104 10608
rect 13196 10546 18104 10552
rect 18272 10552 18346 10556
rect 18272 10496 18281 10552
rect 18337 10496 18346 10552
rect 18272 10492 18346 10496
rect 18277 10408 18351 10412
rect 18277 10352 18286 10408
rect 18342 10352 18351 10408
rect 18277 10348 18351 10352
rect 18278 10256 18352 10260
rect 18278 10200 18287 10256
rect 18343 10200 18352 10256
rect 18278 10196 18352 10200
rect 18278 10086 18352 10090
rect 18278 10030 18287 10086
rect 18343 10030 18352 10086
rect 18278 10026 18352 10030
rect 11855 10009 11911 10018
rect 11855 9944 11911 9953
rect 11986 10008 12042 10017
rect 11986 9943 12042 9952
rect 12130 10009 12186 10018
rect 12130 9944 12186 9953
rect 18277 9929 18351 9933
rect 18277 9873 18286 9929
rect 18342 9873 18351 9929
rect 18277 9869 18351 9873
rect 12122 9644 12130 9696
rect 12182 9644 12188 9696
rect 18572 9695 18646 9699
rect 12122 9643 12188 9644
rect 18195 9687 18269 9691
rect 12140 9567 12186 9643
rect 18195 9631 18204 9687
rect 18260 9631 18269 9687
rect 18572 9639 18581 9695
rect 18637 9639 18646 9695
rect 18572 9635 18646 9639
rect 18772 9695 18846 9699
rect 18772 9639 18781 9695
rect 18837 9639 18846 9695
rect 18772 9635 18846 9639
rect 18195 9627 18269 9631
rect 12140 9521 12379 9567
rect 11873 9463 11929 9472
rect 11873 9398 11929 9407
rect 11993 9463 12049 9472
rect 11993 9398 12049 9407
rect 12136 9463 12192 9472
rect 12136 9398 12192 9407
rect 12136 9118 12201 9119
rect 12136 9066 12142 9118
rect 12194 9115 12201 9118
rect 12333 9115 12379 9521
rect 13679 9428 13758 9429
rect 13906 9428 13985 9429
rect 14891 9428 14970 9429
rect 15118 9428 15197 9429
rect 16103 9428 16182 9429
rect 16330 9428 16409 9429
rect 17315 9428 17394 9429
rect 17542 9428 17621 9429
rect 12947 9425 13026 9426
rect 12944 9361 12954 9425
rect 13018 9361 13027 9425
rect 13676 9364 13686 9428
rect 13750 9364 13759 9428
rect 13905 9364 13914 9428
rect 13978 9364 13988 9428
rect 14888 9364 14898 9428
rect 14962 9364 14971 9428
rect 15117 9364 15126 9428
rect 15190 9364 15200 9428
rect 16100 9364 16110 9428
rect 16174 9364 16183 9428
rect 16329 9364 16338 9428
rect 16402 9364 16412 9428
rect 17312 9364 17322 9428
rect 17386 9364 17395 9428
rect 17541 9364 17550 9428
rect 17614 9364 17624 9428
rect 18283 9426 18357 9430
rect 18283 9370 18292 9426
rect 18348 9370 18357 9426
rect 18283 9366 18357 9370
rect 13301 9162 13310 9226
rect 13374 9162 13383 9226
rect 13301 9161 13383 9162
rect 14033 9162 14042 9226
rect 14106 9162 14115 9226
rect 14033 9161 14115 9162
rect 14251 9162 14260 9226
rect 14324 9162 14333 9226
rect 14251 9161 14333 9162
rect 15245 9162 15254 9226
rect 15318 9162 15327 9226
rect 15245 9161 15327 9162
rect 15463 9162 15472 9226
rect 15536 9162 15545 9226
rect 15463 9161 15545 9162
rect 16583 9162 16592 9226
rect 16656 9162 16665 9226
rect 16583 9161 16665 9162
rect 16801 9162 16810 9226
rect 16874 9162 16883 9226
rect 16801 9161 16883 9162
rect 17535 9162 17544 9226
rect 17608 9162 17617 9226
rect 18283 9223 18357 9227
rect 18283 9167 18292 9223
rect 18348 9167 18357 9223
rect 18283 9163 18357 9167
rect 17535 9161 17617 9162
rect 12623 9115 12630 9118
rect 12194 9069 12630 9115
rect 12194 9066 12201 9069
rect 12623 9066 12630 9069
rect 12682 9066 12688 9118
rect 12623 9065 12688 9066
rect 18383 9053 18457 9057
rect 18383 8997 18392 9053
rect 18448 8997 18457 9053
rect 18383 8993 18457 8997
rect 18192 8961 18266 8965
rect 18192 8905 18201 8961
rect 18257 8905 18266 8961
rect 18192 8901 18266 8905
rect 12449 8036 12523 8040
rect 12449 7980 12458 8036
rect 12514 7980 12523 8036
rect 12449 7976 12523 7980
rect 12984 8039 13316 8043
rect 12984 7983 13000 8039
rect 13056 7983 13080 8039
rect 13136 7983 13160 8039
rect 13216 7983 13240 8039
rect 13296 7983 13316 8039
rect 12984 7975 13316 7983
rect 13716 8039 14048 8043
rect 13716 7983 13732 8039
rect 13788 7983 13812 8039
rect 13868 7983 13892 8039
rect 13948 7983 13972 8039
rect 14028 7983 14048 8039
rect 13716 7975 14048 7983
rect 14318 8039 14650 8043
rect 14318 7983 14338 8039
rect 14394 7983 14418 8039
rect 14474 7983 14498 8039
rect 14554 7983 14578 8039
rect 14634 7983 14650 8039
rect 14318 7975 14650 7983
rect 14928 8039 15260 8043
rect 14928 7983 14944 8039
rect 15000 7983 15024 8039
rect 15080 7983 15104 8039
rect 15160 7983 15184 8039
rect 15240 7983 15260 8039
rect 14928 7975 15260 7983
rect 15530 8039 15862 8043
rect 15530 7983 15550 8039
rect 15606 7983 15630 8039
rect 15686 7983 15710 8039
rect 15766 7983 15790 8039
rect 15846 7983 15862 8039
rect 15530 7975 15862 7983
rect 16266 8039 16598 8043
rect 16266 7983 16282 8039
rect 16338 7983 16362 8039
rect 16418 7983 16442 8039
rect 16498 7983 16522 8039
rect 16578 7983 16598 8039
rect 16266 7975 16598 7983
rect 16868 8039 17200 8043
rect 16868 7983 16888 8039
rect 16944 7983 16968 8039
rect 17024 7983 17048 8039
rect 17104 7983 17128 8039
rect 17184 7983 17200 8039
rect 16868 7975 17200 7983
rect 17602 8039 17934 8043
rect 17602 7983 17622 8039
rect 17678 7983 17702 8039
rect 17758 7983 17782 8039
rect 17838 7983 17862 8039
rect 17918 7983 17934 8039
rect 17602 7975 17934 7983
rect 13409 7655 13415 7707
rect 13467 7655 13473 7707
rect 15803 7655 15809 7707
rect 15861 7655 15867 7707
rect 13428 7370 13456 7655
rect 13496 7535 13505 7591
rect 13561 7535 13571 7591
rect 13496 7534 13571 7535
rect 13670 7534 13679 7590
rect 13735 7534 13745 7590
rect 13895 7536 13904 7592
rect 13960 7536 13970 7592
rect 14096 7538 14105 7594
rect 14161 7538 14171 7594
rect 14096 7537 14171 7538
rect 13895 7535 13970 7536
rect 14319 7536 14328 7592
rect 14384 7536 14394 7592
rect 14528 7541 14537 7597
rect 14593 7541 14603 7597
rect 14528 7540 14603 7541
rect 14319 7535 14394 7536
rect 13670 7533 13745 7534
rect 14756 7534 14765 7590
rect 14821 7534 14831 7590
rect 14946 7538 14955 7594
rect 15011 7538 15021 7594
rect 15151 7541 15160 7597
rect 15216 7541 15226 7597
rect 15151 7540 15226 7541
rect 15350 7541 15359 7597
rect 15415 7541 15425 7597
rect 15350 7540 15425 7541
rect 14946 7537 15021 7538
rect 15566 7536 15575 7592
rect 15631 7536 15641 7592
rect 15566 7535 15641 7536
rect 14756 7533 14831 7534
rect 13406 7364 13458 7370
rect 14854 7348 14863 7404
rect 14919 7348 14929 7404
rect 14854 7347 14929 7348
rect 13406 7306 13458 7312
rect 13428 6721 13456 7306
rect 15239 7297 15248 7353
rect 15304 7297 15314 7353
rect 15822 7328 15850 7655
rect 15954 7541 15963 7597
rect 16019 7541 16029 7597
rect 15954 7540 16029 7541
rect 16189 7536 16198 7592
rect 16254 7536 16264 7592
rect 16431 7538 16440 7594
rect 16496 7538 16506 7594
rect 16663 7539 16672 7595
rect 16728 7539 16738 7595
rect 16892 7542 16901 7598
rect 16957 7542 16967 7598
rect 16892 7541 16967 7542
rect 16663 7538 16738 7539
rect 16431 7537 16506 7538
rect 16189 7535 16264 7536
rect 17141 7534 17150 7590
rect 17206 7534 17216 7590
rect 17359 7538 17368 7594
rect 17424 7538 17434 7594
rect 17359 7537 17434 7538
rect 17141 7533 17216 7534
rect 17588 7534 17597 7590
rect 17653 7534 17663 7590
rect 17809 7536 17818 7592
rect 17874 7536 17884 7592
rect 18025 7541 18034 7597
rect 18090 7541 18100 7597
rect 18025 7540 18100 7541
rect 17809 7535 17884 7536
rect 17588 7533 17663 7534
rect 17249 7347 17258 7403
rect 17314 7347 17324 7403
rect 17249 7346 17324 7347
rect 15239 7296 15314 7297
rect 15798 7322 15850 7328
rect 17634 7298 17643 7354
rect 17699 7298 17709 7354
rect 17634 7297 17709 7298
rect 15798 7264 15850 7270
rect 13498 6952 13507 7008
rect 13563 6952 13573 7008
rect 13498 6951 13573 6952
rect 13673 6950 13682 7006
rect 13738 6950 13748 7006
rect 13870 6952 13879 7008
rect 13935 6952 13945 7008
rect 14089 6955 14098 7011
rect 14154 6955 14164 7011
rect 14089 6954 14164 6955
rect 13870 6951 13945 6952
rect 14321 6951 14330 7007
rect 14386 6951 14396 7007
rect 14321 6950 14396 6951
rect 14505 6958 14554 7014
rect 14610 6958 14620 7014
rect 13673 6949 13748 6950
rect 13401 6715 13456 6721
rect 13453 6663 13456 6715
rect 13401 6657 13456 6663
rect 13428 6106 13456 6657
rect 14505 6905 14620 6958
rect 14757 6946 14766 7002
rect 14822 6946 14832 7002
rect 14757 6945 14832 6946
rect 14979 6942 14988 6998
rect 15044 6942 15054 6998
rect 14979 6941 15054 6942
rect 15201 6995 15289 7000
rect 15201 6939 15211 6995
rect 15267 6939 15289 6995
rect 15201 6919 15289 6939
rect 15412 6939 15421 6995
rect 15477 6939 15487 6995
rect 15412 6938 15487 6939
rect 15625 6939 15634 6995
rect 15690 6939 15700 6995
rect 15625 6938 15700 6939
rect 14505 6576 14549 6905
rect 15253 6640 15289 6919
rect 15822 6679 15850 7264
rect 15942 6932 15951 6988
rect 16007 6932 16017 6988
rect 16144 6935 16153 6991
rect 16209 6935 16219 6991
rect 16345 6936 16354 6992
rect 16410 6936 16420 6992
rect 16524 6937 16533 6993
rect 16589 6937 16599 6993
rect 16716 6941 16725 6997
rect 16781 6941 16791 6997
rect 16716 6940 16791 6941
rect 16889 6994 16977 6998
rect 16524 6936 16599 6937
rect 16889 6938 16910 6994
rect 16966 6938 16977 6994
rect 16345 6935 16420 6936
rect 16144 6934 16219 6935
rect 15942 6931 16017 6932
rect 15797 6673 15850 6679
rect 15242 6588 15248 6640
rect 15300 6588 15306 6640
rect 15849 6621 15850 6673
rect 15797 6615 15850 6621
rect 14484 6524 14490 6576
rect 14542 6559 14549 6576
rect 14542 6524 14548 6559
rect 14484 6523 14548 6524
rect 13525 6303 13534 6359
rect 13590 6303 13600 6359
rect 13741 6308 13750 6364
rect 13806 6308 13816 6364
rect 13947 6309 13956 6365
rect 14012 6309 14022 6365
rect 13947 6308 14022 6309
rect 13741 6307 13816 6308
rect 13525 6302 13600 6303
rect 14149 6301 14158 6357
rect 14214 6301 14224 6357
rect 14345 6303 14354 6359
rect 14410 6303 14420 6359
rect 14570 6305 14579 6361
rect 14635 6305 14645 6361
rect 14570 6304 14645 6305
rect 14345 6302 14420 6303
rect 14149 6300 14224 6301
rect 14785 6301 14794 6357
rect 14850 6301 14860 6357
rect 14785 6300 14860 6301
rect 15020 6301 15029 6357
rect 15085 6301 15095 6357
rect 15228 6304 15237 6360
rect 15293 6304 15303 6360
rect 15228 6303 15303 6304
rect 15470 6304 15479 6360
rect 15535 6304 15545 6360
rect 15668 6305 15677 6361
rect 15733 6305 15743 6361
rect 15668 6304 15743 6305
rect 15470 6303 15545 6304
rect 15020 6300 15095 6301
rect 13409 6100 13461 6106
rect 14859 6074 14868 6130
rect 14924 6074 14934 6130
rect 14859 6073 14934 6074
rect 13409 6042 13461 6048
rect 13428 5346 13456 6042
rect 15242 6015 15251 6071
rect 15307 6015 15317 6071
rect 15822 6063 15850 6615
rect 16889 6923 16977 6938
rect 17133 6937 17142 6993
rect 17198 6937 17208 6993
rect 17338 6939 17347 6995
rect 17403 6939 17413 6995
rect 17544 6941 17553 6997
rect 17609 6941 17619 6997
rect 17544 6940 17619 6941
rect 17649 6940 17655 6992
rect 17707 6940 17713 6992
rect 17752 6948 17761 7004
rect 17817 6948 17827 7004
rect 17974 6949 17983 7005
rect 18039 6949 18049 7005
rect 17974 6948 18049 6949
rect 17752 6947 17827 6948
rect 17338 6938 17413 6939
rect 17133 6936 17208 6937
rect 16889 6576 16933 6923
rect 17649 6641 17699 6940
rect 17635 6589 17641 6641
rect 17693 6589 17699 6641
rect 16879 6524 16885 6576
rect 16937 6524 16943 6576
rect 15975 6305 15984 6361
rect 16040 6305 16050 6361
rect 16200 6306 16209 6362
rect 16265 6306 16275 6362
rect 16200 6305 16275 6306
rect 16429 6305 16438 6361
rect 16494 6305 16504 6361
rect 16645 6309 16654 6365
rect 16710 6309 16720 6365
rect 16868 6312 16877 6368
rect 16933 6312 16943 6368
rect 16868 6311 16943 6312
rect 16645 6308 16720 6309
rect 17092 6308 17101 6364
rect 17157 6308 17167 6364
rect 17092 6307 17167 6308
rect 15975 6304 16050 6305
rect 16429 6304 16504 6305
rect 17319 6297 17328 6353
rect 17384 6297 17394 6353
rect 17319 6296 17394 6297
rect 17532 6296 17541 6352
rect 17597 6296 17607 6352
rect 17743 6300 17752 6356
rect 17808 6300 17818 6356
rect 17970 6301 17979 6357
rect 18035 6301 18045 6357
rect 17970 6300 18045 6301
rect 17743 6299 17818 6300
rect 17532 6295 17607 6296
rect 17251 6076 17260 6132
rect 17316 6076 17326 6132
rect 17251 6075 17326 6076
rect 15242 6014 15317 6015
rect 15796 6057 15850 6063
rect 15848 6005 15850 6057
rect 17628 6022 17637 6078
rect 17693 6022 17703 6078
rect 17628 6021 17703 6022
rect 15796 5999 15850 6005
rect 13551 5658 13560 5714
rect 13616 5658 13626 5714
rect 13776 5667 13785 5723
rect 13841 5667 13851 5723
rect 13776 5666 13851 5667
rect 14053 5664 14062 5720
rect 14118 5664 14128 5720
rect 14274 5667 14283 5723
rect 14339 5667 14349 5723
rect 14274 5666 14349 5667
rect 14490 5720 14558 5722
rect 14053 5663 14128 5664
rect 14490 5664 14528 5720
rect 14584 5664 14594 5720
rect 14745 5668 14754 5724
rect 14810 5668 14820 5724
rect 14745 5667 14820 5668
rect 14957 5666 14966 5722
rect 15022 5666 15032 5722
rect 15177 5672 15186 5728
rect 15242 5725 15252 5728
rect 15242 5672 15291 5725
rect 15415 5674 15424 5730
rect 15480 5674 15490 5730
rect 15628 5676 15637 5732
rect 15693 5676 15703 5732
rect 15628 5675 15703 5676
rect 15415 5673 15490 5674
rect 15177 5671 15291 5672
rect 14957 5665 15032 5666
rect 14490 5663 14594 5664
rect 13551 5657 13626 5658
rect 13404 5340 13456 5346
rect 14507 5296 14543 5663
rect 15246 5362 15291 5671
rect 15822 5376 15850 5999
rect 16015 5666 16024 5722
rect 16080 5666 16090 5722
rect 16362 5667 16371 5723
rect 16427 5667 16437 5723
rect 16779 5720 17096 5726
rect 16779 5718 17030 5720
rect 16362 5666 16437 5667
rect 16015 5665 16090 5666
rect 16598 5662 16607 5718
rect 16663 5662 16673 5718
rect 16598 5661 16673 5662
rect 16779 5662 16791 5718
rect 16847 5664 17030 5718
rect 17086 5664 17096 5720
rect 16847 5662 17096 5664
rect 16779 5651 17096 5662
rect 17224 5660 17233 5716
rect 17289 5660 17299 5716
rect 17224 5659 17299 5660
rect 17409 5657 17418 5713
rect 17474 5657 17484 5713
rect 17600 5659 17609 5715
rect 17665 5712 17675 5715
rect 17665 5659 17688 5712
rect 17791 5663 17800 5719
rect 17856 5663 17866 5719
rect 17791 5662 17866 5663
rect 17600 5658 17688 5659
rect 17977 5659 17986 5715
rect 18042 5659 18052 5715
rect 17977 5658 18052 5659
rect 17409 5656 17484 5657
rect 15797 5370 15850 5376
rect 15242 5361 15307 5362
rect 15242 5309 15248 5361
rect 15300 5309 15307 5361
rect 15849 5318 15850 5370
rect 15797 5312 15850 5318
rect 13404 5282 13456 5288
rect 13428 5281 13456 5282
rect 14490 5257 14499 5296
rect 14491 5244 14499 5257
rect 14551 5257 14558 5296
rect 15822 5294 15850 5312
rect 16900 5296 16936 5651
rect 17651 5363 17688 5658
rect 17634 5362 17698 5363
rect 17634 5310 17640 5362
rect 17692 5310 17698 5362
rect 14551 5244 14557 5257
rect 16882 5244 16889 5296
rect 16942 5244 16949 5296
rect 13424 5076 13433 5132
rect 13489 5076 13499 5132
rect 13424 5075 13499 5076
rect 13629 5072 13638 5128
rect 13694 5072 13704 5128
rect 13815 5077 13824 5133
rect 13880 5077 13890 5133
rect 13815 5076 13890 5077
rect 13629 5071 13704 5072
rect 14009 5070 14018 5126
rect 14074 5070 14084 5126
rect 14228 5075 14237 5131
rect 14293 5075 14303 5131
rect 14228 5074 14303 5075
rect 14438 5075 14447 5131
rect 14503 5075 14513 5131
rect 14438 5074 14513 5075
rect 14667 5072 14676 5128
rect 14732 5072 14742 5128
rect 14667 5071 14742 5072
rect 14913 5072 14922 5128
rect 14978 5072 14988 5128
rect 14913 5071 14988 5072
rect 15187 5072 15196 5128
rect 15252 5072 15262 5128
rect 15187 5071 15262 5072
rect 15462 5072 15471 5128
rect 15527 5072 15537 5128
rect 15462 5071 15537 5072
rect 15698 5072 15707 5128
rect 15763 5072 15773 5128
rect 15921 5075 15930 5131
rect 15986 5075 15996 5131
rect 16139 5078 16148 5134
rect 16204 5078 16214 5134
rect 16139 5077 16214 5078
rect 15921 5074 15996 5075
rect 15698 5071 15773 5072
rect 14009 5069 14084 5070
rect 16317 5069 16326 5125
rect 16382 5069 16392 5125
rect 16556 5071 16565 5127
rect 16621 5071 16631 5127
rect 16556 5070 16631 5071
rect 16753 5071 16762 5127
rect 16818 5071 16828 5127
rect 16753 5070 16828 5071
rect 16951 5071 16960 5127
rect 17016 5071 17026 5127
rect 17164 5072 17173 5128
rect 17229 5072 17239 5128
rect 17164 5071 17239 5072
rect 17387 5071 17396 5127
rect 17452 5071 17462 5127
rect 17584 5076 17593 5132
rect 17649 5076 17659 5132
rect 17584 5075 17659 5076
rect 17800 5074 17809 5130
rect 17865 5074 17875 5130
rect 17800 5073 17875 5074
rect 18009 5074 18018 5130
rect 18074 5074 18084 5130
rect 18009 5073 18084 5074
rect 16951 5070 17026 5071
rect 17387 5070 17462 5071
rect 16317 5068 16392 5069
<< via2 >>
rect 12472 10612 12528 10614
rect 12472 10560 12474 10612
rect 12474 10560 12526 10612
rect 12526 10560 12528 10612
rect 12472 10558 12528 10560
rect 12568 10603 12624 10605
rect 12568 10551 12572 10603
rect 12572 10551 12624 10603
rect 12568 10549 12624 10551
rect 12648 10603 12704 10605
rect 12648 10551 12652 10603
rect 12652 10551 12704 10603
rect 12648 10549 12704 10551
rect 12728 10603 12784 10605
rect 12728 10551 12732 10603
rect 12732 10551 12784 10603
rect 12728 10549 12784 10551
rect 12808 10603 12864 10605
rect 12808 10551 12812 10603
rect 12812 10551 12864 10603
rect 12808 10549 12864 10551
rect 12888 10603 12944 10605
rect 12888 10551 12892 10603
rect 12892 10551 12944 10603
rect 12888 10549 12944 10551
rect 12968 10603 13024 10605
rect 12968 10551 12972 10603
rect 12972 10551 13024 10603
rect 12968 10549 13024 10551
rect 13300 10606 13356 10608
rect 13300 10554 13304 10606
rect 13304 10554 13356 10606
rect 13300 10552 13356 10554
rect 13380 10606 13436 10608
rect 13380 10554 13384 10606
rect 13384 10554 13436 10606
rect 13380 10552 13436 10554
rect 13460 10606 13516 10608
rect 13460 10554 13464 10606
rect 13464 10554 13516 10606
rect 13460 10552 13516 10554
rect 13540 10606 13596 10608
rect 13540 10554 13544 10606
rect 13544 10554 13596 10606
rect 13540 10552 13596 10554
rect 13620 10606 13676 10608
rect 13620 10554 13624 10606
rect 13624 10554 13676 10606
rect 13620 10552 13676 10554
rect 13700 10606 13756 10608
rect 13700 10554 13704 10606
rect 13704 10554 13756 10606
rect 13700 10552 13756 10554
rect 13908 10606 13964 10608
rect 13908 10554 13960 10606
rect 13960 10554 13964 10606
rect 13908 10552 13964 10554
rect 13988 10606 14044 10608
rect 13988 10554 14040 10606
rect 14040 10554 14044 10606
rect 13988 10552 14044 10554
rect 14068 10606 14124 10608
rect 14068 10554 14120 10606
rect 14120 10554 14124 10606
rect 14068 10552 14124 10554
rect 14148 10606 14204 10608
rect 14148 10554 14200 10606
rect 14200 10554 14204 10606
rect 14148 10552 14204 10554
rect 14228 10606 14284 10608
rect 14228 10554 14280 10606
rect 14280 10554 14284 10606
rect 14228 10552 14284 10554
rect 14308 10606 14364 10608
rect 14308 10554 14360 10606
rect 14360 10554 14364 10606
rect 14308 10552 14364 10554
rect 14512 10606 14568 10608
rect 14512 10554 14516 10606
rect 14516 10554 14568 10606
rect 14512 10552 14568 10554
rect 14592 10606 14648 10608
rect 14592 10554 14596 10606
rect 14596 10554 14648 10606
rect 14592 10552 14648 10554
rect 14672 10606 14728 10608
rect 14672 10554 14676 10606
rect 14676 10554 14728 10606
rect 14672 10552 14728 10554
rect 14752 10606 14808 10608
rect 14752 10554 14756 10606
rect 14756 10554 14808 10606
rect 14752 10552 14808 10554
rect 14832 10606 14888 10608
rect 14832 10554 14836 10606
rect 14836 10554 14888 10606
rect 14832 10552 14888 10554
rect 14912 10606 14968 10608
rect 14912 10554 14916 10606
rect 14916 10554 14968 10606
rect 14912 10552 14968 10554
rect 15120 10606 15176 10608
rect 15120 10554 15172 10606
rect 15172 10554 15176 10606
rect 15120 10552 15176 10554
rect 15200 10606 15256 10608
rect 15200 10554 15252 10606
rect 15252 10554 15256 10606
rect 15200 10552 15256 10554
rect 15280 10606 15336 10608
rect 15280 10554 15332 10606
rect 15332 10554 15336 10606
rect 15280 10552 15336 10554
rect 15360 10606 15416 10608
rect 15360 10554 15412 10606
rect 15412 10554 15416 10606
rect 15360 10552 15416 10554
rect 15440 10606 15496 10608
rect 15440 10554 15492 10606
rect 15492 10554 15496 10606
rect 15440 10552 15496 10554
rect 15520 10606 15576 10608
rect 15520 10554 15572 10606
rect 15572 10554 15576 10606
rect 15520 10552 15576 10554
rect 15724 10606 15780 10608
rect 15724 10554 15728 10606
rect 15728 10554 15780 10606
rect 15724 10552 15780 10554
rect 15804 10606 15860 10608
rect 15804 10554 15808 10606
rect 15808 10554 15860 10606
rect 15804 10552 15860 10554
rect 15884 10606 15940 10608
rect 15884 10554 15888 10606
rect 15888 10554 15940 10606
rect 15884 10552 15940 10554
rect 15964 10606 16020 10608
rect 15964 10554 15968 10606
rect 15968 10554 16020 10606
rect 15964 10552 16020 10554
rect 16044 10606 16100 10608
rect 16044 10554 16048 10606
rect 16048 10554 16100 10606
rect 16044 10552 16100 10554
rect 16124 10606 16180 10608
rect 16124 10554 16128 10606
rect 16128 10554 16180 10606
rect 16124 10552 16180 10554
rect 16332 10606 16388 10608
rect 16332 10554 16384 10606
rect 16384 10554 16388 10606
rect 16332 10552 16388 10554
rect 16412 10606 16468 10608
rect 16412 10554 16464 10606
rect 16464 10554 16468 10606
rect 16412 10552 16468 10554
rect 16492 10606 16548 10608
rect 16492 10554 16544 10606
rect 16544 10554 16548 10606
rect 16492 10552 16548 10554
rect 16572 10606 16628 10608
rect 16572 10554 16624 10606
rect 16624 10554 16628 10606
rect 16572 10552 16628 10554
rect 16652 10606 16708 10608
rect 16652 10554 16704 10606
rect 16704 10554 16708 10606
rect 16652 10552 16708 10554
rect 16732 10606 16788 10608
rect 16732 10554 16784 10606
rect 16784 10554 16788 10606
rect 16732 10552 16788 10554
rect 16936 10606 16992 10608
rect 16936 10554 16940 10606
rect 16940 10554 16992 10606
rect 16936 10552 16992 10554
rect 17016 10606 17072 10608
rect 17016 10554 17020 10606
rect 17020 10554 17072 10606
rect 17016 10552 17072 10554
rect 17096 10606 17152 10608
rect 17096 10554 17100 10606
rect 17100 10554 17152 10606
rect 17096 10552 17152 10554
rect 17176 10606 17232 10608
rect 17176 10554 17180 10606
rect 17180 10554 17232 10606
rect 17176 10552 17232 10554
rect 17256 10606 17312 10608
rect 17256 10554 17260 10606
rect 17260 10554 17312 10606
rect 17256 10552 17312 10554
rect 17336 10606 17392 10608
rect 17336 10554 17340 10606
rect 17340 10554 17392 10606
rect 17336 10552 17392 10554
rect 17544 10606 17600 10608
rect 17544 10554 17596 10606
rect 17596 10554 17600 10606
rect 17544 10552 17600 10554
rect 17624 10606 17680 10608
rect 17624 10554 17676 10606
rect 17676 10554 17680 10606
rect 17624 10552 17680 10554
rect 17704 10606 17760 10608
rect 17704 10554 17756 10606
rect 17756 10554 17760 10606
rect 17704 10552 17760 10554
rect 17784 10606 17840 10608
rect 17784 10554 17836 10606
rect 17836 10554 17840 10606
rect 17784 10552 17840 10554
rect 17864 10606 17920 10608
rect 17864 10554 17916 10606
rect 17916 10554 17920 10606
rect 17864 10552 17920 10554
rect 17944 10606 18000 10608
rect 17944 10554 17996 10606
rect 17996 10554 18000 10606
rect 17944 10552 18000 10554
rect 18281 10550 18337 10552
rect 18281 10498 18283 10550
rect 18283 10498 18335 10550
rect 18335 10498 18337 10550
rect 18281 10496 18337 10498
rect 18286 10406 18342 10408
rect 18286 10354 18288 10406
rect 18288 10354 18340 10406
rect 18340 10354 18342 10406
rect 18286 10352 18342 10354
rect 18287 10254 18343 10256
rect 18287 10202 18289 10254
rect 18289 10202 18341 10254
rect 18341 10202 18343 10254
rect 18287 10200 18343 10202
rect 18287 10084 18343 10086
rect 18287 10032 18289 10084
rect 18289 10032 18341 10084
rect 18341 10032 18343 10084
rect 18287 10030 18343 10032
rect 11855 10007 11911 10009
rect 11855 9955 11857 10007
rect 11857 9955 11909 10007
rect 11909 9955 11911 10007
rect 11855 9953 11911 9955
rect 11986 10006 12042 10008
rect 11986 9954 11988 10006
rect 11988 9954 12040 10006
rect 12040 9954 12042 10006
rect 11986 9952 12042 9954
rect 12130 10007 12186 10009
rect 12130 9955 12132 10007
rect 12132 9955 12184 10007
rect 12184 9955 12186 10007
rect 12130 9953 12186 9955
rect 18286 9927 18342 9929
rect 18286 9875 18288 9927
rect 18288 9875 18340 9927
rect 18340 9875 18342 9927
rect 18286 9873 18342 9875
rect 18204 9685 18260 9687
rect 18204 9633 18206 9685
rect 18206 9633 18258 9685
rect 18258 9633 18260 9685
rect 18204 9631 18260 9633
rect 18581 9693 18637 9695
rect 18581 9641 18583 9693
rect 18583 9641 18635 9693
rect 18635 9641 18637 9693
rect 18581 9639 18637 9641
rect 18781 9693 18837 9695
rect 18781 9641 18783 9693
rect 18783 9641 18835 9693
rect 18835 9641 18837 9693
rect 18781 9639 18837 9641
rect 11873 9461 11929 9463
rect 11873 9409 11875 9461
rect 11875 9409 11927 9461
rect 11927 9409 11929 9461
rect 11873 9407 11929 9409
rect 11993 9461 12049 9463
rect 11993 9409 11995 9461
rect 11995 9409 12047 9461
rect 12047 9409 12049 9461
rect 11993 9407 12049 9409
rect 12136 9461 12192 9463
rect 12136 9409 12138 9461
rect 12138 9409 12190 9461
rect 12190 9409 12192 9461
rect 12136 9407 12192 9409
rect 12954 9361 13018 9425
rect 13686 9364 13750 9428
rect 13914 9364 13978 9428
rect 14898 9364 14962 9428
rect 15126 9364 15190 9428
rect 16110 9364 16174 9428
rect 16338 9364 16402 9428
rect 17322 9364 17386 9428
rect 17550 9364 17614 9428
rect 18292 9424 18348 9426
rect 18292 9372 18294 9424
rect 18294 9372 18346 9424
rect 18346 9372 18348 9424
rect 18292 9370 18348 9372
rect 13310 9162 13374 9226
rect 14042 9162 14106 9226
rect 14260 9162 14324 9226
rect 15254 9162 15318 9226
rect 15472 9162 15536 9226
rect 16592 9162 16656 9226
rect 16810 9162 16874 9226
rect 17544 9162 17608 9226
rect 18292 9221 18348 9223
rect 18292 9169 18294 9221
rect 18294 9169 18346 9221
rect 18346 9169 18348 9221
rect 18292 9167 18348 9169
rect 18392 9051 18448 9053
rect 18392 8999 18394 9051
rect 18394 8999 18446 9051
rect 18446 8999 18448 9051
rect 18392 8997 18448 8999
rect 18201 8959 18257 8961
rect 18201 8907 18203 8959
rect 18203 8907 18255 8959
rect 18255 8907 18257 8959
rect 18201 8905 18257 8907
rect 12458 8034 12514 8036
rect 12458 7982 12460 8034
rect 12460 7982 12512 8034
rect 12512 7982 12514 8034
rect 12458 7980 12514 7982
rect 13000 8037 13056 8039
rect 13000 7985 13002 8037
rect 13002 7985 13054 8037
rect 13054 7985 13056 8037
rect 13000 7983 13056 7985
rect 13080 8037 13136 8039
rect 13080 7985 13082 8037
rect 13082 7985 13134 8037
rect 13134 7985 13136 8037
rect 13080 7983 13136 7985
rect 13160 8037 13216 8039
rect 13160 7985 13162 8037
rect 13162 7985 13214 8037
rect 13214 7985 13216 8037
rect 13160 7983 13216 7985
rect 13240 8037 13296 8039
rect 13240 7985 13242 8037
rect 13242 7985 13294 8037
rect 13294 7985 13296 8037
rect 13240 7983 13296 7985
rect 13732 8037 13788 8039
rect 13732 7985 13734 8037
rect 13734 7985 13786 8037
rect 13786 7985 13788 8037
rect 13732 7983 13788 7985
rect 13812 8037 13868 8039
rect 13812 7985 13814 8037
rect 13814 7985 13866 8037
rect 13866 7985 13868 8037
rect 13812 7983 13868 7985
rect 13892 8037 13948 8039
rect 13892 7985 13894 8037
rect 13894 7985 13946 8037
rect 13946 7985 13948 8037
rect 13892 7983 13948 7985
rect 13972 8037 14028 8039
rect 13972 7985 13974 8037
rect 13974 7985 14026 8037
rect 14026 7985 14028 8037
rect 13972 7983 14028 7985
rect 14338 8037 14394 8039
rect 14338 7985 14340 8037
rect 14340 7985 14392 8037
rect 14392 7985 14394 8037
rect 14338 7983 14394 7985
rect 14418 8037 14474 8039
rect 14418 7985 14420 8037
rect 14420 7985 14472 8037
rect 14472 7985 14474 8037
rect 14418 7983 14474 7985
rect 14498 8037 14554 8039
rect 14498 7985 14500 8037
rect 14500 7985 14552 8037
rect 14552 7985 14554 8037
rect 14498 7983 14554 7985
rect 14578 8037 14634 8039
rect 14578 7985 14580 8037
rect 14580 7985 14632 8037
rect 14632 7985 14634 8037
rect 14578 7983 14634 7985
rect 14944 8037 15000 8039
rect 14944 7985 14946 8037
rect 14946 7985 14998 8037
rect 14998 7985 15000 8037
rect 14944 7983 15000 7985
rect 15024 8037 15080 8039
rect 15024 7985 15026 8037
rect 15026 7985 15078 8037
rect 15078 7985 15080 8037
rect 15024 7983 15080 7985
rect 15104 8037 15160 8039
rect 15104 7985 15106 8037
rect 15106 7985 15158 8037
rect 15158 7985 15160 8037
rect 15104 7983 15160 7985
rect 15184 8037 15240 8039
rect 15184 7985 15186 8037
rect 15186 7985 15238 8037
rect 15238 7985 15240 8037
rect 15184 7983 15240 7985
rect 15550 8037 15606 8039
rect 15550 7985 15552 8037
rect 15552 7985 15604 8037
rect 15604 7985 15606 8037
rect 15550 7983 15606 7985
rect 15630 8037 15686 8039
rect 15630 7985 15632 8037
rect 15632 7985 15684 8037
rect 15684 7985 15686 8037
rect 15630 7983 15686 7985
rect 15710 8037 15766 8039
rect 15710 7985 15712 8037
rect 15712 7985 15764 8037
rect 15764 7985 15766 8037
rect 15710 7983 15766 7985
rect 15790 8037 15846 8039
rect 15790 7985 15792 8037
rect 15792 7985 15844 8037
rect 15844 7985 15846 8037
rect 15790 7983 15846 7985
rect 16282 8037 16338 8039
rect 16282 7985 16284 8037
rect 16284 7985 16336 8037
rect 16336 7985 16338 8037
rect 16282 7983 16338 7985
rect 16362 8037 16418 8039
rect 16362 7985 16364 8037
rect 16364 7985 16416 8037
rect 16416 7985 16418 8037
rect 16362 7983 16418 7985
rect 16442 8037 16498 8039
rect 16442 7985 16444 8037
rect 16444 7985 16496 8037
rect 16496 7985 16498 8037
rect 16442 7983 16498 7985
rect 16522 8037 16578 8039
rect 16522 7985 16524 8037
rect 16524 7985 16576 8037
rect 16576 7985 16578 8037
rect 16522 7983 16578 7985
rect 16888 8037 16944 8039
rect 16888 7985 16890 8037
rect 16890 7985 16942 8037
rect 16942 7985 16944 8037
rect 16888 7983 16944 7985
rect 16968 8037 17024 8039
rect 16968 7985 16970 8037
rect 16970 7985 17022 8037
rect 17022 7985 17024 8037
rect 16968 7983 17024 7985
rect 17048 8037 17104 8039
rect 17048 7985 17050 8037
rect 17050 7985 17102 8037
rect 17102 7985 17104 8037
rect 17048 7983 17104 7985
rect 17128 8037 17184 8039
rect 17128 7985 17130 8037
rect 17130 7985 17182 8037
rect 17182 7985 17184 8037
rect 17128 7983 17184 7985
rect 17622 8037 17678 8039
rect 17622 7985 17624 8037
rect 17624 7985 17676 8037
rect 17676 7985 17678 8037
rect 17622 7983 17678 7985
rect 17702 8037 17758 8039
rect 17702 7985 17704 8037
rect 17704 7985 17756 8037
rect 17756 7985 17758 8037
rect 17702 7983 17758 7985
rect 17782 8037 17838 8039
rect 17782 7985 17784 8037
rect 17784 7985 17836 8037
rect 17836 7985 17838 8037
rect 17782 7983 17838 7985
rect 17862 8037 17918 8039
rect 17862 7985 17864 8037
rect 17864 7985 17916 8037
rect 17916 7985 17918 8037
rect 17862 7983 17918 7985
rect 13505 7589 13561 7591
rect 13505 7537 13507 7589
rect 13507 7537 13559 7589
rect 13559 7537 13561 7589
rect 13505 7535 13561 7537
rect 13679 7588 13735 7590
rect 13679 7536 13681 7588
rect 13681 7536 13733 7588
rect 13733 7536 13735 7588
rect 13679 7534 13735 7536
rect 13904 7590 13960 7592
rect 13904 7538 13906 7590
rect 13906 7538 13958 7590
rect 13958 7538 13960 7590
rect 13904 7536 13960 7538
rect 14105 7592 14161 7594
rect 14105 7540 14107 7592
rect 14107 7540 14159 7592
rect 14159 7540 14161 7592
rect 14105 7538 14161 7540
rect 14328 7590 14384 7592
rect 14328 7538 14330 7590
rect 14330 7538 14382 7590
rect 14382 7538 14384 7590
rect 14328 7536 14384 7538
rect 14537 7595 14593 7597
rect 14537 7543 14539 7595
rect 14539 7543 14591 7595
rect 14591 7543 14593 7595
rect 14537 7541 14593 7543
rect 14765 7588 14821 7590
rect 14765 7536 14767 7588
rect 14767 7536 14819 7588
rect 14819 7536 14821 7588
rect 14765 7534 14821 7536
rect 14955 7592 15011 7594
rect 14955 7540 14957 7592
rect 14957 7540 15009 7592
rect 15009 7540 15011 7592
rect 14955 7538 15011 7540
rect 15160 7595 15216 7597
rect 15160 7543 15162 7595
rect 15162 7543 15214 7595
rect 15214 7543 15216 7595
rect 15160 7541 15216 7543
rect 15359 7595 15415 7597
rect 15359 7543 15361 7595
rect 15361 7543 15413 7595
rect 15413 7543 15415 7595
rect 15359 7541 15415 7543
rect 15575 7590 15631 7592
rect 15575 7538 15577 7590
rect 15577 7538 15629 7590
rect 15629 7538 15631 7590
rect 15575 7536 15631 7538
rect 14863 7402 14919 7404
rect 14863 7350 14865 7402
rect 14865 7350 14917 7402
rect 14917 7350 14919 7402
rect 14863 7348 14919 7350
rect 15248 7351 15304 7353
rect 15248 7299 15250 7351
rect 15250 7299 15302 7351
rect 15302 7299 15304 7351
rect 15248 7297 15304 7299
rect 15963 7595 16019 7597
rect 15963 7543 15965 7595
rect 15965 7543 16017 7595
rect 16017 7543 16019 7595
rect 15963 7541 16019 7543
rect 16198 7590 16254 7592
rect 16198 7538 16200 7590
rect 16200 7538 16252 7590
rect 16252 7538 16254 7590
rect 16198 7536 16254 7538
rect 16440 7592 16496 7594
rect 16440 7540 16442 7592
rect 16442 7540 16494 7592
rect 16494 7540 16496 7592
rect 16440 7538 16496 7540
rect 16672 7593 16728 7595
rect 16672 7541 16674 7593
rect 16674 7541 16726 7593
rect 16726 7541 16728 7593
rect 16672 7539 16728 7541
rect 16901 7596 16957 7598
rect 16901 7544 16903 7596
rect 16903 7544 16955 7596
rect 16955 7544 16957 7596
rect 16901 7542 16957 7544
rect 17150 7588 17206 7590
rect 17150 7536 17152 7588
rect 17152 7536 17204 7588
rect 17204 7536 17206 7588
rect 17150 7534 17206 7536
rect 17368 7592 17424 7594
rect 17368 7540 17370 7592
rect 17370 7540 17422 7592
rect 17422 7540 17424 7592
rect 17368 7538 17424 7540
rect 17597 7588 17653 7590
rect 17597 7536 17599 7588
rect 17599 7536 17651 7588
rect 17651 7536 17653 7588
rect 17597 7534 17653 7536
rect 17818 7590 17874 7592
rect 17818 7538 17820 7590
rect 17820 7538 17872 7590
rect 17872 7538 17874 7590
rect 17818 7536 17874 7538
rect 18034 7595 18090 7597
rect 18034 7543 18036 7595
rect 18036 7543 18088 7595
rect 18088 7543 18090 7595
rect 18034 7541 18090 7543
rect 17258 7401 17314 7403
rect 17258 7349 17260 7401
rect 17260 7349 17312 7401
rect 17312 7349 17314 7401
rect 17258 7347 17314 7349
rect 17643 7352 17699 7354
rect 17643 7300 17645 7352
rect 17645 7300 17697 7352
rect 17697 7300 17699 7352
rect 17643 7298 17699 7300
rect 13507 7006 13563 7008
rect 13507 6954 13509 7006
rect 13509 6954 13561 7006
rect 13561 6954 13563 7006
rect 13507 6952 13563 6954
rect 13682 7004 13738 7006
rect 13682 6952 13684 7004
rect 13684 6952 13736 7004
rect 13736 6952 13738 7004
rect 13682 6950 13738 6952
rect 13879 7006 13935 7008
rect 13879 6954 13881 7006
rect 13881 6954 13933 7006
rect 13933 6954 13935 7006
rect 13879 6952 13935 6954
rect 14098 7009 14154 7011
rect 14098 6957 14100 7009
rect 14100 6957 14152 7009
rect 14152 6957 14154 7009
rect 14098 6955 14154 6957
rect 14330 7005 14386 7007
rect 14330 6953 14332 7005
rect 14332 6953 14384 7005
rect 14384 6953 14386 7005
rect 14330 6951 14386 6953
rect 14554 7012 14610 7014
rect 14554 6960 14556 7012
rect 14556 6960 14608 7012
rect 14608 6960 14610 7012
rect 14554 6958 14610 6960
rect 14766 7000 14822 7002
rect 14766 6948 14768 7000
rect 14768 6948 14820 7000
rect 14820 6948 14822 7000
rect 14766 6946 14822 6948
rect 14988 6996 15044 6998
rect 14988 6944 14990 6996
rect 14990 6944 15042 6996
rect 15042 6944 15044 6996
rect 14988 6942 15044 6944
rect 15211 6993 15267 6995
rect 15211 6941 15213 6993
rect 15213 6941 15265 6993
rect 15265 6941 15267 6993
rect 15211 6939 15267 6941
rect 15421 6993 15477 6995
rect 15421 6941 15423 6993
rect 15423 6941 15475 6993
rect 15475 6941 15477 6993
rect 15421 6939 15477 6941
rect 15634 6993 15690 6995
rect 15634 6941 15636 6993
rect 15636 6941 15688 6993
rect 15688 6941 15690 6993
rect 15634 6939 15690 6941
rect 15951 6986 16007 6988
rect 15951 6934 15953 6986
rect 15953 6934 16005 6986
rect 16005 6934 16007 6986
rect 15951 6932 16007 6934
rect 16153 6989 16209 6991
rect 16153 6937 16155 6989
rect 16155 6937 16207 6989
rect 16207 6937 16209 6989
rect 16153 6935 16209 6937
rect 16354 6990 16410 6992
rect 16354 6938 16356 6990
rect 16356 6938 16408 6990
rect 16408 6938 16410 6990
rect 16354 6936 16410 6938
rect 16533 6991 16589 6993
rect 16533 6939 16535 6991
rect 16535 6939 16587 6991
rect 16587 6939 16589 6991
rect 16533 6937 16589 6939
rect 16725 6995 16781 6997
rect 16725 6943 16727 6995
rect 16727 6943 16779 6995
rect 16779 6943 16781 6995
rect 16725 6941 16781 6943
rect 16910 6992 16966 6994
rect 16910 6940 16912 6992
rect 16912 6940 16964 6992
rect 16964 6940 16966 6992
rect 16910 6938 16966 6940
rect 13534 6357 13590 6359
rect 13534 6305 13536 6357
rect 13536 6305 13588 6357
rect 13588 6305 13590 6357
rect 13534 6303 13590 6305
rect 13750 6362 13806 6364
rect 13750 6310 13752 6362
rect 13752 6310 13804 6362
rect 13804 6310 13806 6362
rect 13750 6308 13806 6310
rect 13956 6363 14012 6365
rect 13956 6311 13958 6363
rect 13958 6311 14010 6363
rect 14010 6311 14012 6363
rect 13956 6309 14012 6311
rect 14158 6355 14214 6357
rect 14158 6303 14160 6355
rect 14160 6303 14212 6355
rect 14212 6303 14214 6355
rect 14158 6301 14214 6303
rect 14354 6357 14410 6359
rect 14354 6305 14356 6357
rect 14356 6305 14408 6357
rect 14408 6305 14410 6357
rect 14354 6303 14410 6305
rect 14579 6359 14635 6361
rect 14579 6307 14581 6359
rect 14581 6307 14633 6359
rect 14633 6307 14635 6359
rect 14579 6305 14635 6307
rect 14794 6355 14850 6357
rect 14794 6303 14796 6355
rect 14796 6303 14848 6355
rect 14848 6303 14850 6355
rect 14794 6301 14850 6303
rect 15029 6355 15085 6357
rect 15029 6303 15031 6355
rect 15031 6303 15083 6355
rect 15083 6303 15085 6355
rect 15029 6301 15085 6303
rect 15237 6358 15293 6360
rect 15237 6306 15239 6358
rect 15239 6306 15291 6358
rect 15291 6306 15293 6358
rect 15237 6304 15293 6306
rect 15479 6358 15535 6360
rect 15479 6306 15481 6358
rect 15481 6306 15533 6358
rect 15533 6306 15535 6358
rect 15479 6304 15535 6306
rect 15677 6359 15733 6361
rect 15677 6307 15679 6359
rect 15679 6307 15731 6359
rect 15731 6307 15733 6359
rect 15677 6305 15733 6307
rect 14868 6128 14924 6130
rect 14868 6076 14870 6128
rect 14870 6076 14922 6128
rect 14922 6076 14924 6128
rect 14868 6074 14924 6076
rect 15251 6069 15307 6071
rect 15251 6017 15253 6069
rect 15253 6017 15305 6069
rect 15305 6017 15307 6069
rect 15251 6015 15307 6017
rect 17142 6991 17198 6993
rect 17142 6939 17144 6991
rect 17144 6939 17196 6991
rect 17196 6939 17198 6991
rect 17142 6937 17198 6939
rect 17347 6993 17403 6995
rect 17347 6941 17349 6993
rect 17349 6941 17401 6993
rect 17401 6941 17403 6993
rect 17347 6939 17403 6941
rect 17553 6995 17609 6997
rect 17553 6943 17555 6995
rect 17555 6943 17607 6995
rect 17607 6943 17609 6995
rect 17553 6941 17609 6943
rect 17761 7002 17817 7004
rect 17761 6950 17763 7002
rect 17763 6950 17815 7002
rect 17815 6950 17817 7002
rect 17761 6948 17817 6950
rect 17983 7003 18039 7005
rect 17983 6951 17985 7003
rect 17985 6951 18037 7003
rect 18037 6951 18039 7003
rect 17983 6949 18039 6951
rect 15984 6359 16040 6361
rect 15984 6307 15986 6359
rect 15986 6307 16038 6359
rect 16038 6307 16040 6359
rect 15984 6305 16040 6307
rect 16209 6360 16265 6362
rect 16209 6308 16211 6360
rect 16211 6308 16263 6360
rect 16263 6308 16265 6360
rect 16209 6306 16265 6308
rect 16438 6359 16494 6361
rect 16438 6307 16440 6359
rect 16440 6307 16492 6359
rect 16492 6307 16494 6359
rect 16438 6305 16494 6307
rect 16654 6363 16710 6365
rect 16654 6311 16656 6363
rect 16656 6311 16708 6363
rect 16708 6311 16710 6363
rect 16654 6309 16710 6311
rect 16877 6366 16933 6368
rect 16877 6314 16879 6366
rect 16879 6314 16931 6366
rect 16931 6314 16933 6366
rect 16877 6312 16933 6314
rect 17101 6362 17157 6364
rect 17101 6310 17103 6362
rect 17103 6310 17155 6362
rect 17155 6310 17157 6362
rect 17101 6308 17157 6310
rect 17328 6351 17384 6353
rect 17328 6299 17330 6351
rect 17330 6299 17382 6351
rect 17382 6299 17384 6351
rect 17328 6297 17384 6299
rect 17541 6350 17597 6352
rect 17541 6298 17543 6350
rect 17543 6298 17595 6350
rect 17595 6298 17597 6350
rect 17541 6296 17597 6298
rect 17752 6354 17808 6356
rect 17752 6302 17754 6354
rect 17754 6302 17806 6354
rect 17806 6302 17808 6354
rect 17752 6300 17808 6302
rect 17979 6355 18035 6357
rect 17979 6303 17981 6355
rect 17981 6303 18033 6355
rect 18033 6303 18035 6355
rect 17979 6301 18035 6303
rect 17260 6130 17316 6132
rect 17260 6078 17262 6130
rect 17262 6078 17314 6130
rect 17314 6078 17316 6130
rect 17260 6076 17316 6078
rect 17637 6076 17693 6078
rect 17637 6024 17639 6076
rect 17639 6024 17691 6076
rect 17691 6024 17693 6076
rect 17637 6022 17693 6024
rect 13560 5712 13616 5714
rect 13560 5660 13562 5712
rect 13562 5660 13614 5712
rect 13614 5660 13616 5712
rect 13560 5658 13616 5660
rect 13785 5721 13841 5723
rect 13785 5669 13787 5721
rect 13787 5669 13839 5721
rect 13839 5669 13841 5721
rect 13785 5667 13841 5669
rect 14062 5718 14118 5720
rect 14062 5666 14064 5718
rect 14064 5666 14116 5718
rect 14116 5666 14118 5718
rect 14062 5664 14118 5666
rect 14283 5721 14339 5723
rect 14283 5669 14285 5721
rect 14285 5669 14337 5721
rect 14337 5669 14339 5721
rect 14283 5667 14339 5669
rect 14528 5718 14584 5720
rect 14528 5666 14530 5718
rect 14530 5666 14582 5718
rect 14582 5666 14584 5718
rect 14528 5664 14584 5666
rect 14754 5722 14810 5724
rect 14754 5670 14756 5722
rect 14756 5670 14808 5722
rect 14808 5670 14810 5722
rect 14754 5668 14810 5670
rect 14966 5720 15022 5722
rect 14966 5668 14968 5720
rect 14968 5668 15020 5720
rect 15020 5668 15022 5720
rect 14966 5666 15022 5668
rect 15186 5726 15242 5728
rect 15186 5674 15188 5726
rect 15188 5674 15240 5726
rect 15240 5674 15242 5726
rect 15186 5672 15242 5674
rect 15424 5728 15480 5730
rect 15424 5676 15426 5728
rect 15426 5676 15478 5728
rect 15478 5676 15480 5728
rect 15424 5674 15480 5676
rect 15637 5730 15693 5732
rect 15637 5678 15639 5730
rect 15639 5678 15691 5730
rect 15691 5678 15693 5730
rect 15637 5676 15693 5678
rect 16024 5720 16080 5722
rect 16024 5668 16026 5720
rect 16026 5668 16078 5720
rect 16078 5668 16080 5720
rect 16024 5666 16080 5668
rect 16371 5721 16427 5723
rect 16371 5669 16373 5721
rect 16373 5669 16425 5721
rect 16425 5669 16427 5721
rect 16371 5667 16427 5669
rect 17030 5718 17086 5720
rect 16607 5716 16663 5718
rect 16607 5664 16609 5716
rect 16609 5664 16661 5716
rect 16661 5664 16663 5716
rect 16607 5662 16663 5664
rect 16791 5716 16847 5718
rect 16791 5664 16793 5716
rect 16793 5664 16845 5716
rect 16845 5664 16847 5716
rect 17030 5666 17032 5718
rect 17032 5666 17084 5718
rect 17084 5666 17086 5718
rect 17030 5664 17086 5666
rect 16791 5662 16847 5664
rect 17233 5714 17289 5716
rect 17233 5662 17235 5714
rect 17235 5662 17287 5714
rect 17287 5662 17289 5714
rect 17233 5660 17289 5662
rect 17418 5711 17474 5713
rect 17418 5659 17420 5711
rect 17420 5659 17472 5711
rect 17472 5659 17474 5711
rect 17418 5657 17474 5659
rect 17609 5713 17665 5715
rect 17609 5661 17611 5713
rect 17611 5661 17663 5713
rect 17663 5661 17665 5713
rect 17609 5659 17665 5661
rect 17800 5717 17856 5719
rect 17800 5665 17802 5717
rect 17802 5665 17854 5717
rect 17854 5665 17856 5717
rect 17800 5663 17856 5665
rect 17986 5713 18042 5715
rect 17986 5661 17988 5713
rect 17988 5661 18040 5713
rect 18040 5661 18042 5713
rect 17986 5659 18042 5661
rect 13433 5130 13489 5132
rect 13433 5078 13435 5130
rect 13435 5078 13487 5130
rect 13487 5078 13489 5130
rect 13433 5076 13489 5078
rect 13638 5126 13694 5128
rect 13638 5074 13640 5126
rect 13640 5074 13692 5126
rect 13692 5074 13694 5126
rect 13638 5072 13694 5074
rect 13824 5131 13880 5133
rect 13824 5079 13826 5131
rect 13826 5079 13878 5131
rect 13878 5079 13880 5131
rect 13824 5077 13880 5079
rect 14018 5124 14074 5126
rect 14018 5072 14020 5124
rect 14020 5072 14072 5124
rect 14072 5072 14074 5124
rect 14018 5070 14074 5072
rect 14237 5129 14293 5131
rect 14237 5077 14239 5129
rect 14239 5077 14291 5129
rect 14291 5077 14293 5129
rect 14237 5075 14293 5077
rect 14447 5129 14503 5131
rect 14447 5077 14449 5129
rect 14449 5077 14501 5129
rect 14501 5077 14503 5129
rect 14447 5075 14503 5077
rect 14676 5126 14732 5128
rect 14676 5074 14678 5126
rect 14678 5074 14730 5126
rect 14730 5074 14732 5126
rect 14676 5072 14732 5074
rect 14922 5126 14978 5128
rect 14922 5074 14924 5126
rect 14924 5074 14976 5126
rect 14976 5074 14978 5126
rect 14922 5072 14978 5074
rect 15196 5126 15252 5128
rect 15196 5074 15198 5126
rect 15198 5074 15250 5126
rect 15250 5074 15252 5126
rect 15196 5072 15252 5074
rect 15471 5126 15527 5128
rect 15471 5074 15473 5126
rect 15473 5074 15525 5126
rect 15525 5074 15527 5126
rect 15471 5072 15527 5074
rect 15707 5126 15763 5128
rect 15707 5074 15709 5126
rect 15709 5074 15761 5126
rect 15761 5074 15763 5126
rect 15707 5072 15763 5074
rect 15930 5129 15986 5131
rect 15930 5077 15932 5129
rect 15932 5077 15984 5129
rect 15984 5077 15986 5129
rect 15930 5075 15986 5077
rect 16148 5132 16204 5134
rect 16148 5080 16150 5132
rect 16150 5080 16202 5132
rect 16202 5080 16204 5132
rect 16148 5078 16204 5080
rect 16326 5123 16382 5125
rect 16326 5071 16328 5123
rect 16328 5071 16380 5123
rect 16380 5071 16382 5123
rect 16326 5069 16382 5071
rect 16565 5125 16621 5127
rect 16565 5073 16567 5125
rect 16567 5073 16619 5125
rect 16619 5073 16621 5125
rect 16565 5071 16621 5073
rect 16762 5125 16818 5127
rect 16762 5073 16764 5125
rect 16764 5073 16816 5125
rect 16816 5073 16818 5125
rect 16762 5071 16818 5073
rect 16960 5125 17016 5127
rect 16960 5073 16962 5125
rect 16962 5073 17014 5125
rect 17014 5073 17016 5125
rect 16960 5071 17016 5073
rect 17173 5126 17229 5128
rect 17173 5074 17175 5126
rect 17175 5074 17227 5126
rect 17227 5074 17229 5126
rect 17173 5072 17229 5074
rect 17396 5125 17452 5127
rect 17396 5073 17398 5125
rect 17398 5073 17450 5125
rect 17450 5073 17452 5125
rect 17396 5071 17452 5073
rect 17593 5130 17649 5132
rect 17593 5078 17595 5130
rect 17595 5078 17647 5130
rect 17647 5078 17649 5130
rect 17593 5076 17649 5078
rect 17809 5128 17865 5130
rect 17809 5076 17811 5128
rect 17811 5076 17863 5128
rect 17863 5076 17865 5128
rect 17809 5074 17865 5076
rect 18018 5128 18074 5130
rect 18018 5076 18020 5128
rect 18020 5076 18072 5128
rect 18072 5076 18074 5128
rect 18018 5074 18074 5076
<< metal3 >>
rect 12437 10618 12563 10628
rect 12437 10554 12468 10618
rect 12532 10610 12563 10618
rect 13193 10611 18107 10613
rect 12532 10608 13133 10610
rect 12532 10554 12565 10608
rect 12437 10545 12565 10554
rect 12461 10544 12565 10545
rect 12629 10544 12645 10608
rect 12709 10544 12725 10608
rect 12789 10544 12805 10608
rect 12869 10544 12885 10608
rect 12949 10544 12965 10608
rect 13029 10544 13133 10608
rect 13193 10547 13297 10611
rect 13361 10547 13377 10611
rect 13441 10547 13457 10611
rect 13521 10547 13537 10611
rect 13601 10547 13617 10611
rect 13681 10547 13697 10611
rect 13761 10547 13903 10611
rect 13967 10547 13983 10611
rect 14047 10547 14063 10611
rect 14127 10547 14143 10611
rect 14207 10547 14223 10611
rect 14287 10547 14303 10611
rect 14367 10547 14509 10611
rect 14573 10547 14589 10611
rect 14653 10547 14669 10611
rect 14733 10547 14749 10611
rect 14813 10547 14829 10611
rect 14893 10547 14909 10611
rect 14973 10547 15115 10611
rect 15179 10547 15195 10611
rect 15259 10547 15275 10611
rect 15339 10547 15355 10611
rect 15419 10547 15435 10611
rect 15499 10547 15515 10611
rect 15579 10547 15721 10611
rect 15785 10547 15801 10611
rect 15865 10547 15881 10611
rect 15945 10547 15961 10611
rect 16025 10547 16041 10611
rect 16105 10547 16121 10611
rect 16185 10547 16327 10611
rect 16391 10547 16407 10611
rect 16471 10547 16487 10611
rect 16551 10547 16567 10611
rect 16631 10547 16647 10611
rect 16711 10547 16727 10611
rect 16791 10547 16933 10611
rect 16997 10547 17013 10611
rect 17077 10547 17093 10611
rect 17157 10547 17173 10611
rect 17237 10547 17253 10611
rect 17317 10547 17333 10611
rect 17397 10547 17539 10611
rect 17603 10547 17619 10611
rect 17683 10547 17699 10611
rect 17763 10547 17779 10611
rect 17843 10547 17859 10611
rect 17923 10547 17939 10611
rect 18003 10547 18107 10611
rect 13193 10545 18107 10547
rect 18246 10556 18372 10566
rect 12461 10542 13133 10544
rect 12461 10388 12527 10478
rect 12461 10324 12462 10388
rect 12526 10324 12527 10388
rect 12461 10308 12527 10324
rect 12461 10244 12462 10308
rect 12526 10244 12527 10308
rect 12461 10228 12527 10244
rect 12461 10164 12462 10228
rect 12526 10164 12527 10228
rect 12461 10148 12527 10164
rect 12461 10084 12462 10148
rect 12526 10084 12527 10148
rect 12461 10068 12527 10084
rect 11836 10027 11954 10028
rect 12085 10027 12229 10028
rect 11836 10013 12229 10027
rect 11836 9949 11851 10013
rect 11915 10012 12126 10013
rect 11915 9949 11982 10012
rect 11836 9948 11982 9949
rect 12046 9949 12126 10012
rect 12190 9949 12229 10013
rect 12046 9948 12229 9949
rect 11836 9932 12229 9948
rect 12461 10004 12462 10068
rect 12526 10004 12527 10068
rect 12461 9988 12527 10004
rect 11941 9931 12085 9932
rect 12461 9924 12462 9988
rect 12526 9924 12527 9988
rect 12461 9908 12527 9924
rect 12461 9844 12462 9908
rect 12526 9844 12527 9908
rect 12461 9828 12527 9844
rect 12461 9764 12462 9828
rect 12526 9764 12527 9828
rect 12461 9748 12527 9764
rect 12461 9684 12462 9748
rect 12526 9684 12527 9748
rect 12461 9668 12527 9684
rect 12461 9604 12462 9668
rect 12526 9604 12527 9668
rect 11976 9482 12068 9483
rect 11862 9467 12235 9482
rect 11862 9403 11869 9467
rect 11933 9403 11989 9467
rect 12053 9403 12132 9467
rect 12196 9403 12235 9467
rect 11862 9386 12235 9403
rect 12461 9450 12527 9604
rect 12587 9450 12647 10482
rect 12707 9512 12767 10542
rect 12827 9450 12887 10482
rect 12947 9512 13007 10542
rect 13067 10388 13133 10478
rect 13067 10324 13068 10388
rect 13132 10324 13133 10388
rect 13067 10308 13133 10324
rect 13067 10244 13068 10308
rect 13132 10244 13133 10308
rect 13067 10228 13133 10244
rect 13067 10164 13068 10228
rect 13132 10164 13133 10228
rect 13067 10148 13133 10164
rect 13067 10084 13068 10148
rect 13132 10084 13133 10148
rect 13067 10068 13133 10084
rect 13067 10004 13068 10068
rect 13132 10004 13133 10068
rect 13067 9988 13133 10004
rect 13067 9924 13068 9988
rect 13132 9924 13133 9988
rect 13067 9908 13133 9924
rect 13067 9844 13068 9908
rect 13132 9844 13133 9908
rect 13067 9828 13133 9844
rect 13067 9764 13068 9828
rect 13132 9764 13133 9828
rect 13067 9748 13133 9764
rect 13067 9684 13068 9748
rect 13132 9684 13133 9748
rect 13067 9668 13133 9684
rect 13067 9604 13068 9668
rect 13132 9604 13133 9668
rect 13067 9450 13133 9604
rect 12461 9448 13133 9450
rect 12461 9384 12565 9448
rect 12629 9384 12645 9448
rect 12709 9384 12725 9448
rect 12789 9384 12805 9448
rect 12869 9384 12885 9448
rect 12949 9425 12965 9448
rect 12949 9384 12954 9425
rect 13029 9384 13133 9448
rect 13193 10391 13259 10481
rect 13193 10327 13194 10391
rect 13258 10327 13259 10391
rect 13193 10311 13259 10327
rect 13193 10247 13194 10311
rect 13258 10247 13259 10311
rect 13193 10231 13259 10247
rect 13193 10167 13194 10231
rect 13258 10167 13259 10231
rect 13193 10151 13259 10167
rect 13193 10087 13194 10151
rect 13258 10087 13259 10151
rect 13193 10071 13259 10087
rect 13193 10007 13194 10071
rect 13258 10007 13259 10071
rect 13193 9991 13259 10007
rect 13193 9927 13194 9991
rect 13258 9927 13259 9991
rect 13193 9911 13259 9927
rect 13193 9847 13194 9911
rect 13258 9847 13259 9911
rect 13193 9831 13259 9847
rect 13193 9767 13194 9831
rect 13258 9767 13259 9831
rect 13193 9751 13259 9767
rect 13193 9687 13194 9751
rect 13258 9687 13259 9751
rect 13193 9671 13259 9687
rect 13193 9607 13194 9671
rect 13258 9607 13259 9671
rect 13193 9453 13259 9607
rect 13319 9453 13379 10485
rect 13439 9515 13499 10545
rect 13559 9453 13619 10485
rect 13679 9515 13739 10545
rect 13799 10391 13865 10481
rect 13799 10327 13800 10391
rect 13864 10327 13865 10391
rect 13799 10311 13865 10327
rect 13799 10247 13800 10311
rect 13864 10247 13865 10311
rect 13799 10231 13865 10247
rect 13799 10167 13800 10231
rect 13864 10167 13865 10231
rect 13799 10151 13865 10167
rect 13799 10087 13800 10151
rect 13864 10087 13865 10151
rect 13799 10071 13865 10087
rect 13799 10007 13800 10071
rect 13864 10007 13865 10071
rect 13799 9991 13865 10007
rect 13799 9927 13800 9991
rect 13864 9927 13865 9991
rect 13799 9911 13865 9927
rect 13799 9847 13800 9911
rect 13864 9847 13865 9911
rect 13799 9831 13865 9847
rect 13799 9767 13800 9831
rect 13864 9767 13865 9831
rect 13799 9751 13865 9767
rect 13799 9687 13800 9751
rect 13864 9687 13865 9751
rect 13799 9671 13865 9687
rect 13799 9607 13800 9671
rect 13864 9607 13865 9671
rect 13799 9453 13865 9607
rect 13925 9515 13985 10545
rect 14045 9453 14105 10485
rect 14165 9515 14225 10545
rect 14285 9453 14345 10485
rect 14405 10391 14471 10481
rect 14405 10327 14406 10391
rect 14470 10327 14471 10391
rect 14405 10311 14471 10327
rect 14405 10247 14406 10311
rect 14470 10247 14471 10311
rect 14405 10231 14471 10247
rect 14405 10167 14406 10231
rect 14470 10167 14471 10231
rect 14405 10151 14471 10167
rect 14405 10087 14406 10151
rect 14470 10087 14471 10151
rect 14405 10071 14471 10087
rect 14405 10007 14406 10071
rect 14470 10007 14471 10071
rect 14405 9991 14471 10007
rect 14405 9927 14406 9991
rect 14470 9927 14471 9991
rect 14405 9911 14471 9927
rect 14405 9847 14406 9911
rect 14470 9847 14471 9911
rect 14405 9831 14471 9847
rect 14405 9767 14406 9831
rect 14470 9767 14471 9831
rect 14405 9751 14471 9767
rect 14405 9687 14406 9751
rect 14470 9687 14471 9751
rect 14405 9671 14471 9687
rect 14405 9607 14406 9671
rect 14470 9607 14471 9671
rect 14405 9453 14471 9607
rect 14531 9453 14591 10485
rect 14651 9515 14711 10545
rect 14771 9453 14831 10485
rect 14891 9515 14951 10545
rect 15011 10391 15077 10481
rect 15011 10327 15012 10391
rect 15076 10327 15077 10391
rect 15011 10311 15077 10327
rect 15011 10247 15012 10311
rect 15076 10247 15077 10311
rect 15011 10231 15077 10247
rect 15011 10167 15012 10231
rect 15076 10167 15077 10231
rect 15011 10151 15077 10167
rect 15011 10087 15012 10151
rect 15076 10087 15077 10151
rect 15011 10071 15077 10087
rect 15011 10007 15012 10071
rect 15076 10007 15077 10071
rect 15011 9991 15077 10007
rect 15011 9927 15012 9991
rect 15076 9927 15077 9991
rect 15011 9911 15077 9927
rect 15011 9847 15012 9911
rect 15076 9847 15077 9911
rect 15011 9831 15077 9847
rect 15011 9767 15012 9831
rect 15076 9767 15077 9831
rect 15011 9751 15077 9767
rect 15011 9687 15012 9751
rect 15076 9687 15077 9751
rect 15011 9671 15077 9687
rect 15011 9607 15012 9671
rect 15076 9607 15077 9671
rect 15011 9453 15077 9607
rect 15137 9515 15197 10545
rect 15257 9453 15317 10485
rect 15377 9515 15437 10545
rect 15497 9453 15557 10485
rect 15617 10391 15683 10481
rect 15617 10327 15618 10391
rect 15682 10327 15683 10391
rect 15617 10311 15683 10327
rect 15617 10247 15618 10311
rect 15682 10247 15683 10311
rect 15617 10231 15683 10247
rect 15617 10167 15618 10231
rect 15682 10167 15683 10231
rect 15617 10151 15683 10167
rect 15617 10087 15618 10151
rect 15682 10087 15683 10151
rect 15617 10071 15683 10087
rect 15617 10007 15618 10071
rect 15682 10007 15683 10071
rect 15617 9991 15683 10007
rect 15617 9927 15618 9991
rect 15682 9927 15683 9991
rect 15617 9911 15683 9927
rect 15617 9847 15618 9911
rect 15682 9847 15683 9911
rect 15617 9831 15683 9847
rect 15617 9767 15618 9831
rect 15682 9767 15683 9831
rect 15617 9751 15683 9767
rect 15617 9687 15618 9751
rect 15682 9687 15683 9751
rect 15617 9671 15683 9687
rect 15617 9607 15618 9671
rect 15682 9607 15683 9671
rect 15617 9453 15683 9607
rect 15743 9453 15803 10485
rect 15863 9515 15923 10545
rect 15983 9453 16043 10485
rect 16103 9515 16163 10545
rect 16223 10391 16289 10481
rect 16223 10327 16224 10391
rect 16288 10327 16289 10391
rect 16223 10311 16289 10327
rect 16223 10247 16224 10311
rect 16288 10247 16289 10311
rect 16223 10231 16289 10247
rect 16223 10167 16224 10231
rect 16288 10167 16289 10231
rect 16223 10151 16289 10167
rect 16223 10087 16224 10151
rect 16288 10087 16289 10151
rect 16223 10071 16289 10087
rect 16223 10007 16224 10071
rect 16288 10007 16289 10071
rect 16223 9991 16289 10007
rect 16223 9927 16224 9991
rect 16288 9927 16289 9991
rect 16223 9911 16289 9927
rect 16223 9847 16224 9911
rect 16288 9847 16289 9911
rect 16223 9831 16289 9847
rect 16223 9767 16224 9831
rect 16288 9767 16289 9831
rect 16223 9751 16289 9767
rect 16223 9687 16224 9751
rect 16288 9687 16289 9751
rect 16223 9671 16289 9687
rect 16223 9607 16224 9671
rect 16288 9607 16289 9671
rect 16223 9453 16289 9607
rect 16349 9515 16409 10545
rect 16469 9453 16529 10485
rect 16589 9515 16649 10545
rect 16709 9453 16769 10485
rect 16829 10391 16895 10481
rect 16829 10327 16830 10391
rect 16894 10327 16895 10391
rect 16829 10311 16895 10327
rect 16829 10247 16830 10311
rect 16894 10247 16895 10311
rect 16829 10231 16895 10247
rect 16829 10167 16830 10231
rect 16894 10167 16895 10231
rect 16829 10151 16895 10167
rect 16829 10087 16830 10151
rect 16894 10087 16895 10151
rect 16829 10071 16895 10087
rect 16829 10007 16830 10071
rect 16894 10007 16895 10071
rect 16829 9991 16895 10007
rect 16829 9927 16830 9991
rect 16894 9927 16895 9991
rect 16829 9911 16895 9927
rect 16829 9847 16830 9911
rect 16894 9847 16895 9911
rect 16829 9831 16895 9847
rect 16829 9767 16830 9831
rect 16894 9767 16895 9831
rect 16829 9751 16895 9767
rect 16829 9687 16830 9751
rect 16894 9687 16895 9751
rect 16829 9671 16895 9687
rect 16829 9607 16830 9671
rect 16894 9607 16895 9671
rect 16829 9453 16895 9607
rect 16955 9453 17015 10485
rect 17075 9515 17135 10545
rect 17195 9453 17255 10485
rect 17315 9515 17375 10545
rect 17435 10391 17501 10481
rect 17435 10327 17436 10391
rect 17500 10327 17501 10391
rect 17435 10311 17501 10327
rect 17435 10247 17436 10311
rect 17500 10247 17501 10311
rect 17435 10231 17501 10247
rect 17435 10167 17436 10231
rect 17500 10167 17501 10231
rect 17435 10151 17501 10167
rect 17435 10087 17436 10151
rect 17500 10087 17501 10151
rect 17435 10071 17501 10087
rect 17435 10007 17436 10071
rect 17500 10007 17501 10071
rect 17435 9991 17501 10007
rect 17435 9927 17436 9991
rect 17500 9927 17501 9991
rect 17435 9911 17501 9927
rect 17435 9847 17436 9911
rect 17500 9847 17501 9911
rect 17435 9831 17501 9847
rect 17435 9767 17436 9831
rect 17500 9767 17501 9831
rect 17435 9751 17501 9767
rect 17435 9687 17436 9751
rect 17500 9687 17501 9751
rect 17435 9671 17501 9687
rect 17435 9607 17436 9671
rect 17500 9607 17501 9671
rect 17435 9453 17501 9607
rect 17561 9515 17621 10545
rect 17681 9453 17741 10485
rect 17801 9515 17861 10545
rect 18246 10492 18277 10556
rect 18341 10492 18372 10556
rect 17921 9453 17981 10485
rect 18246 10482 18372 10492
rect 18041 10391 18107 10481
rect 18041 10327 18042 10391
rect 18106 10327 18107 10391
rect 18251 10412 18377 10422
rect 18251 10348 18282 10412
rect 18346 10348 18377 10412
rect 18251 10338 18377 10348
rect 18041 10311 18107 10327
rect 18041 10247 18042 10311
rect 18106 10247 18107 10311
rect 18041 10231 18107 10247
rect 18041 10167 18042 10231
rect 18106 10167 18107 10231
rect 18252 10260 18378 10270
rect 18252 10196 18283 10260
rect 18347 10196 18378 10260
rect 18252 10186 18378 10196
rect 18041 10151 18107 10167
rect 18041 10087 18042 10151
rect 18106 10087 18107 10151
rect 18041 10071 18107 10087
rect 18041 10007 18042 10071
rect 18106 10007 18107 10071
rect 18252 10090 18378 10100
rect 18252 10026 18283 10090
rect 18347 10026 18378 10090
rect 18252 10016 18378 10026
rect 18041 9991 18107 10007
rect 18041 9927 18042 9991
rect 18106 9927 18107 9991
rect 18041 9911 18107 9927
rect 18041 9847 18042 9911
rect 18106 9847 18107 9911
rect 18251 9933 18377 9943
rect 18251 9869 18282 9933
rect 18346 9869 18377 9933
rect 18251 9859 18377 9869
rect 18041 9831 18107 9847
rect 18041 9767 18042 9831
rect 18106 9767 18107 9831
rect 18041 9751 18107 9767
rect 18041 9687 18042 9751
rect 18106 9687 18107 9751
rect 18041 9671 18107 9687
rect 18041 9607 18042 9671
rect 18106 9607 18107 9671
rect 18169 9691 18295 9701
rect 18169 9627 18200 9691
rect 18264 9627 18295 9691
rect 18169 9617 18295 9627
rect 18546 9699 18672 9709
rect 18546 9635 18577 9699
rect 18641 9635 18672 9699
rect 18546 9625 18672 9635
rect 18746 9699 18872 9709
rect 18746 9635 18777 9699
rect 18841 9635 18872 9699
rect 18746 9625 18872 9635
rect 18041 9453 18107 9607
rect 13193 9451 18107 9453
rect 13193 9387 13297 9451
rect 13361 9387 13377 9451
rect 13441 9387 13457 9451
rect 13521 9387 13537 9451
rect 13601 9387 13617 9451
rect 13681 9428 13697 9451
rect 13681 9387 13686 9428
rect 13761 9387 13903 9451
rect 13967 9428 13983 9451
rect 13978 9387 13983 9428
rect 14047 9387 14063 9451
rect 14127 9387 14143 9451
rect 14207 9387 14223 9451
rect 14287 9387 14303 9451
rect 14367 9387 14509 9451
rect 14573 9387 14589 9451
rect 14653 9387 14669 9451
rect 14733 9387 14749 9451
rect 14813 9387 14829 9451
rect 14893 9428 14909 9451
rect 14893 9387 14898 9428
rect 14973 9387 15115 9451
rect 15179 9428 15195 9451
rect 15190 9387 15195 9428
rect 15259 9387 15275 9451
rect 15339 9387 15355 9451
rect 15419 9387 15435 9451
rect 15499 9387 15515 9451
rect 15579 9387 15721 9451
rect 15785 9387 15801 9451
rect 15865 9387 15881 9451
rect 15945 9387 15961 9451
rect 16025 9387 16041 9451
rect 16105 9428 16121 9451
rect 16105 9387 16110 9428
rect 16185 9387 16327 9451
rect 16391 9428 16407 9451
rect 16402 9387 16407 9428
rect 16471 9387 16487 9451
rect 16551 9387 16567 9451
rect 16631 9387 16647 9451
rect 16711 9387 16727 9451
rect 16791 9387 16933 9451
rect 16997 9387 17013 9451
rect 17077 9387 17093 9451
rect 17157 9387 17173 9451
rect 17237 9387 17253 9451
rect 17317 9428 17333 9451
rect 17317 9387 17322 9428
rect 17397 9387 17539 9451
rect 17603 9428 17619 9451
rect 17614 9387 17619 9428
rect 17683 9387 17699 9451
rect 17763 9387 17779 9451
rect 17843 9387 17859 9451
rect 17923 9387 17939 9451
rect 18003 9387 18107 9451
rect 13193 9385 13686 9387
rect 12461 9382 12954 9384
rect 12944 9361 12954 9382
rect 13018 9382 13133 9384
rect 13018 9361 13027 9382
rect 12944 9356 13027 9361
rect 13676 9364 13686 9385
rect 13750 9385 13914 9387
rect 13750 9364 13759 9385
rect 13676 9359 13759 9364
rect 13905 9364 13914 9385
rect 13978 9385 14898 9387
rect 13978 9364 13988 9385
rect 13905 9359 13988 9364
rect 14888 9364 14898 9385
rect 14962 9385 15126 9387
rect 14962 9364 14971 9385
rect 14888 9359 14971 9364
rect 15117 9364 15126 9385
rect 15190 9385 16110 9387
rect 15190 9364 15200 9385
rect 15117 9359 15200 9364
rect 16100 9364 16110 9385
rect 16174 9385 16338 9387
rect 16174 9364 16183 9385
rect 16100 9359 16183 9364
rect 16329 9364 16338 9385
rect 16402 9385 17322 9387
rect 16402 9364 16412 9385
rect 16329 9359 16412 9364
rect 17312 9364 17322 9385
rect 17386 9385 17550 9387
rect 17386 9364 17395 9385
rect 17312 9359 17395 9364
rect 17541 9364 17550 9385
rect 17614 9385 18107 9387
rect 18257 9430 18383 9440
rect 17614 9364 17624 9385
rect 17541 9359 17624 9364
rect 18257 9366 18288 9430
rect 18352 9366 18383 9430
rect 18257 9356 18383 9366
rect 13301 9226 13383 9232
rect 13301 9205 13310 9226
rect 12812 9203 13310 9205
rect 13374 9205 13383 9226
rect 14033 9226 14115 9232
rect 14033 9205 14042 9226
rect 13374 9203 13484 9205
rect 12812 9139 12916 9203
rect 12980 9139 12996 9203
rect 13060 9139 13076 9203
rect 13140 9139 13156 9203
rect 13220 9139 13236 9203
rect 13300 9162 13310 9203
rect 13300 9139 13316 9162
rect 13380 9139 13484 9203
rect 12812 9137 13484 9139
rect 12812 8983 12878 9137
rect 12812 8919 12813 8983
rect 12877 8919 12878 8983
rect 12812 8903 12878 8919
rect 12812 8839 12813 8903
rect 12877 8839 12878 8903
rect 12812 8823 12878 8839
rect 12812 8759 12813 8823
rect 12877 8759 12878 8823
rect 12812 8743 12878 8759
rect 12812 8679 12813 8743
rect 12877 8679 12878 8743
rect 12812 8663 12878 8679
rect 12812 8599 12813 8663
rect 12877 8599 12878 8663
rect 12812 8583 12878 8599
rect 12812 8519 12813 8583
rect 12877 8519 12878 8583
rect 12812 8503 12878 8519
rect 12812 8439 12813 8503
rect 12877 8439 12878 8503
rect 12812 8423 12878 8439
rect 12812 8359 12813 8423
rect 12877 8359 12878 8423
rect 12812 8343 12878 8359
rect 12812 8279 12813 8343
rect 12877 8279 12878 8343
rect 12812 8263 12878 8279
rect 12812 8199 12813 8263
rect 12877 8199 12878 8263
rect 12812 8109 12878 8199
rect 12938 8105 12998 9137
rect 12424 8040 12549 8050
rect 13058 8045 13118 9075
rect 13178 8105 13238 9137
rect 13298 8045 13358 9075
rect 13418 8983 13484 9137
rect 13418 8919 13419 8983
rect 13483 8919 13484 8983
rect 13418 8903 13484 8919
rect 13418 8839 13419 8903
rect 13483 8839 13484 8903
rect 13418 8823 13484 8839
rect 13418 8759 13419 8823
rect 13483 8759 13484 8823
rect 13418 8743 13484 8759
rect 13418 8679 13419 8743
rect 13483 8679 13484 8743
rect 13418 8663 13484 8679
rect 13418 8599 13419 8663
rect 13483 8599 13484 8663
rect 13418 8583 13484 8599
rect 13418 8519 13419 8583
rect 13483 8519 13484 8583
rect 13418 8503 13484 8519
rect 13418 8439 13419 8503
rect 13483 8439 13484 8503
rect 13418 8423 13484 8439
rect 13418 8359 13419 8423
rect 13483 8359 13484 8423
rect 13418 8343 13484 8359
rect 13418 8279 13419 8343
rect 13483 8279 13484 8343
rect 13418 8263 13484 8279
rect 13418 8199 13419 8263
rect 13483 8199 13484 8263
rect 13418 8109 13484 8199
rect 13544 9203 14042 9205
rect 14106 9205 14115 9226
rect 14251 9226 14333 9232
rect 14251 9205 14260 9226
rect 14106 9203 14260 9205
rect 14324 9205 14333 9226
rect 15245 9226 15327 9232
rect 15245 9205 15254 9226
rect 14324 9203 15254 9205
rect 15318 9205 15327 9226
rect 15463 9226 15545 9232
rect 15463 9205 15472 9226
rect 15318 9203 15472 9205
rect 15536 9205 15545 9226
rect 16583 9226 16665 9232
rect 16583 9205 16592 9226
rect 15536 9203 16034 9205
rect 13544 9139 13648 9203
rect 13712 9139 13728 9203
rect 13792 9139 13808 9203
rect 13872 9139 13888 9203
rect 13952 9139 13968 9203
rect 14032 9162 14042 9203
rect 14032 9139 14048 9162
rect 14112 9139 14254 9203
rect 14324 9162 14334 9203
rect 14318 9139 14334 9162
rect 14398 9139 14414 9203
rect 14478 9139 14494 9203
rect 14558 9139 14574 9203
rect 14638 9139 14654 9203
rect 14718 9139 14860 9203
rect 14924 9139 14940 9203
rect 15004 9139 15020 9203
rect 15084 9139 15100 9203
rect 15164 9139 15180 9203
rect 15244 9162 15254 9203
rect 15244 9139 15260 9162
rect 15324 9139 15466 9203
rect 15536 9162 15546 9203
rect 15530 9139 15546 9162
rect 15610 9139 15626 9203
rect 15690 9139 15706 9203
rect 15770 9139 15786 9203
rect 15850 9139 15866 9203
rect 15930 9139 16034 9203
rect 13544 9137 16034 9139
rect 13544 8983 13610 9137
rect 13544 8919 13545 8983
rect 13609 8919 13610 8983
rect 13544 8903 13610 8919
rect 13544 8839 13545 8903
rect 13609 8839 13610 8903
rect 13544 8823 13610 8839
rect 13544 8759 13545 8823
rect 13609 8759 13610 8823
rect 13544 8743 13610 8759
rect 13544 8679 13545 8743
rect 13609 8679 13610 8743
rect 13544 8663 13610 8679
rect 13544 8599 13545 8663
rect 13609 8599 13610 8663
rect 13544 8583 13610 8599
rect 13544 8519 13545 8583
rect 13609 8519 13610 8583
rect 13544 8503 13610 8519
rect 13544 8439 13545 8503
rect 13609 8439 13610 8503
rect 13544 8423 13610 8439
rect 13544 8359 13545 8423
rect 13609 8359 13610 8423
rect 13544 8343 13610 8359
rect 13544 8279 13545 8343
rect 13609 8279 13610 8343
rect 13544 8263 13610 8279
rect 13544 8199 13545 8263
rect 13609 8199 13610 8263
rect 13544 8109 13610 8199
rect 13670 8105 13730 9137
rect 13790 8045 13850 9075
rect 13910 8105 13970 9137
rect 14030 8045 14090 9075
rect 14150 8983 14216 9137
rect 14150 8919 14151 8983
rect 14215 8919 14216 8983
rect 14150 8903 14216 8919
rect 14150 8839 14151 8903
rect 14215 8839 14216 8903
rect 14150 8823 14216 8839
rect 14150 8759 14151 8823
rect 14215 8759 14216 8823
rect 14150 8743 14216 8759
rect 14150 8679 14151 8743
rect 14215 8679 14216 8743
rect 14150 8663 14216 8679
rect 14150 8599 14151 8663
rect 14215 8599 14216 8663
rect 14150 8583 14216 8599
rect 14150 8519 14151 8583
rect 14215 8519 14216 8583
rect 14150 8503 14216 8519
rect 14150 8439 14151 8503
rect 14215 8439 14216 8503
rect 14150 8423 14216 8439
rect 14150 8359 14151 8423
rect 14215 8359 14216 8423
rect 14150 8343 14216 8359
rect 14150 8279 14151 8343
rect 14215 8279 14216 8343
rect 14150 8263 14216 8279
rect 14150 8199 14151 8263
rect 14215 8199 14216 8263
rect 14150 8109 14216 8199
rect 14276 8045 14336 9075
rect 14396 8105 14456 9137
rect 14516 8045 14576 9075
rect 14636 8105 14696 9137
rect 14756 8983 14822 9137
rect 14756 8919 14757 8983
rect 14821 8919 14822 8983
rect 14756 8903 14822 8919
rect 14756 8839 14757 8903
rect 14821 8839 14822 8903
rect 14756 8823 14822 8839
rect 14756 8759 14757 8823
rect 14821 8759 14822 8823
rect 14756 8743 14822 8759
rect 14756 8679 14757 8743
rect 14821 8679 14822 8743
rect 14756 8663 14822 8679
rect 14756 8599 14757 8663
rect 14821 8599 14822 8663
rect 14756 8583 14822 8599
rect 14756 8519 14757 8583
rect 14821 8519 14822 8583
rect 14756 8503 14822 8519
rect 14756 8439 14757 8503
rect 14821 8439 14822 8503
rect 14756 8423 14822 8439
rect 14756 8359 14757 8423
rect 14821 8359 14822 8423
rect 14756 8343 14822 8359
rect 14756 8279 14757 8343
rect 14821 8279 14822 8343
rect 14756 8263 14822 8279
rect 14756 8199 14757 8263
rect 14821 8199 14822 8263
rect 14756 8109 14822 8199
rect 14882 8105 14942 9137
rect 15002 8045 15062 9075
rect 15122 8105 15182 9137
rect 15242 8045 15302 9075
rect 15362 8983 15428 9137
rect 15362 8919 15363 8983
rect 15427 8919 15428 8983
rect 15362 8903 15428 8919
rect 15362 8839 15363 8903
rect 15427 8839 15428 8903
rect 15362 8823 15428 8839
rect 15362 8759 15363 8823
rect 15427 8759 15428 8823
rect 15362 8743 15428 8759
rect 15362 8679 15363 8743
rect 15427 8679 15428 8743
rect 15362 8663 15428 8679
rect 15362 8599 15363 8663
rect 15427 8599 15428 8663
rect 15362 8583 15428 8599
rect 15362 8519 15363 8583
rect 15427 8519 15428 8583
rect 15362 8503 15428 8519
rect 15362 8439 15363 8503
rect 15427 8439 15428 8503
rect 15362 8423 15428 8439
rect 15362 8359 15363 8423
rect 15427 8359 15428 8423
rect 15362 8343 15428 8359
rect 15362 8279 15363 8343
rect 15427 8279 15428 8343
rect 15362 8263 15428 8279
rect 15362 8199 15363 8263
rect 15427 8199 15428 8263
rect 15362 8109 15428 8199
rect 15488 8045 15548 9075
rect 15608 8105 15668 9137
rect 15728 8045 15788 9075
rect 15848 8105 15908 9137
rect 15968 8983 16034 9137
rect 15968 8919 15969 8983
rect 16033 8919 16034 8983
rect 15968 8903 16034 8919
rect 15968 8839 15969 8903
rect 16033 8839 16034 8903
rect 15968 8823 16034 8839
rect 15968 8759 15969 8823
rect 16033 8759 16034 8823
rect 15968 8743 16034 8759
rect 15968 8679 15969 8743
rect 16033 8679 16034 8743
rect 15968 8663 16034 8679
rect 15968 8599 15969 8663
rect 16033 8599 16034 8663
rect 15968 8583 16034 8599
rect 15968 8519 15969 8583
rect 16033 8519 16034 8583
rect 15968 8503 16034 8519
rect 15968 8439 15969 8503
rect 16033 8439 16034 8503
rect 15968 8423 16034 8439
rect 15968 8359 15969 8423
rect 16033 8359 16034 8423
rect 15968 8343 16034 8359
rect 15968 8279 15969 8343
rect 16033 8279 16034 8343
rect 15968 8263 16034 8279
rect 15968 8199 15969 8263
rect 16033 8199 16034 8263
rect 15968 8109 16034 8199
rect 16094 9203 16592 9205
rect 16656 9205 16665 9226
rect 16801 9226 16883 9232
rect 16801 9205 16810 9226
rect 16656 9203 16810 9205
rect 16874 9205 16883 9226
rect 17535 9226 17617 9232
rect 17535 9205 17544 9226
rect 16874 9203 17372 9205
rect 16094 9139 16198 9203
rect 16262 9139 16278 9203
rect 16342 9139 16358 9203
rect 16422 9139 16438 9203
rect 16502 9139 16518 9203
rect 16582 9162 16592 9203
rect 16582 9139 16598 9162
rect 16662 9139 16804 9203
rect 16874 9162 16884 9203
rect 16868 9139 16884 9162
rect 16948 9139 16964 9203
rect 17028 9139 17044 9203
rect 17108 9139 17124 9203
rect 17188 9139 17204 9203
rect 17268 9139 17372 9203
rect 16094 9137 17372 9139
rect 16094 8983 16160 9137
rect 16094 8919 16095 8983
rect 16159 8919 16160 8983
rect 16094 8903 16160 8919
rect 16094 8839 16095 8903
rect 16159 8839 16160 8903
rect 16094 8823 16160 8839
rect 16094 8759 16095 8823
rect 16159 8759 16160 8823
rect 16094 8743 16160 8759
rect 16094 8679 16095 8743
rect 16159 8679 16160 8743
rect 16094 8663 16160 8679
rect 16094 8599 16095 8663
rect 16159 8599 16160 8663
rect 16094 8583 16160 8599
rect 16094 8519 16095 8583
rect 16159 8519 16160 8583
rect 16094 8503 16160 8519
rect 16094 8439 16095 8503
rect 16159 8439 16160 8503
rect 16094 8423 16160 8439
rect 16094 8359 16095 8423
rect 16159 8359 16160 8423
rect 16094 8343 16160 8359
rect 16094 8279 16095 8343
rect 16159 8279 16160 8343
rect 16094 8263 16160 8279
rect 16094 8199 16095 8263
rect 16159 8199 16160 8263
rect 16094 8109 16160 8199
rect 16220 8105 16280 9137
rect 16340 8045 16400 9075
rect 16460 8105 16520 9137
rect 16580 8045 16640 9075
rect 16700 8983 16766 9137
rect 16700 8919 16701 8983
rect 16765 8919 16766 8983
rect 16700 8903 16766 8919
rect 16700 8839 16701 8903
rect 16765 8839 16766 8903
rect 16700 8823 16766 8839
rect 16700 8759 16701 8823
rect 16765 8759 16766 8823
rect 16700 8743 16766 8759
rect 16700 8679 16701 8743
rect 16765 8679 16766 8743
rect 16700 8663 16766 8679
rect 16700 8599 16701 8663
rect 16765 8599 16766 8663
rect 16700 8583 16766 8599
rect 16700 8519 16701 8583
rect 16765 8519 16766 8583
rect 16700 8503 16766 8519
rect 16700 8439 16701 8503
rect 16765 8439 16766 8503
rect 16700 8423 16766 8439
rect 16700 8359 16701 8423
rect 16765 8359 16766 8423
rect 16700 8343 16766 8359
rect 16700 8279 16701 8343
rect 16765 8279 16766 8343
rect 16700 8263 16766 8279
rect 16700 8199 16701 8263
rect 16765 8199 16766 8263
rect 16700 8109 16766 8199
rect 16826 8045 16886 9075
rect 16946 8105 17006 9137
rect 17066 8045 17126 9075
rect 17186 8105 17246 9137
rect 17306 8983 17372 9137
rect 17306 8919 17307 8983
rect 17371 8919 17372 8983
rect 17306 8903 17372 8919
rect 17306 8839 17307 8903
rect 17371 8839 17372 8903
rect 17306 8823 17372 8839
rect 17306 8759 17307 8823
rect 17371 8759 17372 8823
rect 17306 8743 17372 8759
rect 17306 8679 17307 8743
rect 17371 8679 17372 8743
rect 17306 8663 17372 8679
rect 17306 8599 17307 8663
rect 17371 8599 17372 8663
rect 17306 8583 17372 8599
rect 17306 8519 17307 8583
rect 17371 8519 17372 8583
rect 17306 8503 17372 8519
rect 17306 8439 17307 8503
rect 17371 8439 17372 8503
rect 17306 8423 17372 8439
rect 17306 8359 17307 8423
rect 17371 8359 17372 8423
rect 17306 8343 17372 8359
rect 17306 8279 17307 8343
rect 17371 8279 17372 8343
rect 17306 8263 17372 8279
rect 17306 8199 17307 8263
rect 17371 8199 17372 8263
rect 17306 8109 17372 8199
rect 17434 9203 17544 9205
rect 17608 9205 17617 9226
rect 18257 9227 18383 9237
rect 17608 9203 18106 9205
rect 17434 9139 17538 9203
rect 17608 9162 17618 9203
rect 17602 9139 17618 9162
rect 17682 9139 17698 9203
rect 17762 9139 17778 9203
rect 17842 9139 17858 9203
rect 17922 9139 17938 9203
rect 18002 9139 18106 9203
rect 18257 9163 18288 9227
rect 18352 9163 18383 9227
rect 18257 9153 18383 9163
rect 18283 9152 18357 9153
rect 17434 9137 18106 9139
rect 17434 8983 17500 9137
rect 17434 8919 17435 8983
rect 17499 8919 17500 8983
rect 17434 8903 17500 8919
rect 17434 8839 17435 8903
rect 17499 8839 17500 8903
rect 17434 8823 17500 8839
rect 17434 8759 17435 8823
rect 17499 8759 17500 8823
rect 17434 8743 17500 8759
rect 17434 8679 17435 8743
rect 17499 8679 17500 8743
rect 17434 8663 17500 8679
rect 17434 8599 17435 8663
rect 17499 8599 17500 8663
rect 17434 8583 17500 8599
rect 17434 8519 17435 8583
rect 17499 8519 17500 8583
rect 17434 8503 17500 8519
rect 17434 8439 17435 8503
rect 17499 8439 17500 8503
rect 17434 8423 17500 8439
rect 17434 8359 17435 8423
rect 17499 8359 17500 8423
rect 17434 8343 17500 8359
rect 17434 8279 17435 8343
rect 17499 8279 17500 8343
rect 17434 8263 17500 8279
rect 17434 8199 17435 8263
rect 17499 8199 17500 8263
rect 17434 8109 17500 8199
rect 17560 8045 17620 9075
rect 17680 8105 17740 9137
rect 17800 8045 17860 9075
rect 17920 8105 17980 9137
rect 18040 8983 18106 9137
rect 18358 9057 18483 9067
rect 18358 8993 18388 9057
rect 18452 8993 18483 9057
rect 18358 8983 18483 8993
rect 18040 8919 18041 8983
rect 18105 8919 18106 8983
rect 18040 8903 18106 8919
rect 18040 8839 18041 8903
rect 18105 8839 18106 8903
rect 18167 8965 18292 8975
rect 18167 8901 18197 8965
rect 18261 8901 18292 8965
rect 18167 8891 18292 8901
rect 18040 8823 18106 8839
rect 18040 8759 18041 8823
rect 18105 8759 18106 8823
rect 18040 8743 18106 8759
rect 18040 8679 18041 8743
rect 18105 8679 18106 8743
rect 18040 8663 18106 8679
rect 18040 8599 18041 8663
rect 18105 8599 18106 8663
rect 18040 8583 18106 8599
rect 18040 8519 18041 8583
rect 18105 8519 18106 8583
rect 18040 8503 18106 8519
rect 18040 8439 18041 8503
rect 18105 8439 18106 8503
rect 18040 8423 18106 8439
rect 18040 8359 18041 8423
rect 18105 8359 18106 8423
rect 18040 8343 18106 8359
rect 18040 8279 18041 8343
rect 18105 8279 18106 8343
rect 18040 8263 18106 8279
rect 18040 8199 18041 8263
rect 18105 8199 18106 8263
rect 18040 8109 18106 8199
rect 12424 7976 12454 8040
rect 12518 7976 12549 8040
rect 12812 8043 13484 8045
rect 12812 7979 12996 8043
rect 13060 7979 13076 8043
rect 13140 7979 13156 8043
rect 13220 7979 13236 8043
rect 13300 7979 13484 8043
rect 12812 7977 13484 7979
rect 13544 8043 16034 8045
rect 13544 7979 13728 8043
rect 13792 7979 13808 8043
rect 13872 7979 13888 8043
rect 13952 7979 13968 8043
rect 14032 7979 14334 8043
rect 14398 7979 14414 8043
rect 14478 7979 14494 8043
rect 14558 7979 14574 8043
rect 14638 7979 14940 8043
rect 15004 7979 15020 8043
rect 15084 7979 15100 8043
rect 15164 7979 15180 8043
rect 15244 7979 15546 8043
rect 15610 7979 15626 8043
rect 15690 7979 15706 8043
rect 15770 7979 15786 8043
rect 15850 7979 16034 8043
rect 13544 7977 16034 7979
rect 16094 8043 17372 8045
rect 16094 7979 16278 8043
rect 16342 7979 16358 8043
rect 16422 7979 16438 8043
rect 16502 7979 16518 8043
rect 16582 7979 16884 8043
rect 16948 7979 16964 8043
rect 17028 7979 17044 8043
rect 17108 7979 17124 8043
rect 17188 7979 17372 8043
rect 16094 7977 17372 7979
rect 17434 8043 18106 8045
rect 17434 7979 17618 8043
rect 17682 7979 17698 8043
rect 17762 7979 17778 8043
rect 17842 7979 17858 8043
rect 17922 7979 18106 8043
rect 17434 7977 18106 7979
rect 12424 7966 12549 7976
rect 13478 7595 13592 7608
rect 13478 7531 13501 7595
rect 13565 7531 13592 7595
rect 13478 7521 13592 7531
rect 13652 7594 13766 7607
rect 13652 7530 13675 7594
rect 13739 7530 13766 7594
rect 13652 7520 13766 7530
rect 13877 7596 13991 7609
rect 13877 7532 13900 7596
rect 13964 7532 13991 7596
rect 13877 7522 13991 7532
rect 14078 7598 14192 7611
rect 14078 7534 14101 7598
rect 14165 7534 14192 7598
rect 14078 7524 14192 7534
rect 14301 7596 14415 7609
rect 14301 7532 14324 7596
rect 14388 7532 14415 7596
rect 14301 7522 14415 7532
rect 14510 7601 14624 7614
rect 14510 7537 14533 7601
rect 14597 7537 14624 7601
rect 14510 7527 14624 7537
rect 14738 7594 14852 7607
rect 14738 7530 14761 7594
rect 14825 7530 14852 7594
rect 14738 7520 14852 7530
rect 14928 7598 15042 7611
rect 14928 7534 14951 7598
rect 15015 7534 15042 7598
rect 14928 7524 15042 7534
rect 15133 7601 15247 7614
rect 15133 7537 15156 7601
rect 15220 7537 15247 7601
rect 15133 7527 15247 7537
rect 15332 7601 15446 7614
rect 15332 7537 15355 7601
rect 15419 7537 15446 7601
rect 15332 7527 15446 7537
rect 15548 7596 15662 7609
rect 15548 7532 15571 7596
rect 15635 7532 15662 7596
rect 15548 7522 15662 7532
rect 15936 7601 16050 7614
rect 15936 7537 15959 7601
rect 16023 7537 16050 7601
rect 15936 7527 16050 7537
rect 16171 7596 16285 7609
rect 16171 7532 16194 7596
rect 16258 7532 16285 7596
rect 16171 7522 16285 7532
rect 16413 7598 16527 7611
rect 16413 7534 16436 7598
rect 16500 7534 16527 7598
rect 16413 7524 16527 7534
rect 16645 7599 16759 7612
rect 16645 7535 16668 7599
rect 16732 7535 16759 7599
rect 16645 7525 16759 7535
rect 16874 7602 16988 7615
rect 16874 7538 16897 7602
rect 16961 7538 16988 7602
rect 16874 7528 16988 7538
rect 17123 7594 17237 7607
rect 17123 7530 17146 7594
rect 17210 7530 17237 7594
rect 17123 7520 17237 7530
rect 17341 7598 17455 7611
rect 17341 7534 17364 7598
rect 17428 7534 17455 7598
rect 17341 7524 17455 7534
rect 17570 7594 17684 7607
rect 17570 7530 17593 7594
rect 17657 7530 17684 7594
rect 17570 7520 17684 7530
rect 17791 7596 17905 7609
rect 17791 7532 17814 7596
rect 17878 7532 17905 7596
rect 17791 7522 17905 7532
rect 18007 7601 18121 7614
rect 18007 7537 18030 7601
rect 18094 7537 18121 7601
rect 18007 7527 18121 7537
rect 14836 7408 14950 7421
rect 14836 7344 14859 7408
rect 14923 7344 14950 7408
rect 17231 7407 17345 7420
rect 14836 7334 14950 7344
rect 15221 7357 15335 7370
rect 15221 7293 15244 7357
rect 15308 7293 15335 7357
rect 17231 7343 17254 7407
rect 17318 7343 17345 7407
rect 17231 7333 17345 7343
rect 17616 7358 17730 7371
rect 15221 7283 15335 7293
rect 17616 7294 17639 7358
rect 17703 7294 17730 7358
rect 17616 7284 17730 7294
rect 13480 7012 13594 7025
rect 13480 6948 13503 7012
rect 13567 6948 13594 7012
rect 13480 6938 13594 6948
rect 13655 7010 13769 7023
rect 13655 6946 13678 7010
rect 13742 6946 13769 7010
rect 13655 6936 13769 6946
rect 13852 7012 13966 7025
rect 13852 6948 13875 7012
rect 13939 6948 13966 7012
rect 13852 6938 13966 6948
rect 14071 7015 14185 7028
rect 14071 6951 14094 7015
rect 14158 6951 14185 7015
rect 14071 6941 14185 6951
rect 14303 7011 14417 7024
rect 14303 6947 14326 7011
rect 14390 6947 14417 7011
rect 14303 6937 14417 6947
rect 14527 7018 14641 7031
rect 14527 6954 14550 7018
rect 14614 6954 14641 7018
rect 14527 6944 14641 6954
rect 14739 7006 14853 7019
rect 14739 6942 14762 7006
rect 14826 6942 14853 7006
rect 14739 6932 14853 6942
rect 14961 7002 15075 7015
rect 14961 6938 14984 7002
rect 15048 6938 15075 7002
rect 14961 6928 15075 6938
rect 15184 6999 15298 7012
rect 15184 6935 15207 6999
rect 15271 6935 15298 6999
rect 15184 6925 15298 6935
rect 15394 6999 15508 7012
rect 15394 6935 15417 6999
rect 15481 6935 15508 6999
rect 15394 6925 15508 6935
rect 15607 6999 15721 7012
rect 15607 6935 15630 6999
rect 15694 6935 15721 6999
rect 15607 6925 15721 6935
rect 15924 6992 16038 7005
rect 15924 6928 15947 6992
rect 16011 6928 16038 6992
rect 15924 6918 16038 6928
rect 16126 6995 16240 7008
rect 16126 6931 16149 6995
rect 16213 6931 16240 6995
rect 16126 6921 16240 6931
rect 16327 6996 16441 7009
rect 16327 6932 16350 6996
rect 16414 6932 16441 6996
rect 16327 6922 16441 6932
rect 16506 6997 16620 7010
rect 16506 6933 16529 6997
rect 16593 6933 16620 6997
rect 16506 6923 16620 6933
rect 16698 7001 16812 7014
rect 16698 6937 16721 7001
rect 16785 6937 16812 7001
rect 16698 6927 16812 6937
rect 16883 6998 16997 7011
rect 16883 6934 16906 6998
rect 16970 6934 16997 6998
rect 16883 6924 16997 6934
rect 17115 6997 17229 7010
rect 17115 6933 17138 6997
rect 17202 6933 17229 6997
rect 17115 6923 17229 6933
rect 17320 6999 17434 7012
rect 17320 6935 17343 6999
rect 17407 6935 17434 6999
rect 17320 6925 17434 6935
rect 17526 7001 17640 7014
rect 17526 6937 17549 7001
rect 17613 6937 17640 7001
rect 17526 6927 17640 6937
rect 17734 7008 17848 7021
rect 17734 6944 17757 7008
rect 17821 6944 17848 7008
rect 17734 6934 17848 6944
rect 17956 7009 18070 7022
rect 17956 6945 17979 7009
rect 18043 6945 18070 7009
rect 17956 6935 18070 6945
rect 13507 6363 13621 6376
rect 13507 6299 13530 6363
rect 13594 6299 13621 6363
rect 13507 6289 13621 6299
rect 13723 6368 13837 6381
rect 13723 6304 13746 6368
rect 13810 6304 13837 6368
rect 13723 6294 13837 6304
rect 13929 6369 14043 6382
rect 13929 6305 13952 6369
rect 14016 6305 14043 6369
rect 13929 6295 14043 6305
rect 14131 6361 14245 6374
rect 14131 6297 14154 6361
rect 14218 6297 14245 6361
rect 14131 6287 14245 6297
rect 14327 6363 14441 6376
rect 14327 6299 14350 6363
rect 14414 6299 14441 6363
rect 14327 6289 14441 6299
rect 14552 6365 14666 6378
rect 14552 6301 14575 6365
rect 14639 6301 14666 6365
rect 14552 6291 14666 6301
rect 14767 6361 14881 6374
rect 14767 6297 14790 6361
rect 14854 6297 14881 6361
rect 14767 6287 14881 6297
rect 15002 6361 15116 6374
rect 15002 6297 15025 6361
rect 15089 6297 15116 6361
rect 15002 6287 15116 6297
rect 15210 6364 15324 6377
rect 15210 6300 15233 6364
rect 15297 6300 15324 6364
rect 15210 6290 15324 6300
rect 15452 6364 15566 6377
rect 15452 6300 15475 6364
rect 15539 6300 15566 6364
rect 15452 6290 15566 6300
rect 15650 6365 15764 6378
rect 15650 6301 15673 6365
rect 15737 6301 15764 6365
rect 15650 6291 15764 6301
rect 15957 6365 16071 6378
rect 15957 6301 15980 6365
rect 16044 6301 16071 6365
rect 15957 6291 16071 6301
rect 16182 6366 16296 6379
rect 16182 6302 16205 6366
rect 16269 6302 16296 6366
rect 16182 6292 16296 6302
rect 16411 6365 16525 6378
rect 16411 6301 16434 6365
rect 16498 6301 16525 6365
rect 16411 6291 16525 6301
rect 16627 6369 16741 6382
rect 16627 6305 16650 6369
rect 16714 6305 16741 6369
rect 16627 6295 16741 6305
rect 16850 6372 16964 6385
rect 16850 6308 16873 6372
rect 16937 6308 16964 6372
rect 16850 6298 16964 6308
rect 17074 6368 17188 6381
rect 17074 6304 17097 6368
rect 17161 6304 17188 6368
rect 17074 6294 17188 6304
rect 17301 6357 17415 6370
rect 17301 6293 17324 6357
rect 17388 6293 17415 6357
rect 17301 6283 17415 6293
rect 17514 6356 17628 6369
rect 17514 6292 17537 6356
rect 17601 6292 17628 6356
rect 17514 6282 17628 6292
rect 17725 6360 17839 6373
rect 17725 6296 17748 6360
rect 17812 6296 17839 6360
rect 17725 6286 17839 6296
rect 17952 6361 18066 6374
rect 17952 6297 17975 6361
rect 18039 6297 18066 6361
rect 17952 6287 18066 6297
rect 14841 6134 14955 6147
rect 14841 6070 14864 6134
rect 14928 6070 14955 6134
rect 17233 6136 17347 6149
rect 14841 6060 14955 6070
rect 15224 6075 15338 6088
rect 15224 6011 15247 6075
rect 15311 6011 15338 6075
rect 17233 6072 17256 6136
rect 17320 6072 17347 6136
rect 17233 6062 17347 6072
rect 17610 6082 17724 6095
rect 15224 6001 15338 6011
rect 17610 6018 17633 6082
rect 17697 6018 17724 6082
rect 17610 6008 17724 6018
rect 13533 5718 13647 5731
rect 13533 5654 13556 5718
rect 13620 5654 13647 5718
rect 13533 5644 13647 5654
rect 13758 5727 13872 5740
rect 13758 5663 13781 5727
rect 13845 5663 13872 5727
rect 13758 5653 13872 5663
rect 14035 5724 14149 5737
rect 14035 5660 14058 5724
rect 14122 5660 14149 5724
rect 14035 5650 14149 5660
rect 14256 5727 14370 5740
rect 14256 5663 14279 5727
rect 14343 5663 14370 5727
rect 14256 5653 14370 5663
rect 14501 5724 14615 5737
rect 14501 5660 14524 5724
rect 14588 5660 14615 5724
rect 14501 5650 14615 5660
rect 14727 5728 14841 5741
rect 14727 5664 14750 5728
rect 14814 5664 14841 5728
rect 14727 5654 14841 5664
rect 14939 5726 15053 5739
rect 14939 5662 14962 5726
rect 15026 5662 15053 5726
rect 14939 5652 15053 5662
rect 15159 5732 15273 5745
rect 15159 5668 15182 5732
rect 15246 5668 15273 5732
rect 15159 5658 15273 5668
rect 15397 5734 15511 5747
rect 15397 5670 15420 5734
rect 15484 5670 15511 5734
rect 15397 5660 15511 5670
rect 15610 5736 15724 5749
rect 15610 5672 15633 5736
rect 15697 5672 15724 5736
rect 15610 5662 15724 5672
rect 15997 5726 16111 5739
rect 15997 5662 16020 5726
rect 16084 5662 16111 5726
rect 15997 5652 16111 5662
rect 16344 5727 16458 5740
rect 16344 5663 16367 5727
rect 16431 5663 16458 5727
rect 16344 5653 16458 5663
rect 16580 5722 16694 5735
rect 16580 5658 16603 5722
rect 16667 5658 16694 5722
rect 16580 5648 16694 5658
rect 16764 5722 16878 5735
rect 16764 5658 16787 5722
rect 16851 5658 16878 5722
rect 16764 5648 16878 5658
rect 17003 5724 17117 5737
rect 17003 5660 17026 5724
rect 17090 5660 17117 5724
rect 17003 5650 17117 5660
rect 17206 5720 17320 5733
rect 17206 5656 17229 5720
rect 17293 5656 17320 5720
rect 17206 5646 17320 5656
rect 17391 5717 17505 5730
rect 17391 5653 17414 5717
rect 17478 5653 17505 5717
rect 17391 5643 17505 5653
rect 17582 5719 17696 5732
rect 17582 5655 17605 5719
rect 17669 5655 17696 5719
rect 17582 5645 17696 5655
rect 17773 5723 17887 5736
rect 17773 5659 17796 5723
rect 17860 5659 17887 5723
rect 17773 5649 17887 5659
rect 17959 5719 18073 5732
rect 17959 5655 17982 5719
rect 18046 5655 18073 5719
rect 17959 5645 18073 5655
rect 13406 5136 13520 5149
rect 13406 5072 13429 5136
rect 13493 5072 13520 5136
rect 13406 5062 13520 5072
rect 13611 5132 13725 5145
rect 13611 5068 13634 5132
rect 13698 5068 13725 5132
rect 13611 5058 13725 5068
rect 13797 5137 13911 5150
rect 13797 5073 13820 5137
rect 13884 5073 13911 5137
rect 13797 5063 13911 5073
rect 13991 5130 14105 5143
rect 13991 5066 14014 5130
rect 14078 5066 14105 5130
rect 13991 5056 14105 5066
rect 14210 5135 14324 5148
rect 14210 5071 14233 5135
rect 14297 5071 14324 5135
rect 14210 5061 14324 5071
rect 14420 5135 14534 5148
rect 14420 5071 14443 5135
rect 14507 5071 14534 5135
rect 14420 5061 14534 5071
rect 14649 5132 14763 5145
rect 14649 5068 14672 5132
rect 14736 5068 14763 5132
rect 14649 5058 14763 5068
rect 14895 5132 15009 5145
rect 14895 5068 14918 5132
rect 14982 5068 15009 5132
rect 14895 5058 15009 5068
rect 15169 5132 15283 5145
rect 15169 5068 15192 5132
rect 15256 5068 15283 5132
rect 15169 5058 15283 5068
rect 15444 5132 15558 5145
rect 15444 5068 15467 5132
rect 15531 5068 15558 5132
rect 15444 5058 15558 5068
rect 15680 5132 15794 5145
rect 15680 5068 15703 5132
rect 15767 5068 15794 5132
rect 15680 5058 15794 5068
rect 15903 5135 16017 5148
rect 15903 5071 15926 5135
rect 15990 5071 16017 5135
rect 15903 5061 16017 5071
rect 16121 5138 16235 5151
rect 16121 5074 16144 5138
rect 16208 5074 16235 5138
rect 16121 5064 16235 5074
rect 16299 5129 16413 5142
rect 16299 5065 16322 5129
rect 16386 5065 16413 5129
rect 16299 5055 16413 5065
rect 16538 5131 16652 5144
rect 16538 5067 16561 5131
rect 16625 5067 16652 5131
rect 16538 5057 16652 5067
rect 16735 5131 16849 5144
rect 16735 5067 16758 5131
rect 16822 5067 16849 5131
rect 16735 5057 16849 5067
rect 16933 5131 17047 5144
rect 16933 5067 16956 5131
rect 17020 5067 17047 5131
rect 16933 5057 17047 5067
rect 17146 5132 17260 5145
rect 17146 5068 17169 5132
rect 17233 5068 17260 5132
rect 17146 5058 17260 5068
rect 17369 5131 17483 5144
rect 17369 5067 17392 5131
rect 17456 5067 17483 5131
rect 17369 5057 17483 5067
rect 17566 5136 17680 5149
rect 17566 5072 17589 5136
rect 17653 5072 17680 5136
rect 17566 5062 17680 5072
rect 17782 5134 17896 5147
rect 17782 5070 17805 5134
rect 17869 5070 17896 5134
rect 17782 5060 17896 5070
rect 17991 5134 18105 5147
rect 17991 5070 18014 5134
rect 18078 5070 18105 5134
rect 17991 5060 18105 5070
<< via3 >>
rect 12468 10614 12532 10618
rect 12468 10558 12472 10614
rect 12472 10558 12528 10614
rect 12528 10558 12532 10614
rect 12468 10554 12532 10558
rect 12565 10605 12629 10608
rect 12565 10549 12568 10605
rect 12568 10549 12624 10605
rect 12624 10549 12629 10605
rect 12565 10544 12629 10549
rect 12645 10605 12709 10608
rect 12645 10549 12648 10605
rect 12648 10549 12704 10605
rect 12704 10549 12709 10605
rect 12645 10544 12709 10549
rect 12725 10605 12789 10608
rect 12725 10549 12728 10605
rect 12728 10549 12784 10605
rect 12784 10549 12789 10605
rect 12725 10544 12789 10549
rect 12805 10605 12869 10608
rect 12805 10549 12808 10605
rect 12808 10549 12864 10605
rect 12864 10549 12869 10605
rect 12805 10544 12869 10549
rect 12885 10605 12949 10608
rect 12885 10549 12888 10605
rect 12888 10549 12944 10605
rect 12944 10549 12949 10605
rect 12885 10544 12949 10549
rect 12965 10605 13029 10608
rect 12965 10549 12968 10605
rect 12968 10549 13024 10605
rect 13024 10549 13029 10605
rect 12965 10544 13029 10549
rect 13297 10608 13361 10611
rect 13297 10552 13300 10608
rect 13300 10552 13356 10608
rect 13356 10552 13361 10608
rect 13297 10547 13361 10552
rect 13377 10608 13441 10611
rect 13377 10552 13380 10608
rect 13380 10552 13436 10608
rect 13436 10552 13441 10608
rect 13377 10547 13441 10552
rect 13457 10608 13521 10611
rect 13457 10552 13460 10608
rect 13460 10552 13516 10608
rect 13516 10552 13521 10608
rect 13457 10547 13521 10552
rect 13537 10608 13601 10611
rect 13537 10552 13540 10608
rect 13540 10552 13596 10608
rect 13596 10552 13601 10608
rect 13537 10547 13601 10552
rect 13617 10608 13681 10611
rect 13617 10552 13620 10608
rect 13620 10552 13676 10608
rect 13676 10552 13681 10608
rect 13617 10547 13681 10552
rect 13697 10608 13761 10611
rect 13697 10552 13700 10608
rect 13700 10552 13756 10608
rect 13756 10552 13761 10608
rect 13697 10547 13761 10552
rect 13903 10608 13967 10611
rect 13903 10552 13908 10608
rect 13908 10552 13964 10608
rect 13964 10552 13967 10608
rect 13903 10547 13967 10552
rect 13983 10608 14047 10611
rect 13983 10552 13988 10608
rect 13988 10552 14044 10608
rect 14044 10552 14047 10608
rect 13983 10547 14047 10552
rect 14063 10608 14127 10611
rect 14063 10552 14068 10608
rect 14068 10552 14124 10608
rect 14124 10552 14127 10608
rect 14063 10547 14127 10552
rect 14143 10608 14207 10611
rect 14143 10552 14148 10608
rect 14148 10552 14204 10608
rect 14204 10552 14207 10608
rect 14143 10547 14207 10552
rect 14223 10608 14287 10611
rect 14223 10552 14228 10608
rect 14228 10552 14284 10608
rect 14284 10552 14287 10608
rect 14223 10547 14287 10552
rect 14303 10608 14367 10611
rect 14303 10552 14308 10608
rect 14308 10552 14364 10608
rect 14364 10552 14367 10608
rect 14303 10547 14367 10552
rect 14509 10608 14573 10611
rect 14509 10552 14512 10608
rect 14512 10552 14568 10608
rect 14568 10552 14573 10608
rect 14509 10547 14573 10552
rect 14589 10608 14653 10611
rect 14589 10552 14592 10608
rect 14592 10552 14648 10608
rect 14648 10552 14653 10608
rect 14589 10547 14653 10552
rect 14669 10608 14733 10611
rect 14669 10552 14672 10608
rect 14672 10552 14728 10608
rect 14728 10552 14733 10608
rect 14669 10547 14733 10552
rect 14749 10608 14813 10611
rect 14749 10552 14752 10608
rect 14752 10552 14808 10608
rect 14808 10552 14813 10608
rect 14749 10547 14813 10552
rect 14829 10608 14893 10611
rect 14829 10552 14832 10608
rect 14832 10552 14888 10608
rect 14888 10552 14893 10608
rect 14829 10547 14893 10552
rect 14909 10608 14973 10611
rect 14909 10552 14912 10608
rect 14912 10552 14968 10608
rect 14968 10552 14973 10608
rect 14909 10547 14973 10552
rect 15115 10608 15179 10611
rect 15115 10552 15120 10608
rect 15120 10552 15176 10608
rect 15176 10552 15179 10608
rect 15115 10547 15179 10552
rect 15195 10608 15259 10611
rect 15195 10552 15200 10608
rect 15200 10552 15256 10608
rect 15256 10552 15259 10608
rect 15195 10547 15259 10552
rect 15275 10608 15339 10611
rect 15275 10552 15280 10608
rect 15280 10552 15336 10608
rect 15336 10552 15339 10608
rect 15275 10547 15339 10552
rect 15355 10608 15419 10611
rect 15355 10552 15360 10608
rect 15360 10552 15416 10608
rect 15416 10552 15419 10608
rect 15355 10547 15419 10552
rect 15435 10608 15499 10611
rect 15435 10552 15440 10608
rect 15440 10552 15496 10608
rect 15496 10552 15499 10608
rect 15435 10547 15499 10552
rect 15515 10608 15579 10611
rect 15515 10552 15520 10608
rect 15520 10552 15576 10608
rect 15576 10552 15579 10608
rect 15515 10547 15579 10552
rect 15721 10608 15785 10611
rect 15721 10552 15724 10608
rect 15724 10552 15780 10608
rect 15780 10552 15785 10608
rect 15721 10547 15785 10552
rect 15801 10608 15865 10611
rect 15801 10552 15804 10608
rect 15804 10552 15860 10608
rect 15860 10552 15865 10608
rect 15801 10547 15865 10552
rect 15881 10608 15945 10611
rect 15881 10552 15884 10608
rect 15884 10552 15940 10608
rect 15940 10552 15945 10608
rect 15881 10547 15945 10552
rect 15961 10608 16025 10611
rect 15961 10552 15964 10608
rect 15964 10552 16020 10608
rect 16020 10552 16025 10608
rect 15961 10547 16025 10552
rect 16041 10608 16105 10611
rect 16041 10552 16044 10608
rect 16044 10552 16100 10608
rect 16100 10552 16105 10608
rect 16041 10547 16105 10552
rect 16121 10608 16185 10611
rect 16121 10552 16124 10608
rect 16124 10552 16180 10608
rect 16180 10552 16185 10608
rect 16121 10547 16185 10552
rect 16327 10608 16391 10611
rect 16327 10552 16332 10608
rect 16332 10552 16388 10608
rect 16388 10552 16391 10608
rect 16327 10547 16391 10552
rect 16407 10608 16471 10611
rect 16407 10552 16412 10608
rect 16412 10552 16468 10608
rect 16468 10552 16471 10608
rect 16407 10547 16471 10552
rect 16487 10608 16551 10611
rect 16487 10552 16492 10608
rect 16492 10552 16548 10608
rect 16548 10552 16551 10608
rect 16487 10547 16551 10552
rect 16567 10608 16631 10611
rect 16567 10552 16572 10608
rect 16572 10552 16628 10608
rect 16628 10552 16631 10608
rect 16567 10547 16631 10552
rect 16647 10608 16711 10611
rect 16647 10552 16652 10608
rect 16652 10552 16708 10608
rect 16708 10552 16711 10608
rect 16647 10547 16711 10552
rect 16727 10608 16791 10611
rect 16727 10552 16732 10608
rect 16732 10552 16788 10608
rect 16788 10552 16791 10608
rect 16727 10547 16791 10552
rect 16933 10608 16997 10611
rect 16933 10552 16936 10608
rect 16936 10552 16992 10608
rect 16992 10552 16997 10608
rect 16933 10547 16997 10552
rect 17013 10608 17077 10611
rect 17013 10552 17016 10608
rect 17016 10552 17072 10608
rect 17072 10552 17077 10608
rect 17013 10547 17077 10552
rect 17093 10608 17157 10611
rect 17093 10552 17096 10608
rect 17096 10552 17152 10608
rect 17152 10552 17157 10608
rect 17093 10547 17157 10552
rect 17173 10608 17237 10611
rect 17173 10552 17176 10608
rect 17176 10552 17232 10608
rect 17232 10552 17237 10608
rect 17173 10547 17237 10552
rect 17253 10608 17317 10611
rect 17253 10552 17256 10608
rect 17256 10552 17312 10608
rect 17312 10552 17317 10608
rect 17253 10547 17317 10552
rect 17333 10608 17397 10611
rect 17333 10552 17336 10608
rect 17336 10552 17392 10608
rect 17392 10552 17397 10608
rect 17333 10547 17397 10552
rect 17539 10608 17603 10611
rect 17539 10552 17544 10608
rect 17544 10552 17600 10608
rect 17600 10552 17603 10608
rect 17539 10547 17603 10552
rect 17619 10608 17683 10611
rect 17619 10552 17624 10608
rect 17624 10552 17680 10608
rect 17680 10552 17683 10608
rect 17619 10547 17683 10552
rect 17699 10608 17763 10611
rect 17699 10552 17704 10608
rect 17704 10552 17760 10608
rect 17760 10552 17763 10608
rect 17699 10547 17763 10552
rect 17779 10608 17843 10611
rect 17779 10552 17784 10608
rect 17784 10552 17840 10608
rect 17840 10552 17843 10608
rect 17779 10547 17843 10552
rect 17859 10608 17923 10611
rect 17859 10552 17864 10608
rect 17864 10552 17920 10608
rect 17920 10552 17923 10608
rect 17859 10547 17923 10552
rect 17939 10608 18003 10611
rect 17939 10552 17944 10608
rect 17944 10552 18000 10608
rect 18000 10552 18003 10608
rect 17939 10547 18003 10552
rect 12462 10324 12526 10388
rect 12462 10244 12526 10308
rect 12462 10164 12526 10228
rect 12462 10084 12526 10148
rect 11851 10009 11915 10013
rect 11851 9953 11855 10009
rect 11855 9953 11911 10009
rect 11911 9953 11915 10009
rect 11851 9949 11915 9953
rect 11982 10008 12046 10012
rect 11982 9952 11986 10008
rect 11986 9952 12042 10008
rect 12042 9952 12046 10008
rect 11982 9948 12046 9952
rect 12126 10009 12190 10013
rect 12126 9953 12130 10009
rect 12130 9953 12186 10009
rect 12186 9953 12190 10009
rect 12126 9949 12190 9953
rect 12462 10004 12526 10068
rect 12462 9924 12526 9988
rect 12462 9844 12526 9908
rect 12462 9764 12526 9828
rect 12462 9684 12526 9748
rect 12462 9604 12526 9668
rect 11869 9463 11933 9467
rect 11869 9407 11873 9463
rect 11873 9407 11929 9463
rect 11929 9407 11933 9463
rect 11869 9403 11933 9407
rect 11989 9463 12053 9467
rect 11989 9407 11993 9463
rect 11993 9407 12049 9463
rect 12049 9407 12053 9463
rect 11989 9403 12053 9407
rect 12132 9463 12196 9467
rect 12132 9407 12136 9463
rect 12136 9407 12192 9463
rect 12192 9407 12196 9463
rect 12132 9403 12196 9407
rect 13068 10324 13132 10388
rect 13068 10244 13132 10308
rect 13068 10164 13132 10228
rect 13068 10084 13132 10148
rect 13068 10004 13132 10068
rect 13068 9924 13132 9988
rect 13068 9844 13132 9908
rect 13068 9764 13132 9828
rect 13068 9684 13132 9748
rect 13068 9604 13132 9668
rect 12565 9384 12629 9448
rect 12645 9384 12709 9448
rect 12725 9384 12789 9448
rect 12805 9384 12869 9448
rect 12885 9384 12949 9448
rect 12965 9425 13029 9448
rect 12965 9384 13018 9425
rect 13018 9384 13029 9425
rect 13194 10327 13258 10391
rect 13194 10247 13258 10311
rect 13194 10167 13258 10231
rect 13194 10087 13258 10151
rect 13194 10007 13258 10071
rect 13194 9927 13258 9991
rect 13194 9847 13258 9911
rect 13194 9767 13258 9831
rect 13194 9687 13258 9751
rect 13194 9607 13258 9671
rect 13800 10327 13864 10391
rect 13800 10247 13864 10311
rect 13800 10167 13864 10231
rect 13800 10087 13864 10151
rect 13800 10007 13864 10071
rect 13800 9927 13864 9991
rect 13800 9847 13864 9911
rect 13800 9767 13864 9831
rect 13800 9687 13864 9751
rect 13800 9607 13864 9671
rect 14406 10327 14470 10391
rect 14406 10247 14470 10311
rect 14406 10167 14470 10231
rect 14406 10087 14470 10151
rect 14406 10007 14470 10071
rect 14406 9927 14470 9991
rect 14406 9847 14470 9911
rect 14406 9767 14470 9831
rect 14406 9687 14470 9751
rect 14406 9607 14470 9671
rect 15012 10327 15076 10391
rect 15012 10247 15076 10311
rect 15012 10167 15076 10231
rect 15012 10087 15076 10151
rect 15012 10007 15076 10071
rect 15012 9927 15076 9991
rect 15012 9847 15076 9911
rect 15012 9767 15076 9831
rect 15012 9687 15076 9751
rect 15012 9607 15076 9671
rect 15618 10327 15682 10391
rect 15618 10247 15682 10311
rect 15618 10167 15682 10231
rect 15618 10087 15682 10151
rect 15618 10007 15682 10071
rect 15618 9927 15682 9991
rect 15618 9847 15682 9911
rect 15618 9767 15682 9831
rect 15618 9687 15682 9751
rect 15618 9607 15682 9671
rect 16224 10327 16288 10391
rect 16224 10247 16288 10311
rect 16224 10167 16288 10231
rect 16224 10087 16288 10151
rect 16224 10007 16288 10071
rect 16224 9927 16288 9991
rect 16224 9847 16288 9911
rect 16224 9767 16288 9831
rect 16224 9687 16288 9751
rect 16224 9607 16288 9671
rect 16830 10327 16894 10391
rect 16830 10247 16894 10311
rect 16830 10167 16894 10231
rect 16830 10087 16894 10151
rect 16830 10007 16894 10071
rect 16830 9927 16894 9991
rect 16830 9847 16894 9911
rect 16830 9767 16894 9831
rect 16830 9687 16894 9751
rect 16830 9607 16894 9671
rect 17436 10327 17500 10391
rect 17436 10247 17500 10311
rect 17436 10167 17500 10231
rect 17436 10087 17500 10151
rect 17436 10007 17500 10071
rect 17436 9927 17500 9991
rect 17436 9847 17500 9911
rect 17436 9767 17500 9831
rect 17436 9687 17500 9751
rect 17436 9607 17500 9671
rect 18277 10552 18341 10556
rect 18277 10496 18281 10552
rect 18281 10496 18337 10552
rect 18337 10496 18341 10552
rect 18277 10492 18341 10496
rect 18042 10327 18106 10391
rect 18282 10408 18346 10412
rect 18282 10352 18286 10408
rect 18286 10352 18342 10408
rect 18342 10352 18346 10408
rect 18282 10348 18346 10352
rect 18042 10247 18106 10311
rect 18042 10167 18106 10231
rect 18283 10256 18347 10260
rect 18283 10200 18287 10256
rect 18287 10200 18343 10256
rect 18343 10200 18347 10256
rect 18283 10196 18347 10200
rect 18042 10087 18106 10151
rect 18042 10007 18106 10071
rect 18283 10086 18347 10090
rect 18283 10030 18287 10086
rect 18287 10030 18343 10086
rect 18343 10030 18347 10086
rect 18283 10026 18347 10030
rect 18042 9927 18106 9991
rect 18042 9847 18106 9911
rect 18282 9929 18346 9933
rect 18282 9873 18286 9929
rect 18286 9873 18342 9929
rect 18342 9873 18346 9929
rect 18282 9869 18346 9873
rect 18042 9767 18106 9831
rect 18042 9687 18106 9751
rect 18042 9607 18106 9671
rect 18200 9687 18264 9691
rect 18200 9631 18204 9687
rect 18204 9631 18260 9687
rect 18260 9631 18264 9687
rect 18200 9627 18264 9631
rect 18577 9695 18641 9699
rect 18577 9639 18581 9695
rect 18581 9639 18637 9695
rect 18637 9639 18641 9695
rect 18577 9635 18641 9639
rect 18777 9695 18841 9699
rect 18777 9639 18781 9695
rect 18781 9639 18837 9695
rect 18837 9639 18841 9695
rect 18777 9635 18841 9639
rect 13297 9387 13361 9451
rect 13377 9387 13441 9451
rect 13457 9387 13521 9451
rect 13537 9387 13601 9451
rect 13617 9387 13681 9451
rect 13697 9428 13761 9451
rect 13697 9387 13750 9428
rect 13750 9387 13761 9428
rect 13903 9428 13967 9451
rect 13903 9387 13914 9428
rect 13914 9387 13967 9428
rect 13983 9387 14047 9451
rect 14063 9387 14127 9451
rect 14143 9387 14207 9451
rect 14223 9387 14287 9451
rect 14303 9387 14367 9451
rect 14509 9387 14573 9451
rect 14589 9387 14653 9451
rect 14669 9387 14733 9451
rect 14749 9387 14813 9451
rect 14829 9387 14893 9451
rect 14909 9428 14973 9451
rect 14909 9387 14962 9428
rect 14962 9387 14973 9428
rect 15115 9428 15179 9451
rect 15115 9387 15126 9428
rect 15126 9387 15179 9428
rect 15195 9387 15259 9451
rect 15275 9387 15339 9451
rect 15355 9387 15419 9451
rect 15435 9387 15499 9451
rect 15515 9387 15579 9451
rect 15721 9387 15785 9451
rect 15801 9387 15865 9451
rect 15881 9387 15945 9451
rect 15961 9387 16025 9451
rect 16041 9387 16105 9451
rect 16121 9428 16185 9451
rect 16121 9387 16174 9428
rect 16174 9387 16185 9428
rect 16327 9428 16391 9451
rect 16327 9387 16338 9428
rect 16338 9387 16391 9428
rect 16407 9387 16471 9451
rect 16487 9387 16551 9451
rect 16567 9387 16631 9451
rect 16647 9387 16711 9451
rect 16727 9387 16791 9451
rect 16933 9387 16997 9451
rect 17013 9387 17077 9451
rect 17093 9387 17157 9451
rect 17173 9387 17237 9451
rect 17253 9387 17317 9451
rect 17333 9428 17397 9451
rect 17333 9387 17386 9428
rect 17386 9387 17397 9428
rect 17539 9428 17603 9451
rect 17539 9387 17550 9428
rect 17550 9387 17603 9428
rect 17619 9387 17683 9451
rect 17699 9387 17763 9451
rect 17779 9387 17843 9451
rect 17859 9387 17923 9451
rect 17939 9387 18003 9451
rect 18288 9426 18352 9430
rect 18288 9370 18292 9426
rect 18292 9370 18348 9426
rect 18348 9370 18352 9426
rect 18288 9366 18352 9370
rect 12916 9139 12980 9203
rect 12996 9139 13060 9203
rect 13076 9139 13140 9203
rect 13156 9139 13220 9203
rect 13236 9139 13300 9203
rect 13316 9162 13374 9203
rect 13374 9162 13380 9203
rect 13316 9139 13380 9162
rect 12813 8919 12877 8983
rect 12813 8839 12877 8903
rect 12813 8759 12877 8823
rect 12813 8679 12877 8743
rect 12813 8599 12877 8663
rect 12813 8519 12877 8583
rect 12813 8439 12877 8503
rect 12813 8359 12877 8423
rect 12813 8279 12877 8343
rect 12813 8199 12877 8263
rect 13419 8919 13483 8983
rect 13419 8839 13483 8903
rect 13419 8759 13483 8823
rect 13419 8679 13483 8743
rect 13419 8599 13483 8663
rect 13419 8519 13483 8583
rect 13419 8439 13483 8503
rect 13419 8359 13483 8423
rect 13419 8279 13483 8343
rect 13419 8199 13483 8263
rect 13648 9139 13712 9203
rect 13728 9139 13792 9203
rect 13808 9139 13872 9203
rect 13888 9139 13952 9203
rect 13968 9139 14032 9203
rect 14048 9162 14106 9203
rect 14106 9162 14112 9203
rect 14048 9139 14112 9162
rect 14254 9162 14260 9203
rect 14260 9162 14318 9203
rect 14254 9139 14318 9162
rect 14334 9139 14398 9203
rect 14414 9139 14478 9203
rect 14494 9139 14558 9203
rect 14574 9139 14638 9203
rect 14654 9139 14718 9203
rect 14860 9139 14924 9203
rect 14940 9139 15004 9203
rect 15020 9139 15084 9203
rect 15100 9139 15164 9203
rect 15180 9139 15244 9203
rect 15260 9162 15318 9203
rect 15318 9162 15324 9203
rect 15260 9139 15324 9162
rect 15466 9162 15472 9203
rect 15472 9162 15530 9203
rect 15466 9139 15530 9162
rect 15546 9139 15610 9203
rect 15626 9139 15690 9203
rect 15706 9139 15770 9203
rect 15786 9139 15850 9203
rect 15866 9139 15930 9203
rect 13545 8919 13609 8983
rect 13545 8839 13609 8903
rect 13545 8759 13609 8823
rect 13545 8679 13609 8743
rect 13545 8599 13609 8663
rect 13545 8519 13609 8583
rect 13545 8439 13609 8503
rect 13545 8359 13609 8423
rect 13545 8279 13609 8343
rect 13545 8199 13609 8263
rect 14151 8919 14215 8983
rect 14151 8839 14215 8903
rect 14151 8759 14215 8823
rect 14151 8679 14215 8743
rect 14151 8599 14215 8663
rect 14151 8519 14215 8583
rect 14151 8439 14215 8503
rect 14151 8359 14215 8423
rect 14151 8279 14215 8343
rect 14151 8199 14215 8263
rect 14757 8919 14821 8983
rect 14757 8839 14821 8903
rect 14757 8759 14821 8823
rect 14757 8679 14821 8743
rect 14757 8599 14821 8663
rect 14757 8519 14821 8583
rect 14757 8439 14821 8503
rect 14757 8359 14821 8423
rect 14757 8279 14821 8343
rect 14757 8199 14821 8263
rect 15363 8919 15427 8983
rect 15363 8839 15427 8903
rect 15363 8759 15427 8823
rect 15363 8679 15427 8743
rect 15363 8599 15427 8663
rect 15363 8519 15427 8583
rect 15363 8439 15427 8503
rect 15363 8359 15427 8423
rect 15363 8279 15427 8343
rect 15363 8199 15427 8263
rect 15969 8919 16033 8983
rect 15969 8839 16033 8903
rect 15969 8759 16033 8823
rect 15969 8679 16033 8743
rect 15969 8599 16033 8663
rect 15969 8519 16033 8583
rect 15969 8439 16033 8503
rect 15969 8359 16033 8423
rect 15969 8279 16033 8343
rect 15969 8199 16033 8263
rect 16198 9139 16262 9203
rect 16278 9139 16342 9203
rect 16358 9139 16422 9203
rect 16438 9139 16502 9203
rect 16518 9139 16582 9203
rect 16598 9162 16656 9203
rect 16656 9162 16662 9203
rect 16598 9139 16662 9162
rect 16804 9162 16810 9203
rect 16810 9162 16868 9203
rect 16804 9139 16868 9162
rect 16884 9139 16948 9203
rect 16964 9139 17028 9203
rect 17044 9139 17108 9203
rect 17124 9139 17188 9203
rect 17204 9139 17268 9203
rect 16095 8919 16159 8983
rect 16095 8839 16159 8903
rect 16095 8759 16159 8823
rect 16095 8679 16159 8743
rect 16095 8599 16159 8663
rect 16095 8519 16159 8583
rect 16095 8439 16159 8503
rect 16095 8359 16159 8423
rect 16095 8279 16159 8343
rect 16095 8199 16159 8263
rect 16701 8919 16765 8983
rect 16701 8839 16765 8903
rect 16701 8759 16765 8823
rect 16701 8679 16765 8743
rect 16701 8599 16765 8663
rect 16701 8519 16765 8583
rect 16701 8439 16765 8503
rect 16701 8359 16765 8423
rect 16701 8279 16765 8343
rect 16701 8199 16765 8263
rect 17307 8919 17371 8983
rect 17307 8839 17371 8903
rect 17307 8759 17371 8823
rect 17307 8679 17371 8743
rect 17307 8599 17371 8663
rect 17307 8519 17371 8583
rect 17307 8439 17371 8503
rect 17307 8359 17371 8423
rect 17307 8279 17371 8343
rect 17307 8199 17371 8263
rect 17538 9162 17544 9203
rect 17544 9162 17602 9203
rect 17538 9139 17602 9162
rect 17618 9139 17682 9203
rect 17698 9139 17762 9203
rect 17778 9139 17842 9203
rect 17858 9139 17922 9203
rect 17938 9139 18002 9203
rect 18288 9223 18352 9227
rect 18288 9167 18292 9223
rect 18292 9167 18348 9223
rect 18348 9167 18352 9223
rect 18288 9163 18352 9167
rect 17435 8919 17499 8983
rect 17435 8839 17499 8903
rect 17435 8759 17499 8823
rect 17435 8679 17499 8743
rect 17435 8599 17499 8663
rect 17435 8519 17499 8583
rect 17435 8439 17499 8503
rect 17435 8359 17499 8423
rect 17435 8279 17499 8343
rect 17435 8199 17499 8263
rect 18388 9053 18452 9057
rect 18388 8997 18392 9053
rect 18392 8997 18448 9053
rect 18448 8997 18452 9053
rect 18388 8993 18452 8997
rect 18041 8919 18105 8983
rect 18041 8839 18105 8903
rect 18197 8961 18261 8965
rect 18197 8905 18201 8961
rect 18201 8905 18257 8961
rect 18257 8905 18261 8961
rect 18197 8901 18261 8905
rect 18041 8759 18105 8823
rect 18041 8679 18105 8743
rect 18041 8599 18105 8663
rect 18041 8519 18105 8583
rect 18041 8439 18105 8503
rect 18041 8359 18105 8423
rect 18041 8279 18105 8343
rect 18041 8199 18105 8263
rect 12454 8036 12518 8040
rect 12454 7980 12458 8036
rect 12458 7980 12514 8036
rect 12514 7980 12518 8036
rect 12454 7976 12518 7980
rect 12996 8039 13060 8043
rect 12996 7983 13000 8039
rect 13000 7983 13056 8039
rect 13056 7983 13060 8039
rect 12996 7979 13060 7983
rect 13076 8039 13140 8043
rect 13076 7983 13080 8039
rect 13080 7983 13136 8039
rect 13136 7983 13140 8039
rect 13076 7979 13140 7983
rect 13156 8039 13220 8043
rect 13156 7983 13160 8039
rect 13160 7983 13216 8039
rect 13216 7983 13220 8039
rect 13156 7979 13220 7983
rect 13236 8039 13300 8043
rect 13236 7983 13240 8039
rect 13240 7983 13296 8039
rect 13296 7983 13300 8039
rect 13236 7979 13300 7983
rect 13728 8039 13792 8043
rect 13728 7983 13732 8039
rect 13732 7983 13788 8039
rect 13788 7983 13792 8039
rect 13728 7979 13792 7983
rect 13808 8039 13872 8043
rect 13808 7983 13812 8039
rect 13812 7983 13868 8039
rect 13868 7983 13872 8039
rect 13808 7979 13872 7983
rect 13888 8039 13952 8043
rect 13888 7983 13892 8039
rect 13892 7983 13948 8039
rect 13948 7983 13952 8039
rect 13888 7979 13952 7983
rect 13968 8039 14032 8043
rect 13968 7983 13972 8039
rect 13972 7983 14028 8039
rect 14028 7983 14032 8039
rect 13968 7979 14032 7983
rect 14334 8039 14398 8043
rect 14334 7983 14338 8039
rect 14338 7983 14394 8039
rect 14394 7983 14398 8039
rect 14334 7979 14398 7983
rect 14414 8039 14478 8043
rect 14414 7983 14418 8039
rect 14418 7983 14474 8039
rect 14474 7983 14478 8039
rect 14414 7979 14478 7983
rect 14494 8039 14558 8043
rect 14494 7983 14498 8039
rect 14498 7983 14554 8039
rect 14554 7983 14558 8039
rect 14494 7979 14558 7983
rect 14574 8039 14638 8043
rect 14574 7983 14578 8039
rect 14578 7983 14634 8039
rect 14634 7983 14638 8039
rect 14574 7979 14638 7983
rect 14940 8039 15004 8043
rect 14940 7983 14944 8039
rect 14944 7983 15000 8039
rect 15000 7983 15004 8039
rect 14940 7979 15004 7983
rect 15020 8039 15084 8043
rect 15020 7983 15024 8039
rect 15024 7983 15080 8039
rect 15080 7983 15084 8039
rect 15020 7979 15084 7983
rect 15100 8039 15164 8043
rect 15100 7983 15104 8039
rect 15104 7983 15160 8039
rect 15160 7983 15164 8039
rect 15100 7979 15164 7983
rect 15180 8039 15244 8043
rect 15180 7983 15184 8039
rect 15184 7983 15240 8039
rect 15240 7983 15244 8039
rect 15180 7979 15244 7983
rect 15546 8039 15610 8043
rect 15546 7983 15550 8039
rect 15550 7983 15606 8039
rect 15606 7983 15610 8039
rect 15546 7979 15610 7983
rect 15626 8039 15690 8043
rect 15626 7983 15630 8039
rect 15630 7983 15686 8039
rect 15686 7983 15690 8039
rect 15626 7979 15690 7983
rect 15706 8039 15770 8043
rect 15706 7983 15710 8039
rect 15710 7983 15766 8039
rect 15766 7983 15770 8039
rect 15706 7979 15770 7983
rect 15786 8039 15850 8043
rect 15786 7983 15790 8039
rect 15790 7983 15846 8039
rect 15846 7983 15850 8039
rect 15786 7979 15850 7983
rect 16278 8039 16342 8043
rect 16278 7983 16282 8039
rect 16282 7983 16338 8039
rect 16338 7983 16342 8039
rect 16278 7979 16342 7983
rect 16358 8039 16422 8043
rect 16358 7983 16362 8039
rect 16362 7983 16418 8039
rect 16418 7983 16422 8039
rect 16358 7979 16422 7983
rect 16438 8039 16502 8043
rect 16438 7983 16442 8039
rect 16442 7983 16498 8039
rect 16498 7983 16502 8039
rect 16438 7979 16502 7983
rect 16518 8039 16582 8043
rect 16518 7983 16522 8039
rect 16522 7983 16578 8039
rect 16578 7983 16582 8039
rect 16518 7979 16582 7983
rect 16884 8039 16948 8043
rect 16884 7983 16888 8039
rect 16888 7983 16944 8039
rect 16944 7983 16948 8039
rect 16884 7979 16948 7983
rect 16964 8039 17028 8043
rect 16964 7983 16968 8039
rect 16968 7983 17024 8039
rect 17024 7983 17028 8039
rect 16964 7979 17028 7983
rect 17044 8039 17108 8043
rect 17044 7983 17048 8039
rect 17048 7983 17104 8039
rect 17104 7983 17108 8039
rect 17044 7979 17108 7983
rect 17124 8039 17188 8043
rect 17124 7983 17128 8039
rect 17128 7983 17184 8039
rect 17184 7983 17188 8039
rect 17124 7979 17188 7983
rect 17618 8039 17682 8043
rect 17618 7983 17622 8039
rect 17622 7983 17678 8039
rect 17678 7983 17682 8039
rect 17618 7979 17682 7983
rect 17698 8039 17762 8043
rect 17698 7983 17702 8039
rect 17702 7983 17758 8039
rect 17758 7983 17762 8039
rect 17698 7979 17762 7983
rect 17778 8039 17842 8043
rect 17778 7983 17782 8039
rect 17782 7983 17838 8039
rect 17838 7983 17842 8039
rect 17778 7979 17842 7983
rect 17858 8039 17922 8043
rect 17858 7983 17862 8039
rect 17862 7983 17918 8039
rect 17918 7983 17922 8039
rect 17858 7979 17922 7983
rect 13501 7591 13565 7595
rect 13501 7535 13505 7591
rect 13505 7535 13561 7591
rect 13561 7535 13565 7591
rect 13501 7531 13565 7535
rect 13675 7590 13739 7594
rect 13675 7534 13679 7590
rect 13679 7534 13735 7590
rect 13735 7534 13739 7590
rect 13675 7530 13739 7534
rect 13900 7592 13964 7596
rect 13900 7536 13904 7592
rect 13904 7536 13960 7592
rect 13960 7536 13964 7592
rect 13900 7532 13964 7536
rect 14101 7594 14165 7598
rect 14101 7538 14105 7594
rect 14105 7538 14161 7594
rect 14161 7538 14165 7594
rect 14101 7534 14165 7538
rect 14324 7592 14388 7596
rect 14324 7536 14328 7592
rect 14328 7536 14384 7592
rect 14384 7536 14388 7592
rect 14324 7532 14388 7536
rect 14533 7597 14597 7601
rect 14533 7541 14537 7597
rect 14537 7541 14593 7597
rect 14593 7541 14597 7597
rect 14533 7537 14597 7541
rect 14761 7590 14825 7594
rect 14761 7534 14765 7590
rect 14765 7534 14821 7590
rect 14821 7534 14825 7590
rect 14761 7530 14825 7534
rect 14951 7594 15015 7598
rect 14951 7538 14955 7594
rect 14955 7538 15011 7594
rect 15011 7538 15015 7594
rect 14951 7534 15015 7538
rect 15156 7597 15220 7601
rect 15156 7541 15160 7597
rect 15160 7541 15216 7597
rect 15216 7541 15220 7597
rect 15156 7537 15220 7541
rect 15355 7597 15419 7601
rect 15355 7541 15359 7597
rect 15359 7541 15415 7597
rect 15415 7541 15419 7597
rect 15355 7537 15419 7541
rect 15571 7592 15635 7596
rect 15571 7536 15575 7592
rect 15575 7536 15631 7592
rect 15631 7536 15635 7592
rect 15571 7532 15635 7536
rect 15959 7597 16023 7601
rect 15959 7541 15963 7597
rect 15963 7541 16019 7597
rect 16019 7541 16023 7597
rect 15959 7537 16023 7541
rect 16194 7592 16258 7596
rect 16194 7536 16198 7592
rect 16198 7536 16254 7592
rect 16254 7536 16258 7592
rect 16194 7532 16258 7536
rect 16436 7594 16500 7598
rect 16436 7538 16440 7594
rect 16440 7538 16496 7594
rect 16496 7538 16500 7594
rect 16436 7534 16500 7538
rect 16668 7595 16732 7599
rect 16668 7539 16672 7595
rect 16672 7539 16728 7595
rect 16728 7539 16732 7595
rect 16668 7535 16732 7539
rect 16897 7598 16961 7602
rect 16897 7542 16901 7598
rect 16901 7542 16957 7598
rect 16957 7542 16961 7598
rect 16897 7538 16961 7542
rect 17146 7590 17210 7594
rect 17146 7534 17150 7590
rect 17150 7534 17206 7590
rect 17206 7534 17210 7590
rect 17146 7530 17210 7534
rect 17364 7594 17428 7598
rect 17364 7538 17368 7594
rect 17368 7538 17424 7594
rect 17424 7538 17428 7594
rect 17364 7534 17428 7538
rect 17593 7590 17657 7594
rect 17593 7534 17597 7590
rect 17597 7534 17653 7590
rect 17653 7534 17657 7590
rect 17593 7530 17657 7534
rect 17814 7592 17878 7596
rect 17814 7536 17818 7592
rect 17818 7536 17874 7592
rect 17874 7536 17878 7592
rect 17814 7532 17878 7536
rect 18030 7597 18094 7601
rect 18030 7541 18034 7597
rect 18034 7541 18090 7597
rect 18090 7541 18094 7597
rect 18030 7537 18094 7541
rect 14859 7404 14923 7408
rect 14859 7348 14863 7404
rect 14863 7348 14919 7404
rect 14919 7348 14923 7404
rect 14859 7344 14923 7348
rect 15244 7353 15308 7357
rect 15244 7297 15248 7353
rect 15248 7297 15304 7353
rect 15304 7297 15308 7353
rect 15244 7293 15308 7297
rect 17254 7403 17318 7407
rect 17254 7347 17258 7403
rect 17258 7347 17314 7403
rect 17314 7347 17318 7403
rect 17254 7343 17318 7347
rect 17639 7354 17703 7358
rect 17639 7298 17643 7354
rect 17643 7298 17699 7354
rect 17699 7298 17703 7354
rect 17639 7294 17703 7298
rect 13503 7008 13567 7012
rect 13503 6952 13507 7008
rect 13507 6952 13563 7008
rect 13563 6952 13567 7008
rect 13503 6948 13567 6952
rect 13678 7006 13742 7010
rect 13678 6950 13682 7006
rect 13682 6950 13738 7006
rect 13738 6950 13742 7006
rect 13678 6946 13742 6950
rect 13875 7008 13939 7012
rect 13875 6952 13879 7008
rect 13879 6952 13935 7008
rect 13935 6952 13939 7008
rect 13875 6948 13939 6952
rect 14094 7011 14158 7015
rect 14094 6955 14098 7011
rect 14098 6955 14154 7011
rect 14154 6955 14158 7011
rect 14094 6951 14158 6955
rect 14326 7007 14390 7011
rect 14326 6951 14330 7007
rect 14330 6951 14386 7007
rect 14386 6951 14390 7007
rect 14326 6947 14390 6951
rect 14550 7014 14614 7018
rect 14550 6958 14554 7014
rect 14554 6958 14610 7014
rect 14610 6958 14614 7014
rect 14550 6954 14614 6958
rect 14762 7002 14826 7006
rect 14762 6946 14766 7002
rect 14766 6946 14822 7002
rect 14822 6946 14826 7002
rect 14762 6942 14826 6946
rect 14984 6998 15048 7002
rect 14984 6942 14988 6998
rect 14988 6942 15044 6998
rect 15044 6942 15048 6998
rect 14984 6938 15048 6942
rect 15207 6995 15271 6999
rect 15207 6939 15211 6995
rect 15211 6939 15267 6995
rect 15267 6939 15271 6995
rect 15207 6935 15271 6939
rect 15417 6995 15481 6999
rect 15417 6939 15421 6995
rect 15421 6939 15477 6995
rect 15477 6939 15481 6995
rect 15417 6935 15481 6939
rect 15630 6995 15694 6999
rect 15630 6939 15634 6995
rect 15634 6939 15690 6995
rect 15690 6939 15694 6995
rect 15630 6935 15694 6939
rect 15947 6988 16011 6992
rect 15947 6932 15951 6988
rect 15951 6932 16007 6988
rect 16007 6932 16011 6988
rect 15947 6928 16011 6932
rect 16149 6991 16213 6995
rect 16149 6935 16153 6991
rect 16153 6935 16209 6991
rect 16209 6935 16213 6991
rect 16149 6931 16213 6935
rect 16350 6992 16414 6996
rect 16350 6936 16354 6992
rect 16354 6936 16410 6992
rect 16410 6936 16414 6992
rect 16350 6932 16414 6936
rect 16529 6993 16593 6997
rect 16529 6937 16533 6993
rect 16533 6937 16589 6993
rect 16589 6937 16593 6993
rect 16529 6933 16593 6937
rect 16721 6997 16785 7001
rect 16721 6941 16725 6997
rect 16725 6941 16781 6997
rect 16781 6941 16785 6997
rect 16721 6937 16785 6941
rect 16906 6994 16970 6998
rect 16906 6938 16910 6994
rect 16910 6938 16966 6994
rect 16966 6938 16970 6994
rect 16906 6934 16970 6938
rect 17138 6993 17202 6997
rect 17138 6937 17142 6993
rect 17142 6937 17198 6993
rect 17198 6937 17202 6993
rect 17138 6933 17202 6937
rect 17343 6995 17407 6999
rect 17343 6939 17347 6995
rect 17347 6939 17403 6995
rect 17403 6939 17407 6995
rect 17343 6935 17407 6939
rect 17549 6997 17613 7001
rect 17549 6941 17553 6997
rect 17553 6941 17609 6997
rect 17609 6941 17613 6997
rect 17549 6937 17613 6941
rect 17757 7004 17821 7008
rect 17757 6948 17761 7004
rect 17761 6948 17817 7004
rect 17817 6948 17821 7004
rect 17757 6944 17821 6948
rect 17979 7005 18043 7009
rect 17979 6949 17983 7005
rect 17983 6949 18039 7005
rect 18039 6949 18043 7005
rect 17979 6945 18043 6949
rect 13530 6359 13594 6363
rect 13530 6303 13534 6359
rect 13534 6303 13590 6359
rect 13590 6303 13594 6359
rect 13530 6299 13594 6303
rect 13746 6364 13810 6368
rect 13746 6308 13750 6364
rect 13750 6308 13806 6364
rect 13806 6308 13810 6364
rect 13746 6304 13810 6308
rect 13952 6365 14016 6369
rect 13952 6309 13956 6365
rect 13956 6309 14012 6365
rect 14012 6309 14016 6365
rect 13952 6305 14016 6309
rect 14154 6357 14218 6361
rect 14154 6301 14158 6357
rect 14158 6301 14214 6357
rect 14214 6301 14218 6357
rect 14154 6297 14218 6301
rect 14350 6359 14414 6363
rect 14350 6303 14354 6359
rect 14354 6303 14410 6359
rect 14410 6303 14414 6359
rect 14350 6299 14414 6303
rect 14575 6361 14639 6365
rect 14575 6305 14579 6361
rect 14579 6305 14635 6361
rect 14635 6305 14639 6361
rect 14575 6301 14639 6305
rect 14790 6357 14854 6361
rect 14790 6301 14794 6357
rect 14794 6301 14850 6357
rect 14850 6301 14854 6357
rect 14790 6297 14854 6301
rect 15025 6357 15089 6361
rect 15025 6301 15029 6357
rect 15029 6301 15085 6357
rect 15085 6301 15089 6357
rect 15025 6297 15089 6301
rect 15233 6360 15297 6364
rect 15233 6304 15237 6360
rect 15237 6304 15293 6360
rect 15293 6304 15297 6360
rect 15233 6300 15297 6304
rect 15475 6360 15539 6364
rect 15475 6304 15479 6360
rect 15479 6304 15535 6360
rect 15535 6304 15539 6360
rect 15475 6300 15539 6304
rect 15673 6361 15737 6365
rect 15673 6305 15677 6361
rect 15677 6305 15733 6361
rect 15733 6305 15737 6361
rect 15673 6301 15737 6305
rect 15980 6361 16044 6365
rect 15980 6305 15984 6361
rect 15984 6305 16040 6361
rect 16040 6305 16044 6361
rect 15980 6301 16044 6305
rect 16205 6362 16269 6366
rect 16205 6306 16209 6362
rect 16209 6306 16265 6362
rect 16265 6306 16269 6362
rect 16205 6302 16269 6306
rect 16434 6361 16498 6365
rect 16434 6305 16438 6361
rect 16438 6305 16494 6361
rect 16494 6305 16498 6361
rect 16434 6301 16498 6305
rect 16650 6365 16714 6369
rect 16650 6309 16654 6365
rect 16654 6309 16710 6365
rect 16710 6309 16714 6365
rect 16650 6305 16714 6309
rect 16873 6368 16937 6372
rect 16873 6312 16877 6368
rect 16877 6312 16933 6368
rect 16933 6312 16937 6368
rect 16873 6308 16937 6312
rect 17097 6364 17161 6368
rect 17097 6308 17101 6364
rect 17101 6308 17157 6364
rect 17157 6308 17161 6364
rect 17097 6304 17161 6308
rect 17324 6353 17388 6357
rect 17324 6297 17328 6353
rect 17328 6297 17384 6353
rect 17384 6297 17388 6353
rect 17324 6293 17388 6297
rect 17537 6352 17601 6356
rect 17537 6296 17541 6352
rect 17541 6296 17597 6352
rect 17597 6296 17601 6352
rect 17537 6292 17601 6296
rect 17748 6356 17812 6360
rect 17748 6300 17752 6356
rect 17752 6300 17808 6356
rect 17808 6300 17812 6356
rect 17748 6296 17812 6300
rect 17975 6357 18039 6361
rect 17975 6301 17979 6357
rect 17979 6301 18035 6357
rect 18035 6301 18039 6357
rect 17975 6297 18039 6301
rect 14864 6130 14928 6134
rect 14864 6074 14868 6130
rect 14868 6074 14924 6130
rect 14924 6074 14928 6130
rect 14864 6070 14928 6074
rect 15247 6071 15311 6075
rect 15247 6015 15251 6071
rect 15251 6015 15307 6071
rect 15307 6015 15311 6071
rect 15247 6011 15311 6015
rect 17256 6132 17320 6136
rect 17256 6076 17260 6132
rect 17260 6076 17316 6132
rect 17316 6076 17320 6132
rect 17256 6072 17320 6076
rect 17633 6078 17697 6082
rect 17633 6022 17637 6078
rect 17637 6022 17693 6078
rect 17693 6022 17697 6078
rect 17633 6018 17697 6022
rect 13556 5714 13620 5718
rect 13556 5658 13560 5714
rect 13560 5658 13616 5714
rect 13616 5658 13620 5714
rect 13556 5654 13620 5658
rect 13781 5723 13845 5727
rect 13781 5667 13785 5723
rect 13785 5667 13841 5723
rect 13841 5667 13845 5723
rect 13781 5663 13845 5667
rect 14058 5720 14122 5724
rect 14058 5664 14062 5720
rect 14062 5664 14118 5720
rect 14118 5664 14122 5720
rect 14058 5660 14122 5664
rect 14279 5723 14343 5727
rect 14279 5667 14283 5723
rect 14283 5667 14339 5723
rect 14339 5667 14343 5723
rect 14279 5663 14343 5667
rect 14524 5720 14588 5724
rect 14524 5664 14528 5720
rect 14528 5664 14584 5720
rect 14584 5664 14588 5720
rect 14524 5660 14588 5664
rect 14750 5724 14814 5728
rect 14750 5668 14754 5724
rect 14754 5668 14810 5724
rect 14810 5668 14814 5724
rect 14750 5664 14814 5668
rect 14962 5722 15026 5726
rect 14962 5666 14966 5722
rect 14966 5666 15022 5722
rect 15022 5666 15026 5722
rect 14962 5662 15026 5666
rect 15182 5728 15246 5732
rect 15182 5672 15186 5728
rect 15186 5672 15242 5728
rect 15242 5672 15246 5728
rect 15182 5668 15246 5672
rect 15420 5730 15484 5734
rect 15420 5674 15424 5730
rect 15424 5674 15480 5730
rect 15480 5674 15484 5730
rect 15420 5670 15484 5674
rect 15633 5732 15697 5736
rect 15633 5676 15637 5732
rect 15637 5676 15693 5732
rect 15693 5676 15697 5732
rect 15633 5672 15697 5676
rect 16020 5722 16084 5726
rect 16020 5666 16024 5722
rect 16024 5666 16080 5722
rect 16080 5666 16084 5722
rect 16020 5662 16084 5666
rect 16367 5723 16431 5727
rect 16367 5667 16371 5723
rect 16371 5667 16427 5723
rect 16427 5667 16431 5723
rect 16367 5663 16431 5667
rect 16603 5718 16667 5722
rect 16603 5662 16607 5718
rect 16607 5662 16663 5718
rect 16663 5662 16667 5718
rect 16603 5658 16667 5662
rect 16787 5718 16851 5722
rect 16787 5662 16791 5718
rect 16791 5662 16847 5718
rect 16847 5662 16851 5718
rect 16787 5658 16851 5662
rect 17026 5720 17090 5724
rect 17026 5664 17030 5720
rect 17030 5664 17086 5720
rect 17086 5664 17090 5720
rect 17026 5660 17090 5664
rect 17229 5716 17293 5720
rect 17229 5660 17233 5716
rect 17233 5660 17289 5716
rect 17289 5660 17293 5716
rect 17229 5656 17293 5660
rect 17414 5713 17478 5717
rect 17414 5657 17418 5713
rect 17418 5657 17474 5713
rect 17474 5657 17478 5713
rect 17414 5653 17478 5657
rect 17605 5715 17669 5719
rect 17605 5659 17609 5715
rect 17609 5659 17665 5715
rect 17665 5659 17669 5715
rect 17605 5655 17669 5659
rect 17796 5719 17860 5723
rect 17796 5663 17800 5719
rect 17800 5663 17856 5719
rect 17856 5663 17860 5719
rect 17796 5659 17860 5663
rect 17982 5715 18046 5719
rect 17982 5659 17986 5715
rect 17986 5659 18042 5715
rect 18042 5659 18046 5715
rect 17982 5655 18046 5659
rect 13429 5132 13493 5136
rect 13429 5076 13433 5132
rect 13433 5076 13489 5132
rect 13489 5076 13493 5132
rect 13429 5072 13493 5076
rect 13634 5128 13698 5132
rect 13634 5072 13638 5128
rect 13638 5072 13694 5128
rect 13694 5072 13698 5128
rect 13634 5068 13698 5072
rect 13820 5133 13884 5137
rect 13820 5077 13824 5133
rect 13824 5077 13880 5133
rect 13880 5077 13884 5133
rect 13820 5073 13884 5077
rect 14014 5126 14078 5130
rect 14014 5070 14018 5126
rect 14018 5070 14074 5126
rect 14074 5070 14078 5126
rect 14014 5066 14078 5070
rect 14233 5131 14297 5135
rect 14233 5075 14237 5131
rect 14237 5075 14293 5131
rect 14293 5075 14297 5131
rect 14233 5071 14297 5075
rect 14443 5131 14507 5135
rect 14443 5075 14447 5131
rect 14447 5075 14503 5131
rect 14503 5075 14507 5131
rect 14443 5071 14507 5075
rect 14672 5128 14736 5132
rect 14672 5072 14676 5128
rect 14676 5072 14732 5128
rect 14732 5072 14736 5128
rect 14672 5068 14736 5072
rect 14918 5128 14982 5132
rect 14918 5072 14922 5128
rect 14922 5072 14978 5128
rect 14978 5072 14982 5128
rect 14918 5068 14982 5072
rect 15192 5128 15256 5132
rect 15192 5072 15196 5128
rect 15196 5072 15252 5128
rect 15252 5072 15256 5128
rect 15192 5068 15256 5072
rect 15467 5128 15531 5132
rect 15467 5072 15471 5128
rect 15471 5072 15527 5128
rect 15527 5072 15531 5128
rect 15467 5068 15531 5072
rect 15703 5128 15767 5132
rect 15703 5072 15707 5128
rect 15707 5072 15763 5128
rect 15763 5072 15767 5128
rect 15703 5068 15767 5072
rect 15926 5131 15990 5135
rect 15926 5075 15930 5131
rect 15930 5075 15986 5131
rect 15986 5075 15990 5131
rect 15926 5071 15990 5075
rect 16144 5134 16208 5138
rect 16144 5078 16148 5134
rect 16148 5078 16204 5134
rect 16204 5078 16208 5134
rect 16144 5074 16208 5078
rect 16322 5125 16386 5129
rect 16322 5069 16326 5125
rect 16326 5069 16382 5125
rect 16382 5069 16386 5125
rect 16322 5065 16386 5069
rect 16561 5127 16625 5131
rect 16561 5071 16565 5127
rect 16565 5071 16621 5127
rect 16621 5071 16625 5127
rect 16561 5067 16625 5071
rect 16758 5127 16822 5131
rect 16758 5071 16762 5127
rect 16762 5071 16818 5127
rect 16818 5071 16822 5127
rect 16758 5067 16822 5071
rect 16956 5127 17020 5131
rect 16956 5071 16960 5127
rect 16960 5071 17016 5127
rect 17016 5071 17020 5127
rect 16956 5067 17020 5071
rect 17169 5128 17233 5132
rect 17169 5072 17173 5128
rect 17173 5072 17229 5128
rect 17229 5072 17233 5128
rect 17169 5068 17233 5072
rect 17392 5127 17456 5131
rect 17392 5071 17396 5127
rect 17396 5071 17452 5127
rect 17452 5071 17456 5127
rect 17392 5067 17456 5071
rect 17589 5132 17653 5136
rect 17589 5076 17593 5132
rect 17593 5076 17649 5132
rect 17649 5076 17653 5132
rect 17589 5072 17653 5076
rect 17805 5130 17869 5134
rect 17805 5074 17809 5130
rect 17809 5074 17865 5130
rect 17865 5074 17869 5130
rect 17805 5070 17869 5074
rect 18014 5130 18078 5134
rect 18014 5074 18018 5130
rect 18018 5074 18074 5130
rect 18074 5074 18078 5130
rect 18014 5070 18078 5074
<< metal4 >>
rect 12437 10623 12563 10628
rect 11836 10618 19041 10623
rect 11836 10554 12468 10618
rect 12532 10611 19041 10618
rect 12532 10608 13297 10611
rect 12532 10554 12565 10608
rect 11836 10545 12565 10554
rect 11836 10013 12254 10545
rect 12461 10544 12565 10545
rect 12629 10544 12645 10608
rect 12709 10544 12725 10608
rect 12789 10544 12805 10608
rect 12869 10544 12885 10608
rect 12949 10544 12965 10608
rect 13029 10547 13297 10608
rect 13361 10547 13377 10611
rect 13441 10547 13457 10611
rect 13521 10547 13537 10611
rect 13601 10547 13617 10611
rect 13681 10547 13697 10611
rect 13761 10547 13903 10611
rect 13967 10547 13983 10611
rect 14047 10547 14063 10611
rect 14127 10547 14143 10611
rect 14207 10547 14223 10611
rect 14287 10547 14303 10611
rect 14367 10547 14509 10611
rect 14573 10547 14589 10611
rect 14653 10547 14669 10611
rect 14733 10547 14749 10611
rect 14813 10547 14829 10611
rect 14893 10547 14909 10611
rect 14973 10547 15115 10611
rect 15179 10547 15195 10611
rect 15259 10547 15275 10611
rect 15339 10547 15355 10611
rect 15419 10547 15435 10611
rect 15499 10547 15515 10611
rect 15579 10547 15721 10611
rect 15785 10547 15801 10611
rect 15865 10547 15881 10611
rect 15945 10547 15961 10611
rect 16025 10547 16041 10611
rect 16105 10547 16121 10611
rect 16185 10547 16327 10611
rect 16391 10547 16407 10611
rect 16471 10547 16487 10611
rect 16551 10547 16567 10611
rect 16631 10547 16647 10611
rect 16711 10547 16727 10611
rect 16791 10547 16933 10611
rect 16997 10547 17013 10611
rect 17077 10547 17093 10611
rect 17157 10547 17173 10611
rect 17237 10547 17253 10611
rect 17317 10547 17333 10611
rect 17397 10547 17539 10611
rect 17603 10547 17619 10611
rect 17683 10547 17699 10611
rect 17763 10547 17779 10611
rect 17843 10547 17859 10611
rect 17923 10547 17939 10611
rect 18003 10556 19041 10611
rect 18003 10547 18277 10556
rect 13029 10545 18277 10547
rect 13029 10544 13134 10545
rect 12461 10543 13134 10544
rect 12461 10542 13133 10543
rect 11836 9949 11851 10013
rect 11915 10012 12126 10013
rect 11915 9949 11982 10012
rect 11836 9948 11982 9949
rect 12046 9949 12126 10012
rect 12190 10007 12254 10013
rect 12461 10388 12527 10478
rect 12461 10324 12462 10388
rect 12526 10324 12527 10388
rect 12461 10308 12527 10324
rect 12461 10244 12462 10308
rect 12526 10244 12527 10308
rect 12461 10228 12527 10244
rect 12461 10164 12462 10228
rect 12526 10164 12527 10228
rect 12461 10148 12527 10164
rect 12461 10084 12462 10148
rect 12526 10084 12527 10148
rect 12461 10068 12527 10084
rect 12190 9949 12253 10007
rect 12046 9948 12253 9949
rect 11836 9930 12253 9948
rect 12461 10004 12462 10068
rect 12526 10004 12527 10068
rect 12461 9988 12527 10004
rect 12461 9924 12462 9988
rect 12526 9924 12527 9988
rect 12461 9908 12527 9924
rect 12461 9844 12462 9908
rect 12526 9844 12527 9908
rect 12461 9828 12527 9844
rect 12461 9764 12462 9828
rect 12526 9764 12527 9828
rect 12461 9748 12527 9764
rect 12461 9684 12462 9748
rect 12526 9684 12527 9748
rect 12461 9668 12527 9684
rect 12461 9604 12462 9668
rect 12526 9604 12527 9668
rect 11862 9467 12239 9482
rect 11862 9403 11869 9467
rect 11933 9403 11989 9467
rect 12053 9403 12132 9467
rect 12196 9403 12239 9467
rect 12461 9450 12527 9604
rect 12587 9512 12647 10542
rect 12707 9450 12767 10482
rect 12827 9512 12887 10542
rect 12947 9450 13007 10482
rect 13067 10388 13133 10478
rect 13067 10324 13068 10388
rect 13132 10324 13133 10388
rect 13067 10308 13133 10324
rect 13067 10244 13068 10308
rect 13132 10244 13133 10308
rect 13067 10228 13133 10244
rect 13067 10164 13068 10228
rect 13132 10164 13133 10228
rect 13067 10148 13133 10164
rect 13067 10084 13068 10148
rect 13132 10084 13133 10148
rect 13067 10068 13133 10084
rect 13067 10004 13068 10068
rect 13132 10004 13133 10068
rect 13067 9988 13133 10004
rect 13067 9924 13068 9988
rect 13132 9924 13133 9988
rect 13067 9908 13133 9924
rect 13067 9844 13068 9908
rect 13132 9844 13133 9908
rect 13067 9828 13133 9844
rect 13067 9764 13068 9828
rect 13132 9764 13133 9828
rect 13067 9748 13133 9764
rect 13067 9684 13068 9748
rect 13132 9684 13133 9748
rect 13067 9668 13133 9684
rect 13067 9604 13068 9668
rect 13132 9604 13133 9668
rect 13067 9450 13133 9604
rect 12461 9448 13133 9450
rect 11864 8044 12240 9403
rect 12461 9384 12565 9448
rect 12629 9384 12645 9448
rect 12709 9384 12725 9448
rect 12789 9384 12805 9448
rect 12869 9384 12885 9448
rect 12949 9384 12965 9448
rect 13029 9384 13133 9448
rect 13193 10391 13259 10481
rect 13193 10327 13194 10391
rect 13258 10327 13259 10391
rect 13193 10311 13259 10327
rect 13193 10247 13194 10311
rect 13258 10247 13259 10311
rect 13193 10231 13259 10247
rect 13193 10167 13194 10231
rect 13258 10167 13259 10231
rect 13193 10151 13259 10167
rect 13193 10087 13194 10151
rect 13258 10087 13259 10151
rect 13193 10071 13259 10087
rect 13193 10007 13194 10071
rect 13258 10007 13259 10071
rect 13193 9991 13259 10007
rect 13193 9927 13194 9991
rect 13258 9927 13259 9991
rect 13193 9911 13259 9927
rect 13193 9847 13194 9911
rect 13258 9847 13259 9911
rect 13193 9831 13259 9847
rect 13193 9767 13194 9831
rect 13258 9767 13259 9831
rect 13193 9751 13259 9767
rect 13193 9687 13194 9751
rect 13258 9687 13259 9751
rect 13193 9671 13259 9687
rect 13193 9607 13194 9671
rect 13258 9607 13259 9671
rect 13193 9453 13259 9607
rect 13319 9515 13379 10545
rect 13439 9453 13499 10485
rect 13559 9515 13619 10545
rect 13679 9453 13739 10485
rect 13799 10391 13865 10481
rect 13799 10327 13800 10391
rect 13864 10327 13865 10391
rect 13799 10311 13865 10327
rect 13799 10247 13800 10311
rect 13864 10247 13865 10311
rect 13799 10231 13865 10247
rect 13799 10167 13800 10231
rect 13864 10167 13865 10231
rect 13799 10151 13865 10167
rect 13799 10087 13800 10151
rect 13864 10087 13865 10151
rect 13799 10071 13865 10087
rect 13799 10007 13800 10071
rect 13864 10007 13865 10071
rect 13799 9991 13865 10007
rect 13799 9927 13800 9991
rect 13864 9927 13865 9991
rect 13799 9911 13865 9927
rect 13799 9847 13800 9911
rect 13864 9847 13865 9911
rect 13799 9831 13865 9847
rect 13799 9767 13800 9831
rect 13864 9767 13865 9831
rect 13799 9751 13865 9767
rect 13799 9687 13800 9751
rect 13864 9687 13865 9751
rect 13799 9671 13865 9687
rect 13799 9607 13800 9671
rect 13864 9607 13865 9671
rect 13799 9453 13865 9607
rect 13925 9453 13985 10485
rect 14045 9515 14105 10545
rect 14165 9453 14225 10485
rect 14285 9515 14345 10545
rect 14405 10391 14471 10481
rect 14405 10327 14406 10391
rect 14470 10327 14471 10391
rect 14405 10311 14471 10327
rect 14405 10247 14406 10311
rect 14470 10247 14471 10311
rect 14405 10231 14471 10247
rect 14405 10167 14406 10231
rect 14470 10167 14471 10231
rect 14405 10151 14471 10167
rect 14405 10087 14406 10151
rect 14470 10087 14471 10151
rect 14405 10071 14471 10087
rect 14405 10007 14406 10071
rect 14470 10007 14471 10071
rect 14405 9991 14471 10007
rect 14405 9927 14406 9991
rect 14470 9927 14471 9991
rect 14405 9911 14471 9927
rect 14405 9847 14406 9911
rect 14470 9847 14471 9911
rect 14405 9831 14471 9847
rect 14405 9767 14406 9831
rect 14470 9767 14471 9831
rect 14405 9751 14471 9767
rect 14405 9687 14406 9751
rect 14470 9687 14471 9751
rect 14405 9671 14471 9687
rect 14405 9607 14406 9671
rect 14470 9607 14471 9671
rect 14405 9453 14471 9607
rect 14531 9515 14591 10545
rect 14651 9453 14711 10485
rect 14771 9515 14831 10545
rect 14891 9453 14951 10485
rect 15011 10391 15077 10481
rect 15011 10327 15012 10391
rect 15076 10327 15077 10391
rect 15011 10311 15077 10327
rect 15011 10247 15012 10311
rect 15076 10247 15077 10311
rect 15011 10231 15077 10247
rect 15011 10167 15012 10231
rect 15076 10167 15077 10231
rect 15011 10151 15077 10167
rect 15011 10087 15012 10151
rect 15076 10087 15077 10151
rect 15011 10071 15077 10087
rect 15011 10007 15012 10071
rect 15076 10007 15077 10071
rect 15011 9991 15077 10007
rect 15011 9927 15012 9991
rect 15076 9927 15077 9991
rect 15011 9911 15077 9927
rect 15011 9847 15012 9911
rect 15076 9847 15077 9911
rect 15011 9831 15077 9847
rect 15011 9767 15012 9831
rect 15076 9767 15077 9831
rect 15011 9751 15077 9767
rect 15011 9687 15012 9751
rect 15076 9687 15077 9751
rect 15011 9671 15077 9687
rect 15011 9607 15012 9671
rect 15076 9607 15077 9671
rect 15011 9453 15077 9607
rect 15137 9453 15197 10485
rect 15257 9515 15317 10545
rect 15377 9453 15437 10485
rect 15497 9515 15557 10545
rect 15617 10391 15683 10481
rect 15617 10327 15618 10391
rect 15682 10327 15683 10391
rect 15617 10311 15683 10327
rect 15617 10247 15618 10311
rect 15682 10247 15683 10311
rect 15617 10231 15683 10247
rect 15617 10167 15618 10231
rect 15682 10167 15683 10231
rect 15617 10151 15683 10167
rect 15617 10087 15618 10151
rect 15682 10087 15683 10151
rect 15617 10071 15683 10087
rect 15617 10007 15618 10071
rect 15682 10007 15683 10071
rect 15617 9991 15683 10007
rect 15617 9927 15618 9991
rect 15682 9927 15683 9991
rect 15617 9911 15683 9927
rect 15617 9847 15618 9911
rect 15682 9847 15683 9911
rect 15617 9831 15683 9847
rect 15617 9767 15618 9831
rect 15682 9767 15683 9831
rect 15617 9751 15683 9767
rect 15617 9687 15618 9751
rect 15682 9687 15683 9751
rect 15617 9671 15683 9687
rect 15617 9607 15618 9671
rect 15682 9607 15683 9671
rect 15617 9453 15683 9607
rect 15743 9515 15803 10545
rect 15863 9453 15923 10485
rect 15983 9515 16043 10545
rect 16103 9453 16163 10485
rect 16223 10391 16289 10481
rect 16223 10327 16224 10391
rect 16288 10327 16289 10391
rect 16223 10311 16289 10327
rect 16223 10247 16224 10311
rect 16288 10247 16289 10311
rect 16223 10231 16289 10247
rect 16223 10167 16224 10231
rect 16288 10167 16289 10231
rect 16223 10151 16289 10167
rect 16223 10087 16224 10151
rect 16288 10087 16289 10151
rect 16223 10071 16289 10087
rect 16223 10007 16224 10071
rect 16288 10007 16289 10071
rect 16223 9991 16289 10007
rect 16223 9927 16224 9991
rect 16288 9927 16289 9991
rect 16223 9911 16289 9927
rect 16223 9847 16224 9911
rect 16288 9847 16289 9911
rect 16223 9831 16289 9847
rect 16223 9767 16224 9831
rect 16288 9767 16289 9831
rect 16223 9751 16289 9767
rect 16223 9687 16224 9751
rect 16288 9687 16289 9751
rect 16223 9671 16289 9687
rect 16223 9607 16224 9671
rect 16288 9607 16289 9671
rect 16223 9453 16289 9607
rect 16349 9453 16409 10485
rect 16469 9515 16529 10545
rect 16589 9453 16649 10485
rect 16709 9515 16769 10545
rect 16829 10391 16895 10481
rect 16829 10327 16830 10391
rect 16894 10327 16895 10391
rect 16829 10311 16895 10327
rect 16829 10247 16830 10311
rect 16894 10247 16895 10311
rect 16829 10231 16895 10247
rect 16829 10167 16830 10231
rect 16894 10167 16895 10231
rect 16829 10151 16895 10167
rect 16829 10087 16830 10151
rect 16894 10087 16895 10151
rect 16829 10071 16895 10087
rect 16829 10007 16830 10071
rect 16894 10007 16895 10071
rect 16829 9991 16895 10007
rect 16829 9927 16830 9991
rect 16894 9927 16895 9991
rect 16829 9911 16895 9927
rect 16829 9847 16830 9911
rect 16894 9847 16895 9911
rect 16829 9831 16895 9847
rect 16829 9767 16830 9831
rect 16894 9767 16895 9831
rect 16829 9751 16895 9767
rect 16829 9687 16830 9751
rect 16894 9687 16895 9751
rect 16829 9671 16895 9687
rect 16829 9607 16830 9671
rect 16894 9607 16895 9671
rect 16829 9453 16895 9607
rect 16955 9515 17015 10545
rect 17075 9453 17135 10485
rect 17195 9515 17255 10545
rect 17315 9453 17375 10485
rect 17435 10391 17501 10481
rect 17435 10327 17436 10391
rect 17500 10327 17501 10391
rect 17435 10311 17501 10327
rect 17435 10247 17436 10311
rect 17500 10247 17501 10311
rect 17435 10231 17501 10247
rect 17435 10167 17436 10231
rect 17500 10167 17501 10231
rect 17435 10151 17501 10167
rect 17435 10087 17436 10151
rect 17500 10087 17501 10151
rect 17435 10071 17501 10087
rect 17435 10007 17436 10071
rect 17500 10007 17501 10071
rect 17435 9991 17501 10007
rect 17435 9927 17436 9991
rect 17500 9927 17501 9991
rect 17435 9911 17501 9927
rect 17435 9847 17436 9911
rect 17500 9847 17501 9911
rect 17435 9831 17501 9847
rect 17435 9767 17436 9831
rect 17500 9767 17501 9831
rect 17435 9751 17501 9767
rect 17435 9687 17436 9751
rect 17500 9687 17501 9751
rect 17435 9671 17501 9687
rect 17435 9607 17436 9671
rect 17500 9607 17501 9671
rect 17435 9453 17501 9607
rect 17561 9453 17621 10485
rect 17681 9515 17741 10545
rect 17801 9453 17861 10485
rect 17921 9515 17981 10545
rect 18167 10492 18277 10545
rect 18341 10492 19041 10556
rect 18041 10391 18107 10481
rect 18041 10327 18042 10391
rect 18106 10327 18107 10391
rect 18041 10311 18107 10327
rect 18041 10247 18042 10311
rect 18106 10247 18107 10311
rect 18041 10231 18107 10247
rect 18041 10167 18042 10231
rect 18106 10167 18107 10231
rect 18041 10151 18107 10167
rect 18041 10087 18042 10151
rect 18106 10087 18107 10151
rect 18041 10071 18107 10087
rect 18041 10007 18042 10071
rect 18106 10007 18107 10071
rect 18041 9991 18107 10007
rect 18041 9927 18042 9991
rect 18106 9927 18107 9991
rect 18041 9911 18107 9927
rect 18041 9847 18042 9911
rect 18106 9847 18107 9911
rect 18041 9831 18107 9847
rect 18041 9767 18042 9831
rect 18106 9767 18107 9831
rect 18041 9751 18107 9767
rect 18041 9687 18042 9751
rect 18106 9687 18107 9751
rect 18041 9671 18107 9687
rect 18041 9607 18042 9671
rect 18106 9607 18107 9671
rect 18167 10412 18493 10492
rect 18167 10348 18282 10412
rect 18346 10348 18493 10412
rect 18167 10260 18493 10348
rect 18167 10196 18283 10260
rect 18347 10217 18493 10260
rect 18590 10217 19041 10492
rect 18347 10196 19041 10217
rect 18167 10090 19041 10196
rect 18167 10026 18283 10090
rect 18347 10026 19041 10090
rect 18167 9933 19041 10026
rect 18167 9869 18282 9933
rect 18346 9869 19041 9933
rect 18167 9699 19041 9869
rect 18167 9691 18577 9699
rect 18167 9627 18200 9691
rect 18264 9636 18577 9691
rect 18264 9627 18485 9636
rect 18167 9615 18485 9627
rect 18041 9453 18107 9607
rect 13193 9451 18107 9453
rect 13193 9387 13297 9451
rect 13361 9387 13377 9451
rect 13441 9387 13457 9451
rect 13521 9387 13537 9451
rect 13601 9387 13617 9451
rect 13681 9387 13697 9451
rect 13761 9387 13903 9451
rect 13967 9387 13983 9451
rect 14047 9387 14063 9451
rect 14127 9387 14143 9451
rect 14207 9387 14223 9451
rect 14287 9387 14303 9451
rect 14367 9387 14509 9451
rect 14573 9387 14589 9451
rect 14653 9387 14669 9451
rect 14733 9387 14749 9451
rect 14813 9387 14829 9451
rect 14893 9387 14909 9451
rect 14973 9387 15115 9451
rect 15179 9387 15195 9451
rect 15259 9387 15275 9451
rect 15339 9387 15355 9451
rect 15419 9387 15435 9451
rect 15499 9387 15515 9451
rect 15579 9387 15721 9451
rect 15785 9387 15801 9451
rect 15865 9387 15881 9451
rect 15945 9387 15961 9451
rect 16025 9387 16041 9451
rect 16105 9387 16121 9451
rect 16185 9387 16327 9451
rect 16391 9387 16407 9451
rect 16471 9387 16487 9451
rect 16551 9387 16567 9451
rect 16631 9387 16647 9451
rect 16711 9387 16727 9451
rect 16791 9387 16933 9451
rect 16997 9387 17013 9451
rect 17077 9387 17093 9451
rect 17157 9387 17173 9451
rect 17237 9387 17253 9451
rect 17317 9387 17333 9451
rect 17397 9387 17539 9451
rect 17603 9387 17619 9451
rect 17683 9387 17699 9451
rect 17763 9387 17779 9451
rect 17843 9387 17859 9451
rect 17923 9387 17939 9451
rect 18003 9387 18107 9451
rect 13193 9385 18107 9387
rect 18167 9430 18365 9440
rect 12461 9382 13133 9384
rect 18167 9366 18288 9430
rect 18352 9366 18365 9430
rect 18167 9356 18365 9366
rect 12812 9203 13484 9205
rect 12812 9139 12916 9203
rect 12980 9139 12996 9203
rect 13060 9139 13076 9203
rect 13140 9139 13156 9203
rect 13220 9139 13236 9203
rect 13300 9139 13316 9203
rect 13380 9139 13484 9203
rect 12812 9137 13484 9139
rect 12812 8983 12878 9137
rect 12812 8919 12813 8983
rect 12877 8919 12878 8983
rect 12812 8903 12878 8919
rect 12812 8839 12813 8903
rect 12877 8839 12878 8903
rect 12812 8823 12878 8839
rect 12812 8759 12813 8823
rect 12877 8759 12878 8823
rect 12812 8743 12878 8759
rect 12812 8679 12813 8743
rect 12877 8679 12878 8743
rect 12812 8663 12878 8679
rect 12812 8599 12813 8663
rect 12877 8599 12878 8663
rect 12812 8583 12878 8599
rect 12812 8519 12813 8583
rect 12877 8519 12878 8583
rect 12812 8503 12878 8519
rect 12812 8439 12813 8503
rect 12877 8439 12878 8503
rect 12812 8423 12878 8439
rect 12812 8359 12813 8423
rect 12877 8359 12878 8423
rect 12812 8343 12878 8359
rect 12812 8279 12813 8343
rect 12877 8279 12878 8343
rect 12812 8263 12878 8279
rect 12812 8199 12813 8263
rect 12877 8199 12878 8263
rect 12812 8109 12878 8199
rect 12424 8044 12549 8050
rect 12938 8045 12998 9075
rect 13058 8105 13118 9137
rect 13178 8045 13238 9075
rect 13298 8105 13358 9137
rect 13418 8983 13484 9137
rect 13418 8919 13419 8983
rect 13483 8919 13484 8983
rect 13418 8903 13484 8919
rect 13418 8839 13419 8903
rect 13483 8839 13484 8903
rect 13418 8823 13484 8839
rect 13418 8759 13419 8823
rect 13483 8759 13484 8823
rect 13418 8743 13484 8759
rect 13418 8679 13419 8743
rect 13483 8679 13484 8743
rect 13418 8663 13484 8679
rect 13418 8599 13419 8663
rect 13483 8599 13484 8663
rect 13418 8583 13484 8599
rect 13418 8519 13419 8583
rect 13483 8519 13484 8583
rect 13418 8503 13484 8519
rect 13418 8439 13419 8503
rect 13483 8439 13484 8503
rect 13418 8423 13484 8439
rect 13418 8359 13419 8423
rect 13483 8359 13484 8423
rect 13418 8343 13484 8359
rect 13418 8279 13419 8343
rect 13483 8279 13484 8343
rect 13418 8263 13484 8279
rect 13418 8199 13419 8263
rect 13483 8199 13484 8263
rect 13418 8109 13484 8199
rect 13544 9203 16034 9205
rect 13544 9139 13648 9203
rect 13712 9139 13728 9203
rect 13792 9139 13808 9203
rect 13872 9139 13888 9203
rect 13952 9139 13968 9203
rect 14032 9139 14048 9203
rect 14112 9139 14254 9203
rect 14318 9139 14334 9203
rect 14398 9139 14414 9203
rect 14478 9139 14494 9203
rect 14558 9139 14574 9203
rect 14638 9139 14654 9203
rect 14718 9139 14860 9203
rect 14924 9139 14940 9203
rect 15004 9139 15020 9203
rect 15084 9139 15100 9203
rect 15164 9139 15180 9203
rect 15244 9139 15260 9203
rect 15324 9139 15466 9203
rect 15530 9139 15546 9203
rect 15610 9139 15626 9203
rect 15690 9139 15706 9203
rect 15770 9139 15786 9203
rect 15850 9139 15866 9203
rect 15930 9139 16034 9203
rect 13544 9137 16034 9139
rect 13544 8983 13610 9137
rect 13544 8919 13545 8983
rect 13609 8919 13610 8983
rect 13544 8903 13610 8919
rect 13544 8839 13545 8903
rect 13609 8839 13610 8903
rect 13544 8823 13610 8839
rect 13544 8759 13545 8823
rect 13609 8759 13610 8823
rect 13544 8743 13610 8759
rect 13544 8679 13545 8743
rect 13609 8679 13610 8743
rect 13544 8663 13610 8679
rect 13544 8599 13545 8663
rect 13609 8599 13610 8663
rect 13544 8583 13610 8599
rect 13544 8519 13545 8583
rect 13609 8519 13610 8583
rect 13544 8503 13610 8519
rect 13544 8439 13545 8503
rect 13609 8439 13610 8503
rect 13544 8423 13610 8439
rect 13544 8359 13545 8423
rect 13609 8359 13610 8423
rect 13544 8343 13610 8359
rect 13544 8279 13545 8343
rect 13609 8279 13610 8343
rect 13544 8263 13610 8279
rect 13544 8199 13545 8263
rect 13609 8199 13610 8263
rect 13544 8109 13610 8199
rect 13670 8045 13730 9075
rect 13790 8105 13850 9137
rect 13910 8045 13970 9075
rect 14030 8105 14090 9137
rect 14150 8983 14216 9137
rect 14150 8919 14151 8983
rect 14215 8919 14216 8983
rect 14150 8903 14216 8919
rect 14150 8839 14151 8903
rect 14215 8839 14216 8903
rect 14150 8823 14216 8839
rect 14150 8759 14151 8823
rect 14215 8759 14216 8823
rect 14150 8743 14216 8759
rect 14150 8679 14151 8743
rect 14215 8679 14216 8743
rect 14150 8663 14216 8679
rect 14150 8599 14151 8663
rect 14215 8599 14216 8663
rect 14150 8583 14216 8599
rect 14150 8519 14151 8583
rect 14215 8519 14216 8583
rect 14150 8503 14216 8519
rect 14150 8439 14151 8503
rect 14215 8439 14216 8503
rect 14150 8423 14216 8439
rect 14150 8359 14151 8423
rect 14215 8359 14216 8423
rect 14150 8343 14216 8359
rect 14150 8279 14151 8343
rect 14215 8279 14216 8343
rect 14150 8263 14216 8279
rect 14150 8199 14151 8263
rect 14215 8199 14216 8263
rect 14150 8109 14216 8199
rect 14276 8105 14336 9137
rect 14396 8045 14456 9075
rect 14516 8105 14576 9137
rect 14636 8045 14696 9075
rect 14756 8983 14822 9137
rect 14756 8919 14757 8983
rect 14821 8919 14822 8983
rect 14756 8903 14822 8919
rect 14756 8839 14757 8903
rect 14821 8839 14822 8903
rect 14756 8823 14822 8839
rect 14756 8759 14757 8823
rect 14821 8759 14822 8823
rect 14756 8743 14822 8759
rect 14756 8679 14757 8743
rect 14821 8679 14822 8743
rect 14756 8663 14822 8679
rect 14756 8599 14757 8663
rect 14821 8599 14822 8663
rect 14756 8583 14822 8599
rect 14756 8519 14757 8583
rect 14821 8519 14822 8583
rect 14756 8503 14822 8519
rect 14756 8439 14757 8503
rect 14821 8439 14822 8503
rect 14756 8423 14822 8439
rect 14756 8359 14757 8423
rect 14821 8359 14822 8423
rect 14756 8343 14822 8359
rect 14756 8279 14757 8343
rect 14821 8279 14822 8343
rect 14756 8263 14822 8279
rect 14756 8199 14757 8263
rect 14821 8199 14822 8263
rect 14756 8109 14822 8199
rect 14882 8045 14942 9075
rect 15002 8105 15062 9137
rect 15122 8045 15182 9075
rect 15242 8105 15302 9137
rect 15362 8983 15428 9137
rect 15362 8919 15363 8983
rect 15427 8919 15428 8983
rect 15362 8903 15428 8919
rect 15362 8839 15363 8903
rect 15427 8839 15428 8903
rect 15362 8823 15428 8839
rect 15362 8759 15363 8823
rect 15427 8759 15428 8823
rect 15362 8743 15428 8759
rect 15362 8679 15363 8743
rect 15427 8679 15428 8743
rect 15362 8663 15428 8679
rect 15362 8599 15363 8663
rect 15427 8599 15428 8663
rect 15362 8583 15428 8599
rect 15362 8519 15363 8583
rect 15427 8519 15428 8583
rect 15362 8503 15428 8519
rect 15362 8439 15363 8503
rect 15427 8439 15428 8503
rect 15362 8423 15428 8439
rect 15362 8359 15363 8423
rect 15427 8359 15428 8423
rect 15362 8343 15428 8359
rect 15362 8279 15363 8343
rect 15427 8279 15428 8343
rect 15362 8263 15428 8279
rect 15362 8199 15363 8263
rect 15427 8199 15428 8263
rect 15362 8109 15428 8199
rect 15488 8105 15548 9137
rect 15608 8045 15668 9075
rect 15728 8105 15788 9137
rect 15848 8045 15908 9075
rect 15968 8983 16034 9137
rect 15968 8919 15969 8983
rect 16033 8919 16034 8983
rect 15968 8903 16034 8919
rect 15968 8839 15969 8903
rect 16033 8839 16034 8903
rect 15968 8823 16034 8839
rect 15968 8759 15969 8823
rect 16033 8759 16034 8823
rect 15968 8743 16034 8759
rect 15968 8679 15969 8743
rect 16033 8679 16034 8743
rect 15968 8663 16034 8679
rect 15968 8599 15969 8663
rect 16033 8599 16034 8663
rect 15968 8583 16034 8599
rect 15968 8519 15969 8583
rect 16033 8519 16034 8583
rect 15968 8503 16034 8519
rect 15968 8439 15969 8503
rect 16033 8439 16034 8503
rect 15968 8423 16034 8439
rect 15968 8359 15969 8423
rect 16033 8359 16034 8423
rect 15968 8343 16034 8359
rect 15968 8279 15969 8343
rect 16033 8279 16034 8343
rect 15968 8263 16034 8279
rect 15968 8199 15969 8263
rect 16033 8199 16034 8263
rect 15968 8109 16034 8199
rect 16094 9203 17372 9205
rect 16094 9139 16198 9203
rect 16262 9139 16278 9203
rect 16342 9139 16358 9203
rect 16422 9139 16438 9203
rect 16502 9139 16518 9203
rect 16582 9139 16598 9203
rect 16662 9139 16804 9203
rect 16868 9139 16884 9203
rect 16948 9139 16964 9203
rect 17028 9139 17044 9203
rect 17108 9139 17124 9203
rect 17188 9139 17204 9203
rect 17268 9139 17372 9203
rect 16094 9137 17372 9139
rect 16094 8983 16160 9137
rect 16094 8919 16095 8983
rect 16159 8919 16160 8983
rect 16094 8903 16160 8919
rect 16094 8839 16095 8903
rect 16159 8839 16160 8903
rect 16094 8823 16160 8839
rect 16094 8759 16095 8823
rect 16159 8759 16160 8823
rect 16094 8743 16160 8759
rect 16094 8679 16095 8743
rect 16159 8679 16160 8743
rect 16094 8663 16160 8679
rect 16094 8599 16095 8663
rect 16159 8599 16160 8663
rect 16094 8583 16160 8599
rect 16094 8519 16095 8583
rect 16159 8519 16160 8583
rect 16094 8503 16160 8519
rect 16094 8439 16095 8503
rect 16159 8439 16160 8503
rect 16094 8423 16160 8439
rect 16094 8359 16095 8423
rect 16159 8359 16160 8423
rect 16094 8343 16160 8359
rect 16094 8279 16095 8343
rect 16159 8279 16160 8343
rect 16094 8263 16160 8279
rect 16094 8199 16095 8263
rect 16159 8199 16160 8263
rect 16094 8109 16160 8199
rect 16220 8045 16280 9075
rect 16340 8105 16400 9137
rect 16460 8045 16520 9075
rect 16580 8105 16640 9137
rect 16700 8983 16766 9137
rect 16700 8919 16701 8983
rect 16765 8919 16766 8983
rect 16700 8903 16766 8919
rect 16700 8839 16701 8903
rect 16765 8839 16766 8903
rect 16700 8823 16766 8839
rect 16700 8759 16701 8823
rect 16765 8759 16766 8823
rect 16700 8743 16766 8759
rect 16700 8679 16701 8743
rect 16765 8679 16766 8743
rect 16700 8663 16766 8679
rect 16700 8599 16701 8663
rect 16765 8599 16766 8663
rect 16700 8583 16766 8599
rect 16700 8519 16701 8583
rect 16765 8519 16766 8583
rect 16700 8503 16766 8519
rect 16700 8439 16701 8503
rect 16765 8439 16766 8503
rect 16700 8423 16766 8439
rect 16700 8359 16701 8423
rect 16765 8359 16766 8423
rect 16700 8343 16766 8359
rect 16700 8279 16701 8343
rect 16765 8279 16766 8343
rect 16700 8263 16766 8279
rect 16700 8199 16701 8263
rect 16765 8199 16766 8263
rect 16700 8109 16766 8199
rect 16826 8105 16886 9137
rect 16946 8045 17006 9075
rect 17066 8105 17126 9137
rect 17186 8045 17246 9075
rect 17306 8983 17372 9137
rect 17306 8919 17307 8983
rect 17371 8919 17372 8983
rect 17306 8903 17372 8919
rect 17306 8839 17307 8903
rect 17371 8839 17372 8903
rect 17306 8823 17372 8839
rect 17306 8759 17307 8823
rect 17371 8759 17372 8823
rect 17306 8743 17372 8759
rect 17306 8679 17307 8743
rect 17371 8679 17372 8743
rect 17306 8663 17372 8679
rect 17306 8599 17307 8663
rect 17371 8599 17372 8663
rect 17306 8583 17372 8599
rect 17306 8519 17307 8583
rect 17371 8519 17372 8583
rect 17306 8503 17372 8519
rect 17306 8439 17307 8503
rect 17371 8439 17372 8503
rect 17306 8423 17372 8439
rect 17306 8359 17307 8423
rect 17371 8359 17372 8423
rect 17306 8343 17372 8359
rect 17306 8279 17307 8343
rect 17371 8279 17372 8343
rect 17306 8263 17372 8279
rect 17306 8199 17307 8263
rect 17371 8199 17372 8263
rect 17306 8109 17372 8199
rect 17434 9203 18106 9205
rect 17434 9139 17538 9203
rect 17602 9139 17618 9203
rect 17682 9139 17698 9203
rect 17762 9139 17778 9203
rect 17842 9139 17858 9203
rect 17922 9139 17938 9203
rect 18002 9139 18106 9203
rect 17434 9137 18106 9139
rect 17434 8983 17500 9137
rect 17434 8919 17435 8983
rect 17499 8919 17500 8983
rect 17434 8903 17500 8919
rect 17434 8839 17435 8903
rect 17499 8839 17500 8903
rect 17434 8823 17500 8839
rect 17434 8759 17435 8823
rect 17499 8759 17500 8823
rect 17434 8743 17500 8759
rect 17434 8679 17435 8743
rect 17499 8679 17500 8743
rect 17434 8663 17500 8679
rect 17434 8599 17435 8663
rect 17499 8599 17500 8663
rect 17434 8583 17500 8599
rect 17434 8519 17435 8583
rect 17499 8519 17500 8583
rect 17434 8503 17500 8519
rect 17434 8439 17435 8503
rect 17499 8439 17500 8503
rect 17434 8423 17500 8439
rect 17434 8359 17435 8423
rect 17499 8359 17500 8423
rect 17434 8343 17500 8359
rect 17434 8279 17435 8343
rect 17499 8279 17500 8343
rect 17434 8263 17500 8279
rect 17434 8199 17435 8263
rect 17499 8199 17500 8263
rect 17434 8109 17500 8199
rect 17560 8105 17620 9137
rect 17680 8045 17740 9075
rect 17800 8105 17860 9137
rect 17920 8045 17980 9075
rect 18040 8983 18106 9137
rect 18040 8919 18041 8983
rect 18105 8919 18106 8983
rect 18040 8903 18106 8919
rect 18040 8839 18041 8903
rect 18105 8839 18106 8903
rect 18040 8823 18106 8839
rect 18040 8759 18041 8823
rect 18105 8759 18106 8823
rect 18040 8743 18106 8759
rect 18040 8679 18041 8743
rect 18105 8679 18106 8743
rect 18040 8663 18106 8679
rect 18040 8599 18041 8663
rect 18105 8599 18106 8663
rect 18040 8583 18106 8599
rect 18040 8519 18041 8583
rect 18105 8519 18106 8583
rect 18040 8503 18106 8519
rect 18040 8439 18041 8503
rect 18105 8439 18106 8503
rect 18040 8423 18106 8439
rect 18040 8359 18041 8423
rect 18105 8359 18106 8423
rect 18040 8343 18106 8359
rect 18040 8279 18041 8343
rect 18105 8279 18106 8343
rect 18040 8263 18106 8279
rect 18040 8199 18041 8263
rect 18105 8199 18106 8263
rect 18040 8109 18106 8199
rect 18167 9093 18227 9356
rect 18425 9237 18485 9615
rect 18287 9227 18485 9237
rect 18287 9163 18288 9227
rect 18352 9163 18485 9227
rect 18287 9153 18485 9163
rect 18545 9635 18577 9636
rect 18641 9635 18777 9699
rect 18841 9635 19041 9699
rect 18167 9057 18483 9093
rect 18167 8993 18388 9057
rect 18452 8993 18483 9057
rect 18167 8975 18483 8993
rect 18167 8965 18485 8975
rect 18167 8901 18197 8965
rect 18261 8901 18485 8965
rect 12812 8044 13484 8045
rect 13544 8044 16034 8045
rect 16094 8044 17372 8045
rect 17434 8044 18106 8045
rect 18167 8044 18485 8901
rect 11864 8043 18485 8044
rect 11864 8040 12996 8043
rect 11864 7976 12454 8040
rect 12518 7979 12996 8040
rect 13060 7979 13076 8043
rect 13140 7979 13156 8043
rect 13220 7979 13236 8043
rect 13300 7979 13728 8043
rect 13792 7979 13808 8043
rect 13872 7979 13888 8043
rect 13952 7979 13968 8043
rect 14032 7979 14334 8043
rect 14398 7979 14414 8043
rect 14478 7979 14494 8043
rect 14558 7979 14574 8043
rect 14638 7979 14940 8043
rect 15004 7979 15020 8043
rect 15084 7979 15100 8043
rect 15164 7979 15180 8043
rect 15244 7979 15546 8043
rect 15610 7979 15626 8043
rect 15690 7979 15706 8043
rect 15770 7979 15786 8043
rect 15850 7979 16278 8043
rect 16342 7979 16358 8043
rect 16422 7979 16438 8043
rect 16502 7979 16518 8043
rect 16582 7979 16884 8043
rect 16948 7979 16964 8043
rect 17028 7979 17044 8043
rect 17108 7979 17124 8043
rect 17188 7979 17618 8043
rect 17682 7979 17698 8043
rect 17762 7979 17778 8043
rect 17842 7979 17858 8043
rect 17922 7979 18485 8043
rect 12518 7976 18485 7979
rect 11864 7966 18485 7976
rect 11864 7602 18154 7966
rect 11864 7601 16897 7602
rect 11864 7598 14533 7601
rect 11864 7596 14101 7598
rect 11864 7595 13900 7596
rect 11864 7531 13501 7595
rect 13565 7594 13900 7595
rect 13565 7531 13675 7594
rect 11864 7530 13675 7531
rect 13739 7532 13900 7594
rect 13964 7534 14101 7596
rect 14165 7596 14533 7598
rect 14165 7534 14324 7596
rect 13964 7532 14324 7534
rect 14388 7537 14533 7596
rect 14597 7598 15156 7601
rect 14597 7594 14951 7598
rect 14597 7537 14761 7594
rect 14388 7532 14761 7537
rect 13739 7530 14761 7532
rect 14825 7534 14951 7594
rect 15015 7537 15156 7598
rect 15220 7537 15355 7601
rect 15419 7596 15959 7601
rect 15419 7537 15571 7596
rect 15015 7534 15571 7537
rect 14825 7532 15571 7534
rect 15635 7537 15959 7596
rect 16023 7599 16897 7601
rect 16023 7598 16668 7599
rect 16023 7596 16436 7598
rect 16023 7537 16194 7596
rect 15635 7532 16194 7537
rect 16258 7534 16436 7596
rect 16500 7535 16668 7598
rect 16732 7538 16897 7599
rect 16961 7601 18154 7602
rect 16961 7598 18030 7601
rect 16961 7594 17364 7598
rect 16961 7538 17146 7594
rect 16732 7535 17146 7538
rect 16500 7534 17146 7535
rect 16258 7532 17146 7534
rect 14825 7530 17146 7532
rect 17210 7534 17364 7594
rect 17428 7596 18030 7598
rect 17428 7594 17814 7596
rect 17428 7534 17593 7594
rect 17210 7530 17593 7534
rect 17657 7532 17814 7594
rect 17878 7537 18030 7596
rect 18094 7537 18154 7601
rect 17878 7532 18154 7537
rect 17657 7530 18154 7532
rect 11864 7481 18154 7530
rect 12771 6704 13267 7481
rect 14836 7408 14950 7421
rect 14836 7351 14859 7408
rect 13330 7344 14859 7351
rect 14923 7351 14950 7408
rect 17231 7407 17345 7420
rect 15221 7357 15335 7370
rect 15221 7351 15244 7357
rect 14923 7344 15244 7351
rect 13330 7293 15244 7344
rect 15308 7351 15335 7357
rect 17231 7351 17254 7407
rect 15308 7343 17254 7351
rect 17318 7351 17345 7407
rect 17616 7358 17730 7371
rect 17616 7351 17639 7358
rect 17318 7343 17639 7351
rect 15308 7294 17639 7343
rect 17703 7351 17730 7358
rect 18545 7351 19041 9635
rect 17703 7294 19043 7351
rect 15308 7293 19043 7294
rect 13330 7146 19043 7293
rect 13330 7018 19042 7146
rect 13330 7015 14550 7018
rect 13330 7012 14094 7015
rect 13330 6948 13503 7012
rect 13567 7010 13875 7012
rect 13567 6948 13678 7010
rect 13330 6946 13678 6948
rect 13742 6948 13875 7010
rect 13939 6951 14094 7012
rect 14158 7011 14550 7015
rect 14158 6951 14326 7011
rect 13939 6948 14326 6951
rect 13742 6947 14326 6948
rect 14390 6954 14550 7011
rect 14614 7009 19042 7018
rect 14614 7008 17979 7009
rect 14614 7006 17757 7008
rect 14614 6954 14762 7006
rect 14390 6947 14762 6954
rect 13742 6946 14762 6947
rect 13330 6942 14762 6946
rect 14826 7002 17757 7006
rect 14826 6942 14984 7002
rect 13330 6938 14984 6942
rect 15048 7001 17757 7002
rect 15048 6999 16721 7001
rect 15048 6938 15207 6999
rect 13330 6935 15207 6938
rect 15271 6935 15417 6999
rect 15481 6935 15630 6999
rect 15694 6997 16721 6999
rect 15694 6996 16529 6997
rect 15694 6995 16350 6996
rect 15694 6992 16149 6995
rect 15694 6935 15947 6992
rect 13330 6928 15947 6935
rect 16011 6931 16149 6992
rect 16213 6932 16350 6995
rect 16414 6933 16529 6996
rect 16593 6937 16721 6997
rect 16785 6999 17549 7001
rect 16785 6998 17343 6999
rect 16785 6937 16906 6998
rect 16593 6934 16906 6937
rect 16970 6997 17343 6998
rect 16970 6934 17138 6997
rect 16593 6933 17138 6934
rect 17202 6935 17343 6997
rect 17407 6937 17549 6999
rect 17613 6944 17757 7001
rect 17821 6945 17979 7008
rect 18043 6945 19042 7009
rect 17821 6944 19042 6945
rect 17613 6937 19042 6944
rect 17407 6935 19042 6937
rect 17202 6933 19042 6935
rect 16414 6932 19042 6933
rect 16213 6931 19042 6932
rect 16011 6928 19042 6931
rect 13330 6866 19042 6928
rect 12771 6372 18193 6704
rect 12771 6369 16873 6372
rect 12771 6368 13952 6369
rect 12771 6363 13746 6368
rect 12771 6299 13530 6363
rect 13594 6304 13746 6363
rect 13810 6305 13952 6368
rect 14016 6366 16650 6369
rect 14016 6365 16205 6366
rect 14016 6363 14575 6365
rect 14016 6361 14350 6363
rect 14016 6305 14154 6361
rect 13810 6304 14154 6305
rect 13594 6299 14154 6304
rect 12771 6297 14154 6299
rect 14218 6299 14350 6361
rect 14414 6301 14575 6363
rect 14639 6364 15673 6365
rect 14639 6361 15233 6364
rect 14639 6301 14790 6361
rect 14414 6299 14790 6301
rect 14218 6297 14790 6299
rect 14854 6297 15025 6361
rect 15089 6300 15233 6361
rect 15297 6300 15475 6364
rect 15539 6301 15673 6364
rect 15737 6301 15980 6365
rect 16044 6302 16205 6365
rect 16269 6365 16650 6366
rect 16269 6302 16434 6365
rect 16044 6301 16434 6302
rect 16498 6305 16650 6365
rect 16714 6308 16873 6369
rect 16937 6368 18193 6372
rect 16937 6308 17097 6368
rect 16714 6305 17097 6308
rect 16498 6304 17097 6305
rect 17161 6361 18193 6368
rect 17161 6360 17975 6361
rect 17161 6357 17748 6360
rect 17161 6304 17324 6357
rect 16498 6301 17324 6304
rect 15539 6300 17324 6301
rect 15089 6297 17324 6300
rect 12771 6293 17324 6297
rect 17388 6356 17748 6357
rect 17388 6293 17537 6356
rect 12771 6292 17537 6293
rect 17601 6296 17748 6356
rect 17812 6297 17975 6360
rect 18039 6297 18193 6361
rect 17812 6296 18193 6297
rect 17601 6292 18193 6296
rect 12771 6219 18193 6292
rect 12771 5525 13267 6219
rect 14841 6134 14955 6147
rect 14841 6076 14864 6134
rect 13327 6070 14864 6076
rect 14928 6076 14955 6134
rect 17233 6136 17347 6149
rect 15224 6076 15338 6088
rect 17233 6076 17256 6136
rect 14928 6075 17256 6076
rect 14928 6070 15247 6075
rect 13327 6011 15247 6070
rect 15311 6072 17256 6075
rect 17320 6076 17347 6136
rect 17610 6082 17724 6095
rect 17610 6076 17633 6082
rect 17320 6072 17633 6076
rect 15311 6018 17633 6072
rect 17697 6076 17724 6082
rect 18545 6076 19041 6866
rect 17697 6018 19043 6076
rect 15311 6011 19043 6018
rect 13327 5894 19043 6011
rect 13327 5785 19042 5894
rect 13327 5736 19043 5785
rect 13327 5734 15633 5736
rect 13327 5732 15420 5734
rect 13327 5728 15182 5732
rect 13327 5727 14750 5728
rect 13327 5718 13781 5727
rect 13327 5654 13556 5718
rect 13620 5663 13781 5718
rect 13845 5724 14279 5727
rect 13845 5663 14058 5724
rect 13620 5660 14058 5663
rect 14122 5663 14279 5724
rect 14343 5724 14750 5727
rect 14343 5663 14524 5724
rect 14122 5660 14524 5663
rect 14588 5664 14750 5724
rect 14814 5726 15182 5728
rect 14814 5664 14962 5726
rect 14588 5662 14962 5664
rect 15026 5668 15182 5726
rect 15246 5670 15420 5732
rect 15484 5672 15633 5734
rect 15697 5727 19043 5736
rect 15697 5726 16367 5727
rect 15697 5672 16020 5726
rect 15484 5670 16020 5672
rect 15246 5668 16020 5670
rect 15026 5662 16020 5668
rect 16084 5663 16367 5726
rect 16431 5724 19043 5727
rect 16431 5722 17026 5724
rect 16431 5663 16603 5722
rect 16084 5662 16603 5663
rect 14588 5660 16603 5662
rect 13620 5658 16603 5660
rect 16667 5658 16787 5722
rect 16851 5660 17026 5722
rect 17090 5723 19043 5724
rect 17090 5720 17796 5723
rect 17090 5660 17229 5720
rect 16851 5658 17229 5660
rect 13620 5656 17229 5658
rect 17293 5719 17796 5720
rect 17293 5717 17605 5719
rect 17293 5656 17414 5717
rect 13620 5654 17414 5656
rect 13327 5653 17414 5654
rect 17478 5655 17605 5717
rect 17669 5659 17796 5719
rect 17860 5719 19043 5723
rect 17860 5659 17982 5719
rect 17669 5655 17982 5659
rect 18046 5655 19043 5719
rect 17478 5653 19043 5655
rect 13327 5591 19043 5653
rect 12771 5138 18195 5525
rect 12771 5137 16144 5138
rect 12771 5136 13820 5137
rect 12771 5072 13429 5136
rect 13493 5132 13820 5136
rect 13493 5072 13634 5132
rect 12771 5068 13634 5072
rect 13698 5073 13820 5132
rect 13884 5135 16144 5137
rect 13884 5130 14233 5135
rect 13884 5073 14014 5130
rect 13698 5068 14014 5073
rect 12771 5066 14014 5068
rect 14078 5071 14233 5130
rect 14297 5071 14443 5135
rect 14507 5132 15926 5135
rect 14507 5071 14672 5132
rect 14078 5068 14672 5071
rect 14736 5068 14918 5132
rect 14982 5068 15192 5132
rect 15256 5068 15467 5132
rect 15531 5068 15703 5132
rect 15767 5071 15926 5132
rect 15990 5074 16144 5135
rect 16208 5136 18195 5138
rect 16208 5132 17589 5136
rect 16208 5131 17169 5132
rect 16208 5129 16561 5131
rect 16208 5074 16322 5129
rect 15990 5071 16322 5074
rect 15767 5068 16322 5071
rect 14078 5066 16322 5068
rect 12771 5065 16322 5066
rect 16386 5067 16561 5129
rect 16625 5067 16758 5131
rect 16822 5067 16956 5131
rect 17020 5068 17169 5131
rect 17233 5131 17589 5132
rect 17233 5068 17392 5131
rect 17020 5067 17392 5068
rect 17456 5072 17589 5131
rect 17653 5134 18195 5136
rect 17653 5072 17805 5134
rect 17456 5070 17805 5072
rect 17869 5070 18014 5134
rect 18078 5070 18195 5134
rect 17456 5067 18195 5070
rect 16386 5065 18195 5067
rect 12771 5040 18195 5065
<< labels >>
flabel metal4 11864 7966 12240 9403 0 FreeSans 320 0 0 0 VSS
port 5 nsew
flabel metal4 11836 10013 12254 10623 0 FreeSans 320 0 0 0 VDD
port 2 nsew
flabel metal1 11767 9271 11864 9318 0 FreeSans 320 0 0 0 eob
port 4 nsew
flabel metal1 12030 9069 12142 9117 0 FreeSans 320 0 0 0 delay_offset
flabel metal1 13338 7918 14277 7946 0 FreeSans 320 0 0 0 delay_code[2]
port 6 nsew
flabel metal1 13338 7862 16703 7890 0 FreeSans 320 0 0 0 delay_code[1]
port 7 nsew
flabel metal1 13338 7806 17560 7834 0 FreeSans 320 0 0 0 delay_code[0]
port 8 nsew
flabel metal1 11730 9654 11784 9688 0 FreeSans 320 0 0 0 delay_code[3]
port 9 nsew
flabel metal1 13297 7232 13342 7280 0 FreeSans 320 0 0 0 sar_logic[0]
flabel metal1 13289 7438 13334 7486 0 FreeSans 320 0 0 0 sar_logic[1]
port 10 nsew
flabel metal1 13307 6591 13352 6639 0 FreeSans 320 0 0 0 sar_logic[2]
port 11 nsew
flabel metal1 13298 5954 13343 6002 0 FreeSans 320 0 0 0 sar_logic[4]
port 14 nsew
flabel metal1 13297 6157 13342 6205 0 FreeSans 320 0 0 0 sar_logic[5]
port 13 nsew
flabel metal1 18207 7428 18252 7476 0 FreeSans 320 0 0 0 sar_retimer[1]
port 17 nsew
flabel metal1 18207 7098 18252 7146 0 FreeSans 320 0 0 0 sar_retimer[0]
port 18 nsew
flabel metal1 18212 6457 18257 6505 0 FreeSans 320 0 0 0 sar_retimer[3]
port 19 nsew
flabel metal1 18207 6799 18252 6847 0 FreeSans 320 0 0 0 sar_retimer[2]
port 20 nsew
flabel metal1 18203 6147 18248 6195 0 FreeSans 320 0 0 0 sar_retimer[5]
port 21 nsew
flabel metal1 18206 5816 18251 5864 0 FreeSans 320 0 0 0 sar_retimer[4]
port 22 nsew
flabel metal1 18205 5176 18250 5224 0 FreeSans 320 0 0 0 sar_retimer[7]
port 23 nsew
flabel metal1 18209 5520 18254 5568 0 FreeSans 320 0 0 0 sar_retimer[6]
port 25 nsew
flabel metal1 13285 5376 13330 5424 0 FreeSans 320 0 0 0 sar_retimer[6]
port 26 nsew
flabel metal1 13282 5177 13327 5225 0 FreeSans 320 0 0 0 sar_retimer[7]
port 27 nsew
flabel metal1 13310 6457 13355 6505 0 FreeSans 320 0 0 0 sar_logic[3]
port 28 nsew
flabel locali 15233 7299 15308 7345 0 FreeSans 400 0 0 0 x1[0].RESET_B
flabel locali 13400 7547 13434 7581 3 FreeSans 400 0 0 0 x1[0].VGND
flabel locali 13400 7309 13434 7343 0 FreeSans 400 0 0 0 x1[0].CLK
flabel locali 13400 7241 13434 7275 0 FreeSans 400 0 0 0 x1[0].CLK
flabel locali 14136 7377 14170 7411 0 FreeSans 400 0 0 0 x1[0].SET_B
flabel locali 15698 7445 15732 7479 0 FreeSans 400 0 0 0 x1[0].Q
flabel locali 15698 7173 15732 7207 0 FreeSans 400 0 0 0 x1[0].Q
flabel locali 15698 7105 15732 7139 0 FreeSans 400 0 0 0 x1[0].Q
flabel locali 13400 7003 13434 7037 3 FreeSans 400 0 0 0 x1[0].VPWR
flabel locali 13768 7309 13802 7343 0 FreeSans 200 0 0 0 x1[0].D
flabel locali 13768 7241 13802 7275 0 FreeSans 200 0 0 0 x1[0].D
flabel locali 15418 7105 15452 7139 0 FreeSans 400 0 0 0 x1[0].Q_N
flabel locali 15418 7173 15452 7207 0 FreeSans 400 0 0 0 x1[0].Q_N
flabel locali 15418 7445 15452 7479 0 FreeSans 400 0 0 0 x1[0].Q_N
flabel metal1 13400 7547 13434 7581 0 FreeSans 200 0 0 0 x1[0].VGND
flabel metal1 13400 7003 13434 7037 0 FreeSans 200 0 0 0 x1[0].VPWR
flabel nwell 13400 7003 13434 7037 3 FreeSans 400 0 0 0 x1[0].VPB
flabel nwell 13417 7020 13417 7020 0 FreeSans 200 0 0 0 x1[0].VPB
flabel pwell 13400 7547 13434 7581 3 FreeSans 400 0 0 0 x1[0].VNB
flabel pwell 13417 7564 13417 7564 0 FreeSans 200 0 0 0 x1[0].VNB
rlabel comment 13370 7564 13370 7564 2 x1[0].dfbbp_1
rlabel locali 14862 7351 14937 7417 5 x1[0].SET_B
rlabel metal1 14860 7371 14918 7380 5 x1[0].SET_B
rlabel metal1 14860 7408 14918 7417 5 x1[0].SET_B
rlabel metal1 14124 7371 14182 7380 5 x1[0].SET_B
rlabel metal1 14124 7380 14918 7408 5 x1[0].SET_B
rlabel metal1 14124 7408 14182 7417 5 x1[0].SET_B
rlabel metal1 13370 7516 15762 7612 5 x1[0].VGND
rlabel metal1 13370 6972 15762 7068 5 x1[0].VPWR
flabel locali 17625 7299 17700 7345 0 FreeSans 400 0 0 0 x1[1].RESET_B
flabel locali 15792 7547 15826 7581 3 FreeSans 400 0 0 0 x1[1].VGND
flabel locali 15792 7309 15826 7343 0 FreeSans 400 0 0 0 x1[1].CLK
flabel locali 15792 7241 15826 7275 0 FreeSans 400 0 0 0 x1[1].CLK
flabel locali 16528 7377 16562 7411 0 FreeSans 400 0 0 0 x1[1].SET_B
flabel locali 18090 7445 18124 7479 0 FreeSans 400 0 0 0 x1[1].Q
flabel locali 18090 7173 18124 7207 0 FreeSans 400 0 0 0 x1[1].Q
flabel locali 18090 7105 18124 7139 0 FreeSans 400 0 0 0 x1[1].Q
flabel locali 15792 7003 15826 7037 3 FreeSans 400 0 0 0 x1[1].VPWR
flabel locali 16160 7309 16194 7343 0 FreeSans 200 0 0 0 x1[1].D
flabel locali 16160 7241 16194 7275 0 FreeSans 200 0 0 0 x1[1].D
flabel locali 17810 7105 17844 7139 0 FreeSans 400 0 0 0 x1[1].Q_N
flabel locali 17810 7173 17844 7207 0 FreeSans 400 0 0 0 x1[1].Q_N
flabel locali 17810 7445 17844 7479 0 FreeSans 400 0 0 0 x1[1].Q_N
flabel metal1 15792 7547 15826 7581 0 FreeSans 200 0 0 0 x1[1].VGND
flabel metal1 15792 7003 15826 7037 0 FreeSans 200 0 0 0 x1[1].VPWR
flabel nwell 15792 7003 15826 7037 3 FreeSans 400 0 0 0 x1[1].VPB
flabel nwell 15809 7020 15809 7020 0 FreeSans 200 0 0 0 x1[1].VPB
flabel pwell 15792 7547 15826 7581 3 FreeSans 400 0 0 0 x1[1].VNB
flabel pwell 15809 7564 15809 7564 0 FreeSans 200 0 0 0 x1[1].VNB
rlabel comment 15762 7564 15762 7564 2 x1[1].dfbbp_1
rlabel locali 17254 7351 17329 7417 5 x1[1].SET_B
rlabel metal1 17252 7371 17310 7380 5 x1[1].SET_B
rlabel metal1 17252 7408 17310 7417 5 x1[1].SET_B
rlabel metal1 16516 7371 16574 7380 5 x1[1].SET_B
rlabel metal1 16516 7380 17310 7408 5 x1[1].SET_B
rlabel metal1 16516 7408 16574 7417 5 x1[1].SET_B
rlabel metal1 15762 7516 18154 7612 5 x1[1].VGND
rlabel metal1 15762 6972 18154 7068 5 x1[1].VPWR
flabel locali 15233 6599 15308 6645 0 FreeSans 400 0 0 0 x1[2].RESET_B
flabel locali 13400 6363 13434 6397 3 FreeSans 400 0 0 0 x1[2].VGND
flabel locali 13400 6601 13434 6635 0 FreeSans 400 0 0 0 x1[2].CLK
flabel locali 13400 6669 13434 6703 0 FreeSans 400 0 0 0 x1[2].CLK
flabel locali 14136 6533 14170 6567 0 FreeSans 400 0 0 0 x1[2].SET_B
flabel locali 15698 6465 15732 6499 0 FreeSans 400 0 0 0 x1[2].Q
flabel locali 15698 6737 15732 6771 0 FreeSans 400 0 0 0 x1[2].Q
flabel locali 15698 6805 15732 6839 0 FreeSans 400 0 0 0 x1[2].Q
flabel locali 13400 6907 13434 6941 3 FreeSans 400 0 0 0 x1[2].VPWR
flabel locali 13768 6601 13802 6635 0 FreeSans 200 0 0 0 x1[2].D
flabel locali 13768 6669 13802 6703 0 FreeSans 200 0 0 0 x1[2].D
flabel locali 15418 6805 15452 6839 0 FreeSans 400 0 0 0 x1[2].Q_N
flabel locali 15418 6737 15452 6771 0 FreeSans 400 0 0 0 x1[2].Q_N
flabel locali 15418 6465 15452 6499 0 FreeSans 400 0 0 0 x1[2].Q_N
flabel metal1 13400 6363 13434 6397 0 FreeSans 200 0 0 0 x1[2].VGND
flabel metal1 13400 6907 13434 6941 0 FreeSans 200 0 0 0 x1[2].VPWR
flabel nwell 13400 6907 13434 6941 3 FreeSans 400 0 0 0 x1[2].VPB
flabel nwell 13417 6924 13417 6924 0 FreeSans 200 0 0 0 x1[2].VPB
flabel pwell 13400 6363 13434 6397 3 FreeSans 400 0 0 0 x1[2].VNB
flabel pwell 13417 6380 13417 6380 0 FreeSans 200 0 0 0 x1[2].VNB
rlabel comment 13370 6380 13370 6380 4 x1[2].dfbbp_1
rlabel locali 14862 6527 14937 6593 1 x1[2].SET_B
rlabel metal1 14860 6564 14918 6573 1 x1[2].SET_B
rlabel metal1 14860 6527 14918 6536 1 x1[2].SET_B
rlabel metal1 14124 6564 14182 6573 1 x1[2].SET_B
rlabel metal1 14124 6536 14918 6564 1 x1[2].SET_B
rlabel metal1 14124 6527 14182 6536 1 x1[2].SET_B
rlabel metal1 13370 6332 15762 6428 1 x1[2].VGND
rlabel metal1 13370 6876 15762 6972 1 x1[2].VPWR
flabel locali 17625 6599 17700 6645 0 FreeSans 400 0 0 0 x1[3].RESET_B
flabel locali 15792 6363 15826 6397 3 FreeSans 400 0 0 0 x1[3].VGND
flabel locali 15792 6601 15826 6635 0 FreeSans 400 0 0 0 x1[3].CLK
flabel locali 15792 6669 15826 6703 0 FreeSans 400 0 0 0 x1[3].CLK
flabel locali 16528 6533 16562 6567 0 FreeSans 400 0 0 0 x1[3].SET_B
flabel locali 18090 6465 18124 6499 0 FreeSans 400 0 0 0 x1[3].Q
flabel locali 18090 6737 18124 6771 0 FreeSans 400 0 0 0 x1[3].Q
flabel locali 18090 6805 18124 6839 0 FreeSans 400 0 0 0 x1[3].Q
flabel locali 15792 6907 15826 6941 3 FreeSans 400 0 0 0 x1[3].VPWR
flabel locali 16160 6601 16194 6635 0 FreeSans 200 0 0 0 x1[3].D
flabel locali 16160 6669 16194 6703 0 FreeSans 200 0 0 0 x1[3].D
flabel locali 17810 6805 17844 6839 0 FreeSans 400 0 0 0 x1[3].Q_N
flabel locali 17810 6737 17844 6771 0 FreeSans 400 0 0 0 x1[3].Q_N
flabel locali 17810 6465 17844 6499 0 FreeSans 400 0 0 0 x1[3].Q_N
flabel metal1 15792 6363 15826 6397 0 FreeSans 200 0 0 0 x1[3].VGND
flabel metal1 15792 6907 15826 6941 0 FreeSans 200 0 0 0 x1[3].VPWR
flabel nwell 15792 6907 15826 6941 3 FreeSans 400 0 0 0 x1[3].VPB
flabel nwell 15809 6924 15809 6924 0 FreeSans 200 0 0 0 x1[3].VPB
flabel pwell 15792 6363 15826 6397 3 FreeSans 400 0 0 0 x1[3].VNB
flabel pwell 15809 6380 15809 6380 0 FreeSans 200 0 0 0 x1[3].VNB
rlabel comment 15762 6380 15762 6380 4 x1[3].dfbbp_1
rlabel locali 17254 6527 17329 6593 1 x1[3].SET_B
rlabel metal1 17252 6564 17310 6573 1 x1[3].SET_B
rlabel metal1 17252 6527 17310 6536 1 x1[3].SET_B
rlabel metal1 16516 6564 16574 6573 1 x1[3].SET_B
rlabel metal1 16516 6536 17310 6564 1 x1[3].SET_B
rlabel metal1 16516 6527 16574 6536 1 x1[3].SET_B
rlabel metal1 15762 6332 18154 6428 1 x1[3].VGND
rlabel metal1 15762 6876 18154 6972 1 x1[3].VPWR
flabel locali 15233 6019 15308 6065 0 FreeSans 400 0 0 0 x1[4].RESET_B
flabel locali 13400 6267 13434 6301 3 FreeSans 400 0 0 0 x1[4].VGND
flabel locali 13400 6029 13434 6063 0 FreeSans 400 0 0 0 x1[4].CLK
flabel locali 13400 5961 13434 5995 0 FreeSans 400 0 0 0 x1[4].CLK
flabel locali 14136 6097 14170 6131 0 FreeSans 400 0 0 0 x1[4].SET_B
flabel locali 15698 6165 15732 6199 0 FreeSans 400 0 0 0 x1[4].Q
flabel locali 15698 5893 15732 5927 0 FreeSans 400 0 0 0 x1[4].Q
flabel locali 15698 5825 15732 5859 0 FreeSans 400 0 0 0 x1[4].Q
flabel locali 13400 5723 13434 5757 3 FreeSans 400 0 0 0 x1[4].VPWR
flabel locali 13768 6029 13802 6063 0 FreeSans 200 0 0 0 x1[4].D
flabel locali 13768 5961 13802 5995 0 FreeSans 200 0 0 0 x1[4].D
flabel locali 15418 5825 15452 5859 0 FreeSans 400 0 0 0 x1[4].Q_N
flabel locali 15418 5893 15452 5927 0 FreeSans 400 0 0 0 x1[4].Q_N
flabel locali 15418 6165 15452 6199 0 FreeSans 400 0 0 0 x1[4].Q_N
flabel metal1 13400 6267 13434 6301 0 FreeSans 200 0 0 0 x1[4].VGND
flabel metal1 13400 5723 13434 5757 0 FreeSans 200 0 0 0 x1[4].VPWR
flabel nwell 13400 5723 13434 5757 3 FreeSans 400 0 0 0 x1[4].VPB
flabel nwell 13417 5740 13417 5740 0 FreeSans 200 0 0 0 x1[4].VPB
flabel pwell 13400 6267 13434 6301 3 FreeSans 400 0 0 0 x1[4].VNB
flabel pwell 13417 6284 13417 6284 0 FreeSans 200 0 0 0 x1[4].VNB
rlabel comment 13370 6284 13370 6284 2 x1[4].dfbbp_1
rlabel locali 14862 6071 14937 6137 5 x1[4].SET_B
rlabel metal1 14860 6091 14918 6100 5 x1[4].SET_B
rlabel metal1 14860 6128 14918 6137 5 x1[4].SET_B
rlabel metal1 14124 6091 14182 6100 5 x1[4].SET_B
rlabel metal1 14124 6100 14918 6128 5 x1[4].SET_B
rlabel metal1 14124 6128 14182 6137 5 x1[4].SET_B
rlabel metal1 13370 6236 15762 6332 5 x1[4].VGND
rlabel metal1 13370 5692 15762 5788 5 x1[4].VPWR
flabel locali 17625 6019 17700 6065 0 FreeSans 400 0 0 0 x1[5].RESET_B
flabel locali 15792 6267 15826 6301 3 FreeSans 400 0 0 0 x1[5].VGND
flabel locali 15792 6029 15826 6063 0 FreeSans 400 0 0 0 x1[5].CLK
flabel locali 15792 5961 15826 5995 0 FreeSans 400 0 0 0 x1[5].CLK
flabel locali 16528 6097 16562 6131 0 FreeSans 400 0 0 0 x1[5].SET_B
flabel locali 18090 6165 18124 6199 0 FreeSans 400 0 0 0 x1[5].Q
flabel locali 18090 5893 18124 5927 0 FreeSans 400 0 0 0 x1[5].Q
flabel locali 18090 5825 18124 5859 0 FreeSans 400 0 0 0 x1[5].Q
flabel locali 15792 5723 15826 5757 3 FreeSans 400 0 0 0 x1[5].VPWR
flabel locali 16160 6029 16194 6063 0 FreeSans 200 0 0 0 x1[5].D
flabel locali 16160 5961 16194 5995 0 FreeSans 200 0 0 0 x1[5].D
flabel locali 17810 5825 17844 5859 0 FreeSans 400 0 0 0 x1[5].Q_N
flabel locali 17810 5893 17844 5927 0 FreeSans 400 0 0 0 x1[5].Q_N
flabel locali 17810 6165 17844 6199 0 FreeSans 400 0 0 0 x1[5].Q_N
flabel metal1 15792 6267 15826 6301 0 FreeSans 200 0 0 0 x1[5].VGND
flabel metal1 15792 5723 15826 5757 0 FreeSans 200 0 0 0 x1[5].VPWR
flabel nwell 15792 5723 15826 5757 3 FreeSans 400 0 0 0 x1[5].VPB
flabel nwell 15809 5740 15809 5740 0 FreeSans 200 0 0 0 x1[5].VPB
flabel pwell 15792 6267 15826 6301 3 FreeSans 400 0 0 0 x1[5].VNB
flabel pwell 15809 6284 15809 6284 0 FreeSans 200 0 0 0 x1[5].VNB
rlabel comment 15762 6284 15762 6284 2 x1[5].dfbbp_1
rlabel locali 17254 6071 17329 6137 5 x1[5].SET_B
rlabel metal1 17252 6091 17310 6100 5 x1[5].SET_B
rlabel metal1 17252 6128 17310 6137 5 x1[5].SET_B
rlabel metal1 16516 6091 16574 6100 5 x1[5].SET_B
rlabel metal1 16516 6100 17310 6128 5 x1[5].SET_B
rlabel metal1 16516 6128 16574 6137 5 x1[5].SET_B
rlabel metal1 15762 6236 18154 6332 5 x1[5].VGND
rlabel metal1 15762 5692 18154 5788 5 x1[5].VPWR
flabel locali 15233 5319 15308 5365 0 FreeSans 400 0 0 0 x1[6].RESET_B
flabel locali 13400 5083 13434 5117 3 FreeSans 400 0 0 0 x1[6].VGND
flabel locali 13400 5321 13434 5355 0 FreeSans 400 0 0 0 x1[6].CLK
flabel locali 13400 5389 13434 5423 0 FreeSans 400 0 0 0 x1[6].CLK
flabel locali 14136 5253 14170 5287 0 FreeSans 400 0 0 0 x1[6].SET_B
flabel locali 15698 5185 15732 5219 0 FreeSans 400 0 0 0 x1[6].Q
flabel locali 15698 5457 15732 5491 0 FreeSans 400 0 0 0 x1[6].Q
flabel locali 15698 5525 15732 5559 0 FreeSans 400 0 0 0 x1[6].Q
flabel locali 13400 5627 13434 5661 3 FreeSans 400 0 0 0 x1[6].VPWR
flabel locali 13768 5321 13802 5355 0 FreeSans 200 0 0 0 x1[6].D
flabel locali 13768 5389 13802 5423 0 FreeSans 200 0 0 0 x1[6].D
flabel locali 15418 5525 15452 5559 0 FreeSans 400 0 0 0 x1[6].Q_N
flabel locali 15418 5457 15452 5491 0 FreeSans 400 0 0 0 x1[6].Q_N
flabel locali 15418 5185 15452 5219 0 FreeSans 400 0 0 0 x1[6].Q_N
flabel metal1 13400 5083 13434 5117 0 FreeSans 200 0 0 0 x1[6].VGND
flabel metal1 13400 5627 13434 5661 0 FreeSans 200 0 0 0 x1[6].VPWR
flabel nwell 13400 5627 13434 5661 3 FreeSans 400 0 0 0 x1[6].VPB
flabel nwell 13417 5644 13417 5644 0 FreeSans 200 0 0 0 x1[6].VPB
flabel pwell 13400 5083 13434 5117 3 FreeSans 400 0 0 0 x1[6].VNB
flabel pwell 13417 5100 13417 5100 0 FreeSans 200 0 0 0 x1[6].VNB
rlabel comment 13370 5100 13370 5100 4 x1[6].dfbbp_1
rlabel locali 14862 5247 14937 5313 1 x1[6].SET_B
rlabel metal1 14860 5284 14918 5293 1 x1[6].SET_B
rlabel metal1 14860 5247 14918 5256 1 x1[6].SET_B
rlabel metal1 14124 5284 14182 5293 1 x1[6].SET_B
rlabel metal1 14124 5256 14918 5284 1 x1[6].SET_B
rlabel metal1 14124 5247 14182 5256 1 x1[6].SET_B
rlabel metal1 13370 5052 15762 5148 1 x1[6].VGND
rlabel metal1 13370 5596 15762 5692 1 x1[6].VPWR
flabel locali 17625 5319 17700 5365 0 FreeSans 400 0 0 0 x1[7].RESET_B
flabel locali 15792 5083 15826 5117 3 FreeSans 400 0 0 0 x1[7].VGND
flabel locali 15792 5321 15826 5355 0 FreeSans 400 0 0 0 x1[7].CLK
flabel locali 15792 5389 15826 5423 0 FreeSans 400 0 0 0 x1[7].CLK
flabel locali 16528 5253 16562 5287 0 FreeSans 400 0 0 0 x1[7].SET_B
flabel locali 18090 5185 18124 5219 0 FreeSans 400 0 0 0 x1[7].Q
flabel locali 18090 5457 18124 5491 0 FreeSans 400 0 0 0 x1[7].Q
flabel locali 18090 5525 18124 5559 0 FreeSans 400 0 0 0 x1[7].Q
flabel locali 15792 5627 15826 5661 3 FreeSans 400 0 0 0 x1[7].VPWR
flabel locali 16160 5321 16194 5355 0 FreeSans 200 0 0 0 x1[7].D
flabel locali 16160 5389 16194 5423 0 FreeSans 200 0 0 0 x1[7].D
flabel locali 17810 5525 17844 5559 0 FreeSans 400 0 0 0 x1[7].Q_N
flabel locali 17810 5457 17844 5491 0 FreeSans 400 0 0 0 x1[7].Q_N
flabel locali 17810 5185 17844 5219 0 FreeSans 400 0 0 0 x1[7].Q_N
flabel metal1 15792 5083 15826 5117 0 FreeSans 200 0 0 0 x1[7].VGND
flabel metal1 15792 5627 15826 5661 0 FreeSans 200 0 0 0 x1[7].VPWR
flabel nwell 15792 5627 15826 5661 3 FreeSans 400 0 0 0 x1[7].VPB
flabel nwell 15809 5644 15809 5644 0 FreeSans 200 0 0 0 x1[7].VPB
flabel pwell 15792 5083 15826 5117 3 FreeSans 400 0 0 0 x1[7].VNB
flabel pwell 15809 5100 15809 5100 0 FreeSans 200 0 0 0 x1[7].VNB
rlabel comment 15762 5100 15762 5100 4 x1[7].dfbbp_1
rlabel locali 17254 5247 17329 5313 1 x1[7].SET_B
rlabel metal1 17252 5284 17310 5293 1 x1[7].SET_B
rlabel metal1 17252 5247 17310 5256 1 x1[7].SET_B
rlabel metal1 16516 5284 16574 5293 1 x1[7].SET_B
rlabel metal1 16516 5256 17310 5284 1 x1[7].SET_B
rlabel metal1 16516 5247 16574 5256 1 x1[7].SET_B
rlabel metal1 15762 5052 18154 5148 1 x1[7].VGND
rlabel metal1 15762 5596 18154 5692 1 x1[7].VPWR
flabel metal1 11767 9271 12435 9318 0 FreeSans 320 0 0 0 x2.IN
flabel metal1 18243 9269 18425 9315 0 FreeSans 320 0 0 0 x2.OUT
flabel metal1 11730 9654 11868 9688 0 FreeSans 320 0 0 0 x2.code[3]
flabel metal1 16645 7943 16703 9120 0 FreeSans 320 0 0 0 x2.code[1]
flabel metal1 14219 7943 14277 9120 0 FreeSans 320 0 0 0 x2.code[2]
flabel metal4 11836 10013 12254 10623 0 FreeSans 320 0 0 0 x2.VDD
flabel metal4 11864 7966 12240 9403 0 FreeSans 320 0 0 0 x2.VSS
flabel metal2 12194 9069 12630 9115 0 FreeSans 320 0 0 0 x2.code_offset
flabel metal1 17501 7942 17560 9123 0 FreeSans 320 0 0 0 x2.code[0]
flabel metal1 12378 9724 12412 9758 0 FreeSans 320 0 0 0 x2.x8.input_stack
flabel nwell 12422 10507 12456 10567 0 FreeSans 320 0 0 0 x2.x8.vdd
flabel metal1 12416 9805 12462 9817 0 FreeSans 320 0 0 0 x2.x8.output_stack
flabel poly 12355 9067 12457 9097 0 FreeSans 320 0 0 0 x2.x9.input_stack
flabel metal1 12469 8014 12503 8074 0 FreeSans 320 0 0 0 x2.x9.vss
flabel metal1 12463 9040 12509 9052 0 FreeSans 320 0 0 0 x2.x9.output_stack
flabel locali 11956 9724 11990 9758 0 FreeSans 340 0 0 0 x2.x10.Y
flabel locali 11956 9656 11990 9690 0 FreeSans 340 0 0 0 x2.x10.Y
flabel locali 11864 9656 11898 9690 0 FreeSans 340 0 0 0 x2.x10.A
flabel metal1 11821 9418 11855 9452 0 FreeSans 200 0 0 0 x2.x10.VGND
flabel metal1 11821 9962 11855 9996 0 FreeSans 200 0 0 0 x2.x10.VPWR
rlabel comment 11792 9435 11792 9435 4 x2.x10.inv_1
rlabel metal1 11792 9387 12068 9483 1 x2.x10.VGND
rlabel metal1 11792 9931 12068 10027 1 x2.x10.VPWR
flabel pwell 11821 9418 11855 9452 0 FreeSans 200 0 0 0 x2.x10.VNB
flabel nwell 11821 9962 11855 9996 0 FreeSans 200 0 0 0 x2.x10.VPB
flabel locali 12054 9724 12088 9758 0 FreeSans 340 0 0 0 x2.x11.Y
flabel locali 12054 9656 12088 9690 0 FreeSans 340 0 0 0 x2.x11.Y
flabel locali 12146 9656 12180 9690 0 FreeSans 340 0 0 0 x2.x11.A
flabel metal1 12189 9418 12223 9452 0 FreeSans 200 0 0 0 x2.x11.VGND
flabel metal1 12189 9962 12223 9996 0 FreeSans 200 0 0 0 x2.x11.VPWR
rlabel comment 12252 9435 12252 9435 6 x2.x11.inv_1
rlabel metal1 11976 9387 12252 9483 1 x2.x11.VGND
rlabel metal1 11976 9931 12252 10027 1 x2.x11.VPWR
flabel pwell 12189 9418 12223 9452 0 FreeSans 200 0 0 0 x2.x11.VNB
flabel nwell 12189 9962 12223 9996 0 FreeSans 200 0 0 0 x2.x11.VPB
flabel metal1 13020 9481 13054 9515 0 FreeSans 320 0 0 0 x2.x6.SW
flabel nwell 12464 10543 13134 10611 0 FreeSans 320 0 0 0 x2.x6.VDD
flabel pdiff 13052 9350 13110 9434 0 FreeSans 320 0 0 0 x2.x6.delay_signal
flabel metal4 12464 10542 12565 10611 0 FreeSans 320 0 0 0 x2.x6.VDD
flabel via3 12565 9384 12629 9448 0 FreeSans 320 0 0 0 x2.x6.floating
flabel viali 13373 9080 13407 9114 0 FreeSans 320 0 0 0 x2.x7.SW
flabel ndiff 13405 9152 13463 9236 0 FreeSans 320 0 0 0 x2.x7.delay_signal
flabel metal4 12812 7975 13484 8043 0 FreeSans 320 0 0 0 x2.x7.VSS
flabel via3 12916 9139 12980 9203 0 FreeSans 320 0 0 0 x2.x7.floating
flabel viali 14105 9080 14139 9114 0 FreeSans 320 0 0 0 x2.x4[3].SW
flabel ndiff 14137 9152 14195 9236 0 FreeSans 320 0 0 0 x2.x4[3].delay_signal
flabel metal4 13544 7975 14216 8043 0 FreeSans 320 0 0 0 x2.x4[3].VSS
flabel via3 13648 9139 13712 9203 0 FreeSans 320 0 0 0 x2.x4[3].floating
flabel metal1 13878 9484 13912 9518 0 FreeSans 320 0 0 0 x2.x5[6].SW
flabel nwell 13798 10546 14468 10614 0 FreeSans 320 0 0 0 x2.x5[6].VDD
flabel pdiff 13822 9353 13880 9437 0 FreeSans 320 0 0 0 x2.x5[6].delay_signal
flabel metal4 14367 10545 14468 10614 0 FreeSans 320 0 0 0 x2.x5[6].VDD
flabel via3 14303 9387 14367 9451 0 FreeSans 320 0 0 0 x2.x5[6].floating
flabel metal1 13752 9484 13786 9518 0 FreeSans 320 0 0 0 x2.x5[7].SW
flabel nwell 13196 10546 13866 10614 0 FreeSans 320 0 0 0 x2.x5[7].VDD
flabel pdiff 13784 9353 13842 9437 0 FreeSans 320 0 0 0 x2.x5[7].delay_signal
flabel metal4 13196 10545 13297 10614 0 FreeSans 320 0 0 0 x2.x5[7].VDD
flabel via3 13297 9387 13361 9451 0 FreeSans 320 0 0 0 x2.x5[7].floating
flabel viali 14227 9080 14261 9114 0 FreeSans 320 0 0 0 x2.x4[2].SW
flabel ndiff 14171 9152 14229 9236 0 FreeSans 320 0 0 0 x2.x4[2].delay_signal
flabel metal4 14150 7975 14822 8043 0 FreeSans 320 0 0 0 x2.x4[2].VSS
flabel via3 14654 9139 14718 9203 0 FreeSans 320 0 0 0 x2.x4[2].floating
flabel metal1 14964 9484 14998 9518 0 FreeSans 320 0 0 0 x2.x5[5].SW
flabel nwell 14408 10546 15078 10614 0 FreeSans 320 0 0 0 x2.x5[5].VDD
flabel pdiff 14996 9353 15054 9437 0 FreeSans 320 0 0 0 x2.x5[5].delay_signal
flabel metal4 14408 10545 14509 10614 0 FreeSans 320 0 0 0 x2.x5[5].VDD
flabel via3 14509 9387 14573 9451 0 FreeSans 320 0 0 0 x2.x5[5].floating
flabel viali 15317 9080 15351 9114 0 FreeSans 320 0 0 0 x2.x4[1].SW
flabel ndiff 15349 9152 15407 9236 0 FreeSans 320 0 0 0 x2.x4[1].delay_signal
flabel metal4 14756 7975 15428 8043 0 FreeSans 320 0 0 0 x2.x4[1].VSS
flabel via3 14860 9139 14924 9203 0 FreeSans 320 0 0 0 x2.x4[1].floating
flabel metal1 15090 9484 15124 9518 0 FreeSans 320 0 0 0 x2.x5[4].SW
flabel nwell 15010 10546 15680 10614 0 FreeSans 320 0 0 0 x2.x5[4].VDD
flabel pdiff 15034 9353 15092 9437 0 FreeSans 320 0 0 0 x2.x5[4].delay_signal
flabel metal4 15579 10545 15680 10614 0 FreeSans 320 0 0 0 x2.x5[4].VDD
flabel via3 15515 9387 15579 9451 0 FreeSans 320 0 0 0 x2.x5[4].floating
flabel viali 15439 9080 15473 9114 0 FreeSans 320 0 0 0 x2.x4[0].SW
flabel ndiff 15383 9152 15441 9236 0 FreeSans 320 0 0 0 x2.x4[0].delay_signal
flabel metal4 15362 7975 16034 8043 0 FreeSans 320 0 0 0 x2.x4[0].VSS
flabel via3 15866 9139 15930 9203 0 FreeSans 320 0 0 0 x2.x4[0].floating
flabel metal1 16176 9484 16210 9518 0 FreeSans 320 0 0 0 x2.x5[3].SW
flabel nwell 15620 10546 16290 10614 0 FreeSans 320 0 0 0 x2.x5[3].VDD
flabel pdiff 16208 9353 16266 9437 0 FreeSans 320 0 0 0 x2.x5[3].delay_signal
flabel metal4 15620 10545 15721 10614 0 FreeSans 320 0 0 0 x2.x5[3].VDD
flabel via3 15721 9387 15785 9451 0 FreeSans 320 0 0 0 x2.x5[3].floating
flabel viali 16655 9080 16689 9114 0 FreeSans 320 0 0 0 x2.x3[1].SW
flabel ndiff 16687 9152 16745 9236 0 FreeSans 320 0 0 0 x2.x3[1].delay_signal
flabel metal4 16094 7975 16766 8043 0 FreeSans 320 0 0 0 x2.x3[1].VSS
flabel via3 16198 9139 16262 9203 0 FreeSans 320 0 0 0 x2.x3[1].floating
flabel metal1 16302 9484 16336 9518 0 FreeSans 320 0 0 0 x2.x5[2].SW
flabel nwell 16222 10546 16892 10614 0 FreeSans 320 0 0 0 x2.x5[2].VDD
flabel pdiff 16246 9353 16304 9437 0 FreeSans 320 0 0 0 x2.x5[2].delay_signal
flabel metal4 16791 10545 16892 10614 0 FreeSans 320 0 0 0 x2.x5[2].VDD
flabel via3 16727 9387 16791 9451 0 FreeSans 320 0 0 0 x2.x5[2].floating
flabel viali 16777 9080 16811 9114 0 FreeSans 320 0 0 0 x2.x3[0].SW
flabel ndiff 16721 9152 16779 9236 0 FreeSans 320 0 0 0 x2.x3[0].delay_signal
flabel metal4 16700 7975 17372 8043 0 FreeSans 320 0 0 0 x2.x3[0].VSS
flabel via3 17204 9139 17268 9203 0 FreeSans 320 0 0 0 x2.x3[0].floating
flabel metal1 17388 9484 17422 9518 0 FreeSans 320 0 0 0 x2.x5[1].SW
flabel nwell 16832 10546 17502 10614 0 FreeSans 320 0 0 0 x2.x5[1].VDD
flabel pdiff 17420 9353 17478 9437 0 FreeSans 320 0 0 0 x2.x5[1].delay_signal
flabel metal4 16832 10545 16933 10614 0 FreeSans 320 0 0 0 x2.x5[1].VDD
flabel via3 16933 9387 16997 9451 0 FreeSans 320 0 0 0 x2.x5[1].floating
flabel viali 17511 9080 17545 9114 0 FreeSans 320 0 0 0 x2.x2.SW
flabel ndiff 17455 9152 17513 9236 0 FreeSans 320 0 0 0 x2.x2.delay_signal
flabel metal4 17434 7975 18106 8043 0 FreeSans 320 0 0 0 x2.x2.VSS
flabel via3 17938 9139 18002 9203 0 FreeSans 320 0 0 0 x2.x2.floating
flabel metal1 17514 9484 17548 9518 0 FreeSans 320 0 0 0 x2.x5[0].SW
flabel nwell 17434 10546 18104 10614 0 FreeSans 320 0 0 0 x2.x5[0].VDD
flabel pdiff 17458 9353 17516 9437 0 FreeSans 320 0 0 0 x2.x5[0].delay_signal
flabel metal4 18003 10545 18104 10614 0 FreeSans 320 0 0 0 x2.x5[0].VDD
flabel via3 17939 9387 18003 9451 0 FreeSans 320 0 0 0 x2.x5[0].floating
flabel metal1 18501 9585 18535 9619 0 FreeSans 200 0 0 0 x3.VPWR
flabel metal1 18501 9041 18535 9075 0 FreeSans 200 0 0 0 x3.VGND
flabel locali 18501 9585 18535 9619 0 FreeSans 200 0 0 0 x3.VPWR
flabel locali 18501 9041 18535 9075 0 FreeSans 200 0 0 0 x3.VGND
flabel locali 18684 9143 18718 9177 0 FreeSans 200 0 0 0 x3.X
flabel locali 18684 9415 18718 9449 0 FreeSans 200 0 0 0 x3.X
flabel locali 18684 9483 18718 9517 0 FreeSans 200 0 0 0 x3.X
flabel locali 18501 9279 18535 9313 0 FreeSans 200 0 0 0 x3.A
flabel nwell 18501 9585 18535 9619 0 FreeSans 200 0 0 0 x3.VPB
flabel pwell 18501 9041 18535 9075 0 FreeSans 200 0 0 0 x3.VNB
rlabel comment 18472 9058 18472 9058 4 x3.buf_2
rlabel metal1 18472 9010 18840 9106 1 x3.VGND
rlabel metal1 18472 9554 18840 9650 1 x3.VPWR
<< end >>
