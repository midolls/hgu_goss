magic
tech sky130A
magscale 1 2
timestamp 1698804095
<< error_p >>
rect -15 54 15 68
rect -239 -48 -237 12
rect -207 -48 -205 12
rect -15 -68 15 -58
<< nmos >>
rect -15 -42 15 42
<< ndiff >>
rect -73 30 -15 42
rect -245 12 -199 24
rect -245 -48 -239 12
rect -205 -48 -199 12
rect -73 -30 -61 30
rect -27 -30 -15 30
rect -73 -42 -15 -30
rect 15 30 73 42
rect 15 -30 27 30
rect 61 -30 73 30
rect 15 -42 73 -30
rect -245 -60 -199 -48
<< ndiffc >>
rect -239 -48 -205 12
rect -61 -30 -27 30
rect 27 -30 61 30
<< poly >>
rect -15 42 15 54
rect -15 -58 15 -42
<< locali >>
rect -61 30 -27 46
rect -239 12 -205 28
rect -61 -46 -27 -30
rect 27 30 61 46
rect 27 -46 61 -30
rect -239 -64 -205 -48
<< viali >>
rect -239 -48 -205 12
rect -61 -30 -27 30
rect 27 -30 61 30
<< metal1 >>
rect -67 30 -21 42
rect -245 12 -199 24
rect -245 -48 -239 12
rect -205 -48 -199 12
rect -67 -30 -61 30
rect -27 -30 -21 30
rect -67 -42 -21 -30
rect 21 30 67 42
rect 21 -30 27 30
rect 61 -30 67 30
rect 21 -42 67 -30
rect -245 -60 -199 -48
<< properties >>
string FIXED_BBOX -158 -199 158 199
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.420 l 0.150 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
