magic
tech sky130A
magscale 1 2
timestamp 1696942209
<< error_p >>
rect -29 156 29 162
rect -29 122 -17 156
rect -29 116 29 122
rect -29 -122 29 -116
rect -29 -156 -17 -122
rect -29 -162 29 -156
<< pwell >>
rect -211 -294 211 294
<< nmos >>
rect -15 -84 15 84
<< ndiff >>
rect -73 72 -15 84
rect -73 -72 -61 72
rect -27 -72 -15 72
rect -73 -84 -15 -72
rect 15 72 73 84
rect 15 -72 27 72
rect 61 -72 73 72
rect 15 -84 73 -72
<< ndiffc >>
rect -61 -72 -27 72
rect 27 -72 61 72
<< psubdiff >>
rect -175 224 -79 258
rect 79 224 175 258
rect -175 162 -141 224
rect 141 162 175 224
rect -175 -224 -141 -162
rect 141 -224 175 -162
rect -175 -258 -79 -224
rect 79 -258 175 -224
<< psubdiffcont >>
rect -79 224 79 258
rect -175 -162 -141 162
rect 141 -162 175 162
rect -79 -258 79 -224
<< poly >>
rect -33 156 33 172
rect -33 122 -17 156
rect 17 122 33 156
rect -33 106 33 122
rect -15 84 15 106
rect -15 -106 15 -84
rect -33 -122 33 -106
rect -33 -156 -17 -122
rect 17 -156 33 -122
rect -33 -172 33 -156
<< polycont >>
rect -17 122 17 156
rect -17 -156 17 -122
<< locali >>
rect -175 224 -79 258
rect 79 224 175 258
rect -175 162 -141 224
rect 141 162 175 224
rect -33 122 -17 156
rect 17 122 33 156
rect -61 72 -27 88
rect -61 -88 -27 -72
rect 27 72 61 88
rect 27 -88 61 -72
rect -33 -156 -17 -122
rect 17 -156 33 -122
rect -175 -224 -141 -162
rect 141 -224 175 -162
rect -175 -258 -79 -224
rect 79 -258 175 -224
<< viali >>
rect -17 122 17 156
rect -61 -72 -27 72
rect 27 -72 61 72
rect -17 -156 17 -122
<< metal1 >>
rect -29 156 29 162
rect -29 122 -17 156
rect 17 122 29 156
rect -29 116 29 122
rect -67 72 -21 84
rect -67 -72 -61 72
rect -27 -72 -21 72
rect -67 -84 -21 -72
rect 21 72 67 84
rect 21 -72 27 72
rect 61 -72 67 72
rect 21 -84 67 -72
rect -29 -122 29 -116
rect -29 -156 -17 -122
rect 17 -156 29 -122
rect -29 -162 29 -156
<< properties >>
string FIXED_BBOX -158 -241 158 241
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.84 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
