magic
tech sky130A
magscale 1 2
timestamp 1699326276
<< nwell >>
rect 9791 2389 15997 2986
rect 9742 2388 15997 2389
rect 9262 2322 15997 2388
rect 9262 2300 9760 2322
rect 9264 2298 9760 2300
rect 9453 2146 9501 2202
rect 9791 1692 15997 2322
<< ndiff >>
rect 11664 1549 11722 1561
rect 11664 1489 11676 1549
rect 11710 1489 11722 1549
rect 11664 1477 11722 1489
rect 12875 1549 12933 1561
rect 12875 1489 12887 1549
rect 12921 1489 12933 1549
rect 12875 1477 12933 1489
rect 14215 1549 14273 1561
rect 14215 1489 14227 1549
rect 14261 1489 14273 1549
rect 14215 1477 14273 1489
rect 14962 1549 15020 1561
rect 14962 1489 14974 1549
rect 15008 1489 15020 1549
rect 14962 1477 15020 1489
<< pdiff >>
rect 9453 2146 9501 2202
rect 11309 1750 11367 1762
rect 11309 1690 11321 1750
rect 11355 1690 11367 1750
rect 11309 1678 11367 1690
rect 12520 1750 12578 1762
rect 12520 1690 12532 1750
rect 12566 1690 12578 1750
rect 12520 1678 12578 1690
rect 13733 1750 13791 1762
rect 13733 1690 13745 1750
rect 13779 1690 13791 1750
rect 13733 1678 13791 1690
rect 14947 1750 15005 1762
rect 14947 1690 14959 1750
rect 14993 1690 15005 1750
rect 14947 1678 15005 1690
<< ndiffc >>
rect 10927 1489 10961 1549
rect 11676 1489 11710 1549
rect 12887 1489 12921 1549
rect 14227 1489 14261 1549
rect 14974 1489 15008 1549
<< pdiffc >>
rect 10572 1690 10606 1750
rect 11321 1690 11355 1750
rect 12532 1690 12566 1750
rect 13745 1690 13779 1750
rect 14959 1690 14993 1750
<< psubdiff >>
rect 9370 1714 9394 1748
rect 9428 1714 9512 1748
rect 9546 1714 9656 1748
rect 9690 1714 9732 1748
rect 9370 1712 9732 1714
<< nsubdiff >>
rect 15776 2868 15862 2894
rect 15776 2834 15802 2868
rect 15836 2834 15862 2868
rect 15776 2808 15862 2834
rect 15781 2724 15867 2750
rect 15781 2690 15807 2724
rect 15841 2690 15867 2724
rect 15781 2664 15867 2690
rect 15782 2572 15868 2598
rect 15782 2538 15808 2572
rect 15842 2538 15868 2572
rect 15782 2512 15868 2538
rect 15782 2402 15868 2428
rect 15782 2368 15808 2402
rect 15842 2368 15868 2402
rect 9344 2350 9760 2352
rect 9344 2316 9374 2350
rect 9408 2316 9504 2350
rect 9538 2316 9650 2350
rect 9684 2316 9760 2350
rect 15782 2342 15868 2368
rect 9344 2312 9760 2316
rect 15781 2245 15867 2271
rect 15781 2211 15807 2245
rect 15841 2211 15867 2245
rect 15781 2185 15867 2211
<< psubdiffcont >>
rect 9394 1714 9428 1748
rect 9512 1714 9546 1748
rect 9656 1714 9690 1748
<< nsubdiffcont >>
rect 15802 2834 15836 2868
rect 15807 2690 15841 2724
rect 15808 2538 15842 2572
rect 15808 2368 15842 2402
rect 9374 2316 9408 2350
rect 9504 2316 9538 2350
rect 9650 2316 9684 2350
rect 15807 2211 15841 2245
<< poly >>
rect 15544 1636 15703 1656
rect 15544 1602 15556 1636
rect 15590 1602 15703 1636
rect 15544 1583 15703 1602
rect 15765 1577 15891 1656
rect 9881 1449 9947 1465
rect 9881 1422 9897 1449
rect 9863 1415 9897 1422
rect 9931 1422 9947 1449
rect 9931 1415 9965 1422
rect 9863 1392 9965 1415
<< polycont >>
rect 15556 1602 15590 1636
rect 9897 1415 9931 1449
<< locali >>
rect 9938 2868 10053 2908
rect 15776 2868 15862 2894
rect 15776 2834 15802 2868
rect 15836 2834 15862 2868
rect 15776 2808 15862 2834
rect 15781 2724 15867 2750
rect 15781 2690 15807 2724
rect 15841 2690 15867 2724
rect 15781 2664 15867 2690
rect 15782 2572 15868 2598
rect 15782 2538 15808 2572
rect 15842 2538 15868 2572
rect 15782 2512 15868 2538
rect 15782 2402 15868 2428
rect 15782 2368 15808 2402
rect 15842 2368 15868 2402
rect 9358 2316 9374 2350
rect 9408 2316 9424 2350
rect 9488 2316 9504 2350
rect 9538 2316 9558 2350
rect 9634 2318 9650 2350
rect 9684 2318 9704 2350
rect 15782 2342 15868 2368
rect 15781 2245 15867 2271
rect 15781 2211 15807 2245
rect 15841 2211 15867 2245
rect 9453 2178 9501 2202
rect 15781 2185 15867 2211
rect 9453 2146 9457 2178
rect 9491 2146 9501 2178
rect 9647 2012 9681 2021
rect 9780 2013 9829 2025
rect 9647 1987 9650 2012
rect 9780 1979 9789 2013
rect 9823 2008 9829 2013
rect 9823 1979 10112 2008
rect 9780 1973 10112 1979
rect 9780 1966 9829 1973
rect 10077 1950 10112 1973
rect 10077 1938 10126 1950
rect 9818 1920 9867 1932
rect 9818 1886 9827 1920
rect 9861 1886 10028 1920
rect 10077 1904 10086 1938
rect 10120 1904 10126 1938
rect 10077 1891 10126 1904
rect 9818 1873 9867 1886
rect 9987 1844 10028 1886
rect 10078 1845 10127 1857
rect 10078 1844 10087 1845
rect 9987 1811 10087 1844
rect 10121 1811 10127 1845
rect 9987 1810 10127 1811
rect 10078 1798 10127 1810
rect 9378 1748 9454 1756
rect 9378 1714 9394 1748
rect 9428 1714 9454 1748
rect 9496 1748 9572 1756
rect 10572 1750 10606 1766
rect 9496 1714 9512 1748
rect 9546 1714 9572 1748
rect 9638 1714 9656 1744
rect 9690 1714 9706 1744
rect 10572 1674 10606 1690
rect 11321 1750 11355 1766
rect 11321 1674 11355 1690
rect 12532 1750 12566 1766
rect 12532 1674 12566 1690
rect 13745 1750 13779 1766
rect 13745 1674 13779 1690
rect 14959 1750 14993 1766
rect 14959 1674 14993 1690
rect 15540 1602 15556 1636
rect 15590 1602 15606 1636
rect 10927 1549 10961 1565
rect 10927 1473 10961 1489
rect 11676 1549 11710 1565
rect 11676 1473 11710 1489
rect 12887 1549 12921 1565
rect 12887 1473 12921 1489
rect 14227 1549 14261 1565
rect 14227 1473 14261 1489
rect 14974 1549 15008 1565
rect 14974 1473 15008 1489
rect 9881 1415 9897 1449
rect 9931 1415 9947 1449
<< viali >>
rect 15802 2834 15836 2868
rect 15807 2690 15841 2724
rect 15808 2538 15842 2572
rect 15808 2368 15842 2402
rect 15807 2211 15841 2245
rect 9457 2144 9491 2178
rect 9566 2089 9600 2123
rect 9376 1979 9410 2013
rect 9650 1978 9684 2012
rect 9789 1979 9823 2013
rect 9827 1886 9861 1920
rect 10086 1904 10120 1938
rect 10087 1811 10121 1845
rect 10572 1690 10606 1750
rect 11321 1690 11355 1750
rect 12532 1690 12566 1750
rect 13745 1690 13779 1750
rect 14959 1690 14993 1750
rect 15556 1602 15590 1636
rect 10927 1489 10961 1549
rect 11676 1489 11710 1549
rect 12887 1489 12921 1549
rect 14227 1489 14261 1549
rect 14974 1489 15008 1549
rect 9897 1415 9931 1449
<< metal1 >>
rect 9963 2937 10053 2953
rect 9963 2926 9982 2937
rect 9945 2885 9982 2926
rect 10034 2885 10053 2937
rect 9945 2870 10053 2885
rect 15772 2875 15862 2891
rect 9945 2838 9998 2870
rect 15772 2823 15791 2875
rect 15843 2823 15862 2875
rect 15772 2807 15862 2823
rect 15777 2731 15867 2747
rect 15777 2679 15796 2731
rect 15848 2679 15867 2731
rect 15777 2663 15867 2679
rect 15778 2579 15868 2595
rect 15778 2527 15797 2579
rect 15849 2527 15868 2579
rect 15778 2511 15868 2527
rect 15778 2409 15868 2425
rect 15778 2357 15797 2409
rect 15849 2357 15868 2409
rect 9358 2332 9424 2350
rect 9358 2316 9365 2332
rect 9363 2280 9365 2316
rect 9417 2316 9424 2332
rect 9494 2331 9550 2342
rect 9417 2280 9419 2316
rect 9363 2269 9419 2280
rect 9494 2279 9496 2331
rect 9548 2279 9550 2331
rect 9634 2332 9704 2350
rect 15778 2341 15868 2357
rect 9634 2318 9640 2332
rect 9494 2268 9550 2279
rect 9638 2280 9640 2318
rect 9692 2318 9704 2332
rect 9692 2280 9694 2318
rect 9638 2269 9694 2280
rect 15777 2252 15867 2268
rect 9445 2178 9808 2185
rect 9445 2144 9457 2178
rect 9491 2157 9808 2178
rect 9491 2144 9503 2157
rect 9445 2137 9503 2144
rect 9550 2123 9617 2129
rect 9550 2089 9566 2123
rect 9600 2110 9617 2123
rect 9600 2089 9752 2110
rect 9550 2082 9752 2089
rect 9630 2021 9696 2023
rect 9368 2016 9422 2020
rect 9367 2013 9422 2016
rect 9238 1979 9376 2013
rect 9410 1979 9422 2013
rect 9367 1976 9422 1979
rect 9367 1972 9421 1976
rect 9630 1969 9638 2021
rect 9690 1969 9696 2021
rect 9630 1968 9696 1969
rect 9724 1938 9752 2082
rect 9780 2025 9808 2157
rect 9956 2130 10027 2214
rect 15777 2200 15796 2252
rect 15848 2200 15867 2252
rect 15777 2184 15867 2200
rect 9780 2013 9829 2025
rect 9780 1979 9789 2013
rect 9823 1979 9829 2013
rect 9780 1966 9829 1979
rect 9724 1920 9867 1938
rect 9724 1910 9827 1920
rect 9818 1886 9827 1910
rect 9861 1886 9867 1920
rect 9818 1873 9867 1886
rect 9381 1786 9437 1797
rect 9381 1756 9383 1786
rect 9378 1734 9383 1756
rect 9435 1756 9437 1786
rect 9501 1786 9557 1797
rect 9501 1756 9503 1786
rect 9435 1734 9454 1756
rect 9378 1714 9454 1734
rect 9496 1734 9503 1756
rect 9555 1756 9557 1786
rect 9644 1786 9700 1797
rect 9555 1734 9572 1756
rect 9644 1744 9646 1786
rect 9496 1714 9572 1734
rect 9638 1734 9646 1744
rect 9698 1744 9700 1786
rect 9698 1734 9706 1744
rect 9638 1714 9706 1734
rect 9895 1643 9943 2089
rect 9275 1596 9943 1643
rect 9895 1455 9943 1596
rect 9885 1449 9943 1455
rect 9644 1443 9709 1444
rect 9644 1442 9650 1443
rect 9548 1440 9650 1442
rect 9546 1394 9650 1440
rect 9644 1391 9650 1394
rect 9702 1391 9709 1443
rect 9885 1415 9897 1449
rect 9931 1415 9943 1449
rect 9885 1409 9943 1415
rect 9981 1640 10027 2130
rect 15695 2010 15785 2026
rect 15695 1999 15714 2010
rect 15620 1958 15714 1999
rect 15766 1958 15785 2010
rect 10077 1943 10126 1950
rect 10077 1938 10696 1943
rect 10077 1904 10086 1938
rect 10120 1904 10696 1938
rect 10077 1896 10696 1904
rect 10077 1891 10126 1896
rect 10078 1849 10127 1857
rect 10647 1849 10696 1896
rect 15620 1940 15785 1958
rect 15620 1894 15667 1940
rect 10078 1845 10579 1849
rect 10078 1811 10087 1845
rect 10121 1811 10579 1845
rect 10078 1803 10579 1811
rect 10647 1803 15068 1849
rect 10078 1802 10567 1803
rect 10647 1802 11093 1803
rect 10078 1798 10127 1802
rect 15709 1793 15947 1822
rect 10566 1750 10612 1762
rect 10566 1690 10572 1750
rect 10606 1690 10612 1750
rect 10566 1640 10612 1690
rect 11315 1750 11361 1762
rect 11315 1690 11321 1750
rect 11355 1690 11361 1750
rect 11315 1640 11361 1690
rect 12526 1750 12572 1762
rect 12526 1690 12532 1750
rect 12566 1690 12572 1750
rect 12526 1640 12572 1690
rect 13739 1750 13785 1762
rect 13739 1690 13745 1750
rect 13779 1690 13785 1750
rect 13739 1640 13785 1690
rect 14953 1750 14999 1762
rect 15709 1756 15755 1793
rect 14953 1690 14959 1750
rect 14993 1690 14999 1750
rect 14953 1640 14999 1690
rect 15783 1749 15873 1765
rect 15901 1764 15947 1793
rect 15783 1697 15802 1749
rect 15854 1697 15873 1749
rect 15540 1640 15606 1642
rect 9981 1636 15606 1640
rect 9981 1602 15556 1636
rect 15590 1602 15606 1636
rect 9981 1598 15606 1602
rect 9981 1368 10027 1598
rect 10921 1549 10967 1598
rect 10921 1489 10927 1549
rect 10961 1489 10967 1549
rect 10921 1477 10967 1489
rect 11670 1549 11716 1598
rect 11670 1489 11676 1549
rect 11710 1489 11716 1549
rect 11670 1477 11716 1489
rect 12881 1549 12927 1598
rect 12881 1489 12887 1549
rect 12921 1489 12927 1549
rect 12881 1477 12927 1489
rect 14221 1549 14267 1598
rect 14221 1489 14227 1549
rect 14261 1489 14267 1549
rect 14221 1477 14267 1489
rect 14968 1549 15014 1598
rect 15544 1596 15606 1598
rect 15639 1633 15667 1683
rect 15783 1681 15873 1697
rect 15751 1633 15933 1640
rect 15639 1604 15933 1633
rect 15639 1556 15667 1604
rect 15751 1594 15933 1604
rect 14968 1489 14974 1549
rect 15008 1489 15014 1549
rect 14968 1477 15014 1489
rect 15783 1546 15873 1562
rect 15783 1494 15802 1546
rect 15854 1494 15873 1546
rect 15709 1450 15755 1480
rect 15783 1478 15873 1494
rect 15901 1450 15947 1481
rect 10131 1391 10138 1443
rect 10190 1441 10196 1443
rect 10190 1424 10913 1441
rect 10190 1394 10929 1424
rect 11603 1399 12997 1445
rect 14153 1399 14335 1445
rect 10190 1391 10196 1394
rect 10131 1390 10196 1391
rect 10871 1389 10929 1394
rect 10013 1293 10027 1368
rect 9932 359 10039 375
rect 9932 307 9968 359
rect 10020 307 10039 359
rect 9932 291 10039 307
rect 11727 268 11785 1399
rect 14153 268 14211 1399
rect 15009 267 15068 1448
rect 15709 1421 15947 1450
rect 15621 1300 15667 1344
rect 15621 1284 15782 1300
rect 15621 1232 15711 1284
rect 15763 1232 15782 1284
rect 15621 1216 15782 1232
<< via1 >>
rect 9982 2885 10034 2937
rect 15791 2868 15843 2875
rect 15791 2834 15802 2868
rect 15802 2834 15836 2868
rect 15836 2834 15843 2868
rect 15791 2823 15843 2834
rect 15796 2724 15848 2731
rect 15796 2690 15807 2724
rect 15807 2690 15841 2724
rect 15841 2690 15848 2724
rect 15796 2679 15848 2690
rect 15797 2572 15849 2579
rect 15797 2538 15808 2572
rect 15808 2538 15842 2572
rect 15842 2538 15849 2572
rect 15797 2527 15849 2538
rect 15797 2402 15849 2409
rect 15797 2368 15808 2402
rect 15808 2368 15842 2402
rect 15842 2368 15849 2402
rect 15797 2357 15849 2368
rect 9365 2280 9417 2332
rect 9496 2279 9548 2331
rect 9640 2280 9692 2332
rect 9638 2012 9690 2021
rect 9638 1978 9650 2012
rect 9650 1978 9684 2012
rect 9684 1978 9690 2012
rect 9638 1969 9690 1978
rect 15796 2245 15848 2252
rect 15796 2211 15807 2245
rect 15807 2211 15841 2245
rect 15841 2211 15848 2245
rect 15796 2200 15848 2211
rect 9383 1734 9435 1786
rect 9503 1734 9555 1786
rect 9646 1734 9698 1786
rect 9650 1391 9702 1443
rect 15714 1958 15766 2010
rect 15802 1697 15854 1749
rect 15802 1494 15854 1546
rect 10138 1391 10190 1443
rect 9968 307 10020 359
rect 15711 1232 15763 1284
<< metal2 >>
rect 9971 2939 10045 2943
rect 9971 2883 9980 2939
rect 10036 2883 10045 2939
rect 9971 2879 10045 2883
rect 15780 2877 15854 2881
rect 15780 2821 15789 2877
rect 15845 2821 15854 2877
rect 15780 2817 15854 2821
rect 15785 2733 15859 2737
rect 15785 2677 15794 2733
rect 15850 2677 15859 2733
rect 15785 2673 15859 2677
rect 15786 2581 15860 2585
rect 15786 2525 15795 2581
rect 15851 2525 15860 2581
rect 15786 2521 15860 2525
rect 15786 2411 15860 2415
rect 15786 2355 15795 2411
rect 15851 2355 15860 2411
rect 15786 2351 15860 2355
rect 9363 2334 9419 2343
rect 9363 2269 9419 2278
rect 9494 2333 9550 2342
rect 9494 2268 9550 2277
rect 9638 2334 9694 2343
rect 9638 2269 9694 2278
rect 15785 2254 15859 2258
rect 15785 2198 15794 2254
rect 15850 2198 15859 2254
rect 15785 2194 15859 2198
rect 9630 1969 9638 2021
rect 9690 1969 9696 2021
rect 9630 1968 9696 1969
rect 15703 2012 15777 2016
rect 9648 1892 9694 1968
rect 15703 1956 15712 2012
rect 15768 1956 15777 2012
rect 15703 1952 15777 1956
rect 9648 1846 9887 1892
rect 9381 1788 9437 1797
rect 9381 1723 9437 1732
rect 9501 1788 9557 1797
rect 9501 1723 9557 1732
rect 9644 1788 9700 1797
rect 9644 1723 9700 1732
rect 9644 1443 9709 1444
rect 9644 1391 9650 1443
rect 9702 1440 9709 1443
rect 9841 1440 9887 1846
rect 15791 1751 15865 1755
rect 15791 1695 15800 1751
rect 15856 1695 15865 1751
rect 15791 1691 15865 1695
rect 15791 1548 15865 1552
rect 15791 1492 15800 1548
rect 15856 1492 15865 1548
rect 15791 1488 15865 1492
rect 10131 1440 10138 1443
rect 9702 1394 10138 1440
rect 9702 1391 9709 1394
rect 10131 1391 10138 1394
rect 10190 1391 10196 1443
rect 10131 1390 10196 1391
rect 15700 1286 15774 1290
rect 15700 1230 15709 1286
rect 15765 1230 15774 1286
rect 15700 1226 15774 1230
rect 9957 361 10031 365
rect 9957 305 9966 361
rect 10022 305 10031 361
rect 9957 301 10031 305
<< via2 >>
rect 9980 2937 10036 2939
rect 9980 2885 9982 2937
rect 9982 2885 10034 2937
rect 10034 2885 10036 2937
rect 9980 2883 10036 2885
rect 15789 2875 15845 2877
rect 15789 2823 15791 2875
rect 15791 2823 15843 2875
rect 15843 2823 15845 2875
rect 15789 2821 15845 2823
rect 15794 2731 15850 2733
rect 15794 2679 15796 2731
rect 15796 2679 15848 2731
rect 15848 2679 15850 2731
rect 15794 2677 15850 2679
rect 15795 2579 15851 2581
rect 15795 2527 15797 2579
rect 15797 2527 15849 2579
rect 15849 2527 15851 2579
rect 15795 2525 15851 2527
rect 15795 2409 15851 2411
rect 15795 2357 15797 2409
rect 15797 2357 15849 2409
rect 15849 2357 15851 2409
rect 15795 2355 15851 2357
rect 9363 2332 9419 2334
rect 9363 2280 9365 2332
rect 9365 2280 9417 2332
rect 9417 2280 9419 2332
rect 9363 2278 9419 2280
rect 9494 2331 9550 2333
rect 9494 2279 9496 2331
rect 9496 2279 9548 2331
rect 9548 2279 9550 2331
rect 9494 2277 9550 2279
rect 9638 2332 9694 2334
rect 9638 2280 9640 2332
rect 9640 2280 9692 2332
rect 9692 2280 9694 2332
rect 9638 2278 9694 2280
rect 15794 2252 15850 2254
rect 15794 2200 15796 2252
rect 15796 2200 15848 2252
rect 15848 2200 15850 2252
rect 15794 2198 15850 2200
rect 15712 2010 15768 2012
rect 15712 1958 15714 2010
rect 15714 1958 15766 2010
rect 15766 1958 15768 2010
rect 15712 1956 15768 1958
rect 9381 1786 9437 1788
rect 9381 1734 9383 1786
rect 9383 1734 9435 1786
rect 9435 1734 9437 1786
rect 9381 1732 9437 1734
rect 9501 1786 9557 1788
rect 9501 1734 9503 1786
rect 9503 1734 9555 1786
rect 9555 1734 9557 1786
rect 9501 1732 9557 1734
rect 9644 1786 9700 1788
rect 9644 1734 9646 1786
rect 9646 1734 9698 1786
rect 9698 1734 9700 1786
rect 9644 1732 9700 1734
rect 15800 1749 15856 1751
rect 15800 1697 15802 1749
rect 15802 1697 15854 1749
rect 15854 1697 15856 1749
rect 15800 1695 15856 1697
rect 15800 1546 15856 1548
rect 15800 1494 15802 1546
rect 15802 1494 15854 1546
rect 15854 1494 15856 1546
rect 15800 1492 15856 1494
rect 15709 1284 15765 1286
rect 15709 1232 15711 1284
rect 15711 1232 15763 1284
rect 15763 1232 15765 1284
rect 15709 1230 15765 1232
rect 9966 359 10022 361
rect 9966 307 9968 359
rect 9968 307 10020 359
rect 10020 307 10022 359
rect 9966 305 10022 307
<< metal3 >>
rect 9945 2943 10071 2953
rect 9945 2879 9976 2943
rect 10040 2879 10071 2943
rect 9945 2870 10071 2879
rect 15754 2881 15880 2891
rect 15754 2817 15785 2881
rect 15849 2817 15880 2881
rect 15754 2807 15880 2817
rect 15759 2737 15885 2747
rect 15759 2673 15790 2737
rect 15854 2673 15885 2737
rect 15759 2663 15885 2673
rect 15760 2585 15886 2595
rect 15760 2521 15791 2585
rect 15855 2521 15886 2585
rect 15760 2511 15886 2521
rect 15760 2415 15886 2425
rect 9344 2352 9462 2353
rect 9593 2352 9737 2353
rect 9344 2338 9737 2352
rect 15760 2351 15791 2415
rect 15855 2351 15886 2415
rect 15760 2341 15886 2351
rect 9344 2274 9359 2338
rect 9423 2337 9634 2338
rect 9423 2274 9490 2337
rect 9344 2273 9490 2274
rect 9554 2274 9634 2337
rect 9698 2274 9737 2338
rect 9554 2273 9737 2274
rect 9344 2257 9737 2273
rect 15759 2258 15885 2268
rect 9449 2256 9593 2257
rect 15759 2194 15790 2258
rect 15854 2194 15885 2258
rect 15759 2184 15885 2194
rect 15677 2016 15803 2026
rect 15677 1952 15708 2016
rect 15772 1952 15803 2016
rect 15677 1942 15803 1952
rect 9484 1807 9576 1808
rect 9370 1792 9743 1807
rect 9370 1728 9377 1792
rect 9441 1728 9497 1792
rect 9561 1728 9640 1792
rect 9704 1728 9743 1792
rect 9370 1711 9743 1728
rect 15765 1755 15891 1765
rect 15765 1691 15796 1755
rect 15860 1691 15891 1755
rect 15765 1681 15891 1691
rect 15765 1552 15891 1562
rect 15765 1488 15796 1552
rect 15860 1488 15891 1552
rect 15765 1478 15891 1488
rect 15791 1477 15865 1478
rect 15675 1290 15800 1300
rect 15675 1226 15705 1290
rect 15769 1226 15800 1290
rect 15675 1216 15800 1226
rect 9932 365 10057 375
rect 9932 301 9962 365
rect 10026 301 10057 365
rect 9932 291 10057 301
<< via3 >>
rect 9976 2939 10040 2943
rect 9976 2883 9980 2939
rect 9980 2883 10036 2939
rect 10036 2883 10040 2939
rect 9976 2879 10040 2883
rect 15785 2877 15849 2881
rect 15785 2821 15789 2877
rect 15789 2821 15845 2877
rect 15845 2821 15849 2877
rect 15785 2817 15849 2821
rect 15790 2733 15854 2737
rect 15790 2677 15794 2733
rect 15794 2677 15850 2733
rect 15850 2677 15854 2733
rect 15790 2673 15854 2677
rect 15791 2581 15855 2585
rect 15791 2525 15795 2581
rect 15795 2525 15851 2581
rect 15851 2525 15855 2581
rect 15791 2521 15855 2525
rect 15791 2411 15855 2415
rect 15791 2355 15795 2411
rect 15795 2355 15851 2411
rect 15851 2355 15855 2411
rect 15791 2351 15855 2355
rect 9359 2334 9423 2338
rect 9359 2278 9363 2334
rect 9363 2278 9419 2334
rect 9419 2278 9423 2334
rect 9359 2274 9423 2278
rect 9490 2333 9554 2337
rect 9490 2277 9494 2333
rect 9494 2277 9550 2333
rect 9550 2277 9554 2333
rect 9490 2273 9554 2277
rect 9634 2334 9698 2338
rect 9634 2278 9638 2334
rect 9638 2278 9694 2334
rect 9694 2278 9698 2334
rect 9634 2274 9698 2278
rect 15790 2254 15854 2258
rect 15790 2198 15794 2254
rect 15794 2198 15850 2254
rect 15850 2198 15854 2254
rect 15790 2194 15854 2198
rect 15708 2012 15772 2016
rect 15708 1956 15712 2012
rect 15712 1956 15768 2012
rect 15768 1956 15772 2012
rect 15708 1952 15772 1956
rect 9377 1788 9441 1792
rect 9377 1732 9381 1788
rect 9381 1732 9437 1788
rect 9437 1732 9441 1788
rect 9377 1728 9441 1732
rect 9497 1788 9561 1792
rect 9497 1732 9501 1788
rect 9501 1732 9557 1788
rect 9557 1732 9561 1788
rect 9497 1728 9561 1732
rect 9640 1788 9704 1792
rect 9640 1732 9644 1788
rect 9644 1732 9700 1788
rect 9700 1732 9704 1788
rect 9640 1728 9704 1732
rect 15796 1751 15860 1755
rect 15796 1695 15800 1751
rect 15800 1695 15856 1751
rect 15856 1695 15860 1751
rect 15796 1691 15860 1695
rect 15796 1548 15860 1552
rect 15796 1492 15800 1548
rect 15800 1492 15856 1548
rect 15856 1492 15860 1548
rect 15796 1488 15860 1492
rect 15705 1286 15769 1290
rect 15705 1230 15709 1286
rect 15709 1230 15765 1286
rect 15765 1230 15769 1286
rect 15705 1226 15769 1230
rect 9962 361 10026 365
rect 9962 305 9966 361
rect 9966 305 10022 361
rect 10022 305 10026 361
rect 9962 301 10026 305
<< metal4 >>
rect 9945 2948 10071 2953
rect 9344 2943 15993 2948
rect 9344 2879 9976 2943
rect 10040 2881 15993 2943
rect 10040 2879 15785 2881
rect 9344 2870 15785 2879
rect 9344 2338 9762 2870
rect 9344 2274 9359 2338
rect 9423 2337 9634 2338
rect 9423 2274 9490 2337
rect 9344 2273 9490 2274
rect 9554 2274 9634 2337
rect 9698 2332 9762 2338
rect 15675 2817 15785 2870
rect 15849 2817 15993 2881
rect 15675 2737 15993 2817
rect 15675 2673 15790 2737
rect 15854 2673 15993 2737
rect 15675 2585 15993 2673
rect 15675 2521 15791 2585
rect 15855 2521 15993 2585
rect 15675 2415 15993 2521
rect 15675 2351 15791 2415
rect 15855 2351 15993 2415
rect 9698 2274 9761 2332
rect 9554 2273 9761 2274
rect 9344 2255 9761 2273
rect 15675 2258 15993 2351
rect 15675 2194 15790 2258
rect 15854 2194 15993 2258
rect 15675 2016 15993 2194
rect 15675 1952 15708 2016
rect 15772 1952 15993 2016
rect 15675 1940 15993 1952
rect 9370 1792 9747 1807
rect 9370 1728 9377 1792
rect 9441 1728 9497 1792
rect 9561 1728 9640 1792
rect 9704 1728 9747 1792
rect 15675 1755 15873 1765
rect 9372 369 9748 1728
rect 15675 1691 15796 1755
rect 15860 1691 15873 1755
rect 15675 1681 15873 1691
rect 15675 1300 15735 1681
rect 15933 1562 15993 1940
rect 15795 1552 15993 1562
rect 15795 1488 15796 1552
rect 15860 1488 15993 1552
rect 15795 1478 15993 1488
rect 15675 1290 15993 1300
rect 15675 1226 15705 1290
rect 15769 1226 15993 1290
rect 9932 369 10057 375
rect 15675 369 15993 1226
rect 9372 365 15993 369
rect 9372 301 9962 365
rect 10026 301 15993 365
rect 9372 291 15993 301
use hgu_sw_cap_nmos  x2
timestamp 1699326276
transform -1 0 15982 0 1 -246
box 368 546 1040 1833
use hgu_sw_cap_nmos  x3[0]
timestamp 1699326276
transform -1 0 15248 0 1 -246
box 368 546 1040 1833
use hgu_sw_cap_nmos  x3[1]
timestamp 1699326276
transform 1 0 13234 0 1 -246
box 368 546 1040 1833
use hgu_sw_cap_nmos  x4[0]
timestamp 1699326276
transform -1 0 13910 0 1 -246
box 368 546 1040 1833
use hgu_sw_cap_nmos  x4[1]
timestamp 1699326276
transform 1 0 11896 0 1 -246
box 368 546 1040 1833
use hgu_sw_cap_nmos  x4[2]
timestamp 1699326276
transform -1 0 12698 0 1 -246
box 368 546 1040 1833
use hgu_sw_cap_nmos  x4[3]
timestamp 1699326276
transform 1 0 10684 0 1 -246
box 368 546 1040 1833
use hgu_sw_cap_pmos  x5[0]
timestamp 1699325447
transform -1 0 15984 0 -1 3485
box 369 500 1054 1856
use hgu_sw_cap_pmos  x5[1]
timestamp 1699325447
transform 1 0 13968 0 -1 3485
box 369 500 1054 1856
use hgu_sw_cap_pmos  x5[2]
timestamp 1699325447
transform -1 0 14772 0 -1 3485
box 369 500 1054 1856
use hgu_sw_cap_pmos  x5[3]
timestamp 1699325447
transform 1 0 12756 0 -1 3485
box 369 500 1054 1856
use hgu_sw_cap_pmos  x5[4]
timestamp 1699325447
transform -1 0 13560 0 -1 3485
box 369 500 1054 1856
use hgu_sw_cap_pmos  x5[5]
timestamp 1699325447
transform 1 0 11544 0 -1 3485
box 369 500 1054 1856
use hgu_sw_cap_pmos  x5[6]
timestamp 1699325447
transform -1 0 12348 0 -1 3485
box 369 500 1054 1856
use hgu_sw_cap_pmos  x5[7]
timestamp 1699325447
transform 1 0 10332 0 -1 3485
box 369 500 1054 1856
use hgu_sw_cap_pmos  x6
timestamp 1699325447
transform 1 0 9600 0 -1 3482
box 369 500 1054 1856
use hgu_sw_cap_nmos  x7
timestamp 1699326276
transform 1 0 9952 0 1 -246
box 368 546 1040 1833
use hgu_pfet_hvt_stack_in_delay  x8
timestamp 1699184006
transform -1 0 10061 0 -1 2980
box -98 40 268 947
use hgu_nfet_hvt_stack_in_delay  x9
timestamp 1699184006
transform -1 0 10108 0 1 536
box -90 -235 303 886
use sky130_fd_sc_hd__inv_1  x10 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1697965495
transform 1 0 9300 0 1 1760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x11
timestamp 1697965495
transform -1 0 9760 0 1 1760
box -38 -48 314 592
use sky130_fd_pr__nfet_01v8_MVW3GX  XM1
timestamp 1698807554
transform 1 0 15828 0 -1 1520
box -125 -130 125 68
use sky130_fd_pr__nfet_01v8_L7T3GD  XM13
timestamp 1698825334
transform 1 0 15688 0 1 1520
box -73 -69 73 70
use sky130_fd_pr__nfet_01v8_L7T3GD  XM15
timestamp 1698825334
transform 1 0 15688 0 1 1382
box -73 -69 73 70
use sky130_fd_pr__pfet_01v8_hvt_M479BZ  XM46
timestamp 1698807554
transform 1 0 15688 0 1 1723
box -110 -80 109 88
use sky130_fd_pr__pfet_01v8_hvt_M479BZ  XM47
timestamp 1698807554
transform 1 0 15688 0 1 1861
box -110 -80 109 88
use sky130_fd_pr__pfet_01v8_hvt_M433PY  XM48
timestamp 1698807554
transform 1 0 15828 0 1 1723
box -161 -139 161 90
<< labels >>
flabel metal1 9275 1596 9943 1643 0 FreeSans 320 0 0 0 IN
port 1 nsew
flabel metal1 15751 1594 15933 1640 0 FreeSans 320 0 0 0 OUT
port 2 nsew
flabel metal1 9238 1979 9376 2013 0 FreeSans 320 0 0 0 code[3]
port 5 nsew
flabel metal1 14153 268 14211 1445 0 FreeSans 320 0 0 0 code[1]
port 8 nsew
flabel metal1 11727 268 11785 1445 0 FreeSans 320 0 0 0 code[2]
port 10 nsew
flabel metal4 9344 2338 9762 2948 0 FreeSans 320 0 0 0 VDD
port 17 nsew
flabel metal4 9372 291 9748 1728 0 FreeSans 320 0 0 0 VSS
port 19 nsew
flabel metal2 9702 1394 10138 1440 0 FreeSans 320 0 0 0 code_offset
port 21 nsew
flabel metal1 15009 267 15068 1448 0 FreeSans 320 0 0 0 code[0]
port 22 nsew
<< end >>
