magic
tech sky130A
magscale 1 2
timestamp 1699443150
<< error_s >>
rect 1298 898 1380 942
rect 1552 524 1634 898
<< nwell >>
rect 1663 898 2556 1022
rect 1552 524 2556 898
rect 1693 517 2411 524
<< nmos >>
rect 1779 69 1823 449
rect 1881 69 1925 449
rect 1983 69 2027 449
rect 2085 69 2129 449
rect 2187 69 2231 449
rect 2289 69 2333 449
<< pmos >>
rect 1775 606 1819 986
rect 1877 606 1921 986
rect 1979 606 2023 986
rect 2081 606 2125 986
rect 2183 606 2227 986
rect 2285 606 2329 986
<< ndiff >>
rect 1721 437 1779 449
rect 1721 118 1733 437
rect 1767 118 1779 437
rect 1721 69 1779 118
rect 1823 356 1881 449
rect 1823 81 1835 356
rect 1869 81 1881 356
rect 1823 69 1881 81
rect 1925 437 1983 449
rect 1925 81 1937 437
rect 1971 81 1983 437
rect 1925 69 1983 81
rect 2027 363 2085 449
rect 2027 81 2039 363
rect 2073 81 2085 363
rect 2027 69 2085 81
rect 2129 437 2187 449
rect 2129 81 2141 437
rect 2175 81 2187 437
rect 2129 69 2187 81
rect 2231 437 2289 449
rect 2231 81 2243 437
rect 2277 81 2289 437
rect 2231 69 2289 81
rect 2333 437 2392 449
rect 2333 121 2345 437
rect 2379 121 2392 437
rect 2333 69 2392 121
<< pdiff >>
rect 1722 946 1775 986
rect 1722 618 1730 946
rect 1764 618 1775 946
rect 1722 606 1775 618
rect 1819 974 1877 986
rect 1819 618 1831 974
rect 1865 618 1877 974
rect 1819 606 1877 618
rect 1921 974 1979 986
rect 1921 618 1933 974
rect 1967 618 1979 974
rect 1921 606 1979 618
rect 2023 974 2081 986
rect 2023 695 2035 974
rect 2069 695 2081 974
rect 2023 606 2081 695
rect 2125 974 2183 986
rect 2125 618 2137 974
rect 2171 618 2183 974
rect 2125 606 2183 618
rect 2227 974 2285 986
rect 2227 695 2239 974
rect 2273 695 2285 974
rect 2227 606 2285 695
rect 2329 948 2387 986
rect 2329 618 2341 948
rect 2375 618 2387 948
rect 2329 606 2387 618
<< ndiffc >>
rect 1733 118 1767 437
rect 1835 81 1869 356
rect 1937 81 1971 437
rect 2039 81 2073 363
rect 2141 81 2175 437
rect 2243 81 2277 437
rect 2345 121 2379 437
<< pdiffc >>
rect 1730 618 1764 946
rect 1831 618 1865 974
rect 1933 618 1967 974
rect 2035 695 2069 974
rect 2137 618 2171 974
rect 2239 695 2273 974
rect 2341 618 2375 948
<< poly >>
rect 1775 986 1819 1012
rect 1877 986 1921 1012
rect 1979 986 2023 1012
rect 2081 986 2125 1012
rect 2183 986 2227 1012
rect 2285 986 2329 1012
rect 1775 590 1819 606
rect 1877 590 1921 606
rect 1775 556 1921 590
rect 1775 504 1821 556
rect 1886 504 1921 556
rect 1979 591 2023 606
rect 2081 591 2125 606
rect 2183 591 2227 606
rect 2285 591 2329 606
rect 1979 587 2329 591
rect 1979 548 2333 587
rect 1979 536 2220 548
rect 1775 494 1921 504
rect 2187 496 2220 536
rect 2285 496 2333 548
rect 1775 468 2129 494
rect 1779 464 2129 468
rect 1779 449 1823 464
rect 1881 449 1925 464
rect 1983 449 2027 464
rect 2085 449 2129 464
rect 2187 464 2333 496
rect 2187 449 2231 464
rect 2289 449 2333 464
rect 1779 43 1823 69
rect 1881 43 1925 69
rect 1983 43 2027 69
rect 2085 43 2129 69
rect 2187 43 2231 69
rect 2289 43 2333 69
<< polycont >>
rect 1821 504 1886 556
rect 2220 496 2285 548
<< locali >>
rect 1831 974 1865 990
rect 1730 946 1764 971
rect 1764 618 1831 645
rect 1933 974 1967 990
rect 1865 618 1933 645
rect 2035 974 2069 990
rect 2035 679 2069 695
rect 2137 974 2171 990
rect 1967 618 2137 645
rect 2239 974 2273 990
rect 2239 679 2273 695
rect 2341 948 2375 964
rect 2171 618 2341 645
rect 1730 602 2375 618
rect 1804 504 1821 556
rect 1886 504 1902 556
rect 2009 455 2093 602
rect 2204 496 2220 548
rect 2285 496 2301 548
rect 1729 437 2379 455
rect 1729 118 1733 437
rect 1767 414 1937 437
rect 1729 94 1767 118
rect 1835 356 1869 380
rect 1835 65 1869 81
rect 1971 413 2141 437
rect 1937 65 1971 81
rect 2039 363 2073 379
rect 2039 65 2073 81
rect 2175 413 2243 437
rect 2141 65 2175 81
rect 2277 413 2345 437
rect 2344 121 2345 413
rect 2344 104 2379 121
rect 2243 65 2277 81
use adc_array_wafflecap_gate  adc_array_wafflecap_gate_0
timestamp 1671464254
transform 1 0 376 0 1 -62
box 0 0 1004 1004
use adc_gate_switch  adc_gate_switch_0
timestamp 1699443150
transform 1 0 2353 0 1 -81
box 318 245 1399 957
<< end >>
