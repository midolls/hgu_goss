magic
tech sky130A
magscale 1 2
timestamp 1699365206
<< error_p >>
rect 19 114 77 120
rect 19 80 31 114
rect 19 74 77 80
rect -77 -80 -19 -74
rect -77 -114 -65 -80
rect -77 -120 -19 -114
<< pwell >>
rect -263 -252 263 252
<< nmos >>
rect -63 -42 -33 42
rect 33 -42 63 42
<< ndiff >>
rect -125 30 -63 42
rect -125 -30 -113 30
rect -79 -30 -63 30
rect -125 -42 -63 -30
rect -33 30 33 42
rect -33 -30 -17 30
rect 17 -30 33 30
rect -33 -42 33 -30
rect 63 30 125 42
rect 63 -30 79 30
rect 113 -30 125 30
rect 63 -42 125 -30
<< ndiffc >>
rect -113 -30 -79 30
rect -17 -30 17 30
rect 79 -30 113 30
<< psubdiff >>
rect -227 182 -131 216
rect 131 182 227 216
rect -227 120 -193 182
rect 193 120 227 182
rect -227 -182 -193 -120
rect 193 -182 227 -120
rect -227 -216 -131 -182
rect 131 -216 227 -182
<< psubdiffcont >>
rect -131 182 131 216
rect -227 -120 -193 120
rect 193 -120 227 120
rect -131 -216 131 -182
<< poly >>
rect 15 114 81 130
rect 15 80 31 114
rect 65 80 81 114
rect -63 42 -33 68
rect 15 64 81 80
rect 33 42 63 64
rect -63 -64 -33 -42
rect -81 -80 -15 -64
rect 33 -68 63 -42
rect -81 -114 -65 -80
rect -31 -114 -15 -80
rect -81 -130 -15 -114
<< polycont >>
rect 31 80 65 114
rect -65 -114 -31 -80
<< locali >>
rect -227 182 -131 216
rect 131 182 227 216
rect -227 120 -193 182
rect 193 120 227 182
rect 15 80 31 114
rect 65 80 81 114
rect -113 30 -79 46
rect -113 -46 -79 -30
rect -17 30 17 46
rect -17 -46 17 -30
rect 79 30 113 46
rect 79 -46 113 -30
rect -81 -114 -65 -80
rect -31 -114 -15 -80
rect -227 -182 -193 -120
rect 193 -182 227 -120
rect -227 -216 -131 -182
rect 131 -216 227 -182
<< viali >>
rect 31 80 65 114
rect -113 -30 -79 30
rect -17 -30 17 30
rect 79 -30 113 30
rect -65 -114 -31 -80
<< metal1 >>
rect 19 114 77 120
rect 19 80 31 114
rect 65 80 77 114
rect 19 74 77 80
rect -119 30 -73 42
rect -119 -30 -113 30
rect -79 -30 -73 30
rect -119 -42 -73 -30
rect -23 30 23 42
rect -23 -30 -17 30
rect 17 -30 23 30
rect -23 -42 23 -30
rect 73 30 119 42
rect 73 -30 79 30
rect 113 -30 119 30
rect 73 -42 119 -30
rect -77 -80 -19 -74
rect -77 -114 -65 -80
rect -31 -114 -19 -80
rect -77 -120 -19 -114
<< properties >>
string FIXED_BBOX -210 -199 210 199
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.42 l 0.15 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
