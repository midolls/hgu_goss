* NGSPICE file created from hgu_clk_sample_flat.ext - technology: sky130A

.subckt hgu_clk_sample_flat set reset sample_delay_offset CAP_CTRL_CODE0[2] CAP_CTRL_CODE0[1]
+ CAP_CTRL_CODE1[2] CAP_CTRL_CODE1[1] CAP_CTRL_CODE1[0] CAP_CTRL_CODE2[2] CAP_CTRL_CODE2[1]
+ CAP_CTRL_CODE3[2] CAP_CTRL_CODE3[1] CAP_CTRL_CODE3[0] CAP_CTRL_CODE1[3] CAP_CTRL_CODE3[3]
+ sample_clk_b sample_clk clk CAP_CTRL_CODE2[3] CAP_CTRL_CODE0[0] CAP_CTRL_CODE0[3]
+ CAP_CTRL_CODE2[0] vdd vss
X0 a_11371_5456# x2.x1.IN a_11283_5456# vss.t99 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X1 vss.t25 a_3106_6090# a_3041_6494# vss.t24 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X2 x2.x4.x2.floating CAP_CTRL_CODE0[0].t0 x2.x4.x9.output_stack vss.t68 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.124 ps=1.43 w=0.42 l=0.15
X3 a_4687_7397# x3.A a_4599_7535# vdd.t82 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X4 x2.x1.x5[7].floating.t7 x2.x1.x10.Y.t2 x2.x1.x9.output_stack vdd.t4 sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X5 x7.A x2.x3.x9.output_stack a_4047_2819# vdd.t46 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.0651 ps=0.73 w=0.42 l=0.15
X6 a_2325_6090# x1.x3.Y vdd.t36 vdd.t35 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X7 a_10112_1680# x2.x3.IN a_10024_1818# vdd.t29 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X8 x2.x4.x9.output_stack x2.x4.x10.Y.t2 x2.x4.x5[7].floating.t7 vdd.t1 sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X9 a_10472_6534# x2.x4.x9.output_stack x2.x1.IN vdd.t32 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.122 ps=1.42 w=0.42 l=0.15
X10 a_3340_6116# a_2932_6494# a_3106_6090# vdd.t73 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X11 a_10065_3897# x2.x3.IN a_9977_3897# vss.t29 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X12 a_2325_6090# a_2151_6116# a_2465_6482# vss.t55 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X13 a_11396_7121# x2.x1.IN a_11308_6983# vdd.t93 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X14 x2.x1.x10.Y.t0 CAP_CTRL_CODE1[3].t0 vdd.t111 vdd.t110 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X15 x2.x4.x10.Y.t0 CAP_CTRL_CODE0[3].t0 vss.t2 vss.t1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X16 a_2151_6116# a_1870_6122# a_2058_6116# vdd.t70 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X17 a_4734_5594# x3.A a_4662_5594# vss.t92 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X18 x2.x2.x5[7].floating.t7 x2.x2.x10.Y.t2 x2.x2.x9.output_stack vdd.t62 sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X19 vss.t63 a_2678_2626# sample_clk.t2 vss.t60 sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X20 a_16846_3483# x2.x2.IN a_16774_3483# vss.t41 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X21 x2.x2.x6.SW sample_delay_offset.t0 vdd.t127 vdd.t126 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X22 vdd.t18 a_3106_6090# a_3813_6132# vdd.t17 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X23 vdd.t64 x7.Y x3.Y vdd.t44 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X24 x2.x3.x9.output_stack CAP_CTRL_CODE3[2].t0 x2.x3.x4[3].floating vss.t66 sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X25 vdd.t55 a_2678_2626# sample_clk.t5 vdd.t52 sky130_fd_pr__pfet_01v8 ad=0.391 pd=3.14 as=0.208 ps=1.59 w=1.26 l=0.15
X26 a_17181_6534# x2.x1.x9.output_stack x2.x2.IN vdd.t39 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.122 ps=1.42 w=0.42 l=0.15
X27 x3.A a_3813_6132# vdd.t59 vdd.t58 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X28 x2.x2.x7.floating sample_delay_offset.t1 x2.x2.x9.output_stack vss.t67 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X29 x2.x1.x9.output_stack x2.x1.x6.SW x2.x1.x6.floating vdd.t99 sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X30 a_10472_6193# x2.x1.IN vdd.t92 vss.t105 sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X31 vdd.t131 CAP_CTRL_CODE3[3].t0 x2.x3.x10.Y.t1 vdd.t130 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X32 vdd.t12 a_2678_2006# sample_clk_b.t5 vdd.t9 sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.391 ps=3.14 w=1.26 l=0.15
X33 a_4662_5180# x3.A a_4574_5180# vss.t91 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X34 vss.t104 x2.x1.IN a_11371_5180# vss.t100 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X35 a_16846_3759# x2.x2.IN a_16774_3759# vss.t41 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X36 a_4047_3022# x7.A vdd.t48 vss.t54 sky130_fd_pr__nfet_01v8 ad=0.0651 pd=0.73 as=0.0693 ps=0.75 w=0.42 l=0.15
X37 a_11371_5870# x2.x1.IN a_11283_5732# vss.t99 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X38 x2.x1.x9.output_stack x2.x1.x10.Y.t3 x2.x1.x5[7].floating.t6 vdd.t4 sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X39 a_16774_4173# x2.x2.IN vss.t46 vss.t40 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X40 x2.x3.x5[7].floating.t7 x2.x3.x10.Y.t2 x2.x3.x9.output_stack vdd.t0 sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X41 x2.x4.x9.output_stack CAP_CTRL_CODE0[2].t0 x2.x4.x4[3].floating vss.t75 sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X42 a_4662_5456# x3.A a_4574_5456# vss.t91 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X43 a_11443_5318# x2.x1.IN a_11371_5456# vss.t100 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X44 x2.x1.x5[7].floating.t5 x2.x1.x10.Y.t4 x2.x1.x9.output_stack vdd.t4 sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X45 a_16774_3345# x2.x2.IN a_16686_3345# vss.t40 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X46 x2.x3.x9.output_stack x2.x3.x10.Y.t3 x2.x3.x5[7].floating.t6 vdd.t0 sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X47 x2.x4.x5[7].floating.t6 x2.x4.x10.Y.t3 x2.x4.x9.output_stack vdd.t1 sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X48 a_17181_6534# x2.x2.IN vss.t45 vdd.t39 sky130_fd_pr__pfet_01v8_hvt ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X49 x2.x1.x9.output_stack sample_delay_offset.t2 x2.x1.x7.floating vss.t132 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X50 vdd.t61 a_3056_2150# a_2678_2006# vdd.t60 sky130_fd_pr__pfet_01v8 ad=0.365 pd=3.1 as=0.365 ps=3.1 w=1.26 l=0.15
X51 x2.x3.x5[7].floating.t5 x2.x3.x10.Y.t4 x2.x3.x9.output_stack vdd.t0 sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X52 x2.x1.x9.output_stack x2.x1.x10.Y.t5 x2.x1.x5[7].floating.t4 vdd.t4 sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X53 x1.x4.Y reset.t0 vdd.t129 vdd.t128 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X54 a_10137_3759# x2.x3.IN a_10065_3897# vss.t27 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X55 vss.t18 a_2678_2006# sample_clk_b.t2 vss.t17 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X56 x2.x2.x9.output_stack x2.x2.x10.Y.t3 x2.x2.x5[7].floating.t6 vdd.t2 sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X57 x2.x1.x5[7].floating.t3 x2.x1.x10.Y.t6 x2.x1.x9.output_stack vdd.t4 sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X58 a_11371_6146# x2.x1.IN a_11283_6008# vss.t99 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X59 a_4687_7121# x3.A a_4599_6983# vdd.t81 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X60 x2.x2.x4[3].floating CAP_CTRL_CODE2[2].t0 x2.x2.x9.output_stack vss.t124 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X61 vdd.t118 sample_delay_offset.t3 x2.x1.x6.SW vdd.t117 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X62 a_11371_5318# x2.x1.IN a_11283_5180# vss.t99 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X63 a_10112_2232# x2.x3.IN a_10024_2094# vdd.t28 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X64 a_4047_2819# x7.A vss.t53 vdd.t46 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.0693 ps=0.75 w=0.42 l=0.15
X65 x2.x2.x9.output_stack CAP_CTRL_CODE2[2].t1 x2.x2.x4[3].floating vss.t118 sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X66 a_2058_6116# x1.x2.D vss.t10 vss.t9 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X67 a_10065_3483# x2.x3.IN a_9977_3345# vss.t29 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X68 vss.t138 clk.t0 a_1704_6122# vss.t137 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X69 a_10472_6193# x2.x4.x9.output_stack vss.t35 vss.t34 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X70 x2.x1.x9.output_stack CAP_CTRL_CODE1[1].t0 x2.x1.x3[1].floating vss.t47 sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X71 x2.x2.x6.floating x2.x2.x6.SW x2.x2.x9.output_stack vdd.t103 sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X72 vss.t93 x3.A a_4662_5180# vss.t92 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X73 a_4662_5870# x3.A a_4574_5732# vss.t91 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X74 a_11443_5870# x2.x1.IN a_11371_5870# vss.t100 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X75 a_10065_3759# x2.x3.IN a_9977_3621# vss.t29 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X76 x2.x2.x4[3].floating CAP_CTRL_CODE2[2].t2 x2.x2.x9.output_stack vss.t76 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X77 vdd.t51 a_3056_2936# a_2678_2626# vdd.t50 sky130_fd_pr__pfet_01v8 ad=0.365 pd=3.1 as=0.365 ps=3.1 w=1.26 l=0.15
X78 vss.t117 a_2325_6090# a_2259_6494# vss.t116 sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X79 a_3106_6090# x1.x3.Y vdd.t34 vdd.t33 sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X80 x2.x4.x9.output_stack x2.x4.x10.Y.t4 x2.x4.x5[7].floating.t5 vdd.t1 sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X81 a_16846_4035# x2.x2.IN a_16774_4173# vss.t41 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X82 x2.x4.x5[7].floating.t4 x2.x4.x10.Y.t5 x2.x4.x9.output_stack vdd.t1 sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X83 a_17181_6193# x2.x1.x9.output_stack vss.t85 vss.t84 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X84 a_4734_5318# x3.A a_4662_5456# vss.t92 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X85 x2.x3.x6.SW sample_delay_offset.t4 vdd.t109 vdd.t108 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X86 x2.x3.x9.output_stack x2.x3.x10.Y.t5 x2.x3.x5[7].floating.t4 vdd.t0 sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X87 sample_clk.t1 a_2678_2626# vss.t62 vss.t60 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X88 vdd.t16 a_3106_6090# a_3018_6116# vdd.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X89 x2.x4.x9.output_stack sample_delay_offset.t5 x2.x4.x7.floating vss.t129 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X90 a_16846_3207# x2.x2.IN a_16774_3345# vss.t41 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X91 vss.t112 x2.x2.x9.output_stack a_10756_3022# vss.t111 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X92 sample_clk.t4 a_2678_2626# vdd.t54 vdd.t52 sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X93 vss.t52 x7.A x7.Y vss.t51 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X94 a_3106_6090# a_2932_6494# a_3222_6482# vss.t86 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X95 vdd.t91 x2.x1.IN a_10472_6193# vss.t103 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0651 ps=0.73 w=0.42 l=0.15
X96 a_11371_5732# x2.x1.IN a_11283_5732# vss.t99 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X97 x2.x3.x9.output_stack x2.x3.x10.Y.t6 x2.x3.x5[7].floating.t3 vdd.t0 sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X98 vdd.t47 x7.A a_4047_3022# vss.t50 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X99 a_11396_7397# x2.x1.IN a_11308_7259# vdd.t90 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X100 a_3222_6482# x1.x3.Y vss.t39 vss.t38 sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X101 x1.x2.D a_3106_6090# vss.t23 vss.t22 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X102 a_4662_6146# x3.A a_4574_6008# vss.t91 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X103 x2.x1.x9.output_stack x2.x1.IN a_11371_6146# vss.t100 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X104 vdd.t116 a_2619_6316# a_2569_6116# vdd.t115 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X105 x2.x3.x4[3].floating CAP_CTRL_CODE3[2].t1 x2.x3.x9.output_stack vss.t98 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X106 vdd.t66 sample_delay_offset.t6 x2.x4.x6.SW vdd.t65 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X107 a_4662_5318# x3.A a_4574_5180# vss.t91 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X108 a_16774_4035# x2.x2.IN a_16686_3897# vss.t40 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X109 a_11443_5318# x2.x1.IN a_11371_5318# vss.t100 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X110 a_10472_6534# x2.x1.IN vss.t102 vdd.t32 sky130_fd_pr__pfet_01v8_hvt ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X111 x2.x4.x3[1].floating CAP_CTRL_CODE0[1].t0 x2.x4.x9.output_stack vss.t0 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X112 a_10137_3483# x2.x3.IN a_10065_3483# vss.t27 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X113 x2.x2.x9.output_stack CAP_CTRL_CODE2[1].t0 x2.x2.x3[1].floating vss.t69 sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X114 a_16774_3207# x2.x2.IN x2.x2.x9.output_stack vss.t40 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X115 x2.x1.x5[7].floating.t2 x2.x1.x10.Y.t7 x2.x1.x9.output_stack vdd.t4 sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X116 vdd.t41 x2.x2.IN a_17181_6193# vss.t44 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0651 ps=0.73 w=0.42 l=0.15
X117 a_16821_1956# x2.x2.IN a_16733_2094# vdd.t37 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X118 vdd.t101 x2.x2.x9.output_stack a_10756_2819# vdd.t100 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X119 a_2465_6482# a_2619_6316# a_2325_6090# vss.t128 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X120 x2.x4.x9.output_stack CAP_CTRL_CODE0[1].t1 x2.x4.x3[1].floating vss.t8 sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X121 x2.x2.x5[7].floating.t5 x2.x2.x10.Y.t4 x2.x2.x9.output_stack vdd.t94 sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X122 x2.x1.x9.output_stack CAP_CTRL_CODE1[2].t0 x2.x1.x4[3].floating vss.t48 sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X123 x2.x2.x9.output_stack CAP_CTRL_CODE2[0].t0 x2.x2.x2.floating vss.t110 sky130_fd_pr__nfet_01v8 ad=0.124 pd=1.43 as=0.122 ps=1.42 w=0.42 l=0.15
X124 x2.x1.x4[3].floating CAP_CTRL_CODE1[2].t1 x2.x1.x9.output_stack vss.t19 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X125 a_4734_5870# x3.A a_4662_5870# vss.t92 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X126 a_10137_3759# x2.x3.IN a_10065_3759# vss.t27 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X127 a_2235_6116# a_1704_6122# a_2151_6116# vdd.t98 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X128 a_3553_3025# x3.A x3.Y vss.t78 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X129 a_11371_6008# x2.x1.IN a_11283_6008# vss.t99 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X130 a_10065_4173# x2.x3.IN vss.t32 vss.t29 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X131 vss.t49 x7.A a_4047_2819# vdd.t46 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X132 vdd.t114 a_2619_6316# a_3340_6116# vdd.t113 sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X133 a_10065_3345# x2.x3.IN a_9977_3345# vss.t29 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X134 vss.t134 x3.Y a_3056_2936# vss.t133 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X135 a_1870_6122# a_1704_6122# vdd.t97 vdd.t96 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X136 x2.x1.x9.output_stack x2.x1.IN a_11308_6983# vdd.t89 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X137 a_4662_5732# x3.A a_4574_5732# vss.t91 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X138 a_11443_5594# x2.x1.IN a_11371_5732# vss.t100 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X139 a_4687_7397# x3.A a_4599_7259# vdd.t80 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X140 x2.x4.x9.output_stack x3.A a_4662_6146# vss.t92 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X141 x1.x3.Y set.t0 vss.t89 vss.t88 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X142 a_16774_3621# x2.x2.IN a_16686_3621# vss.t40 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X143 vss.t123 CAP_CTRL_CODE2[3].t0 x2.x2.x10.Y.t0 vss.t122 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X144 x2.x4.x9.output_stack x2.x4.x6.SW x2.x4.x6.floating vdd.t102 sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X145 a_16846_4035# x2.x2.IN a_16774_4035# vss.t41 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X146 a_4734_5318# x3.A a_4662_5318# vss.t92 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X147 vss.t61 a_2678_2626# sample_clk.t0 vss.t60 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X148 a_16821_1680# x2.x2.IN vdd.t40 vdd.t37 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X149 x2.x3.x9.output_stack CAP_CTRL_CODE3[1].t0 x2.x3.x3[1].floating vss.t130 sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X150 a_16846_3207# x2.x2.IN a_16774_3207# vss.t41 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X151 x2.x3.IN x2.x2.x9.output_stack a_10756_3022# vss.t111 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0651 ps=0.73 w=0.42 l=0.15
X152 a_2058_6116# x1.x2.D vdd.t6 vdd.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X153 vdd.t53 a_2678_2626# sample_clk.t3 vdd.t52 sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.391 ps=3.14 w=1.26 l=0.15
X154 vss.t59 a_3056_2936# a_2678_2626# vss.t58 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X155 x2.x4.x9.output_stack CAP_CTRL_CODE0[2].t1 x2.x4.x4[3].floating vss.t121 sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X156 x2.x3.x9.output_stack CAP_CTRL_CODE3[0].t0 x2.x3.x2.floating vss.t119 sky130_fd_pr__nfet_01v8 ad=0.124 pd=1.43 as=0.122 ps=1.42 w=0.42 l=0.15
X157 x2.x4.x10.Y.t1 CAP_CTRL_CODE0[3].t1 vdd.t43 vdd.t42 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X158 a_3018_6116# a_1870_6122# a_2932_6494# vdd.t69 sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X159 x2.x4.x4[3].floating CAP_CTRL_CODE0[2].t2 x2.x4.x9.output_stack vss.t33 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X160 a_16821_1956# x2.x2.IN a_16733_1818# vdd.t37 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X161 a_11396_7121# x2.x1.IN a_11308_7259# vdd.t88 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X162 a_2932_6494# a_1870_6122# a_2837_6438# vss.t83 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X163 x2.x3.x5[7].floating.t2 x2.x3.x10.Y.t7 x2.x3.x9.output_stack vdd.t0 sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X164 a_4662_6008# x3.A a_4574_6008# vss.t91 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X165 a_11443_5870# x2.x1.IN a_11371_6008# vss.t100 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X166 vdd.t107 a_2325_6090# a_2235_6116# vdd.t106 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X167 x2.x1.x9.output_stack x2.x1.x10.Y.t8 x2.x1.x5[7].floating.t1 vdd.t4 sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X168 a_10137_4035# x2.x3.IN a_10065_4173# vss.t27 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X169 x2.x3.x7.floating sample_delay_offset.t7 x2.x3.x9.output_stack vss.t77 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X170 vss.t101 x2.x1.IN a_10472_6534# vdd.t32 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0651 ps=0.73 w=0.42 l=0.15
X171 a_10137_3207# x2.x3.IN a_10065_3345# vss.t27 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X172 x2.x1.x10.Y.t1 CAP_CTRL_CODE1[3].t1 vss.t136 vss.t135 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X173 a_3041_6494# a_1704_6122# a_2932_6494# vss.t109 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X174 x2.x4.x9.output_stack x3.A a_4599_6983# vdd.t79 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X175 x2.x1.x2.floating CAP_CTRL_CODE1[0].t0 x2.x1.x9.output_stack vss.t139 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.124 ps=1.43 w=0.42 l=0.15
X176 a_4734_5594# x3.A a_4662_5732# vss.t92 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X177 x2.x2.x9.output_stack CAP_CTRL_CODE2[2].t3 x2.x2.x4[3].floating vss.t4 sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X178 a_16846_3483# x2.x2.IN a_16774_3621# vss.t41 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X179 x2.x2.x9.output_stack x2.x2.x10.Y.t5 x2.x2.x5[7].floating.t4 vdd.t74 sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X180 x2.x3.IN x2.x2.x9.output_stack a_10756_2819# vdd.t100 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.0651 ps=0.73 w=0.42 l=0.15
X181 a_10756_3022# x2.x3.IN vdd.t27 vss.t31 sky130_fd_pr__nfet_01v8 ad=0.0651 pd=0.73 as=0.0693 ps=0.75 w=0.42 l=0.15
X182 a_2151_6116# a_1704_6122# a_2058_6116# vss.t108 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X183 vss.t43 x2.x2.IN a_17181_6534# vdd.t39 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0651 ps=0.73 w=0.42 l=0.15
X184 vdd.t8 x1.x4.Y a_2619_6316# vdd.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X185 a_10065_4035# x2.x3.IN a_9977_3897# vss.t29 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X186 x2.x3.x6.floating x2.x3.x6.SW x2.x3.x9.output_stack vdd.t119 sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X187 a_10065_3207# x2.x3.IN x2.x3.x9.output_stack vss.t29 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X188 vdd.t45 x7.A x7.Y vdd.t44 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X189 vdd.t87 x2.x1.IN a_11308_7535# vdd.t86 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X190 vss.t12 x1.x4.Y a_2619_6316# vss.t11 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X191 x2.x4.x9.output_stack x2.x4.x10.Y.t6 x2.x4.x5[7].floating.t3 vdd.t1 sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X192 a_10112_1956# x2.x3.IN a_10024_2094# vdd.t26 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X193 vdd.t11 a_2678_2006# sample_clk_b.t4 vdd.t9 sky130_fd_pr__pfet_01v8 ad=0.391 pd=3.14 as=0.208 ps=1.59 w=1.26 l=0.15
X194 a_2790_6116# a_2325_6090# vdd.t105 vdd.t104 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X195 x2.x4.x5[7].floating.t2 x2.x4.x10.Y.t7 x2.x4.x9.output_stack vdd.t1 sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X196 x2.x2.x6.SW sample_delay_offset.t8 vss.t97 vss.t96 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X197 a_4687_7121# x3.A a_4599_7259# vdd.t78 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X198 vss.t65 x2.x3.x9.output_stack a_4047_3022# vss.t64 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X199 x2.x2.x5[7].floating.t3 x2.x2.x10.Y.t6 x2.x2.x9.output_stack vdd.t124 sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X200 x3.A a_3813_6132# vss.t71 vss.t70 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X201 a_4734_5870# x3.A a_4662_6008# vss.t92 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X202 vss.t95 CAP_CTRL_CODE3[3].t1 x2.x3.x10.Y.t0 vss.t94 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X203 x2.x3.x9.output_stack CAP_CTRL_CODE3[2].t2 x2.x3.x4[3].floating vss.t7 sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X204 a_16821_2232# x2.x2.IN x2.x2.x9.output_stack vdd.t37 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X205 a_2837_6438# a_2325_6090# vss.t115 vss.t114 sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X206 x1.x4.Y reset.t1 vss.t125 vss.t88 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X207 a_2465_6482# x1.x3.Y vss.t37 vss.t36 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X208 x1.x2.D a_3106_6090# vdd.t14 vdd.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X209 x2.x3.x4[3].floating CAP_CTRL_CODE3[2].t3 x2.x3.x9.output_stack vss.t3 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X210 vss.t79 x7.Y a_3553_3025# vss.t78 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X211 vss.t57 sample_delay_offset.t9 x2.x1.x6.SW vss.t56 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X212 x2.x1.x9.output_stack x2.x1.x10.Y.t9 x2.x1.x5[7].floating.t0 vdd.t4 sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X213 a_10756_2819# x2.x3.IN vss.t30 vdd.t25 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.0693 ps=0.75 w=0.42 l=0.15
X214 a_2569_6116# a_2151_6116# a_2325_6090# vdd.t49 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X215 x2.x1.x9.output_stack CAP_CTRL_CODE1[2].t2 x2.x1.x4[3].floating vss.t74 sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X216 a_16821_1680# x2.x2.IN a_16733_1818# vdd.t37 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X217 vss.t16 a_2678_2006# sample_clk_b.t1 vss.t15 sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X218 x2.x2.x9.output_stack x2.x2.x10.Y.t7 x2.x2.x5[7].floating.t2 vdd.t125 sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X219 a_16774_3897# x2.x2.IN a_16686_3897# vss.t40 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X220 x3.Y x3.A vdd.t77 vdd.t44 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X221 x2.x2.x3[1].floating CAP_CTRL_CODE2[1].t1 x2.x2.x9.output_stack vss.t131 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X222 vss.t21 a_3106_6090# a_3813_6132# vss.t20 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X223 x2.x4.x5[7].floating.t1 x2.x4.x10.Y.t8 x2.x4.x9.output_stack vdd.t1 sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X224 x2.x3.x9.output_stack x2.x3.x10.Y.t8 x2.x3.x5[7].floating.t1 vdd.t0 sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X225 a_10065_3621# x2.x3.IN a_9977_3621# vss.t29 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X226 vdd.t57 x2.x3.x9.output_stack a_4047_2819# vdd.t56 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X227 x2.x3.x5[7].floating.t0 x2.x3.x10.Y.t9 x2.x3.x9.output_stack vdd.t0 sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X228 vdd.t123 x3.Y a_3056_2936# vdd.t122 sky130_fd_pr__pfet_01v8 ad=0.406 pd=3.38 as=0.406 ps=3.38 w=1.4 l=0.15
X229 a_10472_6193# x2.x4.x9.output_stack x2.x1.IN vss.t34 sky130_fd_pr__nfet_01v8 ad=0.0651 pd=0.73 as=0.122 ps=1.42 w=0.42 l=0.15
X230 x2.x1.x4[3].floating CAP_CTRL_CODE1[2].t3 x2.x1.x9.output_stack vss.t87 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X231 a_11371_5594# x2.x1.IN a_11283_5456# vss.t99 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X232 a_10137_4035# x2.x3.IN a_10065_4035# vss.t27 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X233 a_10137_3207# x2.x3.IN a_10065_3207# vss.t27 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X234 a_10112_1680# x2.x3.IN vdd.t24 vdd.t23 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X235 vdd.t76 x3.A a_4599_7535# vdd.t75 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X236 x2.x2.x9.output_stack x2.x2.x10.Y.t8 x2.x2.x5[7].floating.t1 vdd.t112 sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X237 a_10472_6534# x2.x4.x9.output_stack vdd.t31 vdd.t30 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X238 a_1870_6122# a_1704_6122# vss.t107 vss.t106 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X239 a_17181_6193# x2.x1.x9.output_stack x2.x2.IN vss.t84 sky130_fd_pr__nfet_01v8 ad=0.0651 pd=0.73 as=0.122 ps=1.42 w=0.42 l=0.15
X240 a_10112_1956# x2.x3.IN a_10024_1818# vdd.t22 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X241 vdd.t21 x2.x3.IN a_10756_3022# vss.t28 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X242 a_2259_6494# a_1870_6122# a_2151_6116# vss.t82 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X243 vdd.t68 clk.t1 a_1704_6122# vdd.t67 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X244 a_11396_7397# x2.x1.IN a_11308_7535# vdd.t85 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X245 a_17181_6534# x2.x1.x9.output_stack vdd.t72 vdd.t71 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X246 vss.t81 sample_delay_offset.t10 x2.x4.x6.SW vss.t80 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X247 x2.x4.x9.output_stack x2.x4.x10.Y.t9 x2.x4.x5[7].floating.t0 vdd.t1 sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X248 sample_clk_b.t3 a_2678_2006# vdd.t10 vdd.t9 sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X249 x2.x3.x6.SW sample_delay_offset.t11 vss.t6 vss.t5 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X250 x2.x1.x3[1].floating CAP_CTRL_CODE1[1].t1 x2.x1.x9.output_stack vss.t126 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X251 vdd.t121 CAP_CTRL_CODE2[3].t1 x2.x2.x10.Y.t1 vdd.t120 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X252 a_17181_6193# x2.x2.IN vdd.t38 vss.t42 sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X253 a_16846_3759# x2.x2.IN a_16774_3897# vss.t41 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X254 x3.Y vdd.t132 a_3056_2150# vss.t90 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X255 x2.x3.x3[1].floating CAP_CTRL_CODE3[1].t1 x2.x3.x9.output_stack vss.t120 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X256 a_3222_6482# a_2619_6316# a_3106_6090# vss.t127 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X257 x7.A x2.x3.x9.output_stack a_4047_3022# vss.t64 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0651 ps=0.73 w=0.42 l=0.15
X258 a_10137_3483# x2.x3.IN a_10065_3621# vss.t27 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X259 a_16821_2232# x2.x2.IN a_16733_2094# vdd.t37 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X260 x2.x4.x4[3].floating CAP_CTRL_CODE0[2].t3 x2.x4.x9.output_stack vss.t113 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X261 a_4662_5594# x3.A a_4574_5456# vss.t91 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X262 a_11443_5594# x2.x1.IN a_11371_5594# vss.t100 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X263 x3.Y vss.t140 a_3056_2150# vdd.t3 sky130_fd_pr__pfet_01v8 ad=0.551 pd=4.38 as=0.551 ps=4.38 w=1.9 l=0.15
X264 a_16774_3483# x2.x2.IN a_16686_3345# vss.t40 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X265 vss.t73 a_3056_2150# a_2678_2006# vss.t72 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X266 x1.x3.Y set.t1 vdd.t84 vdd.t83 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X267 a_2932_6494# a_1704_6122# a_2790_6116# vdd.t95 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X268 vss.t26 x2.x3.IN a_10756_2819# vdd.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X269 a_11371_5180# x2.x1.IN a_11283_5180# vss.t99 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X270 a_16774_3759# x2.x2.IN a_16686_3621# vss.t40 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X271 sample_clk_b.t0 a_2678_2006# vss.t14 vss.t13 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X272 a_10112_2232# x2.x3.IN x2.x3.x9.output_stack vdd.t19 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X273 x2.x2.x5[7].floating.t0 x2.x2.x10.Y.t9 x2.x2.x9.output_stack vdd.t63 sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
R0 vss.n1171 vss.n1170 808007
R1 vss.n2024 vss.n2023 553784
R2 vss.n2111 vss.n2110 553379
R3 vss.t51 vss.n3185 118558
R4 vss.n1171 vss.n1169 21533.3
R5 vss.n1875 vss.n1874 15644.4
R6 vss.n2843 vss.n169 15644.4
R7 vss vss.t88 15460.2
R8 vss.n496 vss.n495 15155.6
R9 vss.n3186 vss 13072.6
R10 vss.n1170 vss.t90 9378.04
R11 vss vss.n118 8510.53
R12 vss.t17 vss.t133 5109.31
R13 vss.n3186 vss 2172.1
R14 vss.n3187 vss.n3186 2079.76
R15 vss.n3186 vss.n118 1586.32
R16 vss.t72 vss.t15 1302.76
R17 vss.n1203 vss.t96 1270.52
R18 vss vss.n1171 1176.9
R19 vss.n2023 vss.t56 1150.15
R20 vss.n2111 vss.t5 1136.78
R21 vss vss.t51 1100
R22 vss.n2003 vss 1043.16
R23 vss.n1200 vss.t122 1043.16
R24 vss.n2962 vss 984.212
R25 vss.n2943 vss.n2942 922.797
R26 vss.n3184 vss.t80 815.806
R27 vss.n1204 vss.n1142 782.529
R28 vss.n2121 vss 775.684
R29 vss.n1202 vss 775.684
R30 vss.n1170 vss.t72 696.082
R31 vss.t96 vss.n1202 641.946
R32 vss.n1949 vss.n1948 626.532
R33 vss.t15 vss.t13 613.062
R34 vss.t13 vss.t17 613.062
R35 vss.n564 vss 601.824
R36 vss.n1174 vss 601.824
R37 vss.n1199 vss.n1198 585
R38 vss.n1200 vss.n1199 585
R39 vss.n1176 vss.n1175 585
R40 vss.n1175 vss.n1174 585
R41 vss.n1199 vss.n1143 481.557
R42 vss.n3189 vss.n3188 431.957
R43 vss.n1242 vss.t139 424.519
R44 vss.n3204 vss.n3203 403.038
R45 vss.n4 vss.t140 393.514
R46 vss.n1975 vss.t111 360.534
R47 vss.t34 vss.n2109 360.534
R48 vss.n2907 vss 320.974
R49 vss.n609 vss 320.974
R50 vss.n3026 vss.n3025 295.61
R51 vss.n1147 vss.n1146 294.606
R52 vss.n1875 vss.t110 294.416
R53 vss.n2909 vss.n2908 292.5
R54 vss.n2908 vss.n2907 292.5
R55 vss.n2965 vss.n2964 292.5
R56 vss.n2964 vss.n2963 292.5
R57 vss.n3013 vss.n3012 292.5
R58 vss.n3014 vss.n3013 292.5
R59 vss.n3017 vss.n3016 292.5
R60 vss.n3016 vss.n3015 292.5
R61 vss.n3021 vss.n3020 292.5
R62 vss.n3020 vss.n3019 292.5
R63 vss.n3025 vss.n3024 292.5
R64 vss.n3031 vss.n3030 292.5
R65 vss.n3030 vss.n3029 292.5
R66 vss.n3036 vss.n3035 292.5
R67 vss.n3035 vss.n3034 292.5
R68 vss.n3040 vss.n3039 292.5
R69 vss.n3039 vss.n3038 292.5
R70 vss.n3047 vss.n3046 292.5
R71 vss.n3046 vss.n3045 292.5
R72 vss.n3051 vss.n3050 292.5
R73 vss.n3050 vss.n3049 292.5
R74 vss.n3055 vss.n3054 292.5
R75 vss.n3054 vss.n3053 292.5
R76 vss.n3060 vss.n3059 292.5
R77 vss.n3059 vss.n3058 292.5
R78 vss.n3065 vss.n3064 292.5
R79 vss.n3064 vss.n3063 292.5
R80 vss.n3070 vss.n3069 292.5
R81 vss.n3069 vss.n3068 292.5
R82 vss.n3074 vss.n3073 292.5
R83 vss.n3073 vss.n3072 292.5
R84 vss.n3079 vss.n3078 292.5
R85 vss.n3078 vss.n3077 292.5
R86 vss.n3083 vss.n3082 292.5
R87 vss.n3082 vss.n3081 292.5
R88 vss.n3090 vss.n3089 292.5
R89 vss.n3089 vss.n3088 292.5
R90 vss.n3094 vss.n3093 292.5
R91 vss.n3093 vss.n3092 292.5
R92 vss.n3099 vss.n3098 292.5
R93 vss.n3098 vss.n3097 292.5
R94 vss.n3103 vss.n3102 292.5
R95 vss.n3102 vss.n3101 292.5
R96 vss.n3114 vss.n3113 292.5
R97 vss.n3113 vss.n3112 292.5
R98 vss.n3107 vss.n3106 292.5
R99 vss.n3106 vss.n3105 292.5
R100 vss.n3118 vss.n3117 292.5
R101 vss.n3117 vss.n3116 292.5
R102 vss.n3129 vss.n3128 292.5
R103 vss.n3128 vss.n3127 292.5
R104 vss.n3123 vss.n3122 292.5
R105 vss.n3122 vss.n3121 292.5
R106 vss.n2123 vss.n2122 292.5
R107 vss.n2122 vss.n2121 292.5
R108 vss.n611 vss.n610 292.5
R109 vss.n610 vss.n609 292.5
R110 vss.n1201 vss.n1126 292.5
R111 vss.n1173 vss.n1147 292.5
R112 vss.n1142 vss.n1141 292.5
R113 vss.n1202 vss.n1142 292.5
R114 vss.n1126 vss.n1124 292.5
R115 vss.n3228 vss.n3227 292.5
R116 vss.n3218 vss.n3217 292.5
R117 vss.n113 vss.n112 292.5
R118 vss.n3234 vss.n3233 292.5
R119 vss.n1169 vss.n1168 292.168
R120 vss.t119 vss.n2843 289.248
R121 vss.t88 vss 248.185
R122 vss.t105 vss.t28 234.535
R123 vss.n2893 vss.n2892 227.357
R124 vss.n2022 vss.n601 227.357
R125 vss.n600 vss.n599 213.982
R126 vss.n1201 vss.n1200 213.982
R127 vss.n566 vss.n565 187.234
R128 vss.n1173 vss.n1172 187.234
R129 vss.n3062 vss.t115 184.713
R130 vss.t78 vss 182.773
R131 vss.n3185 vss.n3184 178.941
R132 vss.n2945 vss.n2944 173.861
R133 vss.n2005 vss.n2004 173.861
R134 vss.n1084 vss.t47 153.446
R135 vss.n1023 vss.t124 153.446
R136 vss.n1007 vss.t118 153.446
R137 vss.n1392 vss.t19 153.446
R138 vss.n1651 vss.t4 153.446
R139 vss.n1525 vss.t87 153.446
R140 vss.n1540 vss.t48 153.446
R141 vss.n1771 vss.t131 153.446
R142 vss.n2223 vss.t8 153.446
R143 vss.n2531 vss.t98 153.446
R144 vss.n2550 vss.t7 153.446
R145 vss.n2495 vss.t33 153.446
R146 vss.n2669 vss.t66 153.446
R147 vss.n2342 vss.t113 153.446
R148 vss.n2745 vss.t121 153.446
R149 vss.n264 vss.t120 153.446
R150 vss.n3185 vss.n119 149.526
R151 vss.n2945 vss.t1 147.113
R152 vss.n2005 vss.t135 147.113
R153 vss.n3027 vss.t10 144.97
R154 vss.n566 vss.t94 133.739
R155 vss.n2112 vss.n2111 133.739
R156 vss.n2023 vss.n2022 133.739
R157 vss.n1172 vss.t122 133.739
R158 vss.t137 vss 132.565
R159 vss.n3034 vss.t108 126.924
R160 vss.n3127 vss.t70 124.103
R161 vss.n3024 vss.t9 124.103
R162 vss.n3015 vss.t137 124.103
R163 vss.n2942 vss 120.365
R164 vss.n3121 vss.t20 115.641
R165 vss.t84 vss.t44 114.87
R166 vss.t111 vss.t31 114.772
R167 vss.t103 vss.t34 114.772
R168 vss.n846 vss.t67 114.772
R169 vss.n1823 vss.t132 114.772
R170 vss.n2266 vss.t77 114.772
R171 vss.n2818 vss.t129 114.772
R172 vss.n3044 vss.n3043 113.207
R173 vss.n3015 vss.t106 112.822
R174 vss.t64 vss.t54 112.758
R175 vss.n968 vss.t74 112.278
R176 vss.n726 vss.t76 112.278
R177 vss.n369 vss.t75 112.278
R178 vss.n2408 vss.t3 112.278
R179 vss.n3276 vss.t52 111.924
R180 vss.n3227 vss.n3226 110.538
R181 vss.n2909 vss.t81 107.195
R182 vss.n611 vss.t57 107.195
R183 vss.n3225 vss.t125 107.195
R184 vss.n3191 vss.t89 107.195
R185 vss.n1141 vss.t97 107.195
R186 vss.n2937 vss.t2 107.195
R187 vss.n1998 vss.t136 107.195
R188 vss.n1177 vss.t123 107.195
R189 vss.n2123 vss.t6 107.195
R190 vss.n559 vss.t95 107.195
R191 vss.n3092 vss.t86 107.18
R192 vss.n3087 vss.n3086 106.038
R193 vss.n3126 vss.n3125 105.3
R194 vss.n3250 vss.t79 104.666
R195 vss.n3112 vss.t22 104.359
R196 vss.n3009 vss.n3008 103.942
R197 vss.n3111 vss.n3110 103.942
R198 vss.n2110 vss.t105 103.544
R199 vss.t28 vss.n2024 102.297
R200 vss.n3312 vss.n3311 97.3398
R201 vss.n3105 vss.t11 95.8979
R202 vss.n2894 vss.n2891 93.0283
R203 vss.n2021 vss.n602 93.0283
R204 vss.n1199 vss.n1126 87.5561
R205 vss.n598 vss.n597 87.5561
R206 vss.n3038 vss.t82 87.4364
R207 vss.n1240 vss.n1239 87.4012
R208 vss.n1950 vss.n1949 87.3268
R209 vss.n2052 vss.n2051 87.3268
R210 vss.n2845 vss.n2844 85.7944
R211 vss.n3097 vss.t127 84.6159
R212 vss.n1148 vss.t42 82.4069
R213 vss.n3297 vss.t134 77.4275
R214 vss.n773 vss.t45 77.3934
R215 vss.n773 vss.t43 77.3934
R216 vss.n2061 vss.t102 77.3934
R217 vss.n2061 vss.t101 77.3934
R218 vss.n638 vss.t30 77.3934
R219 vss.n638 vss.t26 77.3934
R220 vss.n3254 vss.t53 77.3934
R221 vss.n3254 vss.t49 77.3934
R222 vss.n56 vss.t16 77.2767
R223 vss.n3312 vss.t63 76.9003
R224 vss.n5 vss.t73 76.7239
R225 vss.n1147 vss.n1143 76.6116
R226 vss.n567 vss.n563 76.6116
R227 vss.n3188 vss.n3187 76.5234
R228 vss.n3045 vss.t116 76.1543
R229 vss.n3043 vss.t117 75.7148
R230 vss.n3314 vss.t59 75.7036
R231 vss.n2946 vss.n2941 71.1394
R232 vss.n2006 vss.n2002 71.1394
R233 vss.n1169 vss.t84 68.6725
R234 vss.t139 vss.n1240 66.1753
R235 vss.n1949 vss.t110 66.119
R236 vss.n2051 vss.t68 66.119
R237 vss.n2844 vss.t119 64.9587
R238 vss.t54 vss.n3183 57.605
R239 vss.n1975 vss.t99 57.3864
R240 vss.t126 vss.n845 57.3864
R241 vss.t0 vss.n2265 57.3864
R242 vss.n119 vss.t91 56.3793
R243 vss.t69 vss.n1822 56.1389
R244 vss.t130 vss.n2817 56.1389
R245 vss.n3110 vss.t12 54.2862
R246 vss.n3125 vss.t21 54.2862
R247 vss.n2944 vss.n2943 53.4959
R248 vss.n2004 vss.n2003 53.4959
R249 vss.n1877 vss.n1876 51.1488
R250 vss.n498 vss.n497 51.1488
R251 vss.n2842 vss.n2841 51.1488
R252 vss.n3081 vss.t24 50.7697
R253 vss.n1149 vss.t40 47.4466
R254 vss.n1969 vss.t100 47.4062
R255 vss.n2037 vss.t29 47.4062
R256 vss.n3311 vss.t62 47.1434
R257 vss.n3311 vss.t61 47.1434
R258 vss.n94 vss.t14 47.1434
R259 vss.n94 vss.t18 47.1434
R260 vss.n2864 vss.t92 46.5743
R261 vss.n3014 vss 45.1287
R262 vss.n648 vss.t112 43.7547
R263 vss.n784 vss.t85 43.7547
R264 vss.n2072 vss.t35 43.7547
R265 vss.n3269 vss.t65 43.7547
R266 vss.n1149 vss.t41 42.4523
R267 vss.n2037 vss.t27 42.4162
R268 vss.n3077 vss.t109 42.3082
R269 vss.n129 vss.t93 41.4448
R270 vss.n1948 vss.t104 41.4448
R271 vss.n1218 vss.t46 41.4448
R272 vss.n2137 vss.t32 41.4448
R273 vss.n3086 vss.t25 41.4291
R274 vss.n565 vss.n564 40.1221
R275 vss.n1174 vss.n1173 40.1221
R276 vss.t67 vss.t126 38.6736
R277 vss.t132 vss.t69 38.6736
R278 vss.n1877 vss.n1873 38.6736
R279 vss.t77 vss.t0 38.6736
R280 vss.t129 vss.t130 38.6736
R281 vss.n2819 vss.n2818 38.6736
R282 vss.n2841 vss.n170 38.6736
R283 vss.n3008 vss.t107 38.5719
R284 vss.n3008 vss.t138 38.5719
R285 vss.n3043 vss.t37 38.5719
R286 vss.n3086 vss.t39 38.5719
R287 vss.t44 vss.n1148 37.4579
R288 vss.n3183 vss.n3182 36.7693
R289 vss.n3088 vss.t38 33.8467
R290 vss.n3187 vss 32.7071
R291 vss.n96 vss.n94 30.6282
R292 vss.n3296 vss.n3250 26.3593
R293 vss.n2965 vss.n2961 25.977
R294 vss.n3110 vss.t23 25.9346
R295 vss.n3125 vss.t71 25.9346
R296 vss.n3184 vss.t64 25.7387
R297 vss.n3058 vss.t128 25.3851
R298 vss.n3049 vss.t36 25.3851
R299 vss.n1127 vss.n1125 23.9034
R300 vss.t60 vss.t78 23.0875
R301 vss.t58 vss.t60 23.0875
R302 vss.n1198 vss.n1197 22.6545
R303 vss.n2963 vss.n2962 22.5646
R304 vss.n2941 vss.n2940 21.8894
R305 vss.n2002 vss.n2001 21.8894
R306 vss.n121 vss.t50 20.8362
R307 vss vss.n1177 20.1079
R308 vss.n559 vss 20.1079
R309 vss.n467 vss.n466 17.6397
R310 vss.n2024 vss.t31 17.4658
R311 vss.n1175 vss.n1147 16.4172
R312 vss.n563 vss.n562 16.4172
R313 vss.n2110 vss.t103 16.2182
R314 vss.n1077 vss.n1076 16.2182
R315 vss.n864 vss.n863 16.2182
R316 vss.n1062 vss.n1061 16.2182
R317 vss.n2216 vss.n2215 16.2182
R318 vss.n2203 vss.n2202 16.2182
R319 vss.n2524 vss.n2523 16.2182
R320 vss.t50 vss.n120 15.9336
R321 vss.n3068 vss.t114 14.1031
R322 vss.n2077 vss 14.0497
R323 vss.n2112 vss.n600 13.3744
R324 vss.n1203 vss.n1201 13.3744
R325 vss.n2909 vss.n2906 13.1351
R326 vss.n1141 vss.n1127 13.1351
R327 vss.n612 vss.n611 13.1351
R328 vss.n1228 vss 12.4783
R329 vss.n3276 vss.n3275 11.427
R330 vss.n3277 vss.n3276 10.5417
R331 vss.n2947 vss.n2946 9.3005
R332 vss.n2946 vss.n2945 9.3005
R333 vss.n2934 vss.n2933 9.3005
R334 vss.n2932 vss.n2931 9.3005
R335 vss.n1197 vss.n1196 9.3005
R336 vss.n1125 vss.n1123 9.3005
R337 vss.n1194 vss.n1144 9.3005
R338 vss.n1193 vss.n1192 9.3005
R339 vss.n576 vss.n575 9.3005
R340 vss.n574 vss.n573 9.3005
R341 vss.n2115 vss.n2113 9.3005
R342 vss.n2113 vss.n2112 9.3005
R343 vss.n568 vss.n567 9.3005
R344 vss.n567 vss.n566 9.3005
R345 vss.n2007 vss.n2006 9.3005
R346 vss.n2006 vss.n2005 9.3005
R347 vss.n2014 vss.n2013 9.3005
R348 vss.n2012 vss.n2011 9.3005
R349 vss.n1205 vss.n1204 9.3005
R350 vss.n1204 vss.n1203 9.3005
R351 vss.n1190 vss.n1189 9.3005
R352 vss.n1190 vss.n1143 9.3005
R353 vss.n1172 vss.n1143 9.3005
R354 vss.n2253 vss.n2252 9.15497
R355 vss.n537 vss.n536 9.15497
R356 vss.n2046 vss.n2045 9.15497
R357 vss.n2045 vss.n2044 9.15497
R358 vss.n2054 vss.n2053 9.15497
R359 vss.n2053 vss.n2052 9.15497
R360 vss.n2108 vss.n2107 9.15497
R361 vss.n2109 vss.n2108 9.15497
R362 vss.n2039 vss.n2038 9.15497
R363 vss.n2038 vss.n2037 9.15497
R364 vss.n1959 vss.n1958 9.15497
R365 vss.n1958 vss.n1957 9.15497
R366 vss.n1971 vss.n1970 9.15497
R367 vss.n1970 vss.n1969 9.15497
R368 vss.n1977 vss.n1976 9.15497
R369 vss.n1976 vss.n1975 9.15497
R370 vss.n1952 vss.n1951 9.15497
R371 vss.n1951 vss.n1950 9.15497
R372 vss.n1857 vss.n1856 9.15497
R373 vss.n1887 vss.n1886 9.15497
R374 vss.n1298 vss.n1297 9.15497
R375 vss.n1297 vss.n1296 9.15497
R376 vss.n1305 vss.n1304 9.15497
R377 vss.n1304 vss.n1303 9.15497
R378 vss.n1632 vss.n1631 9.15497
R379 vss.n1631 vss.n1630 9.15497
R380 vss.n1642 vss.n1641 9.15497
R381 vss.n1641 vss.n1640 9.15497
R382 vss.n1635 vss.n1634 9.15497
R383 vss.n1634 vss.n1633 9.15497
R384 vss.n1653 vss.n1652 9.15497
R385 vss.n1652 vss.n1651 9.15497
R386 vss.n700 vss.n699 9.15497
R387 vss.n699 vss.n698 9.15497
R388 vss.n707 vss.n706 9.15497
R389 vss.n706 vss.n705 9.15497
R390 vss.n714 vss.n713 9.15497
R391 vss.n713 vss.n712 9.15497
R392 vss.n970 vss.n969 9.15497
R393 vss.n969 vss.n968 9.15497
R394 vss.n1001 vss.n1000 9.15497
R395 vss.n1000 vss.n999 9.15497
R396 vss.n906 vss.n905 9.15497
R397 vss.n905 vss.n904 9.15497
R398 vss.n918 vss.n917 9.15497
R399 vss.n917 vss.n916 9.15497
R400 vss.n1009 vss.n1008 9.15497
R401 vss.n1008 vss.n1007 9.15497
R402 vss.n866 vss.n865 9.15497
R403 vss.n865 vss.n864 9.15497
R404 vss.n1064 vss.n1063 9.15497
R405 vss.n1063 vss.n1062 9.15497
R406 vss.n1025 vss.n1024 9.15497
R407 vss.n1024 vss.n1023 9.15497
R408 vss.n1075 vss.n1074 9.15497
R409 vss.n1076 vss.n1075 9.15497
R410 vss.n1817 vss.n1816 9.15497
R411 vss.n1825 vss.n1824 9.15497
R412 vss.n1824 vss.n1823 9.15497
R413 vss.n1759 vss.n1758 9.15497
R414 vss.n1758 vss.n1757 9.15497
R415 vss.n1766 vss.n1765 9.15497
R416 vss.n1765 vss.n1764 9.15497
R417 vss.n1773 vss.n1772 9.15497
R418 vss.n1772 vss.n1771 9.15497
R419 vss.n1712 vss.n1711 9.15497
R420 vss.n1711 vss.n1710 9.15497
R421 vss.n1079 vss.n1078 9.15497
R422 vss.n1078 vss.n1077 9.15497
R423 vss.n862 vss.n861 9.15497
R424 vss.n863 vss.n862 9.15497
R425 vss.n1060 vss.n1059 9.15497
R426 vss.n1061 vss.n1060 9.15497
R427 vss.n1086 vss.n1085 9.15497
R428 vss.n1085 vss.n1084 9.15497
R429 vss.n840 vss.n839 9.15497
R430 vss.n839 vss.n838 9.15497
R431 vss.n848 vss.n847 9.15497
R432 vss.n847 vss.n846 9.15497
R433 vss.n1533 vss.n1532 9.15497
R434 vss.n1532 vss.n1531 9.15497
R435 vss.n1576 vss.n1575 9.15497
R436 vss.n1575 vss.n1574 9.15497
R437 vss.n1559 vss.n1558 9.15497
R438 vss.n1558 vss.n1557 9.15497
R439 vss.n1542 vss.n1541 9.15497
R440 vss.n1541 vss.n1540 9.15497
R441 vss.n1513 vss.n1512 9.15497
R442 vss.n1512 vss.n1511 9.15497
R443 vss.n1520 vss.n1519 9.15497
R444 vss.n1519 vss.n1518 9.15497
R445 vss.n1527 vss.n1526 9.15497
R446 vss.n1526 vss.n1525 9.15497
R447 vss.n1506 vss.n1505 9.15497
R448 vss.n1505 vss.n1504 9.15497
R449 vss.n1400 vss.n1399 9.15497
R450 vss.n1399 vss.n1398 9.15497
R451 vss.n1427 vss.n1426 9.15497
R452 vss.n1426 vss.n1425 9.15497
R453 vss.n728 vss.n727 9.15497
R454 vss.n727 vss.n726 9.15497
R455 vss.n1408 vss.n1407 9.15497
R456 vss.n1407 vss.n1406 9.15497
R457 vss.n1380 vss.n1379 9.15497
R458 vss.n1379 vss.n1378 9.15497
R459 vss.n1387 vss.n1386 9.15497
R460 vss.n1386 vss.n1385 9.15497
R461 vss.n1394 vss.n1393 9.15497
R462 vss.n1393 vss.n1392 9.15497
R463 vss.n1373 vss.n1372 9.15497
R464 vss.n1372 vss.n1371 9.15497
R465 vss.n1879 vss.n1878 9.15497
R466 vss.n1878 vss.n1877 9.15497
R467 vss.n1898 vss.n1897 9.15497
R468 vss.n1897 vss.n1896 9.15497
R469 vss.n1263 vss.n1262 9.15497
R470 vss.n1262 vss.n1261 9.15497
R471 vss.n1244 vss.n1243 9.15497
R472 vss.n1243 vss.n1242 9.15497
R473 vss.n1151 vss.n1150 9.15497
R474 vss.n1150 vss.n1149 9.15497
R475 vss.n1156 vss.n1155 9.15497
R476 vss.n1155 vss.n1154 9.15497
R477 vss.n1238 vss.n1237 9.15497
R478 vss.n1239 vss.n1238 9.15497
R479 vss.n1167 vss.n1166 9.15497
R480 vss.n1168 vss.n1167 9.15497
R481 vss.n833 vss.n832 9.15497
R482 vss.n832 vss.n831 9.15497
R483 vss.n826 vss.n825 9.15497
R484 vss.n825 vss.n824 9.15497
R485 vss.n2854 vss.n2853 9.15497
R486 vss.n2853 vss.n2852 9.15497
R487 vss.n2866 vss.n2865 9.15497
R488 vss.n2865 vss.n2864 9.15497
R489 vss.n2871 vss.n2870 9.15497
R490 vss.n2870 vss.n119 9.15497
R491 vss.n2847 vss.n2846 9.15497
R492 vss.n2846 vss.n2845 9.15497
R493 vss.n2732 vss.n2731 9.15497
R494 vss.n2731 vss.n2730 9.15497
R495 vss.n2736 vss.n2735 9.15497
R496 vss.n2735 vss.n2734 9.15497
R497 vss.n2794 vss.n2793 9.15497
R498 vss.n2793 vss.n2792 9.15497
R499 vss.n2747 vss.n2746 9.15497
R500 vss.n2746 vss.n2745 9.15497
R501 vss.n2372 vss.n2371 9.15497
R502 vss.n2371 vss.n2370 9.15497
R503 vss.n2337 vss.n2336 9.15497
R504 vss.n2336 vss.n2335 9.15497
R505 vss.n2344 vss.n2343 9.15497
R506 vss.n2343 vss.n2342 9.15497
R507 vss.n2392 vss.n2391 9.15497
R508 vss.n2391 vss.n2390 9.15497
R509 vss.n2451 vss.n2450 9.15497
R510 vss.n2450 vss.n2449 9.15497
R511 vss.n2427 vss.n2426 9.15497
R512 vss.n2426 vss.n2425 9.15497
R513 vss.n2410 vss.n2409 9.15497
R514 vss.n2409 vss.n2408 9.15497
R515 vss.n2459 vss.n2458 9.15497
R516 vss.n2458 vss.n2457 9.15497
R517 vss.n2490 vss.n2489 9.15497
R518 vss.n2489 vss.n2488 9.15497
R519 vss.n2497 vss.n2496 9.15497
R520 vss.n2496 vss.n2495 9.15497
R521 vss.n2476 vss.n2475 9.15497
R522 vss.n2475 vss.n2474 9.15497
R523 vss.n2483 vss.n2482 9.15497
R524 vss.n2482 vss.n2481 9.15497
R525 vss.n2218 vss.n2217 9.15497
R526 vss.n2217 vss.n2216 9.15497
R527 vss.n2201 vss.n2200 9.15497
R528 vss.n2202 vss.n2201 9.15497
R529 vss.n2522 vss.n2521 9.15497
R530 vss.n2523 vss.n2522 9.15497
R531 vss.n2225 vss.n2224 9.15497
R532 vss.n2224 vss.n2223 9.15497
R533 vss.n2260 vss.n2259 9.15497
R534 vss.n2259 vss.n2258 9.15497
R535 vss.n2268 vss.n2267 9.15497
R536 vss.n2267 vss.n2266 9.15497
R537 vss.n500 vss.n499 9.15497
R538 vss.n499 vss.n498 9.15497
R539 vss.n507 vss.n506 9.15497
R540 vss.n506 vss.n505 9.15497
R541 vss.n2655 vss.n2654 9.15497
R542 vss.n2654 vss.n2653 9.15497
R543 vss.n2660 vss.n2659 9.15497
R544 vss.n2659 vss.n2658 9.15497
R545 vss.n2696 vss.n2695 9.15497
R546 vss.n2695 vss.n2694 9.15497
R547 vss.n2671 vss.n2670 9.15497
R548 vss.n2670 vss.n2669 9.15497
R549 vss.n378 vss.n377 9.15497
R550 vss.n377 vss.n376 9.15497
R551 vss.n385 vss.n384 9.15497
R552 vss.n384 vss.n383 9.15497
R553 vss.n392 vss.n391 9.15497
R554 vss.n391 vss.n390 9.15497
R555 vss.n371 vss.n370 9.15497
R556 vss.n370 vss.n369 9.15497
R557 vss.n2544 vss.n2543 9.15497
R558 vss.n2543 vss.n2542 9.15497
R559 vss.n2579 vss.n2578 9.15497
R560 vss.n2578 vss.n2577 9.15497
R561 vss.n2595 vss.n2594 9.15497
R562 vss.n2594 vss.n2593 9.15497
R563 vss.n2552 vss.n2551 9.15497
R564 vss.n2551 vss.n2550 9.15497
R565 vss.n2205 vss.n2204 9.15497
R566 vss.n2204 vss.n2203 9.15497
R567 vss.n2526 vss.n2525 9.15497
R568 vss.n2525 vss.n2524 9.15497
R569 vss.n2533 vss.n2532 9.15497
R570 vss.n2532 vss.n2531 9.15497
R571 vss.n2214 vss.n2213 9.15497
R572 vss.n2215 vss.n2214 9.15497
R573 vss.n271 vss.n270 9.15497
R574 vss.n270 vss.n170 9.15497
R575 vss.n290 vss.n289 9.15497
R576 vss.n252 vss.n251 9.15497
R577 vss.n251 vss.n250 9.15497
R578 vss.n259 vss.n258 9.15497
R579 vss.n258 vss.n257 9.15497
R580 vss.n266 vss.n265 9.15497
R581 vss.n265 vss.n264 9.15497
R582 vss.n245 vss.n244 9.15497
R583 vss.n244 vss.n243 9.15497
R584 vss.n280 vss.n279 9.15497
R585 vss.n2828 vss.n2827 9.15497
R586 vss.n2821 vss.n2820 9.15497
R587 vss.n2820 vss.n2819 9.15497
R588 vss.n2840 vss.n2839 9.15497
R589 vss.n2841 vss.n2840 9.15497
R590 vss.n2895 vss.n2894 9.01392
R591 vss.n2021 vss.n2020 9.01392
R592 vss.n2022 vss.n2021 9.01392
R593 vss.n2894 vss.n2893 9.01392
R594 vss.n1856 vss.n1855 8.48574
R595 vss.n1886 vss.n1885 8.48574
R596 vss.n279 vss.n278 8.48574
R597 vss.n2827 vss.n2826 8.48523
R598 vss.n2252 vss.n2251 8.48521
R599 vss.n3065 vss.n3062 8.47109
R600 vss.n1141 vss.n1140 8.11658
R601 vss.n2124 vss.n2123 8.11658
R602 vss vss.n2909 7.93155
R603 vss.n611 vss 7.93155
R604 vss.n1177 vss.n1176 7.90638
R605 vss.n560 vss.n559 7.90638
R606 vss.n3228 vss.n3225 7.71815
R607 vss.n3047 vss.n3044 7.71815
R608 vss.n2938 vss.n2937 7.52991
R609 vss.n1999 vss.n1998 7.52991
R610 vss.n1242 vss.n1241 7.49199
R611 vss.n3090 vss.n3087 7.34168
R612 vss.n3313 vss.n3312 6.28259
R613 vss.n1876 vss.n1875 6.2381
R614 vss.n2843 vss.n2842 6.12863
R615 vss.n3072 vss.t83 5.64153
R616 vss.n1204 vss.n1126 5.47272
R617 vss.n2113 vss.n598 5.47272
R618 vss.n3192 vss.n3191 5.45932
R619 vss.n2883 vss 5.28181
R620 vss.n1132 vss.n1116 5.18083
R621 vss.n497 vss.n496 4.99058
R622 vss.n120 vss.n118 4.90301
R623 vss vss.n1115 4.7265
R624 vss.n114 vss.n113 4.6505
R625 vss.n3219 vss.n3218 4.6505
R626 vss.n3235 vss.n3234 4.6505
R627 vss.n3229 vss.n3228 4.6505
R628 vss.n3012 vss.n3011 4.6505
R629 vss.n3022 vss.n3021 4.6505
R630 vss.n3018 vss.n3017 4.6505
R631 vss.n3028 vss.n3027 4.6505
R632 vss.n2906 vss.n2905 4.6505
R633 vss.n2961 vss.n2960 4.6505
R634 vss.n3130 vss.n3129 4.6505
R635 vss.n3124 vss.n3123 4.6505
R636 vss.n3115 vss.n3114 4.6505
R637 vss.n3108 vss.n3107 4.6505
R638 vss.n3100 vss.n3099 4.6505
R639 vss.n3091 vss.n3090 4.6505
R640 vss.n3080 vss.n3079 4.6505
R641 vss.n3071 vss.n3070 4.6505
R642 vss.n3061 vss.n3060 4.6505
R643 vss.n3052 vss.n3051 4.6505
R644 vss.n3041 vss.n3040 4.6505
R645 vss.n3032 vss.n3031 4.6505
R646 vss.n3037 vss.n3036 4.6505
R647 vss.n3048 vss.n3047 4.6505
R648 vss.n3056 vss.n3055 4.6505
R649 vss.n3066 vss.n3065 4.6505
R650 vss.n3075 vss.n3074 4.6505
R651 vss.n3084 vss.n3083 4.6505
R652 vss.n3095 vss.n3094 4.6505
R653 vss.n3104 vss.n3103 4.6505
R654 vss.n3119 vss.n3118 4.6505
R655 vss.n2966 vss.n2965 4.6505
R656 vss.n1129 vss.n1127 4.6505
R657 vss.n2120 vss.n2119 4.6505
R658 vss.n613 vss.n612 4.6505
R659 vss.n3302 vss.n3301 4.6505
R660 vss.n3316 vss.n3315 4.6505
R661 vss.n3300 vss.n3299 4.6505
R662 vss.n3298 vss.n3297 4.6505
R663 vss.n3281 vss.n3277 4.6505
R664 vss.n3280 vss.n3279 4.6505
R665 vss.n3294 vss.n3250 4.6505
R666 vss.n3207 vss.n3206 4.5005
R667 vss.n3221 vss.n3220 4.5005
R668 vss.n3193 vss.n3192 4.5005
R669 vss vss.n2902 4.5005
R670 vss.n2949 vss.n2948 4.5005
R671 vss.n1179 vss.n1178 4.5005
R672 vss.n1186 vss.n1145 4.5005
R673 vss.n1191 vss.n1145 4.5005
R674 vss.n1139 vss.n1138 4.5005
R675 vss.n1195 vss.n1120 4.5005
R676 vss.n1207 vss.n1206 4.5005
R677 vss.n1128 vss.n1122 4.5005
R678 vss.n571 vss.n570 4.5005
R679 vss.n2009 vss.n2008 4.5005
R680 vss vss.n608 4.5005
R681 vss.n2948 vss.n2936 3.76521
R682 vss.n1192 vss.n1191 3.76521
R683 vss.n570 vss.n569 3.76521
R684 vss.n2008 vss.n1997 3.76521
R685 vss.n3315 vss.n3314 3.50366
R686 vss.n1181 vss.n1179 3.45606
R687 vss.n2895 vss.n2890 3.45447
R688 vss.n1205 vss.n1125 3.45447
R689 vss.n2115 vss.n2114 3.45447
R690 vss.n2020 vss.n2019 3.45447
R691 vss.n1186 vss.n1185 3.42401
R692 vss.n1138 vss.n1137 3.42259
R693 vss.n1564 vss 3.42087
R694 vss.n1120 vss.n1117 3.42064
R695 vss.n1122 vss.n1119 3.41895
R696 vss.n1184 vss.n1183 3.4105
R697 vss.n1133 vss.n1116 3.4105
R698 vss.n1136 vss.n1135 3.4105
R699 vss.n1182 vss.n1180 3.4105
R700 vss.n1210 vss.n1209 3.4105
R701 vss.n1225 vss.n1224 3.4105
R702 vss.n2939 vss.n2938 3.38874
R703 vss.n1190 vss.n1146 3.38874
R704 vss.n568 vss.n561 3.38874
R705 vss.n2000 vss.n1999 3.38874
R706 vss.n2896 vss.n2889 3.25129
R707 vss.n1198 vss.n1124 3.25129
R708 vss.n596 vss.n595 3.25129
R709 vss.n2018 vss.n603 3.25129
R710 vss.n3190 vss.n3189 3.19788
R711 vss.n3027 vss.n3026 3.10907
R712 vss.n3205 vss.n3204 3.1005
R713 vss.n253 vss.n252 3.03311
R714 vss.n285 vss.n271 3.03311
R715 vss.n2855 vss.n2854 3.03311
R716 vss.n2897 vss.n2896 3.03311
R717 vss.n1892 vss.n1879 3.03311
R718 vss.n1760 vss.n1759 3.03311
R719 vss.n1381 vss.n1380 3.03311
R720 vss.n1402 vss.n1400 3.03311
R721 vss.n1514 vss.n1513 3.03311
R722 vss.n1536 vss.n1533 3.03311
R723 vss.n1264 vss.n1263 3.03311
R724 vss.n1161 vss.n1151 3.03311
R725 vss.n834 vss.n833 3.03311
R726 vss.n1080 vss.n1079 3.03311
R727 vss.n1069 vss.n866 3.03311
R728 vss.n1003 vss.n1001 3.03311
R729 vss.n701 vss.n700 3.03311
R730 vss.n1647 vss.n1632 3.03311
R731 vss.n1960 vss.n1959 3.03311
R732 vss.n2107 vss.n2106 3.03311
R733 vss.n2219 vss.n2218 3.03311
R734 vss.n2246 vss.n2245 3.03311
R735 vss.n2254 vss.n2253 3.03311
R736 vss.n538 vss.n537 3.03311
R737 vss.n468 vss.n467 3.03311
R738 vss.n2208 vss.n2205 3.03311
R739 vss.n2546 vss.n2544 3.03311
R740 vss.n379 vss.n378 3.03311
R741 vss.n2665 vss.n2655 3.03311
R742 vss.n2477 vss.n2476 3.03311
R743 vss.n2453 vss.n2451 3.03311
R744 vss.n2373 vss.n2372 3.03311
R745 vss.n2741 vss.n2732 3.03311
R746 vss.n2047 vss.n2046 3.03311
R747 vss.n2055 vss.n2054 3.03311
R748 vss.n2040 vss.n2039 3.03311
R749 vss.n1972 vss.n1971 3.03311
R750 vss.n1978 vss.n1977 3.03311
R751 vss.n1953 vss.n1952 3.03311
R752 vss.n2018 vss.n2017 3.03311
R753 vss.n1859 vss.n1857 3.03311
R754 vss.n1806 vss.n1805 3.03311
R755 vss.n1888 vss.n1887 3.03311
R756 vss.n1881 vss.n1880 3.03311
R757 vss.n1299 vss.n1298 3.03311
R758 vss.n1306 vss.n1305 3.03311
R759 vss.n1643 vss.n1642 3.03311
R760 vss.n1636 vss.n1635 3.03311
R761 vss.n1654 vss.n1653 3.03311
R762 vss.n708 vss.n707 3.03311
R763 vss.n715 vss.n714 3.03311
R764 vss.n971 vss.n970 3.03311
R765 vss.n907 vss.n906 3.03311
R766 vss.n919 vss.n918 3.03311
R767 vss.n1010 vss.n1009 3.03311
R768 vss.n1065 vss.n1064 3.03311
R769 vss.n1026 vss.n1025 3.03311
R770 vss.n1074 vss.n1073 3.03311
R771 vss.n1818 vss.n1817 3.03311
R772 vss.n1826 vss.n1825 3.03311
R773 vss.n1767 vss.n1766 3.03311
R774 vss.n1774 vss.n1773 3.03311
R775 vss.n1713 vss.n1712 3.03311
R776 vss.n861 vss.n860 3.03311
R777 vss.n1059 vss.n1058 3.03311
R778 vss.n1087 vss.n1086 3.03311
R779 vss.n841 vss.n840 3.03311
R780 vss.n849 vss.n848 3.03311
R781 vss.n1577 vss.n1576 3.03311
R782 vss.n1560 vss.n1559 3.03311
R783 vss.n1543 vss.n1542 3.03311
R784 vss.n1521 vss.n1520 3.03311
R785 vss.n1528 vss.n1527 3.03311
R786 vss.n1507 vss.n1506 3.03311
R787 vss.n1428 vss.n1427 3.03311
R788 vss.n729 vss.n728 3.03311
R789 vss.n1409 vss.n1408 3.03311
R790 vss.n1388 vss.n1387 3.03311
R791 vss.n1395 vss.n1394 3.03311
R792 vss.n1374 vss.n1373 3.03311
R793 vss.n1899 vss.n1898 3.03311
R794 vss.n1245 vss.n1244 3.03311
R795 vss.n1157 vss.n1156 3.03311
R796 vss.n1237 vss.n1236 3.03311
R797 vss.n1166 vss.n1165 3.03311
R798 vss.n827 vss.n826 3.03311
R799 vss.n2867 vss.n2866 3.03311
R800 vss.n2872 vss.n2871 3.03311
R801 vss.n2848 vss.n2847 3.03311
R802 vss.n2737 vss.n2736 3.03311
R803 vss.n2795 vss.n2794 3.03311
R804 vss.n2748 vss.n2747 3.03311
R805 vss.n2338 vss.n2337 3.03311
R806 vss.n2345 vss.n2344 3.03311
R807 vss.n2393 vss.n2392 3.03311
R808 vss.n2428 vss.n2427 3.03311
R809 vss.n2411 vss.n2410 3.03311
R810 vss.n2460 vss.n2459 3.03311
R811 vss.n2491 vss.n2490 3.03311
R812 vss.n2498 vss.n2497 3.03311
R813 vss.n2484 vss.n2483 3.03311
R814 vss.n2200 vss.n2199 3.03311
R815 vss.n2521 vss.n2520 3.03311
R816 vss.n2226 vss.n2225 3.03311
R817 vss.n2261 vss.n2260 3.03311
R818 vss.n2269 vss.n2268 3.03311
R819 vss.n501 vss.n500 3.03311
R820 vss.n508 vss.n507 3.03311
R821 vss.n2661 vss.n2660 3.03311
R822 vss.n2697 vss.n2696 3.03311
R823 vss.n2672 vss.n2671 3.03311
R824 vss.n386 vss.n385 3.03311
R825 vss.n393 vss.n392 3.03311
R826 vss.n372 vss.n371 3.03311
R827 vss.n2580 vss.n2579 3.03311
R828 vss.n2596 vss.n2595 3.03311
R829 vss.n2553 vss.n2552 3.03311
R830 vss.n2527 vss.n2526 3.03311
R831 vss.n2534 vss.n2533 3.03311
R832 vss.n2213 vss.n2212 3.03311
R833 vss.n291 vss.n290 3.03311
R834 vss.n260 vss.n259 3.03311
R835 vss.n267 vss.n266 3.03311
R836 vss.n246 vss.n245 3.03311
R837 vss.n281 vss.n280 3.03311
R838 vss.n273 vss.n272 3.03311
R839 vss.n2834 vss.n2828 3.03311
R840 vss.n2822 vss.n2821 3.03311
R841 vss.n2830 vss.n2829 3.03311
R842 vss.n2839 vss.n2838 3.03311
R843 vss.n2888 vss 3.01818
R844 vss.n2947 vss.n2939 3.01226
R845 vss.n1176 vss.n1146 3.01226
R846 vss.n561 vss.n560 3.01226
R847 vss.n2007 vss.n2000 3.01226
R848 vss.n3053 vss.t55 2.82101
R849 vss vss.n3014 2.82101
R850 vss vss.n2883 2.44479
R851 vss.n72 vss.n71 2.3255
R852 vss.n60 vss.n59 2.3255
R853 vss.n8 vss.n7 2.3255
R854 vss.n35 vss.n34 2.3255
R855 vss.n2116 vss.n2115 2.28739
R856 vss.n1206 vss.n1205 2.28739
R857 vss.n77 vss.n76 2.2505
R858 vss.n132 vss.n131 2.24031
R859 vss.n1946 vss.n684 2.24031
R860 vss.n3010 vss 2.04217
R861 vss.n3318 vss.n3317 2.01288
R862 vss.n133 vss 1.94963
R863 vss vss.n1945 1.94963
R864 vss.n3195 vss.n3194 1.94045
R865 vss.n3222 vss.n3213 1.94045
R866 vss.n3239 vss.n3237 1.94045
R867 vss.n3076 vss.n2986 1.94045
R868 vss.n3096 vss.n2978 1.94045
R869 vss.n3109 vss.n2974 1.94045
R870 vss.n3120 vss.n2970 1.94045
R871 vss.n3132 vss.n3131 1.94045
R872 vss.n3085 vss.n2982 1.94045
R873 vss.n3067 vss.n2990 1.94045
R874 vss.n3057 vss.n2994 1.94045
R875 vss.n3042 vss.n2998 1.94045
R876 vss.n3033 vss.n3002 1.94045
R877 vss.n3023 vss.n3006 1.94045
R878 vss.n3304 vss.n3303 1.94045
R879 vss.n3283 vss.n3282 1.94045
R880 vss.n3293 vss.n3292 1.94045
R881 vss.n81 vss.n80 1.94045
R882 vss.n100 vss.n99 1.94045
R883 vss.n17 vss.n13 1.94045
R884 vss.n43 vss.n40 1.94045
R885 vss.t133 vss.t58 1.92442
R886 vss.n2948 vss.n2947 1.50638
R887 vss.n1192 vss.n1144 1.50638
R888 vss.n2008 vss.n2007 1.50638
R889 vss.n2863 vss.n2862 1.35607
R890 vss.n2958 vss.n2957 1.35607
R891 vss.n2929 vss.n2928 1.35607
R892 vss.n1968 vss.n1967 1.35607
R893 vss.n557 vss.n556 1.35607
R894 vss.n1995 vss.n1994 1.35607
R895 vss.n2016 vss.n619 1.35607
R896 vss.n1861 vss.n1860 1.35607
R897 vss.n2875 vss.n2873 1.35607
R898 vss.n2913 vss.n2911 1.35607
R899 vss.n1718 vss.n1715 1.35607
R900 vss.n1582 vss.n1578 1.35607
R901 vss.n1563 vss.n1561 1.35607
R902 vss.n1432 vss.n1429 1.35607
R903 vss.n732 vss.n730 1.35607
R904 vss.n1250 vss.n1247 1.35607
R905 vss.n1268 vss.n1265 1.35607
R906 vss.n859 vss.n858 1.35607
R907 vss.n1057 vss.n1056 1.35607
R908 vss.n1188 vss.n1187 1.35607
R909 vss.n1208 vss.n1121 1.35607
R910 vss.n976 vss.n973 1.35607
R911 vss.n911 vss.n908 1.35607
R912 vss.n922 vss.n920 1.35607
R913 vss.n1981 vss.n1979 1.35607
R914 vss.n2105 vss.n2104 1.35607
R915 vss.n2198 vss.n2197 1.35607
R916 vss.n2519 vss.n2518 1.35607
R917 vss.n473 vss.n470 1.35607
R918 vss.n542 vss.n539 1.35607
R919 vss.n2700 vss.n2698 1.35607
R920 vss.n2584 vss.n2581 1.35607
R921 vss.n2599 vss.n2597 1.35607
R922 vss.n2798 vss.n2796 1.35607
R923 vss.n2398 vss.n2395 1.35607
R924 vss.n2379 vss.n2375 1.35607
R925 vss.n2432 vss.n2429 1.35607
R926 vss.n2414 vss.n2412 1.35607
R927 vss.n594 vss.n593 1.35607
R928 vss.n607 vss.n605 1.35607
R929 vss.n1808 vss.n1807 1.35607
R930 vss.n57 vss.n56 1.28807
R931 vss.n29 vss.n28 1.14394
R932 vss.n3317 vss.n3313 1.14386
R933 vss.n786 vss.n785 1.13981
R934 vss.n2074 vss.n2073 1.13981
R935 vss.n650 vss.n649 1.13981
R936 vss.n3271 vss.n3270 1.13981
R937 vss.n2097 vss.n2096 1.13729
R938 vss.n2059 vss.n2058 1.13729
R939 vss.n1209 vss.n1118 1.13717
R940 vss.n1921 vss.n1872 1.13685
R941 vss.n2362 vss.n2355 1.1368
R942 vss.n3242 vss.n3241 1.13462
R943 vss.n1214 vss.n1213 1.13462
R944 vss.n2145 vss.n2144 1.13462
R945 vss.n137 vss.n136 1.13462
R946 vss.n3211 vss.n3199 1.13451
R947 vss.n3198 vss.n3197 1.13451
R948 vss.n2878 vss.n2877 1.13388
R949 vss.n1232 vss.n1231 1.13388
R950 vss.n1054 vss.n1053 1.13388
R951 vss.n1321 vss.n1320 1.13388
R952 vss.n2099 vss.n2098 1.13388
R953 vss.n1191 vss.n1190 1.12991
R954 vss.n1197 vss.n1144 1.12991
R955 vss.n570 vss.n568 1.12991
R956 vss.n1131 vss.n1130 1.04225
R957 vss.n2128 vss.n2126 1.04225
R958 vss.n1221 vss.n1220 1.04145
R959 vss.n2140 vss.n2139 1.04145
R960 vss.n268 vss.n267 1.04008
R961 vss.n1775 vss.n1774 1.04008
R962 vss.n1396 vss.n1395 1.04008
R963 vss.n1529 vss.n1528 1.04008
R964 vss.n1307 vss.n1306 1.04008
R965 vss.n1236 vss.n1235 1.04008
R966 vss.n850 vss.n849 1.04008
R967 vss.n1026 vss.n1022 1.04008
R968 vss.n716 vss.n715 1.04008
R969 vss.n2056 vss.n2055 1.04008
R970 vss.n509 vss.n508 1.04008
R971 vss.n2535 vss.n2534 1.04008
R972 vss.n394 vss.n393 1.04008
R973 vss.n2499 vss.n2498 1.04008
R974 vss.n2346 vss.n2345 1.04008
R975 vss.n292 vss.n291 1.03985
R976 vss.n2848 vss.n168 1.03985
R977 vss.n1827 vss.n1826 1.03985
R978 vss.n1900 vss.n1899 1.03985
R979 vss.n1410 vss.n1409 1.03985
R980 vss.n1544 vss.n1543 1.03985
R981 vss.n1088 vss.n1087 1.03985
R982 vss.n1011 vss.n1010 1.03985
R983 vss.n1655 vss.n1654 1.03985
R984 vss.n1953 vss.n683 1.03985
R985 vss.n2227 vss.n2226 1.03985
R986 vss.n2270 vss.n2269 1.03985
R987 vss.n2554 vss.n2553 1.03985
R988 vss.n2673 vss.n2672 1.03985
R989 vss.n2461 vss.n2460 1.03985
R990 vss.n2749 vss.n2748 1.03985
R991 vss.n2822 vss.n2816 1.03984
R992 vss.n652 vss.n461 1.03084
R993 vss.n3324 vss.n104 0.969015
R994 vss.n3129 vss.n3126 0.941676
R995 vss.n3114 vss.n3111 0.941676
R996 vss.n1183 vss.n1181 0.871022
R997 vss.n1137 vss.n1136 0.870834
R998 vss.n135 vss.n133 0.853
R999 vss.n3213 vss.n3212 0.853
R1000 vss.n3196 vss.n3195 0.853
R1001 vss.n2928 vss.n2927 0.853
R1002 vss.n2957 vss.n2956 0.853
R1003 vss.n1921 vss.n1920 0.853
R1004 vss.n1719 vss.n1718 0.853
R1005 vss.n1473 vss.n1472 0.853
R1006 vss.n1565 vss.n1563 0.853
R1007 vss.n1585 vss.n1582 0.853
R1008 vss.n1599 vss.n1596 0.853
R1009 vss.n1604 vss.n1548 0.853
R1010 vss.n1609 vss.n1530 0.853
R1011 vss.n1495 vss.n1494 0.853
R1012 vss.n1484 vss.n1483 0.853
R1013 vss.n1610 vss.n1609 0.853
R1014 vss.n1604 vss.n1603 0.853
R1015 vss.n1600 vss.n1599 0.853
R1016 vss.n1586 vss.n1585 0.853
R1017 vss.n1566 vss.n1565 0.853
R1018 vss.n1251 vss.n1250 0.853
R1019 vss.n793 vss.n792 0.853
R1020 vss.n1102 vss.n851 0.853
R1021 vss.n815 vss.n814 0.853
R1022 vss.n804 vss.n803 0.853
R1023 vss.n1103 vss.n1102 0.853
R1024 vss.n778 vss.n776 0.853
R1025 vss.n1187 vss.n1115 0.853
R1026 vss.n1209 vss.n1208 0.853
R1027 vss.n1224 vss.n1222 0.853
R1028 vss.n1234 vss.n1233 0.853
R1029 vss.n1252 vss.n1251 0.853
R1030 vss.n1310 vss.n1308 0.853
R1031 vss.n1285 vss.n1282 0.853
R1032 vss.n1271 vss.n1268 0.853
R1033 vss.n1272 vss.n1271 0.853
R1034 vss.n1286 vss.n1285 0.853
R1035 vss.n1311 vss.n1310 0.853
R1036 vss.n1015 vss.n1014 0.853
R1037 vss.n960 vss.n957 0.853
R1038 vss.n979 vss.n976 0.853
R1039 vss.n984 vss.n922 0.853
R1040 vss.n989 vss.n911 0.853
R1041 vss.n994 vss.n898 0.853
R1042 vss.n984 vss.n983 0.853
R1043 vss.n980 vss.n979 0.853
R1044 vss.n961 vss.n960 0.853
R1045 vss.n1021 vss.n1020 0.853
R1046 vss.n889 vss.n888 0.853
R1047 vss.n879 vss.n878 0.853
R1048 vss.n1319 vss.n1318 0.853
R1049 vss.n1056 vss.n1055 0.853
R1050 vss.n1097 vss.n1096 0.853
R1051 vss.n1465 vss.n732 0.853
R1052 vss.n1436 vss.n1432 0.853
R1053 vss.n1441 vss.n1419 0.853
R1054 vss.n1446 vss.n1413 0.853
R1055 vss.n1451 vss.n1397 0.853
R1056 vss.n1362 vss.n1361 0.853
R1057 vss.n1351 vss.n1350 0.853
R1058 vss.n1340 vss.n1339 0.853
R1059 vss.n1452 vss.n1451 0.853
R1060 vss.n1465 vss.n1464 0.853
R1061 vss.n1692 vss.n1660 0.853
R1062 vss.n1625 vss.n717 0.853
R1063 vss.n945 vss.n942 0.853
R1064 vss.n946 vss.n945 0.853
R1065 vss.n1625 vss.n1624 0.853
R1066 vss.n1693 vss.n1692 0.853
R1067 vss.n1677 vss.n1675 0.853
R1068 vss.n1682 vss.n1672 0.853
R1069 vss.n1687 vss.n1666 0.853
R1070 vss.n1720 vss.n1719 0.853
R1071 vss.n1779 vss.n1776 0.853
R1072 vss.n1747 vss.n1744 0.853
R1073 vss.n1733 vss.n1730 0.853
R1074 vss.n1734 vss.n1733 0.853
R1075 vss.n1748 vss.n1747 0.853
R1076 vss.n1780 vss.n1779 0.853
R1077 vss.n1937 vss.n1936 0.853
R1078 vss.n1944 vss.n1943 0.853
R1079 vss.n1945 vss.n1944 0.853
R1080 vss.n2058 vss.n2057 0.853
R1081 vss.n2175 vss.n2174 0.853
R1082 vss.n474 vss.n473 0.853
R1083 vss.n549 vss.n474 0.853
R1084 vss.n512 vss.n510 0.853
R1085 vss.n526 vss.n523 0.853
R1086 vss.n545 vss.n542 0.853
R1087 vss.n546 vss.n545 0.853
R1088 vss.n527 vss.n526 0.853
R1089 vss.n513 vss.n512 0.853
R1090 vss.n2712 vss.n2711 0.853
R1091 vss.n2348 vss.n2347 0.853
R1092 vss.n2362 vss.n2361 0.853
R1093 vss.n2702 vss.n2700 0.853
R1094 vss.n2717 vss.n2692 0.853
R1095 vss.n2680 vss.n2677 0.853
R1096 vss.n2648 vss.n395 0.853
R1097 vss.n2618 vss.n2614 0.853
R1098 vss.n2623 vss.n2608 0.853
R1099 vss.n2628 vss.n2602 0.853
R1100 vss.n2633 vss.n2599 0.853
R1101 vss.n2634 vss.n2633 0.853
R1102 vss.n2648 vss.n2647 0.853
R1103 vss.n2681 vss.n2680 0.853
R1104 vss.n2718 vss.n2717 0.853
R1105 vss.n2537 vss.n2536 0.853
R1106 vss.n428 vss.n427 0.853
R1107 vss.n417 vss.n416 0.853
R1108 vss.n406 vss.n405 0.853
R1109 vss.n2585 vss.n2584 0.853
R1110 vss.n2568 vss.n2567 0.853
R1111 vss.n2558 vss.n2557 0.853
R1112 vss.n2290 vss.n2289 0.853
R1113 vss.n2381 vss.n2380 0.853
R1114 vss.n2380 vss.n2379 0.853
R1115 vss.n2400 vss.n2399 0.853
R1116 vss.n2399 vss.n2398 0.853
R1117 vss.n2433 vss.n2432 0.853
R1118 vss.n2415 vss.n2403 0.853
R1119 vss.n2415 vss.n2414 0.853
R1120 vss.n2444 vss.n2443 0.853
R1121 vss.n2465 vss.n2464 0.853
R1122 vss.n2312 vss.n2311 0.853
R1123 vss.n2502 vss.n2501 0.853
R1124 vss.n2501 vss.n2500 0.853
R1125 vss.n2301 vss.n2300 0.853
R1126 vss.n2164 vss.n2163 0.853
R1127 vss.n2517 vss.n2516 0.853
R1128 vss.n2518 vss.n2517 0.853
R1129 vss.n2236 vss.n2235 0.853
R1130 vss.n2186 vss.n2185 0.853
R1131 vss.n2273 vss.n2272 0.853
R1132 vss.n2272 vss.n2271 0.853
R1133 vss.n2066 vss.n2064 0.853
R1134 vss.n2104 vss.n2103 0.853
R1135 vss.n2096 vss.n2095 0.853
R1136 vss.n2083 vss.n2082 0.853
R1137 vss.n2143 vss.n2141 0.853
R1138 vss.n593 vss.n592 0.853
R1139 vss.n630 vss.n619 0.853
R1140 vss.n1994 vss.n1992 0.853
R1141 vss.n642 vss.n641 0.853
R1142 vss.n1983 vss.n1981 0.853
R1143 vss.n682 vss.n681 0.853
R1144 vss.n1984 vss.n1983 0.853
R1145 vss.n1810 vss.n1809 0.853
R1146 vss.n1863 vss.n1862 0.853
R1147 vss.n1862 vss.n1861 0.853
R1148 vss.n1809 vss.n1808 0.853
R1149 vss.n1841 vss.n1840 0.853
R1150 vss.n1831 vss.n1830 0.853
R1151 vss.n2815 vss.n2814 0.853
R1152 vss.n2814 vss.n2813 0.853
R1153 vss.n2783 vss.n2782 0.853
R1154 vss.n2782 vss.n2781 0.853
R1155 vss.n2800 vss.n2799 0.853
R1156 vss.n2799 vss.n2798 0.853
R1157 vss.n2769 vss.n2768 0.853
R1158 vss.n2768 vss.n2767 0.853
R1159 vss.n2755 vss.n2754 0.853
R1160 vss.n2754 vss.n2753 0.853
R1161 vss.n341 vss.n312 0.853
R1162 vss.n346 vss.n269 0.853
R1163 vss.n234 vss.n233 0.853
R1164 vss.n223 vss.n222 0.853
R1165 vss.n212 vss.n211 0.853
R1166 vss.n347 vss.n346 0.853
R1167 vss.n341 vss.n340 0.853
R1168 vss.n2876 vss.n2875 0.853
R1169 vss.n167 vss.n166 0.853
R1170 vss.n2914 vss.n2913 0.853
R1171 vss.n2956 vss.n2886 0.853
R1172 vss.n3166 vss.n3134 0.853
R1173 vss.n2927 vss.n2926 0.853
R1174 vss.n3258 vss.n3257 0.853
R1175 vss.n3290 vss.n3289 0.853
R1176 vss.n3286 vss.n3285 0.853
R1177 vss.n101 vss.n100 0.853
R1178 vss.n18 vss.n17 0.853
R1179 vss.n82 vss.n81 0.853
R1180 vss.n45 vss.n43 0.853
R1181 vss.n46 vss.n45 0.853
R1182 vss.n102 vss.n101 0.853
R1183 vss.n19 vss.n18 0.853
R1184 vss.n83 vss.n82 0.853
R1185 vss.n3307 vss.n3306 0.853
R1186 vss.n3321 vss.n3320 0.853
R1187 vss.n3240 vss.n3239 0.853
R1188 vss vss.n2882 0.843143
R1189 vss.n2882 vss 0.715571
R1190 vss.n584 vss.n583 0.699777
R1191 vss.n1991 vss.n1990 0.699777
R1192 vss.n2131 vss.n2130 0.699516
R1193 vss.n624 vss.n623 0.699516
R1194 vss.n780 vss.n779 0.698382
R1195 vss.n2068 vss.n2067 0.698382
R1196 vss.n644 vss.n643 0.698382
R1197 vss.n3260 vss.n3259 0.698382
R1198 vss.n97 vss.n96 0.689091
R1199 vss.n649 vss.n648 0.684595
R1200 vss.n785 vss.n784 0.684595
R1201 vss.n2073 vss.n2072 0.684595
R1202 vss.n3270 vss.n3269 0.684595
R1203 vss.n1134 vss.n1131 0.682713
R1204 vss.n2129 vss.n2128 0.682713
R1205 vss.n3006 vss.n3005 0.682697
R1206 vss.n3002 vss.n3001 0.682697
R1207 vss.n2998 vss.n2997 0.682697
R1208 vss.n2994 vss.n2993 0.682697
R1209 vss.n2990 vss.n2989 0.682697
R1210 vss.n2982 vss.n2981 0.682697
R1211 vss.n3133 vss.n3132 0.682697
R1212 vss.n2970 vss.n2969 0.682697
R1213 vss.n2974 vss.n2973 0.682697
R1214 vss.n2978 vss.n2977 0.682697
R1215 vss.n2986 vss.n2985 0.682697
R1216 vss.n3284 vss.n3283 0.682697
R1217 vss.n3305 vss.n3304 0.682697
R1218 vss.n3319 vss.n3318 0.682697
R1219 vss.n3292 vss.n3291 0.682697
R1220 vss.n3218 vss.n3216 0.565206
R1221 vss vss.n1210 0.5645
R1222 vss.n1210 vss.n1116 0.4705
R1223 vss.n2885 vss 0.426857
R1224 vss.n96 vss.n95 0.41184
R1225 vss.n3017 vss.n3009 0.376971
R1226 vss.n2069 vss.n2068 0.354051
R1227 vss.n645 vss.n644 0.354051
R1228 vss.n117 vss 0.353441
R1229 vss.n781 vss.n780 0.352759
R1230 vss.n3261 vss.n3260 0.350986
R1231 vss.n3202 vss 0.339791
R1232 vss.n1855 vss.n1854 0.33661
R1233 vss.n278 vss.n277 0.33661
R1234 vss.n2251 vss.n2250 0.336142
R1235 vss.n3202 vss 0.294692
R1236 vss.n3180 vss.n3179 0.261125
R1237 vss.n2076 vss.n461 0.253125
R1238 vss.n2148 vss.n461 0.249386
R1239 vss.n344 vss.n343 0.212
R1240 vss.n1449 vss.n1448 0.212
R1241 vss.n1468 vss.n1467 0.212
R1242 vss.n1607 vss.n1606 0.212
R1243 vss.n1100 vss.n1099 0.212
R1244 vss.n1018 vss.n1017 0.212
R1245 vss.n965 vss.n964 0.212
R1246 vss.n1628 vss.n1627 0.212
R1247 vss.n2239 vss.n2238 0.212
R1248 vss.n2540 vss.n2539 0.212
R1249 vss.n2631 vss.n2630 0.212
R1250 vss.n2651 vss.n2650 0.212
R1251 vss.n2468 vss.n2467 0.212
R1252 vss.n2385 vss.n2384 0.212
R1253 vss.n2896 vss.n2895 0.203675
R1254 vss.n1205 vss.n1124 0.203675
R1255 vss.n2115 vss.n596 0.203675
R1256 vss.n2020 vss.n2018 0.203675
R1257 vss.n111 vss 0.202323
R1258 vss.n3214 vss 0.202272
R1259 vss.n652 vss.n651 0.183261
R1260 vss.n2884 vss 0.182195
R1261 vss.n1987 vss 0.180125
R1262 vss.n2132 vss 0.170375
R1263 vss vss.n3296 0.167718
R1264 vss.n115 vss 0.157066
R1265 vss.n3298 vss 0.156006
R1266 vss.n3231 vss 0.153278
R1267 vss.n67 vss.n66 0.151979
R1268 vss.n76 vss.n75 0.151979
R1269 vss.n3170 vss.n2885 0.147518
R1270 vss.n3295 vss 0.140344
R1271 vss.n1228 vss.n787 0.127459
R1272 vss.n1211 vss 0.125741
R1273 vss.n3232 vss 0.122593
R1274 vss.n3281 vss.n3280 0.120292
R1275 vss.n2077 vss.n2076 0.119277
R1276 vss.n1986 vss 0.112761
R1277 vss.n3281 vss 0.106981
R1278 vss.n130 vss 0.104812
R1279 vss.n1947 vss 0.104812
R1280 vss.n2514 vss 0.103332
R1281 vss.n3265 vss.n3264 0.102977
R1282 vss.n2076 vss.n2075 0.101141
R1283 vss.n1325 vss 0.0994474
R1284 vss.n2905 vss.n2904 0.0929479
R1285 vss.n614 vss.n613 0.0929479
R1286 vss.n3266 vss.n3265 0.0904594
R1287 vss.n1324 vss 0.0903012
R1288 vss.n1325 vss 0.0897843
R1289 vss vss.n2884 0.0847561
R1290 vss.n3230 vss 0.0825312
R1291 vss.n1196 vss.n1195 0.0825312
R1292 vss.n577 vss.n576 0.0825312
R1293 vss.n2881 vss 0.0801269
R1294 vss.n2132 vss 0.0763587
R1295 vss.n3231 vss.n3230 0.0760208
R1296 vss.n1620 vss 0.0753227
R1297 vss.n3130 vss.n3124 0.0746936
R1298 vss.n3119 vss.n3115 0.0746936
R1299 vss.n3108 vss.n3104 0.0746936
R1300 vss.n3104 vss.n3100 0.0746936
R1301 vss.n3095 vss.n3091 0.0746936
R1302 vss.n3084 vss.n3080 0.0746936
R1303 vss.n3075 vss.n3071 0.0746936
R1304 vss.n3066 vss.n3061 0.0746936
R1305 vss.n3056 vss.n3052 0.0746936
R1306 vss.n3052 vss.n3048 0.0746936
R1307 vss.n3041 vss.n3037 0.0746936
R1308 vss.n3032 vss.n3028 0.0746936
R1309 vss.n3022 vss.n3018 0.0746936
R1310 vss.n2960 vss.n2959 0.0734167
R1311 vss.n621 vss.n620 0.0734167
R1312 vss.n2885 vss 0.0732927
R1313 vss.n3042 vss.n3041 0.0730806
R1314 vss.n3300 vss.n3298 0.0728562
R1315 vss.n2724 vss 0.0724848
R1316 vss.n3033 vss.n3032 0.0722742
R1317 vss.n3023 vss.n3022 0.0714677
R1318 vss.n3288 vss.n3287 0.0711263
R1319 vss.n1211 vss 0.0707673
R1320 vss.n3011 vss.n3007 0.0690484
R1321 vss.n288 vss.n287 0.0685147
R1322 vss.n284 vss.n283 0.0685147
R1323 vss.n276 vss.n275 0.0685147
R1324 vss.n249 vss.n248 0.0685147
R1325 vss.n256 vss.n255 0.0685147
R1326 vss.n263 vss.n262 0.0685147
R1327 vss.n2850 vss.n2849 0.0685147
R1328 vss.n2857 vss.n2856 0.0685147
R1329 vss.n2869 vss.n2868 0.0685147
R1330 vss.n1821 vss.n1820 0.0685147
R1331 vss.n1895 vss.n1894 0.0685147
R1332 vss.n1891 vss.n1890 0.0685147
R1333 vss.n1884 vss.n1883 0.0685147
R1334 vss.n1763 vss.n1762 0.0685147
R1335 vss.n1770 vss.n1769 0.0685147
R1336 vss.n1377 vss.n1376 0.0685147
R1337 vss.n1384 vss.n1383 0.0685147
R1338 vss.n1391 vss.n1390 0.0685147
R1339 vss.n1405 vss.n1404 0.0685147
R1340 vss.n1510 vss.n1509 0.0685147
R1341 vss.n1517 vss.n1516 0.0685147
R1342 vss.n1524 vss.n1523 0.0685147
R1343 vss.n1539 vss.n1538 0.0685147
R1344 vss.n1535 vss.n1534 0.0685147
R1345 vss.n1295 vss.n1294 0.0685147
R1346 vss.n1302 vss.n1301 0.0685147
R1347 vss.n1163 vss.n1162 0.0685147
R1348 vss.n1159 vss.n1158 0.0685147
R1349 vss.n1152 vss.n738 0.0685147
R1350 vss.n830 vss.n829 0.0685147
R1351 vss.n837 vss.n836 0.0685147
R1352 vss.n844 vss.n843 0.0685147
R1353 vss.n1083 vss.n1082 0.0685147
R1354 vss.n853 vss.n852 0.0685147
R1355 vss.n1031 vss.n1030 0.0685147
R1356 vss.n1071 vss.n1070 0.0685147
R1357 vss.n1067 vss.n1066 0.0685147
R1358 vss.n1028 vss.n1027 0.0685147
R1359 vss.n1006 vss.n1005 0.0685147
R1360 vss.n704 vss.n703 0.0685147
R1361 vss.n711 vss.n710 0.0685147
R1362 vss.n1650 vss.n1649 0.0685147
R1363 vss.n1646 vss.n1645 0.0685147
R1364 vss.n1639 vss.n1638 0.0685147
R1365 vss.n1955 vss.n1954 0.0685147
R1366 vss.n1962 vss.n1961 0.0685147
R1367 vss.n1974 vss.n1973 0.0685147
R1368 vss.n2043 vss.n2042 0.0685147
R1369 vss.n2050 vss.n2049 0.0685147
R1370 vss.n2222 vss.n2221 0.0685147
R1371 vss.n2192 vss.n2191 0.0685147
R1372 vss.n439 vss.n438 0.0685147
R1373 vss.n2249 vss.n2248 0.0685147
R1374 vss.n2257 vss.n2256 0.0685147
R1375 vss.n2264 vss.n2263 0.0685147
R1376 vss.n494 vss.n493 0.0685147
R1377 vss.n504 vss.n503 0.0685147
R1378 vss.n2210 vss.n2209 0.0685147
R1379 vss.n2206 vss.n437 0.0685147
R1380 vss.n2530 vss.n2529 0.0685147
R1381 vss.n2549 vss.n2548 0.0685147
R1382 vss.n375 vss.n374 0.0685147
R1383 vss.n382 vss.n381 0.0685147
R1384 vss.n389 vss.n388 0.0685147
R1385 vss.n2668 vss.n2667 0.0685147
R1386 vss.n2664 vss.n2663 0.0685147
R1387 vss.n2657 vss.n2656 0.0685147
R1388 vss.n2480 vss.n2479 0.0685147
R1389 vss.n2487 vss.n2486 0.0685147
R1390 vss.n2494 vss.n2493 0.0685147
R1391 vss.n2456 vss.n2455 0.0685147
R1392 vss.n2341 vss.n2340 0.0685147
R1393 vss.n2744 vss.n2743 0.0685147
R1394 vss.n2740 vss.n2739 0.0685147
R1395 vss.n2824 vss.n2823 0.0685147
R1396 vss.n2837 vss.n2836 0.0685147
R1397 vss.n2833 vss.n2832 0.0685147
R1398 vss.n3131 vss.n3130 0.0682419
R1399 vss.n3296 vss.n3295 0.0670294
R1400 vss.n3325 vss 0.0663531
R1401 vss.n1130 vss.n1129 0.0656042
R1402 vss.n2126 vss.n2120 0.0656042
R1403 vss.n613 vss.n604 0.0643021
R1404 vss.n3170 vss.n3169 0.0639127
R1405 vss.n2723 vss.n357 0.0635421
R1406 vss.n3096 vss.n3095 0.0625968
R1407 vss.n1865 vss.n1864 0.0620273
R1408 vss.n1325 vss.n1324 0.061334
R1409 vss.n3303 vss.n3302 0.0610288
R1410 vss.n3061 vss.n3057 0.0609839
R1411 vss.n1129 vss 0.0603958
R1412 vss.n2120 vss 0.0603958
R1413 vss.n3071 vss.n3067 0.0601774
R1414 vss.n3317 vss.n3316 0.057898
R1415 vss.n358 vss 0.0560168
R1416 vss.n1216 vss 0.0548478
R1417 vss.n2135 vss 0.0548478
R1418 vss.n3115 vss.n3109 0.0545323
R1419 vss.n3275 vss 0.0537407
R1420 vss.n2722 vss.n358 0.0524782
R1421 vss.n3323 vss.n105 0.0523603
R1422 vss.n1136 vss.n1116 0.0518289
R1423 vss.n3172 vss 0.0515286
R1424 vss.n2932 vss 0.0512812
R1425 vss.n1178 vss 0.0512812
R1426 vss vss.n558 0.0512812
R1427 vss vss.n2014 0.0512812
R1428 vss.n2149 vss 0.0506333
R1429 vss.n2722 vss.n2721 0.0505748
R1430 vss.n2724 vss.n2723 0.0496761
R1431 vss.n3239 vss.n3201 0.0493281
R1432 vss vss.n2131 0.0492848
R1433 vss.n1226 vss.n733 0.0491931
R1434 vss.n3282 vss.n3281 0.0483395
R1435 vss.n218 vss.n217 0.0482941
R1436 vss.n229 vss.n228 0.0482941
R1437 vss.n240 vss.n239 0.0482941
R1438 vss.n309 vss.n308 0.0482941
R1439 vss.n303 vss.n302 0.0482941
R1440 vss.n297 vss.n296 0.0482941
R1441 vss.n162 vss.n161 0.0482941
R1442 vss.n2860 vss.n2859 0.0482941
R1443 vss.n156 vss.n155 0.0482941
R1444 vss.n1917 vss.n1916 0.0482941
R1445 vss.n1911 vss.n1910 0.0482941
R1446 vss.n1905 vss.n1904 0.0482941
R1447 vss.n1346 vss.n1345 0.0482941
R1448 vss.n1357 vss.n1356 0.0482941
R1449 vss.n1368 vss.n1367 0.0482941
R1450 vss.n1415 vss.n1414 0.0482941
R1451 vss.n1421 vss.n1420 0.0482941
R1452 vss.n723 vss.n722 0.0482941
R1453 vss.n1479 vss.n1478 0.0482941
R1454 vss.n1490 vss.n1489 0.0482941
R1455 vss.n1501 vss.n1500 0.0482941
R1456 vss.n743 vss.n742 0.0482941
R1457 vss.n749 vss.n748 0.0482941
R1458 vss.n755 vss.n754 0.0482941
R1459 vss.n799 vss.n798 0.0482941
R1460 vss.n810 vss.n809 0.0482941
R1461 vss.n821 vss.n820 0.0482941
R1462 vss.n1093 vss.n1092 0.0482941
R1463 vss.n856 vss.n855 0.0482941
R1464 vss.n1035 vss.n1034 0.0482941
R1465 vss.n884 vss.n883 0.0482941
R1466 vss.n868 vss.n867 0.0482941
R1467 vss.n894 vss.n893 0.0482941
R1468 vss.n900 vss.n899 0.0482941
R1469 vss.n913 vss.n912 0.0482941
R1470 vss.n1657 vss.n1656 0.0482941
R1471 vss.n1663 vss.n1662 0.0482941
R1472 vss.n1669 vss.n1668 0.0482941
R1473 vss.n677 vss.n676 0.0482941
R1474 vss.n1965 vss.n1964 0.0482941
R1475 vss.n671 vss.n670 0.0482941
R1476 vss.n2028 vss.n2027 0.0482941
R1477 vss.n2090 vss.n2089 0.0482941
R1478 vss.n2170 vss.n2169 0.0482941
R1479 vss.n2181 vss.n2180 0.0482941
R1480 vss.n2242 vss.n2241 0.0482941
R1481 vss.n2232 vss.n2231 0.0482941
R1482 vss.n2195 vss.n2194 0.0482941
R1483 vss.n443 vss.n442 0.0482941
R1484 vss.n412 vss.n411 0.0482941
R1485 vss.n423 vss.n422 0.0482941
R1486 vss.n434 vss.n433 0.0482941
R1487 vss.n2563 vss.n2562 0.0482941
R1488 vss.n2573 vss.n2572 0.0482941
R1489 vss.n2590 vss.n2589 0.0482941
R1490 vss.n2604 vss.n2603 0.0482941
R1491 vss.n2610 vss.n2609 0.0482941
R1492 vss.n366 vss.n365 0.0482941
R1493 vss.n2689 vss.n2688 0.0482941
R1494 vss.n2708 vss.n2707 0.0482941
R1495 vss.n2296 vss.n2295 0.0482941
R1496 vss.n2307 vss.n2306 0.0482941
R1497 vss.n2471 vss.n2470 0.0482941
R1498 vss.n2439 vss.n2438 0.0482941
R1499 vss.n2421 vss.n2420 0.0482941
R1500 vss.n2405 vss.n2404 0.0482941
R1501 vss.n2377 vss.n2376 0.0482941
R1502 vss.n2359 vss.n2358 0.0482941
R1503 vss.n1836 vss.n1835 0.0482941
R1504 vss.n1848 vss.n1847 0.0482941
R1505 vss.n187 vss.n186 0.0482941
R1506 vss.n181 vss.n180 0.0482941
R1507 vss.n175 vss.n174 0.0482941
R1508 vss.n3080 vss.n3076 0.0480806
R1509 vss.n3236 vss.n3235 0.0479806
R1510 vss.n949 vss 0.0479063
R1511 vss.n3280 vss.n3278 0.047375
R1512 vss.n1942 vss 0.0471846
R1513 vss.n2721 vss 0.0466376
R1514 vss.n3213 vss.n3209 0.0454219
R1515 vss.n3326 vss.n3325 0.0446573
R1516 vss.n1138 vss.n1131 0.0444189
R1517 vss.n2128 vss.n2127 0.0444189
R1518 vss.n1222 vss.n1215 0.0434688
R1519 vss.n2141 vss.n2134 0.0434688
R1520 vss.n2913 vss.n2902 0.0427297
R1521 vss.n608 vss.n607 0.0427297
R1522 vss.n2147 vss.n550 0.0425162
R1523 vss.n1865 vss.n690 0.0424314
R1524 vss.n3085 vss.n3084 0.041629
R1525 vss.n133 vss.n128 0.0415156
R1526 vss.n3195 vss.n110 0.0415156
R1527 vss.n776 vss.n772 0.0415156
R1528 vss.n1945 vss.n685 0.0415156
R1529 vss.n2064 vss.n2060 0.0415156
R1530 vss.n641 vss.n637 0.0415156
R1531 vss.n3257 vss.n3253 0.0415156
R1532 vss.n100 vss.n91 0.0415156
R1533 vss.n1135 vss.n1133 0.0411354
R1534 vss.n590 vss.n552 0.0411354
R1535 vss.n628 vss.n627 0.0411354
R1536 vss.n116 vss.n115 0.0408226
R1537 vss.n2882 vss.n139 0.0399444
R1538 vss.n3172 vss 0.0398007
R1539 vss.n2150 vss.n2149 0.039647
R1540 vss.n88 vss.n87 0.0395625
R1541 vss.n43 vss.n42 0.0395625
R1542 vss.n1227 vss.n1113 0.039516
R1543 vss.n2802 vss 0.0393305
R1544 vss.n1326 vss.n1325 0.0392005
R1545 vss.n291 vss.n288 0.0391029
R1546 vss.n287 vss.n286 0.0391029
R1547 vss.n285 vss.n284 0.0391029
R1548 vss.n283 vss.n282 0.0391029
R1549 vss.n281 vss.n276 0.0391029
R1550 vss.n275 vss.n274 0.0391029
R1551 vss.n248 vss.n247 0.0391029
R1552 vss.n253 vss.n249 0.0391029
R1553 vss.n255 vss.n254 0.0391029
R1554 vss.n260 vss.n256 0.0391029
R1555 vss.n262 vss.n261 0.0391029
R1556 vss.n267 vss.n263 0.0391029
R1557 vss.n211 vss.n210 0.0391029
R1558 vss.n220 vss.n219 0.0391029
R1559 vss.n222 vss.n221 0.0391029
R1560 vss.n231 vss.n230 0.0391029
R1561 vss.n233 vss.n232 0.0391029
R1562 vss.n242 vss.n241 0.0391029
R1563 vss.n311 vss.n310 0.0391029
R1564 vss.n307 vss.n306 0.0391029
R1565 vss.n305 vss.n304 0.0391029
R1566 vss.n301 vss.n300 0.0391029
R1567 vss.n299 vss.n298 0.0391029
R1568 vss.n295 vss.n294 0.0391029
R1569 vss.n2849 vss.n2848 0.0391029
R1570 vss.n2851 vss.n2850 0.0391029
R1571 vss.n2856 vss.n2855 0.0391029
R1572 vss.n2863 vss.n2857 0.0391029
R1573 vss.n2868 vss.n2867 0.0391029
R1574 vss.n2873 vss.n2869 0.0391029
R1575 vss.n164 vss.n163 0.0391029
R1576 vss.n160 vss.n159 0.0391029
R1577 vss.n2862 vss.n2861 0.0391029
R1578 vss.n154 vss.n153 0.0391029
R1579 vss.n2875 vss.n157 0.0391029
R1580 vss.n1826 vss.n1821 0.0391029
R1581 vss.n1820 vss.n1819 0.0391029
R1582 vss.n1818 vss.n1815 0.0391029
R1583 vss.n1860 vss.n1853 0.0391029
R1584 vss.n1859 vss.n1858 0.0391029
R1585 vss.n1807 vss.n1804 0.0391029
R1586 vss.n1899 vss.n1895 0.0391029
R1587 vss.n1894 vss.n1893 0.0391029
R1588 vss.n1892 vss.n1891 0.0391029
R1589 vss.n1890 vss.n1889 0.0391029
R1590 vss.n1888 vss.n1884 0.0391029
R1591 vss.n1883 vss.n1882 0.0391029
R1592 vss.n1919 vss.n1918 0.0391029
R1593 vss.n1915 vss.n1914 0.0391029
R1594 vss.n1913 vss.n1912 0.0391029
R1595 vss.n1909 vss.n1908 0.0391029
R1596 vss.n1907 vss.n1906 0.0391029
R1597 vss.n1903 vss.n1902 0.0391029
R1598 vss.n1715 vss.n1714 0.0391029
R1599 vss.n1760 vss.n1756 0.0391029
R1600 vss.n1762 vss.n1761 0.0391029
R1601 vss.n1767 vss.n1763 0.0391029
R1602 vss.n1769 vss.n1768 0.0391029
R1603 vss.n1774 vss.n1770 0.0391029
R1604 vss.n1718 vss.n1717 0.0391029
R1605 vss.n1727 vss.n1726 0.0391029
R1606 vss.n1730 vss.n1729 0.0391029
R1607 vss.n1741 vss.n1740 0.0391029
R1608 vss.n1744 vss.n1743 0.0391029
R1609 vss.n1755 vss.n1754 0.0391029
R1610 vss.n1376 vss.n1375 0.0391029
R1611 vss.n1381 vss.n1377 0.0391029
R1612 vss.n1383 vss.n1382 0.0391029
R1613 vss.n1388 vss.n1384 0.0391029
R1614 vss.n1390 vss.n1389 0.0391029
R1615 vss.n1395 vss.n1391 0.0391029
R1616 vss.n1339 vss.n1338 0.0391029
R1617 vss.n1348 vss.n1347 0.0391029
R1618 vss.n1350 vss.n1349 0.0391029
R1619 vss.n1359 vss.n1358 0.0391029
R1620 vss.n1361 vss.n1360 0.0391029
R1621 vss.n1370 vss.n1369 0.0391029
R1622 vss.n1409 vss.n1405 0.0391029
R1623 vss.n1404 vss.n1403 0.0391029
R1624 vss.n1402 vss.n1401 0.0391029
R1625 vss.n1429 vss.n1423 0.0391029
R1626 vss.n1428 vss.n1424 0.0391029
R1627 vss.n730 vss.n725 0.0391029
R1628 vss.n1412 vss.n1411 0.0391029
R1629 vss.n1419 vss.n1416 0.0391029
R1630 vss.n1418 vss.n1417 0.0391029
R1631 vss.n1432 vss.n1422 0.0391029
R1632 vss.n1431 vss.n1430 0.0391029
R1633 vss.n732 vss.n724 0.0391029
R1634 vss.n1509 vss.n1508 0.0391029
R1635 vss.n1514 vss.n1510 0.0391029
R1636 vss.n1516 vss.n1515 0.0391029
R1637 vss.n1521 vss.n1517 0.0391029
R1638 vss.n1523 vss.n1522 0.0391029
R1639 vss.n1528 vss.n1524 0.0391029
R1640 vss.n1472 vss.n1471 0.0391029
R1641 vss.n1481 vss.n1480 0.0391029
R1642 vss.n1483 vss.n1482 0.0391029
R1643 vss.n1492 vss.n1491 0.0391029
R1644 vss.n1494 vss.n1493 0.0391029
R1645 vss.n1503 vss.n1502 0.0391029
R1646 vss.n1543 vss.n1539 0.0391029
R1647 vss.n1538 vss.n1537 0.0391029
R1648 vss.n1536 vss.n1535 0.0391029
R1649 vss.n1577 vss.n1573 0.0391029
R1650 vss.n1561 vss.n1556 0.0391029
R1651 vss.n1547 vss.n1546 0.0391029
R1652 vss.n1596 vss.n1592 0.0391029
R1653 vss.n1595 vss.n1594 0.0391029
R1654 vss.n1582 vss.n1572 0.0391029
R1655 vss.n1581 vss.n1580 0.0391029
R1656 vss.n1563 vss.n1555 0.0391029
R1657 vss.n1247 vss.n1246 0.0391029
R1658 vss.n1264 vss.n1260 0.0391029
R1659 vss.n1299 vss.n1295 0.0391029
R1660 vss.n1301 vss.n1300 0.0391029
R1661 vss.n1306 vss.n1302 0.0391029
R1662 vss.n1250 vss.n1249 0.0391029
R1663 vss.n1259 vss.n1258 0.0391029
R1664 vss.n1268 vss.n1267 0.0391029
R1665 vss.n1279 vss.n1278 0.0391029
R1666 vss.n1282 vss.n1281 0.0391029
R1667 vss.n1293 vss.n1292 0.0391029
R1668 vss.n1164 vss.n1163 0.0391029
R1669 vss.n1162 vss.n1161 0.0391029
R1670 vss.n1160 vss.n1159 0.0391029
R1671 vss.n1158 vss.n1157 0.0391029
R1672 vss.n1153 vss.n1152 0.0391029
R1673 vss.n1236 vss.n738 0.0391029
R1674 vss.n741 vss.n740 0.0391029
R1675 vss.n745 vss.n744 0.0391029
R1676 vss.n747 vss.n746 0.0391029
R1677 vss.n751 vss.n750 0.0391029
R1678 vss.n753 vss.n752 0.0391029
R1679 vss.n757 vss.n756 0.0391029
R1680 vss.n829 vss.n828 0.0391029
R1681 vss.n834 vss.n830 0.0391029
R1682 vss.n836 vss.n835 0.0391029
R1683 vss.n841 vss.n837 0.0391029
R1684 vss.n843 vss.n842 0.0391029
R1685 vss.n849 vss.n844 0.0391029
R1686 vss.n792 vss.n791 0.0391029
R1687 vss.n801 vss.n800 0.0391029
R1688 vss.n803 vss.n802 0.0391029
R1689 vss.n812 vss.n811 0.0391029
R1690 vss.n814 vss.n813 0.0391029
R1691 vss.n823 vss.n822 0.0391029
R1692 vss.n1087 vss.n1083 0.0391029
R1693 vss.n1082 vss.n1081 0.0391029
R1694 vss.n859 vss.n853 0.0391029
R1695 vss.n1057 vss.n1031 0.0391029
R1696 vss.n1095 vss.n1094 0.0391029
R1697 vss.n1091 vss.n1090 0.0391029
R1698 vss.n858 vss.n857 0.0391029
R1699 vss.n1033 vss.n1032 0.0391029
R1700 vss.n1056 vss.n1036 0.0391029
R1701 vss.n1072 vss.n1071 0.0391029
R1702 vss.n1070 vss.n1069 0.0391029
R1703 vss.n1068 vss.n1067 0.0391029
R1704 vss.n1066 vss.n1065 0.0391029
R1705 vss.n1029 vss.n1028 0.0391029
R1706 vss.n1027 vss.n1026 0.0391029
R1707 vss.n1318 vss.n1317 0.0391029
R1708 vss.n876 vss.n875 0.0391029
R1709 vss.n878 vss.n877 0.0391029
R1710 vss.n886 vss.n885 0.0391029
R1711 vss.n888 vss.n887 0.0391029
R1712 vss.n870 vss.n869 0.0391029
R1713 vss.n1010 vss.n1006 0.0391029
R1714 vss.n1005 vss.n1004 0.0391029
R1715 vss.n1003 vss.n1002 0.0391029
R1716 vss.n908 vss.n902 0.0391029
R1717 vss.n907 vss.n903 0.0391029
R1718 vss.n920 vss.n915 0.0391029
R1719 vss.n1013 vss.n1012 0.0391029
R1720 vss.n898 vss.n895 0.0391029
R1721 vss.n897 vss.n896 0.0391029
R1722 vss.n911 vss.n901 0.0391029
R1723 vss.n910 vss.n909 0.0391029
R1724 vss.n922 vss.n914 0.0391029
R1725 vss.n973 vss.n972 0.0391029
R1726 vss.n701 vss.n697 0.0391029
R1727 vss.n703 vss.n702 0.0391029
R1728 vss.n708 vss.n704 0.0391029
R1729 vss.n710 vss.n709 0.0391029
R1730 vss.n715 vss.n711 0.0391029
R1731 vss.n976 vss.n975 0.0391029
R1732 vss.n954 vss.n953 0.0391029
R1733 vss.n957 vss.n956 0.0391029
R1734 vss.n939 vss.n938 0.0391029
R1735 vss.n942 vss.n941 0.0391029
R1736 vss.n696 vss.n695 0.0391029
R1737 vss.n1654 vss.n1650 0.0391029
R1738 vss.n1649 vss.n1648 0.0391029
R1739 vss.n1647 vss.n1646 0.0391029
R1740 vss.n1645 vss.n1644 0.0391029
R1741 vss.n1643 vss.n1639 0.0391029
R1742 vss.n1638 vss.n1637 0.0391029
R1743 vss.n1659 vss.n1658 0.0391029
R1744 vss.n1666 vss.n1661 0.0391029
R1745 vss.n1665 vss.n1664 0.0391029
R1746 vss.n1672 vss.n1667 0.0391029
R1747 vss.n1671 vss.n1670 0.0391029
R1748 vss.n1675 vss.n1673 0.0391029
R1749 vss.n1954 vss.n1953 0.0391029
R1750 vss.n1956 vss.n1955 0.0391029
R1751 vss.n1961 vss.n1960 0.0391029
R1752 vss.n1968 vss.n1962 0.0391029
R1753 vss.n1973 vss.n1972 0.0391029
R1754 vss.n1979 vss.n1974 0.0391029
R1755 vss.n679 vss.n678 0.0391029
R1756 vss.n675 vss.n674 0.0391029
R1757 vss.n1967 vss.n1966 0.0391029
R1758 vss.n669 vss.n668 0.0391029
R1759 vss.n1981 vss.n672 0.0391029
R1760 vss.n2105 vss.n2025 0.0391029
R1761 vss.n2040 vss.n2036 0.0391029
R1762 vss.n2042 vss.n2041 0.0391029
R1763 vss.n2047 vss.n2043 0.0391029
R1764 vss.n2049 vss.n2048 0.0391029
R1765 vss.n2055 vss.n2050 0.0391029
R1766 vss.n2104 vss.n2029 0.0391029
R1767 vss.n2080 vss.n2079 0.0391029
R1768 vss.n2082 vss.n2081 0.0391029
R1769 vss.n2092 vss.n2091 0.0391029
R1770 vss.n2095 vss.n2094 0.0391029
R1771 vss.n2035 vss.n2034 0.0391029
R1772 vss.n2163 vss.n2162 0.0391029
R1773 vss.n2172 vss.n2171 0.0391029
R1774 vss.n2174 vss.n2173 0.0391029
R1775 vss.n2183 vss.n2182 0.0391029
R1776 vss.n2185 vss.n2184 0.0391029
R1777 vss.n2244 vss.n2243 0.0391029
R1778 vss.n2226 vss.n2222 0.0391029
R1779 vss.n2221 vss.n2220 0.0391029
R1780 vss.n2198 vss.n2192 0.0391029
R1781 vss.n2519 vss.n439 0.0391029
R1782 vss.n2234 vss.n2233 0.0391029
R1783 vss.n2230 vss.n2229 0.0391029
R1784 vss.n2197 vss.n2196 0.0391029
R1785 vss.n441 vss.n440 0.0391029
R1786 vss.n2518 vss.n444 0.0391029
R1787 vss.n2248 vss.n2247 0.0391029
R1788 vss.n2254 vss.n2249 0.0391029
R1789 vss.n2256 vss.n2255 0.0391029
R1790 vss.n2261 vss.n2257 0.0391029
R1791 vss.n2263 vss.n2262 0.0391029
R1792 vss.n2269 vss.n2264 0.0391029
R1793 vss.n470 vss.n469 0.0391029
R1794 vss.n538 vss.n535 0.0391029
R1795 vss.n501 vss.n494 0.0391029
R1796 vss.n503 vss.n502 0.0391029
R1797 vss.n508 vss.n504 0.0391029
R1798 vss.n473 vss.n472 0.0391029
R1799 vss.n534 vss.n533 0.0391029
R1800 vss.n542 vss.n541 0.0391029
R1801 vss.n520 vss.n519 0.0391029
R1802 vss.n523 vss.n522 0.0391029
R1803 vss.n492 vss.n491 0.0391029
R1804 vss.n2211 vss.n2210 0.0391029
R1805 vss.n2209 vss.n2208 0.0391029
R1806 vss.n2207 vss.n2206 0.0391029
R1807 vss.n2527 vss.n437 0.0391029
R1808 vss.n2529 vss.n2528 0.0391029
R1809 vss.n2534 vss.n2530 0.0391029
R1810 vss.n405 vss.n404 0.0391029
R1811 vss.n414 vss.n413 0.0391029
R1812 vss.n416 vss.n415 0.0391029
R1813 vss.n425 vss.n424 0.0391029
R1814 vss.n427 vss.n426 0.0391029
R1815 vss.n436 vss.n435 0.0391029
R1816 vss.n2553 vss.n2549 0.0391029
R1817 vss.n2548 vss.n2547 0.0391029
R1818 vss.n2546 vss.n2545 0.0391029
R1819 vss.n2581 vss.n2575 0.0391029
R1820 vss.n2580 vss.n2576 0.0391029
R1821 vss.n2597 vss.n2592 0.0391029
R1822 vss.n2556 vss.n2555 0.0391029
R1823 vss.n2567 vss.n2564 0.0391029
R1824 vss.n2566 vss.n2565 0.0391029
R1825 vss.n2584 vss.n2574 0.0391029
R1826 vss.n2583 vss.n2582 0.0391029
R1827 vss.n2599 vss.n2591 0.0391029
R1828 vss.n374 vss.n373 0.0391029
R1829 vss.n379 vss.n375 0.0391029
R1830 vss.n381 vss.n380 0.0391029
R1831 vss.n386 vss.n382 0.0391029
R1832 vss.n388 vss.n387 0.0391029
R1833 vss.n393 vss.n389 0.0391029
R1834 vss.n2602 vss.n2601 0.0391029
R1835 vss.n2606 vss.n2605 0.0391029
R1836 vss.n2608 vss.n2607 0.0391029
R1837 vss.n2612 vss.n2611 0.0391029
R1838 vss.n2614 vss.n2613 0.0391029
R1839 vss.n368 vss.n367 0.0391029
R1840 vss.n2672 vss.n2668 0.0391029
R1841 vss.n2667 vss.n2666 0.0391029
R1842 vss.n2665 vss.n2664 0.0391029
R1843 vss.n2663 vss.n2662 0.0391029
R1844 vss.n2661 vss.n2657 0.0391029
R1845 vss.n2676 vss.n2675 0.0391029
R1846 vss.n2692 vss.n2687 0.0391029
R1847 vss.n2691 vss.n2690 0.0391029
R1848 vss.n2711 vss.n2706 0.0391029
R1849 vss.n2710 vss.n2709 0.0391029
R1850 vss.n2700 vss.n2693 0.0391029
R1851 vss.n2479 vss.n2478 0.0391029
R1852 vss.n2484 vss.n2480 0.0391029
R1853 vss.n2486 vss.n2485 0.0391029
R1854 vss.n2491 vss.n2487 0.0391029
R1855 vss.n2493 vss.n2492 0.0391029
R1856 vss.n2498 vss.n2494 0.0391029
R1857 vss.n2289 vss.n2288 0.0391029
R1858 vss.n2298 vss.n2297 0.0391029
R1859 vss.n2300 vss.n2299 0.0391029
R1860 vss.n2309 vss.n2308 0.0391029
R1861 vss.n2311 vss.n2310 0.0391029
R1862 vss.n2473 vss.n2472 0.0391029
R1863 vss.n2460 vss.n2456 0.0391029
R1864 vss.n2455 vss.n2454 0.0391029
R1865 vss.n2453 vss.n2452 0.0391029
R1866 vss.n2429 vss.n2423 0.0391029
R1867 vss.n2428 vss.n2424 0.0391029
R1868 vss.n2412 vss.n2407 0.0391029
R1869 vss.n2463 vss.n2462 0.0391029
R1870 vss.n2443 vss.n2440 0.0391029
R1871 vss.n2442 vss.n2441 0.0391029
R1872 vss.n2432 vss.n2422 0.0391029
R1873 vss.n2431 vss.n2430 0.0391029
R1874 vss.n2414 vss.n2406 0.0391029
R1875 vss.n2395 vss.n2394 0.0391029
R1876 vss.n2373 vss.n2369 0.0391029
R1877 vss.n2375 vss.n2374 0.0391029
R1878 vss.n2338 vss.n2334 0.0391029
R1879 vss.n2340 vss.n2339 0.0391029
R1880 vss.n2345 vss.n2341 0.0391029
R1881 vss.n2398 vss.n2397 0.0391029
R1882 vss.n2368 vss.n2367 0.0391029
R1883 vss.n2379 vss.n2378 0.0391029
R1884 vss.n2357 vss.n2356 0.0391029
R1885 vss.n2361 vss.n2360 0.0391029
R1886 vss.n2333 vss.n2332 0.0391029
R1887 vss.n2748 vss.n2744 0.0391029
R1888 vss.n2743 vss.n2742 0.0391029
R1889 vss.n2741 vss.n2740 0.0391029
R1890 vss.n2739 vss.n2738 0.0391029
R1891 vss.n2737 vss.n2733 0.0391029
R1892 vss.n2796 vss.n2791 0.0391029
R1893 vss.n2752 vss.n2751 0.0391029
R1894 vss.n2767 vss.n2763 0.0391029
R1895 vss.n2766 vss.n2765 0.0391029
R1896 vss.n2781 vss.n2777 0.0391029
R1897 vss.n2780 vss.n2779 0.0391029
R1898 vss.n2798 vss.n2790 0.0391029
R1899 vss.n1829 vss.n1828 0.0391029
R1900 vss.n1840 vss.n1837 0.0391029
R1901 vss.n1839 vss.n1838 0.0391029
R1902 vss.n1861 vss.n1849 0.0391029
R1903 vss.n1852 vss.n1851 0.0391029
R1904 vss.n1808 vss.n1802 0.0391029
R1905 vss.n2823 vss.n2822 0.0391029
R1906 vss.n2825 vss.n2824 0.0391029
R1907 vss.n2838 vss.n2837 0.0391029
R1908 vss.n2836 vss.n2835 0.0391029
R1909 vss.n2834 vss.n2833 0.0391029
R1910 vss.n2832 vss.n2831 0.0391029
R1911 vss.n189 vss.n188 0.0391029
R1912 vss.n185 vss.n184 0.0391029
R1913 vss.n183 vss.n182 0.0391029
R1914 vss.n179 vss.n178 0.0391029
R1915 vss.n177 vss.n176 0.0391029
R1916 vss.n173 vss.n172 0.0391029
R1917 vss.n3323 vss.n3247 0.0388652
R1918 vss.n3120 vss.n3119 0.0384032
R1919 vss.n2882 vss.n2881 0.0383889
R1920 vss.n7 vss.n5 0.0383698
R1921 vss.n7 vss.n6 0.0383698
R1922 vss.n28 vss.n26 0.0383698
R1923 vss.n28 vss.n27 0.0383698
R1924 vss.n34 vss.n32 0.0383698
R1925 vss.n34 vss.n33 0.0383698
R1926 vss.n59 vss.n57 0.0383698
R1927 vss.n59 vss.n58 0.0383698
R1928 vss.n68 vss.n67 0.0383698
R1929 vss.n69 vss.n68 0.0383698
R1930 vss.n71 vss.n69 0.0383698
R1931 vss.n71 vss.n70 0.0383698
R1932 vss.n75 vss.n74 0.0383698
R1933 vss.n1140 vss 0.0378217
R1934 vss.n2124 vss 0.0378217
R1935 vss.n23 vss.n22 0.0376094
R1936 vss.n1183 vss.n1182 0.0376053
R1937 vss.n125 vss.n124 0.0375879
R1938 vss.n3173 vss.n3172 0.0369063
R1939 vss.n3124 vss.n3120 0.0367903
R1940 vss.n583 vss.n582 0.0361962
R1941 vss.n1990 vss.n1989 0.0361962
R1942 vss.n2966 vss.n2888 0.0359839
R1943 vss.n2899 vss.n2898 0.035973
R1944 vss.n2928 vss.n2900 0.035973
R1945 vss.n617 vss.n616 0.035973
R1946 vss.n619 vss.n618 0.035973
R1947 vss.n1208 vss.n1120 0.035973
R1948 vss.n1207 vss.n1122 0.035973
R1949 vss.n593 vss.n578 0.035973
R1950 vss.n580 vss.n579 0.035973
R1951 vss.n1227 vss.n1226 0.035918
R1952 vss vss.n486 0.0358842
R1953 vss.n17 vss.n3 0.0356562
R1954 vss.n15 vss.n14 0.0356562
R1955 vss.n81 vss.n53 0.0356562
R1956 vss.n1986 vss.n635 0.0345671
R1957 vss.n1139 vss.n1130 0.0343542
R1958 vss.n2126 vss.n2125 0.0343542
R1959 vss vss.n1796 0.034115
R1960 vss.n1705 vss 0.0338434
R1961 vss.n3091 vss.n3085 0.0335645
R1962 vss.n2911 vss 0.0330521
R1963 vss vss.n1128 0.0330521
R1964 vss vss.n2118 0.0330521
R1965 vss vss.n605 0.0330521
R1966 vss.n3246 vss.n3245 0.032623
R1967 vss.n2957 vss.n2951 0.0325946
R1968 vss.n1994 vss.n622 0.0325946
R1969 vss.n1187 vss.n1186 0.0325946
R1970 vss.n556 vss.n555 0.0325946
R1971 vss.n690 vss 0.0325669
R1972 vss vss.n2930 0.03175
R1973 vss.n2015 vss 0.03175
R1974 vss.n1694 vss 0.0299577
R1975 vss.n62 vss.n61 0.0299384
R1976 vss.n1184 vss.n1180 0.029875
R1977 vss.n588 vss.n587 0.029875
R1978 vss.n633 vss.n632 0.029875
R1979 vss vss.n2285 0.0298356
R1980 vss.n2402 vss 0.0298356
R1981 vss vss.n2274 0.0298356
R1982 vss.n2515 vss 0.0298356
R1983 vss.n2803 vss 0.0298356
R1984 vss vss.n2801 0.0298356
R1985 vss vss.n1941 0.0297375
R1986 vss vss.n720 0.0297375
R1987 vss.n788 vss 0.0297375
R1988 vss vss.n1453 0.0297375
R1989 vss.n1217 vss 0.0285374
R1990 vss.n2136 vss 0.0285374
R1991 vss.n3326 vss 0.0278851
R1992 vss.n2930 vss.n2929 0.0278438
R1993 vss.n1195 vss.n1121 0.0278438
R1994 vss.n594 vss.n577 0.0278438
R1995 vss.n2016 vss.n2015 0.0278438
R1996 vss.n3293 vss 0.0278438
R1997 vss.n3295 vss 0.0278438
R1998 vss.n3171 vss.n3170 0.0272993
R1999 vss.n487 vss 0.0272339
R2000 vss.n2646 vss 0.0272339
R2001 vss vss.n207 0.0272339
R2002 vss vss.n2635 0.0272339
R2003 vss.n330 vss 0.0272339
R2004 vss.n3076 vss.n3075 0.0271129
R2005 vss vss.n1227 0.0269789
R2006 vss.n2514 vss.n2513 0.0266812
R2007 vss.n2881 vss 0.0263989
R2008 vss.n3246 vss 0.0261458
R2009 vss.n131 vss.n130 0.0257686
R2010 vss.n1947 vss.n1946 0.0257686
R2011 vss vss.n1312 0.0256931
R2012 vss.n982 vss 0.0256931
R2013 vss vss.n1704 0.0256931
R2014 vss vss.n1985 0.0256931
R2015 vss.n1797 vss 0.0256931
R2016 vss.n475 vss.n401 0.025078
R2017 vss.n3237 vss.n3207 0.0247248
R2018 vss vss.n652 0.024393
R2019 vss.n1220 vss.n1219 0.0241592
R2020 vss.n2139 vss.n2138 0.0241592
R2021 vss vss.n139 0.0240791
R2022 vss.n774 vss.n773 0.024008
R2023 vss.n2062 vss.n2061 0.024008
R2024 vss.n639 vss.n638 0.024008
R2025 vss.n3255 vss.n3254 0.024008
R2026 vss.n3222 vss.n3221 0.0231378
R2027 vss vss.n3326 0.0229802
R2028 vss.n1867 vss.n1865 0.0227182
R2029 vss.n37 vss.n36 0.022692
R2030 vss.n2916 vss.n2915 0.0226661
R2031 vss.n2917 vss.n2916 0.0226661
R2032 vss.n2960 vss 0.0226354
R2033 vss.n1206 vss.n1123 0.0226354
R2034 vss.n2117 vss.n2116 0.0226354
R2035 vss.n620 vss 0.0226354
R2036 vss.n133 vss.n132 0.0223823
R2037 vss.n1945 vss.n684 0.0223823
R2038 vss vss.n3010 0.0222742
R2039 vss.n3215 vss.n3214 0.0221535
R2040 vss.n211 vss.n209 0.0219755
R2041 vss.n294 vss.n293 0.0219755
R2042 vss.n2875 vss.n2874 0.0219755
R2043 vss.n1902 vss.n1901 0.0219755
R2044 vss.n1718 vss.n1709 0.0219755
R2045 vss.n1339 vss.n1337 0.0219755
R2046 vss.n732 vss.n731 0.0219755
R2047 vss.n1472 vss.n1470 0.0219755
R2048 vss.n1563 vss.n1562 0.0219755
R2049 vss.n1250 vss.n737 0.0219755
R2050 vss.n740 vss.n739 0.0219755
R2051 vss.n792 vss.n790 0.0219755
R2052 vss.n1056 vss.n1037 0.0219755
R2053 vss.n1318 vss.n1315 0.0219755
R2054 vss.n922 vss.n921 0.0219755
R2055 vss.n976 vss.n967 0.0219755
R2056 vss.n1675 vss.n1674 0.0219755
R2057 vss.n1981 vss.n1980 0.0219755
R2058 vss.n2104 vss.n2026 0.0219755
R2059 vss.n2163 vss.n2161 0.0219755
R2060 vss.n2518 vss.n445 0.0219755
R2061 vss.n473 vss.n465 0.0219755
R2062 vss.n405 vss.n403 0.0219755
R2063 vss.n2599 vss.n2598 0.0219755
R2064 vss.n2602 vss.n2600 0.0219755
R2065 vss.n2700 vss.n2699 0.0219755
R2066 vss.n2289 vss.n2287 0.0219755
R2067 vss.n2414 vss.n2413 0.0219755
R2068 vss.n2398 vss.n2389 0.0219755
R2069 vss.n2798 vss.n2797 0.0219755
R2070 vss.n1808 vss.n1803 0.0219755
R2071 vss.n172 vss.n171 0.0219755
R2072 vss.n114 vss.n111 0.0219646
R2073 vss.n3230 vss.n3229 0.0219646
R2074 vss.n49 vss.n48 0.0219591
R2075 vss.n10 vss.n9 0.0217862
R2076 vss.n3194 vss.n3193 0.0216694
R2077 vss.n2903 vss.n2897 0.0213333
R2078 vss.n1189 vss.n1188 0.0213333
R2079 vss.n557 vss.n553 0.0213333
R2080 vss.n2017 vss.n615 0.0213333
R2081 vss.n2884 vss.n105 0.0212995
R2082 vss.n2148 vss.n2147 0.0211532
R2083 vss.n3109 vss.n3108 0.0206613
R2084 vss.n1622 vss 0.0201488
R2085 vss.n2958 vss.n2950 0.0200312
R2086 vss.n1996 vss.n1995 0.0200312
R2087 vss.n2318 vss 0.0194262
R2088 vss vss.n2401 0.0194262
R2089 vss.n2275 vss 0.0194262
R2090 vss.n1551 vss 0.0193629
R2091 vss.n1454 vss 0.0193629
R2092 vss vss.n1621 0.0193629
R2093 vss.n3326 vss.n3324 0.0192184
R2094 vss.n212 vss.n208 0.0191618
R2095 vss.n213 vss.n212 0.0191618
R2096 vss.n223 vss.n216 0.0191618
R2097 vss.n224 vss.n223 0.0191618
R2098 vss.n234 vss.n227 0.0191618
R2099 vss.n235 vss.n234 0.0191618
R2100 vss.n346 vss.n238 0.0191618
R2101 vss.n346 vss.n345 0.0191618
R2102 vss.n342 vss.n341 0.0191618
R2103 vss.n341 vss.n328 0.0191618
R2104 vss.n325 vss.n324 0.0191618
R2105 vss.n324 vss.n323 0.0191618
R2106 vss.n320 vss.n319 0.0191618
R2107 vss.n319 vss.n318 0.0191618
R2108 vss.n315 vss.n314 0.0191618
R2109 vss.n314 vss.n313 0.0191618
R2110 vss.n145 vss.n144 0.0191618
R2111 vss.n146 vss.n145 0.0191618
R2112 vss.n149 vss.n148 0.0191618
R2113 vss.n150 vss.n149 0.0191618
R2114 vss.n2876 vss.n152 0.0191618
R2115 vss.n1921 vss.n689 0.0191618
R2116 vss.n1922 vss.n1921 0.0191618
R2117 vss.n1925 vss.n1924 0.0191618
R2118 vss.n1926 vss.n1925 0.0191618
R2119 vss.n1936 vss.n1929 0.0191618
R2120 vss.n1936 vss.n1935 0.0191618
R2121 vss.n1932 vss.n1931 0.0191618
R2122 vss.n1931 vss.n1930 0.0191618
R2123 vss.n1719 vss.n1706 0.0191618
R2124 vss.n1719 vss.n1708 0.0191618
R2125 vss.n1733 vss.n1724 0.0191618
R2126 vss.n1733 vss.n1732 0.0191618
R2127 vss.n1747 vss.n1738 0.0191618
R2128 vss.n1747 vss.n1746 0.0191618
R2129 vss.n1779 vss.n1752 0.0191618
R2130 vss.n1779 vss.n1778 0.0191618
R2131 vss.n1831 vss.n1814 0.0191618
R2132 vss.n1832 vss.n1831 0.0191618
R2133 vss.n1841 vss.n1834 0.0191618
R2134 vss.n1842 vss.n1841 0.0191618
R2135 vss.n1862 vss.n1844 0.0191618
R2136 vss.n1862 vss.n1846 0.0191618
R2137 vss.n1809 vss.n1799 0.0191618
R2138 vss.n1809 vss.n1800 0.0191618
R2139 vss.n1340 vss.n1336 0.0191618
R2140 vss.n1341 vss.n1340 0.0191618
R2141 vss.n1351 vss.n1344 0.0191618
R2142 vss.n1352 vss.n1351 0.0191618
R2143 vss.n1362 vss.n1355 0.0191618
R2144 vss.n1363 vss.n1362 0.0191618
R2145 vss.n1451 vss.n1366 0.0191618
R2146 vss.n1451 vss.n1450 0.0191618
R2147 vss.n1447 vss.n1446 0.0191618
R2148 vss.n1446 vss.n1445 0.0191618
R2149 vss.n1442 vss.n1441 0.0191618
R2150 vss.n1441 vss.n1440 0.0191618
R2151 vss.n1437 vss.n1436 0.0191618
R2152 vss.n1436 vss.n1435 0.0191618
R2153 vss.n1465 vss.n721 0.0191618
R2154 vss.n1466 vss.n1465 0.0191618
R2155 vss.n1473 vss.n1469 0.0191618
R2156 vss.n1474 vss.n1473 0.0191618
R2157 vss.n1484 vss.n1477 0.0191618
R2158 vss.n1485 vss.n1484 0.0191618
R2159 vss.n1495 vss.n1488 0.0191618
R2160 vss.n1496 vss.n1495 0.0191618
R2161 vss.n1609 vss.n1499 0.0191618
R2162 vss.n1609 vss.n1608 0.0191618
R2163 vss.n1605 vss.n1604 0.0191618
R2164 vss.n1604 vss.n1550 0.0191618
R2165 vss.n1599 vss.n1590 0.0191618
R2166 vss.n1599 vss.n1598 0.0191618
R2167 vss.n1585 vss.n1570 0.0191618
R2168 vss.n1585 vss.n1584 0.0191618
R2169 vss.n1565 vss.n1553 0.0191618
R2170 vss.n1565 vss.n1564 0.0191618
R2171 vss.n1251 vss.n734 0.0191618
R2172 vss.n1251 vss.n736 0.0191618
R2173 vss.n1271 vss.n1256 0.0191618
R2174 vss.n1271 vss.n1270 0.0191618
R2175 vss.n1285 vss.n1276 0.0191618
R2176 vss.n1285 vss.n1284 0.0191618
R2177 vss.n1310 vss.n1290 0.0191618
R2178 vss.n1310 vss.n1309 0.0191618
R2179 vss.n759 vss.n758 0.0191618
R2180 vss.n760 vss.n759 0.0191618
R2181 vss.n763 vss.n762 0.0191618
R2182 vss.n764 vss.n763 0.0191618
R2183 vss.n767 vss.n766 0.0191618
R2184 vss.n768 vss.n767 0.0191618
R2185 vss.n1233 vss.n770 0.0191618
R2186 vss.n793 vss.n789 0.0191618
R2187 vss.n794 vss.n793 0.0191618
R2188 vss.n804 vss.n797 0.0191618
R2189 vss.n805 vss.n804 0.0191618
R2190 vss.n815 vss.n808 0.0191618
R2191 vss.n816 vss.n815 0.0191618
R2192 vss.n1102 vss.n819 0.0191618
R2193 vss.n1102 vss.n1101 0.0191618
R2194 vss.n1098 vss.n1097 0.0191618
R2195 vss.n1041 vss.n1040 0.0191618
R2196 vss.n1042 vss.n1041 0.0191618
R2197 vss.n1045 vss.n1044 0.0191618
R2198 vss.n1046 vss.n1045 0.0191618
R2199 vss.n1055 vss.n1048 0.0191618
R2200 vss.n879 vss.n873 0.0191618
R2201 vss.n880 vss.n879 0.0191618
R2202 vss.n889 vss.n882 0.0191618
R2203 vss.n890 vss.n889 0.0191618
R2204 vss.n1020 vss.n892 0.0191618
R2205 vss.n1020 vss.n1019 0.0191618
R2206 vss.n1016 vss.n1015 0.0191618
R2207 vss.n1015 vss.n998 0.0191618
R2208 vss.n995 vss.n994 0.0191618
R2209 vss.n994 vss.n993 0.0191618
R2210 vss.n990 vss.n989 0.0191618
R2211 vss.n989 vss.n988 0.0191618
R2212 vss.n985 vss.n984 0.0191618
R2213 vss.n984 vss.n923 0.0191618
R2214 vss.n979 vss.n966 0.0191618
R2215 vss.n979 vss.n978 0.0191618
R2216 vss.n960 vss.n951 0.0191618
R2217 vss.n960 vss.n959 0.0191618
R2218 vss.n945 vss.n936 0.0191618
R2219 vss.n945 vss.n944 0.0191618
R2220 vss.n1625 vss.n693 0.0191618
R2221 vss.n1626 vss.n1625 0.0191618
R2222 vss.n1692 vss.n1629 0.0191618
R2223 vss.n1692 vss.n1691 0.0191618
R2224 vss.n1688 vss.n1687 0.0191618
R2225 vss.n1687 vss.n1686 0.0191618
R2226 vss.n1683 vss.n1682 0.0191618
R2227 vss.n1682 vss.n1681 0.0191618
R2228 vss.n1678 vss.n1677 0.0191618
R2229 vss.n1677 vss.n1676 0.0191618
R2230 vss.n681 vss.n680 0.0191618
R2231 vss.n658 vss.n657 0.0191618
R2232 vss.n659 vss.n658 0.0191618
R2233 vss.n663 vss.n662 0.0191618
R2234 vss.n664 vss.n663 0.0191618
R2235 vss.n1983 vss.n667 0.0191618
R2236 vss.n1983 vss.n1982 0.0191618
R2237 vss.n2103 vss.n2102 0.0191618
R2238 vss.n2084 vss.n2083 0.0191618
R2239 vss.n2096 vss.n2086 0.0191618
R2240 vss.n2096 vss.n2088 0.0191618
R2241 vss.n2058 vss.n2031 0.0191618
R2242 vss.n2058 vss.n2032 0.0191618
R2243 vss.n2164 vss.n2160 0.0191618
R2244 vss.n2165 vss.n2164 0.0191618
R2245 vss.n2175 vss.n2168 0.0191618
R2246 vss.n2176 vss.n2175 0.0191618
R2247 vss.n2186 vss.n2179 0.0191618
R2248 vss.n2187 vss.n2186 0.0191618
R2249 vss.n2272 vss.n2190 0.0191618
R2250 vss.n2272 vss.n2240 0.0191618
R2251 vss.n2237 vss.n2236 0.0191618
R2252 vss.n450 vss.n449 0.0191618
R2253 vss.n451 vss.n450 0.0191618
R2254 vss.n455 vss.n454 0.0191618
R2255 vss.n456 vss.n455 0.0191618
R2256 vss.n2517 vss.n459 0.0191618
R2257 vss.n2517 vss.n460 0.0191618
R2258 vss.n474 vss.n462 0.0191618
R2259 vss.n474 vss.n464 0.0191618
R2260 vss.n545 vss.n531 0.0191618
R2261 vss.n545 vss.n544 0.0191618
R2262 vss.n526 vss.n517 0.0191618
R2263 vss.n526 vss.n525 0.0191618
R2264 vss.n512 vss.n489 0.0191618
R2265 vss.n512 vss.n511 0.0191618
R2266 vss.n406 vss.n402 0.0191618
R2267 vss.n407 vss.n406 0.0191618
R2268 vss.n417 vss.n410 0.0191618
R2269 vss.n418 vss.n417 0.0191618
R2270 vss.n428 vss.n421 0.0191618
R2271 vss.n429 vss.n428 0.0191618
R2272 vss.n2537 vss.n432 0.0191618
R2273 vss.n2538 vss.n2537 0.0191618
R2274 vss.n2558 vss.n2541 0.0191618
R2275 vss.n2559 vss.n2558 0.0191618
R2276 vss.n2568 vss.n2561 0.0191618
R2277 vss.n2569 vss.n2568 0.0191618
R2278 vss.n2585 vss.n2571 0.0191618
R2279 vss.n2586 vss.n2585 0.0191618
R2280 vss.n2633 vss.n2588 0.0191618
R2281 vss.n2633 vss.n2632 0.0191618
R2282 vss.n2629 vss.n2628 0.0191618
R2283 vss.n2628 vss.n2627 0.0191618
R2284 vss.n2624 vss.n2623 0.0191618
R2285 vss.n2623 vss.n2622 0.0191618
R2286 vss.n2619 vss.n2618 0.0191618
R2287 vss.n2618 vss.n2617 0.0191618
R2288 vss.n2648 vss.n364 0.0191618
R2289 vss.n2649 vss.n2648 0.0191618
R2290 vss.n2680 vss.n2652 0.0191618
R2291 vss.n2680 vss.n2679 0.0191618
R2292 vss.n2717 vss.n2685 0.0191618
R2293 vss.n2717 vss.n2716 0.0191618
R2294 vss.n2713 vss.n2712 0.0191618
R2295 vss.n2712 vss.n2705 0.0191618
R2296 vss.n2703 vss.n2702 0.0191618
R2297 vss.n2290 vss.n2286 0.0191618
R2298 vss.n2291 vss.n2290 0.0191618
R2299 vss.n2301 vss.n2294 0.0191618
R2300 vss.n2302 vss.n2301 0.0191618
R2301 vss.n2312 vss.n2305 0.0191618
R2302 vss.n2313 vss.n2312 0.0191618
R2303 vss.n2501 vss.n2316 0.0191618
R2304 vss.n2501 vss.n2469 0.0191618
R2305 vss.n2466 vss.n2465 0.0191618
R2306 vss.n2465 vss.n2448 0.0191618
R2307 vss.n2445 vss.n2444 0.0191618
R2308 vss.n2444 vss.n2437 0.0191618
R2309 vss.n2434 vss.n2433 0.0191618
R2310 vss.n2433 vss.n2419 0.0191618
R2311 vss.n2416 vss.n2415 0.0191618
R2312 vss.n2415 vss.n2317 0.0191618
R2313 vss.n2399 vss.n2386 0.0191618
R2314 vss.n2399 vss.n2388 0.0191618
R2315 vss.n2380 vss.n2329 0.0191618
R2316 vss.n2380 vss.n2365 0.0191618
R2317 vss.n2363 vss.n2362 0.0191618
R2318 vss.n2362 vss.n2351 0.0191618
R2319 vss.n2349 vss.n2348 0.0191618
R2320 vss.n2348 vss.n2331 0.0191618
R2321 vss.n2754 vss.n2727 0.0191618
R2322 vss.n2754 vss.n2729 0.0191618
R2323 vss.n2768 vss.n2759 0.0191618
R2324 vss.n2768 vss.n2761 0.0191618
R2325 vss.n2782 vss.n2773 0.0191618
R2326 vss.n2782 vss.n2775 0.0191618
R2327 vss.n2799 vss.n2787 0.0191618
R2328 vss.n2799 vss.n2788 0.0191618
R2329 vss.n2814 vss.n190 0.0191618
R2330 vss.n2814 vss.n206 0.0191618
R2331 vss.n203 vss.n202 0.0191618
R2332 vss.n202 vss.n201 0.0191618
R2333 vss.n198 vss.n197 0.0191618
R2334 vss.n197 vss.n196 0.0191618
R2335 vss.n193 vss.n192 0.0191618
R2336 vss.n192 vss.n191 0.0191618
R2337 vss.n1182 vss.n1118 0.0190526
R2338 vss.n1118 vss.n1116 0.0190526
R2339 vss vss.n690 0.0189314
R2340 vss.n2149 vss.n2148 0.0186413
R2341 vss.n1324 vss 0.0185144
R2342 vss.n582 vss.n581 0.0183481
R2343 vss.n581 vss.n551 0.0183481
R2344 vss.n1988 vss.n1987 0.0183481
R2345 vss.n1989 vss.n1988 0.0183481
R2346 vss.n115 vss.n114 0.0181768
R2347 vss.n2636 vss 0.0177477
R2348 vss vss.n363 0.0177477
R2349 vss.n329 vss 0.0177477
R2350 vss.n117 vss 0.0176371
R2351 vss.n3263 vss.n3248 0.0175415
R2352 vss.n1219 vss.n1218 0.0173735
R2353 vss.n2138 vss.n2137 0.0173735
R2354 vss.n3207 vss.n3205 0.0169729
R2355 vss.n924 vss 0.0167536
R2356 vss vss.n981 0.0167536
R2357 vss.n3190 vss 0.016562
R2358 vss.n81 vss.n54 0.016125
R2359 vss.n18 vss.n1 0.0157892
R2360 vss.n18 vss.n2 0.0157892
R2361 vss.n3159 vss.n3158 0.0156732
R2362 vss.n135 vss.n134 0.0156071
R2363 vss.n3212 vss.n3210 0.0156071
R2364 vss.n3196 vss.n108 0.0156071
R2365 vss.n3240 vss.n3200 0.0156071
R2366 vss.n3004 vss.n3003 0.0156071
R2367 vss.n3000 vss.n2999 0.0156071
R2368 vss.n2996 vss.n2995 0.0156071
R2369 vss.n2992 vss.n2991 0.0156071
R2370 vss.n2988 vss.n2987 0.0156071
R2371 vss.n2980 vss.n2979 0.0156071
R2372 vss.n3134 vss.n2887 0.0156071
R2373 vss.n2968 vss.n2967 0.0156071
R2374 vss.n2972 vss.n2971 0.0156071
R2375 vss.n2976 vss.n2975 0.0156071
R2376 vss.n2984 vss.n2983 0.0156071
R2377 vss.n647 vss.n646 0.0156071
R2378 vss.n1224 vss.n1223 0.0156071
R2379 vss.n783 vss.n782 0.0156071
R2380 vss.n778 vss.n777 0.0156071
R2381 vss.n1944 vss.n686 0.0156071
R2382 vss.n1944 vss.n687 0.0156071
R2383 vss.n2143 vss.n2142 0.0156071
R2384 vss.n2071 vss.n2070 0.0156071
R2385 vss.n2066 vss.n2065 0.0156071
R2386 vss.n642 vss.n636 0.0156071
R2387 vss.n3268 vss.n3267 0.0156071
R2388 vss.n3258 vss.n3252 0.0156071
R2389 vss.n3285 vss.n3274 0.0156071
R2390 vss.n3306 vss.n3249 0.0156071
R2391 vss.n3320 vss.n3310 0.0156071
R2392 vss.n3290 vss.n3251 0.0156071
R2393 vss.n101 vss.n84 0.0156071
R2394 vss.n101 vss.n85 0.0156071
R2395 vss.n82 vss.n51 0.0156071
R2396 vss.n82 vss.n52 0.0156071
R2397 vss.n45 vss.n20 0.0156071
R2398 vss.n45 vss.n44 0.0156071
R2399 vss.n3324 vss.n3323 0.0155019
R2400 vss.n3165 vss.n3164 0.0153957
R2401 vss.n3067 vss.n3066 0.0150161
R2402 vss.n2721 vss.n362 0.0149953
R2403 vss.n3193 vss.n3190 0.0146702
R2404 vss.n3156 vss.n3155 0.014378
R2405 vss.n215 vss.n214 0.0143235
R2406 vss.n226 vss.n225 0.0143235
R2407 vss.n237 vss.n236 0.0143235
R2408 vss.n327 vss.n326 0.0143235
R2409 vss.n322 vss.n321 0.0143235
R2410 vss.n317 vss.n316 0.0143235
R2411 vss.n1928 vss.n1927 0.0143235
R2412 vss.n1934 vss.n1933 0.0143235
R2413 vss.n1343 vss.n1342 0.0143235
R2414 vss.n1354 vss.n1353 0.0143235
R2415 vss.n1365 vss.n1364 0.0143235
R2416 vss.n1444 vss.n1443 0.0143235
R2417 vss.n1439 vss.n1438 0.0143235
R2418 vss.n1434 vss.n1433 0.0143235
R2419 vss.n1476 vss.n1475 0.0143235
R2420 vss.n1487 vss.n1486 0.0143235
R2421 vss.n1498 vss.n1497 0.0143235
R2422 vss.n796 vss.n795 0.0143235
R2423 vss.n807 vss.n806 0.0143235
R2424 vss.n818 vss.n817 0.0143235
R2425 vss.n997 vss.n996 0.0143235
R2426 vss.n992 vss.n991 0.0143235
R2427 vss.n987 vss.n986 0.0143235
R2428 vss.n1690 vss.n1689 0.0143235
R2429 vss.n1685 vss.n1684 0.0143235
R2430 vss.n1680 vss.n1679 0.0143235
R2431 vss.n656 vss.n655 0.0143235
R2432 vss.n661 vss.n660 0.0143235
R2433 vss.n666 vss.n665 0.0143235
R2434 vss.n2167 vss.n2166 0.0143235
R2435 vss.n2178 vss.n2177 0.0143235
R2436 vss.n2189 vss.n2188 0.0143235
R2437 vss.n448 vss.n447 0.0143235
R2438 vss.n453 vss.n452 0.0143235
R2439 vss.n458 vss.n457 0.0143235
R2440 vss.n409 vss.n408 0.0143235
R2441 vss.n420 vss.n419 0.0143235
R2442 vss.n431 vss.n430 0.0143235
R2443 vss.n2626 vss.n2625 0.0143235
R2444 vss.n2621 vss.n2620 0.0143235
R2445 vss.n2616 vss.n2615 0.0143235
R2446 vss.n2715 vss.n2714 0.0143235
R2447 vss.n2293 vss.n2292 0.0143235
R2448 vss.n2304 vss.n2303 0.0143235
R2449 vss.n2315 vss.n2314 0.0143235
R2450 vss.n2447 vss.n2446 0.0143235
R2451 vss.n2436 vss.n2435 0.0143235
R2452 vss.n2418 vss.n2417 0.0143235
R2453 vss.n205 vss.n204 0.0143235
R2454 vss.n200 vss.n199 0.0143235
R2455 vss.n195 vss.n194 0.0143235
R2456 vss.n130 vss.n129 0.0142993
R2457 vss.n1948 vss.n1947 0.0142993
R2458 vss.n3221 vss.n3219 0.0142795
R2459 vss.n3057 vss.n3056 0.0142097
R2460 vss.n3162 vss.n3161 0.0140079
R2461 vss.n1864 vss.n1787 0.0138065
R2462 vss.n3144 vss.n3143 0.0137303
R2463 vss.n775 vss.n774 0.0137243
R2464 vss.n2063 vss.n2062 0.0137243
R2465 vss.n640 vss.n639 0.0137243
R2466 vss.n3256 vss.n3255 0.0137243
R2467 vss.n2915 vss.n2914 0.0137188
R2468 vss.n2927 vss.n2917 0.0137188
R2469 vss.n2927 vss.n2919 0.0137188
R2470 vss.n2956 vss.n2954 0.0137188
R2471 vss.n2956 vss.n2955 0.0137188
R2472 vss.n1185 vss.n1115 0.0137188
R2473 vss.n1209 vss.n1117 0.0137188
R2474 vss.n1209 vss.n1119 0.0137188
R2475 vss.n586 vss.n585 0.0137188
R2476 vss.n592 vss.n589 0.0137188
R2477 vss.n592 vss.n591 0.0137188
R2478 vss.n626 vss.n625 0.0137188
R2479 vss.n630 vss.n629 0.0137188
R2480 vss.n631 vss.n630 0.0137188
R2481 vss.n1992 vss.n634 0.0137188
R2482 vss.n3153 vss.n3152 0.0136378
R2483 vss.n3275 vss 0.0136173
R2484 vss.n2949 vss.n2935 0.0135208
R2485 vss.n1193 vss.n1145 0.0135208
R2486 vss.n572 vss.n571 0.0135208
R2487 vss.n2010 vss.n2009 0.0135208
R2488 vss.n3278 vss 0.0135208
R2489 vss vss.n105 0.0134853
R2490 vss.n3011 vss 0.0134032
R2491 vss.n1864 vss 0.0133674
R2492 vss.n3150 vss.n3149 0.0133602
R2493 vss vss.n2514 0.0131493
R2494 vss.n3229 vss.n3224 0.0131263
R2495 vss.n1135 vss.n1134 0.0130393
R2496 vss.n2129 vss.n552 0.0130393
R2497 vss vss.n3294 0.013
R2498 vss.n1864 vss.n1782 0.0128256
R2499 vss vss.n117 0.0125968
R2500 vss.n3100 vss.n3096 0.0125968
R2501 vss.n2957 vss.n2952 0.0123243
R2502 vss.n1994 vss.n1993 0.0123243
R2503 vss.n1187 vss.n1179 0.0123243
R2504 vss.n556 vss.n554 0.0123243
R2505 vss.n17 vss.n16 0.0122188
R2506 vss.n131 vss 0.0121822
R2507 vss.n1946 vss 0.0121822
R2508 vss.n401 vss.n400 0.0121325
R2509 vss.n3235 vss.n3232 0.0121279
R2510 vss vss.n358 0.012067
R2511 vss.n3147 vss.n3146 0.012065
R2512 vss.n3141 vss.n3140 0.012065
R2513 vss.n3138 vss.n3137 0.012065
R2514 vss.n139 vss.n138 0.0118873
R2515 vss.n127 vss.n126 0.0116721
R2516 vss.n308 vss.n307 0.0115294
R2517 vss.n302 vss.n301 0.0115294
R2518 vss.n296 vss.n295 0.0115294
R2519 vss.n161 vss.n160 0.0115294
R2520 vss.n2861 vss.n2860 0.0115294
R2521 vss.n157 vss.n156 0.0115294
R2522 vss.n1916 vss.n1915 0.0115294
R2523 vss.n1910 vss.n1909 0.0115294
R2524 vss.n1904 vss.n1903 0.0115294
R2525 vss.n1717 vss.n1716 0.0115294
R2526 vss.n1729 vss.n1728 0.0115294
R2527 vss.n1743 vss.n1742 0.0115294
R2528 vss.n1416 vss.n1415 0.0115294
R2529 vss.n1422 vss.n1421 0.0115294
R2530 vss.n724 vss.n723 0.0115294
R2531 vss.n1592 vss.n1591 0.0115294
R2532 vss.n1572 vss.n1571 0.0115294
R2533 vss.n1555 vss.n1554 0.0115294
R2534 vss.n1249 vss.n1248 0.0115294
R2535 vss.n1267 vss.n1266 0.0115294
R2536 vss.n1281 vss.n1280 0.0115294
R2537 vss.n742 vss.n741 0.0115294
R2538 vss.n748 vss.n747 0.0115294
R2539 vss.n754 vss.n753 0.0115294
R2540 vss.n1092 vss.n1091 0.0115294
R2541 vss.n857 vss.n856 0.0115294
R2542 vss.n1036 vss.n1035 0.0115294
R2543 vss.n1317 vss.n1316 0.0115294
R2544 vss.n895 vss.n894 0.0115294
R2545 vss.n901 vss.n900 0.0115294
R2546 vss.n914 vss.n913 0.0115294
R2547 vss.n975 vss.n974 0.0115294
R2548 vss.n956 vss.n955 0.0115294
R2549 vss.n941 vss.n940 0.0115294
R2550 vss.n676 vss.n675 0.0115294
R2551 vss.n1966 vss.n1965 0.0115294
R2552 vss.n672 vss.n671 0.0115294
R2553 vss.n2029 vss.n2028 0.0115294
R2554 vss.n2094 vss.n2093 0.0115294
R2555 vss.n2231 vss.n2230 0.0115294
R2556 vss.n2196 vss.n2195 0.0115294
R2557 vss.n444 vss.n443 0.0115294
R2558 vss.n472 vss.n471 0.0115294
R2559 vss.n541 vss.n540 0.0115294
R2560 vss.n522 vss.n521 0.0115294
R2561 vss.n2564 vss.n2563 0.0115294
R2562 vss.n2574 vss.n2573 0.0115294
R2563 vss.n2591 vss.n2590 0.0115294
R2564 vss.n2687 vss.n2686 0.0115294
R2565 vss.n2440 vss.n2439 0.0115294
R2566 vss.n2422 vss.n2421 0.0115294
R2567 vss.n2406 vss.n2405 0.0115294
R2568 vss.n2397 vss.n2396 0.0115294
R2569 vss.n2378 vss.n2377 0.0115294
R2570 vss.n2360 vss.n2359 0.0115294
R2571 vss.n2763 vss.n2762 0.0115294
R2572 vss.n2777 vss.n2776 0.0115294
R2573 vss.n2790 vss.n2789 0.0115294
R2574 vss.n1837 vss.n1836 0.0115294
R2575 vss.n1849 vss.n1848 0.0115294
R2576 vss.n1802 vss.n1801 0.0115294
R2577 vss.n186 vss.n185 0.0115294
R2578 vss.n180 vss.n179 0.0115294
R2579 vss.n174 vss.n173 0.0115294
R2580 vss.n3289 vss.n3288 0.0115156
R2581 vss.n2881 vss.n2880 0.0115
R2582 vss.n1217 vss.n1216 0.0113696
R2583 vss.n2136 vss.n2135 0.0113696
R2584 vss.n3287 vss.n3286 0.0113462
R2585 vss.n1222 vss.n1221 0.0107133
R2586 vss.n2141 vss.n2140 0.0107133
R2587 vss.n3282 vss 0.0105309
R2588 vss.n269 vss.n268 0.0104679
R2589 vss.n1776 vss.n1775 0.0104679
R2590 vss.n1397 vss.n1396 0.0104679
R2591 vss.n1530 vss.n1529 0.0104679
R2592 vss.n1308 vss.n1307 0.0104679
R2593 vss.n1235 vss.n1234 0.0104679
R2594 vss.n851 vss.n850 0.0104679
R2595 vss.n1022 vss.n1021 0.0104679
R2596 vss.n717 vss.n716 0.0104679
R2597 vss.n2057 vss.n2056 0.0104679
R2598 vss.n510 vss.n509 0.0104679
R2599 vss.n2536 vss.n2535 0.0104679
R2600 vss.n395 vss.n394 0.0104679
R2601 vss.n2500 vss.n2499 0.0104679
R2602 vss.n2347 vss.n2346 0.0104679
R2603 vss vss.n1867 0.0102662
R2604 vss.n3195 vss.n109 0.0102656
R2605 vss.n1324 vss.n1323 0.010166
R2606 vss.n1622 vss.n719 0.0100886
R2607 vss.n2816 vss.n2815 0.0100486
R2608 vss.n99 vss.n98 0.0100109
R2609 vss.n143 vss.n142 0.00997131
R2610 vss.n144 vss.n143 0.00997131
R2611 vss.n147 vss.n146 0.00997131
R2612 vss.n148 vss.n147 0.00997131
R2613 vss.n151 vss.n150 0.00997131
R2614 vss.n152 vss.n151 0.00997131
R2615 vss.n1923 vss.n1922 0.00997131
R2616 vss.n1924 vss.n1923 0.00997131
R2617 vss.n1833 vss.n1832 0.00997131
R2618 vss.n1834 vss.n1833 0.00997131
R2619 vss.n1843 vss.n1842 0.00997131
R2620 vss.n1844 vss.n1843 0.00997131
R2621 vss.n761 vss.n760 0.00997131
R2622 vss.n762 vss.n761 0.00997131
R2623 vss.n765 vss.n764 0.00997131
R2624 vss.n766 vss.n765 0.00997131
R2625 vss.n769 vss.n768 0.00997131
R2626 vss.n770 vss.n769 0.00997131
R2627 vss.n1039 vss.n1038 0.00997131
R2628 vss.n1040 vss.n1039 0.00997131
R2629 vss.n1043 vss.n1042 0.00997131
R2630 vss.n1044 vss.n1043 0.00997131
R2631 vss.n1047 vss.n1046 0.00997131
R2632 vss.n1048 vss.n1047 0.00997131
R2633 vss.n872 vss.n871 0.00997131
R2634 vss.n873 vss.n872 0.00997131
R2635 vss.n881 vss.n880 0.00997131
R2636 vss.n882 vss.n881 0.00997131
R2637 vss.n891 vss.n890 0.00997131
R2638 vss.n892 vss.n891 0.00997131
R2639 vss.n2102 vss.n2101 0.00997131
R2640 vss.n2101 vss.n2100 0.00997131
R2641 vss.n2085 vss.n2084 0.00997131
R2642 vss.n2086 vss.n2085 0.00997131
R2643 vss.n2088 vss.n2087 0.00997131
R2644 vss.n2560 vss.n2559 0.00997131
R2645 vss.n2561 vss.n2560 0.00997131
R2646 vss.n2570 vss.n2569 0.00997131
R2647 vss.n2571 vss.n2570 0.00997131
R2648 vss.n2587 vss.n2586 0.00997131
R2649 vss.n2588 vss.n2587 0.00997131
R2650 vss.n2705 vss.n2704 0.00997131
R2651 vss.n2704 vss.n2703 0.00997131
R2652 vss.n2365 vss.n2364 0.00997131
R2653 vss.n2364 vss.n2363 0.00997131
R2654 vss.n2351 vss.n2350 0.00997131
R2655 vss.n2350 vss.n2349 0.00997131
R2656 vss.n1324 vss 0.00986931
R2657 vss.n312 vss.n292 0.0098203
R2658 vss.n168 vss.n167 0.0098203
R2659 vss.n1920 vss.n1900 0.0098203
R2660 vss.n1548 vss.n1544 0.0098203
R2661 vss.n1413 vss.n1410 0.0098203
R2662 vss.n1096 vss.n1088 0.0098203
R2663 vss.n1660 vss.n1655 0.0098203
R2664 vss.n1014 vss.n1011 0.0098203
R2665 vss.n683 vss.n682 0.0098203
R2666 vss.n2235 vss.n2227 0.0098203
R2667 vss.n2271 vss.n2270 0.0098203
R2668 vss.n2677 vss.n2673 0.0098203
R2669 vss.n2557 vss.n2554 0.0098203
R2670 vss.n2753 vss.n2749 0.0098203
R2671 vss.n2464 vss.n2461 0.0098203
R2672 vss.n1830 vss.n1827 0.0098203
R2673 vss.n2723 vss.n2722 0.00977288
R2674 vss.n219 vss.n218 0.00969118
R2675 vss.n230 vss.n229 0.00969118
R2676 vss.n241 vss.n240 0.00969118
R2677 vss.n310 vss.n309 0.00969118
R2678 vss.n304 vss.n303 0.00969118
R2679 vss.n298 vss.n297 0.00969118
R2680 vss.n163 vss.n162 0.00969118
R2681 vss.n2859 vss.n2858 0.00969118
R2682 vss.n155 vss.n154 0.00969118
R2683 vss.n1918 vss.n1917 0.00969118
R2684 vss.n1912 vss.n1911 0.00969118
R2685 vss.n1906 vss.n1905 0.00969118
R2686 vss.n1726 vss.n1725 0.00969118
R2687 vss.n1740 vss.n1739 0.00969118
R2688 vss.n1754 vss.n1753 0.00969118
R2689 vss.n1347 vss.n1346 0.00969118
R2690 vss.n1358 vss.n1357 0.00969118
R2691 vss.n1369 vss.n1368 0.00969118
R2692 vss.n1480 vss.n1479 0.00969118
R2693 vss.n1491 vss.n1490 0.00969118
R2694 vss.n1502 vss.n1501 0.00969118
R2695 vss.n1546 vss.n1545 0.00969118
R2696 vss.n1594 vss.n1593 0.00969118
R2697 vss.n1580 vss.n1579 0.00969118
R2698 vss.n1258 vss.n1257 0.00969118
R2699 vss.n1278 vss.n1277 0.00969118
R2700 vss.n1292 vss.n1291 0.00969118
R2701 vss.n744 vss.n743 0.00969118
R2702 vss.n750 vss.n749 0.00969118
R2703 vss.n756 vss.n755 0.00969118
R2704 vss.n800 vss.n799 0.00969118
R2705 vss.n811 vss.n810 0.00969118
R2706 vss.n822 vss.n821 0.00969118
R2707 vss.n1094 vss.n1093 0.00969118
R2708 vss.n855 vss.n854 0.00969118
R2709 vss.n1034 vss.n1033 0.00969118
R2710 vss.n875 vss.n874 0.00969118
R2711 vss.n885 vss.n884 0.00969118
R2712 vss.n869 vss.n868 0.00969118
R2713 vss.n953 vss.n952 0.00969118
R2714 vss.n938 vss.n937 0.00969118
R2715 vss.n695 vss.n694 0.00969118
R2716 vss.n1658 vss.n1657 0.00969118
R2717 vss.n1664 vss.n1663 0.00969118
R2718 vss.n1670 vss.n1669 0.00969118
R2719 vss.n678 vss.n677 0.00969118
R2720 vss.n1964 vss.n1963 0.00969118
R2721 vss.n670 vss.n669 0.00969118
R2722 vss.n2091 vss.n2090 0.00969118
R2723 vss.n2034 vss.n2033 0.00969118
R2724 vss.n2171 vss.n2170 0.00969118
R2725 vss.n2182 vss.n2181 0.00969118
R2726 vss.n2243 vss.n2242 0.00969118
R2727 vss.n2233 vss.n2232 0.00969118
R2728 vss.n2194 vss.n2193 0.00969118
R2729 vss.n442 vss.n441 0.00969118
R2730 vss.n533 vss.n532 0.00969118
R2731 vss.n519 vss.n518 0.00969118
R2732 vss.n491 vss.n490 0.00969118
R2733 vss.n413 vss.n412 0.00969118
R2734 vss.n424 vss.n423 0.00969118
R2735 vss.n435 vss.n434 0.00969118
R2736 vss.n2605 vss.n2604 0.00969118
R2737 vss.n2611 vss.n2610 0.00969118
R2738 vss.n367 vss.n366 0.00969118
R2739 vss.n2675 vss.n2674 0.00969118
R2740 vss.n2690 vss.n2689 0.00969118
R2741 vss.n2709 vss.n2708 0.00969118
R2742 vss.n2297 vss.n2296 0.00969118
R2743 vss.n2308 vss.n2307 0.00969118
R2744 vss.n2472 vss.n2471 0.00969118
R2745 vss.n2367 vss.n2366 0.00969118
R2746 vss.n2751 vss.n2750 0.00969118
R2747 vss.n2765 vss.n2764 0.00969118
R2748 vss.n2779 vss.n2778 0.00969118
R2749 vss.n1851 vss.n1850 0.00969118
R2750 vss.n188 vss.n187 0.00969118
R2751 vss.n182 vss.n181 0.00969118
R2752 vss.n176 vss.n175 0.00969118
R2753 vss.n2959 vss.n2958 0.00961458
R2754 vss.n1188 vss.n1178 0.00961458
R2755 vss.n558 vss.n557 0.00961458
R2756 vss.n1995 vss.n621 0.00961458
R2757 vss vss.n3167 0.00938189
R2758 vss vss.n1986 0.009375
R2759 vss.n3224 vss 0.00933838
R2760 vss.n3294 vss.n3293 0.00909375
R2761 vss vss.n691 0.00844366
R2762 vss.n3278 vss 0.0083125
R2763 vss.n3309 vss.n3308 0.00829556
R2764 vss.n40 vss.n39 0.00819928
R2765 vss.n2074 vss.n2069 0.00816304
R2766 vss.n2075 vss.n2074 0.00816304
R2767 vss.n651 vss.n650 0.00816304
R2768 vss.n650 vss.n645 0.00816304
R2769 vss.n1140 vss.n1139 0.00811225
R2770 vss.n2125 vss.n2124 0.00811225
R2771 vss.n1219 vss.n1217 0.00809436
R2772 vss.n2138 vss.n2136 0.00809436
R2773 vss.n2914 vss.n2901 0.00759517
R2774 vss.n1325 vss 0.00759434
R2775 vss.n166 vss.n165 0.0075272
R2776 vss.n1233 vss.n1232 0.0075272
R2777 vss.n1320 vss.n1319 0.0075272
R2778 vss.n1055 vss.n1054 0.0075272
R2779 vss.n2103 vss.n2099 0.0075272
R2780 vss.n2702 vss.n2701 0.0075272
R2781 vss.n2877 vss.n2876 0.0075272
R2782 vss.n3224 vss 0.00738976
R2783 vss.n3286 vss.n3273 0.00736923
R2784 vss.n2923 vss.n2921 0.00709146
R2785 vss.n2904 vss.n2903 0.00701042
R2786 vss.n615 vss.n614 0.00701042
R2787 vss.n3131 vss.n2966 0.00695161
R2788 vss.n13 vss.n12 0.00684058
R2789 vss.n3232 vss.n3231 0.00681313
R2790 vss.n2130 vss.n2129 0.00673148
R2791 vss.n1622 vss 0.00672253
R2792 vss.n1623 vss.n1622 0.00659014
R2793 vss.n1325 vss 0.00647324
R2794 vss vss.n3223 0.00640551
R2795 vss.n80 vss.n79 0.00638768
R2796 vss.n3213 vss.n3208 0.00635938
R2797 vss.n136 vss.n135 0.00635126
R2798 vss.n1224 vss.n1214 0.00635126
R2799 vss.n2144 vss.n2143 0.00635126
R2800 vss.n3241 vss.n3240 0.00635126
R2801 vss.n3018 vss.n3007 0.00614516
R2802 vss.n2925 vss.n2924 0.00605118
R2803 vss.n1226 vss.n1225 0.00603245
R2804 vss.n3197 vss.n3196 0.00601924
R2805 vss.n3212 vss.n3211 0.00601924
R2806 vss.n2147 vss.n2146 0.00591449
R2807 vss.n3273 vss.n3272 0.00577551
R2808 vss.n2934 vss.n2932 0.00570833
R2809 vss.n2950 vss.n2949 0.00570833
R2810 vss.n1194 vss.n1193 0.00570833
R2811 vss.n1128 vss.n1123 0.00570833
R2812 vss.n574 vss.n572 0.00570833
R2813 vss.n2118 vss.n2117 0.00570833
R2814 vss.n2014 vss.n2012 0.00570833
R2815 vss.n2009 vss.n1996 0.00570833
R2816 vss.n3194 vss.n116 0.00554032
R2817 vss.n2725 vss.n2724 0.00531433
R2818 vss.n1943 vss.n1942 0.00523154
R2819 vss.n1943 vss.n635 0.00523154
R2820 vss.n2513 vss.n2512 0.00523154
R2821 vss.n2509 vss.n2508 0.00523154
R2822 vss.n2508 vss.n2507 0.00523154
R2823 vss.n2506 vss.n2505 0.00523154
R2824 vss.n2505 vss.n2504 0.00523154
R2825 vss.n2503 vss.n2502 0.00523154
R2826 vss.n2502 vss.n2285 0.00523154
R2827 vss.n2319 vss.n2318 0.00523154
R2828 vss.n2320 vss.n2319 0.00523154
R2829 vss.n2322 vss.n2321 0.00523154
R2830 vss.n2323 vss.n2322 0.00523154
R2831 vss.n2325 vss.n2324 0.00523154
R2832 vss.n2326 vss.n2325 0.00523154
R2833 vss.n2403 vss.n2327 0.00523154
R2834 vss.n2403 vss.n2402 0.00523154
R2835 vss.n2401 vss.n2400 0.00523154
R2836 vss.n2400 vss.n2383 0.00523154
R2837 vss.n2382 vss.n2381 0.00523154
R2838 vss.n2151 vss.n2150 0.00523154
R2839 vss.n2152 vss.n2151 0.00523154
R2840 vss.n2154 vss.n2153 0.00523154
R2841 vss.n2155 vss.n2154 0.00523154
R2842 vss.n2157 vss.n2156 0.00523154
R2843 vss.n2158 vss.n2157 0.00523154
R2844 vss.n2273 vss.n2159 0.00523154
R2845 vss.n2274 vss.n2273 0.00523154
R2846 vss.n2276 vss.n2275 0.00523154
R2847 vss.n2277 vss.n2276 0.00523154
R2848 vss.n2279 vss.n2278 0.00523154
R2849 vss.n2280 vss.n2279 0.00523154
R2850 vss.n2282 vss.n2281 0.00523154
R2851 vss.n2283 vss.n2282 0.00523154
R2852 vss.n2516 vss.n2284 0.00523154
R2853 vss.n2516 vss.n2515 0.00523154
R2854 vss.n2813 vss.n2802 0.00523154
R2855 vss.n2813 vss.n2812 0.00523154
R2856 vss.n2811 vss.n2810 0.00523154
R2857 vss.n2810 vss.n2809 0.00523154
R2858 vss.n2808 vss.n2807 0.00523154
R2859 vss.n2807 vss.n2806 0.00523154
R2860 vss.n2805 vss.n2804 0.00523154
R2861 vss.n2804 vss.n2803 0.00523154
R2862 vss.n2755 vss.n2725 0.00523154
R2863 vss.n2756 vss.n2755 0.00523154
R2864 vss.n2769 vss.n2757 0.00523154
R2865 vss.n2770 vss.n2769 0.00523154
R2866 vss.n2783 vss.n2771 0.00523154
R2867 vss.n2784 vss.n2783 0.00523154
R2868 vss.n2800 vss.n2785 0.00523154
R2869 vss.n2801 vss.n2800 0.00523154
R2870 vss.n1619 vss.n1618 0.00521572
R2871 vss.n1617 vss.n1616 0.00521572
R2872 vss.n1616 vss.n1615 0.00521572
R2873 vss.n1614 vss.n1613 0.00521572
R2874 vss.n1613 vss.n1612 0.00521572
R2875 vss.n1611 vss.n1610 0.00521572
R2876 vss.n1610 vss.n720 0.00521572
R2877 vss.n1603 vss.n1551 0.00521572
R2878 vss.n1603 vss.n1602 0.00521572
R2879 vss.n1601 vss.n1600 0.00521572
R2880 vss.n1600 vss.n1588 0.00521572
R2881 vss.n1587 vss.n1586 0.00521572
R2882 vss.n1586 vss.n1568 0.00521572
R2883 vss.n1567 vss.n1566 0.00521572
R2884 vss.n1113 vss.n1112 0.00521572
R2885 vss.n1112 vss.n1111 0.00521572
R2886 vss.n1110 vss.n1109 0.00521572
R2887 vss.n1109 vss.n1108 0.00521572
R2888 vss.n1107 vss.n1106 0.00521572
R2889 vss.n1106 vss.n1105 0.00521572
R2890 vss.n1104 vss.n1103 0.00521572
R2891 vss.n1103 vss.n788 0.00521572
R2892 vss.n1327 vss.n1326 0.00521572
R2893 vss.n1328 vss.n1327 0.00521572
R2894 vss.n1330 vss.n1329 0.00521572
R2895 vss.n1331 vss.n1330 0.00521572
R2896 vss.n1333 vss.n1332 0.00521572
R2897 vss.n1334 vss.n1333 0.00521572
R2898 vss.n1452 vss.n1335 0.00521572
R2899 vss.n1453 vss.n1452 0.00521572
R2900 vss.n1455 vss.n1454 0.00521572
R2901 vss.n1456 vss.n1455 0.00521572
R2902 vss.n1458 vss.n1457 0.00521572
R2903 vss.n1459 vss.n1458 0.00521572
R2904 vss.n1461 vss.n1460 0.00521572
R2905 vss.n1462 vss.n1461 0.00521572
R2906 vss.n1464 vss.n1463 0.00521572
R2907 vss.n1464 vss.n719 0.00521572
R2908 vss.n1937 vss.n688 0.00521572
R2909 vss.n1938 vss.n1937 0.00521572
R2910 vss.n1940 vss.n1939 0.00521572
R2911 vss.n1941 vss.n1940 0.00521572
R2912 vss.n2149 vss 0.00496556
R2913 vss.n786 vss.n781 0.00493396
R2914 vss.n787 vss.n786 0.00493396
R2915 vss.n1181 vss.n1115 0.00490287
R2916 vss.n779 vss.n778 0.00489326
R2917 vss.n2067 vss.n2066 0.00489326
R2918 vss.n643 vss.n642 0.00489326
R2919 vss.n3259 vss.n3258 0.00489326
R2920 vss.n362 vss.n361 0.00489252
R2921 vss.n550 vss.n549 0.00481193
R2922 vss.n549 vss.n548 0.00481193
R2923 vss.n547 vss.n546 0.00481193
R2924 vss.n546 vss.n529 0.00481193
R2925 vss.n528 vss.n527 0.00481193
R2926 vss.n527 vss.n515 0.00481193
R2927 vss.n514 vss.n513 0.00481193
R2928 vss.n513 vss.n487 0.00481193
R2929 vss.n2635 vss.n2634 0.00481193
R2930 vss.n2637 vss.n2636 0.00481193
R2931 vss.n2638 vss.n2637 0.00481193
R2932 vss.n2640 vss.n2639 0.00481193
R2933 vss.n2641 vss.n2640 0.00481193
R2934 vss.n2643 vss.n2642 0.00481193
R2935 vss.n2644 vss.n2643 0.00481193
R2936 vss.n2647 vss.n2645 0.00481193
R2937 vss.n2647 vss.n2646 0.00481193
R2938 vss.n2681 vss.n363 0.00481193
R2939 vss.n2682 vss.n2681 0.00481193
R2940 vss.n2718 vss.n2683 0.00481193
R2941 vss.n2719 vss.n2718 0.00481193
R2942 vss.n486 vss.n485 0.00481193
R2943 vss.n485 vss.n484 0.00481193
R2944 vss.n483 vss.n482 0.00481193
R2945 vss.n482 vss.n481 0.00481193
R2946 vss.n480 vss.n479 0.00481193
R2947 vss.n479 vss.n478 0.00481193
R2948 vss.n477 vss.n476 0.00481193
R2949 vss.n476 vss.n475 0.00481193
R2950 vss.n357 vss.n356 0.00481193
R2951 vss.n356 vss.n355 0.00481193
R2952 vss.n354 vss.n353 0.00481193
R2953 vss.n353 vss.n352 0.00481193
R2954 vss.n351 vss.n350 0.00481193
R2955 vss.n350 vss.n349 0.00481193
R2956 vss.n348 vss.n347 0.00481193
R2957 vss.n347 vss.n207 0.00481193
R2958 vss.n340 vss.n329 0.00481193
R2959 vss.n340 vss.n339 0.00481193
R2960 vss.n338 vss.n337 0.00481193
R2961 vss.n337 vss.n336 0.00481193
R2962 vss.n335 vss.n334 0.00481193
R2963 vss.n334 vss.n333 0.00481193
R2964 vss.n332 vss.n331 0.00481193
R2965 vss.n331 vss.n330 0.00481193
R2966 vss.n1227 vss 0.00463641
R2967 vss.n2511 vss.n2510 0.00460067
R2968 vss.n77 vss.n73 0.00457609
R2969 vss.n1252 vss.n733 0.0045634
R2970 vss.n1253 vss.n1252 0.0045634
R2971 vss.n1272 vss.n1254 0.0045634
R2972 vss.n1273 vss.n1272 0.0045634
R2973 vss.n1286 vss.n1274 0.0045634
R2974 vss.n1287 vss.n1286 0.0045634
R2975 vss.n1311 vss.n1288 0.0045634
R2976 vss.n1312 vss.n1311 0.0045634
R2977 vss.n925 vss.n924 0.0045634
R2978 vss.n926 vss.n925 0.0045634
R2979 vss.n928 vss.n927 0.0045634
R2980 vss.n929 vss.n928 0.0045634
R2981 vss.n931 vss.n930 0.0045634
R2982 vss.n932 vss.n931 0.0045634
R2983 vss.n983 vss.n933 0.0045634
R2984 vss.n983 vss.n982 0.0045634
R2985 vss.n981 vss.n980 0.0045634
R2986 vss.n980 vss.n963 0.0045634
R2987 vss.n962 vss.n961 0.0045634
R2988 vss.n1697 vss.n1696 0.0045634
R2989 vss.n1698 vss.n1697 0.0045634
R2990 vss.n1700 vss.n1699 0.0045634
R2991 vss.n1701 vss.n1700 0.0045634
R2992 vss.n1703 vss.n1702 0.0045634
R2993 vss.n1704 vss.n1703 0.0045634
R2994 vss.n1720 vss.n1705 0.0045634
R2995 vss.n1721 vss.n1720 0.0045634
R2996 vss.n1734 vss.n1722 0.0045634
R2997 vss.n1735 vss.n1734 0.0045634
R2998 vss.n1748 vss.n1736 0.0045634
R2999 vss.n1749 vss.n1748 0.0045634
R3000 vss.n1780 vss.n1750 0.0045634
R3001 vss.n1796 vss.n1795 0.0045634
R3002 vss.n1795 vss.n1794 0.0045634
R3003 vss.n1793 vss.n1792 0.0045634
R3004 vss.n1792 vss.n1791 0.0045634
R3005 vss.n1790 vss.n1789 0.0045634
R3006 vss.n1789 vss.n1788 0.0045634
R3007 vss.n1984 vss.n653 0.0045634
R3008 vss.n1985 vss.n1984 0.0045634
R3009 vss.n1863 vss.n1812 0.0045634
R3010 vss.n1811 vss.n1810 0.0045634
R3011 vss.n1810 vss.n1797 0.0045634
R3012 vss.n585 vss.n584 0.00451955
R3013 vss.n1992 vss.n1991 0.00451955
R3014 vss.n2935 vss.n2934 0.00440625
R3015 vss.n1189 vss.n1145 0.00440625
R3016 vss.n1196 vss.n1194 0.00440625
R3017 vss.n571 vss.n553 0.00440625
R3018 vss.n576 vss.n574 0.00440625
R3019 vss.n2012 vss.n2010 0.00440625
R3020 vss.n100 vss.n89 0.00440625
R3021 vss.n43 vss.n24 0.00440625
R3022 vss.n2381 vss.n358 0.00428523
R3023 vss.n1137 vss.n1132 0.0042807
R3024 vss.n3271 vss.n3266 0.00415285
R3025 vss.n1787 vss.n1786 0.00410644
R3026 vss.n1784 vss.n1783 0.00410644
R3027 vss.n1870 vss.n1869 0.00410644
R3028 vss.n961 vss.n949 0.00402161
R3029 vss.n400 vss.n399 0.00401501
R3030 vss.n3005 vss.n3004 0.00397409
R3031 vss.n3001 vss.n3000 0.00397409
R3032 vss.n2997 vss.n2996 0.00397409
R3033 vss.n2993 vss.n2992 0.00397409
R3034 vss.n2989 vss.n2988 0.00397409
R3035 vss.n2981 vss.n2980 0.00397409
R3036 vss.n3134 vss.n3133 0.00397409
R3037 vss.n2969 vss.n2968 0.00397409
R3038 vss.n2973 vss.n2972 0.00397409
R3039 vss.n2977 vss.n2976 0.00397409
R3040 vss.n2985 vss.n2984 0.00397409
R3041 vss.n3285 vss.n3284 0.00397409
R3042 vss.n3306 vss.n3305 0.00397409
R3043 vss.n3320 vss.n3319 0.00397409
R3044 vss.n3291 vss.n3290 0.00397409
R3045 vss.n2353 vss.n2352 0.00392584
R3046 vss.n360 vss.n359 0.00392584
R3047 vss.n2880 vss.n2879 0.0038874
R3048 vss.n2883 vss 0.00385714
R3049 vss.n3323 vss.n3322 0.00385391
R3050 vss.n3028 vss.n3023 0.00372581
R3051 vss.n3273 vss.n3271 0.0036658
R3052 vss.n2510 vss.n2509 0.00365436
R3053 vss.n2507 vss.n2506 0.00365436
R3054 vss.n2504 vss.n2503 0.00365436
R3055 vss.n2321 vss.n2320 0.00365436
R3056 vss.n2324 vss.n2323 0.00365436
R3057 vss.n2327 vss.n2326 0.00365436
R3058 vss.n2383 vss.n2382 0.00365436
R3059 vss.n2153 vss.n2152 0.00365436
R3060 vss.n2156 vss.n2155 0.00365436
R3061 vss.n2159 vss.n2158 0.00365436
R3062 vss.n2278 vss.n2277 0.00365436
R3063 vss.n2281 vss.n2280 0.00365436
R3064 vss.n2284 vss.n2283 0.00365436
R3065 vss.n2812 vss.n2811 0.00365436
R3066 vss.n2809 vss.n2808 0.00365436
R3067 vss.n2806 vss.n2805 0.00365436
R3068 vss.n2757 vss.n2756 0.00365436
R3069 vss.n2771 vss.n2770 0.00365436
R3070 vss.n2785 vss.n2784 0.00365436
R3071 vss.n1620 vss.n1619 0.00364381
R3072 vss.n1618 vss.n1617 0.00364381
R3073 vss.n1615 vss.n1614 0.00364381
R3074 vss.n1612 vss.n1611 0.00364381
R3075 vss.n1602 vss.n1601 0.00364381
R3076 vss.n1588 vss.n1587 0.00364381
R3077 vss.n1568 vss.n1567 0.00364381
R3078 vss.n1111 vss.n1110 0.00364381
R3079 vss.n1108 vss.n1107 0.00364381
R3080 vss.n1105 vss.n1104 0.00364381
R3081 vss.n1329 vss.n1328 0.00364381
R3082 vss.n1332 vss.n1331 0.00364381
R3083 vss.n1335 vss.n1334 0.00364381
R3084 vss.n1457 vss.n1456 0.00364381
R3085 vss.n1460 vss.n1459 0.00364381
R3086 vss.n1463 vss.n1462 0.00364381
R3087 vss.n1866 vss.n688 0.00364381
R3088 vss.n1939 vss.n1938 0.00364381
R3089 vss.n625 vss.n624 0.00362372
R3090 vss.n1134 vss.n1132 0.00360776
R3091 vss.n3223 vss.n3222 0.00345276
R3092 vss.n3219 vss.n3215 0.00345276
R3093 vss.n1872 vss.n1868 0.00343981
R3094 vss.n1052 vss.n1051 0.0034393
R3095 vss.n1323 vss.n1322 0.0034393
R3096 vss.n3205 vss.n3202 0.00340698
R3097 vss.n548 vss.n547 0.00337462
R3098 vss.n529 vss.n528 0.00337462
R3099 vss.n515 vss.n514 0.00337462
R3100 vss.n2639 vss.n2638 0.00337462
R3101 vss.n2642 vss.n2641 0.00337462
R3102 vss.n2645 vss.n2644 0.00337462
R3103 vss.n2683 vss.n2682 0.00337462
R3104 vss.n2720 vss.n2719 0.00337462
R3105 vss.n484 vss.n483 0.00337462
R3106 vss.n481 vss.n480 0.00337462
R3107 vss.n478 vss.n477 0.00337462
R3108 vss.n355 vss.n354 0.00337462
R3109 vss.n352 vss.n351 0.00337462
R3110 vss.n349 vss.n348 0.00337462
R3111 vss.n339 vss.n338 0.00337462
R3112 vss.n336 vss.n335 0.00337462
R3113 vss.n333 vss.n332 0.00337462
R3114 vss.n397 vss.n396 0.00334838
R3115 vss.n2926 vss.n2925 0.00327559
R3116 vss.n2924 vss.n2886 0.00327559
R3117 vss.n3167 vss.n3166 0.00327559
R3118 vss.n3166 vss.n3165 0.00327559
R3119 vss.n3164 vss.n3163 0.00327559
R3120 vss.n3163 vss.n3162 0.00327559
R3121 vss.n3161 vss.n3160 0.00327559
R3122 vss.n3160 vss.n3159 0.00327559
R3123 vss.n3158 vss.n3157 0.00327559
R3124 vss.n3157 vss.n3156 0.00327559
R3125 vss.n3155 vss.n3154 0.00327559
R3126 vss.n3154 vss.n3153 0.00327559
R3127 vss.n3152 vss.n3151 0.00327559
R3128 vss.n3151 vss.n3150 0.00327559
R3129 vss.n3149 vss.n3148 0.00327559
R3130 vss.n3148 vss.n3147 0.00327559
R3131 vss.n3146 vss.n3145 0.00327559
R3132 vss.n3145 vss.n3144 0.00327559
R3133 vss.n3143 vss.n3142 0.00327559
R3134 vss.n3142 vss.n3141 0.00327559
R3135 vss.n3140 vss.n3139 0.00327559
R3136 vss.n3139 vss.n3138 0.00327559
R3137 vss.n3137 vss.n3136 0.00327559
R3138 vss.n3136 vss.n3135 0.00327559
R3139 vss.n3176 vss.n125 0.00324725
R3140 vss.n141 vss.n140 0.00322077
R3141 vss.n1254 vss.n1253 0.00320893
R3142 vss.n1274 vss.n1273 0.00320893
R3143 vss.n1288 vss.n1287 0.00320893
R3144 vss.n927 vss.n926 0.00320893
R3145 vss.n930 vss.n929 0.00320893
R3146 vss.n933 vss.n932 0.00320893
R3147 vss.n963 vss.n962 0.00320893
R3148 vss.n1696 vss.n1695 0.00320893
R3149 vss.n1699 vss.n1698 0.00320893
R3150 vss.n1702 vss.n1701 0.00320893
R3151 vss.n1722 vss.n1721 0.00320893
R3152 vss.n1736 vss.n1735 0.00320893
R3153 vss.n1750 vss.n1749 0.00320893
R3154 vss.n1794 vss.n1793 0.00320893
R3155 vss.n1791 vss.n1790 0.00320893
R3156 vss.n1788 vss.n653 0.00320893
R3157 vss.n1864 vss.n1863 0.00320893
R3158 vss.n1812 vss.n1811 0.00320893
R3159 vss.n1695 vss.n1694 0.00307349
R3160 vss.n1781 vss.n1780 0.00307349
R3161 vss.n19 vss.n0 0.00306576
R3162 vss.n47 vss.n46 0.00306576
R3163 vss vss.n2888 0.00302525
R3164 vss.n2926 vss.n2923 0.00299803
R3165 vss.n3303 vss.n3300 0.00293507
R3166 vss.n3037 vss.n3033 0.00291935
R3167 vss.n3010 vss 0.00291935
R3168 vss.n3198 vss.n107 0.00286895
R3169 vss.n3243 vss.n3242 0.00286895
R3170 vss.n83 vss.n50 0.00283251
R3171 vss.n2355 vss.n2354 0.00279583
R3172 vss.n1314 vss.n1313 0.00277266
R3173 vss.n1050 vss.n1049 0.00277266
R3174 vss.n1230 vss.n1229 0.00270045
R3175 vss.n138 vss.n137 0.00266667
R3176 vss.n401 vss 0.00265596
R3177 vss.n214 vss.n213 0.00257353
R3178 vss.n216 vss.n215 0.00257353
R3179 vss.n225 vss.n224 0.00257353
R3180 vss.n227 vss.n226 0.00257353
R3181 vss.n236 vss.n235 0.00257353
R3182 vss.n238 vss.n237 0.00257353
R3183 vss.n345 vss.n344 0.00257353
R3184 vss.n343 vss.n342 0.00257353
R3185 vss.n328 vss.n327 0.00257353
R3186 vss.n326 vss.n325 0.00257353
R3187 vss.n323 vss.n322 0.00257353
R3188 vss.n321 vss.n320 0.00257353
R3189 vss.n318 vss.n317 0.00257353
R3190 vss.n316 vss.n315 0.00257353
R3191 vss.n1927 vss.n1926 0.00257353
R3192 vss.n1929 vss.n1928 0.00257353
R3193 vss.n1935 vss.n1934 0.00257353
R3194 vss.n1933 vss.n1932 0.00257353
R3195 vss.n1708 vss.n1707 0.00257353
R3196 vss.n1724 vss.n1723 0.00257353
R3197 vss.n1732 vss.n1731 0.00257353
R3198 vss.n1738 vss.n1737 0.00257353
R3199 vss.n1746 vss.n1745 0.00257353
R3200 vss.n1752 vss.n1751 0.00257353
R3201 vss.n1778 vss.n1777 0.00257353
R3202 vss.n1814 vss.n1813 0.00257353
R3203 vss.n1846 vss.n1845 0.00257353
R3204 vss.n1799 vss.n1798 0.00257353
R3205 vss.n1342 vss.n1341 0.00257353
R3206 vss.n1344 vss.n1343 0.00257353
R3207 vss.n1353 vss.n1352 0.00257353
R3208 vss.n1355 vss.n1354 0.00257353
R3209 vss.n1364 vss.n1363 0.00257353
R3210 vss.n1366 vss.n1365 0.00257353
R3211 vss.n1450 vss.n1449 0.00257353
R3212 vss.n1448 vss.n1447 0.00257353
R3213 vss.n1445 vss.n1444 0.00257353
R3214 vss.n1443 vss.n1442 0.00257353
R3215 vss.n1440 vss.n1439 0.00257353
R3216 vss.n1438 vss.n1437 0.00257353
R3217 vss.n1435 vss.n1434 0.00257353
R3218 vss.n1433 vss.n721 0.00257353
R3219 vss.n1467 vss.n1466 0.00257353
R3220 vss.n1469 vss.n1468 0.00257353
R3221 vss.n1475 vss.n1474 0.00257353
R3222 vss.n1477 vss.n1476 0.00257353
R3223 vss.n1486 vss.n1485 0.00257353
R3224 vss.n1488 vss.n1487 0.00257353
R3225 vss.n1497 vss.n1496 0.00257353
R3226 vss.n1499 vss.n1498 0.00257353
R3227 vss.n1608 vss.n1607 0.00257353
R3228 vss.n1606 vss.n1605 0.00257353
R3229 vss.n1550 vss.n1549 0.00257353
R3230 vss.n1590 vss.n1589 0.00257353
R3231 vss.n1598 vss.n1597 0.00257353
R3232 vss.n1570 vss.n1569 0.00257353
R3233 vss.n1584 vss.n1583 0.00257353
R3234 vss.n1553 vss.n1552 0.00257353
R3235 vss.n736 vss.n735 0.00257353
R3236 vss.n1256 vss.n1255 0.00257353
R3237 vss.n1270 vss.n1269 0.00257353
R3238 vss.n1276 vss.n1275 0.00257353
R3239 vss.n1284 vss.n1283 0.00257353
R3240 vss.n1290 vss.n1289 0.00257353
R3241 vss.n795 vss.n794 0.00257353
R3242 vss.n797 vss.n796 0.00257353
R3243 vss.n806 vss.n805 0.00257353
R3244 vss.n808 vss.n807 0.00257353
R3245 vss.n817 vss.n816 0.00257353
R3246 vss.n819 vss.n818 0.00257353
R3247 vss.n1101 vss.n1100 0.00257353
R3248 vss.n1099 vss.n1098 0.00257353
R3249 vss.n1019 vss.n1018 0.00257353
R3250 vss.n1017 vss.n1016 0.00257353
R3251 vss.n998 vss.n997 0.00257353
R3252 vss.n996 vss.n995 0.00257353
R3253 vss.n993 vss.n992 0.00257353
R3254 vss.n991 vss.n990 0.00257353
R3255 vss.n988 vss.n987 0.00257353
R3256 vss.n986 vss.n985 0.00257353
R3257 vss.n964 vss.n923 0.00257353
R3258 vss.n966 vss.n965 0.00257353
R3259 vss.n978 vss.n977 0.00257353
R3260 vss.n951 vss.n950 0.00257353
R3261 vss.n959 vss.n958 0.00257353
R3262 vss.n936 vss.n935 0.00257353
R3263 vss.n944 vss.n943 0.00257353
R3264 vss.n693 vss.n692 0.00257353
R3265 vss.n1627 vss.n1626 0.00257353
R3266 vss.n1629 vss.n1628 0.00257353
R3267 vss.n1691 vss.n1690 0.00257353
R3268 vss.n1689 vss.n1688 0.00257353
R3269 vss.n1686 vss.n1685 0.00257353
R3270 vss.n1684 vss.n1683 0.00257353
R3271 vss.n1681 vss.n1680 0.00257353
R3272 vss.n1679 vss.n1678 0.00257353
R3273 vss.n655 vss.n654 0.00257353
R3274 vss.n657 vss.n656 0.00257353
R3275 vss.n660 vss.n659 0.00257353
R3276 vss.n662 vss.n661 0.00257353
R3277 vss.n665 vss.n664 0.00257353
R3278 vss.n667 vss.n666 0.00257353
R3279 vss.n2166 vss.n2165 0.00257353
R3280 vss.n2168 vss.n2167 0.00257353
R3281 vss.n2177 vss.n2176 0.00257353
R3282 vss.n2179 vss.n2178 0.00257353
R3283 vss.n2188 vss.n2187 0.00257353
R3284 vss.n2190 vss.n2189 0.00257353
R3285 vss.n2240 vss.n2239 0.00257353
R3286 vss.n2238 vss.n2237 0.00257353
R3287 vss.n447 vss.n446 0.00257353
R3288 vss.n449 vss.n448 0.00257353
R3289 vss.n452 vss.n451 0.00257353
R3290 vss.n454 vss.n453 0.00257353
R3291 vss.n457 vss.n456 0.00257353
R3292 vss.n459 vss.n458 0.00257353
R3293 vss.n464 vss.n463 0.00257353
R3294 vss.n531 vss.n530 0.00257353
R3295 vss.n544 vss.n543 0.00257353
R3296 vss.n517 vss.n516 0.00257353
R3297 vss.n525 vss.n524 0.00257353
R3298 vss.n489 vss.n488 0.00257353
R3299 vss.n408 vss.n407 0.00257353
R3300 vss.n410 vss.n409 0.00257353
R3301 vss.n419 vss.n418 0.00257353
R3302 vss.n421 vss.n420 0.00257353
R3303 vss.n430 vss.n429 0.00257353
R3304 vss.n432 vss.n431 0.00257353
R3305 vss.n2539 vss.n2538 0.00257353
R3306 vss.n2541 vss.n2540 0.00257353
R3307 vss.n2632 vss.n2631 0.00257353
R3308 vss.n2630 vss.n2629 0.00257353
R3309 vss.n2627 vss.n2626 0.00257353
R3310 vss.n2625 vss.n2624 0.00257353
R3311 vss.n2622 vss.n2621 0.00257353
R3312 vss.n2620 vss.n2619 0.00257353
R3313 vss.n2617 vss.n2616 0.00257353
R3314 vss.n2615 vss.n364 0.00257353
R3315 vss.n2650 vss.n2649 0.00257353
R3316 vss.n2652 vss.n2651 0.00257353
R3317 vss.n2679 vss.n2678 0.00257353
R3318 vss.n2685 vss.n2684 0.00257353
R3319 vss.n2716 vss.n2715 0.00257353
R3320 vss.n2714 vss.n2713 0.00257353
R3321 vss.n2292 vss.n2291 0.00257353
R3322 vss.n2294 vss.n2293 0.00257353
R3323 vss.n2303 vss.n2302 0.00257353
R3324 vss.n2305 vss.n2304 0.00257353
R3325 vss.n2314 vss.n2313 0.00257353
R3326 vss.n2316 vss.n2315 0.00257353
R3327 vss.n2469 vss.n2468 0.00257353
R3328 vss.n2467 vss.n2466 0.00257353
R3329 vss.n2448 vss.n2447 0.00257353
R3330 vss.n2446 vss.n2445 0.00257353
R3331 vss.n2437 vss.n2436 0.00257353
R3332 vss.n2435 vss.n2434 0.00257353
R3333 vss.n2419 vss.n2418 0.00257353
R3334 vss.n2417 vss.n2416 0.00257353
R3335 vss.n2384 vss.n2317 0.00257353
R3336 vss.n2386 vss.n2385 0.00257353
R3337 vss.n2388 vss.n2387 0.00257353
R3338 vss.n2329 vss.n2328 0.00257353
R3339 vss.n2331 vss.n2330 0.00257353
R3340 vss.n2727 vss.n2726 0.00257353
R3341 vss.n2729 vss.n2728 0.00257353
R3342 vss.n2759 vss.n2758 0.00257353
R3343 vss.n2761 vss.n2760 0.00257353
R3344 vss.n2773 vss.n2772 0.00257353
R3345 vss.n2775 vss.n2774 0.00257353
R3346 vss.n2787 vss.n2786 0.00257353
R3347 vss.n206 vss.n205 0.00257353
R3348 vss.n204 vss.n203 0.00257353
R3349 vss.n201 vss.n200 0.00257353
R3350 vss.n199 vss.n198 0.00257353
R3351 vss.n196 vss.n195 0.00257353
R3352 vss.n194 vss.n193 0.00257353
R3353 vss.n1871 vss.n1870 0.00255288
R3354 vss.n1785 vss.n1784 0.00255288
R3355 vss.n1786 vss.n1785 0.00255288
R3356 vss.n399 vss.n398 0.00250717
R3357 vss.n2923 vss.n2922 0.0025061
R3358 vss.n947 vss.n946 0.00248592
R3359 vss.n1624 vss.n718 0.00248592
R3360 vss.n1624 vss.n1623 0.00248592
R3361 vss.n1693 vss.n691 0.00248592
R3362 vss.n946 vss.n934 0.00248592
R3363 vss.n2354 vss.n2353 0.00246292
R3364 vss.n361 vss.n360 0.00246292
R3365 vss.n3239 vss.n3238 0.00245312
R3366 vss.n87 vss.n86 0.00245312
R3367 vss.n89 vss.n88 0.00245312
R3368 vss.n91 vss.n90 0.00245312
R3369 vss.n16 vss.n15 0.00245312
R3370 vss.n22 vss.n21 0.00245312
R3371 vss.n24 vss.n23 0.00245312
R3372 vss.n42 vss.n41 0.00245312
R3373 vss.n3175 vss.n3174 0.00244755
R3374 vss.n2879 vss.n2878 0.00244338
R3375 vss.n1566 vss.n690 0.00238629
R3376 vss.n286 vss.n285 0.00233824
R3377 vss.n282 vss.n281 0.00233824
R3378 vss.n274 vss.n273 0.00233824
R3379 vss.n247 vss.n246 0.00233824
R3380 vss.n254 vss.n253 0.00233824
R3381 vss.n261 vss.n260 0.00233824
R3382 vss.n222 vss.n220 0.00233824
R3383 vss.n233 vss.n231 0.00233824
R3384 vss.n269 vss.n242 0.00233824
R3385 vss.n312 vss.n311 0.00233824
R3386 vss.n306 vss.n305 0.00233824
R3387 vss.n300 vss.n299 0.00233824
R3388 vss.n2855 vss.n2851 0.00233824
R3389 vss.n2867 vss.n2863 0.00233824
R3390 vss.n2873 vss.n2872 0.00233824
R3391 vss.n167 vss.n164 0.00233824
R3392 vss.n159 vss.n158 0.00233824
R3393 vss.n1819 vss.n1818 0.00233824
R3394 vss.n1860 vss.n1859 0.00233824
R3395 vss.n1807 vss.n1806 0.00233824
R3396 vss.n1893 vss.n1892 0.00233824
R3397 vss.n1889 vss.n1888 0.00233824
R3398 vss.n1882 vss.n1881 0.00233824
R3399 vss.n1920 vss.n1919 0.00233824
R3400 vss.n1914 vss.n1913 0.00233824
R3401 vss.n1908 vss.n1907 0.00233824
R3402 vss.n1715 vss.n1713 0.00233824
R3403 vss.n1761 vss.n1760 0.00233824
R3404 vss.n1768 vss.n1767 0.00233824
R3405 vss.n1730 vss.n1727 0.00233824
R3406 vss.n1744 vss.n1741 0.00233824
R3407 vss.n1776 vss.n1755 0.00233824
R3408 vss.n1375 vss.n1374 0.00233824
R3409 vss.n1382 vss.n1381 0.00233824
R3410 vss.n1389 vss.n1388 0.00233824
R3411 vss.n1350 vss.n1348 0.00233824
R3412 vss.n1361 vss.n1359 0.00233824
R3413 vss.n1397 vss.n1370 0.00233824
R3414 vss.n1403 vss.n1402 0.00233824
R3415 vss.n1429 vss.n1428 0.00233824
R3416 vss.n730 vss.n729 0.00233824
R3417 vss.n1413 vss.n1412 0.00233824
R3418 vss.n1419 vss.n1418 0.00233824
R3419 vss.n1432 vss.n1431 0.00233824
R3420 vss.n1508 vss.n1507 0.00233824
R3421 vss.n1515 vss.n1514 0.00233824
R3422 vss.n1522 vss.n1521 0.00233824
R3423 vss.n1483 vss.n1481 0.00233824
R3424 vss.n1494 vss.n1492 0.00233824
R3425 vss.n1530 vss.n1503 0.00233824
R3426 vss.n1537 vss.n1536 0.00233824
R3427 vss.n1578 vss.n1577 0.00233824
R3428 vss.n1561 vss.n1560 0.00233824
R3429 vss.n1548 vss.n1547 0.00233824
R3430 vss.n1596 vss.n1595 0.00233824
R3431 vss.n1582 vss.n1581 0.00233824
R3432 vss.n1247 vss.n1245 0.00233824
R3433 vss.n1265 vss.n1264 0.00233824
R3434 vss.n1300 vss.n1299 0.00233824
R3435 vss.n1268 vss.n1259 0.00233824
R3436 vss.n1282 vss.n1279 0.00233824
R3437 vss.n1308 vss.n1293 0.00233824
R3438 vss.n1165 vss.n1164 0.00233824
R3439 vss.n1161 vss.n1160 0.00233824
R3440 vss.n1157 vss.n1153 0.00233824
R3441 vss.n746 vss.n745 0.00233824
R3442 vss.n752 vss.n751 0.00233824
R3443 vss.n1234 vss.n757 0.00233824
R3444 vss.n828 vss.n827 0.00233824
R3445 vss.n835 vss.n834 0.00233824
R3446 vss.n842 vss.n841 0.00233824
R3447 vss.n803 vss.n801 0.00233824
R3448 vss.n814 vss.n812 0.00233824
R3449 vss.n851 vss.n823 0.00233824
R3450 vss.n1081 vss.n1080 0.00233824
R3451 vss.n860 vss.n859 0.00233824
R3452 vss.n1058 vss.n1057 0.00233824
R3453 vss.n1096 vss.n1095 0.00233824
R3454 vss.n1090 vss.n1089 0.00233824
R3455 vss.n1073 vss.n1072 0.00233824
R3456 vss.n1069 vss.n1068 0.00233824
R3457 vss.n1065 vss.n1029 0.00233824
R3458 vss.n878 vss.n876 0.00233824
R3459 vss.n888 vss.n886 0.00233824
R3460 vss.n1021 vss.n870 0.00233824
R3461 vss.n1004 vss.n1003 0.00233824
R3462 vss.n908 vss.n907 0.00233824
R3463 vss.n920 vss.n919 0.00233824
R3464 vss.n1014 vss.n1013 0.00233824
R3465 vss.n898 vss.n897 0.00233824
R3466 vss.n911 vss.n910 0.00233824
R3467 vss.n973 vss.n971 0.00233824
R3468 vss.n702 vss.n701 0.00233824
R3469 vss.n709 vss.n708 0.00233824
R3470 vss.n957 vss.n954 0.00233824
R3471 vss.n942 vss.n939 0.00233824
R3472 vss.n717 vss.n696 0.00233824
R3473 vss.n1648 vss.n1647 0.00233824
R3474 vss.n1644 vss.n1643 0.00233824
R3475 vss.n1637 vss.n1636 0.00233824
R3476 vss.n1660 vss.n1659 0.00233824
R3477 vss.n1666 vss.n1665 0.00233824
R3478 vss.n1672 vss.n1671 0.00233824
R3479 vss.n1960 vss.n1956 0.00233824
R3480 vss.n1972 vss.n1968 0.00233824
R3481 vss.n1979 vss.n1978 0.00233824
R3482 vss.n682 vss.n679 0.00233824
R3483 vss.n674 vss.n673 0.00233824
R3484 vss.n2106 vss.n2105 0.00233824
R3485 vss.n2041 vss.n2040 0.00233824
R3486 vss.n2048 vss.n2047 0.00233824
R3487 vss.n2082 vss.n2080 0.00233824
R3488 vss.n2095 vss.n2092 0.00233824
R3489 vss.n2057 vss.n2035 0.00233824
R3490 vss.n2174 vss.n2172 0.00233824
R3491 vss.n2185 vss.n2183 0.00233824
R3492 vss.n2271 vss.n2244 0.00233824
R3493 vss.n2220 vss.n2219 0.00233824
R3494 vss.n2199 vss.n2198 0.00233824
R3495 vss.n2520 vss.n2519 0.00233824
R3496 vss.n2235 vss.n2234 0.00233824
R3497 vss.n2229 vss.n2228 0.00233824
R3498 vss.n2247 vss.n2246 0.00233824
R3499 vss.n2255 vss.n2254 0.00233824
R3500 vss.n2262 vss.n2261 0.00233824
R3501 vss.n470 vss.n468 0.00233824
R3502 vss.n539 vss.n538 0.00233824
R3503 vss.n502 vss.n501 0.00233824
R3504 vss.n542 vss.n534 0.00233824
R3505 vss.n523 vss.n520 0.00233824
R3506 vss.n510 vss.n492 0.00233824
R3507 vss.n2212 vss.n2211 0.00233824
R3508 vss.n2208 vss.n2207 0.00233824
R3509 vss.n2528 vss.n2527 0.00233824
R3510 vss.n416 vss.n414 0.00233824
R3511 vss.n427 vss.n425 0.00233824
R3512 vss.n2536 vss.n436 0.00233824
R3513 vss.n2547 vss.n2546 0.00233824
R3514 vss.n2581 vss.n2580 0.00233824
R3515 vss.n2597 vss.n2596 0.00233824
R3516 vss.n2557 vss.n2556 0.00233824
R3517 vss.n2567 vss.n2566 0.00233824
R3518 vss.n2584 vss.n2583 0.00233824
R3519 vss.n373 vss.n372 0.00233824
R3520 vss.n380 vss.n379 0.00233824
R3521 vss.n387 vss.n386 0.00233824
R3522 vss.n2608 vss.n2606 0.00233824
R3523 vss.n2614 vss.n2612 0.00233824
R3524 vss.n395 vss.n368 0.00233824
R3525 vss.n2666 vss.n2665 0.00233824
R3526 vss.n2662 vss.n2661 0.00233824
R3527 vss.n2698 vss.n2697 0.00233824
R3528 vss.n2677 vss.n2676 0.00233824
R3529 vss.n2692 vss.n2691 0.00233824
R3530 vss.n2711 vss.n2710 0.00233824
R3531 vss.n2478 vss.n2477 0.00233824
R3532 vss.n2485 vss.n2484 0.00233824
R3533 vss.n2492 vss.n2491 0.00233824
R3534 vss.n2300 vss.n2298 0.00233824
R3535 vss.n2311 vss.n2309 0.00233824
R3536 vss.n2500 vss.n2473 0.00233824
R3537 vss.n2454 vss.n2453 0.00233824
R3538 vss.n2429 vss.n2428 0.00233824
R3539 vss.n2412 vss.n2411 0.00233824
R3540 vss.n2464 vss.n2463 0.00233824
R3541 vss.n2443 vss.n2442 0.00233824
R3542 vss.n2432 vss.n2431 0.00233824
R3543 vss.n2395 vss.n2393 0.00233824
R3544 vss.n2375 vss.n2373 0.00233824
R3545 vss.n2339 vss.n2338 0.00233824
R3546 vss.n2379 vss.n2368 0.00233824
R3547 vss.n2361 vss.n2357 0.00233824
R3548 vss.n2347 vss.n2333 0.00233824
R3549 vss.n2742 vss.n2741 0.00233824
R3550 vss.n2738 vss.n2737 0.00233824
R3551 vss.n2796 vss.n2795 0.00233824
R3552 vss.n2753 vss.n2752 0.00233824
R3553 vss.n2767 vss.n2766 0.00233824
R3554 vss.n2781 vss.n2780 0.00233824
R3555 vss.n1830 vss.n1829 0.00233824
R3556 vss.n1840 vss.n1839 0.00233824
R3557 vss.n1861 vss.n1852 0.00233824
R3558 vss.n2838 vss.n2825 0.00233824
R3559 vss.n2835 vss.n2834 0.00233824
R3560 vss.n2831 vss.n2830 0.00233824
R3561 vss.n2815 vss.n189 0.00233824
R3562 vss.n184 vss.n183 0.00233824
R3563 vss.n178 vss.n177 0.00233824
R3564 vss.n63 vss.n62 0.00231159
R3565 vss.n78 vss.n77 0.00231159
R3566 vss.n3169 vss.n3168 0.00225787
R3567 vss.n1872 vss.n1871 0.00221991
R3568 vss.n1053 vss.n1052 0.00221938
R3569 vss.n1322 vss.n1321 0.00221938
R3570 vss.n3182 vss.n3181 0.00219508
R3571 vss.n2928 vss.n2899 0.00218919
R3572 vss.n2913 vss.n2912 0.00218919
R3573 vss.n619 vss.n617 0.00218919
R3574 vss.n1208 vss.n1207 0.00218919
R3575 vss.n593 vss.n580 0.00218919
R3576 vss.n607 vss.n606 0.00218919
R3577 vss.n2146 vss.n2145 0.00217458
R3578 vss.n2145 vss.n2133 0.00217458
R3579 vss.n398 vss.n397 0.00217419
R3580 vss.n785 vss.n783 0.0021514
R3581 vss.n2073 vss.n2071 0.0021514
R3582 vss.n649 vss.n647 0.0021514
R3583 vss.n3270 vss.n3268 0.0021514
R3584 vss.n2097 vss.n2078 0.00211602
R3585 vss.n2059 vss.n2030 0.00211602
R3586 vss.n3048 vss.n3042 0.0021129
R3587 vss.n2878 vss.n141 0.00211039
R3588 vss.n1621 vss.n1620 0.00207191
R3589 vss.n1213 vss.n1212 0.00205116
R3590 vss.n1114 vss.n771 0.00203379
R3591 vss.n2921 vss.n2920 0.00200179
R3592 vss.n1782 vss.n1781 0.00198991
R3593 vss.n2919 vss.n2918 0.00196875
R3594 vss.n2954 vss.n2953 0.00196875
R3595 vss.n1185 vss.n1184 0.00196875
R3596 vss.n1180 vss.n1117 0.00196875
R3597 vss.n1133 vss.n1119 0.00196875
R3598 vss.n587 vss.n586 0.00196875
R3599 vss.n589 vss.n588 0.00196875
R3600 vss.n591 vss.n590 0.00196875
R3601 vss.n627 vss.n626 0.00196875
R3602 vss.n629 vss.n628 0.00196875
R3603 vss.n632 vss.n631 0.00196875
R3604 vss.n634 vss.n633 0.00196875
R3605 vss.n3262 vss.n3261 0.00196114
R3606 vss.n3178 vss.n3177 0.00188889
R3607 vss.n1053 vss.n1050 0.00188633
R3608 vss.n1321 vss.n1314 0.00188633
R3609 vss.n3307 vss.n3248 0.00185969
R3610 vss.n3308 vss.n3307 0.00185969
R3611 vss.n3321 vss.n3309 0.00185969
R3612 vss.n3322 vss.n3321 0.00185969
R3613 vss.n11 vss.n10 0.0018587
R3614 vss.n39 vss.n38 0.0018587
R3615 vss.n1231 vss.n1230 0.00185004
R3616 vss.n948 vss.n947 0.00182394
R3617 vss.n934 vss.n718 0.00182394
R3618 vss.n2911 vss.n2910 0.00180208
R3619 vss.n2929 vss.n2897 0.00180208
R3620 vss.n1206 vss.n1121 0.00180208
R3621 vss.n2116 vss.n594 0.00180208
R3622 vss.n605 vss.n604 0.00180208
R3623 vss.n2017 vss.n2016 0.00180208
R3624 vss.n1213 vss 0.00174092
R3625 vss.n3173 vss.n3171 0.00170184
R3626 vss.n50 vss.n49 0.00166625
R3627 vss.n102 vss.n83 0.00166625
R3628 vss.n104 vss.n102 0.00166625
R3629 vss.n104 vss.n103 0.00166625
R3630 vss.n2098 vss.n2059 0.00155801
R3631 vss.n2098 vss.n2097 0.00155801
R3632 vss.n3169 vss.n2886 0.00151772
R3633 vss.n1231 vss.n771 0.00151689
R3634 vss.n3176 vss.n3175 0.00150004
R3635 vss.n3237 vss.n3236 0.00146899
R3636 vss.n3174 vss.n3173 0.00146875
R3637 vss.n46 vss.n19 0.001433
R3638 vss.n48 vss.n47 0.001433
R3639 vss.n99 vss.n93 0.0014058
R3640 vss.n2352 vss 0.0013785
R3641 vss.n1868 vss 0.00123247
R3642 vss.n1694 vss.n1693 0.00122817
R3643 vss.n2634 vss.n401 0.00121865
R3644 vss.n2721 vss.n2720 0.00121865
R3645 vss.n3181 vss.n3180 0.00115602
R3646 vss.n3168 vss 0.00114764
R3647 vss.n3264 vss.n3263 0.00113452
R3648 vss.n2512 vss.n2511 0.00113087
R3649 vss.n776 vss.n775 0.0011215
R3650 vss.n2064 vss.n2063 0.0011215
R3651 vss.n641 vss.n640 0.0011215
R3652 vss.n3257 vss.n3256 0.0011215
R3653 vss vss.n551 0.00109494
R3654 vss.n3179 vss.n123 0.00104413
R3655 vss.n1049 vss 0.00103208
R3656 vss.n123 vss.n122 0.00100447
R3657 vss.n3273 vss.n3262 0.000987047
R3658 vss.n8 vss.n4 0.000952899
R3659 vss.n9 vss.n8 0.000952899
R3660 vss.n12 vss.n11 0.000952899
R3661 vss.n29 vss.n25 0.000952899
R3662 vss.n30 vss.n29 0.000952899
R3663 vss.n40 vss.n30 0.000952899
R3664 vss.n38 vss.n37 0.000952899
R3665 vss.n36 vss.n35 0.000952899
R3666 vss.n35 vss.n31 0.000952899
R3667 vss.n60 vss.n55 0.000952899
R3668 vss.n61 vss.n60 0.000952899
R3669 vss.n64 vss.n63 0.000952899
R3670 vss.n65 vss.n64 0.000952899
R3671 vss.n72 vss.n65 0.000952899
R3672 vss.n73 vss.n72 0.000952899
R3673 vss.n79 vss.n78 0.000952899
R3674 vss.n93 vss.n92 0.000952899
R3675 vss.n98 vss.n97 0.000952899
R3676 vss.n3174 vss.n127 0.000885246
R3677 vss.n2030 vss 0.000834917
R3678 vss.n2133 vss.n2132 0.000834917
R3679 vss vss.n1114 0.000810231
R3680 vss.n1225 vss 0.000810231
R3681 vss.n1212 vss.n1211 0.000810231
R3682 vss.n359 vss 0.000792835
R3683 vss.n3199 vss.n3198 0.000784274
R3684 vss.n3244 vss.n3243 0.000784274
R3685 vss.n949 vss.n948 0.000764789
R3686 vss.n1783 vss 0.000744156
R3687 vss.n396 vss 0.000735
R3688 vss.n140 vss 0.000722222
R3689 vss.n107 vss.n106 0.000689516
R3690 vss.n3242 vss.n3199 0.000689516
R3691 vss.n3245 vss.n3244 0.000689516
R3692 vss.n3177 vss.n3176 0.000677523
R3693 vss.n1313 vss 0.000677358
R3694 vss.n2078 vss.n2077 0.000667458
R3695 vss.n1867 vss.n1866 0.000657191
R3696 vss.n1229 vss.n1228 0.000655116
R3697 vss.n3247 vss.n3246 0.00060341
R3698 vss.n122 vss.n121 0.000548599
R3699 vss.n3179 vss.n3178 0.000518408
R3700 CAP_CTRL_CODE0[0] CAP_CTRL_CODE0[0].t0 140.376
R3701 CAP_CTRL_CODE0[0] CAP_CTRL_CODE0[0].n0 24.5005
R3702 CAP_CTRL_CODE0[0].n0 CAP_CTRL_CODE0[0] 4.42631
R3703 CAP_CTRL_CODE0[0].n0 CAP_CTRL_CODE0[0] 0.0238871
R3704 vdd.n3977 vdd.n3946 76633.3
R3705 vdd.n4644 vdd.n250 3782.21
R3706 vdd.n3922 vdd.t20 1820.83
R3707 vdd.n4005 vdd 1670.22
R3708 vdd vdd.n3835 1492.86
R3709 vdd.n7483 vdd.n212 1116.08
R3710 vdd.n3822 vdd.n3821 870.486
R3711 vdd.n49 vdd.t114 500.865
R3712 vdd.n2171 vdd.t9 470.389
R3713 vdd.n39 vdd.n38 440.25
R3714 vdd.n7485 vdd.n195 426
R3715 vdd.n7465 vdd.n226 426
R3716 vdd.n4003 vdd.n3837 423
R3717 vdd.n4619 vdd.n4585 423
R3718 vdd.n3820 vdd.t3 403.856
R3719 vdd.n2170 vdd.n2069 389.976
R3720 vdd.n172 vdd.t6 371
R3721 vdd.n3835 vdd 368.283
R3722 vdd.n3834 vdd.n2069 355.967
R3723 vdd.n3981 vdd.n3867 354
R3724 vdd.n4623 vdd.n847 354
R3725 vdd.n7510 vdd.n193 351
R3726 vdd.n7481 vdd.n214 351
R3727 vdd.n2171 vdd.n2170 344.63
R3728 vdd.t56 vdd.t46 312.889
R3729 vdd.n16 vdd.n15 308.598
R3730 vdd.n150 vdd.n149 304.122
R3731 vdd.n101 vdd.n100 302.438
R3732 vdd.n3836 vdd 288.394
R3733 vdd.n4620 vdd.t126 256.267
R3734 vdd vdd.t37 237.195
R3735 vdd.n3921 vdd.n3920 198.234
R3736 vdd.n1002 vdd.n988 198.234
R3737 vdd.n7060 vdd.n7059 198.118
R3738 vdd.n6833 vdd.n6832 198.118
R3739 vdd.n6606 vdd.n6605 198.118
R3740 vdd.n5802 vdd.n5790 198.118
R3741 vdd.n6608 vdd.n6607 198.118
R3742 vdd.n6835 vdd.n6834 198.118
R3743 vdd.n7062 vdd.n7061 198.118
R3744 vdd.n5729 vdd.n5728 198.118
R3745 vdd.n5360 vdd.n5359 198.118
R3746 vdd.n5132 vdd.n5131 198.118
R3747 vdd.n4904 vdd.n4903 198.118
R3748 vdd.n4024 vdd.n4023 198.118
R3749 vdd.n3586 vdd.n3585 198.118
R3750 vdd.n3358 vdd.n3357 198.118
R3751 vdd.n3130 vdd.n3129 198.118
R3752 vdd.n4622 vdd.t120 191.554
R3753 vdd.n7504 vdd.n193 185
R3754 vdd.n7508 vdd.n193 185
R3755 vdd.n7318 vdd.n7317 185
R3756 vdd.n5848 vdd.n5847 185
R3757 vdd.n5837 vdd.n5836 185
R3758 vdd.n5826 vdd.n5825 185
R3759 vdd.n5814 vdd.n5813 185
R3760 vdd.n7337 vdd.n7336 185
R3761 vdd.n7337 vdd.n5812 185
R3762 vdd.n7356 vdd.n7355 185
R3763 vdd.n7356 vdd.n5812 185
R3764 vdd.n7375 vdd.n7374 185
R3765 vdd.n7375 vdd.n5812 185
R3766 vdd.n7398 vdd.n7397 185
R3767 vdd.n5801 vdd.n5800 185
R3768 vdd.n7299 vdd.n5859 185
R3769 vdd.n6410 vdd.n6409 185
R3770 vdd.n6360 vdd.n6359 185
R3771 vdd.n6459 vdd.n6458 185
R3772 vdd.n6478 vdd.n6347 185
R3773 vdd.n6496 vdd.n6495 185
R3774 vdd.n6516 vdd.n6313 185
R3775 vdd.n6515 vdd.n6316 185
R3776 vdd.n6519 vdd.n6315 185
R3777 vdd.n6314 vdd.n6299 185
R3778 vdd.n6555 vdd.n6554 185
R3779 vdd.n6552 vdd.n6298 185
R3780 vdd.n6582 vdd.n6581 185
R3781 vdd.n6584 vdd.n6280 185
R3782 vdd.n6603 vdd.n6602 185
R3783 vdd.n6270 vdd.n6269 185
R3784 vdd.n6609 vdd.n6268 185
R3785 vdd.n6242 vdd.n6241 185
R3786 vdd.n6227 vdd.n6226 185
R3787 vdd.n6686 vdd.n6685 185
R3788 vdd.n6705 vdd.n6214 185
R3789 vdd.n6723 vdd.n6722 185
R3790 vdd.n6743 vdd.n6180 185
R3791 vdd.n6742 vdd.n6183 185
R3792 vdd.n6746 vdd.n6182 185
R3793 vdd.n6181 vdd.n6166 185
R3794 vdd.n6782 vdd.n6781 185
R3795 vdd.n6779 vdd.n6165 185
R3796 vdd.n6809 vdd.n6808 185
R3797 vdd.n6811 vdd.n6147 185
R3798 vdd.n6830 vdd.n6829 185
R3799 vdd.n6137 vdd.n6136 185
R3800 vdd.n6836 vdd.n6135 185
R3801 vdd.n6109 vdd.n6108 185
R3802 vdd.n6094 vdd.n6093 185
R3803 vdd.n6913 vdd.n6912 185
R3804 vdd.n6932 vdd.n6081 185
R3805 vdd.n6950 vdd.n6949 185
R3806 vdd.n6970 vdd.n6047 185
R3807 vdd.n6969 vdd.n6050 185
R3808 vdd.n6973 vdd.n6049 185
R3809 vdd.n6048 vdd.n6033 185
R3810 vdd.n7009 vdd.n7008 185
R3811 vdd.n7006 vdd.n6032 185
R3812 vdd.n7036 vdd.n7035 185
R3813 vdd.n7038 vdd.n6014 185
R3814 vdd.n7057 vdd.n7056 185
R3815 vdd.n6004 vdd.n6003 185
R3816 vdd.n7063 vdd.n6002 185
R3817 vdd.n5976 vdd.n5975 185
R3818 vdd.n5961 vdd.n5960 185
R3819 vdd.n7140 vdd.n7139 185
R3820 vdd.n7159 vdd.n5948 185
R3821 vdd.n7177 vdd.n7176 185
R3822 vdd.n7197 vdd.n5914 185
R3823 vdd.n7196 vdd.n5917 185
R3824 vdd.n7200 vdd.n5916 185
R3825 vdd.n5915 vdd.n5900 185
R3826 vdd.n7236 vdd.n7235 185
R3827 vdd.n7233 vdd.n5899 185
R3828 vdd.n7263 vdd.n7262 185
R3829 vdd.n7265 vdd.n5881 185
R3830 vdd.n7289 vdd.n7288 185
R3831 vdd.n5870 vdd.n5869 185
R3832 vdd.n7157 vdd.n7156 185
R3833 vdd.n7137 vdd.n5959 185
R3834 vdd.n7112 vdd.n7111 185
R3835 vdd.n7091 vdd.n7090 185
R3836 vdd.n7178 vdd.n5928 185
R3837 vdd.n5987 vdd.n5986 185
R3838 vdd.n6930 vdd.n6929 185
R3839 vdd.n6910 vdd.n6092 185
R3840 vdd.n6885 vdd.n6884 185
R3841 vdd.n6864 vdd.n6863 185
R3842 vdd.n6951 vdd.n6061 185
R3843 vdd.n6120 vdd.n6119 185
R3844 vdd.n6703 vdd.n6702 185
R3845 vdd.n6683 vdd.n6225 185
R3846 vdd.n6658 vdd.n6657 185
R3847 vdd.n6637 vdd.n6636 185
R3848 vdd.n6724 vdd.n6194 185
R3849 vdd.n6253 vdd.n6252 185
R3850 vdd.n6476 vdd.n6475 185
R3851 vdd.n6456 vdd.n6358 185
R3852 vdd.n6431 vdd.n6430 185
R3853 vdd.n6497 vdd.n6327 185
R3854 vdd.n6408 vdd.n6375 185
R3855 vdd.n2169 vdd.n2167 185
R3856 vdd.n2923 vdd.n2773 185
R3857 vdd.n2952 vdd.n2951 185
R3858 vdd.n2746 vdd.n2745 185
R3859 vdd.n2986 vdd.n2985 185
R3860 vdd.n3004 vdd.n3003 185
R3861 vdd.n2719 vdd.n2701 185
R3862 vdd.n3035 vdd.n2700 185
R3863 vdd.n3065 vdd.n3064 185
R3864 vdd.n2668 vdd.n2667 185
R3865 vdd.n3093 vdd.n3092 185
R3866 vdd.n3151 vdd.n2638 185
R3867 vdd.n3180 vdd.n3179 185
R3868 vdd.n2611 vdd.n2610 185
R3869 vdd.n3214 vdd.n3213 185
R3870 vdd.n3232 vdd.n3231 185
R3871 vdd.n2584 vdd.n2566 185
R3872 vdd.n3263 vdd.n2565 185
R3873 vdd.n3293 vdd.n3292 185
R3874 vdd.n2533 vdd.n2532 185
R3875 vdd.n3321 vdd.n3320 185
R3876 vdd.n3379 vdd.n2503 185
R3877 vdd.n3408 vdd.n3407 185
R3878 vdd.n2476 vdd.n2475 185
R3879 vdd.n3442 vdd.n3441 185
R3880 vdd.n3460 vdd.n3459 185
R3881 vdd.n2449 vdd.n2431 185
R3882 vdd.n3491 vdd.n2430 185
R3883 vdd.n3521 vdd.n3520 185
R3884 vdd.n2398 vdd.n2397 185
R3885 vdd.n3549 vdd.n3548 185
R3886 vdd.n3607 vdd.n2368 185
R3887 vdd.n3636 vdd.n3635 185
R3888 vdd.n2341 vdd.n2340 185
R3889 vdd.n3670 vdd.n3669 185
R3890 vdd.n3687 vdd.n3686 185
R3891 vdd.n3708 vdd.n2298 185
R3892 vdd.n3727 vdd.n2297 185
R3893 vdd.n2296 vdd.n2294 185
R3894 vdd.n3762 vdd.n2277 185
R3895 vdd.n3796 vdd.n3795 185
R3896 vdd.n3798 vdd.n2257 185
R3897 vdd.n3765 vdd.n3764 185
R3898 vdd.n2293 vdd.n2278 185
R3899 vdd.n3728 vdd.n2292 185
R3900 vdd.n3707 vdd.n3706 185
R3901 vdd.n3667 vdd.n2339 185
R3902 vdd.n3641 vdd.n3640 185
R3903 vdd.n3634 vdd.n2356 185
R3904 vdd.n3605 vdd.n3604 185
R3905 vdd.n3689 vdd.n2319 185
R3906 vdd.n3588 vdd.n3587 185
R3907 vdd.n3550 vdd.n2380 185
R3908 vdd.n3544 vdd.n3543 185
R3909 vdd.n3523 vdd.n2412 185
R3910 vdd.n3494 vdd.n3493 185
R3911 vdd.n3584 vdd.n3583 185
R3912 vdd.n3583 vdd.n2065 185
R3913 vdd.n3582 vdd.n2379 185
R3914 vdd.n2452 vdd.n2450 185
R3915 vdd.n3439 vdd.n2474 185
R3916 vdd.n3413 vdd.n3412 185
R3917 vdd.n3406 vdd.n2491 185
R3918 vdd.n3377 vdd.n3376 185
R3919 vdd.n3462 vdd.n2445 185
R3920 vdd.n3360 vdd.n3359 185
R3921 vdd.n3322 vdd.n2515 185
R3922 vdd.n3316 vdd.n3315 185
R3923 vdd.n3295 vdd.n2547 185
R3924 vdd.n3266 vdd.n3265 185
R3925 vdd.n3356 vdd.n3355 185
R3926 vdd.n3355 vdd.n2065 185
R3927 vdd.n3354 vdd.n2514 185
R3928 vdd.n2587 vdd.n2585 185
R3929 vdd.n3211 vdd.n2609 185
R3930 vdd.n3185 vdd.n3184 185
R3931 vdd.n3178 vdd.n2626 185
R3932 vdd.n3149 vdd.n3148 185
R3933 vdd.n3234 vdd.n2580 185
R3934 vdd.n3132 vdd.n3131 185
R3935 vdd.n3094 vdd.n2650 185
R3936 vdd.n3088 vdd.n3087 185
R3937 vdd.n3067 vdd.n2682 185
R3938 vdd.n3038 vdd.n3037 185
R3939 vdd.n3128 vdd.n3127 185
R3940 vdd.n3127 vdd.n2065 185
R3941 vdd.n3126 vdd.n2649 185
R3942 vdd.n2722 vdd.n2720 185
R3943 vdd.n2983 vdd.n2744 185
R3944 vdd.n2957 vdd.n2956 185
R3945 vdd.n2921 vdd.n2920 185
R3946 vdd.n2950 vdd.n2761 185
R3947 vdd.n3006 vdd.n2715 185
R3948 vdd.n4015 vdd.n4014 185
R3949 vdd.n2826 vdd.n2057 185
R3950 vdd.n2852 vdd.n2851 185
R3951 vdd.n2872 vdd.n2871 185
R3952 vdd.n2881 vdd.n2880 185
R3953 vdd.n4022 vdd.n2067 185
R3954 vdd.n2056 vdd.n2054 185
R3955 vdd.n2807 vdd.n2806 185
R3956 vdd.n2854 vdd.n2853 185
R3957 vdd.n2874 vdd.n2873 185
R3958 vdd.n2879 vdd.n2878 185
R3959 vdd.n3982 vdd.n3981 185
R3960 vdd.n3981 vdd.n3980 185
R3961 vdd.n4521 vdd.n4520 185
R3962 vdd.n4522 vdd.n4521 185
R3963 vdd.n1061 vdd.n1060 185
R3964 vdd.n1060 vdd.n1059 185
R3965 vdd.n1051 vdd.n1049 185
R3966 vdd.n1071 vdd.n1051 185
R3967 vdd.n4494 vdd.n4493 185
R3968 vdd.n4495 vdd.n4494 185
R3969 vdd.n1125 vdd.n1124 185
R3970 vdd.n1124 vdd.n1123 185
R3971 vdd.n4469 vdd.n4468 185
R3972 vdd.n4470 vdd.n4469 185
R3973 vdd.n1181 vdd.n1180 185
R3974 vdd.n1182 vdd.n1181 185
R3975 vdd.n1170 vdd.n1168 185
R3976 vdd.n4449 vdd.n1170 185
R3977 vdd.n1223 vdd.n1222 185
R3978 vdd.n1224 vdd.n1223 185
R3979 vdd.n1212 vdd.n1210 185
R3980 vdd.n4427 vdd.n1212 185
R3981 vdd.n1269 vdd.n1268 185
R3982 vdd.n1270 vdd.n1269 185
R3983 vdd.n4400 vdd.n4399 185
R3984 vdd.n4401 vdd.n4400 185
R3985 vdd.n1325 vdd.n1324 185
R3986 vdd.n1324 vdd.n1323 185
R3987 vdd.n1315 vdd.n1313 185
R3988 vdd.n1335 vdd.n1315 185
R3989 vdd.n4373 vdd.n4372 185
R3990 vdd.n4374 vdd.n4373 185
R3991 vdd.n1389 vdd.n1388 185
R3992 vdd.n1388 vdd.n1387 185
R3993 vdd.n4348 vdd.n4347 185
R3994 vdd.n4349 vdd.n4348 185
R3995 vdd.n1445 vdd.n1444 185
R3996 vdd.n1446 vdd.n1445 185
R3997 vdd.n1434 vdd.n1432 185
R3998 vdd.n4328 vdd.n1434 185
R3999 vdd.n1487 vdd.n1486 185
R4000 vdd.n1488 vdd.n1487 185
R4001 vdd.n1476 vdd.n1474 185
R4002 vdd.n4306 vdd.n1476 185
R4003 vdd.n1533 vdd.n1532 185
R4004 vdd.n1534 vdd.n1533 185
R4005 vdd.n4279 vdd.n4278 185
R4006 vdd.n4280 vdd.n4279 185
R4007 vdd.n1589 vdd.n1588 185
R4008 vdd.n1588 vdd.n1587 185
R4009 vdd.n1579 vdd.n1577 185
R4010 vdd.n1599 vdd.n1579 185
R4011 vdd.n4252 vdd.n4251 185
R4012 vdd.n4253 vdd.n4252 185
R4013 vdd.n1653 vdd.n1652 185
R4014 vdd.n1652 vdd.n1651 185
R4015 vdd.n4227 vdd.n4226 185
R4016 vdd.n4228 vdd.n4227 185
R4017 vdd.n1709 vdd.n1708 185
R4018 vdd.n1710 vdd.n1709 185
R4019 vdd.n1698 vdd.n1696 185
R4020 vdd.n4207 vdd.n1698 185
R4021 vdd.n1751 vdd.n1750 185
R4022 vdd.n1752 vdd.n1751 185
R4023 vdd.n1740 vdd.n1738 185
R4024 vdd.n4185 vdd.n1740 185
R4025 vdd.n1797 vdd.n1796 185
R4026 vdd.n1798 vdd.n1797 185
R4027 vdd.n4158 vdd.n4157 185
R4028 vdd.n4159 vdd.n4158 185
R4029 vdd.n1853 vdd.n1852 185
R4030 vdd.n1852 vdd.n1851 185
R4031 vdd.n1843 vdd.n1841 185
R4032 vdd.n1863 vdd.n1843 185
R4033 vdd.n4131 vdd.n4130 185
R4034 vdd.n4132 vdd.n4131 185
R4035 vdd.n1917 vdd.n1916 185
R4036 vdd.n1916 vdd.n1915 185
R4037 vdd.n4106 vdd.n4105 185
R4038 vdd.n4107 vdd.n4106 185
R4039 vdd.n1973 vdd.n1972 185
R4040 vdd.n1974 vdd.n1973 185
R4041 vdd.n1962 vdd.n1960 185
R4042 vdd.n4086 vdd.n1962 185
R4043 vdd.n2015 vdd.n2014 185
R4044 vdd.n2016 vdd.n2015 185
R4045 vdd.n2004 vdd.n2002 185
R4046 vdd.n4064 vdd.n2004 185
R4047 vdd.n4062 vdd.n4061 185
R4048 vdd.n4063 vdd.n4062 185
R4049 vdd.n2013 vdd.n2003 185
R4050 vdd.n2017 vdd.n2003 185
R4051 vdd.n4084 vdd.n4083 185
R4052 vdd.n4085 vdd.n4084 185
R4053 vdd.n1971 vdd.n1961 185
R4054 vdd.n1975 vdd.n1961 185
R4055 vdd.n3918 vdd.n3917 185
R4056 vdd.n1911 vdd.n1910 185
R4057 vdd.n4108 vdd.n1911 185
R4058 vdd.n1866 vdd.n1844 185
R4059 vdd.n4133 vdd.n1844 185
R4060 vdd.n1861 vdd.n1860 185
R4061 vdd.n1862 vdd.n1861 185
R4062 vdd.n1849 vdd.n1848 185
R4063 vdd.n1850 vdd.n1849 185
R4064 vdd.n1802 vdd.n1788 185
R4065 vdd.n4160 vdd.n1788 185
R4066 vdd.n1918 vdd.n1913 185
R4067 vdd.n1913 vdd.n1912 185
R4068 vdd.n1787 vdd.n1785 185
R4069 vdd.n1799 vdd.n1787 185
R4070 vdd.n4183 vdd.n4182 185
R4071 vdd.n4184 vdd.n4183 185
R4072 vdd.n1749 vdd.n1739 185
R4073 vdd.n1753 vdd.n1739 185
R4074 vdd.n4205 vdd.n4204 185
R4075 vdd.n4206 vdd.n4205 185
R4076 vdd.n1707 vdd.n1697 185
R4077 vdd.n1711 vdd.n1697 185
R4078 vdd.n1795 vdd.n1794 185
R4079 vdd.n1794 vdd.n1793 185
R4080 vdd.n1791 vdd.n1790 185
R4081 vdd.n1792 vdd.n1791 185
R4082 vdd.n1647 vdd.n1646 185
R4083 vdd.n4229 vdd.n1647 185
R4084 vdd.n1602 vdd.n1580 185
R4085 vdd.n4254 vdd.n1580 185
R4086 vdd.n1597 vdd.n1596 185
R4087 vdd.n1598 vdd.n1597 185
R4088 vdd.n1585 vdd.n1584 185
R4089 vdd.n1586 vdd.n1585 185
R4090 vdd.n1538 vdd.n1524 185
R4091 vdd.n4281 vdd.n1524 185
R4092 vdd.n1654 vdd.n1649 185
R4093 vdd.n1649 vdd.n1648 185
R4094 vdd.n1523 vdd.n1521 185
R4095 vdd.n1535 vdd.n1523 185
R4096 vdd.n4304 vdd.n4303 185
R4097 vdd.n4305 vdd.n4304 185
R4098 vdd.n1485 vdd.n1475 185
R4099 vdd.n1489 vdd.n1475 185
R4100 vdd.n4326 vdd.n4325 185
R4101 vdd.n4327 vdd.n4326 185
R4102 vdd.n1443 vdd.n1433 185
R4103 vdd.n1447 vdd.n1433 185
R4104 vdd.n1531 vdd.n1530 185
R4105 vdd.n1530 vdd.n1529 185
R4106 vdd.n1527 vdd.n1526 185
R4107 vdd.n1528 vdd.n1527 185
R4108 vdd.n1383 vdd.n1382 185
R4109 vdd.n4350 vdd.n1383 185
R4110 vdd.n1338 vdd.n1316 185
R4111 vdd.n4375 vdd.n1316 185
R4112 vdd.n1333 vdd.n1332 185
R4113 vdd.n1334 vdd.n1333 185
R4114 vdd.n1321 vdd.n1320 185
R4115 vdd.n1322 vdd.n1321 185
R4116 vdd.n1274 vdd.n1260 185
R4117 vdd.n4402 vdd.n1260 185
R4118 vdd.n1390 vdd.n1385 185
R4119 vdd.n1385 vdd.n1384 185
R4120 vdd.n1259 vdd.n1257 185
R4121 vdd.n1271 vdd.n1259 185
R4122 vdd.n4425 vdd.n4424 185
R4123 vdd.n4426 vdd.n4425 185
R4124 vdd.n1221 vdd.n1211 185
R4125 vdd.n1225 vdd.n1211 185
R4126 vdd.n4447 vdd.n4446 185
R4127 vdd.n4448 vdd.n4447 185
R4128 vdd.n1179 vdd.n1169 185
R4129 vdd.n1183 vdd.n1169 185
R4130 vdd.n1267 vdd.n1266 185
R4131 vdd.n1266 vdd.n1265 185
R4132 vdd.n1263 vdd.n1262 185
R4133 vdd.n1264 vdd.n1263 185
R4134 vdd.n1119 vdd.n1118 185
R4135 vdd.n4471 vdd.n1119 185
R4136 vdd.n1074 vdd.n1052 185
R4137 vdd.n4496 vdd.n1052 185
R4138 vdd.n1069 vdd.n1068 185
R4139 vdd.n1070 vdd.n1069 185
R4140 vdd.n1006 vdd.n991 185
R4141 vdd.n4523 vdd.n991 185
R4142 vdd.n1057 vdd.n1056 185
R4143 vdd.n1058 vdd.n1057 185
R4144 vdd.n1126 vdd.n1121 185
R4145 vdd.n1121 vdd.n1120 185
R4146 vdd.n1003 vdd.n990 185
R4147 vdd.n4581 vdd.n4580 185
R4148 vdd.n4582 vdd.n4581 185
R4149 vdd.n858 vdd.n855 185
R4150 vdd.n4575 vdd.n855 185
R4151 vdd.n930 vdd.n929 185
R4152 vdd.n931 vdd.n930 185
R4153 vdd.n942 vdd.n941 185
R4154 vdd.n943 vdd.n942 185
R4155 vdd.n947 vdd.n925 185
R4156 vdd.n4548 vdd.n925 185
R4157 vdd.n997 vdd.n996 185
R4158 vdd.n996 vdd.n995 185
R4159 vdd.n4579 vdd.n852 185
R4160 vdd.n852 vdd.n851 185
R4161 vdd.n4573 vdd.n4572 185
R4162 vdd.n4574 vdd.n4573 185
R4163 vdd.n934 vdd.n933 185
R4164 vdd.n933 vdd.n932 185
R4165 vdd.n924 vdd.n922 185
R4166 vdd.n944 vdd.n924 185
R4167 vdd.n4546 vdd.n4545 185
R4168 vdd.n4547 vdd.n4546 185
R4169 vdd.n998 vdd.n993 185
R4170 vdd.n993 vdd.n992 185
R4171 vdd.n4624 vdd.n4623 185
R4172 vdd.n4623 vdd.n4622 185
R4173 vdd.n4697 vdd.n797 185
R4174 vdd.n4726 vdd.n4725 185
R4175 vdd.n770 vdd.n769 185
R4176 vdd.n4760 vdd.n4759 185
R4177 vdd.n4778 vdd.n4777 185
R4178 vdd.n743 vdd.n725 185
R4179 vdd.n4809 vdd.n724 185
R4180 vdd.n4839 vdd.n4838 185
R4181 vdd.n692 vdd.n691 185
R4182 vdd.n4867 vdd.n4866 185
R4183 vdd.n4925 vdd.n662 185
R4184 vdd.n4954 vdd.n4953 185
R4185 vdd.n635 vdd.n634 185
R4186 vdd.n4988 vdd.n4987 185
R4187 vdd.n5006 vdd.n5005 185
R4188 vdd.n608 vdd.n590 185
R4189 vdd.n5037 vdd.n589 185
R4190 vdd.n5067 vdd.n5066 185
R4191 vdd.n557 vdd.n556 185
R4192 vdd.n5095 vdd.n5094 185
R4193 vdd.n5153 vdd.n527 185
R4194 vdd.n5182 vdd.n5181 185
R4195 vdd.n500 vdd.n499 185
R4196 vdd.n5216 vdd.n5215 185
R4197 vdd.n5234 vdd.n5233 185
R4198 vdd.n473 vdd.n455 185
R4199 vdd.n5265 vdd.n454 185
R4200 vdd.n5295 vdd.n5294 185
R4201 vdd.n422 vdd.n421 185
R4202 vdd.n5323 vdd.n5322 185
R4203 vdd.n5381 vdd.n392 185
R4204 vdd.n5410 vdd.n5409 185
R4205 vdd.n365 vdd.n364 185
R4206 vdd.n5444 vdd.n5443 185
R4207 vdd.n5461 vdd.n5460 185
R4208 vdd.n5483 vdd.n324 185
R4209 vdd.n5503 vdd.n323 185
R4210 vdd.n322 vdd.n320 185
R4211 vdd.n5538 vdd.n303 185
R4212 vdd.n5572 vdd.n5571 185
R4213 vdd.n5574 vdd.n283 185
R4214 vdd.n5541 vdd.n5540 185
R4215 vdd.n319 vdd.n304 185
R4216 vdd.n5504 vdd.n318 185
R4217 vdd.n5482 vdd.n5481 185
R4218 vdd.n5441 vdd.n363 185
R4219 vdd.n5415 vdd.n5414 185
R4220 vdd.n5408 vdd.n380 185
R4221 vdd.n5379 vdd.n5378 185
R4222 vdd.n5463 vdd.n343 185
R4223 vdd.n5362 vdd.n5361 185
R4224 vdd.n5324 vdd.n404 185
R4225 vdd.n5318 vdd.n5317 185
R4226 vdd.n5297 vdd.n436 185
R4227 vdd.n5268 vdd.n5267 185
R4228 vdd.n5358 vdd.n5357 185
R4229 vdd.n5357 vdd.n250 185
R4230 vdd.n5356 vdd.n403 185
R4231 vdd.n476 vdd.n474 185
R4232 vdd.n5213 vdd.n498 185
R4233 vdd.n5187 vdd.n5186 185
R4234 vdd.n5180 vdd.n515 185
R4235 vdd.n5151 vdd.n5150 185
R4236 vdd.n5236 vdd.n469 185
R4237 vdd.n5134 vdd.n5133 185
R4238 vdd.n5096 vdd.n539 185
R4239 vdd.n5090 vdd.n5089 185
R4240 vdd.n5069 vdd.n571 185
R4241 vdd.n5040 vdd.n5039 185
R4242 vdd.n5130 vdd.n5129 185
R4243 vdd.n5129 vdd.n250 185
R4244 vdd.n5128 vdd.n538 185
R4245 vdd.n611 vdd.n609 185
R4246 vdd.n4985 vdd.n633 185
R4247 vdd.n4959 vdd.n4958 185
R4248 vdd.n4952 vdd.n650 185
R4249 vdd.n4923 vdd.n4922 185
R4250 vdd.n5008 vdd.n604 185
R4251 vdd.n4906 vdd.n4905 185
R4252 vdd.n4868 vdd.n674 185
R4253 vdd.n4862 vdd.n4861 185
R4254 vdd.n4841 vdd.n706 185
R4255 vdd.n4812 vdd.n4811 185
R4256 vdd.n4902 vdd.n4901 185
R4257 vdd.n4901 vdd.n250 185
R4258 vdd.n4900 vdd.n673 185
R4259 vdd.n746 vdd.n744 185
R4260 vdd.n4757 vdd.n768 185
R4261 vdd.n4731 vdd.n4730 185
R4262 vdd.n4695 vdd.n4694 185
R4263 vdd.n4724 vdd.n785 185
R4264 vdd.n4780 vdd.n739 185
R4265 vdd.n5723 vdd.n5722 185
R4266 vdd.n265 vdd.n264 185
R4267 vdd.n5621 vdd.n5620 185
R4268 vdd.n5698 vdd.n5697 185
R4269 vdd.n5668 vdd.n5667 185
R4270 vdd.n5670 vdd.n5669 185
R4271 vdd.n5696 vdd.n253 185
R4272 vdd.n5727 vdd.n253 185
R4273 vdd.n5622 vdd.n257 185
R4274 vdd.n5727 vdd.n257 185
R4275 vdd.n5612 vdd.n251 185
R4276 vdd.n5727 vdd.n251 185
R4277 vdd.n249 vdd.n248 185
R4278 vdd.n5724 vdd.n260 185
R4279 vdd.n224 vdd.n214 185
R4280 vdd.n7462 vdd.n214 185
R4281 vdd.n4584 vdd 165.668
R4282 vdd.n25 vdd.n24 165.252
R4283 vdd.n55 vdd.n54 160.918
R4284 vdd.n2101 vdd.t45 158.06
R4285 vdd.n7512 vdd.t43 152.88
R4286 vdd.n7479 vdd.t111 152.88
R4287 vdd.n7 vdd.t84 152.88
R4288 vdd.n164 vdd.t129 152.88
R4289 vdd.n211 vdd.t66 152.879
R4290 vdd.n3854 vdd.t131 152.879
R4291 vdd.n4001 vdd.t109 152.879
R4292 vdd.n844 vdd.t121 152.879
R4293 vdd.n4609 vdd.t127 152.879
R4294 vdd.n5752 vdd.t118 152.879
R4295 vdd.n2206 vdd.t77 151.633
R4296 vdd.n2171 vdd.t52 150.648
R4297 vdd.n2212 vdd.t64 149.696
R4298 vdd.n2105 vdd.t132 140.375
R4299 vdd.n2172 vdd 135.256
R4300 vdd.n1002 vdd 131.415
R4301 vdd.t120 vdd.n849 113.897
R4302 vdd.n5575 vdd.n5574 111.234
R4303 vdd.n3799 vdd.n3798 111.234
R4304 vdd.n4695 vdd.n798 111.234
R4305 vdd.n2921 vdd.n2774 111.234
R4306 vdd.n7231 vdd.n5900 111.177
R4307 vdd.n7267 vdd.n7265 111.177
R4308 vdd.n7090 vdd.n7088 111.177
R4309 vdd.n7111 vdd.n7109 111.177
R4310 vdd.n7137 vdd.n7136 111.177
R4311 vdd.n7157 vdd.n5949 111.177
R4312 vdd.n7004 vdd.n6033 111.177
R4313 vdd.n7040 vdd.n7038 111.177
R4314 vdd.n6863 vdd.n6861 111.177
R4315 vdd.n6884 vdd.n6882 111.177
R4316 vdd.n6910 vdd.n6909 111.177
R4317 vdd.n6930 vdd.n6082 111.177
R4318 vdd.n6777 vdd.n6166 111.177
R4319 vdd.n6813 vdd.n6811 111.177
R4320 vdd.n6636 vdd.n6634 111.177
R4321 vdd.n6657 vdd.n6655 111.177
R4322 vdd.n6683 vdd.n6682 111.177
R4323 vdd.n6703 vdd.n6215 111.177
R4324 vdd.n6550 vdd.n6299 111.177
R4325 vdd.n6586 vdd.n6584 111.177
R4326 vdd.n6430 vdd.n6428 111.177
R4327 vdd.n6456 vdd.n6455 111.177
R4328 vdd.n6476 vdd.n6348 111.177
R4329 vdd.n7320 vdd.n7318 111.177
R4330 vdd.n7339 vdd.n7337 111.177
R4331 vdd.n7358 vdd.n7356 111.177
R4332 vdd.n7377 vdd.n7375 111.177
R4333 vdd.n5722 vdd.n5721 111.177
R4334 vdd.n5618 vdd.n251 111.177
R4335 vdd.n5699 vdd.n257 111.177
R4336 vdd.n5665 vdd.n253 111.177
R4337 vdd.n5501 vdd.n324 111.177
R4338 vdd.n5536 vdd.n304 111.177
R4339 vdd.n5379 vdd.n393 111.177
R4340 vdd.n5414 vdd.n5412 111.177
R4341 vdd.n5461 vdd.n353 111.177
R4342 vdd.n5263 vdd.n455 111.177
R4343 vdd.n5299 vdd.n5297 111.177
R4344 vdd.n5354 vdd.n404 111.177
R4345 vdd.n5151 vdd.n528 111.177
R4346 vdd.n5186 vdd.n5184 111.177
R4347 vdd.n5234 vdd.n488 111.177
R4348 vdd.n5035 vdd.n590 111.177
R4349 vdd.n5071 vdd.n5069 111.177
R4350 vdd.n5126 vdd.n539 111.177
R4351 vdd.n4923 vdd.n663 111.177
R4352 vdd.n4958 vdd.n4956 111.177
R4353 vdd.n5006 vdd.n623 111.177
R4354 vdd.n4807 vdd.n725 111.177
R4355 vdd.n4843 vdd.n4841 111.177
R4356 vdd.n4898 vdd.n674 111.177
R4357 vdd.n4730 vdd.n4728 111.177
R4358 vdd.n4778 vdd.n758 111.177
R4359 vdd.n4577 vdd.n855 111.177
R4360 vdd.n930 vdd.n857 111.177
R4361 vdd.n942 vdd.n927 111.177
R4362 vdd.n4550 vdd.n925 111.177
R4363 vdd.n996 vdd.n946 111.177
R4364 vdd.n4106 vdd.n1935 111.177
R4365 vdd.n4088 vdd.n1961 111.177
R4366 vdd.n4084 vdd.n1977 111.177
R4367 vdd.n4066 vdd.n2003 111.177
R4368 vdd.n4062 vdd.n2019 111.177
R4369 vdd.n4162 vdd.n1788 111.177
R4370 vdd.n1849 vdd.n1801 111.177
R4371 vdd.n1861 vdd.n1846 111.177
R4372 vdd.n4135 vdd.n1844 111.177
R4373 vdd.n1916 vdd.n1865 111.177
R4374 vdd.n4227 vdd.n1671 111.177
R4375 vdd.n4209 vdd.n1697 111.177
R4376 vdd.n4205 vdd.n1713 111.177
R4377 vdd.n4187 vdd.n1739 111.177
R4378 vdd.n4183 vdd.n1755 111.177
R4379 vdd.n4283 vdd.n1524 111.177
R4380 vdd.n1585 vdd.n1537 111.177
R4381 vdd.n1597 vdd.n1582 111.177
R4382 vdd.n4256 vdd.n1580 111.177
R4383 vdd.n1652 vdd.n1601 111.177
R4384 vdd.n4348 vdd.n1407 111.177
R4385 vdd.n4330 vdd.n1433 111.177
R4386 vdd.n4326 vdd.n1449 111.177
R4387 vdd.n4308 vdd.n1475 111.177
R4388 vdd.n4304 vdd.n1491 111.177
R4389 vdd.n4404 vdd.n1260 111.177
R4390 vdd.n1321 vdd.n1273 111.177
R4391 vdd.n1333 vdd.n1318 111.177
R4392 vdd.n4377 vdd.n1316 111.177
R4393 vdd.n1388 vdd.n1337 111.177
R4394 vdd.n4469 vdd.n1143 111.177
R4395 vdd.n4451 vdd.n1169 111.177
R4396 vdd.n4447 vdd.n1185 111.177
R4397 vdd.n4429 vdd.n1211 111.177
R4398 vdd.n4425 vdd.n1227 111.177
R4399 vdd.n4525 vdd.n991 111.177
R4400 vdd.n1057 vdd.n1005 111.177
R4401 vdd.n1069 vdd.n1054 111.177
R4402 vdd.n4498 vdd.n1052 111.177
R4403 vdd.n1124 vdd.n1073 111.177
R4404 vdd.n4014 vdd.n2066 111.177
R4405 vdd.n2851 vdd.n2850 111.177
R4406 vdd.n2882 vdd.n2881 111.177
R4407 vdd.n3725 vdd.n2298 111.177
R4408 vdd.n3760 vdd.n2278 111.177
R4409 vdd.n3605 vdd.n2369 111.177
R4410 vdd.n3640 vdd.n3638 111.177
R4411 vdd.n3687 vdd.n2329 111.177
R4412 vdd.n3489 vdd.n2431 111.177
R4413 vdd.n3525 vdd.n3523 111.177
R4414 vdd.n3580 vdd.n2380 111.177
R4415 vdd.n3377 vdd.n2504 111.177
R4416 vdd.n3412 vdd.n3410 111.177
R4417 vdd.n3460 vdd.n2464 111.177
R4418 vdd.n3261 vdd.n2566 111.177
R4419 vdd.n3297 vdd.n3295 111.177
R4420 vdd.n3352 vdd.n2515 111.177
R4421 vdd.n3149 vdd.n2639 111.177
R4422 vdd.n3184 vdd.n3182 111.177
R4423 vdd.n3232 vdd.n2599 111.177
R4424 vdd.n3033 vdd.n2701 111.177
R4425 vdd.n3069 vdd.n3067 111.177
R4426 vdd.n3124 vdd.n2650 111.177
R4427 vdd.n2956 vdd.n2954 111.177
R4428 vdd.n3004 vdd.n2734 111.177
R4429 vdd.n4584 vdd.t126 108.719
R4430 vdd vdd.n168 105.715
R4431 vdd.n26 vdd.t58 102.957
R4432 vdd.n2171 vdd.t122 99.1309
R4433 vdd.n2182 vdd.t51 99.0968
R4434 vdd.t65 vdd.n194 98.5482
R4435 vdd.n2171 vdd.t56 97.4945
R4436 vdd.n30 vdd.t17 95.9365
R4437 vdd vdd.n7483 92.6353
R4438 vdd.n7506 vdd.n7505 92.5005
R4439 vdd.n7507 vdd.n7506 92.5005
R4440 vdd.n7511 vdd.n7510 92.5005
R4441 vdd.n7510 vdd.n7509 92.5005
R4442 vdd.n7486 vdd.n7485 92.5005
R4443 vdd.n7485 vdd.n7484 92.5005
R4444 vdd.n3868 vdd.n3866 92.5005
R4445 vdd.n3979 vdd.n3868 92.5005
R4446 vdd.n4003 vdd.n4002 92.5005
R4447 vdd.n4004 vdd.n4003 92.5005
R4448 vdd.n3867 vdd.n3855 92.5005
R4449 vdd.n3945 vdd.n3867 92.5005
R4450 vdd.n847 vdd.n845 92.5005
R4451 vdd.n849 vdd.n847 92.5005
R4452 vdd.n4621 vdd.n848 92.5005
R4453 vdd.n848 vdd.n846 92.5005
R4454 vdd.n4610 vdd.n4585 92.5005
R4455 vdd.n4585 vdd.n4584 92.5005
R4456 vdd.n7481 vdd.n7480 92.5005
R4457 vdd.n7482 vdd.n7481 92.5005
R4458 vdd.n5753 vdd.n226 92.5005
R4459 vdd.n4643 vdd.n226 92.5005
R4460 vdd.n227 vdd.n225 92.5005
R4461 vdd.n7463 vdd.n227 92.5005
R4462 vdd.n161 vdd.n160 92.5005
R4463 vdd.n160 vdd.n159 92.5005
R4464 vdd.n176 vdd.n175 92.5005
R4465 vdd.n175 vdd.n174 92.5005
R4466 vdd.n171 vdd.n170 92.5005
R4467 vdd.n170 vdd.n169 92.5005
R4468 vdd.n167 vdd.n166 92.5005
R4469 vdd.n168 vdd.n167 92.5005
R4470 vdd.n14 vdd.n13 92.5005
R4471 vdd.n13 vdd.n12 92.5005
R4472 vdd.n10 vdd.n9 92.5005
R4473 vdd.n11 vdd.n10 92.5005
R4474 vdd.n157 vdd.n156 92.5005
R4475 vdd.n156 vdd.n155 92.5005
R4476 vdd.n112 vdd.n111 92.5005
R4477 vdd.n111 vdd.n110 92.5005
R4478 vdd.n108 vdd.n107 92.5005
R4479 vdd.n107 vdd.n106 92.5005
R4480 vdd.n104 vdd.n103 92.5005
R4481 vdd.n103 vdd.n102 92.5005
R4482 vdd.n91 vdd.n90 92.5005
R4483 vdd.n90 vdd.n89 92.5005
R4484 vdd.n87 vdd.n86 92.5005
R4485 vdd.n86 vdd.n85 92.5005
R4486 vdd.n75 vdd.t95 92.5005
R4487 vdd.n76 vdd.n75 92.5005
R4488 vdd.n73 vdd.n72 92.5005
R4489 vdd.n72 vdd.n71 92.5005
R4490 vdd.n62 vdd.n61 92.5005
R4491 vdd.n61 vdd.n60 92.5005
R4492 vdd.n58 vdd.n57 92.5005
R4493 vdd.n57 vdd.n56 92.5005
R4494 vdd.n136 vdd.n135 92.5005
R4495 vdd.n135 vdd.n134 92.5005
R4496 vdd.n132 vdd.n131 92.5005
R4497 vdd.n131 vdd.n130 92.5005
R4498 vdd.n153 vdd.n152 92.5005
R4499 vdd.n152 vdd.n151 92.5005
R4500 vdd.n42 vdd.n41 92.5005
R4501 vdd.n41 vdd.n40 92.5005
R4502 vdd.n46 vdd.n45 92.5005
R4503 vdd.n45 vdd.n44 92.5005
R4504 vdd.n52 vdd.n51 92.5005
R4505 vdd.n51 vdd.n50 92.5005
R4506 vdd.n23 vdd.n22 92.5005
R4507 vdd.n28 vdd.n27 92.5005
R4508 vdd.n27 vdd.n26 92.5005
R4509 vdd.n32 vdd.n31 92.5005
R4510 vdd.n31 vdd.n30 92.5005
R4511 vdd.n36 vdd.n35 92.5005
R4512 vdd.n35 vdd.n34 92.5005
R4513 vdd.n100 vdd.t34 91.4648
R4514 vdd.n100 vdd.t16 91.4648
R4515 vdd.n149 vdd.t36 91.4648
R4516 vdd.n4644 vdd 89.6591
R4517 vdd.n3946 vdd.n3944 88.3561
R4518 vdd.n2172 vdd.n2168 88.0097
R4519 vdd.n2193 vdd.t55 87.5415
R4520 vdd.n2193 vdd.t11 87.5415
R4521 vdd.n2181 vdd.t61 87.0498
R4522 vdd.n4526 vdd.n988 86.9025
R4523 vdd.n3920 vdd.n3919 86.9025
R4524 vdd.n54 vdd.t105 86.7743
R4525 vdd.n149 vdd.t107 86.7743
R4526 vdd.n5858 vdd.n5812 85.9427
R4527 vdd.n5812 vdd.n5802 85.9427
R4528 vdd.n6429 vdd.n212 85.9427
R4529 vdd.n6457 vdd.n212 85.9427
R4530 vdd.n6477 vdd.n212 85.9427
R4531 vdd.n6518 vdd.n212 85.9427
R4532 vdd.n6583 vdd.n212 85.9427
R4533 vdd.n6608 vdd.n212 85.9427
R4534 vdd.n6605 vdd.n212 85.9427
R4535 vdd.n6635 vdd.n212 85.9427
R4536 vdd.n6656 vdd.n212 85.9427
R4537 vdd.n6684 vdd.n212 85.9427
R4538 vdd.n6704 vdd.n212 85.9427
R4539 vdd.n6745 vdd.n212 85.9427
R4540 vdd.n6810 vdd.n212 85.9427
R4541 vdd.n6835 vdd.n212 85.9427
R4542 vdd.n6832 vdd.n212 85.9427
R4543 vdd.n6862 vdd.n212 85.9427
R4544 vdd.n6883 vdd.n212 85.9427
R4545 vdd.n6911 vdd.n212 85.9427
R4546 vdd.n6931 vdd.n212 85.9427
R4547 vdd.n6972 vdd.n212 85.9427
R4548 vdd.n7037 vdd.n212 85.9427
R4549 vdd.n7062 vdd.n212 85.9427
R4550 vdd.n7059 vdd.n212 85.9427
R4551 vdd.n7089 vdd.n212 85.9427
R4552 vdd.n7110 vdd.n212 85.9427
R4553 vdd.n7138 vdd.n212 85.9427
R4554 vdd.n7158 vdd.n212 85.9427
R4555 vdd.n7199 vdd.n212 85.9427
R4556 vdd.n7264 vdd.n212 85.9427
R4557 vdd.n3005 vdd.n2065 85.9427
R4558 vdd.n2721 vdd.n2065 85.9427
R4559 vdd.n3066 vdd.n2065 85.9427
R4560 vdd.n3091 vdd.n2065 85.9427
R4561 vdd.n3130 vdd.n2065 85.9427
R4562 vdd.n3233 vdd.n2065 85.9427
R4563 vdd.n2586 vdd.n2065 85.9427
R4564 vdd.n3294 vdd.n2065 85.9427
R4565 vdd.n3319 vdd.n2065 85.9427
R4566 vdd.n3358 vdd.n2065 85.9427
R4567 vdd.n3461 vdd.n2065 85.9427
R4568 vdd.n2451 vdd.n2065 85.9427
R4569 vdd.n3522 vdd.n2065 85.9427
R4570 vdd.n3547 vdd.n2065 85.9427
R4571 vdd.n3586 vdd.n2065 85.9427
R4572 vdd.n3688 vdd.n2065 85.9427
R4573 vdd.n3705 vdd.n2065 85.9427
R4574 vdd.n2295 vdd.n2065 85.9427
R4575 vdd.n3797 vdd.n2065 85.9427
R4576 vdd.n3639 vdd.n2065 85.9427
R4577 vdd.n3606 vdd.n2065 85.9427
R4578 vdd.n3411 vdd.n2065 85.9427
R4579 vdd.n3378 vdd.n2065 85.9427
R4580 vdd.n3183 vdd.n2065 85.9427
R4581 vdd.n3150 vdd.n2065 85.9427
R4582 vdd.n2955 vdd.n2065 85.9427
R4583 vdd.n2922 vdd.n2065 85.9427
R4584 vdd.n4025 vdd.n4024 85.9427
R4585 vdd.n4025 vdd.n2058 85.9427
R4586 vdd.n4025 vdd.n2060 85.9427
R4587 vdd.n4025 vdd.n2063 85.9427
R4588 vdd.n4779 vdd.n250 85.9427
R4589 vdd.n745 vdd.n250 85.9427
R4590 vdd.n4840 vdd.n250 85.9427
R4591 vdd.n4865 vdd.n250 85.9427
R4592 vdd.n4904 vdd.n250 85.9427
R4593 vdd.n5007 vdd.n250 85.9427
R4594 vdd.n610 vdd.n250 85.9427
R4595 vdd.n5068 vdd.n250 85.9427
R4596 vdd.n5093 vdd.n250 85.9427
R4597 vdd.n5132 vdd.n250 85.9427
R4598 vdd.n5235 vdd.n250 85.9427
R4599 vdd.n475 vdd.n250 85.9427
R4600 vdd.n5296 vdd.n250 85.9427
R4601 vdd.n5321 vdd.n250 85.9427
R4602 vdd.n5360 vdd.n250 85.9427
R4603 vdd.n5462 vdd.n250 85.9427
R4604 vdd.n5480 vdd.n250 85.9427
R4605 vdd.n321 vdd.n250 85.9427
R4606 vdd.n5573 vdd.n250 85.9427
R4607 vdd.n5413 vdd.n250 85.9427
R4608 vdd.n5380 vdd.n250 85.9427
R4609 vdd.n5185 vdd.n250 85.9427
R4610 vdd.n5152 vdd.n250 85.9427
R4611 vdd.n4957 vdd.n250 85.9427
R4612 vdd.n4924 vdd.n250 85.9427
R4613 vdd.n4729 vdd.n250 85.9427
R4614 vdd.n4696 vdd.n250 85.9427
R4615 vdd.n5727 vdd.n259 85.9427
R4616 vdd.n5728 vdd.n5727 85.9427
R4617 vdd.n1265 vdd 85.8969
R4618 vdd.n1529 vdd 85.8969
R4619 vdd.n1793 vdd 85.8969
R4620 vdd vdd.n3921 85.8969
R4621 vdd.n3976 vdd.t108 85.2946
R4622 vdd.n3835 vdd.n3834 79.3561
R4623 vdd vdd.n4583 79.2895
R4624 vdd.n3946 vdd 73.5299
R4625 vdd.n3980 vdd.t130 72.5495
R4626 vdd.n849 vdd 72.4801
R4627 vdd.t42 vdd.n7508 71.9403
R4628 vdd vdd.t103 71.2138
R4629 vdd.n4006 vdd 71.1459
R4630 vdd.n6392 vdd.t31 70.3649
R4631 vdd.n4670 vdd.t72 70.3649
R4632 vdd.n2223 vdd.t57 70.3628
R4633 vdd.n3889 vdd.t101 70.3628
R4634 vdd.n7462 vdd.t110 69.629
R4635 vdd.n7422 vdd.t76 68.0287
R4636 vdd.n5731 vdd.t87 68.0287
R4637 vdd.n4010 vdd.t24 68.0287
R4638 vdd.n876 vdd.t40 68.0287
R4639 vdd.n1141 vdd.t63 67.9081
R4640 vdd.n1405 vdd.t94 67.9081
R4641 vdd.n1669 vdd.t124 67.9081
R4642 vdd.n1933 vdd.t62 67.9081
R4643 vdd.n6409 vdd.n6407 67.5405
R4644 vdd.n7290 vdd.n7289 67.5405
R4645 vdd.n7177 vdd.n5938 67.3307
R4646 vdd.n6950 vdd.n6071 67.3307
R4647 vdd.n6723 vdd.n6204 67.3307
R4648 vdd.n6496 vdd.n6337 67.3307
R4649 vdd.n7399 vdd.n7398 67.3307
R4650 vdd.n6517 vdd.n6516 67.3307
R4651 vdd.n6554 vdd.n6553 67.3307
R4652 vdd.n6604 vdd.n6603 67.3307
R4653 vdd.n6744 vdd.n6743 67.3307
R4654 vdd.n6781 vdd.n6780 67.3307
R4655 vdd.n6831 vdd.n6830 67.3307
R4656 vdd.n6971 vdd.n6970 67.3307
R4657 vdd.n7008 vdd.n7007 67.3307
R4658 vdd.n7058 vdd.n7057 67.3307
R4659 vdd.n7198 vdd.n7197 67.3307
R4660 vdd.n7235 vdd.n7234 67.3307
R4661 vdd.n5669 vdd.n255 67.3307
R4662 vdd.n5505 vdd.n5504 67.3307
R4663 vdd.n5540 vdd.n5539 67.3307
R4664 vdd.n5267 vdd.n5266 67.3307
R4665 vdd.n5319 vdd.n5318 67.3307
R4666 vdd.n5039 vdd.n5038 67.3307
R4667 vdd.n5091 vdd.n5090 67.3307
R4668 vdd.n4811 vdd.n4810 67.3307
R4669 vdd.n4863 vdd.n4862 67.3307
R4670 vdd.n3729 vdd.n3728 67.3307
R4671 vdd.n3764 vdd.n3763 67.3307
R4672 vdd.n3493 vdd.n3492 67.3307
R4673 vdd.n3545 vdd.n3544 67.3307
R4674 vdd.n3265 vdd.n3264 67.3307
R4675 vdd.n3317 vdd.n3316 67.3307
R4676 vdd.n3037 vdd.n3036 67.3307
R4677 vdd.n3089 vdd.n3088 67.3307
R4678 vdd.n3667 vdd.n3666 67.3307
R4679 vdd.n3608 vdd.n2356 67.3307
R4680 vdd.n3439 vdd.n3438 67.3307
R4681 vdd.n3380 vdd.n2491 67.3307
R4682 vdd.n3211 vdd.n3210 67.3307
R4683 vdd.n3152 vdd.n2626 67.3307
R4684 vdd.n2983 vdd.n2982 67.3307
R4685 vdd.n2924 vdd.n2761 67.3307
R4686 vdd.n4026 vdd.n2057 67.3307
R4687 vdd.n2872 vdd.n2061 67.3307
R4688 vdd.n5441 vdd.n5440 67.3307
R4689 vdd.n5382 vdd.n380 67.3307
R4690 vdd.n5213 vdd.n5212 67.3307
R4691 vdd.n5154 vdd.n515 67.3307
R4692 vdd.n4985 vdd.n4984 67.3307
R4693 vdd.n4926 vdd.n650 67.3307
R4694 vdd.n4757 vdd.n4756 67.3307
R4695 vdd.n4698 vdd.n785 67.3307
R4696 vdd.t67 vdd 67.1434
R4697 vdd.n2178 vdd.n2177 67.0123
R4698 vdd.t25 vdd.t100 65.1272
R4699 vdd.n3835 vdd.n2068 64.8683
R4700 vdd.n169 vdd.t5 64.2862
R4701 vdd.n38 vdd.t8 63.1021
R4702 vdd vdd.n4004 62.7456
R4703 vdd.n2192 vdd.n2190 61.7439
R4704 vdd.n2192 vdd.n2191 61.7439
R4705 vdd.n174 vdd.t70 61.4291
R4706 vdd.n7509 vdd 61.1001
R4707 vdd vdd.n7482 59.137
R4708 vdd.n4005 vdd 58.824
R4709 vdd.t83 vdd.t67 58.5719
R4710 vdd.n24 vdd.t18 58.4849
R4711 vdd.n2173 vdd.n2169 57.9274
R4712 vdd.n60 vdd.t104 57.1434
R4713 vdd.t100 vdd 55.7965
R4714 vdd.n12 vdd.t96 55.7148
R4715 vdd.n2170 vdd.t0 55.1586
R4716 vdd.n106 vdd.t73 54.2862
R4717 vdd.n40 vdd.t13 52.8576
R4718 vdd.n159 vdd.t98 51.4291
R4719 vdd.n7464 vdd.n7461 48.6451
R4720 vdd.n102 vdd.t33 48.5719
R4721 vdd.t122 vdd.t44 48.3856
R4722 vdd.t79 vdd.t30 47.6077
R4723 vdd.t89 vdd.t71 47.6077
R4724 vdd.n2125 vdd.t48 47.1434
R4725 vdd.n2125 vdd.t47 47.1434
R4726 vdd.n3896 vdd.t27 47.1434
R4727 vdd.n3896 vdd.t21 47.1434
R4728 vdd.n833 vdd.t38 47.1434
R4729 vdd.n833 vdd.t41 47.1434
R4730 vdd.n5768 vdd.t92 47.1434
R4731 vdd.n5768 vdd.t91 47.1434
R4732 vdd.n4576 vdd.n4575 46.2524
R4733 vdd.n931 vdd.n856 46.2524
R4734 vdd.n943 vdd.n926 46.2524
R4735 vdd.n4549 vdd.n4548 46.2524
R4736 vdd.n995 vdd.n945 46.2524
R4737 vdd.n4524 vdd.n4523 46.2524
R4738 vdd.n1058 vdd.n1004 46.2524
R4739 vdd.n1070 vdd.n1053 46.2524
R4740 vdd.n4497 vdd.n4496 46.2524
R4741 vdd.n1123 vdd.n1072 46.2524
R4742 vdd.n4470 vdd.n1142 46.2524
R4743 vdd.n4450 vdd.n1183 46.2524
R4744 vdd.n4448 vdd.n1184 46.2524
R4745 vdd.n4428 vdd.n1225 46.2524
R4746 vdd.n4426 vdd.n1226 46.2524
R4747 vdd.n4403 vdd.n4402 46.2524
R4748 vdd.n1322 vdd.n1272 46.2524
R4749 vdd.n1334 vdd.n1317 46.2524
R4750 vdd.n4376 vdd.n4375 46.2524
R4751 vdd.n1387 vdd.n1336 46.2524
R4752 vdd.n4349 vdd.n1406 46.2524
R4753 vdd.n4329 vdd.n1447 46.2524
R4754 vdd.n4327 vdd.n1448 46.2524
R4755 vdd.n4307 vdd.n1489 46.2524
R4756 vdd.n4305 vdd.n1490 46.2524
R4757 vdd.n4282 vdd.n4281 46.2524
R4758 vdd.n1586 vdd.n1536 46.2524
R4759 vdd.n1598 vdd.n1581 46.2524
R4760 vdd.n4255 vdd.n4254 46.2524
R4761 vdd.n1651 vdd.n1600 46.2524
R4762 vdd.n4228 vdd.n1670 46.2524
R4763 vdd.n4208 vdd.n1711 46.2524
R4764 vdd.n4206 vdd.n1712 46.2524
R4765 vdd.n4186 vdd.n1753 46.2524
R4766 vdd.n4184 vdd.n1754 46.2524
R4767 vdd.n4161 vdd.n4160 46.2524
R4768 vdd.n1850 vdd.n1800 46.2524
R4769 vdd.n1862 vdd.n1845 46.2524
R4770 vdd.n4134 vdd.n4133 46.2524
R4771 vdd.n1915 vdd.n1864 46.2524
R4772 vdd.n4107 vdd.n1934 46.2524
R4773 vdd.n4087 vdd.n1975 46.2524
R4774 vdd.n4085 vdd.n1976 46.2524
R4775 vdd.n4065 vdd.n2017 46.2524
R4776 vdd.n4063 vdd.n2018 46.2524
R4777 vdd vdd.n2171 46.0253
R4778 vdd.n44 vdd.t7 45.7148
R4779 vdd.t37 vdd 44.7841
R4780 vdd.n7509 vdd.t42 43.3615
R4781 vdd.n3945 vdd.t130 43.1378
R4782 vdd.n7482 vdd.t110 41.9684
R4783 vdd.n1270 vdd 41.8475
R4784 vdd.n1534 vdd 41.8475
R4785 vdd.n1798 vdd 41.8475
R4786 vdd.n15 vdd.t97 41.5552
R4787 vdd.n15 vdd.t68 41.5552
R4788 vdd.n7484 vdd.t65 41.3905
R4789 vdd.n4004 vdd.t108 41.177
R4790 vdd.n4643 vdd.t117 40.0607
R4791 vdd.n7483 vdd 39.1069
R4792 vdd.n7506 vdd.n193 39.0005
R4793 vdd.n227 vdd.n214 39.0005
R4794 vdd.n54 vdd.t116 38.6969
R4795 vdd.n151 vdd.t106 38.5719
R4796 vdd.n3944 vdd.n3943 37.3561
R4797 vdd.t117 vdd.n228 36.2455
R4798 vdd.n3981 vdd.n3868 36.0005
R4799 vdd.n4623 vdd.n848 36.0005
R4800 vdd.n2214 vdd.n2213 34.6358
R4801 vdd.n6607 vdd.n6606 33.746
R4802 vdd.n6834 vdd.n6833 33.746
R4803 vdd.n7061 vdd.n7060 33.746
R4804 vdd.n3129 vdd.n3128 33.746
R4805 vdd.n3357 vdd.n3356 33.746
R4806 vdd.n3585 vdd.n3584 33.746
R4807 vdd.n1268 vdd.n1267 33.746
R4808 vdd.n1532 vdd.n1531 33.746
R4809 vdd.n1796 vdd.n1795 33.746
R4810 vdd.n4903 vdd.n4902 33.746
R4811 vdd.n5131 vdd.n5130 33.746
R4812 vdd.n5359 vdd.n5358 33.746
R4813 vdd.n6335 vdd.n6328 32.9702
R4814 vdd.n6202 vdd.n6195 32.9702
R4815 vdd.n6069 vdd.n6062 32.9702
R4816 vdd.n5936 vdd.n5929 32.9702
R4817 vdd.n2732 vdd.n2716 32.9702
R4818 vdd.n2597 vdd.n2581 32.9702
R4819 vdd.n2462 vdd.n2446 32.9702
R4820 vdd.n2327 vdd.n2320 32.9702
R4821 vdd.n1130 vdd.n1127 32.9702
R4822 vdd.n1394 vdd.n1391 32.9702
R4823 vdd.n1658 vdd.n1655 32.9702
R4824 vdd.n1922 vdd.n1919 32.9702
R4825 vdd.n756 vdd.n740 32.9702
R4826 vdd.n621 vdd.n605 32.9702
R4827 vdd.n486 vdd.n470 32.9702
R4828 vdd.n351 vdd.n344 32.9702
R4829 vdd.n2193 vdd.n2192 32.3373
R4830 vdd.n24 vdd.t59 31.831
R4831 vdd.n4622 vdd.n4621 31.0632
R4832 vdd.n7484 vdd 29.5648
R4833 vdd.n7424 vdd.n7423 29.4128
R4834 vdd.n5730 vdd.n247 29.4128
R4835 vdd.n4008 vdd.n4007 29.2586
R4836 vdd.n4583 vdd.n850 29.2586
R4837 vdd.t103 vdd.n1001 28.6326
R4838 vdd.t63 vdd.n1140 28.6326
R4839 vdd.n4472 vdd.t74 28.6326
R4840 vdd.t94 vdd.n1404 28.6326
R4841 vdd.n4351 vdd.t125 28.6326
R4842 vdd.t124 vdd.n1668 28.6326
R4843 vdd.n4230 vdd.t112 28.6326
R4844 vdd.t62 vdd.n1932 28.6326
R4845 vdd.n4109 vdd.t2 28.6326
R4846 vdd vdd.n4643 28.615
R4847 vdd.n7197 vdd.n7196 28.2358
R4848 vdd.n7235 vdd.n7233 28.2358
R4849 vdd.n7289 vdd.n5869 28.2358
R4850 vdd.n7178 vdd.n7177 28.2358
R4851 vdd.n6970 vdd.n6969 28.2358
R4852 vdd.n7008 vdd.n7006 28.2358
R4853 vdd.n7057 vdd.n6003 28.2358
R4854 vdd.n6951 vdd.n6950 28.2358
R4855 vdd.n6743 vdd.n6742 28.2358
R4856 vdd.n6781 vdd.n6779 28.2358
R4857 vdd.n6830 vdd.n6136 28.2358
R4858 vdd.n6724 vdd.n6723 28.2358
R4859 vdd.n6516 vdd.n6515 28.2358
R4860 vdd.n6554 vdd.n6552 28.2358
R4861 vdd.n6603 vdd.n6269 28.2358
R4862 vdd.n6409 vdd.n6408 28.2358
R4863 vdd.n6497 vdd.n6496 28.2358
R4864 vdd.n7337 vdd.n5847 28.2358
R4865 vdd.n7356 vdd.n5836 28.2358
R4866 vdd.n7375 vdd.n5825 28.2358
R4867 vdd.n7398 vdd.n5813 28.2358
R4868 vdd.n264 vdd.n251 28.2358
R4869 vdd.n5620 vdd.n257 28.2358
R4870 vdd.n5697 vdd.n253 28.2358
R4871 vdd.n5669 vdd.n5668 28.2358
R4872 vdd.n5504 vdd.n5503 28.2358
R4873 vdd.n5540 vdd.n5538 28.2358
R4874 vdd.n5410 vdd.n380 28.2358
R4875 vdd.n5443 vdd.n5441 28.2358
R4876 vdd.n5267 vdd.n5265 28.2358
R4877 vdd.n5318 vdd.n421 28.2358
R4878 vdd.n5357 vdd.n5356 28.2358
R4879 vdd.n5182 vdd.n515 28.2358
R4880 vdd.n5215 vdd.n5213 28.2358
R4881 vdd.n5039 vdd.n5037 28.2358
R4882 vdd.n5090 vdd.n556 28.2358
R4883 vdd.n5129 vdd.n5128 28.2358
R4884 vdd.n4954 vdd.n650 28.2358
R4885 vdd.n4987 vdd.n4985 28.2358
R4886 vdd.n4811 vdd.n4809 28.2358
R4887 vdd.n4862 vdd.n691 28.2358
R4888 vdd.n4901 vdd.n4900 28.2358
R4889 vdd.n4726 vdd.n785 28.2358
R4890 vdd.n4759 vdd.n4757 28.2358
R4891 vdd.n4581 vdd.n852 28.2358
R4892 vdd.n4573 vdd.n855 28.2358
R4893 vdd.n933 vdd.n930 28.2358
R4894 vdd.n942 vdd.n924 28.2358
R4895 vdd.n4546 vdd.n925 28.2358
R4896 vdd.n996 vdd.n993 28.2358
R4897 vdd.n4106 vdd.n1911 28.2358
R4898 vdd.n1973 vdd.n1961 28.2358
R4899 vdd.n4084 vdd.n1962 28.2358
R4900 vdd.n2015 vdd.n2003 28.2358
R4901 vdd.n4062 vdd.n2004 28.2358
R4902 vdd.n1797 vdd.n1787 28.2358
R4903 vdd.n4158 vdd.n1788 28.2358
R4904 vdd.n1852 vdd.n1849 28.2358
R4905 vdd.n1861 vdd.n1843 28.2358
R4906 vdd.n4131 vdd.n1844 28.2358
R4907 vdd.n1916 vdd.n1913 28.2358
R4908 vdd.n4227 vdd.n1647 28.2358
R4909 vdd.n1709 vdd.n1697 28.2358
R4910 vdd.n4205 vdd.n1698 28.2358
R4911 vdd.n1751 vdd.n1739 28.2358
R4912 vdd.n4183 vdd.n1740 28.2358
R4913 vdd.n1794 vdd.n1791 28.2358
R4914 vdd.n1533 vdd.n1523 28.2358
R4915 vdd.n4279 vdd.n1524 28.2358
R4916 vdd.n1588 vdd.n1585 28.2358
R4917 vdd.n1597 vdd.n1579 28.2358
R4918 vdd.n4252 vdd.n1580 28.2358
R4919 vdd.n1652 vdd.n1649 28.2358
R4920 vdd.n4348 vdd.n1383 28.2358
R4921 vdd.n1445 vdd.n1433 28.2358
R4922 vdd.n4326 vdd.n1434 28.2358
R4923 vdd.n1487 vdd.n1475 28.2358
R4924 vdd.n4304 vdd.n1476 28.2358
R4925 vdd.n1530 vdd.n1527 28.2358
R4926 vdd.n1269 vdd.n1259 28.2358
R4927 vdd.n4400 vdd.n1260 28.2358
R4928 vdd.n1324 vdd.n1321 28.2358
R4929 vdd.n1333 vdd.n1315 28.2358
R4930 vdd.n4373 vdd.n1316 28.2358
R4931 vdd.n1388 vdd.n1385 28.2358
R4932 vdd.n4469 vdd.n1119 28.2358
R4933 vdd.n1181 vdd.n1169 28.2358
R4934 vdd.n4447 vdd.n1170 28.2358
R4935 vdd.n1223 vdd.n1211 28.2358
R4936 vdd.n4425 vdd.n1212 28.2358
R4937 vdd.n1266 vdd.n1263 28.2358
R4938 vdd.n4521 vdd.n991 28.2358
R4939 vdd.n1060 vdd.n1057 28.2358
R4940 vdd.n1069 vdd.n1051 28.2358
R4941 vdd.n4494 vdd.n1052 28.2358
R4942 vdd.n1124 vdd.n1121 28.2358
R4943 vdd.n2806 vdd.n2057 28.2358
R4944 vdd.n2873 vdd.n2872 28.2358
R4945 vdd.n3728 vdd.n3727 28.2358
R4946 vdd.n3764 vdd.n3762 28.2358
R4947 vdd.n3636 vdd.n2356 28.2358
R4948 vdd.n3669 vdd.n3667 28.2358
R4949 vdd.n3493 vdd.n3491 28.2358
R4950 vdd.n3544 vdd.n2397 28.2358
R4951 vdd.n3583 vdd.n3582 28.2358
R4952 vdd.n3408 vdd.n2491 28.2358
R4953 vdd.n3441 vdd.n3439 28.2358
R4954 vdd.n3265 vdd.n3263 28.2358
R4955 vdd.n3316 vdd.n2532 28.2358
R4956 vdd.n3355 vdd.n3354 28.2358
R4957 vdd.n3180 vdd.n2626 28.2358
R4958 vdd.n3213 vdd.n3211 28.2358
R4959 vdd.n3037 vdd.n3035 28.2358
R4960 vdd.n3088 vdd.n2667 28.2358
R4961 vdd.n3127 vdd.n3126 28.2358
R4962 vdd.n2952 vdd.n2761 28.2358
R4963 vdd.n2985 vdd.n2983 28.2358
R4964 vdd.n38 vdd.t14 28.0332
R4965 vdd vdd.n3945 27.4515
R4966 vdd.n7489 vdd.n7488 27.3454
R4967 vdd.n5755 vdd.n5754 27.3454
R4968 vdd.n3858 vdd.n3838 27.1422
R4969 vdd.n4611 vdd.n4607 27.1422
R4970 vdd.n2191 vdd.t10 25.7981
R4971 vdd.n2191 vdd.t12 25.7981
R4972 vdd.n2190 vdd.t54 25.7981
R4973 vdd.n2190 vdd.t53 25.7981
R4974 vdd.n110 vdd.t113 25.7148
R4975 vdd.n89 vdd.t15 25.7148
R4976 vdd.n3923 vdd.n3922 25.696
R4977 vdd.n2175 vdd.n2169 24.2862
R4978 vdd.n2213 vdd.n2212 23.7181
R4979 vdd.n2212 vdd.n2211 23.3417
R4980 vdd.n3983 vdd.n3982 23.0907
R4981 vdd.n4625 vdd.n4624 23.0907
R4982 vdd.n7504 vdd.n192 22.8875
R4983 vdd.n224 vdd.n215 22.8875
R4984 vdd.n169 vdd 22.8576
R4985 vdd.n11 vdd 22.8576
R4986 vdd.t19 vdd.t28 22.6547
R4987 vdd.t28 vdd.t26 22.6547
R4988 vdd.t29 vdd.t23 22.6547
R4989 vdd.t30 vdd.t32 21.1252
R4990 vdd.t71 vdd.t39 21.1252
R4991 vdd.n7461 vdd.n7460 20.7428
R4992 vdd.n7461 vdd.n229 20.7428
R4993 vdd.n5743 vdd.n228 20.7428
R4994 vdd.n7437 vdd.n7436 20.7428
R4995 vdd.n7444 vdd.n5777 20.7428
R4996 vdd.n5783 vdd.n213 20.7428
R4997 vdd.n7426 vdd.n7425 20.7428
R4998 vdd.n5811 vdd.n5810 20.7428
R4999 vdd.n3808 vdd.n2068 20.7428
R5000 vdd.n3820 vdd.n3819 20.7428
R5001 vdd.n3821 vdd.n2080 20.7428
R5002 vdd.n3823 vdd.n3822 20.7428
R5003 vdd.n2243 vdd.n2079 20.7428
R5004 vdd.n3834 vdd.n3833 20.7428
R5005 vdd.n2232 vdd.n2069 20.7428
R5006 vdd.n3976 vdd.n3975 20.7428
R5007 vdd.n3976 vdd.n3948 20.7428
R5008 vdd.n3976 vdd.n3947 20.7428
R5009 vdd.n3932 vdd.n3869 20.7428
R5010 vdd.n3943 vdd.n3942 20.7428
R5011 vdd.n3943 vdd.n3870 20.7428
R5012 vdd.n3884 vdd.n3869 20.7428
R5013 vdd.n3924 vdd.n3923 20.7428
R5014 vdd.n827 vdd.n826 20.7428
R5015 vdd.n4642 vdd.n4641 20.7428
R5016 vdd.n4656 vdd.n4654 20.7428
R5017 vdd.n4653 vdd.n4651 20.7428
R5018 vdd.n4664 vdd.n812 20.7428
R5019 vdd.n2207 vdd.n2206 20.7064
R5020 vdd.n2178 vdd.t123 20.406
R5021 vdd.t74 vdd.n1141 20.3031
R5022 vdd.t125 vdd.n1405 20.3031
R5023 vdd.t112 vdd.n1669 20.3031
R5024 vdd.t2 vdd.n1933 20.3031
R5025 vdd.n2170 vdd.t19 19.0432
R5026 vdd.n130 vdd.t35 18.5719
R5027 vdd.n7425 vdd.t80 18.5229
R5028 vdd.t90 vdd.n827 18.5229
R5029 vdd.n7415 vdd 16.8265
R5030 vdd.n3821 vdd.n3820 16.7406
R5031 vdd vdd.t82 16.5329
R5032 vdd vdd.t85 16.5329
R5033 vdd.n2181 vdd.n2180 15.6903
R5034 vdd.n3854 vdd 15.4887
R5035 vdd.n844 vdd 15.4887
R5036 vdd.n7513 vdd.n7512 15.4666
R5037 vdd.n7479 vdd.n7478 15.4666
R5038 vdd.n211 vdd 15.1421
R5039 vdd.n5752 vdd 15.1421
R5040 vdd.n4001 vdd.n4000 15.12
R5041 vdd.n4609 vdd.n4608 15.12
R5042 vdd.n3868 vdd.n3837 15.0005
R5043 vdd.n4619 vdd.n848 15.0005
R5044 vdd.n2194 vdd.n2193 14.0645
R5045 vdd.n4010 vdd.n4008 13.7917
R5046 vdd.n876 vdd.n850 13.7917
R5047 vdd.t22 vdd.n4005 13.4617
R5048 vdd.n7423 vdd.n7422 13.3673
R5049 vdd.n5731 vdd.n5730 13.3673
R5050 vdd.n7200 vdd.n7199 13.1177
R5051 vdd.n7264 vdd.n7263 13.1177
R5052 vdd.n7089 vdd.n5975 13.1177
R5053 vdd.n7110 vdd.n5960 13.1177
R5054 vdd.n7139 vdd.n7138 13.1177
R5055 vdd.n7159 vdd.n7158 13.1177
R5056 vdd.n6973 vdd.n6972 13.1177
R5057 vdd.n7037 vdd.n7036 13.1177
R5058 vdd.n7063 vdd.n7062 13.1177
R5059 vdd.n6862 vdd.n6108 13.1177
R5060 vdd.n6883 vdd.n6093 13.1177
R5061 vdd.n6912 vdd.n6911 13.1177
R5062 vdd.n6932 vdd.n6931 13.1177
R5063 vdd.n6746 vdd.n6745 13.1177
R5064 vdd.n6810 vdd.n6809 13.1177
R5065 vdd.n6836 vdd.n6835 13.1177
R5066 vdd.n6635 vdd.n6241 13.1177
R5067 vdd.n6656 vdd.n6226 13.1177
R5068 vdd.n6685 vdd.n6684 13.1177
R5069 vdd.n6705 vdd.n6704 13.1177
R5070 vdd.n6519 vdd.n6518 13.1177
R5071 vdd.n6583 vdd.n6582 13.1177
R5072 vdd.n6609 vdd.n6608 13.1177
R5073 vdd.n6429 vdd.n6359 13.1177
R5074 vdd.n6458 vdd.n6457 13.1177
R5075 vdd.n6478 vdd.n6477 13.1177
R5076 vdd.n7318 vdd.n5858 13.1177
R5077 vdd.n5802 vdd.n5801 13.1177
R5078 vdd.n7299 vdd.n5858 13.1177
R5079 vdd.n6518 vdd.n6299 13.1177
R5080 vdd.n6584 vdd.n6583 13.1177
R5081 vdd.n6745 vdd.n6166 13.1177
R5082 vdd.n6811 vdd.n6810 13.1177
R5083 vdd.n6972 vdd.n6033 13.1177
R5084 vdd.n7038 vdd.n7037 13.1177
R5085 vdd.n7199 vdd.n5900 13.1177
R5086 vdd.n7265 vdd.n7264 13.1177
R5087 vdd.n7158 vdd.n7157 13.1177
R5088 vdd.n7138 vdd.n7137 13.1177
R5089 vdd.n7111 vdd.n7110 13.1177
R5090 vdd.n7090 vdd.n7089 13.1177
R5091 vdd.n7059 vdd.n5986 13.1177
R5092 vdd.n6931 vdd.n6930 13.1177
R5093 vdd.n6911 vdd.n6910 13.1177
R5094 vdd.n6884 vdd.n6883 13.1177
R5095 vdd.n6863 vdd.n6862 13.1177
R5096 vdd.n6832 vdd.n6119 13.1177
R5097 vdd.n6704 vdd.n6703 13.1177
R5098 vdd.n6684 vdd.n6683 13.1177
R5099 vdd.n6657 vdd.n6656 13.1177
R5100 vdd.n6636 vdd.n6635 13.1177
R5101 vdd.n6605 vdd.n6252 13.1177
R5102 vdd.n6477 vdd.n6476 13.1177
R5103 vdd.n6457 vdd.n6456 13.1177
R5104 vdd.n6430 vdd.n6429 13.1177
R5105 vdd.n5722 vdd.n259 13.1177
R5106 vdd.n5480 vdd.n324 13.1177
R5107 vdd.n322 vdd.n321 13.1177
R5108 vdd.n5573 vdd.n5572 13.1177
R5109 vdd.n5380 vdd.n5379 13.1177
R5110 vdd.n5414 vdd.n5413 13.1177
R5111 vdd.n5462 vdd.n5461 13.1177
R5112 vdd.n475 vdd.n455 13.1177
R5113 vdd.n5296 vdd.n5295 13.1177
R5114 vdd.n5322 vdd.n5321 13.1177
R5115 vdd.n5152 vdd.n5151 13.1177
R5116 vdd.n5186 vdd.n5185 13.1177
R5117 vdd.n5235 vdd.n5234 13.1177
R5118 vdd.n610 vdd.n590 13.1177
R5119 vdd.n5068 vdd.n5067 13.1177
R5120 vdd.n5094 vdd.n5093 13.1177
R5121 vdd.n4924 vdd.n4923 13.1177
R5122 vdd.n4958 vdd.n4957 13.1177
R5123 vdd.n5007 vdd.n5006 13.1177
R5124 vdd.n745 vdd.n725 13.1177
R5125 vdd.n4840 vdd.n4839 13.1177
R5126 vdd.n4866 vdd.n4865 13.1177
R5127 vdd.n4696 vdd.n4695 13.1177
R5128 vdd.n4730 vdd.n4729 13.1177
R5129 vdd.n4779 vdd.n4778 13.1177
R5130 vdd.n4014 vdd.n2058 13.1177
R5131 vdd.n2851 vdd.n2060 13.1177
R5132 vdd.n2881 vdd.n2063 13.1177
R5133 vdd.n3705 vdd.n2298 13.1177
R5134 vdd.n2296 vdd.n2295 13.1177
R5135 vdd.n3797 vdd.n3796 13.1177
R5136 vdd.n3606 vdd.n3605 13.1177
R5137 vdd.n3640 vdd.n3639 13.1177
R5138 vdd.n3688 vdd.n3687 13.1177
R5139 vdd.n2451 vdd.n2431 13.1177
R5140 vdd.n3522 vdd.n3521 13.1177
R5141 vdd.n3548 vdd.n3547 13.1177
R5142 vdd.n3378 vdd.n3377 13.1177
R5143 vdd.n3412 vdd.n3411 13.1177
R5144 vdd.n3461 vdd.n3460 13.1177
R5145 vdd.n2586 vdd.n2566 13.1177
R5146 vdd.n3294 vdd.n3293 13.1177
R5147 vdd.n3320 vdd.n3319 13.1177
R5148 vdd.n3150 vdd.n3149 13.1177
R5149 vdd.n3184 vdd.n3183 13.1177
R5150 vdd.n3233 vdd.n3232 13.1177
R5151 vdd.n2721 vdd.n2701 13.1177
R5152 vdd.n3066 vdd.n3065 13.1177
R5153 vdd.n3092 vdd.n3091 13.1177
R5154 vdd.n2922 vdd.n2921 13.1177
R5155 vdd.n2956 vdd.n2955 13.1177
R5156 vdd.n3005 vdd.n3004 13.1177
R5157 vdd.n2923 vdd.n2922 13.1177
R5158 vdd.n2955 vdd.n2745 13.1177
R5159 vdd.n3151 vdd.n3150 13.1177
R5160 vdd.n3183 vdd.n2610 13.1177
R5161 vdd.n3379 vdd.n3378 13.1177
R5162 vdd.n3411 vdd.n2475 13.1177
R5163 vdd.n3607 vdd.n3606 13.1177
R5164 vdd.n3639 vdd.n2340 13.1177
R5165 vdd.n3798 vdd.n3797 13.1177
R5166 vdd.n2295 vdd.n2278 13.1177
R5167 vdd.n3706 vdd.n3705 13.1177
R5168 vdd.n3689 vdd.n3688 13.1177
R5169 vdd.n3587 vdd.n3586 13.1177
R5170 vdd.n3547 vdd.n2380 13.1177
R5171 vdd.n3523 vdd.n3522 13.1177
R5172 vdd.n2452 vdd.n2451 13.1177
R5173 vdd.n3462 vdd.n3461 13.1177
R5174 vdd.n3359 vdd.n3358 13.1177
R5175 vdd.n3319 vdd.n2515 13.1177
R5176 vdd.n3295 vdd.n3294 13.1177
R5177 vdd.n2587 vdd.n2586 13.1177
R5178 vdd.n3234 vdd.n3233 13.1177
R5179 vdd.n3131 vdd.n3130 13.1177
R5180 vdd.n3091 vdd.n2650 13.1177
R5181 vdd.n3067 vdd.n3066 13.1177
R5182 vdd.n2722 vdd.n2721 13.1177
R5183 vdd.n3006 vdd.n3005 13.1177
R5184 vdd.n4024 vdd.n2067 13.1177
R5185 vdd.n2058 vdd.n2056 13.1177
R5186 vdd.n2854 vdd.n2060 13.1177
R5187 vdd.n2878 vdd.n2063 13.1177
R5188 vdd.n4697 vdd.n4696 13.1177
R5189 vdd.n4729 vdd.n769 13.1177
R5190 vdd.n4925 vdd.n4924 13.1177
R5191 vdd.n4957 vdd.n634 13.1177
R5192 vdd.n5153 vdd.n5152 13.1177
R5193 vdd.n5185 vdd.n499 13.1177
R5194 vdd.n5381 vdd.n5380 13.1177
R5195 vdd.n5413 vdd.n364 13.1177
R5196 vdd.n5574 vdd.n5573 13.1177
R5197 vdd.n321 vdd.n304 13.1177
R5198 vdd.n5481 vdd.n5480 13.1177
R5199 vdd.n5463 vdd.n5462 13.1177
R5200 vdd.n5361 vdd.n5360 13.1177
R5201 vdd.n5321 vdd.n404 13.1177
R5202 vdd.n5297 vdd.n5296 13.1177
R5203 vdd.n476 vdd.n475 13.1177
R5204 vdd.n5236 vdd.n5235 13.1177
R5205 vdd.n5133 vdd.n5132 13.1177
R5206 vdd.n5093 vdd.n539 13.1177
R5207 vdd.n5069 vdd.n5068 13.1177
R5208 vdd.n611 vdd.n610 13.1177
R5209 vdd.n5008 vdd.n5007 13.1177
R5210 vdd.n4905 vdd.n4904 13.1177
R5211 vdd.n4865 vdd.n674 13.1177
R5212 vdd.n4841 vdd.n4840 13.1177
R5213 vdd.n746 vdd.n745 13.1177
R5214 vdd.n4780 vdd.n4779 13.1177
R5215 vdd.n5728 vdd.n249 13.1177
R5216 vdd.n260 vdd.n259 13.1177
R5217 vdd.n3920 vdd.n3918 13.0163
R5218 vdd.n990 vdd.n988 13.0163
R5219 vdd.n4621 vdd.n4620 12.9433
R5220 vdd.n7508 vdd.n7507 12.8117
R5221 vdd.n7436 vdd.t81 12.5529
R5222 vdd.t93 vdd.n4653 12.5529
R5223 vdd.n4583 vdd.n4582 12.4812
R5224 vdd.n7463 vdd.n7462 12.4001
R5225 vdd.n4007 vdd.n4006 12.1484
R5226 vdd.n2182 vdd.n2181 12.0476
R5227 vdd.n7506 vdd.n195 12.0005
R5228 vdd.n7465 vdd.n227 12.0005
R5229 vdd.n7511 vdd.n192 11.9758
R5230 vdd.n3983 vdd.n3855 11.9758
R5231 vdd.n4625 vdd.n845 11.9758
R5232 vdd.n7480 vdd.n215 11.9758
R5233 vdd.n3980 vdd.n3979 11.7652
R5234 vdd.n4582 vdd.n851 11.747
R5235 vdd.n4575 vdd.n4574 11.747
R5236 vdd.n932 vdd.n931 11.747
R5237 vdd.n944 vdd.n943 11.747
R5238 vdd.n4548 vdd.n4547 11.747
R5239 vdd.n995 vdd.n992 11.747
R5240 vdd.n1003 vdd.n1002 11.747
R5241 vdd.n4523 vdd.n4522 11.747
R5242 vdd.n1059 vdd.n1058 11.747
R5243 vdd.n1071 vdd.n1070 11.747
R5244 vdd.n4496 vdd.n4495 11.747
R5245 vdd.n1123 vdd.n1120 11.747
R5246 vdd.n4471 vdd.n4470 11.747
R5247 vdd.n1183 vdd.n1182 11.747
R5248 vdd.n4449 vdd.n4448 11.747
R5249 vdd.n1225 vdd.n1224 11.747
R5250 vdd.n4427 vdd.n4426 11.747
R5251 vdd.n1265 vdd.n1264 11.747
R5252 vdd.n1271 vdd.n1270 11.747
R5253 vdd.n4402 vdd.n4401 11.747
R5254 vdd.n1323 vdd.n1322 11.747
R5255 vdd.n1335 vdd.n1334 11.747
R5256 vdd.n4375 vdd.n4374 11.747
R5257 vdd.n1387 vdd.n1384 11.747
R5258 vdd.n4350 vdd.n4349 11.747
R5259 vdd.n1447 vdd.n1446 11.747
R5260 vdd.n4328 vdd.n4327 11.747
R5261 vdd.n1489 vdd.n1488 11.747
R5262 vdd.n4306 vdd.n4305 11.747
R5263 vdd.n1529 vdd.n1528 11.747
R5264 vdd.n1535 vdd.n1534 11.747
R5265 vdd.n4281 vdd.n4280 11.747
R5266 vdd.n1587 vdd.n1586 11.747
R5267 vdd.n1599 vdd.n1598 11.747
R5268 vdd.n4254 vdd.n4253 11.747
R5269 vdd.n1651 vdd.n1648 11.747
R5270 vdd.n4229 vdd.n4228 11.747
R5271 vdd.n1711 vdd.n1710 11.747
R5272 vdd.n4207 vdd.n4206 11.747
R5273 vdd.n1753 vdd.n1752 11.747
R5274 vdd.n4185 vdd.n4184 11.747
R5275 vdd.n1793 vdd.n1792 11.747
R5276 vdd.n1799 vdd.n1798 11.747
R5277 vdd.n4160 vdd.n4159 11.747
R5278 vdd.n1851 vdd.n1850 11.747
R5279 vdd.n1863 vdd.n1862 11.747
R5280 vdd.n4133 vdd.n4132 11.747
R5281 vdd.n1915 vdd.n1912 11.747
R5282 vdd.n4108 vdd.n4107 11.747
R5283 vdd.n1975 vdd.n1974 11.747
R5284 vdd.n4086 vdd.n4085 11.747
R5285 vdd.n2017 vdd.n2016 11.747
R5286 vdd.n4064 vdd.n4063 11.747
R5287 vdd.n3921 vdd.n3917 11.747
R5288 vdd.n7291 vdd.n7290 11.5452
R5289 vdd.n6407 vdd.n6406 11.5452
R5290 vdd.t81 vdd.n5777 11.4813
R5291 vdd.n4654 vdd.t93 11.4813
R5292 vdd.n85 vdd.t69 11.4291
R5293 vdd vdd.n7415 11.3275
R5294 vdd.n7489 vdd.n7486 11.2229
R5295 vdd.n4002 vdd.n3838 11.2229
R5296 vdd.n4611 vdd.n4610 11.2229
R5297 vdd.n5754 vdd.n5753 11.2229
R5298 vdd.n2214 vdd.n2101 10.5417
R5299 vdd.n7461 vdd.n228 10.4925
R5300 vdd.n2079 vdd.n2068 10.4631
R5301 vdd.n2174 vdd.n2172 10.1637
R5302 vdd.n4006 vdd.t22 10.0143
R5303 vdd.n2194 vdd.n2183 9.75971
R5304 vdd.n5777 vdd.t78 9.64439
R5305 vdd.n4654 vdd.t88 9.64439
R5306 vdd.n7195 vdd.n7194 9.38471
R5307 vdd.n7180 vdd.n7179 9.38471
R5308 vdd.n6968 vdd.n6967 9.38471
R5309 vdd.n6953 vdd.n6952 9.38471
R5310 vdd.n6741 vdd.n6740 9.38471
R5311 vdd.n6726 vdd.n6725 9.38471
R5312 vdd.n6514 vdd.n6513 9.38471
R5313 vdd.n6499 vdd.n6498 9.38471
R5314 vdd.n7488 vdd.n7487 9.3005
R5315 vdd.n7503 vdd.n7502 9.3005
R5316 vdd.n7503 vdd.n195 9.3005
R5317 vdd.n195 vdd.n194 9.3005
R5318 vdd.n6335 vdd.n6334 9.3005
R5319 vdd.n6601 vdd.n6600 9.3005
R5320 vdd.n6557 vdd.n6556 9.3005
R5321 vdd.n6524 vdd.n6523 9.3005
R5322 vdd.n6329 vdd.n6328 9.3005
R5323 vdd.n6301 vdd.n6300 9.3005
R5324 vdd.n6286 vdd.n6285 9.3005
R5325 vdd.n6202 vdd.n6201 9.3005
R5326 vdd.n6828 vdd.n6827 9.3005
R5327 vdd.n6784 vdd.n6783 9.3005
R5328 vdd.n6751 vdd.n6750 9.3005
R5329 vdd.n6196 vdd.n6195 9.3005
R5330 vdd.n6168 vdd.n6167 9.3005
R5331 vdd.n6153 vdd.n6152 9.3005
R5332 vdd.n6069 vdd.n6068 9.3005
R5333 vdd.n7055 vdd.n7054 9.3005
R5334 vdd.n7011 vdd.n7010 9.3005
R5335 vdd.n6978 vdd.n6977 9.3005
R5336 vdd.n6063 vdd.n6062 9.3005
R5337 vdd.n6035 vdd.n6034 9.3005
R5338 vdd.n6020 vdd.n6019 9.3005
R5339 vdd.n5936 vdd.n5935 9.3005
R5340 vdd.n7287 vdd.n7286 9.3005
R5341 vdd.n7238 vdd.n7237 9.3005
R5342 vdd.n7205 vdd.n7204 9.3005
R5343 vdd.n5930 vdd.n5929 9.3005
R5344 vdd.n5902 vdd.n5901 9.3005
R5345 vdd.n5887 vdd.n5886 9.3005
R5346 vdd.n7175 vdd.n7174 9.3005
R5347 vdd.n7155 vdd.n7154 9.3005
R5348 vdd.n5966 vdd.n5965 9.3005
R5349 vdd.n7114 vdd.n7113 9.3005
R5350 vdd.n7093 vdd.n7092 9.3005
R5351 vdd.n6948 vdd.n6947 9.3005
R5352 vdd.n6928 vdd.n6927 9.3005
R5353 vdd.n6099 vdd.n6098 9.3005
R5354 vdd.n6887 vdd.n6886 9.3005
R5355 vdd.n6866 vdd.n6865 9.3005
R5356 vdd.n6721 vdd.n6720 9.3005
R5357 vdd.n6701 vdd.n6700 9.3005
R5358 vdd.n6232 vdd.n6231 9.3005
R5359 vdd.n6660 vdd.n6659 9.3005
R5360 vdd.n6639 vdd.n6638 9.3005
R5361 vdd.n6494 vdd.n6493 9.3005
R5362 vdd.n6474 vdd.n6473 9.3005
R5363 vdd.n6365 vdd.n6364 9.3005
R5364 vdd.n6412 vdd.n6411 9.3005
R5365 vdd.n6433 vdd.n6432 9.3005
R5366 vdd.n7316 vdd.n7315 9.3005
R5367 vdd.n7335 vdd.n7334 9.3005
R5368 vdd.n7354 vdd.n7353 9.3005
R5369 vdd.n7373 vdd.n7372 9.3005
R5370 vdd.n7396 vdd.n7395 9.3005
R5371 vdd.n7322 vdd.n7321 9.3005
R5372 vdd.n7321 vdd.n7320 9.3005
R5373 vdd.n7341 vdd.n7340 9.3005
R5374 vdd.n7340 vdd.n7339 9.3005
R5375 vdd.n7360 vdd.n7359 9.3005
R5376 vdd.n7359 vdd.n7358 9.3005
R5377 vdd.n7379 vdd.n7378 9.3005
R5378 vdd.n7378 vdd.n7377 9.3005
R5379 vdd.n7402 vdd.n7401 9.3005
R5380 vdd.n7401 vdd.n7400 9.3005
R5381 vdd.n7301 vdd.n7300 9.3005
R5382 vdd.n7300 vdd.n5812 9.3005
R5383 vdd.n6612 vdd.n6611 9.3005
R5384 vdd.n6611 vdd.n6610 9.3005
R5385 vdd.n6580 vdd.n6579 9.3005
R5386 vdd.n6580 vdd.n6281 9.3005
R5387 vdd.n6521 vdd.n6303 9.3005
R5388 vdd.n6521 vdd.n6520 9.3005
R5389 vdd.n6513 vdd.n6512 9.3005
R5390 vdd.n6549 vdd.n6297 9.3005
R5391 vdd.n6550 vdd.n6549 9.3005
R5392 vdd.n6588 vdd.n6587 9.3005
R5393 vdd.n6587 vdd.n6586 9.3005
R5394 vdd.n6839 vdd.n6838 9.3005
R5395 vdd.n6838 vdd.n6837 9.3005
R5396 vdd.n6807 vdd.n6806 9.3005
R5397 vdd.n6807 vdd.n6148 9.3005
R5398 vdd.n6748 vdd.n6170 9.3005
R5399 vdd.n6748 vdd.n6747 9.3005
R5400 vdd.n6740 vdd.n6739 9.3005
R5401 vdd.n6776 vdd.n6164 9.3005
R5402 vdd.n6777 vdd.n6776 9.3005
R5403 vdd.n6815 vdd.n6814 9.3005
R5404 vdd.n6814 vdd.n6813 9.3005
R5405 vdd.n7066 vdd.n7065 9.3005
R5406 vdd.n7065 vdd.n7064 9.3005
R5407 vdd.n7034 vdd.n7033 9.3005
R5408 vdd.n7034 vdd.n6015 9.3005
R5409 vdd.n6975 vdd.n6037 9.3005
R5410 vdd.n6975 vdd.n6974 9.3005
R5411 vdd.n6967 vdd.n6966 9.3005
R5412 vdd.n7003 vdd.n6031 9.3005
R5413 vdd.n7004 vdd.n7003 9.3005
R5414 vdd.n7042 vdd.n7041 9.3005
R5415 vdd.n7041 vdd.n7040 9.3005
R5416 vdd.n7261 vdd.n7260 9.3005
R5417 vdd.n7261 vdd.n5882 9.3005
R5418 vdd.n7202 vdd.n5904 9.3005
R5419 vdd.n7202 vdd.n7201 9.3005
R5420 vdd.n7194 vdd.n7193 9.3005
R5421 vdd.n7230 vdd.n5898 9.3005
R5422 vdd.n7231 vdd.n7230 9.3005
R5423 vdd.n7269 vdd.n7268 9.3005
R5424 vdd.n7268 vdd.n7267 9.3005
R5425 vdd.n7292 vdd.n7291 9.3005
R5426 vdd.n7162 vdd.n7161 9.3005
R5427 vdd.n7161 vdd.n7160 9.3005
R5428 vdd.n7142 vdd.n7141 9.3005
R5429 vdd.n7141 vdd.n5949 9.3005
R5430 vdd.n5949 vdd.n212 9.3005
R5431 vdd.n7135 vdd.n7134 9.3005
R5432 vdd.n7136 vdd.n7135 9.3005
R5433 vdd.n7136 vdd.n212 9.3005
R5434 vdd.n7108 vdd.n7107 9.3005
R5435 vdd.n7109 vdd.n7108 9.3005
R5436 vdd.n7109 vdd.n212 9.3005
R5437 vdd.n7181 vdd.n7180 9.3005
R5438 vdd.n7087 vdd.n7086 9.3005
R5439 vdd.n7088 vdd.n7087 9.3005
R5440 vdd.n7088 vdd.n212 9.3005
R5441 vdd.n6935 vdd.n6934 9.3005
R5442 vdd.n6934 vdd.n6933 9.3005
R5443 vdd.n6915 vdd.n6914 9.3005
R5444 vdd.n6914 vdd.n6082 9.3005
R5445 vdd.n6082 vdd.n212 9.3005
R5446 vdd.n6908 vdd.n6907 9.3005
R5447 vdd.n6909 vdd.n6908 9.3005
R5448 vdd.n6909 vdd.n212 9.3005
R5449 vdd.n6881 vdd.n6880 9.3005
R5450 vdd.n6882 vdd.n6881 9.3005
R5451 vdd.n6882 vdd.n212 9.3005
R5452 vdd.n6954 vdd.n6953 9.3005
R5453 vdd.n6860 vdd.n6859 9.3005
R5454 vdd.n6861 vdd.n6860 9.3005
R5455 vdd.n6861 vdd.n212 9.3005
R5456 vdd.n6708 vdd.n6707 9.3005
R5457 vdd.n6707 vdd.n6706 9.3005
R5458 vdd.n6688 vdd.n6687 9.3005
R5459 vdd.n6687 vdd.n6215 9.3005
R5460 vdd.n6215 vdd.n212 9.3005
R5461 vdd.n6681 vdd.n6680 9.3005
R5462 vdd.n6682 vdd.n6681 9.3005
R5463 vdd.n6682 vdd.n212 9.3005
R5464 vdd.n6654 vdd.n6653 9.3005
R5465 vdd.n6655 vdd.n6654 9.3005
R5466 vdd.n6655 vdd.n212 9.3005
R5467 vdd.n6727 vdd.n6726 9.3005
R5468 vdd.n6633 vdd.n6632 9.3005
R5469 vdd.n6634 vdd.n6633 9.3005
R5470 vdd.n6634 vdd.n212 9.3005
R5471 vdd.n6481 vdd.n6480 9.3005
R5472 vdd.n6480 vdd.n6479 9.3005
R5473 vdd.n6461 vdd.n6460 9.3005
R5474 vdd.n6460 vdd.n6348 9.3005
R5475 vdd.n6348 vdd.n212 9.3005
R5476 vdd.n6454 vdd.n6453 9.3005
R5477 vdd.n6455 vdd.n6454 9.3005
R5478 vdd.n6455 vdd.n212 9.3005
R5479 vdd.n6500 vdd.n6499 9.3005
R5480 vdd.n6406 vdd.n6405 9.3005
R5481 vdd.n6427 vdd.n6426 9.3005
R5482 vdd.n6428 vdd.n6427 9.3005
R5483 vdd.n5677 vdd.n5676 9.3005
R5484 vdd.n5695 vdd.n5694 9.3005
R5485 vdd.n5623 vdd.n5609 9.3005
R5486 vdd.n5587 vdd.n262 9.3005
R5487 vdd.n5614 vdd.n5613 9.3005
R5488 vdd.n2211 vdd.n2210 9.3005
R5489 vdd.n2732 vdd.n2731 9.3005
R5490 vdd.n2718 vdd.n2716 9.3005
R5491 vdd.n3096 vdd.n3095 9.3005
R5492 vdd.n2597 vdd.n2596 9.3005
R5493 vdd.n2583 vdd.n2581 9.3005
R5494 vdd.n3324 vdd.n3323 9.3005
R5495 vdd.n2462 vdd.n2461 9.3005
R5496 vdd.n2448 vdd.n2446 9.3005
R5497 vdd.n3552 vdd.n3551 9.3005
R5498 vdd.n2327 vdd.n2326 9.3005
R5499 vdd.n2321 vdd.n2320 9.3005
R5500 vdd.n2263 vdd.n2262 9.3005
R5501 vdd.n3767 vdd.n3766 9.3005
R5502 vdd.n2280 vdd.n2279 9.3005
R5503 vdd.n3734 vdd.n3733 9.3005
R5504 vdd.n3710 vdd.n3709 9.3005
R5505 vdd.n3685 vdd.n3684 9.3005
R5506 vdd.n2346 vdd.n2345 9.3005
R5507 vdd.n3643 vdd.n3642 9.3005
R5508 vdd.n3633 vdd.n3632 9.3005
R5509 vdd.n3603 vdd.n3602 9.3005
R5510 vdd.n3542 vdd.n3541 9.3005
R5511 vdd.n2418 vdd.n2417 9.3005
R5512 vdd.n3496 vdd.n3495 9.3005
R5513 vdd.n2433 vdd.n2432 9.3005
R5514 vdd.n3458 vdd.n3457 9.3005
R5515 vdd.n2481 vdd.n2480 9.3005
R5516 vdd.n3415 vdd.n3414 9.3005
R5517 vdd.n3405 vdd.n3404 9.3005
R5518 vdd.n3375 vdd.n3374 9.3005
R5519 vdd.n3314 vdd.n3313 9.3005
R5520 vdd.n2553 vdd.n2552 9.3005
R5521 vdd.n3268 vdd.n3267 9.3005
R5522 vdd.n2568 vdd.n2567 9.3005
R5523 vdd.n3230 vdd.n3229 9.3005
R5524 vdd.n2616 vdd.n2615 9.3005
R5525 vdd.n3187 vdd.n3186 9.3005
R5526 vdd.n3177 vdd.n3176 9.3005
R5527 vdd.n3147 vdd.n3146 9.3005
R5528 vdd.n3086 vdd.n3085 9.3005
R5529 vdd.n2688 vdd.n2687 9.3005
R5530 vdd.n3040 vdd.n3039 9.3005
R5531 vdd.n2703 vdd.n2702 9.3005
R5532 vdd.n3002 vdd.n3001 9.3005
R5533 vdd.n2751 vdd.n2750 9.3005
R5534 vdd.n2949 vdd.n2948 9.3005
R5535 vdd.n2959 vdd.n2958 9.3005
R5536 vdd.n2919 vdd.n2918 9.3005
R5537 vdd.n4017 vdd.n4016 9.3005
R5538 vdd.n2828 vdd.n2827 9.3005
R5539 vdd.n2811 vdd.n2805 9.3005
R5540 vdd.n2870 vdd.n2869 9.3005
R5541 vdd.n2877 vdd.n2876 9.3005
R5542 vdd.n1128 vdd.n1127 9.3005
R5543 vdd.n1131 vdd.n1130 9.3005
R5544 vdd.n4423 vdd.n4422 9.3005
R5545 vdd.n1392 vdd.n1391 9.3005
R5546 vdd.n1395 vdd.n1394 9.3005
R5547 vdd.n4302 vdd.n4301 9.3005
R5548 vdd.n1656 vdd.n1655 9.3005
R5549 vdd.n1659 vdd.n1658 9.3005
R5550 vdd.n4181 vdd.n4180 9.3005
R5551 vdd.n1920 vdd.n1919 9.3005
R5552 vdd.n1923 vdd.n1922 9.3005
R5553 vdd.n4060 vdd.n4059 9.3005
R5554 vdd.n2012 vdd.n2011 9.3005
R5555 vdd.n4082 vdd.n4081 9.3005
R5556 vdd.n1970 vdd.n1969 9.3005
R5557 vdd.n4104 vdd.n4103 9.3005
R5558 vdd.n1914 vdd.n1870 9.3005
R5559 vdd.n1886 vdd.n1885 9.3005
R5560 vdd.n1859 vdd.n1858 9.3005
R5561 vdd.n1847 vdd.n1806 9.3005
R5562 vdd.n1817 vdd.n1816 9.3005
R5563 vdd.n1748 vdd.n1747 9.3005
R5564 vdd.n4203 vdd.n4202 9.3005
R5565 vdd.n1706 vdd.n1705 9.3005
R5566 vdd.n4225 vdd.n4224 9.3005
R5567 vdd.n1650 vdd.n1606 9.3005
R5568 vdd.n1622 vdd.n1621 9.3005
R5569 vdd.n1595 vdd.n1594 9.3005
R5570 vdd.n1583 vdd.n1542 9.3005
R5571 vdd.n1553 vdd.n1552 9.3005
R5572 vdd.n1484 vdd.n1483 9.3005
R5573 vdd.n4324 vdd.n4323 9.3005
R5574 vdd.n1442 vdd.n1441 9.3005
R5575 vdd.n4346 vdd.n4345 9.3005
R5576 vdd.n1386 vdd.n1342 9.3005
R5577 vdd.n1358 vdd.n1357 9.3005
R5578 vdd.n1331 vdd.n1330 9.3005
R5579 vdd.n1319 vdd.n1278 9.3005
R5580 vdd.n1289 vdd.n1288 9.3005
R5581 vdd.n1220 vdd.n1219 9.3005
R5582 vdd.n4445 vdd.n4444 9.3005
R5583 vdd.n1178 vdd.n1177 9.3005
R5584 vdd.n4467 vdd.n4466 9.3005
R5585 vdd.n1122 vdd.n1078 9.3005
R5586 vdd.n1094 vdd.n1093 9.3005
R5587 vdd.n1055 vdd.n1010 9.3005
R5588 vdd.n1067 vdd.n1066 9.3005
R5589 vdd.n1025 vdd.n1024 9.3005
R5590 vdd.n898 vdd.n897 9.3005
R5591 vdd.n928 vdd.n862 9.3005
R5592 vdd.n940 vdd.n939 9.3005
R5593 vdd.n967 vdd.n966 9.3005
R5594 vdd.n994 vdd.n951 9.3005
R5595 vdd.n3859 vdd.n3858 9.3005
R5596 vdd.n3794 vdd.n3793 9.3005
R5597 vdd.n3794 vdd.n2258 9.3005
R5598 vdd.n3759 vdd.n2276 9.3005
R5599 vdd.n3760 vdd.n3759 9.3005
R5600 vdd.n3731 vdd.n2282 9.3005
R5601 vdd.n3731 vdd.n3730 9.3005
R5602 vdd.n3724 vdd.n3723 9.3005
R5603 vdd.n3725 vdd.n3724 9.3005
R5604 vdd.n3801 vdd.n3800 9.3005
R5605 vdd.n3703 vdd.n3702 9.3005
R5606 vdd.n3704 vdd.n3703 9.3005
R5607 vdd.n3704 vdd.n2065 9.3005
R5608 vdd.n3672 vdd.n3671 9.3005
R5609 vdd.n3671 vdd.n2329 9.3005
R5610 vdd.n3664 vdd.n3663 9.3005
R5611 vdd.n3665 vdd.n3664 9.3005
R5612 vdd.n3624 vdd.n2355 9.3005
R5613 vdd.n3638 vdd.n2355 9.3005
R5614 vdd.n3611 vdd.n3610 9.3005
R5615 vdd.n3610 vdd.n3609 9.3005
R5616 vdd.n3692 vdd.n3691 9.3005
R5617 vdd.n3691 vdd.n3690 9.3005
R5618 vdd.n3690 vdd.n2065 9.3005
R5619 vdd.n3590 vdd.n3589 9.3005
R5620 vdd.n3589 vdd.n2369 9.3005
R5621 vdd.n2369 vdd.n2065 9.3005
R5622 vdd.n2396 vdd.n2395 9.3005
R5623 vdd.n3546 vdd.n2396 9.3005
R5624 vdd.n3527 vdd.n3526 9.3005
R5625 vdd.n3526 vdd.n3525 9.3005
R5626 vdd.n3519 vdd.n3518 9.3005
R5627 vdd.n3519 vdd.n2413 9.3005
R5628 vdd.n3488 vdd.n2429 9.3005
R5629 vdd.n3489 vdd.n3488 9.3005
R5630 vdd.n3579 vdd.n3578 9.3005
R5631 vdd.n3580 vdd.n3579 9.3005
R5632 vdd.n2454 vdd.n2435 9.3005
R5633 vdd.n2454 vdd.n2453 9.3005
R5634 vdd.n2453 vdd.n2065 9.3005
R5635 vdd.n3444 vdd.n3443 9.3005
R5636 vdd.n3443 vdd.n2464 9.3005
R5637 vdd.n3436 vdd.n3435 9.3005
R5638 vdd.n3437 vdd.n3436 9.3005
R5639 vdd.n3396 vdd.n2490 9.3005
R5640 vdd.n3410 vdd.n2490 9.3005
R5641 vdd.n3383 vdd.n3382 9.3005
R5642 vdd.n3382 vdd.n3381 9.3005
R5643 vdd.n3465 vdd.n3464 9.3005
R5644 vdd.n3464 vdd.n3463 9.3005
R5645 vdd.n3463 vdd.n2065 9.3005
R5646 vdd.n3362 vdd.n3361 9.3005
R5647 vdd.n3361 vdd.n2504 9.3005
R5648 vdd.n2504 vdd.n2065 9.3005
R5649 vdd.n2531 vdd.n2530 9.3005
R5650 vdd.n3318 vdd.n2531 9.3005
R5651 vdd.n3299 vdd.n3298 9.3005
R5652 vdd.n3298 vdd.n3297 9.3005
R5653 vdd.n3291 vdd.n3290 9.3005
R5654 vdd.n3291 vdd.n2548 9.3005
R5655 vdd.n3260 vdd.n2564 9.3005
R5656 vdd.n3261 vdd.n3260 9.3005
R5657 vdd.n3351 vdd.n3350 9.3005
R5658 vdd.n3352 vdd.n3351 9.3005
R5659 vdd.n2589 vdd.n2570 9.3005
R5660 vdd.n2589 vdd.n2588 9.3005
R5661 vdd.n2588 vdd.n2065 9.3005
R5662 vdd.n3216 vdd.n3215 9.3005
R5663 vdd.n3215 vdd.n2599 9.3005
R5664 vdd.n3208 vdd.n3207 9.3005
R5665 vdd.n3209 vdd.n3208 9.3005
R5666 vdd.n3168 vdd.n2625 9.3005
R5667 vdd.n3182 vdd.n2625 9.3005
R5668 vdd.n3155 vdd.n3154 9.3005
R5669 vdd.n3154 vdd.n3153 9.3005
R5670 vdd.n3237 vdd.n3236 9.3005
R5671 vdd.n3236 vdd.n3235 9.3005
R5672 vdd.n3235 vdd.n2065 9.3005
R5673 vdd.n3134 vdd.n3133 9.3005
R5674 vdd.n3133 vdd.n2639 9.3005
R5675 vdd.n2639 vdd.n2065 9.3005
R5676 vdd.n2666 vdd.n2665 9.3005
R5677 vdd.n3090 vdd.n2666 9.3005
R5678 vdd.n3071 vdd.n3070 9.3005
R5679 vdd.n3070 vdd.n3069 9.3005
R5680 vdd.n3063 vdd.n3062 9.3005
R5681 vdd.n3063 vdd.n2683 9.3005
R5682 vdd.n3032 vdd.n2699 9.3005
R5683 vdd.n3033 vdd.n3032 9.3005
R5684 vdd.n3123 vdd.n3122 9.3005
R5685 vdd.n3124 vdd.n3123 9.3005
R5686 vdd.n2724 vdd.n2705 9.3005
R5687 vdd.n2724 vdd.n2723 9.3005
R5688 vdd.n2723 vdd.n2065 9.3005
R5689 vdd.n2988 vdd.n2987 9.3005
R5690 vdd.n2987 vdd.n2734 9.3005
R5691 vdd.n2980 vdd.n2979 9.3005
R5692 vdd.n2981 vdd.n2980 9.3005
R5693 vdd.n2927 vdd.n2926 9.3005
R5694 vdd.n2926 vdd.n2925 9.3005
R5695 vdd.n2940 vdd.n2760 9.3005
R5696 vdd.n2954 vdd.n2760 9.3005
R5697 vdd.n3009 vdd.n3008 9.3005
R5698 vdd.n3008 vdd.n3007 9.3005
R5699 vdd.n3007 vdd.n2065 9.3005
R5700 vdd.n2906 vdd.n2905 9.3005
R5701 vdd.n4021 vdd.n4020 9.3005
R5702 vdd.n4021 vdd.n2066 9.3005
R5703 vdd.n4025 vdd.n2066 9.3005
R5704 vdd.n4029 vdd.n4028 9.3005
R5705 vdd.n4028 vdd.n4027 9.3005
R5706 vdd.n2849 vdd.n2848 9.3005
R5707 vdd.n2850 vdd.n2849 9.3005
R5708 vdd.n2857 vdd.n2856 9.3005
R5709 vdd.n2856 vdd.n2855 9.3005
R5710 vdd.n2884 vdd.n2883 9.3005
R5711 vdd.n2883 vdd.n2882 9.3005
R5712 vdd.n2786 vdd.n2064 9.3005
R5713 vdd.n4025 vdd.n2064 9.3005
R5714 vdd.n3865 vdd.n3864 9.3005
R5715 vdd.n3865 vdd.n3837 9.3005
R5716 vdd.n3978 vdd.n3837 9.3005
R5717 vdd.n4068 vdd.n4067 9.3005
R5718 vdd.n4067 vdd.n4066 9.3005
R5719 vdd.n4066 vdd.n4065 9.3005
R5720 vdd.n2005 vdd.n1980 9.3005
R5721 vdd.n2005 vdd.n1977 9.3005
R5722 vdd.n1977 vdd.n1976 9.3005
R5723 vdd.n4090 vdd.n4089 9.3005
R5724 vdd.n4089 vdd.n4088 9.3005
R5725 vdd.n4088 vdd.n4087 9.3005
R5726 vdd.n1963 vdd.n1938 9.3005
R5727 vdd.n1963 vdd.n1935 9.3005
R5728 vdd.n1935 vdd.n1934 9.3005
R5729 vdd.n3919 vdd.n2022 9.3005
R5730 vdd.n3919 vdd.n2019 9.3005
R5731 vdd.n2019 vdd.n2018 9.3005
R5732 vdd.n4112 vdd.n4111 9.3005
R5733 vdd.n4111 vdd.n4110 9.3005
R5734 vdd.n4110 vdd.n4109 9.3005
R5735 vdd.n4129 vdd.n4128 9.3005
R5736 vdd.n4129 vdd.n1865 9.3005
R5737 vdd.n1865 vdd.n1864 9.3005
R5738 vdd.n4137 vdd.n4136 9.3005
R5739 vdd.n4136 vdd.n4135 9.3005
R5740 vdd.n4135 vdd.n4134 9.3005
R5741 vdd.n1854 vdd.n1808 9.3005
R5742 vdd.n1854 vdd.n1846 9.3005
R5743 vdd.n1846 vdd.n1845 9.3005
R5744 vdd.n4156 vdd.n4155 9.3005
R5745 vdd.n4156 vdd.n1801 9.3005
R5746 vdd.n1801 vdd.n1800 9.3005
R5747 vdd.n1930 vdd.n1872 9.3005
R5748 vdd.n1931 vdd.n1930 9.3005
R5749 vdd.n1932 vdd.n1931 9.3005
R5750 vdd.n4164 vdd.n4163 9.3005
R5751 vdd.n4163 vdd.n4162 9.3005
R5752 vdd.n4162 vdd.n4161 9.3005
R5753 vdd.n4189 vdd.n4188 9.3005
R5754 vdd.n4188 vdd.n4187 9.3005
R5755 vdd.n4187 vdd.n4186 9.3005
R5756 vdd.n1741 vdd.n1716 9.3005
R5757 vdd.n1741 vdd.n1713 9.3005
R5758 vdd.n1713 vdd.n1712 9.3005
R5759 vdd.n4211 vdd.n4210 9.3005
R5760 vdd.n4210 vdd.n4209 9.3005
R5761 vdd.n4209 vdd.n4208 9.3005
R5762 vdd.n1699 vdd.n1674 9.3005
R5763 vdd.n1699 vdd.n1671 9.3005
R5764 vdd.n1671 vdd.n1670 9.3005
R5765 vdd.n1789 vdd.n1758 9.3005
R5766 vdd.n1789 vdd.n1755 9.3005
R5767 vdd.n1755 vdd.n1754 9.3005
R5768 vdd.n4233 vdd.n4232 9.3005
R5769 vdd.n4232 vdd.n4231 9.3005
R5770 vdd.n4231 vdd.n4230 9.3005
R5771 vdd.n4250 vdd.n4249 9.3005
R5772 vdd.n4250 vdd.n1601 9.3005
R5773 vdd.n1601 vdd.n1600 9.3005
R5774 vdd.n4258 vdd.n4257 9.3005
R5775 vdd.n4257 vdd.n4256 9.3005
R5776 vdd.n4256 vdd.n4255 9.3005
R5777 vdd.n1590 vdd.n1544 9.3005
R5778 vdd.n1590 vdd.n1582 9.3005
R5779 vdd.n1582 vdd.n1581 9.3005
R5780 vdd.n4277 vdd.n4276 9.3005
R5781 vdd.n4277 vdd.n1537 9.3005
R5782 vdd.n1537 vdd.n1536 9.3005
R5783 vdd.n1666 vdd.n1608 9.3005
R5784 vdd.n1667 vdd.n1666 9.3005
R5785 vdd.n1668 vdd.n1667 9.3005
R5786 vdd.n4285 vdd.n4284 9.3005
R5787 vdd.n4284 vdd.n4283 9.3005
R5788 vdd.n4283 vdd.n4282 9.3005
R5789 vdd.n4310 vdd.n4309 9.3005
R5790 vdd.n4309 vdd.n4308 9.3005
R5791 vdd.n4308 vdd.n4307 9.3005
R5792 vdd.n1477 vdd.n1452 9.3005
R5793 vdd.n1477 vdd.n1449 9.3005
R5794 vdd.n1449 vdd.n1448 9.3005
R5795 vdd.n4332 vdd.n4331 9.3005
R5796 vdd.n4331 vdd.n4330 9.3005
R5797 vdd.n4330 vdd.n4329 9.3005
R5798 vdd.n1435 vdd.n1410 9.3005
R5799 vdd.n1435 vdd.n1407 9.3005
R5800 vdd.n1407 vdd.n1406 9.3005
R5801 vdd.n1525 vdd.n1494 9.3005
R5802 vdd.n1525 vdd.n1491 9.3005
R5803 vdd.n1491 vdd.n1490 9.3005
R5804 vdd.n4354 vdd.n4353 9.3005
R5805 vdd.n4353 vdd.n4352 9.3005
R5806 vdd.n4352 vdd.n4351 9.3005
R5807 vdd.n4371 vdd.n4370 9.3005
R5808 vdd.n4371 vdd.n1337 9.3005
R5809 vdd.n1337 vdd.n1336 9.3005
R5810 vdd.n4379 vdd.n4378 9.3005
R5811 vdd.n4378 vdd.n4377 9.3005
R5812 vdd.n4377 vdd.n4376 9.3005
R5813 vdd.n1326 vdd.n1280 9.3005
R5814 vdd.n1326 vdd.n1318 9.3005
R5815 vdd.n1318 vdd.n1317 9.3005
R5816 vdd.n4398 vdd.n4397 9.3005
R5817 vdd.n4398 vdd.n1273 9.3005
R5818 vdd.n1273 vdd.n1272 9.3005
R5819 vdd.n1402 vdd.n1344 9.3005
R5820 vdd.n1403 vdd.n1402 9.3005
R5821 vdd.n1404 vdd.n1403 9.3005
R5822 vdd.n4406 vdd.n4405 9.3005
R5823 vdd.n4405 vdd.n4404 9.3005
R5824 vdd.n4404 vdd.n4403 9.3005
R5825 vdd.n4431 vdd.n4430 9.3005
R5826 vdd.n4430 vdd.n4429 9.3005
R5827 vdd.n4429 vdd.n4428 9.3005
R5828 vdd.n1213 vdd.n1188 9.3005
R5829 vdd.n1213 vdd.n1185 9.3005
R5830 vdd.n1185 vdd.n1184 9.3005
R5831 vdd.n4453 vdd.n4452 9.3005
R5832 vdd.n4452 vdd.n4451 9.3005
R5833 vdd.n4451 vdd.n4450 9.3005
R5834 vdd.n1171 vdd.n1146 9.3005
R5835 vdd.n1171 vdd.n1143 9.3005
R5836 vdd.n1143 vdd.n1142 9.3005
R5837 vdd.n1261 vdd.n1230 9.3005
R5838 vdd.n1261 vdd.n1227 9.3005
R5839 vdd.n1227 vdd.n1226 9.3005
R5840 vdd.n4475 vdd.n4474 9.3005
R5841 vdd.n4474 vdd.n4473 9.3005
R5842 vdd.n4473 vdd.n4472 9.3005
R5843 vdd.n4492 vdd.n4491 9.3005
R5844 vdd.n4492 vdd.n1073 9.3005
R5845 vdd.n1073 vdd.n1072 9.3005
R5846 vdd.n4500 vdd.n4499 9.3005
R5847 vdd.n4499 vdd.n4498 9.3005
R5848 vdd.n4498 vdd.n4497 9.3005
R5849 vdd.n4519 vdd.n4518 9.3005
R5850 vdd.n4519 vdd.n1005 9.3005
R5851 vdd.n1005 vdd.n1004 9.3005
R5852 vdd.n1062 vdd.n1012 9.3005
R5853 vdd.n1062 vdd.n1054 9.3005
R5854 vdd.n1054 vdd.n1053 9.3005
R5855 vdd.n1138 vdd.n1080 9.3005
R5856 vdd.n1139 vdd.n1138 9.3005
R5857 vdd.n1140 vdd.n1139 9.3005
R5858 vdd.n4527 vdd.n4526 9.3005
R5859 vdd.n4526 vdd.n4525 9.3005
R5860 vdd.n4525 vdd.n4524 9.3005
R5861 vdd.n4578 vdd.n854 9.3005
R5862 vdd.n4578 vdd.n4577 9.3005
R5863 vdd.n4577 vdd.n4576 9.3005
R5864 vdd.n4571 vdd.n4570 9.3005
R5865 vdd.n4571 vdd.n857 9.3005
R5866 vdd.n857 vdd.n856 9.3005
R5867 vdd.n935 vdd.n864 9.3005
R5868 vdd.n935 vdd.n927 9.3005
R5869 vdd.n927 vdd.n926 9.3005
R5870 vdd.n4552 vdd.n4551 9.3005
R5871 vdd.n4551 vdd.n4550 9.3005
R5872 vdd.n4550 vdd.n4549 9.3005
R5873 vdd.n4544 vdd.n4543 9.3005
R5874 vdd.n4544 vdd.n946 9.3005
R5875 vdd.n946 vdd.n945 9.3005
R5876 vdd.n1000 vdd.n999 9.3005
R5877 vdd.n1001 vdd.n1000 9.3005
R5878 vdd.n4618 vdd.n4617 9.3005
R5879 vdd.n4619 vdd.n4618 9.3005
R5880 vdd.n4620 vdd.n4619 9.3005
R5881 vdd.n4607 vdd.n4588 9.3005
R5882 vdd.n756 vdd.n755 9.3005
R5883 vdd.n742 vdd.n740 9.3005
R5884 vdd.n4870 vdd.n4869 9.3005
R5885 vdd.n621 vdd.n620 9.3005
R5886 vdd.n607 vdd.n605 9.3005
R5887 vdd.n5098 vdd.n5097 9.3005
R5888 vdd.n486 vdd.n485 9.3005
R5889 vdd.n472 vdd.n470 9.3005
R5890 vdd.n5326 vdd.n5325 9.3005
R5891 vdd.n351 vdd.n350 9.3005
R5892 vdd.n345 vdd.n344 9.3005
R5893 vdd.n289 vdd.n288 9.3005
R5894 vdd.n5543 vdd.n5542 9.3005
R5895 vdd.n306 vdd.n305 9.3005
R5896 vdd.n5510 vdd.n5509 9.3005
R5897 vdd.n5485 vdd.n5484 9.3005
R5898 vdd.n5459 vdd.n5458 9.3005
R5899 vdd.n370 vdd.n369 9.3005
R5900 vdd.n5417 vdd.n5416 9.3005
R5901 vdd.n5407 vdd.n5406 9.3005
R5902 vdd.n5377 vdd.n5376 9.3005
R5903 vdd.n5316 vdd.n5315 9.3005
R5904 vdd.n442 vdd.n441 9.3005
R5905 vdd.n5270 vdd.n5269 9.3005
R5906 vdd.n457 vdd.n456 9.3005
R5907 vdd.n5232 vdd.n5231 9.3005
R5908 vdd.n505 vdd.n504 9.3005
R5909 vdd.n5189 vdd.n5188 9.3005
R5910 vdd.n5179 vdd.n5178 9.3005
R5911 vdd.n5149 vdd.n5148 9.3005
R5912 vdd.n5088 vdd.n5087 9.3005
R5913 vdd.n577 vdd.n576 9.3005
R5914 vdd.n5042 vdd.n5041 9.3005
R5915 vdd.n592 vdd.n591 9.3005
R5916 vdd.n5004 vdd.n5003 9.3005
R5917 vdd.n640 vdd.n639 9.3005
R5918 vdd.n4961 vdd.n4960 9.3005
R5919 vdd.n4951 vdd.n4950 9.3005
R5920 vdd.n4921 vdd.n4920 9.3005
R5921 vdd.n4860 vdd.n4859 9.3005
R5922 vdd.n712 vdd.n711 9.3005
R5923 vdd.n4814 vdd.n4813 9.3005
R5924 vdd.n727 vdd.n726 9.3005
R5925 vdd.n4776 vdd.n4775 9.3005
R5926 vdd.n775 vdd.n774 9.3005
R5927 vdd.n4723 vdd.n4722 9.3005
R5928 vdd.n4733 vdd.n4732 9.3005
R5929 vdd.n4693 vdd.n4692 9.3005
R5930 vdd.n5570 vdd.n5569 9.3005
R5931 vdd.n5570 vdd.n284 9.3005
R5932 vdd.n5535 vdd.n302 9.3005
R5933 vdd.n5536 vdd.n5535 9.3005
R5934 vdd.n5507 vdd.n308 9.3005
R5935 vdd.n5507 vdd.n5506 9.3005
R5936 vdd.n5500 vdd.n5499 9.3005
R5937 vdd.n5501 vdd.n5500 9.3005
R5938 vdd.n5577 vdd.n5576 9.3005
R5939 vdd.n5478 vdd.n5477 9.3005
R5940 vdd.n5479 vdd.n5478 9.3005
R5941 vdd.n5479 vdd.n250 9.3005
R5942 vdd.n5446 vdd.n5445 9.3005
R5943 vdd.n5445 vdd.n353 9.3005
R5944 vdd.n5438 vdd.n5437 9.3005
R5945 vdd.n5439 vdd.n5438 9.3005
R5946 vdd.n5398 vdd.n379 9.3005
R5947 vdd.n5412 vdd.n379 9.3005
R5948 vdd.n5385 vdd.n5384 9.3005
R5949 vdd.n5384 vdd.n5383 9.3005
R5950 vdd.n5466 vdd.n5465 9.3005
R5951 vdd.n5465 vdd.n5464 9.3005
R5952 vdd.n5464 vdd.n250 9.3005
R5953 vdd.n5364 vdd.n5363 9.3005
R5954 vdd.n5363 vdd.n393 9.3005
R5955 vdd.n393 vdd.n250 9.3005
R5956 vdd.n420 vdd.n419 9.3005
R5957 vdd.n5320 vdd.n420 9.3005
R5958 vdd.n5301 vdd.n5300 9.3005
R5959 vdd.n5300 vdd.n5299 9.3005
R5960 vdd.n5293 vdd.n5292 9.3005
R5961 vdd.n5293 vdd.n437 9.3005
R5962 vdd.n5262 vdd.n453 9.3005
R5963 vdd.n5263 vdd.n5262 9.3005
R5964 vdd.n5353 vdd.n5352 9.3005
R5965 vdd.n5354 vdd.n5353 9.3005
R5966 vdd.n478 vdd.n459 9.3005
R5967 vdd.n478 vdd.n477 9.3005
R5968 vdd.n477 vdd.n250 9.3005
R5969 vdd.n5218 vdd.n5217 9.3005
R5970 vdd.n5217 vdd.n488 9.3005
R5971 vdd.n5210 vdd.n5209 9.3005
R5972 vdd.n5211 vdd.n5210 9.3005
R5973 vdd.n5170 vdd.n514 9.3005
R5974 vdd.n5184 vdd.n514 9.3005
R5975 vdd.n5157 vdd.n5156 9.3005
R5976 vdd.n5156 vdd.n5155 9.3005
R5977 vdd.n5239 vdd.n5238 9.3005
R5978 vdd.n5238 vdd.n5237 9.3005
R5979 vdd.n5237 vdd.n250 9.3005
R5980 vdd.n5136 vdd.n5135 9.3005
R5981 vdd.n5135 vdd.n528 9.3005
R5982 vdd.n528 vdd.n250 9.3005
R5983 vdd.n555 vdd.n554 9.3005
R5984 vdd.n5092 vdd.n555 9.3005
R5985 vdd.n5073 vdd.n5072 9.3005
R5986 vdd.n5072 vdd.n5071 9.3005
R5987 vdd.n5065 vdd.n5064 9.3005
R5988 vdd.n5065 vdd.n572 9.3005
R5989 vdd.n5034 vdd.n588 9.3005
R5990 vdd.n5035 vdd.n5034 9.3005
R5991 vdd.n5125 vdd.n5124 9.3005
R5992 vdd.n5126 vdd.n5125 9.3005
R5993 vdd.n613 vdd.n594 9.3005
R5994 vdd.n613 vdd.n612 9.3005
R5995 vdd.n612 vdd.n250 9.3005
R5996 vdd.n4990 vdd.n4989 9.3005
R5997 vdd.n4989 vdd.n623 9.3005
R5998 vdd.n4982 vdd.n4981 9.3005
R5999 vdd.n4983 vdd.n4982 9.3005
R6000 vdd.n4942 vdd.n649 9.3005
R6001 vdd.n4956 vdd.n649 9.3005
R6002 vdd.n4929 vdd.n4928 9.3005
R6003 vdd.n4928 vdd.n4927 9.3005
R6004 vdd.n5011 vdd.n5010 9.3005
R6005 vdd.n5010 vdd.n5009 9.3005
R6006 vdd.n5009 vdd.n250 9.3005
R6007 vdd.n4908 vdd.n4907 9.3005
R6008 vdd.n4907 vdd.n663 9.3005
R6009 vdd.n663 vdd.n250 9.3005
R6010 vdd.n690 vdd.n689 9.3005
R6011 vdd.n4864 vdd.n690 9.3005
R6012 vdd.n4845 vdd.n4844 9.3005
R6013 vdd.n4844 vdd.n4843 9.3005
R6014 vdd.n4837 vdd.n4836 9.3005
R6015 vdd.n4837 vdd.n707 9.3005
R6016 vdd.n4806 vdd.n723 9.3005
R6017 vdd.n4807 vdd.n4806 9.3005
R6018 vdd.n4897 vdd.n4896 9.3005
R6019 vdd.n4898 vdd.n4897 9.3005
R6020 vdd.n748 vdd.n729 9.3005
R6021 vdd.n748 vdd.n747 9.3005
R6022 vdd.n747 vdd.n250 9.3005
R6023 vdd.n4762 vdd.n4761 9.3005
R6024 vdd.n4761 vdd.n758 9.3005
R6025 vdd.n4754 vdd.n4753 9.3005
R6026 vdd.n4755 vdd.n4754 9.3005
R6027 vdd.n4701 vdd.n4700 9.3005
R6028 vdd.n4700 vdd.n4699 9.3005
R6029 vdd.n4714 vdd.n784 9.3005
R6030 vdd.n4728 vdd.n784 9.3005
R6031 vdd.n4783 vdd.n4782 9.3005
R6032 vdd.n4782 vdd.n4781 9.3005
R6033 vdd.n4781 vdd.n250 9.3005
R6034 vdd.n4680 vdd.n4679 9.3005
R6035 vdd.n5666 vdd.n5626 9.3005
R6036 vdd.n5666 vdd.n5665 9.3005
R6037 vdd.n5700 vdd.n5611 9.3005
R6038 vdd.n5700 vdd.n5699 9.3005
R6039 vdd.n5720 vdd.n5719 9.3005
R6040 vdd.n5721 vdd.n5720 9.3005
R6041 vdd.n5619 vdd.n5608 9.3005
R6042 vdd.n5619 vdd.n5618 9.3005
R6043 vdd.n5681 vdd.n5680 9.3005
R6044 vdd.n5680 vdd.n5679 9.3005
R6045 vdd.n5726 vdd.n5725 9.3005
R6046 vdd.n5727 vdd.n5726 9.3005
R6047 vdd.n5756 vdd.n5755 9.3005
R6048 vdd.n7467 vdd.n7466 9.3005
R6049 vdd.n7466 vdd.n7465 9.3005
R6050 vdd.n7465 vdd.n7464 9.3005
R6051 vdd.n4005 vdd.t26 9.19352
R6052 vdd.n6411 vdd.n6410 8.92171
R6053 vdd.n6432 vdd.n6431 8.92171
R6054 vdd.n6364 vdd.n6358 8.92171
R6055 vdd.n6475 vdd.n6474 8.92171
R6056 vdd.n6495 vdd.n6494 8.92171
R6057 vdd.n6523 vdd.n6313 8.92171
R6058 vdd.n6314 vdd.n6300 8.92171
R6059 vdd.n6556 vdd.n6555 8.92171
R6060 vdd.n6285 vdd.n6280 8.92171
R6061 vdd.n6602 vdd.n6601 8.92171
R6062 vdd.n6638 vdd.n6637 8.92171
R6063 vdd.n6659 vdd.n6658 8.92171
R6064 vdd.n6231 vdd.n6225 8.92171
R6065 vdd.n6702 vdd.n6701 8.92171
R6066 vdd.n6722 vdd.n6721 8.92171
R6067 vdd.n6750 vdd.n6180 8.92171
R6068 vdd.n6181 vdd.n6167 8.92171
R6069 vdd.n6783 vdd.n6782 8.92171
R6070 vdd.n6152 vdd.n6147 8.92171
R6071 vdd.n6829 vdd.n6828 8.92171
R6072 vdd.n6865 vdd.n6864 8.92171
R6073 vdd.n6886 vdd.n6885 8.92171
R6074 vdd.n6098 vdd.n6092 8.92171
R6075 vdd.n6929 vdd.n6928 8.92171
R6076 vdd.n6949 vdd.n6948 8.92171
R6077 vdd.n6977 vdd.n6047 8.92171
R6078 vdd.n6048 vdd.n6034 8.92171
R6079 vdd.n7010 vdd.n7009 8.92171
R6080 vdd.n6019 vdd.n6014 8.92171
R6081 vdd.n7056 vdd.n7055 8.92171
R6082 vdd.n7092 vdd.n7091 8.92171
R6083 vdd.n7113 vdd.n7112 8.92171
R6084 vdd.n5965 vdd.n5959 8.92171
R6085 vdd.n7156 vdd.n7155 8.92171
R6086 vdd.n7176 vdd.n7175 8.92171
R6087 vdd.n7204 vdd.n5914 8.92171
R6088 vdd.n5915 vdd.n5901 8.92171
R6089 vdd.n7237 vdd.n7236 8.92171
R6090 vdd.n5886 vdd.n5881 8.92171
R6091 vdd.n7288 vdd.n7287 8.92171
R6092 vdd.n7317 vdd.n7316 8.92171
R6093 vdd.n7336 vdd.n7335 8.92171
R6094 vdd.n7355 vdd.n7354 8.92171
R6095 vdd.n7374 vdd.n7373 8.92171
R6096 vdd.n7397 vdd.n7396 8.92171
R6097 vdd.n5723 vdd.n262 8.92171
R6098 vdd.n5613 vdd.n5612 8.92171
R6099 vdd.n5623 vdd.n5622 8.92171
R6100 vdd.n5696 vdd.n5695 8.92171
R6101 vdd.n5677 vdd.n5670 8.92171
R6102 vdd.n2920 vdd.n2919 8.92171
R6103 vdd.n2950 vdd.n2949 8.92171
R6104 vdd.n2958 vdd.n2957 8.92171
R6105 vdd.n2750 vdd.n2744 8.92171
R6106 vdd.n3003 vdd.n3002 8.92171
R6107 vdd.n2719 vdd.n2702 8.92171
R6108 vdd.n3039 vdd.n3038 8.92171
R6109 vdd.n2687 vdd.n2682 8.92171
R6110 vdd.n3087 vdd.n3086 8.92171
R6111 vdd.n3095 vdd.n3094 8.92171
R6112 vdd.n3148 vdd.n3147 8.92171
R6113 vdd.n3178 vdd.n3177 8.92171
R6114 vdd.n3186 vdd.n3185 8.92171
R6115 vdd.n2615 vdd.n2609 8.92171
R6116 vdd.n3231 vdd.n3230 8.92171
R6117 vdd.n2584 vdd.n2567 8.92171
R6118 vdd.n3267 vdd.n3266 8.92171
R6119 vdd.n2552 vdd.n2547 8.92171
R6120 vdd.n3315 vdd.n3314 8.92171
R6121 vdd.n3323 vdd.n3322 8.92171
R6122 vdd.n3376 vdd.n3375 8.92171
R6123 vdd.n3406 vdd.n3405 8.92171
R6124 vdd.n3414 vdd.n3413 8.92171
R6125 vdd.n2480 vdd.n2474 8.92171
R6126 vdd.n3459 vdd.n3458 8.92171
R6127 vdd.n2449 vdd.n2432 8.92171
R6128 vdd.n3495 vdd.n3494 8.92171
R6129 vdd.n2417 vdd.n2412 8.92171
R6130 vdd.n3543 vdd.n3542 8.92171
R6131 vdd.n3551 vdd.n3550 8.92171
R6132 vdd.n3604 vdd.n3603 8.92171
R6133 vdd.n3634 vdd.n3633 8.92171
R6134 vdd.n3642 vdd.n3641 8.92171
R6135 vdd.n2345 vdd.n2339 8.92171
R6136 vdd.n3686 vdd.n3685 8.92171
R6137 vdd.n3709 vdd.n3708 8.92171
R6138 vdd.n3733 vdd.n2292 8.92171
R6139 vdd.n2293 vdd.n2279 8.92171
R6140 vdd.n3766 vdd.n3765 8.92171
R6141 vdd.n2262 vdd.n2257 8.92171
R6142 vdd.n4016 vdd.n4015 8.92171
R6143 vdd.n2827 vdd.n2826 8.92171
R6144 vdd.n2852 vdd.n2805 8.92171
R6145 vdd.n2871 vdd.n2870 8.92171
R6146 vdd.n2880 vdd.n2877 8.92171
R6147 vdd.n1024 vdd.n1006 8.92171
R6148 vdd.n1056 vdd.n1055 8.92171
R6149 vdd.n1068 vdd.n1067 8.92171
R6150 vdd.n1093 vdd.n1074 8.92171
R6151 vdd.n1125 vdd.n1122 8.92171
R6152 vdd.n4468 vdd.n4467 8.92171
R6153 vdd.n1179 vdd.n1178 8.92171
R6154 vdd.n4446 vdd.n4445 8.92171
R6155 vdd.n1221 vdd.n1220 8.92171
R6156 vdd.n4424 vdd.n4423 8.92171
R6157 vdd.n1288 vdd.n1274 8.92171
R6158 vdd.n1320 vdd.n1319 8.92171
R6159 vdd.n1332 vdd.n1331 8.92171
R6160 vdd.n1357 vdd.n1338 8.92171
R6161 vdd.n1389 vdd.n1386 8.92171
R6162 vdd.n4347 vdd.n4346 8.92171
R6163 vdd.n1443 vdd.n1442 8.92171
R6164 vdd.n4325 vdd.n4324 8.92171
R6165 vdd.n1485 vdd.n1484 8.92171
R6166 vdd.n4303 vdd.n4302 8.92171
R6167 vdd.n1552 vdd.n1538 8.92171
R6168 vdd.n1584 vdd.n1583 8.92171
R6169 vdd.n1596 vdd.n1595 8.92171
R6170 vdd.n1621 vdd.n1602 8.92171
R6171 vdd.n1653 vdd.n1650 8.92171
R6172 vdd.n4226 vdd.n4225 8.92171
R6173 vdd.n1707 vdd.n1706 8.92171
R6174 vdd.n4204 vdd.n4203 8.92171
R6175 vdd.n1749 vdd.n1748 8.92171
R6176 vdd.n4182 vdd.n4181 8.92171
R6177 vdd.n1816 vdd.n1802 8.92171
R6178 vdd.n1848 vdd.n1847 8.92171
R6179 vdd.n1860 vdd.n1859 8.92171
R6180 vdd.n1885 vdd.n1866 8.92171
R6181 vdd.n1917 vdd.n1914 8.92171
R6182 vdd.n4105 vdd.n4104 8.92171
R6183 vdd.n1971 vdd.n1970 8.92171
R6184 vdd.n4083 vdd.n4082 8.92171
R6185 vdd.n2013 vdd.n2012 8.92171
R6186 vdd.n4061 vdd.n4060 8.92171
R6187 vdd.n897 vdd.n858 8.92171
R6188 vdd.n929 vdd.n928 8.92171
R6189 vdd.n941 vdd.n940 8.92171
R6190 vdd.n966 vdd.n947 8.92171
R6191 vdd.n997 vdd.n994 8.92171
R6192 vdd.n4694 vdd.n4693 8.92171
R6193 vdd.n4724 vdd.n4723 8.92171
R6194 vdd.n4732 vdd.n4731 8.92171
R6195 vdd.n774 vdd.n768 8.92171
R6196 vdd.n4777 vdd.n4776 8.92171
R6197 vdd.n743 vdd.n726 8.92171
R6198 vdd.n4813 vdd.n4812 8.92171
R6199 vdd.n711 vdd.n706 8.92171
R6200 vdd.n4861 vdd.n4860 8.92171
R6201 vdd.n4869 vdd.n4868 8.92171
R6202 vdd.n4922 vdd.n4921 8.92171
R6203 vdd.n4952 vdd.n4951 8.92171
R6204 vdd.n4960 vdd.n4959 8.92171
R6205 vdd.n639 vdd.n633 8.92171
R6206 vdd.n5005 vdd.n5004 8.92171
R6207 vdd.n608 vdd.n591 8.92171
R6208 vdd.n5041 vdd.n5040 8.92171
R6209 vdd.n576 vdd.n571 8.92171
R6210 vdd.n5089 vdd.n5088 8.92171
R6211 vdd.n5097 vdd.n5096 8.92171
R6212 vdd.n5150 vdd.n5149 8.92171
R6213 vdd.n5180 vdd.n5179 8.92171
R6214 vdd.n5188 vdd.n5187 8.92171
R6215 vdd.n504 vdd.n498 8.92171
R6216 vdd.n5233 vdd.n5232 8.92171
R6217 vdd.n473 vdd.n456 8.92171
R6218 vdd.n5269 vdd.n5268 8.92171
R6219 vdd.n441 vdd.n436 8.92171
R6220 vdd.n5317 vdd.n5316 8.92171
R6221 vdd.n5325 vdd.n5324 8.92171
R6222 vdd.n5378 vdd.n5377 8.92171
R6223 vdd.n5408 vdd.n5407 8.92171
R6224 vdd.n5416 vdd.n5415 8.92171
R6225 vdd.n369 vdd.n363 8.92171
R6226 vdd.n5460 vdd.n5459 8.92171
R6227 vdd.n5484 vdd.n5483 8.92171
R6228 vdd.n5509 vdd.n318 8.92171
R6229 vdd.n319 vdd.n305 8.92171
R6230 vdd.n5542 vdd.n5541 8.92171
R6231 vdd.n288 vdd.n283 8.92171
R6232 vdd.n2176 vdd.n2175 8.85536
R6233 vdd.n2175 vdd.n2174 8.85536
R6234 vdd.n7319 vdd.n5812 8.77616
R6235 vdd.n7338 vdd.n5812 8.77616
R6236 vdd.n7357 vdd.n5812 8.77616
R6237 vdd.n7376 vdd.n5812 8.77616
R6238 vdd.n6514 vdd.n212 8.77616
R6239 vdd.n6551 vdd.n212 8.77616
R6240 vdd.n6585 vdd.n212 8.77616
R6241 vdd.n6741 vdd.n212 8.77616
R6242 vdd.n6778 vdd.n212 8.77616
R6243 vdd.n6812 vdd.n212 8.77616
R6244 vdd.n6968 vdd.n212 8.77616
R6245 vdd.n7005 vdd.n212 8.77616
R6246 vdd.n7039 vdd.n212 8.77616
R6247 vdd.n7195 vdd.n212 8.77616
R6248 vdd.n7232 vdd.n212 8.77616
R6249 vdd.n7266 vdd.n212 8.77616
R6250 vdd.n7179 vdd.n212 8.77616
R6251 vdd.n6952 vdd.n212 8.77616
R6252 vdd.n6725 vdd.n212 8.77616
R6253 vdd.n6498 vdd.n212 8.77616
R6254 vdd.n6374 vdd.n212 8.77616
R6255 vdd.n2953 vdd.n2065 8.77616
R6256 vdd.n2984 vdd.n2065 8.77616
R6257 vdd.n3181 vdd.n2065 8.77616
R6258 vdd.n3212 vdd.n2065 8.77616
R6259 vdd.n3409 vdd.n2065 8.77616
R6260 vdd.n3440 vdd.n2065 8.77616
R6261 vdd.n3637 vdd.n2065 8.77616
R6262 vdd.n3668 vdd.n2065 8.77616
R6263 vdd.n3761 vdd.n2065 8.77616
R6264 vdd.n3726 vdd.n2065 8.77616
R6265 vdd.n3524 vdd.n2065 8.77616
R6266 vdd.n3490 vdd.n2065 8.77616
R6267 vdd.n3581 vdd.n2065 8.77616
R6268 vdd.n3296 vdd.n2065 8.77616
R6269 vdd.n3262 vdd.n2065 8.77616
R6270 vdd.n3353 vdd.n2065 8.77616
R6271 vdd.n3068 vdd.n2065 8.77616
R6272 vdd.n3034 vdd.n2065 8.77616
R6273 vdd.n3125 vdd.n2065 8.77616
R6274 vdd.n4025 vdd.n2059 8.77616
R6275 vdd.n4025 vdd.n2062 8.77616
R6276 vdd.n4727 vdd.n250 8.77616
R6277 vdd.n4758 vdd.n250 8.77616
R6278 vdd.n4955 vdd.n250 8.77616
R6279 vdd.n4986 vdd.n250 8.77616
R6280 vdd.n5183 vdd.n250 8.77616
R6281 vdd.n5214 vdd.n250 8.77616
R6282 vdd.n5411 vdd.n250 8.77616
R6283 vdd.n5442 vdd.n250 8.77616
R6284 vdd.n5537 vdd.n250 8.77616
R6285 vdd.n5502 vdd.n250 8.77616
R6286 vdd.n5298 vdd.n250 8.77616
R6287 vdd.n5264 vdd.n250 8.77616
R6288 vdd.n5355 vdd.n250 8.77616
R6289 vdd.n5070 vdd.n250 8.77616
R6290 vdd.n5036 vdd.n250 8.77616
R6291 vdd.n5127 vdd.n250 8.77616
R6292 vdd.n4842 vdd.n250 8.77616
R6293 vdd.n4808 vdd.n250 8.77616
R6294 vdd.n4899 vdd.n250 8.77616
R6295 vdd.n5727 vdd.n258 8.77616
R6296 vdd.n5727 vdd.n252 8.77616
R6297 vdd.n5727 vdd.n256 8.77616
R6298 vdd.n5727 vdd.n254 8.77616
R6299 vdd.n7436 vdd.t79 8.57285
R6300 vdd.n4653 vdd.t89 8.57285
R6301 vdd.n4679 vdd.n798 8.45943
R6302 vdd.n2905 vdd.n2774 8.45943
R6303 vdd.n3800 vdd.n3799 8.4584
R6304 vdd.n5576 vdd.n5575 8.4584
R6305 vdd.n5575 vdd.n250 8.45416
R6306 vdd.n3799 vdd.n2065 8.45416
R6307 vdd.n2774 vdd.n2065 8.45226
R6308 vdd.n798 vdd.n250 8.45226
R6309 vdd.n2180 vdd.n2168 8.45089
R6310 vdd.n7483 vdd.t78 8.41977
R6311 vdd.t88 vdd.n4644 8.41977
R6312 vdd.n7483 vdd.n213 7.96054
R6313 vdd.n4644 vdd.n4642 7.96054
R6314 vdd.n2180 vdd.n2179 7.89809
R6315 vdd.n3977 vdd.n3976 7.84364
R6316 vdd.n56 vdd.t115 7.14336
R6317 vdd.n174 vdd.t128 7.14336
R6318 vdd.n2180 vdd.n2167 7.02351
R6319 vdd.n2136 vdd.n2101 6.94993
R6320 vdd.n2174 vdd.n2173 6.08327
R6321 vdd.n2183 vdd.n2182 5.81188
R6322 vdd.n12 vdd.t83 5.71479
R6323 vdd.n58 vdd.n55 5.67473
R6324 vdd.n7399 vdd.n5812 5.63319
R6325 vdd.n6337 vdd.n212 5.63319
R6326 vdd.n6604 vdd.n212 5.63319
R6327 vdd.n6553 vdd.n212 5.63319
R6328 vdd.n6517 vdd.n212 5.63319
R6329 vdd.n6204 vdd.n212 5.63319
R6330 vdd.n6831 vdd.n212 5.63319
R6331 vdd.n6780 vdd.n212 5.63319
R6332 vdd.n6744 vdd.n212 5.63319
R6333 vdd.n6071 vdd.n212 5.63319
R6334 vdd.n7058 vdd.n212 5.63319
R6335 vdd.n7007 vdd.n212 5.63319
R6336 vdd.n6971 vdd.n212 5.63319
R6337 vdd.n5938 vdd.n212 5.63319
R6338 vdd.n7234 vdd.n212 5.63319
R6339 vdd.n7198 vdd.n212 5.63319
R6340 vdd.n3763 vdd.n2065 5.63319
R6341 vdd.n3729 vdd.n2065 5.63319
R6342 vdd.n3666 vdd.n2065 5.63319
R6343 vdd.n3608 vdd.n2065 5.63319
R6344 vdd.n3545 vdd.n2065 5.63319
R6345 vdd.n3492 vdd.n2065 5.63319
R6346 vdd.n3438 vdd.n2065 5.63319
R6347 vdd.n3380 vdd.n2065 5.63319
R6348 vdd.n3317 vdd.n2065 5.63319
R6349 vdd.n3264 vdd.n2065 5.63319
R6350 vdd.n3210 vdd.n2065 5.63319
R6351 vdd.n3152 vdd.n2065 5.63319
R6352 vdd.n3089 vdd.n2065 5.63319
R6353 vdd.n3036 vdd.n2065 5.63319
R6354 vdd.n2982 vdd.n2065 5.63319
R6355 vdd.n2924 vdd.n2065 5.63319
R6356 vdd.n4026 vdd.n4025 5.63319
R6357 vdd.n4025 vdd.n2061 5.63319
R6358 vdd.n5539 vdd.n250 5.63319
R6359 vdd.n5505 vdd.n250 5.63319
R6360 vdd.n5440 vdd.n250 5.63319
R6361 vdd.n5382 vdd.n250 5.63319
R6362 vdd.n5319 vdd.n250 5.63319
R6363 vdd.n5266 vdd.n250 5.63319
R6364 vdd.n5212 vdd.n250 5.63319
R6365 vdd.n5154 vdd.n250 5.63319
R6366 vdd.n5091 vdd.n250 5.63319
R6367 vdd.n5038 vdd.n250 5.63319
R6368 vdd.n4984 vdd.n250 5.63319
R6369 vdd.n4926 vdd.n250 5.63319
R6370 vdd.n4863 vdd.n250 5.63319
R6371 vdd.n4810 vdd.n250 5.63319
R6372 vdd.n4756 vdd.n250 5.63319
R6373 vdd.n4698 vdd.n250 5.63319
R6374 vdd.n5727 vdd.n255 5.63319
R6375 vdd.n2207 vdd.n2103 5.27109
R6376 vdd.n6407 vdd.n212 5.1329
R6377 vdd.n7290 vdd.n212 5.1329
R6378 vdd.n4633 vdd 5.06361
R6379 vdd.t23 vdd 4.92533
R6380 vdd.n3979 vdd.n3978 4.90246
R6381 vdd.n29 vdd.n23 4.77029
R6382 vdd.t80 vdd.n213 4.74591
R6383 vdd.n4642 vdd.t90 4.74591
R6384 vdd.n192 vdd.n191 4.6505
R6385 vdd.n7490 vdd.n7489 4.6505
R6386 vdd.n2212 vdd.n2102 4.6505
R6387 vdd.n2206 vdd.n2205 4.6505
R6388 vdd.n2209 vdd.n2103 4.6505
R6389 vdd.n2213 vdd.n2100 4.6505
R6390 vdd.n2215 vdd.n2214 4.6505
R6391 vdd.n3984 vdd.n3983 4.6505
R6392 vdd.n3839 vdd.n3838 4.6505
R6393 vdd.n4626 vdd.n4625 4.6505
R6394 vdd.n4612 vdd.n4611 4.6505
R6395 vdd.n216 vdd.n215 4.6505
R6396 vdd.n5754 vdd.n241 4.6505
R6397 vdd.n47 vdd.n46 4.6505
R6398 vdd.n43 vdd.n42 4.6505
R6399 vdd.n37 vdd.n36 4.6505
R6400 vdd.n33 vdd.n32 4.6505
R6401 vdd.n29 vdd.n28 4.6505
R6402 vdd.n154 vdd.n153 4.6505
R6403 vdd.n133 vdd.n132 4.6505
R6404 vdd.n137 vdd.n136 4.6505
R6405 vdd.n59 vdd.n58 4.6505
R6406 vdd.n63 vdd.n62 4.6505
R6407 vdd.n74 vdd.n73 4.6505
R6408 vdd.n77 vdd.n76 4.6505
R6409 vdd.n88 vdd.n87 4.6505
R6410 vdd.n92 vdd.n91 4.6505
R6411 vdd.n105 vdd.n104 4.6505
R6412 vdd.n109 vdd.n108 4.6505
R6413 vdd.n113 vdd.n112 4.6505
R6414 vdd.n53 vdd.n52 4.6505
R6415 vdd.n158 vdd.n157 4.6505
R6416 vdd.n3836 vdd.n2065 4.59701
R6417 vdd.n6405 vdd.n6385 4.54027
R6418 vdd.n7293 vdd.n7292 4.54027
R6419 vdd.n4680 vdd.n4678 4.54027
R6420 vdd.n5578 vdd.n5577 4.54027
R6421 vdd.n2906 vdd.n2904 4.54027
R6422 vdd.n3802 vdd.n3801 4.54027
R6423 vdd.n4528 vdd.n4527 4.54027
R6424 vdd.n4049 vdd.n2022 4.54027
R6425 vdd.n2127 vdd.n2126 4.52882
R6426 vdd.n3898 vdd.n3897 4.52882
R6427 vdd.n835 vdd.n834 4.52882
R6428 vdd.n5770 vdd.n5769 4.52882
R6429 vdd.n210 vdd.n209 4.5005
R6430 vdd.n7499 vdd.n198 4.5005
R6431 vdd.n199 vdd.n197 4.5005
R6432 vdd.n6414 vdd.n6413 4.5005
R6433 vdd.n6435 vdd.n6434 4.5005
R6434 vdd.n6333 vdd.n6332 4.5005
R6435 vdd.n6341 vdd.n6325 4.5005
R6436 vdd.n6622 vdd.n6254 4.5005
R6437 vdd.n6266 vdd.n6259 4.5005
R6438 vdd.n6599 vdd.n6598 4.5005
R6439 vdd.n6578 vdd.n6577 4.5005
R6440 vdd.n6560 vdd.n6559 4.5005
R6441 vdd.n6543 vdd.n6542 4.5005
R6442 vdd.n6526 vdd.n6525 4.5005
R6443 vdd.n6311 vdd.n6309 4.5005
R6444 vdd.n6331 vdd.n6330 4.5005
R6445 vdd.n6562 vdd.n6561 4.5005
R6446 vdd.n6545 vdd.n6544 4.5005
R6447 vdd.n6272 vdd.n6271 4.5005
R6448 vdd.n6289 vdd.n6287 4.5005
R6449 vdd.n6200 vdd.n6199 4.5005
R6450 vdd.n6208 vdd.n6192 4.5005
R6451 vdd.n6849 vdd.n6121 4.5005
R6452 vdd.n6133 vdd.n6126 4.5005
R6453 vdd.n6826 vdd.n6825 4.5005
R6454 vdd.n6805 vdd.n6804 4.5005
R6455 vdd.n6787 vdd.n6786 4.5005
R6456 vdd.n6770 vdd.n6769 4.5005
R6457 vdd.n6753 vdd.n6752 4.5005
R6458 vdd.n6178 vdd.n6176 4.5005
R6459 vdd.n6198 vdd.n6197 4.5005
R6460 vdd.n6789 vdd.n6788 4.5005
R6461 vdd.n6772 vdd.n6771 4.5005
R6462 vdd.n6139 vdd.n6138 4.5005
R6463 vdd.n6156 vdd.n6154 4.5005
R6464 vdd.n6067 vdd.n6066 4.5005
R6465 vdd.n6075 vdd.n6059 4.5005
R6466 vdd.n7076 vdd.n5988 4.5005
R6467 vdd.n6000 vdd.n5993 4.5005
R6468 vdd.n7053 vdd.n7052 4.5005
R6469 vdd.n7032 vdd.n7031 4.5005
R6470 vdd.n7014 vdd.n7013 4.5005
R6471 vdd.n6997 vdd.n6996 4.5005
R6472 vdd.n6980 vdd.n6979 4.5005
R6473 vdd.n6045 vdd.n6043 4.5005
R6474 vdd.n6065 vdd.n6064 4.5005
R6475 vdd.n7016 vdd.n7015 4.5005
R6476 vdd.n6999 vdd.n6998 4.5005
R6477 vdd.n6006 vdd.n6005 4.5005
R6478 vdd.n6023 vdd.n6021 4.5005
R6479 vdd.n5934 vdd.n5933 4.5005
R6480 vdd.n5942 vdd.n5926 4.5005
R6481 vdd.n7285 vdd.n7284 4.5005
R6482 vdd.n7259 vdd.n7258 4.5005
R6483 vdd.n7241 vdd.n7240 4.5005
R6484 vdd.n7224 vdd.n7223 4.5005
R6485 vdd.n7207 vdd.n7206 4.5005
R6486 vdd.n5912 vdd.n5910 4.5005
R6487 vdd.n5932 vdd.n5931 4.5005
R6488 vdd.n7243 vdd.n7242 4.5005
R6489 vdd.n7226 vdd.n7225 4.5005
R6490 vdd.n5872 vdd.n5871 4.5005
R6491 vdd.n5890 vdd.n5888 4.5005
R6492 vdd.n7096 vdd.n5977 4.5005
R6493 vdd.n7173 vdd.n7172 4.5005
R6494 vdd.n5953 vdd.n5947 4.5005
R6495 vdd.n7153 vdd.n7152 4.5005
R6496 vdd.n5967 vdd.n5958 4.5005
R6497 vdd.n7131 vdd.n7130 4.5005
R6498 vdd.n7118 vdd.n5963 4.5005
R6499 vdd.n7116 vdd.n7115 4.5005
R6500 vdd.n7095 vdd.n7094 4.5005
R6501 vdd.n6869 vdd.n6110 4.5005
R6502 vdd.n6946 vdd.n6945 4.5005
R6503 vdd.n6086 vdd.n6080 4.5005
R6504 vdd.n6926 vdd.n6925 4.5005
R6505 vdd.n6100 vdd.n6091 4.5005
R6506 vdd.n6904 vdd.n6903 4.5005
R6507 vdd.n6891 vdd.n6096 4.5005
R6508 vdd.n6889 vdd.n6888 4.5005
R6509 vdd.n6868 vdd.n6867 4.5005
R6510 vdd.n6642 vdd.n6243 4.5005
R6511 vdd.n6719 vdd.n6718 4.5005
R6512 vdd.n6219 vdd.n6213 4.5005
R6513 vdd.n6699 vdd.n6698 4.5005
R6514 vdd.n6233 vdd.n6224 4.5005
R6515 vdd.n6677 vdd.n6676 4.5005
R6516 vdd.n6664 vdd.n6229 4.5005
R6517 vdd.n6662 vdd.n6661 4.5005
R6518 vdd.n6641 vdd.n6640 4.5005
R6519 vdd.n6437 vdd.n6362 4.5005
R6520 vdd.n6492 vdd.n6491 4.5005
R6521 vdd.n6352 vdd.n6346 4.5005
R6522 vdd.n6472 vdd.n6471 4.5005
R6523 vdd.n6366 vdd.n6357 4.5005
R6524 vdd.n6450 vdd.n6449 4.5005
R6525 vdd.n6415 vdd.n6376 4.5005
R6526 vdd.n6383 vdd.n6382 4.5005
R6527 vdd.n6384 vdd.n6383 4.5005
R6528 vdd.n6265 vdd.n6263 4.5005
R6529 vdd.n6267 vdd.n6265 4.5005
R6530 vdd.n6558 vdd.n6283 4.5005
R6531 vdd.n6283 vdd.n6282 4.5005
R6532 vdd.n6312 vdd.n6310 4.5005
R6533 vdd.n6522 vdd.n6312 4.5005
R6534 vdd.n6319 vdd.n6318 4.5005
R6535 vdd.n6318 vdd.n6317 4.5005
R6536 vdd.n6547 vdd.n6546 4.5005
R6537 vdd.n6548 vdd.n6547 4.5005
R6538 vdd.n6278 vdd.n6276 4.5005
R6539 vdd.n6279 vdd.n6278 4.5005
R6540 vdd.n6132 vdd.n6130 4.5005
R6541 vdd.n6134 vdd.n6132 4.5005
R6542 vdd.n6785 vdd.n6150 4.5005
R6543 vdd.n6150 vdd.n6149 4.5005
R6544 vdd.n6179 vdd.n6177 4.5005
R6545 vdd.n6749 vdd.n6179 4.5005
R6546 vdd.n6186 vdd.n6185 4.5005
R6547 vdd.n6185 vdd.n6184 4.5005
R6548 vdd.n6774 vdd.n6773 4.5005
R6549 vdd.n6775 vdd.n6774 4.5005
R6550 vdd.n6145 vdd.n6143 4.5005
R6551 vdd.n6146 vdd.n6145 4.5005
R6552 vdd.n5999 vdd.n5997 4.5005
R6553 vdd.n6001 vdd.n5999 4.5005
R6554 vdd.n7012 vdd.n6017 4.5005
R6555 vdd.n6017 vdd.n6016 4.5005
R6556 vdd.n6046 vdd.n6044 4.5005
R6557 vdd.n6976 vdd.n6046 4.5005
R6558 vdd.n6053 vdd.n6052 4.5005
R6559 vdd.n6052 vdd.n6051 4.5005
R6560 vdd.n7001 vdd.n7000 4.5005
R6561 vdd.n7002 vdd.n7001 4.5005
R6562 vdd.n6012 vdd.n6010 4.5005
R6563 vdd.n6013 vdd.n6012 4.5005
R6564 vdd.n7239 vdd.n5884 4.5005
R6565 vdd.n5884 vdd.n5883 4.5005
R6566 vdd.n5913 vdd.n5911 4.5005
R6567 vdd.n7203 vdd.n5913 4.5005
R6568 vdd.n5920 vdd.n5919 4.5005
R6569 vdd.n5919 vdd.n5918 4.5005
R6570 vdd.n7228 vdd.n7227 4.5005
R6571 vdd.n7229 vdd.n7228 4.5005
R6572 vdd.n5879 vdd.n5877 4.5005
R6573 vdd.n5880 vdd.n5879 4.5005
R6574 vdd.n7283 vdd.n5866 4.5005
R6575 vdd.n5868 vdd.n5866 4.5005
R6576 vdd.n5941 vdd.n5940 4.5005
R6577 vdd.n5940 vdd.n5939 4.5005
R6578 vdd.n5952 vdd.n5951 4.5005
R6579 vdd.n5951 vdd.n5950 4.5005
R6580 vdd.n7133 vdd.n7132 4.5005
R6581 vdd.n7133 vdd.n5962 4.5005
R6582 vdd.n5973 vdd.n5972 4.5005
R6583 vdd.n5974 vdd.n5973 4.5005
R6584 vdd.n5927 vdd.n5925 4.5005
R6585 vdd.n5937 vdd.n5927 4.5005
R6586 vdd.n5984 vdd.n5983 4.5005
R6587 vdd.n5985 vdd.n5984 4.5005
R6588 vdd.n6074 vdd.n6073 4.5005
R6589 vdd.n6073 vdd.n6072 4.5005
R6590 vdd.n6085 vdd.n6084 4.5005
R6591 vdd.n6084 vdd.n6083 4.5005
R6592 vdd.n6906 vdd.n6905 4.5005
R6593 vdd.n6906 vdd.n6095 4.5005
R6594 vdd.n6106 vdd.n6105 4.5005
R6595 vdd.n6107 vdd.n6106 4.5005
R6596 vdd.n6060 vdd.n6058 4.5005
R6597 vdd.n6070 vdd.n6060 4.5005
R6598 vdd.n6117 vdd.n6116 4.5005
R6599 vdd.n6118 vdd.n6117 4.5005
R6600 vdd.n6207 vdd.n6206 4.5005
R6601 vdd.n6206 vdd.n6205 4.5005
R6602 vdd.n6218 vdd.n6217 4.5005
R6603 vdd.n6217 vdd.n6216 4.5005
R6604 vdd.n6679 vdd.n6678 4.5005
R6605 vdd.n6679 vdd.n6228 4.5005
R6606 vdd.n6239 vdd.n6238 4.5005
R6607 vdd.n6240 vdd.n6239 4.5005
R6608 vdd.n6193 vdd.n6191 4.5005
R6609 vdd.n6203 vdd.n6193 4.5005
R6610 vdd.n6250 vdd.n6249 4.5005
R6611 vdd.n6251 vdd.n6250 4.5005
R6612 vdd.n6340 vdd.n6339 4.5005
R6613 vdd.n6339 vdd.n6338 4.5005
R6614 vdd.n6351 vdd.n6350 4.5005
R6615 vdd.n6350 vdd.n6349 4.5005
R6616 vdd.n6452 vdd.n6451 4.5005
R6617 vdd.n6452 vdd.n6361 4.5005
R6618 vdd.n6326 vdd.n6324 4.5005
R6619 vdd.n6336 vdd.n6326 4.5005
R6620 vdd.n6372 vdd.n6371 4.5005
R6621 vdd.n6373 vdd.n6372 4.5005
R6622 vdd.n7394 vdd.n7393 4.5005
R6623 vdd.n7405 vdd.n5791 4.5005
R6624 vdd.n5861 vdd.n5860 4.5005
R6625 vdd.n5850 vdd.n5849 4.5005
R6626 vdd.n7314 vdd.n7313 4.5005
R6627 vdd.n5839 vdd.n5838 4.5005
R6628 vdd.n7333 vdd.n7332 4.5005
R6629 vdd.n5828 vdd.n5827 4.5005
R6630 vdd.n7352 vdd.n7351 4.5005
R6631 vdd.n5816 vdd.n5815 4.5005
R6632 vdd.n7371 vdd.n7370 4.5005
R6633 vdd.n5798 vdd.n5796 4.5005
R6634 vdd.n5799 vdd.n5798 4.5005
R6635 vdd.n5856 vdd.n5854 4.5005
R6636 vdd.n5857 vdd.n5856 4.5005
R6637 vdd.n5845 vdd.n5843 4.5005
R6638 vdd.n5846 vdd.n5845 4.5005
R6639 vdd.n5834 vdd.n5832 4.5005
R6640 vdd.n5835 vdd.n5834 4.5005
R6641 vdd.n5823 vdd.n5821 4.5005
R6642 vdd.n5824 vdd.n5823 4.5005
R6643 vdd.n5590 vdd.n5589 4.5005
R6644 vdd.n5588 vdd.n266 4.5005
R6645 vdd.n266 vdd.n263 4.5005
R6646 vdd.n5718 vdd.n5717 4.5005
R6647 vdd.n5592 vdd.n5591 4.5005
R6648 vdd.n5652 vdd.n246 4.5005
R6649 vdd.n5672 vdd.n5671 4.5005
R6650 vdd.n5627 vdd.n5625 4.5005
R6651 vdd.n5693 vdd.n5692 4.5005
R6652 vdd.n5693 vdd.n5624 4.5005
R6653 vdd.n5642 vdd.n5641 4.5005
R6654 vdd.n5705 vdd.n5704 4.5005
R6655 vdd.n5703 vdd.n5702 4.5005
R6656 vdd.n5702 vdd.n5701 4.5005
R6657 vdd.n5707 vdd.n5706 4.5005
R6658 vdd.n270 vdd.n268 4.5005
R6659 vdd.n5616 vdd.n5615 4.5005
R6660 vdd.n5617 vdd.n5616 4.5005
R6661 vdd.n5675 vdd.n5674 4.5005
R6662 vdd.n5664 vdd.n5651 4.5005
R6663 vdd.n5678 vdd.n5664 4.5005
R6664 vdd.n2198 vdd.n2197 4.5005
R6665 vdd.n2195 vdd.n2189 4.5005
R6666 vdd.n2208 vdd.n2106 4.5005
R6667 vdd.n2208 vdd.n2207 4.5005
R6668 vdd.n2156 vdd.n2107 4.5005
R6669 vdd.n2136 vdd.n2134 4.5005
R6670 vdd.n2135 vdd.n2099 4.5005
R6671 vdd.n2778 vdd.n2772 4.5005
R6672 vdd.n2765 vdd.n2763 4.5005
R6673 vdd.n2763 vdd.n2762 4.5005
R6674 vdd.n2947 vdd.n2946 4.5005
R6675 vdd.n2917 vdd.n2916 4.5005
R6676 vdd.n2730 vdd.n2729 4.5005
R6677 vdd.n2728 vdd.n2717 4.5005
R6678 vdd.n3026 vdd.n3025 4.5005
R6679 vdd.n3121 vdd.n3120 4.5005
R6680 vdd.n2655 vdd.n2648 4.5005
R6681 vdd.n3145 vdd.n3144 4.5005
R6682 vdd.n2595 vdd.n2594 4.5005
R6683 vdd.n2593 vdd.n2582 4.5005
R6684 vdd.n3254 vdd.n3253 4.5005
R6685 vdd.n3349 vdd.n3348 4.5005
R6686 vdd.n2520 vdd.n2513 4.5005
R6687 vdd.n3373 vdd.n3372 4.5005
R6688 vdd.n2460 vdd.n2459 4.5005
R6689 vdd.n2458 vdd.n2447 4.5005
R6690 vdd.n3482 vdd.n3481 4.5005
R6691 vdd.n3577 vdd.n3576 4.5005
R6692 vdd.n2385 vdd.n2378 4.5005
R6693 vdd.n3601 vdd.n3600 4.5005
R6694 vdd.n2325 vdd.n2324 4.5005
R6695 vdd.n2323 vdd.n2322 4.5005
R6696 vdd.n2307 vdd.n2306 4.5005
R6697 vdd.n3792 vdd.n3791 4.5005
R6698 vdd.n3770 vdd.n3769 4.5005
R6699 vdd.n3768 vdd.n2260 4.5005
R6700 vdd.n2260 vdd.n2259 4.5005
R6701 vdd.n3772 vdd.n3771 4.5005
R6702 vdd.n3755 vdd.n3754 4.5005
R6703 vdd.n3757 vdd.n3756 4.5005
R6704 vdd.n3758 vdd.n3757 4.5005
R6705 vdd.n3753 vdd.n3752 4.5005
R6706 vdd.n3736 vdd.n3735 4.5005
R6707 vdd.n2291 vdd.n2289 4.5005
R6708 vdd.n3732 vdd.n2291 4.5005
R6709 vdd.n2290 vdd.n2288 4.5005
R6710 vdd.n3712 vdd.n3711 4.5005
R6711 vdd.n2301 vdd.n2300 4.5005
R6712 vdd.n2300 vdd.n2299 4.5005
R6713 vdd.n2267 vdd.n2264 4.5005
R6714 vdd.n2266 vdd.n2254 4.5005
R6715 vdd.n2256 vdd.n2254 4.5005
R6716 vdd.n2310 vdd.n2309 4.5005
R6717 vdd.n2309 vdd.n2308 4.5005
R6718 vdd.n3683 vdd.n3682 4.5005
R6719 vdd.n2347 vdd.n2338 4.5005
R6720 vdd.n2332 vdd.n2331 4.5005
R6721 vdd.n2331 vdd.n2330 4.5005
R6722 vdd.n3660 vdd.n3659 4.5005
R6723 vdd.n3647 vdd.n2343 4.5005
R6724 vdd.n3662 vdd.n3661 4.5005
R6725 vdd.n3662 vdd.n2342 4.5005
R6726 vdd.n3645 vdd.n3644 4.5005
R6727 vdd.n2361 vdd.n2359 4.5005
R6728 vdd.n2353 vdd.n2352 4.5005
R6729 vdd.n2354 vdd.n2353 4.5005
R6730 vdd.n3631 vdd.n3630 4.5005
R6731 vdd.n2373 vdd.n2367 4.5005
R6732 vdd.n2360 vdd.n2358 4.5005
R6733 vdd.n2358 vdd.n2357 4.5005
R6734 vdd.n2333 vdd.n2317 4.5005
R6735 vdd.n2318 vdd.n2316 4.5005
R6736 vdd.n2328 vdd.n2318 4.5005
R6737 vdd.n2372 vdd.n2371 4.5005
R6738 vdd.n2371 vdd.n2370 4.5005
R6739 vdd.n3557 vdd.n3556 4.5005
R6740 vdd.n3538 vdd.n2400 4.5005
R6741 vdd.n3540 vdd.n3539 4.5005
R6742 vdd.n3540 vdd.n2399 4.5005
R6743 vdd.n2410 vdd.n2401 4.5005
R6744 vdd.n2421 vdd.n2419 4.5005
R6745 vdd.n2409 vdd.n2407 4.5005
R6746 vdd.n2411 vdd.n2409 4.5005
R6747 vdd.n3517 vdd.n3516 4.5005
R6748 vdd.n3499 vdd.n3498 4.5005
R6749 vdd.n3497 vdd.n2415 4.5005
R6750 vdd.n2415 vdd.n2414 4.5005
R6751 vdd.n3501 vdd.n3500 4.5005
R6752 vdd.n3484 vdd.n3483 4.5005
R6753 vdd.n3486 vdd.n3485 4.5005
R6754 vdd.n3487 vdd.n3486 4.5005
R6755 vdd.n3555 vdd.n3554 4.5005
R6756 vdd.n3553 vdd.n2382 4.5005
R6757 vdd.n2382 vdd.n2381 4.5005
R6758 vdd.n2457 vdd.n2456 4.5005
R6759 vdd.n2456 vdd.n2455 4.5005
R6760 vdd.n3456 vdd.n3455 4.5005
R6761 vdd.n2482 vdd.n2473 4.5005
R6762 vdd.n2467 vdd.n2466 4.5005
R6763 vdd.n2466 vdd.n2465 4.5005
R6764 vdd.n3432 vdd.n3431 4.5005
R6765 vdd.n3419 vdd.n2478 4.5005
R6766 vdd.n3434 vdd.n3433 4.5005
R6767 vdd.n3434 vdd.n2477 4.5005
R6768 vdd.n3417 vdd.n3416 4.5005
R6769 vdd.n2496 vdd.n2494 4.5005
R6770 vdd.n2488 vdd.n2487 4.5005
R6771 vdd.n2489 vdd.n2488 4.5005
R6772 vdd.n3403 vdd.n3402 4.5005
R6773 vdd.n2508 vdd.n2502 4.5005
R6774 vdd.n2495 vdd.n2493 4.5005
R6775 vdd.n2493 vdd.n2492 4.5005
R6776 vdd.n2468 vdd.n2443 4.5005
R6777 vdd.n2444 vdd.n2442 4.5005
R6778 vdd.n2463 vdd.n2444 4.5005
R6779 vdd.n2507 vdd.n2506 4.5005
R6780 vdd.n2506 vdd.n2505 4.5005
R6781 vdd.n3329 vdd.n3328 4.5005
R6782 vdd.n3310 vdd.n2535 4.5005
R6783 vdd.n3312 vdd.n3311 4.5005
R6784 vdd.n3312 vdd.n2534 4.5005
R6785 vdd.n2545 vdd.n2536 4.5005
R6786 vdd.n2556 vdd.n2554 4.5005
R6787 vdd.n2544 vdd.n2542 4.5005
R6788 vdd.n2546 vdd.n2544 4.5005
R6789 vdd.n3289 vdd.n3288 4.5005
R6790 vdd.n3271 vdd.n3270 4.5005
R6791 vdd.n3269 vdd.n2550 4.5005
R6792 vdd.n2550 vdd.n2549 4.5005
R6793 vdd.n3273 vdd.n3272 4.5005
R6794 vdd.n3256 vdd.n3255 4.5005
R6795 vdd.n3258 vdd.n3257 4.5005
R6796 vdd.n3259 vdd.n3258 4.5005
R6797 vdd.n3327 vdd.n3326 4.5005
R6798 vdd.n3325 vdd.n2517 4.5005
R6799 vdd.n2517 vdd.n2516 4.5005
R6800 vdd.n2592 vdd.n2591 4.5005
R6801 vdd.n2591 vdd.n2590 4.5005
R6802 vdd.n3228 vdd.n3227 4.5005
R6803 vdd.n2617 vdd.n2608 4.5005
R6804 vdd.n2602 vdd.n2601 4.5005
R6805 vdd.n2601 vdd.n2600 4.5005
R6806 vdd.n3204 vdd.n3203 4.5005
R6807 vdd.n3191 vdd.n2613 4.5005
R6808 vdd.n3206 vdd.n3205 4.5005
R6809 vdd.n3206 vdd.n2612 4.5005
R6810 vdd.n3189 vdd.n3188 4.5005
R6811 vdd.n2631 vdd.n2629 4.5005
R6812 vdd.n2623 vdd.n2622 4.5005
R6813 vdd.n2624 vdd.n2623 4.5005
R6814 vdd.n3175 vdd.n3174 4.5005
R6815 vdd.n2643 vdd.n2637 4.5005
R6816 vdd.n2630 vdd.n2628 4.5005
R6817 vdd.n2628 vdd.n2627 4.5005
R6818 vdd.n2603 vdd.n2578 4.5005
R6819 vdd.n2579 vdd.n2577 4.5005
R6820 vdd.n2598 vdd.n2579 4.5005
R6821 vdd.n2642 vdd.n2641 4.5005
R6822 vdd.n2641 vdd.n2640 4.5005
R6823 vdd.n3101 vdd.n3100 4.5005
R6824 vdd.n3082 vdd.n2670 4.5005
R6825 vdd.n3084 vdd.n3083 4.5005
R6826 vdd.n3084 vdd.n2669 4.5005
R6827 vdd.n2680 vdd.n2671 4.5005
R6828 vdd.n2691 vdd.n2689 4.5005
R6829 vdd.n2679 vdd.n2677 4.5005
R6830 vdd.n2681 vdd.n2679 4.5005
R6831 vdd.n3061 vdd.n3060 4.5005
R6832 vdd.n3043 vdd.n3042 4.5005
R6833 vdd.n3041 vdd.n2685 4.5005
R6834 vdd.n2685 vdd.n2684 4.5005
R6835 vdd.n3045 vdd.n3044 4.5005
R6836 vdd.n3028 vdd.n3027 4.5005
R6837 vdd.n3030 vdd.n3029 4.5005
R6838 vdd.n3031 vdd.n3030 4.5005
R6839 vdd.n3099 vdd.n3098 4.5005
R6840 vdd.n3097 vdd.n2652 4.5005
R6841 vdd.n2652 vdd.n2651 4.5005
R6842 vdd.n2727 vdd.n2726 4.5005
R6843 vdd.n2726 vdd.n2725 4.5005
R6844 vdd.n3000 vdd.n2999 4.5005
R6845 vdd.n2752 vdd.n2743 4.5005
R6846 vdd.n2737 vdd.n2736 4.5005
R6847 vdd.n2736 vdd.n2735 4.5005
R6848 vdd.n2976 vdd.n2975 4.5005
R6849 vdd.n2963 vdd.n2748 4.5005
R6850 vdd.n2978 vdd.n2977 4.5005
R6851 vdd.n2978 vdd.n2747 4.5005
R6852 vdd.n2961 vdd.n2960 4.5005
R6853 vdd.n2766 vdd.n2764 4.5005
R6854 vdd.n2758 vdd.n2757 4.5005
R6855 vdd.n2759 vdd.n2758 4.5005
R6856 vdd.n2738 vdd.n2713 4.5005
R6857 vdd.n2714 vdd.n2712 4.5005
R6858 vdd.n2733 vdd.n2714 4.5005
R6859 vdd.n2777 vdd.n2776 4.5005
R6860 vdd.n2776 vdd.n2775 4.5005
R6861 vdd.n2895 vdd.n2894 4.5005
R6862 vdd.n2788 vdd.n2787 4.5005
R6863 vdd.n2799 vdd.n2794 4.5005
R6864 vdd.n2795 vdd.n2793 4.5005
R6865 vdd.n2875 vdd.n2795 4.5005
R6866 vdd.n2868 vdd.n2867 4.5005
R6867 vdd.n2812 vdd.n2804 4.5005
R6868 vdd.n2798 vdd.n2797 4.5005
R6869 vdd.n2797 vdd.n2796 4.5005
R6870 vdd.n2845 vdd.n2844 4.5005
R6871 vdd.n2832 vdd.n2809 4.5005
R6872 vdd.n2847 vdd.n2846 4.5005
R6873 vdd.n2847 vdd.n2808 4.5005
R6874 vdd.n2830 vdd.n2829 4.5005
R6875 vdd.n4031 vdd.n4030 4.5005
R6876 vdd.n2825 vdd.n2053 4.5005
R6877 vdd.n2055 vdd.n2053 4.5005
R6878 vdd.n2051 vdd.n2049 4.5005
R6879 vdd.n4012 vdd.n2040 4.5005
R6880 vdd.n4019 vdd.n4018 4.5005
R6881 vdd.n4019 vdd.n4009 4.5005
R6882 vdd.n1029 vdd.n1008 4.5005
R6883 vdd.n4517 vdd.n4516 4.5005
R6884 vdd.n4517 vdd.n1007 4.5005
R6885 vdd.n4515 vdd.n4514 4.5005
R6886 vdd.n1027 vdd.n1026 4.5005
R6887 vdd.n1134 vdd.n1133 4.5005
R6888 vdd.n1132 vdd.n1129 4.5005
R6889 vdd.n1154 vdd.n1116 4.5005
R6890 vdd.n1254 vdd.n1253 4.5005
R6891 vdd.n1255 vdd.n1248 4.5005
R6892 vdd.n1291 vdd.n1290 4.5005
R6893 vdd.n1398 vdd.n1397 4.5005
R6894 vdd.n1396 vdd.n1393 4.5005
R6895 vdd.n1418 vdd.n1380 4.5005
R6896 vdd.n1518 vdd.n1517 4.5005
R6897 vdd.n1519 vdd.n1512 4.5005
R6898 vdd.n1555 vdd.n1554 4.5005
R6899 vdd.n1662 vdd.n1661 4.5005
R6900 vdd.n1660 vdd.n1657 4.5005
R6901 vdd.n1682 vdd.n1644 4.5005
R6902 vdd.n1782 vdd.n1781 4.5005
R6903 vdd.n1783 vdd.n1776 4.5005
R6904 vdd.n1819 vdd.n1818 4.5005
R6905 vdd.n1926 vdd.n1925 4.5005
R6906 vdd.n1924 vdd.n1921 4.5005
R6907 vdd.n1946 vdd.n1908 4.5005
R6908 vdd.n2030 vdd.n2000 4.5005
R6909 vdd.n2010 vdd.n2009 4.5005
R6910 vdd.n1999 vdd.n1997 4.5005
R6911 vdd.n2001 vdd.n1999 4.5005
R6912 vdd.n2007 vdd.n2006 4.5005
R6913 vdd.n1981 vdd.n1979 4.5005
R6914 vdd.n4080 vdd.n4079 4.5005
R6915 vdd.n4080 vdd.n1978 4.5005
R6916 vdd.n1988 vdd.n1958 4.5005
R6917 vdd.n1968 vdd.n1967 4.5005
R6918 vdd.n1957 vdd.n1955 4.5005
R6919 vdd.n1959 vdd.n1957 4.5005
R6920 vdd.n1965 vdd.n1964 4.5005
R6921 vdd.n1939 vdd.n1937 4.5005
R6922 vdd.n4102 vdd.n4101 4.5005
R6923 vdd.n4102 vdd.n1936 4.5005
R6924 vdd.n2023 vdd.n2021 4.5005
R6925 vdd.n4058 vdd.n4057 4.5005
R6926 vdd.n4058 vdd.n2020 4.5005
R6927 vdd.n1907 vdd.n1905 4.5005
R6928 vdd.n1909 vdd.n1907 4.5005
R6929 vdd.n4125 vdd.n4124 4.5005
R6930 vdd.n1890 vdd.n1868 4.5005
R6931 vdd.n4127 vdd.n4126 4.5005
R6932 vdd.n4127 vdd.n1867 4.5005
R6933 vdd.n1888 vdd.n1887 4.5005
R6934 vdd.n4139 vdd.n4138 4.5005
R6935 vdd.n1884 vdd.n1840 4.5005
R6936 vdd.n1842 vdd.n1840 4.5005
R6937 vdd.n1838 vdd.n1836 4.5005
R6938 vdd.n4150 vdd.n4149 4.5005
R6939 vdd.n1857 vdd.n1856 4.5005
R6940 vdd.n1857 vdd.n1855 4.5005
R6941 vdd.n4152 vdd.n4151 4.5005
R6942 vdd.n1821 vdd.n1804 4.5005
R6943 vdd.n4154 vdd.n4153 4.5005
R6944 vdd.n4154 vdd.n1803 4.5005
R6945 vdd.n4123 vdd.n4122 4.5005
R6946 vdd.n1928 vdd.n1927 4.5005
R6947 vdd.n1929 vdd.n1928 4.5005
R6948 vdd.n1784 vdd.n1777 4.5005
R6949 vdd.n1786 vdd.n1784 4.5005
R6950 vdd.n1766 vdd.n1736 4.5005
R6951 vdd.n1746 vdd.n1745 4.5005
R6952 vdd.n1735 vdd.n1733 4.5005
R6953 vdd.n1737 vdd.n1735 4.5005
R6954 vdd.n1743 vdd.n1742 4.5005
R6955 vdd.n1717 vdd.n1715 4.5005
R6956 vdd.n4201 vdd.n4200 4.5005
R6957 vdd.n4201 vdd.n1714 4.5005
R6958 vdd.n1724 vdd.n1694 4.5005
R6959 vdd.n1704 vdd.n1703 4.5005
R6960 vdd.n1693 vdd.n1691 4.5005
R6961 vdd.n1695 vdd.n1693 4.5005
R6962 vdd.n1701 vdd.n1700 4.5005
R6963 vdd.n1675 vdd.n1673 4.5005
R6964 vdd.n4223 vdd.n4222 4.5005
R6965 vdd.n4223 vdd.n1672 4.5005
R6966 vdd.n1759 vdd.n1757 4.5005
R6967 vdd.n4179 vdd.n4178 4.5005
R6968 vdd.n4179 vdd.n1756 4.5005
R6969 vdd.n1643 vdd.n1641 4.5005
R6970 vdd.n1645 vdd.n1643 4.5005
R6971 vdd.n4246 vdd.n4245 4.5005
R6972 vdd.n1626 vdd.n1604 4.5005
R6973 vdd.n4248 vdd.n4247 4.5005
R6974 vdd.n4248 vdd.n1603 4.5005
R6975 vdd.n1624 vdd.n1623 4.5005
R6976 vdd.n4260 vdd.n4259 4.5005
R6977 vdd.n1620 vdd.n1576 4.5005
R6978 vdd.n1578 vdd.n1576 4.5005
R6979 vdd.n1574 vdd.n1572 4.5005
R6980 vdd.n4271 vdd.n4270 4.5005
R6981 vdd.n1593 vdd.n1592 4.5005
R6982 vdd.n1593 vdd.n1591 4.5005
R6983 vdd.n4273 vdd.n4272 4.5005
R6984 vdd.n1557 vdd.n1540 4.5005
R6985 vdd.n4275 vdd.n4274 4.5005
R6986 vdd.n4275 vdd.n1539 4.5005
R6987 vdd.n4244 vdd.n4243 4.5005
R6988 vdd.n1664 vdd.n1663 4.5005
R6989 vdd.n1665 vdd.n1664 4.5005
R6990 vdd.n1520 vdd.n1513 4.5005
R6991 vdd.n1522 vdd.n1520 4.5005
R6992 vdd.n1502 vdd.n1472 4.5005
R6993 vdd.n1482 vdd.n1481 4.5005
R6994 vdd.n1471 vdd.n1469 4.5005
R6995 vdd.n1473 vdd.n1471 4.5005
R6996 vdd.n1479 vdd.n1478 4.5005
R6997 vdd.n1453 vdd.n1451 4.5005
R6998 vdd.n4322 vdd.n4321 4.5005
R6999 vdd.n4322 vdd.n1450 4.5005
R7000 vdd.n1460 vdd.n1430 4.5005
R7001 vdd.n1440 vdd.n1439 4.5005
R7002 vdd.n1429 vdd.n1427 4.5005
R7003 vdd.n1431 vdd.n1429 4.5005
R7004 vdd.n1437 vdd.n1436 4.5005
R7005 vdd.n1411 vdd.n1409 4.5005
R7006 vdd.n4344 vdd.n4343 4.5005
R7007 vdd.n4344 vdd.n1408 4.5005
R7008 vdd.n1495 vdd.n1493 4.5005
R7009 vdd.n4300 vdd.n4299 4.5005
R7010 vdd.n4300 vdd.n1492 4.5005
R7011 vdd.n1379 vdd.n1377 4.5005
R7012 vdd.n1381 vdd.n1379 4.5005
R7013 vdd.n4367 vdd.n4366 4.5005
R7014 vdd.n1362 vdd.n1340 4.5005
R7015 vdd.n4369 vdd.n4368 4.5005
R7016 vdd.n4369 vdd.n1339 4.5005
R7017 vdd.n1360 vdd.n1359 4.5005
R7018 vdd.n4381 vdd.n4380 4.5005
R7019 vdd.n1356 vdd.n1312 4.5005
R7020 vdd.n1314 vdd.n1312 4.5005
R7021 vdd.n1310 vdd.n1308 4.5005
R7022 vdd.n4392 vdd.n4391 4.5005
R7023 vdd.n1329 vdd.n1328 4.5005
R7024 vdd.n1329 vdd.n1327 4.5005
R7025 vdd.n4394 vdd.n4393 4.5005
R7026 vdd.n1293 vdd.n1276 4.5005
R7027 vdd.n4396 vdd.n4395 4.5005
R7028 vdd.n4396 vdd.n1275 4.5005
R7029 vdd.n4365 vdd.n4364 4.5005
R7030 vdd.n1400 vdd.n1399 4.5005
R7031 vdd.n1401 vdd.n1400 4.5005
R7032 vdd.n1256 vdd.n1249 4.5005
R7033 vdd.n1258 vdd.n1256 4.5005
R7034 vdd.n1238 vdd.n1208 4.5005
R7035 vdd.n1218 vdd.n1217 4.5005
R7036 vdd.n1207 vdd.n1205 4.5005
R7037 vdd.n1209 vdd.n1207 4.5005
R7038 vdd.n1215 vdd.n1214 4.5005
R7039 vdd.n1189 vdd.n1187 4.5005
R7040 vdd.n4443 vdd.n4442 4.5005
R7041 vdd.n4443 vdd.n1186 4.5005
R7042 vdd.n1196 vdd.n1166 4.5005
R7043 vdd.n1176 vdd.n1175 4.5005
R7044 vdd.n1165 vdd.n1163 4.5005
R7045 vdd.n1167 vdd.n1165 4.5005
R7046 vdd.n1173 vdd.n1172 4.5005
R7047 vdd.n1147 vdd.n1145 4.5005
R7048 vdd.n4465 vdd.n4464 4.5005
R7049 vdd.n4465 vdd.n1144 4.5005
R7050 vdd.n1231 vdd.n1229 4.5005
R7051 vdd.n4421 vdd.n4420 4.5005
R7052 vdd.n4421 vdd.n1228 4.5005
R7053 vdd.n1115 vdd.n1113 4.5005
R7054 vdd.n1117 vdd.n1115 4.5005
R7055 vdd.n4488 vdd.n4487 4.5005
R7056 vdd.n1098 vdd.n1076 4.5005
R7057 vdd.n4490 vdd.n4489 4.5005
R7058 vdd.n4490 vdd.n1075 4.5005
R7059 vdd.n1096 vdd.n1095 4.5005
R7060 vdd.n4502 vdd.n4501 4.5005
R7061 vdd.n1092 vdd.n1048 4.5005
R7062 vdd.n1050 vdd.n1048 4.5005
R7063 vdd.n1046 vdd.n1044 4.5005
R7064 vdd.n4513 vdd.n4512 4.5005
R7065 vdd.n1065 vdd.n1064 4.5005
R7066 vdd.n1065 vdd.n1063 4.5005
R7067 vdd.n4486 vdd.n4485 4.5005
R7068 vdd.n1136 vdd.n1135 4.5005
R7069 vdd.n1137 vdd.n1136 4.5005
R7070 vdd.n1023 vdd.n987 4.5005
R7071 vdd.n989 vdd.n987 4.5005
R7072 vdd.n4538 vdd.n4537 4.5005
R7073 vdd.n4540 vdd.n4539 4.5005
R7074 vdd.n971 vdd.n949 4.5005
R7075 vdd.n4542 vdd.n4541 4.5005
R7076 vdd.n4542 vdd.n948 4.5005
R7077 vdd.n969 vdd.n968 4.5005
R7078 vdd.n4554 vdd.n4553 4.5005
R7079 vdd.n965 vdd.n921 4.5005
R7080 vdd.n923 vdd.n921 4.5005
R7081 vdd.n919 vdd.n917 4.5005
R7082 vdd.n4565 vdd.n4564 4.5005
R7083 vdd.n938 vdd.n937 4.5005
R7084 vdd.n938 vdd.n936 4.5005
R7085 vdd.n4567 vdd.n4566 4.5005
R7086 vdd.n902 vdd.n860 4.5005
R7087 vdd.n4569 vdd.n4568 4.5005
R7088 vdd.n4569 vdd.n859 4.5005
R7089 vdd.n900 vdd.n899 4.5005
R7090 vdd.n885 vdd.n884 4.5005
R7091 vdd.n896 vdd.n895 4.5005
R7092 vdd.n896 vdd.n853 4.5005
R7093 vdd.n3853 vdd.n3852 4.5005
R7094 vdd.n3863 vdd.n3862 4.5005
R7095 vdd.n3861 vdd.n3860 4.5005
R7096 vdd.n4596 vdd.n843 4.5005
R7097 vdd.n4616 vdd.n4615 4.5005
R7098 vdd.n4614 vdd.n4613 4.5005
R7099 vdd.n802 vdd.n796 4.5005
R7100 vdd.n4721 vdd.n4720 4.5005
R7101 vdd.n4691 vdd.n4690 4.5005
R7102 vdd.n754 vdd.n753 4.5005
R7103 vdd.n752 vdd.n741 4.5005
R7104 vdd.n4800 vdd.n4799 4.5005
R7105 vdd.n4895 vdd.n4894 4.5005
R7106 vdd.n679 vdd.n672 4.5005
R7107 vdd.n4919 vdd.n4918 4.5005
R7108 vdd.n619 vdd.n618 4.5005
R7109 vdd.n617 vdd.n606 4.5005
R7110 vdd.n5028 vdd.n5027 4.5005
R7111 vdd.n5123 vdd.n5122 4.5005
R7112 vdd.n544 vdd.n537 4.5005
R7113 vdd.n5147 vdd.n5146 4.5005
R7114 vdd.n484 vdd.n483 4.5005
R7115 vdd.n482 vdd.n471 4.5005
R7116 vdd.n5256 vdd.n5255 4.5005
R7117 vdd.n5351 vdd.n5350 4.5005
R7118 vdd.n409 vdd.n402 4.5005
R7119 vdd.n5375 vdd.n5374 4.5005
R7120 vdd.n349 vdd.n348 4.5005
R7121 vdd.n347 vdd.n346 4.5005
R7122 vdd.n332 vdd.n331 4.5005
R7123 vdd.n5568 vdd.n5567 4.5005
R7124 vdd.n5546 vdd.n5545 4.5005
R7125 vdd.n5548 vdd.n5547 4.5005
R7126 vdd.n5531 vdd.n5530 4.5005
R7127 vdd.n5529 vdd.n5528 4.5005
R7128 vdd.n5512 vdd.n5511 4.5005
R7129 vdd.n316 vdd.n314 4.5005
R7130 vdd.n5487 vdd.n5486 4.5005
R7131 vdd.n293 vdd.n290 4.5005
R7132 vdd.n5457 vdd.n5456 4.5005
R7133 vdd.n371 vdd.n362 4.5005
R7134 vdd.n5434 vdd.n5433 4.5005
R7135 vdd.n5421 vdd.n367 4.5005
R7136 vdd.n5419 vdd.n5418 4.5005
R7137 vdd.n385 vdd.n383 4.5005
R7138 vdd.n5405 vdd.n5404 4.5005
R7139 vdd.n397 vdd.n391 4.5005
R7140 vdd.n357 vdd.n341 4.5005
R7141 vdd.n5331 vdd.n5330 4.5005
R7142 vdd.n5312 vdd.n424 4.5005
R7143 vdd.n434 vdd.n425 4.5005
R7144 vdd.n445 vdd.n443 4.5005
R7145 vdd.n5291 vdd.n5290 4.5005
R7146 vdd.n5273 vdd.n5272 4.5005
R7147 vdd.n5275 vdd.n5274 4.5005
R7148 vdd.n5258 vdd.n5257 4.5005
R7149 vdd.n5329 vdd.n5328 4.5005
R7150 vdd.n5230 vdd.n5229 4.5005
R7151 vdd.n506 vdd.n497 4.5005
R7152 vdd.n5206 vdd.n5205 4.5005
R7153 vdd.n5193 vdd.n502 4.5005
R7154 vdd.n5191 vdd.n5190 4.5005
R7155 vdd.n520 vdd.n518 4.5005
R7156 vdd.n5177 vdd.n5176 4.5005
R7157 vdd.n532 vdd.n526 4.5005
R7158 vdd.n492 vdd.n467 4.5005
R7159 vdd.n5103 vdd.n5102 4.5005
R7160 vdd.n5084 vdd.n559 4.5005
R7161 vdd.n569 vdd.n560 4.5005
R7162 vdd.n580 vdd.n578 4.5005
R7163 vdd.n5063 vdd.n5062 4.5005
R7164 vdd.n5045 vdd.n5044 4.5005
R7165 vdd.n5047 vdd.n5046 4.5005
R7166 vdd.n5030 vdd.n5029 4.5005
R7167 vdd.n5101 vdd.n5100 4.5005
R7168 vdd.n5002 vdd.n5001 4.5005
R7169 vdd.n641 vdd.n632 4.5005
R7170 vdd.n4978 vdd.n4977 4.5005
R7171 vdd.n4965 vdd.n637 4.5005
R7172 vdd.n4963 vdd.n4962 4.5005
R7173 vdd.n655 vdd.n653 4.5005
R7174 vdd.n4949 vdd.n4948 4.5005
R7175 vdd.n667 vdd.n661 4.5005
R7176 vdd.n627 vdd.n602 4.5005
R7177 vdd.n4875 vdd.n4874 4.5005
R7178 vdd.n4856 vdd.n694 4.5005
R7179 vdd.n704 vdd.n695 4.5005
R7180 vdd.n715 vdd.n713 4.5005
R7181 vdd.n4835 vdd.n4834 4.5005
R7182 vdd.n4817 vdd.n4816 4.5005
R7183 vdd.n4819 vdd.n4818 4.5005
R7184 vdd.n4802 vdd.n4801 4.5005
R7185 vdd.n4873 vdd.n4872 4.5005
R7186 vdd.n4774 vdd.n4773 4.5005
R7187 vdd.n776 vdd.n767 4.5005
R7188 vdd.n4750 vdd.n4749 4.5005
R7189 vdd.n4737 vdd.n772 4.5005
R7190 vdd.n4735 vdd.n4734 4.5005
R7191 vdd.n790 vdd.n788 4.5005
R7192 vdd.n762 vdd.n737 4.5005
R7193 vdd.n789 vdd.n787 4.5005
R7194 vdd.n787 vdd.n786 4.5005
R7195 vdd.n5544 vdd.n286 4.5005
R7196 vdd.n286 vdd.n285 4.5005
R7197 vdd.n5533 vdd.n5532 4.5005
R7198 vdd.n5534 vdd.n5533 4.5005
R7199 vdd.n317 vdd.n315 4.5005
R7200 vdd.n5508 vdd.n317 4.5005
R7201 vdd.n327 vdd.n326 4.5005
R7202 vdd.n326 vdd.n325 4.5005
R7203 vdd.n292 vdd.n280 4.5005
R7204 vdd.n282 vdd.n280 4.5005
R7205 vdd.n335 vdd.n334 4.5005
R7206 vdd.n334 vdd.n333 4.5005
R7207 vdd.n356 vdd.n355 4.5005
R7208 vdd.n355 vdd.n354 4.5005
R7209 vdd.n5436 vdd.n5435 4.5005
R7210 vdd.n5436 vdd.n366 4.5005
R7211 vdd.n377 vdd.n376 4.5005
R7212 vdd.n378 vdd.n377 4.5005
R7213 vdd.n384 vdd.n382 4.5005
R7214 vdd.n382 vdd.n381 4.5005
R7215 vdd.n342 vdd.n340 4.5005
R7216 vdd.n352 vdd.n342 4.5005
R7217 vdd.n396 vdd.n395 4.5005
R7218 vdd.n395 vdd.n394 4.5005
R7219 vdd.n5314 vdd.n5313 4.5005
R7220 vdd.n5314 vdd.n423 4.5005
R7221 vdd.n433 vdd.n431 4.5005
R7222 vdd.n435 vdd.n433 4.5005
R7223 vdd.n5271 vdd.n439 4.5005
R7224 vdd.n439 vdd.n438 4.5005
R7225 vdd.n5260 vdd.n5259 4.5005
R7226 vdd.n5261 vdd.n5260 4.5005
R7227 vdd.n5327 vdd.n406 4.5005
R7228 vdd.n406 vdd.n405 4.5005
R7229 vdd.n481 vdd.n480 4.5005
R7230 vdd.n480 vdd.n479 4.5005
R7231 vdd.n491 vdd.n490 4.5005
R7232 vdd.n490 vdd.n489 4.5005
R7233 vdd.n5208 vdd.n5207 4.5005
R7234 vdd.n5208 vdd.n501 4.5005
R7235 vdd.n512 vdd.n511 4.5005
R7236 vdd.n513 vdd.n512 4.5005
R7237 vdd.n519 vdd.n517 4.5005
R7238 vdd.n517 vdd.n516 4.5005
R7239 vdd.n468 vdd.n466 4.5005
R7240 vdd.n487 vdd.n468 4.5005
R7241 vdd.n531 vdd.n530 4.5005
R7242 vdd.n530 vdd.n529 4.5005
R7243 vdd.n5086 vdd.n5085 4.5005
R7244 vdd.n5086 vdd.n558 4.5005
R7245 vdd.n568 vdd.n566 4.5005
R7246 vdd.n570 vdd.n568 4.5005
R7247 vdd.n5043 vdd.n574 4.5005
R7248 vdd.n574 vdd.n573 4.5005
R7249 vdd.n5032 vdd.n5031 4.5005
R7250 vdd.n5033 vdd.n5032 4.5005
R7251 vdd.n5099 vdd.n541 4.5005
R7252 vdd.n541 vdd.n540 4.5005
R7253 vdd.n616 vdd.n615 4.5005
R7254 vdd.n615 vdd.n614 4.5005
R7255 vdd.n626 vdd.n625 4.5005
R7256 vdd.n625 vdd.n624 4.5005
R7257 vdd.n4980 vdd.n4979 4.5005
R7258 vdd.n4980 vdd.n636 4.5005
R7259 vdd.n647 vdd.n646 4.5005
R7260 vdd.n648 vdd.n647 4.5005
R7261 vdd.n654 vdd.n652 4.5005
R7262 vdd.n652 vdd.n651 4.5005
R7263 vdd.n603 vdd.n601 4.5005
R7264 vdd.n622 vdd.n603 4.5005
R7265 vdd.n666 vdd.n665 4.5005
R7266 vdd.n665 vdd.n664 4.5005
R7267 vdd.n4858 vdd.n4857 4.5005
R7268 vdd.n4858 vdd.n693 4.5005
R7269 vdd.n703 vdd.n701 4.5005
R7270 vdd.n705 vdd.n703 4.5005
R7271 vdd.n4815 vdd.n709 4.5005
R7272 vdd.n709 vdd.n708 4.5005
R7273 vdd.n4804 vdd.n4803 4.5005
R7274 vdd.n4805 vdd.n4804 4.5005
R7275 vdd.n4871 vdd.n676 4.5005
R7276 vdd.n676 vdd.n675 4.5005
R7277 vdd.n751 vdd.n750 4.5005
R7278 vdd.n750 vdd.n749 4.5005
R7279 vdd.n761 vdd.n760 4.5005
R7280 vdd.n760 vdd.n759 4.5005
R7281 vdd.n4752 vdd.n4751 4.5005
R7282 vdd.n4752 vdd.n771 4.5005
R7283 vdd.n782 vdd.n781 4.5005
R7284 vdd.n783 vdd.n782 4.5005
R7285 vdd.n738 vdd.n736 4.5005
R7286 vdd.n757 vdd.n738 4.5005
R7287 vdd.n801 vdd.n800 4.5005
R7288 vdd.n800 vdd.n799 4.5005
R7289 vdd.n5758 vdd.n5757 4.5005
R7290 vdd.n240 vdd.n222 4.5005
R7291 vdd.n7470 vdd.n7469 4.5005
R7292 vdd.n5812 vdd 4.28667
R7293 vdd.n5727 vdd 4.28667
R7294 vdd.n134 vdd.t49 4.28621
R7295 vdd.n172 vdd.n164 4.23435
R7296 vdd.n9 vdd.n7 4.23435
R7297 vdd.n153 vdd.n150 3.95926
R7298 vdd.n7507 vdd.n194 3.94241
R7299 vdd.n3978 vdd.n3977 3.92207
R7300 vdd.n7464 vdd.n7463 3.81576
R7301 vdd.n3923 vdd.n3869 3.67129
R7302 vdd.n5750 vdd.n242 3.46788
R7303 vdd.n3998 vdd.n3997 3.46651
R7304 vdd.n3986 vdd.n3848 3.46651
R7305 vdd.n4605 vdd.n4604 3.46651
R7306 vdd.n4628 vdd.n841 3.46651
R7307 vdd.n7476 vdd.n7475 3.46651
R7308 vdd.n7492 vdd.n204 3.46607
R7309 vdd.n2160 vdd.n2109 3.46583
R7310 vdd.n2098 vdd.n2096 3.46583
R7311 vdd.n2118 vdd.n2117 3.46583
R7312 vdd.n2242 vdd.n2240 3.46575
R7313 vdd.n2078 vdd.n2075 3.46575
R7314 vdd.n2231 vdd.n2228 3.46575
R7315 vdd.n3829 vdd.n2070 3.46575
R7316 vdd.n2088 vdd.n2086 3.46575
R7317 vdd.n3815 vdd.n2081 3.46575
R7318 vdd.n3960 vdd.n3959 3.46575
R7319 vdd.n3954 vdd.n3953 3.46575
R7320 vdd.n3971 vdd.n3949 3.46575
R7321 vdd.n3916 vdd.n3914 3.46575
R7322 vdd.n3883 vdd.n3881 3.46575
R7323 vdd.n3876 vdd.n3875 3.46575
R7324 vdd.n3938 vdd.n3871 3.46575
R7325 vdd.n3931 vdd.n3912 3.46575
R7326 vdd.n6393 vdd.n6392 3.46323
R7327 vdd.n4671 vdd.n4670 3.46323
R7328 vdd.n2224 vdd.n2223 3.46323
R7329 vdd.n3890 vdd.n3889 3.46323
R7330 vdd.n2128 vdd.n2122 3.46321
R7331 vdd.n3899 vdd.n3893 3.46321
R7332 vdd.n836 vdd.n830 3.46321
R7333 vdd.n5771 vdd.n5765 3.46321
R7334 vdd.n2157 vdd.n2156 3.45968
R7335 vdd.n7515 vdd.n190 3.45611
R7336 vdd.n3810 vdd.n3809 3.45454
R7337 vdd.n7459 vdd.n231 3.45407
R7338 vdd.n7454 vdd.n7453 3.45407
R7339 vdd.n5742 vdd.n5741 3.45407
R7340 vdd.n7439 vdd.n7438 3.45407
R7341 vdd.n7443 vdd.n7442 3.45407
R7342 vdd.n5784 vdd.n5779 3.45407
R7343 vdd.n7427 vdd.n5780 3.45407
R7344 vdd.n5809 vdd.n5804 3.45407
R7345 vdd.n4666 vdd.n4665 3.45407
R7346 vdd.n4650 vdd.n4646 3.45407
R7347 vdd.n4658 vdd.n4657 3.45407
R7348 vdd.n4640 vdd.n4638 3.45407
R7349 vdd.n825 vdd.n821 3.45407
R7350 vdd.n2135 vdd.n2132 3.45353
R7351 vdd.n232 vdd.n230 3.44028
R7352 vdd.n236 vdd.n235 3.44028
R7353 vdd.n5745 vdd.n5744 3.44028
R7354 vdd.n7434 vdd.n7433 3.44028
R7355 vdd.n7446 vdd.n7445 3.44028
R7356 vdd.n5782 vdd.n5773 3.44028
R7357 vdd.n5789 vdd.n5788 3.44028
R7358 vdd.n5806 vdd.n5803 3.44028
R7359 vdd.n4663 vdd.n4662 3.44028
R7360 vdd.n4647 vdd.n4645 3.44028
R7361 vdd.n4655 vdd.n816 3.44028
R7362 vdd.n4637 vdd.n4636 3.44028
R7363 vdd.n822 vdd.n820 3.44028
R7364 vdd.n2245 vdd.n2244 3.4393
R7365 vdd.n3825 vdd.n3824 3.4393
R7366 vdd.n2234 vdd.n2233 3.4393
R7367 vdd.n3832 vdd.n3831 3.4393
R7368 vdd.n2091 vdd.n2090 3.4393
R7369 vdd.n3818 vdd.n3817 3.4393
R7370 vdd.n3963 vdd.n3962 3.4393
R7371 vdd.n3957 vdd.n3956 3.4393
R7372 vdd.n3974 vdd.n3973 3.4393
R7373 vdd.n3926 vdd.n3925 3.4393
R7374 vdd.n3886 vdd.n3885 3.4393
R7375 vdd.n3879 vdd.n3878 3.4393
R7376 vdd.n3941 vdd.n3940 3.4393
R7377 vdd.n3934 vdd.n3933 3.4393
R7378 vdd.n3807 vdd.n2250 3.4393
R7379 vdd.n2899 vdd.n2898 3.43054
R7380 vdd.n4532 vdd.n4531 3.43054
R7381 vdd.n7305 vdd.n7298 3.42985
R7382 vdd.n5584 vdd.n5583 3.42985
R7383 vdd.n2202 vdd.n2201 3.42753
R7384 vdd.n2149 vdd.n2148 3.42753
R7385 vdd.n3852 vdd.n3845 3.42739
R7386 vdd.n4597 vdd.n4596 3.42739
R7387 vdd.n7419 vdd.n7418 3.42653
R7388 vdd.n7471 vdd.n7470 3.4257
R7389 vdd.n7499 vdd.n7498 3.4257
R7390 vdd.n7517 vdd.n7516 3.42514
R7391 vdd.n2134 vdd.n2131 3.42484
R7392 vdd.n6391 vdd.n6390 3.42476
R7393 vdd.n4669 vdd.n4668 3.42476
R7394 vdd.n5735 vdd.n5734 3.42443
R7395 vdd.n4046 vdd.n4045 3.42443
R7396 vdd.n881 vdd.n838 3.42443
R7397 vdd.n6397 vdd.n6385 3.42376
R7398 vdd.n7294 vdd.n7293 3.42376
R7399 vdd.n2904 vdd.n2903 3.42376
R7400 vdd.n3803 vdd.n3802 3.42376
R7401 vdd.n4529 vdd.n4528 3.42376
R7402 vdd.n4050 vdd.n4049 3.42376
R7403 vdd.n4678 vdd.n4677 3.42376
R7404 vdd.n5579 vdd.n5578 3.42376
R7405 vdd.n2199 vdd.n2198 3.42075
R7406 vdd.n2113 vdd.n2106 3.4187
R7407 vdd.n2189 vdd.n2188 3.4187
R7408 vdd.n832 vdd.n829 3.41853
R7409 vdd.n5767 vdd.n5764 3.41853
R7410 vdd.n2188 vdd.n2187 3.41443
R7411 vdd.n7495 vdd.n7494 3.41405
R7412 vdd.n5759 vdd.n5758 3.41388
R7413 vdd.n209 vdd.n208 3.41388
R7414 vdd.n7295 vdd.n7294 3.41326
R7415 vdd.n5580 vdd.n5579 3.41326
R7416 vdd.n3804 vdd.n3803 3.41326
R7417 vdd.n4051 vdd.n4050 3.41326
R7418 vdd.n6397 vdd.n6396 3.41257
R7419 vdd.n4677 vdd.n4674 3.41257
R7420 vdd.n2903 vdd.n2900 3.41257
R7421 vdd.n4530 vdd.n4529 3.41257
R7422 vdd.n2160 vdd.n2159 3.41222
R7423 vdd.n2219 vdd.n2096 3.41222
R7424 vdd.n2141 vdd.n2131 3.41222
R7425 vdd.n2114 vdd.n2113 3.41222
R7426 vdd.n2200 vdd.n2199 3.41222
R7427 vdd.n2117 vdd.n2095 3.41222
R7428 vdd.n3861 vdd.n3843 3.41219
R7429 vdd.n4614 vdd.n4590 3.41219
R7430 vdd.n6394 vdd.n6393 3.41218
R7431 vdd.n5738 vdd.n232 3.41218
R7432 vdd.n7452 vdd.n231 3.41218
R7433 vdd.n5738 vdd.n235 3.41218
R7434 vdd.n7454 vdd.n7452 3.41218
R7435 vdd.n5746 vdd.n5745 3.41218
R7436 vdd.n5741 vdd.n234 3.41218
R7437 vdd.n7433 vdd.n5774 3.41218
R7438 vdd.n7440 vdd.n7439 3.41218
R7439 vdd.n7447 vdd.n7446 3.41218
R7440 vdd.n7442 vdd.n7441 3.41218
R7441 vdd.n7447 vdd.n5773 3.41218
R7442 vdd.n7441 vdd.n5779 3.41218
R7443 vdd.n5788 vdd.n5774 3.41218
R7444 vdd.n7440 vdd.n5780 3.41218
R7445 vdd.n5806 vdd.n5805 3.41218
R7446 vdd.n5804 vdd.n5781 3.41218
R7447 vdd.n4662 vdd.n4661 3.41218
R7448 vdd.n4667 vdd.n4666 3.41218
R7449 vdd.n4672 vdd.n4671 3.41218
R7450 vdd.n4647 vdd.n813 3.41218
R7451 vdd.n4646 vdd.n809 3.41218
R7452 vdd.n4635 vdd.n816 3.41218
R7453 vdd.n4658 vdd.n819 3.41218
R7454 vdd.n4636 vdd.n4635 3.41218
R7455 vdd.n4638 vdd.n819 3.41218
R7456 vdd.n822 vdd.n813 3.41218
R7457 vdd.n821 vdd.n809 3.41218
R7458 vdd.n2245 vdd.n2239 3.41218
R7459 vdd.n3825 vdd.n2074 3.41218
R7460 vdd.n2224 vdd.n2221 3.41218
R7461 vdd.n2234 vdd.n2227 3.41218
R7462 vdd.n3831 vdd.n3830 3.41218
R7463 vdd.n2091 vdd.n2085 3.41218
R7464 vdd.n3817 vdd.n3816 3.41218
R7465 vdd.n3963 vdd.n3958 3.41218
R7466 vdd.n3957 vdd.n3952 3.41218
R7467 vdd.n3973 vdd.n3972 3.41218
R7468 vdd.n3926 vdd.n3913 3.41218
R7469 vdd.n3890 vdd.n3887 3.41218
R7470 vdd.n3886 vdd.n3880 3.41218
R7471 vdd.n3879 vdd.n3874 3.41218
R7472 vdd.n3940 vdd.n3939 3.41218
R7473 vdd.n3934 vdd.n3911 3.41218
R7474 vdd.n3811 vdd.n3810 3.41218
R7475 vdd.n3811 vdd.n2250 3.41218
R7476 vdd.n2141 vdd.n2132 3.41165
R7477 vdd.n2158 vdd.n2157 3.41165
R7478 vdd.n2121 vdd.n2120 3.41162
R7479 vdd.n2123 vdd.n2120 3.41162
R7480 vdd.n3892 vdd.n3891 3.41162
R7481 vdd.n3894 vdd.n3891 3.41162
R7482 vdd.n831 vdd.n828 3.41162
R7483 vdd.n5766 vdd.n5763 3.41162
R7484 vdd.n6417 vdd.n6416 3.4105
R7485 vdd.n6425 vdd.n6424 3.4105
R7486 vdd.n6511 vdd.n6509 3.4105
R7487 vdd.n6530 vdd.n6304 3.4105
R7488 vdd.n6535 vdd.n6295 3.4105
R7489 vdd.n6569 vdd.n6284 3.4105
R7490 vdd.n6590 vdd.n6589 3.4105
R7491 vdd.n6614 vdd.n6613 3.4105
R7492 vdd.n6624 vdd.n6623 3.4105
R7493 vdd.n6738 vdd.n6736 3.4105
R7494 vdd.n6757 vdd.n6171 3.4105
R7495 vdd.n6762 vdd.n6162 3.4105
R7496 vdd.n6796 vdd.n6151 3.4105
R7497 vdd.n6817 vdd.n6816 3.4105
R7498 vdd.n6841 vdd.n6840 3.4105
R7499 vdd.n6851 vdd.n6850 3.4105
R7500 vdd.n6965 vdd.n6963 3.4105
R7501 vdd.n6984 vdd.n6038 3.4105
R7502 vdd.n6989 vdd.n6029 3.4105
R7503 vdd.n7023 vdd.n6018 3.4105
R7504 vdd.n7044 vdd.n7043 3.4105
R7505 vdd.n7068 vdd.n7067 3.4105
R7506 vdd.n7078 vdd.n7077 3.4105
R7507 vdd.n7192 vdd.n7190 3.4105
R7508 vdd.n7211 vdd.n5905 3.4105
R7509 vdd.n7216 vdd.n5896 3.4105
R7510 vdd.n7250 vdd.n5885 3.4105
R7511 vdd.n7271 vdd.n7270 3.4105
R7512 vdd.n7275 vdd.n5867 3.4105
R7513 vdd.n7282 vdd.n7281 3.4105
R7514 vdd.n7257 vdd.n7256 3.4105
R7515 vdd.n5897 vdd.n5893 3.4105
R7516 vdd.n5907 vdd.n5903 3.4105
R7517 vdd.n7209 vdd.n7208 3.4105
R7518 vdd.n7164 vdd.n7163 3.4105
R7519 vdd.n7151 vdd.n7150 3.4105
R7520 vdd.n7144 vdd.n7143 3.4105
R7521 vdd.n7129 vdd.n7128 3.4105
R7522 vdd.n7122 vdd.n5964 3.4105
R7523 vdd.n7117 vdd.n5970 3.4105
R7524 vdd.n7106 vdd.n7105 3.4105
R7525 vdd.n7098 vdd.n7097 3.4105
R7526 vdd.n7171 vdd.n7170 3.4105
R7527 vdd.n7183 vdd.n7182 3.4105
R7528 vdd.n7085 vdd.n7084 3.4105
R7529 vdd.n7075 vdd.n7074 3.4105
R7530 vdd.n7051 vdd.n7050 3.4105
R7531 vdd.n7030 vdd.n7029 3.4105
R7532 vdd.n6030 vdd.n6026 3.4105
R7533 vdd.n6040 vdd.n6036 3.4105
R7534 vdd.n6982 vdd.n6981 3.4105
R7535 vdd.n6937 vdd.n6936 3.4105
R7536 vdd.n6924 vdd.n6923 3.4105
R7537 vdd.n6917 vdd.n6916 3.4105
R7538 vdd.n6902 vdd.n6901 3.4105
R7539 vdd.n6895 vdd.n6097 3.4105
R7540 vdd.n6890 vdd.n6103 3.4105
R7541 vdd.n6879 vdd.n6878 3.4105
R7542 vdd.n6871 vdd.n6870 3.4105
R7543 vdd.n6944 vdd.n6943 3.4105
R7544 vdd.n6956 vdd.n6955 3.4105
R7545 vdd.n6858 vdd.n6857 3.4105
R7546 vdd.n6848 vdd.n6847 3.4105
R7547 vdd.n6824 vdd.n6823 3.4105
R7548 vdd.n6803 vdd.n6802 3.4105
R7549 vdd.n6163 vdd.n6159 3.4105
R7550 vdd.n6173 vdd.n6169 3.4105
R7551 vdd.n6755 vdd.n6754 3.4105
R7552 vdd.n6710 vdd.n6709 3.4105
R7553 vdd.n6697 vdd.n6696 3.4105
R7554 vdd.n6690 vdd.n6689 3.4105
R7555 vdd.n6675 vdd.n6674 3.4105
R7556 vdd.n6668 vdd.n6230 3.4105
R7557 vdd.n6663 vdd.n6236 3.4105
R7558 vdd.n6652 vdd.n6651 3.4105
R7559 vdd.n6644 vdd.n6643 3.4105
R7560 vdd.n6717 vdd.n6716 3.4105
R7561 vdd.n6729 vdd.n6728 3.4105
R7562 vdd.n6631 vdd.n6630 3.4105
R7563 vdd.n6621 vdd.n6620 3.4105
R7564 vdd.n6597 vdd.n6596 3.4105
R7565 vdd.n6576 vdd.n6575 3.4105
R7566 vdd.n6296 vdd.n6292 3.4105
R7567 vdd.n6306 vdd.n6302 3.4105
R7568 vdd.n6528 vdd.n6527 3.4105
R7569 vdd.n6483 vdd.n6482 3.4105
R7570 vdd.n6470 vdd.n6469 3.4105
R7571 vdd.n6463 vdd.n6462 3.4105
R7572 vdd.n6448 vdd.n6447 3.4105
R7573 vdd.n6441 vdd.n6363 3.4105
R7574 vdd.n6436 vdd.n6369 3.4105
R7575 vdd.n6490 vdd.n6489 3.4105
R7576 vdd.n6502 vdd.n6501 3.4105
R7577 vdd.n6404 vdd.n6403 3.4105
R7578 vdd.n7409 vdd.n5792 3.4105
R7579 vdd.n7407 vdd.n7406 3.4105
R7580 vdd.n7305 vdd.n7304 3.4105
R7581 vdd.n7312 vdd.n7311 3.4105
R7582 vdd.n7392 vdd.n7391 3.4105
R7583 vdd.n7381 vdd.n7380 3.4105
R7584 vdd.n7369 vdd.n7368 3.4105
R7585 vdd.n7362 vdd.n7361 3.4105
R7586 vdd.n7350 vdd.n7349 3.4105
R7587 vdd.n7343 vdd.n7342 3.4105
R7588 vdd.n7331 vdd.n7330 3.4105
R7589 vdd.n7324 vdd.n7323 3.4105
R7590 vdd.n7403 vdd.n5797 3.4105
R7591 vdd.n5585 vdd.n5584 3.4105
R7592 vdd.n5586 vdd.n274 3.4105
R7593 vdd.n5716 vdd.n5715 3.4105
R7594 vdd.n5607 vdd.n5605 3.4105
R7595 vdd.n5606 vdd.n5604 3.4105
R7596 vdd.n5644 vdd.n5643 3.4105
R7597 vdd.n5632 vdd.n5610 3.4105
R7598 vdd.n5673 vdd.n5649 3.4105
R7599 vdd.n5691 vdd.n5690 3.4105
R7600 vdd.n5654 vdd.n5653 3.4105
R7601 vdd.n5683 vdd.n5682 3.4105
R7602 vdd.n5599 vdd.n267 3.4105
R7603 vdd.n5657 vdd.n245 3.4105
R7604 vdd.n5658 vdd.n5656 3.4105
R7605 vdd.n5662 vdd.n5661 3.4105
R7606 vdd.n5647 vdd.n5629 3.4105
R7607 vdd.n5687 vdd.n5630 3.4105
R7608 vdd.n5686 vdd.n5685 3.4105
R7609 vdd.n5684 vdd.n5648 3.4105
R7610 vdd.n5646 vdd.n5645 3.4105
R7611 vdd.n5636 vdd.n5635 3.4105
R7612 vdd.n5639 vdd.n5631 3.4105
R7613 vdd.n5712 vdd.n272 3.4105
R7614 vdd.n5709 vdd.n5603 3.4105
R7615 vdd.n5634 vdd.n5633 3.4105
R7616 vdd.n5714 vdd.n5713 3.4105
R7617 vdd.n5598 vdd.n273 3.4105
R7618 vdd.n5602 vdd.n271 3.4105
R7619 vdd.n5595 vdd.n5594 3.4105
R7620 vdd.n5597 vdd.n5596 3.4105
R7621 vdd.n5660 vdd.n5659 3.4105
R7622 vdd.n2187 vdd.n2186 3.4105
R7623 vdd.n2147 vdd.n2146 3.4105
R7624 vdd.n2163 vdd.n2110 3.4105
R7625 vdd.n2152 vdd.n2111 3.4105
R7626 vdd.n2124 vdd.n2121 3.4105
R7627 vdd.n2124 vdd.n2123 3.4105
R7628 vdd.n2084 vdd.n2083 3.4105
R7629 vdd.n3814 vdd.n2083 3.4105
R7630 vdd.n2093 vdd.n2092 3.4105
R7631 vdd.n2092 vdd.n2087 3.4105
R7632 vdd.n2143 vdd.n2094 3.4105
R7633 vdd.n2130 vdd.n2119 3.4105
R7634 vdd.n2141 vdd.n2140 3.4105
R7635 vdd.n2908 vdd.n2907 3.4105
R7636 vdd.n3738 vdd.n3737 3.4105
R7637 vdd.n3722 vdd.n3721 3.4105
R7638 vdd.n2285 vdd.n2281 3.4105
R7639 vdd.n3740 vdd.n2283 3.4105
R7640 vdd.n2275 vdd.n2271 3.4105
R7641 vdd.n3745 vdd.n2274 3.4105
R7642 vdd.n3790 vdd.n3789 3.4105
R7643 vdd.n3779 vdd.n2261 3.4105
R7644 vdd.n3783 vdd.n2255 3.4105
R7645 vdd.n3714 vdd.n3713 3.4105
R7646 vdd.n3701 vdd.n3700 3.4105
R7647 vdd.n3599 vdd.n3598 3.4105
R7648 vdd.n3613 vdd.n3612 3.4105
R7649 vdd.n3629 vdd.n3628 3.4105
R7650 vdd.n3625 vdd.n3623 3.4105
R7651 vdd.n3646 vdd.n2350 3.4105
R7652 vdd.n3651 vdd.n2344 3.4105
R7653 vdd.n3658 vdd.n3657 3.4105
R7654 vdd.n3674 vdd.n3673 3.4105
R7655 vdd.n3681 vdd.n3680 3.4105
R7656 vdd.n3694 vdd.n3693 3.4105
R7657 vdd.n3568 vdd.n2386 3.4105
R7658 vdd.n3592 vdd.n3591 3.4105
R7659 vdd.n2428 vdd.n2424 3.4105
R7660 vdd.n3474 vdd.n2427 3.4105
R7661 vdd.n3515 vdd.n3514 3.4105
R7662 vdd.n3508 vdd.n2416 3.4105
R7663 vdd.n3537 vdd.n3536 3.4105
R7664 vdd.n3529 vdd.n3528 3.4105
R7665 vdd.n2394 vdd.n2390 3.4105
R7666 vdd.n2403 vdd.n2393 3.4105
R7667 vdd.n3575 vdd.n3574 3.4105
R7668 vdd.n3564 vdd.n2383 3.4105
R7669 vdd.n2438 vdd.n2434 3.4105
R7670 vdd.n3469 vdd.n2436 3.4105
R7671 vdd.n3371 vdd.n3370 3.4105
R7672 vdd.n3385 vdd.n3384 3.4105
R7673 vdd.n3401 vdd.n3400 3.4105
R7674 vdd.n3397 vdd.n3395 3.4105
R7675 vdd.n3418 vdd.n2485 3.4105
R7676 vdd.n3423 vdd.n2479 3.4105
R7677 vdd.n3430 vdd.n3429 3.4105
R7678 vdd.n3446 vdd.n3445 3.4105
R7679 vdd.n3454 vdd.n3453 3.4105
R7680 vdd.n3467 vdd.n3466 3.4105
R7681 vdd.n3340 vdd.n2521 3.4105
R7682 vdd.n3364 vdd.n3363 3.4105
R7683 vdd.n2563 vdd.n2559 3.4105
R7684 vdd.n3246 vdd.n2562 3.4105
R7685 vdd.n3287 vdd.n3286 3.4105
R7686 vdd.n3280 vdd.n2551 3.4105
R7687 vdd.n3309 vdd.n3308 3.4105
R7688 vdd.n3301 vdd.n3300 3.4105
R7689 vdd.n2529 vdd.n2525 3.4105
R7690 vdd.n2538 vdd.n2528 3.4105
R7691 vdd.n3347 vdd.n3346 3.4105
R7692 vdd.n3336 vdd.n2518 3.4105
R7693 vdd.n2573 vdd.n2569 3.4105
R7694 vdd.n3241 vdd.n2571 3.4105
R7695 vdd.n3143 vdd.n3142 3.4105
R7696 vdd.n3157 vdd.n3156 3.4105
R7697 vdd.n3173 vdd.n3172 3.4105
R7698 vdd.n3169 vdd.n3167 3.4105
R7699 vdd.n3190 vdd.n2620 3.4105
R7700 vdd.n3195 vdd.n2614 3.4105
R7701 vdd.n3202 vdd.n3201 3.4105
R7702 vdd.n3218 vdd.n3217 3.4105
R7703 vdd.n3226 vdd.n3225 3.4105
R7704 vdd.n3239 vdd.n3238 3.4105
R7705 vdd.n3112 vdd.n2656 3.4105
R7706 vdd.n3136 vdd.n3135 3.4105
R7707 vdd.n2698 vdd.n2694 3.4105
R7708 vdd.n3018 vdd.n2697 3.4105
R7709 vdd.n3059 vdd.n3058 3.4105
R7710 vdd.n3052 vdd.n2686 3.4105
R7711 vdd.n3081 vdd.n3080 3.4105
R7712 vdd.n3073 vdd.n3072 3.4105
R7713 vdd.n2664 vdd.n2660 3.4105
R7714 vdd.n2673 vdd.n2663 3.4105
R7715 vdd.n3119 vdd.n3118 3.4105
R7716 vdd.n3108 vdd.n2653 3.4105
R7717 vdd.n2708 vdd.n2704 3.4105
R7718 vdd.n3013 vdd.n2706 3.4105
R7719 vdd.n2945 vdd.n2944 3.4105
R7720 vdd.n2941 vdd.n2939 3.4105
R7721 vdd.n2962 vdd.n2755 3.4105
R7722 vdd.n2967 vdd.n2749 3.4105
R7723 vdd.n2974 vdd.n2973 3.4105
R7724 vdd.n2990 vdd.n2989 3.4105
R7725 vdd.n2998 vdd.n2997 3.4105
R7726 vdd.n3011 vdd.n3010 3.4105
R7727 vdd.n2929 vdd.n2928 3.4105
R7728 vdd.n2915 vdd.n2914 3.4105
R7729 vdd.n4041 vdd.n4040 3.4105
R7730 vdd.n2893 vdd.n2892 3.4105
R7731 vdd.n4013 vdd.n2047 3.4105
R7732 vdd.n4033 vdd.n4032 3.4105
R7733 vdd.n2820 vdd.n2052 3.4105
R7734 vdd.n2831 vdd.n2815 3.4105
R7735 vdd.n2836 vdd.n2810 3.4105
R7736 vdd.n2843 vdd.n2842 3.4105
R7737 vdd.n2859 vdd.n2858 3.4105
R7738 vdd.n2866 vdd.n2865 3.4105
R7739 vdd.n2886 vdd.n2885 3.4105
R7740 vdd.n2898 vdd.n2897 3.4105
R7741 vdd.n4043 vdd.n4042 3.4105
R7742 vdd.n1021 vdd.n986 3.4105
R7743 vdd.n1966 vdd.n1953 3.4105
R7744 vdd.n4100 vdd.n4099 3.4105
R7745 vdd.n1990 vdd.n1989 3.4105
R7746 vdd.n4092 vdd.n4091 3.4105
R7747 vdd.n2008 vdd.n1995 3.4105
R7748 vdd.n4078 vdd.n4077 3.4105
R7749 vdd.n2032 vdd.n2031 3.4105
R7750 vdd.n4070 vdd.n4069 3.4105
R7751 vdd.n4056 vdd.n4055 3.4105
R7752 vdd.n1948 vdd.n1947 3.4105
R7753 vdd.n4114 vdd.n4113 3.4105
R7754 vdd.n1823 vdd.n1822 3.4105
R7755 vdd.n1829 vdd.n1805 3.4105
R7756 vdd.n1810 vdd.n1807 3.4105
R7757 vdd.n1834 vdd.n1809 3.4105
R7758 vdd.n4141 vdd.n4140 3.4105
R7759 vdd.n1882 vdd.n1839 3.4105
R7760 vdd.n1892 vdd.n1891 3.4105
R7761 vdd.n1898 vdd.n1869 3.4105
R7762 vdd.n1874 vdd.n1871 3.4105
R7763 vdd.n1903 vdd.n1873 3.4105
R7764 vdd.n1779 vdd.n1773 3.4105
R7765 vdd.n4165 vdd.n1778 3.4105
R7766 vdd.n1702 vdd.n1689 3.4105
R7767 vdd.n4221 vdd.n4220 3.4105
R7768 vdd.n1726 vdd.n1725 3.4105
R7769 vdd.n4213 vdd.n4212 3.4105
R7770 vdd.n1744 vdd.n1731 3.4105
R7771 vdd.n4199 vdd.n4198 3.4105
R7772 vdd.n1768 vdd.n1767 3.4105
R7773 vdd.n4191 vdd.n4190 3.4105
R7774 vdd.n1780 vdd.n1772 3.4105
R7775 vdd.n4177 vdd.n4176 3.4105
R7776 vdd.n1684 vdd.n1683 3.4105
R7777 vdd.n4235 vdd.n4234 3.4105
R7778 vdd.n1559 vdd.n1558 3.4105
R7779 vdd.n1565 vdd.n1541 3.4105
R7780 vdd.n1546 vdd.n1543 3.4105
R7781 vdd.n1570 vdd.n1545 3.4105
R7782 vdd.n4262 vdd.n4261 3.4105
R7783 vdd.n1618 vdd.n1575 3.4105
R7784 vdd.n1628 vdd.n1627 3.4105
R7785 vdd.n1634 vdd.n1605 3.4105
R7786 vdd.n1610 vdd.n1607 3.4105
R7787 vdd.n1639 vdd.n1609 3.4105
R7788 vdd.n1515 vdd.n1509 3.4105
R7789 vdd.n4286 vdd.n1514 3.4105
R7790 vdd.n1438 vdd.n1425 3.4105
R7791 vdd.n4342 vdd.n4341 3.4105
R7792 vdd.n1462 vdd.n1461 3.4105
R7793 vdd.n4334 vdd.n4333 3.4105
R7794 vdd.n1480 vdd.n1467 3.4105
R7795 vdd.n4320 vdd.n4319 3.4105
R7796 vdd.n1504 vdd.n1503 3.4105
R7797 vdd.n4312 vdd.n4311 3.4105
R7798 vdd.n1516 vdd.n1508 3.4105
R7799 vdd.n4298 vdd.n4297 3.4105
R7800 vdd.n1420 vdd.n1419 3.4105
R7801 vdd.n4356 vdd.n4355 3.4105
R7802 vdd.n1295 vdd.n1294 3.4105
R7803 vdd.n1301 vdd.n1277 3.4105
R7804 vdd.n1282 vdd.n1279 3.4105
R7805 vdd.n1306 vdd.n1281 3.4105
R7806 vdd.n4383 vdd.n4382 3.4105
R7807 vdd.n1354 vdd.n1311 3.4105
R7808 vdd.n1364 vdd.n1363 3.4105
R7809 vdd.n1370 vdd.n1341 3.4105
R7810 vdd.n1346 vdd.n1343 3.4105
R7811 vdd.n1375 vdd.n1345 3.4105
R7812 vdd.n1251 vdd.n1245 3.4105
R7813 vdd.n4407 vdd.n1250 3.4105
R7814 vdd.n1174 vdd.n1161 3.4105
R7815 vdd.n4463 vdd.n4462 3.4105
R7816 vdd.n1198 vdd.n1197 3.4105
R7817 vdd.n4455 vdd.n4454 3.4105
R7818 vdd.n1216 vdd.n1203 3.4105
R7819 vdd.n4441 vdd.n4440 3.4105
R7820 vdd.n1240 vdd.n1239 3.4105
R7821 vdd.n4433 vdd.n4432 3.4105
R7822 vdd.n1252 vdd.n1244 3.4105
R7823 vdd.n4419 vdd.n4418 3.4105
R7824 vdd.n1156 vdd.n1155 3.4105
R7825 vdd.n4477 vdd.n4476 3.4105
R7826 vdd.n1014 vdd.n1011 3.4105
R7827 vdd.n1042 vdd.n1013 3.4105
R7828 vdd.n4504 vdd.n4503 3.4105
R7829 vdd.n1090 vdd.n1047 3.4105
R7830 vdd.n1100 vdd.n1099 3.4105
R7831 vdd.n1106 vdd.n1077 3.4105
R7832 vdd.n1082 vdd.n1079 3.4105
R7833 vdd.n1111 vdd.n1081 3.4105
R7834 vdd.n1037 vdd.n1009 3.4105
R7835 vdd.n1031 vdd.n1030 3.4105
R7836 vdd.n887 vdd.n886 3.4105
R7837 vdd.n955 vdd.n952 3.4105
R7838 vdd.n894 vdd.n893 3.4105
R7839 vdd.n904 vdd.n903 3.4105
R7840 vdd.n910 vdd.n861 3.4105
R7841 vdd.n866 vdd.n863 3.4105
R7842 vdd.n915 vdd.n865 3.4105
R7843 vdd.n4556 vdd.n4555 3.4105
R7844 vdd.n963 vdd.n920 3.4105
R7845 vdd.n973 vdd.n972 3.4105
R7846 vdd.n979 vdd.n950 3.4105
R7847 vdd.n4531 vdd.n954 3.4105
R7848 vdd.n877 vdd.n875 3.4105
R7849 vdd.n982 vdd.n981 3.4105
R7850 vdd.n4535 vdd.n4534 3.4105
R7851 vdd.n980 vdd.n957 3.4105
R7852 vdd.n975 vdd.n974 3.4105
R7853 vdd.n976 vdd.n958 3.4105
R7854 vdd.n964 vdd.n959 3.4105
R7855 vdd.n4557 vdd.n914 3.4105
R7856 vdd.n960 vdd.n916 3.4105
R7857 vdd.n4559 vdd.n4558 3.4105
R7858 vdd.n913 vdd.n912 3.4105
R7859 vdd.n4562 vdd.n4561 3.4105
R7860 vdd.n911 vdd.n868 3.4105
R7861 vdd.n906 vdd.n905 3.4105
R7862 vdd.n907 vdd.n869 3.4105
R7863 vdd.n871 vdd.n870 3.4105
R7864 vdd.n889 vdd.n888 3.4105
R7865 vdd.n890 vdd.n873 3.4105
R7866 vdd.n878 vdd.n874 3.4105
R7867 vdd.n2035 vdd.n2025 3.4105
R7868 vdd.n4052 vdd.n2026 3.4105
R7869 vdd.n2034 vdd.n2033 3.4105
R7870 vdd.n4071 vdd.n1994 3.4105
R7871 vdd.n2029 vdd.n2028 3.4105
R7872 vdd.n1993 vdd.n1983 3.4105
R7873 vdd.n4074 vdd.n1984 3.4105
R7874 vdd.n4073 vdd.n4072 3.4105
R7875 vdd.n1992 vdd.n1991 3.4105
R7876 vdd.n4093 vdd.n1952 3.4105
R7877 vdd.n1987 vdd.n1986 3.4105
R7878 vdd.n1951 vdd.n1941 3.4105
R7879 vdd.n4096 vdd.n1942 3.4105
R7880 vdd.n4095 vdd.n4094 3.4105
R7881 vdd.n1950 vdd.n1949 3.4105
R7882 vdd.n4115 vdd.n1902 3.4105
R7883 vdd.n1945 vdd.n1944 3.4105
R7884 vdd.n1901 vdd.n1900 3.4105
R7885 vdd.n4120 vdd.n4119 3.4105
R7886 vdd.n4117 vdd.n4116 3.4105
R7887 vdd.n1899 vdd.n1876 3.4105
R7888 vdd.n1894 vdd.n1893 3.4105
R7889 vdd.n1895 vdd.n1877 3.4105
R7890 vdd.n4142 vdd.n1833 3.4105
R7891 vdd.n1879 vdd.n1835 3.4105
R7892 vdd.n1883 vdd.n1878 3.4105
R7893 vdd.n4144 vdd.n4143 3.4105
R7894 vdd.n1832 vdd.n1831 3.4105
R7895 vdd.n4147 vdd.n4146 3.4105
R7896 vdd.n1825 vdd.n1824 3.4105
R7897 vdd.n1826 vdd.n1813 3.4105
R7898 vdd.n1830 vdd.n1812 3.4105
R7899 vdd.n1815 vdd.n1814 3.4105
R7900 vdd.n4170 vdd.n4169 3.4105
R7901 vdd.n4168 vdd.n4167 3.4105
R7902 vdd.n1771 vdd.n1761 3.4105
R7903 vdd.n4173 vdd.n1762 3.4105
R7904 vdd.n4172 vdd.n4171 3.4105
R7905 vdd.n1770 vdd.n1769 3.4105
R7906 vdd.n4192 vdd.n1730 3.4105
R7907 vdd.n1765 vdd.n1764 3.4105
R7908 vdd.n1729 vdd.n1719 3.4105
R7909 vdd.n4195 vdd.n1720 3.4105
R7910 vdd.n4194 vdd.n4193 3.4105
R7911 vdd.n1728 vdd.n1727 3.4105
R7912 vdd.n4214 vdd.n1688 3.4105
R7913 vdd.n1723 vdd.n1722 3.4105
R7914 vdd.n1687 vdd.n1677 3.4105
R7915 vdd.n4217 vdd.n1678 3.4105
R7916 vdd.n4216 vdd.n4215 3.4105
R7917 vdd.n1686 vdd.n1685 3.4105
R7918 vdd.n4236 vdd.n1638 3.4105
R7919 vdd.n1681 vdd.n1680 3.4105
R7920 vdd.n1637 vdd.n1636 3.4105
R7921 vdd.n4241 vdd.n4240 3.4105
R7922 vdd.n4238 vdd.n4237 3.4105
R7923 vdd.n1635 vdd.n1612 3.4105
R7924 vdd.n1630 vdd.n1629 3.4105
R7925 vdd.n1631 vdd.n1613 3.4105
R7926 vdd.n4263 vdd.n1569 3.4105
R7927 vdd.n1615 vdd.n1571 3.4105
R7928 vdd.n1619 vdd.n1614 3.4105
R7929 vdd.n4265 vdd.n4264 3.4105
R7930 vdd.n1568 vdd.n1567 3.4105
R7931 vdd.n4268 vdd.n4267 3.4105
R7932 vdd.n1561 vdd.n1560 3.4105
R7933 vdd.n1562 vdd.n1549 3.4105
R7934 vdd.n1566 vdd.n1548 3.4105
R7935 vdd.n1551 vdd.n1550 3.4105
R7936 vdd.n4291 vdd.n4290 3.4105
R7937 vdd.n4289 vdd.n4288 3.4105
R7938 vdd.n1507 vdd.n1497 3.4105
R7939 vdd.n4294 vdd.n1498 3.4105
R7940 vdd.n4293 vdd.n4292 3.4105
R7941 vdd.n1506 vdd.n1505 3.4105
R7942 vdd.n4313 vdd.n1466 3.4105
R7943 vdd.n1501 vdd.n1500 3.4105
R7944 vdd.n1465 vdd.n1455 3.4105
R7945 vdd.n4316 vdd.n1456 3.4105
R7946 vdd.n4315 vdd.n4314 3.4105
R7947 vdd.n1464 vdd.n1463 3.4105
R7948 vdd.n4335 vdd.n1424 3.4105
R7949 vdd.n1459 vdd.n1458 3.4105
R7950 vdd.n1423 vdd.n1413 3.4105
R7951 vdd.n4338 vdd.n1414 3.4105
R7952 vdd.n4337 vdd.n4336 3.4105
R7953 vdd.n1422 vdd.n1421 3.4105
R7954 vdd.n4357 vdd.n1374 3.4105
R7955 vdd.n1417 vdd.n1416 3.4105
R7956 vdd.n1373 vdd.n1372 3.4105
R7957 vdd.n4362 vdd.n4361 3.4105
R7958 vdd.n4359 vdd.n4358 3.4105
R7959 vdd.n1371 vdd.n1348 3.4105
R7960 vdd.n1366 vdd.n1365 3.4105
R7961 vdd.n1367 vdd.n1349 3.4105
R7962 vdd.n4384 vdd.n1305 3.4105
R7963 vdd.n1351 vdd.n1307 3.4105
R7964 vdd.n1355 vdd.n1350 3.4105
R7965 vdd.n4386 vdd.n4385 3.4105
R7966 vdd.n1304 vdd.n1303 3.4105
R7967 vdd.n4389 vdd.n4388 3.4105
R7968 vdd.n1297 vdd.n1296 3.4105
R7969 vdd.n1298 vdd.n1285 3.4105
R7970 vdd.n1302 vdd.n1284 3.4105
R7971 vdd.n1287 vdd.n1286 3.4105
R7972 vdd.n4412 vdd.n4411 3.4105
R7973 vdd.n4410 vdd.n4409 3.4105
R7974 vdd.n1243 vdd.n1233 3.4105
R7975 vdd.n4415 vdd.n1234 3.4105
R7976 vdd.n4414 vdd.n4413 3.4105
R7977 vdd.n1242 vdd.n1241 3.4105
R7978 vdd.n4434 vdd.n1202 3.4105
R7979 vdd.n1237 vdd.n1236 3.4105
R7980 vdd.n1201 vdd.n1191 3.4105
R7981 vdd.n4437 vdd.n1192 3.4105
R7982 vdd.n4436 vdd.n4435 3.4105
R7983 vdd.n1200 vdd.n1199 3.4105
R7984 vdd.n4456 vdd.n1160 3.4105
R7985 vdd.n1195 vdd.n1194 3.4105
R7986 vdd.n1159 vdd.n1149 3.4105
R7987 vdd.n4459 vdd.n1150 3.4105
R7988 vdd.n4458 vdd.n4457 3.4105
R7989 vdd.n1158 vdd.n1157 3.4105
R7990 vdd.n4478 vdd.n1110 3.4105
R7991 vdd.n1153 vdd.n1152 3.4105
R7992 vdd.n1109 vdd.n1108 3.4105
R7993 vdd.n4483 vdd.n4482 3.4105
R7994 vdd.n4480 vdd.n4479 3.4105
R7995 vdd.n1107 vdd.n1084 3.4105
R7996 vdd.n1102 vdd.n1101 3.4105
R7997 vdd.n1103 vdd.n1085 3.4105
R7998 vdd.n4505 vdd.n1041 3.4105
R7999 vdd.n1087 vdd.n1043 3.4105
R8000 vdd.n1091 vdd.n1086 3.4105
R8001 vdd.n4507 vdd.n4506 3.4105
R8002 vdd.n1040 vdd.n1039 3.4105
R8003 vdd.n4510 vdd.n4509 3.4105
R8004 vdd.n1033 vdd.n1032 3.4105
R8005 vdd.n1034 vdd.n1017 3.4105
R8006 vdd.n1038 vdd.n1016 3.4105
R8007 vdd.n1022 vdd.n1018 3.4105
R8008 vdd.n984 vdd.n983 3.4105
R8009 vdd.n3895 vdd.n3892 3.4105
R8010 vdd.n3895 vdd.n3894 3.4105
R8011 vdd.n3936 vdd.n3935 3.4105
R8012 vdd.n3935 vdd.n3929 3.4105
R8013 vdd.n3910 vdd.n3873 3.4105
R8014 vdd.n3937 vdd.n3873 3.4105
R8015 vdd.n3908 vdd.n3907 3.4105
R8016 vdd.n3909 vdd.n3908 3.4105
R8017 vdd.n3905 vdd.n3904 3.4105
R8018 vdd.n3906 vdd.n3905 3.4105
R8019 vdd.n3902 vdd.n3901 3.4105
R8020 vdd.n3903 vdd.n3902 3.4105
R8021 vdd.n3928 vdd.n3927 3.4105
R8022 vdd.n3927 vdd.n2036 3.4105
R8023 vdd.n3849 vdd.n3844 3.4105
R8024 vdd.n3994 vdd.n3993 3.4105
R8025 vdd.n3851 vdd.n3850 3.4105
R8026 vdd.n3996 vdd.n3995 3.4105
R8027 vdd.n3969 vdd.n3951 3.4105
R8028 vdd.n3970 vdd.n3951 3.4105
R8029 vdd.n3967 vdd.n3966 3.4105
R8030 vdd.n3968 vdd.n3967 3.4105
R8031 vdd.n3964 vdd.n3847 3.4105
R8032 vdd.n3965 vdd.n3964 3.4105
R8033 vdd.n3989 vdd.n3841 3.4105
R8034 vdd.n3989 vdd.n3988 3.4105
R8035 vdd.n3991 vdd.n3990 3.4105
R8036 vdd.n2889 vdd.n2789 3.4105
R8037 vdd.n2891 vdd.n2890 3.4105
R8038 vdd.n2888 vdd.n2887 3.4105
R8039 vdd.n2862 vdd.n2800 3.4105
R8040 vdd.n2864 vdd.n2863 3.4105
R8041 vdd.n2839 vdd.n2813 3.4105
R8042 vdd.n2841 vdd.n2840 3.4105
R8043 vdd.n2861 vdd.n2860 3.4105
R8044 vdd.n2838 vdd.n2837 3.4105
R8045 vdd.n2823 vdd.n2822 3.4105
R8046 vdd.n2834 vdd.n2824 3.4105
R8047 vdd.n4034 vdd.n2046 3.4105
R8048 vdd.n2817 vdd.n2048 3.4105
R8049 vdd.n2821 vdd.n2816 3.4105
R8050 vdd.n4036 vdd.n4035 3.4105
R8051 vdd.n2045 vdd.n2041 3.4105
R8052 vdd.n4039 vdd.n4038 3.4105
R8053 vdd.n2044 vdd.n2039 3.4105
R8054 vdd.n3786 vdd.n2269 3.4105
R8055 vdd.n2252 vdd.n2251 3.4105
R8056 vdd.n3788 vdd.n3787 3.4105
R8057 vdd.n3778 vdd.n2270 3.4105
R8058 vdd.n3782 vdd.n2268 3.4105
R8059 vdd.n3777 vdd.n3776 3.4105
R8060 vdd.n3746 vdd.n3744 3.4105
R8061 vdd.n3775 vdd.n3774 3.4105
R8062 vdd.n3748 vdd.n3747 3.4105
R8063 vdd.n3742 vdd.n3741 3.4105
R8064 vdd.n3750 vdd.n3749 3.4105
R8065 vdd.n3739 vdd.n2286 3.4105
R8066 vdd.n3717 vdd.n2303 3.4105
R8067 vdd.n3718 vdd.n2287 3.4105
R8068 vdd.n3716 vdd.n3715 3.4105
R8069 vdd.n3697 vdd.n2312 3.4105
R8070 vdd.n2305 vdd.n2304 3.4105
R8071 vdd.n3696 vdd.n3695 3.4105
R8072 vdd.n3677 vdd.n2334 3.4105
R8073 vdd.n3679 vdd.n3678 3.4105
R8074 vdd.n3676 vdd.n3675 3.4105
R8075 vdd.n3654 vdd.n2348 3.4105
R8076 vdd.n3656 vdd.n3655 3.4105
R8077 vdd.n3653 vdd.n3652 3.4105
R8078 vdd.n3620 vdd.n3618 3.4105
R8079 vdd.n3649 vdd.n2351 3.4105
R8080 vdd.n3622 vdd.n3621 3.4105
R8081 vdd.n3616 vdd.n2362 3.4105
R8082 vdd.n3627 vdd.n3617 3.4105
R8083 vdd.n3615 vdd.n3614 3.4105
R8084 vdd.n3595 vdd.n2374 3.4105
R8085 vdd.n3597 vdd.n3596 3.4105
R8086 vdd.n3594 vdd.n3593 3.4105
R8087 vdd.n3571 vdd.n2388 3.4105
R8088 vdd.n3570 vdd.n3569 3.4105
R8089 vdd.n3573 vdd.n3572 3.4105
R8090 vdd.n3563 vdd.n2389 3.4105
R8091 vdd.n3567 vdd.n2387 3.4105
R8092 vdd.n3562 vdd.n3561 3.4105
R8093 vdd.n3533 vdd.n2404 3.4105
R8094 vdd.n3560 vdd.n3559 3.4105
R8095 vdd.n3535 vdd.n3534 3.4105
R8096 vdd.n2406 vdd.n2405 3.4105
R8097 vdd.n3532 vdd.n2402 3.4105
R8098 vdd.n3513 vdd.n3512 3.4105
R8099 vdd.n3507 vdd.n2423 3.4105
R8100 vdd.n3511 vdd.n2422 3.4105
R8101 vdd.n3506 vdd.n3505 3.4105
R8102 vdd.n3475 vdd.n3473 3.4105
R8103 vdd.n3504 vdd.n3503 3.4105
R8104 vdd.n3477 vdd.n3476 3.4105
R8105 vdd.n3471 vdd.n3470 3.4105
R8106 vdd.n3479 vdd.n3478 3.4105
R8107 vdd.n3468 vdd.n2439 3.4105
R8108 vdd.n3449 vdd.n2469 3.4105
R8109 vdd.n3452 vdd.n3451 3.4105
R8110 vdd.n3448 vdd.n3447 3.4105
R8111 vdd.n3426 vdd.n2483 3.4105
R8112 vdd.n3428 vdd.n3427 3.4105
R8113 vdd.n3425 vdd.n3424 3.4105
R8114 vdd.n3392 vdd.n3390 3.4105
R8115 vdd.n3421 vdd.n2486 3.4105
R8116 vdd.n3394 vdd.n3393 3.4105
R8117 vdd.n3388 vdd.n2497 3.4105
R8118 vdd.n3399 vdd.n3389 3.4105
R8119 vdd.n3387 vdd.n3386 3.4105
R8120 vdd.n3367 vdd.n2509 3.4105
R8121 vdd.n3369 vdd.n3368 3.4105
R8122 vdd.n3366 vdd.n3365 3.4105
R8123 vdd.n3343 vdd.n2523 3.4105
R8124 vdd.n3342 vdd.n3341 3.4105
R8125 vdd.n3345 vdd.n3344 3.4105
R8126 vdd.n3335 vdd.n2524 3.4105
R8127 vdd.n3339 vdd.n2522 3.4105
R8128 vdd.n3334 vdd.n3333 3.4105
R8129 vdd.n3305 vdd.n2539 3.4105
R8130 vdd.n3332 vdd.n3331 3.4105
R8131 vdd.n3307 vdd.n3306 3.4105
R8132 vdd.n2541 vdd.n2540 3.4105
R8133 vdd.n3304 vdd.n2537 3.4105
R8134 vdd.n3285 vdd.n3284 3.4105
R8135 vdd.n3279 vdd.n2558 3.4105
R8136 vdd.n3283 vdd.n2557 3.4105
R8137 vdd.n3278 vdd.n3277 3.4105
R8138 vdd.n3247 vdd.n3245 3.4105
R8139 vdd.n3276 vdd.n3275 3.4105
R8140 vdd.n3249 vdd.n3248 3.4105
R8141 vdd.n3243 vdd.n3242 3.4105
R8142 vdd.n3251 vdd.n3250 3.4105
R8143 vdd.n3240 vdd.n2574 3.4105
R8144 vdd.n3221 vdd.n2604 3.4105
R8145 vdd.n3224 vdd.n3223 3.4105
R8146 vdd.n3220 vdd.n3219 3.4105
R8147 vdd.n3198 vdd.n2618 3.4105
R8148 vdd.n3200 vdd.n3199 3.4105
R8149 vdd.n3197 vdd.n3196 3.4105
R8150 vdd.n3164 vdd.n3162 3.4105
R8151 vdd.n3193 vdd.n2621 3.4105
R8152 vdd.n3166 vdd.n3165 3.4105
R8153 vdd.n3160 vdd.n2632 3.4105
R8154 vdd.n3171 vdd.n3161 3.4105
R8155 vdd.n3159 vdd.n3158 3.4105
R8156 vdd.n3139 vdd.n2644 3.4105
R8157 vdd.n3141 vdd.n3140 3.4105
R8158 vdd.n3138 vdd.n3137 3.4105
R8159 vdd.n3115 vdd.n2658 3.4105
R8160 vdd.n3114 vdd.n3113 3.4105
R8161 vdd.n3117 vdd.n3116 3.4105
R8162 vdd.n3107 vdd.n2659 3.4105
R8163 vdd.n3111 vdd.n2657 3.4105
R8164 vdd.n3106 vdd.n3105 3.4105
R8165 vdd.n3077 vdd.n2674 3.4105
R8166 vdd.n3104 vdd.n3103 3.4105
R8167 vdd.n3079 vdd.n3078 3.4105
R8168 vdd.n2676 vdd.n2675 3.4105
R8169 vdd.n3076 vdd.n2672 3.4105
R8170 vdd.n3057 vdd.n3056 3.4105
R8171 vdd.n3051 vdd.n2693 3.4105
R8172 vdd.n3055 vdd.n2692 3.4105
R8173 vdd.n3050 vdd.n3049 3.4105
R8174 vdd.n3019 vdd.n3017 3.4105
R8175 vdd.n3048 vdd.n3047 3.4105
R8176 vdd.n3021 vdd.n3020 3.4105
R8177 vdd.n3015 vdd.n3014 3.4105
R8178 vdd.n3023 vdd.n3022 3.4105
R8179 vdd.n3012 vdd.n2709 3.4105
R8180 vdd.n2993 vdd.n2739 3.4105
R8181 vdd.n2996 vdd.n2995 3.4105
R8182 vdd.n2992 vdd.n2991 3.4105
R8183 vdd.n2970 vdd.n2753 3.4105
R8184 vdd.n2972 vdd.n2971 3.4105
R8185 vdd.n2969 vdd.n2968 3.4105
R8186 vdd.n2936 vdd.n2934 3.4105
R8187 vdd.n2965 vdd.n2756 3.4105
R8188 vdd.n2938 vdd.n2937 3.4105
R8189 vdd.n2932 vdd.n2767 3.4105
R8190 vdd.n2943 vdd.n2933 3.4105
R8191 vdd.n2931 vdd.n2930 3.4105
R8192 vdd.n2911 vdd.n2779 3.4105
R8193 vdd.n2913 vdd.n2912 3.4105
R8194 vdd.n2910 vdd.n2909 3.4105
R8195 vdd.n2902 vdd.n2901 3.4105
R8196 vdd.n2073 vdd.n2072 3.4105
R8197 vdd.n3828 vdd.n2072 3.4105
R8198 vdd.n2236 vdd.n2235 3.4105
R8199 vdd.n2235 vdd.n2229 3.4105
R8200 vdd.n3827 vdd.n3826 3.4105
R8201 vdd.n3826 vdd.n2076 3.4105
R8202 vdd.n2247 vdd.n2246 3.4105
R8203 vdd.n2248 vdd.n2247 3.4105
R8204 vdd.n3805 vdd.n2249 3.4105
R8205 vdd.n4595 vdd.n4594 3.4105
R8206 vdd.n4601 vdd.n4600 3.4105
R8207 vdd.n4593 vdd.n842 3.4105
R8208 vdd.n4603 vdd.n4602 3.4105
R8209 vdd.n4631 vdd.n840 3.4105
R8210 vdd.n4631 vdd.n4630 3.4105
R8211 vdd.n4598 vdd.n839 3.4105
R8212 vdd.n832 vdd.n831 3.4105
R8213 vdd.n837 vdd.n836 3.4105
R8214 vdd.n5562 vdd.n295 3.4105
R8215 vdd.n5564 vdd.n5563 3.4105
R8216 vdd.n5554 vdd.n296 3.4105
R8217 vdd.n5553 vdd.n5552 3.4105
R8218 vdd.n5522 vdd.n5520 3.4105
R8219 vdd.n5524 vdd.n5523 3.4105
R8220 vdd.n5518 vdd.n5517 3.4105
R8221 vdd.n5515 vdd.n312 3.4105
R8222 vdd.n5492 vdd.n328 3.4105
R8223 vdd.n5491 vdd.n5490 3.4105
R8224 vdd.n5471 vdd.n336 3.4105
R8225 vdd.n5470 vdd.n5469 3.4105
R8226 vdd.n5451 vdd.n358 3.4105
R8227 vdd.n5450 vdd.n5449 3.4105
R8228 vdd.n5428 vdd.n372 3.4105
R8229 vdd.n5427 vdd.n5426 3.4105
R8230 vdd.n5394 vdd.n5392 3.4105
R8231 vdd.n5396 vdd.n5395 3.4105
R8232 vdd.n5390 vdd.n386 3.4105
R8233 vdd.n5389 vdd.n5388 3.4105
R8234 vdd.n5369 vdd.n398 3.4105
R8235 vdd.n5368 vdd.n5367 3.4105
R8236 vdd.n5345 vdd.n412 3.4105
R8237 vdd.n5347 vdd.n5346 3.4105
R8238 vdd.n5337 vdd.n413 3.4105
R8239 vdd.n5336 vdd.n5335 3.4105
R8240 vdd.n5307 vdd.n428 3.4105
R8241 vdd.n5309 vdd.n5308 3.4105
R8242 vdd.n430 vdd.n429 3.4105
R8243 vdd.n5287 vdd.n5286 3.4105
R8244 vdd.n5281 vdd.n447 3.4105
R8245 vdd.n5280 vdd.n5279 3.4105
R8246 vdd.n5249 vdd.n5247 3.4105
R8247 vdd.n5251 vdd.n5250 3.4105
R8248 vdd.n5245 vdd.n5244 3.4105
R8249 vdd.n5242 vdd.n463 3.4105
R8250 vdd.n5223 vdd.n493 3.4105
R8251 vdd.n5222 vdd.n5221 3.4105
R8252 vdd.n5200 vdd.n507 3.4105
R8253 vdd.n5199 vdd.n5198 3.4105
R8254 vdd.n5166 vdd.n5164 3.4105
R8255 vdd.n5168 vdd.n5167 3.4105
R8256 vdd.n5162 vdd.n521 3.4105
R8257 vdd.n5161 vdd.n5160 3.4105
R8258 vdd.n5141 vdd.n533 3.4105
R8259 vdd.n5140 vdd.n5139 3.4105
R8260 vdd.n5117 vdd.n547 3.4105
R8261 vdd.n5119 vdd.n5118 3.4105
R8262 vdd.n5109 vdd.n548 3.4105
R8263 vdd.n5108 vdd.n5107 3.4105
R8264 vdd.n5079 vdd.n563 3.4105
R8265 vdd.n5081 vdd.n5080 3.4105
R8266 vdd.n565 vdd.n564 3.4105
R8267 vdd.n5059 vdd.n5058 3.4105
R8268 vdd.n5053 vdd.n582 3.4105
R8269 vdd.n5052 vdd.n5051 3.4105
R8270 vdd.n5021 vdd.n5019 3.4105
R8271 vdd.n5023 vdd.n5022 3.4105
R8272 vdd.n5017 vdd.n5016 3.4105
R8273 vdd.n5014 vdd.n598 3.4105
R8274 vdd.n4995 vdd.n628 3.4105
R8275 vdd.n4994 vdd.n4993 3.4105
R8276 vdd.n4972 vdd.n642 3.4105
R8277 vdd.n4971 vdd.n4970 3.4105
R8278 vdd.n4938 vdd.n4936 3.4105
R8279 vdd.n4940 vdd.n4939 3.4105
R8280 vdd.n4934 vdd.n656 3.4105
R8281 vdd.n4933 vdd.n4932 3.4105
R8282 vdd.n4913 vdd.n668 3.4105
R8283 vdd.n4912 vdd.n4911 3.4105
R8284 vdd.n4889 vdd.n682 3.4105
R8285 vdd.n4891 vdd.n4890 3.4105
R8286 vdd.n4881 vdd.n683 3.4105
R8287 vdd.n4880 vdd.n4879 3.4105
R8288 vdd.n4851 vdd.n698 3.4105
R8289 vdd.n4853 vdd.n4852 3.4105
R8290 vdd.n700 vdd.n699 3.4105
R8291 vdd.n4831 vdd.n4830 3.4105
R8292 vdd.n4825 vdd.n717 3.4105
R8293 vdd.n4824 vdd.n4823 3.4105
R8294 vdd.n4793 vdd.n4791 3.4105
R8295 vdd.n4795 vdd.n4794 3.4105
R8296 vdd.n4789 vdd.n4788 3.4105
R8297 vdd.n4786 vdd.n733 3.4105
R8298 vdd.n4767 vdd.n763 3.4105
R8299 vdd.n4766 vdd.n4765 3.4105
R8300 vdd.n4744 vdd.n777 3.4105
R8301 vdd.n4743 vdd.n4742 3.4105
R8302 vdd.n4710 vdd.n4708 3.4105
R8303 vdd.n4712 vdd.n4711 3.4105
R8304 vdd.n4706 vdd.n791 3.4105
R8305 vdd.n4705 vdd.n4704 3.4105
R8306 vdd.n4685 vdd.n803 3.4105
R8307 vdd.n4684 vdd.n4683 3.4105
R8308 vdd.n278 vdd.n277 3.4105
R8309 vdd.n5558 vdd.n294 3.4105
R8310 vdd.n5551 vdd.n5550 3.4105
R8311 vdd.n5526 vdd.n5525 3.4105
R8312 vdd.n5493 vdd.n313 3.4105
R8313 vdd.n330 vdd.n329 3.4105
R8314 vdd.n5453 vdd.n5452 3.4105
R8315 vdd.n5430 vdd.n5429 3.4105
R8316 vdd.n5423 vdd.n375 3.4105
R8317 vdd.n5401 vdd.n5391 3.4105
R8318 vdd.n5371 vdd.n5370 3.4105
R8319 vdd.n5344 vdd.n5343 3.4105
R8320 vdd.n5341 vdd.n411 3.4105
R8321 vdd.n5334 vdd.n5333 3.4105
R8322 vdd.n5306 vdd.n426 3.4105
R8323 vdd.n5285 vdd.n446 3.4105
R8324 vdd.n5278 vdd.n5277 3.4105
R8325 vdd.n5253 vdd.n5252 3.4105
R8326 vdd.n5226 vdd.n5225 3.4105
R8327 vdd.n5202 vdd.n5201 3.4105
R8328 vdd.n5195 vdd.n510 3.4105
R8329 vdd.n5173 vdd.n5163 3.4105
R8330 vdd.n5143 vdd.n5142 3.4105
R8331 vdd.n5116 vdd.n5115 3.4105
R8332 vdd.n5113 vdd.n546 3.4105
R8333 vdd.n5106 vdd.n5105 3.4105
R8334 vdd.n5078 vdd.n561 3.4105
R8335 vdd.n5057 vdd.n581 3.4105
R8336 vdd.n5050 vdd.n5049 3.4105
R8337 vdd.n5025 vdd.n5024 3.4105
R8338 vdd.n4998 vdd.n4997 3.4105
R8339 vdd.n4974 vdd.n4973 3.4105
R8340 vdd.n4967 vdd.n645 3.4105
R8341 vdd.n4945 vdd.n4935 3.4105
R8342 vdd.n4915 vdd.n4914 3.4105
R8343 vdd.n4888 vdd.n4887 3.4105
R8344 vdd.n4885 vdd.n681 3.4105
R8345 vdd.n4878 vdd.n4877 3.4105
R8346 vdd.n4850 vdd.n696 3.4105
R8347 vdd.n4829 vdd.n716 3.4105
R8348 vdd.n4822 vdd.n4821 3.4105
R8349 vdd.n4797 vdd.n4796 3.4105
R8350 vdd.n4770 vdd.n4769 3.4105
R8351 vdd.n4746 vdd.n4745 3.4105
R8352 vdd.n4739 vdd.n780 3.4105
R8353 vdd.n4717 vdd.n4707 3.4105
R8354 vdd.n4687 vdd.n4686 3.4105
R8355 vdd.n4682 vdd.n4681 3.4105
R8356 vdd.n5514 vdd.n5513 3.4105
R8357 vdd.n5498 vdd.n5496 3.4105
R8358 vdd.n311 vdd.n307 3.4105
R8359 vdd.n5516 vdd.n309 3.4105
R8360 vdd.n301 vdd.n297 3.4105
R8361 vdd.n5521 vdd.n300 3.4105
R8362 vdd.n5566 vdd.n5565 3.4105
R8363 vdd.n5555 vdd.n287 3.4105
R8364 vdd.n5559 vdd.n281 3.4105
R8365 vdd.n5489 vdd.n5488 3.4105
R8366 vdd.n5476 vdd.n5474 3.4105
R8367 vdd.n5373 vdd.n5372 3.4105
R8368 vdd.n5387 vdd.n5386 3.4105
R8369 vdd.n5403 vdd.n5402 3.4105
R8370 vdd.n5399 vdd.n5397 3.4105
R8371 vdd.n5420 vdd.n374 3.4105
R8372 vdd.n5425 vdd.n368 3.4105
R8373 vdd.n5432 vdd.n5431 3.4105
R8374 vdd.n5448 vdd.n5447 3.4105
R8375 vdd.n5455 vdd.n5454 3.4105
R8376 vdd.n5468 vdd.n5467 3.4105
R8377 vdd.n5342 vdd.n410 3.4105
R8378 vdd.n5366 vdd.n5365 3.4105
R8379 vdd.n452 vdd.n448 3.4105
R8380 vdd.n5248 vdd.n451 3.4105
R8381 vdd.n5289 vdd.n5288 3.4105
R8382 vdd.n5282 vdd.n440 3.4105
R8383 vdd.n5311 vdd.n5310 3.4105
R8384 vdd.n5303 vdd.n5302 3.4105
R8385 vdd.n418 vdd.n414 3.4105
R8386 vdd.n427 vdd.n417 3.4105
R8387 vdd.n5349 vdd.n5348 3.4105
R8388 vdd.n5338 vdd.n407 3.4105
R8389 vdd.n462 vdd.n458 3.4105
R8390 vdd.n5243 vdd.n460 3.4105
R8391 vdd.n5145 vdd.n5144 3.4105
R8392 vdd.n5159 vdd.n5158 3.4105
R8393 vdd.n5175 vdd.n5174 3.4105
R8394 vdd.n5171 vdd.n5169 3.4105
R8395 vdd.n5192 vdd.n509 3.4105
R8396 vdd.n5197 vdd.n503 3.4105
R8397 vdd.n5204 vdd.n5203 3.4105
R8398 vdd.n5220 vdd.n5219 3.4105
R8399 vdd.n5228 vdd.n5227 3.4105
R8400 vdd.n5241 vdd.n5240 3.4105
R8401 vdd.n5114 vdd.n545 3.4105
R8402 vdd.n5138 vdd.n5137 3.4105
R8403 vdd.n587 vdd.n583 3.4105
R8404 vdd.n5020 vdd.n586 3.4105
R8405 vdd.n5061 vdd.n5060 3.4105
R8406 vdd.n5054 vdd.n575 3.4105
R8407 vdd.n5083 vdd.n5082 3.4105
R8408 vdd.n5075 vdd.n5074 3.4105
R8409 vdd.n553 vdd.n549 3.4105
R8410 vdd.n562 vdd.n552 3.4105
R8411 vdd.n5121 vdd.n5120 3.4105
R8412 vdd.n5110 vdd.n542 3.4105
R8413 vdd.n597 vdd.n593 3.4105
R8414 vdd.n5015 vdd.n595 3.4105
R8415 vdd.n4917 vdd.n4916 3.4105
R8416 vdd.n4931 vdd.n4930 3.4105
R8417 vdd.n4947 vdd.n4946 3.4105
R8418 vdd.n4943 vdd.n4941 3.4105
R8419 vdd.n4964 vdd.n644 3.4105
R8420 vdd.n4969 vdd.n638 3.4105
R8421 vdd.n4976 vdd.n4975 3.4105
R8422 vdd.n4992 vdd.n4991 3.4105
R8423 vdd.n5000 vdd.n4999 3.4105
R8424 vdd.n5013 vdd.n5012 3.4105
R8425 vdd.n4886 vdd.n680 3.4105
R8426 vdd.n4910 vdd.n4909 3.4105
R8427 vdd.n722 vdd.n718 3.4105
R8428 vdd.n4792 vdd.n721 3.4105
R8429 vdd.n4833 vdd.n4832 3.4105
R8430 vdd.n4826 vdd.n710 3.4105
R8431 vdd.n4855 vdd.n4854 3.4105
R8432 vdd.n4847 vdd.n4846 3.4105
R8433 vdd.n688 vdd.n684 3.4105
R8434 vdd.n697 vdd.n687 3.4105
R8435 vdd.n4893 vdd.n4892 3.4105
R8436 vdd.n4882 vdd.n677 3.4105
R8437 vdd.n732 vdd.n728 3.4105
R8438 vdd.n4787 vdd.n730 3.4105
R8439 vdd.n4719 vdd.n4718 3.4105
R8440 vdd.n4715 vdd.n4713 3.4105
R8441 vdd.n4736 vdd.n779 3.4105
R8442 vdd.n4741 vdd.n773 3.4105
R8443 vdd.n4748 vdd.n4747 3.4105
R8444 vdd.n4764 vdd.n4763 3.4105
R8445 vdd.n4772 vdd.n4771 3.4105
R8446 vdd.n4785 vdd.n4784 3.4105
R8447 vdd.n4703 vdd.n4702 3.4105
R8448 vdd.n4689 vdd.n4688 3.4105
R8449 vdd.n4676 vdd.n4675 3.4105
R8450 vdd.n5762 vdd.n5760 3.4105
R8451 vdd.n7472 vdd.n219 3.4105
R8452 vdd.n7474 vdd.n7473 3.4105
R8453 vdd.n239 vdd.n238 3.4105
R8454 vdd.n7450 vdd.n218 3.4105
R8455 vdd.n7451 vdd.n220 3.4105
R8456 vdd.n5748 vdd.n5747 3.4105
R8457 vdd.n5767 vdd.n5766 3.4105
R8458 vdd.n5772 vdd.n5771 3.4105
R8459 vdd.n6399 vdd.n6398 3.4105
R8460 vdd.n6402 vdd.n6401 3.4105
R8461 vdd.n6423 vdd.n6422 3.4105
R8462 vdd.n7278 vdd.n5874 3.4105
R8463 vdd.n5864 vdd.n5863 3.4105
R8464 vdd.n7280 vdd.n7279 3.4105
R8465 vdd.n5876 vdd.n5875 3.4105
R8466 vdd.n7274 vdd.n5873 3.4105
R8467 vdd.n7255 vdd.n7254 3.4105
R8468 vdd.n7249 vdd.n5892 3.4105
R8469 vdd.n7253 vdd.n5891 3.4105
R8470 vdd.n7248 vdd.n7247 3.4105
R8471 vdd.n7217 vdd.n7215 3.4105
R8472 vdd.n7246 vdd.n7245 3.4105
R8473 vdd.n7219 vdd.n7218 3.4105
R8474 vdd.n7213 vdd.n7212 3.4105
R8475 vdd.n7221 vdd.n7220 3.4105
R8476 vdd.n7210 vdd.n5908 3.4105
R8477 vdd.n7186 vdd.n5921 3.4105
R8478 vdd.n7187 vdd.n5909 3.4105
R8479 vdd.n7104 vdd.n7103 3.4105
R8480 vdd.n5982 vdd.n5981 3.4105
R8481 vdd.n7100 vdd.n7099 3.4105
R8482 vdd.n7124 vdd.n7123 3.4105
R8483 vdd.n7102 vdd.n5980 3.4105
R8484 vdd.n7120 vdd.n5971 3.4105
R8485 vdd.n7146 vdd.n7145 3.4105
R8486 vdd.n7125 vdd.n5968 3.4105
R8487 vdd.n7127 vdd.n7126 3.4105
R8488 vdd.n7166 vdd.n7165 3.4105
R8489 vdd.n7147 vdd.n5954 3.4105
R8490 vdd.n7149 vdd.n7148 3.4105
R8491 vdd.n7185 vdd.n7184 3.4105
R8492 vdd.n7167 vdd.n5943 3.4105
R8493 vdd.n7169 vdd.n7168 3.4105
R8494 vdd.n7083 vdd.n7082 3.4105
R8495 vdd.n5992 vdd.n5991 3.4105
R8496 vdd.n7080 vdd.n7079 3.4105
R8497 vdd.n7073 vdd.n7072 3.4105
R8498 vdd.n5996 vdd.n5995 3.4105
R8499 vdd.n7071 vdd.n5994 3.4105
R8500 vdd.n7049 vdd.n7048 3.4105
R8501 vdd.n6009 vdd.n6008 3.4105
R8502 vdd.n7047 vdd.n6007 3.4105
R8503 vdd.n7028 vdd.n7027 3.4105
R8504 vdd.n7022 vdd.n6025 3.4105
R8505 vdd.n7026 vdd.n6024 3.4105
R8506 vdd.n7021 vdd.n7020 3.4105
R8507 vdd.n6990 vdd.n6988 3.4105
R8508 vdd.n7019 vdd.n7018 3.4105
R8509 vdd.n6992 vdd.n6991 3.4105
R8510 vdd.n6986 vdd.n6985 3.4105
R8511 vdd.n6994 vdd.n6993 3.4105
R8512 vdd.n6983 vdd.n6041 3.4105
R8513 vdd.n6959 vdd.n6054 3.4105
R8514 vdd.n6960 vdd.n6042 3.4105
R8515 vdd.n6877 vdd.n6876 3.4105
R8516 vdd.n6115 vdd.n6114 3.4105
R8517 vdd.n6873 vdd.n6872 3.4105
R8518 vdd.n6897 vdd.n6896 3.4105
R8519 vdd.n6875 vdd.n6113 3.4105
R8520 vdd.n6893 vdd.n6104 3.4105
R8521 vdd.n6919 vdd.n6918 3.4105
R8522 vdd.n6898 vdd.n6101 3.4105
R8523 vdd.n6900 vdd.n6899 3.4105
R8524 vdd.n6939 vdd.n6938 3.4105
R8525 vdd.n6920 vdd.n6087 3.4105
R8526 vdd.n6922 vdd.n6921 3.4105
R8527 vdd.n6958 vdd.n6957 3.4105
R8528 vdd.n6940 vdd.n6076 3.4105
R8529 vdd.n6942 vdd.n6941 3.4105
R8530 vdd.n6856 vdd.n6855 3.4105
R8531 vdd.n6125 vdd.n6124 3.4105
R8532 vdd.n6853 vdd.n6852 3.4105
R8533 vdd.n6846 vdd.n6845 3.4105
R8534 vdd.n6129 vdd.n6128 3.4105
R8535 vdd.n6844 vdd.n6127 3.4105
R8536 vdd.n6822 vdd.n6821 3.4105
R8537 vdd.n6142 vdd.n6141 3.4105
R8538 vdd.n6820 vdd.n6140 3.4105
R8539 vdd.n6801 vdd.n6800 3.4105
R8540 vdd.n6795 vdd.n6158 3.4105
R8541 vdd.n6799 vdd.n6157 3.4105
R8542 vdd.n6794 vdd.n6793 3.4105
R8543 vdd.n6763 vdd.n6761 3.4105
R8544 vdd.n6792 vdd.n6791 3.4105
R8545 vdd.n6765 vdd.n6764 3.4105
R8546 vdd.n6759 vdd.n6758 3.4105
R8547 vdd.n6767 vdd.n6766 3.4105
R8548 vdd.n6756 vdd.n6174 3.4105
R8549 vdd.n6732 vdd.n6187 3.4105
R8550 vdd.n6733 vdd.n6175 3.4105
R8551 vdd.n6650 vdd.n6649 3.4105
R8552 vdd.n6248 vdd.n6247 3.4105
R8553 vdd.n6646 vdd.n6645 3.4105
R8554 vdd.n6670 vdd.n6669 3.4105
R8555 vdd.n6648 vdd.n6246 3.4105
R8556 vdd.n6666 vdd.n6237 3.4105
R8557 vdd.n6692 vdd.n6691 3.4105
R8558 vdd.n6671 vdd.n6234 3.4105
R8559 vdd.n6673 vdd.n6672 3.4105
R8560 vdd.n6712 vdd.n6711 3.4105
R8561 vdd.n6693 vdd.n6220 3.4105
R8562 vdd.n6695 vdd.n6694 3.4105
R8563 vdd.n6731 vdd.n6730 3.4105
R8564 vdd.n6713 vdd.n6209 3.4105
R8565 vdd.n6715 vdd.n6714 3.4105
R8566 vdd.n6629 vdd.n6628 3.4105
R8567 vdd.n6258 vdd.n6257 3.4105
R8568 vdd.n6626 vdd.n6625 3.4105
R8569 vdd.n6619 vdd.n6618 3.4105
R8570 vdd.n6262 vdd.n6261 3.4105
R8571 vdd.n6617 vdd.n6260 3.4105
R8572 vdd.n6595 vdd.n6594 3.4105
R8573 vdd.n6275 vdd.n6274 3.4105
R8574 vdd.n6593 vdd.n6273 3.4105
R8575 vdd.n6574 vdd.n6573 3.4105
R8576 vdd.n6568 vdd.n6291 3.4105
R8577 vdd.n6572 vdd.n6290 3.4105
R8578 vdd.n6567 vdd.n6566 3.4105
R8579 vdd.n6536 vdd.n6534 3.4105
R8580 vdd.n6565 vdd.n6564 3.4105
R8581 vdd.n6538 vdd.n6537 3.4105
R8582 vdd.n6532 vdd.n6531 3.4105
R8583 vdd.n6540 vdd.n6539 3.4105
R8584 vdd.n6529 vdd.n6307 3.4105
R8585 vdd.n6505 vdd.n6320 3.4105
R8586 vdd.n6506 vdd.n6308 3.4105
R8587 vdd.n6443 vdd.n6442 3.4105
R8588 vdd.n6421 vdd.n6379 3.4105
R8589 vdd.n6439 vdd.n6370 3.4105
R8590 vdd.n6465 vdd.n6464 3.4105
R8591 vdd.n6444 vdd.n6367 3.4105
R8592 vdd.n6446 vdd.n6445 3.4105
R8593 vdd.n6485 vdd.n6484 3.4105
R8594 vdd.n6466 vdd.n6353 3.4105
R8595 vdd.n6468 vdd.n6467 3.4105
R8596 vdd.n6504 vdd.n6503 3.4105
R8597 vdd.n6486 vdd.n6342 3.4105
R8598 vdd.n6488 vdd.n6487 3.4105
R8599 vdd.n6419 vdd.n6418 3.4105
R8600 vdd.n6381 vdd.n6380 3.4105
R8601 vdd.n7408 vdd.n5794 3.4105
R8602 vdd.n7388 vdd.n5818 3.4105
R8603 vdd.n5820 vdd.n5819 3.4105
R8604 vdd.n7384 vdd.n5817 3.4105
R8605 vdd.n7390 vdd.n7389 3.4105
R8606 vdd.n7367 vdd.n7366 3.4105
R8607 vdd.n5831 vdd.n5830 3.4105
R8608 vdd.n7365 vdd.n5829 3.4105
R8609 vdd.n5842 vdd.n5841 3.4105
R8610 vdd.n7346 vdd.n5840 3.4105
R8611 vdd.n7348 vdd.n7347 3.4105
R8612 vdd.n7329 vdd.n7328 3.4105
R8613 vdd.n5853 vdd.n5852 3.4105
R8614 vdd.n7327 vdd.n5851 3.4105
R8615 vdd.n7411 vdd.n7410 3.4105
R8616 vdd.n7308 vdd.n5862 3.4105
R8617 vdd.n7310 vdd.n7309 3.4105
R8618 vdd.n7385 vdd.n5795 3.4105
R8619 vdd.n7496 vdd.n203 3.4105
R8620 vdd.n7497 vdd.n7496 3.4105
R8621 vdd.n205 vdd.n200 3.4105
R8622 vdd.n7494 vdd.n206 3.4105
R8623 vdd.n207 vdd.n202 3.4105
R8624 vdd.n7413 vdd.n201 3.4105
R8625 vdd.n7201 vdd.n7198 3.38568
R8626 vdd.n7234 vdd.n5882 3.38568
R8627 vdd.n6974 vdd.n6971 3.38568
R8628 vdd.n7007 vdd.n6015 3.38568
R8629 vdd.n7064 vdd.n7058 3.38568
R8630 vdd.n6747 vdd.n6744 3.38568
R8631 vdd.n6780 vdd.n6148 3.38568
R8632 vdd.n6837 vdd.n6831 3.38568
R8633 vdd.n6520 vdd.n6517 3.38568
R8634 vdd.n6553 vdd.n6281 3.38568
R8635 vdd.n6610 vdd.n6604 3.38568
R8636 vdd.n7400 vdd.n7399 3.38568
R8637 vdd.n7160 vdd.n5938 3.38568
R8638 vdd.n6933 vdd.n6071 3.38568
R8639 vdd.n6706 vdd.n6204 3.38568
R8640 vdd.n6479 vdd.n6337 3.38568
R8641 vdd.n5383 vdd.n5382 3.38568
R8642 vdd.n5440 vdd.n5439 3.38568
R8643 vdd.n5155 vdd.n5154 3.38568
R8644 vdd.n5212 vdd.n5211 3.38568
R8645 vdd.n4927 vdd.n4926 3.38568
R8646 vdd.n4984 vdd.n4983 3.38568
R8647 vdd.n4699 vdd.n4698 3.38568
R8648 vdd.n4756 vdd.n4755 3.38568
R8649 vdd.n4027 vdd.n4026 3.38568
R8650 vdd.n2855 vdd.n2061 3.38568
R8651 vdd.n3609 vdd.n3608 3.38568
R8652 vdd.n3666 vdd.n3665 3.38568
R8653 vdd.n3381 vdd.n3380 3.38568
R8654 vdd.n3438 vdd.n3437 3.38568
R8655 vdd.n3153 vdd.n3152 3.38568
R8656 vdd.n3210 vdd.n3209 3.38568
R8657 vdd.n2925 vdd.n2924 3.38568
R8658 vdd.n2982 vdd.n2981 3.38568
R8659 vdd.n3763 vdd.n2258 3.38568
R8660 vdd.n3730 vdd.n3729 3.38568
R8661 vdd.n3546 vdd.n3545 3.38568
R8662 vdd.n3492 vdd.n2413 3.38568
R8663 vdd.n3318 vdd.n3317 3.38568
R8664 vdd.n3264 vdd.n2548 3.38568
R8665 vdd.n3090 vdd.n3089 3.38568
R8666 vdd.n3036 vdd.n2683 3.38568
R8667 vdd.n5539 vdd.n284 3.38568
R8668 vdd.n5506 vdd.n5505 3.38568
R8669 vdd.n5320 vdd.n5319 3.38568
R8670 vdd.n5266 vdd.n437 3.38568
R8671 vdd.n5092 vdd.n5091 3.38568
R8672 vdd.n5038 vdd.n572 3.38568
R8673 vdd.n4864 vdd.n4863 3.38568
R8674 vdd.n4810 vdd.n707 3.38568
R8675 vdd.n5679 vdd.n255 3.38568
R8676 vdd.n2176 vdd.n2108 3.35453
R8677 vdd.n6411 vdd.n6384 3.10353
R8678 vdd.n6410 vdd.n6375 3.10353
R8679 vdd.n6432 vdd.n6373 3.10353
R8680 vdd.n6431 vdd.n6360 3.10353
R8681 vdd.n6364 vdd.n6361 3.10353
R8682 vdd.n6459 vdd.n6358 3.10353
R8683 vdd.n6474 vdd.n6349 3.10353
R8684 vdd.n6475 vdd.n6347 3.10353
R8685 vdd.n6494 vdd.n6338 3.10353
R8686 vdd.n6495 vdd.n6327 3.10353
R8687 vdd.n6336 vdd.n6335 3.10353
R8688 vdd.n6328 vdd.n6317 3.10353
R8689 vdd.n6316 vdd.n6313 3.10353
R8690 vdd.n6523 vdd.n6522 3.10353
R8691 vdd.n6315 vdd.n6314 3.10353
R8692 vdd.n6548 vdd.n6300 3.10353
R8693 vdd.n6555 vdd.n6298 3.10353
R8694 vdd.n6556 vdd.n6282 3.10353
R8695 vdd.n6581 vdd.n6280 3.10353
R8696 vdd.n6285 vdd.n6279 3.10353
R8697 vdd.n6602 vdd.n6270 3.10353
R8698 vdd.n6601 vdd.n6267 3.10353
R8699 vdd.n6607 vdd.n6268 3.10353
R8700 vdd.n6606 vdd.n6253 3.10353
R8701 vdd.n6638 vdd.n6251 3.10353
R8702 vdd.n6637 vdd.n6242 3.10353
R8703 vdd.n6659 vdd.n6240 3.10353
R8704 vdd.n6658 vdd.n6227 3.10353
R8705 vdd.n6231 vdd.n6228 3.10353
R8706 vdd.n6686 vdd.n6225 3.10353
R8707 vdd.n6701 vdd.n6216 3.10353
R8708 vdd.n6702 vdd.n6214 3.10353
R8709 vdd.n6721 vdd.n6205 3.10353
R8710 vdd.n6722 vdd.n6194 3.10353
R8711 vdd.n6203 vdd.n6202 3.10353
R8712 vdd.n6195 vdd.n6184 3.10353
R8713 vdd.n6183 vdd.n6180 3.10353
R8714 vdd.n6750 vdd.n6749 3.10353
R8715 vdd.n6182 vdd.n6181 3.10353
R8716 vdd.n6775 vdd.n6167 3.10353
R8717 vdd.n6782 vdd.n6165 3.10353
R8718 vdd.n6783 vdd.n6149 3.10353
R8719 vdd.n6808 vdd.n6147 3.10353
R8720 vdd.n6152 vdd.n6146 3.10353
R8721 vdd.n6829 vdd.n6137 3.10353
R8722 vdd.n6828 vdd.n6134 3.10353
R8723 vdd.n6834 vdd.n6135 3.10353
R8724 vdd.n6833 vdd.n6120 3.10353
R8725 vdd.n6865 vdd.n6118 3.10353
R8726 vdd.n6864 vdd.n6109 3.10353
R8727 vdd.n6886 vdd.n6107 3.10353
R8728 vdd.n6885 vdd.n6094 3.10353
R8729 vdd.n6098 vdd.n6095 3.10353
R8730 vdd.n6913 vdd.n6092 3.10353
R8731 vdd.n6928 vdd.n6083 3.10353
R8732 vdd.n6929 vdd.n6081 3.10353
R8733 vdd.n6948 vdd.n6072 3.10353
R8734 vdd.n6949 vdd.n6061 3.10353
R8735 vdd.n6070 vdd.n6069 3.10353
R8736 vdd.n6062 vdd.n6051 3.10353
R8737 vdd.n6050 vdd.n6047 3.10353
R8738 vdd.n6977 vdd.n6976 3.10353
R8739 vdd.n6049 vdd.n6048 3.10353
R8740 vdd.n7002 vdd.n6034 3.10353
R8741 vdd.n7009 vdd.n6032 3.10353
R8742 vdd.n7010 vdd.n6016 3.10353
R8743 vdd.n7035 vdd.n6014 3.10353
R8744 vdd.n6019 vdd.n6013 3.10353
R8745 vdd.n7056 vdd.n6004 3.10353
R8746 vdd.n7055 vdd.n6001 3.10353
R8747 vdd.n7061 vdd.n6002 3.10353
R8748 vdd.n7060 vdd.n5987 3.10353
R8749 vdd.n7092 vdd.n5985 3.10353
R8750 vdd.n7091 vdd.n5976 3.10353
R8751 vdd.n7113 vdd.n5974 3.10353
R8752 vdd.n7112 vdd.n5961 3.10353
R8753 vdd.n5965 vdd.n5962 3.10353
R8754 vdd.n7140 vdd.n5959 3.10353
R8755 vdd.n7155 vdd.n5950 3.10353
R8756 vdd.n7156 vdd.n5948 3.10353
R8757 vdd.n7175 vdd.n5939 3.10353
R8758 vdd.n7176 vdd.n5928 3.10353
R8759 vdd.n5937 vdd.n5936 3.10353
R8760 vdd.n5929 vdd.n5918 3.10353
R8761 vdd.n5917 vdd.n5914 3.10353
R8762 vdd.n7204 vdd.n7203 3.10353
R8763 vdd.n5916 vdd.n5915 3.10353
R8764 vdd.n7229 vdd.n5901 3.10353
R8765 vdd.n7236 vdd.n5899 3.10353
R8766 vdd.n7237 vdd.n5883 3.10353
R8767 vdd.n7262 vdd.n5881 3.10353
R8768 vdd.n5886 vdd.n5880 3.10353
R8769 vdd.n7288 vdd.n5870 3.10353
R8770 vdd.n7287 vdd.n5868 3.10353
R8771 vdd.n7317 vdd.n5859 3.10353
R8772 vdd.n7316 vdd.n5857 3.10353
R8773 vdd.n7336 vdd.n5848 3.10353
R8774 vdd.n7335 vdd.n5846 3.10353
R8775 vdd.n7355 vdd.n5837 3.10353
R8776 vdd.n7354 vdd.n5835 3.10353
R8777 vdd.n7374 vdd.n5826 3.10353
R8778 vdd.n7373 vdd.n5824 3.10353
R8779 vdd.n7397 vdd.n5814 3.10353
R8780 vdd.n7396 vdd.n5799 3.10353
R8781 vdd.n5724 vdd.n5723 3.10353
R8782 vdd.n263 vdd.n262 3.10353
R8783 vdd.n5612 vdd.n265 3.10353
R8784 vdd.n5617 vdd.n5613 3.10353
R8785 vdd.n5622 vdd.n5621 3.10353
R8786 vdd.n5701 vdd.n5623 3.10353
R8787 vdd.n5698 vdd.n5696 3.10353
R8788 vdd.n5695 vdd.n5624 3.10353
R8789 vdd.n5670 vdd.n5667 3.10353
R8790 vdd.n5678 vdd.n5677 3.10353
R8791 vdd.n2919 vdd.n2775 3.10353
R8792 vdd.n2920 vdd.n2773 3.10353
R8793 vdd.n2949 vdd.n2762 3.10353
R8794 vdd.n2951 vdd.n2950 3.10353
R8795 vdd.n2958 vdd.n2759 3.10353
R8796 vdd.n2957 vdd.n2746 3.10353
R8797 vdd.n2750 vdd.n2747 3.10353
R8798 vdd.n2986 vdd.n2744 3.10353
R8799 vdd.n3002 vdd.n2735 3.10353
R8800 vdd.n3003 vdd.n2715 3.10353
R8801 vdd.n2733 vdd.n2732 3.10353
R8802 vdd.n2725 vdd.n2716 3.10353
R8803 vdd.n2720 vdd.n2719 3.10353
R8804 vdd.n3031 vdd.n2702 3.10353
R8805 vdd.n3038 vdd.n2700 3.10353
R8806 vdd.n3039 vdd.n2684 3.10353
R8807 vdd.n3064 vdd.n2682 3.10353
R8808 vdd.n2687 vdd.n2681 3.10353
R8809 vdd.n3087 vdd.n2668 3.10353
R8810 vdd.n3086 vdd.n2669 3.10353
R8811 vdd.n3094 vdd.n3093 3.10353
R8812 vdd.n3095 vdd.n2651 3.10353
R8813 vdd.n3128 vdd.n2649 3.10353
R8814 vdd.n3132 vdd.n3129 3.10353
R8815 vdd.n3147 vdd.n2640 3.10353
R8816 vdd.n3148 vdd.n2638 3.10353
R8817 vdd.n3177 vdd.n2627 3.10353
R8818 vdd.n3179 vdd.n3178 3.10353
R8819 vdd.n3186 vdd.n2624 3.10353
R8820 vdd.n3185 vdd.n2611 3.10353
R8821 vdd.n2615 vdd.n2612 3.10353
R8822 vdd.n3214 vdd.n2609 3.10353
R8823 vdd.n3230 vdd.n2600 3.10353
R8824 vdd.n3231 vdd.n2580 3.10353
R8825 vdd.n2598 vdd.n2597 3.10353
R8826 vdd.n2590 vdd.n2581 3.10353
R8827 vdd.n2585 vdd.n2584 3.10353
R8828 vdd.n3259 vdd.n2567 3.10353
R8829 vdd.n3266 vdd.n2565 3.10353
R8830 vdd.n3267 vdd.n2549 3.10353
R8831 vdd.n3292 vdd.n2547 3.10353
R8832 vdd.n2552 vdd.n2546 3.10353
R8833 vdd.n3315 vdd.n2533 3.10353
R8834 vdd.n3314 vdd.n2534 3.10353
R8835 vdd.n3322 vdd.n3321 3.10353
R8836 vdd.n3323 vdd.n2516 3.10353
R8837 vdd.n3356 vdd.n2514 3.10353
R8838 vdd.n3360 vdd.n3357 3.10353
R8839 vdd.n3375 vdd.n2505 3.10353
R8840 vdd.n3376 vdd.n2503 3.10353
R8841 vdd.n3405 vdd.n2492 3.10353
R8842 vdd.n3407 vdd.n3406 3.10353
R8843 vdd.n3414 vdd.n2489 3.10353
R8844 vdd.n3413 vdd.n2476 3.10353
R8845 vdd.n2480 vdd.n2477 3.10353
R8846 vdd.n3442 vdd.n2474 3.10353
R8847 vdd.n3458 vdd.n2465 3.10353
R8848 vdd.n3459 vdd.n2445 3.10353
R8849 vdd.n2463 vdd.n2462 3.10353
R8850 vdd.n2455 vdd.n2446 3.10353
R8851 vdd.n2450 vdd.n2449 3.10353
R8852 vdd.n3487 vdd.n2432 3.10353
R8853 vdd.n3494 vdd.n2430 3.10353
R8854 vdd.n3495 vdd.n2414 3.10353
R8855 vdd.n3520 vdd.n2412 3.10353
R8856 vdd.n2417 vdd.n2411 3.10353
R8857 vdd.n3543 vdd.n2398 3.10353
R8858 vdd.n3542 vdd.n2399 3.10353
R8859 vdd.n3550 vdd.n3549 3.10353
R8860 vdd.n3551 vdd.n2381 3.10353
R8861 vdd.n3584 vdd.n2379 3.10353
R8862 vdd.n3588 vdd.n3585 3.10353
R8863 vdd.n3603 vdd.n2370 3.10353
R8864 vdd.n3604 vdd.n2368 3.10353
R8865 vdd.n3633 vdd.n2357 3.10353
R8866 vdd.n3635 vdd.n3634 3.10353
R8867 vdd.n3642 vdd.n2354 3.10353
R8868 vdd.n3641 vdd.n2341 3.10353
R8869 vdd.n2345 vdd.n2342 3.10353
R8870 vdd.n3670 vdd.n2339 3.10353
R8871 vdd.n3685 vdd.n2330 3.10353
R8872 vdd.n3686 vdd.n2319 3.10353
R8873 vdd.n2328 vdd.n2327 3.10353
R8874 vdd.n2320 vdd.n2308 3.10353
R8875 vdd.n3708 vdd.n3707 3.10353
R8876 vdd.n3709 vdd.n2299 3.10353
R8877 vdd.n2297 vdd.n2292 3.10353
R8878 vdd.n3733 vdd.n3732 3.10353
R8879 vdd.n2294 vdd.n2293 3.10353
R8880 vdd.n3758 vdd.n2279 3.10353
R8881 vdd.n3765 vdd.n2277 3.10353
R8882 vdd.n3766 vdd.n2259 3.10353
R8883 vdd.n3795 vdd.n2257 3.10353
R8884 vdd.n2262 vdd.n2256 3.10353
R8885 vdd.n4016 vdd.n4009 3.10353
R8886 vdd.n4015 vdd.n2054 3.10353
R8887 vdd.n2827 vdd.n2055 3.10353
R8888 vdd.n2826 vdd.n2807 3.10353
R8889 vdd.n2808 vdd.n2805 3.10353
R8890 vdd.n2853 vdd.n2852 3.10353
R8891 vdd.n2870 vdd.n2796 3.10353
R8892 vdd.n2874 vdd.n2871 3.10353
R8893 vdd.n2877 vdd.n2875 3.10353
R8894 vdd.n2880 vdd.n2879 3.10353
R8895 vdd.n1024 vdd.n989 3.10353
R8896 vdd.n4520 vdd.n1006 3.10353
R8897 vdd.n1055 vdd.n1007 3.10353
R8898 vdd.n1061 vdd.n1056 3.10353
R8899 vdd.n1067 vdd.n1063 3.10353
R8900 vdd.n1068 vdd.n1049 3.10353
R8901 vdd.n1093 vdd.n1050 3.10353
R8902 vdd.n4493 vdd.n1074 3.10353
R8903 vdd.n1122 vdd.n1075 3.10353
R8904 vdd.n1126 vdd.n1125 3.10353
R8905 vdd.n1137 vdd.n1127 3.10353
R8906 vdd.n1130 vdd.n1117 3.10353
R8907 vdd.n4468 vdd.n1118 3.10353
R8908 vdd.n4467 vdd.n1144 3.10353
R8909 vdd.n1180 vdd.n1179 3.10353
R8910 vdd.n1178 vdd.n1167 3.10353
R8911 vdd.n4446 vdd.n1168 3.10353
R8912 vdd.n4445 vdd.n1186 3.10353
R8913 vdd.n1222 vdd.n1221 3.10353
R8914 vdd.n1220 vdd.n1209 3.10353
R8915 vdd.n4424 vdd.n1210 3.10353
R8916 vdd.n4423 vdd.n1228 3.10353
R8917 vdd.n1267 vdd.n1262 3.10353
R8918 vdd.n1268 vdd.n1257 3.10353
R8919 vdd.n1288 vdd.n1258 3.10353
R8920 vdd.n4399 vdd.n1274 3.10353
R8921 vdd.n1319 vdd.n1275 3.10353
R8922 vdd.n1325 vdd.n1320 3.10353
R8923 vdd.n1331 vdd.n1327 3.10353
R8924 vdd.n1332 vdd.n1313 3.10353
R8925 vdd.n1357 vdd.n1314 3.10353
R8926 vdd.n4372 vdd.n1338 3.10353
R8927 vdd.n1386 vdd.n1339 3.10353
R8928 vdd.n1390 vdd.n1389 3.10353
R8929 vdd.n1401 vdd.n1391 3.10353
R8930 vdd.n1394 vdd.n1381 3.10353
R8931 vdd.n4347 vdd.n1382 3.10353
R8932 vdd.n4346 vdd.n1408 3.10353
R8933 vdd.n1444 vdd.n1443 3.10353
R8934 vdd.n1442 vdd.n1431 3.10353
R8935 vdd.n4325 vdd.n1432 3.10353
R8936 vdd.n4324 vdd.n1450 3.10353
R8937 vdd.n1486 vdd.n1485 3.10353
R8938 vdd.n1484 vdd.n1473 3.10353
R8939 vdd.n4303 vdd.n1474 3.10353
R8940 vdd.n4302 vdd.n1492 3.10353
R8941 vdd.n1531 vdd.n1526 3.10353
R8942 vdd.n1532 vdd.n1521 3.10353
R8943 vdd.n1552 vdd.n1522 3.10353
R8944 vdd.n4278 vdd.n1538 3.10353
R8945 vdd.n1583 vdd.n1539 3.10353
R8946 vdd.n1589 vdd.n1584 3.10353
R8947 vdd.n1595 vdd.n1591 3.10353
R8948 vdd.n1596 vdd.n1577 3.10353
R8949 vdd.n1621 vdd.n1578 3.10353
R8950 vdd.n4251 vdd.n1602 3.10353
R8951 vdd.n1650 vdd.n1603 3.10353
R8952 vdd.n1654 vdd.n1653 3.10353
R8953 vdd.n1665 vdd.n1655 3.10353
R8954 vdd.n1658 vdd.n1645 3.10353
R8955 vdd.n4226 vdd.n1646 3.10353
R8956 vdd.n4225 vdd.n1672 3.10353
R8957 vdd.n1708 vdd.n1707 3.10353
R8958 vdd.n1706 vdd.n1695 3.10353
R8959 vdd.n4204 vdd.n1696 3.10353
R8960 vdd.n4203 vdd.n1714 3.10353
R8961 vdd.n1750 vdd.n1749 3.10353
R8962 vdd.n1748 vdd.n1737 3.10353
R8963 vdd.n4182 vdd.n1738 3.10353
R8964 vdd.n4181 vdd.n1756 3.10353
R8965 vdd.n1795 vdd.n1790 3.10353
R8966 vdd.n1796 vdd.n1785 3.10353
R8967 vdd.n1816 vdd.n1786 3.10353
R8968 vdd.n4157 vdd.n1802 3.10353
R8969 vdd.n1847 vdd.n1803 3.10353
R8970 vdd.n1853 vdd.n1848 3.10353
R8971 vdd.n1859 vdd.n1855 3.10353
R8972 vdd.n1860 vdd.n1841 3.10353
R8973 vdd.n1885 vdd.n1842 3.10353
R8974 vdd.n4130 vdd.n1866 3.10353
R8975 vdd.n1914 vdd.n1867 3.10353
R8976 vdd.n1918 vdd.n1917 3.10353
R8977 vdd.n1929 vdd.n1919 3.10353
R8978 vdd.n1922 vdd.n1909 3.10353
R8979 vdd.n4105 vdd.n1910 3.10353
R8980 vdd.n4104 vdd.n1936 3.10353
R8981 vdd.n1972 vdd.n1971 3.10353
R8982 vdd.n1970 vdd.n1959 3.10353
R8983 vdd.n4083 vdd.n1960 3.10353
R8984 vdd.n4082 vdd.n1978 3.10353
R8985 vdd.n2014 vdd.n2013 3.10353
R8986 vdd.n2012 vdd.n2001 3.10353
R8987 vdd.n4061 vdd.n2002 3.10353
R8988 vdd.n4060 vdd.n2020 3.10353
R8989 vdd.n897 vdd.n853 3.10353
R8990 vdd.n4572 vdd.n858 3.10353
R8991 vdd.n928 vdd.n859 3.10353
R8992 vdd.n934 vdd.n929 3.10353
R8993 vdd.n940 vdd.n936 3.10353
R8994 vdd.n941 vdd.n922 3.10353
R8995 vdd.n966 vdd.n923 3.10353
R8996 vdd.n4545 vdd.n947 3.10353
R8997 vdd.n994 vdd.n948 3.10353
R8998 vdd.n998 vdd.n997 3.10353
R8999 vdd.n4693 vdd.n799 3.10353
R9000 vdd.n4694 vdd.n797 3.10353
R9001 vdd.n4723 vdd.n786 3.10353
R9002 vdd.n4725 vdd.n4724 3.10353
R9003 vdd.n4732 vdd.n783 3.10353
R9004 vdd.n4731 vdd.n770 3.10353
R9005 vdd.n774 vdd.n771 3.10353
R9006 vdd.n4760 vdd.n768 3.10353
R9007 vdd.n4776 vdd.n759 3.10353
R9008 vdd.n4777 vdd.n739 3.10353
R9009 vdd.n757 vdd.n756 3.10353
R9010 vdd.n749 vdd.n740 3.10353
R9011 vdd.n744 vdd.n743 3.10353
R9012 vdd.n4805 vdd.n726 3.10353
R9013 vdd.n4812 vdd.n724 3.10353
R9014 vdd.n4813 vdd.n708 3.10353
R9015 vdd.n4838 vdd.n706 3.10353
R9016 vdd.n711 vdd.n705 3.10353
R9017 vdd.n4861 vdd.n692 3.10353
R9018 vdd.n4860 vdd.n693 3.10353
R9019 vdd.n4868 vdd.n4867 3.10353
R9020 vdd.n4869 vdd.n675 3.10353
R9021 vdd.n4902 vdd.n673 3.10353
R9022 vdd.n4906 vdd.n4903 3.10353
R9023 vdd.n4921 vdd.n664 3.10353
R9024 vdd.n4922 vdd.n662 3.10353
R9025 vdd.n4951 vdd.n651 3.10353
R9026 vdd.n4953 vdd.n4952 3.10353
R9027 vdd.n4960 vdd.n648 3.10353
R9028 vdd.n4959 vdd.n635 3.10353
R9029 vdd.n639 vdd.n636 3.10353
R9030 vdd.n4988 vdd.n633 3.10353
R9031 vdd.n5004 vdd.n624 3.10353
R9032 vdd.n5005 vdd.n604 3.10353
R9033 vdd.n622 vdd.n621 3.10353
R9034 vdd.n614 vdd.n605 3.10353
R9035 vdd.n609 vdd.n608 3.10353
R9036 vdd.n5033 vdd.n591 3.10353
R9037 vdd.n5040 vdd.n589 3.10353
R9038 vdd.n5041 vdd.n573 3.10353
R9039 vdd.n5066 vdd.n571 3.10353
R9040 vdd.n576 vdd.n570 3.10353
R9041 vdd.n5089 vdd.n557 3.10353
R9042 vdd.n5088 vdd.n558 3.10353
R9043 vdd.n5096 vdd.n5095 3.10353
R9044 vdd.n5097 vdd.n540 3.10353
R9045 vdd.n5130 vdd.n538 3.10353
R9046 vdd.n5134 vdd.n5131 3.10353
R9047 vdd.n5149 vdd.n529 3.10353
R9048 vdd.n5150 vdd.n527 3.10353
R9049 vdd.n5179 vdd.n516 3.10353
R9050 vdd.n5181 vdd.n5180 3.10353
R9051 vdd.n5188 vdd.n513 3.10353
R9052 vdd.n5187 vdd.n500 3.10353
R9053 vdd.n504 vdd.n501 3.10353
R9054 vdd.n5216 vdd.n498 3.10353
R9055 vdd.n5232 vdd.n489 3.10353
R9056 vdd.n5233 vdd.n469 3.10353
R9057 vdd.n487 vdd.n486 3.10353
R9058 vdd.n479 vdd.n470 3.10353
R9059 vdd.n474 vdd.n473 3.10353
R9060 vdd.n5261 vdd.n456 3.10353
R9061 vdd.n5268 vdd.n454 3.10353
R9062 vdd.n5269 vdd.n438 3.10353
R9063 vdd.n5294 vdd.n436 3.10353
R9064 vdd.n441 vdd.n435 3.10353
R9065 vdd.n5317 vdd.n422 3.10353
R9066 vdd.n5316 vdd.n423 3.10353
R9067 vdd.n5324 vdd.n5323 3.10353
R9068 vdd.n5325 vdd.n405 3.10353
R9069 vdd.n5358 vdd.n403 3.10353
R9070 vdd.n5362 vdd.n5359 3.10353
R9071 vdd.n5377 vdd.n394 3.10353
R9072 vdd.n5378 vdd.n392 3.10353
R9073 vdd.n5407 vdd.n381 3.10353
R9074 vdd.n5409 vdd.n5408 3.10353
R9075 vdd.n5416 vdd.n378 3.10353
R9076 vdd.n5415 vdd.n365 3.10353
R9077 vdd.n369 vdd.n366 3.10353
R9078 vdd.n5444 vdd.n363 3.10353
R9079 vdd.n5459 vdd.n354 3.10353
R9080 vdd.n5460 vdd.n343 3.10353
R9081 vdd.n352 vdd.n351 3.10353
R9082 vdd.n344 vdd.n333 3.10353
R9083 vdd.n5483 vdd.n5482 3.10353
R9084 vdd.n5484 vdd.n325 3.10353
R9085 vdd.n323 vdd.n318 3.10353
R9086 vdd.n5509 vdd.n5508 3.10353
R9087 vdd.n320 vdd.n319 3.10353
R9088 vdd.n5534 vdd.n305 3.10353
R9089 vdd.n5541 vdd.n303 3.10353
R9090 vdd.n5542 vdd.n285 3.10353
R9091 vdd.n5571 vdd.n283 3.10353
R9092 vdd.n288 vdd.n282 3.10353
R9093 vdd.n197 vdd.n196 3.03311
R9094 vdd.n3863 vdd.n3856 3.03311
R9095 vdd.n4616 vdd.n4586 3.03311
R9096 vdd.n223 vdd.n222 3.03311
R9097 vdd.n2173 vdd.n2168 2.91297
R9098 vdd.n5811 vdd 2.90898
R9099 vdd.n812 vdd 2.90898
R9100 vdd.n3922 vdd.t25 2.83209
R9101 vdd.n7505 vdd.n7504 2.64177
R9102 vdd.n3858 vdd.n3856 2.64177
R9103 vdd.n4607 vdd.n4586 2.64177
R9104 vdd.n225 vdd.n224 2.64177
R9105 vdd.n5725 vdd.n261 2.54483
R9106 vdd.n2896 vdd.n2786 2.54336
R9107 vdd.n999 vdd.n953 2.54336
R9108 vdd.n7302 vdd.n7301 2.5429
R9109 vdd.n7449 vdd 2.54117
R9110 vdd.n7488 vdd.n196 2.4386
R9111 vdd.n3982 vdd.n3866 2.4386
R9112 vdd.n4624 vdd.n846 2.4386
R9113 vdd.n5755 vdd.n223 2.4386
R9114 vdd.n48 vdd 2.39764
R9115 vdd.n52 vdd.n49 2.36813
R9116 vdd.n163 vdd.n162 2.3255
R9117 vdd.n178 vdd.n177 2.3255
R9118 vdd.n173 vdd.n172 2.3255
R9119 vdd.n165 vdd.n19 2.3255
R9120 vdd.n18 vdd.n17 2.3255
R9121 vdd.n9 vdd.n8 2.3255
R9122 vdd.n5800 vdd.n5790 2.28608
R9123 vdd.n5729 vdd.n248 2.28608
R9124 vdd.n4023 vdd.n4022 2.28608
R9125 vdd.n4580 vdd.n4579 2.28608
R9126 vdd.n7460 vdd.n230 2.24869
R9127 vdd.n236 vdd.n229 2.24869
R9128 vdd.n5744 vdd.n5743 2.24869
R9129 vdd.n7437 vdd.n7434 2.24869
R9130 vdd.n7445 vdd.n7444 2.24869
R9131 vdd.n5783 vdd.n5782 2.24869
R9132 vdd.n7426 vdd.n5789 2.24869
R9133 vdd.n5810 vdd.n5803 2.24869
R9134 vdd.n4664 vdd.n4663 2.24869
R9135 vdd.n4651 vdd.n4645 2.24869
R9136 vdd.n4656 vdd.n4655 2.24869
R9137 vdd.n4641 vdd.n4637 2.24869
R9138 vdd.n826 vdd.n820 2.24869
R9139 vdd.n3808 vdd.n3807 2.24858
R9140 vdd.n2244 vdd.n2243 2.24858
R9141 vdd.n3824 vdd.n3823 2.24858
R9142 vdd.n2233 vdd.n2232 2.24858
R9143 vdd.n3833 vdd.n3832 2.24858
R9144 vdd.n2090 vdd.n2080 2.24858
R9145 vdd.n3819 vdd.n3818 2.24858
R9146 vdd.n3962 vdd.n3947 2.24858
R9147 vdd.n3956 vdd.n3948 2.24858
R9148 vdd.n3975 vdd.n3974 2.24858
R9149 vdd.n3925 vdd.n3924 2.24858
R9150 vdd.n3885 vdd.n3884 2.24858
R9151 vdd.n3878 vdd.n3870 2.24858
R9152 vdd.n3942 vdd.n3941 2.24858
R9153 vdd.n3933 vdd.n3932 2.24858
R9154 vdd.n7423 vdd.n5790 2.15377
R9155 vdd.n5730 vdd.n5729 2.15377
R9156 vdd.n3822 vdd.n2079 2.09301
R9157 vdd.n4023 vdd.n4008 2.03414
R9158 vdd.n4580 vdd.n850 2.03414
R9159 vdd.n7425 vdd.n7424 1.99051
R9160 vdd.n827 vdd.n247 1.99051
R9161 vdd.n5581 vdd 1.98118
R9162 vdd.n104 vdd.n101 1.97988
R9163 vdd.n5582 vdd 1.9603
R9164 vdd.n7492 vdd.n7491 1.94045
R9165 vdd.n7515 vdd.n7514 1.94045
R9166 vdd.n7421 vdd.n7420 1.94045
R9167 vdd.n5733 vdd.n5732 1.94045
R9168 vdd.n4011 vdd.n2038 1.94045
R9169 vdd.n883 vdd.n882 1.94045
R9170 vdd.n3986 vdd.n3985 1.94045
R9171 vdd.n3999 vdd.n3998 1.94045
R9172 vdd.n4628 vdd.n4627 1.94045
R9173 vdd.n4606 vdd.n4605 1.94045
R9174 vdd.n7477 vdd.n7476 1.94045
R9175 vdd.n5751 vdd.n5750 1.94045
R9176 vdd.n5736 vdd 1.7865
R9177 vdd.n7201 vdd.n7200 1.76521
R9178 vdd.n7263 vdd.n5882 1.76521
R9179 vdd.n7088 vdd.n5986 1.76521
R9180 vdd.n7109 vdd.n5975 1.76521
R9181 vdd.n7136 vdd.n5960 1.76521
R9182 vdd.n7139 vdd.n5949 1.76521
R9183 vdd.n7160 vdd.n7159 1.76521
R9184 vdd.n6974 vdd.n6973 1.76521
R9185 vdd.n7036 vdd.n6015 1.76521
R9186 vdd.n7064 vdd.n7063 1.76521
R9187 vdd.n6861 vdd.n6119 1.76521
R9188 vdd.n6882 vdd.n6108 1.76521
R9189 vdd.n6909 vdd.n6093 1.76521
R9190 vdd.n6912 vdd.n6082 1.76521
R9191 vdd.n6933 vdd.n6932 1.76521
R9192 vdd.n6747 vdd.n6746 1.76521
R9193 vdd.n6809 vdd.n6148 1.76521
R9194 vdd.n6837 vdd.n6836 1.76521
R9195 vdd.n6634 vdd.n6252 1.76521
R9196 vdd.n6655 vdd.n6241 1.76521
R9197 vdd.n6682 vdd.n6226 1.76521
R9198 vdd.n6685 vdd.n6215 1.76521
R9199 vdd.n6706 vdd.n6705 1.76521
R9200 vdd.n6520 vdd.n6519 1.76521
R9201 vdd.n6582 vdd.n6281 1.76521
R9202 vdd.n6610 vdd.n6609 1.76521
R9203 vdd.n6455 vdd.n6359 1.76521
R9204 vdd.n6458 vdd.n6348 1.76521
R9205 vdd.n6479 vdd.n6478 1.76521
R9206 vdd.n7300 vdd.n7299 1.76521
R9207 vdd.n7400 vdd.n5801 1.76521
R9208 vdd.n5726 vdd.n260 1.76521
R9209 vdd.n5679 vdd.n249 1.76521
R9210 vdd.n5481 vdd.n5479 1.76521
R9211 vdd.n5506 vdd.n322 1.76521
R9212 vdd.n5572 vdd.n284 1.76521
R9213 vdd.n5361 vdd.n393 1.76521
R9214 vdd.n5383 vdd.n5381 1.76521
R9215 vdd.n5439 vdd.n364 1.76521
R9216 vdd.n5464 vdd.n5463 1.76521
R9217 vdd.n477 vdd.n476 1.76521
R9218 vdd.n5295 vdd.n437 1.76521
R9219 vdd.n5322 vdd.n5320 1.76521
R9220 vdd.n5133 vdd.n528 1.76521
R9221 vdd.n5155 vdd.n5153 1.76521
R9222 vdd.n5211 vdd.n499 1.76521
R9223 vdd.n5237 vdd.n5236 1.76521
R9224 vdd.n612 vdd.n611 1.76521
R9225 vdd.n5067 vdd.n572 1.76521
R9226 vdd.n5094 vdd.n5092 1.76521
R9227 vdd.n4905 vdd.n663 1.76521
R9228 vdd.n4927 vdd.n4925 1.76521
R9229 vdd.n4983 vdd.n634 1.76521
R9230 vdd.n5009 vdd.n5008 1.76521
R9231 vdd.n747 vdd.n746 1.76521
R9232 vdd.n4839 vdd.n707 1.76521
R9233 vdd.n4866 vdd.n4864 1.76521
R9234 vdd.n4699 vdd.n4697 1.76521
R9235 vdd.n4755 vdd.n769 1.76521
R9236 vdd.n4781 vdd.n4780 1.76521
R9237 vdd.n4577 vdd.n852 1.76521
R9238 vdd.n4573 vdd.n857 1.76521
R9239 vdd.n933 vdd.n927 1.76521
R9240 vdd.n4550 vdd.n924 1.76521
R9241 vdd.n4546 vdd.n946 1.76521
R9242 vdd.n1000 vdd.n993 1.76521
R9243 vdd.n4110 vdd.n1911 1.76521
R9244 vdd.n1973 vdd.n1935 1.76521
R9245 vdd.n4088 vdd.n1962 1.76521
R9246 vdd.n2015 vdd.n1977 1.76521
R9247 vdd.n4066 vdd.n2004 1.76521
R9248 vdd.n3918 vdd.n2019 1.76521
R9249 vdd.n4162 vdd.n1787 1.76521
R9250 vdd.n4158 vdd.n1801 1.76521
R9251 vdd.n1852 vdd.n1846 1.76521
R9252 vdd.n4135 vdd.n1843 1.76521
R9253 vdd.n4131 vdd.n1865 1.76521
R9254 vdd.n1931 vdd.n1913 1.76521
R9255 vdd.n4231 vdd.n1647 1.76521
R9256 vdd.n1709 vdd.n1671 1.76521
R9257 vdd.n4209 vdd.n1698 1.76521
R9258 vdd.n1751 vdd.n1713 1.76521
R9259 vdd.n4187 vdd.n1740 1.76521
R9260 vdd.n1791 vdd.n1755 1.76521
R9261 vdd.n4283 vdd.n1523 1.76521
R9262 vdd.n4279 vdd.n1537 1.76521
R9263 vdd.n1588 vdd.n1582 1.76521
R9264 vdd.n4256 vdd.n1579 1.76521
R9265 vdd.n4252 vdd.n1601 1.76521
R9266 vdd.n1667 vdd.n1649 1.76521
R9267 vdd.n4352 vdd.n1383 1.76521
R9268 vdd.n1445 vdd.n1407 1.76521
R9269 vdd.n4330 vdd.n1434 1.76521
R9270 vdd.n1487 vdd.n1449 1.76521
R9271 vdd.n4308 vdd.n1476 1.76521
R9272 vdd.n1527 vdd.n1491 1.76521
R9273 vdd.n4404 vdd.n1259 1.76521
R9274 vdd.n4400 vdd.n1273 1.76521
R9275 vdd.n1324 vdd.n1318 1.76521
R9276 vdd.n4377 vdd.n1315 1.76521
R9277 vdd.n4373 vdd.n1337 1.76521
R9278 vdd.n1403 vdd.n1385 1.76521
R9279 vdd.n4473 vdd.n1119 1.76521
R9280 vdd.n1181 vdd.n1143 1.76521
R9281 vdd.n4451 vdd.n1170 1.76521
R9282 vdd.n1223 vdd.n1185 1.76521
R9283 vdd.n4429 vdd.n1212 1.76521
R9284 vdd.n1263 vdd.n1227 1.76521
R9285 vdd.n4525 vdd.n990 1.76521
R9286 vdd.n4521 vdd.n1005 1.76521
R9287 vdd.n1060 vdd.n1054 1.76521
R9288 vdd.n4498 vdd.n1051 1.76521
R9289 vdd.n4494 vdd.n1073 1.76521
R9290 vdd.n1139 vdd.n1121 1.76521
R9291 vdd.n2067 vdd.n2066 1.76521
R9292 vdd.n4027 vdd.n2056 1.76521
R9293 vdd.n2855 vdd.n2854 1.76521
R9294 vdd.n2878 vdd.n2064 1.76521
R9295 vdd.n3706 vdd.n3704 1.76521
R9296 vdd.n3730 vdd.n2296 1.76521
R9297 vdd.n3796 vdd.n2258 1.76521
R9298 vdd.n3587 vdd.n2369 1.76521
R9299 vdd.n3609 vdd.n3607 1.76521
R9300 vdd.n3665 vdd.n2340 1.76521
R9301 vdd.n3690 vdd.n3689 1.76521
R9302 vdd.n2453 vdd.n2452 1.76521
R9303 vdd.n3521 vdd.n2413 1.76521
R9304 vdd.n3548 vdd.n3546 1.76521
R9305 vdd.n3359 vdd.n2504 1.76521
R9306 vdd.n3381 vdd.n3379 1.76521
R9307 vdd.n3437 vdd.n2475 1.76521
R9308 vdd.n3463 vdd.n3462 1.76521
R9309 vdd.n2588 vdd.n2587 1.76521
R9310 vdd.n3293 vdd.n2548 1.76521
R9311 vdd.n3320 vdd.n3318 1.76521
R9312 vdd.n3131 vdd.n2639 1.76521
R9313 vdd.n3153 vdd.n3151 1.76521
R9314 vdd.n3209 vdd.n2610 1.76521
R9315 vdd.n3235 vdd.n3234 1.76521
R9316 vdd.n2723 vdd.n2722 1.76521
R9317 vdd.n3065 vdd.n2683 1.76521
R9318 vdd.n3092 vdd.n3090 1.76521
R9319 vdd.n2925 vdd.n2923 1.76521
R9320 vdd.n2981 vdd.n2745 1.76521
R9321 vdd.n3007 vdd.n3006 1.76521
R9322 vdd.n5737 vdd 1.76349
R9323 vdd.n2197 vdd.n2183 1.75828
R9324 vdd.n2195 vdd.n2194 1.75828
R9325 vdd.n2219 vdd.n2218 1.70997
R9326 vdd.n2226 vdd.n2225 1.706
R9327 vdd.n2220 vdd.n2094 1.70524
R9328 vdd.n2142 vdd.n2119 1.70524
R9329 vdd.t75 vdd.n5811 1.68435
R9330 vdd.n812 vdd.t86 1.68435
R9331 vdd.n7319 vdd.n5847 1.66612
R9332 vdd.n7338 vdd.n5836 1.66612
R9333 vdd.n7357 vdd.n5825 1.66612
R9334 vdd.n7376 vdd.n5813 1.66612
R9335 vdd.n6515 vdd.n6514 1.66612
R9336 vdd.n6552 vdd.n6551 1.66612
R9337 vdd.n6585 vdd.n6269 1.66612
R9338 vdd.n6742 vdd.n6741 1.66612
R9339 vdd.n6779 vdd.n6778 1.66612
R9340 vdd.n6812 vdd.n6136 1.66612
R9341 vdd.n6969 vdd.n6968 1.66612
R9342 vdd.n7006 vdd.n7005 1.66612
R9343 vdd.n7039 vdd.n6003 1.66612
R9344 vdd.n7196 vdd.n7195 1.66612
R9345 vdd.n7233 vdd.n7232 1.66612
R9346 vdd.n7266 vdd.n5869 1.66612
R9347 vdd.n7179 vdd.n7178 1.66612
R9348 vdd.n6952 vdd.n6951 1.66612
R9349 vdd.n6725 vdd.n6724 1.66612
R9350 vdd.n6498 vdd.n6497 1.66612
R9351 vdd.n6408 vdd.n6374 1.66612
R9352 vdd.n264 vdd.n258 1.66612
R9353 vdd.n5620 vdd.n252 1.66612
R9354 vdd.n5697 vdd.n256 1.66612
R9355 vdd.n5668 vdd.n254 1.66612
R9356 vdd.n5411 vdd.n5410 1.66612
R9357 vdd.n5443 vdd.n5442 1.66612
R9358 vdd.n5183 vdd.n5182 1.66612
R9359 vdd.n5215 vdd.n5214 1.66612
R9360 vdd.n4955 vdd.n4954 1.66612
R9361 vdd.n4987 vdd.n4986 1.66612
R9362 vdd.n4727 vdd.n4726 1.66612
R9363 vdd.n4759 vdd.n4758 1.66612
R9364 vdd.n2806 vdd.n2059 1.66612
R9365 vdd.n2873 vdd.n2062 1.66612
R9366 vdd.n3637 vdd.n3636 1.66612
R9367 vdd.n3669 vdd.n3668 1.66612
R9368 vdd.n3409 vdd.n3408 1.66612
R9369 vdd.n3441 vdd.n3440 1.66612
R9370 vdd.n3181 vdd.n3180 1.66612
R9371 vdd.n3213 vdd.n3212 1.66612
R9372 vdd.n2953 vdd.n2952 1.66612
R9373 vdd.n2985 vdd.n2984 1.66612
R9374 vdd.n3035 vdd.n3034 1.66612
R9375 vdd.n3068 vdd.n2667 1.66612
R9376 vdd.n3263 vdd.n3262 1.66612
R9377 vdd.n3296 vdd.n2532 1.66612
R9378 vdd.n3491 vdd.n3490 1.66612
R9379 vdd.n3524 vdd.n2397 1.66612
R9380 vdd.n3727 vdd.n3726 1.66612
R9381 vdd.n3762 vdd.n3761 1.66612
R9382 vdd.n3582 vdd.n3581 1.66612
R9383 vdd.n3354 vdd.n3353 1.66612
R9384 vdd.n3126 vdd.n3125 1.66612
R9385 vdd.n4809 vdd.n4808 1.66612
R9386 vdd.n4842 vdd.n691 1.66612
R9387 vdd.n5037 vdd.n5036 1.66612
R9388 vdd.n5070 vdd.n556 1.66612
R9389 vdd.n5265 vdd.n5264 1.66612
R9390 vdd.n5298 vdd.n421 1.66612
R9391 vdd.n5503 vdd.n5502 1.66612
R9392 vdd.n5538 vdd.n5537 1.66612
R9393 vdd.n5356 vdd.n5355 1.66612
R9394 vdd.n5128 vdd.n5127 1.66612
R9395 vdd.n4900 vdd.n4899 1.66612
R9396 vdd.t52 vdd.t50 1.53772
R9397 vdd.t9 vdd.t60 1.53772
R9398 vdd vdd.n11 1.42907
R9399 vdd.n7501 vdd.n7500 1.35607
R9400 vdd.n6613 vdd.n6612 1.35607
R9401 vdd.n6579 vdd.n6284 1.35607
R9402 vdd.n6304 vdd.n6303 1.35607
R9403 vdd.n6512 vdd.n6511 1.35607
R9404 vdd.n6297 vdd.n6295 1.35607
R9405 vdd.n6589 vdd.n6588 1.35607
R9406 vdd.n6840 vdd.n6839 1.35607
R9407 vdd.n6806 vdd.n6151 1.35607
R9408 vdd.n6171 vdd.n6170 1.35607
R9409 vdd.n6739 vdd.n6738 1.35607
R9410 vdd.n6164 vdd.n6162 1.35607
R9411 vdd.n6816 vdd.n6815 1.35607
R9412 vdd.n7067 vdd.n7066 1.35607
R9413 vdd.n7033 vdd.n6018 1.35607
R9414 vdd.n6038 vdd.n6037 1.35607
R9415 vdd.n6966 vdd.n6965 1.35607
R9416 vdd.n6031 vdd.n6029 1.35607
R9417 vdd.n7043 vdd.n7042 1.35607
R9418 vdd.n7260 vdd.n5885 1.35607
R9419 vdd.n5905 vdd.n5904 1.35607
R9420 vdd.n7193 vdd.n7192 1.35607
R9421 vdd.n5898 vdd.n5896 1.35607
R9422 vdd.n7270 vdd.n7269 1.35607
R9423 vdd.n7163 vdd.n7162 1.35607
R9424 vdd.n7143 vdd.n7142 1.35607
R9425 vdd.n7134 vdd.n5964 1.35607
R9426 vdd.n6936 vdd.n6935 1.35607
R9427 vdd.n6916 vdd.n6915 1.35607
R9428 vdd.n6907 vdd.n6097 1.35607
R9429 vdd.n6709 vdd.n6708 1.35607
R9430 vdd.n6689 vdd.n6688 1.35607
R9431 vdd.n6680 vdd.n6230 1.35607
R9432 vdd.n6482 vdd.n6481 1.35607
R9433 vdd.n6462 vdd.n6461 1.35607
R9434 vdd.n7403 vdd.n7402 1.35607
R9435 vdd.n3857 vdd.n3846 1.35607
R9436 vdd.n4589 vdd.n4587 1.35607
R9437 vdd.n5499 vdd.n5498 1.35607
R9438 vdd.n309 vdd.n308 1.35607
R9439 vdd.n302 vdd.n300 1.35607
R9440 vdd.n5569 vdd.n287 1.35607
R9441 vdd.n5477 vdd.n5476 1.35607
R9442 vdd.n5386 vdd.n5385 1.35607
R9443 vdd.n5399 vdd.n5398 1.35607
R9444 vdd.n5437 vdd.n368 1.35607
R9445 vdd.n5447 vdd.n5446 1.35607
R9446 vdd.n5365 vdd.n5364 1.35607
R9447 vdd.n453 vdd.n451 1.35607
R9448 vdd.n5292 vdd.n440 1.35607
R9449 vdd.n5302 vdd.n5301 1.35607
R9450 vdd.n419 vdd.n417 1.35607
R9451 vdd.n460 vdd.n459 1.35607
R9452 vdd.n5158 vdd.n5157 1.35607
R9453 vdd.n5171 vdd.n5170 1.35607
R9454 vdd.n5209 vdd.n503 1.35607
R9455 vdd.n5219 vdd.n5218 1.35607
R9456 vdd.n5137 vdd.n5136 1.35607
R9457 vdd.n588 vdd.n586 1.35607
R9458 vdd.n5064 vdd.n575 1.35607
R9459 vdd.n5074 vdd.n5073 1.35607
R9460 vdd.n554 vdd.n552 1.35607
R9461 vdd.n595 vdd.n594 1.35607
R9462 vdd.n4930 vdd.n4929 1.35607
R9463 vdd.n4943 vdd.n4942 1.35607
R9464 vdd.n4981 vdd.n638 1.35607
R9465 vdd.n4991 vdd.n4990 1.35607
R9466 vdd.n4909 vdd.n4908 1.35607
R9467 vdd.n723 vdd.n721 1.35607
R9468 vdd.n4836 vdd.n710 1.35607
R9469 vdd.n4846 vdd.n4845 1.35607
R9470 vdd.n689 vdd.n687 1.35607
R9471 vdd.n730 vdd.n729 1.35607
R9472 vdd.n4715 vdd.n4714 1.35607
R9473 vdd.n4753 vdd.n773 1.35607
R9474 vdd.n4763 vdd.n4762 1.35607
R9475 vdd.n6426 vdd.n6425 1.35607
R9476 vdd.n7292 vdd.n5867 1.35607
R9477 vdd.n7107 vdd.n7106 1.35607
R9478 vdd.n7182 vdd.n7181 1.35607
R9479 vdd.n7086 vdd.n7085 1.35607
R9480 vdd.n6880 vdd.n6879 1.35607
R9481 vdd.n6955 vdd.n6954 1.35607
R9482 vdd.n6859 vdd.n6858 1.35607
R9483 vdd.n6653 vdd.n6652 1.35607
R9484 vdd.n6728 vdd.n6727 1.35607
R9485 vdd.n6632 vdd.n6631 1.35607
R9486 vdd.n6453 vdd.n6363 1.35607
R9487 vdd.n6501 vdd.n6500 1.35607
R9488 vdd.n6405 vdd.n6404 1.35607
R9489 vdd.n7380 vdd.n7379 1.35607
R9490 vdd.n7361 vdd.n7360 1.35607
R9491 vdd.n7342 vdd.n7341 1.35607
R9492 vdd.n7323 vdd.n7322 1.35607
R9493 vdd.n5608 vdd.n5606 1.35607
R9494 vdd.n5611 vdd.n5610 1.35607
R9495 vdd.n5691 vdd.n5626 1.35607
R9496 vdd.n5682 vdd.n5681 1.35607
R9497 vdd.n5719 vdd.n267 1.35607
R9498 vdd.n2907 vdd.n2906 1.35607
R9499 vdd.n3723 vdd.n3722 1.35607
R9500 vdd.n2283 vdd.n2282 1.35607
R9501 vdd.n2276 vdd.n2274 1.35607
R9502 vdd.n3793 vdd.n2261 1.35607
R9503 vdd.n3801 vdd.n2255 1.35607
R9504 vdd.n3702 vdd.n3701 1.35607
R9505 vdd.n3612 vdd.n3611 1.35607
R9506 vdd.n3625 vdd.n3624 1.35607
R9507 vdd.n3663 vdd.n2344 1.35607
R9508 vdd.n3673 vdd.n3672 1.35607
R9509 vdd.n3693 vdd.n3692 1.35607
R9510 vdd.n3591 vdd.n3590 1.35607
R9511 vdd.n2429 vdd.n2427 1.35607
R9512 vdd.n3518 vdd.n2416 1.35607
R9513 vdd.n3528 vdd.n3527 1.35607
R9514 vdd.n2395 vdd.n2393 1.35607
R9515 vdd.n3578 vdd.n2383 1.35607
R9516 vdd.n2436 vdd.n2435 1.35607
R9517 vdd.n3384 vdd.n3383 1.35607
R9518 vdd.n3397 vdd.n3396 1.35607
R9519 vdd.n3435 vdd.n2479 1.35607
R9520 vdd.n3445 vdd.n3444 1.35607
R9521 vdd.n3466 vdd.n3465 1.35607
R9522 vdd.n3363 vdd.n3362 1.35607
R9523 vdd.n2564 vdd.n2562 1.35607
R9524 vdd.n3290 vdd.n2551 1.35607
R9525 vdd.n3300 vdd.n3299 1.35607
R9526 vdd.n2530 vdd.n2528 1.35607
R9527 vdd.n3350 vdd.n2518 1.35607
R9528 vdd.n2571 vdd.n2570 1.35607
R9529 vdd.n3156 vdd.n3155 1.35607
R9530 vdd.n3169 vdd.n3168 1.35607
R9531 vdd.n3207 vdd.n2614 1.35607
R9532 vdd.n3217 vdd.n3216 1.35607
R9533 vdd.n3238 vdd.n3237 1.35607
R9534 vdd.n3135 vdd.n3134 1.35607
R9535 vdd.n2699 vdd.n2697 1.35607
R9536 vdd.n3062 vdd.n2686 1.35607
R9537 vdd.n3072 vdd.n3071 1.35607
R9538 vdd.n2665 vdd.n2663 1.35607
R9539 vdd.n3122 vdd.n2653 1.35607
R9540 vdd.n2706 vdd.n2705 1.35607
R9541 vdd.n2941 vdd.n2940 1.35607
R9542 vdd.n2979 vdd.n2749 1.35607
R9543 vdd.n2989 vdd.n2988 1.35607
R9544 vdd.n3010 vdd.n3009 1.35607
R9545 vdd.n2928 vdd.n2927 1.35607
R9546 vdd.n4020 vdd.n4013 1.35607
R9547 vdd.n4029 vdd.n2052 1.35607
R9548 vdd.n2848 vdd.n2810 1.35607
R9549 vdd.n2858 vdd.n2857 1.35607
R9550 vdd.n2885 vdd.n2884 1.35607
R9551 vdd.n4527 vdd.n986 1.35607
R9552 vdd.n4100 vdd.n1938 1.35607
R9553 vdd.n4091 vdd.n4090 1.35607
R9554 vdd.n4078 vdd.n1980 1.35607
R9555 vdd.n4069 vdd.n4068 1.35607
R9556 vdd.n4056 vdd.n2022 1.35607
R9557 vdd.n4113 vdd.n4112 1.35607
R9558 vdd.n4155 vdd.n1805 1.35607
R9559 vdd.n1809 vdd.n1808 1.35607
R9560 vdd.n4137 vdd.n1839 1.35607
R9561 vdd.n4128 vdd.n1869 1.35607
R9562 vdd.n1873 vdd.n1872 1.35607
R9563 vdd.n4165 vdd.n4164 1.35607
R9564 vdd.n4221 vdd.n1674 1.35607
R9565 vdd.n4212 vdd.n4211 1.35607
R9566 vdd.n4199 vdd.n1716 1.35607
R9567 vdd.n4190 vdd.n4189 1.35607
R9568 vdd.n4177 vdd.n1758 1.35607
R9569 vdd.n4234 vdd.n4233 1.35607
R9570 vdd.n4276 vdd.n1541 1.35607
R9571 vdd.n1545 vdd.n1544 1.35607
R9572 vdd.n4258 vdd.n1575 1.35607
R9573 vdd.n4249 vdd.n1605 1.35607
R9574 vdd.n1609 vdd.n1608 1.35607
R9575 vdd.n4286 vdd.n4285 1.35607
R9576 vdd.n4342 vdd.n1410 1.35607
R9577 vdd.n4333 vdd.n4332 1.35607
R9578 vdd.n4320 vdd.n1452 1.35607
R9579 vdd.n4311 vdd.n4310 1.35607
R9580 vdd.n4298 vdd.n1494 1.35607
R9581 vdd.n4355 vdd.n4354 1.35607
R9582 vdd.n4397 vdd.n1277 1.35607
R9583 vdd.n1281 vdd.n1280 1.35607
R9584 vdd.n4379 vdd.n1311 1.35607
R9585 vdd.n4370 vdd.n1341 1.35607
R9586 vdd.n1345 vdd.n1344 1.35607
R9587 vdd.n4407 vdd.n4406 1.35607
R9588 vdd.n4463 vdd.n1146 1.35607
R9589 vdd.n4454 vdd.n4453 1.35607
R9590 vdd.n4441 vdd.n1188 1.35607
R9591 vdd.n4432 vdd.n4431 1.35607
R9592 vdd.n4419 vdd.n1230 1.35607
R9593 vdd.n4476 vdd.n4475 1.35607
R9594 vdd.n1013 vdd.n1012 1.35607
R9595 vdd.n4500 vdd.n1047 1.35607
R9596 vdd.n4491 vdd.n1077 1.35607
R9597 vdd.n1081 vdd.n1080 1.35607
R9598 vdd.n4518 vdd.n1009 1.35607
R9599 vdd.n894 vdd.n854 1.35607
R9600 vdd.n4570 vdd.n861 1.35607
R9601 vdd.n865 vdd.n864 1.35607
R9602 vdd.n4552 vdd.n920 1.35607
R9603 vdd.n4543 vdd.n950 1.35607
R9604 vdd.n4681 vdd.n4680 1.35607
R9605 vdd.n5577 vdd.n281 1.35607
R9606 vdd.n5467 vdd.n5466 1.35607
R9607 vdd.n5352 vdd.n407 1.35607
R9608 vdd.n5240 vdd.n5239 1.35607
R9609 vdd.n5124 vdd.n542 1.35607
R9610 vdd.n5012 vdd.n5011 1.35607
R9611 vdd.n4896 vdd.n677 1.35607
R9612 vdd.n4784 vdd.n4783 1.35607
R9613 vdd.n4702 vdd.n4701 1.35607
R9614 vdd.n7468 vdd.n221 1.35607
R9615 vdd.n7416 vdd 1.3165
R9616 vdd.n4025 vdd 1.14963
R9617 vdd.n3888 vdd.n3887 1.13981
R9618 vdd.n2222 vdd.n2221 1.13981
R9619 vdd.n5663 vdd.n5662 1.13717
R9620 vdd.n5630 vdd.n5628 1.13717
R9621 vdd.n5640 vdd.n5639 1.13717
R9622 vdd.n5709 vdd.n5708 1.13717
R9623 vdd.n271 vdd.n269 1.13717
R9624 vdd.n5594 vdd.n5593 1.13717
R9625 vdd.n276 vdd.n275 1.13717
R9626 vdd.n5601 vdd.n5600 1.13717
R9627 vdd.n5711 vdd.n5710 1.13717
R9628 vdd.n5638 vdd.n5637 1.13717
R9629 vdd.n5689 vdd.n5688 1.13717
R9630 vdd.n5655 vdd.n5650 1.13717
R9631 vdd.n2110 vdd.n2109 1.13717
R9632 vdd.n2098 vdd.n2097 1.13717
R9633 vdd.n2140 vdd.n2139 1.13717
R9634 vdd.n2186 vdd.n2166 1.13717
R9635 vdd.n2147 vdd.n2118 1.13717
R9636 vdd.n2145 vdd.n2116 1.13717
R9637 vdd.n2165 vdd.n2164 1.13717
R9638 vdd.n2162 vdd.n2161 1.13717
R9639 vdd.n2153 vdd.n2152 1.13717
R9640 vdd.n2151 vdd.n2150 1.13717
R9641 vdd.n4039 vdd.n2043 1.13717
R9642 vdd.n873 vdd.n872 1.13717
R9643 vdd.n4536 vdd.n4535 1.13717
R9644 vdd.n970 vdd.n958 1.13717
R9645 vdd.n918 vdd.n916 1.13717
R9646 vdd.n4563 vdd.n4562 1.13717
R9647 vdd.n901 vdd.n869 1.13717
R9648 vdd.n892 vdd.n891 1.13717
R9649 vdd.n909 vdd.n908 1.13717
R9650 vdd.n4560 vdd.n867 1.13717
R9651 vdd.n962 vdd.n961 1.13717
R9652 vdd.n978 vdd.n977 1.13717
R9653 vdd.n4533 vdd.n956 1.13717
R9654 vdd.n2026 vdd.n2024 1.13717
R9655 vdd.n2029 vdd.n1998 1.13717
R9656 vdd.n1984 vdd.n1982 1.13717
R9657 vdd.n1987 vdd.n1956 1.13717
R9658 vdd.n1942 vdd.n1940 1.13717
R9659 vdd.n1945 vdd.n1906 1.13717
R9660 vdd.n4121 vdd.n4120 1.13717
R9661 vdd.n1889 vdd.n1877 1.13717
R9662 vdd.n1837 vdd.n1835 1.13717
R9663 vdd.n4148 vdd.n4147 1.13717
R9664 vdd.n1820 vdd.n1813 1.13717
R9665 vdd.n4167 vdd.n4166 1.13717
R9666 vdd.n1762 vdd.n1760 1.13717
R9667 vdd.n1765 vdd.n1734 1.13717
R9668 vdd.n1720 vdd.n1718 1.13717
R9669 vdd.n1723 vdd.n1692 1.13717
R9670 vdd.n1678 vdd.n1676 1.13717
R9671 vdd.n1681 vdd.n1642 1.13717
R9672 vdd.n4242 vdd.n4241 1.13717
R9673 vdd.n1625 vdd.n1613 1.13717
R9674 vdd.n1573 vdd.n1571 1.13717
R9675 vdd.n4269 vdd.n4268 1.13717
R9676 vdd.n1556 vdd.n1549 1.13717
R9677 vdd.n4288 vdd.n4287 1.13717
R9678 vdd.n1498 vdd.n1496 1.13717
R9679 vdd.n1501 vdd.n1470 1.13717
R9680 vdd.n1456 vdd.n1454 1.13717
R9681 vdd.n1459 vdd.n1428 1.13717
R9682 vdd.n1414 vdd.n1412 1.13717
R9683 vdd.n1417 vdd.n1378 1.13717
R9684 vdd.n4363 vdd.n4362 1.13717
R9685 vdd.n1361 vdd.n1349 1.13717
R9686 vdd.n1309 vdd.n1307 1.13717
R9687 vdd.n4390 vdd.n4389 1.13717
R9688 vdd.n1292 vdd.n1285 1.13717
R9689 vdd.n4409 vdd.n4408 1.13717
R9690 vdd.n1234 vdd.n1232 1.13717
R9691 vdd.n1237 vdd.n1206 1.13717
R9692 vdd.n1192 vdd.n1190 1.13717
R9693 vdd.n1195 vdd.n1164 1.13717
R9694 vdd.n1150 vdd.n1148 1.13717
R9695 vdd.n1153 vdd.n1114 1.13717
R9696 vdd.n4484 vdd.n4483 1.13717
R9697 vdd.n1097 vdd.n1085 1.13717
R9698 vdd.n1045 vdd.n1043 1.13717
R9699 vdd.n4511 vdd.n4510 1.13717
R9700 vdd.n1028 vdd.n1017 1.13717
R9701 vdd.n985 vdd.n984 1.13717
R9702 vdd.n1020 vdd.n1019 1.13717
R9703 vdd.n1036 vdd.n1035 1.13717
R9704 vdd.n4508 vdd.n1015 1.13717
R9705 vdd.n1089 vdd.n1088 1.13717
R9706 vdd.n1105 vdd.n1104 1.13717
R9707 vdd.n4481 vdd.n1083 1.13717
R9708 vdd.n1151 vdd.n1112 1.13717
R9709 vdd.n4461 vdd.n4460 1.13717
R9710 vdd.n1193 vdd.n1162 1.13717
R9711 vdd.n4439 vdd.n4438 1.13717
R9712 vdd.n1235 vdd.n1204 1.13717
R9713 vdd.n4417 vdd.n4416 1.13717
R9714 vdd.n1247 vdd.n1246 1.13717
R9715 vdd.n1300 vdd.n1299 1.13717
R9716 vdd.n4387 vdd.n1283 1.13717
R9717 vdd.n1353 vdd.n1352 1.13717
R9718 vdd.n1369 vdd.n1368 1.13717
R9719 vdd.n4360 vdd.n1347 1.13717
R9720 vdd.n1415 vdd.n1376 1.13717
R9721 vdd.n4340 vdd.n4339 1.13717
R9722 vdd.n1457 vdd.n1426 1.13717
R9723 vdd.n4318 vdd.n4317 1.13717
R9724 vdd.n1499 vdd.n1468 1.13717
R9725 vdd.n4296 vdd.n4295 1.13717
R9726 vdd.n1511 vdd.n1510 1.13717
R9727 vdd.n1564 vdd.n1563 1.13717
R9728 vdd.n4266 vdd.n1547 1.13717
R9729 vdd.n1617 vdd.n1616 1.13717
R9730 vdd.n1633 vdd.n1632 1.13717
R9731 vdd.n4239 vdd.n1611 1.13717
R9732 vdd.n1679 vdd.n1640 1.13717
R9733 vdd.n4219 vdd.n4218 1.13717
R9734 vdd.n1721 vdd.n1690 1.13717
R9735 vdd.n4197 vdd.n4196 1.13717
R9736 vdd.n1763 vdd.n1732 1.13717
R9737 vdd.n4175 vdd.n4174 1.13717
R9738 vdd.n1775 vdd.n1774 1.13717
R9739 vdd.n1828 vdd.n1827 1.13717
R9740 vdd.n4145 vdd.n1811 1.13717
R9741 vdd.n1881 vdd.n1880 1.13717
R9742 vdd.n1897 vdd.n1896 1.13717
R9743 vdd.n4118 vdd.n1875 1.13717
R9744 vdd.n1943 vdd.n1904 1.13717
R9745 vdd.n4098 vdd.n4097 1.13717
R9746 vdd.n1985 vdd.n1954 1.13717
R9747 vdd.n4076 vdd.n4075 1.13717
R9748 vdd.n2027 vdd.n1996 1.13717
R9749 vdd.n4054 vdd.n4053 1.13717
R9750 vdd.n3992 vdd.n3991 1.13717
R9751 vdd.n2891 vdd.n2785 1.13717
R9752 vdd.n2864 vdd.n2792 1.13717
R9753 vdd.n2841 vdd.n2803 1.13717
R9754 vdd.n2834 vdd.n2833 1.13717
R9755 vdd.n2050 vdd.n2048 1.13717
R9756 vdd.n4037 vdd.n2042 1.13717
R9757 vdd.n2819 vdd.n2818 1.13717
R9758 vdd.n2835 vdd.n2814 1.13717
R9759 vdd.n2802 vdd.n2801 1.13717
R9760 vdd.n2791 vdd.n2790 1.13717
R9761 vdd.n2784 vdd.n2783 1.13717
R9762 vdd.n2781 vdd.n2780 1.13717
R9763 vdd.n2253 vdd.n2252 1.13717
R9764 vdd.n2268 vdd.n2265 1.13717
R9765 vdd.n3774 vdd.n3773 1.13717
R9766 vdd.n3751 vdd.n3750 1.13717
R9767 vdd.n2302 vdd.n2287 1.13717
R9768 vdd.n2311 vdd.n2305 1.13717
R9769 vdd.n3679 vdd.n2315 1.13717
R9770 vdd.n3656 vdd.n2337 1.13717
R9771 vdd.n3649 vdd.n3648 1.13717
R9772 vdd.n3627 vdd.n3626 1.13717
R9773 vdd.n3597 vdd.n2366 1.13717
R9774 vdd.n3569 vdd.n2377 1.13717
R9775 vdd.n2387 vdd.n2384 1.13717
R9776 vdd.n3559 vdd.n3558 1.13717
R9777 vdd.n2408 vdd.n2402 1.13717
R9778 vdd.n2422 vdd.n2420 1.13717
R9779 vdd.n3503 vdd.n3502 1.13717
R9780 vdd.n3480 vdd.n3479 1.13717
R9781 vdd.n3452 vdd.n2441 1.13717
R9782 vdd.n3428 vdd.n2472 1.13717
R9783 vdd.n3421 vdd.n3420 1.13717
R9784 vdd.n3399 vdd.n3398 1.13717
R9785 vdd.n3369 vdd.n2501 1.13717
R9786 vdd.n3341 vdd.n2512 1.13717
R9787 vdd.n2522 vdd.n2519 1.13717
R9788 vdd.n3331 vdd.n3330 1.13717
R9789 vdd.n2543 vdd.n2537 1.13717
R9790 vdd.n2557 vdd.n2555 1.13717
R9791 vdd.n3275 vdd.n3274 1.13717
R9792 vdd.n3252 vdd.n3251 1.13717
R9793 vdd.n3224 vdd.n2576 1.13717
R9794 vdd.n3200 vdd.n2607 1.13717
R9795 vdd.n3193 vdd.n3192 1.13717
R9796 vdd.n3171 vdd.n3170 1.13717
R9797 vdd.n3141 vdd.n2636 1.13717
R9798 vdd.n3113 vdd.n2647 1.13717
R9799 vdd.n2657 vdd.n2654 1.13717
R9800 vdd.n3103 vdd.n3102 1.13717
R9801 vdd.n2678 vdd.n2672 1.13717
R9802 vdd.n2692 vdd.n2690 1.13717
R9803 vdd.n3047 vdd.n3046 1.13717
R9804 vdd.n3024 vdd.n3023 1.13717
R9805 vdd.n2996 vdd.n2711 1.13717
R9806 vdd.n2972 vdd.n2742 1.13717
R9807 vdd.n2965 vdd.n2964 1.13717
R9808 vdd.n2943 vdd.n2942 1.13717
R9809 vdd.n2913 vdd.n2771 1.13717
R9810 vdd.n2902 vdd.n2782 1.13717
R9811 vdd.n2770 vdd.n2769 1.13717
R9812 vdd.n2935 vdd.n2768 1.13717
R9813 vdd.n2966 vdd.n2754 1.13717
R9814 vdd.n2741 vdd.n2740 1.13717
R9815 vdd.n2994 vdd.n2710 1.13717
R9816 vdd.n3016 vdd.n2707 1.13717
R9817 vdd.n2696 vdd.n2695 1.13717
R9818 vdd.n3054 vdd.n3053 1.13717
R9819 vdd.n3075 vdd.n3074 1.13717
R9820 vdd.n2662 vdd.n2661 1.13717
R9821 vdd.n3110 vdd.n3109 1.13717
R9822 vdd.n2646 vdd.n2645 1.13717
R9823 vdd.n2635 vdd.n2634 1.13717
R9824 vdd.n3163 vdd.n2633 1.13717
R9825 vdd.n3194 vdd.n2619 1.13717
R9826 vdd.n2606 vdd.n2605 1.13717
R9827 vdd.n3222 vdd.n2575 1.13717
R9828 vdd.n3244 vdd.n2572 1.13717
R9829 vdd.n2561 vdd.n2560 1.13717
R9830 vdd.n3282 vdd.n3281 1.13717
R9831 vdd.n3303 vdd.n3302 1.13717
R9832 vdd.n2527 vdd.n2526 1.13717
R9833 vdd.n3338 vdd.n3337 1.13717
R9834 vdd.n2511 vdd.n2510 1.13717
R9835 vdd.n2500 vdd.n2499 1.13717
R9836 vdd.n3391 vdd.n2498 1.13717
R9837 vdd.n3422 vdd.n2484 1.13717
R9838 vdd.n2471 vdd.n2470 1.13717
R9839 vdd.n3450 vdd.n2440 1.13717
R9840 vdd.n3472 vdd.n2437 1.13717
R9841 vdd.n2426 vdd.n2425 1.13717
R9842 vdd.n3510 vdd.n3509 1.13717
R9843 vdd.n3531 vdd.n3530 1.13717
R9844 vdd.n2392 vdd.n2391 1.13717
R9845 vdd.n3566 vdd.n3565 1.13717
R9846 vdd.n2376 vdd.n2375 1.13717
R9847 vdd.n2365 vdd.n2364 1.13717
R9848 vdd.n3619 vdd.n2363 1.13717
R9849 vdd.n3650 vdd.n2349 1.13717
R9850 vdd.n2336 vdd.n2335 1.13717
R9851 vdd.n2314 vdd.n2313 1.13717
R9852 vdd.n3699 vdd.n3698 1.13717
R9853 vdd.n3720 vdd.n3719 1.13717
R9854 vdd.n3743 vdd.n2284 1.13717
R9855 vdd.n2273 vdd.n2272 1.13717
R9856 vdd.n3781 vdd.n3780 1.13717
R9857 vdd.n3785 vdd.n3784 1.13717
R9858 vdd.n4599 vdd.n4598 1.13717
R9859 vdd.n805 vdd.n804 1.13717
R9860 vdd.n794 vdd.n793 1.13717
R9861 vdd.n4709 vdd.n792 1.13717
R9862 vdd.n4740 vdd.n778 1.13717
R9863 vdd.n765 vdd.n764 1.13717
R9864 vdd.n4768 vdd.n734 1.13717
R9865 vdd.n4790 vdd.n731 1.13717
R9866 vdd.n720 vdd.n719 1.13717
R9867 vdd.n4828 vdd.n4827 1.13717
R9868 vdd.n4849 vdd.n4848 1.13717
R9869 vdd.n686 vdd.n685 1.13717
R9870 vdd.n4884 vdd.n4883 1.13717
R9871 vdd.n670 vdd.n669 1.13717
R9872 vdd.n659 vdd.n658 1.13717
R9873 vdd.n4937 vdd.n657 1.13717
R9874 vdd.n4968 vdd.n643 1.13717
R9875 vdd.n630 vdd.n629 1.13717
R9876 vdd.n4996 vdd.n599 1.13717
R9877 vdd.n5018 vdd.n596 1.13717
R9878 vdd.n585 vdd.n584 1.13717
R9879 vdd.n5056 vdd.n5055 1.13717
R9880 vdd.n5077 vdd.n5076 1.13717
R9881 vdd.n551 vdd.n550 1.13717
R9882 vdd.n5112 vdd.n5111 1.13717
R9883 vdd.n535 vdd.n534 1.13717
R9884 vdd.n524 vdd.n523 1.13717
R9885 vdd.n5165 vdd.n522 1.13717
R9886 vdd.n5196 vdd.n508 1.13717
R9887 vdd.n495 vdd.n494 1.13717
R9888 vdd.n5224 vdd.n464 1.13717
R9889 vdd.n5246 vdd.n461 1.13717
R9890 vdd.n450 vdd.n449 1.13717
R9891 vdd.n5284 vdd.n5283 1.13717
R9892 vdd.n5305 vdd.n5304 1.13717
R9893 vdd.n416 vdd.n415 1.13717
R9894 vdd.n5340 vdd.n5339 1.13717
R9895 vdd.n400 vdd.n399 1.13717
R9896 vdd.n389 vdd.n388 1.13717
R9897 vdd.n5393 vdd.n387 1.13717
R9898 vdd.n5424 vdd.n373 1.13717
R9899 vdd.n360 vdd.n359 1.13717
R9900 vdd.n338 vdd.n337 1.13717
R9901 vdd.n5473 vdd.n5472 1.13717
R9902 vdd.n5495 vdd.n5494 1.13717
R9903 vdd.n5519 vdd.n310 1.13717
R9904 vdd.n299 vdd.n298 1.13717
R9905 vdd.n5557 vdd.n5556 1.13717
R9906 vdd.n5561 vdd.n5560 1.13717
R9907 vdd.n5497 vdd.n313 1.13717
R9908 vdd.n5527 vdd.n5526 1.13717
R9909 vdd.n5550 vdd.n5549 1.13717
R9910 vdd.n294 vdd.n291 1.13717
R9911 vdd.n279 vdd.n278 1.13717
R9912 vdd.n5475 vdd.n330 1.13717
R9913 vdd.n5371 vdd.n390 1.13717
R9914 vdd.n5401 vdd.n5400 1.13717
R9915 vdd.n5423 vdd.n5422 1.13717
R9916 vdd.n5430 vdd.n361 1.13717
R9917 vdd.n5453 vdd.n339 1.13717
R9918 vdd.n5343 vdd.n401 1.13717
R9919 vdd.n5277 vdd.n5276 1.13717
R9920 vdd.n446 vdd.n444 1.13717
R9921 vdd.n432 vdd.n426 1.13717
R9922 vdd.n5333 vdd.n5332 1.13717
R9923 vdd.n411 vdd.n408 1.13717
R9924 vdd.n5254 vdd.n5253 1.13717
R9925 vdd.n5143 vdd.n525 1.13717
R9926 vdd.n5173 vdd.n5172 1.13717
R9927 vdd.n5195 vdd.n5194 1.13717
R9928 vdd.n5202 vdd.n496 1.13717
R9929 vdd.n5226 vdd.n465 1.13717
R9930 vdd.n5115 vdd.n536 1.13717
R9931 vdd.n5049 vdd.n5048 1.13717
R9932 vdd.n581 vdd.n579 1.13717
R9933 vdd.n567 vdd.n561 1.13717
R9934 vdd.n5105 vdd.n5104 1.13717
R9935 vdd.n546 vdd.n543 1.13717
R9936 vdd.n5026 vdd.n5025 1.13717
R9937 vdd.n4915 vdd.n660 1.13717
R9938 vdd.n4945 vdd.n4944 1.13717
R9939 vdd.n4967 vdd.n4966 1.13717
R9940 vdd.n4974 vdd.n631 1.13717
R9941 vdd.n4998 vdd.n600 1.13717
R9942 vdd.n4887 vdd.n671 1.13717
R9943 vdd.n4821 vdd.n4820 1.13717
R9944 vdd.n716 vdd.n714 1.13717
R9945 vdd.n702 vdd.n696 1.13717
R9946 vdd.n4877 vdd.n4876 1.13717
R9947 vdd.n681 vdd.n678 1.13717
R9948 vdd.n4798 vdd.n4797 1.13717
R9949 vdd.n4717 vdd.n4716 1.13717
R9950 vdd.n4739 vdd.n4738 1.13717
R9951 vdd.n4746 vdd.n766 1.13717
R9952 vdd.n4770 vdd.n735 1.13717
R9953 vdd.n4687 vdd.n795 1.13717
R9954 vdd.n4676 vdd.n806 1.13717
R9955 vdd.n5761 vdd.n220 1.13717
R9956 vdd.n6398 vdd.n6386 1.13717
R9957 vdd.n7277 vdd.n7276 1.13717
R9958 vdd.n5865 vdd.n5864 1.13717
R9959 vdd.n7273 vdd.n7272 1.13717
R9960 vdd.n5878 vdd.n5873 1.13717
R9961 vdd.n7252 vdd.n7251 1.13717
R9962 vdd.n5891 vdd.n5889 1.13717
R9963 vdd.n5895 vdd.n5894 1.13717
R9964 vdd.n7245 vdd.n7244 1.13717
R9965 vdd.n7214 vdd.n5906 1.13717
R9966 vdd.n7222 vdd.n7221 1.13717
R9967 vdd.n7189 vdd.n7188 1.13717
R9968 vdd.n7191 vdd.n5909 1.13717
R9969 vdd.n7101 vdd.n5979 1.13717
R9970 vdd.n7099 vdd.n5978 1.13717
R9971 vdd.n7121 vdd.n5969 1.13717
R9972 vdd.n7120 vdd.n7119 1.13717
R9973 vdd.n5956 vdd.n5955 1.13717
R9974 vdd.n7127 vdd.n5957 1.13717
R9975 vdd.n5945 vdd.n5944 1.13717
R9976 vdd.n7149 vdd.n5946 1.13717
R9977 vdd.n5923 vdd.n5922 1.13717
R9978 vdd.n7169 vdd.n5924 1.13717
R9979 vdd.n7081 vdd.n5990 1.13717
R9980 vdd.n7079 vdd.n5989 1.13717
R9981 vdd.n7070 vdd.n7069 1.13717
R9982 vdd.n5998 vdd.n5994 1.13717
R9983 vdd.n7046 vdd.n7045 1.13717
R9984 vdd.n6011 vdd.n6007 1.13717
R9985 vdd.n7025 vdd.n7024 1.13717
R9986 vdd.n6024 vdd.n6022 1.13717
R9987 vdd.n6028 vdd.n6027 1.13717
R9988 vdd.n7018 vdd.n7017 1.13717
R9989 vdd.n6987 vdd.n6039 1.13717
R9990 vdd.n6995 vdd.n6994 1.13717
R9991 vdd.n6962 vdd.n6961 1.13717
R9992 vdd.n6964 vdd.n6042 1.13717
R9993 vdd.n6874 vdd.n6112 1.13717
R9994 vdd.n6872 vdd.n6111 1.13717
R9995 vdd.n6894 vdd.n6102 1.13717
R9996 vdd.n6893 vdd.n6892 1.13717
R9997 vdd.n6089 vdd.n6088 1.13717
R9998 vdd.n6900 vdd.n6090 1.13717
R9999 vdd.n6078 vdd.n6077 1.13717
R10000 vdd.n6922 vdd.n6079 1.13717
R10001 vdd.n6056 vdd.n6055 1.13717
R10002 vdd.n6942 vdd.n6057 1.13717
R10003 vdd.n6854 vdd.n6123 1.13717
R10004 vdd.n6852 vdd.n6122 1.13717
R10005 vdd.n6843 vdd.n6842 1.13717
R10006 vdd.n6131 vdd.n6127 1.13717
R10007 vdd.n6819 vdd.n6818 1.13717
R10008 vdd.n6144 vdd.n6140 1.13717
R10009 vdd.n6798 vdd.n6797 1.13717
R10010 vdd.n6157 vdd.n6155 1.13717
R10011 vdd.n6161 vdd.n6160 1.13717
R10012 vdd.n6791 vdd.n6790 1.13717
R10013 vdd.n6760 vdd.n6172 1.13717
R10014 vdd.n6768 vdd.n6767 1.13717
R10015 vdd.n6735 vdd.n6734 1.13717
R10016 vdd.n6737 vdd.n6175 1.13717
R10017 vdd.n6647 vdd.n6245 1.13717
R10018 vdd.n6645 vdd.n6244 1.13717
R10019 vdd.n6667 vdd.n6235 1.13717
R10020 vdd.n6666 vdd.n6665 1.13717
R10021 vdd.n6222 vdd.n6221 1.13717
R10022 vdd.n6673 vdd.n6223 1.13717
R10023 vdd.n6211 vdd.n6210 1.13717
R10024 vdd.n6695 vdd.n6212 1.13717
R10025 vdd.n6189 vdd.n6188 1.13717
R10026 vdd.n6715 vdd.n6190 1.13717
R10027 vdd.n6627 vdd.n6256 1.13717
R10028 vdd.n6625 vdd.n6255 1.13717
R10029 vdd.n6616 vdd.n6615 1.13717
R10030 vdd.n6264 vdd.n6260 1.13717
R10031 vdd.n6592 vdd.n6591 1.13717
R10032 vdd.n6277 vdd.n6273 1.13717
R10033 vdd.n6571 vdd.n6570 1.13717
R10034 vdd.n6290 vdd.n6288 1.13717
R10035 vdd.n6294 vdd.n6293 1.13717
R10036 vdd.n6564 vdd.n6563 1.13717
R10037 vdd.n6533 vdd.n6305 1.13717
R10038 vdd.n6541 vdd.n6540 1.13717
R10039 vdd.n6508 vdd.n6507 1.13717
R10040 vdd.n6510 vdd.n6308 1.13717
R10041 vdd.n6440 vdd.n6368 1.13717
R10042 vdd.n6439 vdd.n6438 1.13717
R10043 vdd.n6355 vdd.n6354 1.13717
R10044 vdd.n6446 vdd.n6356 1.13717
R10045 vdd.n6344 vdd.n6343 1.13717
R10046 vdd.n6468 vdd.n6345 1.13717
R10047 vdd.n6322 vdd.n6321 1.13717
R10048 vdd.n6488 vdd.n6323 1.13717
R10049 vdd.n6418 vdd.n6377 1.13717
R10050 vdd.n6420 vdd.n6378 1.13717
R10051 vdd.n6400 vdd.n6387 1.13717
R10052 vdd.n5822 vdd.n5817 1.13717
R10053 vdd.n5833 vdd.n5829 1.13717
R10054 vdd.n5844 vdd.n5840 1.13717
R10055 vdd.n5855 vdd.n5851 1.13717
R10056 vdd.n7303 vdd.n5862 1.13717
R10057 vdd.n7307 vdd.n7306 1.13717
R10058 vdd.n7326 vdd.n7325 1.13717
R10059 vdd.n7345 vdd.n7344 1.13717
R10060 vdd.n7364 vdd.n7363 1.13717
R10061 vdd.n7383 vdd.n7382 1.13717
R10062 vdd.n7387 vdd.n7386 1.13717
R10063 vdd.n7404 vdd.n5795 1.13717
R10064 vdd.n7526 vdd.n7525 1.13717
R10065 vdd.n184 vdd.n183 1.13717
R10066 vdd.n143 vdd.n142 1.13717
R10067 vdd.n7495 vdd.n200 1.13667
R10068 vdd.n3812 vdd.n2249 1.13645
R10069 vdd.n204 vdd.n202 1.13501
R10070 vdd.n3816 vdd.n3815 1.13462
R10071 vdd.n2086 vdd.n2085 1.13462
R10072 vdd.n3912 vdd.n3911 1.13462
R10073 vdd.n3939 vdd.n3938 1.13462
R10074 vdd.n3875 vdd.n3874 1.13462
R10075 vdd.n3881 vdd.n3880 1.13462
R10076 vdd.n3914 vdd.n3913 1.13462
R10077 vdd.n3972 vdd.n3971 1.13462
R10078 vdd.n3953 vdd.n3952 1.13462
R10079 vdd.n3959 vdd.n3958 1.13462
R10080 vdd.n3830 vdd.n3829 1.13462
R10081 vdd.n2228 vdd.n2227 1.13462
R10082 vdd.n2075 vdd.n2074 1.13462
R10083 vdd.n2240 vdd.n2239 1.13462
R10084 vdd.n2128 vdd.n2127 1.13005
R10085 vdd.n3899 vdd.n3898 1.13005
R10086 vdd.n836 vdd.n835 1.13005
R10087 vdd.n5771 vdd.n5770 1.13005
R10088 vdd.n2211 vdd.n2103 1.12991
R10089 vdd.n3809 vdd.n3808 1.04044
R10090 vdd.n2243 vdd.n2242 1.04044
R10091 vdd.n3823 vdd.n2078 1.04044
R10092 vdd.n2232 vdd.n2231 1.04044
R10093 vdd.n3833 vdd.n2070 1.04044
R10094 vdd.n2088 vdd.n2080 1.04044
R10095 vdd.n3819 vdd.n2081 1.04044
R10096 vdd.n3960 vdd.n3947 1.04044
R10097 vdd.n3954 vdd.n3948 1.04044
R10098 vdd.n3975 vdd.n3949 1.04044
R10099 vdd.n3924 vdd.n3916 1.04044
R10100 vdd.n3884 vdd.n3883 1.04044
R10101 vdd.n3876 vdd.n3870 1.04044
R10102 vdd.n3942 vdd.n3871 1.04044
R10103 vdd.n3932 vdd.n3931 1.04044
R10104 vdd.n7460 vdd.n7459 1.04017
R10105 vdd.n7453 vdd.n229 1.04017
R10106 vdd.n5743 vdd.n5742 1.04017
R10107 vdd.n7438 vdd.n7437 1.04017
R10108 vdd.n7444 vdd.n7443 1.04017
R10109 vdd.n5784 vdd.n5783 1.04017
R10110 vdd.n7427 vdd.n7426 1.04017
R10111 vdd.n5810 vdd.n5809 1.04017
R10112 vdd.n4665 vdd.n4664 1.04017
R10113 vdd.n4651 vdd.n4650 1.04017
R10114 vdd.n4657 vdd.n4656 1.04017
R10115 vdd.n4641 vdd.n4640 1.04017
R10116 vdd.n826 vdd.n825 1.04017
R10117 vdd.n2177 vdd.n2176 1.01997
R10118 vdd.n7503 vdd.n196 1.01637
R10119 vdd.n3866 vdd.n3865 1.01637
R10120 vdd.n4618 vdd.n846 1.01637
R10121 vdd.n7466 vdd.n223 1.01637
R10122 vdd vdd.n3836 0.985466
R10123 vdd.n4633 vdd.n4632 0.936863
R10124 vdd vdd.t75 0.918966
R10125 vdd.t86 vdd 0.918966
R10126 vdd.n2177 vdd.n2167 0.906695
R10127 vdd.n242 vdd.n238 0.870766
R10128 vdd.n3850 vdd.n3848 0.870578
R10129 vdd.n3997 vdd.n3996 0.870578
R10130 vdd.n4593 vdd.n841 0.870578
R10131 vdd.n4604 vdd.n4603 0.870578
R10132 vdd.n7475 vdd.n7474 0.870578
R10133 vdd.n829 vdd.n828 0.853291
R10134 vdd.n5764 vdd.n5763 0.853291
R10135 vdd.n7500 vdd.n200 0.853
R10136 vdd.n244 vdd.n243 0.853
R10137 vdd.n2083 vdd.n2082 0.853
R10138 vdd.n2092 vdd.n2089 0.853
R10139 vdd.n880 vdd.n879 0.853
R10140 vdd.n3935 vdd.n3930 0.853
R10141 vdd.n3873 vdd.n3872 0.853
R10142 vdd.n3908 vdd.n3877 0.853
R10143 vdd.n3905 vdd.n3882 0.853
R10144 vdd.n3927 vdd.n3915 0.853
R10145 vdd.n3991 vdd.n3846 0.853
R10146 vdd.n3951 vdd.n3950 0.853
R10147 vdd.n3967 vdd.n3955 0.853
R10148 vdd.n3964 vdd.n3961 0.853
R10149 vdd.n4044 vdd.n2037 0.853
R10150 vdd.n2072 vdd.n2071 0.853
R10151 vdd.n2235 vdd.n2230 0.853
R10152 vdd.n3826 vdd.n2077 0.853
R10153 vdd.n2247 vdd.n2241 0.853
R10154 vdd.n3806 vdd.n2249 0.853
R10155 vdd.n4598 vdd.n4589 0.853
R10156 vdd.n824 vdd.n823 0.853
R10157 vdd.n823 vdd.n814 0.853
R10158 vdd.n4639 vdd.n815 0.853
R10159 vdd.n4660 vdd.n815 0.853
R10160 vdd.n4659 vdd.n817 0.853
R10161 vdd.n4660 vdd.n4659 0.853
R10162 vdd.n4649 vdd.n4648 0.853
R10163 vdd.n4648 vdd.n814 0.853
R10164 vdd.n808 vdd.n807 0.853
R10165 vdd.n811 vdd.n810 0.853
R10166 vdd.n818 vdd.n810 0.853
R10167 vdd.n221 vdd.n220 0.853
R10168 vdd.n5740 vdd.n5739 0.853
R10169 vdd.n5739 vdd.n233 0.853
R10170 vdd.n7455 vdd.n237 0.853
R10171 vdd.n7456 vdd.n7455 0.853
R10172 vdd.n7458 vdd.n7457 0.853
R10173 vdd.n7457 vdd.n7456 0.853
R10174 vdd.n5808 vdd.n5807 0.853
R10175 vdd.n5807 vdd.n5778 0.853
R10176 vdd.n7429 vdd.n7428 0.853
R10177 vdd.n7430 vdd.n7429 0.853
R10178 vdd.n5786 vdd.n5785 0.853
R10179 vdd.n5787 vdd.n5786 0.853
R10180 vdd.n5776 vdd.n5775 0.853
R10181 vdd.n5787 vdd.n5775 0.853
R10182 vdd.n7432 vdd.n7431 0.853
R10183 vdd.n7431 vdd.n7430 0.853
R10184 vdd.n6389 vdd.n6388 0.853
R10185 vdd.n7412 vdd.n5793 0.853
R10186 vdd.n189 vdd.n188 0.853
R10187 vdd.n2129 vdd.n2128 0.851407
R10188 vdd.n3900 vdd.n3899 0.851407
R10189 vdd.n7304 vdd.n7302 0.849366
R10190 vdd.n2897 vdd.n2896 0.84923
R10191 vdd.n954 vdd.n953 0.84923
R10192 vdd.n5585 vdd.n261 0.849012
R10193 vdd.n7486 vdd.n211 0.813198
R10194 vdd.n7505 vdd.n7503 0.813198
R10195 vdd.n3865 vdd.n3856 0.813198
R10196 vdd.n4002 vdd.n4001 0.813198
R10197 vdd.n4618 vdd.n4586 0.813198
R10198 vdd.n4610 vdd.n4609 0.813198
R10199 vdd.n5753 vdd.n5752 0.813198
R10200 vdd.n7466 vdd.n225 0.813198
R10201 vdd.n4576 vdd.n851 0.734658
R10202 vdd.n4574 vdd.n856 0.734658
R10203 vdd.n932 vdd.n926 0.734658
R10204 vdd.n4549 vdd.n944 0.734658
R10205 vdd.n4547 vdd.n945 0.734658
R10206 vdd.n1001 vdd.n992 0.734658
R10207 vdd.n4524 vdd.n1003 0.734658
R10208 vdd.n4522 vdd.n1004 0.734658
R10209 vdd.n1059 vdd.n1053 0.734658
R10210 vdd.n4497 vdd.n1071 0.734658
R10211 vdd.n4495 vdd.n1072 0.734658
R10212 vdd.n1140 vdd.n1120 0.734658
R10213 vdd.n4472 vdd.n4471 0.734658
R10214 vdd.n1182 vdd.n1142 0.734658
R10215 vdd.n4450 vdd.n4449 0.734658
R10216 vdd.n1224 vdd.n1184 0.734658
R10217 vdd.n4428 vdd.n4427 0.734658
R10218 vdd.n1264 vdd.n1226 0.734658
R10219 vdd.n4403 vdd.n1271 0.734658
R10220 vdd.n4401 vdd.n1272 0.734658
R10221 vdd.n1323 vdd.n1317 0.734658
R10222 vdd.n4376 vdd.n1335 0.734658
R10223 vdd.n4374 vdd.n1336 0.734658
R10224 vdd.n1404 vdd.n1384 0.734658
R10225 vdd.n4351 vdd.n4350 0.734658
R10226 vdd.n1446 vdd.n1406 0.734658
R10227 vdd.n4329 vdd.n4328 0.734658
R10228 vdd.n1488 vdd.n1448 0.734658
R10229 vdd.n4307 vdd.n4306 0.734658
R10230 vdd.n1528 vdd.n1490 0.734658
R10231 vdd.n4282 vdd.n1535 0.734658
R10232 vdd.n4280 vdd.n1536 0.734658
R10233 vdd.n1587 vdd.n1581 0.734658
R10234 vdd.n4255 vdd.n1599 0.734658
R10235 vdd.n4253 vdd.n1600 0.734658
R10236 vdd.n1668 vdd.n1648 0.734658
R10237 vdd.n4230 vdd.n4229 0.734658
R10238 vdd.n1710 vdd.n1670 0.734658
R10239 vdd.n4208 vdd.n4207 0.734658
R10240 vdd.n1752 vdd.n1712 0.734658
R10241 vdd.n4186 vdd.n4185 0.734658
R10242 vdd.n1792 vdd.n1754 0.734658
R10243 vdd.n4161 vdd.n1799 0.734658
R10244 vdd.n4159 vdd.n1800 0.734658
R10245 vdd.n1851 vdd.n1845 0.734658
R10246 vdd.n4134 vdd.n1863 0.734658
R10247 vdd.n4132 vdd.n1864 0.734658
R10248 vdd.n1932 vdd.n1912 0.734658
R10249 vdd.n4109 vdd.n4108 0.734658
R10250 vdd.n1974 vdd.n1934 0.734658
R10251 vdd.n4087 vdd.n4086 0.734658
R10252 vdd.n2016 vdd.n1976 0.734658
R10253 vdd.n4065 vdd.n4064 0.734658
R10254 vdd.n3917 vdd.n2018 0.734658
R10255 vdd.n3943 vdd.n3869 0.734658
R10256 vdd.n2223 vdd.n2222 0.684595
R10257 vdd.n3889 vdd.n3888 0.684595
R10258 vdd.n7516 vdd.n7515 0.682973
R10259 vdd.n7476 vdd.n217 0.682713
R10260 vdd.n7493 vdd.n7492 0.682713
R10261 vdd.n3998 vdd.n3840 0.682713
R10262 vdd.n3987 vdd.n3986 0.682713
R10263 vdd.n4605 vdd.n4591 0.682713
R10264 vdd.n4629 vdd.n4628 0.682713
R10265 vdd.n5750 vdd.n5749 0.682713
R10266 vdd.n7420 vdd.n7419 0.682707
R10267 vdd.n6392 vdd.n6391 0.682697
R10268 vdd.n4670 vdd.n4669 0.682697
R10269 vdd.n5734 vdd.n5733 0.682447
R10270 vdd.n4045 vdd.n2038 0.682447
R10271 vdd.n882 vdd.n881 0.682447
R10272 vdd.n28 vdd.n25 0.660294
R10273 vdd.n7424 vdd.t82 0.612811
R10274 vdd.t85 vdd.n247 0.612811
R10275 vdd.n115 vdd.n114 0.600276
R10276 vdd.n4673 vdd 0.547714
R10277 vdd.n1141 vdd 0.534441
R10278 vdd.n1405 vdd 0.534441
R10279 vdd.n1669 vdd 0.534441
R10280 vdd.n1933 vdd 0.534441
R10281 vdd.n4007 vdd.t29 0.492983
R10282 vdd.n4025 vdd.n2065 0.492983
R10283 vdd.t0 vdd.t119 0.491014
R10284 vdd.n5812 vdd.n212 0.459733
R10285 vdd.n5727 vdd.n250 0.459733
R10286 vdd.t32 vdd.n7435 0.454532
R10287 vdd.t39 vdd.n4652 0.454532
R10288 vdd.n7435 vdd.t102 0.45205
R10289 vdd.n4652 vdd.t99 0.45205
R10290 vdd.n7512 vdd.n7511 0.406849
R10291 vdd.n3855 vdd.n3854 0.406849
R10292 vdd.n845 vdd.n844 0.406849
R10293 vdd.n7480 vdd.n7479 0.406849
R10294 vdd.n3901 vdd.n3900 0.370457
R10295 vdd.n42 vdd.n39 0.370442
R10296 vdd.n4634 vdd.n837 0.35535
R10297 vdd.n7448 vdd.n5772 0.35535
R10298 vdd.n7296 vdd 0.321584
R10299 vdd.n7297 vdd 0.317995
R10300 vdd.n6266 vdd.n6254 0.314894
R10301 vdd.n6133 vdd.n6121 0.314894
R10302 vdd.n6000 vdd.n5988 0.314894
R10303 vdd.n4895 vdd.n672 0.314894
R10304 vdd.n5123 vdd.n537 0.314894
R10305 vdd.n5351 vdd.n402 0.314894
R10306 vdd.n3121 vdd.n2648 0.314894
R10307 vdd.n3349 vdd.n2513 0.314894
R10308 vdd.n3577 vdd.n2378 0.314894
R10309 vdd.n1255 vdd.n1254 0.314894
R10310 vdd.n1519 vdd.n1518 0.314894
R10311 vdd.n1783 vdd.n1782 0.314894
R10312 vdd.n6333 vdd.n6330 0.30353
R10313 vdd.n6200 vdd.n6197 0.30353
R10314 vdd.n6067 vdd.n6064 0.30353
R10315 vdd.n5934 vdd.n5931 0.30353
R10316 vdd.n6332 vdd.n6331 0.30353
R10317 vdd.n6199 vdd.n6198 0.30353
R10318 vdd.n6066 vdd.n6065 0.30353
R10319 vdd.n5933 vdd.n5932 0.30353
R10320 vdd.n754 vdd.n741 0.30353
R10321 vdd.n619 vdd.n606 0.30353
R10322 vdd.n484 vdd.n471 0.30353
R10323 vdd.n349 vdd.n346 0.30353
R10324 vdd.n2730 vdd.n2717 0.30353
R10325 vdd.n2595 vdd.n2582 0.30353
R10326 vdd.n2460 vdd.n2447 0.30353
R10327 vdd.n2325 vdd.n2322 0.30353
R10328 vdd.n2729 vdd.n2728 0.30353
R10329 vdd.n2594 vdd.n2593 0.30353
R10330 vdd.n2459 vdd.n2458 0.30353
R10331 vdd.n2324 vdd.n2323 0.30353
R10332 vdd.n1133 vdd.n1132 0.30353
R10333 vdd.n1397 vdd.n1396 0.30353
R10334 vdd.n1661 vdd.n1660 0.30353
R10335 vdd.n1925 vdd.n1924 0.30353
R10336 vdd.n1134 vdd.n1129 0.30353
R10337 vdd.n1398 vdd.n1393 0.30353
R10338 vdd.n1662 vdd.n1657 0.30353
R10339 vdd.n1926 vdd.n1921 0.30353
R10340 vdd.n753 vdd.n752 0.30353
R10341 vdd.n618 vdd.n617 0.30353
R10342 vdd.n483 vdd.n482 0.30353
R10343 vdd.n348 vdd.n347 0.30353
R10344 vdd.n6623 vdd.n6621 0.288379
R10345 vdd.n6850 vdd.n6848 0.288379
R10346 vdd.n7077 vdd.n7075 0.288379
R10347 vdd.n3119 vdd.n2656 0.288379
R10348 vdd.n3347 vdd.n2521 0.288379
R10349 vdd.n3575 vdd.n2386 0.288379
R10350 vdd.n1252 vdd.n1251 0.288379
R10351 vdd.n1516 vdd.n1515 0.288379
R10352 vdd.n1780 vdd.n1779 0.288379
R10353 vdd.n4893 vdd.n680 0.288379
R10354 vdd.n5121 vdd.n545 0.288379
R10355 vdd.n5349 vdd.n410 0.288379
R10356 vdd.n6395 vdd 0.266176
R10357 vdd.n3813 vdd.n2238 0.243205
R10358 vdd.n3814 vdd.n3813 0.214242
R10359 vdd.n7519 vdd.n7518 0.199638
R10360 vdd.n177 vdd.n176 0.197423
R10361 vdd.n17 vdd.n16 0.197423
R10362 vdd.n6406 vdd.n6384 0.194439
R10363 vdd.n6427 vdd.n6375 0.194439
R10364 vdd.n6427 vdd.n6373 0.194439
R10365 vdd.n6454 vdd.n6360 0.194439
R10366 vdd.n6454 vdd.n6361 0.194439
R10367 vdd.n6460 vdd.n6459 0.194439
R10368 vdd.n6460 vdd.n6349 0.194439
R10369 vdd.n6480 vdd.n6347 0.194439
R10370 vdd.n6480 vdd.n6338 0.194439
R10371 vdd.n6499 vdd.n6327 0.194439
R10372 vdd.n6499 vdd.n6336 0.194439
R10373 vdd.n6513 vdd.n6317 0.194439
R10374 vdd.n6513 vdd.n6316 0.194439
R10375 vdd.n6522 vdd.n6521 0.194439
R10376 vdd.n6521 vdd.n6315 0.194439
R10377 vdd.n6549 vdd.n6548 0.194439
R10378 vdd.n6549 vdd.n6298 0.194439
R10379 vdd.n6580 vdd.n6282 0.194439
R10380 vdd.n6581 vdd.n6580 0.194439
R10381 vdd.n6587 vdd.n6279 0.194439
R10382 vdd.n6587 vdd.n6270 0.194439
R10383 vdd.n6611 vdd.n6267 0.194439
R10384 vdd.n6611 vdd.n6268 0.194439
R10385 vdd.n6633 vdd.n6253 0.194439
R10386 vdd.n6633 vdd.n6251 0.194439
R10387 vdd.n6654 vdd.n6242 0.194439
R10388 vdd.n6654 vdd.n6240 0.194439
R10389 vdd.n6681 vdd.n6227 0.194439
R10390 vdd.n6681 vdd.n6228 0.194439
R10391 vdd.n6687 vdd.n6686 0.194439
R10392 vdd.n6687 vdd.n6216 0.194439
R10393 vdd.n6707 vdd.n6214 0.194439
R10394 vdd.n6707 vdd.n6205 0.194439
R10395 vdd.n6726 vdd.n6194 0.194439
R10396 vdd.n6726 vdd.n6203 0.194439
R10397 vdd.n6740 vdd.n6184 0.194439
R10398 vdd.n6740 vdd.n6183 0.194439
R10399 vdd.n6749 vdd.n6748 0.194439
R10400 vdd.n6748 vdd.n6182 0.194439
R10401 vdd.n6776 vdd.n6775 0.194439
R10402 vdd.n6776 vdd.n6165 0.194439
R10403 vdd.n6807 vdd.n6149 0.194439
R10404 vdd.n6808 vdd.n6807 0.194439
R10405 vdd.n6814 vdd.n6146 0.194439
R10406 vdd.n6814 vdd.n6137 0.194439
R10407 vdd.n6838 vdd.n6134 0.194439
R10408 vdd.n6838 vdd.n6135 0.194439
R10409 vdd.n6860 vdd.n6120 0.194439
R10410 vdd.n6860 vdd.n6118 0.194439
R10411 vdd.n6881 vdd.n6109 0.194439
R10412 vdd.n6881 vdd.n6107 0.194439
R10413 vdd.n6908 vdd.n6094 0.194439
R10414 vdd.n6908 vdd.n6095 0.194439
R10415 vdd.n6914 vdd.n6913 0.194439
R10416 vdd.n6914 vdd.n6083 0.194439
R10417 vdd.n6934 vdd.n6081 0.194439
R10418 vdd.n6934 vdd.n6072 0.194439
R10419 vdd.n6953 vdd.n6061 0.194439
R10420 vdd.n6953 vdd.n6070 0.194439
R10421 vdd.n6967 vdd.n6051 0.194439
R10422 vdd.n6967 vdd.n6050 0.194439
R10423 vdd.n6976 vdd.n6975 0.194439
R10424 vdd.n6975 vdd.n6049 0.194439
R10425 vdd.n7003 vdd.n7002 0.194439
R10426 vdd.n7003 vdd.n6032 0.194439
R10427 vdd.n7034 vdd.n6016 0.194439
R10428 vdd.n7035 vdd.n7034 0.194439
R10429 vdd.n7041 vdd.n6013 0.194439
R10430 vdd.n7041 vdd.n6004 0.194439
R10431 vdd.n7065 vdd.n6001 0.194439
R10432 vdd.n7065 vdd.n6002 0.194439
R10433 vdd.n7087 vdd.n5987 0.194439
R10434 vdd.n7087 vdd.n5985 0.194439
R10435 vdd.n7108 vdd.n5976 0.194439
R10436 vdd.n7108 vdd.n5974 0.194439
R10437 vdd.n7135 vdd.n5961 0.194439
R10438 vdd.n7135 vdd.n5962 0.194439
R10439 vdd.n7141 vdd.n7140 0.194439
R10440 vdd.n7141 vdd.n5950 0.194439
R10441 vdd.n7161 vdd.n5948 0.194439
R10442 vdd.n7161 vdd.n5939 0.194439
R10443 vdd.n7180 vdd.n5928 0.194439
R10444 vdd.n7180 vdd.n5937 0.194439
R10445 vdd.n7194 vdd.n5918 0.194439
R10446 vdd.n7194 vdd.n5917 0.194439
R10447 vdd.n7203 vdd.n7202 0.194439
R10448 vdd.n7202 vdd.n5916 0.194439
R10449 vdd.n7230 vdd.n7229 0.194439
R10450 vdd.n7230 vdd.n5899 0.194439
R10451 vdd.n7261 vdd.n5883 0.194439
R10452 vdd.n7262 vdd.n7261 0.194439
R10453 vdd.n7268 vdd.n5880 0.194439
R10454 vdd.n7268 vdd.n5870 0.194439
R10455 vdd.n7291 vdd.n5868 0.194439
R10456 vdd.n7301 vdd.n5859 0.194439
R10457 vdd.n7321 vdd.n5857 0.194439
R10458 vdd.n7321 vdd.n5848 0.194439
R10459 vdd.n7340 vdd.n5846 0.194439
R10460 vdd.n7340 vdd.n5837 0.194439
R10461 vdd.n7359 vdd.n5835 0.194439
R10462 vdd.n7359 vdd.n5826 0.194439
R10463 vdd.n7378 vdd.n5824 0.194439
R10464 vdd.n7378 vdd.n5814 0.194439
R10465 vdd.n7401 vdd.n5799 0.194439
R10466 vdd.n7401 vdd.n5800 0.194439
R10467 vdd.n5725 vdd.n5724 0.194439
R10468 vdd.n5720 vdd.n263 0.194439
R10469 vdd.n5720 vdd.n265 0.194439
R10470 vdd.n5619 vdd.n5617 0.194439
R10471 vdd.n5621 vdd.n5619 0.194439
R10472 vdd.n5701 vdd.n5700 0.194439
R10473 vdd.n5700 vdd.n5698 0.194439
R10474 vdd.n5666 vdd.n5624 0.194439
R10475 vdd.n5667 vdd.n5666 0.194439
R10476 vdd.n5680 vdd.n5678 0.194439
R10477 vdd.n5680 vdd.n248 0.194439
R10478 vdd.n2905 vdd.n2775 0.194439
R10479 vdd.n2926 vdd.n2773 0.194439
R10480 vdd.n2926 vdd.n2762 0.194439
R10481 vdd.n2951 vdd.n2760 0.194439
R10482 vdd.n2760 vdd.n2759 0.194439
R10483 vdd.n2980 vdd.n2746 0.194439
R10484 vdd.n2980 vdd.n2747 0.194439
R10485 vdd.n2987 vdd.n2986 0.194439
R10486 vdd.n2987 vdd.n2735 0.194439
R10487 vdd.n3008 vdd.n2715 0.194439
R10488 vdd.n3008 vdd.n2733 0.194439
R10489 vdd.n2725 vdd.n2724 0.194439
R10490 vdd.n2724 vdd.n2720 0.194439
R10491 vdd.n3032 vdd.n3031 0.194439
R10492 vdd.n3032 vdd.n2700 0.194439
R10493 vdd.n3063 vdd.n2684 0.194439
R10494 vdd.n3064 vdd.n3063 0.194439
R10495 vdd.n3070 vdd.n2681 0.194439
R10496 vdd.n3070 vdd.n2668 0.194439
R10497 vdd.n2669 vdd.n2666 0.194439
R10498 vdd.n3093 vdd.n2666 0.194439
R10499 vdd.n3123 vdd.n2651 0.194439
R10500 vdd.n3123 vdd.n2649 0.194439
R10501 vdd.n3133 vdd.n3132 0.194439
R10502 vdd.n3133 vdd.n2640 0.194439
R10503 vdd.n3154 vdd.n2638 0.194439
R10504 vdd.n3154 vdd.n2627 0.194439
R10505 vdd.n3179 vdd.n2625 0.194439
R10506 vdd.n2625 vdd.n2624 0.194439
R10507 vdd.n3208 vdd.n2611 0.194439
R10508 vdd.n3208 vdd.n2612 0.194439
R10509 vdd.n3215 vdd.n3214 0.194439
R10510 vdd.n3215 vdd.n2600 0.194439
R10511 vdd.n3236 vdd.n2580 0.194439
R10512 vdd.n3236 vdd.n2598 0.194439
R10513 vdd.n2590 vdd.n2589 0.194439
R10514 vdd.n2589 vdd.n2585 0.194439
R10515 vdd.n3260 vdd.n3259 0.194439
R10516 vdd.n3260 vdd.n2565 0.194439
R10517 vdd.n3291 vdd.n2549 0.194439
R10518 vdd.n3292 vdd.n3291 0.194439
R10519 vdd.n3298 vdd.n2546 0.194439
R10520 vdd.n3298 vdd.n2533 0.194439
R10521 vdd.n2534 vdd.n2531 0.194439
R10522 vdd.n3321 vdd.n2531 0.194439
R10523 vdd.n3351 vdd.n2516 0.194439
R10524 vdd.n3351 vdd.n2514 0.194439
R10525 vdd.n3361 vdd.n3360 0.194439
R10526 vdd.n3361 vdd.n2505 0.194439
R10527 vdd.n3382 vdd.n2503 0.194439
R10528 vdd.n3382 vdd.n2492 0.194439
R10529 vdd.n3407 vdd.n2490 0.194439
R10530 vdd.n2490 vdd.n2489 0.194439
R10531 vdd.n3436 vdd.n2476 0.194439
R10532 vdd.n3436 vdd.n2477 0.194439
R10533 vdd.n3443 vdd.n3442 0.194439
R10534 vdd.n3443 vdd.n2465 0.194439
R10535 vdd.n3464 vdd.n2445 0.194439
R10536 vdd.n3464 vdd.n2463 0.194439
R10537 vdd.n2455 vdd.n2454 0.194439
R10538 vdd.n2454 vdd.n2450 0.194439
R10539 vdd.n3488 vdd.n3487 0.194439
R10540 vdd.n3488 vdd.n2430 0.194439
R10541 vdd.n3519 vdd.n2414 0.194439
R10542 vdd.n3520 vdd.n3519 0.194439
R10543 vdd.n3526 vdd.n2411 0.194439
R10544 vdd.n3526 vdd.n2398 0.194439
R10545 vdd.n2399 vdd.n2396 0.194439
R10546 vdd.n3549 vdd.n2396 0.194439
R10547 vdd.n3579 vdd.n2381 0.194439
R10548 vdd.n3579 vdd.n2379 0.194439
R10549 vdd.n3589 vdd.n3588 0.194439
R10550 vdd.n3589 vdd.n2370 0.194439
R10551 vdd.n3610 vdd.n2368 0.194439
R10552 vdd.n3610 vdd.n2357 0.194439
R10553 vdd.n3635 vdd.n2355 0.194439
R10554 vdd.n2355 vdd.n2354 0.194439
R10555 vdd.n3664 vdd.n2341 0.194439
R10556 vdd.n3664 vdd.n2342 0.194439
R10557 vdd.n3671 vdd.n3670 0.194439
R10558 vdd.n3671 vdd.n2330 0.194439
R10559 vdd.n3691 vdd.n2319 0.194439
R10560 vdd.n3691 vdd.n2328 0.194439
R10561 vdd.n3703 vdd.n2308 0.194439
R10562 vdd.n3707 vdd.n3703 0.194439
R10563 vdd.n3724 vdd.n2299 0.194439
R10564 vdd.n3724 vdd.n2297 0.194439
R10565 vdd.n3732 vdd.n3731 0.194439
R10566 vdd.n3731 vdd.n2294 0.194439
R10567 vdd.n3759 vdd.n3758 0.194439
R10568 vdd.n3759 vdd.n2277 0.194439
R10569 vdd.n3794 vdd.n2259 0.194439
R10570 vdd.n3795 vdd.n3794 0.194439
R10571 vdd.n3800 vdd.n2256 0.194439
R10572 vdd.n4022 vdd.n4021 0.194439
R10573 vdd.n4021 vdd.n4009 0.194439
R10574 vdd.n4028 vdd.n2054 0.194439
R10575 vdd.n4028 vdd.n2055 0.194439
R10576 vdd.n2849 vdd.n2807 0.194439
R10577 vdd.n2849 vdd.n2808 0.194439
R10578 vdd.n2856 vdd.n2853 0.194439
R10579 vdd.n2856 vdd.n2796 0.194439
R10580 vdd.n2883 vdd.n2874 0.194439
R10581 vdd.n2883 vdd.n2875 0.194439
R10582 vdd.n2879 vdd.n2786 0.194439
R10583 vdd.n4526 vdd.n989 0.194439
R10584 vdd.n4520 vdd.n4519 0.194439
R10585 vdd.n4519 vdd.n1007 0.194439
R10586 vdd.n1062 vdd.n1061 0.194439
R10587 vdd.n1063 vdd.n1062 0.194439
R10588 vdd.n4499 vdd.n1049 0.194439
R10589 vdd.n4499 vdd.n1050 0.194439
R10590 vdd.n4493 vdd.n4492 0.194439
R10591 vdd.n4492 vdd.n1075 0.194439
R10592 vdd.n1138 vdd.n1126 0.194439
R10593 vdd.n1138 vdd.n1137 0.194439
R10594 vdd.n4474 vdd.n1117 0.194439
R10595 vdd.n4474 vdd.n1118 0.194439
R10596 vdd.n1171 vdd.n1144 0.194439
R10597 vdd.n1180 vdd.n1171 0.194439
R10598 vdd.n4452 vdd.n1167 0.194439
R10599 vdd.n4452 vdd.n1168 0.194439
R10600 vdd.n1213 vdd.n1186 0.194439
R10601 vdd.n1222 vdd.n1213 0.194439
R10602 vdd.n4430 vdd.n1209 0.194439
R10603 vdd.n4430 vdd.n1210 0.194439
R10604 vdd.n1261 vdd.n1228 0.194439
R10605 vdd.n1262 vdd.n1261 0.194439
R10606 vdd.n4405 vdd.n1257 0.194439
R10607 vdd.n4405 vdd.n1258 0.194439
R10608 vdd.n4399 vdd.n4398 0.194439
R10609 vdd.n4398 vdd.n1275 0.194439
R10610 vdd.n1326 vdd.n1325 0.194439
R10611 vdd.n1327 vdd.n1326 0.194439
R10612 vdd.n4378 vdd.n1313 0.194439
R10613 vdd.n4378 vdd.n1314 0.194439
R10614 vdd.n4372 vdd.n4371 0.194439
R10615 vdd.n4371 vdd.n1339 0.194439
R10616 vdd.n1402 vdd.n1390 0.194439
R10617 vdd.n1402 vdd.n1401 0.194439
R10618 vdd.n4353 vdd.n1381 0.194439
R10619 vdd.n4353 vdd.n1382 0.194439
R10620 vdd.n1435 vdd.n1408 0.194439
R10621 vdd.n1444 vdd.n1435 0.194439
R10622 vdd.n4331 vdd.n1431 0.194439
R10623 vdd.n4331 vdd.n1432 0.194439
R10624 vdd.n1477 vdd.n1450 0.194439
R10625 vdd.n1486 vdd.n1477 0.194439
R10626 vdd.n4309 vdd.n1473 0.194439
R10627 vdd.n4309 vdd.n1474 0.194439
R10628 vdd.n1525 vdd.n1492 0.194439
R10629 vdd.n1526 vdd.n1525 0.194439
R10630 vdd.n4284 vdd.n1521 0.194439
R10631 vdd.n4284 vdd.n1522 0.194439
R10632 vdd.n4278 vdd.n4277 0.194439
R10633 vdd.n4277 vdd.n1539 0.194439
R10634 vdd.n1590 vdd.n1589 0.194439
R10635 vdd.n1591 vdd.n1590 0.194439
R10636 vdd.n4257 vdd.n1577 0.194439
R10637 vdd.n4257 vdd.n1578 0.194439
R10638 vdd.n4251 vdd.n4250 0.194439
R10639 vdd.n4250 vdd.n1603 0.194439
R10640 vdd.n1666 vdd.n1654 0.194439
R10641 vdd.n1666 vdd.n1665 0.194439
R10642 vdd.n4232 vdd.n1645 0.194439
R10643 vdd.n4232 vdd.n1646 0.194439
R10644 vdd.n1699 vdd.n1672 0.194439
R10645 vdd.n1708 vdd.n1699 0.194439
R10646 vdd.n4210 vdd.n1695 0.194439
R10647 vdd.n4210 vdd.n1696 0.194439
R10648 vdd.n1741 vdd.n1714 0.194439
R10649 vdd.n1750 vdd.n1741 0.194439
R10650 vdd.n4188 vdd.n1737 0.194439
R10651 vdd.n4188 vdd.n1738 0.194439
R10652 vdd.n1789 vdd.n1756 0.194439
R10653 vdd.n1790 vdd.n1789 0.194439
R10654 vdd.n4163 vdd.n1785 0.194439
R10655 vdd.n4163 vdd.n1786 0.194439
R10656 vdd.n4157 vdd.n4156 0.194439
R10657 vdd.n4156 vdd.n1803 0.194439
R10658 vdd.n1854 vdd.n1853 0.194439
R10659 vdd.n1855 vdd.n1854 0.194439
R10660 vdd.n4136 vdd.n1841 0.194439
R10661 vdd.n4136 vdd.n1842 0.194439
R10662 vdd.n4130 vdd.n4129 0.194439
R10663 vdd.n4129 vdd.n1867 0.194439
R10664 vdd.n1930 vdd.n1918 0.194439
R10665 vdd.n1930 vdd.n1929 0.194439
R10666 vdd.n4111 vdd.n1909 0.194439
R10667 vdd.n4111 vdd.n1910 0.194439
R10668 vdd.n1963 vdd.n1936 0.194439
R10669 vdd.n1972 vdd.n1963 0.194439
R10670 vdd.n4089 vdd.n1959 0.194439
R10671 vdd.n4089 vdd.n1960 0.194439
R10672 vdd.n2005 vdd.n1978 0.194439
R10673 vdd.n2014 vdd.n2005 0.194439
R10674 vdd.n4067 vdd.n2001 0.194439
R10675 vdd.n4067 vdd.n2002 0.194439
R10676 vdd.n3919 vdd.n2020 0.194439
R10677 vdd.n4579 vdd.n4578 0.194439
R10678 vdd.n4578 vdd.n853 0.194439
R10679 vdd.n4572 vdd.n4571 0.194439
R10680 vdd.n4571 vdd.n859 0.194439
R10681 vdd.n935 vdd.n934 0.194439
R10682 vdd.n936 vdd.n935 0.194439
R10683 vdd.n4551 vdd.n922 0.194439
R10684 vdd.n4551 vdd.n923 0.194439
R10685 vdd.n4545 vdd.n4544 0.194439
R10686 vdd.n4544 vdd.n948 0.194439
R10687 vdd.n999 vdd.n998 0.194439
R10688 vdd.n4679 vdd.n799 0.194439
R10689 vdd.n4700 vdd.n797 0.194439
R10690 vdd.n4700 vdd.n786 0.194439
R10691 vdd.n4725 vdd.n784 0.194439
R10692 vdd.n784 vdd.n783 0.194439
R10693 vdd.n4754 vdd.n770 0.194439
R10694 vdd.n4754 vdd.n771 0.194439
R10695 vdd.n4761 vdd.n4760 0.194439
R10696 vdd.n4761 vdd.n759 0.194439
R10697 vdd.n4782 vdd.n739 0.194439
R10698 vdd.n4782 vdd.n757 0.194439
R10699 vdd.n749 vdd.n748 0.194439
R10700 vdd.n748 vdd.n744 0.194439
R10701 vdd.n4806 vdd.n4805 0.194439
R10702 vdd.n4806 vdd.n724 0.194439
R10703 vdd.n4837 vdd.n708 0.194439
R10704 vdd.n4838 vdd.n4837 0.194439
R10705 vdd.n4844 vdd.n705 0.194439
R10706 vdd.n4844 vdd.n692 0.194439
R10707 vdd.n693 vdd.n690 0.194439
R10708 vdd.n4867 vdd.n690 0.194439
R10709 vdd.n4897 vdd.n675 0.194439
R10710 vdd.n4897 vdd.n673 0.194439
R10711 vdd.n4907 vdd.n4906 0.194439
R10712 vdd.n4907 vdd.n664 0.194439
R10713 vdd.n4928 vdd.n662 0.194439
R10714 vdd.n4928 vdd.n651 0.194439
R10715 vdd.n4953 vdd.n649 0.194439
R10716 vdd.n649 vdd.n648 0.194439
R10717 vdd.n4982 vdd.n635 0.194439
R10718 vdd.n4982 vdd.n636 0.194439
R10719 vdd.n4989 vdd.n4988 0.194439
R10720 vdd.n4989 vdd.n624 0.194439
R10721 vdd.n5010 vdd.n604 0.194439
R10722 vdd.n5010 vdd.n622 0.194439
R10723 vdd.n614 vdd.n613 0.194439
R10724 vdd.n613 vdd.n609 0.194439
R10725 vdd.n5034 vdd.n5033 0.194439
R10726 vdd.n5034 vdd.n589 0.194439
R10727 vdd.n5065 vdd.n573 0.194439
R10728 vdd.n5066 vdd.n5065 0.194439
R10729 vdd.n5072 vdd.n570 0.194439
R10730 vdd.n5072 vdd.n557 0.194439
R10731 vdd.n558 vdd.n555 0.194439
R10732 vdd.n5095 vdd.n555 0.194439
R10733 vdd.n5125 vdd.n540 0.194439
R10734 vdd.n5125 vdd.n538 0.194439
R10735 vdd.n5135 vdd.n5134 0.194439
R10736 vdd.n5135 vdd.n529 0.194439
R10737 vdd.n5156 vdd.n527 0.194439
R10738 vdd.n5156 vdd.n516 0.194439
R10739 vdd.n5181 vdd.n514 0.194439
R10740 vdd.n514 vdd.n513 0.194439
R10741 vdd.n5210 vdd.n500 0.194439
R10742 vdd.n5210 vdd.n501 0.194439
R10743 vdd.n5217 vdd.n5216 0.194439
R10744 vdd.n5217 vdd.n489 0.194439
R10745 vdd.n5238 vdd.n469 0.194439
R10746 vdd.n5238 vdd.n487 0.194439
R10747 vdd.n479 vdd.n478 0.194439
R10748 vdd.n478 vdd.n474 0.194439
R10749 vdd.n5262 vdd.n5261 0.194439
R10750 vdd.n5262 vdd.n454 0.194439
R10751 vdd.n5293 vdd.n438 0.194439
R10752 vdd.n5294 vdd.n5293 0.194439
R10753 vdd.n5300 vdd.n435 0.194439
R10754 vdd.n5300 vdd.n422 0.194439
R10755 vdd.n423 vdd.n420 0.194439
R10756 vdd.n5323 vdd.n420 0.194439
R10757 vdd.n5353 vdd.n405 0.194439
R10758 vdd.n5353 vdd.n403 0.194439
R10759 vdd.n5363 vdd.n5362 0.194439
R10760 vdd.n5363 vdd.n394 0.194439
R10761 vdd.n5384 vdd.n392 0.194439
R10762 vdd.n5384 vdd.n381 0.194439
R10763 vdd.n5409 vdd.n379 0.194439
R10764 vdd.n379 vdd.n378 0.194439
R10765 vdd.n5438 vdd.n365 0.194439
R10766 vdd.n5438 vdd.n366 0.194439
R10767 vdd.n5445 vdd.n5444 0.194439
R10768 vdd.n5445 vdd.n354 0.194439
R10769 vdd.n5465 vdd.n343 0.194439
R10770 vdd.n5465 vdd.n352 0.194439
R10771 vdd.n5478 vdd.n333 0.194439
R10772 vdd.n5482 vdd.n5478 0.194439
R10773 vdd.n5500 vdd.n325 0.194439
R10774 vdd.n5500 vdd.n323 0.194439
R10775 vdd.n5508 vdd.n5507 0.194439
R10776 vdd.n5507 vdd.n320 0.194439
R10777 vdd.n5535 vdd.n5534 0.194439
R10778 vdd.n5535 vdd.n303 0.194439
R10779 vdd.n5570 vdd.n285 0.194439
R10780 vdd.n5571 vdd.n5570 0.194439
R10781 vdd.n5576 vdd.n282 0.194439
R10782 vdd.n2179 vdd.n2178 0.172719
R10783 vdd.n7417 vdd 0.152702
R10784 vdd.n2130 vdd.n2129 0.132423
R10785 vdd.n7422 vdd.n7421 0.132407
R10786 vdd.n5732 vdd.n5731 0.132407
R10787 vdd.n4011 vdd.n4010 0.13107
R10788 vdd.n883 vdd.n876 0.13107
R10789 vdd.n7421 vdd.n5791 0.127283
R10790 vdd.n5732 vdd.n246 0.127283
R10791 vdd.n4012 vdd.n4011 0.127283
R10792 vdd.n884 vdd.n883 0.127283
R10793 vdd.n7518 vdd 0.123643
R10794 vdd.n33 vdd.n29 0.120292
R10795 vdd.n37 vdd.n33 0.120292
R10796 vdd.n43 vdd.n37 0.120292
R10797 vdd.n47 vdd.n43 0.120292
R10798 vdd.n7416 vdd 0.1039
R10799 vdd.n6503 vdd.n6320 0.102103
R10800 vdd.n6730 vdd.n6187 0.102103
R10801 vdd.n6957 vdd.n6054 0.102103
R10802 vdd.n7184 vdd.n5921 0.102103
R10803 vdd.n4788 vdd.n4786 0.102103
R10804 vdd.n5016 vdd.n5014 0.102103
R10805 vdd.n5244 vdd.n5242 0.102103
R10806 vdd.n5469 vdd.n336 0.102103
R10807 vdd.n3014 vdd.n3012 0.102103
R10808 vdd.n3242 vdd.n3240 0.102103
R10809 vdd.n3470 vdd.n3468 0.102103
R10810 vdd.n3695 vdd.n2312 0.102103
R10811 vdd.n4479 vdd.n4478 0.102103
R10812 vdd.n4358 vdd.n4357 0.102103
R10813 vdd.n4237 vdd.n4236 0.102103
R10814 vdd.n4116 vdd.n4115 0.102103
R10815 vdd.n6619 vdd.n6258 0.100721
R10816 vdd.n6846 vdd.n6125 0.100721
R10817 vdd.n7073 vdd.n5992 0.100721
R10818 vdd.n4891 vdd.n682 0.100721
R10819 vdd.n5119 vdd.n547 0.100721
R10820 vdd.n5347 vdd.n412 0.100721
R10821 vdd.n3117 vdd.n2658 0.100721
R10822 vdd.n3345 vdd.n2523 0.100721
R10823 vdd.n3573 vdd.n2388 0.100721
R10824 vdd.n4413 vdd.n4412 0.100721
R10825 vdd.n4292 vdd.n4291 0.100721
R10826 vdd.n4171 vdd.n4170 0.100721
R10827 vdd.n162 vdd.n161 0.0989615
R10828 vdd.n172 vdd.n171 0.0989615
R10829 vdd.n166 vdd.n165 0.0989615
R10830 vdd.n17 vdd.n14 0.0989615
R10831 vdd.n7490 vdd.n210 0.0981562
R10832 vdd.n5757 vdd.n241 0.0981562
R10833 vdd.n3984 vdd.n3853 0.0877396
R10834 vdd.n4626 vdd.n843 0.0877396
R10835 vdd.n7232 vdd.n7231 0.0847059
R10836 vdd.n7267 vdd.n7266 0.0847059
R10837 vdd.n7005 vdd.n7004 0.0847059
R10838 vdd.n7040 vdd.n7039 0.0847059
R10839 vdd.n6778 vdd.n6777 0.0847059
R10840 vdd.n6813 vdd.n6812 0.0847059
R10841 vdd.n6551 vdd.n6550 0.0847059
R10842 vdd.n6586 vdd.n6585 0.0847059
R10843 vdd.n6428 vdd.n6374 0.0847059
R10844 vdd.n7320 vdd.n7319 0.0847059
R10845 vdd.n7339 vdd.n7338 0.0847059
R10846 vdd.n7358 vdd.n7357 0.0847059
R10847 vdd.n7377 vdd.n7376 0.0847059
R10848 vdd.n5502 vdd.n5501 0.0847059
R10849 vdd.n5537 vdd.n5536 0.0847059
R10850 vdd.n5264 vdd.n5263 0.0847059
R10851 vdd.n5299 vdd.n5298 0.0847059
R10852 vdd.n5355 vdd.n5354 0.0847059
R10853 vdd.n5036 vdd.n5035 0.0847059
R10854 vdd.n5071 vdd.n5070 0.0847059
R10855 vdd.n5127 vdd.n5126 0.0847059
R10856 vdd.n4808 vdd.n4807 0.0847059
R10857 vdd.n4843 vdd.n4842 0.0847059
R10858 vdd.n4899 vdd.n4898 0.0847059
R10859 vdd.n3726 vdd.n3725 0.0847059
R10860 vdd.n3761 vdd.n3760 0.0847059
R10861 vdd.n3490 vdd.n3489 0.0847059
R10862 vdd.n3525 vdd.n3524 0.0847059
R10863 vdd.n3581 vdd.n3580 0.0847059
R10864 vdd.n3262 vdd.n3261 0.0847059
R10865 vdd.n3297 vdd.n3296 0.0847059
R10866 vdd.n3353 vdd.n3352 0.0847059
R10867 vdd.n3034 vdd.n3033 0.0847059
R10868 vdd.n3069 vdd.n3068 0.0847059
R10869 vdd.n3125 vdd.n3124 0.0847059
R10870 vdd.n3668 vdd.n2329 0.0847059
R10871 vdd.n3638 vdd.n3637 0.0847059
R10872 vdd.n3440 vdd.n2464 0.0847059
R10873 vdd.n3410 vdd.n3409 0.0847059
R10874 vdd.n3212 vdd.n2599 0.0847059
R10875 vdd.n3182 vdd.n3181 0.0847059
R10876 vdd.n2984 vdd.n2734 0.0847059
R10877 vdd.n2954 vdd.n2953 0.0847059
R10878 vdd.n2850 vdd.n2059 0.0847059
R10879 vdd.n2882 vdd.n2062 0.0847059
R10880 vdd.n5442 vdd.n353 0.0847059
R10881 vdd.n5412 vdd.n5411 0.0847059
R10882 vdd.n5214 vdd.n488 0.0847059
R10883 vdd.n5184 vdd.n5183 0.0847059
R10884 vdd.n4986 vdd.n623 0.0847059
R10885 vdd.n4956 vdd.n4955 0.0847059
R10886 vdd.n4758 vdd.n758 0.0847059
R10887 vdd.n4728 vdd.n4727 0.0847059
R10888 vdd.n5665 vdd.n254 0.0847059
R10889 vdd.n5699 vdd.n256 0.0847059
R10890 vdd.n5721 vdd.n258 0.0847059
R10891 vdd.n5618 vdd.n252 0.0847059
R10892 vdd.n7406 vdd.n5792 0.0796667
R10893 vdd.n5653 vdd.n245 0.0796667
R10894 vdd.n4042 vdd.n4041 0.0796667
R10895 vdd.n886 vdd.n875 0.0796667
R10896 vdd.n3944 vdd.t20 0.074533
R10897 vdd.n6413 vdd.n6376 0.0705758
R10898 vdd.n6434 vdd.n6362 0.0705758
R10899 vdd.n6449 vdd.n6357 0.0705758
R10900 vdd.n6472 vdd.n6346 0.0705758
R10901 vdd.n6492 vdd.n6325 0.0705758
R10902 vdd.n6525 vdd.n6311 0.0705758
R10903 vdd.n6544 vdd.n6543 0.0705758
R10904 vdd.n6561 vdd.n6560 0.0705758
R10905 vdd.n6578 vdd.n6287 0.0705758
R10906 vdd.n6599 vdd.n6271 0.0705758
R10907 vdd.n6640 vdd.n6243 0.0705758
R10908 vdd.n6661 vdd.n6229 0.0705758
R10909 vdd.n6676 vdd.n6224 0.0705758
R10910 vdd.n6699 vdd.n6213 0.0705758
R10911 vdd.n6719 vdd.n6192 0.0705758
R10912 vdd.n6752 vdd.n6178 0.0705758
R10913 vdd.n6771 vdd.n6770 0.0705758
R10914 vdd.n6788 vdd.n6787 0.0705758
R10915 vdd.n6805 vdd.n6154 0.0705758
R10916 vdd.n6826 vdd.n6138 0.0705758
R10917 vdd.n6867 vdd.n6110 0.0705758
R10918 vdd.n6888 vdd.n6096 0.0705758
R10919 vdd.n6903 vdd.n6091 0.0705758
R10920 vdd.n6926 vdd.n6080 0.0705758
R10921 vdd.n6946 vdd.n6059 0.0705758
R10922 vdd.n6979 vdd.n6045 0.0705758
R10923 vdd.n6998 vdd.n6997 0.0705758
R10924 vdd.n7015 vdd.n7014 0.0705758
R10925 vdd.n7032 vdd.n6021 0.0705758
R10926 vdd.n7053 vdd.n6005 0.0705758
R10927 vdd.n7094 vdd.n5977 0.0705758
R10928 vdd.n7115 vdd.n5963 0.0705758
R10929 vdd.n7130 vdd.n5958 0.0705758
R10930 vdd.n7153 vdd.n5947 0.0705758
R10931 vdd.n7173 vdd.n5926 0.0705758
R10932 vdd.n7206 vdd.n5912 0.0705758
R10933 vdd.n7225 vdd.n7224 0.0705758
R10934 vdd.n7242 vdd.n7241 0.0705758
R10935 vdd.n7259 vdd.n5888 0.0705758
R10936 vdd.n7285 vdd.n5871 0.0705758
R10937 vdd.n7314 vdd.n5860 0.0705758
R10938 vdd.n7333 vdd.n5849 0.0705758
R10939 vdd.n7352 vdd.n5838 0.0705758
R10940 vdd.n7371 vdd.n5827 0.0705758
R10941 vdd.n7394 vdd.n5815 0.0705758
R10942 vdd.n4691 vdd.n796 0.0705758
R10943 vdd.n4721 vdd.n788 0.0705758
R10944 vdd.n4734 vdd.n772 0.0705758
R10945 vdd.n4749 vdd.n767 0.0705758
R10946 vdd.n4774 vdd.n737 0.0705758
R10947 vdd.n4801 vdd.n4800 0.0705758
R10948 vdd.n4818 vdd.n4817 0.0705758
R10949 vdd.n4835 vdd.n713 0.0705758
R10950 vdd.n704 vdd.n694 0.0705758
R10951 vdd.n4874 vdd.n4873 0.0705758
R10952 vdd.n4919 vdd.n661 0.0705758
R10953 vdd.n4949 vdd.n653 0.0705758
R10954 vdd.n4962 vdd.n637 0.0705758
R10955 vdd.n4977 vdd.n632 0.0705758
R10956 vdd.n5002 vdd.n602 0.0705758
R10957 vdd.n5029 vdd.n5028 0.0705758
R10958 vdd.n5046 vdd.n5045 0.0705758
R10959 vdd.n5063 vdd.n578 0.0705758
R10960 vdd.n569 vdd.n559 0.0705758
R10961 vdd.n5102 vdd.n5101 0.0705758
R10962 vdd.n5147 vdd.n526 0.0705758
R10963 vdd.n5177 vdd.n518 0.0705758
R10964 vdd.n5190 vdd.n502 0.0705758
R10965 vdd.n5205 vdd.n497 0.0705758
R10966 vdd.n5230 vdd.n467 0.0705758
R10967 vdd.n5257 vdd.n5256 0.0705758
R10968 vdd.n5274 vdd.n5273 0.0705758
R10969 vdd.n5291 vdd.n443 0.0705758
R10970 vdd.n434 vdd.n424 0.0705758
R10971 vdd.n5330 vdd.n5329 0.0705758
R10972 vdd.n5375 vdd.n391 0.0705758
R10973 vdd.n5405 vdd.n383 0.0705758
R10974 vdd.n5418 vdd.n367 0.0705758
R10975 vdd.n5433 vdd.n362 0.0705758
R10976 vdd.n5457 vdd.n341 0.0705758
R10977 vdd.n5486 vdd.n332 0.0705758
R10978 vdd.n5511 vdd.n316 0.0705758
R10979 vdd.n5530 vdd.n5529 0.0705758
R10980 vdd.n5547 vdd.n5546 0.0705758
R10981 vdd.n5568 vdd.n290 0.0705758
R10982 vdd.n5591 vdd.n5590 0.0705758
R10983 vdd.n5718 vdd.n268 0.0705758
R10984 vdd.n5706 vdd.n5705 0.0705758
R10985 vdd.n5641 vdd.n5625 0.0705758
R10986 vdd.n5675 vdd.n5671 0.0705758
R10987 vdd.n2917 vdd.n2772 0.0705758
R10988 vdd.n2947 vdd.n2764 0.0705758
R10989 vdd.n2960 vdd.n2748 0.0705758
R10990 vdd.n2975 vdd.n2743 0.0705758
R10991 vdd.n3000 vdd.n2713 0.0705758
R10992 vdd.n3027 vdd.n3026 0.0705758
R10993 vdd.n3044 vdd.n3043 0.0705758
R10994 vdd.n3061 vdd.n2689 0.0705758
R10995 vdd.n2680 vdd.n2670 0.0705758
R10996 vdd.n3100 vdd.n3099 0.0705758
R10997 vdd.n3145 vdd.n2637 0.0705758
R10998 vdd.n3175 vdd.n2629 0.0705758
R10999 vdd.n3188 vdd.n2613 0.0705758
R11000 vdd.n3203 vdd.n2608 0.0705758
R11001 vdd.n3228 vdd.n2578 0.0705758
R11002 vdd.n3255 vdd.n3254 0.0705758
R11003 vdd.n3272 vdd.n3271 0.0705758
R11004 vdd.n3289 vdd.n2554 0.0705758
R11005 vdd.n2545 vdd.n2535 0.0705758
R11006 vdd.n3328 vdd.n3327 0.0705758
R11007 vdd.n3373 vdd.n2502 0.0705758
R11008 vdd.n3403 vdd.n2494 0.0705758
R11009 vdd.n3416 vdd.n2478 0.0705758
R11010 vdd.n3431 vdd.n2473 0.0705758
R11011 vdd.n3456 vdd.n2443 0.0705758
R11012 vdd.n3483 vdd.n3482 0.0705758
R11013 vdd.n3500 vdd.n3499 0.0705758
R11014 vdd.n3517 vdd.n2419 0.0705758
R11015 vdd.n2410 vdd.n2400 0.0705758
R11016 vdd.n3556 vdd.n3555 0.0705758
R11017 vdd.n3601 vdd.n2367 0.0705758
R11018 vdd.n3631 vdd.n2359 0.0705758
R11019 vdd.n3644 vdd.n2343 0.0705758
R11020 vdd.n3659 vdd.n2338 0.0705758
R11021 vdd.n3683 vdd.n2317 0.0705758
R11022 vdd.n3711 vdd.n2307 0.0705758
R11023 vdd.n3735 vdd.n2290 0.0705758
R11024 vdd.n3754 vdd.n3753 0.0705758
R11025 vdd.n3771 vdd.n3770 0.0705758
R11026 vdd.n3792 vdd.n2264 0.0705758
R11027 vdd.n4030 vdd.n2051 0.0705758
R11028 vdd.n2829 vdd.n2809 0.0705758
R11029 vdd.n2844 vdd.n2804 0.0705758
R11030 vdd.n2868 vdd.n2794 0.0705758
R11031 vdd.n2895 vdd.n2787 0.0705758
R11032 vdd.n1026 vdd.n1008 0.0705758
R11033 vdd.n4514 vdd.n4513 0.0705758
R11034 vdd.n4501 vdd.n1046 0.0705758
R11035 vdd.n1095 vdd.n1076 0.0705758
R11036 vdd.n4487 vdd.n4486 0.0705758
R11037 vdd.n1145 vdd.n1116 0.0705758
R11038 vdd.n1176 vdd.n1172 0.0705758
R11039 vdd.n1187 vdd.n1166 0.0705758
R11040 vdd.n1218 vdd.n1214 0.0705758
R11041 vdd.n1229 vdd.n1208 0.0705758
R11042 vdd.n1290 vdd.n1276 0.0705758
R11043 vdd.n4393 vdd.n4392 0.0705758
R11044 vdd.n4380 vdd.n1310 0.0705758
R11045 vdd.n1359 vdd.n1340 0.0705758
R11046 vdd.n4366 vdd.n4365 0.0705758
R11047 vdd.n1409 vdd.n1380 0.0705758
R11048 vdd.n1440 vdd.n1436 0.0705758
R11049 vdd.n1451 vdd.n1430 0.0705758
R11050 vdd.n1482 vdd.n1478 0.0705758
R11051 vdd.n1493 vdd.n1472 0.0705758
R11052 vdd.n1554 vdd.n1540 0.0705758
R11053 vdd.n4272 vdd.n4271 0.0705758
R11054 vdd.n4259 vdd.n1574 0.0705758
R11055 vdd.n1623 vdd.n1604 0.0705758
R11056 vdd.n4245 vdd.n4244 0.0705758
R11057 vdd.n1673 vdd.n1644 0.0705758
R11058 vdd.n1704 vdd.n1700 0.0705758
R11059 vdd.n1715 vdd.n1694 0.0705758
R11060 vdd.n1746 vdd.n1742 0.0705758
R11061 vdd.n1757 vdd.n1736 0.0705758
R11062 vdd.n1818 vdd.n1804 0.0705758
R11063 vdd.n4151 vdd.n4150 0.0705758
R11064 vdd.n4138 vdd.n1838 0.0705758
R11065 vdd.n1887 vdd.n1868 0.0705758
R11066 vdd.n4124 vdd.n4123 0.0705758
R11067 vdd.n1937 vdd.n1908 0.0705758
R11068 vdd.n1968 vdd.n1964 0.0705758
R11069 vdd.n1979 vdd.n1958 0.0705758
R11070 vdd.n2010 vdd.n2006 0.0705758
R11071 vdd.n2021 vdd.n2000 0.0705758
R11072 vdd.n899 vdd.n860 0.0705758
R11073 vdd.n4566 vdd.n4565 0.0705758
R11074 vdd.n4553 vdd.n919 0.0705758
R11075 vdd.n968 vdd.n949 0.0705758
R11076 vdd.n4539 vdd.n4538 0.0705758
R11077 vdd vdd.n4631 0.0693134
R11078 vdd.n4532 vdd 0.066192
R11079 vdd vdd.n2899 0.066192
R11080 vdd.n4000 vdd.n3999 0.063
R11081 vdd.n4608 vdd.n4606 0.063
R11082 vdd.n7514 vdd.n191 0.0616979
R11083 vdd.n3985 vdd.n3984 0.0616979
R11084 vdd.n4627 vdd.n4626 0.0616979
R11085 vdd.n7477 vdd.n216 0.0616979
R11086 vdd vdd.n191 0.0603958
R11087 vdd vdd.n3839 0.0603958
R11088 vdd vdd.n4612 0.0603958
R11089 vdd vdd.n216 0.0603958
R11090 vdd.n113 vdd.n109 0.0603958
R11091 vdd.n109 vdd.n105 0.0603958
R11092 vdd.n92 vdd.n88 0.0603958
R11093 vdd.n77 vdd.n74 0.0603958
R11094 vdd.n63 vdd.n59 0.0603958
R11095 vdd.n137 vdd.n133 0.0603958
R11096 vdd.n158 vdd.n154 0.0603958
R11097 vdd.n163 vdd.n158 0.0603958
R11098 vdd.n178 vdd.n173 0.0603958
R11099 vdd.n19 vdd.n18 0.0603958
R11100 vdd.n7514 vdd.n7513 0.0590938
R11101 vdd.n7478 vdd.n7477 0.0590938
R11102 vdd.n48 vdd.n47 0.0590938
R11103 vdd.n7491 vdd.n7490 0.0577917
R11104 vdd.n3999 vdd.n3839 0.0577917
R11105 vdd.n4612 vdd.n4606 0.0577917
R11106 vdd.n5751 vdd.n241 0.0577917
R11107 vdd.n6416 vdd.n6414 0.0573182
R11108 vdd.n6436 vdd.n6435 0.0573182
R11109 vdd.n6450 vdd.n6448 0.0573182
R11110 vdd.n6471 vdd.n6470 0.0573182
R11111 vdd.n6491 vdd.n6490 0.0573182
R11112 vdd.n6527 vdd.n6526 0.0573182
R11113 vdd.n6545 vdd.n6302 0.0573182
R11114 vdd.n6559 vdd.n6296 0.0573182
R11115 vdd.n6576 vdd.n6289 0.0573182
R11116 vdd.n6598 vdd.n6597 0.0573182
R11117 vdd.n6643 vdd.n6641 0.0573182
R11118 vdd.n6663 vdd.n6662 0.0573182
R11119 vdd.n6677 vdd.n6675 0.0573182
R11120 vdd.n6698 vdd.n6697 0.0573182
R11121 vdd.n6718 vdd.n6717 0.0573182
R11122 vdd.n6754 vdd.n6753 0.0573182
R11123 vdd.n6772 vdd.n6169 0.0573182
R11124 vdd.n6786 vdd.n6163 0.0573182
R11125 vdd.n6803 vdd.n6156 0.0573182
R11126 vdd.n6825 vdd.n6824 0.0573182
R11127 vdd.n6870 vdd.n6868 0.0573182
R11128 vdd.n6890 vdd.n6889 0.0573182
R11129 vdd.n6904 vdd.n6902 0.0573182
R11130 vdd.n6925 vdd.n6924 0.0573182
R11131 vdd.n6945 vdd.n6944 0.0573182
R11132 vdd.n6981 vdd.n6980 0.0573182
R11133 vdd.n6999 vdd.n6036 0.0573182
R11134 vdd.n7013 vdd.n6030 0.0573182
R11135 vdd.n7030 vdd.n6023 0.0573182
R11136 vdd.n7052 vdd.n7051 0.0573182
R11137 vdd.n7097 vdd.n7095 0.0573182
R11138 vdd.n7117 vdd.n7116 0.0573182
R11139 vdd.n7131 vdd.n7129 0.0573182
R11140 vdd.n7152 vdd.n7151 0.0573182
R11141 vdd.n7172 vdd.n7171 0.0573182
R11142 vdd.n7208 vdd.n7207 0.0573182
R11143 vdd.n7226 vdd.n5903 0.0573182
R11144 vdd.n7240 vdd.n5897 0.0573182
R11145 vdd.n7257 vdd.n5890 0.0573182
R11146 vdd.n7284 vdd.n7282 0.0573182
R11147 vdd.n7313 vdd.n7312 0.0573182
R11148 vdd.n7332 vdd.n7331 0.0573182
R11149 vdd.n7351 vdd.n7350 0.0573182
R11150 vdd.n7370 vdd.n7369 0.0573182
R11151 vdd.n7393 vdd.n7392 0.0573182
R11152 vdd.n5589 vdd.n5586 0.0573182
R11153 vdd.n5716 vdd.n270 0.0573182
R11154 vdd.n5704 vdd.n5607 0.0573182
R11155 vdd.n5643 vdd.n5627 0.0573182
R11156 vdd.n5674 vdd.n5673 0.0573182
R11157 vdd.n2916 vdd.n2915 0.0573182
R11158 vdd.n2946 vdd.n2945 0.0573182
R11159 vdd.n2962 vdd.n2961 0.0573182
R11160 vdd.n2976 vdd.n2974 0.0573182
R11161 vdd.n2999 vdd.n2998 0.0573182
R11162 vdd.n3028 vdd.n2704 0.0573182
R11163 vdd.n3042 vdd.n2698 0.0573182
R11164 vdd.n3059 vdd.n2691 0.0573182
R11165 vdd.n3082 vdd.n3081 0.0573182
R11166 vdd.n3098 vdd.n2664 0.0573182
R11167 vdd.n3144 vdd.n3143 0.0573182
R11168 vdd.n3174 vdd.n3173 0.0573182
R11169 vdd.n3190 vdd.n3189 0.0573182
R11170 vdd.n3204 vdd.n3202 0.0573182
R11171 vdd.n3227 vdd.n3226 0.0573182
R11172 vdd.n3256 vdd.n2569 0.0573182
R11173 vdd.n3270 vdd.n2563 0.0573182
R11174 vdd.n3287 vdd.n2556 0.0573182
R11175 vdd.n3310 vdd.n3309 0.0573182
R11176 vdd.n3326 vdd.n2529 0.0573182
R11177 vdd.n3372 vdd.n3371 0.0573182
R11178 vdd.n3402 vdd.n3401 0.0573182
R11179 vdd.n3418 vdd.n3417 0.0573182
R11180 vdd.n3432 vdd.n3430 0.0573182
R11181 vdd.n3455 vdd.n3454 0.0573182
R11182 vdd.n3484 vdd.n2434 0.0573182
R11183 vdd.n3498 vdd.n2428 0.0573182
R11184 vdd.n3515 vdd.n2421 0.0573182
R11185 vdd.n3538 vdd.n3537 0.0573182
R11186 vdd.n3554 vdd.n2394 0.0573182
R11187 vdd.n3600 vdd.n3599 0.0573182
R11188 vdd.n3630 vdd.n3629 0.0573182
R11189 vdd.n3646 vdd.n3645 0.0573182
R11190 vdd.n3660 vdd.n3658 0.0573182
R11191 vdd.n3682 vdd.n3681 0.0573182
R11192 vdd.n3713 vdd.n3712 0.0573182
R11193 vdd.n3737 vdd.n3736 0.0573182
R11194 vdd.n3755 vdd.n2281 0.0573182
R11195 vdd.n3769 vdd.n2275 0.0573182
R11196 vdd.n3790 vdd.n2267 0.0573182
R11197 vdd.n4032 vdd.n2049 0.0573182
R11198 vdd.n2831 vdd.n2830 0.0573182
R11199 vdd.n2845 vdd.n2843 0.0573182
R11200 vdd.n2867 vdd.n2866 0.0573182
R11201 vdd.n2893 vdd.n2788 0.0573182
R11202 vdd.n1030 vdd.n1027 0.0573182
R11203 vdd.n4515 vdd.n1011 0.0573182
R11204 vdd.n4503 vdd.n1044 0.0573182
R11205 vdd.n1099 vdd.n1096 0.0573182
R11206 vdd.n4488 vdd.n1079 0.0573182
R11207 vdd.n1155 vdd.n1147 0.0573182
R11208 vdd.n1175 vdd.n1174 0.0573182
R11209 vdd.n1197 vdd.n1189 0.0573182
R11210 vdd.n1217 vdd.n1216 0.0573182
R11211 vdd.n1239 vdd.n1231 0.0573182
R11212 vdd.n1294 vdd.n1291 0.0573182
R11213 vdd.n4394 vdd.n1279 0.0573182
R11214 vdd.n4382 vdd.n1308 0.0573182
R11215 vdd.n1363 vdd.n1360 0.0573182
R11216 vdd.n4367 vdd.n1343 0.0573182
R11217 vdd.n1419 vdd.n1411 0.0573182
R11218 vdd.n1439 vdd.n1438 0.0573182
R11219 vdd.n1461 vdd.n1453 0.0573182
R11220 vdd.n1481 vdd.n1480 0.0573182
R11221 vdd.n1503 vdd.n1495 0.0573182
R11222 vdd.n1558 vdd.n1555 0.0573182
R11223 vdd.n4273 vdd.n1543 0.0573182
R11224 vdd.n4261 vdd.n1572 0.0573182
R11225 vdd.n1627 vdd.n1624 0.0573182
R11226 vdd.n4246 vdd.n1607 0.0573182
R11227 vdd.n1683 vdd.n1675 0.0573182
R11228 vdd.n1703 vdd.n1702 0.0573182
R11229 vdd.n1725 vdd.n1717 0.0573182
R11230 vdd.n1745 vdd.n1744 0.0573182
R11231 vdd.n1767 vdd.n1759 0.0573182
R11232 vdd.n1822 vdd.n1819 0.0573182
R11233 vdd.n4152 vdd.n1807 0.0573182
R11234 vdd.n4140 vdd.n1836 0.0573182
R11235 vdd.n1891 vdd.n1888 0.0573182
R11236 vdd.n4125 vdd.n1871 0.0573182
R11237 vdd.n1947 vdd.n1939 0.0573182
R11238 vdd.n1967 vdd.n1966 0.0573182
R11239 vdd.n1989 vdd.n1981 0.0573182
R11240 vdd.n2009 vdd.n2008 0.0573182
R11241 vdd.n2031 vdd.n2023 0.0573182
R11242 vdd.n903 vdd.n900 0.0573182
R11243 vdd.n4567 vdd.n863 0.0573182
R11244 vdd.n4555 vdd.n917 0.0573182
R11245 vdd.n972 vdd.n969 0.0573182
R11246 vdd.n4540 vdd.n952 0.0573182
R11247 vdd.n4690 vdd.n4689 0.0573182
R11248 vdd.n4720 vdd.n4719 0.0573182
R11249 vdd.n4736 vdd.n4735 0.0573182
R11250 vdd.n4750 vdd.n4748 0.0573182
R11251 vdd.n4773 vdd.n4772 0.0573182
R11252 vdd.n4802 vdd.n728 0.0573182
R11253 vdd.n4816 vdd.n722 0.0573182
R11254 vdd.n4833 vdd.n715 0.0573182
R11255 vdd.n4856 vdd.n4855 0.0573182
R11256 vdd.n4872 vdd.n688 0.0573182
R11257 vdd.n4918 vdd.n4917 0.0573182
R11258 vdd.n4948 vdd.n4947 0.0573182
R11259 vdd.n4964 vdd.n4963 0.0573182
R11260 vdd.n4978 vdd.n4976 0.0573182
R11261 vdd.n5001 vdd.n5000 0.0573182
R11262 vdd.n5030 vdd.n593 0.0573182
R11263 vdd.n5044 vdd.n587 0.0573182
R11264 vdd.n5061 vdd.n580 0.0573182
R11265 vdd.n5084 vdd.n5083 0.0573182
R11266 vdd.n5100 vdd.n553 0.0573182
R11267 vdd.n5146 vdd.n5145 0.0573182
R11268 vdd.n5176 vdd.n5175 0.0573182
R11269 vdd.n5192 vdd.n5191 0.0573182
R11270 vdd.n5206 vdd.n5204 0.0573182
R11271 vdd.n5229 vdd.n5228 0.0573182
R11272 vdd.n5258 vdd.n458 0.0573182
R11273 vdd.n5272 vdd.n452 0.0573182
R11274 vdd.n5289 vdd.n445 0.0573182
R11275 vdd.n5312 vdd.n5311 0.0573182
R11276 vdd.n5328 vdd.n418 0.0573182
R11277 vdd.n5374 vdd.n5373 0.0573182
R11278 vdd.n5404 vdd.n5403 0.0573182
R11279 vdd.n5420 vdd.n5419 0.0573182
R11280 vdd.n5434 vdd.n5432 0.0573182
R11281 vdd.n5456 vdd.n5455 0.0573182
R11282 vdd.n5488 vdd.n5487 0.0573182
R11283 vdd.n5513 vdd.n5512 0.0573182
R11284 vdd.n5531 vdd.n307 0.0573182
R11285 vdd.n5545 vdd.n301 0.0573182
R11286 vdd.n5566 vdd.n293 0.0573182
R11287 vdd.n179 vdd.n178 0.0545365
R11288 vdd.n99 vdd.n92 0.0538854
R11289 vdd.n4632 vdd.n838 0.0533411
R11290 vdd.n4047 vdd.n4046 0.0533411
R11291 vdd.n5762 vdd.n238 0.0517727
R11292 vdd.n5737 vdd.n5736 0.0517053
R11293 vdd.n7417 vdd.n7416 0.0517053
R11294 vdd.n3996 vdd.n3842 0.0511623
R11295 vdd.n4603 vdd.n4592 0.0511623
R11296 vdd.n7414 vdd 0.0508121
R11297 vdd.n18 vdd.n6 0.0506302
R11298 vdd.n84 vdd.n77 0.0493281
R11299 vdd.n114 vdd.n53 0.048026
R11300 vdd.n70 vdd.n63 0.048026
R11301 vdd.n2153 vdd.n2106 0.0476312
R11302 vdd.n2189 vdd.n2184 0.0476312
R11303 vdd.n2198 vdd.n2166 0.045582
R11304 vdd.n7420 vdd.n5792 0.0455
R11305 vdd.n5733 vdd.n245 0.0455
R11306 vdd.n4042 vdd.n2038 0.0455
R11307 vdd.n882 vdd.n875 0.0455
R11308 vdd.n3850 vdd.n3844 0.0438377
R11309 vdd.n4594 vdd.n4593 0.0438377
R11310 vdd.n7474 vdd.n219 0.0438377
R11311 vdd.n5591 vdd.n261 0.0434423
R11312 vdd.n2896 vdd.n2895 0.0429349
R11313 vdd.n4538 vdd.n953 0.0429349
R11314 vdd.n7302 vdd.n5860 0.0429036
R11315 vdd.n207 vdd.n203 0.041625
R11316 vdd.n3995 vdd.n3994 0.041625
R11317 vdd.n4602 vdd.n4601 0.041625
R11318 vdd.n5760 vdd.n239 0.041625
R11319 vdd.n2139 vdd.n2134 0.0414836
R11320 vdd vdd.n4673 0.0410684
R11321 vdd vdd.n6395 0.0410684
R11322 vdd.n7491 vdd 0.0408646
R11323 vdd vdd.n5751 0.0408646
R11324 vdd.n6426 vdd.n6376 0.0402727
R11325 vdd.n6453 vdd.n6362 0.0402727
R11326 vdd.n6461 vdd.n6357 0.0402727
R11327 vdd.n6481 vdd.n6346 0.0402727
R11328 vdd.n6500 vdd.n6325 0.0402727
R11329 vdd.n6512 vdd.n6311 0.0402727
R11330 vdd.n6543 vdd.n6303 0.0402727
R11331 vdd.n6561 vdd.n6297 0.0402727
R11332 vdd.n6579 vdd.n6578 0.0402727
R11333 vdd.n6588 vdd.n6271 0.0402727
R11334 vdd.n6612 vdd.n6266 0.0402727
R11335 vdd.n6632 vdd.n6254 0.0402727
R11336 vdd.n6653 vdd.n6243 0.0402727
R11337 vdd.n6680 vdd.n6229 0.0402727
R11338 vdd.n6688 vdd.n6224 0.0402727
R11339 vdd.n6708 vdd.n6213 0.0402727
R11340 vdd.n6727 vdd.n6192 0.0402727
R11341 vdd.n6739 vdd.n6178 0.0402727
R11342 vdd.n6770 vdd.n6170 0.0402727
R11343 vdd.n6788 vdd.n6164 0.0402727
R11344 vdd.n6806 vdd.n6805 0.0402727
R11345 vdd.n6815 vdd.n6138 0.0402727
R11346 vdd.n6839 vdd.n6133 0.0402727
R11347 vdd.n6859 vdd.n6121 0.0402727
R11348 vdd.n6880 vdd.n6110 0.0402727
R11349 vdd.n6907 vdd.n6096 0.0402727
R11350 vdd.n6915 vdd.n6091 0.0402727
R11351 vdd.n6935 vdd.n6080 0.0402727
R11352 vdd.n6954 vdd.n6059 0.0402727
R11353 vdd.n6966 vdd.n6045 0.0402727
R11354 vdd.n6997 vdd.n6037 0.0402727
R11355 vdd.n7015 vdd.n6031 0.0402727
R11356 vdd.n7033 vdd.n7032 0.0402727
R11357 vdd.n7042 vdd.n6005 0.0402727
R11358 vdd.n7066 vdd.n6000 0.0402727
R11359 vdd.n7086 vdd.n5988 0.0402727
R11360 vdd.n7107 vdd.n5977 0.0402727
R11361 vdd.n7134 vdd.n5963 0.0402727
R11362 vdd.n7142 vdd.n5958 0.0402727
R11363 vdd.n7162 vdd.n5947 0.0402727
R11364 vdd.n7181 vdd.n5926 0.0402727
R11365 vdd.n7193 vdd.n5912 0.0402727
R11366 vdd.n7224 vdd.n5904 0.0402727
R11367 vdd.n7242 vdd.n5898 0.0402727
R11368 vdd.n7260 vdd.n7259 0.0402727
R11369 vdd.n7269 vdd.n5871 0.0402727
R11370 vdd.n6414 vdd.n6382 0.0402727
R11371 vdd.n6435 vdd.n6371 0.0402727
R11372 vdd.n6451 vdd.n6450 0.0402727
R11373 vdd.n6471 vdd.n6351 0.0402727
R11374 vdd.n6491 vdd.n6340 0.0402727
R11375 vdd.n6332 vdd.n6324 0.0402727
R11376 vdd.n6331 vdd.n6319 0.0402727
R11377 vdd.n6526 vdd.n6310 0.0402727
R11378 vdd.n6546 vdd.n6545 0.0402727
R11379 vdd.n6559 vdd.n6558 0.0402727
R11380 vdd.n6289 vdd.n6276 0.0402727
R11381 vdd.n6598 vdd.n6263 0.0402727
R11382 vdd.n6641 vdd.n6249 0.0402727
R11383 vdd.n6662 vdd.n6238 0.0402727
R11384 vdd.n6678 vdd.n6677 0.0402727
R11385 vdd.n6698 vdd.n6218 0.0402727
R11386 vdd.n6718 vdd.n6207 0.0402727
R11387 vdd.n6199 vdd.n6191 0.0402727
R11388 vdd.n6198 vdd.n6186 0.0402727
R11389 vdd.n6753 vdd.n6177 0.0402727
R11390 vdd.n6773 vdd.n6772 0.0402727
R11391 vdd.n6786 vdd.n6785 0.0402727
R11392 vdd.n6156 vdd.n6143 0.0402727
R11393 vdd.n6825 vdd.n6130 0.0402727
R11394 vdd.n6868 vdd.n6116 0.0402727
R11395 vdd.n6889 vdd.n6105 0.0402727
R11396 vdd.n6905 vdd.n6904 0.0402727
R11397 vdd.n6925 vdd.n6085 0.0402727
R11398 vdd.n6945 vdd.n6074 0.0402727
R11399 vdd.n6066 vdd.n6058 0.0402727
R11400 vdd.n6065 vdd.n6053 0.0402727
R11401 vdd.n6980 vdd.n6044 0.0402727
R11402 vdd.n7000 vdd.n6999 0.0402727
R11403 vdd.n7013 vdd.n7012 0.0402727
R11404 vdd.n6023 vdd.n6010 0.0402727
R11405 vdd.n7052 vdd.n5997 0.0402727
R11406 vdd.n7095 vdd.n5983 0.0402727
R11407 vdd.n7116 vdd.n5972 0.0402727
R11408 vdd.n7132 vdd.n7131 0.0402727
R11409 vdd.n7152 vdd.n5952 0.0402727
R11410 vdd.n7172 vdd.n5941 0.0402727
R11411 vdd.n5933 vdd.n5925 0.0402727
R11412 vdd.n5932 vdd.n5920 0.0402727
R11413 vdd.n7207 vdd.n5911 0.0402727
R11414 vdd.n7227 vdd.n7226 0.0402727
R11415 vdd.n7240 vdd.n7239 0.0402727
R11416 vdd.n5890 vdd.n5877 0.0402727
R11417 vdd.n7284 vdd.n7283 0.0402727
R11418 vdd.n7322 vdd.n5849 0.0402727
R11419 vdd.n7341 vdd.n5838 0.0402727
R11420 vdd.n7360 vdd.n5827 0.0402727
R11421 vdd.n7379 vdd.n5815 0.0402727
R11422 vdd.n7402 vdd.n5791 0.0402727
R11423 vdd.n7313 vdd.n5854 0.0402727
R11424 vdd.n7332 vdd.n5843 0.0402727
R11425 vdd.n7351 vdd.n5832 0.0402727
R11426 vdd.n7370 vdd.n5821 0.0402727
R11427 vdd.n7393 vdd.n5796 0.0402727
R11428 vdd.n4701 vdd.n796 0.0402727
R11429 vdd.n4714 vdd.n788 0.0402727
R11430 vdd.n4753 vdd.n772 0.0402727
R11431 vdd.n4762 vdd.n767 0.0402727
R11432 vdd.n4783 vdd.n737 0.0402727
R11433 vdd.n4800 vdd.n729 0.0402727
R11434 vdd.n4818 vdd.n723 0.0402727
R11435 vdd.n4836 vdd.n4835 0.0402727
R11436 vdd.n4845 vdd.n704 0.0402727
R11437 vdd.n4874 vdd.n689 0.0402727
R11438 vdd.n4896 vdd.n4895 0.0402727
R11439 vdd.n4908 vdd.n672 0.0402727
R11440 vdd.n4929 vdd.n661 0.0402727
R11441 vdd.n4942 vdd.n653 0.0402727
R11442 vdd.n4981 vdd.n637 0.0402727
R11443 vdd.n4990 vdd.n632 0.0402727
R11444 vdd.n5011 vdd.n602 0.0402727
R11445 vdd.n5028 vdd.n594 0.0402727
R11446 vdd.n5046 vdd.n588 0.0402727
R11447 vdd.n5064 vdd.n5063 0.0402727
R11448 vdd.n5073 vdd.n569 0.0402727
R11449 vdd.n5102 vdd.n554 0.0402727
R11450 vdd.n5124 vdd.n5123 0.0402727
R11451 vdd.n5136 vdd.n537 0.0402727
R11452 vdd.n5157 vdd.n526 0.0402727
R11453 vdd.n5170 vdd.n518 0.0402727
R11454 vdd.n5209 vdd.n502 0.0402727
R11455 vdd.n5218 vdd.n497 0.0402727
R11456 vdd.n5239 vdd.n467 0.0402727
R11457 vdd.n5256 vdd.n459 0.0402727
R11458 vdd.n5274 vdd.n453 0.0402727
R11459 vdd.n5292 vdd.n5291 0.0402727
R11460 vdd.n5301 vdd.n434 0.0402727
R11461 vdd.n5330 vdd.n419 0.0402727
R11462 vdd.n5352 vdd.n5351 0.0402727
R11463 vdd.n5364 vdd.n402 0.0402727
R11464 vdd.n5385 vdd.n391 0.0402727
R11465 vdd.n5398 vdd.n383 0.0402727
R11466 vdd.n5437 vdd.n367 0.0402727
R11467 vdd.n5446 vdd.n362 0.0402727
R11468 vdd.n5466 vdd.n341 0.0402727
R11469 vdd.n5477 vdd.n332 0.0402727
R11470 vdd.n5499 vdd.n316 0.0402727
R11471 vdd.n5529 vdd.n308 0.0402727
R11472 vdd.n5547 vdd.n302 0.0402727
R11473 vdd.n5569 vdd.n5568 0.0402727
R11474 vdd.n5719 vdd.n5718 0.0402727
R11475 vdd.n5706 vdd.n5608 0.0402727
R11476 vdd.n5641 vdd.n5611 0.0402727
R11477 vdd.n5671 vdd.n5626 0.0402727
R11478 vdd.n5681 vdd.n246 0.0402727
R11479 vdd.n5589 vdd.n5588 0.0402727
R11480 vdd.n5615 vdd.n270 0.0402727
R11481 vdd.n5704 vdd.n5703 0.0402727
R11482 vdd.n5692 vdd.n5627 0.0402727
R11483 vdd.n5674 vdd.n5651 0.0402727
R11484 vdd.n2927 vdd.n2772 0.0402727
R11485 vdd.n2940 vdd.n2764 0.0402727
R11486 vdd.n2979 vdd.n2748 0.0402727
R11487 vdd.n2988 vdd.n2743 0.0402727
R11488 vdd.n3009 vdd.n2713 0.0402727
R11489 vdd.n3026 vdd.n2705 0.0402727
R11490 vdd.n3044 vdd.n2699 0.0402727
R11491 vdd.n3062 vdd.n3061 0.0402727
R11492 vdd.n3071 vdd.n2680 0.0402727
R11493 vdd.n3100 vdd.n2665 0.0402727
R11494 vdd.n3122 vdd.n3121 0.0402727
R11495 vdd.n3134 vdd.n2648 0.0402727
R11496 vdd.n3155 vdd.n2637 0.0402727
R11497 vdd.n3168 vdd.n2629 0.0402727
R11498 vdd.n3207 vdd.n2613 0.0402727
R11499 vdd.n3216 vdd.n2608 0.0402727
R11500 vdd.n3237 vdd.n2578 0.0402727
R11501 vdd.n3254 vdd.n2570 0.0402727
R11502 vdd.n3272 vdd.n2564 0.0402727
R11503 vdd.n3290 vdd.n3289 0.0402727
R11504 vdd.n3299 vdd.n2545 0.0402727
R11505 vdd.n3328 vdd.n2530 0.0402727
R11506 vdd.n3350 vdd.n3349 0.0402727
R11507 vdd.n3362 vdd.n2513 0.0402727
R11508 vdd.n3383 vdd.n2502 0.0402727
R11509 vdd.n3396 vdd.n2494 0.0402727
R11510 vdd.n3435 vdd.n2478 0.0402727
R11511 vdd.n3444 vdd.n2473 0.0402727
R11512 vdd.n3465 vdd.n2443 0.0402727
R11513 vdd.n3482 vdd.n2435 0.0402727
R11514 vdd.n3500 vdd.n2429 0.0402727
R11515 vdd.n3518 vdd.n3517 0.0402727
R11516 vdd.n3527 vdd.n2410 0.0402727
R11517 vdd.n3556 vdd.n2395 0.0402727
R11518 vdd.n3578 vdd.n3577 0.0402727
R11519 vdd.n3590 vdd.n2378 0.0402727
R11520 vdd.n3611 vdd.n2367 0.0402727
R11521 vdd.n3624 vdd.n2359 0.0402727
R11522 vdd.n3663 vdd.n2343 0.0402727
R11523 vdd.n3672 vdd.n2338 0.0402727
R11524 vdd.n3692 vdd.n2317 0.0402727
R11525 vdd.n3702 vdd.n2307 0.0402727
R11526 vdd.n3723 vdd.n2290 0.0402727
R11527 vdd.n3753 vdd.n2282 0.0402727
R11528 vdd.n3771 vdd.n2276 0.0402727
R11529 vdd.n3793 vdd.n3792 0.0402727
R11530 vdd.n2916 vdd.n2777 0.0402727
R11531 vdd.n2946 vdd.n2765 0.0402727
R11532 vdd.n2961 vdd.n2757 0.0402727
R11533 vdd.n2977 vdd.n2976 0.0402727
R11534 vdd.n2999 vdd.n2737 0.0402727
R11535 vdd.n2729 vdd.n2712 0.0402727
R11536 vdd.n2728 vdd.n2727 0.0402727
R11537 vdd.n3029 vdd.n3028 0.0402727
R11538 vdd.n3042 vdd.n3041 0.0402727
R11539 vdd.n2691 vdd.n2677 0.0402727
R11540 vdd.n3083 vdd.n3082 0.0402727
R11541 vdd.n3098 vdd.n3097 0.0402727
R11542 vdd.n3144 vdd.n2642 0.0402727
R11543 vdd.n3174 vdd.n2630 0.0402727
R11544 vdd.n3189 vdd.n2622 0.0402727
R11545 vdd.n3205 vdd.n3204 0.0402727
R11546 vdd.n3227 vdd.n2602 0.0402727
R11547 vdd.n2594 vdd.n2577 0.0402727
R11548 vdd.n2593 vdd.n2592 0.0402727
R11549 vdd.n3257 vdd.n3256 0.0402727
R11550 vdd.n3270 vdd.n3269 0.0402727
R11551 vdd.n2556 vdd.n2542 0.0402727
R11552 vdd.n3311 vdd.n3310 0.0402727
R11553 vdd.n3326 vdd.n3325 0.0402727
R11554 vdd.n3372 vdd.n2507 0.0402727
R11555 vdd.n3402 vdd.n2495 0.0402727
R11556 vdd.n3417 vdd.n2487 0.0402727
R11557 vdd.n3433 vdd.n3432 0.0402727
R11558 vdd.n3455 vdd.n2467 0.0402727
R11559 vdd.n2459 vdd.n2442 0.0402727
R11560 vdd.n2458 vdd.n2457 0.0402727
R11561 vdd.n3485 vdd.n3484 0.0402727
R11562 vdd.n3498 vdd.n3497 0.0402727
R11563 vdd.n2421 vdd.n2407 0.0402727
R11564 vdd.n3539 vdd.n3538 0.0402727
R11565 vdd.n3554 vdd.n3553 0.0402727
R11566 vdd.n3600 vdd.n2372 0.0402727
R11567 vdd.n3630 vdd.n2360 0.0402727
R11568 vdd.n3645 vdd.n2352 0.0402727
R11569 vdd.n3661 vdd.n3660 0.0402727
R11570 vdd.n3682 vdd.n2332 0.0402727
R11571 vdd.n2324 vdd.n2316 0.0402727
R11572 vdd.n2323 vdd.n2310 0.0402727
R11573 vdd.n3712 vdd.n2301 0.0402727
R11574 vdd.n3736 vdd.n2289 0.0402727
R11575 vdd.n3756 vdd.n3755 0.0402727
R11576 vdd.n3769 vdd.n3768 0.0402727
R11577 vdd.n2267 vdd.n2266 0.0402727
R11578 vdd.n4020 vdd.n4012 0.0402727
R11579 vdd.n4030 vdd.n4029 0.0402727
R11580 vdd.n2848 vdd.n2809 0.0402727
R11581 vdd.n2857 vdd.n2804 0.0402727
R11582 vdd.n2884 vdd.n2794 0.0402727
R11583 vdd.n4018 vdd.n2049 0.0402727
R11584 vdd.n2830 vdd.n2825 0.0402727
R11585 vdd.n2846 vdd.n2845 0.0402727
R11586 vdd.n2867 vdd.n2798 0.0402727
R11587 vdd.n2793 vdd.n2788 0.0402727
R11588 vdd.n4518 vdd.n1008 0.0402727
R11589 vdd.n4513 vdd.n1012 0.0402727
R11590 vdd.n4501 vdd.n4500 0.0402727
R11591 vdd.n4491 vdd.n1076 0.0402727
R11592 vdd.n4486 vdd.n1080 0.0402727
R11593 vdd.n4475 vdd.n1116 0.0402727
R11594 vdd.n1172 vdd.n1146 0.0402727
R11595 vdd.n4453 vdd.n1166 0.0402727
R11596 vdd.n1214 vdd.n1188 0.0402727
R11597 vdd.n4431 vdd.n1208 0.0402727
R11598 vdd.n1254 vdd.n1230 0.0402727
R11599 vdd.n4406 vdd.n1255 0.0402727
R11600 vdd.n4397 vdd.n1276 0.0402727
R11601 vdd.n4392 vdd.n1280 0.0402727
R11602 vdd.n4380 vdd.n4379 0.0402727
R11603 vdd.n4370 vdd.n1340 0.0402727
R11604 vdd.n4365 vdd.n1344 0.0402727
R11605 vdd.n4354 vdd.n1380 0.0402727
R11606 vdd.n1436 vdd.n1410 0.0402727
R11607 vdd.n4332 vdd.n1430 0.0402727
R11608 vdd.n1478 vdd.n1452 0.0402727
R11609 vdd.n4310 vdd.n1472 0.0402727
R11610 vdd.n1518 vdd.n1494 0.0402727
R11611 vdd.n4285 vdd.n1519 0.0402727
R11612 vdd.n4276 vdd.n1540 0.0402727
R11613 vdd.n4271 vdd.n1544 0.0402727
R11614 vdd.n4259 vdd.n4258 0.0402727
R11615 vdd.n4249 vdd.n1604 0.0402727
R11616 vdd.n4244 vdd.n1608 0.0402727
R11617 vdd.n4233 vdd.n1644 0.0402727
R11618 vdd.n1700 vdd.n1674 0.0402727
R11619 vdd.n4211 vdd.n1694 0.0402727
R11620 vdd.n1742 vdd.n1716 0.0402727
R11621 vdd.n4189 vdd.n1736 0.0402727
R11622 vdd.n1782 vdd.n1758 0.0402727
R11623 vdd.n4164 vdd.n1783 0.0402727
R11624 vdd.n4155 vdd.n1804 0.0402727
R11625 vdd.n4150 vdd.n1808 0.0402727
R11626 vdd.n4138 vdd.n4137 0.0402727
R11627 vdd.n4128 vdd.n1868 0.0402727
R11628 vdd.n4123 vdd.n1872 0.0402727
R11629 vdd.n4112 vdd.n1908 0.0402727
R11630 vdd.n1964 vdd.n1938 0.0402727
R11631 vdd.n4090 vdd.n1958 0.0402727
R11632 vdd.n2006 vdd.n1980 0.0402727
R11633 vdd.n4068 vdd.n2000 0.0402727
R11634 vdd.n1027 vdd.n1023 0.0402727
R11635 vdd.n4516 vdd.n4515 0.0402727
R11636 vdd.n1064 vdd.n1044 0.0402727
R11637 vdd.n1096 vdd.n1092 0.0402727
R11638 vdd.n4489 vdd.n4488 0.0402727
R11639 vdd.n1135 vdd.n1134 0.0402727
R11640 vdd.n1129 vdd.n1113 0.0402727
R11641 vdd.n4464 vdd.n1147 0.0402727
R11642 vdd.n1175 vdd.n1163 0.0402727
R11643 vdd.n4442 vdd.n1189 0.0402727
R11644 vdd.n1217 vdd.n1205 0.0402727
R11645 vdd.n4420 vdd.n1231 0.0402727
R11646 vdd.n1291 vdd.n1249 0.0402727
R11647 vdd.n4395 vdd.n4394 0.0402727
R11648 vdd.n1328 vdd.n1308 0.0402727
R11649 vdd.n1360 vdd.n1356 0.0402727
R11650 vdd.n4368 vdd.n4367 0.0402727
R11651 vdd.n1399 vdd.n1398 0.0402727
R11652 vdd.n1393 vdd.n1377 0.0402727
R11653 vdd.n4343 vdd.n1411 0.0402727
R11654 vdd.n1439 vdd.n1427 0.0402727
R11655 vdd.n4321 vdd.n1453 0.0402727
R11656 vdd.n1481 vdd.n1469 0.0402727
R11657 vdd.n4299 vdd.n1495 0.0402727
R11658 vdd.n1555 vdd.n1513 0.0402727
R11659 vdd.n4274 vdd.n4273 0.0402727
R11660 vdd.n1592 vdd.n1572 0.0402727
R11661 vdd.n1624 vdd.n1620 0.0402727
R11662 vdd.n4247 vdd.n4246 0.0402727
R11663 vdd.n1663 vdd.n1662 0.0402727
R11664 vdd.n1657 vdd.n1641 0.0402727
R11665 vdd.n4222 vdd.n1675 0.0402727
R11666 vdd.n1703 vdd.n1691 0.0402727
R11667 vdd.n4200 vdd.n1717 0.0402727
R11668 vdd.n1745 vdd.n1733 0.0402727
R11669 vdd.n4178 vdd.n1759 0.0402727
R11670 vdd.n1819 vdd.n1777 0.0402727
R11671 vdd.n4153 vdd.n4152 0.0402727
R11672 vdd.n1856 vdd.n1836 0.0402727
R11673 vdd.n1888 vdd.n1884 0.0402727
R11674 vdd.n4126 vdd.n4125 0.0402727
R11675 vdd.n1927 vdd.n1926 0.0402727
R11676 vdd.n1921 vdd.n1905 0.0402727
R11677 vdd.n4101 vdd.n1939 0.0402727
R11678 vdd.n1967 vdd.n1955 0.0402727
R11679 vdd.n4079 vdd.n1981 0.0402727
R11680 vdd.n2009 vdd.n1997 0.0402727
R11681 vdd.n4057 vdd.n2023 0.0402727
R11682 vdd.n884 vdd.n854 0.0402727
R11683 vdd.n4570 vdd.n860 0.0402727
R11684 vdd.n4565 vdd.n864 0.0402727
R11685 vdd.n4553 vdd.n4552 0.0402727
R11686 vdd.n4543 vdd.n949 0.0402727
R11687 vdd.n900 vdd.n895 0.0402727
R11688 vdd.n4568 vdd.n4567 0.0402727
R11689 vdd.n937 vdd.n917 0.0402727
R11690 vdd.n969 vdd.n965 0.0402727
R11691 vdd.n4541 vdd.n4540 0.0402727
R11692 vdd.n4690 vdd.n801 0.0402727
R11693 vdd.n4720 vdd.n789 0.0402727
R11694 vdd.n4735 vdd.n781 0.0402727
R11695 vdd.n4751 vdd.n4750 0.0402727
R11696 vdd.n4773 vdd.n761 0.0402727
R11697 vdd.n753 vdd.n736 0.0402727
R11698 vdd.n752 vdd.n751 0.0402727
R11699 vdd.n4803 vdd.n4802 0.0402727
R11700 vdd.n4816 vdd.n4815 0.0402727
R11701 vdd.n715 vdd.n701 0.0402727
R11702 vdd.n4857 vdd.n4856 0.0402727
R11703 vdd.n4872 vdd.n4871 0.0402727
R11704 vdd.n4918 vdd.n666 0.0402727
R11705 vdd.n4948 vdd.n654 0.0402727
R11706 vdd.n4963 vdd.n646 0.0402727
R11707 vdd.n4979 vdd.n4978 0.0402727
R11708 vdd.n5001 vdd.n626 0.0402727
R11709 vdd.n618 vdd.n601 0.0402727
R11710 vdd.n617 vdd.n616 0.0402727
R11711 vdd.n5031 vdd.n5030 0.0402727
R11712 vdd.n5044 vdd.n5043 0.0402727
R11713 vdd.n580 vdd.n566 0.0402727
R11714 vdd.n5085 vdd.n5084 0.0402727
R11715 vdd.n5100 vdd.n5099 0.0402727
R11716 vdd.n5146 vdd.n531 0.0402727
R11717 vdd.n5176 vdd.n519 0.0402727
R11718 vdd.n5191 vdd.n511 0.0402727
R11719 vdd.n5207 vdd.n5206 0.0402727
R11720 vdd.n5229 vdd.n491 0.0402727
R11721 vdd.n483 vdd.n466 0.0402727
R11722 vdd.n482 vdd.n481 0.0402727
R11723 vdd.n5259 vdd.n5258 0.0402727
R11724 vdd.n5272 vdd.n5271 0.0402727
R11725 vdd.n445 vdd.n431 0.0402727
R11726 vdd.n5313 vdd.n5312 0.0402727
R11727 vdd.n5328 vdd.n5327 0.0402727
R11728 vdd.n5374 vdd.n396 0.0402727
R11729 vdd.n5404 vdd.n384 0.0402727
R11730 vdd.n5419 vdd.n376 0.0402727
R11731 vdd.n5435 vdd.n5434 0.0402727
R11732 vdd.n5456 vdd.n356 0.0402727
R11733 vdd.n348 vdd.n340 0.0402727
R11734 vdd.n347 vdd.n335 0.0402727
R11735 vdd.n5487 vdd.n327 0.0402727
R11736 vdd.n5512 vdd.n315 0.0402727
R11737 vdd.n5532 vdd.n5531 0.0402727
R11738 vdd.n5545 vdd.n5544 0.0402727
R11739 vdd.n293 vdd.n292 0.0402727
R11740 vdd.n7415 vdd 0.0385101
R11741 vdd.n2197 vdd.n2196 0.0383289
R11742 vdd.n2196 vdd.n2195 0.0383289
R11743 vdd.n2215 vdd.n2100 0.037359
R11744 vdd.n3985 vdd 0.0369583
R11745 vdd.n3860 vdd 0.0369583
R11746 vdd.n4627 vdd 0.0369583
R11747 vdd.n4613 vdd 0.0369583
R11748 vdd.n138 vdd.n137 0.0369583
R11749 vdd.n4789 vdd.n733 0.0368632
R11750 vdd.n5017 vdd.n598 0.0368632
R11751 vdd.n5245 vdd.n463 0.0368632
R11752 vdd.n5471 vdd.n5470 0.0368632
R11753 vdd.n6505 vdd.n6504 0.0368632
R11754 vdd.n6732 vdd.n6731 0.0368632
R11755 vdd.n6959 vdd.n6958 0.0368632
R11756 vdd.n7186 vdd.n7185 0.0368632
R11757 vdd.n6386 vdd.n6385 0.0364848
R11758 vdd.n6415 vdd.n6377 0.0364848
R11759 vdd.n6438 vdd.n6437 0.0364848
R11760 vdd.n6366 vdd.n6356 0.0364848
R11761 vdd.n6352 vdd.n6345 0.0364848
R11762 vdd.n6341 vdd.n6323 0.0364848
R11763 vdd.n6510 vdd.n6309 0.0364848
R11764 vdd.n6542 vdd.n6541 0.0364848
R11765 vdd.n6563 vdd.n6562 0.0364848
R11766 vdd.n6577 vdd.n6288 0.0364848
R11767 vdd.n6277 vdd.n6272 0.0364848
R11768 vdd.n6264 vdd.n6259 0.0364848
R11769 vdd.n6622 vdd.n6255 0.0364848
R11770 vdd.n6642 vdd.n6244 0.0364848
R11771 vdd.n6665 vdd.n6664 0.0364848
R11772 vdd.n6233 vdd.n6223 0.0364848
R11773 vdd.n6219 vdd.n6212 0.0364848
R11774 vdd.n6208 vdd.n6190 0.0364848
R11775 vdd.n6737 vdd.n6176 0.0364848
R11776 vdd.n6769 vdd.n6768 0.0364848
R11777 vdd.n6790 vdd.n6789 0.0364848
R11778 vdd.n6804 vdd.n6155 0.0364848
R11779 vdd.n6144 vdd.n6139 0.0364848
R11780 vdd.n6131 vdd.n6126 0.0364848
R11781 vdd.n6849 vdd.n6122 0.0364848
R11782 vdd.n6869 vdd.n6111 0.0364848
R11783 vdd.n6892 vdd.n6891 0.0364848
R11784 vdd.n6100 vdd.n6090 0.0364848
R11785 vdd.n6086 vdd.n6079 0.0364848
R11786 vdd.n6075 vdd.n6057 0.0364848
R11787 vdd.n6964 vdd.n6043 0.0364848
R11788 vdd.n6996 vdd.n6995 0.0364848
R11789 vdd.n7017 vdd.n7016 0.0364848
R11790 vdd.n7031 vdd.n6022 0.0364848
R11791 vdd.n6011 vdd.n6006 0.0364848
R11792 vdd.n5998 vdd.n5993 0.0364848
R11793 vdd.n7076 vdd.n5989 0.0364848
R11794 vdd.n7096 vdd.n5978 0.0364848
R11795 vdd.n7119 vdd.n7118 0.0364848
R11796 vdd.n5967 vdd.n5957 0.0364848
R11797 vdd.n5953 vdd.n5946 0.0364848
R11798 vdd.n5942 vdd.n5924 0.0364848
R11799 vdd.n7191 vdd.n5910 0.0364848
R11800 vdd.n7223 vdd.n7222 0.0364848
R11801 vdd.n7244 vdd.n7243 0.0364848
R11802 vdd.n7258 vdd.n5889 0.0364848
R11803 vdd.n5878 vdd.n5872 0.0364848
R11804 vdd.n7293 vdd.n5865 0.0364848
R11805 vdd.n7303 vdd.n5861 0.0364848
R11806 vdd.n5855 vdd.n5850 0.0364848
R11807 vdd.n5844 vdd.n5839 0.0364848
R11808 vdd.n5833 vdd.n5828 0.0364848
R11809 vdd.n5822 vdd.n5816 0.0364848
R11810 vdd.n7405 vdd.n7404 0.0364848
R11811 vdd.n5593 vdd.n5592 0.0364848
R11812 vdd.n5717 vdd.n269 0.0364848
R11813 vdd.n5708 vdd.n5707 0.0364848
R11814 vdd.n5642 vdd.n5640 0.0364848
R11815 vdd.n5672 vdd.n5628 0.0364848
R11816 vdd.n5663 vdd.n5652 0.0364848
R11817 vdd.n2904 vdd.n2782 0.0364848
R11818 vdd.n2778 vdd.n2771 0.0364848
R11819 vdd.n2942 vdd.n2766 0.0364848
R11820 vdd.n2964 vdd.n2963 0.0364848
R11821 vdd.n2752 vdd.n2742 0.0364848
R11822 vdd.n2738 vdd.n2711 0.0364848
R11823 vdd.n3025 vdd.n3024 0.0364848
R11824 vdd.n3046 vdd.n3045 0.0364848
R11825 vdd.n3060 vdd.n2690 0.0364848
R11826 vdd.n2678 vdd.n2671 0.0364848
R11827 vdd.n3102 vdd.n3101 0.0364848
R11828 vdd.n3120 vdd.n2654 0.0364848
R11829 vdd.n2655 vdd.n2647 0.0364848
R11830 vdd.n2643 vdd.n2636 0.0364848
R11831 vdd.n3170 vdd.n2631 0.0364848
R11832 vdd.n3192 vdd.n3191 0.0364848
R11833 vdd.n2617 vdd.n2607 0.0364848
R11834 vdd.n2603 vdd.n2576 0.0364848
R11835 vdd.n3253 vdd.n3252 0.0364848
R11836 vdd.n3274 vdd.n3273 0.0364848
R11837 vdd.n3288 vdd.n2555 0.0364848
R11838 vdd.n2543 vdd.n2536 0.0364848
R11839 vdd.n3330 vdd.n3329 0.0364848
R11840 vdd.n3348 vdd.n2519 0.0364848
R11841 vdd.n2520 vdd.n2512 0.0364848
R11842 vdd.n2508 vdd.n2501 0.0364848
R11843 vdd.n3398 vdd.n2496 0.0364848
R11844 vdd.n3420 vdd.n3419 0.0364848
R11845 vdd.n2482 vdd.n2472 0.0364848
R11846 vdd.n2468 vdd.n2441 0.0364848
R11847 vdd.n3481 vdd.n3480 0.0364848
R11848 vdd.n3502 vdd.n3501 0.0364848
R11849 vdd.n3516 vdd.n2420 0.0364848
R11850 vdd.n2408 vdd.n2401 0.0364848
R11851 vdd.n3558 vdd.n3557 0.0364848
R11852 vdd.n3576 vdd.n2384 0.0364848
R11853 vdd.n2385 vdd.n2377 0.0364848
R11854 vdd.n2373 vdd.n2366 0.0364848
R11855 vdd.n3626 vdd.n2361 0.0364848
R11856 vdd.n3648 vdd.n3647 0.0364848
R11857 vdd.n2347 vdd.n2337 0.0364848
R11858 vdd.n2333 vdd.n2315 0.0364848
R11859 vdd.n2311 vdd.n2306 0.0364848
R11860 vdd.n2302 vdd.n2288 0.0364848
R11861 vdd.n3752 vdd.n3751 0.0364848
R11862 vdd.n3773 vdd.n3772 0.0364848
R11863 vdd.n3791 vdd.n2265 0.0364848
R11864 vdd.n3802 vdd.n2253 0.0364848
R11865 vdd.n2043 vdd.n2040 0.0364848
R11866 vdd.n4031 vdd.n2050 0.0364848
R11867 vdd.n2833 vdd.n2832 0.0364848
R11868 vdd.n2812 vdd.n2803 0.0364848
R11869 vdd.n2799 vdd.n2792 0.0364848
R11870 vdd.n2894 vdd.n2785 0.0364848
R11871 vdd.n4528 vdd.n985 0.0364848
R11872 vdd.n1029 vdd.n1028 0.0364848
R11873 vdd.n4512 vdd.n4511 0.0364848
R11874 vdd.n4502 vdd.n1045 0.0364848
R11875 vdd.n1098 vdd.n1097 0.0364848
R11876 vdd.n4485 vdd.n4484 0.0364848
R11877 vdd.n1154 vdd.n1114 0.0364848
R11878 vdd.n1173 vdd.n1148 0.0364848
R11879 vdd.n1196 vdd.n1164 0.0364848
R11880 vdd.n1215 vdd.n1190 0.0364848
R11881 vdd.n1238 vdd.n1206 0.0364848
R11882 vdd.n1253 vdd.n1232 0.0364848
R11883 vdd.n4408 vdd.n1248 0.0364848
R11884 vdd.n1293 vdd.n1292 0.0364848
R11885 vdd.n4391 vdd.n4390 0.0364848
R11886 vdd.n4381 vdd.n1309 0.0364848
R11887 vdd.n1362 vdd.n1361 0.0364848
R11888 vdd.n4364 vdd.n4363 0.0364848
R11889 vdd.n1418 vdd.n1378 0.0364848
R11890 vdd.n1437 vdd.n1412 0.0364848
R11891 vdd.n1460 vdd.n1428 0.0364848
R11892 vdd.n1479 vdd.n1454 0.0364848
R11893 vdd.n1502 vdd.n1470 0.0364848
R11894 vdd.n1517 vdd.n1496 0.0364848
R11895 vdd.n4287 vdd.n1512 0.0364848
R11896 vdd.n1557 vdd.n1556 0.0364848
R11897 vdd.n4270 vdd.n4269 0.0364848
R11898 vdd.n4260 vdd.n1573 0.0364848
R11899 vdd.n1626 vdd.n1625 0.0364848
R11900 vdd.n4243 vdd.n4242 0.0364848
R11901 vdd.n1682 vdd.n1642 0.0364848
R11902 vdd.n1701 vdd.n1676 0.0364848
R11903 vdd.n1724 vdd.n1692 0.0364848
R11904 vdd.n1743 vdd.n1718 0.0364848
R11905 vdd.n1766 vdd.n1734 0.0364848
R11906 vdd.n1781 vdd.n1760 0.0364848
R11907 vdd.n4166 vdd.n1776 0.0364848
R11908 vdd.n1821 vdd.n1820 0.0364848
R11909 vdd.n4149 vdd.n4148 0.0364848
R11910 vdd.n4139 vdd.n1837 0.0364848
R11911 vdd.n1890 vdd.n1889 0.0364848
R11912 vdd.n4122 vdd.n4121 0.0364848
R11913 vdd.n1946 vdd.n1906 0.0364848
R11914 vdd.n1965 vdd.n1940 0.0364848
R11915 vdd.n1988 vdd.n1956 0.0364848
R11916 vdd.n2007 vdd.n1982 0.0364848
R11917 vdd.n2030 vdd.n1998 0.0364848
R11918 vdd.n4049 vdd.n2024 0.0364848
R11919 vdd.n885 vdd.n872 0.0364848
R11920 vdd.n902 vdd.n901 0.0364848
R11921 vdd.n4564 vdd.n4563 0.0364848
R11922 vdd.n4554 vdd.n918 0.0364848
R11923 vdd.n971 vdd.n970 0.0364848
R11924 vdd.n4537 vdd.n4536 0.0364848
R11925 vdd.n4678 vdd.n806 0.0364848
R11926 vdd.n802 vdd.n795 0.0364848
R11927 vdd.n4716 vdd.n790 0.0364848
R11928 vdd.n4738 vdd.n4737 0.0364848
R11929 vdd.n776 vdd.n766 0.0364848
R11930 vdd.n762 vdd.n735 0.0364848
R11931 vdd.n4799 vdd.n4798 0.0364848
R11932 vdd.n4820 vdd.n4819 0.0364848
R11933 vdd.n4834 vdd.n714 0.0364848
R11934 vdd.n702 vdd.n695 0.0364848
R11935 vdd.n4876 vdd.n4875 0.0364848
R11936 vdd.n4894 vdd.n678 0.0364848
R11937 vdd.n679 vdd.n671 0.0364848
R11938 vdd.n667 vdd.n660 0.0364848
R11939 vdd.n4944 vdd.n655 0.0364848
R11940 vdd.n4966 vdd.n4965 0.0364848
R11941 vdd.n641 vdd.n631 0.0364848
R11942 vdd.n627 vdd.n600 0.0364848
R11943 vdd.n5027 vdd.n5026 0.0364848
R11944 vdd.n5048 vdd.n5047 0.0364848
R11945 vdd.n5062 vdd.n579 0.0364848
R11946 vdd.n567 vdd.n560 0.0364848
R11947 vdd.n5104 vdd.n5103 0.0364848
R11948 vdd.n5122 vdd.n543 0.0364848
R11949 vdd.n544 vdd.n536 0.0364848
R11950 vdd.n532 vdd.n525 0.0364848
R11951 vdd.n5172 vdd.n520 0.0364848
R11952 vdd.n5194 vdd.n5193 0.0364848
R11953 vdd.n506 vdd.n496 0.0364848
R11954 vdd.n492 vdd.n465 0.0364848
R11955 vdd.n5255 vdd.n5254 0.0364848
R11956 vdd.n5276 vdd.n5275 0.0364848
R11957 vdd.n5290 vdd.n444 0.0364848
R11958 vdd.n432 vdd.n425 0.0364848
R11959 vdd.n5332 vdd.n5331 0.0364848
R11960 vdd.n5350 vdd.n408 0.0364848
R11961 vdd.n409 vdd.n401 0.0364848
R11962 vdd.n397 vdd.n390 0.0364848
R11963 vdd.n5400 vdd.n385 0.0364848
R11964 vdd.n5422 vdd.n5421 0.0364848
R11965 vdd.n371 vdd.n361 0.0364848
R11966 vdd.n357 vdd.n339 0.0364848
R11967 vdd.n5475 vdd.n331 0.0364848
R11968 vdd.n5497 vdd.n314 0.0364848
R11969 vdd.n5528 vdd.n5527 0.0364848
R11970 vdd.n5549 vdd.n5548 0.0364848
R11971 vdd.n5567 vdd.n291 0.0364848
R11972 vdd.n5578 vdd.n279 0.0364848
R11973 vdd.n4480 vdd.n1110 0.0364844
R11974 vdd.n4359 vdd.n1374 0.0364844
R11975 vdd.n4238 vdd.n1638 0.0364844
R11976 vdd.n4117 vdd.n1902 0.0364844
R11977 vdd.n3015 vdd.n2709 0.0364844
R11978 vdd.n3243 vdd.n2574 0.0364844
R11979 vdd.n3471 vdd.n2439 0.0364844
R11980 vdd.n3697 vdd.n3696 0.0364844
R11981 vdd.n146 vdd.n145 0.0361321
R11982 vdd.n7497 vdd.n201 0.0351948
R11983 vdd.n3851 vdd.n3849 0.0351948
R11984 vdd.n4595 vdd.n842 0.0351948
R11985 vdd.n7473 vdd.n7472 0.0351948
R11986 vdd.n2237 vdd.n2226 0.0350615
R11987 vdd.n3805 vdd 0.0317707
R11988 vdd.n53 vdd.n48 0.031099
R11989 vdd.n7470 vdd.n221 0.0309054
R11990 vdd.n7500 vdd.n7499 0.0309054
R11991 vdd.n3862 vdd.n3861 0.0309054
R11992 vdd.n4615 vdd.n4614 0.0309054
R11993 vdd.n6412 vdd.n6383 0.030803
R11994 vdd.n6433 vdd.n6372 0.030803
R11995 vdd.n6452 vdd.n6365 0.030803
R11996 vdd.n6473 vdd.n6350 0.030803
R11997 vdd.n6493 vdd.n6339 0.030803
R11998 vdd.n6334 vdd.n6326 0.030803
R11999 vdd.n6329 vdd.n6318 0.030803
R12000 vdd.n6524 vdd.n6312 0.030803
R12001 vdd.n6547 vdd.n6301 0.030803
R12002 vdd.n6557 vdd.n6283 0.030803
R12003 vdd.n6286 vdd.n6278 0.030803
R12004 vdd.n6600 vdd.n6265 0.030803
R12005 vdd.n6639 vdd.n6250 0.030803
R12006 vdd.n6660 vdd.n6239 0.030803
R12007 vdd.n6679 vdd.n6232 0.030803
R12008 vdd.n6700 vdd.n6217 0.030803
R12009 vdd.n6720 vdd.n6206 0.030803
R12010 vdd.n6201 vdd.n6193 0.030803
R12011 vdd.n6196 vdd.n6185 0.030803
R12012 vdd.n6751 vdd.n6179 0.030803
R12013 vdd.n6774 vdd.n6168 0.030803
R12014 vdd.n6784 vdd.n6150 0.030803
R12015 vdd.n6153 vdd.n6145 0.030803
R12016 vdd.n6827 vdd.n6132 0.030803
R12017 vdd.n6866 vdd.n6117 0.030803
R12018 vdd.n6887 vdd.n6106 0.030803
R12019 vdd.n6906 vdd.n6099 0.030803
R12020 vdd.n6927 vdd.n6084 0.030803
R12021 vdd.n6947 vdd.n6073 0.030803
R12022 vdd.n6068 vdd.n6060 0.030803
R12023 vdd.n6063 vdd.n6052 0.030803
R12024 vdd.n6978 vdd.n6046 0.030803
R12025 vdd.n7001 vdd.n6035 0.030803
R12026 vdd.n7011 vdd.n6017 0.030803
R12027 vdd.n6020 vdd.n6012 0.030803
R12028 vdd.n7054 vdd.n5999 0.030803
R12029 vdd.n7093 vdd.n5984 0.030803
R12030 vdd.n7114 vdd.n5973 0.030803
R12031 vdd.n7133 vdd.n5966 0.030803
R12032 vdd.n7154 vdd.n5951 0.030803
R12033 vdd.n7174 vdd.n5940 0.030803
R12034 vdd.n5935 vdd.n5927 0.030803
R12035 vdd.n5930 vdd.n5919 0.030803
R12036 vdd.n7205 vdd.n5913 0.030803
R12037 vdd.n7228 vdd.n5902 0.030803
R12038 vdd.n7238 vdd.n5884 0.030803
R12039 vdd.n5887 vdd.n5879 0.030803
R12040 vdd.n7286 vdd.n5866 0.030803
R12041 vdd.n7315 vdd.n5856 0.030803
R12042 vdd.n7334 vdd.n5845 0.030803
R12043 vdd.n7353 vdd.n5834 0.030803
R12044 vdd.n7372 vdd.n5823 0.030803
R12045 vdd.n7395 vdd.n5798 0.030803
R12046 vdd.n4692 vdd.n800 0.030803
R12047 vdd.n4722 vdd.n787 0.030803
R12048 vdd.n4733 vdd.n782 0.030803
R12049 vdd.n4752 vdd.n775 0.030803
R12050 vdd.n4775 vdd.n760 0.030803
R12051 vdd.n755 vdd.n738 0.030803
R12052 vdd.n750 vdd.n742 0.030803
R12053 vdd.n4804 vdd.n727 0.030803
R12054 vdd.n4814 vdd.n709 0.030803
R12055 vdd.n712 vdd.n703 0.030803
R12056 vdd.n4859 vdd.n4858 0.030803
R12057 vdd.n4870 vdd.n676 0.030803
R12058 vdd.n4920 vdd.n665 0.030803
R12059 vdd.n4950 vdd.n652 0.030803
R12060 vdd.n4961 vdd.n647 0.030803
R12061 vdd.n4980 vdd.n640 0.030803
R12062 vdd.n5003 vdd.n625 0.030803
R12063 vdd.n620 vdd.n603 0.030803
R12064 vdd.n615 vdd.n607 0.030803
R12065 vdd.n5032 vdd.n592 0.030803
R12066 vdd.n5042 vdd.n574 0.030803
R12067 vdd.n577 vdd.n568 0.030803
R12068 vdd.n5087 vdd.n5086 0.030803
R12069 vdd.n5098 vdd.n541 0.030803
R12070 vdd.n5148 vdd.n530 0.030803
R12071 vdd.n5178 vdd.n517 0.030803
R12072 vdd.n5189 vdd.n512 0.030803
R12073 vdd.n5208 vdd.n505 0.030803
R12074 vdd.n5231 vdd.n490 0.030803
R12075 vdd.n485 vdd.n468 0.030803
R12076 vdd.n480 vdd.n472 0.030803
R12077 vdd.n5260 vdd.n457 0.030803
R12078 vdd.n5270 vdd.n439 0.030803
R12079 vdd.n442 vdd.n433 0.030803
R12080 vdd.n5315 vdd.n5314 0.030803
R12081 vdd.n5326 vdd.n406 0.030803
R12082 vdd.n5376 vdd.n395 0.030803
R12083 vdd.n5406 vdd.n382 0.030803
R12084 vdd.n5417 vdd.n377 0.030803
R12085 vdd.n5436 vdd.n370 0.030803
R12086 vdd.n5458 vdd.n355 0.030803
R12087 vdd.n350 vdd.n342 0.030803
R12088 vdd.n345 vdd.n334 0.030803
R12089 vdd.n5485 vdd.n326 0.030803
R12090 vdd.n5510 vdd.n317 0.030803
R12091 vdd.n5533 vdd.n306 0.030803
R12092 vdd.n5543 vdd.n286 0.030803
R12093 vdd.n289 vdd.n280 0.030803
R12094 vdd.n5587 vdd.n266 0.030803
R12095 vdd.n5616 vdd.n5614 0.030803
R12096 vdd.n5702 vdd.n5609 0.030803
R12097 vdd.n5694 vdd.n5693 0.030803
R12098 vdd.n5676 vdd.n5664 0.030803
R12099 vdd.n2918 vdd.n2776 0.030803
R12100 vdd.n2948 vdd.n2763 0.030803
R12101 vdd.n2959 vdd.n2758 0.030803
R12102 vdd.n2978 vdd.n2751 0.030803
R12103 vdd.n3001 vdd.n2736 0.030803
R12104 vdd.n2731 vdd.n2714 0.030803
R12105 vdd.n2726 vdd.n2718 0.030803
R12106 vdd.n3030 vdd.n2703 0.030803
R12107 vdd.n3040 vdd.n2685 0.030803
R12108 vdd.n2688 vdd.n2679 0.030803
R12109 vdd.n3085 vdd.n3084 0.030803
R12110 vdd.n3096 vdd.n2652 0.030803
R12111 vdd.n3146 vdd.n2641 0.030803
R12112 vdd.n3176 vdd.n2628 0.030803
R12113 vdd.n3187 vdd.n2623 0.030803
R12114 vdd.n3206 vdd.n2616 0.030803
R12115 vdd.n3229 vdd.n2601 0.030803
R12116 vdd.n2596 vdd.n2579 0.030803
R12117 vdd.n2591 vdd.n2583 0.030803
R12118 vdd.n3258 vdd.n2568 0.030803
R12119 vdd.n3268 vdd.n2550 0.030803
R12120 vdd.n2553 vdd.n2544 0.030803
R12121 vdd.n3313 vdd.n3312 0.030803
R12122 vdd.n3324 vdd.n2517 0.030803
R12123 vdd.n3374 vdd.n2506 0.030803
R12124 vdd.n3404 vdd.n2493 0.030803
R12125 vdd.n3415 vdd.n2488 0.030803
R12126 vdd.n3434 vdd.n2481 0.030803
R12127 vdd.n3457 vdd.n2466 0.030803
R12128 vdd.n2461 vdd.n2444 0.030803
R12129 vdd.n2456 vdd.n2448 0.030803
R12130 vdd.n3486 vdd.n2433 0.030803
R12131 vdd.n3496 vdd.n2415 0.030803
R12132 vdd.n2418 vdd.n2409 0.030803
R12133 vdd.n3541 vdd.n3540 0.030803
R12134 vdd.n3552 vdd.n2382 0.030803
R12135 vdd.n3602 vdd.n2371 0.030803
R12136 vdd.n3632 vdd.n2358 0.030803
R12137 vdd.n3643 vdd.n2353 0.030803
R12138 vdd.n3662 vdd.n2346 0.030803
R12139 vdd.n3684 vdd.n2331 0.030803
R12140 vdd.n2326 vdd.n2318 0.030803
R12141 vdd.n2321 vdd.n2309 0.030803
R12142 vdd.n3710 vdd.n2300 0.030803
R12143 vdd.n3734 vdd.n2291 0.030803
R12144 vdd.n3757 vdd.n2280 0.030803
R12145 vdd.n3767 vdd.n2260 0.030803
R12146 vdd.n2263 vdd.n2254 0.030803
R12147 vdd.n4019 vdd.n4017 0.030803
R12148 vdd.n2828 vdd.n2053 0.030803
R12149 vdd.n2847 vdd.n2811 0.030803
R12150 vdd.n2869 vdd.n2797 0.030803
R12151 vdd.n2876 vdd.n2795 0.030803
R12152 vdd.n1025 vdd.n987 0.030803
R12153 vdd.n4517 vdd.n1010 0.030803
R12154 vdd.n1066 vdd.n1065 0.030803
R12155 vdd.n1094 vdd.n1048 0.030803
R12156 vdd.n4490 vdd.n1078 0.030803
R12157 vdd.n1136 vdd.n1128 0.030803
R12158 vdd.n1131 vdd.n1115 0.030803
R12159 vdd.n4466 vdd.n4465 0.030803
R12160 vdd.n1177 vdd.n1165 0.030803
R12161 vdd.n4444 vdd.n4443 0.030803
R12162 vdd.n1219 vdd.n1207 0.030803
R12163 vdd.n4422 vdd.n4421 0.030803
R12164 vdd.n1289 vdd.n1256 0.030803
R12165 vdd.n4396 vdd.n1278 0.030803
R12166 vdd.n1330 vdd.n1329 0.030803
R12167 vdd.n1358 vdd.n1312 0.030803
R12168 vdd.n4369 vdd.n1342 0.030803
R12169 vdd.n1400 vdd.n1392 0.030803
R12170 vdd.n1395 vdd.n1379 0.030803
R12171 vdd.n4345 vdd.n4344 0.030803
R12172 vdd.n1441 vdd.n1429 0.030803
R12173 vdd.n4323 vdd.n4322 0.030803
R12174 vdd.n1483 vdd.n1471 0.030803
R12175 vdd.n4301 vdd.n4300 0.030803
R12176 vdd.n1553 vdd.n1520 0.030803
R12177 vdd.n4275 vdd.n1542 0.030803
R12178 vdd.n1594 vdd.n1593 0.030803
R12179 vdd.n1622 vdd.n1576 0.030803
R12180 vdd.n4248 vdd.n1606 0.030803
R12181 vdd.n1664 vdd.n1656 0.030803
R12182 vdd.n1659 vdd.n1643 0.030803
R12183 vdd.n4224 vdd.n4223 0.030803
R12184 vdd.n1705 vdd.n1693 0.030803
R12185 vdd.n4202 vdd.n4201 0.030803
R12186 vdd.n1747 vdd.n1735 0.030803
R12187 vdd.n4180 vdd.n4179 0.030803
R12188 vdd.n1817 vdd.n1784 0.030803
R12189 vdd.n4154 vdd.n1806 0.030803
R12190 vdd.n1858 vdd.n1857 0.030803
R12191 vdd.n1886 vdd.n1840 0.030803
R12192 vdd.n4127 vdd.n1870 0.030803
R12193 vdd.n1928 vdd.n1920 0.030803
R12194 vdd.n1923 vdd.n1907 0.030803
R12195 vdd.n4103 vdd.n4102 0.030803
R12196 vdd.n1969 vdd.n1957 0.030803
R12197 vdd.n4081 vdd.n4080 0.030803
R12198 vdd.n2011 vdd.n1999 0.030803
R12199 vdd.n4059 vdd.n4058 0.030803
R12200 vdd.n898 vdd.n896 0.030803
R12201 vdd.n4569 vdd.n862 0.030803
R12202 vdd.n939 vdd.n938 0.030803
R12203 vdd.n967 vdd.n921 0.030803
R12204 vdd.n4542 vdd.n951 0.030803
R12205 vdd.n5758 vdd.n240 0.0292162
R12206 vdd.n209 vdd.n199 0.0292162
R12207 vdd.n3852 vdd.n3846 0.0292162
R12208 vdd.n4596 vdd.n4589 0.0292162
R12209 vdd.n2201 vdd.n2200 0.028087
R12210 vdd.n2104 vdd 0.0277436
R12211 vdd.n3904 vdd.n3903 0.0273994
R12212 vdd.n5583 vdd.n5582 0.026557
R12213 vdd.n7298 vdd.n7297 0.026557
R12214 vdd.n198 vdd 0.0265417
R12215 vdd.n7469 vdd 0.0265417
R12216 vdd.n2238 vdd.n2237 0.0263658
R12217 vdd.n4048 vdd.n4047 0.0263291
R12218 vdd.n4890 vdd 0.0257316
R12219 vdd.n5118 vdd 0.0257316
R12220 vdd.n5346 vdd 0.0257316
R12221 vdd vdd.n5580 0.0257316
R12222 vdd.n6618 vdd 0.0257316
R12223 vdd.n6845 vdd 0.0257316
R12224 vdd.n7072 vdd 0.0257316
R12225 vdd vdd.n7295 0.0257316
R12226 vdd.n4414 vdd 0.0254688
R12227 vdd.n4293 vdd 0.0254688
R12228 vdd.n4172 vdd 0.0254688
R12229 vdd.n4051 vdd 0.0254688
R12230 vdd.n3116 vdd 0.0254688
R12231 vdd.n3344 vdd 0.0254688
R12232 vdd.n3572 vdd 0.0254688
R12233 vdd vdd.n3804 0.0254688
R12234 vdd.n2244 vdd.n2241 0.0252507
R12235 vdd.n3824 vdd.n2077 0.0252507
R12236 vdd.n2233 vdd.n2230 0.0252507
R12237 vdd.n3832 vdd.n2071 0.0252507
R12238 vdd.n2090 vdd.n2089 0.0252507
R12239 vdd.n3818 vdd.n2082 0.0252507
R12240 vdd.n3962 vdd.n3961 0.0252507
R12241 vdd.n3956 vdd.n3955 0.0252507
R12242 vdd.n3974 vdd.n3950 0.0252507
R12243 vdd.n3925 vdd.n3915 0.0252507
R12244 vdd.n3885 vdd.n3882 0.0252507
R12245 vdd.n3878 vdd.n3877 0.0252507
R12246 vdd.n3941 vdd.n3872 0.0252507
R12247 vdd.n3933 vdd.n3930 0.0252507
R12248 vdd.n3807 vdd.n3806 0.0252507
R12249 vdd.n2087 vdd.n2084 0.0249156
R12250 vdd.n2204 vdd.n2108 0.0248273
R12251 vdd.n7458 vdd.n230 0.0242893
R12252 vdd.n237 vdd.n236 0.0242893
R12253 vdd.n5744 vdd.n5740 0.0242893
R12254 vdd.n7434 vdd.n7432 0.0242893
R12255 vdd.n7445 vdd.n5776 0.0242893
R12256 vdd.n5785 vdd.n5782 0.0242893
R12257 vdd.n7428 vdd.n5789 0.0242893
R12258 vdd.n5808 vdd.n5803 0.0242893
R12259 vdd.n4663 vdd.n811 0.0242893
R12260 vdd.n4649 vdd.n4645 0.0242893
R12261 vdd.n4655 vdd.n817 0.0242893
R12262 vdd.n4639 vdd.n4637 0.0242893
R12263 vdd.n824 vdd.n820 0.0242893
R12264 vdd.n7501 vdd.n198 0.0239375
R12265 vdd.n7469 vdd.n7468 0.0239375
R12266 vdd.n2126 vdd.n2125 0.0234759
R12267 vdd.n3897 vdd.n3896 0.0234759
R12268 vdd.n834 vdd.n833 0.0234759
R12269 vdd.n5769 vdd.n5768 0.0234759
R12270 vdd vdd.n7449 0.0234268
R12271 vdd.n7513 vdd 0.0226354
R12272 vdd.n3857 vdd.n3853 0.0226354
R12273 vdd.n4000 vdd 0.0226354
R12274 vdd.n4587 vdd.n843 0.0226354
R12275 vdd.n4608 vdd 0.0226354
R12276 vdd.n7478 vdd 0.0226354
R12277 vdd.n2041 vdd.n2039 0.0212996
R12278 vdd.n888 vdd.n874 0.0212996
R12279 vdd.n2205 vdd.n2107 0.0209327
R12280 vdd.n7530 vdd.n19 0.0206823
R12281 vdd.n7410 vdd.n7408 0.0206084
R12282 vdd.n5659 vdd.n5658 0.0206084
R12283 vdd.n6403 vdd.n6402 0.0205441
R12284 vdd.n6424 vdd.n6423 0.0205441
R12285 vdd.n6442 vdd.n6441 0.0205441
R12286 vdd.n6464 vdd.n6463 0.0205441
R12287 vdd.n6484 vdd.n6483 0.0205441
R12288 vdd.n6503 vdd.n6502 0.0205441
R12289 vdd.n6630 vdd.n6629 0.0205441
R12290 vdd.n6651 vdd.n6650 0.0205441
R12291 vdd.n6669 vdd.n6668 0.0205441
R12292 vdd.n6691 vdd.n6690 0.0205441
R12293 vdd.n6711 vdd.n6710 0.0205441
R12294 vdd.n6730 vdd.n6729 0.0205441
R12295 vdd.n6857 vdd.n6856 0.0205441
R12296 vdd.n6878 vdd.n6877 0.0205441
R12297 vdd.n6896 vdd.n6895 0.0205441
R12298 vdd.n6918 vdd.n6917 0.0205441
R12299 vdd.n6938 vdd.n6937 0.0205441
R12300 vdd.n6957 vdd.n6956 0.0205441
R12301 vdd.n7084 vdd.n7083 0.0205441
R12302 vdd.n7105 vdd.n7104 0.0205441
R12303 vdd.n7123 vdd.n7122 0.0205441
R12304 vdd.n7145 vdd.n7144 0.0205441
R12305 vdd.n7165 vdd.n7164 0.0205441
R12306 vdd.n7184 vdd.n7183 0.0205441
R12307 vdd.n4683 vdd.n4682 0.0205441
R12308 vdd.n4704 vdd.n4703 0.0205441
R12309 vdd.n4713 vdd.n4712 0.0205441
R12310 vdd.n4742 vdd.n4741 0.0205441
R12311 vdd.n4765 vdd.n4764 0.0205441
R12312 vdd.n4786 vdd.n4785 0.0205441
R12313 vdd.n4911 vdd.n4910 0.0205441
R12314 vdd.n4932 vdd.n4931 0.0205441
R12315 vdd.n4941 vdd.n4940 0.0205441
R12316 vdd.n4970 vdd.n4969 0.0205441
R12317 vdd.n4993 vdd.n4992 0.0205441
R12318 vdd.n5014 vdd.n5013 0.0205441
R12319 vdd.n5139 vdd.n5138 0.0205441
R12320 vdd.n5160 vdd.n5159 0.0205441
R12321 vdd.n5169 vdd.n5168 0.0205441
R12322 vdd.n5198 vdd.n5197 0.0205441
R12323 vdd.n5221 vdd.n5220 0.0205441
R12324 vdd.n5242 vdd.n5241 0.0205441
R12325 vdd.n5367 vdd.n5366 0.0205441
R12326 vdd.n5388 vdd.n5387 0.0205441
R12327 vdd.n5397 vdd.n5396 0.0205441
R12328 vdd.n5426 vdd.n5425 0.0205441
R12329 vdd.n5449 vdd.n5448 0.0205441
R12330 vdd.n5469 vdd.n5468 0.0205441
R12331 vdd.n2909 vdd.n2908 0.0205441
R12332 vdd.n2930 vdd.n2929 0.0205441
R12333 vdd.n2939 vdd.n2938 0.0205441
R12334 vdd.n2968 vdd.n2967 0.0205441
R12335 vdd.n2991 vdd.n2990 0.0205441
R12336 vdd.n3012 vdd.n3011 0.0205441
R12337 vdd.n3137 vdd.n3136 0.0205441
R12338 vdd.n3158 vdd.n3157 0.0205441
R12339 vdd.n3167 vdd.n3166 0.0205441
R12340 vdd.n3196 vdd.n3195 0.0205441
R12341 vdd.n3219 vdd.n3218 0.0205441
R12342 vdd.n3240 vdd.n3239 0.0205441
R12343 vdd.n3365 vdd.n3364 0.0205441
R12344 vdd.n3386 vdd.n3385 0.0205441
R12345 vdd.n3395 vdd.n3394 0.0205441
R12346 vdd.n3424 vdd.n3423 0.0205441
R12347 vdd.n3447 vdd.n3446 0.0205441
R12348 vdd.n3468 vdd.n3467 0.0205441
R12349 vdd.n3593 vdd.n3592 0.0205441
R12350 vdd.n3614 vdd.n3613 0.0205441
R12351 vdd.n3623 vdd.n3622 0.0205441
R12352 vdd.n3652 vdd.n3651 0.0205441
R12353 vdd.n3675 vdd.n3674 0.0205441
R12354 vdd.n3695 vdd.n3694 0.0205441
R12355 vdd.n4035 vdd.n2047 0.0205441
R12356 vdd.n2821 vdd.n2820 0.0205441
R12357 vdd.n2837 vdd.n2836 0.0205441
R12358 vdd.n2860 vdd.n2859 0.0205441
R12359 vdd.n2887 vdd.n2886 0.0205441
R12360 vdd.n1022 vdd.n1021 0.0205441
R12361 vdd.n1038 vdd.n1037 0.0205441
R12362 vdd.n4506 vdd.n1042 0.0205441
R12363 vdd.n1091 vdd.n1090 0.0205441
R12364 vdd.n1107 vdd.n1106 0.0205441
R12365 vdd.n4479 vdd.n1111 0.0205441
R12366 vdd.n1287 vdd.n1250 0.0205441
R12367 vdd.n1302 vdd.n1301 0.0205441
R12368 vdd.n4385 vdd.n1306 0.0205441
R12369 vdd.n1355 vdd.n1354 0.0205441
R12370 vdd.n1371 vdd.n1370 0.0205441
R12371 vdd.n4358 vdd.n1375 0.0205441
R12372 vdd.n1551 vdd.n1514 0.0205441
R12373 vdd.n1566 vdd.n1565 0.0205441
R12374 vdd.n4264 vdd.n1570 0.0205441
R12375 vdd.n1619 vdd.n1618 0.0205441
R12376 vdd.n1635 vdd.n1634 0.0205441
R12377 vdd.n4237 vdd.n1639 0.0205441
R12378 vdd.n1815 vdd.n1778 0.0205441
R12379 vdd.n1830 vdd.n1829 0.0205441
R12380 vdd.n4143 vdd.n1834 0.0205441
R12381 vdd.n1883 vdd.n1882 0.0205441
R12382 vdd.n1899 vdd.n1898 0.0205441
R12383 vdd.n4116 vdd.n1903 0.0205441
R12384 vdd.n893 vdd.n871 0.0205441
R12385 vdd.n911 vdd.n910 0.0205441
R12386 vdd.n4558 vdd.n915 0.0205441
R12387 vdd.n964 vdd.n963 0.0205441
R12388 vdd.n980 vdd.n979 0.0205441
R12389 vdd.n3828 vdd.n3827 0.0205388
R12390 vdd.n6509 vdd.n6320 0.0198529
R12391 vdd.n6531 vdd.n6530 0.0198529
R12392 vdd.n6536 vdd.n6535 0.0198529
R12393 vdd.n6569 vdd.n6568 0.0198529
R12394 vdd.n6590 vdd.n6275 0.0198529
R12395 vdd.n6614 vdd.n6262 0.0198529
R12396 vdd.n6736 vdd.n6187 0.0198529
R12397 vdd.n6758 vdd.n6757 0.0198529
R12398 vdd.n6763 vdd.n6762 0.0198529
R12399 vdd.n6796 vdd.n6795 0.0198529
R12400 vdd.n6817 vdd.n6142 0.0198529
R12401 vdd.n6841 vdd.n6129 0.0198529
R12402 vdd.n6963 vdd.n6054 0.0198529
R12403 vdd.n6985 vdd.n6984 0.0198529
R12404 vdd.n6990 vdd.n6989 0.0198529
R12405 vdd.n7023 vdd.n7022 0.0198529
R12406 vdd.n7044 vdd.n6009 0.0198529
R12407 vdd.n7068 vdd.n5996 0.0198529
R12408 vdd.n7190 vdd.n5921 0.0198529
R12409 vdd.n7212 vdd.n7211 0.0198529
R12410 vdd.n7217 vdd.n7216 0.0198529
R12411 vdd.n7250 vdd.n7249 0.0198529
R12412 vdd.n7271 vdd.n5876 0.0198529
R12413 vdd.n7275 vdd.n5874 0.0198529
R12414 vdd.n7324 vdd.n5853 0.0198529
R12415 vdd.n7343 vdd.n5842 0.0198529
R12416 vdd.n7362 vdd.n5831 0.0198529
R12417 vdd.n7381 vdd.n5820 0.0198529
R12418 vdd.n5818 vdd.n5797 0.0198529
R12419 vdd.n4788 vdd.n4787 0.0198529
R12420 vdd.n4793 vdd.n4792 0.0198529
R12421 vdd.n4826 vdd.n4825 0.0198529
R12422 vdd.n4847 vdd.n700 0.0198529
R12423 vdd.n698 vdd.n697 0.0198529
R12424 vdd.n4882 vdd.n4881 0.0198529
R12425 vdd.n5016 vdd.n5015 0.0198529
R12426 vdd.n5021 vdd.n5020 0.0198529
R12427 vdd.n5054 vdd.n5053 0.0198529
R12428 vdd.n5075 vdd.n565 0.0198529
R12429 vdd.n563 vdd.n562 0.0198529
R12430 vdd.n5110 vdd.n5109 0.0198529
R12431 vdd.n5244 vdd.n5243 0.0198529
R12432 vdd.n5249 vdd.n5248 0.0198529
R12433 vdd.n5282 vdd.n5281 0.0198529
R12434 vdd.n5303 vdd.n430 0.0198529
R12435 vdd.n428 vdd.n427 0.0198529
R12436 vdd.n5338 vdd.n5337 0.0198529
R12437 vdd.n5474 vdd.n336 0.0198529
R12438 vdd.n5496 vdd.n328 0.0198529
R12439 vdd.n5517 vdd.n5516 0.0198529
R12440 vdd.n5522 vdd.n5521 0.0198529
R12441 vdd.n5555 vdd.n5554 0.0198529
R12442 vdd.n5559 vdd.n295 0.0198529
R12443 vdd.n5599 vdd.n5598 0.0198529
R12444 vdd.n5604 vdd.n272 0.0198529
R12445 vdd.n5635 vdd.n5632 0.0198529
R12446 vdd.n5690 vdd.n5629 0.0198529
R12447 vdd.n5684 vdd.n5683 0.0198529
R12448 vdd.n3014 vdd.n3013 0.0198529
R12449 vdd.n3019 vdd.n3018 0.0198529
R12450 vdd.n3052 vdd.n3051 0.0198529
R12451 vdd.n3073 vdd.n2676 0.0198529
R12452 vdd.n2674 vdd.n2673 0.0198529
R12453 vdd.n3108 vdd.n3107 0.0198529
R12454 vdd.n3242 vdd.n3241 0.0198529
R12455 vdd.n3247 vdd.n3246 0.0198529
R12456 vdd.n3280 vdd.n3279 0.0198529
R12457 vdd.n3301 vdd.n2541 0.0198529
R12458 vdd.n2539 vdd.n2538 0.0198529
R12459 vdd.n3336 vdd.n3335 0.0198529
R12460 vdd.n3470 vdd.n3469 0.0198529
R12461 vdd.n3475 vdd.n3474 0.0198529
R12462 vdd.n3508 vdd.n3507 0.0198529
R12463 vdd.n3529 vdd.n2406 0.0198529
R12464 vdd.n2404 vdd.n2403 0.0198529
R12465 vdd.n3564 vdd.n3563 0.0198529
R12466 vdd.n3700 vdd.n2312 0.0198529
R12467 vdd.n3721 vdd.n2303 0.0198529
R12468 vdd.n3741 vdd.n3740 0.0198529
R12469 vdd.n3746 vdd.n3745 0.0198529
R12470 vdd.n3779 vdd.n3778 0.0198529
R12471 vdd.n3783 vdd.n2269 0.0198529
R12472 vdd.n4478 vdd.n4477 0.0198529
R12473 vdd.n4462 vdd.n1149 0.0198529
R12474 vdd.n4456 vdd.n4455 0.0198529
R12475 vdd.n4440 vdd.n1191 0.0198529
R12476 vdd.n4434 vdd.n4433 0.0198529
R12477 vdd.n4418 vdd.n1233 0.0198529
R12478 vdd.n4357 vdd.n4356 0.0198529
R12479 vdd.n4341 vdd.n1413 0.0198529
R12480 vdd.n4335 vdd.n4334 0.0198529
R12481 vdd.n4319 vdd.n1455 0.0198529
R12482 vdd.n4313 vdd.n4312 0.0198529
R12483 vdd.n4297 vdd.n1497 0.0198529
R12484 vdd.n4236 vdd.n4235 0.0198529
R12485 vdd.n4220 vdd.n1677 0.0198529
R12486 vdd.n4214 vdd.n4213 0.0198529
R12487 vdd.n4198 vdd.n1719 0.0198529
R12488 vdd.n4192 vdd.n4191 0.0198529
R12489 vdd.n4176 vdd.n1761 0.0198529
R12490 vdd.n4115 vdd.n4114 0.0198529
R12491 vdd.n4099 vdd.n1941 0.0198529
R12492 vdd.n4093 vdd.n4092 0.0198529
R12493 vdd.n4077 vdd.n1983 0.0198529
R12494 vdd.n4071 vdd.n4070 0.0198529
R12495 vdd.n4055 vdd.n2025 0.0198529
R12496 vdd vdd.n2100 0.0189295
R12497 vdd.n2102 vdd 0.0189295
R12498 vdd.n2205 vdd 0.0189295
R12499 vdd.n3992 vdd.n3844 0.0188117
R12500 vdd.n3993 vdd.n3992 0.0188117
R12501 vdd.n4599 vdd.n4594 0.0188117
R12502 vdd.n4600 vdd.n4599 0.0188117
R12503 vdd.n5762 vdd.n5761 0.0188117
R12504 vdd.n5761 vdd.n219 0.0188117
R12505 vdd.n6398 vdd.n6397 0.0184706
R12506 vdd.n6418 vdd.n6417 0.0184706
R12507 vdd.n6439 vdd.n6369 0.0184706
R12508 vdd.n6447 vdd.n6446 0.0184706
R12509 vdd.n6469 vdd.n6468 0.0184706
R12510 vdd.n6489 vdd.n6488 0.0184706
R12511 vdd.n6528 vdd.n6308 0.0184706
R12512 vdd.n6540 vdd.n6306 0.0184706
R12513 vdd.n6564 vdd.n6292 0.0184706
R12514 vdd.n6575 vdd.n6290 0.0184706
R12515 vdd.n6596 vdd.n6273 0.0184706
R12516 vdd.n6620 vdd.n6260 0.0184706
R12517 vdd.n6625 vdd.n6624 0.0184706
R12518 vdd.n6645 vdd.n6644 0.0184706
R12519 vdd.n6666 vdd.n6236 0.0184706
R12520 vdd.n6674 vdd.n6673 0.0184706
R12521 vdd.n6696 vdd.n6695 0.0184706
R12522 vdd.n6716 vdd.n6715 0.0184706
R12523 vdd.n6755 vdd.n6175 0.0184706
R12524 vdd.n6767 vdd.n6173 0.0184706
R12525 vdd.n6791 vdd.n6159 0.0184706
R12526 vdd.n6802 vdd.n6157 0.0184706
R12527 vdd.n6823 vdd.n6140 0.0184706
R12528 vdd.n6847 vdd.n6127 0.0184706
R12529 vdd.n6852 vdd.n6851 0.0184706
R12530 vdd.n6872 vdd.n6871 0.0184706
R12531 vdd.n6893 vdd.n6103 0.0184706
R12532 vdd.n6901 vdd.n6900 0.0184706
R12533 vdd.n6923 vdd.n6922 0.0184706
R12534 vdd.n6943 vdd.n6942 0.0184706
R12535 vdd.n6982 vdd.n6042 0.0184706
R12536 vdd.n6994 vdd.n6040 0.0184706
R12537 vdd.n7018 vdd.n6026 0.0184706
R12538 vdd.n7029 vdd.n6024 0.0184706
R12539 vdd.n7050 vdd.n6007 0.0184706
R12540 vdd.n7074 vdd.n5994 0.0184706
R12541 vdd.n7079 vdd.n7078 0.0184706
R12542 vdd.n7099 vdd.n7098 0.0184706
R12543 vdd.n7120 vdd.n5970 0.0184706
R12544 vdd.n7128 vdd.n7127 0.0184706
R12545 vdd.n7150 vdd.n7149 0.0184706
R12546 vdd.n7170 vdd.n7169 0.0184706
R12547 vdd.n7209 vdd.n5909 0.0184706
R12548 vdd.n7221 vdd.n5907 0.0184706
R12549 vdd.n7245 vdd.n5893 0.0184706
R12550 vdd.n7256 vdd.n5891 0.0184706
R12551 vdd.n7281 vdd.n5873 0.0184706
R12552 vdd.n7294 vdd.n5864 0.0184706
R12553 vdd.n7311 vdd.n5862 0.0184706
R12554 vdd.n7330 vdd.n5851 0.0184706
R12555 vdd.n7349 vdd.n5840 0.0184706
R12556 vdd.n7368 vdd.n5829 0.0184706
R12557 vdd.n7391 vdd.n5817 0.0184706
R12558 vdd.n7407 vdd.n5795 0.0184706
R12559 vdd.n4677 vdd.n4676 0.0184706
R12560 vdd.n4688 vdd.n4687 0.0184706
R12561 vdd.n4718 vdd.n4717 0.0184706
R12562 vdd.n4739 vdd.n779 0.0184706
R12563 vdd.n4747 vdd.n4746 0.0184706
R12564 vdd.n4771 vdd.n4770 0.0184706
R12565 vdd.n4797 vdd.n732 0.0184706
R12566 vdd.n4821 vdd.n718 0.0184706
R12567 vdd.n4832 vdd.n716 0.0184706
R12568 vdd.n4854 vdd.n696 0.0184706
R12569 vdd.n4877 vdd.n684 0.0184706
R12570 vdd.n4892 vdd.n681 0.0184706
R12571 vdd.n4887 vdd.n4886 0.0184706
R12572 vdd.n4916 vdd.n4915 0.0184706
R12573 vdd.n4946 vdd.n4945 0.0184706
R12574 vdd.n4967 vdd.n644 0.0184706
R12575 vdd.n4975 vdd.n4974 0.0184706
R12576 vdd.n4999 vdd.n4998 0.0184706
R12577 vdd.n5025 vdd.n597 0.0184706
R12578 vdd.n5049 vdd.n583 0.0184706
R12579 vdd.n5060 vdd.n581 0.0184706
R12580 vdd.n5082 vdd.n561 0.0184706
R12581 vdd.n5105 vdd.n549 0.0184706
R12582 vdd.n5120 vdd.n546 0.0184706
R12583 vdd.n5115 vdd.n5114 0.0184706
R12584 vdd.n5144 vdd.n5143 0.0184706
R12585 vdd.n5174 vdd.n5173 0.0184706
R12586 vdd.n5195 vdd.n509 0.0184706
R12587 vdd.n5203 vdd.n5202 0.0184706
R12588 vdd.n5227 vdd.n5226 0.0184706
R12589 vdd.n5253 vdd.n462 0.0184706
R12590 vdd.n5277 vdd.n448 0.0184706
R12591 vdd.n5288 vdd.n446 0.0184706
R12592 vdd.n5310 vdd.n426 0.0184706
R12593 vdd.n5333 vdd.n414 0.0184706
R12594 vdd.n5348 vdd.n411 0.0184706
R12595 vdd.n5343 vdd.n5342 0.0184706
R12596 vdd.n5372 vdd.n5371 0.0184706
R12597 vdd.n5402 vdd.n5401 0.0184706
R12598 vdd.n5423 vdd.n374 0.0184706
R12599 vdd.n5431 vdd.n5430 0.0184706
R12600 vdd.n5454 vdd.n5453 0.0184706
R12601 vdd.n5489 vdd.n330 0.0184706
R12602 vdd.n5514 vdd.n313 0.0184706
R12603 vdd.n5526 vdd.n311 0.0184706
R12604 vdd.n5550 vdd.n297 0.0184706
R12605 vdd.n5565 vdd.n294 0.0184706
R12606 vdd.n5579 vdd.n278 0.0184706
R12607 vdd.n5594 vdd.n274 0.0184706
R12608 vdd.n5715 vdd.n271 0.0184706
R12609 vdd.n5709 vdd.n5605 0.0184706
R12610 vdd.n5644 vdd.n5639 0.0184706
R12611 vdd.n5649 vdd.n5630 0.0184706
R12612 vdd.n5662 vdd.n5654 0.0184706
R12613 vdd.n2903 vdd.n2902 0.0184706
R12614 vdd.n2914 vdd.n2913 0.0184706
R12615 vdd.n2944 vdd.n2943 0.0184706
R12616 vdd.n2965 vdd.n2755 0.0184706
R12617 vdd.n2973 vdd.n2972 0.0184706
R12618 vdd.n2997 vdd.n2996 0.0184706
R12619 vdd.n3023 vdd.n2708 0.0184706
R12620 vdd.n3047 vdd.n2694 0.0184706
R12621 vdd.n3058 vdd.n2692 0.0184706
R12622 vdd.n3080 vdd.n2672 0.0184706
R12623 vdd.n3103 vdd.n2660 0.0184706
R12624 vdd.n3118 vdd.n2657 0.0184706
R12625 vdd.n3113 vdd.n3112 0.0184706
R12626 vdd.n3142 vdd.n3141 0.0184706
R12627 vdd.n3172 vdd.n3171 0.0184706
R12628 vdd.n3193 vdd.n2620 0.0184706
R12629 vdd.n3201 vdd.n3200 0.0184706
R12630 vdd.n3225 vdd.n3224 0.0184706
R12631 vdd.n3251 vdd.n2573 0.0184706
R12632 vdd.n3275 vdd.n2559 0.0184706
R12633 vdd.n3286 vdd.n2557 0.0184706
R12634 vdd.n3308 vdd.n2537 0.0184706
R12635 vdd.n3331 vdd.n2525 0.0184706
R12636 vdd.n3346 vdd.n2522 0.0184706
R12637 vdd.n3341 vdd.n3340 0.0184706
R12638 vdd.n3370 vdd.n3369 0.0184706
R12639 vdd.n3400 vdd.n3399 0.0184706
R12640 vdd.n3421 vdd.n2485 0.0184706
R12641 vdd.n3429 vdd.n3428 0.0184706
R12642 vdd.n3453 vdd.n3452 0.0184706
R12643 vdd.n3479 vdd.n2438 0.0184706
R12644 vdd.n3503 vdd.n2424 0.0184706
R12645 vdd.n3514 vdd.n2422 0.0184706
R12646 vdd.n3536 vdd.n2402 0.0184706
R12647 vdd.n3559 vdd.n2390 0.0184706
R12648 vdd.n3574 vdd.n2387 0.0184706
R12649 vdd.n3569 vdd.n3568 0.0184706
R12650 vdd.n3598 vdd.n3597 0.0184706
R12651 vdd.n3628 vdd.n3627 0.0184706
R12652 vdd.n3649 vdd.n2350 0.0184706
R12653 vdd.n3657 vdd.n3656 0.0184706
R12654 vdd.n3680 vdd.n3679 0.0184706
R12655 vdd.n3714 vdd.n2305 0.0184706
R12656 vdd.n3738 vdd.n2287 0.0184706
R12657 vdd.n3750 vdd.n2285 0.0184706
R12658 vdd.n3774 vdd.n2271 0.0184706
R12659 vdd.n3789 vdd.n2268 0.0184706
R12660 vdd.n3803 vdd.n2252 0.0184706
R12661 vdd.n4040 vdd.n4039 0.0184706
R12662 vdd.n4033 vdd.n2048 0.0184706
R12663 vdd.n2834 vdd.n2815 0.0184706
R12664 vdd.n2842 vdd.n2841 0.0184706
R12665 vdd.n2865 vdd.n2864 0.0184706
R12666 vdd.n2892 vdd.n2891 0.0184706
R12667 vdd.n4529 vdd.n984 0.0184706
R12668 vdd.n1031 vdd.n1017 0.0184706
R12669 vdd.n4510 vdd.n1014 0.0184706
R12670 vdd.n4504 vdd.n1043 0.0184706
R12671 vdd.n1100 vdd.n1085 0.0184706
R12672 vdd.n4483 vdd.n1082 0.0184706
R12673 vdd.n1156 vdd.n1153 0.0184706
R12674 vdd.n1161 vdd.n1150 0.0184706
R12675 vdd.n1198 vdd.n1195 0.0184706
R12676 vdd.n1203 vdd.n1192 0.0184706
R12677 vdd.n1240 vdd.n1237 0.0184706
R12678 vdd.n1244 vdd.n1234 0.0184706
R12679 vdd.n4409 vdd.n1245 0.0184706
R12680 vdd.n1295 vdd.n1285 0.0184706
R12681 vdd.n4389 vdd.n1282 0.0184706
R12682 vdd.n4383 vdd.n1307 0.0184706
R12683 vdd.n1364 vdd.n1349 0.0184706
R12684 vdd.n4362 vdd.n1346 0.0184706
R12685 vdd.n1420 vdd.n1417 0.0184706
R12686 vdd.n1425 vdd.n1414 0.0184706
R12687 vdd.n1462 vdd.n1459 0.0184706
R12688 vdd.n1467 vdd.n1456 0.0184706
R12689 vdd.n1504 vdd.n1501 0.0184706
R12690 vdd.n1508 vdd.n1498 0.0184706
R12691 vdd.n4288 vdd.n1509 0.0184706
R12692 vdd.n1559 vdd.n1549 0.0184706
R12693 vdd.n4268 vdd.n1546 0.0184706
R12694 vdd.n4262 vdd.n1571 0.0184706
R12695 vdd.n1628 vdd.n1613 0.0184706
R12696 vdd.n4241 vdd.n1610 0.0184706
R12697 vdd.n1684 vdd.n1681 0.0184706
R12698 vdd.n1689 vdd.n1678 0.0184706
R12699 vdd.n1726 vdd.n1723 0.0184706
R12700 vdd.n1731 vdd.n1720 0.0184706
R12701 vdd.n1768 vdd.n1765 0.0184706
R12702 vdd.n1772 vdd.n1762 0.0184706
R12703 vdd.n4167 vdd.n1773 0.0184706
R12704 vdd.n1823 vdd.n1813 0.0184706
R12705 vdd.n4147 vdd.n1810 0.0184706
R12706 vdd.n4141 vdd.n1835 0.0184706
R12707 vdd.n1892 vdd.n1877 0.0184706
R12708 vdd.n4120 vdd.n1874 0.0184706
R12709 vdd.n1948 vdd.n1945 0.0184706
R12710 vdd.n1953 vdd.n1942 0.0184706
R12711 vdd.n1990 vdd.n1987 0.0184706
R12712 vdd.n1995 vdd.n1984 0.0184706
R12713 vdd.n2032 vdd.n2029 0.0184706
R12714 vdd.n4050 vdd.n2026 0.0184706
R12715 vdd.n887 vdd.n873 0.0184706
R12716 vdd.n904 vdd.n869 0.0184706
R12717 vdd.n4562 vdd.n866 0.0184706
R12718 vdd.n4556 vdd.n916 0.0184706
R12719 vdd.n973 vdd.n958 0.0184706
R12720 vdd.n4535 vdd.n955 0.0184706
R12721 vdd.n2229 vdd.n2073 0.0181705
R12722 vdd.n3813 vdd.n3812 0.0177558
R12723 vdd.n3863 vdd.n3859 0.0174271
R12724 vdd.n4616 vdd.n4588 0.0174271
R12725 vdd.n187 vdd.n186 0.017313
R12726 vdd.n837 vdd.n828 0.0172857
R12727 vdd.n5772 vdd.n5763 0.0172857
R12728 vdd.n2246 vdd.n2076 0.0172597
R12729 vdd.n3910 vdd.n3909 0.0167579
R12730 vdd.n7487 vdd.n197 0.016125
R12731 vdd.n5756 vdd.n222 0.016125
R12732 vdd.n2133 vdd.n2132 0.0159756
R12733 vdd.n2157 vdd.n2112 0.0159756
R12734 vdd.n2188 vdd.n2185 0.0159756
R12735 vdd vdd.n4048 0.0159219
R12736 vdd.n5581 vdd 0.0158368
R12737 vdd.n7296 vdd 0.0158368
R12738 vdd.n3966 vdd.n3965 0.0157919
R12739 vdd vdd.n2204 0.0157244
R12740 vdd.n6393 vdd.n6389 0.0156071
R12741 vdd.n7457 vdd.n232 0.0156071
R12742 vdd.n7457 vdd.n231 0.0156071
R12743 vdd.n7455 vdd.n235 0.0156071
R12744 vdd.n7455 vdd.n7454 0.0156071
R12745 vdd.n5745 vdd.n5739 0.0156071
R12746 vdd.n5741 vdd.n5739 0.0156071
R12747 vdd.n7433 vdd.n7431 0.0156071
R12748 vdd.n7439 vdd.n7431 0.0156071
R12749 vdd.n7446 vdd.n5775 0.0156071
R12750 vdd.n7442 vdd.n5775 0.0156071
R12751 vdd.n5786 vdd.n5773 0.0156071
R12752 vdd.n5786 vdd.n5779 0.0156071
R12753 vdd.n7429 vdd.n5788 0.0156071
R12754 vdd.n7429 vdd.n5780 0.0156071
R12755 vdd.n5807 vdd.n5806 0.0156071
R12756 vdd.n5807 vdd.n5804 0.0156071
R12757 vdd.n4662 vdd.n810 0.0156071
R12758 vdd.n4666 vdd.n810 0.0156071
R12759 vdd.n4671 vdd.n808 0.0156071
R12760 vdd.n4648 vdd.n4647 0.0156071
R12761 vdd.n4648 vdd.n4646 0.0156071
R12762 vdd.n4659 vdd.n816 0.0156071
R12763 vdd.n4659 vdd.n4658 0.0156071
R12764 vdd.n4636 vdd.n815 0.0156071
R12765 vdd.n4638 vdd.n815 0.0156071
R12766 vdd.n823 vdd.n822 0.0156071
R12767 vdd.n823 vdd.n821 0.0156071
R12768 vdd.n2247 vdd.n2245 0.0156071
R12769 vdd.n3826 vdd.n3825 0.0156071
R12770 vdd.n2225 vdd.n2224 0.0156071
R12771 vdd.n2235 vdd.n2234 0.0156071
R12772 vdd.n3831 vdd.n2072 0.0156071
R12773 vdd.n2092 vdd.n2091 0.0156071
R12774 vdd.n3817 vdd.n2083 0.0156071
R12775 vdd.n3964 vdd.n3963 0.0156071
R12776 vdd.n3967 vdd.n3957 0.0156071
R12777 vdd.n3973 vdd.n3951 0.0156071
R12778 vdd.n3927 vdd.n3926 0.0156071
R12779 vdd.n3902 vdd.n3890 0.0156071
R12780 vdd.n3905 vdd.n3886 0.0156071
R12781 vdd.n3908 vdd.n3879 0.0156071
R12782 vdd.n3940 vdd.n3873 0.0156071
R12783 vdd.n3935 vdd.n3934 0.0156071
R12784 vdd.n3810 vdd.n2249 0.0156071
R12785 vdd.n2250 vdd.n2249 0.0156071
R12786 vdd.n2161 vdd.n2160 0.0154024
R12787 vdd.n2096 vdd.n2094 0.0154024
R12788 vdd.n2131 vdd.n2119 0.0154024
R12789 vdd.n2151 vdd.n2113 0.0154024
R12790 vdd.n2199 vdd.n2165 0.0154024
R12791 vdd.n2117 vdd.n2116 0.0154024
R12792 vdd.n2 vdd.n1 0.0154024
R12793 vdd.n142 vdd.n128 0.0154024
R12794 vdd.n80 vdd.n79 0.0154024
R12795 vdd.n95 vdd.n94 0.0154024
R12796 vdd.n66 vdd.n65 0.0154024
R12797 vdd.n183 vdd.n147 0.0154024
R12798 vdd.n7526 vdd.n21 0.0154024
R12799 vdd.n7409 vdd.n5793 0.0152558
R12800 vdd.n5657 vdd.n244 0.0152558
R12801 vdd.n4044 vdd.n4043 0.0152558
R12802 vdd.n880 vdd.n877 0.0152558
R12803 vdd.n2127 vdd.n2124 0.0148621
R12804 vdd.n3898 vdd.n3895 0.0148621
R12805 vdd.n835 vdd.n832 0.0148621
R12806 vdd.n5770 vdd.n5767 0.0148621
R12807 vdd.n3907 vdd.n3906 0.0148365
R12808 vdd.n6402 vdd.n6381 0.0143235
R12809 vdd.n6423 vdd.n6379 0.0143235
R12810 vdd.n6442 vdd.n6367 0.0143235
R12811 vdd.n6464 vdd.n6353 0.0143235
R12812 vdd.n6484 vdd.n6342 0.0143235
R12813 vdd.n6531 vdd.n6529 0.0143235
R12814 vdd.n6537 vdd.n6536 0.0143235
R12815 vdd.n6568 vdd.n6567 0.0143235
R12816 vdd.n6574 vdd.n6275 0.0143235
R12817 vdd.n6595 vdd.n6262 0.0143235
R12818 vdd.n6629 vdd.n6248 0.0143235
R12819 vdd.n6650 vdd.n6246 0.0143235
R12820 vdd.n6669 vdd.n6234 0.0143235
R12821 vdd.n6691 vdd.n6220 0.0143235
R12822 vdd.n6711 vdd.n6209 0.0143235
R12823 vdd.n6758 vdd.n6756 0.0143235
R12824 vdd.n6764 vdd.n6763 0.0143235
R12825 vdd.n6795 vdd.n6794 0.0143235
R12826 vdd.n6801 vdd.n6142 0.0143235
R12827 vdd.n6822 vdd.n6129 0.0143235
R12828 vdd.n6856 vdd.n6115 0.0143235
R12829 vdd.n6877 vdd.n6113 0.0143235
R12830 vdd.n6896 vdd.n6101 0.0143235
R12831 vdd.n6918 vdd.n6087 0.0143235
R12832 vdd.n6938 vdd.n6076 0.0143235
R12833 vdd.n6985 vdd.n6983 0.0143235
R12834 vdd.n6991 vdd.n6990 0.0143235
R12835 vdd.n7022 vdd.n7021 0.0143235
R12836 vdd.n7028 vdd.n6009 0.0143235
R12837 vdd.n7049 vdd.n5996 0.0143235
R12838 vdd.n7083 vdd.n5982 0.0143235
R12839 vdd.n7104 vdd.n5980 0.0143235
R12840 vdd.n7123 vdd.n5968 0.0143235
R12841 vdd.n7145 vdd.n5954 0.0143235
R12842 vdd.n7165 vdd.n5943 0.0143235
R12843 vdd.n7212 vdd.n7210 0.0143235
R12844 vdd.n7218 vdd.n7217 0.0143235
R12845 vdd.n7249 vdd.n7248 0.0143235
R12846 vdd.n7255 vdd.n5876 0.0143235
R12847 vdd.n7280 vdd.n5874 0.0143235
R12848 vdd.n7310 vdd.n5853 0.0143235
R12849 vdd.n7329 vdd.n5842 0.0143235
R12850 vdd.n7348 vdd.n5831 0.0143235
R12851 vdd.n7367 vdd.n5820 0.0143235
R12852 vdd.n7390 vdd.n5818 0.0143235
R12853 vdd.n4683 vdd.n803 0.0143235
R12854 vdd.n4704 vdd.n791 0.0143235
R12855 vdd.n4712 vdd.n4708 0.0143235
R12856 vdd.n4742 vdd.n777 0.0143235
R12857 vdd.n4765 vdd.n763 0.0143235
R12858 vdd.n4794 vdd.n4793 0.0143235
R12859 vdd.n4825 vdd.n4824 0.0143235
R12860 vdd.n4831 vdd.n700 0.0143235
R12861 vdd.n4853 vdd.n698 0.0143235
R12862 vdd.n4881 vdd.n4880 0.0143235
R12863 vdd.n4911 vdd.n668 0.0143235
R12864 vdd.n4932 vdd.n656 0.0143235
R12865 vdd.n4940 vdd.n4936 0.0143235
R12866 vdd.n4970 vdd.n642 0.0143235
R12867 vdd.n4993 vdd.n628 0.0143235
R12868 vdd.n5022 vdd.n5021 0.0143235
R12869 vdd.n5053 vdd.n5052 0.0143235
R12870 vdd.n5059 vdd.n565 0.0143235
R12871 vdd.n5081 vdd.n563 0.0143235
R12872 vdd.n5109 vdd.n5108 0.0143235
R12873 vdd.n5139 vdd.n533 0.0143235
R12874 vdd.n5160 vdd.n521 0.0143235
R12875 vdd.n5168 vdd.n5164 0.0143235
R12876 vdd.n5198 vdd.n507 0.0143235
R12877 vdd.n5221 vdd.n493 0.0143235
R12878 vdd.n5250 vdd.n5249 0.0143235
R12879 vdd.n5281 vdd.n5280 0.0143235
R12880 vdd.n5287 vdd.n430 0.0143235
R12881 vdd.n5309 vdd.n428 0.0143235
R12882 vdd.n5337 vdd.n5336 0.0143235
R12883 vdd.n5367 vdd.n398 0.0143235
R12884 vdd.n5388 vdd.n386 0.0143235
R12885 vdd.n5396 vdd.n5392 0.0143235
R12886 vdd.n5426 vdd.n372 0.0143235
R12887 vdd.n5449 vdd.n358 0.0143235
R12888 vdd.n5490 vdd.n328 0.0143235
R12889 vdd.n5517 vdd.n5515 0.0143235
R12890 vdd.n5523 vdd.n5522 0.0143235
R12891 vdd.n5554 vdd.n5553 0.0143235
R12892 vdd.n5564 vdd.n295 0.0143235
R12893 vdd.n5598 vdd.n5597 0.0143235
R12894 vdd.n5714 vdd.n272 0.0143235
R12895 vdd.n5635 vdd.n5634 0.0143235
R12896 vdd.n5645 vdd.n5629 0.0143235
R12897 vdd.n5685 vdd.n5684 0.0143235
R12898 vdd.n2909 vdd.n2779 0.0143235
R12899 vdd.n2930 vdd.n2767 0.0143235
R12900 vdd.n2938 vdd.n2934 0.0143235
R12901 vdd.n2968 vdd.n2753 0.0143235
R12902 vdd.n2991 vdd.n2739 0.0143235
R12903 vdd.n3020 vdd.n3019 0.0143235
R12904 vdd.n3051 vdd.n3050 0.0143235
R12905 vdd.n3057 vdd.n2676 0.0143235
R12906 vdd.n3079 vdd.n2674 0.0143235
R12907 vdd.n3107 vdd.n3106 0.0143235
R12908 vdd.n3137 vdd.n2644 0.0143235
R12909 vdd.n3158 vdd.n2632 0.0143235
R12910 vdd.n3166 vdd.n3162 0.0143235
R12911 vdd.n3196 vdd.n2618 0.0143235
R12912 vdd.n3219 vdd.n2604 0.0143235
R12913 vdd.n3248 vdd.n3247 0.0143235
R12914 vdd.n3279 vdd.n3278 0.0143235
R12915 vdd.n3285 vdd.n2541 0.0143235
R12916 vdd.n3307 vdd.n2539 0.0143235
R12917 vdd.n3335 vdd.n3334 0.0143235
R12918 vdd.n3365 vdd.n2509 0.0143235
R12919 vdd.n3386 vdd.n2497 0.0143235
R12920 vdd.n3394 vdd.n3390 0.0143235
R12921 vdd.n3424 vdd.n2483 0.0143235
R12922 vdd.n3447 vdd.n2469 0.0143235
R12923 vdd.n3476 vdd.n3475 0.0143235
R12924 vdd.n3507 vdd.n3506 0.0143235
R12925 vdd.n3513 vdd.n2406 0.0143235
R12926 vdd.n3535 vdd.n2404 0.0143235
R12927 vdd.n3563 vdd.n3562 0.0143235
R12928 vdd.n3593 vdd.n2374 0.0143235
R12929 vdd.n3614 vdd.n2362 0.0143235
R12930 vdd.n3622 vdd.n3618 0.0143235
R12931 vdd.n3652 vdd.n2348 0.0143235
R12932 vdd.n3675 vdd.n2334 0.0143235
R12933 vdd.n3715 vdd.n2303 0.0143235
R12934 vdd.n3741 vdd.n3739 0.0143235
R12935 vdd.n3747 vdd.n3746 0.0143235
R12936 vdd.n3778 vdd.n3777 0.0143235
R12937 vdd.n3788 vdd.n2269 0.0143235
R12938 vdd.n4035 vdd.n4034 0.0143235
R12939 vdd.n2822 vdd.n2821 0.0143235
R12940 vdd.n2837 vdd.n2813 0.0143235
R12941 vdd.n2860 vdd.n2800 0.0143235
R12942 vdd.n2887 vdd.n2789 0.0143235
R12943 vdd.n1032 vdd.n1022 0.0143235
R12944 vdd.n1039 vdd.n1038 0.0143235
R12945 vdd.n4506 vdd.n4505 0.0143235
R12946 vdd.n1101 vdd.n1091 0.0143235
R12947 vdd.n1108 vdd.n1107 0.0143235
R12948 vdd.n1157 vdd.n1149 0.0143235
R12949 vdd.n4457 vdd.n4456 0.0143235
R12950 vdd.n1199 vdd.n1191 0.0143235
R12951 vdd.n4435 vdd.n4434 0.0143235
R12952 vdd.n1241 vdd.n1233 0.0143235
R12953 vdd.n1296 vdd.n1287 0.0143235
R12954 vdd.n1303 vdd.n1302 0.0143235
R12955 vdd.n4385 vdd.n4384 0.0143235
R12956 vdd.n1365 vdd.n1355 0.0143235
R12957 vdd.n1372 vdd.n1371 0.0143235
R12958 vdd.n1421 vdd.n1413 0.0143235
R12959 vdd.n4336 vdd.n4335 0.0143235
R12960 vdd.n1463 vdd.n1455 0.0143235
R12961 vdd.n4314 vdd.n4313 0.0143235
R12962 vdd.n1505 vdd.n1497 0.0143235
R12963 vdd.n1560 vdd.n1551 0.0143235
R12964 vdd.n1567 vdd.n1566 0.0143235
R12965 vdd.n4264 vdd.n4263 0.0143235
R12966 vdd.n1629 vdd.n1619 0.0143235
R12967 vdd.n1636 vdd.n1635 0.0143235
R12968 vdd.n1685 vdd.n1677 0.0143235
R12969 vdd.n4215 vdd.n4214 0.0143235
R12970 vdd.n1727 vdd.n1719 0.0143235
R12971 vdd.n4193 vdd.n4192 0.0143235
R12972 vdd.n1769 vdd.n1761 0.0143235
R12973 vdd.n1824 vdd.n1815 0.0143235
R12974 vdd.n1831 vdd.n1830 0.0143235
R12975 vdd.n4143 vdd.n4142 0.0143235
R12976 vdd.n1893 vdd.n1883 0.0143235
R12977 vdd.n1900 vdd.n1899 0.0143235
R12978 vdd.n1949 vdd.n1941 0.0143235
R12979 vdd.n4094 vdd.n4093 0.0143235
R12980 vdd.n1991 vdd.n1983 0.0143235
R12981 vdd.n4072 vdd.n4071 0.0143235
R12982 vdd.n2033 vdd.n2025 0.0143235
R12983 vdd.n905 vdd.n871 0.0143235
R12984 vdd.n912 vdd.n911 0.0143235
R12985 vdd.n4558 vdd.n4557 0.0143235
R12986 vdd.n974 vdd.n964 0.0143235
R12987 vdd.n981 vdd.n980 0.0143235
R12988 vdd.n2216 vdd.n2215 0.0141218
R12989 vdd.n3937 vdd.n3936 0.0140975
R12990 vdd.n240 vdd.n221 0.0140135
R12991 vdd.n7500 vdd.n199 0.0140135
R12992 vdd.n3862 vdd.n3846 0.0140135
R12993 vdd.n4615 vdd.n4589 0.0140135
R12994 vdd.n127 vdd.n126 0.0139695
R12995 vdd.n7523 vdd.n7522 0.013874
R12996 vdd.n6416 vdd.n6415 0.0137576
R12997 vdd.n6437 vdd.n6436 0.0137576
R12998 vdd.n6448 vdd.n6366 0.0137576
R12999 vdd.n6470 vdd.n6352 0.0137576
R13000 vdd.n6490 vdd.n6341 0.0137576
R13001 vdd.n6527 vdd.n6309 0.0137576
R13002 vdd.n6542 vdd.n6302 0.0137576
R13003 vdd.n6562 vdd.n6296 0.0137576
R13004 vdd.n6577 vdd.n6576 0.0137576
R13005 vdd.n6597 vdd.n6272 0.0137576
R13006 vdd.n6621 vdd.n6259 0.0137576
R13007 vdd.n6623 vdd.n6622 0.0137576
R13008 vdd.n6643 vdd.n6642 0.0137576
R13009 vdd.n6664 vdd.n6663 0.0137576
R13010 vdd.n6675 vdd.n6233 0.0137576
R13011 vdd.n6697 vdd.n6219 0.0137576
R13012 vdd.n6717 vdd.n6208 0.0137576
R13013 vdd.n6754 vdd.n6176 0.0137576
R13014 vdd.n6769 vdd.n6169 0.0137576
R13015 vdd.n6789 vdd.n6163 0.0137576
R13016 vdd.n6804 vdd.n6803 0.0137576
R13017 vdd.n6824 vdd.n6139 0.0137576
R13018 vdd.n6848 vdd.n6126 0.0137576
R13019 vdd.n6850 vdd.n6849 0.0137576
R13020 vdd.n6870 vdd.n6869 0.0137576
R13021 vdd.n6891 vdd.n6890 0.0137576
R13022 vdd.n6902 vdd.n6100 0.0137576
R13023 vdd.n6924 vdd.n6086 0.0137576
R13024 vdd.n6944 vdd.n6075 0.0137576
R13025 vdd.n6981 vdd.n6043 0.0137576
R13026 vdd.n6996 vdd.n6036 0.0137576
R13027 vdd.n7016 vdd.n6030 0.0137576
R13028 vdd.n7031 vdd.n7030 0.0137576
R13029 vdd.n7051 vdd.n6006 0.0137576
R13030 vdd.n7075 vdd.n5993 0.0137576
R13031 vdd.n7077 vdd.n7076 0.0137576
R13032 vdd.n7097 vdd.n7096 0.0137576
R13033 vdd.n7118 vdd.n7117 0.0137576
R13034 vdd.n7129 vdd.n5967 0.0137576
R13035 vdd.n7151 vdd.n5953 0.0137576
R13036 vdd.n7171 vdd.n5942 0.0137576
R13037 vdd.n7208 vdd.n5910 0.0137576
R13038 vdd.n7223 vdd.n5903 0.0137576
R13039 vdd.n7243 vdd.n5897 0.0137576
R13040 vdd.n7258 vdd.n7257 0.0137576
R13041 vdd.n7282 vdd.n5872 0.0137576
R13042 vdd.n7312 vdd.n5861 0.0137576
R13043 vdd.n7331 vdd.n5850 0.0137576
R13044 vdd.n7350 vdd.n5839 0.0137576
R13045 vdd.n7369 vdd.n5828 0.0137576
R13046 vdd.n7392 vdd.n5816 0.0137576
R13047 vdd.n7406 vdd.n7405 0.0137576
R13048 vdd.n5592 vdd.n5586 0.0137576
R13049 vdd.n5717 vdd.n5716 0.0137576
R13050 vdd.n5707 vdd.n5607 0.0137576
R13051 vdd.n5643 vdd.n5642 0.0137576
R13052 vdd.n5673 vdd.n5672 0.0137576
R13053 vdd.n5653 vdd.n5652 0.0137576
R13054 vdd.n2915 vdd.n2778 0.0137576
R13055 vdd.n2945 vdd.n2766 0.0137576
R13056 vdd.n2963 vdd.n2962 0.0137576
R13057 vdd.n2974 vdd.n2752 0.0137576
R13058 vdd.n2998 vdd.n2738 0.0137576
R13059 vdd.n3025 vdd.n2704 0.0137576
R13060 vdd.n3045 vdd.n2698 0.0137576
R13061 vdd.n3060 vdd.n3059 0.0137576
R13062 vdd.n3081 vdd.n2671 0.0137576
R13063 vdd.n3101 vdd.n2664 0.0137576
R13064 vdd.n3120 vdd.n3119 0.0137576
R13065 vdd.n2656 vdd.n2655 0.0137576
R13066 vdd.n3143 vdd.n2643 0.0137576
R13067 vdd.n3173 vdd.n2631 0.0137576
R13068 vdd.n3191 vdd.n3190 0.0137576
R13069 vdd.n3202 vdd.n2617 0.0137576
R13070 vdd.n3226 vdd.n2603 0.0137576
R13071 vdd.n3253 vdd.n2569 0.0137576
R13072 vdd.n3273 vdd.n2563 0.0137576
R13073 vdd.n3288 vdd.n3287 0.0137576
R13074 vdd.n3309 vdd.n2536 0.0137576
R13075 vdd.n3329 vdd.n2529 0.0137576
R13076 vdd.n3348 vdd.n3347 0.0137576
R13077 vdd.n2521 vdd.n2520 0.0137576
R13078 vdd.n3371 vdd.n2508 0.0137576
R13079 vdd.n3401 vdd.n2496 0.0137576
R13080 vdd.n3419 vdd.n3418 0.0137576
R13081 vdd.n3430 vdd.n2482 0.0137576
R13082 vdd.n3454 vdd.n2468 0.0137576
R13083 vdd.n3481 vdd.n2434 0.0137576
R13084 vdd.n3501 vdd.n2428 0.0137576
R13085 vdd.n3516 vdd.n3515 0.0137576
R13086 vdd.n3537 vdd.n2401 0.0137576
R13087 vdd.n3557 vdd.n2394 0.0137576
R13088 vdd.n3576 vdd.n3575 0.0137576
R13089 vdd.n2386 vdd.n2385 0.0137576
R13090 vdd.n3599 vdd.n2373 0.0137576
R13091 vdd.n3629 vdd.n2361 0.0137576
R13092 vdd.n3647 vdd.n3646 0.0137576
R13093 vdd.n3658 vdd.n2347 0.0137576
R13094 vdd.n3681 vdd.n2333 0.0137576
R13095 vdd.n3713 vdd.n2306 0.0137576
R13096 vdd.n3737 vdd.n2288 0.0137576
R13097 vdd.n3752 vdd.n2281 0.0137576
R13098 vdd.n3772 vdd.n2275 0.0137576
R13099 vdd.n3791 vdd.n3790 0.0137576
R13100 vdd.n4041 vdd.n2040 0.0137576
R13101 vdd.n4032 vdd.n4031 0.0137576
R13102 vdd.n2832 vdd.n2831 0.0137576
R13103 vdd.n2843 vdd.n2812 0.0137576
R13104 vdd.n2866 vdd.n2799 0.0137576
R13105 vdd.n2894 vdd.n2893 0.0137576
R13106 vdd.n1030 vdd.n1029 0.0137576
R13107 vdd.n4512 vdd.n1011 0.0137576
R13108 vdd.n4503 vdd.n4502 0.0137576
R13109 vdd.n1099 vdd.n1098 0.0137576
R13110 vdd.n4485 vdd.n1079 0.0137576
R13111 vdd.n1155 vdd.n1154 0.0137576
R13112 vdd.n1174 vdd.n1173 0.0137576
R13113 vdd.n1197 vdd.n1196 0.0137576
R13114 vdd.n1216 vdd.n1215 0.0137576
R13115 vdd.n1239 vdd.n1238 0.0137576
R13116 vdd.n1253 vdd.n1252 0.0137576
R13117 vdd.n1251 vdd.n1248 0.0137576
R13118 vdd.n1294 vdd.n1293 0.0137576
R13119 vdd.n4391 vdd.n1279 0.0137576
R13120 vdd.n4382 vdd.n4381 0.0137576
R13121 vdd.n1363 vdd.n1362 0.0137576
R13122 vdd.n4364 vdd.n1343 0.0137576
R13123 vdd.n1419 vdd.n1418 0.0137576
R13124 vdd.n1438 vdd.n1437 0.0137576
R13125 vdd.n1461 vdd.n1460 0.0137576
R13126 vdd.n1480 vdd.n1479 0.0137576
R13127 vdd.n1503 vdd.n1502 0.0137576
R13128 vdd.n1517 vdd.n1516 0.0137576
R13129 vdd.n1515 vdd.n1512 0.0137576
R13130 vdd.n1558 vdd.n1557 0.0137576
R13131 vdd.n4270 vdd.n1543 0.0137576
R13132 vdd.n4261 vdd.n4260 0.0137576
R13133 vdd.n1627 vdd.n1626 0.0137576
R13134 vdd.n4243 vdd.n1607 0.0137576
R13135 vdd.n1683 vdd.n1682 0.0137576
R13136 vdd.n1702 vdd.n1701 0.0137576
R13137 vdd.n1725 vdd.n1724 0.0137576
R13138 vdd.n1744 vdd.n1743 0.0137576
R13139 vdd.n1767 vdd.n1766 0.0137576
R13140 vdd.n1781 vdd.n1780 0.0137576
R13141 vdd.n1779 vdd.n1776 0.0137576
R13142 vdd.n1822 vdd.n1821 0.0137576
R13143 vdd.n4149 vdd.n1807 0.0137576
R13144 vdd.n4140 vdd.n4139 0.0137576
R13145 vdd.n1891 vdd.n1890 0.0137576
R13146 vdd.n4122 vdd.n1871 0.0137576
R13147 vdd.n1947 vdd.n1946 0.0137576
R13148 vdd.n1966 vdd.n1965 0.0137576
R13149 vdd.n1989 vdd.n1988 0.0137576
R13150 vdd.n2008 vdd.n2007 0.0137576
R13151 vdd.n2031 vdd.n2030 0.0137576
R13152 vdd.n886 vdd.n885 0.0137576
R13153 vdd.n903 vdd.n902 0.0137576
R13154 vdd.n4564 vdd.n863 0.0137576
R13155 vdd.n4555 vdd.n4554 0.0137576
R13156 vdd.n972 vdd.n971 0.0137576
R13157 vdd.n4537 vdd.n952 0.0137576
R13158 vdd.n4689 vdd.n802 0.0137576
R13159 vdd.n4719 vdd.n790 0.0137576
R13160 vdd.n4737 vdd.n4736 0.0137576
R13161 vdd.n4748 vdd.n776 0.0137576
R13162 vdd.n4772 vdd.n762 0.0137576
R13163 vdd.n4799 vdd.n728 0.0137576
R13164 vdd.n4819 vdd.n722 0.0137576
R13165 vdd.n4834 vdd.n4833 0.0137576
R13166 vdd.n4855 vdd.n695 0.0137576
R13167 vdd.n4875 vdd.n688 0.0137576
R13168 vdd.n4894 vdd.n4893 0.0137576
R13169 vdd.n680 vdd.n679 0.0137576
R13170 vdd.n4917 vdd.n667 0.0137576
R13171 vdd.n4947 vdd.n655 0.0137576
R13172 vdd.n4965 vdd.n4964 0.0137576
R13173 vdd.n4976 vdd.n641 0.0137576
R13174 vdd.n5000 vdd.n627 0.0137576
R13175 vdd.n5027 vdd.n593 0.0137576
R13176 vdd.n5047 vdd.n587 0.0137576
R13177 vdd.n5062 vdd.n5061 0.0137576
R13178 vdd.n5083 vdd.n560 0.0137576
R13179 vdd.n5103 vdd.n553 0.0137576
R13180 vdd.n5122 vdd.n5121 0.0137576
R13181 vdd.n545 vdd.n544 0.0137576
R13182 vdd.n5145 vdd.n532 0.0137576
R13183 vdd.n5175 vdd.n520 0.0137576
R13184 vdd.n5193 vdd.n5192 0.0137576
R13185 vdd.n5204 vdd.n506 0.0137576
R13186 vdd.n5228 vdd.n492 0.0137576
R13187 vdd.n5255 vdd.n458 0.0137576
R13188 vdd.n5275 vdd.n452 0.0137576
R13189 vdd.n5290 vdd.n5289 0.0137576
R13190 vdd.n5311 vdd.n425 0.0137576
R13191 vdd.n5331 vdd.n418 0.0137576
R13192 vdd.n5350 vdd.n5349 0.0137576
R13193 vdd.n410 vdd.n409 0.0137576
R13194 vdd.n5373 vdd.n397 0.0137576
R13195 vdd.n5403 vdd.n385 0.0137576
R13196 vdd.n5421 vdd.n5420 0.0137576
R13197 vdd.n5432 vdd.n371 0.0137576
R13198 vdd.n5455 vdd.n357 0.0137576
R13199 vdd.n5488 vdd.n331 0.0137576
R13200 vdd.n5513 vdd.n314 0.0137576
R13201 vdd.n5528 vdd.n307 0.0137576
R13202 vdd.n5548 vdd.n301 0.0137576
R13203 vdd.n5567 vdd.n5566 0.0137576
R13204 vdd.n2126 vdd.n2122 0.0137243
R13205 vdd.n3897 vdd.n3893 0.0137243
R13206 vdd.n834 vdd.n830 0.0137243
R13207 vdd.n5769 vdd.n5765 0.0137243
R13208 vdd.n190 vdd.n189 0.0137188
R13209 vdd.n208 vdd.n200 0.0137188
R13210 vdd.n7498 vdd.n200 0.0137188
R13211 vdd.n3991 vdd.n3845 0.0137188
R13212 vdd.n3991 vdd.n3843 0.0137188
R13213 vdd.n4598 vdd.n4597 0.0137188
R13214 vdd.n4598 vdd.n4590 0.0137188
R13215 vdd.n5759 vdd.n220 0.0137188
R13216 vdd.n7471 vdd.n220 0.0137188
R13217 vdd.n3969 vdd.n3968 0.0134306
R13218 vdd.n4048 vdd.n2036 0.0133585
R13219 vdd.n7493 vdd.n207 0.0130393
R13220 vdd.n3995 vdd.n3840 0.0130393
R13221 vdd.n3987 vdd.n3851 0.0130393
R13222 vdd.n4602 vdd.n4591 0.0130393
R13223 vdd.n4629 vdd.n842 0.0130393
R13224 vdd.n5749 vdd.n239 0.0130393
R13225 vdd.n7473 vdd.n217 0.0130393
R13226 vdd.n119 vdd.n118 0.0130142
R13227 vdd.n3929 vdd.n3928 0.0129151
R13228 vdd.n114 vdd.n113 0.0128698
R13229 vdd.n74 vdd.n70 0.0128698
R13230 vdd.n2138 vdd.n2135 0.0127951
R13231 vdd.n123 vdd.n122 0.0125366
R13232 vdd.n2144 vdd.n2142 0.0118819
R13233 vdd.n88 vdd.n84 0.0115677
R13234 vdd.n173 vdd 0.0115677
R13235 vdd.n8 vdd 0.0109167
R13236 vdd.n3970 vdd 0.0108445
R13237 vdd.n2128 vdd.n2121 0.0105714
R13238 vdd.n2128 vdd.n2123 0.0105714
R13239 vdd.n3899 vdd.n3892 0.0105714
R13240 vdd.n3899 vdd.n3894 0.0105714
R13241 vdd.n836 vdd.n831 0.0105714
R13242 vdd.n5771 vdd.n5766 0.0105714
R13243 vdd.n3989 vdd.n3847 0.0105072
R13244 vdd.n7459 vdd.n7458 0.0103794
R13245 vdd.n7453 vdd.n237 0.0103794
R13246 vdd.n5742 vdd.n5740 0.0103794
R13247 vdd.n7438 vdd.n7432 0.0103794
R13248 vdd.n7443 vdd.n5776 0.0103794
R13249 vdd.n5785 vdd.n5784 0.0103794
R13250 vdd.n7428 vdd.n7427 0.0103794
R13251 vdd.n5809 vdd.n5808 0.0103794
R13252 vdd.n4665 vdd.n811 0.0103794
R13253 vdd.n4650 vdd.n4649 0.0103794
R13254 vdd.n4657 vdd.n817 0.0103794
R13255 vdd.n4640 vdd.n4639 0.0103794
R13256 vdd.n825 vdd.n824 0.0103794
R13257 vdd vdd.n7530 0.0102656
R13258 vdd.n8 vdd.n6 0.0102656
R13259 vdd.n6413 vdd.n6412 0.0099697
R13260 vdd.n6434 vdd.n6433 0.0099697
R13261 vdd.n6449 vdd.n6365 0.0099697
R13262 vdd.n6473 vdd.n6472 0.0099697
R13263 vdd.n6493 vdd.n6492 0.0099697
R13264 vdd.n6334 vdd.n6333 0.0099697
R13265 vdd.n6330 vdd.n6329 0.0099697
R13266 vdd.n6525 vdd.n6524 0.0099697
R13267 vdd.n6544 vdd.n6301 0.0099697
R13268 vdd.n6560 vdd.n6557 0.0099697
R13269 vdd.n6287 vdd.n6286 0.0099697
R13270 vdd.n6600 vdd.n6599 0.0099697
R13271 vdd.n6640 vdd.n6639 0.0099697
R13272 vdd.n6661 vdd.n6660 0.0099697
R13273 vdd.n6676 vdd.n6232 0.0099697
R13274 vdd.n6700 vdd.n6699 0.0099697
R13275 vdd.n6720 vdd.n6719 0.0099697
R13276 vdd.n6201 vdd.n6200 0.0099697
R13277 vdd.n6197 vdd.n6196 0.0099697
R13278 vdd.n6752 vdd.n6751 0.0099697
R13279 vdd.n6771 vdd.n6168 0.0099697
R13280 vdd.n6787 vdd.n6784 0.0099697
R13281 vdd.n6154 vdd.n6153 0.0099697
R13282 vdd.n6827 vdd.n6826 0.0099697
R13283 vdd.n6867 vdd.n6866 0.0099697
R13284 vdd.n6888 vdd.n6887 0.0099697
R13285 vdd.n6903 vdd.n6099 0.0099697
R13286 vdd.n6927 vdd.n6926 0.0099697
R13287 vdd.n6947 vdd.n6946 0.0099697
R13288 vdd.n6068 vdd.n6067 0.0099697
R13289 vdd.n6064 vdd.n6063 0.0099697
R13290 vdd.n6979 vdd.n6978 0.0099697
R13291 vdd.n6998 vdd.n6035 0.0099697
R13292 vdd.n7014 vdd.n7011 0.0099697
R13293 vdd.n6021 vdd.n6020 0.0099697
R13294 vdd.n7054 vdd.n7053 0.0099697
R13295 vdd.n7094 vdd.n7093 0.0099697
R13296 vdd.n7115 vdd.n7114 0.0099697
R13297 vdd.n7130 vdd.n5966 0.0099697
R13298 vdd.n7154 vdd.n7153 0.0099697
R13299 vdd.n7174 vdd.n7173 0.0099697
R13300 vdd.n5935 vdd.n5934 0.0099697
R13301 vdd.n5931 vdd.n5930 0.0099697
R13302 vdd.n7206 vdd.n7205 0.0099697
R13303 vdd.n7225 vdd.n5902 0.0099697
R13304 vdd.n7241 vdd.n7238 0.0099697
R13305 vdd.n5888 vdd.n5887 0.0099697
R13306 vdd.n7286 vdd.n7285 0.0099697
R13307 vdd.n7315 vdd.n7314 0.0099697
R13308 vdd.n7334 vdd.n7333 0.0099697
R13309 vdd.n7353 vdd.n7352 0.0099697
R13310 vdd.n7372 vdd.n7371 0.0099697
R13311 vdd.n7395 vdd.n7394 0.0099697
R13312 vdd.n4692 vdd.n4691 0.0099697
R13313 vdd.n4722 vdd.n4721 0.0099697
R13314 vdd.n4734 vdd.n4733 0.0099697
R13315 vdd.n4749 vdd.n775 0.0099697
R13316 vdd.n4775 vdd.n4774 0.0099697
R13317 vdd.n755 vdd.n754 0.0099697
R13318 vdd.n742 vdd.n741 0.0099697
R13319 vdd.n4801 vdd.n727 0.0099697
R13320 vdd.n4817 vdd.n4814 0.0099697
R13321 vdd.n713 vdd.n712 0.0099697
R13322 vdd.n4859 vdd.n694 0.0099697
R13323 vdd.n4873 vdd.n4870 0.0099697
R13324 vdd.n4920 vdd.n4919 0.0099697
R13325 vdd.n4950 vdd.n4949 0.0099697
R13326 vdd.n4962 vdd.n4961 0.0099697
R13327 vdd.n4977 vdd.n640 0.0099697
R13328 vdd.n5003 vdd.n5002 0.0099697
R13329 vdd.n620 vdd.n619 0.0099697
R13330 vdd.n607 vdd.n606 0.0099697
R13331 vdd.n5029 vdd.n592 0.0099697
R13332 vdd.n5045 vdd.n5042 0.0099697
R13333 vdd.n578 vdd.n577 0.0099697
R13334 vdd.n5087 vdd.n559 0.0099697
R13335 vdd.n5101 vdd.n5098 0.0099697
R13336 vdd.n5148 vdd.n5147 0.0099697
R13337 vdd.n5178 vdd.n5177 0.0099697
R13338 vdd.n5190 vdd.n5189 0.0099697
R13339 vdd.n5205 vdd.n505 0.0099697
R13340 vdd.n5231 vdd.n5230 0.0099697
R13341 vdd.n485 vdd.n484 0.0099697
R13342 vdd.n472 vdd.n471 0.0099697
R13343 vdd.n5257 vdd.n457 0.0099697
R13344 vdd.n5273 vdd.n5270 0.0099697
R13345 vdd.n443 vdd.n442 0.0099697
R13346 vdd.n5315 vdd.n424 0.0099697
R13347 vdd.n5329 vdd.n5326 0.0099697
R13348 vdd.n5376 vdd.n5375 0.0099697
R13349 vdd.n5406 vdd.n5405 0.0099697
R13350 vdd.n5418 vdd.n5417 0.0099697
R13351 vdd.n5433 vdd.n370 0.0099697
R13352 vdd.n5458 vdd.n5457 0.0099697
R13353 vdd.n350 vdd.n349 0.0099697
R13354 vdd.n346 vdd.n345 0.0099697
R13355 vdd.n5486 vdd.n5485 0.0099697
R13356 vdd.n5511 vdd.n5510 0.0099697
R13357 vdd.n5530 vdd.n306 0.0099697
R13358 vdd.n5546 vdd.n5543 0.0099697
R13359 vdd.n290 vdd.n289 0.0099697
R13360 vdd.n5590 vdd.n5587 0.0099697
R13361 vdd.n5614 vdd.n268 0.0099697
R13362 vdd.n5705 vdd.n5609 0.0099697
R13363 vdd.n5694 vdd.n5625 0.0099697
R13364 vdd.n5676 vdd.n5675 0.0099697
R13365 vdd.n2918 vdd.n2917 0.0099697
R13366 vdd.n2948 vdd.n2947 0.0099697
R13367 vdd.n2960 vdd.n2959 0.0099697
R13368 vdd.n2975 vdd.n2751 0.0099697
R13369 vdd.n3001 vdd.n3000 0.0099697
R13370 vdd.n2731 vdd.n2730 0.0099697
R13371 vdd.n2718 vdd.n2717 0.0099697
R13372 vdd.n3027 vdd.n2703 0.0099697
R13373 vdd.n3043 vdd.n3040 0.0099697
R13374 vdd.n2689 vdd.n2688 0.0099697
R13375 vdd.n3085 vdd.n2670 0.0099697
R13376 vdd.n3099 vdd.n3096 0.0099697
R13377 vdd.n3146 vdd.n3145 0.0099697
R13378 vdd.n3176 vdd.n3175 0.0099697
R13379 vdd.n3188 vdd.n3187 0.0099697
R13380 vdd.n3203 vdd.n2616 0.0099697
R13381 vdd.n3229 vdd.n3228 0.0099697
R13382 vdd.n2596 vdd.n2595 0.0099697
R13383 vdd.n2583 vdd.n2582 0.0099697
R13384 vdd.n3255 vdd.n2568 0.0099697
R13385 vdd.n3271 vdd.n3268 0.0099697
R13386 vdd.n2554 vdd.n2553 0.0099697
R13387 vdd.n3313 vdd.n2535 0.0099697
R13388 vdd.n3327 vdd.n3324 0.0099697
R13389 vdd.n3374 vdd.n3373 0.0099697
R13390 vdd.n3404 vdd.n3403 0.0099697
R13391 vdd.n3416 vdd.n3415 0.0099697
R13392 vdd.n3431 vdd.n2481 0.0099697
R13393 vdd.n3457 vdd.n3456 0.0099697
R13394 vdd.n2461 vdd.n2460 0.0099697
R13395 vdd.n2448 vdd.n2447 0.0099697
R13396 vdd.n3483 vdd.n2433 0.0099697
R13397 vdd.n3499 vdd.n3496 0.0099697
R13398 vdd.n2419 vdd.n2418 0.0099697
R13399 vdd.n3541 vdd.n2400 0.0099697
R13400 vdd.n3555 vdd.n3552 0.0099697
R13401 vdd.n3602 vdd.n3601 0.0099697
R13402 vdd.n3632 vdd.n3631 0.0099697
R13403 vdd.n3644 vdd.n3643 0.0099697
R13404 vdd.n3659 vdd.n2346 0.0099697
R13405 vdd.n3684 vdd.n3683 0.0099697
R13406 vdd.n2326 vdd.n2325 0.0099697
R13407 vdd.n2322 vdd.n2321 0.0099697
R13408 vdd.n3711 vdd.n3710 0.0099697
R13409 vdd.n3735 vdd.n3734 0.0099697
R13410 vdd.n3754 vdd.n2280 0.0099697
R13411 vdd.n3770 vdd.n3767 0.0099697
R13412 vdd.n2264 vdd.n2263 0.0099697
R13413 vdd.n4017 vdd.n2051 0.0099697
R13414 vdd.n2829 vdd.n2828 0.0099697
R13415 vdd.n2844 vdd.n2811 0.0099697
R13416 vdd.n2869 vdd.n2868 0.0099697
R13417 vdd.n2876 vdd.n2787 0.0099697
R13418 vdd.n1026 vdd.n1025 0.0099697
R13419 vdd.n4514 vdd.n1010 0.0099697
R13420 vdd.n1066 vdd.n1046 0.0099697
R13421 vdd.n1095 vdd.n1094 0.0099697
R13422 vdd.n4487 vdd.n1078 0.0099697
R13423 vdd.n1133 vdd.n1128 0.0099697
R13424 vdd.n1132 vdd.n1131 0.0099697
R13425 vdd.n4466 vdd.n1145 0.0099697
R13426 vdd.n1177 vdd.n1176 0.0099697
R13427 vdd.n4444 vdd.n1187 0.0099697
R13428 vdd.n1219 vdd.n1218 0.0099697
R13429 vdd.n4422 vdd.n1229 0.0099697
R13430 vdd.n1290 vdd.n1289 0.0099697
R13431 vdd.n4393 vdd.n1278 0.0099697
R13432 vdd.n1330 vdd.n1310 0.0099697
R13433 vdd.n1359 vdd.n1358 0.0099697
R13434 vdd.n4366 vdd.n1342 0.0099697
R13435 vdd.n1397 vdd.n1392 0.0099697
R13436 vdd.n1396 vdd.n1395 0.0099697
R13437 vdd.n4345 vdd.n1409 0.0099697
R13438 vdd.n1441 vdd.n1440 0.0099697
R13439 vdd.n4323 vdd.n1451 0.0099697
R13440 vdd.n1483 vdd.n1482 0.0099697
R13441 vdd.n4301 vdd.n1493 0.0099697
R13442 vdd.n1554 vdd.n1553 0.0099697
R13443 vdd.n4272 vdd.n1542 0.0099697
R13444 vdd.n1594 vdd.n1574 0.0099697
R13445 vdd.n1623 vdd.n1622 0.0099697
R13446 vdd.n4245 vdd.n1606 0.0099697
R13447 vdd.n1661 vdd.n1656 0.0099697
R13448 vdd.n1660 vdd.n1659 0.0099697
R13449 vdd.n4224 vdd.n1673 0.0099697
R13450 vdd.n1705 vdd.n1704 0.0099697
R13451 vdd.n4202 vdd.n1715 0.0099697
R13452 vdd.n1747 vdd.n1746 0.0099697
R13453 vdd.n4180 vdd.n1757 0.0099697
R13454 vdd.n1818 vdd.n1817 0.0099697
R13455 vdd.n4151 vdd.n1806 0.0099697
R13456 vdd.n1858 vdd.n1838 0.0099697
R13457 vdd.n1887 vdd.n1886 0.0099697
R13458 vdd.n4124 vdd.n1870 0.0099697
R13459 vdd.n1925 vdd.n1920 0.0099697
R13460 vdd.n1924 vdd.n1923 0.0099697
R13461 vdd.n4103 vdd.n1937 0.0099697
R13462 vdd.n1969 vdd.n1968 0.0099697
R13463 vdd.n4081 vdd.n1979 0.0099697
R13464 vdd.n2011 vdd.n2010 0.0099697
R13465 vdd.n4059 vdd.n2021 0.0099697
R13466 vdd.n899 vdd.n898 0.0099697
R13467 vdd.n4566 vdd.n862 0.0099697
R13468 vdd.n939 vdd.n919 0.0099697
R13469 vdd.n968 vdd.n967 0.0099697
R13470 vdd.n4539 vdd.n951 0.0099697
R13471 vdd.n2242 vdd.n2241 0.00993793
R13472 vdd.n2078 vdd.n2077 0.00993793
R13473 vdd.n2231 vdd.n2230 0.00993793
R13474 vdd.n2071 vdd.n2070 0.00993793
R13475 vdd.n2089 vdd.n2088 0.00993793
R13476 vdd.n2082 vdd.n2081 0.00993793
R13477 vdd.n3961 vdd.n3960 0.00993793
R13478 vdd.n3955 vdd.n3954 0.00993793
R13479 vdd.n3950 vdd.n3949 0.00993793
R13480 vdd.n3916 vdd.n3915 0.00993793
R13481 vdd.n3883 vdd.n3882 0.00993793
R13482 vdd.n3877 vdd.n3876 0.00993793
R13483 vdd.n3872 vdd.n3871 0.00993793
R13484 vdd.n3931 vdd.n3930 0.00993793
R13485 vdd.n3809 vdd.n3806 0.00993793
R13486 vdd.n2237 vdd.n2220 0.00935838
R13487 vdd.n2208 vdd.n2105 0.0093141
R13488 vdd.n5660 vdd.n5656 0.00926684
R13489 vdd.n7411 vdd.n5794 0.00926684
R13490 vdd.n7451 vdd.n7450 0.00895742
R13491 vdd.n878 vdd 0.0089359
R13492 vdd vdd.n2044 0.0089359
R13493 vdd.n2238 vdd.n2093 0.00889286
R13494 vdd.n2216 vdd.n2099 0.00851282
R13495 vdd.n4684 vdd.n804 0.00792105
R13496 vdd.n4743 vdd.n778 0.00792105
R13497 vdd.n4912 vdd.n669 0.00792105
R13498 vdd.n4971 vdd.n643 0.00792105
R13499 vdd.n5140 vdd.n534 0.00792105
R13500 vdd.n5199 vdd.n508 0.00792105
R13501 vdd.n5368 vdd.n399 0.00792105
R13502 vdd.n5427 vdd.n373 0.00792105
R13503 vdd.n6401 vdd.n6400 0.00792105
R13504 vdd.n6465 vdd.n6354 0.00792105
R13505 vdd.n6628 vdd.n6627 0.00792105
R13506 vdd.n6692 vdd.n6221 0.00792105
R13507 vdd.n6855 vdd.n6854 0.00792105
R13508 vdd.n6919 vdd.n6088 0.00792105
R13509 vdd.n7082 vdd.n7081 0.00792105
R13510 vdd.n7146 vdd.n5955 0.00792105
R13511 vdd.n4705 vdd.n793 0.00792105
R13512 vdd.n4711 vdd.n4709 0.00792105
R13513 vdd.n4766 vdd.n764 0.00792105
R13514 vdd.n4768 vdd.n733 0.00792105
R13515 vdd.n4796 vdd.n4795 0.00792105
R13516 vdd.n4823 vdd.n4822 0.00792105
R13517 vdd.n4830 vdd.n4829 0.00792105
R13518 vdd.n4852 vdd.n4850 0.00792105
R13519 vdd.n4879 vdd.n4878 0.00792105
R13520 vdd.n4890 vdd.n4885 0.00792105
R13521 vdd.n4933 vdd.n658 0.00792105
R13522 vdd.n4939 vdd.n4937 0.00792105
R13523 vdd.n4994 vdd.n629 0.00792105
R13524 vdd.n4996 vdd.n598 0.00792105
R13525 vdd.n5024 vdd.n5023 0.00792105
R13526 vdd.n5051 vdd.n5050 0.00792105
R13527 vdd.n5058 vdd.n5057 0.00792105
R13528 vdd.n5080 vdd.n5078 0.00792105
R13529 vdd.n5107 vdd.n5106 0.00792105
R13530 vdd.n5118 vdd.n5113 0.00792105
R13531 vdd.n5161 vdd.n523 0.00792105
R13532 vdd.n5167 vdd.n5165 0.00792105
R13533 vdd.n5222 vdd.n494 0.00792105
R13534 vdd.n5224 vdd.n463 0.00792105
R13535 vdd.n5252 vdd.n5251 0.00792105
R13536 vdd.n5279 vdd.n5278 0.00792105
R13537 vdd.n5286 vdd.n5285 0.00792105
R13538 vdd.n5308 vdd.n5306 0.00792105
R13539 vdd.n5335 vdd.n5334 0.00792105
R13540 vdd.n5346 vdd.n5341 0.00792105
R13541 vdd.n5389 vdd.n388 0.00792105
R13542 vdd.n5395 vdd.n5393 0.00792105
R13543 vdd.n5450 vdd.n359 0.00792105
R13544 vdd.n5470 vdd.n337 0.00792105
R13545 vdd.n5491 vdd.n329 0.00792105
R13546 vdd.n5493 vdd.n312 0.00792105
R13547 vdd.n5525 vdd.n5524 0.00792105
R13548 vdd.n5552 vdd.n5551 0.00792105
R13549 vdd.n5563 vdd.n5558 0.00792105
R13550 vdd.n5580 vdd.n277 0.00792105
R13551 vdd.n6422 vdd.n6420 0.00792105
R13552 vdd.n6443 vdd.n6368 0.00792105
R13553 vdd.n6485 vdd.n6343 0.00792105
R13554 vdd.n6504 vdd.n6321 0.00792105
R13555 vdd.n6506 vdd.n6307 0.00792105
R13556 vdd.n6539 vdd.n6538 0.00792105
R13557 vdd.n6566 vdd.n6565 0.00792105
R13558 vdd.n6573 vdd.n6572 0.00792105
R13559 vdd.n6594 vdd.n6593 0.00792105
R13560 vdd.n6618 vdd.n6617 0.00792105
R13561 vdd.n6649 vdd.n6647 0.00792105
R13562 vdd.n6670 vdd.n6235 0.00792105
R13563 vdd.n6712 vdd.n6210 0.00792105
R13564 vdd.n6731 vdd.n6188 0.00792105
R13565 vdd.n6733 vdd.n6174 0.00792105
R13566 vdd.n6766 vdd.n6765 0.00792105
R13567 vdd.n6793 vdd.n6792 0.00792105
R13568 vdd.n6800 vdd.n6799 0.00792105
R13569 vdd.n6821 vdd.n6820 0.00792105
R13570 vdd.n6845 vdd.n6844 0.00792105
R13571 vdd.n6876 vdd.n6874 0.00792105
R13572 vdd.n6897 vdd.n6102 0.00792105
R13573 vdd.n6939 vdd.n6077 0.00792105
R13574 vdd.n6958 vdd.n6055 0.00792105
R13575 vdd.n6960 vdd.n6041 0.00792105
R13576 vdd.n6993 vdd.n6992 0.00792105
R13577 vdd.n7020 vdd.n7019 0.00792105
R13578 vdd.n7027 vdd.n7026 0.00792105
R13579 vdd.n7048 vdd.n7047 0.00792105
R13580 vdd.n7072 vdd.n7071 0.00792105
R13581 vdd.n7103 vdd.n7101 0.00792105
R13582 vdd.n7124 vdd.n5969 0.00792105
R13583 vdd.n7166 vdd.n5944 0.00792105
R13584 vdd.n7185 vdd.n5922 0.00792105
R13585 vdd.n7187 vdd.n5908 0.00792105
R13586 vdd.n7220 vdd.n7219 0.00792105
R13587 vdd.n7247 vdd.n7246 0.00792105
R13588 vdd.n7254 vdd.n7253 0.00792105
R13589 vdd.n7279 vdd.n7274 0.00792105
R13590 vdd.n7295 vdd.n5863 0.00792105
R13591 vdd.n1019 vdd.n1018 0.00784375
R13592 vdd.n1035 vdd.n1016 0.00784375
R13593 vdd.n4508 vdd.n4507 0.00784375
R13594 vdd.n1088 vdd.n1086 0.00784375
R13595 vdd.n1104 vdd.n1084 0.00784375
R13596 vdd.n4481 vdd.n4480 0.00784375
R13597 vdd.n1158 vdd.n1152 0.00784375
R13598 vdd.n4459 vdd.n4458 0.00784375
R13599 vdd.n1200 vdd.n1194 0.00784375
R13600 vdd.n4437 vdd.n4436 0.00784375
R13601 vdd.n1242 vdd.n1236 0.00784375
R13602 vdd.n4415 vdd.n4414 0.00784375
R13603 vdd.n1286 vdd.n1246 0.00784375
R13604 vdd.n1299 vdd.n1284 0.00784375
R13605 vdd.n4387 vdd.n4386 0.00784375
R13606 vdd.n1352 vdd.n1350 0.00784375
R13607 vdd.n1368 vdd.n1348 0.00784375
R13608 vdd.n4360 vdd.n4359 0.00784375
R13609 vdd.n1422 vdd.n1416 0.00784375
R13610 vdd.n4338 vdd.n4337 0.00784375
R13611 vdd.n1464 vdd.n1458 0.00784375
R13612 vdd.n4316 vdd.n4315 0.00784375
R13613 vdd.n1506 vdd.n1500 0.00784375
R13614 vdd.n4294 vdd.n4293 0.00784375
R13615 vdd.n1550 vdd.n1510 0.00784375
R13616 vdd.n1563 vdd.n1548 0.00784375
R13617 vdd.n4266 vdd.n4265 0.00784375
R13618 vdd.n1616 vdd.n1614 0.00784375
R13619 vdd.n1632 vdd.n1612 0.00784375
R13620 vdd.n4239 vdd.n4238 0.00784375
R13621 vdd.n1686 vdd.n1680 0.00784375
R13622 vdd.n4217 vdd.n4216 0.00784375
R13623 vdd.n1728 vdd.n1722 0.00784375
R13624 vdd.n4195 vdd.n4194 0.00784375
R13625 vdd.n1770 vdd.n1764 0.00784375
R13626 vdd.n4173 vdd.n4172 0.00784375
R13627 vdd.n1814 vdd.n1774 0.00784375
R13628 vdd.n1827 vdd.n1812 0.00784375
R13629 vdd.n4145 vdd.n4144 0.00784375
R13630 vdd.n1880 vdd.n1878 0.00784375
R13631 vdd.n1896 vdd.n1876 0.00784375
R13632 vdd.n4118 vdd.n4117 0.00784375
R13633 vdd.n1950 vdd.n1944 0.00784375
R13634 vdd.n4096 vdd.n4095 0.00784375
R13635 vdd.n1992 vdd.n1986 0.00784375
R13636 vdd.n4074 vdd.n4073 0.00784375
R13637 vdd.n2034 vdd.n2028 0.00784375
R13638 vdd.n4052 vdd.n4051 0.00784375
R13639 vdd.n2910 vdd.n2780 0.00784375
R13640 vdd.n2931 vdd.n2769 0.00784375
R13641 vdd.n2937 vdd.n2935 0.00784375
R13642 vdd.n2969 vdd.n2754 0.00784375
R13643 vdd.n2992 vdd.n2740 0.00784375
R13644 vdd.n2994 vdd.n2709 0.00784375
R13645 vdd.n3022 vdd.n3021 0.00784375
R13646 vdd.n3049 vdd.n3048 0.00784375
R13647 vdd.n3056 vdd.n3055 0.00784375
R13648 vdd.n3078 vdd.n3076 0.00784375
R13649 vdd.n3105 vdd.n3104 0.00784375
R13650 vdd.n3116 vdd.n3111 0.00784375
R13651 vdd.n3138 vdd.n2645 0.00784375
R13652 vdd.n3159 vdd.n2634 0.00784375
R13653 vdd.n3165 vdd.n3163 0.00784375
R13654 vdd.n3197 vdd.n2619 0.00784375
R13655 vdd.n3220 vdd.n2605 0.00784375
R13656 vdd.n3222 vdd.n2574 0.00784375
R13657 vdd.n3250 vdd.n3249 0.00784375
R13658 vdd.n3277 vdd.n3276 0.00784375
R13659 vdd.n3284 vdd.n3283 0.00784375
R13660 vdd.n3306 vdd.n3304 0.00784375
R13661 vdd.n3333 vdd.n3332 0.00784375
R13662 vdd.n3344 vdd.n3339 0.00784375
R13663 vdd.n3366 vdd.n2510 0.00784375
R13664 vdd.n3387 vdd.n2499 0.00784375
R13665 vdd.n3393 vdd.n3391 0.00784375
R13666 vdd.n3425 vdd.n2484 0.00784375
R13667 vdd.n3448 vdd.n2470 0.00784375
R13668 vdd.n3450 vdd.n2439 0.00784375
R13669 vdd.n3478 vdd.n3477 0.00784375
R13670 vdd.n3505 vdd.n3504 0.00784375
R13671 vdd.n3512 vdd.n3511 0.00784375
R13672 vdd.n3534 vdd.n3532 0.00784375
R13673 vdd.n3561 vdd.n3560 0.00784375
R13674 vdd.n3572 vdd.n3567 0.00784375
R13675 vdd.n3594 vdd.n2375 0.00784375
R13676 vdd.n3615 vdd.n2364 0.00784375
R13677 vdd.n3621 vdd.n3619 0.00784375
R13678 vdd.n3653 vdd.n2349 0.00784375
R13679 vdd.n3676 vdd.n2335 0.00784375
R13680 vdd.n3696 vdd.n2313 0.00784375
R13681 vdd.n3716 vdd.n2304 0.00784375
R13682 vdd.n3718 vdd.n2286 0.00784375
R13683 vdd.n3749 vdd.n3748 0.00784375
R13684 vdd.n3776 vdd.n3775 0.00784375
R13685 vdd.n3787 vdd.n3782 0.00784375
R13686 vdd.n3804 vdd.n2251 0.00784375
R13687 vdd.n5596 vdd.n5595 0.0078057
R13688 vdd.n5713 vdd.n5602 0.0078057
R13689 vdd.n5633 vdd.n5603 0.0078057
R13690 vdd.n5646 vdd.n5631 0.0078057
R13691 vdd.n5687 vdd.n5686 0.0078057
R13692 vdd.n5661 vdd.n5660 0.0078057
R13693 vdd.n5656 vdd.n243 0.0078057
R13694 vdd.n5735 vdd.n243 0.0078057
R13695 vdd.n7309 vdd.n7308 0.0078057
R13696 vdd.n7328 vdd.n7327 0.0078057
R13697 vdd.n7347 vdd.n7346 0.0078057
R13698 vdd.n7366 vdd.n7365 0.0078057
R13699 vdd.n7389 vdd.n7384 0.0078057
R13700 vdd.n7385 vdd.n5794 0.0078057
R13701 vdd.n7412 vdd.n7411 0.0078057
R13702 vdd.n7418 vdd.n7412 0.0078057
R13703 vdd.n2159 vdd.n2158 0.00774506
R13704 vdd.n879 vdd.n838 0.00773077
R13705 vdd.n879 vdd.n878 0.00773077
R13706 vdd.n891 vdd.n870 0.00773077
R13707 vdd.n908 vdd.n868 0.00773077
R13708 vdd.n4560 vdd.n4559 0.00773077
R13709 vdd.n961 vdd.n959 0.00773077
R13710 vdd.n977 vdd.n957 0.00773077
R13711 vdd.n4533 vdd.n4532 0.00773077
R13712 vdd.n4046 vdd.n2037 0.00773077
R13713 vdd.n2044 vdd.n2037 0.00773077
R13714 vdd.n4037 vdd.n4036 0.00773077
R13715 vdd.n2818 vdd.n2816 0.00773077
R13716 vdd.n2838 vdd.n2814 0.00773077
R13717 vdd.n2861 vdd.n2801 0.00773077
R13718 vdd.n2888 vdd.n2790 0.00773077
R13719 vdd.n2899 vdd.n2783 0.00773077
R13720 vdd.n4675 vdd.n4674 0.00767368
R13721 vdd.n4686 vdd.n4685 0.00767368
R13722 vdd.n4707 vdd.n4706 0.00767368
R13723 vdd.n4710 vdd.n780 0.00767368
R13724 vdd.n4745 vdd.n4744 0.00767368
R13725 vdd.n4769 vdd.n4767 0.00767368
R13726 vdd.n4790 vdd.n4789 0.00767368
R13727 vdd.n4791 vdd.n719 0.00767368
R13728 vdd.n4828 vdd.n717 0.00767368
R13729 vdd.n4849 vdd.n699 0.00767368
R13730 vdd.n4851 vdd.n685 0.00767368
R13731 vdd.n4884 vdd.n683 0.00767368
R13732 vdd.n4889 vdd.n4888 0.00767368
R13733 vdd.n4914 vdd.n4913 0.00767368
R13734 vdd.n4935 vdd.n4934 0.00767368
R13735 vdd.n4938 vdd.n645 0.00767368
R13736 vdd.n4973 vdd.n4972 0.00767368
R13737 vdd.n4997 vdd.n4995 0.00767368
R13738 vdd.n5018 vdd.n5017 0.00767368
R13739 vdd.n5019 vdd.n584 0.00767368
R13740 vdd.n5056 vdd.n582 0.00767368
R13741 vdd.n5077 vdd.n564 0.00767368
R13742 vdd.n5079 vdd.n550 0.00767368
R13743 vdd.n5112 vdd.n548 0.00767368
R13744 vdd.n5117 vdd.n5116 0.00767368
R13745 vdd.n5142 vdd.n5141 0.00767368
R13746 vdd.n5163 vdd.n5162 0.00767368
R13747 vdd.n5166 vdd.n510 0.00767368
R13748 vdd.n5201 vdd.n5200 0.00767368
R13749 vdd.n5225 vdd.n5223 0.00767368
R13750 vdd.n5246 vdd.n5245 0.00767368
R13751 vdd.n5247 vdd.n449 0.00767368
R13752 vdd.n5284 vdd.n447 0.00767368
R13753 vdd.n5305 vdd.n429 0.00767368
R13754 vdd.n5307 vdd.n415 0.00767368
R13755 vdd.n5340 vdd.n413 0.00767368
R13756 vdd.n5345 vdd.n5344 0.00767368
R13757 vdd.n5370 vdd.n5369 0.00767368
R13758 vdd.n5391 vdd.n5390 0.00767368
R13759 vdd.n5394 vdd.n375 0.00767368
R13760 vdd.n5429 vdd.n5428 0.00767368
R13761 vdd.n5452 vdd.n5451 0.00767368
R13762 vdd.n5472 vdd.n5471 0.00767368
R13763 vdd.n5494 vdd.n5492 0.00767368
R13764 vdd.n5519 vdd.n5518 0.00767368
R13765 vdd.n5520 vdd.n298 0.00767368
R13766 vdd.n5557 vdd.n296 0.00767368
R13767 vdd.n5562 vdd.n5561 0.00767368
R13768 vdd.n6399 vdd.n6396 0.00767368
R13769 vdd.n6419 vdd.n6380 0.00767368
R13770 vdd.n6421 vdd.n6370 0.00767368
R13771 vdd.n6445 vdd.n6444 0.00767368
R13772 vdd.n6467 vdd.n6466 0.00767368
R13773 vdd.n6487 vdd.n6486 0.00767368
R13774 vdd.n6507 vdd.n6505 0.00767368
R13775 vdd.n6533 vdd.n6532 0.00767368
R13776 vdd.n6534 vdd.n6293 0.00767368
R13777 vdd.n6571 vdd.n6291 0.00767368
R13778 vdd.n6592 vdd.n6274 0.00767368
R13779 vdd.n6616 vdd.n6261 0.00767368
R13780 vdd.n6626 vdd.n6257 0.00767368
R13781 vdd.n6646 vdd.n6247 0.00767368
R13782 vdd.n6648 vdd.n6237 0.00767368
R13783 vdd.n6672 vdd.n6671 0.00767368
R13784 vdd.n6694 vdd.n6693 0.00767368
R13785 vdd.n6714 vdd.n6713 0.00767368
R13786 vdd.n6734 vdd.n6732 0.00767368
R13787 vdd.n6760 vdd.n6759 0.00767368
R13788 vdd.n6761 vdd.n6160 0.00767368
R13789 vdd.n6798 vdd.n6158 0.00767368
R13790 vdd.n6819 vdd.n6141 0.00767368
R13791 vdd.n6843 vdd.n6128 0.00767368
R13792 vdd.n6853 vdd.n6124 0.00767368
R13793 vdd.n6873 vdd.n6114 0.00767368
R13794 vdd.n6875 vdd.n6104 0.00767368
R13795 vdd.n6899 vdd.n6898 0.00767368
R13796 vdd.n6921 vdd.n6920 0.00767368
R13797 vdd.n6941 vdd.n6940 0.00767368
R13798 vdd.n6961 vdd.n6959 0.00767368
R13799 vdd.n6987 vdd.n6986 0.00767368
R13800 vdd.n6988 vdd.n6027 0.00767368
R13801 vdd.n7025 vdd.n6025 0.00767368
R13802 vdd.n7046 vdd.n6008 0.00767368
R13803 vdd.n7070 vdd.n5995 0.00767368
R13804 vdd.n7080 vdd.n5991 0.00767368
R13805 vdd.n7100 vdd.n5981 0.00767368
R13806 vdd.n7102 vdd.n5971 0.00767368
R13807 vdd.n7126 vdd.n7125 0.00767368
R13808 vdd.n7148 vdd.n7147 0.00767368
R13809 vdd.n7168 vdd.n7167 0.00767368
R13810 vdd.n7188 vdd.n7186 0.00767368
R13811 vdd.n7214 vdd.n7213 0.00767368
R13812 vdd.n7215 vdd.n5894 0.00767368
R13813 vdd.n7252 vdd.n5892 0.00767368
R13814 vdd.n7273 vdd.n5875 0.00767368
R13815 vdd.n7278 vdd.n7277 0.00767368
R13816 vdd.n4530 vdd.n983 0.00759896
R13817 vdd.n1034 vdd.n1033 0.00759896
R13818 vdd.n4509 vdd.n1040 0.00759896
R13819 vdd.n1087 vdd.n1041 0.00759896
R13820 vdd.n1103 vdd.n1102 0.00759896
R13821 vdd.n4482 vdd.n1109 0.00759896
R13822 vdd.n1151 vdd.n1110 0.00759896
R13823 vdd.n4460 vdd.n1159 0.00759896
R13824 vdd.n1193 vdd.n1160 0.00759896
R13825 vdd.n4438 vdd.n1201 0.00759896
R13826 vdd.n1235 vdd.n1202 0.00759896
R13827 vdd.n4416 vdd.n1243 0.00759896
R13828 vdd.n4411 vdd.n4410 0.00759896
R13829 vdd.n1298 vdd.n1297 0.00759896
R13830 vdd.n4388 vdd.n1304 0.00759896
R13831 vdd.n1351 vdd.n1305 0.00759896
R13832 vdd.n1367 vdd.n1366 0.00759896
R13833 vdd.n4361 vdd.n1373 0.00759896
R13834 vdd.n1415 vdd.n1374 0.00759896
R13835 vdd.n4339 vdd.n1423 0.00759896
R13836 vdd.n1457 vdd.n1424 0.00759896
R13837 vdd.n4317 vdd.n1465 0.00759896
R13838 vdd.n1499 vdd.n1466 0.00759896
R13839 vdd.n4295 vdd.n1507 0.00759896
R13840 vdd.n4290 vdd.n4289 0.00759896
R13841 vdd.n1562 vdd.n1561 0.00759896
R13842 vdd.n4267 vdd.n1568 0.00759896
R13843 vdd.n1615 vdd.n1569 0.00759896
R13844 vdd.n1631 vdd.n1630 0.00759896
R13845 vdd.n4240 vdd.n1637 0.00759896
R13846 vdd.n1679 vdd.n1638 0.00759896
R13847 vdd.n4218 vdd.n1687 0.00759896
R13848 vdd.n1721 vdd.n1688 0.00759896
R13849 vdd.n4196 vdd.n1729 0.00759896
R13850 vdd.n1763 vdd.n1730 0.00759896
R13851 vdd.n4174 vdd.n1771 0.00759896
R13852 vdd.n4169 vdd.n4168 0.00759896
R13853 vdd.n1826 vdd.n1825 0.00759896
R13854 vdd.n4146 vdd.n1832 0.00759896
R13855 vdd.n1879 vdd.n1833 0.00759896
R13856 vdd.n1895 vdd.n1894 0.00759896
R13857 vdd.n4119 vdd.n1901 0.00759896
R13858 vdd.n1943 vdd.n1902 0.00759896
R13859 vdd.n4097 vdd.n1951 0.00759896
R13860 vdd.n1985 vdd.n1952 0.00759896
R13861 vdd.n4075 vdd.n1993 0.00759896
R13862 vdd.n2027 vdd.n1994 0.00759896
R13863 vdd.n4053 vdd.n2035 0.00759896
R13864 vdd.n2901 vdd.n2900 0.00759896
R13865 vdd.n2912 vdd.n2911 0.00759896
R13866 vdd.n2933 vdd.n2932 0.00759896
R13867 vdd.n2936 vdd.n2756 0.00759896
R13868 vdd.n2971 vdd.n2970 0.00759896
R13869 vdd.n2995 vdd.n2993 0.00759896
R13870 vdd.n3016 vdd.n3015 0.00759896
R13871 vdd.n3017 vdd.n2695 0.00759896
R13872 vdd.n3054 vdd.n2693 0.00759896
R13873 vdd.n3075 vdd.n2675 0.00759896
R13874 vdd.n3077 vdd.n2661 0.00759896
R13875 vdd.n3110 vdd.n2659 0.00759896
R13876 vdd.n3115 vdd.n3114 0.00759896
R13877 vdd.n3140 vdd.n3139 0.00759896
R13878 vdd.n3161 vdd.n3160 0.00759896
R13879 vdd.n3164 vdd.n2621 0.00759896
R13880 vdd.n3199 vdd.n3198 0.00759896
R13881 vdd.n3223 vdd.n3221 0.00759896
R13882 vdd.n3244 vdd.n3243 0.00759896
R13883 vdd.n3245 vdd.n2560 0.00759896
R13884 vdd.n3282 vdd.n2558 0.00759896
R13885 vdd.n3303 vdd.n2540 0.00759896
R13886 vdd.n3305 vdd.n2526 0.00759896
R13887 vdd.n3338 vdd.n2524 0.00759896
R13888 vdd.n3343 vdd.n3342 0.00759896
R13889 vdd.n3368 vdd.n3367 0.00759896
R13890 vdd.n3389 vdd.n3388 0.00759896
R13891 vdd.n3392 vdd.n2486 0.00759896
R13892 vdd.n3427 vdd.n3426 0.00759896
R13893 vdd.n3451 vdd.n3449 0.00759896
R13894 vdd.n3472 vdd.n3471 0.00759896
R13895 vdd.n3473 vdd.n2425 0.00759896
R13896 vdd.n3510 vdd.n2423 0.00759896
R13897 vdd.n3531 vdd.n2405 0.00759896
R13898 vdd.n3533 vdd.n2391 0.00759896
R13899 vdd.n3566 vdd.n2389 0.00759896
R13900 vdd.n3571 vdd.n3570 0.00759896
R13901 vdd.n3596 vdd.n3595 0.00759896
R13902 vdd.n3617 vdd.n3616 0.00759896
R13903 vdd.n3620 vdd.n2351 0.00759896
R13904 vdd.n3655 vdd.n3654 0.00759896
R13905 vdd.n3678 vdd.n3677 0.00759896
R13906 vdd.n3698 vdd.n3697 0.00759896
R13907 vdd.n3719 vdd.n3717 0.00759896
R13908 vdd.n3743 vdd.n3742 0.00759896
R13909 vdd.n3744 vdd.n2272 0.00759896
R13910 vdd.n3781 vdd.n2270 0.00759896
R13911 vdd.n3786 vdd.n3785 0.00759896
R13912 vdd.n5583 vdd.n275 0.00756218
R13913 vdd.n5601 vdd.n273 0.00756218
R13914 vdd.n5637 vdd.n5636 0.00756218
R13915 vdd.n5688 vdd.n5647 0.00756218
R13916 vdd.n7307 vdd.n7298 0.00756218
R13917 vdd.n7326 vdd.n5852 0.00756218
R13918 vdd.n7364 vdd.n5830 0.00756218
R13919 vdd.n7383 vdd.n5819 0.00756218
R13920 vdd.n5712 vdd.n5711 0.00756218
R13921 vdd.n5655 vdd.n5648 0.00756218
R13922 vdd.n7345 vdd.n5841 0.00756218
R13923 vdd.n7388 vdd.n7387 0.00756218
R13924 vdd.n890 vdd.n889 0.00748974
R13925 vdd.n907 vdd.n906 0.00748974
R13926 vdd.n4561 vdd.n913 0.00748974
R13927 vdd.n960 vdd.n914 0.00748974
R13928 vdd.n976 vdd.n975 0.00748974
R13929 vdd.n4534 vdd.n982 0.00748974
R13930 vdd.n4038 vdd.n2045 0.00748974
R13931 vdd.n2817 vdd.n2046 0.00748974
R13932 vdd.n2824 vdd.n2823 0.00748974
R13933 vdd.n2840 vdd.n2839 0.00748974
R13934 vdd.n2863 vdd.n2862 0.00748974
R13935 vdd.n2890 vdd.n2889 0.00748974
R13936 vdd.n2218 vdd.n2217 0.00747321
R13937 vdd.n7487 vdd.n210 0.00701042
R13938 vdd.n7502 vdd.n197 0.00701042
R13939 vdd.n3860 vdd.n3859 0.00701042
R13940 vdd.n4613 vdd.n4588 0.00701042
R13941 vdd.n5757 vdd.n5756 0.00701042
R13942 vdd.n7467 vdd.n222 0.00701042
R13943 vdd.n105 vdd.n99 0.00701042
R13944 vdd vdd.n2102 0.00691026
R13945 vdd.n2179 vdd.n2108 0.00680401
R13946 vdd.n5747 vdd.n5737 0.0066978
R13947 vdd.n7415 vdd.n7414 0.00665101
R13948 vdd.n2156 vdd.n2155 0.00664754
R13949 vdd.n2137 vdd 0.00650962
R13950 vdd.n2203 vdd.n2202 0.00642324
R13951 vdd.n2148 vdd.n2115 0.00642324
R13952 vdd.n181 vdd.n180 0.00642324
R13953 vdd.n69 vdd.n68 0.00642324
R13954 vdd.n98 vdd.n97 0.00642324
R13955 vdd.n83 vdd.n82 0.00642324
R13956 vdd.n140 vdd.n139 0.00642324
R13957 vdd.n5 vdd.n4 0.00642324
R13958 vdd.n7529 vdd.n7528 0.00642324
R13959 vdd.n179 vdd.n163 0.00635938
R13960 vdd.n2247 vdd.n2240 0.00635126
R13961 vdd.n3826 vdd.n2075 0.00635126
R13962 vdd.n2235 vdd.n2228 0.00635126
R13963 vdd.n3829 vdd.n2072 0.00635126
R13964 vdd.n2092 vdd.n2086 0.00635126
R13965 vdd.n3815 vdd.n2083 0.00635126
R13966 vdd.n3964 vdd.n3959 0.00635126
R13967 vdd.n3967 vdd.n3953 0.00635126
R13968 vdd.n3971 vdd.n3951 0.00635126
R13969 vdd.n3927 vdd.n3914 0.00635126
R13970 vdd.n3905 vdd.n3881 0.00635126
R13971 vdd.n3908 vdd.n3875 0.00635126
R13972 vdd.n3938 vdd.n3873 0.00635126
R13973 vdd.n3935 vdd.n3912 0.00635126
R13974 vdd.n2209 vdd.n2208 0.00610897
R13975 vdd.n2236 vdd.n2227 0.00596512
R13976 vdd.n2229 vdd.n2227 0.00596512
R13977 vdd.n3830 vdd.n2073 0.00596512
R13978 vdd.n3830 vdd.n3828 0.00596512
R13979 vdd.n3827 vdd.n2074 0.00596512
R13980 vdd.n2076 vdd.n2074 0.00596512
R13981 vdd.n2246 vdd.n2239 0.00596512
R13982 vdd.n2248 vdd.n2239 0.00596512
R13983 vdd.n3811 vdd.n3805 0.00596512
R13984 vdd.n2185 vdd.n2184 0.005956
R13985 vdd.n2138 vdd.n2133 0.005956
R13986 vdd.n2155 vdd.n2112 0.005956
R13987 vdd.n2138 vdd.n2137 0.00594939
R13988 vdd.n2155 vdd.n2154 0.00594939
R13989 vdd.n2196 vdd.n2184 0.00593623
R13990 vdd.n7494 vdd.n204 0.00572581
R13991 vdd.n3864 vdd.n3857 0.00570833
R13992 vdd.n3864 vdd.n3863 0.00570833
R13993 vdd.n4617 vdd.n4587 0.00570833
R13994 vdd.n4617 vdd.n4616 0.00570833
R13995 vdd.n4685 vdd.n4684 0.00544737
R13996 vdd.n4706 vdd.n4705 0.00544737
R13997 vdd.n4711 vdd.n4710 0.00544737
R13998 vdd.n4744 vdd.n4743 0.00544737
R13999 vdd.n4767 vdd.n4766 0.00544737
R14000 vdd.n4795 vdd.n4791 0.00544737
R14001 vdd.n4823 vdd.n717 0.00544737
R14002 vdd.n4830 vdd.n699 0.00544737
R14003 vdd.n4852 vdd.n4851 0.00544737
R14004 vdd.n4879 vdd.n683 0.00544737
R14005 vdd.n4913 vdd.n4912 0.00544737
R14006 vdd.n4934 vdd.n4933 0.00544737
R14007 vdd.n4939 vdd.n4938 0.00544737
R14008 vdd.n4972 vdd.n4971 0.00544737
R14009 vdd.n4995 vdd.n4994 0.00544737
R14010 vdd.n5023 vdd.n5019 0.00544737
R14011 vdd.n5051 vdd.n582 0.00544737
R14012 vdd.n5058 vdd.n564 0.00544737
R14013 vdd.n5080 vdd.n5079 0.00544737
R14014 vdd.n5107 vdd.n548 0.00544737
R14015 vdd.n5141 vdd.n5140 0.00544737
R14016 vdd.n5162 vdd.n5161 0.00544737
R14017 vdd.n5167 vdd.n5166 0.00544737
R14018 vdd.n5200 vdd.n5199 0.00544737
R14019 vdd.n5223 vdd.n5222 0.00544737
R14020 vdd.n5251 vdd.n5247 0.00544737
R14021 vdd.n5279 vdd.n447 0.00544737
R14022 vdd.n5286 vdd.n429 0.00544737
R14023 vdd.n5308 vdd.n5307 0.00544737
R14024 vdd.n5335 vdd.n413 0.00544737
R14025 vdd.n5369 vdd.n5368 0.00544737
R14026 vdd.n5390 vdd.n5389 0.00544737
R14027 vdd.n5395 vdd.n5394 0.00544737
R14028 vdd.n5428 vdd.n5427 0.00544737
R14029 vdd.n5451 vdd.n5450 0.00544737
R14030 vdd.n5492 vdd.n5491 0.00544737
R14031 vdd.n5518 vdd.n312 0.00544737
R14032 vdd.n5524 vdd.n5520 0.00544737
R14033 vdd.n5552 vdd.n296 0.00544737
R14034 vdd.n5563 vdd.n5562 0.00544737
R14035 vdd.n6401 vdd.n6380 0.00544737
R14036 vdd.n6422 vdd.n6421 0.00544737
R14037 vdd.n6444 vdd.n6443 0.00544737
R14038 vdd.n6466 vdd.n6465 0.00544737
R14039 vdd.n6486 vdd.n6485 0.00544737
R14040 vdd.n6532 vdd.n6307 0.00544737
R14041 vdd.n6538 vdd.n6534 0.00544737
R14042 vdd.n6566 vdd.n6291 0.00544737
R14043 vdd.n6573 vdd.n6274 0.00544737
R14044 vdd.n6594 vdd.n6261 0.00544737
R14045 vdd.n6628 vdd.n6247 0.00544737
R14046 vdd.n6649 vdd.n6648 0.00544737
R14047 vdd.n6671 vdd.n6670 0.00544737
R14048 vdd.n6693 vdd.n6692 0.00544737
R14049 vdd.n6713 vdd.n6712 0.00544737
R14050 vdd.n6759 vdd.n6174 0.00544737
R14051 vdd.n6765 vdd.n6761 0.00544737
R14052 vdd.n6793 vdd.n6158 0.00544737
R14053 vdd.n6800 vdd.n6141 0.00544737
R14054 vdd.n6821 vdd.n6128 0.00544737
R14055 vdd.n6855 vdd.n6114 0.00544737
R14056 vdd.n6876 vdd.n6875 0.00544737
R14057 vdd.n6898 vdd.n6897 0.00544737
R14058 vdd.n6920 vdd.n6919 0.00544737
R14059 vdd.n6940 vdd.n6939 0.00544737
R14060 vdd.n6986 vdd.n6041 0.00544737
R14061 vdd.n6992 vdd.n6988 0.00544737
R14062 vdd.n7020 vdd.n6025 0.00544737
R14063 vdd.n7027 vdd.n6008 0.00544737
R14064 vdd.n7048 vdd.n5995 0.00544737
R14065 vdd.n7082 vdd.n5981 0.00544737
R14066 vdd.n7103 vdd.n7102 0.00544737
R14067 vdd.n7125 vdd.n7124 0.00544737
R14068 vdd.n7147 vdd.n7146 0.00544737
R14069 vdd.n7167 vdd.n7166 0.00544737
R14070 vdd.n7213 vdd.n5908 0.00544737
R14071 vdd.n7219 vdd.n7215 0.00544737
R14072 vdd.n7247 vdd.n5892 0.00544737
R14073 vdd.n7254 vdd.n5875 0.00544737
R14074 vdd.n7279 vdd.n7278 0.00544737
R14075 vdd.n1033 vdd.n1018 0.00539583
R14076 vdd.n1040 vdd.n1016 0.00539583
R14077 vdd.n4507 vdd.n1041 0.00539583
R14078 vdd.n1102 vdd.n1086 0.00539583
R14079 vdd.n1109 vdd.n1084 0.00539583
R14080 vdd.n1159 vdd.n1158 0.00539583
R14081 vdd.n4458 vdd.n1160 0.00539583
R14082 vdd.n1201 vdd.n1200 0.00539583
R14083 vdd.n4436 vdd.n1202 0.00539583
R14084 vdd.n1243 vdd.n1242 0.00539583
R14085 vdd.n1297 vdd.n1286 0.00539583
R14086 vdd.n1304 vdd.n1284 0.00539583
R14087 vdd.n4386 vdd.n1305 0.00539583
R14088 vdd.n1366 vdd.n1350 0.00539583
R14089 vdd.n1373 vdd.n1348 0.00539583
R14090 vdd.n1423 vdd.n1422 0.00539583
R14091 vdd.n4337 vdd.n1424 0.00539583
R14092 vdd.n1465 vdd.n1464 0.00539583
R14093 vdd.n4315 vdd.n1466 0.00539583
R14094 vdd.n1507 vdd.n1506 0.00539583
R14095 vdd.n1561 vdd.n1550 0.00539583
R14096 vdd.n1568 vdd.n1548 0.00539583
R14097 vdd.n4265 vdd.n1569 0.00539583
R14098 vdd.n1630 vdd.n1614 0.00539583
R14099 vdd.n1637 vdd.n1612 0.00539583
R14100 vdd.n1687 vdd.n1686 0.00539583
R14101 vdd.n4216 vdd.n1688 0.00539583
R14102 vdd.n1729 vdd.n1728 0.00539583
R14103 vdd.n4194 vdd.n1730 0.00539583
R14104 vdd.n1771 vdd.n1770 0.00539583
R14105 vdd.n1825 vdd.n1814 0.00539583
R14106 vdd.n1832 vdd.n1812 0.00539583
R14107 vdd.n4144 vdd.n1833 0.00539583
R14108 vdd.n1894 vdd.n1878 0.00539583
R14109 vdd.n1901 vdd.n1876 0.00539583
R14110 vdd.n1951 vdd.n1950 0.00539583
R14111 vdd.n4095 vdd.n1952 0.00539583
R14112 vdd.n1993 vdd.n1992 0.00539583
R14113 vdd.n4073 vdd.n1994 0.00539583
R14114 vdd.n2035 vdd.n2034 0.00539583
R14115 vdd.n2911 vdd.n2910 0.00539583
R14116 vdd.n2932 vdd.n2931 0.00539583
R14117 vdd.n2937 vdd.n2936 0.00539583
R14118 vdd.n2970 vdd.n2969 0.00539583
R14119 vdd.n2993 vdd.n2992 0.00539583
R14120 vdd.n3021 vdd.n3017 0.00539583
R14121 vdd.n3049 vdd.n2693 0.00539583
R14122 vdd.n3056 vdd.n2675 0.00539583
R14123 vdd.n3078 vdd.n3077 0.00539583
R14124 vdd.n3105 vdd.n2659 0.00539583
R14125 vdd.n3139 vdd.n3138 0.00539583
R14126 vdd.n3160 vdd.n3159 0.00539583
R14127 vdd.n3165 vdd.n3164 0.00539583
R14128 vdd.n3198 vdd.n3197 0.00539583
R14129 vdd.n3221 vdd.n3220 0.00539583
R14130 vdd.n3249 vdd.n3245 0.00539583
R14131 vdd.n3277 vdd.n2558 0.00539583
R14132 vdd.n3284 vdd.n2540 0.00539583
R14133 vdd.n3306 vdd.n3305 0.00539583
R14134 vdd.n3333 vdd.n2524 0.00539583
R14135 vdd.n3367 vdd.n3366 0.00539583
R14136 vdd.n3388 vdd.n3387 0.00539583
R14137 vdd.n3393 vdd.n3392 0.00539583
R14138 vdd.n3426 vdd.n3425 0.00539583
R14139 vdd.n3449 vdd.n3448 0.00539583
R14140 vdd.n3477 vdd.n3473 0.00539583
R14141 vdd.n3505 vdd.n2423 0.00539583
R14142 vdd.n3512 vdd.n2405 0.00539583
R14143 vdd.n3534 vdd.n3533 0.00539583
R14144 vdd.n3561 vdd.n2389 0.00539583
R14145 vdd.n3595 vdd.n3594 0.00539583
R14146 vdd.n3616 vdd.n3615 0.00539583
R14147 vdd.n3621 vdd.n3620 0.00539583
R14148 vdd.n3654 vdd.n3653 0.00539583
R14149 vdd.n3677 vdd.n3676 0.00539583
R14150 vdd.n3717 vdd.n3716 0.00539583
R14151 vdd.n3742 vdd.n2286 0.00539583
R14152 vdd.n3748 vdd.n3744 0.00539583
R14153 vdd.n3776 vdd.n2270 0.00539583
R14154 vdd.n3787 vdd.n3786 0.00539583
R14155 vdd.n5596 vdd.n273 0.00537047
R14156 vdd.n5713 vdd.n5712 0.00537047
R14157 vdd.n5636 vdd.n5633 0.00537047
R14158 vdd.n5647 vdd.n5646 0.00537047
R14159 vdd.n5686 vdd.n5648 0.00537047
R14160 vdd.n7309 vdd.n5852 0.00537047
R14161 vdd.n7328 vdd.n5841 0.00537047
R14162 vdd.n7347 vdd.n5830 0.00537047
R14163 vdd.n7366 vdd.n5819 0.00537047
R14164 vdd.n7389 vdd.n7388 0.00537047
R14165 vdd.n906 vdd.n870 0.00532051
R14166 vdd.n913 vdd.n868 0.00532051
R14167 vdd.n4559 vdd.n914 0.00532051
R14168 vdd.n975 vdd.n959 0.00532051
R14169 vdd.n982 vdd.n957 0.00532051
R14170 vdd.n4036 vdd.n2046 0.00532051
R14171 vdd.n2823 vdd.n2816 0.00532051
R14172 vdd.n2839 vdd.n2838 0.00532051
R14173 vdd.n2862 vdd.n2861 0.00532051
R14174 vdd.n2889 vdd.n2888 0.00532051
R14175 vdd.n2129 vdd.n2120 0.00518613
R14176 vdd.n3900 vdd.n3891 0.00518613
R14177 vdd.n4635 vdd.n4634 0.00511607
R14178 vdd.n7448 vdd.n7447 0.00511607
R14179 vdd.n2093 vdd.n2085 0.00507792
R14180 vdd.n2087 vdd.n2085 0.00507792
R14181 vdd.n3816 vdd.n2084 0.00507792
R14182 vdd.n3816 vdd.n3814 0.00507792
R14183 vdd.n205 vdd.n202 0.00507383
R14184 vdd.n3901 vdd.n3887 0.00493396
R14185 vdd.n3903 vdd.n3887 0.00493396
R14186 vdd.n3904 vdd.n3880 0.00493396
R14187 vdd.n3906 vdd.n3880 0.00493396
R14188 vdd.n3907 vdd.n3874 0.00493396
R14189 vdd.n3909 vdd.n3874 0.00493396
R14190 vdd.n3939 vdd.n3910 0.00493396
R14191 vdd.n3939 vdd.n3937 0.00493396
R14192 vdd.n3936 vdd.n3911 0.00493396
R14193 vdd.n3929 vdd.n3911 0.00493396
R14194 vdd.n3928 vdd.n3913 0.00493396
R14195 vdd.n3913 vdd.n2036 0.00493396
R14196 vdd.n5748 vdd.n242 0.00490305
R14197 vdd.n7419 vdd.n5793 0.00480499
R14198 vdd.n7518 vdd 0.00464286
R14199 vdd.n7516 vdd.n189 0.0045027
R14200 vdd.n7502 vdd.n7501 0.00440625
R14201 vdd.n7468 vdd.n7467 0.00440625
R14202 vdd.n7435 vdd.t1 0.00429204
R14203 vdd.n4652 vdd.t4 0.00429204
R14204 vdd.n6404 vdd.n6386 0.00428788
R14205 vdd.n6425 vdd.n6377 0.00428788
R14206 vdd.n6438 vdd.n6363 0.00428788
R14207 vdd.n6462 vdd.n6356 0.00428788
R14208 vdd.n6482 vdd.n6345 0.00428788
R14209 vdd.n6501 vdd.n6323 0.00428788
R14210 vdd.n6511 vdd.n6510 0.00428788
R14211 vdd.n6541 vdd.n6304 0.00428788
R14212 vdd.n6563 vdd.n6295 0.00428788
R14213 vdd.n6288 vdd.n6284 0.00428788
R14214 vdd.n6589 vdd.n6277 0.00428788
R14215 vdd.n6613 vdd.n6264 0.00428788
R14216 vdd.n6631 vdd.n6255 0.00428788
R14217 vdd.n6652 vdd.n6244 0.00428788
R14218 vdd.n6665 vdd.n6230 0.00428788
R14219 vdd.n6689 vdd.n6223 0.00428788
R14220 vdd.n6709 vdd.n6212 0.00428788
R14221 vdd.n6728 vdd.n6190 0.00428788
R14222 vdd.n6738 vdd.n6737 0.00428788
R14223 vdd.n6768 vdd.n6171 0.00428788
R14224 vdd.n6790 vdd.n6162 0.00428788
R14225 vdd.n6155 vdd.n6151 0.00428788
R14226 vdd.n6816 vdd.n6144 0.00428788
R14227 vdd.n6840 vdd.n6131 0.00428788
R14228 vdd.n6858 vdd.n6122 0.00428788
R14229 vdd.n6879 vdd.n6111 0.00428788
R14230 vdd.n6892 vdd.n6097 0.00428788
R14231 vdd.n6916 vdd.n6090 0.00428788
R14232 vdd.n6936 vdd.n6079 0.00428788
R14233 vdd.n6955 vdd.n6057 0.00428788
R14234 vdd.n6965 vdd.n6964 0.00428788
R14235 vdd.n6995 vdd.n6038 0.00428788
R14236 vdd.n7017 vdd.n6029 0.00428788
R14237 vdd.n6022 vdd.n6018 0.00428788
R14238 vdd.n7043 vdd.n6011 0.00428788
R14239 vdd.n7067 vdd.n5998 0.00428788
R14240 vdd.n7085 vdd.n5989 0.00428788
R14241 vdd.n7106 vdd.n5978 0.00428788
R14242 vdd.n7119 vdd.n5964 0.00428788
R14243 vdd.n7143 vdd.n5957 0.00428788
R14244 vdd.n7163 vdd.n5946 0.00428788
R14245 vdd.n7182 vdd.n5924 0.00428788
R14246 vdd.n7192 vdd.n7191 0.00428788
R14247 vdd.n7222 vdd.n5905 0.00428788
R14248 vdd.n7244 vdd.n5896 0.00428788
R14249 vdd.n5889 vdd.n5885 0.00428788
R14250 vdd.n7270 vdd.n5878 0.00428788
R14251 vdd.n5867 vdd.n5865 0.00428788
R14252 vdd.n7304 vdd.n7303 0.00428788
R14253 vdd.n7323 vdd.n5855 0.00428788
R14254 vdd.n7342 vdd.n5844 0.00428788
R14255 vdd.n7361 vdd.n5833 0.00428788
R14256 vdd.n7380 vdd.n5822 0.00428788
R14257 vdd.n7404 vdd.n7403 0.00428788
R14258 vdd.n5593 vdd.n5585 0.00428788
R14259 vdd.n269 vdd.n267 0.00428788
R14260 vdd.n5708 vdd.n5606 0.00428788
R14261 vdd.n5640 vdd.n5610 0.00428788
R14262 vdd.n5691 vdd.n5628 0.00428788
R14263 vdd.n5682 vdd.n5663 0.00428788
R14264 vdd.n2907 vdd.n2782 0.00428788
R14265 vdd.n2928 vdd.n2771 0.00428788
R14266 vdd.n2942 vdd.n2941 0.00428788
R14267 vdd.n2964 vdd.n2749 0.00428788
R14268 vdd.n2989 vdd.n2742 0.00428788
R14269 vdd.n3010 vdd.n2711 0.00428788
R14270 vdd.n3024 vdd.n2706 0.00428788
R14271 vdd.n3046 vdd.n2697 0.00428788
R14272 vdd.n2690 vdd.n2686 0.00428788
R14273 vdd.n3072 vdd.n2678 0.00428788
R14274 vdd.n3102 vdd.n2663 0.00428788
R14275 vdd.n2654 vdd.n2653 0.00428788
R14276 vdd.n3135 vdd.n2647 0.00428788
R14277 vdd.n3156 vdd.n2636 0.00428788
R14278 vdd.n3170 vdd.n3169 0.00428788
R14279 vdd.n3192 vdd.n2614 0.00428788
R14280 vdd.n3217 vdd.n2607 0.00428788
R14281 vdd.n3238 vdd.n2576 0.00428788
R14282 vdd.n3252 vdd.n2571 0.00428788
R14283 vdd.n3274 vdd.n2562 0.00428788
R14284 vdd.n2555 vdd.n2551 0.00428788
R14285 vdd.n3300 vdd.n2543 0.00428788
R14286 vdd.n3330 vdd.n2528 0.00428788
R14287 vdd.n2519 vdd.n2518 0.00428788
R14288 vdd.n3363 vdd.n2512 0.00428788
R14289 vdd.n3384 vdd.n2501 0.00428788
R14290 vdd.n3398 vdd.n3397 0.00428788
R14291 vdd.n3420 vdd.n2479 0.00428788
R14292 vdd.n3445 vdd.n2472 0.00428788
R14293 vdd.n3466 vdd.n2441 0.00428788
R14294 vdd.n3480 vdd.n2436 0.00428788
R14295 vdd.n3502 vdd.n2427 0.00428788
R14296 vdd.n2420 vdd.n2416 0.00428788
R14297 vdd.n3528 vdd.n2408 0.00428788
R14298 vdd.n3558 vdd.n2393 0.00428788
R14299 vdd.n2384 vdd.n2383 0.00428788
R14300 vdd.n3591 vdd.n2377 0.00428788
R14301 vdd.n3612 vdd.n2366 0.00428788
R14302 vdd.n3626 vdd.n3625 0.00428788
R14303 vdd.n3648 vdd.n2344 0.00428788
R14304 vdd.n3673 vdd.n2337 0.00428788
R14305 vdd.n3693 vdd.n2315 0.00428788
R14306 vdd.n3701 vdd.n2311 0.00428788
R14307 vdd.n3722 vdd.n2302 0.00428788
R14308 vdd.n3751 vdd.n2283 0.00428788
R14309 vdd.n3773 vdd.n2274 0.00428788
R14310 vdd.n2265 vdd.n2261 0.00428788
R14311 vdd.n2255 vdd.n2253 0.00428788
R14312 vdd.n4013 vdd.n2043 0.00428788
R14313 vdd.n2052 vdd.n2050 0.00428788
R14314 vdd.n2833 vdd.n2810 0.00428788
R14315 vdd.n2858 vdd.n2803 0.00428788
R14316 vdd.n2885 vdd.n2792 0.00428788
R14317 vdd.n2897 vdd.n2785 0.00428788
R14318 vdd.n986 vdd.n985 0.00428788
R14319 vdd.n1028 vdd.n1009 0.00428788
R14320 vdd.n4511 vdd.n1013 0.00428788
R14321 vdd.n1047 vdd.n1045 0.00428788
R14322 vdd.n1097 vdd.n1077 0.00428788
R14323 vdd.n4484 vdd.n1081 0.00428788
R14324 vdd.n4476 vdd.n1114 0.00428788
R14325 vdd.n4463 vdd.n1148 0.00428788
R14326 vdd.n4454 vdd.n1164 0.00428788
R14327 vdd.n4441 vdd.n1190 0.00428788
R14328 vdd.n4432 vdd.n1206 0.00428788
R14329 vdd.n4419 vdd.n1232 0.00428788
R14330 vdd.n4408 vdd.n4407 0.00428788
R14331 vdd.n1292 vdd.n1277 0.00428788
R14332 vdd.n4390 vdd.n1281 0.00428788
R14333 vdd.n1311 vdd.n1309 0.00428788
R14334 vdd.n1361 vdd.n1341 0.00428788
R14335 vdd.n4363 vdd.n1345 0.00428788
R14336 vdd.n4355 vdd.n1378 0.00428788
R14337 vdd.n4342 vdd.n1412 0.00428788
R14338 vdd.n4333 vdd.n1428 0.00428788
R14339 vdd.n4320 vdd.n1454 0.00428788
R14340 vdd.n4311 vdd.n1470 0.00428788
R14341 vdd.n4298 vdd.n1496 0.00428788
R14342 vdd.n4287 vdd.n4286 0.00428788
R14343 vdd.n1556 vdd.n1541 0.00428788
R14344 vdd.n4269 vdd.n1545 0.00428788
R14345 vdd.n1575 vdd.n1573 0.00428788
R14346 vdd.n1625 vdd.n1605 0.00428788
R14347 vdd.n4242 vdd.n1609 0.00428788
R14348 vdd.n4234 vdd.n1642 0.00428788
R14349 vdd.n4221 vdd.n1676 0.00428788
R14350 vdd.n4212 vdd.n1692 0.00428788
R14351 vdd.n4199 vdd.n1718 0.00428788
R14352 vdd.n4190 vdd.n1734 0.00428788
R14353 vdd.n4177 vdd.n1760 0.00428788
R14354 vdd.n4166 vdd.n4165 0.00428788
R14355 vdd.n1820 vdd.n1805 0.00428788
R14356 vdd.n4148 vdd.n1809 0.00428788
R14357 vdd.n1839 vdd.n1837 0.00428788
R14358 vdd.n1889 vdd.n1869 0.00428788
R14359 vdd.n4121 vdd.n1873 0.00428788
R14360 vdd.n4113 vdd.n1906 0.00428788
R14361 vdd.n4100 vdd.n1940 0.00428788
R14362 vdd.n4091 vdd.n1956 0.00428788
R14363 vdd.n4078 vdd.n1982 0.00428788
R14364 vdd.n4069 vdd.n1998 0.00428788
R14365 vdd.n4056 vdd.n2024 0.00428788
R14366 vdd.n894 vdd.n872 0.00428788
R14367 vdd.n901 vdd.n861 0.00428788
R14368 vdd.n4563 vdd.n865 0.00428788
R14369 vdd.n920 vdd.n918 0.00428788
R14370 vdd.n970 vdd.n950 0.00428788
R14371 vdd.n4536 vdd.n954 0.00428788
R14372 vdd.n4681 vdd.n806 0.00428788
R14373 vdd.n4702 vdd.n795 0.00428788
R14374 vdd.n4716 vdd.n4715 0.00428788
R14375 vdd.n4738 vdd.n773 0.00428788
R14376 vdd.n4763 vdd.n766 0.00428788
R14377 vdd.n4784 vdd.n735 0.00428788
R14378 vdd.n4798 vdd.n730 0.00428788
R14379 vdd.n4820 vdd.n721 0.00428788
R14380 vdd.n714 vdd.n710 0.00428788
R14381 vdd.n4846 vdd.n702 0.00428788
R14382 vdd.n4876 vdd.n687 0.00428788
R14383 vdd.n678 vdd.n677 0.00428788
R14384 vdd.n4909 vdd.n671 0.00428788
R14385 vdd.n4930 vdd.n660 0.00428788
R14386 vdd.n4944 vdd.n4943 0.00428788
R14387 vdd.n4966 vdd.n638 0.00428788
R14388 vdd.n4991 vdd.n631 0.00428788
R14389 vdd.n5012 vdd.n600 0.00428788
R14390 vdd.n5026 vdd.n595 0.00428788
R14391 vdd.n5048 vdd.n586 0.00428788
R14392 vdd.n579 vdd.n575 0.00428788
R14393 vdd.n5074 vdd.n567 0.00428788
R14394 vdd.n5104 vdd.n552 0.00428788
R14395 vdd.n543 vdd.n542 0.00428788
R14396 vdd.n5137 vdd.n536 0.00428788
R14397 vdd.n5158 vdd.n525 0.00428788
R14398 vdd.n5172 vdd.n5171 0.00428788
R14399 vdd.n5194 vdd.n503 0.00428788
R14400 vdd.n5219 vdd.n496 0.00428788
R14401 vdd.n5240 vdd.n465 0.00428788
R14402 vdd.n5254 vdd.n460 0.00428788
R14403 vdd.n5276 vdd.n451 0.00428788
R14404 vdd.n444 vdd.n440 0.00428788
R14405 vdd.n5302 vdd.n432 0.00428788
R14406 vdd.n5332 vdd.n417 0.00428788
R14407 vdd.n408 vdd.n407 0.00428788
R14408 vdd.n5365 vdd.n401 0.00428788
R14409 vdd.n5386 vdd.n390 0.00428788
R14410 vdd.n5400 vdd.n5399 0.00428788
R14411 vdd.n5422 vdd.n368 0.00428788
R14412 vdd.n5447 vdd.n361 0.00428788
R14413 vdd.n5467 vdd.n339 0.00428788
R14414 vdd.n5476 vdd.n5475 0.00428788
R14415 vdd.n5498 vdd.n5497 0.00428788
R14416 vdd.n5527 vdd.n309 0.00428788
R14417 vdd.n5549 vdd.n300 0.00428788
R14418 vdd.n291 vdd.n287 0.00428788
R14419 vdd.n281 vdd.n279 0.00428788
R14420 vdd.n3988 vdd.n3848 0.00428087
R14421 vdd.n3997 vdd.n3841 0.00428087
R14422 vdd.n4630 vdd.n841 0.00428087
R14423 vdd.n4604 vdd.n840 0.00428087
R14424 vdd.n7475 vdd.n218 0.00428087
R14425 vdd.n4669 vdd.n808 0.00397409
R14426 vdd.n6391 vdd.n6389 0.00397409
R14427 vdd.n5734 vdd.n244 0.00391036
R14428 vdd.n4045 vdd.n4044 0.00391036
R14429 vdd.n881 vdd.n880 0.00391036
R14430 vdd.n3958 vdd.n3847 0.00387321
R14431 vdd.n3965 vdd.n3958 0.00387321
R14432 vdd.n3966 vdd.n3952 0.00387321
R14433 vdd.n3968 vdd.n3952 0.00387321
R14434 vdd.n3972 vdd.n3969 0.00387321
R14435 vdd.n3972 vdd.n3970 0.00387321
R14436 vdd.n5747 vdd.n5746 0.00379258
R14437 vdd.n2226 vdd.n2221 0.00373256
R14438 vdd.n7494 vdd.n7493 0.00360776
R14439 vdd.n3988 vdd.n3987 0.00360776
R14440 vdd.n3841 vdd.n3840 0.00360776
R14441 vdd.n4630 vdd.n4629 0.00360776
R14442 vdd.n4591 vdd.n840 0.00360776
R14443 vdd.n5749 vdd.n5748 0.00360776
R14444 vdd.n218 vdd.n217 0.00360776
R14445 vdd.n2217 vdd.n2216 0.00360392
R14446 vdd.n2204 vdd.n2203 0.00360392
R14447 vdd.n2115 vdd.n2104 0.00360392
R14448 vdd.n180 vdd.n179 0.00360392
R14449 vdd.n70 vdd.n69 0.00360392
R14450 vdd.n99 vdd.n98 0.00360392
R14451 vdd.n84 vdd.n83 0.00360392
R14452 vdd.n139 vdd.n138 0.00360392
R14453 vdd.n6 vdd.n5 0.00360392
R14454 vdd.n7530 vdd.n7529 0.00360392
R14455 vdd.n2141 vdd.n2130 0.00354922
R14456 vdd.n7450 vdd 0.00353434
R14457 vdd.n836 vdd.n829 0.00351641
R14458 vdd.n5771 vdd.n5764 0.00351641
R14459 vdd.n118 vdd.n117 0.00336585
R14460 vdd.n122 vdd.n121 0.00336585
R14461 vdd.n126 vdd.n125 0.00336585
R14462 vdd.n145 vdd.n144 0.00336585
R14463 vdd.n186 vdd.n185 0.00336585
R14464 vdd.n7524 vdd.n7523 0.00336585
R14465 vdd.n7520 vdd.n7519 0.00336585
R14466 vdd.n2158 vdd.n2111 0.00328656
R14467 vdd.n2201 vdd.n2163 0.00328656
R14468 vdd.n116 vdd.n115 0.00327033
R14469 vdd.n120 vdd.n119 0.00327033
R14470 vdd.n124 vdd.n123 0.00327033
R14471 vdd.n143 vdd.n127 0.00327033
R14472 vdd.n184 vdd.n146 0.00327033
R14473 vdd.n7525 vdd.n187 0.00327033
R14474 vdd.n7522 vdd.n7521 0.00327033
R14475 vdd.n6529 vdd.n6528 0.00326471
R14476 vdd.n6537 vdd.n6306 0.00326471
R14477 vdd.n6567 vdd.n6292 0.00326471
R14478 vdd.n6575 vdd.n6574 0.00326471
R14479 vdd.n6596 vdd.n6595 0.00326471
R14480 vdd.n6620 vdd.n6619 0.00326471
R14481 vdd.n6756 vdd.n6755 0.00326471
R14482 vdd.n6764 vdd.n6173 0.00326471
R14483 vdd.n6794 vdd.n6159 0.00326471
R14484 vdd.n6802 vdd.n6801 0.00326471
R14485 vdd.n6823 vdd.n6822 0.00326471
R14486 vdd.n6847 vdd.n6846 0.00326471
R14487 vdd.n6983 vdd.n6982 0.00326471
R14488 vdd.n6991 vdd.n6040 0.00326471
R14489 vdd.n7021 vdd.n6026 0.00326471
R14490 vdd.n7029 vdd.n7028 0.00326471
R14491 vdd.n7050 vdd.n7049 0.00326471
R14492 vdd.n7074 vdd.n7073 0.00326471
R14493 vdd.n7210 vdd.n7209 0.00326471
R14494 vdd.n7218 vdd.n5907 0.00326471
R14495 vdd.n7248 vdd.n5893 0.00326471
R14496 vdd.n7256 vdd.n7255 0.00326471
R14497 vdd.n7281 vdd.n7280 0.00326471
R14498 vdd.n7311 vdd.n7310 0.00326471
R14499 vdd.n7330 vdd.n7329 0.00326471
R14500 vdd.n7349 vdd.n7348 0.00326471
R14501 vdd.n7368 vdd.n7367 0.00326471
R14502 vdd.n7391 vdd.n7390 0.00326471
R14503 vdd.n7408 vdd.n7407 0.00326471
R14504 vdd.n4794 vdd.n732 0.00326471
R14505 vdd.n4824 vdd.n718 0.00326471
R14506 vdd.n4832 vdd.n4831 0.00326471
R14507 vdd.n4854 vdd.n4853 0.00326471
R14508 vdd.n4880 vdd.n684 0.00326471
R14509 vdd.n4892 vdd.n4891 0.00326471
R14510 vdd.n5022 vdd.n597 0.00326471
R14511 vdd.n5052 vdd.n583 0.00326471
R14512 vdd.n5060 vdd.n5059 0.00326471
R14513 vdd.n5082 vdd.n5081 0.00326471
R14514 vdd.n5108 vdd.n549 0.00326471
R14515 vdd.n5120 vdd.n5119 0.00326471
R14516 vdd.n5250 vdd.n462 0.00326471
R14517 vdd.n5280 vdd.n448 0.00326471
R14518 vdd.n5288 vdd.n5287 0.00326471
R14519 vdd.n5310 vdd.n5309 0.00326471
R14520 vdd.n5336 vdd.n414 0.00326471
R14521 vdd.n5348 vdd.n5347 0.00326471
R14522 vdd.n5490 vdd.n5489 0.00326471
R14523 vdd.n5515 vdd.n5514 0.00326471
R14524 vdd.n5523 vdd.n311 0.00326471
R14525 vdd.n5553 vdd.n297 0.00326471
R14526 vdd.n5565 vdd.n5564 0.00326471
R14527 vdd.n5597 vdd.n274 0.00326471
R14528 vdd.n5715 vdd.n5714 0.00326471
R14529 vdd.n5634 vdd.n5605 0.00326471
R14530 vdd.n5645 vdd.n5644 0.00326471
R14531 vdd.n5685 vdd.n5649 0.00326471
R14532 vdd.n5659 vdd.n5654 0.00326471
R14533 vdd.n3020 vdd.n2708 0.00326471
R14534 vdd.n3050 vdd.n2694 0.00326471
R14535 vdd.n3058 vdd.n3057 0.00326471
R14536 vdd.n3080 vdd.n3079 0.00326471
R14537 vdd.n3106 vdd.n2660 0.00326471
R14538 vdd.n3118 vdd.n3117 0.00326471
R14539 vdd.n3248 vdd.n2573 0.00326471
R14540 vdd.n3278 vdd.n2559 0.00326471
R14541 vdd.n3286 vdd.n3285 0.00326471
R14542 vdd.n3308 vdd.n3307 0.00326471
R14543 vdd.n3334 vdd.n2525 0.00326471
R14544 vdd.n3346 vdd.n3345 0.00326471
R14545 vdd.n3476 vdd.n2438 0.00326471
R14546 vdd.n3506 vdd.n2424 0.00326471
R14547 vdd.n3514 vdd.n3513 0.00326471
R14548 vdd.n3536 vdd.n3535 0.00326471
R14549 vdd.n3562 vdd.n2390 0.00326471
R14550 vdd.n3574 vdd.n3573 0.00326471
R14551 vdd.n3715 vdd.n3714 0.00326471
R14552 vdd.n3739 vdd.n3738 0.00326471
R14553 vdd.n3747 vdd.n2285 0.00326471
R14554 vdd.n3777 vdd.n2271 0.00326471
R14555 vdd.n3789 vdd.n3788 0.00326471
R14556 vdd.n1157 vdd.n1156 0.00326471
R14557 vdd.n4457 vdd.n1161 0.00326471
R14558 vdd.n1199 vdd.n1198 0.00326471
R14559 vdd.n4435 vdd.n1203 0.00326471
R14560 vdd.n1241 vdd.n1240 0.00326471
R14561 vdd.n4413 vdd.n1244 0.00326471
R14562 vdd.n1421 vdd.n1420 0.00326471
R14563 vdd.n4336 vdd.n1425 0.00326471
R14564 vdd.n1463 vdd.n1462 0.00326471
R14565 vdd.n4314 vdd.n1467 0.00326471
R14566 vdd.n1505 vdd.n1504 0.00326471
R14567 vdd.n4292 vdd.n1508 0.00326471
R14568 vdd.n1685 vdd.n1684 0.00326471
R14569 vdd.n4215 vdd.n1689 0.00326471
R14570 vdd.n1727 vdd.n1726 0.00326471
R14571 vdd.n4193 vdd.n1731 0.00326471
R14572 vdd.n1769 vdd.n1768 0.00326471
R14573 vdd.n4171 vdd.n1772 0.00326471
R14574 vdd.n1949 vdd.n1948 0.00326471
R14575 vdd.n4094 vdd.n1953 0.00326471
R14576 vdd.n1991 vdd.n1990 0.00326471
R14577 vdd.n4072 vdd.n1995 0.00326471
R14578 vdd.n2033 vdd.n2032 0.00326471
R14579 vdd.n2162 vdd.n2159 0.00319368
R14580 vdd.n2200 vdd.n2164 0.00319368
R14581 vdd.n2145 vdd.n2144 0.00310079
R14582 vdd.n2143 vdd.n2095 0.00291834
R14583 vdd vdd.n2136 0.00290385
R14584 vdd.n2137 vdd.n2099 0.00290385
R14585 vdd.n3812 vdd.n3811 0.00281976
R14586 vdd.n2142 vdd.n2141 0.00273422
R14587 vdd.n2220 vdd.n2219 0.00273422
R14588 vdd.n3813 vdd.n2248 0.00268605
R14589 vdd.n6417 vdd.n6381 0.00257353
R14590 vdd.n6379 vdd.n6369 0.00257353
R14591 vdd.n6447 vdd.n6367 0.00257353
R14592 vdd.n6469 vdd.n6353 0.00257353
R14593 vdd.n6489 vdd.n6342 0.00257353
R14594 vdd.n6624 vdd.n6258 0.00257353
R14595 vdd.n6644 vdd.n6248 0.00257353
R14596 vdd.n6246 vdd.n6236 0.00257353
R14597 vdd.n6674 vdd.n6234 0.00257353
R14598 vdd.n6696 vdd.n6220 0.00257353
R14599 vdd.n6716 vdd.n6209 0.00257353
R14600 vdd.n6851 vdd.n6125 0.00257353
R14601 vdd.n6871 vdd.n6115 0.00257353
R14602 vdd.n6113 vdd.n6103 0.00257353
R14603 vdd.n6901 vdd.n6101 0.00257353
R14604 vdd.n6923 vdd.n6087 0.00257353
R14605 vdd.n6943 vdd.n6076 0.00257353
R14606 vdd.n7078 vdd.n5992 0.00257353
R14607 vdd.n7098 vdd.n5982 0.00257353
R14608 vdd.n5980 vdd.n5970 0.00257353
R14609 vdd.n7128 vdd.n5968 0.00257353
R14610 vdd.n7150 vdd.n5954 0.00257353
R14611 vdd.n7170 vdd.n5943 0.00257353
R14612 vdd.n4688 vdd.n803 0.00257353
R14613 vdd.n4718 vdd.n791 0.00257353
R14614 vdd.n4708 vdd.n779 0.00257353
R14615 vdd.n4747 vdd.n777 0.00257353
R14616 vdd.n4771 vdd.n763 0.00257353
R14617 vdd.n4886 vdd.n682 0.00257353
R14618 vdd.n4916 vdd.n668 0.00257353
R14619 vdd.n4946 vdd.n656 0.00257353
R14620 vdd.n4936 vdd.n644 0.00257353
R14621 vdd.n4975 vdd.n642 0.00257353
R14622 vdd.n4999 vdd.n628 0.00257353
R14623 vdd.n5114 vdd.n547 0.00257353
R14624 vdd.n5144 vdd.n533 0.00257353
R14625 vdd.n5174 vdd.n521 0.00257353
R14626 vdd.n5164 vdd.n509 0.00257353
R14627 vdd.n5203 vdd.n507 0.00257353
R14628 vdd.n5227 vdd.n493 0.00257353
R14629 vdd.n5342 vdd.n412 0.00257353
R14630 vdd.n5372 vdd.n398 0.00257353
R14631 vdd.n5402 vdd.n386 0.00257353
R14632 vdd.n5392 vdd.n374 0.00257353
R14633 vdd.n5431 vdd.n372 0.00257353
R14634 vdd.n5454 vdd.n358 0.00257353
R14635 vdd.n2914 vdd.n2779 0.00257353
R14636 vdd.n2944 vdd.n2767 0.00257353
R14637 vdd.n2934 vdd.n2755 0.00257353
R14638 vdd.n2973 vdd.n2753 0.00257353
R14639 vdd.n2997 vdd.n2739 0.00257353
R14640 vdd.n3112 vdd.n2658 0.00257353
R14641 vdd.n3142 vdd.n2644 0.00257353
R14642 vdd.n3172 vdd.n2632 0.00257353
R14643 vdd.n3162 vdd.n2620 0.00257353
R14644 vdd.n3201 vdd.n2618 0.00257353
R14645 vdd.n3225 vdd.n2604 0.00257353
R14646 vdd.n3340 vdd.n2523 0.00257353
R14647 vdd.n3370 vdd.n2509 0.00257353
R14648 vdd.n3400 vdd.n2497 0.00257353
R14649 vdd.n3390 vdd.n2485 0.00257353
R14650 vdd.n3429 vdd.n2483 0.00257353
R14651 vdd.n3453 vdd.n2469 0.00257353
R14652 vdd.n3568 vdd.n2388 0.00257353
R14653 vdd.n3598 vdd.n2374 0.00257353
R14654 vdd.n3628 vdd.n2362 0.00257353
R14655 vdd.n3618 vdd.n2350 0.00257353
R14656 vdd.n3657 vdd.n2348 0.00257353
R14657 vdd.n3680 vdd.n2334 0.00257353
R14658 vdd.n4040 vdd.n2041 0.00257353
R14659 vdd.n4034 vdd.n4033 0.00257353
R14660 vdd.n2822 vdd.n2815 0.00257353
R14661 vdd.n2842 vdd.n2813 0.00257353
R14662 vdd.n2865 vdd.n2800 0.00257353
R14663 vdd.n2892 vdd.n2789 0.00257353
R14664 vdd.n1032 vdd.n1031 0.00257353
R14665 vdd.n1039 vdd.n1014 0.00257353
R14666 vdd.n4505 vdd.n4504 0.00257353
R14667 vdd.n1101 vdd.n1100 0.00257353
R14668 vdd.n1108 vdd.n1082 0.00257353
R14669 vdd.n4412 vdd.n1245 0.00257353
R14670 vdd.n1296 vdd.n1295 0.00257353
R14671 vdd.n1303 vdd.n1282 0.00257353
R14672 vdd.n4384 vdd.n4383 0.00257353
R14673 vdd.n1365 vdd.n1364 0.00257353
R14674 vdd.n1372 vdd.n1346 0.00257353
R14675 vdd.n4291 vdd.n1509 0.00257353
R14676 vdd.n1560 vdd.n1559 0.00257353
R14677 vdd.n1567 vdd.n1546 0.00257353
R14678 vdd.n4263 vdd.n4262 0.00257353
R14679 vdd.n1629 vdd.n1628 0.00257353
R14680 vdd.n1636 vdd.n1610 0.00257353
R14681 vdd.n4170 vdd.n1773 0.00257353
R14682 vdd.n1824 vdd.n1823 0.00257353
R14683 vdd.n1831 vdd.n1810 0.00257353
R14684 vdd.n4142 vdd.n4141 0.00257353
R14685 vdd.n1893 vdd.n1892 0.00257353
R14686 vdd.n1900 vdd.n1874 0.00257353
R14687 vdd.n888 vdd.n887 0.00257353
R14688 vdd.n905 vdd.n904 0.00257353
R14689 vdd.n912 vdd.n866 0.00257353
R14690 vdd.n4557 vdd.n4556 0.00257353
R14691 vdd.n974 vdd.n973 0.00257353
R14692 vdd.n981 vdd.n955 0.00257353
R14693 vdd.n2203 vdd.n2109 0.00254918
R14694 vdd.n2217 vdd.n2098 0.00254918
R14695 vdd.n2139 vdd.n2138 0.00254918
R14696 vdd.n2155 vdd.n2153 0.00254918
R14697 vdd.n2184 vdd.n2166 0.00254918
R14698 vdd.n2118 vdd.n2115 0.00254918
R14699 vdd.n5 vdd.n0 0.00254918
R14700 vdd.n139 vdd.n129 0.00254918
R14701 vdd.n83 vdd.n78 0.00254918
R14702 vdd.n98 vdd.n93 0.00254918
R14703 vdd.n69 vdd.n64 0.00254918
R14704 vdd.n180 vdd.n148 0.00254918
R14705 vdd.n7529 vdd.n20 0.00254918
R14706 vdd.n4047 vdd 0.00252392
R14707 vdd.n4632 vdd 0.00252392
R14708 vdd.n7496 vdd.n7495 0.0025232
R14709 vdd.n2210 vdd.n2104 0.00250321
R14710 vdd.n7414 vdd.n7413 0.00249596
R14711 vdd.n6405 vdd.n6383 0.00239394
R14712 vdd.n6426 vdd.n6372 0.00239394
R14713 vdd.n6453 vdd.n6452 0.00239394
R14714 vdd.n6461 vdd.n6350 0.00239394
R14715 vdd.n6481 vdd.n6339 0.00239394
R14716 vdd.n6500 vdd.n6326 0.00239394
R14717 vdd.n6512 vdd.n6318 0.00239394
R14718 vdd.n6312 vdd.n6303 0.00239394
R14719 vdd.n6547 vdd.n6297 0.00239394
R14720 vdd.n6579 vdd.n6283 0.00239394
R14721 vdd.n6588 vdd.n6278 0.00239394
R14722 vdd.n6612 vdd.n6265 0.00239394
R14723 vdd.n6632 vdd.n6250 0.00239394
R14724 vdd.n6653 vdd.n6239 0.00239394
R14725 vdd.n6680 vdd.n6679 0.00239394
R14726 vdd.n6688 vdd.n6217 0.00239394
R14727 vdd.n6708 vdd.n6206 0.00239394
R14728 vdd.n6727 vdd.n6193 0.00239394
R14729 vdd.n6739 vdd.n6185 0.00239394
R14730 vdd.n6179 vdd.n6170 0.00239394
R14731 vdd.n6774 vdd.n6164 0.00239394
R14732 vdd.n6806 vdd.n6150 0.00239394
R14733 vdd.n6815 vdd.n6145 0.00239394
R14734 vdd.n6839 vdd.n6132 0.00239394
R14735 vdd.n6859 vdd.n6117 0.00239394
R14736 vdd.n6880 vdd.n6106 0.00239394
R14737 vdd.n6907 vdd.n6906 0.00239394
R14738 vdd.n6915 vdd.n6084 0.00239394
R14739 vdd.n6935 vdd.n6073 0.00239394
R14740 vdd.n6954 vdd.n6060 0.00239394
R14741 vdd.n6966 vdd.n6052 0.00239394
R14742 vdd.n6046 vdd.n6037 0.00239394
R14743 vdd.n7001 vdd.n6031 0.00239394
R14744 vdd.n7033 vdd.n6017 0.00239394
R14745 vdd.n7042 vdd.n6012 0.00239394
R14746 vdd.n7066 vdd.n5999 0.00239394
R14747 vdd.n7086 vdd.n5984 0.00239394
R14748 vdd.n7107 vdd.n5973 0.00239394
R14749 vdd.n7134 vdd.n7133 0.00239394
R14750 vdd.n7142 vdd.n5951 0.00239394
R14751 vdd.n7162 vdd.n5940 0.00239394
R14752 vdd.n7181 vdd.n5927 0.00239394
R14753 vdd.n7193 vdd.n5919 0.00239394
R14754 vdd.n5913 vdd.n5904 0.00239394
R14755 vdd.n7228 vdd.n5898 0.00239394
R14756 vdd.n7260 vdd.n5884 0.00239394
R14757 vdd.n7269 vdd.n5879 0.00239394
R14758 vdd.n7292 vdd.n5866 0.00239394
R14759 vdd.n6404 vdd.n6382 0.00239394
R14760 vdd.n6425 vdd.n6371 0.00239394
R14761 vdd.n6451 vdd.n6363 0.00239394
R14762 vdd.n6462 vdd.n6351 0.00239394
R14763 vdd.n6482 vdd.n6340 0.00239394
R14764 vdd.n6501 vdd.n6324 0.00239394
R14765 vdd.n6511 vdd.n6319 0.00239394
R14766 vdd.n6310 vdd.n6304 0.00239394
R14767 vdd.n6546 vdd.n6295 0.00239394
R14768 vdd.n6558 vdd.n6284 0.00239394
R14769 vdd.n6589 vdd.n6276 0.00239394
R14770 vdd.n6613 vdd.n6263 0.00239394
R14771 vdd.n6631 vdd.n6249 0.00239394
R14772 vdd.n6652 vdd.n6238 0.00239394
R14773 vdd.n6678 vdd.n6230 0.00239394
R14774 vdd.n6689 vdd.n6218 0.00239394
R14775 vdd.n6709 vdd.n6207 0.00239394
R14776 vdd.n6728 vdd.n6191 0.00239394
R14777 vdd.n6738 vdd.n6186 0.00239394
R14778 vdd.n6177 vdd.n6171 0.00239394
R14779 vdd.n6773 vdd.n6162 0.00239394
R14780 vdd.n6785 vdd.n6151 0.00239394
R14781 vdd.n6816 vdd.n6143 0.00239394
R14782 vdd.n6840 vdd.n6130 0.00239394
R14783 vdd.n6858 vdd.n6116 0.00239394
R14784 vdd.n6879 vdd.n6105 0.00239394
R14785 vdd.n6905 vdd.n6097 0.00239394
R14786 vdd.n6916 vdd.n6085 0.00239394
R14787 vdd.n6936 vdd.n6074 0.00239394
R14788 vdd.n6955 vdd.n6058 0.00239394
R14789 vdd.n6965 vdd.n6053 0.00239394
R14790 vdd.n6044 vdd.n6038 0.00239394
R14791 vdd.n7000 vdd.n6029 0.00239394
R14792 vdd.n7012 vdd.n6018 0.00239394
R14793 vdd.n7043 vdd.n6010 0.00239394
R14794 vdd.n7067 vdd.n5997 0.00239394
R14795 vdd.n7085 vdd.n5983 0.00239394
R14796 vdd.n7106 vdd.n5972 0.00239394
R14797 vdd.n7132 vdd.n5964 0.00239394
R14798 vdd.n7143 vdd.n5952 0.00239394
R14799 vdd.n7163 vdd.n5941 0.00239394
R14800 vdd.n7182 vdd.n5925 0.00239394
R14801 vdd.n7192 vdd.n5920 0.00239394
R14802 vdd.n5911 vdd.n5905 0.00239394
R14803 vdd.n7227 vdd.n5896 0.00239394
R14804 vdd.n7239 vdd.n5885 0.00239394
R14805 vdd.n7270 vdd.n5877 0.00239394
R14806 vdd.n7283 vdd.n5867 0.00239394
R14807 vdd.n7322 vdd.n5856 0.00239394
R14808 vdd.n7341 vdd.n5845 0.00239394
R14809 vdd.n7360 vdd.n5834 0.00239394
R14810 vdd.n7379 vdd.n5823 0.00239394
R14811 vdd.n7402 vdd.n5798 0.00239394
R14812 vdd.n7323 vdd.n5854 0.00239394
R14813 vdd.n7342 vdd.n5843 0.00239394
R14814 vdd.n7361 vdd.n5832 0.00239394
R14815 vdd.n7380 vdd.n5821 0.00239394
R14816 vdd.n7403 vdd.n5796 0.00239394
R14817 vdd.n4680 vdd.n800 0.00239394
R14818 vdd.n4701 vdd.n787 0.00239394
R14819 vdd.n4714 vdd.n782 0.00239394
R14820 vdd.n4753 vdd.n4752 0.00239394
R14821 vdd.n4762 vdd.n760 0.00239394
R14822 vdd.n4783 vdd.n738 0.00239394
R14823 vdd.n750 vdd.n729 0.00239394
R14824 vdd.n4804 vdd.n723 0.00239394
R14825 vdd.n4836 vdd.n709 0.00239394
R14826 vdd.n4845 vdd.n703 0.00239394
R14827 vdd.n4858 vdd.n689 0.00239394
R14828 vdd.n4896 vdd.n676 0.00239394
R14829 vdd.n4908 vdd.n665 0.00239394
R14830 vdd.n4929 vdd.n652 0.00239394
R14831 vdd.n4942 vdd.n647 0.00239394
R14832 vdd.n4981 vdd.n4980 0.00239394
R14833 vdd.n4990 vdd.n625 0.00239394
R14834 vdd.n5011 vdd.n603 0.00239394
R14835 vdd.n615 vdd.n594 0.00239394
R14836 vdd.n5032 vdd.n588 0.00239394
R14837 vdd.n5064 vdd.n574 0.00239394
R14838 vdd.n5073 vdd.n568 0.00239394
R14839 vdd.n5086 vdd.n554 0.00239394
R14840 vdd.n5124 vdd.n541 0.00239394
R14841 vdd.n5136 vdd.n530 0.00239394
R14842 vdd.n5157 vdd.n517 0.00239394
R14843 vdd.n5170 vdd.n512 0.00239394
R14844 vdd.n5209 vdd.n5208 0.00239394
R14845 vdd.n5218 vdd.n490 0.00239394
R14846 vdd.n5239 vdd.n468 0.00239394
R14847 vdd.n480 vdd.n459 0.00239394
R14848 vdd.n5260 vdd.n453 0.00239394
R14849 vdd.n5292 vdd.n439 0.00239394
R14850 vdd.n5301 vdd.n433 0.00239394
R14851 vdd.n5314 vdd.n419 0.00239394
R14852 vdd.n5352 vdd.n406 0.00239394
R14853 vdd.n5364 vdd.n395 0.00239394
R14854 vdd.n5385 vdd.n382 0.00239394
R14855 vdd.n5398 vdd.n377 0.00239394
R14856 vdd.n5437 vdd.n5436 0.00239394
R14857 vdd.n5446 vdd.n355 0.00239394
R14858 vdd.n5466 vdd.n342 0.00239394
R14859 vdd.n5477 vdd.n334 0.00239394
R14860 vdd.n5499 vdd.n326 0.00239394
R14861 vdd.n317 vdd.n308 0.00239394
R14862 vdd.n5533 vdd.n302 0.00239394
R14863 vdd.n5569 vdd.n286 0.00239394
R14864 vdd.n5577 vdd.n280 0.00239394
R14865 vdd.n5719 vdd.n266 0.00239394
R14866 vdd.n5616 vdd.n5608 0.00239394
R14867 vdd.n5702 vdd.n5611 0.00239394
R14868 vdd.n5693 vdd.n5626 0.00239394
R14869 vdd.n5681 vdd.n5664 0.00239394
R14870 vdd.n5588 vdd.n267 0.00239394
R14871 vdd.n5615 vdd.n5606 0.00239394
R14872 vdd.n5703 vdd.n5610 0.00239394
R14873 vdd.n5692 vdd.n5691 0.00239394
R14874 vdd.n5682 vdd.n5651 0.00239394
R14875 vdd.n2906 vdd.n2776 0.00239394
R14876 vdd.n2927 vdd.n2763 0.00239394
R14877 vdd.n2940 vdd.n2758 0.00239394
R14878 vdd.n2979 vdd.n2978 0.00239394
R14879 vdd.n2988 vdd.n2736 0.00239394
R14880 vdd.n3009 vdd.n2714 0.00239394
R14881 vdd.n2726 vdd.n2705 0.00239394
R14882 vdd.n3030 vdd.n2699 0.00239394
R14883 vdd.n3062 vdd.n2685 0.00239394
R14884 vdd.n3071 vdd.n2679 0.00239394
R14885 vdd.n3084 vdd.n2665 0.00239394
R14886 vdd.n3122 vdd.n2652 0.00239394
R14887 vdd.n3134 vdd.n2641 0.00239394
R14888 vdd.n3155 vdd.n2628 0.00239394
R14889 vdd.n3168 vdd.n2623 0.00239394
R14890 vdd.n3207 vdd.n3206 0.00239394
R14891 vdd.n3216 vdd.n2601 0.00239394
R14892 vdd.n3237 vdd.n2579 0.00239394
R14893 vdd.n2591 vdd.n2570 0.00239394
R14894 vdd.n3258 vdd.n2564 0.00239394
R14895 vdd.n3290 vdd.n2550 0.00239394
R14896 vdd.n3299 vdd.n2544 0.00239394
R14897 vdd.n3312 vdd.n2530 0.00239394
R14898 vdd.n3350 vdd.n2517 0.00239394
R14899 vdd.n3362 vdd.n2506 0.00239394
R14900 vdd.n3383 vdd.n2493 0.00239394
R14901 vdd.n3396 vdd.n2488 0.00239394
R14902 vdd.n3435 vdd.n3434 0.00239394
R14903 vdd.n3444 vdd.n2466 0.00239394
R14904 vdd.n3465 vdd.n2444 0.00239394
R14905 vdd.n2456 vdd.n2435 0.00239394
R14906 vdd.n3486 vdd.n2429 0.00239394
R14907 vdd.n3518 vdd.n2415 0.00239394
R14908 vdd.n3527 vdd.n2409 0.00239394
R14909 vdd.n3540 vdd.n2395 0.00239394
R14910 vdd.n3578 vdd.n2382 0.00239394
R14911 vdd.n3590 vdd.n2371 0.00239394
R14912 vdd.n3611 vdd.n2358 0.00239394
R14913 vdd.n3624 vdd.n2353 0.00239394
R14914 vdd.n3663 vdd.n3662 0.00239394
R14915 vdd.n3672 vdd.n2331 0.00239394
R14916 vdd.n3692 vdd.n2318 0.00239394
R14917 vdd.n3702 vdd.n2309 0.00239394
R14918 vdd.n3723 vdd.n2300 0.00239394
R14919 vdd.n2291 vdd.n2282 0.00239394
R14920 vdd.n3757 vdd.n2276 0.00239394
R14921 vdd.n3793 vdd.n2260 0.00239394
R14922 vdd.n3801 vdd.n2254 0.00239394
R14923 vdd.n2907 vdd.n2777 0.00239394
R14924 vdd.n2928 vdd.n2765 0.00239394
R14925 vdd.n2941 vdd.n2757 0.00239394
R14926 vdd.n2977 vdd.n2749 0.00239394
R14927 vdd.n2989 vdd.n2737 0.00239394
R14928 vdd.n3010 vdd.n2712 0.00239394
R14929 vdd.n2727 vdd.n2706 0.00239394
R14930 vdd.n3029 vdd.n2697 0.00239394
R14931 vdd.n3041 vdd.n2686 0.00239394
R14932 vdd.n3072 vdd.n2677 0.00239394
R14933 vdd.n3083 vdd.n2663 0.00239394
R14934 vdd.n3097 vdd.n2653 0.00239394
R14935 vdd.n3135 vdd.n2642 0.00239394
R14936 vdd.n3156 vdd.n2630 0.00239394
R14937 vdd.n3169 vdd.n2622 0.00239394
R14938 vdd.n3205 vdd.n2614 0.00239394
R14939 vdd.n3217 vdd.n2602 0.00239394
R14940 vdd.n3238 vdd.n2577 0.00239394
R14941 vdd.n2592 vdd.n2571 0.00239394
R14942 vdd.n3257 vdd.n2562 0.00239394
R14943 vdd.n3269 vdd.n2551 0.00239394
R14944 vdd.n3300 vdd.n2542 0.00239394
R14945 vdd.n3311 vdd.n2528 0.00239394
R14946 vdd.n3325 vdd.n2518 0.00239394
R14947 vdd.n3363 vdd.n2507 0.00239394
R14948 vdd.n3384 vdd.n2495 0.00239394
R14949 vdd.n3397 vdd.n2487 0.00239394
R14950 vdd.n3433 vdd.n2479 0.00239394
R14951 vdd.n3445 vdd.n2467 0.00239394
R14952 vdd.n3466 vdd.n2442 0.00239394
R14953 vdd.n2457 vdd.n2436 0.00239394
R14954 vdd.n3485 vdd.n2427 0.00239394
R14955 vdd.n3497 vdd.n2416 0.00239394
R14956 vdd.n3528 vdd.n2407 0.00239394
R14957 vdd.n3539 vdd.n2393 0.00239394
R14958 vdd.n3553 vdd.n2383 0.00239394
R14959 vdd.n3591 vdd.n2372 0.00239394
R14960 vdd.n3612 vdd.n2360 0.00239394
R14961 vdd.n3625 vdd.n2352 0.00239394
R14962 vdd.n3661 vdd.n2344 0.00239394
R14963 vdd.n3673 vdd.n2332 0.00239394
R14964 vdd.n3693 vdd.n2316 0.00239394
R14965 vdd.n3701 vdd.n2310 0.00239394
R14966 vdd.n3722 vdd.n2301 0.00239394
R14967 vdd.n2289 vdd.n2283 0.00239394
R14968 vdd.n3756 vdd.n2274 0.00239394
R14969 vdd.n3768 vdd.n2261 0.00239394
R14970 vdd.n2266 vdd.n2255 0.00239394
R14971 vdd.n4020 vdd.n4019 0.00239394
R14972 vdd.n4029 vdd.n2053 0.00239394
R14973 vdd.n2848 vdd.n2847 0.00239394
R14974 vdd.n2857 vdd.n2797 0.00239394
R14975 vdd.n2884 vdd.n2795 0.00239394
R14976 vdd.n4018 vdd.n4013 0.00239394
R14977 vdd.n2825 vdd.n2052 0.00239394
R14978 vdd.n2846 vdd.n2810 0.00239394
R14979 vdd.n2858 vdd.n2798 0.00239394
R14980 vdd.n2885 vdd.n2793 0.00239394
R14981 vdd.n4527 vdd.n987 0.00239394
R14982 vdd.n4518 vdd.n4517 0.00239394
R14983 vdd.n1065 vdd.n1012 0.00239394
R14984 vdd.n4500 vdd.n1048 0.00239394
R14985 vdd.n4491 vdd.n4490 0.00239394
R14986 vdd.n1136 vdd.n1080 0.00239394
R14987 vdd.n4475 vdd.n1115 0.00239394
R14988 vdd.n4465 vdd.n1146 0.00239394
R14989 vdd.n4453 vdd.n1165 0.00239394
R14990 vdd.n4443 vdd.n1188 0.00239394
R14991 vdd.n4431 vdd.n1207 0.00239394
R14992 vdd.n4421 vdd.n1230 0.00239394
R14993 vdd.n4406 vdd.n1256 0.00239394
R14994 vdd.n4397 vdd.n4396 0.00239394
R14995 vdd.n1329 vdd.n1280 0.00239394
R14996 vdd.n4379 vdd.n1312 0.00239394
R14997 vdd.n4370 vdd.n4369 0.00239394
R14998 vdd.n1400 vdd.n1344 0.00239394
R14999 vdd.n4354 vdd.n1379 0.00239394
R15000 vdd.n4344 vdd.n1410 0.00239394
R15001 vdd.n4332 vdd.n1429 0.00239394
R15002 vdd.n4322 vdd.n1452 0.00239394
R15003 vdd.n4310 vdd.n1471 0.00239394
R15004 vdd.n4300 vdd.n1494 0.00239394
R15005 vdd.n4285 vdd.n1520 0.00239394
R15006 vdd.n4276 vdd.n4275 0.00239394
R15007 vdd.n1593 vdd.n1544 0.00239394
R15008 vdd.n4258 vdd.n1576 0.00239394
R15009 vdd.n4249 vdd.n4248 0.00239394
R15010 vdd.n1664 vdd.n1608 0.00239394
R15011 vdd.n4233 vdd.n1643 0.00239394
R15012 vdd.n4223 vdd.n1674 0.00239394
R15013 vdd.n4211 vdd.n1693 0.00239394
R15014 vdd.n4201 vdd.n1716 0.00239394
R15015 vdd.n4189 vdd.n1735 0.00239394
R15016 vdd.n4179 vdd.n1758 0.00239394
R15017 vdd.n4164 vdd.n1784 0.00239394
R15018 vdd.n4155 vdd.n4154 0.00239394
R15019 vdd.n1857 vdd.n1808 0.00239394
R15020 vdd.n4137 vdd.n1840 0.00239394
R15021 vdd.n4128 vdd.n4127 0.00239394
R15022 vdd.n1928 vdd.n1872 0.00239394
R15023 vdd.n4112 vdd.n1907 0.00239394
R15024 vdd.n4102 vdd.n1938 0.00239394
R15025 vdd.n4090 vdd.n1957 0.00239394
R15026 vdd.n4080 vdd.n1980 0.00239394
R15027 vdd.n4068 vdd.n1999 0.00239394
R15028 vdd.n4058 vdd.n2022 0.00239394
R15029 vdd.n1023 vdd.n986 0.00239394
R15030 vdd.n4516 vdd.n1009 0.00239394
R15031 vdd.n1064 vdd.n1013 0.00239394
R15032 vdd.n1092 vdd.n1047 0.00239394
R15033 vdd.n4489 vdd.n1077 0.00239394
R15034 vdd.n1135 vdd.n1081 0.00239394
R15035 vdd.n4476 vdd.n1113 0.00239394
R15036 vdd.n4464 vdd.n4463 0.00239394
R15037 vdd.n4454 vdd.n1163 0.00239394
R15038 vdd.n4442 vdd.n4441 0.00239394
R15039 vdd.n4432 vdd.n1205 0.00239394
R15040 vdd.n4420 vdd.n4419 0.00239394
R15041 vdd.n4407 vdd.n1249 0.00239394
R15042 vdd.n4395 vdd.n1277 0.00239394
R15043 vdd.n1328 vdd.n1281 0.00239394
R15044 vdd.n1356 vdd.n1311 0.00239394
R15045 vdd.n4368 vdd.n1341 0.00239394
R15046 vdd.n1399 vdd.n1345 0.00239394
R15047 vdd.n4355 vdd.n1377 0.00239394
R15048 vdd.n4343 vdd.n4342 0.00239394
R15049 vdd.n4333 vdd.n1427 0.00239394
R15050 vdd.n4321 vdd.n4320 0.00239394
R15051 vdd.n4311 vdd.n1469 0.00239394
R15052 vdd.n4299 vdd.n4298 0.00239394
R15053 vdd.n4286 vdd.n1513 0.00239394
R15054 vdd.n4274 vdd.n1541 0.00239394
R15055 vdd.n1592 vdd.n1545 0.00239394
R15056 vdd.n1620 vdd.n1575 0.00239394
R15057 vdd.n4247 vdd.n1605 0.00239394
R15058 vdd.n1663 vdd.n1609 0.00239394
R15059 vdd.n4234 vdd.n1641 0.00239394
R15060 vdd.n4222 vdd.n4221 0.00239394
R15061 vdd.n4212 vdd.n1691 0.00239394
R15062 vdd.n4200 vdd.n4199 0.00239394
R15063 vdd.n4190 vdd.n1733 0.00239394
R15064 vdd.n4178 vdd.n4177 0.00239394
R15065 vdd.n4165 vdd.n1777 0.00239394
R15066 vdd.n4153 vdd.n1805 0.00239394
R15067 vdd.n1856 vdd.n1809 0.00239394
R15068 vdd.n1884 vdd.n1839 0.00239394
R15069 vdd.n4126 vdd.n1869 0.00239394
R15070 vdd.n1927 vdd.n1873 0.00239394
R15071 vdd.n4113 vdd.n1905 0.00239394
R15072 vdd.n4101 vdd.n4100 0.00239394
R15073 vdd.n4091 vdd.n1955 0.00239394
R15074 vdd.n4079 vdd.n4078 0.00239394
R15075 vdd.n4069 vdd.n1997 0.00239394
R15076 vdd.n4057 vdd.n4056 0.00239394
R15077 vdd.n896 vdd.n854 0.00239394
R15078 vdd.n4570 vdd.n4569 0.00239394
R15079 vdd.n938 vdd.n864 0.00239394
R15080 vdd.n4552 vdd.n921 0.00239394
R15081 vdd.n4543 vdd.n4542 0.00239394
R15082 vdd.n895 vdd.n894 0.00239394
R15083 vdd.n4568 vdd.n861 0.00239394
R15084 vdd.n937 vdd.n865 0.00239394
R15085 vdd.n965 vdd.n920 0.00239394
R15086 vdd.n4541 vdd.n950 0.00239394
R15087 vdd.n4681 vdd.n801 0.00239394
R15088 vdd.n4702 vdd.n789 0.00239394
R15089 vdd.n4715 vdd.n781 0.00239394
R15090 vdd.n4751 vdd.n773 0.00239394
R15091 vdd.n4763 vdd.n761 0.00239394
R15092 vdd.n4784 vdd.n736 0.00239394
R15093 vdd.n751 vdd.n730 0.00239394
R15094 vdd.n4803 vdd.n721 0.00239394
R15095 vdd.n4815 vdd.n710 0.00239394
R15096 vdd.n4846 vdd.n701 0.00239394
R15097 vdd.n4857 vdd.n687 0.00239394
R15098 vdd.n4871 vdd.n677 0.00239394
R15099 vdd.n4909 vdd.n666 0.00239394
R15100 vdd.n4930 vdd.n654 0.00239394
R15101 vdd.n4943 vdd.n646 0.00239394
R15102 vdd.n4979 vdd.n638 0.00239394
R15103 vdd.n4991 vdd.n626 0.00239394
R15104 vdd.n5012 vdd.n601 0.00239394
R15105 vdd.n616 vdd.n595 0.00239394
R15106 vdd.n5031 vdd.n586 0.00239394
R15107 vdd.n5043 vdd.n575 0.00239394
R15108 vdd.n5074 vdd.n566 0.00239394
R15109 vdd.n5085 vdd.n552 0.00239394
R15110 vdd.n5099 vdd.n542 0.00239394
R15111 vdd.n5137 vdd.n531 0.00239394
R15112 vdd.n5158 vdd.n519 0.00239394
R15113 vdd.n5171 vdd.n511 0.00239394
R15114 vdd.n5207 vdd.n503 0.00239394
R15115 vdd.n5219 vdd.n491 0.00239394
R15116 vdd.n5240 vdd.n466 0.00239394
R15117 vdd.n481 vdd.n460 0.00239394
R15118 vdd.n5259 vdd.n451 0.00239394
R15119 vdd.n5271 vdd.n440 0.00239394
R15120 vdd.n5302 vdd.n431 0.00239394
R15121 vdd.n5313 vdd.n417 0.00239394
R15122 vdd.n5327 vdd.n407 0.00239394
R15123 vdd.n5365 vdd.n396 0.00239394
R15124 vdd.n5386 vdd.n384 0.00239394
R15125 vdd.n5399 vdd.n376 0.00239394
R15126 vdd.n5435 vdd.n368 0.00239394
R15127 vdd.n5447 vdd.n356 0.00239394
R15128 vdd.n5467 vdd.n340 0.00239394
R15129 vdd.n5476 vdd.n335 0.00239394
R15130 vdd.n5498 vdd.n327 0.00239394
R15131 vdd.n315 vdd.n309 0.00239394
R15132 vdd.n5532 vdd.n300 0.00239394
R15133 vdd.n5544 vdd.n287 0.00239394
R15134 vdd.n292 vdd.n281 0.00239394
R15135 vdd.n2237 vdd.n2236 0.00232171
R15136 vdd.n3902 vdd.n3888 0.0021514
R15137 vdd.n2225 vdd.n2222 0.0021514
R15138 vdd.n7410 vdd.n7409 0.00213953
R15139 vdd.n5658 vdd.n5657 0.00213953
R15140 vdd.n4043 vdd.n2039 0.00213953
R15141 vdd.n877 vdd.n874 0.00213953
R15142 vdd.n2146 vdd.n2114 0.00198617
R15143 vdd.n201 vdd.n190 0.00196875
R15144 vdd.n208 vdd.n203 0.00196875
R15145 vdd.n7498 vdd.n7497 0.00196875
R15146 vdd.n3849 vdd.n3845 0.00196875
R15147 vdd.n3994 vdd.n3843 0.00196875
R15148 vdd.n4597 vdd.n4595 0.00196875
R15149 vdd.n4601 vdd.n4590 0.00196875
R15150 vdd.n4673 vdd.n4672 0.00196875
R15151 vdd.n5760 vdd.n5759 0.00196875
R15152 vdd.n7472 vdd.n7471 0.00196875
R15153 vdd.n6395 vdd.n6394 0.00196875
R15154 vdd vdd.n5735 0.00196114
R15155 vdd.n7418 vdd 0.00196114
R15156 vdd.n7413 vdd.n188 0.00192568
R15157 vdd.n7517 vdd.n188 0.00192568
R15158 vdd.n7452 vdd.n7451 0.00192033
R15159 vdd.n2150 vdd.n2149 0.00189328
R15160 vdd.n2149 vdd.n2114 0.0018004
R15161 vdd.n4634 vdd.n4633 0.00175893
R15162 vdd.n4668 vdd.n807 0.00175893
R15163 vdd.n4672 vdd.n807 0.00175893
R15164 vdd.n7449 vdd.n7448 0.00175893
R15165 vdd.n6390 vdd.n6388 0.00175893
R15166 vdd.n6394 vdd.n6388 0.00175893
R15167 vdd.n5738 vdd.n233 0.00172665
R15168 vdd.n7456 vdd.n234 0.00172665
R15169 vdd.n2210 vdd.n2209 0.00170192
R15170 vdd.n2154 vdd.n2107 0.00170192
R15171 vdd.n2202 vdd.n2110 0.00159739
R15172 vdd.n2148 vdd.n2147 0.00159739
R15173 vdd.n4 vdd.n3 0.00159739
R15174 vdd.n141 vdd.n140 0.00159739
R15175 vdd.n82 vdd.n81 0.00159739
R15176 vdd.n97 vdd.n96 0.00159739
R15177 vdd.n68 vdd.n67 0.00159739
R15178 vdd.n182 vdd.n181 0.00159739
R15179 vdd.n7528 vdd.n7527 0.00159739
R15180 vdd.n2218 vdd.n2097 0.00154724
R15181 vdd.n4661 vdd.n4660 0.00150714
R15182 vdd.n819 vdd.n818 0.00150714
R15183 vdd.n5805 vdd.n5787 0.00150714
R15184 vdd.n7441 vdd.n5778 0.00150714
R15185 vdd vdd.n7517 0.00130789
R15186 vdd.n2154 vdd.n2105 0.00130128
R15187 vdd.n5736 vdd 0.00123057
R15188 vdd vdd.n7417 0.00123057
R15189 vdd.n4668 vdd.n4667 0.00121339
R15190 vdd.n6390 vdd.n5781 0.00121339
R15191 vdd.n5746 vdd.n5738 0.00121017
R15192 vdd.n7456 vdd.n233 0.00121017
R15193 vdd.n6398 vdd.n6387 0.00119118
R15194 vdd.n6403 vdd.n6387 0.00119118
R15195 vdd.n6418 vdd.n6378 0.00119118
R15196 vdd.n6424 vdd.n6378 0.00119118
R15197 vdd.n6440 vdd.n6439 0.00119118
R15198 vdd.n6441 vdd.n6440 0.00119118
R15199 vdd.n6446 vdd.n6355 0.00119118
R15200 vdd.n6463 vdd.n6355 0.00119118
R15201 vdd.n6468 vdd.n6344 0.00119118
R15202 vdd.n6483 vdd.n6344 0.00119118
R15203 vdd.n6488 vdd.n6322 0.00119118
R15204 vdd.n6502 vdd.n6322 0.00119118
R15205 vdd.n6509 vdd.n6508 0.00119118
R15206 vdd.n6508 vdd.n6308 0.00119118
R15207 vdd.n6530 vdd.n6305 0.00119118
R15208 vdd.n6540 vdd.n6305 0.00119118
R15209 vdd.n6535 vdd.n6294 0.00119118
R15210 vdd.n6564 vdd.n6294 0.00119118
R15211 vdd.n6570 vdd.n6569 0.00119118
R15212 vdd.n6570 vdd.n6290 0.00119118
R15213 vdd.n6591 vdd.n6590 0.00119118
R15214 vdd.n6591 vdd.n6273 0.00119118
R15215 vdd.n6615 vdd.n6614 0.00119118
R15216 vdd.n6615 vdd.n6260 0.00119118
R15217 vdd.n6625 vdd.n6256 0.00119118
R15218 vdd.n6630 vdd.n6256 0.00119118
R15219 vdd.n6645 vdd.n6245 0.00119118
R15220 vdd.n6651 vdd.n6245 0.00119118
R15221 vdd.n6667 vdd.n6666 0.00119118
R15222 vdd.n6668 vdd.n6667 0.00119118
R15223 vdd.n6673 vdd.n6222 0.00119118
R15224 vdd.n6690 vdd.n6222 0.00119118
R15225 vdd.n6695 vdd.n6211 0.00119118
R15226 vdd.n6710 vdd.n6211 0.00119118
R15227 vdd.n6715 vdd.n6189 0.00119118
R15228 vdd.n6729 vdd.n6189 0.00119118
R15229 vdd.n6736 vdd.n6735 0.00119118
R15230 vdd.n6735 vdd.n6175 0.00119118
R15231 vdd.n6757 vdd.n6172 0.00119118
R15232 vdd.n6767 vdd.n6172 0.00119118
R15233 vdd.n6762 vdd.n6161 0.00119118
R15234 vdd.n6791 vdd.n6161 0.00119118
R15235 vdd.n6797 vdd.n6796 0.00119118
R15236 vdd.n6797 vdd.n6157 0.00119118
R15237 vdd.n6818 vdd.n6817 0.00119118
R15238 vdd.n6818 vdd.n6140 0.00119118
R15239 vdd.n6842 vdd.n6841 0.00119118
R15240 vdd.n6842 vdd.n6127 0.00119118
R15241 vdd.n6852 vdd.n6123 0.00119118
R15242 vdd.n6857 vdd.n6123 0.00119118
R15243 vdd.n6872 vdd.n6112 0.00119118
R15244 vdd.n6878 vdd.n6112 0.00119118
R15245 vdd.n6894 vdd.n6893 0.00119118
R15246 vdd.n6895 vdd.n6894 0.00119118
R15247 vdd.n6900 vdd.n6089 0.00119118
R15248 vdd.n6917 vdd.n6089 0.00119118
R15249 vdd.n6922 vdd.n6078 0.00119118
R15250 vdd.n6937 vdd.n6078 0.00119118
R15251 vdd.n6942 vdd.n6056 0.00119118
R15252 vdd.n6956 vdd.n6056 0.00119118
R15253 vdd.n6963 vdd.n6962 0.00119118
R15254 vdd.n6962 vdd.n6042 0.00119118
R15255 vdd.n6984 vdd.n6039 0.00119118
R15256 vdd.n6994 vdd.n6039 0.00119118
R15257 vdd.n6989 vdd.n6028 0.00119118
R15258 vdd.n7018 vdd.n6028 0.00119118
R15259 vdd.n7024 vdd.n7023 0.00119118
R15260 vdd.n7024 vdd.n6024 0.00119118
R15261 vdd.n7045 vdd.n7044 0.00119118
R15262 vdd.n7045 vdd.n6007 0.00119118
R15263 vdd.n7069 vdd.n7068 0.00119118
R15264 vdd.n7069 vdd.n5994 0.00119118
R15265 vdd.n7079 vdd.n5990 0.00119118
R15266 vdd.n7084 vdd.n5990 0.00119118
R15267 vdd.n7099 vdd.n5979 0.00119118
R15268 vdd.n7105 vdd.n5979 0.00119118
R15269 vdd.n7121 vdd.n7120 0.00119118
R15270 vdd.n7122 vdd.n7121 0.00119118
R15271 vdd.n7127 vdd.n5956 0.00119118
R15272 vdd.n7144 vdd.n5956 0.00119118
R15273 vdd.n7149 vdd.n5945 0.00119118
R15274 vdd.n7164 vdd.n5945 0.00119118
R15275 vdd.n7169 vdd.n5923 0.00119118
R15276 vdd.n7183 vdd.n5923 0.00119118
R15277 vdd.n7190 vdd.n7189 0.00119118
R15278 vdd.n7189 vdd.n5909 0.00119118
R15279 vdd.n7211 vdd.n5906 0.00119118
R15280 vdd.n7221 vdd.n5906 0.00119118
R15281 vdd.n7216 vdd.n5895 0.00119118
R15282 vdd.n7245 vdd.n5895 0.00119118
R15283 vdd.n7251 vdd.n7250 0.00119118
R15284 vdd.n7251 vdd.n5891 0.00119118
R15285 vdd.n7272 vdd.n7271 0.00119118
R15286 vdd.n7272 vdd.n5873 0.00119118
R15287 vdd.n7276 vdd.n7275 0.00119118
R15288 vdd.n7276 vdd.n5864 0.00119118
R15289 vdd.n7306 vdd.n7305 0.00119118
R15290 vdd.n7306 vdd.n5862 0.00119118
R15291 vdd.n7325 vdd.n7324 0.00119118
R15292 vdd.n7325 vdd.n5851 0.00119118
R15293 vdd.n7344 vdd.n7343 0.00119118
R15294 vdd.n7344 vdd.n5840 0.00119118
R15295 vdd.n7363 vdd.n7362 0.00119118
R15296 vdd.n7363 vdd.n5829 0.00119118
R15297 vdd.n7382 vdd.n7381 0.00119118
R15298 vdd.n7382 vdd.n5817 0.00119118
R15299 vdd.n7386 vdd.n5797 0.00119118
R15300 vdd.n7386 vdd.n5795 0.00119118
R15301 vdd.n4676 vdd.n805 0.00119118
R15302 vdd.n4682 vdd.n805 0.00119118
R15303 vdd.n4687 vdd.n794 0.00119118
R15304 vdd.n4703 vdd.n794 0.00119118
R15305 vdd.n4717 vdd.n792 0.00119118
R15306 vdd.n4713 vdd.n792 0.00119118
R15307 vdd.n4740 vdd.n4739 0.00119118
R15308 vdd.n4741 vdd.n4740 0.00119118
R15309 vdd.n4746 vdd.n765 0.00119118
R15310 vdd.n4764 vdd.n765 0.00119118
R15311 vdd.n4770 vdd.n734 0.00119118
R15312 vdd.n4785 vdd.n734 0.00119118
R15313 vdd.n4787 vdd.n731 0.00119118
R15314 vdd.n4797 vdd.n731 0.00119118
R15315 vdd.n4792 vdd.n720 0.00119118
R15316 vdd.n4821 vdd.n720 0.00119118
R15317 vdd.n4827 vdd.n4826 0.00119118
R15318 vdd.n4827 vdd.n716 0.00119118
R15319 vdd.n4848 vdd.n4847 0.00119118
R15320 vdd.n4848 vdd.n696 0.00119118
R15321 vdd.n697 vdd.n686 0.00119118
R15322 vdd.n4877 vdd.n686 0.00119118
R15323 vdd.n4883 vdd.n4882 0.00119118
R15324 vdd.n4883 vdd.n681 0.00119118
R15325 vdd.n4887 vdd.n670 0.00119118
R15326 vdd.n4910 vdd.n670 0.00119118
R15327 vdd.n4915 vdd.n659 0.00119118
R15328 vdd.n4931 vdd.n659 0.00119118
R15329 vdd.n4945 vdd.n657 0.00119118
R15330 vdd.n4941 vdd.n657 0.00119118
R15331 vdd.n4968 vdd.n4967 0.00119118
R15332 vdd.n4969 vdd.n4968 0.00119118
R15333 vdd.n4974 vdd.n630 0.00119118
R15334 vdd.n4992 vdd.n630 0.00119118
R15335 vdd.n4998 vdd.n599 0.00119118
R15336 vdd.n5013 vdd.n599 0.00119118
R15337 vdd.n5015 vdd.n596 0.00119118
R15338 vdd.n5025 vdd.n596 0.00119118
R15339 vdd.n5020 vdd.n585 0.00119118
R15340 vdd.n5049 vdd.n585 0.00119118
R15341 vdd.n5055 vdd.n5054 0.00119118
R15342 vdd.n5055 vdd.n581 0.00119118
R15343 vdd.n5076 vdd.n5075 0.00119118
R15344 vdd.n5076 vdd.n561 0.00119118
R15345 vdd.n562 vdd.n551 0.00119118
R15346 vdd.n5105 vdd.n551 0.00119118
R15347 vdd.n5111 vdd.n5110 0.00119118
R15348 vdd.n5111 vdd.n546 0.00119118
R15349 vdd.n5115 vdd.n535 0.00119118
R15350 vdd.n5138 vdd.n535 0.00119118
R15351 vdd.n5143 vdd.n524 0.00119118
R15352 vdd.n5159 vdd.n524 0.00119118
R15353 vdd.n5173 vdd.n522 0.00119118
R15354 vdd.n5169 vdd.n522 0.00119118
R15355 vdd.n5196 vdd.n5195 0.00119118
R15356 vdd.n5197 vdd.n5196 0.00119118
R15357 vdd.n5202 vdd.n495 0.00119118
R15358 vdd.n5220 vdd.n495 0.00119118
R15359 vdd.n5226 vdd.n464 0.00119118
R15360 vdd.n5241 vdd.n464 0.00119118
R15361 vdd.n5243 vdd.n461 0.00119118
R15362 vdd.n5253 vdd.n461 0.00119118
R15363 vdd.n5248 vdd.n450 0.00119118
R15364 vdd.n5277 vdd.n450 0.00119118
R15365 vdd.n5283 vdd.n5282 0.00119118
R15366 vdd.n5283 vdd.n446 0.00119118
R15367 vdd.n5304 vdd.n5303 0.00119118
R15368 vdd.n5304 vdd.n426 0.00119118
R15369 vdd.n427 vdd.n416 0.00119118
R15370 vdd.n5333 vdd.n416 0.00119118
R15371 vdd.n5339 vdd.n5338 0.00119118
R15372 vdd.n5339 vdd.n411 0.00119118
R15373 vdd.n5343 vdd.n400 0.00119118
R15374 vdd.n5366 vdd.n400 0.00119118
R15375 vdd.n5371 vdd.n389 0.00119118
R15376 vdd.n5387 vdd.n389 0.00119118
R15377 vdd.n5401 vdd.n387 0.00119118
R15378 vdd.n5397 vdd.n387 0.00119118
R15379 vdd.n5424 vdd.n5423 0.00119118
R15380 vdd.n5425 vdd.n5424 0.00119118
R15381 vdd.n5430 vdd.n360 0.00119118
R15382 vdd.n5448 vdd.n360 0.00119118
R15383 vdd.n5453 vdd.n338 0.00119118
R15384 vdd.n5468 vdd.n338 0.00119118
R15385 vdd.n5474 vdd.n5473 0.00119118
R15386 vdd.n5473 vdd.n330 0.00119118
R15387 vdd.n5496 vdd.n5495 0.00119118
R15388 vdd.n5495 vdd.n313 0.00119118
R15389 vdd.n5516 vdd.n310 0.00119118
R15390 vdd.n5526 vdd.n310 0.00119118
R15391 vdd.n5521 vdd.n299 0.00119118
R15392 vdd.n5550 vdd.n299 0.00119118
R15393 vdd.n5556 vdd.n5555 0.00119118
R15394 vdd.n5556 vdd.n294 0.00119118
R15395 vdd.n5560 vdd.n5559 0.00119118
R15396 vdd.n5560 vdd.n278 0.00119118
R15397 vdd.n5584 vdd.n276 0.00119118
R15398 vdd.n5594 vdd.n276 0.00119118
R15399 vdd.n5600 vdd.n5599 0.00119118
R15400 vdd.n5600 vdd.n271 0.00119118
R15401 vdd.n5710 vdd.n5604 0.00119118
R15402 vdd.n5710 vdd.n5709 0.00119118
R15403 vdd.n5638 vdd.n5632 0.00119118
R15404 vdd.n5639 vdd.n5638 0.00119118
R15405 vdd.n5690 vdd.n5689 0.00119118
R15406 vdd.n5689 vdd.n5630 0.00119118
R15407 vdd.n5683 vdd.n5650 0.00119118
R15408 vdd.n5662 vdd.n5650 0.00119118
R15409 vdd.n2902 vdd.n2781 0.00119118
R15410 vdd.n2908 vdd.n2781 0.00119118
R15411 vdd.n2913 vdd.n2770 0.00119118
R15412 vdd.n2929 vdd.n2770 0.00119118
R15413 vdd.n2943 vdd.n2768 0.00119118
R15414 vdd.n2939 vdd.n2768 0.00119118
R15415 vdd.n2966 vdd.n2965 0.00119118
R15416 vdd.n2967 vdd.n2966 0.00119118
R15417 vdd.n2972 vdd.n2741 0.00119118
R15418 vdd.n2990 vdd.n2741 0.00119118
R15419 vdd.n2996 vdd.n2710 0.00119118
R15420 vdd.n3011 vdd.n2710 0.00119118
R15421 vdd.n3013 vdd.n2707 0.00119118
R15422 vdd.n3023 vdd.n2707 0.00119118
R15423 vdd.n3018 vdd.n2696 0.00119118
R15424 vdd.n3047 vdd.n2696 0.00119118
R15425 vdd.n3053 vdd.n3052 0.00119118
R15426 vdd.n3053 vdd.n2692 0.00119118
R15427 vdd.n3074 vdd.n3073 0.00119118
R15428 vdd.n3074 vdd.n2672 0.00119118
R15429 vdd.n2673 vdd.n2662 0.00119118
R15430 vdd.n3103 vdd.n2662 0.00119118
R15431 vdd.n3109 vdd.n3108 0.00119118
R15432 vdd.n3109 vdd.n2657 0.00119118
R15433 vdd.n3113 vdd.n2646 0.00119118
R15434 vdd.n3136 vdd.n2646 0.00119118
R15435 vdd.n3141 vdd.n2635 0.00119118
R15436 vdd.n3157 vdd.n2635 0.00119118
R15437 vdd.n3171 vdd.n2633 0.00119118
R15438 vdd.n3167 vdd.n2633 0.00119118
R15439 vdd.n3194 vdd.n3193 0.00119118
R15440 vdd.n3195 vdd.n3194 0.00119118
R15441 vdd.n3200 vdd.n2606 0.00119118
R15442 vdd.n3218 vdd.n2606 0.00119118
R15443 vdd.n3224 vdd.n2575 0.00119118
R15444 vdd.n3239 vdd.n2575 0.00119118
R15445 vdd.n3241 vdd.n2572 0.00119118
R15446 vdd.n3251 vdd.n2572 0.00119118
R15447 vdd.n3246 vdd.n2561 0.00119118
R15448 vdd.n3275 vdd.n2561 0.00119118
R15449 vdd.n3281 vdd.n3280 0.00119118
R15450 vdd.n3281 vdd.n2557 0.00119118
R15451 vdd.n3302 vdd.n3301 0.00119118
R15452 vdd.n3302 vdd.n2537 0.00119118
R15453 vdd.n2538 vdd.n2527 0.00119118
R15454 vdd.n3331 vdd.n2527 0.00119118
R15455 vdd.n3337 vdd.n3336 0.00119118
R15456 vdd.n3337 vdd.n2522 0.00119118
R15457 vdd.n3341 vdd.n2511 0.00119118
R15458 vdd.n3364 vdd.n2511 0.00119118
R15459 vdd.n3369 vdd.n2500 0.00119118
R15460 vdd.n3385 vdd.n2500 0.00119118
R15461 vdd.n3399 vdd.n2498 0.00119118
R15462 vdd.n3395 vdd.n2498 0.00119118
R15463 vdd.n3422 vdd.n3421 0.00119118
R15464 vdd.n3423 vdd.n3422 0.00119118
R15465 vdd.n3428 vdd.n2471 0.00119118
R15466 vdd.n3446 vdd.n2471 0.00119118
R15467 vdd.n3452 vdd.n2440 0.00119118
R15468 vdd.n3467 vdd.n2440 0.00119118
R15469 vdd.n3469 vdd.n2437 0.00119118
R15470 vdd.n3479 vdd.n2437 0.00119118
R15471 vdd.n3474 vdd.n2426 0.00119118
R15472 vdd.n3503 vdd.n2426 0.00119118
R15473 vdd.n3509 vdd.n3508 0.00119118
R15474 vdd.n3509 vdd.n2422 0.00119118
R15475 vdd.n3530 vdd.n3529 0.00119118
R15476 vdd.n3530 vdd.n2402 0.00119118
R15477 vdd.n2403 vdd.n2392 0.00119118
R15478 vdd.n3559 vdd.n2392 0.00119118
R15479 vdd.n3565 vdd.n3564 0.00119118
R15480 vdd.n3565 vdd.n2387 0.00119118
R15481 vdd.n3569 vdd.n2376 0.00119118
R15482 vdd.n3592 vdd.n2376 0.00119118
R15483 vdd.n3597 vdd.n2365 0.00119118
R15484 vdd.n3613 vdd.n2365 0.00119118
R15485 vdd.n3627 vdd.n2363 0.00119118
R15486 vdd.n3623 vdd.n2363 0.00119118
R15487 vdd.n3650 vdd.n3649 0.00119118
R15488 vdd.n3651 vdd.n3650 0.00119118
R15489 vdd.n3656 vdd.n2336 0.00119118
R15490 vdd.n3674 vdd.n2336 0.00119118
R15491 vdd.n3679 vdd.n2314 0.00119118
R15492 vdd.n3694 vdd.n2314 0.00119118
R15493 vdd.n3700 vdd.n3699 0.00119118
R15494 vdd.n3699 vdd.n2305 0.00119118
R15495 vdd.n3721 vdd.n3720 0.00119118
R15496 vdd.n3720 vdd.n2287 0.00119118
R15497 vdd.n3740 vdd.n2284 0.00119118
R15498 vdd.n3750 vdd.n2284 0.00119118
R15499 vdd.n3745 vdd.n2273 0.00119118
R15500 vdd.n3774 vdd.n2273 0.00119118
R15501 vdd.n3780 vdd.n3779 0.00119118
R15502 vdd.n3780 vdd.n2268 0.00119118
R15503 vdd.n3784 vdd.n3783 0.00119118
R15504 vdd.n3784 vdd.n2252 0.00119118
R15505 vdd.n4039 vdd.n2042 0.00119118
R15506 vdd.n2047 vdd.n2042 0.00119118
R15507 vdd.n2819 vdd.n2048 0.00119118
R15508 vdd.n2820 vdd.n2819 0.00119118
R15509 vdd.n2835 vdd.n2834 0.00119118
R15510 vdd.n2836 vdd.n2835 0.00119118
R15511 vdd.n2841 vdd.n2802 0.00119118
R15512 vdd.n2859 vdd.n2802 0.00119118
R15513 vdd.n2864 vdd.n2791 0.00119118
R15514 vdd.n2886 vdd.n2791 0.00119118
R15515 vdd.n2891 vdd.n2784 0.00119118
R15516 vdd.n2898 vdd.n2784 0.00119118
R15517 vdd.n1020 vdd.n984 0.00119118
R15518 vdd.n1021 vdd.n1020 0.00119118
R15519 vdd.n1036 vdd.n1017 0.00119118
R15520 vdd.n1037 vdd.n1036 0.00119118
R15521 vdd.n4510 vdd.n1015 0.00119118
R15522 vdd.n1042 vdd.n1015 0.00119118
R15523 vdd.n1089 vdd.n1043 0.00119118
R15524 vdd.n1090 vdd.n1089 0.00119118
R15525 vdd.n1105 vdd.n1085 0.00119118
R15526 vdd.n1106 vdd.n1105 0.00119118
R15527 vdd.n4483 vdd.n1083 0.00119118
R15528 vdd.n1111 vdd.n1083 0.00119118
R15529 vdd.n4477 vdd.n1112 0.00119118
R15530 vdd.n1153 vdd.n1112 0.00119118
R15531 vdd.n4462 vdd.n4461 0.00119118
R15532 vdd.n4461 vdd.n1150 0.00119118
R15533 vdd.n4455 vdd.n1162 0.00119118
R15534 vdd.n1195 vdd.n1162 0.00119118
R15535 vdd.n4440 vdd.n4439 0.00119118
R15536 vdd.n4439 vdd.n1192 0.00119118
R15537 vdd.n4433 vdd.n1204 0.00119118
R15538 vdd.n1237 vdd.n1204 0.00119118
R15539 vdd.n4418 vdd.n4417 0.00119118
R15540 vdd.n4417 vdd.n1234 0.00119118
R15541 vdd.n4409 vdd.n1247 0.00119118
R15542 vdd.n1250 vdd.n1247 0.00119118
R15543 vdd.n1300 vdd.n1285 0.00119118
R15544 vdd.n1301 vdd.n1300 0.00119118
R15545 vdd.n4389 vdd.n1283 0.00119118
R15546 vdd.n1306 vdd.n1283 0.00119118
R15547 vdd.n1353 vdd.n1307 0.00119118
R15548 vdd.n1354 vdd.n1353 0.00119118
R15549 vdd.n1369 vdd.n1349 0.00119118
R15550 vdd.n1370 vdd.n1369 0.00119118
R15551 vdd.n4362 vdd.n1347 0.00119118
R15552 vdd.n1375 vdd.n1347 0.00119118
R15553 vdd.n4356 vdd.n1376 0.00119118
R15554 vdd.n1417 vdd.n1376 0.00119118
R15555 vdd.n4341 vdd.n4340 0.00119118
R15556 vdd.n4340 vdd.n1414 0.00119118
R15557 vdd.n4334 vdd.n1426 0.00119118
R15558 vdd.n1459 vdd.n1426 0.00119118
R15559 vdd.n4319 vdd.n4318 0.00119118
R15560 vdd.n4318 vdd.n1456 0.00119118
R15561 vdd.n4312 vdd.n1468 0.00119118
R15562 vdd.n1501 vdd.n1468 0.00119118
R15563 vdd.n4297 vdd.n4296 0.00119118
R15564 vdd.n4296 vdd.n1498 0.00119118
R15565 vdd.n4288 vdd.n1511 0.00119118
R15566 vdd.n1514 vdd.n1511 0.00119118
R15567 vdd.n1564 vdd.n1549 0.00119118
R15568 vdd.n1565 vdd.n1564 0.00119118
R15569 vdd.n4268 vdd.n1547 0.00119118
R15570 vdd.n1570 vdd.n1547 0.00119118
R15571 vdd.n1617 vdd.n1571 0.00119118
R15572 vdd.n1618 vdd.n1617 0.00119118
R15573 vdd.n1633 vdd.n1613 0.00119118
R15574 vdd.n1634 vdd.n1633 0.00119118
R15575 vdd.n4241 vdd.n1611 0.00119118
R15576 vdd.n1639 vdd.n1611 0.00119118
R15577 vdd.n4235 vdd.n1640 0.00119118
R15578 vdd.n1681 vdd.n1640 0.00119118
R15579 vdd.n4220 vdd.n4219 0.00119118
R15580 vdd.n4219 vdd.n1678 0.00119118
R15581 vdd.n4213 vdd.n1690 0.00119118
R15582 vdd.n1723 vdd.n1690 0.00119118
R15583 vdd.n4198 vdd.n4197 0.00119118
R15584 vdd.n4197 vdd.n1720 0.00119118
R15585 vdd.n4191 vdd.n1732 0.00119118
R15586 vdd.n1765 vdd.n1732 0.00119118
R15587 vdd.n4176 vdd.n4175 0.00119118
R15588 vdd.n4175 vdd.n1762 0.00119118
R15589 vdd.n4167 vdd.n1775 0.00119118
R15590 vdd.n1778 vdd.n1775 0.00119118
R15591 vdd.n1828 vdd.n1813 0.00119118
R15592 vdd.n1829 vdd.n1828 0.00119118
R15593 vdd.n4147 vdd.n1811 0.00119118
R15594 vdd.n1834 vdd.n1811 0.00119118
R15595 vdd.n1881 vdd.n1835 0.00119118
R15596 vdd.n1882 vdd.n1881 0.00119118
R15597 vdd.n1897 vdd.n1877 0.00119118
R15598 vdd.n1898 vdd.n1897 0.00119118
R15599 vdd.n4120 vdd.n1875 0.00119118
R15600 vdd.n1903 vdd.n1875 0.00119118
R15601 vdd.n4114 vdd.n1904 0.00119118
R15602 vdd.n1945 vdd.n1904 0.00119118
R15603 vdd.n4099 vdd.n4098 0.00119118
R15604 vdd.n4098 vdd.n1942 0.00119118
R15605 vdd.n4092 vdd.n1954 0.00119118
R15606 vdd.n1987 vdd.n1954 0.00119118
R15607 vdd.n4077 vdd.n4076 0.00119118
R15608 vdd.n4076 vdd.n1984 0.00119118
R15609 vdd.n4070 vdd.n1996 0.00119118
R15610 vdd.n2029 vdd.n1996 0.00119118
R15611 vdd.n4055 vdd.n4054 0.00119118
R15612 vdd.n4054 vdd.n2026 0.00119118
R15613 vdd.n892 vdd.n873 0.00119118
R15614 vdd.n893 vdd.n892 0.00119118
R15615 vdd.n909 vdd.n869 0.00119118
R15616 vdd.n910 vdd.n909 0.00119118
R15617 vdd.n4562 vdd.n867 0.00119118
R15618 vdd.n915 vdd.n867 0.00119118
R15619 vdd.n962 vdd.n916 0.00119118
R15620 vdd.n963 vdd.n962 0.00119118
R15621 vdd.n978 vdd.n958 0.00119118
R15622 vdd.n979 vdd.n978 0.00119118
R15623 vdd.n4535 vdd.n956 0.00119118
R15624 vdd.n4531 vdd.n956 0.00119118
R15625 vdd.n2219 vdd.n2095 0.00113087
R15626 vdd.n2124 vdd.n2122 0.0011215
R15627 vdd.n3895 vdd.n3893 0.0011215
R15628 vdd.n832 vdd.n830 0.0011215
R15629 vdd.n5767 vdd.n5765 0.0011215
R15630 vdd.n3993 vdd.n3842 0.00111039
R15631 vdd.n4600 vdd.n4592 0.00111039
R15632 vdd.n2161 vdd.n2110 0.00107317
R15633 vdd.n2097 vdd.n2094 0.00107317
R15634 vdd.n2140 vdd.n2119 0.00107317
R15635 vdd.n2140 vdd.n2133 0.00107317
R15636 vdd.n2152 vdd.n2151 0.00107317
R15637 vdd.n2152 vdd.n2112 0.00107317
R15638 vdd.n2186 vdd.n2165 0.00107317
R15639 vdd.n2186 vdd.n2185 0.00107317
R15640 vdd.n2147 vdd.n2116 0.00107317
R15641 vdd.n3 vdd.n2 0.00107317
R15642 vdd.n142 vdd.n141 0.00107317
R15643 vdd.n81 vdd.n80 0.00107317
R15644 vdd.n96 vdd.n95 0.00107317
R15645 vdd.n67 vdd.n66 0.00107317
R15646 vdd.n183 vdd.n182 0.00107317
R15647 vdd.n7527 vdd.n7526 0.00107317
R15648 vdd.n7452 vdd.n5762 0.00101648
R15649 vdd.n4674 vdd 0.000994737
R15650 vdd vdd.n4889 0.000994737
R15651 vdd vdd.n5117 0.000994737
R15652 vdd vdd.n5345 0.000994737
R15653 vdd.n6396 vdd 0.000994737
R15654 vdd vdd.n6257 0.000994737
R15655 vdd vdd.n6124 0.000994737
R15656 vdd vdd.n5991 0.000994737
R15657 vdd vdd.n4530 0.000989583
R15658 vdd.n4411 vdd 0.000989583
R15659 vdd.n4290 vdd 0.000989583
R15660 vdd.n4169 vdd 0.000989583
R15661 vdd.n2900 vdd 0.000989583
R15662 vdd vdd.n3115 0.000989583
R15663 vdd vdd.n3343 0.000989583
R15664 vdd vdd.n3571 0.000989583
R15665 vdd.n889 vdd 0.000982051
R15666 vdd.n2045 vdd 0.000982051
R15667 vdd.n3990 vdd.n3842 0.000837321
R15668 vdd.n4592 vdd.n839 0.000837321
R15669 vdd.n2144 vdd.n2143 0.000815436
R15670 vdd vdd.n206 0.000815436
R15671 vdd.n4675 vdd.n804 0.000747368
R15672 vdd.n4686 vdd.n793 0.000747368
R15673 vdd.n4709 vdd.n4707 0.000747368
R15674 vdd.n780 vdd.n778 0.000747368
R15675 vdd.n4745 vdd.n764 0.000747368
R15676 vdd.n4769 vdd.n4768 0.000747368
R15677 vdd.n4796 vdd.n4790 0.000747368
R15678 vdd.n4822 vdd.n719 0.000747368
R15679 vdd.n4829 vdd.n4828 0.000747368
R15680 vdd.n4850 vdd.n4849 0.000747368
R15681 vdd.n4878 vdd.n685 0.000747368
R15682 vdd.n4885 vdd.n4884 0.000747368
R15683 vdd.n4888 vdd.n669 0.000747368
R15684 vdd.n4914 vdd.n658 0.000747368
R15685 vdd.n4937 vdd.n4935 0.000747368
R15686 vdd.n645 vdd.n643 0.000747368
R15687 vdd.n4973 vdd.n629 0.000747368
R15688 vdd.n4997 vdd.n4996 0.000747368
R15689 vdd.n5024 vdd.n5018 0.000747368
R15690 vdd.n5050 vdd.n584 0.000747368
R15691 vdd.n5057 vdd.n5056 0.000747368
R15692 vdd.n5078 vdd.n5077 0.000747368
R15693 vdd.n5106 vdd.n550 0.000747368
R15694 vdd.n5113 vdd.n5112 0.000747368
R15695 vdd.n5116 vdd.n534 0.000747368
R15696 vdd.n5142 vdd.n523 0.000747368
R15697 vdd.n5165 vdd.n5163 0.000747368
R15698 vdd.n510 vdd.n508 0.000747368
R15699 vdd.n5201 vdd.n494 0.000747368
R15700 vdd.n5225 vdd.n5224 0.000747368
R15701 vdd.n5252 vdd.n5246 0.000747368
R15702 vdd.n5278 vdd.n449 0.000747368
R15703 vdd.n5285 vdd.n5284 0.000747368
R15704 vdd.n5306 vdd.n5305 0.000747368
R15705 vdd.n5334 vdd.n415 0.000747368
R15706 vdd.n5341 vdd.n5340 0.000747368
R15707 vdd.n5344 vdd.n399 0.000747368
R15708 vdd.n5370 vdd.n388 0.000747368
R15709 vdd.n5393 vdd.n5391 0.000747368
R15710 vdd.n375 vdd.n373 0.000747368
R15711 vdd.n5429 vdd.n359 0.000747368
R15712 vdd.n5452 vdd.n337 0.000747368
R15713 vdd.n5472 vdd.n329 0.000747368
R15714 vdd.n5494 vdd.n5493 0.000747368
R15715 vdd.n5525 vdd.n5519 0.000747368
R15716 vdd.n5551 vdd.n298 0.000747368
R15717 vdd.n5558 vdd.n5557 0.000747368
R15718 vdd.n5561 vdd.n277 0.000747368
R15719 vdd.n6400 vdd.n6399 0.000747368
R15720 vdd.n6420 vdd.n6419 0.000747368
R15721 vdd.n6370 vdd.n6368 0.000747368
R15722 vdd.n6445 vdd.n6354 0.000747368
R15723 vdd.n6467 vdd.n6343 0.000747368
R15724 vdd.n6487 vdd.n6321 0.000747368
R15725 vdd.n6507 vdd.n6506 0.000747368
R15726 vdd.n6539 vdd.n6533 0.000747368
R15727 vdd.n6565 vdd.n6293 0.000747368
R15728 vdd.n6572 vdd.n6571 0.000747368
R15729 vdd.n6593 vdd.n6592 0.000747368
R15730 vdd.n6617 vdd.n6616 0.000747368
R15731 vdd.n6627 vdd.n6626 0.000747368
R15732 vdd.n6647 vdd.n6646 0.000747368
R15733 vdd.n6237 vdd.n6235 0.000747368
R15734 vdd.n6672 vdd.n6221 0.000747368
R15735 vdd.n6694 vdd.n6210 0.000747368
R15736 vdd.n6714 vdd.n6188 0.000747368
R15737 vdd.n6734 vdd.n6733 0.000747368
R15738 vdd.n6766 vdd.n6760 0.000747368
R15739 vdd.n6792 vdd.n6160 0.000747368
R15740 vdd.n6799 vdd.n6798 0.000747368
R15741 vdd.n6820 vdd.n6819 0.000747368
R15742 vdd.n6844 vdd.n6843 0.000747368
R15743 vdd.n6854 vdd.n6853 0.000747368
R15744 vdd.n6874 vdd.n6873 0.000747368
R15745 vdd.n6104 vdd.n6102 0.000747368
R15746 vdd.n6899 vdd.n6088 0.000747368
R15747 vdd.n6921 vdd.n6077 0.000747368
R15748 vdd.n6941 vdd.n6055 0.000747368
R15749 vdd.n6961 vdd.n6960 0.000747368
R15750 vdd.n6993 vdd.n6987 0.000747368
R15751 vdd.n7019 vdd.n6027 0.000747368
R15752 vdd.n7026 vdd.n7025 0.000747368
R15753 vdd.n7047 vdd.n7046 0.000747368
R15754 vdd.n7071 vdd.n7070 0.000747368
R15755 vdd.n7081 vdd.n7080 0.000747368
R15756 vdd.n7101 vdd.n7100 0.000747368
R15757 vdd.n5971 vdd.n5969 0.000747368
R15758 vdd.n7126 vdd.n5955 0.000747368
R15759 vdd.n7148 vdd.n5944 0.000747368
R15760 vdd.n7168 vdd.n5922 0.000747368
R15761 vdd.n7188 vdd.n7187 0.000747368
R15762 vdd.n7220 vdd.n7214 0.000747368
R15763 vdd.n7246 vdd.n5894 0.000747368
R15764 vdd.n7253 vdd.n7252 0.000747368
R15765 vdd.n7274 vdd.n7273 0.000747368
R15766 vdd.n7277 vdd.n5863 0.000747368
R15767 vdd.n5582 vdd.n5581 0.000744792
R15768 vdd.n1019 vdd.n983 0.000744792
R15769 vdd.n1035 vdd.n1034 0.000744792
R15770 vdd.n4509 vdd.n4508 0.000744792
R15771 vdd.n1088 vdd.n1087 0.000744792
R15772 vdd.n1104 vdd.n1103 0.000744792
R15773 vdd.n4482 vdd.n4481 0.000744792
R15774 vdd.n1152 vdd.n1151 0.000744792
R15775 vdd.n4460 vdd.n4459 0.000744792
R15776 vdd.n1194 vdd.n1193 0.000744792
R15777 vdd.n4438 vdd.n4437 0.000744792
R15778 vdd.n1236 vdd.n1235 0.000744792
R15779 vdd.n4416 vdd.n4415 0.000744792
R15780 vdd.n4410 vdd.n1246 0.000744792
R15781 vdd.n1299 vdd.n1298 0.000744792
R15782 vdd.n4388 vdd.n4387 0.000744792
R15783 vdd.n1352 vdd.n1351 0.000744792
R15784 vdd.n1368 vdd.n1367 0.000744792
R15785 vdd.n4361 vdd.n4360 0.000744792
R15786 vdd.n1416 vdd.n1415 0.000744792
R15787 vdd.n4339 vdd.n4338 0.000744792
R15788 vdd.n1458 vdd.n1457 0.000744792
R15789 vdd.n4317 vdd.n4316 0.000744792
R15790 vdd.n1500 vdd.n1499 0.000744792
R15791 vdd.n4295 vdd.n4294 0.000744792
R15792 vdd.n4289 vdd.n1510 0.000744792
R15793 vdd.n1563 vdd.n1562 0.000744792
R15794 vdd.n4267 vdd.n4266 0.000744792
R15795 vdd.n1616 vdd.n1615 0.000744792
R15796 vdd.n1632 vdd.n1631 0.000744792
R15797 vdd.n4240 vdd.n4239 0.000744792
R15798 vdd.n1680 vdd.n1679 0.000744792
R15799 vdd.n4218 vdd.n4217 0.000744792
R15800 vdd.n1722 vdd.n1721 0.000744792
R15801 vdd.n4196 vdd.n4195 0.000744792
R15802 vdd.n1764 vdd.n1763 0.000744792
R15803 vdd.n4174 vdd.n4173 0.000744792
R15804 vdd.n4168 vdd.n1774 0.000744792
R15805 vdd.n1827 vdd.n1826 0.000744792
R15806 vdd.n4146 vdd.n4145 0.000744792
R15807 vdd.n1880 vdd.n1879 0.000744792
R15808 vdd.n1896 vdd.n1895 0.000744792
R15809 vdd.n4119 vdd.n4118 0.000744792
R15810 vdd.n1944 vdd.n1943 0.000744792
R15811 vdd.n4097 vdd.n4096 0.000744792
R15812 vdd.n1986 vdd.n1985 0.000744792
R15813 vdd.n4075 vdd.n4074 0.000744792
R15814 vdd.n2028 vdd.n2027 0.000744792
R15815 vdd.n4053 vdd.n4052 0.000744792
R15816 vdd.n2901 vdd.n2780 0.000744792
R15817 vdd.n2912 vdd.n2769 0.000744792
R15818 vdd.n2935 vdd.n2933 0.000744792
R15819 vdd.n2756 vdd.n2754 0.000744792
R15820 vdd.n2971 vdd.n2740 0.000744792
R15821 vdd.n2995 vdd.n2994 0.000744792
R15822 vdd.n3022 vdd.n3016 0.000744792
R15823 vdd.n3048 vdd.n2695 0.000744792
R15824 vdd.n3055 vdd.n3054 0.000744792
R15825 vdd.n3076 vdd.n3075 0.000744792
R15826 vdd.n3104 vdd.n2661 0.000744792
R15827 vdd.n3111 vdd.n3110 0.000744792
R15828 vdd.n3114 vdd.n2645 0.000744792
R15829 vdd.n3140 vdd.n2634 0.000744792
R15830 vdd.n3163 vdd.n3161 0.000744792
R15831 vdd.n2621 vdd.n2619 0.000744792
R15832 vdd.n3199 vdd.n2605 0.000744792
R15833 vdd.n3223 vdd.n3222 0.000744792
R15834 vdd.n3250 vdd.n3244 0.000744792
R15835 vdd.n3276 vdd.n2560 0.000744792
R15836 vdd.n3283 vdd.n3282 0.000744792
R15837 vdd.n3304 vdd.n3303 0.000744792
R15838 vdd.n3332 vdd.n2526 0.000744792
R15839 vdd.n3339 vdd.n3338 0.000744792
R15840 vdd.n3342 vdd.n2510 0.000744792
R15841 vdd.n3368 vdd.n2499 0.000744792
R15842 vdd.n3391 vdd.n3389 0.000744792
R15843 vdd.n2486 vdd.n2484 0.000744792
R15844 vdd.n3427 vdd.n2470 0.000744792
R15845 vdd.n3451 vdd.n3450 0.000744792
R15846 vdd.n3478 vdd.n3472 0.000744792
R15847 vdd.n3504 vdd.n2425 0.000744792
R15848 vdd.n3511 vdd.n3510 0.000744792
R15849 vdd.n3532 vdd.n3531 0.000744792
R15850 vdd.n3560 vdd.n2391 0.000744792
R15851 vdd.n3567 vdd.n3566 0.000744792
R15852 vdd.n3570 vdd.n2375 0.000744792
R15853 vdd.n3596 vdd.n2364 0.000744792
R15854 vdd.n3619 vdd.n3617 0.000744792
R15855 vdd.n2351 vdd.n2349 0.000744792
R15856 vdd.n3655 vdd.n2335 0.000744792
R15857 vdd.n3678 vdd.n2313 0.000744792
R15858 vdd.n3698 vdd.n2304 0.000744792
R15859 vdd.n3719 vdd.n3718 0.000744792
R15860 vdd.n3749 vdd.n3743 0.000744792
R15861 vdd.n3775 vdd.n2272 0.000744792
R15862 vdd.n3782 vdd.n3781 0.000744792
R15863 vdd.n3785 vdd.n2251 0.000744792
R15864 vdd.n7297 vdd.n7296 0.000744792
R15865 vdd.n5595 vdd.n275 0.000743523
R15866 vdd.n5602 vdd.n5601 0.000743523
R15867 vdd.n5711 vdd.n5603 0.000743523
R15868 vdd.n5637 vdd.n5631 0.000743523
R15869 vdd.n5688 vdd.n5687 0.000743523
R15870 vdd.n5661 vdd.n5655 0.000743523
R15871 vdd.n7308 vdd.n7307 0.000743523
R15872 vdd.n7327 vdd.n7326 0.000743523
R15873 vdd.n7346 vdd.n7345 0.000743523
R15874 vdd.n7365 vdd.n7364 0.000743523
R15875 vdd.n7384 vdd.n7383 0.000743523
R15876 vdd.n7387 vdd.n7385 0.000743523
R15877 vdd.n891 vdd.n890 0.000741026
R15878 vdd.n908 vdd.n907 0.000741026
R15879 vdd.n4561 vdd.n4560 0.000741026
R15880 vdd.n961 vdd.n960 0.000741026
R15881 vdd.n977 vdd.n976 0.000741026
R15882 vdd.n4534 vdd.n4533 0.000741026
R15883 vdd.n4038 vdd.n4037 0.000741026
R15884 vdd.n2818 vdd.n2817 0.000741026
R15885 vdd.n2824 vdd.n2814 0.000741026
R15886 vdd.n2840 vdd.n2801 0.000741026
R15887 vdd.n2863 vdd.n2790 0.000741026
R15888 vdd.n2890 vdd.n2783 0.000741026
R15889 vdd.n4661 vdd.n813 0.000709821
R15890 vdd.n818 vdd.n814 0.000709821
R15891 vdd.n4667 vdd.n809 0.000709821
R15892 vdd.n5805 vdd.n5774 0.000709821
R15893 vdd.n7430 vdd.n5778 0.000709821
R15894 vdd.n7440 vdd.n5781 0.000709821
R15895 vdd.n5762 vdd.n234 0.000693681
R15896 vdd.n206 vdd.n205 0.000657718
R15897 vdd.n7496 vdd.n202 0.000657718
R15898 vdd.n3990 vdd.n3989 0.00061244
R15899 vdd.n4631 vdd.n839 0.00061244
R15900 vdd.n117 vdd.n116 0.000595528
R15901 vdd.n121 vdd.n120 0.000595528
R15902 vdd.n125 vdd.n124 0.000595528
R15903 vdd.n144 vdd.n143 0.000595528
R15904 vdd.n185 vdd.n184 0.000595528
R15905 vdd.n7525 vdd.n7524 0.000595528
R15906 vdd.n7521 vdd.n7520 0.000595528
R15907 vdd.n2146 vdd.n2145 0.000592885
R15908 vdd.n2150 vdd.n2111 0.000592885
R15909 vdd.n2163 vdd.n2162 0.000592885
R15910 vdd.n2187 vdd.n2164 0.000592885
R15911 vdd.n4635 vdd.n813 0.000541964
R15912 vdd.n4660 vdd.n814 0.000541964
R15913 vdd.n819 vdd.n809 0.000541964
R15914 vdd.n7447 vdd.n5774 0.000541964
R15915 vdd.n7430 vdd.n5787 0.000541964
R15916 vdd.n7441 vdd.n7440 0.000541964
R15917 x2.x1.x10.Y x2.x1.x10.Y.t7 154.847
R15918 x2.x1.x10.Y x2.x1.x10.Y.t9 154.8
R15919 x2.x1.x10.Y x2.x1.x10.Y.t2 154.8
R15920 x2.x1.x10.Y x2.x1.x10.Y.t3 154.8
R15921 x2.x1.x10.Y x2.x1.x10.Y.t4 154.8
R15922 x2.x1.x10.Y x2.x1.x10.Y.t5 154.8
R15923 x2.x1.x10.Y x2.x1.x10.Y.t6 154.8
R15924 x2.x1.x10.Y x2.x1.x10.Y.t8 154.8
R15925 x2.x1.x10.Y.n0 x2.x1.x10.Y 134.239
R15926 x2.x1.x10.Y x2.x1.x10.Y.t1 106.635
R15927 x2.x1.x10.Y.n2 x2.x1.x10.Y.t0 24.6567
R15928 x2.x1.x10.Y.n5 x2.x1.x10.Y.n4 12.4089
R15929 x2.x1.x10.Y.n3 x2.x1.x10.Y.n2 9.12522
R15930 x2.x1.x10.Y.n4 x2.x1.x10.Y.n3 7.34048
R15931 x2.x1.x10.Y.n5 x2.x1.x10.Y 2.22659
R15932 x2.x1.x10.Y.n2 x2.x1.x10.Y.n1 1.93377
R15933 x2.x1.x10.Y x2.x1.x10.Y.n5 1.55202
R15934 x2.x1.x10.Y.n3 x2.x1.x10.Y.n0 0.69928
R15935 x2.x1.x5[7].floating.n154 x2.x1.x5[7].floating.t1 68.0345
R15936 x2.x1.x5[7].floating.n142 x2.x1.x5[7].floating.t3 68.0345
R15937 x2.x1.x5[7].floating.n12 x2.x1.x5[7].floating.t4 68.0345
R15938 x2.x1.x5[7].floating.n24 x2.x1.x5[7].floating.t5 68.0345
R15939 x2.x1.x5[7].floating.n54 x2.x1.x5[7].floating.t7 68.0345
R15940 x2.x1.x5[7].floating.n72 x2.x1.x5[7].floating.t0 68.0345
R15941 x2.x1.x5[7].floating.n84 x2.x1.x5[7].floating.t2 68.0345
R15942 x2.x1.x5[7].floating.n42 x2.x1.x5[7].floating.t6 68.0345
R15943 x2.x1.x5[7].floating.n103 x2.x1.x5[7].floating.n65 0.660401
R15944 x2.x1.x5[7].floating.n112 x2.x1.x5[7].floating.n50 0.660401
R15945 x2.x1.x5[7].floating.n121 x2.x1.x5[7].floating.n35 0.660401
R15946 x2.x1.x5[7].floating.n130 x2.x1.x5[7].floating.n20 0.660401
R15947 x2.x1.x5[7].floating.n139 x2.x1.x5[7].floating.n5 0.660401
R15948 x2.x1.x5[7].floating.n90 x2.x1.x5[7].floating.n89 0.320345
R15949 x2.x1.x5[7].floating.n160 x2.x1.x5[7].floating.n159 0.308269
R15950 x2.x1.x5[7].floating.n161 x2.x1.x5[7].floating.n160 0.173084
R15951 x2.x1.x5[7].floating.n91 x2.x1.x5[7].floating.n90 0.162103
R15952 x2.x1.x5[7].floating.n160 x2.x1.x5[7].floating 0.100688
R15953 x2.x1.x5[7].floating.n90 x2.x1.x5[7].floating 0.0755007
R15954 x2.x1.x5[7].floating.n66 x2.x1.x5[7].floating.n65 0.0716912
R15955 x2.x1.x5[7].floating.n65 x2.x1.x5[7].floating.n64 0.0716912
R15956 x2.x1.x5[7].floating.n36 x2.x1.x5[7].floating.n35 0.0716912
R15957 x2.x1.x5[7].floating.n35 x2.x1.x5[7].floating.n34 0.0716912
R15958 x2.x1.x5[7].floating.n6 x2.x1.x5[7].floating.n5 0.0716912
R15959 x2.x1.x5[7].floating.n5 x2.x1.x5[7].floating.n4 0.0716912
R15960 x2.x1.x5[7].floating.n104 x2.x1.x5[7].floating.n103 0.0716912
R15961 x2.x1.x5[7].floating.n122 x2.x1.x5[7].floating.n121 0.0716912
R15962 x2.x1.x5[7].floating.n140 x2.x1.x5[7].floating.n139 0.0716912
R15963 x2.x1.x5[7].floating.n70 x2.x1.x5[7].floating.n69 0.0557941
R15964 x2.x1.x5[7].floating.n69 x2.x1.x5[7].floating.n68 0.0557941
R15965 x2.x1.x5[7].floating.n68 x2.x1.x5[7].floating.n67 0.0557941
R15966 x2.x1.x5[7].floating.n67 x2.x1.x5[7].floating.n66 0.0557941
R15967 x2.x1.x5[7].floating.n64 x2.x1.x5[7].floating.n63 0.0557941
R15968 x2.x1.x5[7].floating.n63 x2.x1.x5[7].floating.n62 0.0557941
R15969 x2.x1.x5[7].floating.n62 x2.x1.x5[7].floating.n61 0.0557941
R15970 x2.x1.x5[7].floating.n61 x2.x1.x5[7].floating.n60 0.0557941
R15971 x2.x1.x5[7].floating.n40 x2.x1.x5[7].floating.n39 0.0557941
R15972 x2.x1.x5[7].floating.n39 x2.x1.x5[7].floating.n38 0.0557941
R15973 x2.x1.x5[7].floating.n38 x2.x1.x5[7].floating.n37 0.0557941
R15974 x2.x1.x5[7].floating.n37 x2.x1.x5[7].floating.n36 0.0557941
R15975 x2.x1.x5[7].floating.n34 x2.x1.x5[7].floating.n33 0.0557941
R15976 x2.x1.x5[7].floating.n33 x2.x1.x5[7].floating.n32 0.0557941
R15977 x2.x1.x5[7].floating.n32 x2.x1.x5[7].floating.n31 0.0557941
R15978 x2.x1.x5[7].floating.n31 x2.x1.x5[7].floating.n30 0.0557941
R15979 x2.x1.x5[7].floating.n10 x2.x1.x5[7].floating.n9 0.0557941
R15980 x2.x1.x5[7].floating.n9 x2.x1.x5[7].floating.n8 0.0557941
R15981 x2.x1.x5[7].floating.n8 x2.x1.x5[7].floating.n7 0.0557941
R15982 x2.x1.x5[7].floating.n7 x2.x1.x5[7].floating.n6 0.0557941
R15983 x2.x1.x5[7].floating.n4 x2.x1.x5[7].floating.n3 0.0557941
R15984 x2.x1.x5[7].floating.n3 x2.x1.x5[7].floating.n2 0.0557941
R15985 x2.x1.x5[7].floating.n2 x2.x1.x5[7].floating.n1 0.0557941
R15986 x2.x1.x5[7].floating.n1 x2.x1.x5[7].floating.n0 0.0557941
R15987 x2.x1.x5[7].floating.n99 x2.x1.x5[7].floating.n98 0.0557941
R15988 x2.x1.x5[7].floating.n100 x2.x1.x5[7].floating.n99 0.0557941
R15989 x2.x1.x5[7].floating.n101 x2.x1.x5[7].floating.n100 0.0557941
R15990 x2.x1.x5[7].floating.n102 x2.x1.x5[7].floating.n101 0.0557941
R15991 x2.x1.x5[7].floating.n106 x2.x1.x5[7].floating.n105 0.0557941
R15992 x2.x1.x5[7].floating.n107 x2.x1.x5[7].floating.n106 0.0557941
R15993 x2.x1.x5[7].floating.n108 x2.x1.x5[7].floating.n107 0.0557941
R15994 x2.x1.x5[7].floating.n117 x2.x1.x5[7].floating.n116 0.0557941
R15995 x2.x1.x5[7].floating.n118 x2.x1.x5[7].floating.n117 0.0557941
R15996 x2.x1.x5[7].floating.n119 x2.x1.x5[7].floating.n118 0.0557941
R15997 x2.x1.x5[7].floating.n120 x2.x1.x5[7].floating.n119 0.0557941
R15998 x2.x1.x5[7].floating.n124 x2.x1.x5[7].floating.n123 0.0557941
R15999 x2.x1.x5[7].floating.n125 x2.x1.x5[7].floating.n124 0.0557941
R16000 x2.x1.x5[7].floating.n126 x2.x1.x5[7].floating.n125 0.0557941
R16001 x2.x1.x5[7].floating.n135 x2.x1.x5[7].floating.n134 0.0557941
R16002 x2.x1.x5[7].floating.n136 x2.x1.x5[7].floating.n135 0.0557941
R16003 x2.x1.x5[7].floating.n137 x2.x1.x5[7].floating.n136 0.0557941
R16004 x2.x1.x5[7].floating.n138 x2.x1.x5[7].floating.n137 0.0557941
R16005 x2.x1.x5[7].floating.n171 x2.x1.x5[7].floating.n170 0.0557941
R16006 x2.x1.x5[7].floating.n170 x2.x1.x5[7].floating.n169 0.0557941
R16007 x2.x1.x5[7].floating.n169 x2.x1.x5[7].floating.n168 0.0557941
R16008 x2.x1.x5[7].floating.n95 x2.x1.x5[7].floating.n94 0.0537206
R16009 x2.x1.x5[7].floating.n113 x2.x1.x5[7].floating.n112 0.0537206
R16010 x2.x1.x5[7].floating.n131 x2.x1.x5[7].floating.n130 0.0537206
R16011 x2.x1.x5[7].floating.n164 x2.x1.x5[7].floating.n163 0.0537206
R16012 x2.x1.x5[7].floating.n94 x2.x1.x5[7].floating.n93 0.0530294
R16013 x2.x1.x5[7].floating.n112 x2.x1.x5[7].floating.n111 0.0530294
R16014 x2.x1.x5[7].floating.n130 x2.x1.x5[7].floating.n129 0.0530294
R16015 x2.x1.x5[7].floating.n165 x2.x1.x5[7].floating.n164 0.0530294
R16016 x2.x1.x5[7].floating.n80 x2.x1.x5[7].floating.n79 0.0529559
R16017 x2.x1.x5[7].floating.n50 x2.x1.x5[7].floating.n49 0.0529559
R16018 x2.x1.x5[7].floating.n20 x2.x1.x5[7].floating.n19 0.0529559
R16019 x2.x1.x5[7].floating.n151 x2.x1.x5[7].floating.n150 0.0529559
R16020 x2.x1.x5[7].floating.n81 x2.x1.x5[7].floating.n80 0.0524559
R16021 x2.x1.x5[7].floating.n51 x2.x1.x5[7].floating.n50 0.0524559
R16022 x2.x1.x5[7].floating.n21 x2.x1.x5[7].floating.n20 0.0524559
R16023 x2.x1.x5[7].floating.n150 x2.x1.x5[7].floating.n149 0.0524559
R16024 x2.x1.x5[7].floating.n109 x2.x1.x5[7].floating.n108 0.0523382
R16025 x2.x1.x5[7].floating.n127 x2.x1.x5[7].floating.n126 0.0523382
R16026 x2.x1.x5[7].floating.n168 x2.x1.x5[7].floating.n167 0.0523382
R16027 x2.x1.x5[7].floating.n98 x2.x1.x5[7].floating.n97 0.0516471
R16028 x2.x1.x5[7].floating.n116 x2.x1.x5[7].floating.n115 0.0516471
R16029 x2.x1.x5[7].floating.n134 x2.x1.x5[7].floating.n133 0.0516471
R16030 x2.x1.x5[7].floating.n103 x2.x1.x5[7].floating 0.0495735
R16031 x2.x1.x5[7].floating.n121 x2.x1.x5[7].floating 0.0495735
R16032 x2.x1.x5[7].floating.n139 x2.x1.x5[7].floating 0.0495735
R16033 x2.x1.x5[7].floating.n157 x2.x1.x5[7].floating.n156 0.0408846
R16034 x2.x1.x5[7].floating.n15 x2.x1.x5[7].floating.n14 0.0408846
R16035 x2.x1.x5[7].floating.n75 x2.x1.x5[7].floating.n74 0.0408846
R16036 x2.x1.x5[7].floating.n45 x2.x1.x5[7].floating.n44 0.0408846
R16037 x2.x1.x5[7].floating.n105 x2.x1.x5[7].floating 0.0336765
R16038 x2.x1.x5[7].floating.n123 x2.x1.x5[7].floating 0.0336765
R16039 x2.x1.x5[7].floating x2.x1.x5[7].floating.n171 0.0336765
R16040 x2.x1.x5[7].floating.n60 x2.x1.x5[7].floating.n59 0.0271618
R16041 x2.x1.x5[7].floating.n30 x2.x1.x5[7].floating.n29 0.0271618
R16042 x2.x1.x5[7].floating.n71 x2.x1.x5[7].floating.n70 0.0266618
R16043 x2.x1.x5[7].floating.n41 x2.x1.x5[7].floating.n40 0.0266618
R16044 x2.x1.x5[7].floating.n11 x2.x1.x5[7].floating.n10 0.0266618
R16045 x2.x1.x5[7].floating x2.x1.x5[7].floating.n102 0.0226176
R16046 x2.x1.x5[7].floating x2.x1.x5[7].floating.n104 0.0226176
R16047 x2.x1.x5[7].floating x2.x1.x5[7].floating.n120 0.0226176
R16048 x2.x1.x5[7].floating x2.x1.x5[7].floating.n122 0.0226176
R16049 x2.x1.x5[7].floating x2.x1.x5[7].floating.n138 0.0226176
R16050 x2.x1.x5[7].floating x2.x1.x5[7].floating.n140 0.0226176
R16051 x2.x1.x5[7].floating.n93 x2.x1.x5[7].floating.n92 0.0191618
R16052 x2.x1.x5[7].floating.n111 x2.x1.x5[7].floating.n110 0.0191618
R16053 x2.x1.x5[7].floating.n129 x2.x1.x5[7].floating.n128 0.0191618
R16054 x2.x1.x5[7].floating.n166 x2.x1.x5[7].floating.n165 0.0191618
R16055 x2.x1.x5[7].floating.n96 x2.x1.x5[7].floating.n95 0.0184706
R16056 x2.x1.x5[7].floating.n114 x2.x1.x5[7].floating.n113 0.0184706
R16057 x2.x1.x5[7].floating.n132 x2.x1.x5[7].floating.n131 0.0184706
R16058 x2.x1.x5[7].floating.n163 x2.x1.x5[7].floating.n162 0.0184706
R16059 x2.x1.x5[7].floating.n82 x2.x1.x5[7].floating.n81 0.014
R16060 x2.x1.x5[7].floating.n76 x2.x1.x5[7].floating.n71 0.014
R16061 x2.x1.x5[7].floating.n52 x2.x1.x5[7].floating.n51 0.014
R16062 x2.x1.x5[7].floating.n46 x2.x1.x5[7].floating.n41 0.014
R16063 x2.x1.x5[7].floating.n22 x2.x1.x5[7].floating.n21 0.014
R16064 x2.x1.x5[7].floating.n16 x2.x1.x5[7].floating.n11 0.014
R16065 x2.x1.x5[7].floating.n149 x2.x1.x5[7].floating.n148 0.014
R16066 x2.x1.x5[7].floating.n159 x2.x1.x5[7].floating.n158 0.014
R16067 x2.x1.x5[7].floating.n89 x2.x1.x5[7].floating.n88 0.0135
R16068 x2.x1.x5[7].floating.n79 x2.x1.x5[7].floating.n78 0.0135
R16069 x2.x1.x5[7].floating.n59 x2.x1.x5[7].floating.n58 0.0135
R16070 x2.x1.x5[7].floating.n49 x2.x1.x5[7].floating.n48 0.0135
R16071 x2.x1.x5[7].floating.n29 x2.x1.x5[7].floating.n28 0.0135
R16072 x2.x1.x5[7].floating.n19 x2.x1.x5[7].floating.n18 0.0135
R16073 x2.x1.x5[7].floating.n146 x2.x1.x5[7].floating.n141 0.0135
R16074 x2.x1.x5[7].floating.n152 x2.x1.x5[7].floating.n151 0.0135
R16075 x2.x1.x5[7].floating.n145 x2.x1.x5[7].floating.n144 0.0120385
R16076 x2.x1.x5[7].floating.n27 x2.x1.x5[7].floating.n26 0.0120385
R16077 x2.x1.x5[7].floating.n57 x2.x1.x5[7].floating.n56 0.0120385
R16078 x2.x1.x5[7].floating.n87 x2.x1.x5[7].floating.n86 0.0120385
R16079 x2.x1.x5[7].floating.n97 x2.x1.x5[7].floating.n96 0.00464706
R16080 x2.x1.x5[7].floating.n115 x2.x1.x5[7].floating.n114 0.00464706
R16081 x2.x1.x5[7].floating.n133 x2.x1.x5[7].floating.n132 0.00464706
R16082 x2.x1.x5[7].floating.n162 x2.x1.x5[7].floating.n161 0.00464706
R16083 x2.x1.x5[7].floating.n92 x2.x1.x5[7].floating.n91 0.00395588
R16084 x2.x1.x5[7].floating.n110 x2.x1.x5[7].floating.n109 0.00395588
R16085 x2.x1.x5[7].floating.n128 x2.x1.x5[7].floating.n127 0.00395588
R16086 x2.x1.x5[7].floating.n167 x2.x1.x5[7].floating.n166 0.00395588
R16087 x2.x1.x5[7].floating.n143 x2.x1.x5[7].floating.n142 0.00359614
R16088 x2.x1.x5[7].floating.n25 x2.x1.x5[7].floating.n24 0.00359614
R16089 x2.x1.x5[7].floating.n55 x2.x1.x5[7].floating.n54 0.00359614
R16090 x2.x1.x5[7].floating.n85 x2.x1.x5[7].floating.n84 0.00359614
R16091 x2.x1.x5[7].floating.n88 x2.x1.x5[7].floating.n83 0.0035
R16092 x2.x1.x5[7].floating.n78 x2.x1.x5[7].floating.n77 0.0035
R16093 x2.x1.x5[7].floating.n58 x2.x1.x5[7].floating.n53 0.0035
R16094 x2.x1.x5[7].floating.n48 x2.x1.x5[7].floating.n47 0.0035
R16095 x2.x1.x5[7].floating.n28 x2.x1.x5[7].floating.n23 0.0035
R16096 x2.x1.x5[7].floating.n18 x2.x1.x5[7].floating.n17 0.0035
R16097 x2.x1.x5[7].floating.n147 x2.x1.x5[7].floating.n146 0.0035
R16098 x2.x1.x5[7].floating.n153 x2.x1.x5[7].floating.n152 0.0035
R16099 x2.x1.x5[7].floating.n83 x2.x1.x5[7].floating.n82 0.003
R16100 x2.x1.x5[7].floating.n77 x2.x1.x5[7].floating.n76 0.003
R16101 x2.x1.x5[7].floating.n53 x2.x1.x5[7].floating.n52 0.003
R16102 x2.x1.x5[7].floating.n47 x2.x1.x5[7].floating.n46 0.003
R16103 x2.x1.x5[7].floating.n23 x2.x1.x5[7].floating.n22 0.003
R16104 x2.x1.x5[7].floating.n17 x2.x1.x5[7].floating.n16 0.003
R16105 x2.x1.x5[7].floating.n148 x2.x1.x5[7].floating.n147 0.003
R16106 x2.x1.x5[7].floating.n158 x2.x1.x5[7].floating.n153 0.003
R16107 x2.x1.x5[7].floating.n155 x2.x1.x5[7].floating.n154 0.00277942
R16108 x2.x1.x5[7].floating.n43 x2.x1.x5[7].floating.n42 0.0023396
R16109 x2.x1.x5[7].floating.n13 x2.x1.x5[7].floating.n12 0.0023396
R16110 x2.x1.x5[7].floating.n73 x2.x1.x5[7].floating.n72 0.0023396
R16111 x2.x1.x5[7].floating.n157 x2.x1.x5[7].floating.n155 0.00233747
R16112 x2.x1.x5[7].floating.n15 x2.x1.x5[7].floating.n13 0.00200689
R16113 x2.x1.x5[7].floating.n75 x2.x1.x5[7].floating.n73 0.00200689
R16114 x2.x1.x5[7].floating.n45 x2.x1.x5[7].floating.n43 0.00200689
R16115 x2.x1.x5[7].floating.n145 x2.x1.x5[7].floating.n143 0.0010233
R16116 x2.x1.x5[7].floating.n27 x2.x1.x5[7].floating.n25 0.0010233
R16117 x2.x1.x5[7].floating.n57 x2.x1.x5[7].floating.n55 0.0010233
R16118 x2.x1.x5[7].floating.n87 x2.x1.x5[7].floating.n85 0.0010233
R16119 x2.x1.x5[7].floating.n88 x2.x1.x5[7].floating.n87 0.00053972
R16120 x2.x1.x5[7].floating.n76 x2.x1.x5[7].floating.n75 0.00053972
R16121 x2.x1.x5[7].floating.n58 x2.x1.x5[7].floating.n57 0.00053972
R16122 x2.x1.x5[7].floating.n28 x2.x1.x5[7].floating.n27 0.00053972
R16123 x2.x1.x5[7].floating.n16 x2.x1.x5[7].floating.n15 0.00053972
R16124 x2.x1.x5[7].floating.n146 x2.x1.x5[7].floating.n145 0.00053972
R16125 x2.x1.x5[7].floating.n158 x2.x1.x5[7].floating.n157 0.00053972
R16126 x2.x1.x5[7].floating.n46 x2.x1.x5[7].floating.n45 0.00053972
R16127 x2.x4.x10.Y x2.x4.x10.Y.t8 154.847
R16128 x2.x4.x10.Y x2.x4.x10.Y.t9 154.8
R16129 x2.x4.x10.Y x2.x4.x10.Y.t3 154.8
R16130 x2.x4.x10.Y x2.x4.x10.Y.t4 154.8
R16131 x2.x4.x10.Y x2.x4.x10.Y.t5 154.8
R16132 x2.x4.x10.Y x2.x4.x10.Y.t6 154.8
R16133 x2.x4.x10.Y x2.x4.x10.Y.t7 154.8
R16134 x2.x4.x10.Y x2.x4.x10.Y.t2 154.8
R16135 x2.x4.x10.Y.n0 x2.x4.x10.Y 134.239
R16136 x2.x4.x10.Y x2.x4.x10.Y.t0 106.635
R16137 x2.x4.x10.Y.n2 x2.x4.x10.Y.t1 24.6567
R16138 x2.x4.x10.Y.n5 x2.x4.x10.Y.n4 12.4089
R16139 x2.x4.x10.Y.n3 x2.x4.x10.Y.n2 9.12522
R16140 x2.x4.x10.Y.n4 x2.x4.x10.Y.n3 7.34048
R16141 x2.x4.x10.Y.n5 x2.x4.x10.Y 2.22659
R16142 x2.x4.x10.Y.n2 x2.x4.x10.Y.n1 1.93377
R16143 x2.x4.x10.Y x2.x4.x10.Y.n5 1.55202
R16144 x2.x4.x10.Y.n3 x2.x4.x10.Y.n0 0.69928
R16145 x2.x4.x5[7].floating.n77 x2.x4.x5[7].floating.t0 68.0345
R16146 x2.x4.x5[7].floating.n65 x2.x4.x5[7].floating.t1 68.0345
R16147 x2.x4.x5[7].floating.n154 x2.x4.x5[7].floating.t7 68.0345
R16148 x2.x4.x5[7].floating.n142 x2.x4.x5[7].floating.t2 68.0345
R16149 x2.x4.x5[7].floating.n12 x2.x4.x5[7].floating.t3 68.0345
R16150 x2.x4.x5[7].floating.n24 x2.x4.x5[7].floating.t4 68.0345
R16151 x2.x4.x5[7].floating.n42 x2.x4.x5[7].floating.t5 68.0345
R16152 x2.x4.x5[7].floating.n91 x2.x4.x5[7].floating.t6 68.0345
R16153 x2.x4.x5[7].floating.n112 x2.x4.x5[7].floating.n50 0.660401
R16154 x2.x4.x5[7].floating.n121 x2.x4.x5[7].floating.n35 0.660401
R16155 x2.x4.x5[7].floating.n130 x2.x4.x5[7].floating.n20 0.660401
R16156 x2.x4.x5[7].floating.n139 x2.x4.x5[7].floating.n5 0.660401
R16157 x2.x4.x5[7].floating.n103 x2.x4.x5[7].floating.n102 0.660401
R16158 x2.x4.x5[7].floating.n64 x2.x4.x5[7].floating.n63 0.320345
R16159 x2.x4.x5[7].floating.n160 x2.x4.x5[7].floating.n159 0.308269
R16160 x2.x4.x5[7].floating.n161 x2.x4.x5[7].floating.n160 0.173084
R16161 x2.x4.x5[7].floating.n63 x2.x4.x5[7].floating.n62 0.162103
R16162 x2.x4.x5[7].floating.n160 x2.x4.x5[7].floating 0.100688
R16163 x2.x4.x5[7].floating.n63 x2.x4.x5[7].floating 0.0755007
R16164 x2.x4.x5[7].floating.n36 x2.x4.x5[7].floating.n35 0.0716912
R16165 x2.x4.x5[7].floating.n35 x2.x4.x5[7].floating.n34 0.0716912
R16166 x2.x4.x5[7].floating.n6 x2.x4.x5[7].floating.n5 0.0716912
R16167 x2.x4.x5[7].floating.n5 x2.x4.x5[7].floating.n4 0.0716912
R16168 x2.x4.x5[7].floating.n104 x2.x4.x5[7].floating.n103 0.0716912
R16169 x2.x4.x5[7].floating.n122 x2.x4.x5[7].floating.n121 0.0716912
R16170 x2.x4.x5[7].floating.n140 x2.x4.x5[7].floating.n139 0.0716912
R16171 x2.x4.x5[7].floating.n102 x2.x4.x5[7].floating.n87 0.0716912
R16172 x2.x4.x5[7].floating.n102 x2.x4.x5[7].floating.n101 0.0716912
R16173 x2.x4.x5[7].floating.n40 x2.x4.x5[7].floating.n39 0.0557941
R16174 x2.x4.x5[7].floating.n39 x2.x4.x5[7].floating.n38 0.0557941
R16175 x2.x4.x5[7].floating.n38 x2.x4.x5[7].floating.n37 0.0557941
R16176 x2.x4.x5[7].floating.n37 x2.x4.x5[7].floating.n36 0.0557941
R16177 x2.x4.x5[7].floating.n34 x2.x4.x5[7].floating.n33 0.0557941
R16178 x2.x4.x5[7].floating.n33 x2.x4.x5[7].floating.n32 0.0557941
R16179 x2.x4.x5[7].floating.n32 x2.x4.x5[7].floating.n31 0.0557941
R16180 x2.x4.x5[7].floating.n31 x2.x4.x5[7].floating.n30 0.0557941
R16181 x2.x4.x5[7].floating.n10 x2.x4.x5[7].floating.n9 0.0557941
R16182 x2.x4.x5[7].floating.n9 x2.x4.x5[7].floating.n8 0.0557941
R16183 x2.x4.x5[7].floating.n8 x2.x4.x5[7].floating.n7 0.0557941
R16184 x2.x4.x5[7].floating.n7 x2.x4.x5[7].floating.n6 0.0557941
R16185 x2.x4.x5[7].floating.n4 x2.x4.x5[7].floating.n3 0.0557941
R16186 x2.x4.x5[7].floating.n3 x2.x4.x5[7].floating.n2 0.0557941
R16187 x2.x4.x5[7].floating.n2 x2.x4.x5[7].floating.n1 0.0557941
R16188 x2.x4.x5[7].floating.n1 x2.x4.x5[7].floating.n0 0.0557941
R16189 x2.x4.x5[7].floating.n55 x2.x4.x5[7].floating.n54 0.0557941
R16190 x2.x4.x5[7].floating.n54 x2.x4.x5[7].floating.n53 0.0557941
R16191 x2.x4.x5[7].floating.n53 x2.x4.x5[7].floating.n52 0.0557941
R16192 x2.x4.x5[7].floating.n52 x2.x4.x5[7].floating.n51 0.0557941
R16193 x2.x4.x5[7].floating.n106 x2.x4.x5[7].floating.n105 0.0557941
R16194 x2.x4.x5[7].floating.n107 x2.x4.x5[7].floating.n106 0.0557941
R16195 x2.x4.x5[7].floating.n108 x2.x4.x5[7].floating.n107 0.0557941
R16196 x2.x4.x5[7].floating.n117 x2.x4.x5[7].floating.n116 0.0557941
R16197 x2.x4.x5[7].floating.n118 x2.x4.x5[7].floating.n117 0.0557941
R16198 x2.x4.x5[7].floating.n119 x2.x4.x5[7].floating.n118 0.0557941
R16199 x2.x4.x5[7].floating.n120 x2.x4.x5[7].floating.n119 0.0557941
R16200 x2.x4.x5[7].floating.n124 x2.x4.x5[7].floating.n123 0.0557941
R16201 x2.x4.x5[7].floating.n125 x2.x4.x5[7].floating.n124 0.0557941
R16202 x2.x4.x5[7].floating.n126 x2.x4.x5[7].floating.n125 0.0557941
R16203 x2.x4.x5[7].floating.n135 x2.x4.x5[7].floating.n134 0.0557941
R16204 x2.x4.x5[7].floating.n136 x2.x4.x5[7].floating.n135 0.0557941
R16205 x2.x4.x5[7].floating.n137 x2.x4.x5[7].floating.n136 0.0557941
R16206 x2.x4.x5[7].floating.n138 x2.x4.x5[7].floating.n137 0.0557941
R16207 x2.x4.x5[7].floating.n171 x2.x4.x5[7].floating.n170 0.0557941
R16208 x2.x4.x5[7].floating.n170 x2.x4.x5[7].floating.n169 0.0557941
R16209 x2.x4.x5[7].floating.n169 x2.x4.x5[7].floating.n168 0.0557941
R16210 x2.x4.x5[7].floating.n84 x2.x4.x5[7].floating.n83 0.0557941
R16211 x2.x4.x5[7].floating.n85 x2.x4.x5[7].floating.n84 0.0557941
R16212 x2.x4.x5[7].floating.n86 x2.x4.x5[7].floating.n85 0.0557941
R16213 x2.x4.x5[7].floating.n87 x2.x4.x5[7].floating.n86 0.0557941
R16214 x2.x4.x5[7].floating.n101 x2.x4.x5[7].floating.n100 0.0557941
R16215 x2.x4.x5[7].floating.n100 x2.x4.x5[7].floating.n99 0.0557941
R16216 x2.x4.x5[7].floating.n99 x2.x4.x5[7].floating.n98 0.0557941
R16217 x2.x4.x5[7].floating.n98 x2.x4.x5[7].floating.n97 0.0557941
R16218 x2.x4.x5[7].floating.n59 x2.x4.x5[7].floating.n58 0.0537206
R16219 x2.x4.x5[7].floating.n113 x2.x4.x5[7].floating.n112 0.0537206
R16220 x2.x4.x5[7].floating.n131 x2.x4.x5[7].floating.n130 0.0537206
R16221 x2.x4.x5[7].floating.n164 x2.x4.x5[7].floating.n163 0.0537206
R16222 x2.x4.x5[7].floating.n60 x2.x4.x5[7].floating.n59 0.0530294
R16223 x2.x4.x5[7].floating.n112 x2.x4.x5[7].floating.n111 0.0530294
R16224 x2.x4.x5[7].floating.n130 x2.x4.x5[7].floating.n129 0.0530294
R16225 x2.x4.x5[7].floating.n165 x2.x4.x5[7].floating.n164 0.0530294
R16226 x2.x4.x5[7].floating.n74 x2.x4.x5[7].floating.n73 0.0529559
R16227 x2.x4.x5[7].floating.n50 x2.x4.x5[7].floating.n49 0.0529559
R16228 x2.x4.x5[7].floating.n20 x2.x4.x5[7].floating.n19 0.0529559
R16229 x2.x4.x5[7].floating.n151 x2.x4.x5[7].floating.n150 0.0529559
R16230 x2.x4.x5[7].floating.n73 x2.x4.x5[7].floating.n72 0.0524559
R16231 x2.x4.x5[7].floating.n88 x2.x4.x5[7].floating.n50 0.0524559
R16232 x2.x4.x5[7].floating.n21 x2.x4.x5[7].floating.n20 0.0524559
R16233 x2.x4.x5[7].floating.n150 x2.x4.x5[7].floating.n149 0.0524559
R16234 x2.x4.x5[7].floating.n109 x2.x4.x5[7].floating.n108 0.0523382
R16235 x2.x4.x5[7].floating.n127 x2.x4.x5[7].floating.n126 0.0523382
R16236 x2.x4.x5[7].floating.n168 x2.x4.x5[7].floating.n167 0.0523382
R16237 x2.x4.x5[7].floating.n56 x2.x4.x5[7].floating.n55 0.0516471
R16238 x2.x4.x5[7].floating.n116 x2.x4.x5[7].floating.n115 0.0516471
R16239 x2.x4.x5[7].floating.n134 x2.x4.x5[7].floating.n133 0.0516471
R16240 x2.x4.x5[7].floating.n103 x2.x4.x5[7].floating 0.0495735
R16241 x2.x4.x5[7].floating.n121 x2.x4.x5[7].floating 0.0495735
R16242 x2.x4.x5[7].floating.n139 x2.x4.x5[7].floating 0.0495735
R16243 x2.x4.x5[7].floating.n80 x2.x4.x5[7].floating.n79 0.0408846
R16244 x2.x4.x5[7].floating.n157 x2.x4.x5[7].floating.n156 0.0408846
R16245 x2.x4.x5[7].floating.n15 x2.x4.x5[7].floating.n14 0.0408846
R16246 x2.x4.x5[7].floating.n45 x2.x4.x5[7].floating.n44 0.0408846
R16247 x2.x4.x5[7].floating.n105 x2.x4.x5[7].floating 0.0336765
R16248 x2.x4.x5[7].floating.n123 x2.x4.x5[7].floating 0.0336765
R16249 x2.x4.x5[7].floating x2.x4.x5[7].floating.n171 0.0336765
R16250 x2.x4.x5[7].floating.n30 x2.x4.x5[7].floating.n29 0.0271618
R16251 x2.x4.x5[7].floating.n97 x2.x4.x5[7].floating.n96 0.0271618
R16252 x2.x4.x5[7].floating.n83 x2.x4.x5[7].floating.n82 0.0266618
R16253 x2.x4.x5[7].floating.n41 x2.x4.x5[7].floating.n40 0.0266618
R16254 x2.x4.x5[7].floating.n11 x2.x4.x5[7].floating.n10 0.0266618
R16255 x2.x4.x5[7].floating.n51 x2.x4.x5[7].floating 0.0226176
R16256 x2.x4.x5[7].floating x2.x4.x5[7].floating.n104 0.0226176
R16257 x2.x4.x5[7].floating x2.x4.x5[7].floating.n120 0.0226176
R16258 x2.x4.x5[7].floating x2.x4.x5[7].floating.n122 0.0226176
R16259 x2.x4.x5[7].floating x2.x4.x5[7].floating.n138 0.0226176
R16260 x2.x4.x5[7].floating x2.x4.x5[7].floating.n140 0.0226176
R16261 x2.x4.x5[7].floating.n61 x2.x4.x5[7].floating.n60 0.0191618
R16262 x2.x4.x5[7].floating.n111 x2.x4.x5[7].floating.n110 0.0191618
R16263 x2.x4.x5[7].floating.n129 x2.x4.x5[7].floating.n128 0.0191618
R16264 x2.x4.x5[7].floating.n166 x2.x4.x5[7].floating.n165 0.0191618
R16265 x2.x4.x5[7].floating.n58 x2.x4.x5[7].floating.n57 0.0184706
R16266 x2.x4.x5[7].floating.n114 x2.x4.x5[7].floating.n113 0.0184706
R16267 x2.x4.x5[7].floating.n132 x2.x4.x5[7].floating.n131 0.0184706
R16268 x2.x4.x5[7].floating.n163 x2.x4.x5[7].floating.n162 0.0184706
R16269 x2.x4.x5[7].floating.n82 x2.x4.x5[7].floating.n81 0.014
R16270 x2.x4.x5[7].floating.n72 x2.x4.x5[7].floating.n71 0.014
R16271 x2.x4.x5[7].floating.n46 x2.x4.x5[7].floating.n41 0.014
R16272 x2.x4.x5[7].floating.n22 x2.x4.x5[7].floating.n21 0.014
R16273 x2.x4.x5[7].floating.n16 x2.x4.x5[7].floating.n11 0.014
R16274 x2.x4.x5[7].floating.n149 x2.x4.x5[7].floating.n148 0.014
R16275 x2.x4.x5[7].floating.n159 x2.x4.x5[7].floating.n158 0.014
R16276 x2.x4.x5[7].floating.n89 x2.x4.x5[7].floating.n88 0.014
R16277 x2.x4.x5[7].floating.n75 x2.x4.x5[7].floating.n74 0.0135
R16278 x2.x4.x5[7].floating.n69 x2.x4.x5[7].floating.n64 0.0135
R16279 x2.x4.x5[7].floating.n49 x2.x4.x5[7].floating.n48 0.0135
R16280 x2.x4.x5[7].floating.n29 x2.x4.x5[7].floating.n28 0.0135
R16281 x2.x4.x5[7].floating.n19 x2.x4.x5[7].floating.n18 0.0135
R16282 x2.x4.x5[7].floating.n146 x2.x4.x5[7].floating.n141 0.0135
R16283 x2.x4.x5[7].floating.n152 x2.x4.x5[7].floating.n151 0.0135
R16284 x2.x4.x5[7].floating.n96 x2.x4.x5[7].floating.n95 0.0135
R16285 x2.x4.x5[7].floating.n68 x2.x4.x5[7].floating.n67 0.0120385
R16286 x2.x4.x5[7].floating.n145 x2.x4.x5[7].floating.n144 0.0120385
R16287 x2.x4.x5[7].floating.n27 x2.x4.x5[7].floating.n26 0.0120385
R16288 x2.x4.x5[7].floating.n94 x2.x4.x5[7].floating.n93 0.0120385
R16289 x2.x4.x5[7].floating.n57 x2.x4.x5[7].floating.n56 0.00464706
R16290 x2.x4.x5[7].floating.n115 x2.x4.x5[7].floating.n114 0.00464706
R16291 x2.x4.x5[7].floating.n133 x2.x4.x5[7].floating.n132 0.00464706
R16292 x2.x4.x5[7].floating.n162 x2.x4.x5[7].floating.n161 0.00464706
R16293 x2.x4.x5[7].floating.n62 x2.x4.x5[7].floating.n61 0.00395588
R16294 x2.x4.x5[7].floating.n110 x2.x4.x5[7].floating.n109 0.00395588
R16295 x2.x4.x5[7].floating.n128 x2.x4.x5[7].floating.n127 0.00395588
R16296 x2.x4.x5[7].floating.n167 x2.x4.x5[7].floating.n166 0.00395588
R16297 x2.x4.x5[7].floating.n92 x2.x4.x5[7].floating.n91 0.00359614
R16298 x2.x4.x5[7].floating.n66 x2.x4.x5[7].floating.n65 0.00359614
R16299 x2.x4.x5[7].floating.n143 x2.x4.x5[7].floating.n142 0.00359614
R16300 x2.x4.x5[7].floating.n25 x2.x4.x5[7].floating.n24 0.00359614
R16301 x2.x4.x5[7].floating.n76 x2.x4.x5[7].floating.n75 0.0035
R16302 x2.x4.x5[7].floating.n70 x2.x4.x5[7].floating.n69 0.0035
R16303 x2.x4.x5[7].floating.n48 x2.x4.x5[7].floating.n47 0.0035
R16304 x2.x4.x5[7].floating.n28 x2.x4.x5[7].floating.n23 0.0035
R16305 x2.x4.x5[7].floating.n18 x2.x4.x5[7].floating.n17 0.0035
R16306 x2.x4.x5[7].floating.n147 x2.x4.x5[7].floating.n146 0.0035
R16307 x2.x4.x5[7].floating.n153 x2.x4.x5[7].floating.n152 0.0035
R16308 x2.x4.x5[7].floating.n95 x2.x4.x5[7].floating.n90 0.0035
R16309 x2.x4.x5[7].floating.n81 x2.x4.x5[7].floating.n76 0.003
R16310 x2.x4.x5[7].floating.n71 x2.x4.x5[7].floating.n70 0.003
R16311 x2.x4.x5[7].floating.n47 x2.x4.x5[7].floating.n46 0.003
R16312 x2.x4.x5[7].floating.n23 x2.x4.x5[7].floating.n22 0.003
R16313 x2.x4.x5[7].floating.n17 x2.x4.x5[7].floating.n16 0.003
R16314 x2.x4.x5[7].floating.n148 x2.x4.x5[7].floating.n147 0.003
R16315 x2.x4.x5[7].floating.n158 x2.x4.x5[7].floating.n153 0.003
R16316 x2.x4.x5[7].floating.n90 x2.x4.x5[7].floating.n89 0.003
R16317 x2.x4.x5[7].floating.n155 x2.x4.x5[7].floating.n154 0.00277942
R16318 x2.x4.x5[7].floating.n78 x2.x4.x5[7].floating.n77 0.0023396
R16319 x2.x4.x5[7].floating.n13 x2.x4.x5[7].floating.n12 0.0023396
R16320 x2.x4.x5[7].floating.n43 x2.x4.x5[7].floating.n42 0.0023396
R16321 x2.x4.x5[7].floating.n157 x2.x4.x5[7].floating.n155 0.00233747
R16322 x2.x4.x5[7].floating.n80 x2.x4.x5[7].floating.n78 0.00200689
R16323 x2.x4.x5[7].floating.n15 x2.x4.x5[7].floating.n13 0.00200689
R16324 x2.x4.x5[7].floating.n45 x2.x4.x5[7].floating.n43 0.00200689
R16325 x2.x4.x5[7].floating.n68 x2.x4.x5[7].floating.n66 0.0010233
R16326 x2.x4.x5[7].floating.n145 x2.x4.x5[7].floating.n143 0.0010233
R16327 x2.x4.x5[7].floating.n27 x2.x4.x5[7].floating.n25 0.0010233
R16328 x2.x4.x5[7].floating.n94 x2.x4.x5[7].floating.n92 0.0010233
R16329 x2.x4.x5[7].floating.n81 x2.x4.x5[7].floating.n80 0.00053972
R16330 x2.x4.x5[7].floating.n69 x2.x4.x5[7].floating.n68 0.00053972
R16331 x2.x4.x5[7].floating.n46 x2.x4.x5[7].floating.n45 0.00053972
R16332 x2.x4.x5[7].floating.n28 x2.x4.x5[7].floating.n27 0.00053972
R16333 x2.x4.x5[7].floating.n16 x2.x4.x5[7].floating.n15 0.00053972
R16334 x2.x4.x5[7].floating.n146 x2.x4.x5[7].floating.n145 0.00053972
R16335 x2.x4.x5[7].floating.n158 x2.x4.x5[7].floating.n157 0.00053972
R16336 x2.x4.x5[7].floating.n95 x2.x4.x5[7].floating.n94 0.00053972
R16337 CAP_CTRL_CODE1[3].n0 CAP_CTRL_CODE1[3].t0 229.971
R16338 CAP_CTRL_CODE1[3].n0 CAP_CTRL_CODE1[3].t1 158.35
R16339 CAP_CTRL_CODE1[3].n1 CAP_CTRL_CODE1[3].n0 8.50845
R16340 CAP_CTRL_CODE1[3].n1 CAP_CTRL_CODE1[3] 3.95275
R16341 CAP_CTRL_CODE1[3].n2 CAP_CTRL_CODE1[3].n1 1.73287
R16342 CAP_CTRL_CODE1[3] CAP_CTRL_CODE1[3].n3 0.474765
R16343 CAP_CTRL_CODE1[3].n3 CAP_CTRL_CODE1[3] 0.366977
R16344 CAP_CTRL_CODE1[3].n2 CAP_CTRL_CODE1[3] 0.339042
R16345 CAP_CTRL_CODE1[3].n3 CAP_CTRL_CODE1[3].n2 0.00334091
R16346 CAP_CTRL_CODE0[3].n0 CAP_CTRL_CODE0[3].t1 229.971
R16347 CAP_CTRL_CODE0[3].n0 CAP_CTRL_CODE0[3].t0 158.35
R16348 CAP_CTRL_CODE0[3].n1 CAP_CTRL_CODE0[3].n0 8.50845
R16349 CAP_CTRL_CODE0[3].n1 CAP_CTRL_CODE0[3] 3.95275
R16350 CAP_CTRL_CODE0[3].n2 CAP_CTRL_CODE0[3].n1 1.73287
R16351 CAP_CTRL_CODE0[3] CAP_CTRL_CODE0[3].n3 0.474765
R16352 CAP_CTRL_CODE0[3].n3 CAP_CTRL_CODE0[3] 0.366977
R16353 CAP_CTRL_CODE0[3].n2 CAP_CTRL_CODE0[3] 0.339042
R16354 CAP_CTRL_CODE0[3].n3 CAP_CTRL_CODE0[3].n2 0.00334091
R16355 x2.x2.x10.Y.n5 x2.x2.x10.Y.n0 304.151
R16356 x2.x2.x10.Y x2.x2.x10.Y.t3 154.8
R16357 x2.x2.x10.Y x2.x2.x10.Y.t2 154.8
R16358 x2.x2.x10.Y x2.x2.x10.Y.t8 154.8
R16359 x2.x2.x10.Y x2.x2.x10.Y.t6 154.8
R16360 x2.x2.x10.Y x2.x2.x10.Y.t7 154.8
R16361 x2.x2.x10.Y x2.x2.x10.Y.t4 154.8
R16362 x2.x2.x10.Y x2.x2.x10.Y.t5 154.8
R16363 x2.x2.x10.Y x2.x2.x10.Y.t9 154.8
R16364 x2.x2.x10.Y.n2 x2.x2.x10.Y.n0 143.207
R16365 x2.x2.x10.Y x2.x2.x10.Y.n5 134.663
R16366 x2.x2.x10.Y x2.x2.x10.Y.t0 116.097
R16367 x2.x2.x10.Y.n3 x2.x2.x10.Y.t1 25.626
R16368 x2.x2.x10.Y.n1 x2.x2.x10.Y 11.6875
R16369 x2.x2.x10.Y.n4 x2.x2.x10.Y.n3 9.14446
R16370 x2.x2.x10.Y.n2 x2.x2.x10.Y 7.45722
R16371 x2.x2.x10.Y.n4 x2.x2.x10.Y.n2 7.43775
R16372 x2.x2.x10.Y.n1 x2.x2.x10.Y 7.23528
R16373 x2.x2.x10.Y x2.x2.x10.Y.n1 5.04292
R16374 x2.x2.x10.Y.n3 x2.x2.x10.Y.n0 0.969421
R16375 x2.x2.x10.Y.n5 x2.x2.x10.Y.n4 0.652645
R16376 x2.x2.x5[7].floating.n6 x2.x2.x5[7].floating.t0 68.0345
R16377 x2.x2.x5[7].floating.n27 x2.x2.x5[7].floating.t4 68.0345
R16378 x2.x2.x5[7].floating.n45 x2.x2.x5[7].floating.t5 68.0345
R16379 x2.x2.x5[7].floating.n57 x2.x2.x5[7].floating.t2 68.0345
R16380 x2.x2.x5[7].floating.n75 x2.x2.x5[7].floating.t3 68.0345
R16381 x2.x2.x5[7].floating.n87 x2.x2.x5[7].floating.t1 68.0345
R16382 x2.x2.x5[7].floating.n105 x2.x2.x5[7].floating.t7 68.0345
R16383 x2.x2.x5[7].floating.n116 x2.x2.x5[7].floating.t6 68.0345
R16384 x2.x2.x5[7].floating.n135 x2.x2.x5[7].floating.n97 0.660401
R16385 x2.x2.x5[7].floating.n144 x2.x2.x5[7].floating.n82 0.660401
R16386 x2.x2.x5[7].floating.n153 x2.x2.x5[7].floating.n67 0.660401
R16387 x2.x2.x5[7].floating.n162 x2.x2.x5[7].floating.n52 0.660401
R16388 x2.x2.x5[7].floating.n171 x2.x2.x5[7].floating.n37 0.660401
R16389 x2.x2.x5[7].floating.n11 x2.x2.x5[7].floating.n10 0.320345
R16390 x2.x2.x5[7].floating.n122 x2.x2.x5[7].floating.n121 0.308269
R16391 x2.x2.x5[7].floating.n123 x2.x2.x5[7].floating.n122 0.173084
R16392 x2.x2.x5[7].floating.n12 x2.x2.x5[7].floating.n11 0.162103
R16393 x2.x2.x5[7].floating.n122 x2.x2.x5[7].floating 0.100688
R16394 x2.x2.x5[7].floating.n11 x2.x2.x5[7].floating 0.0755007
R16395 x2.x2.x5[7].floating.n97 x2.x2.x5[7].floating.n96 0.0716912
R16396 x2.x2.x5[7].floating.n98 x2.x2.x5[7].floating.n97 0.0716912
R16397 x2.x2.x5[7].floating.n67 x2.x2.x5[7].floating.n66 0.0716912
R16398 x2.x2.x5[7].floating.n68 x2.x2.x5[7].floating.n67 0.0716912
R16399 x2.x2.x5[7].floating.n37 x2.x2.x5[7].floating.n36 0.0716912
R16400 x2.x2.x5[7].floating.n38 x2.x2.x5[7].floating.n37 0.0716912
R16401 x2.x2.x5[7].floating.n171 x2.x2.x5[7].floating.n170 0.0716912
R16402 x2.x2.x5[7].floating.n153 x2.x2.x5[7].floating.n152 0.0716912
R16403 x2.x2.x5[7].floating.n135 x2.x2.x5[7].floating.n134 0.0716912
R16404 x2.x2.x5[7].floating.n93 x2.x2.x5[7].floating.n92 0.0557941
R16405 x2.x2.x5[7].floating.n94 x2.x2.x5[7].floating.n93 0.0557941
R16406 x2.x2.x5[7].floating.n95 x2.x2.x5[7].floating.n94 0.0557941
R16407 x2.x2.x5[7].floating.n96 x2.x2.x5[7].floating.n95 0.0557941
R16408 x2.x2.x5[7].floating.n99 x2.x2.x5[7].floating.n98 0.0557941
R16409 x2.x2.x5[7].floating.n100 x2.x2.x5[7].floating.n99 0.0557941
R16410 x2.x2.x5[7].floating.n101 x2.x2.x5[7].floating.n100 0.0557941
R16411 x2.x2.x5[7].floating.n102 x2.x2.x5[7].floating.n101 0.0557941
R16412 x2.x2.x5[7].floating.n63 x2.x2.x5[7].floating.n62 0.0557941
R16413 x2.x2.x5[7].floating.n64 x2.x2.x5[7].floating.n63 0.0557941
R16414 x2.x2.x5[7].floating.n65 x2.x2.x5[7].floating.n64 0.0557941
R16415 x2.x2.x5[7].floating.n66 x2.x2.x5[7].floating.n65 0.0557941
R16416 x2.x2.x5[7].floating.n69 x2.x2.x5[7].floating.n68 0.0557941
R16417 x2.x2.x5[7].floating.n70 x2.x2.x5[7].floating.n69 0.0557941
R16418 x2.x2.x5[7].floating.n71 x2.x2.x5[7].floating.n70 0.0557941
R16419 x2.x2.x5[7].floating.n72 x2.x2.x5[7].floating.n71 0.0557941
R16420 x2.x2.x5[7].floating.n33 x2.x2.x5[7].floating.n32 0.0557941
R16421 x2.x2.x5[7].floating.n34 x2.x2.x5[7].floating.n33 0.0557941
R16422 x2.x2.x5[7].floating.n35 x2.x2.x5[7].floating.n34 0.0557941
R16423 x2.x2.x5[7].floating.n36 x2.x2.x5[7].floating.n35 0.0557941
R16424 x2.x2.x5[7].floating.n39 x2.x2.x5[7].floating.n38 0.0557941
R16425 x2.x2.x5[7].floating.n40 x2.x2.x5[7].floating.n39 0.0557941
R16426 x2.x2.x5[7].floating.n41 x2.x2.x5[7].floating.n40 0.0557941
R16427 x2.x2.x5[7].floating.n42 x2.x2.x5[7].floating.n41 0.0557941
R16428 x2.x2.x5[7].floating.n20 x2.x2.x5[7].floating.n19 0.0557941
R16429 x2.x2.x5[7].floating.n21 x2.x2.x5[7].floating.n20 0.0557941
R16430 x2.x2.x5[7].floating.n22 x2.x2.x5[7].floating.n21 0.0557941
R16431 x2.x2.x5[7].floating.n23 x2.x2.x5[7].floating.n22 0.0557941
R16432 x2.x2.x5[7].floating.n169 x2.x2.x5[7].floating.n168 0.0557941
R16433 x2.x2.x5[7].floating.n168 x2.x2.x5[7].floating.n167 0.0557941
R16434 x2.x2.x5[7].floating.n167 x2.x2.x5[7].floating.n166 0.0557941
R16435 x2.x2.x5[7].floating.n158 x2.x2.x5[7].floating.n157 0.0557941
R16436 x2.x2.x5[7].floating.n157 x2.x2.x5[7].floating.n156 0.0557941
R16437 x2.x2.x5[7].floating.n156 x2.x2.x5[7].floating.n155 0.0557941
R16438 x2.x2.x5[7].floating.n155 x2.x2.x5[7].floating.n154 0.0557941
R16439 x2.x2.x5[7].floating.n151 x2.x2.x5[7].floating.n150 0.0557941
R16440 x2.x2.x5[7].floating.n150 x2.x2.x5[7].floating.n149 0.0557941
R16441 x2.x2.x5[7].floating.n149 x2.x2.x5[7].floating.n148 0.0557941
R16442 x2.x2.x5[7].floating.n140 x2.x2.x5[7].floating.n139 0.0557941
R16443 x2.x2.x5[7].floating.n139 x2.x2.x5[7].floating.n138 0.0557941
R16444 x2.x2.x5[7].floating.n138 x2.x2.x5[7].floating.n137 0.0557941
R16445 x2.x2.x5[7].floating.n137 x2.x2.x5[7].floating.n136 0.0557941
R16446 x2.x2.x5[7].floating.n133 x2.x2.x5[7].floating.n132 0.0557941
R16447 x2.x2.x5[7].floating.n132 x2.x2.x5[7].floating.n131 0.0557941
R16448 x2.x2.x5[7].floating.n131 x2.x2.x5[7].floating.n130 0.0557941
R16449 x2.x2.x5[7].floating.n16 x2.x2.x5[7].floating.n15 0.0537206
R16450 x2.x2.x5[7].floating.n162 x2.x2.x5[7].floating.n161 0.0537206
R16451 x2.x2.x5[7].floating.n144 x2.x2.x5[7].floating.n143 0.0537206
R16452 x2.x2.x5[7].floating.n126 x2.x2.x5[7].floating.n125 0.0537206
R16453 x2.x2.x5[7].floating.n15 x2.x2.x5[7].floating.n14 0.0530294
R16454 x2.x2.x5[7].floating.n163 x2.x2.x5[7].floating.n162 0.0530294
R16455 x2.x2.x5[7].floating.n145 x2.x2.x5[7].floating.n144 0.0530294
R16456 x2.x2.x5[7].floating.n127 x2.x2.x5[7].floating.n126 0.0530294
R16457 x2.x2.x5[7].floating.n83 x2.x2.x5[7].floating.n82 0.0529559
R16458 x2.x2.x5[7].floating.n53 x2.x2.x5[7].floating.n52 0.0529559
R16459 x2.x2.x5[7].floating.n1 x2.x2.x5[7].floating.n0 0.0529559
R16460 x2.x2.x5[7].floating.n113 x2.x2.x5[7].floating.n112 0.0529559
R16461 x2.x2.x5[7].floating.n112 x2.x2.x5[7].floating.n111 0.0524559
R16462 x2.x2.x5[7].floating.n82 x2.x2.x5[7].floating.n81 0.0524559
R16463 x2.x2.x5[7].floating.n52 x2.x2.x5[7].floating.n51 0.0524559
R16464 x2.x2.x5[7].floating.n2 x2.x2.x5[7].floating.n1 0.0524559
R16465 x2.x2.x5[7].floating.n166 x2.x2.x5[7].floating.n165 0.0523382
R16466 x2.x2.x5[7].floating.n148 x2.x2.x5[7].floating.n147 0.0523382
R16467 x2.x2.x5[7].floating.n130 x2.x2.x5[7].floating.n129 0.0523382
R16468 x2.x2.x5[7].floating.n19 x2.x2.x5[7].floating.n18 0.0516471
R16469 x2.x2.x5[7].floating.n159 x2.x2.x5[7].floating.n158 0.0516471
R16470 x2.x2.x5[7].floating.n141 x2.x2.x5[7].floating.n140 0.0516471
R16471 x2.x2.x5[7].floating x2.x2.x5[7].floating.n171 0.0495735
R16472 x2.x2.x5[7].floating x2.x2.x5[7].floating.n153 0.0495735
R16473 x2.x2.x5[7].floating x2.x2.x5[7].floating.n135 0.0495735
R16474 x2.x2.x5[7].floating.n8 x2.x2.x5[7].floating.n5 0.0408846
R16475 x2.x2.x5[7].floating.n47 x2.x2.x5[7].floating.n44 0.0408846
R16476 x2.x2.x5[7].floating.n77 x2.x2.x5[7].floating.n74 0.0408846
R16477 x2.x2.x5[7].floating.n107 x2.x2.x5[7].floating.n104 0.0408846
R16478 x2.x2.x5[7].floating x2.x2.x5[7].floating.n169 0.0336765
R16479 x2.x2.x5[7].floating x2.x2.x5[7].floating.n151 0.0336765
R16480 x2.x2.x5[7].floating x2.x2.x5[7].floating.n133 0.0336765
R16481 x2.x2.x5[7].floating.n103 x2.x2.x5[7].floating.n102 0.0271618
R16482 x2.x2.x5[7].floating.n73 x2.x2.x5[7].floating.n72 0.0271618
R16483 x2.x2.x5[7].floating.n43 x2.x2.x5[7].floating.n42 0.0271618
R16484 x2.x2.x5[7].floating.n92 x2.x2.x5[7].floating.n91 0.0266618
R16485 x2.x2.x5[7].floating.n62 x2.x2.x5[7].floating.n61 0.0266618
R16486 x2.x2.x5[7].floating.n32 x2.x2.x5[7].floating.n31 0.0266618
R16487 x2.x2.x5[7].floating x2.x2.x5[7].floating.n23 0.0226176
R16488 x2.x2.x5[7].floating.n170 x2.x2.x5[7].floating 0.0226176
R16489 x2.x2.x5[7].floating.n154 x2.x2.x5[7].floating 0.0226176
R16490 x2.x2.x5[7].floating.n152 x2.x2.x5[7].floating 0.0226176
R16491 x2.x2.x5[7].floating.n136 x2.x2.x5[7].floating 0.0226176
R16492 x2.x2.x5[7].floating.n134 x2.x2.x5[7].floating 0.0226176
R16493 x2.x2.x5[7].floating.n119 x2.x2.x5[7].floating.n118 0.021208
R16494 x2.x2.x5[7].floating.n14 x2.x2.x5[7].floating.n13 0.0191618
R16495 x2.x2.x5[7].floating.n164 x2.x2.x5[7].floating.n163 0.0191618
R16496 x2.x2.x5[7].floating.n146 x2.x2.x5[7].floating.n145 0.0191618
R16497 x2.x2.x5[7].floating.n128 x2.x2.x5[7].floating.n127 0.0191618
R16498 x2.x2.x5[7].floating.n17 x2.x2.x5[7].floating.n16 0.0184706
R16499 x2.x2.x5[7].floating.n161 x2.x2.x5[7].floating.n160 0.0184706
R16500 x2.x2.x5[7].floating.n143 x2.x2.x5[7].floating.n142 0.0184706
R16501 x2.x2.x5[7].floating.n125 x2.x2.x5[7].floating.n124 0.0184706
R16502 x2.x2.x5[7].floating.n111 x2.x2.x5[7].floating.n110 0.014
R16503 x2.x2.x5[7].floating.n91 x2.x2.x5[7].floating.n90 0.014
R16504 x2.x2.x5[7].floating.n81 x2.x2.x5[7].floating.n80 0.014
R16505 x2.x2.x5[7].floating.n61 x2.x2.x5[7].floating.n60 0.014
R16506 x2.x2.x5[7].floating.n51 x2.x2.x5[7].floating.n50 0.014
R16507 x2.x2.x5[7].floating.n31 x2.x2.x5[7].floating.n30 0.014
R16508 x2.x2.x5[7].floating.n3 x2.x2.x5[7].floating.n2 0.014
R16509 x2.x2.x5[7].floating.n121 x2.x2.x5[7].floating.n120 0.014
R16510 x2.x2.x5[7].floating.n108 x2.x2.x5[7].floating.n103 0.0135
R16511 x2.x2.x5[7].floating.n84 x2.x2.x5[7].floating.n83 0.0135
R16512 x2.x2.x5[7].floating.n78 x2.x2.x5[7].floating.n73 0.0135
R16513 x2.x2.x5[7].floating.n54 x2.x2.x5[7].floating.n53 0.0135
R16514 x2.x2.x5[7].floating.n48 x2.x2.x5[7].floating.n43 0.0135
R16515 x2.x2.x5[7].floating.n10 x2.x2.x5[7].floating.n9 0.0135
R16516 x2.x2.x5[7].floating.n114 x2.x2.x5[7].floating.n113 0.0135
R16517 x2.x2.x5[7].floating.n29 x2.x2.x5[7].floating.n26 0.0101154
R16518 x2.x2.x5[7].floating.n59 x2.x2.x5[7].floating.n56 0.0101154
R16519 x2.x2.x5[7].floating.n89 x2.x2.x5[7].floating.n86 0.0101154
R16520 x2.x2.x5[7].floating.n18 x2.x2.x5[7].floating.n17 0.00464706
R16521 x2.x2.x5[7].floating.n160 x2.x2.x5[7].floating.n159 0.00464706
R16522 x2.x2.x5[7].floating.n142 x2.x2.x5[7].floating.n141 0.00464706
R16523 x2.x2.x5[7].floating.n124 x2.x2.x5[7].floating.n123 0.00464706
R16524 x2.x2.x5[7].floating.n13 x2.x2.x5[7].floating.n12 0.00395588
R16525 x2.x2.x5[7].floating.n165 x2.x2.x5[7].floating.n164 0.00395588
R16526 x2.x2.x5[7].floating.n147 x2.x2.x5[7].floating.n146 0.00395588
R16527 x2.x2.x5[7].floating.n129 x2.x2.x5[7].floating.n128 0.00395588
R16528 x2.x2.x5[7].floating.n109 x2.x2.x5[7].floating.n108 0.0035
R16529 x2.x2.x5[7].floating.n85 x2.x2.x5[7].floating.n84 0.0035
R16530 x2.x2.x5[7].floating.n79 x2.x2.x5[7].floating.n78 0.0035
R16531 x2.x2.x5[7].floating.n55 x2.x2.x5[7].floating.n54 0.0035
R16532 x2.x2.x5[7].floating.n49 x2.x2.x5[7].floating.n48 0.0035
R16533 x2.x2.x5[7].floating.n25 x2.x2.x5[7].floating.n24 0.0035
R16534 x2.x2.x5[7].floating.n9 x2.x2.x5[7].floating.n4 0.0035
R16535 x2.x2.x5[7].floating.n115 x2.x2.x5[7].floating.n114 0.0035
R16536 x2.x2.x5[7].floating.n110 x2.x2.x5[7].floating.n109 0.003
R16537 x2.x2.x5[7].floating.n90 x2.x2.x5[7].floating.n85 0.003
R16538 x2.x2.x5[7].floating.n80 x2.x2.x5[7].floating.n79 0.003
R16539 x2.x2.x5[7].floating.n60 x2.x2.x5[7].floating.n55 0.003
R16540 x2.x2.x5[7].floating.n50 x2.x2.x5[7].floating.n49 0.003
R16541 x2.x2.x5[7].floating.n30 x2.x2.x5[7].floating.n25 0.003
R16542 x2.x2.x5[7].floating.n4 x2.x2.x5[7].floating.n3 0.003
R16543 x2.x2.x5[7].floating.n120 x2.x2.x5[7].floating.n115 0.003
R16544 x2.x2.x5[7].floating.n28 x2.x2.x5[7].floating.n27 0.00260608
R16545 x2.x2.x5[7].floating.n58 x2.x2.x5[7].floating.n57 0.00260608
R16546 x2.x2.x5[7].floating.n88 x2.x2.x5[7].floating.n87 0.00260608
R16547 x2.x2.x5[7].floating.n117 x2.x2.x5[7].floating.n116 0.00234008
R16548 x2.x2.x5[7].floating.n119 x2.x2.x5[7].floating.n117 0.00200725
R16549 x2.x2.x5[7].floating.n7 x2.x2.x5[7].floating.n6 0.00177054
R16550 x2.x2.x5[7].floating.n46 x2.x2.x5[7].floating.n45 0.00177054
R16551 x2.x2.x5[7].floating.n76 x2.x2.x5[7].floating.n75 0.00177054
R16552 x2.x2.x5[7].floating.n106 x2.x2.x5[7].floating.n105 0.00177054
R16553 x2.x2.x5[7].floating.n8 x2.x2.x5[7].floating.n7 0.00174992
R16554 x2.x2.x5[7].floating.n47 x2.x2.x5[7].floating.n46 0.00174992
R16555 x2.x2.x5[7].floating.n77 x2.x2.x5[7].floating.n76 0.00174992
R16556 x2.x2.x5[7].floating.n107 x2.x2.x5[7].floating.n106 0.00174992
R16557 x2.x2.x5[7].floating.n29 x2.x2.x5[7].floating.n28 0.00101477
R16558 x2.x2.x5[7].floating.n59 x2.x2.x5[7].floating.n58 0.00101477
R16559 x2.x2.x5[7].floating.n89 x2.x2.x5[7].floating.n88 0.00101477
R16560 x2.x2.x5[7].floating.n108 x2.x2.x5[7].floating.n107 0.00053972
R16561 x2.x2.x5[7].floating.n90 x2.x2.x5[7].floating.n89 0.00053972
R16562 x2.x2.x5[7].floating.n78 x2.x2.x5[7].floating.n77 0.00053972
R16563 x2.x2.x5[7].floating.n60 x2.x2.x5[7].floating.n59 0.00053972
R16564 x2.x2.x5[7].floating.n48 x2.x2.x5[7].floating.n47 0.00053972
R16565 x2.x2.x5[7].floating.n30 x2.x2.x5[7].floating.n29 0.00053972
R16566 x2.x2.x5[7].floating.n9 x2.x2.x5[7].floating.n8 0.00053972
R16567 x2.x2.x5[7].floating.n120 x2.x2.x5[7].floating.n119 0.00053972
R16568 sample_clk.n3 sample_clk.t0 47.1678
R16569 sample_clk.n2 sample_clk.t2 47.1434
R16570 sample_clk.n2 sample_clk.t1 47.1434
R16571 sample_clk.n1 sample_clk.t3 25.8015
R16572 sample_clk.n0 sample_clk.t5 25.7981
R16573 sample_clk.n0 sample_clk.t4 25.7981
R16574 sample_clk.n1 sample_clk.n0 1.46997
R16575 sample_clk.n3 sample_clk.n2 1.03455
R16576 sample_clk sample_clk.n3 0.498236
R16577 sample_clk sample_clk.n1 0.299413
R16578 sample_delay_offset.n34 sample_delay_offset.t6 230.016
R16579 sample_delay_offset.n13 sample_delay_offset.t3 230.016
R16580 sample_delay_offset.n21 sample_delay_offset.t4 229.971
R16581 sample_delay_offset.n1 sample_delay_offset.t0 229.971
R16582 sample_delay_offset.n21 sample_delay_offset.t11 158.351
R16583 sample_delay_offset.n1 sample_delay_offset.t8 158.351
R16584 sample_delay_offset.n33 sample_delay_offset.t10 153.665
R16585 sample_delay_offset.n12 sample_delay_offset.t9 153.665
R16586 sample_delay_offset.n34 sample_delay_offset 153.601
R16587 sample_delay_offset.n13 sample_delay_offset 153.601
R16588 sample_delay_offset sample_delay_offset.t5 140.379
R16589 sample_delay_offset sample_delay_offset.t2 140.379
R16590 sample_delay_offset.n29 sample_delay_offset.t7 140.34
R16591 sample_delay_offset.n9 sample_delay_offset.t1 140.34
R16592 sample_delay_offset.n35 sample_delay_offset.n34 9.3005
R16593 sample_delay_offset.n14 sample_delay_offset.n13 9.3005
R16594 sample_delay_offset.n19 sample_delay_offset.n10 9.14466
R16595 sample_delay_offset.n22 sample_delay_offset.n21 7.39809
R16596 sample_delay_offset.n2 sample_delay_offset.n1 7.39809
R16597 sample_delay_offset.n40 sample_delay_offset.n39 5.90325
R16598 sample_delay_offset.n40 sample_delay_offset.n31 5.46925
R16599 sample_delay_offset.n34 sample_delay_offset.n33 4.91671
R16600 sample_delay_offset.n13 sample_delay_offset.n12 4.91671
R16601 sample_delay_offset.n16 sample_delay_offset.n14 4.90192
R16602 sample_delay_offset.n37 sample_delay_offset.n35 4.9013
R16603 sample_delay_offset.n30 sample_delay_offset.n29 4.18104
R16604 sample_delay_offset.n10 sample_delay_offset.n9 4.18104
R16605 sample_delay_offset.n39 sample_delay_offset 4.14309
R16606 sample_delay_offset.n18 sample_delay_offset 4.14309
R16607 sample_delay_offset.n24 sample_delay_offset.n23 4.0005
R16608 sample_delay_offset.n4 sample_delay_offset.n3 4.0005
R16609 sample_delay_offset.n19 sample_delay_offset.n18 3.76287
R16610 sample_delay_offset.n31 sample_delay_offset.n30 3.75602
R16611 sample_delay_offset.n25 sample_delay_offset.n24 3.03311
R16612 sample_delay_offset.n5 sample_delay_offset.n4 3.03311
R16613 sample_delay_offset sample_delay_offset.n32 2.4005
R16614 sample_delay_offset sample_delay_offset.n11 2.4005
R16615 sample_delay_offset.n31 sample_delay_offset.n19 2.01947
R16616 sample_delay_offset.n28 sample_delay_offset.n27 1.87694
R16617 sample_delay_offset.n8 sample_delay_offset.n7 1.87694
R16618 sample_delay_offset.n23 sample_delay_offset 1.6005
R16619 sample_delay_offset.n3 sample_delay_offset 1.6005
R16620 sample_delay_offset.n28 sample_delay_offset 1.43349
R16621 sample_delay_offset.n8 sample_delay_offset 1.43349
R16622 sample_delay_offset.n27 sample_delay_offset.n26 1.12626
R16623 sample_delay_offset.n7 sample_delay_offset.n6 1.12626
R16624 sample_delay_offset.n38 sample_delay_offset 1.01229
R16625 sample_delay_offset.n17 sample_delay_offset 1.01229
R16626 sample_delay_offset.n38 sample_delay_offset.n37 0.726043
R16627 sample_delay_offset.n30 sample_delay_offset.n28 0.726043
R16628 sample_delay_offset.n10 sample_delay_offset.n8 0.726043
R16629 sample_delay_offset.n17 sample_delay_offset.n16 0.726043
R16630 sample_delay_offset sample_delay_offset.n40 0.718134
R16631 sample_delay_offset.n35 sample_delay_offset.n32 0.533833
R16632 sample_delay_offset.n24 sample_delay_offset.n22 0.533833
R16633 sample_delay_offset.n4 sample_delay_offset.n2 0.533833
R16634 sample_delay_offset.n14 sample_delay_offset.n11 0.533833
R16635 sample_delay_offset.n37 sample_delay_offset.n36 0.421696
R16636 sample_delay_offset.n16 sample_delay_offset.n15 0.421696
R16637 sample_delay_offset.n39 sample_delay_offset.n38 0.0783302
R16638 sample_delay_offset.n18 sample_delay_offset.n17 0.0783302
R16639 sample_delay_offset.n30 sample_delay_offset 0.0447308
R16640 sample_delay_offset.n10 sample_delay_offset 0.0447308
R16641 sample_delay_offset.n29 sample_delay_offset 0.0384464
R16642 sample_delay_offset.n9 sample_delay_offset 0.0384464
R16643 sample_delay_offset.n36 sample_delay_offset 0.0195217
R16644 sample_delay_offset.n30 sample_delay_offset 0.0195217
R16645 sample_delay_offset.n10 sample_delay_offset 0.0195217
R16646 sample_delay_offset.n15 sample_delay_offset 0.0195217
R16647 sample_delay_offset.n25 sample_delay_offset.n20 0.0179598
R16648 sample_delay_offset.n5 sample_delay_offset.n0 0.0179598
R16649 sample_delay_offset.n36 sample_delay_offset 0.0170094
R16650 sample_delay_offset.n15 sample_delay_offset 0.0170094
R16651 sample_delay_offset.n26 sample_delay_offset.n25 0.00504545
R16652 sample_delay_offset.n6 sample_delay_offset.n5 0.00504545
R16653 CAP_CTRL_CODE3[2] CAP_CTRL_CODE3[2].t1 140.387
R16654 CAP_CTRL_CODE3[2].n2 CAP_CTRL_CODE3[2].t2 140.34
R16655 CAP_CTRL_CODE3[2].n0 CAP_CTRL_CODE3[2].t0 140.34
R16656 CAP_CTRL_CODE3[2].n1 CAP_CTRL_CODE3[2].t3 140.34
R16657 CAP_CTRL_CODE3[2] CAP_CTRL_CODE3[2].n1 2.87278
R16658 CAP_CTRL_CODE3[2] CAP_CTRL_CODE3[2].n0 0.285826
R16659 CAP_CTRL_CODE3[2].n2 CAP_CTRL_CODE3[2] 0.220255
R16660 CAP_CTRL_CODE3[2].n1 CAP_CTRL_CODE3[2] 0.0466957
R16661 CAP_CTRL_CODE3[2].n0 CAP_CTRL_CODE3[2] 0.0466957
R16662 CAP_CTRL_CODE3[2] CAP_CTRL_CODE3[2].n2 0.00210741
R16663 CAP_CTRL_CODE3[3].n0 CAP_CTRL_CODE3[3].t0 229.964
R16664 CAP_CTRL_CODE3[3].n0 CAP_CTRL_CODE3[3].t1 158.363
R16665 CAP_CTRL_CODE3[3].n1 CAP_CTRL_CODE3[3].n0 8.13263
R16666 CAP_CTRL_CODE3[3].n1 CAP_CTRL_CODE3[3] 2.67916
R16667 CAP_CTRL_CODE3[3].n2 CAP_CTRL_CODE3[3] 2.1255
R16668 CAP_CTRL_CODE3[3] CAP_CTRL_CODE3[3].n1 1.84241
R16669 CAP_CTRL_CODE3[3].n2 CAP_CTRL_CODE3[3] 0.434324
R16670 CAP_CTRL_CODE3[3].n2 CAP_CTRL_CODE3[3] 0.271333
R16671 CAP_CTRL_CODE3[3] CAP_CTRL_CODE3[3].n2 0.0335882
R16672 x2.x3.x10.Y.n5 x2.x3.x10.Y.n0 304.151
R16673 x2.x3.x10.Y x2.x3.x10.Y.t6 154.8
R16674 x2.x3.x10.Y x2.x3.x10.Y.t7 154.8
R16675 x2.x3.x10.Y x2.x3.x10.Y.t5 154.8
R16676 x2.x3.x10.Y x2.x3.x10.Y.t4 154.8
R16677 x2.x3.x10.Y x2.x3.x10.Y.t3 154.8
R16678 x2.x3.x10.Y x2.x3.x10.Y.t9 154.8
R16679 x2.x3.x10.Y x2.x3.x10.Y.t8 154.8
R16680 x2.x3.x10.Y x2.x3.x10.Y.t2 154.8
R16681 x2.x3.x10.Y.n2 x2.x3.x10.Y.n0 143.207
R16682 x2.x3.x10.Y x2.x3.x10.Y.n5 134.663
R16683 x2.x3.x10.Y x2.x3.x10.Y.t0 116.097
R16684 x2.x3.x10.Y.n3 x2.x3.x10.Y.t1 25.626
R16685 x2.x3.x10.Y.n1 x2.x3.x10.Y 11.6875
R16686 x2.x3.x10.Y.n4 x2.x3.x10.Y.n3 9.14446
R16687 x2.x3.x10.Y.n2 x2.x3.x10.Y 7.45722
R16688 x2.x3.x10.Y.n4 x2.x3.x10.Y.n2 7.43775
R16689 x2.x3.x10.Y.n1 x2.x3.x10.Y 7.23528
R16690 x2.x3.x10.Y x2.x3.x10.Y.n1 5.04292
R16691 x2.x3.x10.Y.n3 x2.x3.x10.Y.n0 0.969421
R16692 x2.x3.x10.Y.n5 x2.x3.x10.Y.n4 0.652645
R16693 sample_clk_b.n3 sample_clk_b.t2 47.1678
R16694 sample_clk_b.n2 sample_clk_b.t1 47.1434
R16695 sample_clk_b.n2 sample_clk_b.t0 47.1434
R16696 sample_clk_b.n1 sample_clk_b.t5 25.8015
R16697 sample_clk_b.n0 sample_clk_b.t4 25.7981
R16698 sample_clk_b.n0 sample_clk_b.t3 25.7981
R16699 sample_clk_b.n1 sample_clk_b.n0 1.46997
R16700 sample_clk_b.n3 sample_clk_b.n2 1.03455
R16701 sample_clk_b sample_clk_b.n1 0.731478
R16702 sample_clk_b sample_clk_b.n3 0.0847391
R16703 x2.x3.x5[7].floating.n67 x2.x3.x5[7].floating.t5 68.0345
R16704 x2.x3.x5[7].floating.n79 x2.x3.x5[7].floating.t4 68.0345
R16705 x2.x3.x5[7].floating.n97 x2.x3.x5[7].floating.t2 68.0345
R16706 x2.x3.x5[7].floating.n109 x2.x3.x5[7].floating.t3 68.0345
R16707 x2.x3.x5[7].floating.n6 x2.x3.x5[7].floating.t7 68.0345
R16708 x2.x3.x5[7].floating.n27 x2.x3.x5[7].floating.t1 68.0345
R16709 x2.x3.x5[7].floating.n46 x2.x3.x5[7].floating.t0 68.0345
R16710 x2.x3.x5[7].floating.n154 x2.x3.x5[7].floating.t6 68.0345
R16711 x2.x3.x5[7].floating.n127 x2.x3.x5[7].floating.n89 0.660401
R16712 x2.x3.x5[7].floating.n136 x2.x3.x5[7].floating.n74 0.660401
R16713 x2.x3.x5[7].floating.n146 x2.x3.x5[7].floating.n145 0.660401
R16714 x2.x3.x5[7].floating.n171 x2.x3.x5[7].floating.n37 0.660401
R16715 x2.x3.x5[7].floating.n162 x2.x3.x5[7].floating.n161 0.660401
R16716 x2.x3.x5[7].floating.n11 x2.x3.x5[7].floating.n10 0.320345
R16717 x2.x3.x5[7].floating.n114 x2.x3.x5[7].floating.n113 0.308269
R16718 x2.x3.x5[7].floating.n115 x2.x3.x5[7].floating.n114 0.173084
R16719 x2.x3.x5[7].floating.n12 x2.x3.x5[7].floating.n11 0.162103
R16720 x2.x3.x5[7].floating.n114 x2.x3.x5[7].floating 0.100688
R16721 x2.x3.x5[7].floating.n11 x2.x3.x5[7].floating 0.0755007
R16722 x2.x3.x5[7].floating.n89 x2.x3.x5[7].floating.n88 0.0716912
R16723 x2.x3.x5[7].floating.n90 x2.x3.x5[7].floating.n89 0.0716912
R16724 x2.x3.x5[7].floating.n147 x2.x3.x5[7].floating.n146 0.0716912
R16725 x2.x3.x5[7].floating.n146 x2.x3.x5[7].floating.n53 0.0716912
R16726 x2.x3.x5[7].floating.n37 x2.x3.x5[7].floating.n36 0.0716912
R16727 x2.x3.x5[7].floating.n39 x2.x3.x5[7].floating.n37 0.0716912
R16728 x2.x3.x5[7].floating.n171 x2.x3.x5[7].floating.n170 0.0716912
R16729 x2.x3.x5[7].floating.n145 x2.x3.x5[7].floating.n144 0.0716912
R16730 x2.x3.x5[7].floating.n127 x2.x3.x5[7].floating.n126 0.0716912
R16731 x2.x3.x5[7].floating.n85 x2.x3.x5[7].floating.n84 0.0557941
R16732 x2.x3.x5[7].floating.n86 x2.x3.x5[7].floating.n85 0.0557941
R16733 x2.x3.x5[7].floating.n87 x2.x3.x5[7].floating.n86 0.0557941
R16734 x2.x3.x5[7].floating.n88 x2.x3.x5[7].floating.n87 0.0557941
R16735 x2.x3.x5[7].floating.n91 x2.x3.x5[7].floating.n90 0.0557941
R16736 x2.x3.x5[7].floating.n92 x2.x3.x5[7].floating.n91 0.0557941
R16737 x2.x3.x5[7].floating.n93 x2.x3.x5[7].floating.n92 0.0557941
R16738 x2.x3.x5[7].floating.n94 x2.x3.x5[7].floating.n93 0.0557941
R16739 x2.x3.x5[7].floating.n151 x2.x3.x5[7].floating.n150 0.0557941
R16740 x2.x3.x5[7].floating.n150 x2.x3.x5[7].floating.n149 0.0557941
R16741 x2.x3.x5[7].floating.n149 x2.x3.x5[7].floating.n148 0.0557941
R16742 x2.x3.x5[7].floating.n148 x2.x3.x5[7].floating.n147 0.0557941
R16743 x2.x3.x5[7].floating.n61 x2.x3.x5[7].floating.n53 0.0557941
R16744 x2.x3.x5[7].floating.n62 x2.x3.x5[7].floating.n61 0.0557941
R16745 x2.x3.x5[7].floating.n63 x2.x3.x5[7].floating.n62 0.0557941
R16746 x2.x3.x5[7].floating.n64 x2.x3.x5[7].floating.n63 0.0557941
R16747 x2.x3.x5[7].floating.n33 x2.x3.x5[7].floating.n32 0.0557941
R16748 x2.x3.x5[7].floating.n34 x2.x3.x5[7].floating.n33 0.0557941
R16749 x2.x3.x5[7].floating.n35 x2.x3.x5[7].floating.n34 0.0557941
R16750 x2.x3.x5[7].floating.n36 x2.x3.x5[7].floating.n35 0.0557941
R16751 x2.x3.x5[7].floating.n40 x2.x3.x5[7].floating.n39 0.0557941
R16752 x2.x3.x5[7].floating.n41 x2.x3.x5[7].floating.n40 0.0557941
R16753 x2.x3.x5[7].floating.n42 x2.x3.x5[7].floating.n41 0.0557941
R16754 x2.x3.x5[7].floating.n43 x2.x3.x5[7].floating.n42 0.0557941
R16755 x2.x3.x5[7].floating.n20 x2.x3.x5[7].floating.n19 0.0557941
R16756 x2.x3.x5[7].floating.n21 x2.x3.x5[7].floating.n20 0.0557941
R16757 x2.x3.x5[7].floating.n22 x2.x3.x5[7].floating.n21 0.0557941
R16758 x2.x3.x5[7].floating.n23 x2.x3.x5[7].floating.n22 0.0557941
R16759 x2.x3.x5[7].floating.n169 x2.x3.x5[7].floating.n168 0.0557941
R16760 x2.x3.x5[7].floating.n168 x2.x3.x5[7].floating.n167 0.0557941
R16761 x2.x3.x5[7].floating.n167 x2.x3.x5[7].floating.n166 0.0557941
R16762 x2.x3.x5[7].floating.n57 x2.x3.x5[7].floating.n56 0.0557941
R16763 x2.x3.x5[7].floating.n58 x2.x3.x5[7].floating.n57 0.0557941
R16764 x2.x3.x5[7].floating.n59 x2.x3.x5[7].floating.n58 0.0557941
R16765 x2.x3.x5[7].floating.n60 x2.x3.x5[7].floating.n59 0.0557941
R16766 x2.x3.x5[7].floating.n143 x2.x3.x5[7].floating.n142 0.0557941
R16767 x2.x3.x5[7].floating.n142 x2.x3.x5[7].floating.n141 0.0557941
R16768 x2.x3.x5[7].floating.n141 x2.x3.x5[7].floating.n140 0.0557941
R16769 x2.x3.x5[7].floating.n132 x2.x3.x5[7].floating.n131 0.0557941
R16770 x2.x3.x5[7].floating.n131 x2.x3.x5[7].floating.n130 0.0557941
R16771 x2.x3.x5[7].floating.n130 x2.x3.x5[7].floating.n129 0.0557941
R16772 x2.x3.x5[7].floating.n129 x2.x3.x5[7].floating.n128 0.0557941
R16773 x2.x3.x5[7].floating.n125 x2.x3.x5[7].floating.n124 0.0557941
R16774 x2.x3.x5[7].floating.n124 x2.x3.x5[7].floating.n123 0.0557941
R16775 x2.x3.x5[7].floating.n123 x2.x3.x5[7].floating.n122 0.0557941
R16776 x2.x3.x5[7].floating.n16 x2.x3.x5[7].floating.n15 0.0537206
R16777 x2.x3.x5[7].floating.n162 x2.x3.x5[7].floating.n38 0.0537206
R16778 x2.x3.x5[7].floating.n136 x2.x3.x5[7].floating.n135 0.0537206
R16779 x2.x3.x5[7].floating.n118 x2.x3.x5[7].floating.n117 0.0537206
R16780 x2.x3.x5[7].floating.n15 x2.x3.x5[7].floating.n14 0.0530294
R16781 x2.x3.x5[7].floating.n163 x2.x3.x5[7].floating.n162 0.0530294
R16782 x2.x3.x5[7].floating.n137 x2.x3.x5[7].floating.n136 0.0530294
R16783 x2.x3.x5[7].floating.n119 x2.x3.x5[7].floating.n118 0.0530294
R16784 x2.x3.x5[7].floating.n105 x2.x3.x5[7].floating.n104 0.0529559
R16785 x2.x3.x5[7].floating.n75 x2.x3.x5[7].floating.n74 0.0529559
R16786 x2.x3.x5[7].floating.n1 x2.x3.x5[7].floating.n0 0.0529559
R16787 x2.x3.x5[7].floating.n161 x2.x3.x5[7].floating.n160 0.0529559
R16788 x2.x3.x5[7].floating.n104 x2.x3.x5[7].floating.n103 0.0524559
R16789 x2.x3.x5[7].floating.n74 x2.x3.x5[7].floating.n73 0.0524559
R16790 x2.x3.x5[7].floating.n161 x2.x3.x5[7].floating.n52 0.0524559
R16791 x2.x3.x5[7].floating.n2 x2.x3.x5[7].floating.n1 0.0524559
R16792 x2.x3.x5[7].floating.n166 x2.x3.x5[7].floating.n165 0.0523382
R16793 x2.x3.x5[7].floating.n140 x2.x3.x5[7].floating.n139 0.0523382
R16794 x2.x3.x5[7].floating.n122 x2.x3.x5[7].floating.n121 0.0523382
R16795 x2.x3.x5[7].floating.n19 x2.x3.x5[7].floating.n18 0.0516471
R16796 x2.x3.x5[7].floating.n56 x2.x3.x5[7].floating.n55 0.0516471
R16797 x2.x3.x5[7].floating.n133 x2.x3.x5[7].floating.n132 0.0516471
R16798 x2.x3.x5[7].floating x2.x3.x5[7].floating.n171 0.0495735
R16799 x2.x3.x5[7].floating.n145 x2.x3.x5[7].floating 0.0495735
R16800 x2.x3.x5[7].floating x2.x3.x5[7].floating.n127 0.0495735
R16801 x2.x3.x5[7].floating.n69 x2.x3.x5[7].floating.n66 0.0408846
R16802 x2.x3.x5[7].floating.n99 x2.x3.x5[7].floating.n96 0.0408846
R16803 x2.x3.x5[7].floating.n8 x2.x3.x5[7].floating.n5 0.0408846
R16804 x2.x3.x5[7].floating.n48 x2.x3.x5[7].floating.n45 0.0408846
R16805 x2.x3.x5[7].floating x2.x3.x5[7].floating.n169 0.0336765
R16806 x2.x3.x5[7].floating x2.x3.x5[7].floating.n143 0.0336765
R16807 x2.x3.x5[7].floating x2.x3.x5[7].floating.n125 0.0336765
R16808 x2.x3.x5[7].floating.n95 x2.x3.x5[7].floating.n94 0.0271618
R16809 x2.x3.x5[7].floating.n65 x2.x3.x5[7].floating.n64 0.0271618
R16810 x2.x3.x5[7].floating.n44 x2.x3.x5[7].floating.n43 0.0271618
R16811 x2.x3.x5[7].floating.n84 x2.x3.x5[7].floating.n83 0.0266618
R16812 x2.x3.x5[7].floating.n152 x2.x3.x5[7].floating.n151 0.0266618
R16813 x2.x3.x5[7].floating.n32 x2.x3.x5[7].floating.n31 0.0266618
R16814 x2.x3.x5[7].floating x2.x3.x5[7].floating.n23 0.0226176
R16815 x2.x3.x5[7].floating.n170 x2.x3.x5[7].floating 0.0226176
R16816 x2.x3.x5[7].floating x2.x3.x5[7].floating.n60 0.0226176
R16817 x2.x3.x5[7].floating.n144 x2.x3.x5[7].floating 0.0226176
R16818 x2.x3.x5[7].floating.n128 x2.x3.x5[7].floating 0.0226176
R16819 x2.x3.x5[7].floating.n126 x2.x3.x5[7].floating 0.0226176
R16820 x2.x3.x5[7].floating.n14 x2.x3.x5[7].floating.n13 0.0191618
R16821 x2.x3.x5[7].floating.n164 x2.x3.x5[7].floating.n163 0.0191618
R16822 x2.x3.x5[7].floating.n138 x2.x3.x5[7].floating.n137 0.0191618
R16823 x2.x3.x5[7].floating.n120 x2.x3.x5[7].floating.n119 0.0191618
R16824 x2.x3.x5[7].floating.n17 x2.x3.x5[7].floating.n16 0.0184706
R16825 x2.x3.x5[7].floating.n54 x2.x3.x5[7].floating.n38 0.0184706
R16826 x2.x3.x5[7].floating.n135 x2.x3.x5[7].floating.n134 0.0184706
R16827 x2.x3.x5[7].floating.n117 x2.x3.x5[7].floating.n116 0.0184706
R16828 x2.x3.x5[7].floating.n113 x2.x3.x5[7].floating.n112 0.014
R16829 x2.x3.x5[7].floating.n103 x2.x3.x5[7].floating.n102 0.014
R16830 x2.x3.x5[7].floating.n83 x2.x3.x5[7].floating.n82 0.014
R16831 x2.x3.x5[7].floating.n73 x2.x3.x5[7].floating.n72 0.014
R16832 x2.x3.x5[7].floating.n52 x2.x3.x5[7].floating.n51 0.014
R16833 x2.x3.x5[7].floating.n31 x2.x3.x5[7].floating.n30 0.014
R16834 x2.x3.x5[7].floating.n3 x2.x3.x5[7].floating.n2 0.014
R16835 x2.x3.x5[7].floating.n157 x2.x3.x5[7].floating.n152 0.014
R16836 x2.x3.x5[7].floating.n106 x2.x3.x5[7].floating.n105 0.0135
R16837 x2.x3.x5[7].floating.n100 x2.x3.x5[7].floating.n95 0.0135
R16838 x2.x3.x5[7].floating.n76 x2.x3.x5[7].floating.n75 0.0135
R16839 x2.x3.x5[7].floating.n70 x2.x3.x5[7].floating.n65 0.0135
R16840 x2.x3.x5[7].floating.n49 x2.x3.x5[7].floating.n44 0.0135
R16841 x2.x3.x5[7].floating.n10 x2.x3.x5[7].floating.n9 0.0135
R16842 x2.x3.x5[7].floating.n160 x2.x3.x5[7].floating.n159 0.0135
R16843 x2.x3.x5[7].floating.n81 x2.x3.x5[7].floating.n78 0.0101154
R16844 x2.x3.x5[7].floating.n111 x2.x3.x5[7].floating.n108 0.0101154
R16845 x2.x3.x5[7].floating.n29 x2.x3.x5[7].floating.n26 0.0101154
R16846 x2.x3.x5[7].floating.n156 x2.x3.x5[7].floating.n153 0.0101154
R16847 x2.x3.x5[7].floating.n18 x2.x3.x5[7].floating.n17 0.00464706
R16848 x2.x3.x5[7].floating.n55 x2.x3.x5[7].floating.n54 0.00464706
R16849 x2.x3.x5[7].floating.n134 x2.x3.x5[7].floating.n133 0.00464706
R16850 x2.x3.x5[7].floating.n116 x2.x3.x5[7].floating.n115 0.00464706
R16851 x2.x3.x5[7].floating.n13 x2.x3.x5[7].floating.n12 0.00395588
R16852 x2.x3.x5[7].floating.n165 x2.x3.x5[7].floating.n164 0.00395588
R16853 x2.x3.x5[7].floating.n139 x2.x3.x5[7].floating.n138 0.00395588
R16854 x2.x3.x5[7].floating.n121 x2.x3.x5[7].floating.n120 0.00395588
R16855 x2.x3.x5[7].floating.n107 x2.x3.x5[7].floating.n106 0.0035
R16856 x2.x3.x5[7].floating.n101 x2.x3.x5[7].floating.n100 0.0035
R16857 x2.x3.x5[7].floating.n77 x2.x3.x5[7].floating.n76 0.0035
R16858 x2.x3.x5[7].floating.n71 x2.x3.x5[7].floating.n70 0.0035
R16859 x2.x3.x5[7].floating.n50 x2.x3.x5[7].floating.n49 0.0035
R16860 x2.x3.x5[7].floating.n25 x2.x3.x5[7].floating.n24 0.0035
R16861 x2.x3.x5[7].floating.n9 x2.x3.x5[7].floating.n4 0.0035
R16862 x2.x3.x5[7].floating.n159 x2.x3.x5[7].floating.n158 0.0035
R16863 x2.x3.x5[7].floating.n112 x2.x3.x5[7].floating.n107 0.003
R16864 x2.x3.x5[7].floating.n102 x2.x3.x5[7].floating.n101 0.003
R16865 x2.x3.x5[7].floating.n82 x2.x3.x5[7].floating.n77 0.003
R16866 x2.x3.x5[7].floating.n72 x2.x3.x5[7].floating.n71 0.003
R16867 x2.x3.x5[7].floating.n51 x2.x3.x5[7].floating.n50 0.003
R16868 x2.x3.x5[7].floating.n30 x2.x3.x5[7].floating.n25 0.003
R16869 x2.x3.x5[7].floating.n4 x2.x3.x5[7].floating.n3 0.003
R16870 x2.x3.x5[7].floating.n158 x2.x3.x5[7].floating.n157 0.003
R16871 x2.x3.x5[7].floating.n155 x2.x3.x5[7].floating.n154 0.00260608
R16872 x2.x3.x5[7].floating.n80 x2.x3.x5[7].floating.n79 0.00260608
R16873 x2.x3.x5[7].floating.n110 x2.x3.x5[7].floating.n109 0.00260608
R16874 x2.x3.x5[7].floating.n28 x2.x3.x5[7].floating.n27 0.00260608
R16875 x2.x3.x5[7].floating.n68 x2.x3.x5[7].floating.n67 0.00177054
R16876 x2.x3.x5[7].floating.n98 x2.x3.x5[7].floating.n97 0.00177054
R16877 x2.x3.x5[7].floating.n7 x2.x3.x5[7].floating.n6 0.00177054
R16878 x2.x3.x5[7].floating.n47 x2.x3.x5[7].floating.n46 0.00177054
R16879 x2.x3.x5[7].floating.n69 x2.x3.x5[7].floating.n68 0.00174992
R16880 x2.x3.x5[7].floating.n99 x2.x3.x5[7].floating.n98 0.00174992
R16881 x2.x3.x5[7].floating.n8 x2.x3.x5[7].floating.n7 0.00174992
R16882 x2.x3.x5[7].floating.n48 x2.x3.x5[7].floating.n47 0.00174992
R16883 x2.x3.x5[7].floating.n156 x2.x3.x5[7].floating.n155 0.00101477
R16884 x2.x3.x5[7].floating.n81 x2.x3.x5[7].floating.n80 0.00101477
R16885 x2.x3.x5[7].floating.n111 x2.x3.x5[7].floating.n110 0.00101477
R16886 x2.x3.x5[7].floating.n29 x2.x3.x5[7].floating.n28 0.00101477
R16887 x2.x3.x5[7].floating.n112 x2.x3.x5[7].floating.n111 0.00053972
R16888 x2.x3.x5[7].floating.n100 x2.x3.x5[7].floating.n99 0.00053972
R16889 x2.x3.x5[7].floating.n82 x2.x3.x5[7].floating.n81 0.00053972
R16890 x2.x3.x5[7].floating.n70 x2.x3.x5[7].floating.n69 0.00053972
R16891 x2.x3.x5[7].floating.n49 x2.x3.x5[7].floating.n48 0.00053972
R16892 x2.x3.x5[7].floating.n30 x2.x3.x5[7].floating.n29 0.00053972
R16893 x2.x3.x5[7].floating.n9 x2.x3.x5[7].floating.n8 0.00053972
R16894 x2.x3.x5[7].floating.n157 x2.x3.x5[7].floating.n156 0.00053972
R16895 CAP_CTRL_CODE0[2] CAP_CTRL_CODE0[2].t2 140.387
R16896 CAP_CTRL_CODE0[2].n2 CAP_CTRL_CODE0[2].t3 140.34
R16897 CAP_CTRL_CODE0[2].n1 CAP_CTRL_CODE0[2].t0 140.34
R16898 CAP_CTRL_CODE0[2].n0 CAP_CTRL_CODE0[2].t1 140.34
R16899 CAP_CTRL_CODE0[2].n2 CAP_CTRL_CODE0[2] 2.82997
R16900 CAP_CTRL_CODE0[2].n1 CAP_CTRL_CODE0[2] 0.285826
R16901 CAP_CTRL_CODE0[2] CAP_CTRL_CODE0[2].n0 0.264087
R16902 CAP_CTRL_CODE0[2] CAP_CTRL_CODE0[2].n1 0.0466957
R16903 CAP_CTRL_CODE0[2].n0 CAP_CTRL_CODE0[2] 0.0466957
R16904 CAP_CTRL_CODE0[2] CAP_CTRL_CODE0[2].n2 0.00224038
R16905 reset.n0 reset.t0 230.499
R16906 reset.n0 reset.t1 157.826
R16907 reset.n1 reset.n0 8.91078
R16908 reset.n1 reset 2.92854
R16909 reset.n2 reset.n1 1.73973
R16910 reset.n2 reset 0.435954
R16911 reset reset.n2 0.00849921
R16912 CAP_CTRL_CODE2[2] CAP_CTRL_CODE2[2].t0 140.387
R16913 CAP_CTRL_CODE2[2].n2 CAP_CTRL_CODE2[2].t1 140.34
R16914 CAP_CTRL_CODE2[2].n0 CAP_CTRL_CODE2[2].t3 140.34
R16915 CAP_CTRL_CODE2[2].n1 CAP_CTRL_CODE2[2].t2 140.34
R16916 CAP_CTRL_CODE2[2] CAP_CTRL_CODE2[2].n1 2.87278
R16917 CAP_CTRL_CODE2[2] CAP_CTRL_CODE2[2].n0 0.285826
R16918 CAP_CTRL_CODE2[2].n2 CAP_CTRL_CODE2[2] 0.219989
R16919 CAP_CTRL_CODE2[2].n1 CAP_CTRL_CODE2[2] 0.0466957
R16920 CAP_CTRL_CODE2[2].n0 CAP_CTRL_CODE2[2] 0.0466957
R16921 CAP_CTRL_CODE2[2] CAP_CTRL_CODE2[2].n2 0.00192617
R16922 clk.n0 clk.t1 269.779
R16923 clk.n0 clk.t0 233.476
R16924 clk.n3 clk 10.4568
R16925 clk.n4 clk.n3 9.3005
R16926 clk.n1 clk.n0 7.17622
R16927 clk.n5 clk.n1 4.6438
R16928 clk.n3 clk 1.80332
R16929 clk clk.n2 1.08219
R16930 clk.n2 clk.n1 0.180782
R16931 clk clk.n5 0.0875115
R16932 clk.n5 clk.n4 0.0163608
R16933 CAP_CTRL_CODE1[1] CAP_CTRL_CODE1[1].t1 140.387
R16934 CAP_CTRL_CODE1[1].n0 CAP_CTRL_CODE1[1].t0 140.34
R16935 CAP_CTRL_CODE1[1].n0 CAP_CTRL_CODE1[1] 0.204269
R16936 CAP_CTRL_CODE1[1] CAP_CTRL_CODE1[1].n0 0.00197059
R16937 CAP_CTRL_CODE0[1] CAP_CTRL_CODE0[1].t0 140.387
R16938 CAP_CTRL_CODE0[1].n0 CAP_CTRL_CODE0[1].t1 140.34
R16939 CAP_CTRL_CODE0[1].n0 CAP_CTRL_CODE0[1] 0.204621
R16940 CAP_CTRL_CODE0[1] CAP_CTRL_CODE0[1].n0 0.00216406
R16941 CAP_CTRL_CODE2[1] CAP_CTRL_CODE2[1].t1 140.343
R16942 CAP_CTRL_CODE2[1].n0 CAP_CTRL_CODE2[1].t0 140.34
R16943 CAP_CTRL_CODE2[1] CAP_CTRL_CODE2[1].n0 0.247783
R16944 CAP_CTRL_CODE2[1].n0 CAP_CTRL_CODE2[1] 0.0466957
R16945 CAP_CTRL_CODE1[2] CAP_CTRL_CODE1[2].t1 140.387
R16946 CAP_CTRL_CODE1[2].n2 CAP_CTRL_CODE1[2].t3 140.34
R16947 CAP_CTRL_CODE1[2].n1 CAP_CTRL_CODE1[2].t2 140.34
R16948 CAP_CTRL_CODE1[2].n0 CAP_CTRL_CODE1[2].t0 140.34
R16949 CAP_CTRL_CODE1[2].n2 CAP_CTRL_CODE1[2] 2.82956
R16950 CAP_CTRL_CODE1[2].n1 CAP_CTRL_CODE1[2] 0.285826
R16951 CAP_CTRL_CODE1[2] CAP_CTRL_CODE1[2].n0 0.264087
R16952 CAP_CTRL_CODE1[2] CAP_CTRL_CODE1[2].n1 0.0466957
R16953 CAP_CTRL_CODE1[2].n0 CAP_CTRL_CODE1[2] 0.0466957
R16954 CAP_CTRL_CODE1[2] CAP_CTRL_CODE1[2].n2 0.00202988
R16955 CAP_CTRL_CODE2[0].n0 CAP_CTRL_CODE2[0].t0 140.34
R16956 CAP_CTRL_CODE2[0] CAP_CTRL_CODE2[0].n1 32.8219
R16957 CAP_CTRL_CODE2[0].n1 CAP_CTRL_CODE2[0] 4.5955
R16958 CAP_CTRL_CODE2[0].n1 CAP_CTRL_CODE2[0].n0 2.46566
R16959 CAP_CTRL_CODE2[0].n0 CAP_CTRL_CODE2[0] 0.0365169
R16960 set.n0 set.t1 228.9
R16961 set.n0 set.t0 159.406
R16962 set.n1 set.n0 8.47022
R16963 set.n1 set 3.68707
R16964 set set.n1 1.76402
R16965 CAP_CTRL_CODE2[3].n0 CAP_CTRL_CODE2[3].t1 229.964
R16966 CAP_CTRL_CODE2[3].n0 CAP_CTRL_CODE2[3].t0 158.363
R16967 CAP_CTRL_CODE2[3].n1 CAP_CTRL_CODE2[3].n0 8.13263
R16968 CAP_CTRL_CODE2[3].n1 CAP_CTRL_CODE2[3] 2.67916
R16969 CAP_CTRL_CODE2[3].n2 CAP_CTRL_CODE2[3] 2.1255
R16970 CAP_CTRL_CODE2[3] CAP_CTRL_CODE2[3].n1 1.84241
R16971 CAP_CTRL_CODE2[3].n2 CAP_CTRL_CODE2[3] 0.412265
R16972 CAP_CTRL_CODE2[3].n2 CAP_CTRL_CODE2[3] 0.271333
R16973 CAP_CTRL_CODE2[3] CAP_CTRL_CODE2[3].n2 0.0335882
R16974 CAP_CTRL_CODE3[1] CAP_CTRL_CODE3[1].t1 140.343
R16975 CAP_CTRL_CODE3[1].n0 CAP_CTRL_CODE3[1].t0 140.34
R16976 CAP_CTRL_CODE3[1] CAP_CTRL_CODE3[1].n0 0.247783
R16977 CAP_CTRL_CODE3[1].n0 CAP_CTRL_CODE3[1] 0.0466957
R16978 CAP_CTRL_CODE3[0].n0 CAP_CTRL_CODE3[0].t0 140.34
R16979 CAP_CTRL_CODE3[0] CAP_CTRL_CODE3[0].n0 2.45601
R16980 CAP_CTRL_CODE3[0].n0 CAP_CTRL_CODE3[0] 0.0365169
R16981 CAP_CTRL_CODE1[0] CAP_CTRL_CODE1[0].t0 140.376
R16982 CAP_CTRL_CODE1[0] CAP_CTRL_CODE1[0].n0 54.4514
R16983 CAP_CTRL_CODE1[0].n0 CAP_CTRL_CODE1[0] 4.7207
R16984 CAP_CTRL_CODE1[0].n0 CAP_CTRL_CODE1[0] 0.0117229
C0 a_11371_5318# CAP_CTRL_CODE1[2] 5.02e-19
C1 x2.x2.x5[7].floating a_10024_1818# 8.4e-20
C2 sample_delay_offset a_1870_6122# 3.45e-20
C3 x7.A a_4047_2819# 0.146f
C4 CAP_CTRL_CODE1[1] x2.x1.x2.floating 0.0027f
C5 x1.x3.Y x1.x4.Y 0.261f
C6 a_16686_3621# a_16686_3345# 0.0316f
C7 vdd a_2235_6116# 0.00381f
C8 vdd a_2678_2006# 0.708f
C9 x2.x1.x5[7].floating CAP_CTRL_CODE1[0] 0.00119f
C10 x2.x3.IN a_10065_3621# 5.05e-19
C11 sample_delay_offset a_10756_3022# 0.00652f
C12 x2.x3.x4[3].floating x2.x3.x10.Y 0.00668f
C13 CAP_CTRL_CODE2[1] x2.x2.x4[3].floating 0.00929f
C14 sample_delay_offset a_10112_1956# 6.38e-19
C15 a_4574_5732# a_4574_6008# 0.0316f
C16 a_4662_5456# CAP_CTRL_CODE0[2] 5.52e-19
C17 vdd a_2619_6316# 0.271f
C18 a_16686_3897# x2.x2.x6.SW 7.9e-20
C19 vdd x1.x2.D 1.22f
C20 x2.x4.x6.floating CAP_CTRL_CODE0[0] 1.18e-19
C21 x2.x1.x9.output_stack a_11283_6008# 0.0388f
C22 sample_delay_offset a_4047_3022# 8.56e-21
C23 sample_delay_offset a_11283_6008# 0.0189f
C24 x2.x3.x9.output_stack a_3056_2936# 1.29e-19
C25 x2.x4.x10.Y CAP_CTRL_CODE0[1] 6.94e-19
C26 x2.x1.IN CAP_CTRL_CODE1[0] 1.38e-19
C27 x2.x3.IN x2.x2.x10.Y 1.23e-19
C28 x2.x4.x9.output_stack x2.x4.x5[7].floating 1.19f
C29 a_10137_3759# CAP_CTRL_CODE2[0] 0.00672f
C30 vdd x2.x3.x2.floating 0.0335f
C31 vdd x3.Y 1.6f
C32 x2.x3.x7.floating CAP_CTRL_CODE2[2] 1.63e-20
C33 a_11371_5594# x2.x1.x7.floating 8.52e-19
C34 x2.x3.x3[1].floating CAP_CTRL_CODE2[1] 3.52e-20
C35 a_11283_5456# x2.x1.x4[3].floating 1.17e-19
C36 a_11283_5732# a_11283_5456# 0.0316f
C37 x2.x2.x10.Y x2.x2.IN 0.0967f
C38 x2.x4.x7.floating CAP_CTRL_CODE1[1] 1.73e-20
C39 a_10065_3897# x2.x3.x7.floating 8.52e-19
C40 reset a_1704_6122# 2.51e-21
C41 a_11283_5180# CAP_CTRL_CODE1[0] 6.54e-20
C42 a_10472_6534# x2.x1.x6.floating 0.0013f
C43 vdd CAP_CTRL_CODE1[3] 0.199f
C44 sample_delay_offset a_9977_3621# 0.0128f
C45 CAP_CTRL_CODE2[0] x2.x3.x4[3].floating 0.00915f
C46 x2.x4.x9.output_stack a_4574_6008# 0.0388f
C47 sample_delay_offset a_11371_5456# 0.00103f
C48 vdd a_3018_6116# 0.0036f
C49 x2.x3.x6.floating a_10112_2232# 0.00996f
C50 CAP_CTRL_CODE3[0] CAP_CTRL_CODE3[1] 0.465f
C51 x2.x3.x6.floating a_10756_2819# 0.0013f
C52 x2.x2.x4[3].floating x2.x2.x10.Y 0.00668f
C53 x2.x1.IN CAP_CTRL_CODE0[1] 5.47e-22
C54 x3.A sample_clk 9.97e-19
C55 x3.A x2.x4.x6.floating 0.0308f
C56 CAP_CTRL_CODE3[2] x2.x3.x2.floating 2.06e-20
C57 a_11371_5732# CAP_CTRL_CODE1[2] 1.7e-19
C58 a_10137_3207# x2.x3.x6.SW 0.00179f
C59 x2.x4.x6.SW x2.x4.x7.floating 9.72e-19
C60 CAP_CTRL_CODE0[0] x2.x4.x4[3].floating 8.34e-20
C61 a_10065_3345# CAP_CTRL_CODE2[0] 1.03e-19
C62 sample_delay_offset a_10065_3207# 0.00166f
C63 x2.x3.x9.output_stack a_10024_2094# 0.032f
C64 sample_delay_offset a_3813_6132# 0.00346f
C65 a_16846_4035# x2.x2.IN 0.029f
C66 x3.A x1.x4.Y 0.0439f
C67 a_2932_6494# a_2465_6482# 0.00316f
C68 a_2619_6316# a_3041_6494# 2.87e-21
C69 sample_delay_offset x2.x3.x10.Y 0.0402f
C70 a_4687_7121# x2.x4.x6.floating 0.0194f
C71 sample_delay_offset a_16846_3207# 0.0189f
C72 a_11308_7259# x2.x4.x5[7].floating 4.61e-19
C73 a_4662_5318# x2.x4.x7.floating 8.52e-19
C74 a_4574_5180# x2.x4.x4[3].floating 7.17e-20
C75 a_1704_6122# a_2151_6116# 0.14f
C76 a_1870_6122# a_2325_6090# 0.153f
C77 x2.x4.x10.Y x2.x4.x6.floating 0.0865f
C78 a_11308_6983# x2.x4.x5[7].floating 1.79e-19
C79 a_4599_7259# sample_delay_offset 6.38e-19
C80 x2.x3.x6.SW a_10112_1956# 9.98e-20
C81 a_11443_5870# a_11371_5870# 0.00227f
C82 a_16846_4035# x2.x2.x4[3].floating 7.17e-20
C83 x2.x4.x5[7].floating x2.x1.x6.floating 0.0269f
C84 x2.x1.x9.output_stack x2.x1.x7.floating 0.185f
C85 x3.Y a_4047_2819# 0.00933f
C86 a_11371_5180# CAP_CTRL_CODE1[2] 7.9e-19
C87 a_2678_2626# x2.x3.x5[7].floating 7.05e-19
C88 x2.x2.x5[7].floating a_10112_1680# 3.13e-19
C89 sample_delay_offset x1.x3.Y 2.41e-19
C90 a_10137_3483# a_10065_3483# 0.00227f
C91 vdd a_10112_2232# 0.11f
C92 vdd a_2790_6116# 0.0184f
C93 clk a_2058_6116# 6.72e-19
C94 sample_delay_offset x2.x1.x7.floating 0.259f
C95 sample_delay_offset CAP_CTRL_CODE2[0] 0.0609f
C96 vdd a_10756_2819# 0.21f
C97 sample_delay_offset a_4662_5870# 0.00138f
C98 a_4047_3022# CAP_CTRL_CODE3[0] 0.00169f
C99 CAP_CTRL_CODE2[1] x2.x2.x5[7].floating 0.0022f
C100 x2.x4.x5[7].floating x2.x4.x3[1].floating 0.8f
C101 a_4687_7397# x2.x4.x9.output_stack 1.5e-19
C102 x3.A x2.x4.x4[3].floating 6.65e-19
C103 a_16774_3621# x2.x2.IN 5.05e-19
C104 sample_delay_offset a_10024_1818# 1.9e-19
C105 x7.A x2.x3.x2.floating 0.0195f
C106 a_4734_5870# x2.x4.x7.floating 0.00959f
C107 a_10065_3483# x2.x2.x2.floating 2.21e-19
C108 vdd a_2932_6494# 0.186f
C109 x7.A x3.Y 0.00394f
C110 x2.x1.IN a_11443_5870# 0.0135f
C111 x2.x4.x6.SW x2.x4.x5[7].floating 0.00138f
C112 x3.A a_3553_3025# 2.66e-19
C113 a_4047_3022# x7.Y 0.00318f
C114 vdd x2.x1.x2.floating 0.0486f
C115 a_11443_5594# x2.x1.x6.SW 1.28e-19
C116 a_4599_7535# x2.x4.x5[7].floating 2.14e-19
C117 x2.x1.x10.Y CAP_CTRL_CODE1[2] 0.00201f
C118 CAP_CTRL_CODE1[2] x2.x1.x3[1].floating 0.00115f
C119 a_11371_6008# x2.x4.x2.floating 1.6e-19
C120 sample_delay_offset a_4662_6008# 0.00155f
C121 a_10137_4035# a_10137_3759# 0.0316f
C122 a_9977_3621# x2.x3.x6.SW 1.28e-19
C123 a_16846_4035# a_16774_4035# 0.00227f
C124 x2.x3.x9.output_stack CAP_CTRL_CODE3[1] 0.0715f
C125 sample_delay_offset CAP_CTRL_CODE0[0] 0.0313f
C126 a_11283_6008# a_11371_6146# 0.00227f
C127 vdd CAP_CTRL_CODE2[2] 0.0375f
C128 a_10137_3207# x2.x2.x9.output_stack 5.22e-20
C129 a_4734_5594# a_4662_5594# 0.00227f
C130 a_10472_6193# CAP_CTRL_CODE1[0] 8.82e-21
C131 x2.x4.x6.SW a_4574_6008# 0.00179f
C132 a_16846_3207# x2.x2.x7.floating 0.00409f
C133 x2.x4.x10.Y x2.x4.x4[3].floating 0.00668f
C134 a_10137_4035# x2.x3.x4[3].floating 7.17e-20
C135 a_16774_3345# a_16846_3207# 0.00227f
C136 a_10137_3207# x2.x3.x9.output_stack 0.0388f
C137 a_17181_6534# x2.x1.x5[7].floating 0.0132f
C138 sample_delay_offset a_16686_3621# 0.0132f
C139 x2.x4.x9.output_stack a_11283_6008# 5.22e-20
C140 a_4662_5732# x2.x4.x7.floating 8.52e-19
C141 sample_delay_offset a_4574_5180# 0.0025f
C142 vdd a_10472_6534# 0.211f
C143 x2.x3.IN x2.x3.x5[7].floating 0.00127f
C144 x2.x2.x3[1].floating x2.x2.x4[3].floating 1.19f
C145 x2.x1.x10.Y x2.x1.x3[1].floating 0.00302f
C146 x2.x3.x4[3].floating CAP_CTRL_CODE2[1] 7.03e-20
C147 vdd x2.x4.x7.floating 0.0369f
C148 x2.x3.x6.floating a_10024_2094# 0.0194f
C149 x2.x2.x10.Y a_16821_2232# 0.039f
C150 a_1870_6122# a_2058_6116# 0.163f
C151 x2.x2.x10.Y x2.x2.x5[7].floating 1.01f
C152 x2.x1.IN a_11371_5594# 3.4e-19
C153 x2.x2.x9.output_stack a_10756_3022# 0.00892f
C154 x2.x3.x10.Y x2.x3.x6.SW 0.788f
C155 vdd a_3056_2936# 0.614f
C156 CAP_CTRL_CODE3[0] x2.x3.x10.Y 0.0124f
C157 CAP_CTRL_CODE3[2] CAP_CTRL_CODE2[2] 7.54e-19
C158 a_11283_5456# x2.x4.x2.floating 0.00177f
C159 a_9977_3621# a_10065_3759# 0.00227f
C160 a_16846_3759# a_16686_3621# 0.0388f
C161 CAP_CTRL_CODE0[1] a_10472_6193# 3.4e-20
C162 x2.x3.IN a_10065_4035# 1.8e-19
C163 a_16846_3207# a_16774_3207# 0.00227f
C164 x2.x3.x9.output_stack a_10756_3022# 6.54e-19
C165 a_11371_5456# a_11443_5318# 0.00227f
C166 a_4734_5318# a_4574_5180# 0.0388f
C167 CAP_CTRL_CODE2[2] x2.x2.x2.floating 1.63e-20
C168 x3.A sample_delay_offset 0.343f
C169 x7.Y x2.x3.x10.Y 3.72e-20
C170 a_1704_6122# a_2569_6116# 0.00114f
C171 a_3106_6090# a_3222_6482# 0.0397f
C172 a_2932_6494# a_3041_6494# 0.00707f
C173 x1.x2.D a_2235_6116# 0.00271f
C174 a_16686_3897# x2.x2.x6.floating 0.00109f
C175 x2.x3.x5[7].floating a_3056_2150# 0.00132f
C176 a_4662_5870# CAP_CTRL_CODE0[2] 1.81e-19
C177 a_10137_3207# x2.x3.x7.floating 0.00409f
C178 a_10065_3897# x2.x2.x2.floating 2.21e-19
C179 x3.A a_4662_6146# 0.00225f
C180 a_11396_7121# x2.x4.x5[7].floating 4.88e-20
C181 a_11308_7535# x2.x1.x5[7].floating 2.14e-19
C182 a_4599_6983# x2.x4.x6.floating 0.00996f
C183 x2.x3.x9.output_stack a_4047_3022# 0.00892f
C184 a_4734_5870# a_4574_6008# 0.0388f
C185 a_2151_6116# a_3106_6090# 4.7e-22
C186 a_2325_6090# x1.x3.Y 0.192f
C187 a_1704_6122# a_3106_6090# 0.0492f
C188 x1.x2.D a_2619_6316# 0.177f
C189 x3.Y a_2678_2006# 0.00253f
C190 a_2678_2626# a_3056_2150# 9.31e-20
C191 x2.x4.x9.output_stack a_3813_6132# 1.59e-19
C192 a_4687_7121# sample_delay_offset 3.64e-19
C193 CAP_CTRL_CODE2[0] x2.x3.x6.SW 3.98e-21
C194 CAP_CTRL_CODE3[0] CAP_CTRL_CODE2[0] 1.74e-20
C195 CAP_CTRL_CODE1[3] x2.x1.x10.Y 0.0519f
C196 CAP_CTRL_CODE0[2] a_4662_6008# 1.36e-19
C197 a_4574_5732# a_4662_5870# 0.00227f
C198 a_16686_3621# x2.x2.x7.floating 0.00959f
C199 x3.A a_4734_5318# 0.014f
C200 a_4734_5594# x2.x4.x6.floating 0.00167f
C201 CAP_CTRL_CODE0[2] CAP_CTRL_CODE0[0] 7.44e-20
C202 sample_delay_offset x2.x4.x10.Y 0.0403f
C203 x2.x3.x3[1].floating x2.x3.x5[7].floating 0.8f
C204 vdd set 0.125f
C205 a_9977_3621# x2.x3.x9.output_stack 1.74e-19
C206 a_4599_7535# a_4687_7397# 0.0704f
C207 x2.x1.IN a_11308_7535# 0.00832f
C208 a_10756_3022# x2.x3.x7.floating 7.29e-19
C209 sample_delay_offset a_10137_4035# 0.00246f
C210 x2.x1.x9.output_stack x2.x1.x5[7].floating 1.19f
C211 vdd a_10024_2094# 0.0801f
C212 x2.x3.IN a_9977_3345# 0.0135f
C213 vdd x2.x4.x5[7].floating 44f
C214 sample_delay_offset a_11371_5870# 0.00138f
C215 sample_delay_offset x2.x1.x5[7].floating 0.00308f
C216 x2.x1.x7.floating a_11371_6146# 8.52e-19
C217 x2.x1.x4[3].floating a_11283_6008# 1.17e-19
C218 sample_delay_offset a_10112_1680# 3.28e-19
C219 a_11283_5732# a_11283_6008# 0.0316f
C220 a_4574_5180# CAP_CTRL_CODE0[2] 0.0177f
C221 x3.Y x2.x3.x2.floating 3.67e-19
C222 sample_delay_offset CAP_CTRL_CODE2[1] 0.0313f
C223 a_1704_6122# a_3340_6116# 1.25e-19
C224 vdd a_4574_6008# 0.0171f
C225 a_2619_6316# a_3018_6116# 3.13e-19
C226 x2.x4.x9.output_stack x1.x3.Y 1.29e-20
C227 x1.x2.D a_3018_6116# 0.00218f
C228 x2.x2.x9.output_stack x2.x3.x10.Y 1.93e-19
C229 x2.x4.x9.output_stack x2.x1.x7.floating 3.32e-19
C230 a_11371_6008# CAP_CTRL_CODE1[2] 1.01e-19
C231 a_9977_3897# a_10065_3897# 0.00227f
C232 x2.x1.IN x2.x1.x9.output_stack 0.371f
C233 x2.x4.x5[7].floating x2.x4.x2.floating 0.441f
C234 a_10065_3759# CAP_CTRL_CODE2[0] 2.39e-19
C235 x2.x3.x9.output_stack a_10065_3207# 0.00227f
C236 a_16846_3207# x2.x2.x9.output_stack 0.0388f
C237 a_3056_2936# a_4047_2819# 3.92e-21
C238 a_11443_5318# x2.x1.x7.floating 0.00925f
C239 x2.x1.IN sample_delay_offset 0.258f
C240 a_4574_5180# CAP_CTRL_CODE3[0] 1.29e-20
C241 x2.x3.x9.output_stack x2.x3.x10.Y 1.01f
C242 a_9977_3621# x2.x3.x7.floating 0.00959f
C243 reset x1.x4.Y 0.0529f
C244 x2.x3.IN CAP_CTRL_CODE1[0] 6.06e-20
C245 x3.A CAP_CTRL_CODE0[2] 0.0143f
C246 sample_delay_offset a_10065_3621# 0.00122f
C247 a_4734_5594# x2.x4.x4[3].floating 8.29e-19
C248 sample_delay_offset a_11283_5180# 0.0025f
C249 x2.x2.x4[3].floating x2.x2.IN 6.65e-19
C250 x2.x4.x9.output_stack CAP_CTRL_CODE0[0] 0.0321f
C251 x2.x2.IN CAP_CTRL_CODE1[0] 0.0555f
C252 x7.A a_3056_2936# 0.00243f
C253 x2.x2.x3[1].floating x2.x2.x5[7].floating 0.8f
C254 vdd clk 0.129f
C255 a_1870_6122# a_2465_6482# 0.00118f
C256 x1.x3.Y a_2058_6116# 0.0013f
C257 x2.x2.x10.Y a_16733_2094# 4.2e-19
C258 x2.x3.x6.floating a_10112_1956# 0.00996f
C259 x3.A a_2325_6090# 8.24e-20
C260 x2.x2.x9.output_stack CAP_CTRL_CODE2[0] 0.028f
C261 x3.A a_4574_5732# 0.0146f
C262 x3.A CAP_CTRL_CODE3[0] 0.00498f
C263 a_3222_6482# x2.x4.x6.floating 2.8e-20
C264 vdd CAP_CTRL_CODE3[1] 0.0182f
C265 a_11283_5456# CAP_CTRL_CODE1[2] 1.74e-19
C266 sample_delay_offset x2.x2.x10.Y 0.0403f
C267 a_10065_3207# x2.x3.x7.floating 8.52e-19
C268 x2.x3.x9.output_stack CAP_CTRL_CODE2[0] 0.0111f
C269 x2.x4.x10.Y CAP_CTRL_CODE0[2] 0.00203f
C270 x2.x1.x10.Y x2.x1.x2.floating 0.00202f
C271 x2.x3.x9.output_stack a_10024_1818# 1.5e-19
C272 x2.x3.x7.floating x2.x3.x10.Y 0.00345f
C273 x3.A x7.Y 0.0642f
C274 x2.x3.x5[7].floating sample_clk 2.13e-19
C275 x2.x1.x3[1].floating x2.x1.x2.floating 1.17f
C276 x1.x4.Y a_3222_6482# 3.78e-20
C277 x1.x2.D a_2790_6116# 0.00646f
C278 a_16774_4035# x2.x2.IN 1.8e-19
C279 a_2619_6316# a_2790_6116# 0.00652f
C280 x2.x4.x7.floating CAP_CTRL_CODE1[2] 1.87e-20
C281 vdd a_10137_3207# 0.00115f
C282 a_11396_7397# x2.x1.x5[7].floating 0.00154f
C283 x2.x4.x6.SW a_3813_6132# 7e-21
C284 a_11443_5870# x2.x1.x6.SW 2.44e-19
C285 CAP_CTRL_CODE1[1] x2.x1.x7.floating 1.73e-20
C286 a_2151_6116# x1.x4.Y 5.14e-19
C287 a_2619_6316# a_2932_6494# 0.119f
C288 a_1704_6122# x1.x4.Y 0.00163f
C289 x1.x2.D a_2932_6494# 0.0358f
C290 x2.x4.x10.Y a_4574_5732# 6.65e-20
C291 a_9977_3621# x2.x3.x6.floating 0.00167f
C292 a_16846_3759# x2.x2.x10.Y 4.07e-20
C293 a_2678_2626# sample_clk 0.109f
C294 vdd a_4687_7397# 0.134f
C295 a_10137_4035# x2.x3.x6.SW 3.1e-20
C296 a_4599_6983# sample_delay_offset 0.00273f
C297 x3.A x2.x4.x9.output_stack 0.371f
C298 a_10065_4173# CAP_CTRL_CODE2[0] 8.2e-19
C299 a_16686_3621# x2.x2.x9.output_stack 1.74e-19
C300 a_11283_5456# x2.x1.x10.Y 4.07e-20
C301 a_11283_5732# x2.x1.x7.floating 0.00409f
C302 x2.x1.x7.floating x2.x1.x4[3].floating 1.18f
C303 a_11443_5870# a_11443_5594# 0.0316f
C304 x2.x3.x6.SW a_10112_1680# 5.11e-20
C305 CAP_CTRL_CODE3[1] CAP_CTRL_CODE3[2] 0.889f
C306 x2.x1.x6.floating x2.x1.x7.floating 0.202f
C307 vdd a_1870_6122# 0.303f
C308 x2.x1.x10.Y a_10472_6534# 6.93e-19
C309 a_4599_7259# x2.x4.x6.SW 9.98e-20
C310 a_16846_3483# a_16774_3483# 0.00227f
C311 vdd a_10756_3022# 0.235f
C312 x2.x1.IN a_11396_7397# 0.00847f
C313 a_4599_7535# a_4599_7259# 0.0316f
C314 CAP_CTRL_CODE2[0] x2.x3.x7.floating 0.0075f
C315 a_10137_3483# a_10137_3207# 0.0316f
C316 CAP_CTRL_CODE3[0] CAP_CTRL_CODE2[1] 1.6e-20
C317 sample_delay_offset a_16846_4035# 0.00232f
C318 CAP_CTRL_CODE0[1] CAP_CTRL_CODE1[0] 2.91e-20
C319 CAP_CTRL_CODE0[0] CAP_CTRL_CODE1[1] 1.58e-20
C320 vdd a_10112_1956# 0.0945f
C321 sample_delay_offset a_4734_5594# 0.0133f
C322 a_4687_7121# x2.x4.x9.output_stack 0.032f
C323 a_16686_3345# x2.x2.IN 0.0166f
C324 x2.x3.x2.floating CAP_CTRL_CODE2[2] 1.63e-20
C325 vdd a_4047_3022# 0.236f
C326 a_11283_5732# CAP_CTRL_CODE0[0] 0.00654f
C327 a_10137_3207# x2.x2.x2.floating 8.75e-19
C328 x2.x2.x7.floating x2.x2.x10.Y 0.00345f
C329 x2.x4.x10.Y x2.x4.x9.output_stack 1.01f
C330 x2.x3.x10.Y x2.x3.x6.floating 0.0881f
C331 a_3056_2936# a_2678_2006# 9.31e-20
C332 x1.x2.D x2.x4.x7.floating 6.71e-19
C333 a_2932_6494# a_3018_6116# 0.00976f
C334 x2.x3.x4[3].floating x2.x3.x5[7].floating 1.55f
C335 a_3106_6090# a_3340_6116# 0.00945f
C336 a_2619_6316# x2.x4.x7.floating 1.58e-19
C337 vdd a_11283_6008# 0.00115f
C338 a_4574_5180# CAP_CTRL_CODE1[1] 8.94e-20
C339 a_2058_6116# a_2259_6494# 3.67e-19
C340 a_16846_4035# a_16846_3759# 0.0316f
C341 CAP_CTRL_CODE0[0] x2.x4.x3[1].floating 0.0424f
C342 x2.x4.x5[7].floating CAP_CTRL_CODE1[2] 3.3e-21
C343 a_4734_5870# a_3813_6132# 1.39e-21
C344 x2.x1.x9.output_stack a_10472_6193# 6.54e-19
C345 a_11443_5594# a_11371_5594# 0.00227f
C346 a_4734_5594# a_4734_5318# 0.0316f
C347 x3.A x2.x3.x9.output_stack 0.00106f
C348 x2.x4.x9.output_stack CAP_CTRL_CODE2[1] 9.58e-22
C349 a_16686_3345# x2.x2.x4[3].floating 8.29e-19
C350 x2.x4.x6.SW CAP_CTRL_CODE0[0] 4.21e-21
C351 x2.x1.IN a_11371_6146# 0.00196f
C352 x2.x3.IN x2.x2.x5[7].floating 0.0216f
C353 sample_delay_offset a_10472_6193# 0.00651f
C354 sample_delay_offset a_16774_3621# 0.00123f
C355 a_16821_2232# x2.x2.IN 0.0175f
C356 CAP_CTRL_CODE1[3] a_10472_6534# 0.00241f
C357 x2.x2.x5[7].floating x2.x2.IN 0.00127f
C358 x2.x4.x2.floating a_11283_6008# 8.75e-19
C359 a_10756_3022# x2.x2.x2.floating 0.0104f
C360 a_4574_5456# x2.x4.x7.floating 0.00409f
C361 sample_delay_offset a_4662_5180# 5.69e-19
C362 a_3056_2936# x2.x3.x2.floating 4.15e-20
C363 x3.Y a_3056_2936# 0.0957f
C364 a_2678_2626# a_3553_3025# 6.88e-22
C365 x7.A CAP_CTRL_CODE3[1] 5.47e-22
C366 x2.x3.x6.SW x2.x2.x10.Y 1.5e-20
C367 a_4047_3022# CAP_CTRL_CODE3[2] 1.69e-21
C368 x3.A CAP_CTRL_CODE1[1] 0.0017f
C369 CAP_CTRL_CODE2[0] x2.x3.x6.floating 1.3e-21
C370 x2.x1.IN x2.x4.x9.output_stack 0.127f
C371 x1.x3.Y a_2465_6482# 0.0351f
C372 x2.x2.x10.Y a_16821_1956# 2.35e-19
C373 a_16846_3207# x2.x2.x6.SW 0.00179f
C374 a_2325_6090# a_2837_6438# 9.75e-19
C375 x2.x3.x6.floating a_10024_1818# 0.0191f
C376 x2.x4.x6.SW a_4574_5180# 3.1e-20
C377 sample_delay_offset x2.x2.x3[1].floating 7.23e-20
C378 x2.x1.x10.Y x2.x4.x5[7].floating 0.00422f
C379 x2.x2.IN a_17181_6193# 0.244f
C380 x2.x1.IN a_11443_5318# 0.0135f
C381 a_16846_4035# x2.x2.x7.floating 0.00218f
C382 a_11371_5456# x2.x4.x2.floating 2.21e-19
C383 vdd a_10065_3207# 1.29e-19
C384 a_9977_3621# a_10137_3483# 0.0388f
C385 a_4734_5870# a_4662_5870# 0.00227f
C386 x2.x2.x9.output_stack CAP_CTRL_CODE2[1] 0.0705f
C387 a_16686_3621# a_16774_3759# 0.00227f
C388 vdd a_3813_6132# 0.194f
C389 a_11308_7535# x2.x1.x6.SW 5.11e-20
C390 x2.x2.x4[3].floating x2.x2.x5[7].floating 1.55f
C391 x2.x3.IN a_10137_3759# 0.0136f
C392 vdd x2.x3.x10.Y 2.73f
C393 a_11443_5318# a_11283_5180# 0.0388f
C394 a_4574_5180# a_4662_5318# 0.00227f
C395 sample_delay_offset a_3222_6482# 5.28e-19
C396 x1.x4.Y a_2569_6116# 2.07e-19
C397 a_2932_6494# a_2790_6116# 0.00412f
C398 a_3106_6090# x2.x4.x6.floating 1.28e-19
C399 x2.x3.x9.output_stack CAP_CTRL_CODE2[1] 4.73e-20
C400 vdd a_16846_3207# 0.00163f
C401 a_9977_3345# x2.x3.x4[3].floating 8.29e-19
C402 a_9977_3621# x2.x2.x2.floating 6.88e-19
C403 x2.x3.IN x2.x3.x4[3].floating 6.65e-19
C404 a_11308_7259# x2.x1.x5[7].floating 2.76e-19
C405 a_10137_4035# CAP_CTRL_CODE1[1] 2.46e-20
C406 x3.A x2.x4.x6.SW 0.0928f
C407 sample_delay_offset a_1704_6122# 6.22e-19
C408 a_17181_6534# x2.x2.IN 0.145f
C409 CAP_CTRL_CODE1[0] a_17181_6193# 0.00169f
C410 a_4734_5870# a_4662_6008# 0.00227f
C411 sample_delay_offset x2.x3.x5[7].floating 0.00308f
C412 x3.A a_4599_7535# 0.00832f
C413 a_4047_3022# a_4047_2819# 0.0121f
C414 a_3106_6090# x1.x4.Y 0.117f
C415 vdd a_4599_7259# 0.0712f
C416 x2.x1.x5[7].floating CAP_CTRL_CODE1[1] 0.0022f
C417 x2.x1.x6.SW x2.x1.x9.output_stack 0.164f
C418 a_2619_6316# a_4574_6008# 1.75e-20
C419 a_10065_4173# a_10137_4035# 0.0022f
C420 x1.x2.D a_4574_6008# 9.67e-19
C421 a_11308_6983# x2.x1.x5[7].floating 2.76e-19
C422 sample_delay_offset x2.x1.x6.SW 0.19f
C423 a_11283_5732# a_11371_5870# 0.00227f
C424 a_4574_5732# a_4734_5594# 0.0388f
C425 x2.x1.x5[7].floating x2.x1.x4[3].floating 1.55f
C426 x2.x4.x10.Y x2.x4.x3[1].floating 0.00302f
C427 x3.A a_4662_5318# 5.17e-19
C428 vdd x1.x3.Y 0.834f
C429 a_16774_3621# x2.x2.x7.floating 8.52e-19
C430 a_10137_3483# x2.x3.x10.Y 6.65e-20
C431 a_4047_3022# x7.A 0.151f
C432 x2.x1.x6.floating x2.x1.x5[7].floating 1.18f
C433 x2.x4.x6.floating CAP_CTRL_CODE0[1] 1.27e-19
C434 a_10137_4035# x2.x3.x7.floating 0.00218f
C435 CAP_CTRL_CODE1[3] x2.x4.x5[7].floating 0.00291f
C436 a_11443_5594# x2.x1.x9.output_stack 1.74e-19
C437 vdd CAP_CTRL_CODE2[0] 0.00338f
C438 vdd x2.x1.x7.floating 0.0315f
C439 a_9977_3345# a_10065_3345# 0.00227f
C440 CAP_CTRL_CODE3[2] x2.x3.x10.Y 0.00203f
C441 x2.x3.x5[7].floating sample_clk_b 2.37e-19
C442 x2.x1.IN a_11308_7259# 0.00866f
C443 sample_delay_offset a_10065_4035# 9.64e-19
C444 a_10065_3207# x2.x2.x2.floating 2.02e-19
C445 x2.x3.IN a_10065_3345# 0.0013f
C446 vdd a_10024_1818# 0.138f
C447 sample_delay_offset a_11443_5594# 0.0133f
C448 x2.x1.IN CAP_CTRL_CODE1[1] 1.86e-19
C449 x2.x4.x10.Y x2.x4.x6.SW 0.788f
C450 a_4599_6983# x2.x4.x9.output_stack 0.0702f
C451 a_4599_7535# x2.x4.x10.Y 1.02e-19
C452 x2.x1.IN a_11308_6983# 0.0175f
C453 x2.x3.x7.floating CAP_CTRL_CODE2[1] 1.76e-20
C454 x2.x2.x9.output_stack x2.x2.x10.Y 1.01f
C455 a_4662_5180# CAP_CTRL_CODE0[2] 0.0013f
C456 a_16686_3621# x2.x2.x6.SW 1.28e-19
C457 x2.x4.x4[3].floating CAP_CTRL_CODE1[0] 6.43e-20
C458 clk a_2619_6316# 3.33e-20
C459 clk x1.x2.D 0.007f
C460 a_2678_2626# sample_clk_b 0.00102f
C461 x2.x1.IN x2.x1.x4[3].floating 6.65e-19
C462 x2.x1.IN a_11283_5732# 0.0136f
C463 vdd a_4662_6008# 9.37e-20
C464 x1.x4.Y a_3340_6116# 7.54e-19
C465 x2.x1.IN x2.x1.x6.floating 0.03f
C466 a_11283_5180# CAP_CTRL_CODE1[1] 8.94e-20
C467 vdd CAP_CTRL_CODE0[0] 0.00321f
C468 x3.A a_2465_6482# 6.9e-20
C469 x2.x4.x2.floating x2.x1.x7.floating 0.0475f
C470 a_3018_6116# a_4574_6008# 2.23e-20
C471 x2.x4.x9.output_stack a_4734_5594# 1.74e-19
C472 a_16686_3897# a_16774_3897# 0.00227f
C473 a_9977_3897# a_9977_3621# 0.0316f
C474 a_10137_3483# CAP_CTRL_CODE2[0] 0.00663f
C475 x3.A a_4734_5870# 0.014f
C476 a_11283_5180# x2.x1.x4[3].floating 7.17e-20
C477 a_4574_5456# a_4662_5456# 0.00227f
C478 a_11371_5318# x2.x1.x7.floating 8.52e-19
C479 x2.x3.x3[1].floating x2.x3.x4[3].floating 1.19f
C480 CAP_CTRL_CODE3[2] CAP_CTRL_CODE2[0] 2.26f
C481 a_10065_3621# x2.x3.x7.floating 8.52e-19
C482 x2.x3.x10.Y a_4047_2819# 0.00127f
C483 CAP_CTRL_CODE2[0] x2.x2.x2.floating 0.167f
C484 a_16733_2094# x2.x2.IN 0.00921f
C485 sample_delay_offset a_9977_3345# 0.015f
C486 CAP_CTRL_CODE1[2] a_11283_6008# 5.6e-20
C487 sample_delay_offset x2.x3.IN 0.258f
C488 CAP_CTRL_CODE3[1] x2.x3.x2.floating 0.00656f
C489 x2.x1.x9.output_stack x2.x2.IN 0.127f
C490 CAP_CTRL_CODE0[0] x2.x4.x2.floating 0.164f
C491 CAP_CTRL_CODE0[1] x2.x4.x4[3].floating 0.0296f
C492 sample_delay_offset x2.x2.IN 0.27f
C493 x1.x3.Y a_3041_6494# 7.87e-19
C494 x7.A x2.x3.x10.Y 1.13e-19
C495 x2.x3.x6.floating a_10112_1680# 0.00578f
C496 x2.x2.x10.Y a_16733_1818# 1.49e-19
C497 a_1870_6122# a_2235_6116# 4.45e-20
C498 x2.x4.x9.output_stack a_10472_6193# 0.00892f
C499 x3.A a_4662_5732# 6.73e-19
C500 a_10112_2232# a_10024_2094# 0.0704f
C501 a_11371_5456# CAP_CTRL_CODE1[2] 3.33e-19
C502 x2.x2.x5[7].floating a_16821_2232# 2.76e-19
C503 a_2325_6090# a_2151_6116# 0.205f
C504 a_1870_6122# a_2619_6316# 0.139f
C505 vdd x3.A 0.748f
C506 x1.x2.D a_1870_6122# 0.127f
C507 a_1704_6122# a_2325_6090# 0.111f
C508 x2.x3.x6.SW x2.x3.x5[7].floating 0.00138f
C509 x2.x1.x10.Y a_11283_6008# 1.69e-19
C510 a_4574_5180# CAP_CTRL_CODE3[2] 1.71e-20
C511 CAP_CTRL_CODE3[0] x2.x3.x5[7].floating 0.00121f
C512 x2.x1.x9.output_stack CAP_CTRL_CODE1[0] 0.0244f
C513 x1.x4.Y x2.x4.x6.floating 1.28e-20
C514 a_16846_3759# x2.x2.IN 0.0299f
C515 sample_delay_offset x2.x2.x4[3].floating 0.0137f
C516 sample_delay_offset CAP_CTRL_CODE1[0] 6.99f
C517 a_11396_7121# x2.x1.x5[7].floating 0.00169f
C518 sample_delay_offset a_3106_6090# 0.00255f
C519 x7.Y x2.x3.x5[7].floating 0.00134f
C520 vdd a_4687_7121# 0.0761f
C521 a_2932_6494# a_4574_6008# 3.99e-20
C522 reset a_2058_6116# 6.52e-19
C523 a_3056_2150# sample_clk_b 0.00457f
C524 a_11371_5732# x2.x1.x7.floating 8.52e-19
C525 vdd x2.x4.x10.Y 2.71f
C526 a_4047_3022# x2.x3.x2.floating 0.0104f
C527 sample_delay_offset x2.x3.x3[1].floating 4.68e-20
C528 a_16846_3759# x2.x2.x4[3].floating 1.17e-19
C529 x7.Y a_2678_2626# 1.93e-20
C530 a_4047_3022# x3.Y 0.00115f
C531 x3.A CAP_CTRL_CODE3[2] 0.00186f
C532 a_4599_6983# x2.x4.x6.SW 0.00707f
C533 a_1870_6122# a_3018_6116# 2.13e-19
C534 x2.x1.IN a_11396_7121# 0.00921f
C535 a_16846_3483# a_16846_3207# 0.0316f
C536 sample_delay_offset a_16774_4035# 9.67e-19
C537 x2.x2.x9.output_stack x2.x2.x3[1].floating 0.341f
C538 a_10472_6534# x2.x4.x5[7].floating 0.0132f
C539 x2.x2.x7.floating x2.x2.IN 0.0261f
C540 vdd x2.x1.x5[7].floating 44f
C541 vdd a_10112_1680# 0.171f
C542 sample_delay_offset a_4662_5594# 0.00111f
C543 x2.x4.x5[7].floating x2.x4.x7.floating 0.182f
C544 sample_delay_offset CAP_CTRL_CODE0[1] 0.029f
C545 a_16774_3345# x2.x2.IN 0.0013f
C546 vdd CAP_CTRL_CODE2[1] 0.0183f
C547 x2.x4.x9.output_stack x2.x1.x6.SW 3.62e-19
C548 a_10472_6193# CAP_CTRL_CODE1[1] 9.55e-21
C549 x2.x4.x6.SW a_4734_5594# 1.28e-19
C550 a_3553_3025# sample_clk 2.11e-20
C551 x2.x4.x10.Y x2.x4.x2.floating 0.00202f
C552 a_17181_6534# a_17181_6193# 0.0121f
C553 sample_delay_offset a_3340_6116# 3.81e-20
C554 a_11443_5318# x2.x1.x6.SW 7.9e-20
C555 CAP_CTRL_CODE1[2] x2.x1.x7.floating 0.0129f
C556 x3.A a_3041_6494# 3.6e-20
C557 a_2465_6482# a_2837_6438# 3.34e-19
C558 x2.x4.x7.floating a_4574_6008# 0.00409f
C559 a_11371_5870# x2.x4.x2.floating 2.21e-19
C560 a_9977_3345# x2.x3.x6.SW 2.44e-19
C561 vdd x2.x1.IN 0.613f
C562 x2.x3.IN x2.x3.x6.SW 0.0933f
C563 x2.x2.x4[3].floating x2.x2.x7.floating 1.18f
C564 a_11443_5594# a_11443_5318# 0.0316f
C565 x1.x2.D a_3813_6132# 0.183f
C566 a_2151_6116# a_2058_6116# 0.0367f
C567 a_2619_6316# a_3813_6132# 6.04e-19
C568 a_1704_6122# a_2058_6116# 0.0661f
C569 x3.A a_4047_2819# 3.02e-19
C570 x2.x4.x3[1].floating a_10472_6193# 3.09e-19
C571 x2.x2.x10.Y x2.x2.x6.SW 0.788f
C572 a_16774_3207# x2.x2.IN 0.00196f
C573 a_10137_3759# x2.x3.x4[3].floating 1.17e-19
C574 a_10137_4035# x2.x2.x2.floating 9.24e-19
C575 a_16821_1956# x2.x2.IN 0.00866f
C576 sample_delay_offset a_16686_3345# 0.0153f
C577 x3.A CAP_CTRL_CODE0[3] 6.16e-19
C578 CAP_CTRL_CODE3[2] CAP_CTRL_CODE2[1] 7.21e-19
C579 CAP_CTRL_CODE3[1] CAP_CTRL_CODE2[2] 2.96e-20
C580 a_4662_5456# x2.x4.x7.floating 8.52e-19
C581 x2.x3.x9.output_stack x2.x3.x5[7].floating 1.19f
C582 CAP_CTRL_CODE0[2] CAP_CTRL_CODE1[0] 5.83e-20
C583 CAP_CTRL_CODE0[0] CAP_CTRL_CODE1[2] 3.13f
C584 x2.x1.IN x2.x4.x2.floating 0.0257f
C585 x2.x3.x2.floating x2.x3.x10.Y 0.00202f
C586 CAP_CTRL_CODE2[1] x2.x2.x2.floating 0.00516f
C587 x2.x1.x10.Y x2.x1.x7.floating 0.00345f
C588 x3.Y x2.x3.x10.Y 1.94e-19
C589 x3.A x7.A 0.0116f
C590 a_1870_6122# a_2790_6116# 1.09e-19
C591 x1.x3.Y a_2235_6116# 5.36e-19
C592 x2.x2.x10.Y a_16821_1680# 1.02e-19
C593 a_2325_6090# a_2569_6116# 0.0104f
C594 x2.x1.IN a_11371_5318# 1.8e-19
C595 vdd x2.x2.x10.Y 2.71f
C596 a_16774_4035# x2.x2.x7.floating 8.52e-19
C597 x2.x3.x9.output_stack a_2678_2626# 1.57e-19
C598 a_10756_3022# a_10756_2819# 0.0121f
C599 a_11443_5870# x2.x1.x9.output_stack 0.032f
C600 a_4574_5180# CAP_CTRL_CODE1[2] 1.29e-19
C601 a_16821_2232# a_16733_2094# 0.0704f
C602 a_10112_2232# a_10112_1956# 0.0316f
C603 a_11283_5180# x2.x4.x2.floating 9.24e-19
C604 x2.x2.x5[7].floating a_16733_2094# 0.00169f
C605 a_10065_3621# a_10137_3483# 0.00227f
C606 a_4734_5870# a_4734_5594# 0.0316f
C607 a_16686_3621# a_16846_3483# 0.0388f
C608 a_1870_6122# a_2932_6494# 0.137f
C609 x1.x3.Y a_2619_6316# 0.0972f
C610 vdd a_2837_6438# 0.00126f
C611 a_11308_7259# x2.x1.x6.SW 9.98e-20
C612 x1.x2.D x1.x3.Y 0.0589f
C613 sample_delay_offset a_11443_5870# 0.0155f
C614 x2.x3.IN a_10065_3759# 3.4e-19
C615 a_11283_5180# a_11371_5318# 0.00227f
C616 CAP_CTRL_CODE0[3] x2.x4.x10.Y 0.0519f
C617 sample_delay_offset x2.x4.x6.floating 0.0683f
C618 sample_delay_offset a_16821_2232# 0.00273f
C619 a_11371_6008# a_11283_6008# 0.00227f
C620 sample_delay_offset x2.x2.x5[7].floating 0.00542f
C621 a_11308_6983# x2.x1.x6.SW 0.00707f
C622 a_16686_3621# x2.x2.x6.floating 0.00167f
C623 a_4662_5594# CAP_CTRL_CODE0[2] 3.62e-19
C624 a_10065_3621# x2.x2.x2.floating 2.21e-19
C625 a_16846_4035# x2.x2.x6.SW 3.1e-20
C626 CAP_CTRL_CODE0[2] CAP_CTRL_CODE0[1] 1.31f
C627 x2.x3.x7.floating x2.x3.x5[7].floating 0.182f
C628 x2.x1.x9.output_stack a_17181_6193# 0.00892f
C629 a_11283_5732# x2.x1.x6.SW 8.11e-20
C630 sample_delay_offset x1.x4.Y 0.00954f
C631 CAP_CTRL_CODE2[0] x2.x3.x2.floating 1.9e-20
C632 a_10756_3022# CAP_CTRL_CODE2[2] 8.96e-21
C633 CAP_CTRL_CODE3[0] x2.x3.x3[1].floating 0.0326f
C634 x2.x1.x6.SW x2.x1.x6.floating 0.13f
C635 vdd a_4599_6983# 0.106f
C636 sample_clk sample_clk_b 0.141f
C637 x1.x4.Y a_4662_6146# 2.16e-20
C638 a_10137_4035# a_9977_3897# 0.0388f
C639 a_16774_4173# a_16846_4035# 0.0022f
C640 x3.A CAP_CTRL_CODE1[2] 0.00176f
C641 a_11443_5594# x2.x1.x4[3].floating 8.29e-19
C642 x2.x3.IN x2.x2.x9.output_stack 0.127f
C643 a_4662_5732# a_4734_5594# 0.00227f
C644 a_11283_5732# a_11443_5594# 0.0388f
C645 a_4047_3022# CAP_CTRL_CODE2[2] 1.3e-21
C646 x2.x4.x9.output_stack CAP_CTRL_CODE1[0] 2.42e-20
C647 a_4734_5318# x2.x4.x6.floating 0.00109f
C648 a_11443_5594# x2.x1.x6.floating 0.00167f
C649 a_16686_3345# x2.x2.x7.floating 0.00959f
C650 vdd a_16846_4035# 4.84e-19
C651 x2.x2.x2.floating x2.x2.x10.Y 0.00202f
C652 a_10065_4035# x2.x3.x7.floating 8.52e-19
C653 x2.x2.x9.output_stack x2.x2.IN 0.371f
C654 set clk 0.00167f
C655 x2.x4.x9.output_stack a_3106_6090# 2.52e-19
C656 x1.x3.Y a_3018_6116# 2.23e-19
C657 a_16686_3345# a_16774_3345# 0.00227f
C658 a_9977_3345# x2.x3.x9.output_stack 0.032f
C659 sample_delay_offset a_10137_3759# 0.00294f
C660 x2.x3.IN x2.x3.x9.output_stack 0.371f
C661 sample_delay_offset a_11371_5594# 0.00111f
C662 x2.x1.x9.output_stack a_17181_6534# 0.00887f
C663 sample_delay_offset x2.x3.x4[3].floating 0.00736f
C664 x2.x4.x10.Y CAP_CTRL_CODE1[2] 2.74e-20
C665 x2.x1.IN a_11371_5732# 5.05e-19
C666 sample_delay_offset x2.x4.x4[3].floating 0.00732f
C667 x2.x3.IN CAP_CTRL_CODE1[1] 5.1e-20
C668 a_10137_4035# CAP_CTRL_CODE1[2] 2.07e-20
C669 a_11371_5870# CAP_CTRL_CODE1[2] 1.29e-19
C670 x2.x2.x9.output_stack x2.x2.x4[3].floating 0.636f
C671 a_16686_3897# a_16686_3621# 0.0316f
C672 x2.x3.x10.Y a_10112_2232# 0.039f
C673 x2.x2.x9.output_stack CAP_CTRL_CODE1[0] 4.11e-21
C674 x2.x2.IN CAP_CTRL_CODE1[1] 5.47e-22
C675 x2.x4.x9.output_stack CAP_CTRL_CODE0[1] 0.0744f
C676 x2.x3.x10.Y a_10756_2819# 6.93e-19
C677 a_4047_3022# a_3056_2936# 8.77e-20
C678 x2.x1.x5[7].floating CAP_CTRL_CODE1[2] 0.0056f
C679 x2.x3.x5[7].floating x2.x3.x6.floating 1.18f
C680 x2.x2.x7.floating x2.x2.x5[7].floating 0.182f
C681 x2.x3.IN a_10065_4173# 1.34e-19
C682 a_10065_3483# CAP_CTRL_CODE2[0] 1.32e-19
C683 a_4574_5456# a_4574_5180# 0.0316f
C684 a_11283_5456# a_11371_5456# 0.00227f
C685 vdd reset 0.105f
C686 vdd a_10472_6193# 0.235f
C687 a_2151_6116# a_2465_6482# 0.0258f
C688 x3.A a_2619_6316# 0.00211f
C689 a_1704_6122# a_2465_6482# 6.04e-20
C690 x3.A x1.x2.D 0.00992f
C691 x2.x4.x9.output_stack a_3340_6116# 6.72e-21
C692 x2.x3.x9.output_stack CAP_CTRL_CODE1[0] 4.11e-21
C693 a_9977_3345# x2.x3.x7.floating 0.00959f
C694 x2.x4.x6.floating CAP_CTRL_CODE0[2] 1.36e-19
C695 a_16733_1818# x2.x2.IN 0.00847f
C696 sample_delay_offset a_10065_3345# 0.00154f
C697 x2.x3.IN x2.x3.x7.floating 0.0242f
C698 a_4687_7397# x2.x4.x5[7].floating 0.00154f
C699 a_4734_5318# x2.x4.x4[3].floating 7.47e-19
C700 x2.x4.x10.Y x2.x1.x10.Y 1.79e-20
C701 x3.A x2.x3.x2.floating 0.00544f
C702 x3.A x3.Y 0.211f
C703 x2.x1.IN CAP_CTRL_CODE1[2] 0.0169f
C704 vdd x2.x2.x3[1].floating 0.0301f
C705 a_11308_7535# sample_delay_offset 3.28e-19
C706 CAP_CTRL_CODE1[1] CAP_CTRL_CODE1[0] 6.51f
C707 x1.x3.Y a_2790_6116# 0.0015f
C708 a_11371_6008# x2.x1.x7.floating 8.52e-19
C709 x2.x4.x2.floating a_10472_6193# 0.0104f
C710 x2.x1.x10.Y x2.x1.x5[7].floating 1.01f
C711 x2.x1.x5[7].floating x2.x1.x3[1].floating 0.8f
C712 x2.x3.x6.SW x2.x2.x5[7].floating 0.00313f
C713 x2.x1.IN a_11371_5180# 1.34e-19
C714 x3.A a_4574_5456# 0.0148f
C715 x2.x3.x9.output_stack x2.x3.x3[1].floating 0.341f
C716 a_4599_6983# CAP_CTRL_CODE0[3] 2.69e-19
C717 a_16821_2232# a_16821_1956# 0.0316f
C718 a_11283_5180# CAP_CTRL_CODE1[2] 0.00747f
C719 a_10024_2094# a_10112_1956# 0.0704f
C720 x2.x2.x5[7].floating a_16821_1956# 2.76e-19
C721 CAP_CTRL_CODE1[0] x2.x1.x4[3].floating 6.66e-20
C722 a_2325_6090# x1.x4.Y 0.00131f
C723 x1.x3.Y a_2932_6494# 0.162f
C724 vdd a_3222_6482# 0.00235f
C725 x7.Y sample_clk 9.3e-20
C726 a_1870_6122# a_4574_6008# 9.42e-21
C727 a_4574_5732# x1.x4.Y 0.00234f
C728 a_11283_5180# a_11371_5180# 0.0022f
C729 a_3813_6132# x2.x4.x7.floating 0.00173f
C730 sample_delay_offset a_16733_2094# 3.64e-19
C731 a_16774_3759# x2.x2.IN 3.4e-19
C732 x2.x4.x3[1].floating CAP_CTRL_CODE1[0] 3.21e-20
C733 sample_delay_offset x2.x1.x9.output_stack 0.262f
C734 vdd a_2151_6116# 0.182f
C735 x2.x1.IN x2.x1.x10.Y 0.0967f
C736 vdd x2.x3.x5[7].floating 44f
C737 vdd a_1704_6122# 0.595f
C738 CAP_CTRL_CODE2[0] CAP_CTRL_CODE2[2] 1.48e-20
C739 x2.x4.x10.Y a_4574_5456# 4.07e-20
C740 sample_delay_offset a_4662_6146# 0.00167f
C741 a_16846_3483# x2.x2.x10.Y 6.65e-20
C742 CAP_CTRL_CODE0[1] CAP_CTRL_CODE1[1] 3.15e-20
C743 a_9977_3345# x2.x3.x6.floating 0.00278f
C744 CAP_CTRL_CODE0[2] x2.x4.x4[3].floating 0.532f
C745 a_10137_3759# x2.x3.x6.SW 4.74e-20
C746 x2.x3.IN x2.x3.x6.floating 0.03f
C747 x2.x4.x9.output_stack x2.x4.x6.floating 0.229f
C748 a_11283_5180# x2.x1.x10.Y 2.2e-20
C749 vdd x2.x1.x6.SW 0.452f
C750 a_10065_3897# CAP_CTRL_CODE2[0] 3.43e-19
C751 x2.x2.x2.floating x2.x2.x3[1].floating 1.17f
C752 a_16686_3345# x2.x2.x9.output_stack 0.032f
C753 vdd a_2678_2626# 0.7f
C754 a_11283_5456# x2.x1.x7.floating 0.00409f
C755 x2.x3.x2.floating CAP_CTRL_CODE2[1] 1.76e-20
C756 x2.x2.x10.Y x2.x2.x6.floating 0.0881f
C757 clk a_1870_6122# 0.00626f
C758 x2.x4.x9.output_stack x1.x4.Y 4.23e-20
C759 sample_delay_offset a_16846_3759# 0.00298f
C760 a_4574_5732# x2.x4.x4[3].floating 1.17e-19
C761 a_4662_5870# x2.x4.x7.floating 8.52e-19
C762 CAP_CTRL_CODE3[0] x2.x3.x4[3].floating 2.28e-21
C763 sample_delay_offset a_4734_5318# 0.0126f
C764 CAP_CTRL_CODE0[1] x2.x4.x3[1].floating 0.227f
C765 CAP_CTRL_CODE3[2] x2.x3.x5[7].floating 0.00568f
C766 a_11283_5456# CAP_CTRL_CODE0[0] 0.00654f
C767 x2.x4.x6.SW CAP_CTRL_CODE0[1] 5.52e-21
C768 x2.x1.IN CAP_CTRL_CODE1[3] 0.00868f
C769 x2.x2.x9.output_stack a_16821_2232# 0.0702f
C770 a_4574_5180# CAP_CTRL_CODE2[2] 2.86e-20
C771 x2.x2.x9.output_stack x2.x2.x5[7].floating 1.19f
C772 x2.x2.x6.SW x2.x2.IN 0.0928f
C773 x2.x4.x7.floating a_4662_6008# 8.52e-19
C774 x3.A a_2790_6116# 2.16e-20
C775 a_11308_7535# a_11396_7397# 0.0704f
C776 a_3813_6132# x2.x4.x5[7].floating 2.06e-20
C777 a_3041_6494# a_3222_6482# 4.11e-20
C778 a_11443_5594# x2.x4.x2.floating 6.88e-19
C779 a_10137_3759# a_10065_3759# 0.00227f
C780 x2.x3.x10.Y a_10024_2094# 4.2e-19
C781 a_4047_3022# CAP_CTRL_CODE3[1] 3.52e-20
C782 CAP_CTRL_CODE0[0] x2.x4.x7.floating 2.03e-20
C783 x2.x3.x9.output_stack sample_clk 1.49e-20
C784 a_10137_3207# a_10756_3022# 0.00348f
C785 x3.A a_2932_6494# 2.67e-19
C786 x2.x3.x9.output_stack x2.x2.x5[7].floating 1.33e-19
C787 a_2619_6316# a_2837_6438# 3.73e-19
C788 a_16774_4173# x2.x2.IN 1.34e-19
C789 x1.x4.Y a_2058_6116# 3.34e-21
C790 sample_delay_offset x2.x2.x7.floating 0.264f
C791 x2.x4.x9.output_stack x2.x4.x4[3].floating 0.636f
C792 a_3813_6132# a_4574_6008# 2.47e-19
C793 a_10065_4035# x2.x2.x2.floating 2.21e-19
C794 vdd x2.x3.IN 0.612f
C795 a_4599_7259# x2.x4.x5[7].floating 2.76e-19
C796 sample_delay_offset a_16774_3345# 0.00155f
C797 a_16821_1680# x2.x2.IN 0.00832f
C798 a_4574_5180# x2.x4.x7.floating 0.00218f
C799 a_11396_7397# x2.x1.x9.output_stack 1.5e-19
C800 vdd x2.x2.IN 0.707f
C801 a_4047_2819# x2.x3.x5[7].floating 0.0132f
C802 x3.A CAP_CTRL_CODE2[2] 0.00188f
C803 sample_delay_offset CAP_CTRL_CODE0[2] 0.0696f
C804 set x1.x3.Y 0.0536f
C805 a_11396_7397# sample_delay_offset 1.9e-19
C806 a_10472_6193# CAP_CTRL_CODE1[2] 0.00525f
C807 CAP_CTRL_CODE0[2] a_4662_6146# 1.06e-19
C808 a_11443_5870# x2.x1.x4[3].floating 8.29e-19
C809 a_11443_5870# a_11283_5732# 0.0388f
C810 a_16846_3759# x2.x2.x7.floating 0.00409f
C811 a_11443_5870# x2.x1.x6.floating 0.00278f
C812 a_16733_2094# a_16821_1956# 0.0704f
C813 a_10024_2094# a_10024_1818# 0.0316f
C814 CAP_CTRL_CODE1[1] a_17181_6193# 3.4e-20
C815 a_16774_3621# a_16846_3483# 0.00227f
C816 x2.x2.x5[7].floating a_16733_1818# 0.00154f
C817 x7.A x2.x3.x5[7].floating 0.0208f
C818 sample_delay_offset a_2325_6090# 8.22e-21
C819 a_10137_3483# a_9977_3345# 0.0388f
C820 sample_delay_offset x2.x3.x6.SW 0.19f
C821 x2.x3.IN a_10137_3483# 0.0136f
C822 vdd a_3056_2150# 0.293f
C823 vdd a_2569_6116# 0.0112f
C824 sample_delay_offset a_16774_3207# 0.00167f
C825 sample_delay_offset a_4574_5732# 0.00384f
C826 sample_delay_offset CAP_CTRL_CODE3[0] 0.00152f
C827 x1.x3.Y a_4574_6008# 2.23e-20
C828 vdd x2.x2.x4[3].floating 0.0565f
C829 x3.A x2.x4.x7.floating 0.0275f
C830 sample_delay_offset a_16821_1956# 6.38e-19
C831 vdd CAP_CTRL_CODE1[0] 0.00346f
C832 x2.x1.x5[7].floating x2.x1.x2.floating 0.441f
C833 a_9977_3345# x2.x2.x2.floating 6.24e-19
C834 vdd a_3106_6090# 0.567f
C835 x7.A a_2678_2626# 2.12e-20
C836 x2.x3.x9.output_stack x2.x3.x4[3].floating 0.636f
C837 x2.x3.IN x2.x2.x2.floating 0.0257f
C838 x3.A a_3056_2936# 0.00499f
C839 a_10137_4035# CAP_CTRL_CODE2[2] 6.93e-20
C840 x2.x4.x6.SW x2.x4.x6.floating 0.128f
C841 x2.x1.IN a_11371_6008# 0.0013f
C842 x2.x1.x9.output_stack a_11371_6146# 0.00227f
C843 x2.x4.x5[7].floating CAP_CTRL_CODE0[0] 0.00131f
C844 CAP_CTRL_CODE3[1] x2.x3.x10.Y 6.71e-19
C845 a_4599_7535# x2.x4.x6.floating 0.00578f
C846 sample_delay_offset a_11371_6146# 0.00167f
C847 a_9977_3897# a_10065_4035# 0.00227f
C848 a_16846_4035# a_16686_3897# 0.0388f
C849 a_4574_6008# a_4662_6008# 0.00227f
C850 CAP_CTRL_CODE2[1] CAP_CTRL_CODE2[2] 4.67f
C851 vdd x2.x3.x3[1].floating 0.0301f
C852 a_10137_3207# a_10065_3207# 0.00227f
C853 a_4734_5594# a_4574_5456# 0.0388f
C854 a_11371_5732# a_11443_5594# 0.00227f
C855 x2.x4.x9.output_stack x2.x1.x9.output_stack 2.93e-20
C856 x2.x4.x10.Y a_10472_6534# 0.00127f
C857 x2.x4.x2.floating CAP_CTRL_CODE1[0] 1.61e-20
C858 a_16774_3345# x2.x2.x7.floating 8.52e-19
C859 x2.x4.x4[3].floating CAP_CTRL_CODE1[1] 6.93e-20
C860 a_10137_3207# x2.x3.x10.Y 1.69e-19
C861 clk x1.x3.Y 4.05e-19
C862 x2.x4.x10.Y x2.x4.x7.floating 0.00345f
C863 a_10137_3759# x2.x3.x7.floating 0.00409f
C864 a_11443_5318# x2.x1.x9.output_stack 8.05e-20
C865 sample_delay_offset x2.x4.x9.output_stack 0.263f
C866 reset x1.x2.D 0.00215f
C867 sample_delay_offset a_10065_3759# 0.00111f
C868 vdd CAP_CTRL_CODE0[1] 0.0182f
C869 x2.x4.x9.output_stack a_4662_6146# 0.00227f
C870 sample_delay_offset a_11443_5318# 0.0126f
C871 x2.x1.IN CAP_CTRL_CODE2[2] 5.86e-20
C872 x2.x1.x6.SW CAP_CTRL_CODE1[2] 3.93e-21
C873 x2.x3.x4[3].floating x2.x3.x7.floating 1.18f
C874 vdd a_3340_6116# 0.0055f
C875 a_16686_3345# x2.x2.x6.SW 2.44e-19
C876 CAP_CTRL_CODE3[1] CAP_CTRL_CODE2[0] 3.47e-20
C877 a_1870_6122# a_3813_6132# 9.65e-21
C878 x2.x4.x4[3].floating x2.x4.x3[1].floating 1.19f
C879 x2.x3.x6.floating x2.x2.x5[7].floating 0.0231f
C880 x2.x2.x10.Y a_10756_2819# 0.00127f
C881 x2.x1.IN a_11283_5456# 0.0136f
C882 x2.x2.x9.output_stack a_16733_2094# 0.032f
C883 a_11283_5180# CAP_CTRL_CODE2[2] 2.86e-20
C884 a_16774_3207# x2.x2.x7.floating 8.52e-19
C885 a_4687_7397# a_4599_7259# 0.0704f
C886 x3.A x2.x4.x5[7].floating 0.00127f
C887 a_11308_7535# a_11308_7259# 0.0316f
C888 CAP_CTRL_CODE3[2] x2.x3.x3[1].floating 0.00838f
C889 x2.x4.x9.output_stack a_4734_5318# 8.05e-20
C890 x2.x3.x10.Y a_10112_1956# 2.35e-19
C891 x2.x1.IN a_10472_6534# 0.15f
C892 CAP_CTRL_CODE0[1] x2.x4.x2.floating 0.0027f
C893 a_10137_3207# CAP_CTRL_CODE2[0] 0.00186f
C894 a_4734_5870# x2.x4.x6.floating 0.00278f
C895 x2.x3.IN a_9977_3897# 0.0135f
C896 sample_delay_offset x2.x2.x9.output_stack 0.264f
C897 a_11283_5456# a_11283_5180# 0.0316f
C898 a_1704_6122# a_2235_6116# 5.76e-19
C899 a_2932_6494# a_2837_6438# 0.00276f
C900 a_2619_6316# a_3222_6482# 0.0552f
C901 a_2151_6116# a_2235_6116# 0.00972f
C902 a_3106_6090# a_3041_6494# 4.2e-20
C903 x2.x3.x5[7].floating a_2678_2006# 8.78e-19
C904 a_4574_5732# CAP_CTRL_CODE0[2] 1.33e-19
C905 a_10065_3345# x2.x3.x7.floating 8.52e-19
C906 x3.A a_4574_6008# 0.0311f
C907 x2.x1.x10.Y x2.x1.x6.SW 0.788f
C908 CAP_CTRL_CODE2[2] x2.x2.x10.Y 0.00201f
C909 a_4734_5870# x1.x4.Y 1.29e-20
C910 a_4687_7121# x2.x4.x5[7].floating 0.00169f
C911 sample_delay_offset x2.x3.x9.output_stack 0.261f
C912 a_11308_7535# x2.x1.x6.floating 0.00578f
C913 x2.x2.x6.SW a_16821_2232# 0.00707f
C914 a_1704_6122# a_2619_6316# 0.124f
C915 a_2151_6116# a_2619_6316# 0.0633f
C916 a_1870_6122# x1.x3.Y 0.346f
C917 x2.x2.x6.SW x2.x2.x5[7].floating 0.00138f
C918 x1.x2.D a_2151_6116# 0.0392f
C919 a_1704_6122# x1.x2.D 0.647f
C920 a_2678_2626# a_2678_2006# 0.0231f
C921 x2.x4.x10.Y x2.x4.x5[7].floating 1.01f
C922 a_11308_7259# sample_delay_offset 6.38e-19
C923 x2.x1.x9.output_stack CAP_CTRL_CODE1[1] 0.0731f
C924 a_4574_5180# CAP_CTRL_CODE3[1] 1.48e-20
C925 a_10756_3022# CAP_CTRL_CODE2[0] 0.00699f
C926 a_11308_6983# x2.x1.x9.output_stack 0.0702f
C927 sample_delay_offset CAP_CTRL_CODE1[1] 0.0596f
C928 x3.A a_4662_5456# 5.79e-19
C929 x2.x3.x2.floating x2.x3.x5[7].floating 0.441f
C930 x2.x1.x9.output_stack x2.x1.x4[3].floating 0.636f
C931 sample_delay_offset a_11308_6983# 0.00273f
C932 a_10112_1956# a_10024_1818# 0.0704f
C933 x2.x3.IN CAP_CTRL_CODE1[2] 4.34e-20
C934 x3.Y x2.x3.x5[7].floating 0.00713f
C935 a_16733_2094# a_16733_1818# 0.0316f
C936 x2.x2.x5[7].floating a_16821_1680# 2.14e-19
C937 vdd sample_clk 0.708f
C938 x2.x1.x9.output_stack x2.x1.x6.floating 0.229f
C939 sample_delay_offset a_10065_4173# 5.66e-19
C940 vdd a_16821_2232# 0.104f
C941 x2.x4.x10.Y a_4574_6008# 1.69e-19
C942 vdd x2.x4.x6.floating 5.79f
C943 vdd x2.x2.x5[7].floating 44f
C944 sample_delay_offset x2.x1.x4[3].floating 0.00732f
C945 sample_delay_offset a_11283_5732# 0.00384f
C946 a_4047_3022# CAP_CTRL_CODE2[0] 6.85e-22
C947 x7.Y CAP_CTRL_CODE3[0] 8.54e-21
C948 x2.x4.x9.output_stack CAP_CTRL_CODE0[2] 0.334f
C949 sample_delay_offset x2.x1.x6.floating 0.0706f
C950 a_16846_3483# x2.x2.IN 0.03f
C951 sample_delay_offset a_16733_1818# 1.9e-19
C952 x2.x1.x7.floating a_11283_6008# 0.00409f
C953 a_2678_2626# x2.x3.x2.floating 8.88e-20
C954 a_2678_2626# x3.Y 0.00609f
C955 a_4734_5870# x2.x4.x4[3].floating 8.29e-19
C956 sample_delay_offset x2.x3.x7.floating 0.261f
C957 vdd x1.x4.Y 1.47f
C958 sample_delay_offset x2.x4.x3[1].floating 6.03e-20
C959 x3.A CAP_CTRL_CODE3[1] 0.00183f
C960 vdd a_17181_6193# 0.237f
C961 x2.x2.x6.floating x2.x2.IN 0.0299f
C962 x2.x1.IN x2.x4.x5[7].floating 0.0218f
C963 x2.x2.x9.output_stack x2.x2.x7.floating 0.185f
C964 CAP_CTRL_CODE1[3] x2.x1.x6.SW 0.00466f
C965 a_11443_5870# x2.x4.x2.floating 6.24e-19
C966 sample_delay_offset x2.x4.x6.SW 0.19f
C967 a_11371_5456# x2.x1.x7.floating 8.52e-19
C968 a_4599_7535# sample_delay_offset 3.28e-19
C969 CAP_CTRL_CODE0[0] a_11283_6008# 0.00181f
C970 CAP_CTRL_CODE1[2] CAP_CTRL_CODE1[0] 3.87e-19
C971 x2.x1.x10.Y x2.x2.IN 1.13e-19
C972 a_16846_3483# x2.x2.x4[3].floating 1.17e-19
C973 x3.A a_4687_7397# 0.00847f
C974 sample_delay_offset a_16774_3759# 0.00111f
C975 a_4734_5594# x2.x4.x7.floating 0.00959f
C976 sample_delay_offset a_4662_5318# 9.69e-19
C977 x2.x2.x2.floating x2.x2.x5[7].floating 0.441f
C978 vdd a_17181_6534# 0.217f
C979 vdd x2.x3.x4[3].floating 0.0565f
C980 vdd x2.x4.x4[3].floating 0.0565f
C981 x2.x2.x9.output_stack x2.x3.x6.SW 3.62e-19
C982 CAP_CTRL_CODE2[2] a_10472_6193# 3.71e-21
C983 a_1870_6122# a_2259_6494# 0.0019f
C984 x2.x4.x6.SW a_4734_5318# 7.9e-20
C985 a_2325_6090# a_2058_6116# 6.99e-20
C986 x1.x3.Y a_3813_6132# 4.86e-19
C987 x2.x2.x9.output_stack a_16774_3207# 0.00227f
C988 x3.A a_1870_6122# 4.92e-20
C989 a_10065_3207# CAP_CTRL_CODE2[0] 8.23e-20
C990 x2.x1.x10.Y CAP_CTRL_CODE1[0] 0.0124f
C991 CAP_CTRL_CODE2[0] x2.x3.x10.Y 2.78e-20
C992 a_11396_7397# a_11308_7259# 0.0704f
C993 a_2678_2006# a_3056_2150# 0.0895f
C994 CAP_CTRL_CODE1[0] x2.x1.x3[1].floating 0.0394f
C995 a_4687_7397# a_4687_7121# 0.0316f
C996 vdd a_3553_3025# 5.6e-19
C997 sample_delay_offset x2.x3.x6.floating 0.0706f
C998 a_11371_5594# x2.x4.x2.floating 2.21e-19
C999 CAP_CTRL_CODE3[1] CAP_CTRL_CODE2[1] 3.2e-20
C1000 a_10137_3759# a_10137_3483# 0.0316f
C1001 x2.x3.x10.Y a_10024_1818# 1.49e-19
C1002 x2.x3.x9.output_stack x2.x3.x6.SW 0.164f
C1003 a_16846_3759# a_16774_3759# 0.00227f
C1004 CAP_CTRL_CODE0[1] CAP_CTRL_CODE1[2] 3.42e-20
C1005 CAP_CTRL_CODE0[2] CAP_CTRL_CODE1[1] 6.3e-20
C1006 x2.x3.x9.output_stack CAP_CTRL_CODE3[0] 0.0285f
C1007 a_10472_6534# a_10472_6193# 0.0121f
C1008 CAP_CTRL_CODE2[2] x2.x2.x3[1].floating 0.00624f
C1009 a_4734_5318# a_4662_5318# 0.00227f
C1010 a_4687_7397# x2.x4.x10.Y 1.49e-19
C1011 x3.A a_4047_3022# 0.00142f
C1012 x1.x2.D a_2569_6116# 0.00306f
C1013 a_16686_3897# x2.x2.IN 0.0166f
C1014 a_1704_6122# a_2790_6116# 0.00566f
C1015 a_2932_6494# a_3222_6482# 0.0282f
C1016 a_2619_6316# a_2569_6116# 1.21e-20
C1017 x2.x3.x5[7].floating a_10112_2232# 2.76e-19
C1018 sample_delay_offset a_4734_5870# 0.0155f
C1019 a_10137_3759# x2.x2.x2.floating 0.00177f
C1020 a_10137_3483# x2.x3.x4[3].floating 1.17e-19
C1021 a_4599_6983# x2.x4.x5[7].floating 2.76e-19
C1022 a_11396_7397# x2.x1.x6.floating 0.0191f
C1023 x2.x3.x9.output_stack x7.Y 4.33e-19
C1024 CAP_CTRL_CODE0[3] x2.x4.x6.floating 0.00405f
C1025 CAP_CTRL_CODE3[2] x2.x3.x4[3].floating 0.536f
C1026 a_2619_6316# a_3106_6090# 0.27f
C1027 a_11396_7121# x2.x1.x9.output_stack 0.032f
C1028 x1.x2.D a_3106_6090# 0.208f
C1029 a_1704_6122# a_2932_6494# 0.0322f
C1030 vdd a_11308_7535# 0.179f
C1031 CAP_CTRL_CODE0[2] x2.x4.x3[1].floating 0.00115f
C1032 x7.A sample_clk 4.05e-20
C1033 x3.Y a_3056_2150# 0.432f
C1034 a_11396_7121# sample_delay_offset 3.64e-19
C1035 sample_delay_offset x2.x2.x6.SW 0.19f
C1036 a_16774_3759# x2.x2.x7.floating 8.52e-19
C1037 a_16686_3897# x2.x2.x4[3].floating 7.47e-19
C1038 x2.x4.x6.SW CAP_CTRL_CODE0[2] 9.76e-21
C1039 x2.x3.x7.floating x2.x3.x6.SW 9.72e-19
C1040 a_10112_1956# a_10112_1680# 0.0316f
C1041 a_16821_1956# a_16733_1818# 0.0704f
C1042 a_9977_3345# a_10065_3483# 0.00227f
C1043 a_16846_3483# a_16686_3345# 0.0388f
C1044 a_10756_3022# CAP_CTRL_CODE2[1] 4.37e-20
C1045 sample_delay_offset a_16774_4173# 5.68e-19
C1046 x2.x3.IN a_10065_3483# 7.93e-19
C1047 vdd a_16733_2094# 0.0737f
C1048 sample_delay_offset a_4662_5732# 0.00123f
C1049 vdd x2.x1.x9.output_stack 0.596f
C1050 sample_delay_offset a_16821_1680# 3.28e-19
C1051 x2.x3.x2.floating x2.x3.x3[1].floating 1.17f
C1052 a_4662_5318# CAP_CTRL_CODE0[2] 8.73e-19
C1053 a_16686_3345# x2.x2.x6.floating 0.00278f
C1054 x2.x4.x9.output_stack CAP_CTRL_CODE1[1] 4.64e-20
C1055 vdd sample_delay_offset 0.928f
C1056 a_4047_3022# CAP_CTRL_CODE2[1] 9.41e-22
C1057 a_16846_3759# x2.x2.x6.SW 4.74e-20
C1058 x2.x4.x6.SW a_4574_5732# 8.11e-20
C1059 a_10065_3345# x2.x2.x2.floating 1.6e-19
C1060 x1.x2.D a_3340_6116# 0.00273f
C1061 a_3106_6090# a_3018_6116# 7.71e-20
C1062 a_11283_5456# x2.x1.x6.SW 4.74e-20
C1063 vdd a_4662_6146# 1.29e-19
C1064 a_2619_6316# a_3340_6116# 7.61e-19
C1065 x3.A a_3813_6132# 0.0827f
C1066 set reset 0.0236f
C1067 a_16686_3897# a_16774_4035# 0.00227f
C1068 a_9977_3897# a_10137_3759# 0.0388f
C1069 x2.x4.x6.floating CAP_CTRL_CODE1[2] 3.95e-22
C1070 x2.x1.x6.SW a_10472_6534# 0.00208f
C1071 x2.x4.x9.output_stack x2.x1.x6.floating 4.17e-19
C1072 x2.x3.x9.output_stack x2.x2.x9.output_stack 2.93e-20
C1073 a_11443_5594# a_11283_5456# 0.0388f
C1074 a_3056_2936# x2.x3.x5[7].floating 7.35e-19
C1075 a_11443_5318# x2.x1.x4[3].floating 7.47e-19
C1076 a_4574_5180# CAP_CTRL_CODE2[0] 2e-20
C1077 x2.x1.x9.output_stack x2.x4.x2.floating 2.95e-19
C1078 a_4574_5456# a_4662_5594# 0.00227f
C1079 vdd sample_clk_b 0.716f
C1080 a_11443_5318# x2.x1.x6.floating 0.00109f
C1081 x2.x4.x9.output_stack x2.x4.x3[1].floating 0.341f
C1082 x2.x3.IN a_10112_2232# 0.0175f
C1083 vdd a_16846_3759# 4.84e-19
C1084 sample_delay_offset x2.x4.x2.floating 0.0039f
C1085 x2.x1.IN a_11283_6008# 0.0217f
C1086 x2.x3.IN a_10756_2819# 0.15f
C1087 a_10065_3759# x2.x3.x7.floating 8.52e-19
C1088 a_9977_3897# x2.x3.x4[3].floating 7.47e-19
C1089 sample_delay_offset a_10137_3483# 0.00378f
C1090 x2.x2.x6.floating a_16821_2232# 0.00996f
C1091 x3.A a_4599_7259# 0.00866f
C1092 sample_delay_offset a_11371_5318# 9.69e-19
C1093 x2.x2.x5[7].floating x2.x2.x6.floating 1.18f
C1094 a_2678_2626# a_3056_2936# 0.0969f
C1095 x2.x2.x9.output_stack CAP_CTRL_CODE1[1] 2.48e-21
C1096 x2.x3.x6.SW x2.x3.x6.floating 0.13f
C1097 x2.x4.x6.SW x2.x4.x9.output_stack 0.164f
C1098 x2.x2.x7.floating x2.x2.x6.SW 9.72e-19
C1099 sample_delay_offset CAP_CTRL_CODE3[2] 0.00886f
C1100 a_2325_6090# a_2465_6482# 0.07f
C1101 x3.A x1.x3.Y 0.0052f
C1102 a_1870_6122# a_2837_6438# 0.00126f
C1103 a_4574_5180# CAP_CTRL_CODE0[0] 1.99e-19
C1104 x2.x2.IN x2.x1.x2.floating 0.0392f
C1105 sample_delay_offset x2.x2.x2.floating 0.00558f
C1106 x2.x1.IN a_11371_5456# 2.42e-19
C1107 x2.x3.x9.output_stack CAP_CTRL_CODE1[1] 2.48e-21
C1108 a_10137_4035# x2.x3.x10.Y 2.2e-20
C1109 x3.A CAP_CTRL_CODE2[0] 0.00182f
C1110 x2.x2.x9.output_stack a_16733_1818# 1.5e-19
C1111 x2.x3.IN CAP_CTRL_CODE2[2] 1.46e-19
C1112 a_2678_2006# sample_clk 0.00102f
C1113 x3.A a_4662_5870# 0.00113f
C1114 a_4599_7259# a_4687_7121# 0.0704f
C1115 a_11396_7397# a_11396_7121# 0.0316f
C1116 a_11371_5594# CAP_CTRL_CODE1[2] 2.32e-19
C1117 a_9977_3621# a_10065_3621# 0.00227f
C1118 a_4734_5870# a_4574_5732# 0.0388f
C1119 x2.x3.x10.Y a_10112_1680# 1.02e-19
C1120 x2.x2.x9.output_stack x2.x3.x7.floating 3.32e-19
C1121 x2.x3.IN a_10065_3897# 2.42e-19
C1122 vdd x2.x2.x7.floating 0.0321f
C1123 a_4599_7259# x2.x4.x10.Y 2.35e-19
C1124 set a_1704_6122# 0.00161f
C1125 a_11308_7259# a_11308_6983# 0.0316f
C1126 sample_delay_offset a_3041_6494# 4.25e-20
C1127 x2.x1.x3[1].floating a_17181_6193# 3.09e-19
C1128 x1.x2.D x2.x4.x6.floating 6.74e-20
C1129 a_2619_6316# x2.x4.x6.floating 1.55e-20
C1130 x2.x3.x5[7].floating a_10024_2094# 0.00169f
C1131 x2.x4.x4[3].floating CAP_CTRL_CODE1[2] 7.49e-20
C1132 x2.x3.x9.output_stack x2.x3.x7.floating 0.185f
C1133 a_4662_5732# CAP_CTRL_CODE0[2] 2.5e-19
C1134 x3.A a_4662_6008# 0.00163f
C1135 a_11308_7259# x2.x1.x6.floating 0.00996f
C1136 x3.A CAP_CTRL_CODE0[0] 0.00183f
C1137 CAP_CTRL_CODE1[1] x2.x1.x4[3].floating 0.0226f
C1138 CAP_CTRL_CODE1[0] x2.x1.x2.floating 0.163f
C1139 x2.x2.x6.SW a_16821_1956# 9.98e-20
C1140 a_2619_6316# x1.x4.Y 0.107f
C1141 a_3106_6090# a_2932_6494# 0.197f
C1142 x2.x1.x6.SW x2.x4.x5[7].floating 0.00313f
C1143 x1.x2.D x1.x4.Y 0.0552f
C1144 vdd CAP_CTRL_CODE0[2] 0.0374f
C1145 x2.x3.x2.floating sample_clk 9.72e-20
C1146 x3.Y sample_clk 0.00198f
C1147 vdd a_11396_7397# 0.138f
C1148 a_11308_6983# x2.x1.x6.floating 0.00996f
C1149 CAP_CTRL_CODE2[2] x2.x2.x4[3].floating 0.53f
C1150 CAP_CTRL_CODE0[3] sample_delay_offset 0.0294f
C1151 a_10137_4035# CAP_CTRL_CODE2[0] 0.0131f
C1152 a_11283_5732# x2.x1.x4[3].floating 1.17e-19
C1153 a_11371_5870# x2.x1.x7.floating 8.52e-19
C1154 a_4574_5732# a_4662_5732# 0.00227f
C1155 x2.x4.x3[1].floating CAP_CTRL_CODE1[1] 3.46e-20
C1156 x2.x1.x5[7].floating x2.x1.x7.floating 0.182f
C1157 x3.A a_4574_5180# 0.014f
C1158 vdd a_2325_6090# 0.323f
C1159 x2.x4.x9.output_stack a_4734_5870# 0.032f
C1160 vdd x2.x3.x6.SW 0.45f
C1161 x2.x1.x10.Y a_17181_6534# 0.00127f
C1162 a_10024_1818# a_10112_1680# 0.0704f
C1163 a_16821_1956# a_16821_1680# 0.0316f
C1164 vdd a_16774_3207# 1.29e-19
C1165 vdd a_4574_5732# 0.00849f
C1166 CAP_CTRL_CODE2[0] CAP_CTRL_CODE2[1] 4.26f
C1167 vdd CAP_CTRL_CODE3[0] 0.00327f
C1168 sample_delay_offset a_9977_3897# 0.0121f
C1169 vdd a_16821_1956# 0.0343f
C1170 sample_delay_offset a_11371_5732# 0.00123f
C1171 x2.x4.x10.Y CAP_CTRL_CODE0[0] 0.0125f
C1172 a_16774_3483# x2.x2.IN 7.93e-19
C1173 x2.x2.x9.output_stack x2.x3.x6.floating 4.17e-19
C1174 x2.x3.x3[1].floating CAP_CTRL_CODE2[2] 3.26e-20
C1175 vdd x7.Y 0.326f
C1176 x2.x4.x7.floating CAP_CTRL_CODE1[0] 1.61e-20
C1177 clk a_1704_6122# 0.246f
C1178 x2.x1.IN x2.x1.x7.floating 0.0242f
C1179 x2.x1.IN CAP_CTRL_CODE2[0] 4.21e-20
C1180 x2.x3.x10.Y x2.x2.x10.Y 1.79e-20
C1181 a_3056_2936# a_3056_2150# 0.00995f
C1182 x1.x4.Y a_3018_6116# 2.7e-19
C1183 vdd a_11371_6146# 1.29e-19
C1184 a_3106_6090# x2.x4.x7.floating 0.00116f
C1185 reset a_1870_6122# 2.47e-20
C1186 x2.x4.x10.Y a_4574_5180# 2.2e-20
C1187 x2.x3.x9.output_stack x2.x3.x6.floating 0.229f
C1188 a_16846_3207# x2.x2.x10.Y 1.69e-19
C1189 a_10137_3483# x2.x3.x6.SW 8.11e-20
C1190 a_10065_3621# CAP_CTRL_CODE2[0] 1.74e-19
C1191 a_11283_5180# CAP_CTRL_CODE2[0] 2e-20
C1192 CAP_CTRL_CODE3[1] x2.x3.x5[7].floating 0.00224f
C1193 a_11283_5180# x2.x1.x7.floating 0.00218f
C1194 x2.x1.x9.output_stack CAP_CTRL_CODE1[2] 0.333f
C1195 vdd x2.x4.x9.output_stack 0.595f
C1196 a_11308_7535# x2.x1.x10.Y 1.02e-19
C1197 CAP_CTRL_CODE3[0] CAP_CTRL_CODE3[2] 1.89e-20
C1198 x2.x3.IN a_10024_2094# 0.00921f
C1199 sample_delay_offset CAP_CTRL_CODE1[2] 0.0969f
C1200 x2.x1.IN CAP_CTRL_CODE0[0] 8.71e-19
C1201 a_4574_5180# CAP_CTRL_CODE2[1] 2.37e-20
C1202 a_4599_7535# x2.x4.x6.SW 5.11e-20
C1203 sample_delay_offset a_16846_3483# 0.00382f
C1204 x2.x4.x2.floating a_11371_6146# 2.02e-19
C1205 x2.x2.x9.output_stack x2.x2.x6.SW 0.164f
C1206 a_10472_6193# a_11283_6008# 0.00348f
C1207 x2.x2.x6.floating a_16733_2094# 0.0194f
C1208 x3.A a_4687_7121# 0.00921f
C1209 a_4574_5456# x2.x4.x4[3].floating 1.17e-19
C1210 sample_delay_offset a_11371_5180# 5.69e-19
C1211 a_3553_3025# x2.x3.x2.floating 4.02e-20
C1212 a_10756_3022# x2.x2.x3[1].floating 3.09e-19
C1213 a_4662_5594# x2.x4.x7.floating 8.52e-19
C1214 x3.Y a_3553_3025# 0.00962f
C1215 CAP_CTRL_CODE0[1] x2.x4.x7.floating 2.21e-20
C1216 CAP_CTRL_CODE2[0] x2.x2.x10.Y 0.0124f
C1217 x3.A x2.x4.x10.Y 0.0967f
C1218 sample_delay_offset x2.x2.x6.floating 0.0706f
C1219 x1.x3.Y a_2837_6438# 0.00408f
C1220 a_11283_5180# CAP_CTRL_CODE0[0] 0.00533f
C1221 a_11371_6008# a_11443_5870# 0.00227f
C1222 x2.x4.x9.output_stack x2.x4.x2.floating 0.193f
C1223 x2.x3.x7.floating x2.x3.x6.floating 0.202f
C1224 x2.x1.x10.Y x2.x1.x9.output_stack 1.01f
C1225 x2.x1.x9.output_stack x2.x1.x3[1].floating 0.341f
C1226 a_4599_7259# a_4599_6983# 0.0316f
C1227 a_11308_7259# a_11396_7121# 0.0704f
C1228 x2.x2.x5[7].floating a_10112_2232# 1.79e-19
C1229 vdd x2.x2.x9.output_stack 0.595f
C1230 a_11443_5318# x2.x4.x2.floating 6.88e-19
C1231 a_16846_3759# a_16846_3483# 0.0316f
C1232 sample_delay_offset x2.x1.x10.Y 0.0402f
C1233 a_1870_6122# a_2151_6116# 0.155f
C1234 a_10756_2819# x2.x2.x5[7].floating 0.0132f
C1235 vdd a_2058_6116# 0.109f
C1236 sample_delay_offset x2.x1.x3[1].floating 3.48e-20
C1237 a_1704_6122# a_1870_6122# 0.782f
C1238 x3.A CAP_CTRL_CODE2[1] 0.00184f
C1239 a_4687_7121# x2.x4.x10.Y 4.2e-19
C1240 a_11396_7121# a_11308_6983# 0.0704f
C1241 a_11443_5318# a_11371_5318# 0.00227f
C1242 x1.x4.Y a_2790_6116# 7.18e-19
C1243 a_2932_6494# x2.x4.x6.floating 4.63e-21
C1244 a_16774_3897# x2.x2.IN 2.42e-19
C1245 x2.x3.x5[7].floating a_10112_1956# 2.76e-19
C1246 vdd x2.x3.x9.output_stack 0.599f
C1247 a_10065_3759# x2.x2.x2.floating 2.21e-19
C1248 a_11396_7121# x2.x1.x6.floating 0.0194f
C1249 sample_delay_offset a_2619_6316# 0.00134f
C1250 x7.Y a_4047_2819# 0.00365f
C1251 sample_delay_offset x1.x2.D 0.00127f
C1252 a_2932_6494# x1.x4.Y 0.00621f
C1253 vdd a_11308_7259# 0.0923f
C1254 a_9977_3897# x2.x3.x6.SW 7.9e-20
C1255 x7.A CAP_CTRL_CODE3[0] 4.4e-19
C1256 x2.x4.x6.SW a_4734_5870# 2.44e-19
C1257 CAP_CTRL_CODE2[2] x2.x2.x5[7].floating 0.0056f
C1258 a_3106_6090# a_4574_6008# 3e-19
C1259 a_2678_2006# sample_clk_b 0.109f
C1260 x2.x1.x2.floating a_17181_6193# 0.0104f
C1261 vdd CAP_CTRL_CODE1[1] 0.0183f
C1262 vdd a_11308_6983# 0.11f
C1263 sample_delay_offset x2.x3.x2.floating 0.00186f
C1264 a_16846_3483# x2.x2.x7.floating 0.00409f
C1265 a_4047_3022# a_2678_2626# 8.79e-20
C1266 x7.Y x7.A 0.0744f
C1267 x2.x4.x5[7].floating CAP_CTRL_CODE0[1] 0.00228f
C1268 a_10137_4035# CAP_CTRL_CODE2[1] 9.56e-20
C1269 x2.x1.x6.SW a_11283_6008# 0.00179f
C1270 a_16733_1818# a_16821_1680# 0.0704f
C1271 vdd x2.x1.x4[3].floating 0.0565f
C1272 a_16686_3345# a_16774_3483# 0.00227f
C1273 a_9977_3345# a_10137_3207# 0.0388f
C1274 sample_delay_offset a_16686_3897# 0.0124f
C1275 x2.x2.x9.output_stack x2.x2.x2.floating 0.193f
C1276 vdd a_16733_1818# 0.129f
C1277 vdd x2.x1.x6.floating 5.87f
C1278 x2.x3.IN a_10137_3207# 0.0217f
C1279 x2.x2.x7.floating x2.x2.x6.floating 0.202f
C1280 sample_delay_offset a_4574_5456# 0.00299f
C1281 CAP_CTRL_CODE0[2] CAP_CTRL_CODE1[2] 6.83e-20
C1282 x2.x3.x9.output_stack CAP_CTRL_CODE3[2] 0.334f
C1283 x2.x4.x6.floating x2.x4.x7.floating 0.202f
C1284 sample_delay_offset CAP_CTRL_CODE1[3] 0.0294f
C1285 vdd x2.x3.x7.floating 0.0315f
C1286 x2.x1.IN x2.x4.x10.Y 1.23e-19
C1287 vdd x2.x4.x3[1].floating 0.0301f
C1288 x2.x4.x2.floating CAP_CTRL_CODE1[1] 1.73e-20
C1289 a_3056_2936# sample_clk 0.00366f
C1290 x2.x3.x9.output_stack x2.x2.x2.floating 2.95e-19
C1291 x3.Y sample_clk_b 8.9e-19
C1292 x2.x1.IN a_11371_5870# 7.93e-19
C1293 x1.x4.Y x2.x4.x7.floating 3.62e-19
C1294 reset x1.x3.Y 0.0461f
C1295 x2.x1.IN x2.x1.x5[7].floating 0.00127f
C1296 x3.A a_2837_6438# 6.08e-20
C1297 vdd x2.x4.x6.SW 0.427f
C1298 a_11283_5732# x2.x4.x2.floating 0.00177f
C1299 a_10472_6193# x2.x1.x7.floating 7.29e-19
C1300 a_3340_6116# a_4574_6008# 3.49e-20
C1301 a_10065_3897# a_10137_3759# 0.00227f
C1302 vdd a_4599_7535# 0.149f
C1303 a_16686_3897# a_16846_3759# 0.0388f
C1304 x2.x1.IN CAP_CTRL_CODE2[1] 4.93e-20
C1305 a_11283_5456# a_11371_5594# 0.00227f
C1306 a_4574_5456# a_4734_5318# 0.0388f
C1307 x2.x3.x4[3].floating CAP_CTRL_CODE2[2] 6.52e-20
C1308 x2.x3.IN a_10756_3022# 0.157f
C1309 a_1704_6122# a_3813_6132# 1.03e-19
C1310 x2.x3.IN a_10112_1956# 0.00866f
C1311 a_11396_7397# x2.x1.x10.Y 1.49e-19
C1312 x2.x4.x3[1].floating x2.x4.x2.floating 1.17f
C1313 a_10137_3483# x2.x3.x7.floating 0.00409f
C1314 x2.x3.x10.Y x2.x3.x5[7].floating 1.01f
C1315 sample_delay_offset a_10065_3483# 0.00138f
C1316 CAP_CTRL_CODE2[0] x2.x2.x3[1].floating 0.0326f
C1317 a_11283_5180# CAP_CTRL_CODE2[1] 2.37e-20
C1318 x2.x2.x6.floating a_16821_1956# 0.00996f
C1319 CAP_CTRL_CODE3[2] x2.x3.x7.floating 0.0056f
C1320 CAP_CTRL_CODE1[2] a_11371_6146# 8.1e-20
C1321 x3.A a_4599_6983# 0.0175f
C1322 x2.x3.x9.output_stack a_4047_2819# 0.00887f
C1323 CAP_CTRL_CODE3[1] x2.x3.x3[1].floating 0.23f
C1324 CAP_CTRL_CODE0[0] a_10472_6193# 0.00169f
C1325 x2.x3.x7.floating x2.x2.x2.floating 0.0475f
C1326 x1.x3.Y a_3222_6482# 0.00974f
C1327 a_2325_6090# a_2235_6116# 6.69e-20
C1328 a_1870_6122# a_2569_6116# 2.46e-19
C1329 x2.x4.x7.floating x2.x4.x4[3].floating 1.18f
C1330 x2.x1.IN a_11283_5180# 0.0127f
C1331 x2.x4.x9.output_stack CAP_CTRL_CODE1[2] 0.00469f
C1332 vdd x2.x3.x6.floating 5.87f
C1333 a_16686_3897# x2.x2.x7.floating 0.00925f
C1334 x3.A a_4734_5594# 0.0138f
C1335 CAP_CTRL_CODE2[1] x2.x2.x10.Y 6.64e-19
C1336 x2.x4.x6.floating x2.x4.x5[7].floating 1.18f
C1337 x2.x3.x9.output_stack x7.A 0.127f
C1338 a_4687_7121# a_4599_6983# 0.0704f
C1339 a_9977_3897# x2.x3.x9.output_stack 8.05e-20
C1340 a_16686_3621# a_16774_3621# 0.00227f
C1341 a_10756_3022# CAP_CTRL_CODE1[0] 3.76e-21
C1342 a_1870_6122# a_3106_6090# 0.0264f
C1343 x1.x3.Y a_2151_6116# 0.152f
C1344 a_2325_6090# a_2619_6316# 0.199f
C1345 a_9977_3621# a_9977_3345# 0.0316f
C1346 x1.x2.D a_2325_6090# 0.0326f
C1347 a_1704_6122# x1.x3.Y 0.0445f
C1348 vdd a_2465_6482# 0.00118f
C1349 sample_delay_offset a_11371_6008# 0.00155f
C1350 x2.x3.IN a_9977_3621# 0.0135f
C1351 set x1.x4.Y 2.95e-19
C1352 CAP_CTRL_CODE2[0] x2.x3.x5[7].floating 1.4e-20
C1353 a_4574_5180# a_4662_5180# 0.0022f
C1354 a_4599_6983# x2.x4.x10.Y 0.039f
C1355 sample_delay_offset a_2790_6116# 1.82e-20
C1356 sample_delay_offset a_10112_2232# 0.00273f
C1357 vdd a_4734_5870# 0.00378f
C1358 sample_delay_offset a_10756_2819# 0.00117f
C1359 x2.x3.x5[7].floating a_10024_1818# 0.00154f
C1360 a_4574_5456# CAP_CTRL_CODE0[2] 2.81e-19
C1361 a_4047_3022# CAP_CTRL_CODE1[0] 5.53e-22
C1362 x2.x1.x9.output_stack x2.x1.x2.floating 0.193f
C1363 x2.x1.x6.SW x2.x1.x7.floating 9.72e-19
C1364 x2.x2.x6.SW a_16821_1680# 5.11e-20
C1365 sample_delay_offset a_2932_6494# 2.62e-19
C1366 CAP_CTRL_CODE3[0] x2.x3.x2.floating 0.17f
C1367 x2.x4.x9.output_stack x2.x1.x10.Y 1.93e-19
C1368 vdd a_11396_7121# 0.0797f
C1369 sample_delay_offset x2.x1.x2.floating 0.00286f
C1370 x1.x4.Y a_4574_6008# 5e-20
C1371 vdd x2.x2.x6.SW 0.43f
C1372 a_10065_4035# CAP_CTRL_CODE2[0] 5.2e-19
C1373 a_11443_5594# x2.x1.x7.floating 0.00959f
C1374 x2.x3.IN a_10065_3207# 0.00196f
C1375 a_4574_5732# a_4574_5456# 0.0316f
C1376 a_11283_5732# a_11371_5732# 0.00227f
C1377 sample_delay_offset CAP_CTRL_CODE2[2] 6.09f
C1378 x7.Y x2.x3.x2.floating 6.51e-19
C1379 x3.A a_4662_5180# 4.57e-19
C1380 a_4047_3022# x2.x3.x3[1].floating 3.09e-19
C1381 x7.Y x3.Y 0.0851f
C1382 a_9977_3897# x2.x3.x7.floating 0.00925f
C1383 CAP_CTRL_CODE0[3] x2.x4.x6.SW 0.00466f
C1384 x2.x3.IN x2.x3.x10.Y 0.0967f
C1385 x2.x2.x9.output_stack x2.x2.x6.floating 0.229f
C1386 x2.x4.x9.output_stack a_2619_6316# 2.26e-20
C1387 x2.x4.x9.output_stack x1.x2.D 1.79e-20
C1388 sample_delay_offset a_10065_3897# 0.00102f
C1389 vdd a_16821_1680# 0.112f
C1390 sample_delay_offset a_11283_5456# 0.00299f
C1391 x2.x4.x5[7].floating x2.x4.x4[3].floating 1.55f
C1392 x2.x1.x9.output_stack a_10472_6534# 1.18e-20
C1393 a_16846_3207# x2.x2.IN 0.038f
C1394 sample_delay_offset a_10472_6534# 0.00117f
C1395 CAP_CTRL_CODE1[2] CAP_CTRL_CODE1[1] 5.09f
C1396 sample_delay_offset x2.x4.x7.floating 0.259f
C1397 x2.x4.x7.floating a_4662_6146# 8.52e-19
C1398 x2.x4.x4[3].floating a_4574_6008# 1.17e-19
C1399 x3.A a_3222_6482# 6.54e-19
C1400 a_2465_6482# a_3041_6494# 2.46e-21
C1401 a_2058_6116# a_2235_6116# 8.94e-19
C1402 CAP_CTRL_CODE1[2] x2.x1.x4[3].floating 0.527f
C1403 a_11283_5732# CAP_CTRL_CODE1[2] 9.19e-20
C1404 x2.x1.x6.floating CAP_CTRL_CODE1[2] 3.95e-22
C1405 CAP_CTRL_CODE1[3] x2.x4.x9.output_stack 4.13e-19
C1406 x2.x3.IN CAP_CTRL_CODE2[0] 0.018f
C1407 vdd x2.x4.x2.floating 0.0334f
C1408 a_2151_6116# a_2259_6494# 0.00812f
C1409 x3.A a_2151_6116# 1.73e-20
C1410 a_2619_6316# a_2058_6116# 2.06e-20
C1411 a_3106_6090# a_3813_6132# 0.0968f
C1412 x1.x2.D a_2058_6116# 0.164f
C1413 x2.x3.IN a_10024_1818# 0.00847f
C1414 x2.x4.x3[1].floating CAP_CTRL_CODE1[2] 3.74e-20
C1415 a_11308_7259# x2.x1.x10.Y 2.35e-19
C1416 a_16846_3207# x2.x2.x4[3].floating 1.17e-19
C1417 x3.A a_1704_6122# 2.34e-19
C1418 x3.A x2.x3.x5[7].floating 2.66e-19
C1419 sample_delay_offset a_16774_3483# 0.00138f
C1420 a_4687_7397# x2.x4.x6.floating 0.0191f
C1421 a_11308_7535# x2.x4.x5[7].floating 4.6e-19
C1422 vdd CAP_CTRL_CODE3[2] 0.0374f
C1423 x2.x2.x6.floating a_16733_1818# 0.0191f
C1424 CAP_CTRL_CODE1[1] x2.x1.x3[1].floating 0.224f
C1425 x2.x1.x10.Y CAP_CTRL_CODE1[1] 6.64e-19
C1426 a_4734_5318# x2.x4.x7.floating 0.00925f
C1427 a_11308_6983# x2.x1.x10.Y 0.039f
C1428 a_16846_4035# x2.x2.x10.Y 2.2e-20
C1429 x2.x4.x6.SW CAP_CTRL_CODE1[2] 3.93e-21
C1430 a_9977_3897# x2.x3.x6.floating 0.00109f
C1431 x2.x1.IN a_10472_6193# 0.158f
C1432 CAP_CTRL_CODE2[1] x2.x2.x3[1].floating 0.226f
C1433 CAP_CTRL_CODE2[2] x2.x2.x7.floating 0.0056f
C1434 x2.x3.x3[1].floating x2.x3.x10.Y 0.00302f
C1435 x2.x1.x10.Y x2.x1.x4[3].floating 0.00668f
C1436 vdd x2.x2.x2.floating 0.0334f
C1437 x3.A a_2678_2626# 0.00228f
C1438 x2.x1.x4[3].floating x2.x1.x3[1].floating 1.19f
C1439 a_16686_3897# x2.x2.x9.output_stack 8.05e-20
C1440 a_11283_5732# x2.x1.x10.Y 6.65e-20
C1441 x1.x3.Y a_2569_6116# 9.85e-19
C1442 a_2325_6090# a_2790_6116# 9.46e-19
C1443 x2.x3.x6.SW a_10112_2232# 0.00707f
C1444 x2.x1.x10.Y x2.x1.x6.floating 0.0881f
C1445 x2.x3.x6.SW a_10756_2819# 0.00208f
C1446 x2.x3.x9.output_stack x2.x3.x2.floating 0.193f
C1447 x2.x3.x9.output_stack x3.Y 8.42e-19
C1448 CAP_CTRL_CODE2[0] x2.x2.x4[3].floating 2.28e-21
C1449 a_11371_5318# x2.x4.x2.floating 2.21e-19
C1450 CAP_CTRL_CODE3[1] x2.x3.x4[3].floating 0.00929f
C1451 CAP_CTRL_CODE1[0] x2.x1.x7.floating 1.61e-20
C1452 x2.x2.x5[7].floating a_10112_1956# 1.94e-19
C1453 a_1870_6122# x1.x4.Y 0.00621f
C1454 x1.x3.Y a_3106_6090# 0.143f
C1455 a_2325_6090# a_2932_6494# 0.00187f
C1456 x2.x1.x9.output_stack x2.x4.x5[7].floating 1.33e-19
C1457 vdd a_3041_6494# 7.35e-20
C1458 a_4047_3022# sample_clk 0.00117f
C1459 sample_delay_offset x2.x4.x5[7].floating 0.00542f
C1460 sample_delay_offset a_10024_2094# 3.64e-19
C1461 a_16686_3621# x2.x2.IN 0.0166f
C1462 a_11443_5870# a_11283_6008# 0.0388f
C1463 x2.x3.x5[7].floating a_10112_1680# 2.14e-19
C1464 x2.x4.x10.Y x2.x1.x6.SW 1.5e-20
C1465 a_10137_3483# x2.x2.x2.floating 0.00177f
C1466 a_10137_3207# x2.x3.x4[3].floating 1.17e-19
C1467 vdd a_4047_2819# 0.264f
C1468 CAP_CTRL_CODE2[0] x2.x3.x3[1].floating 3.8e-20
C1469 CAP_CTRL_CODE3[0] CAP_CTRL_CODE2[2] 1.48e-20
C1470 x2.x1.x6.SW x2.x1.x5[7].floating 0.00138f
C1471 vdd CAP_CTRL_CODE0[3] 0.139f
C1472 sample_delay_offset a_4574_6008# 0.0189f
C1473 CAP_CTRL_CODE0[0] CAP_CTRL_CODE1[0] 1.46e-20
C1474 CAP_CTRL_CODE0[2] x2.x4.x7.floating 0.0173f
C1475 a_11308_6983# CAP_CTRL_CODE1[3] 2.69e-19
C1476 a_10137_4035# a_10065_4035# 0.00227f
C1477 a_4574_6008# a_4662_6146# 0.00227f
C1478 x2.x4.x6.SW x1.x2.D 5.6e-21
C1479 vdd x7.A 0.408f
C1480 a_16774_3483# x2.x2.x7.floating 8.52e-19
C1481 a_16686_3621# x2.x2.x4[3].floating 8.29e-19
C1482 x2.x2.x3[1].floating x2.x2.x10.Y 0.00302f
C1483 CAP_CTRL_CODE1[3] x2.x1.x6.floating 0.00506f
C1484 x2.x4.x9.output_stack a_2932_6494# 6.7e-21
C1485 x1.x3.Y a_3340_6116# 2.04e-19
C1486 a_4574_5180# CAP_CTRL_CODE1[0] 6.54e-20
C1487 a_10065_3345# a_10137_3207# 0.00227f
C1488 a_16686_3345# a_16846_3207# 0.0388f
C1489 sample_delay_offset a_16774_3897# 0.00103f
C1490 a_4574_5732# x2.x4.x7.floating 0.00409f
C1491 x2.x1.IN x2.x1.x6.SW 0.0933f
C1492 sample_delay_offset a_4662_5456# 0.00103f
C1493 x2.x4.x6.SW a_4574_5456# 4.74e-20
C1494 a_16846_3483# x2.x2.x6.SW 8.11e-20
C1495 x2.x4.x9.output_stack CAP_CTRL_CODE2[2] 4.06e-21
C1496 CAP_CTRL_CODE0[1] CAP_CTRL_CODE0[0] 2.72f
C1497 x2.x1.IN a_11443_5594# 0.0135f
C1498 a_11283_5180# x2.x1.x6.SW 3.1e-20
C1499 x2.x2.x9.output_stack a_10756_2819# 0.00887f
C1500 a_3813_6132# x2.x4.x6.floating 3.23e-19
C1501 x3.A a_2569_6116# 7.05e-21
C1502 x3.A a_3056_2150# 2.93e-19
C1503 a_11371_5732# x2.x4.x2.floating 2.21e-19
C1504 x2.x2.x6.SW x2.x2.x6.floating 0.13f
C1505 a_10137_3759# a_9977_3621# 0.0388f
C1506 a_16774_3897# a_16846_3759# 0.00227f
C1507 a_4047_3022# a_3553_3025# 1.45e-19
C1508 x7.Y a_3056_2936# 4.39e-19
C1509 sample_delay_offset CAP_CTRL_CODE3[1] 4.51e-19
C1510 x2.x3.x10.Y x2.x2.x5[7].floating 0.00422f
C1511 x2.x3.IN a_10137_4035# 0.0127f
C1512 x3.A CAP_CTRL_CODE1[0] 0.00168f
C1513 a_11283_5456# a_11443_5318# 0.0388f
C1514 a_4662_5456# a_4734_5318# 0.00227f
C1515 x2.x3.x9.output_stack a_10112_2232# 0.0702f
C1516 vdd CAP_CTRL_CODE1[2] 0.0376f
C1517 x2.x4.x9.output_stack a_10472_6534# 0.00887f
C1518 a_2619_6316# a_2465_6482# 0.00943f
C1519 x3.A a_3106_6090# 0.0108f
C1520 x2.x3.x9.output_stack a_10756_2819# 1.18e-20
C1521 x1.x4.Y a_3813_6132# 0.0103f
C1522 a_4574_5180# CAP_CTRL_CODE0[1] 3.36e-19
C1523 a_1704_6122# a_2837_6438# 2.56e-19
C1524 a_11396_7121# x2.x1.x10.Y 4.2e-19
C1525 x2.x3.IN a_10112_1680# 0.00832f
C1526 x2.x4.x9.output_stack x2.x4.x7.floating 0.185f
C1527 vdd a_16846_3483# 4.84e-19
C1528 a_10065_3483# x2.x3.x7.floating 8.52e-19
C1529 a_9977_3897# x2.x2.x2.floating 6.88e-19
C1530 a_9977_3621# x2.x3.x4[3].floating 8.29e-19
C1531 x2.x4.x5[7].floating CAP_CTRL_CODE0[2] 0.00564f
C1532 x2.x2.IN x2.x1.x5[7].floating 0.0199f
C1533 x2.x3.IN CAP_CTRL_CODE2[1] 1.94e-19
C1534 a_4599_7259# x2.x4.x6.floating 0.00996f
C1535 a_11396_7397# x2.x4.x5[7].floating 1.78e-19
C1536 sample_delay_offset a_10137_3207# 0.0189f
C1537 x2.x2.x6.floating a_16821_1680# 0.00578f
C1538 x2.x2.x9.output_stack CAP_CTRL_CODE2[2] 0.322f
C1539 vdd x2.x2.x6.floating 5.78f
C1540 x3.A x2.x3.x3[1].floating 2.07e-20
C1541 a_4687_7397# sample_delay_offset 1.9e-19
C1542 x1.x3.Y x2.x4.x6.floating 8.13e-21
C1543 x2.x4.x2.floating CAP_CTRL_CODE1[2] 0.00611f
C1544 a_11443_5870# x2.x1.x7.floating 0.00959f
C1545 CAP_CTRL_CODE0[2] a_4574_6008# 7.47e-20
C1546 x2.x3.x9.output_stack CAP_CTRL_CODE2[2] 2.46e-20
C1547 a_16774_3897# x2.x2.x7.floating 8.52e-19
C1548 x3.A a_4662_5594# 6.77e-19
C1549 a_10137_3759# x2.x3.x10.Y 4.07e-20
C1550 CAP_CTRL_CODE2[0] x2.x2.x5[7].floating 0.00119f
C1551 vdd x2.x1.x3[1].floating 0.0301f
C1552 vdd x2.x1.x10.Y 2.73f
C1553 x3.A CAP_CTRL_CODE0[1] 0.00191f
C1554 a_10137_4035# CAP_CTRL_CODE1[0] 2.97e-20
C1555 sample_clk_b vss 0.655f
C1556 sample_clk vss 0.615f
C1557 a_16821_1680# vss 0.0953f
C1558 a_10112_1680# vss 0.0334f
C1559 a_16733_1818# vss 0.032f
C1560 a_10024_1818# vss 0.0233f
C1561 a_16821_1956# vss 0.0815f
C1562 a_10112_1956# vss 0.018f
C1563 a_16733_2094# vss 0.0402f
C1564 a_10024_2094# vss 0.0348f
C1565 a_16821_2232# vss 0.0147f
C1566 a_10112_2232# vss 0.00895f
C1567 a_3056_2150# vss 0.531f
C1568 a_2678_2006# vss 0.668f
C1569 x2.x2.x6.floating vss 0.353f
C1570 x2.x2.x5[7].floating vss 0.107p
C1571 a_10756_2819# vss 0.333f
C1572 x2.x2.x6.SW vss 0.299f
C1573 x2.x2.x10.Y vss 2.77f
C1574 x2.x3.x6.floating vss 0.218f
C1575 x2.x3.x5[7].floating vss 0.107p
C1576 a_4047_2819# vss 0.257f
C1577 x2.x3.x6.SW vss 0.282f
C1578 x2.x3.x10.Y vss 2.75f
C1579 x2.x2.x7.floating vss 5.89f
C1580 x2.x2.x4[3].floating vss 21.7f
C1581 x2.x2.x3[1].floating vss 10.9f
C1582 x2.x2.x2.floating vss 6.35f
C1583 CAP_CTRL_CODE2[2] vss 11.3f
C1584 CAP_CTRL_CODE2[1] vss 10.4f
C1585 x2.x3.x7.floating vss 5.82f
C1586 x2.x3.x4[3].floating vss 21.7f
C1587 x2.x3.x3[1].floating vss 10.9f
C1588 x2.x3.x2.floating vss 6.43f
C1589 CAP_CTRL_CODE2[0] vss -12f
C1590 a_16774_3207# vss 6.32e-19
C1591 CAP_CTRL_CODE3[2] vss 3.99f
C1592 CAP_CTRL_CODE3[1] vss 1.27f
C1593 a_3553_3025# vss 0.00235f
C1594 a_3056_2936# vss 0.423f
C1595 x3.Y vss 0.742f
C1596 a_2678_2626# vss 0.664f
C1597 CAP_CTRL_CODE3[0] vss 1.08f
C1598 a_10756_3022# vss 0.275f
C1599 x2.x2.x9.output_stack vss 1.54f
C1600 a_10065_3207# vss 6.56e-19
C1601 x7.A vss 0.618f
C1602 x7.Y vss 0.357f
C1603 a_4047_3022# vss 0.293f
C1604 x2.x3.x9.output_stack vss 1.51f
C1605 a_16846_3207# vss 0.103f
C1606 a_16774_3345# vss 6.69e-19
C1607 a_10137_3207# vss 0.114f
C1608 a_10065_3345# vss 7.81e-19
C1609 a_16774_3483# vss 7.52e-19
C1610 a_16686_3345# vss 0.108f
C1611 a_10065_3483# vss 7.43e-19
C1612 a_9977_3345# vss 0.112f
C1613 a_16846_3483# vss 0.0982f
C1614 a_16774_3621# vss 0.00106f
C1615 a_10137_3483# vss 0.11f
C1616 a_10065_3621# vss 9.98e-19
C1617 a_16774_3759# vss 0.00116f
C1618 a_16686_3621# vss 0.111f
C1619 a_10065_3759# vss 0.00109f
C1620 a_9977_3621# vss 0.114f
C1621 a_16846_3759# vss 0.0991f
C1622 a_16774_3897# vss 0.00129f
C1623 a_10137_3759# vss 0.111f
C1624 a_10065_3897# vss 0.00121f
C1625 a_16774_4035# vss 0.00145f
C1626 a_16686_3897# vss 0.161f
C1627 a_10065_4035# vss 0.00134f
C1628 a_9977_3897# vss 0.165f
C1629 a_16846_4035# vss 0.164f
C1630 a_16774_4173# vss 0.0049f
C1631 a_10137_4035# vss 0.17f
C1632 a_10065_4173# vss 0.005f
C1633 x2.x3.IN vss 1.77f
C1634 a_11371_5180# vss 0.005f
C1635 a_4662_5180# vss 0.00476f
C1636 a_11371_5318# vss 0.00134f
C1637 a_11283_5180# vss 0.17f
C1638 a_4662_5318# vss 0.00134f
C1639 a_4574_5180# vss 0.178f
C1640 a_11443_5318# vss 0.165f
C1641 a_11371_5456# vss 0.00121f
C1642 a_4734_5318# vss 0.165f
C1643 a_4662_5456# vss 0.00121f
C1644 a_11371_5594# vss 0.00109f
C1645 a_11283_5456# vss 0.111f
C1646 a_4662_5594# vss 0.00114f
C1647 a_4574_5456# vss 0.117f
C1648 a_11443_5594# vss 0.114f
C1649 a_11371_5732# vss 9.98e-19
C1650 a_4734_5594# vss 0.115f
C1651 a_4662_5732# vss 0.00157f
C1652 a_11371_5870# vss 7.43e-19
C1653 a_11283_5732# vss 0.11f
C1654 a_4662_5870# vss 7.43e-19
C1655 a_4574_5732# vss 0.106f
C1656 reset vss 0.218f
C1657 set vss 0.239f
C1658 a_11443_5870# vss 0.112f
C1659 a_11371_6008# vss 7.81e-19
C1660 a_4734_5870# vss 0.108f
C1661 a_4662_6008# vss 6.69e-19
C1662 a_11371_6146# vss 6.56e-19
C1663 a_11283_6008# vss 0.114f
C1664 a_4662_6146# vss 6.32e-19
C1665 a_4574_6008# vss 0.0874f
C1666 a_17181_6193# vss 0.256f
C1667 x2.x1.x2.floating vss 6.41f
C1668 x2.x1.x3[1].floating vss 10.9f
C1669 x2.x1.x4[3].floating vss 21.7f
C1670 x2.x1.x7.floating vss 5.82f
C1671 CAP_CTRL_CODE1[0] vss -50.7f
C1672 CAP_CTRL_CODE1[1] vss 12f
C1673 CAP_CTRL_CODE1[2] vss 8.98f
C1674 a_10472_6193# vss 0.276f
C1675 x2.x4.x2.floating vss 6.35f
C1676 x2.x4.x3[1].floating vss 10.9f
C1677 x2.x4.x4[3].floating vss 21.7f
C1678 x2.x4.x7.floating vss 5.88f
C1679 a_3340_6116# vss 0.00104f
C1680 a_3018_6116# vss 8.58e-20
C1681 CAP_CTRL_CODE0[0] vss -4.97f
C1682 CAP_CTRL_CODE0[1] vss 3.9f
C1683 CAP_CTRL_CODE0[2] vss 2.4f
C1684 x2.x1.x5[7].floating vss 0.107p
C1685 x2.x1.x6.floating vss 0.218f
C1686 x2.x2.IN vss 3.33f
C1687 x2.x4.x5[7].floating vss 0.107p
C1688 x2.x4.x6.floating vss 0.379f
C1689 a_2790_6116# vss 0.00109f
C1690 a_2569_6116# vss 9.34e-19
C1691 a_2235_6116# vss 1.36e-19
C1692 a_3222_6482# vss 0.166f
C1693 a_3041_6494# vss 0.00253f
C1694 a_2837_6438# vss 0.0109f
C1695 a_2465_6482# vss 0.189f
C1696 a_2259_6494# vss 0.00244f
C1697 a_2058_6116# vss 0.109f
C1698 a_3813_6132# vss 0.272f
C1699 x1.x4.Y vss 0.632f
C1700 a_2932_6494# vss 0.268f
C1701 a_3106_6090# vss 0.489f
C1702 a_2619_6316# vss 0.422f
C1703 a_2151_6116# vss 0.284f
C1704 x1.x3.Y vss 0.956f
C1705 a_2325_6090# vss 0.303f
C1706 a_1870_6122# vss 0.588f
C1707 x1.x2.D vss 0.354f
C1708 a_1704_6122# vss 0.61f
C1709 clk vss 0.251f
C1710 a_17181_6534# vss 0.319f
C1711 a_10472_6534# vss 0.333f
C1712 x2.x1.x9.output_stack vss 1.53f
C1713 x2.x1.x6.SW vss 0.282f
C1714 x2.x1.x10.Y vss 2.75f
C1715 x2.x4.x9.output_stack vss 1.51f
C1716 CAP_CTRL_CODE1[3] vss 0.211f
C1717 x2.x4.x6.SW vss 0.313f
C1718 x2.x4.x10.Y vss 2.77f
C1719 a_11308_6983# vss 0.00895f
C1720 sample_delay_offset vss 10.5f
C1721 CAP_CTRL_CODE0[3] vss 0.294f
C1722 a_4599_6983# vss 0.0147f
C1723 a_11396_7121# vss 0.0348f
C1724 a_4687_7121# vss 0.0386f
C1725 a_11308_7259# vss 0.0226f
C1726 a_4599_7259# vss 0.049f
C1727 a_11396_7397# vss 0.0236f
C1728 a_4687_7397# vss 0.027f
C1729 a_11308_7535# vss 0.0292f
C1730 x2.x1.IN vss 1.77f
C1731 a_4599_7535# vss 0.0628f
C1732 x3.A vss 3.73f
C1733 vdd vss 0.111p
C1734 CAP_CTRL_CODE1[0].t0 vss 0.0731f
C1735 CAP_CTRL_CODE1[0].n0 vss 66f
C1736 CAP_CTRL_CODE2[0].t0 vss 0.0529f
C1737 CAP_CTRL_CODE2[0].n0 vss 0.923f
C1738 CAP_CTRL_CODE2[0].n1 vss 19.7f
C1739 CAP_CTRL_CODE1[2].t0 vss 0.0455f
C1740 CAP_CTRL_CODE1[2].n0 vss 0.177f
C1741 CAP_CTRL_CODE1[2].t1 vss 0.0455f
C1742 CAP_CTRL_CODE1[2].t2 vss 0.0455f
C1743 CAP_CTRL_CODE1[2].n1 vss 0.181f
C1744 CAP_CTRL_CODE1[2].t3 vss 0.0455f
C1745 CAP_CTRL_CODE1[2].n2 vss 1.69f
C1746 CAP_CTRL_CODE2[1].t0 vss 0.0634f
C1747 CAP_CTRL_CODE2[1].n0 vss 0.243f
C1748 CAP_CTRL_CODE2[1].t1 vss 0.0634f
C1749 CAP_CTRL_CODE0[1].t0 vss 0.0282f
C1750 CAP_CTRL_CODE0[1].t1 vss 0.0281f
C1751 CAP_CTRL_CODE0[1].n0 vss 0.693f
C1752 CAP_CTRL_CODE1[1].t1 vss 0.0648f
C1753 CAP_CTRL_CODE1[1].t0 vss 0.0648f
C1754 CAP_CTRL_CODE1[1].n0 vss 1.78f
C1755 CAP_CTRL_CODE2[2].t2 vss 0.0532f
C1756 CAP_CTRL_CODE2[2].t3 vss 0.0532f
C1757 CAP_CTRL_CODE2[2].n0 vss 0.211f
C1758 CAP_CTRL_CODE2[2].n1 vss 0.702f
C1759 CAP_CTRL_CODE2[2].t0 vss 0.0532f
C1760 CAP_CTRL_CODE2[2].t1 vss 0.0532f
C1761 CAP_CTRL_CODE2[2].n2 vss 1.3f
C1762 x2.x3.x5[7].floating.n0 vss 2.8f
C1763 x2.x3.x5[7].floating.n1 vss 51.4f
C1764 x2.x3.x5[7].floating.n2 vss 2.79f
C1765 x2.x3.x5[7].floating.n3 vss 1.06f
C1766 x2.x3.x5[7].floating.n4 vss 0.367f
C1767 x2.x3.x5[7].floating.n5 vss 1.17f
C1768 x2.x3.x5[7].floating.t7 vss 0.859f
C1769 x2.x3.x5[7].floating.n6 vss 6.5f
C1770 x2.x3.x5[7].floating.n7 vss 1.36f
C1771 x2.x3.x5[7].floating.n8 vss 2.19f
C1772 x2.x3.x5[7].floating.n9 vss 1.06f
C1773 x2.x3.x5[7].floating.n10 vss -15.2f
C1774 x2.x3.x5[7].floating.n11 vss -15.2f
C1775 x2.x3.x5[7].floating.n12 vss -41.6f
C1776 x2.x3.x5[7].floating.n13 vss 0.766f
C1777 x2.x3.x5[7].floating.n14 vss 2.47f
C1778 x2.x3.x5[7].floating.n15 vss 51.5f
C1779 x2.x3.x5[7].floating.n16 vss 2.47f
C1780 x2.x3.x5[7].floating.n17 vss 0.766f
C1781 x2.x3.x5[7].floating.n18 vss -33.5f
C1782 x2.x3.x5[7].floating.n19 vss -4.56f
C1783 x2.x3.x5[7].floating.n20 vss 3.83f
C1784 x2.x3.x5[7].floating.n21 vss -28.9f
C1785 x2.x3.x5[7].floating.n22 vss -7.07f
C1786 x2.x3.x5[7].floating.n23 vss 2.68f
C1787 x2.x3.x5[7].floating.n24 vss 1.06f
C1788 x2.x3.x5[7].floating.n25 vss 0.364f
C1789 x2.x3.x5[7].floating.n26 vss 1.21f
C1790 x2.x3.x5[7].floating.t1 vss 0.859f
C1791 x2.x3.x5[7].floating.n27 vss 6.67f
C1792 x2.x3.x5[7].floating.n28 vss 1.15f
C1793 x2.x3.x5[7].floating.n29 vss 2.17f
C1794 x2.x3.x5[7].floating.n30 vss 1.06f
C1795 x2.x3.x5[7].floating.n31 vss 2.22f
C1796 x2.x3.x5[7].floating.n32 vss -8.01f
C1797 x2.x3.x5[7].floating.n33 vss -28.9f
C1798 x2.x3.x5[7].floating.n34 vss 3.83f
C1799 x2.x3.x5[7].floating.n35 vss -7.07f
C1800 x2.x3.x5[7].floating.n36 vss -28.3f
C1801 x2.x3.x5[7].floating.n37 vss 52.7f
C1802 x2.x3.x5[7].floating.n38 vss 2.47f
C1803 x2.x3.x5[7].floating.n39 vss -28.3f
C1804 x2.x3.x5[7].floating.n40 vss -7.07f
C1805 x2.x3.x5[7].floating.n41 vss 3.83f
C1806 x2.x3.x5[7].floating.n42 vss -28.9f
C1807 x2.x3.x5[7].floating.n43 vss -7.99f
C1808 x2.x3.x5[7].floating.n44 vss 2.22f
C1809 x2.x3.x5[7].floating.n45 vss 1.17f
C1810 x2.x3.x5[7].floating.t0 vss 0.859f
C1811 x2.x3.x5[7].floating.n46 vss 6.5f
C1812 x2.x3.x5[7].floating.n47 vss 1.36f
C1813 x2.x3.x5[7].floating.n48 vss 2.19f
C1814 x2.x3.x5[7].floating.n49 vss 1.06f
C1815 x2.x3.x5[7].floating.n50 vss 0.367f
C1816 x2.x3.x5[7].floating.n51 vss 1.06f
C1817 x2.x3.x5[7].floating.n52 vss 2.79f
C1818 x2.x3.x5[7].floating.n53 vss -28.3f
C1819 x2.x3.x5[7].floating.n54 vss 0.766f
C1820 x2.x3.x5[7].floating.n55 vss -33.5f
C1821 x2.x3.x5[7].floating.n56 vss -4.56f
C1822 x2.x3.x5[7].floating.n57 vss 3.83f
C1823 x2.x3.x5[7].floating.n58 vss -28.9f
C1824 x2.x3.x5[7].floating.n59 vss -7.07f
C1825 x2.x3.x5[7].floating.n60 vss 2.68f
C1826 x2.x3.x5[7].floating.n61 vss -7.07f
C1827 x2.x3.x5[7].floating.n62 vss 3.83f
C1828 x2.x3.x5[7].floating.n63 vss -28.9f
C1829 x2.x3.x5[7].floating.n64 vss -7.99f
C1830 x2.x3.x5[7].floating.n65 vss 2.22f
C1831 x2.x3.x5[7].floating.n66 vss 1.17f
C1832 x2.x3.x5[7].floating.t5 vss 0.859f
C1833 x2.x3.x5[7].floating.n67 vss 6.5f
C1834 x2.x3.x5[7].floating.n68 vss 1.36f
C1835 x2.x3.x5[7].floating.n69 vss 2.19f
C1836 x2.x3.x5[7].floating.n70 vss 1.06f
C1837 x2.x3.x5[7].floating.n71 vss 0.367f
C1838 x2.x3.x5[7].floating.n72 vss 1.06f
C1839 x2.x3.x5[7].floating.n73 vss 2.79f
C1840 x2.x3.x5[7].floating.n74 vss 51.4f
C1841 x2.x3.x5[7].floating.n75 vss 2.8f
C1842 x2.x3.x5[7].floating.n76 vss 1.06f
C1843 x2.x3.x5[7].floating.n77 vss 0.364f
C1844 x2.x3.x5[7].floating.n78 vss 1.21f
C1845 x2.x3.x5[7].floating.t4 vss 0.859f
C1846 x2.x3.x5[7].floating.n79 vss 6.67f
C1847 x2.x3.x5[7].floating.n80 vss 1.15f
C1848 x2.x3.x5[7].floating.n81 vss 2.17f
C1849 x2.x3.x5[7].floating.n82 vss 1.06f
C1850 x2.x3.x5[7].floating.n83 vss 2.22f
C1851 x2.x3.x5[7].floating.n84 vss -8.01f
C1852 x2.x3.x5[7].floating.n85 vss -28.9f
C1853 x2.x3.x5[7].floating.n86 vss 3.83f
C1854 x2.x3.x5[7].floating.n87 vss -7.07f
C1855 x2.x3.x5[7].floating.n88 vss -28.3f
C1856 x2.x3.x5[7].floating.n89 vss 52.7f
C1857 x2.x3.x5[7].floating.n90 vss -28.3f
C1858 x2.x3.x5[7].floating.n91 vss -7.07f
C1859 x2.x3.x5[7].floating.n92 vss 3.83f
C1860 x2.x3.x5[7].floating.n93 vss -28.9f
C1861 x2.x3.x5[7].floating.n94 vss -7.99f
C1862 x2.x3.x5[7].floating.n95 vss 2.22f
C1863 x2.x3.x5[7].floating.n96 vss 1.17f
C1864 x2.x3.x5[7].floating.t2 vss 0.859f
C1865 x2.x3.x5[7].floating.n97 vss 6.5f
C1866 x2.x3.x5[7].floating.n98 vss 1.36f
C1867 x2.x3.x5[7].floating.n99 vss 2.19f
C1868 x2.x3.x5[7].floating.n100 vss 1.06f
C1869 x2.x3.x5[7].floating.n101 vss 0.367f
C1870 x2.x3.x5[7].floating.n102 vss 1.06f
C1871 x2.x3.x5[7].floating.n103 vss 2.79f
C1872 x2.x3.x5[7].floating.n104 vss 51.4f
C1873 x2.x3.x5[7].floating.n105 vss 2.8f
C1874 x2.x3.x5[7].floating.n106 vss 1.06f
C1875 x2.x3.x5[7].floating.n107 vss 0.364f
C1876 x2.x3.x5[7].floating.n108 vss 1.21f
C1877 x2.x3.x5[7].floating.t3 vss 0.859f
C1878 x2.x3.x5[7].floating.n109 vss 6.67f
C1879 x2.x3.x5[7].floating.n110 vss 1.15f
C1880 x2.x3.x5[7].floating.n111 vss 2.17f
C1881 x2.x3.x5[7].floating.n112 vss 1.06f
C1882 x2.x3.x5[7].floating.n113 vss -17.4f
C1883 x2.x3.x5[7].floating.n114 vss -17.2f
C1884 x2.x3.x5[7].floating.n115 vss -43.6f
C1885 x2.x3.x5[7].floating.n116 vss 0.766f
C1886 x2.x3.x5[7].floating.n117 vss 2.47f
C1887 x2.x3.x5[7].floating.n118 vss 51.5f
C1888 x2.x3.x5[7].floating.n119 vss 2.47f
C1889 x2.x3.x5[7].floating.n120 vss 0.766f
C1890 x2.x3.x5[7].floating.n121 vss -33f
C1891 x2.x3.x5[7].floating.n122 vss -5.01f
C1892 x2.x3.x5[7].floating.n123 vss 3.83f
C1893 x2.x3.x5[7].floating.n124 vss -28.9f
C1894 x2.x3.x5[7].floating.n125 vss -7.84f
C1895 x2.x3.x5[7].floating.n126 vss 3.23f
C1896 x2.x3.x5[7].floating.n127 vss 52f
C1897 x2.x3.x5[7].floating.n128 vss 2.68f
C1898 x2.x3.x5[7].floating.n129 vss -7.07f
C1899 x2.x3.x5[7].floating.n130 vss -28.9f
C1900 x2.x3.x5[7].floating.n131 vss 3.83f
C1901 x2.x3.x5[7].floating.n132 vss -4.56f
C1902 x2.x3.x5[7].floating.n133 vss -33.5f
C1903 x2.x3.x5[7].floating.n134 vss 0.766f
C1904 x2.x3.x5[7].floating.n135 vss 2.47f
C1905 x2.x3.x5[7].floating.n136 vss 51.5f
C1906 x2.x3.x5[7].floating.n137 vss 2.47f
C1907 x2.x3.x5[7].floating.n138 vss 0.766f
C1908 x2.x3.x5[7].floating.n139 vss -33f
C1909 x2.x3.x5[7].floating.n140 vss -5.01f
C1910 x2.x3.x5[7].floating.n141 vss 3.83f
C1911 x2.x3.x5[7].floating.n142 vss -28.9f
C1912 x2.x3.x5[7].floating.n143 vss -7.84f
C1913 x2.x3.x5[7].floating.n144 vss 3.23f
C1914 x2.x3.x5[7].floating.n145 vss 52f
C1915 x2.x3.x5[7].floating.n146 vss 52.7f
C1916 x2.x3.x5[7].floating.n147 vss -28.3f
C1917 x2.x3.x5[7].floating.n148 vss -7.07f
C1918 x2.x3.x5[7].floating.n149 vss 3.83f
C1919 x2.x3.x5[7].floating.n150 vss -28.9f
C1920 x2.x3.x5[7].floating.n151 vss -8.01f
C1921 x2.x3.x5[7].floating.n152 vss 2.22f
C1922 x2.x3.x5[7].floating.n153 vss 1.21f
C1923 x2.x3.x5[7].floating.t6 vss 0.859f
C1924 x2.x3.x5[7].floating.n154 vss 6.67f
C1925 x2.x3.x5[7].floating.n155 vss 1.15f
C1926 x2.x3.x5[7].floating.n156 vss 2.17f
C1927 x2.x3.x5[7].floating.n157 vss 1.06f
C1928 x2.x3.x5[7].floating.n158 vss 0.364f
C1929 x2.x3.x5[7].floating.n159 vss 1.06f
C1930 x2.x3.x5[7].floating.n160 vss 2.8f
C1931 x2.x3.x5[7].floating.n161 vss 51.4f
C1932 x2.x3.x5[7].floating.n162 vss 51.5f
C1933 x2.x3.x5[7].floating.n163 vss 2.47f
C1934 x2.x3.x5[7].floating.n164 vss 0.766f
C1935 x2.x3.x5[7].floating.n165 vss -33f
C1936 x2.x3.x5[7].floating.n166 vss -5.01f
C1937 x2.x3.x5[7].floating.n167 vss 3.83f
C1938 x2.x3.x5[7].floating.n168 vss -28.9f
C1939 x2.x3.x5[7].floating.n169 vss -7.84f
C1940 x2.x3.x5[7].floating.n170 vss 3.23f
C1941 x2.x3.x5[7].floating.n171 vss 52f
C1942 x2.x3.x10.Y.n0 vss 0.0359f
C1943 x2.x3.x10.Y.t0 vss 0.0526f
C1944 x2.x3.x10.Y.n1 vss 0.0169f
C1945 x2.x3.x10.Y.n2 vss 0.00704f
C1946 x2.x3.x10.Y.t1 vss 0.0181f
C1947 x2.x3.x10.Y.n3 vss 0.0188f
C1948 x2.x3.x10.Y.n4 vss 0.019f
C1949 x2.x3.x10.Y.n5 vss 0.221f
C1950 x2.x3.x10.Y.t2 vss 0.0167f
C1951 x2.x3.x10.Y.t8 vss 0.0167f
C1952 x2.x3.x10.Y.t9 vss 0.0167f
C1953 x2.x3.x10.Y.t3 vss 0.0167f
C1954 x2.x3.x10.Y.t4 vss 0.0167f
C1955 x2.x3.x10.Y.t5 vss 0.0167f
C1956 x2.x3.x10.Y.t7 vss 0.0167f
C1957 x2.x3.x10.Y.t6 vss 0.0167f
C1958 CAP_CTRL_CODE3[2].t3 vss 0.0192f
C1959 CAP_CTRL_CODE3[2].t0 vss 0.0192f
C1960 CAP_CTRL_CODE3[2].n0 vss 0.0762f
C1961 CAP_CTRL_CODE3[2].n1 vss 0.253f
C1962 CAP_CTRL_CODE3[2].t1 vss 0.0192f
C1963 CAP_CTRL_CODE3[2].t2 vss 0.0192f
C1964 CAP_CTRL_CODE3[2].n2 vss 0.425f
C1965 sample_delay_offset.n0 vss 0.00686f
C1966 sample_delay_offset.t0 vss 0.0258f
C1967 sample_delay_offset.t8 vss 0.0162f
C1968 sample_delay_offset.n1 vss 0.0486f
C1969 sample_delay_offset.n2 vss 0.00969f
C1970 sample_delay_offset.n3 vss 0.00292f
C1971 sample_delay_offset.n4 vss 0.00236f
C1972 sample_delay_offset.n5 vss 0.0027f
C1973 sample_delay_offset.n6 vss 0.0114f
C1974 sample_delay_offset.n7 vss 0.117f
C1975 sample_delay_offset.n8 vss 0.258f
C1976 sample_delay_offset.t1 vss 0.0137f
C1977 sample_delay_offset.n9 vss 0.202f
C1978 sample_delay_offset.n10 vss 1.44f
C1979 sample_delay_offset.n11 vss 0.00152f
C1980 sample_delay_offset.t3 vss 0.0258f
C1981 sample_delay_offset.t9 vss 0.0156f
C1982 sample_delay_offset.n12 vss 0.0191f
C1983 sample_delay_offset.n13 vss 0.0299f
C1984 sample_delay_offset.n14 vss 0.0634f
C1985 sample_delay_offset.n15 vss 0.0226f
C1986 sample_delay_offset.n16 vss 0.234f
C1987 sample_delay_offset.n17 vss 0.106f
C1988 sample_delay_offset.t2 vss 0.0137f
C1989 sample_delay_offset.n18 vss 0.3f
C1990 sample_delay_offset.n19 vss 3.15f
C1991 sample_delay_offset.n20 vss 0.00686f
C1992 sample_delay_offset.t4 vss 0.0258f
C1993 sample_delay_offset.t11 vss 0.0162f
C1994 sample_delay_offset.n21 vss 0.0486f
C1995 sample_delay_offset.n22 vss 0.00969f
C1996 sample_delay_offset.n23 vss 0.00292f
C1997 sample_delay_offset.n24 vss 0.00236f
C1998 sample_delay_offset.n25 vss 0.0027f
C1999 sample_delay_offset.n26 vss 0.0114f
C2000 sample_delay_offset.n27 vss 0.117f
C2001 sample_delay_offset.n28 vss 0.258f
C2002 sample_delay_offset.t7 vss 0.0137f
C2003 sample_delay_offset.n29 vss 0.202f
C2004 sample_delay_offset.n30 vss 0.33f
C2005 sample_delay_offset.n31 vss 2.41f
C2006 sample_delay_offset.n32 vss 0.00152f
C2007 sample_delay_offset.t6 vss 0.0258f
C2008 sample_delay_offset.t10 vss 0.0156f
C2009 sample_delay_offset.n33 vss 0.0191f
C2010 sample_delay_offset.n34 vss 0.0299f
C2011 sample_delay_offset.n35 vss 0.0634f
C2012 sample_delay_offset.n36 vss 0.0226f
C2013 sample_delay_offset.n37 vss 0.234f
C2014 sample_delay_offset.n38 vss 0.106f
C2015 sample_delay_offset.t5 vss 0.0137f
C2016 sample_delay_offset.n39 vss 0.387f
C2017 sample_delay_offset.n40 vss 1.94f
C2018 x2.x2.x5[7].floating.n0 vss 2.8f
C2019 x2.x2.x5[7].floating.n1 vss 51.4f
C2020 x2.x2.x5[7].floating.n2 vss 2.79f
C2021 x2.x2.x5[7].floating.n3 vss 1.06f
C2022 x2.x2.x5[7].floating.n4 vss 0.367f
C2023 x2.x2.x5[7].floating.n5 vss 1.17f
C2024 x2.x2.x5[7].floating.t0 vss 0.859f
C2025 x2.x2.x5[7].floating.n6 vss 6.5f
C2026 x2.x2.x5[7].floating.n7 vss 1.36f
C2027 x2.x2.x5[7].floating.n8 vss 2.19f
C2028 x2.x2.x5[7].floating.n9 vss 1.06f
C2029 x2.x2.x5[7].floating.n10 vss -15.2f
C2030 x2.x2.x5[7].floating.n11 vss -15.2f
C2031 x2.x2.x5[7].floating.n12 vss -41.6f
C2032 x2.x2.x5[7].floating.n13 vss 0.766f
C2033 x2.x2.x5[7].floating.n14 vss 2.47f
C2034 x2.x2.x5[7].floating.n15 vss 51.5f
C2035 x2.x2.x5[7].floating.n16 vss 2.47f
C2036 x2.x2.x5[7].floating.n17 vss 0.766f
C2037 x2.x2.x5[7].floating.n18 vss -33.5f
C2038 x2.x2.x5[7].floating.n19 vss -4.56f
C2039 x2.x2.x5[7].floating.n20 vss 3.83f
C2040 x2.x2.x5[7].floating.n21 vss -28.9f
C2041 x2.x2.x5[7].floating.n22 vss -7.07f
C2042 x2.x2.x5[7].floating.n23 vss 2.68f
C2043 x2.x2.x5[7].floating.n24 vss 1.06f
C2044 x2.x2.x5[7].floating.n25 vss 0.364f
C2045 x2.x2.x5[7].floating.n26 vss 1.21f
C2046 x2.x2.x5[7].floating.t4 vss 0.859f
C2047 x2.x2.x5[7].floating.n27 vss 6.67f
C2048 x2.x2.x5[7].floating.n28 vss 1.15f
C2049 x2.x2.x5[7].floating.n29 vss 2.17f
C2050 x2.x2.x5[7].floating.n30 vss 1.06f
C2051 x2.x2.x5[7].floating.n31 vss 2.22f
C2052 x2.x2.x5[7].floating.n32 vss -8.01f
C2053 x2.x2.x5[7].floating.n33 vss -28.9f
C2054 x2.x2.x5[7].floating.n34 vss 3.83f
C2055 x2.x2.x5[7].floating.n35 vss -7.07f
C2056 x2.x2.x5[7].floating.n36 vss -28.3f
C2057 x2.x2.x5[7].floating.n37 vss 52.7f
C2058 x2.x2.x5[7].floating.n38 vss -28.3f
C2059 x2.x2.x5[7].floating.n39 vss -7.07f
C2060 x2.x2.x5[7].floating.n40 vss 3.83f
C2061 x2.x2.x5[7].floating.n41 vss -28.9f
C2062 x2.x2.x5[7].floating.n42 vss -7.99f
C2063 x2.x2.x5[7].floating.n43 vss 2.22f
C2064 x2.x2.x5[7].floating.n44 vss 1.17f
C2065 x2.x2.x5[7].floating.t5 vss 0.859f
C2066 x2.x2.x5[7].floating.n45 vss 6.5f
C2067 x2.x2.x5[7].floating.n46 vss 1.36f
C2068 x2.x2.x5[7].floating.n47 vss 2.19f
C2069 x2.x2.x5[7].floating.n48 vss 1.06f
C2070 x2.x2.x5[7].floating.n49 vss 0.367f
C2071 x2.x2.x5[7].floating.n50 vss 1.06f
C2072 x2.x2.x5[7].floating.n51 vss 2.79f
C2073 x2.x2.x5[7].floating.n52 vss 51.4f
C2074 x2.x2.x5[7].floating.n53 vss 2.8f
C2075 x2.x2.x5[7].floating.n54 vss 1.06f
C2076 x2.x2.x5[7].floating.n55 vss 0.364f
C2077 x2.x2.x5[7].floating.n56 vss 1.21f
C2078 x2.x2.x5[7].floating.t2 vss 0.859f
C2079 x2.x2.x5[7].floating.n57 vss 6.67f
C2080 x2.x2.x5[7].floating.n58 vss 1.15f
C2081 x2.x2.x5[7].floating.n59 vss 2.17f
C2082 x2.x2.x5[7].floating.n60 vss 1.06f
C2083 x2.x2.x5[7].floating.n61 vss 2.22f
C2084 x2.x2.x5[7].floating.n62 vss -8.01f
C2085 x2.x2.x5[7].floating.n63 vss -28.9f
C2086 x2.x2.x5[7].floating.n64 vss 3.83f
C2087 x2.x2.x5[7].floating.n65 vss -7.07f
C2088 x2.x2.x5[7].floating.n66 vss -28.3f
C2089 x2.x2.x5[7].floating.n67 vss 52.7f
C2090 x2.x2.x5[7].floating.n68 vss -28.3f
C2091 x2.x2.x5[7].floating.n69 vss -7.07f
C2092 x2.x2.x5[7].floating.n70 vss 3.83f
C2093 x2.x2.x5[7].floating.n71 vss -28.9f
C2094 x2.x2.x5[7].floating.n72 vss -7.99f
C2095 x2.x2.x5[7].floating.n73 vss 2.22f
C2096 x2.x2.x5[7].floating.n74 vss 1.17f
C2097 x2.x2.x5[7].floating.t3 vss 0.859f
C2098 x2.x2.x5[7].floating.n75 vss 6.5f
C2099 x2.x2.x5[7].floating.n76 vss 1.36f
C2100 x2.x2.x5[7].floating.n77 vss 2.19f
C2101 x2.x2.x5[7].floating.n78 vss 1.06f
C2102 x2.x2.x5[7].floating.n79 vss 0.367f
C2103 x2.x2.x5[7].floating.n80 vss 1.06f
C2104 x2.x2.x5[7].floating.n81 vss 2.79f
C2105 x2.x2.x5[7].floating.n82 vss 51.4f
C2106 x2.x2.x5[7].floating.n83 vss 2.8f
C2107 x2.x2.x5[7].floating.n84 vss 1.06f
C2108 x2.x2.x5[7].floating.n85 vss 0.364f
C2109 x2.x2.x5[7].floating.n86 vss 1.21f
C2110 x2.x2.x5[7].floating.t1 vss 0.859f
C2111 x2.x2.x5[7].floating.n87 vss 6.67f
C2112 x2.x2.x5[7].floating.n88 vss 1.15f
C2113 x2.x2.x5[7].floating.n89 vss 2.17f
C2114 x2.x2.x5[7].floating.n90 vss 1.06f
C2115 x2.x2.x5[7].floating.n91 vss 2.22f
C2116 x2.x2.x5[7].floating.n92 vss -8.01f
C2117 x2.x2.x5[7].floating.n93 vss -28.9f
C2118 x2.x2.x5[7].floating.n94 vss 3.83f
C2119 x2.x2.x5[7].floating.n95 vss -7.07f
C2120 x2.x2.x5[7].floating.n96 vss -28.3f
C2121 x2.x2.x5[7].floating.n97 vss 52.7f
C2122 x2.x2.x5[7].floating.n98 vss -28.3f
C2123 x2.x2.x5[7].floating.n99 vss -7.07f
C2124 x2.x2.x5[7].floating.n100 vss 3.83f
C2125 x2.x2.x5[7].floating.n101 vss -28.9f
C2126 x2.x2.x5[7].floating.n102 vss -7.99f
C2127 x2.x2.x5[7].floating.n103 vss 2.22f
C2128 x2.x2.x5[7].floating.n104 vss 1.17f
C2129 x2.x2.x5[7].floating.t7 vss 0.859f
C2130 x2.x2.x5[7].floating.n105 vss 6.5f
C2131 x2.x2.x5[7].floating.n106 vss 1.36f
C2132 x2.x2.x5[7].floating.n107 vss 2.19f
C2133 x2.x2.x5[7].floating.n108 vss 1.06f
C2134 x2.x2.x5[7].floating.n109 vss 0.367f
C2135 x2.x2.x5[7].floating.n110 vss 1.06f
C2136 x2.x2.x5[7].floating.n111 vss 2.79f
C2137 x2.x2.x5[7].floating.n112 vss 51.4f
C2138 x2.x2.x5[7].floating.n113 vss 2.8f
C2139 x2.x2.x5[7].floating.n114 vss 1.06f
C2140 x2.x2.x5[7].floating.n115 vss 0.366f
C2141 x2.x2.x5[7].floating.t6 vss 0.859f
C2142 x2.x2.x5[7].floating.n116 vss 7.13f
C2143 x2.x2.x5[7].floating.n117 vss 1.21f
C2144 x2.x2.x5[7].floating.n118 vss 1.16f
C2145 x2.x2.x5[7].floating.n119 vss 1.7f
C2146 x2.x2.x5[7].floating.n120 vss 1.06f
C2147 x2.x2.x5[7].floating.n121 vss -17.4f
C2148 x2.x2.x5[7].floating.n122 vss -17.2f
C2149 x2.x2.x5[7].floating.n123 vss -43.6f
C2150 x2.x2.x5[7].floating.n124 vss 0.766f
C2151 x2.x2.x5[7].floating.n125 vss 2.47f
C2152 x2.x2.x5[7].floating.n126 vss 51.5f
C2153 x2.x2.x5[7].floating.n127 vss 2.47f
C2154 x2.x2.x5[7].floating.n128 vss 0.766f
C2155 x2.x2.x5[7].floating.n129 vss -33f
C2156 x2.x2.x5[7].floating.n130 vss -5.01f
C2157 x2.x2.x5[7].floating.n131 vss 3.83f
C2158 x2.x2.x5[7].floating.n132 vss -28.9f
C2159 x2.x2.x5[7].floating.n133 vss -7.84f
C2160 x2.x2.x5[7].floating.n134 vss 3.23f
C2161 x2.x2.x5[7].floating.n135 vss 52f
C2162 x2.x2.x5[7].floating.n136 vss 2.68f
C2163 x2.x2.x5[7].floating.n137 vss -7.07f
C2164 x2.x2.x5[7].floating.n138 vss -28.9f
C2165 x2.x2.x5[7].floating.n139 vss 3.83f
C2166 x2.x2.x5[7].floating.n140 vss -4.56f
C2167 x2.x2.x5[7].floating.n141 vss -33.5f
C2168 x2.x2.x5[7].floating.n142 vss 0.766f
C2169 x2.x2.x5[7].floating.n143 vss 2.47f
C2170 x2.x2.x5[7].floating.n144 vss 51.5f
C2171 x2.x2.x5[7].floating.n145 vss 2.47f
C2172 x2.x2.x5[7].floating.n146 vss 0.766f
C2173 x2.x2.x5[7].floating.n147 vss -33f
C2174 x2.x2.x5[7].floating.n148 vss -5.01f
C2175 x2.x2.x5[7].floating.n149 vss 3.83f
C2176 x2.x2.x5[7].floating.n150 vss -28.9f
C2177 x2.x2.x5[7].floating.n151 vss -7.84f
C2178 x2.x2.x5[7].floating.n152 vss 3.23f
C2179 x2.x2.x5[7].floating.n153 vss 52f
C2180 x2.x2.x5[7].floating.n154 vss 2.68f
C2181 x2.x2.x5[7].floating.n155 vss -7.07f
C2182 x2.x2.x5[7].floating.n156 vss -28.9f
C2183 x2.x2.x5[7].floating.n157 vss 3.83f
C2184 x2.x2.x5[7].floating.n158 vss -4.56f
C2185 x2.x2.x5[7].floating.n159 vss -33.5f
C2186 x2.x2.x5[7].floating.n160 vss 0.766f
C2187 x2.x2.x5[7].floating.n161 vss 2.47f
C2188 x2.x2.x5[7].floating.n162 vss 51.5f
C2189 x2.x2.x5[7].floating.n163 vss 2.47f
C2190 x2.x2.x5[7].floating.n164 vss 0.766f
C2191 x2.x2.x5[7].floating.n165 vss -33f
C2192 x2.x2.x5[7].floating.n166 vss -5.01f
C2193 x2.x2.x5[7].floating.n167 vss 3.83f
C2194 x2.x2.x5[7].floating.n168 vss -28.9f
C2195 x2.x2.x5[7].floating.n169 vss -7.84f
C2196 x2.x2.x5[7].floating.n170 vss 3.23f
C2197 x2.x2.x5[7].floating.n171 vss 52f
C2198 x2.x2.x10.Y.n0 vss 0.0359f
C2199 x2.x2.x10.Y.t0 vss 0.0526f
C2200 x2.x2.x10.Y.n1 vss 0.0169f
C2201 x2.x2.x10.Y.n2 vss 0.00704f
C2202 x2.x2.x10.Y.t1 vss 0.0181f
C2203 x2.x2.x10.Y.n3 vss 0.0188f
C2204 x2.x2.x10.Y.n4 vss 0.019f
C2205 x2.x2.x10.Y.n5 vss 0.221f
C2206 x2.x2.x10.Y.t9 vss 0.0167f
C2207 x2.x2.x10.Y.t5 vss 0.0167f
C2208 x2.x2.x10.Y.t4 vss 0.0167f
C2209 x2.x2.x10.Y.t7 vss 0.0167f
C2210 x2.x2.x10.Y.t6 vss 0.0167f
C2211 x2.x2.x10.Y.t8 vss 0.0167f
C2212 x2.x2.x10.Y.t2 vss 0.0167f
C2213 x2.x2.x10.Y.t3 vss 0.0167f
C2214 x2.x4.x5[7].floating.n0 vss -7.99f
C2215 x2.x4.x5[7].floating.n1 vss -28.9f
C2216 x2.x4.x5[7].floating.n2 vss 3.83f
C2217 x2.x4.x5[7].floating.n3 vss -7.07f
C2218 x2.x4.x5[7].floating.n4 vss -28.3f
C2219 x2.x4.x5[7].floating.n5 vss 52.7f
C2220 x2.x4.x5[7].floating.n6 vss -28.3f
C2221 x2.x4.x5[7].floating.n7 vss -7.07f
C2222 x2.x4.x5[7].floating.n8 vss 3.83f
C2223 x2.x4.x5[7].floating.n9 vss -28.9f
C2224 x2.x4.x5[7].floating.n10 vss -8.01f
C2225 x2.x4.x5[7].floating.n11 vss 2.21f
C2226 x2.x4.x5[7].floating.t3 vss 0.859f
C2227 x2.x4.x5[7].floating.n12 vss 6.65f
C2228 x2.x4.x5[7].floating.n13 vss 1.21f
C2229 x2.x4.x5[7].floating.n14 vss 1.17f
C2230 x2.x4.x5[7].floating.n15 vss 2.18f
C2231 x2.x4.x5[7].floating.n16 vss 1.06f
C2232 x2.x4.x5[7].floating.n17 vss 0.366f
C2233 x2.x4.x5[7].floating.n18 vss 1.06f
C2234 x2.x4.x5[7].floating.n19 vss 2.8f
C2235 x2.x4.x5[7].floating.n20 vss 51.4f
C2236 x2.x4.x5[7].floating.n21 vss 2.79f
C2237 x2.x4.x5[7].floating.n22 vss 1.06f
C2238 x2.x4.x5[7].floating.n23 vss 0.364f
C2239 x2.x4.x5[7].floating.t4 vss 0.859f
C2240 x2.x4.x5[7].floating.n24 vss 6.48f
C2241 x2.x4.x5[7].floating.n25 vss 1.15f
C2242 x2.x4.x5[7].floating.n26 vss 1.36f
C2243 x2.x4.x5[7].floating.n27 vss 2.2f
C2244 x2.x4.x5[7].floating.n28 vss 1.06f
C2245 x2.x4.x5[7].floating.n29 vss 2.23f
C2246 x2.x4.x5[7].floating.n30 vss -7.99f
C2247 x2.x4.x5[7].floating.n31 vss -28.9f
C2248 x2.x4.x5[7].floating.n32 vss 3.83f
C2249 x2.x4.x5[7].floating.n33 vss -7.07f
C2250 x2.x4.x5[7].floating.n34 vss -28.3f
C2251 x2.x4.x5[7].floating.n35 vss 52.7f
C2252 x2.x4.x5[7].floating.n36 vss -28.3f
C2253 x2.x4.x5[7].floating.n37 vss -7.07f
C2254 x2.x4.x5[7].floating.n38 vss 3.83f
C2255 x2.x4.x5[7].floating.n39 vss -28.9f
C2256 x2.x4.x5[7].floating.n40 vss -8.01f
C2257 x2.x4.x5[7].floating.n41 vss 2.21f
C2258 x2.x4.x5[7].floating.t5 vss 0.859f
C2259 x2.x4.x5[7].floating.n42 vss 6.65f
C2260 x2.x4.x5[7].floating.n43 vss 1.21f
C2261 x2.x4.x5[7].floating.n44 vss 1.17f
C2262 x2.x4.x5[7].floating.n45 vss 2.18f
C2263 x2.x4.x5[7].floating.n46 vss 1.06f
C2264 x2.x4.x5[7].floating.n47 vss 0.366f
C2265 x2.x4.x5[7].floating.n48 vss 1.06f
C2266 x2.x4.x5[7].floating.n49 vss 2.8f
C2267 x2.x4.x5[7].floating.n50 vss 51.4f
C2268 x2.x4.x5[7].floating.n51 vss 2.68f
C2269 x2.x4.x5[7].floating.n52 vss -7.07f
C2270 x2.x4.x5[7].floating.n53 vss -28.9f
C2271 x2.x4.x5[7].floating.n54 vss 3.83f
C2272 x2.x4.x5[7].floating.n55 vss -4.56f
C2273 x2.x4.x5[7].floating.n56 vss -33.5f
C2274 x2.x4.x5[7].floating.n57 vss 0.766f
C2275 x2.x4.x5[7].floating.n58 vss 2.47f
C2276 x2.x4.x5[7].floating.n59 vss 51.5f
C2277 x2.x4.x5[7].floating.n60 vss 2.47f
C2278 x2.x4.x5[7].floating.n61 vss 0.766f
C2279 x2.x4.x5[7].floating.n62 vss -41.6f
C2280 x2.x4.x5[7].floating.n63 vss -15.2f
C2281 x2.x4.x5[7].floating.n64 vss -15.2f
C2282 x2.x4.x5[7].floating.t1 vss 0.859f
C2283 x2.x4.x5[7].floating.n65 vss 6.48f
C2284 x2.x4.x5[7].floating.n66 vss 1.15f
C2285 x2.x4.x5[7].floating.n67 vss 1.36f
C2286 x2.x4.x5[7].floating.n68 vss 2.2f
C2287 x2.x4.x5[7].floating.n69 vss 1.06f
C2288 x2.x4.x5[7].floating.n70 vss 0.364f
C2289 x2.x4.x5[7].floating.n71 vss 1.06f
C2290 x2.x4.x5[7].floating.n72 vss 2.79f
C2291 x2.x4.x5[7].floating.n73 vss 51.4f
C2292 x2.x4.x5[7].floating.n74 vss 2.8f
C2293 x2.x4.x5[7].floating.n75 vss 1.06f
C2294 x2.x4.x5[7].floating.n76 vss 0.366f
C2295 x2.x4.x5[7].floating.t0 vss 0.859f
C2296 x2.x4.x5[7].floating.n77 vss 6.65f
C2297 x2.x4.x5[7].floating.n78 vss 1.21f
C2298 x2.x4.x5[7].floating.n79 vss 1.17f
C2299 x2.x4.x5[7].floating.n80 vss 2.18f
C2300 x2.x4.x5[7].floating.n81 vss 1.06f
C2301 x2.x4.x5[7].floating.n82 vss 2.21f
C2302 x2.x4.x5[7].floating.n83 vss -8.01f
C2303 x2.x4.x5[7].floating.n84 vss -28.9f
C2304 x2.x4.x5[7].floating.n85 vss 3.83f
C2305 x2.x4.x5[7].floating.n86 vss -7.07f
C2306 x2.x4.x5[7].floating.n87 vss -28.3f
C2307 x2.x4.x5[7].floating.n88 vss 2.79f
C2308 x2.x4.x5[7].floating.n89 vss 1.06f
C2309 x2.x4.x5[7].floating.n90 vss 0.364f
C2310 x2.x4.x5[7].floating.t6 vss 0.859f
C2311 x2.x4.x5[7].floating.n91 vss 6.48f
C2312 x2.x4.x5[7].floating.n92 vss 1.15f
C2313 x2.x4.x5[7].floating.n93 vss 1.36f
C2314 x2.x4.x5[7].floating.n94 vss 2.2f
C2315 x2.x4.x5[7].floating.n95 vss 1.06f
C2316 x2.x4.x5[7].floating.n96 vss 2.23f
C2317 x2.x4.x5[7].floating.n97 vss -7.99f
C2318 x2.x4.x5[7].floating.n98 vss -28.9f
C2319 x2.x4.x5[7].floating.n99 vss 3.83f
C2320 x2.x4.x5[7].floating.n100 vss -7.07f
C2321 x2.x4.x5[7].floating.n101 vss -28.3f
C2322 x2.x4.x5[7].floating.n102 vss 52.7f
C2323 x2.x4.x5[7].floating.n103 vss 52f
C2324 x2.x4.x5[7].floating.n104 vss 3.23f
C2325 x2.x4.x5[7].floating.n105 vss -7.84f
C2326 x2.x4.x5[7].floating.n106 vss -28.9f
C2327 x2.x4.x5[7].floating.n107 vss 3.83f
C2328 x2.x4.x5[7].floating.n108 vss -5.01f
C2329 x2.x4.x5[7].floating.n109 vss -33f
C2330 x2.x4.x5[7].floating.n110 vss 0.766f
C2331 x2.x4.x5[7].floating.n111 vss 2.47f
C2332 x2.x4.x5[7].floating.n112 vss 51.5f
C2333 x2.x4.x5[7].floating.n113 vss 2.47f
C2334 x2.x4.x5[7].floating.n114 vss 0.766f
C2335 x2.x4.x5[7].floating.n115 vss -33.5f
C2336 x2.x4.x5[7].floating.n116 vss -4.56f
C2337 x2.x4.x5[7].floating.n117 vss 3.83f
C2338 x2.x4.x5[7].floating.n118 vss -28.9f
C2339 x2.x4.x5[7].floating.n119 vss -7.07f
C2340 x2.x4.x5[7].floating.n120 vss 2.68f
C2341 x2.x4.x5[7].floating.n121 vss 52f
C2342 x2.x4.x5[7].floating.n122 vss 3.23f
C2343 x2.x4.x5[7].floating.n123 vss -7.84f
C2344 x2.x4.x5[7].floating.n124 vss -28.9f
C2345 x2.x4.x5[7].floating.n125 vss 3.83f
C2346 x2.x4.x5[7].floating.n126 vss -5.01f
C2347 x2.x4.x5[7].floating.n127 vss -33f
C2348 x2.x4.x5[7].floating.n128 vss 0.766f
C2349 x2.x4.x5[7].floating.n129 vss 2.47f
C2350 x2.x4.x5[7].floating.n130 vss 51.5f
C2351 x2.x4.x5[7].floating.n131 vss 2.47f
C2352 x2.x4.x5[7].floating.n132 vss 0.766f
C2353 x2.x4.x5[7].floating.n133 vss -33.5f
C2354 x2.x4.x5[7].floating.n134 vss -4.56f
C2355 x2.x4.x5[7].floating.n135 vss 3.83f
C2356 x2.x4.x5[7].floating.n136 vss -28.9f
C2357 x2.x4.x5[7].floating.n137 vss -7.07f
C2358 x2.x4.x5[7].floating.n138 vss 2.68f
C2359 x2.x4.x5[7].floating.n139 vss 52f
C2360 x2.x4.x5[7].floating.n140 vss 3.23f
C2361 x2.x4.x5[7].floating.n141 vss 2.23f
C2362 x2.x4.x5[7].floating.t2 vss 0.859f
C2363 x2.x4.x5[7].floating.n142 vss 6.48f
C2364 x2.x4.x5[7].floating.n143 vss 1.15f
C2365 x2.x4.x5[7].floating.n144 vss 1.36f
C2366 x2.x4.x5[7].floating.n145 vss 2.2f
C2367 x2.x4.x5[7].floating.n146 vss 1.06f
C2368 x2.x4.x5[7].floating.n147 vss 0.364f
C2369 x2.x4.x5[7].floating.n148 vss 1.06f
C2370 x2.x4.x5[7].floating.n149 vss 2.79f
C2371 x2.x4.x5[7].floating.n150 vss 51.4f
C2372 x2.x4.x5[7].floating.n151 vss 2.8f
C2373 x2.x4.x5[7].floating.n152 vss 1.06f
C2374 x2.x4.x5[7].floating.n153 vss 0.366f
C2375 x2.x4.x5[7].floating.t7 vss 0.859f
C2376 x2.x4.x5[7].floating.n154 vss 7.16f
C2377 x2.x4.x5[7].floating.n155 vss 1.21f
C2378 x2.x4.x5[7].floating.n156 vss 1.17f
C2379 x2.x4.x5[7].floating.n157 vss 1.67f
C2380 x2.x4.x5[7].floating.n158 vss 1.06f
C2381 x2.x4.x5[7].floating.n159 vss -17.4f
C2382 x2.x4.x5[7].floating.n160 vss -17.2f
C2383 x2.x4.x5[7].floating.n161 vss -43.6f
C2384 x2.x4.x5[7].floating.n162 vss 0.766f
C2385 x2.x4.x5[7].floating.n163 vss 2.47f
C2386 x2.x4.x5[7].floating.n164 vss 51.5f
C2387 x2.x4.x5[7].floating.n165 vss 2.47f
C2388 x2.x4.x5[7].floating.n166 vss 0.766f
C2389 x2.x4.x5[7].floating.n167 vss -33f
C2390 x2.x4.x5[7].floating.n168 vss -5.01f
C2391 x2.x4.x5[7].floating.n169 vss 3.83f
C2392 x2.x4.x5[7].floating.n170 vss -28.9f
C2393 x2.x4.x5[7].floating.n171 vss -7.84f
C2394 x2.x4.x10.Y.t0 vss 0.0462f
C2395 x2.x4.x10.Y.t8 vss 0.0167f
C2396 x2.x4.x10.Y.t9 vss 0.0167f
C2397 x2.x4.x10.Y.t3 vss 0.0167f
C2398 x2.x4.x10.Y.t4 vss 0.0167f
C2399 x2.x4.x10.Y.t5 vss 0.0167f
C2400 x2.x4.x10.Y.t6 vss 0.0167f
C2401 x2.x4.x10.Y.t7 vss 0.0167f
C2402 x2.x4.x10.Y.t2 vss 0.0167f
C2403 x2.x4.x10.Y.n0 vss 0.222f
C2404 x2.x4.x10.Y.n1 vss 0.0366f
C2405 x2.x4.x10.Y.t1 vss 0.0174f
C2406 x2.x4.x10.Y.n2 vss 0.0188f
C2407 x2.x4.x10.Y.n3 vss 0.0186f
C2408 x2.x4.x10.Y.n4 vss 0.0151f
C2409 x2.x4.x10.Y.n5 vss 0.0211f
C2410 x2.x1.x5[7].floating.n0 vss -7.99f
C2411 x2.x1.x5[7].floating.n1 vss -28.9f
C2412 x2.x1.x5[7].floating.n2 vss 3.83f
C2413 x2.x1.x5[7].floating.n3 vss -7.07f
C2414 x2.x1.x5[7].floating.n4 vss -28.3f
C2415 x2.x1.x5[7].floating.n5 vss 52.7f
C2416 x2.x1.x5[7].floating.n6 vss -28.3f
C2417 x2.x1.x5[7].floating.n7 vss -7.07f
C2418 x2.x1.x5[7].floating.n8 vss 3.83f
C2419 x2.x1.x5[7].floating.n9 vss -28.9f
C2420 x2.x1.x5[7].floating.n10 vss -8.01f
C2421 x2.x1.x5[7].floating.n11 vss 2.21f
C2422 x2.x1.x5[7].floating.t4 vss 0.859f
C2423 x2.x1.x5[7].floating.n12 vss 6.65f
C2424 x2.x1.x5[7].floating.n13 vss 1.21f
C2425 x2.x1.x5[7].floating.n14 vss 1.17f
C2426 x2.x1.x5[7].floating.n15 vss 2.18f
C2427 x2.x1.x5[7].floating.n16 vss 1.06f
C2428 x2.x1.x5[7].floating.n17 vss 0.366f
C2429 x2.x1.x5[7].floating.n18 vss 1.06f
C2430 x2.x1.x5[7].floating.n19 vss 2.8f
C2431 x2.x1.x5[7].floating.n20 vss 51.4f
C2432 x2.x1.x5[7].floating.n21 vss 2.79f
C2433 x2.x1.x5[7].floating.n22 vss 1.06f
C2434 x2.x1.x5[7].floating.n23 vss 0.364f
C2435 x2.x1.x5[7].floating.t5 vss 0.859f
C2436 x2.x1.x5[7].floating.n24 vss 6.48f
C2437 x2.x1.x5[7].floating.n25 vss 1.15f
C2438 x2.x1.x5[7].floating.n26 vss 1.36f
C2439 x2.x1.x5[7].floating.n27 vss 2.2f
C2440 x2.x1.x5[7].floating.n28 vss 1.06f
C2441 x2.x1.x5[7].floating.n29 vss 2.23f
C2442 x2.x1.x5[7].floating.n30 vss -7.99f
C2443 x2.x1.x5[7].floating.n31 vss -28.9f
C2444 x2.x1.x5[7].floating.n32 vss 3.83f
C2445 x2.x1.x5[7].floating.n33 vss -7.07f
C2446 x2.x1.x5[7].floating.n34 vss -28.3f
C2447 x2.x1.x5[7].floating.n35 vss 52.7f
C2448 x2.x1.x5[7].floating.n36 vss -28.3f
C2449 x2.x1.x5[7].floating.n37 vss -7.07f
C2450 x2.x1.x5[7].floating.n38 vss 3.83f
C2451 x2.x1.x5[7].floating.n39 vss -28.9f
C2452 x2.x1.x5[7].floating.n40 vss -8.01f
C2453 x2.x1.x5[7].floating.n41 vss 2.21f
C2454 x2.x1.x5[7].floating.t6 vss 0.859f
C2455 x2.x1.x5[7].floating.n42 vss 6.65f
C2456 x2.x1.x5[7].floating.n43 vss 1.21f
C2457 x2.x1.x5[7].floating.n44 vss 1.17f
C2458 x2.x1.x5[7].floating.n45 vss 2.18f
C2459 x2.x1.x5[7].floating.n46 vss 1.06f
C2460 x2.x1.x5[7].floating.n47 vss 0.366f
C2461 x2.x1.x5[7].floating.n48 vss 1.06f
C2462 x2.x1.x5[7].floating.n49 vss 2.8f
C2463 x2.x1.x5[7].floating.n50 vss 51.4f
C2464 x2.x1.x5[7].floating.n51 vss 2.79f
C2465 x2.x1.x5[7].floating.n52 vss 1.06f
C2466 x2.x1.x5[7].floating.n53 vss 0.364f
C2467 x2.x1.x5[7].floating.t7 vss 0.859f
C2468 x2.x1.x5[7].floating.n54 vss 6.48f
C2469 x2.x1.x5[7].floating.n55 vss 1.15f
C2470 x2.x1.x5[7].floating.n56 vss 1.36f
C2471 x2.x1.x5[7].floating.n57 vss 2.2f
C2472 x2.x1.x5[7].floating.n58 vss 1.06f
C2473 x2.x1.x5[7].floating.n59 vss 2.23f
C2474 x2.x1.x5[7].floating.n60 vss -7.99f
C2475 x2.x1.x5[7].floating.n61 vss -28.9f
C2476 x2.x1.x5[7].floating.n62 vss 3.83f
C2477 x2.x1.x5[7].floating.n63 vss -7.07f
C2478 x2.x1.x5[7].floating.n64 vss -28.3f
C2479 x2.x1.x5[7].floating.n65 vss 52.7f
C2480 x2.x1.x5[7].floating.n66 vss -28.3f
C2481 x2.x1.x5[7].floating.n67 vss -7.07f
C2482 x2.x1.x5[7].floating.n68 vss 3.83f
C2483 x2.x1.x5[7].floating.n69 vss -28.9f
C2484 x2.x1.x5[7].floating.n70 vss -8.01f
C2485 x2.x1.x5[7].floating.n71 vss 2.21f
C2486 x2.x1.x5[7].floating.t0 vss 0.859f
C2487 x2.x1.x5[7].floating.n72 vss 6.65f
C2488 x2.x1.x5[7].floating.n73 vss 1.21f
C2489 x2.x1.x5[7].floating.n74 vss 1.17f
C2490 x2.x1.x5[7].floating.n75 vss 2.18f
C2491 x2.x1.x5[7].floating.n76 vss 1.06f
C2492 x2.x1.x5[7].floating.n77 vss 0.366f
C2493 x2.x1.x5[7].floating.n78 vss 1.06f
C2494 x2.x1.x5[7].floating.n79 vss 2.8f
C2495 x2.x1.x5[7].floating.n80 vss 51.4f
C2496 x2.x1.x5[7].floating.n81 vss 2.79f
C2497 x2.x1.x5[7].floating.n82 vss 1.06f
C2498 x2.x1.x5[7].floating.n83 vss 0.364f
C2499 x2.x1.x5[7].floating.t2 vss 0.859f
C2500 x2.x1.x5[7].floating.n84 vss 6.48f
C2501 x2.x1.x5[7].floating.n85 vss 1.15f
C2502 x2.x1.x5[7].floating.n86 vss 1.36f
C2503 x2.x1.x5[7].floating.n87 vss 2.2f
C2504 x2.x1.x5[7].floating.n88 vss 1.06f
C2505 x2.x1.x5[7].floating.n89 vss -15.2f
C2506 x2.x1.x5[7].floating.n90 vss -15.2f
C2507 x2.x1.x5[7].floating.n91 vss -41.6f
C2508 x2.x1.x5[7].floating.n92 vss 0.766f
C2509 x2.x1.x5[7].floating.n93 vss 2.47f
C2510 x2.x1.x5[7].floating.n94 vss 51.5f
C2511 x2.x1.x5[7].floating.n95 vss 2.47f
C2512 x2.x1.x5[7].floating.n96 vss 0.766f
C2513 x2.x1.x5[7].floating.n97 vss -33.5f
C2514 x2.x1.x5[7].floating.n98 vss -4.56f
C2515 x2.x1.x5[7].floating.n99 vss 3.83f
C2516 x2.x1.x5[7].floating.n100 vss -28.9f
C2517 x2.x1.x5[7].floating.n101 vss -7.07f
C2518 x2.x1.x5[7].floating.n102 vss 2.68f
C2519 x2.x1.x5[7].floating.n103 vss 52f
C2520 x2.x1.x5[7].floating.n104 vss 3.23f
C2521 x2.x1.x5[7].floating.n105 vss -7.84f
C2522 x2.x1.x5[7].floating.n106 vss -28.9f
C2523 x2.x1.x5[7].floating.n107 vss 3.83f
C2524 x2.x1.x5[7].floating.n108 vss -5.01f
C2525 x2.x1.x5[7].floating.n109 vss -33f
C2526 x2.x1.x5[7].floating.n110 vss 0.766f
C2527 x2.x1.x5[7].floating.n111 vss 2.47f
C2528 x2.x1.x5[7].floating.n112 vss 51.5f
C2529 x2.x1.x5[7].floating.n113 vss 2.47f
C2530 x2.x1.x5[7].floating.n114 vss 0.766f
C2531 x2.x1.x5[7].floating.n115 vss -33.5f
C2532 x2.x1.x5[7].floating.n116 vss -4.56f
C2533 x2.x1.x5[7].floating.n117 vss 3.83f
C2534 x2.x1.x5[7].floating.n118 vss -28.9f
C2535 x2.x1.x5[7].floating.n119 vss -7.07f
C2536 x2.x1.x5[7].floating.n120 vss 2.68f
C2537 x2.x1.x5[7].floating.n121 vss 52f
C2538 x2.x1.x5[7].floating.n122 vss 3.23f
C2539 x2.x1.x5[7].floating.n123 vss -7.84f
C2540 x2.x1.x5[7].floating.n124 vss -28.9f
C2541 x2.x1.x5[7].floating.n125 vss 3.83f
C2542 x2.x1.x5[7].floating.n126 vss -5.01f
C2543 x2.x1.x5[7].floating.n127 vss -33f
C2544 x2.x1.x5[7].floating.n128 vss 0.766f
C2545 x2.x1.x5[7].floating.n129 vss 2.47f
C2546 x2.x1.x5[7].floating.n130 vss 51.5f
C2547 x2.x1.x5[7].floating.n131 vss 2.47f
C2548 x2.x1.x5[7].floating.n132 vss 0.766f
C2549 x2.x1.x5[7].floating.n133 vss -33.5f
C2550 x2.x1.x5[7].floating.n134 vss -4.56f
C2551 x2.x1.x5[7].floating.n135 vss 3.83f
C2552 x2.x1.x5[7].floating.n136 vss -28.9f
C2553 x2.x1.x5[7].floating.n137 vss -7.07f
C2554 x2.x1.x5[7].floating.n138 vss 2.68f
C2555 x2.x1.x5[7].floating.n139 vss 52f
C2556 x2.x1.x5[7].floating.n140 vss 3.23f
C2557 x2.x1.x5[7].floating.n141 vss 2.23f
C2558 x2.x1.x5[7].floating.t3 vss 0.859f
C2559 x2.x1.x5[7].floating.n142 vss 6.48f
C2560 x2.x1.x5[7].floating.n143 vss 1.15f
C2561 x2.x1.x5[7].floating.n144 vss 1.36f
C2562 x2.x1.x5[7].floating.n145 vss 2.2f
C2563 x2.x1.x5[7].floating.n146 vss 1.06f
C2564 x2.x1.x5[7].floating.n147 vss 0.364f
C2565 x2.x1.x5[7].floating.n148 vss 1.06f
C2566 x2.x1.x5[7].floating.n149 vss 2.79f
C2567 x2.x1.x5[7].floating.n150 vss 51.4f
C2568 x2.x1.x5[7].floating.n151 vss 2.8f
C2569 x2.x1.x5[7].floating.n152 vss 1.06f
C2570 x2.x1.x5[7].floating.n153 vss 0.366f
C2571 x2.x1.x5[7].floating.t1 vss 0.859f
C2572 x2.x1.x5[7].floating.n154 vss 7.16f
C2573 x2.x1.x5[7].floating.n155 vss 1.21f
C2574 x2.x1.x5[7].floating.n156 vss 1.17f
C2575 x2.x1.x5[7].floating.n157 vss 1.67f
C2576 x2.x1.x5[7].floating.n158 vss 1.06f
C2577 x2.x1.x5[7].floating.n159 vss -17.4f
C2578 x2.x1.x5[7].floating.n160 vss -17.2f
C2579 x2.x1.x5[7].floating.n161 vss -43.6f
C2580 x2.x1.x5[7].floating.n162 vss 0.766f
C2581 x2.x1.x5[7].floating.n163 vss 2.47f
C2582 x2.x1.x5[7].floating.n164 vss 51.5f
C2583 x2.x1.x5[7].floating.n165 vss 2.47f
C2584 x2.x1.x5[7].floating.n166 vss 0.766f
C2585 x2.x1.x5[7].floating.n167 vss -33f
C2586 x2.x1.x5[7].floating.n168 vss -5.01f
C2587 x2.x1.x5[7].floating.n169 vss 3.83f
C2588 x2.x1.x5[7].floating.n170 vss -28.9f
C2589 x2.x1.x5[7].floating.n171 vss -7.84f
C2590 x2.x1.x10.Y.t1 vss 0.0462f
C2591 x2.x1.x10.Y.t7 vss 0.0167f
C2592 x2.x1.x10.Y.t9 vss 0.0167f
C2593 x2.x1.x10.Y.t2 vss 0.0167f
C2594 x2.x1.x10.Y.t3 vss 0.0167f
C2595 x2.x1.x10.Y.t4 vss 0.0167f
C2596 x2.x1.x10.Y.t5 vss 0.0167f
C2597 x2.x1.x10.Y.t6 vss 0.0167f
C2598 x2.x1.x10.Y.t8 vss 0.0167f
C2599 x2.x1.x10.Y.n0 vss 0.222f
C2600 x2.x1.x10.Y.n1 vss 0.0366f
C2601 x2.x1.x10.Y.t0 vss 0.0174f
C2602 x2.x1.x10.Y.n2 vss 0.0188f
C2603 x2.x1.x10.Y.n3 vss 0.0186f
C2604 x2.x1.x10.Y.n4 vss 0.0151f
C2605 x2.x1.x10.Y.n5 vss 0.0211f
C2606 vdd.n0 vss 0.00885f
C2607 vdd.n1 vss 0.0158f
C2608 vdd.n2 vss 0.00433f
C2609 vdd.n3 vss 0.00246f
C2610 vdd.n4 vss 0.0163f
C2611 vdd.n5 vss 0.00885f
C2612 vdd.n6 vss 0.0345f
C2613 vdd.t96 vss 0.12f
C2614 vdd.t84 vss 0.0416f
C2615 vdd.n7 vss 0.0594f
C2616 vdd.n8 vss 0.0116f
C2617 vdd.n9 vss 0.0335f
C2618 vdd.n10 vss 0.021f
C2619 vdd.n11 vss 0.0221f
C2620 vdd.t67 vss 0.114f
C2621 vdd.t83 vss 0.0585f
C2622 vdd.n12 vss 0.0559f
C2623 vdd.n13 vss 0.0217f
C2624 vdd.n14 vss 0.0234f
C2625 vdd.t97 vss 0.00676f
C2626 vdd.t68 vss 0.00676f
C2627 vdd.n15 vss 0.0143f
C2628 vdd.n16 vss 0.0375f
C2629 vdd.n17 vss 7.62e-19
C2630 vdd.n18 vss 0.0634f
C2631 vdd.n19 vss 0.0462f
C2632 vdd.n20 vss 0.00885f
C2633 vdd.n21 vss 0.0158f
C2634 vdd.n22 vss 0.116f
C2635 vdd.n23 vss 0.0348f
C2636 vdd.t59 vss -0.00303f
C2637 vdd.t18 vss 0.00951f
C2638 vdd.n24 vss 0.0438f
C2639 vdd.n25 vss 0.0539f
C2640 vdd.t58 vss 0.15f
C2641 vdd.n26 vss 0.0754f
C2642 vdd.n27 vss 0.0216f
C2643 vdd.n28 vss 0.0184f
C2644 vdd.n29 vss 0.0682f
C2645 vdd.t17 vss 0.073f
C2646 vdd.n30 vss 0.106f
C2647 vdd.n31 vss 0.0216f
C2648 vdd.n32 vss 0.0349f
C2649 vdd.n33 vss 0.0345f
C2650 vdd.n34 vss 0.121f
C2651 vdd.n35 vss 0.0216f
C2652 vdd.n36 vss 0.0338f
C2653 vdd.n37 vss 0.0345f
C2654 vdd.t14 vss -0.00568f
C2655 vdd.t8 vss 0.0103f
C2656 vdd.n38 vss 0.0402f
C2657 vdd.n39 vss 0.0344f
C2658 vdd.t13 vss 0.123f
C2659 vdd.n40 vss 0.126f
C2660 vdd.n41 vss 0.0216f
C2661 vdd.n42 vss 0.0285f
C2662 vdd.n43 vss 0.0345f
C2663 vdd.t7 vss 0.12f
C2664 vdd.n44 vss 0.161f
C2665 vdd.n45 vss 0.0216f
C2666 vdd.n46 vss 0.0605f
C2667 vdd.n47 vss 0.0257f
C2668 vdd.n48 vss 0.372f
C2669 vdd.t114 vss 0.0294f
C2670 vdd.n49 vss 0.0364f
C2671 vdd.n50 vss 0.216f
C2672 vdd.n51 vss 0.0216f
C2673 vdd.n52 vss 0.0419f
C2674 vdd.n53 vss 0.045f
C2675 vdd.t105 vss 0.0243f
C2676 vdd.t116 vss 0.0108f
C2677 vdd.n54 vss 0.0378f
C2678 vdd.n55 vss 0.052f
C2679 vdd.t115 vss 0.116f
C2680 vdd.n56 vss 0.126f
C2681 vdd.n57 vss 0.0216f
C2682 vdd.n58 vss 0.0256f
C2683 vdd.n59 vss 0.048f
C2684 vdd.t104 vss 0.12f
C2685 vdd.n60 vss 0.172f
C2686 vdd.n61 vss 0.0216f
C2687 vdd.n62 vss 0.0267f
C2688 vdd.n63 vss 0.0619f
C2689 vdd.n64 vss 0.00885f
C2690 vdd.n65 vss 0.0158f
C2691 vdd.n66 vss 0.00433f
C2692 vdd.n67 vss 0.00246f
C2693 vdd.n68 vss 0.0163f
C2694 vdd.n69 vss 0.00885f
C2695 vdd.n70 vss 0.0345f
C2696 vdd.n71 vss 0.187f
C2697 vdd.n72 vss 0.0216f
C2698 vdd.n73 vss 0.0349f
C2699 vdd.n74 vss 0.0417f
C2700 vdd.t95 vss 0.229f
C2701 vdd.n75 vss 0.0216f
C2702 vdd.n76 vss 0.0349f
C2703 vdd.n77 vss 0.0627f
C2704 vdd.n78 vss 0.00885f
C2705 vdd.n79 vss 0.0158f
C2706 vdd.n80 vss 0.00433f
C2707 vdd.n81 vss 0.00246f
C2708 vdd.n82 vss 0.0163f
C2709 vdd.n83 vss 0.00885f
C2710 vdd.n84 vss 0.0345f
C2711 vdd.t69 vss 0.12f
C2712 vdd.n85 vss 0.13f
C2713 vdd.n86 vss 0.0216f
C2714 vdd.n87 vss 0.0349f
C2715 vdd.n88 vss 0.0409f
C2716 vdd.t15 vss 0.12f
C2717 vdd.n89 vss 0.143f
C2718 vdd.n90 vss 0.0216f
C2719 vdd.n91 vss 0.032f
C2720 vdd.n92 vss 0.0653f
C2721 vdd.n93 vss 0.00885f
C2722 vdd.n94 vss 0.0158f
C2723 vdd.n95 vss 0.00433f
C2724 vdd.n96 vss 0.00246f
C2725 vdd.n97 vss 0.0163f
C2726 vdd.n98 vss 0.00885f
C2727 vdd.n99 vss 0.0345f
C2728 vdd.t34 vss 0.0064f
C2729 vdd.t16 vss 0.0064f
C2730 vdd.n100 vss 0.0133f
C2731 vdd.n101 vss 0.0396f
C2732 vdd.t33 vss 0.12f
C2733 vdd.n102 vss 0.14f
C2734 vdd.n103 vss 0.0216f
C2735 vdd.n104 vss 0.0203f
C2736 vdd.n105 vss 0.0383f
C2737 vdd.t73 vss 0.12f
C2738 vdd.n106 vss 0.125f
C2739 vdd.n107 vss 0.0216f
C2740 vdd.n108 vss 0.0349f
C2741 vdd.n109 vss 0.0691f
C2742 vdd.t113 vss 0.12f
C2743 vdd.n110 vss 0.0936f
C2744 vdd.n111 vss 0.0216f
C2745 vdd.n112 vss 0.0292f
C2746 vdd.n113 vss 0.0417f
C2747 vdd.n114 vss 0.121f
C2748 vdd.n115 vss 1.24f
C2749 vdd.n116 vss 0.0289f
C2750 vdd.n117 vss 0.0298f
C2751 vdd.n118 vss 0.155f
C2752 vdd.n119 vss 0.154f
C2753 vdd.n120 vss 0.0289f
C2754 vdd.n121 vss 0.0298f
C2755 vdd.n122 vss 0.15f
C2756 vdd.n123 vss 0.149f
C2757 vdd.n124 vss 0.0289f
C2758 vdd.n125 vss 0.0298f
C2759 vdd.n126 vss 0.165f
C2760 vdd.n127 vss 0.164f
C2761 vdd.n128 vss 0.0158f
C2762 vdd.n129 vss 0.00885f
C2763 vdd.t35 vss 0.12f
C2764 vdd.n130 vss 0.136f
C2765 vdd.n131 vss 0.0216f
C2766 vdd.n132 vss 0.0292f
C2767 vdd.n133 vss 0.0691f
C2768 vdd.t49 vss 0.113f
C2769 vdd.n134 vss 0.123f
C2770 vdd.n135 vss 0.0216f
C2771 vdd.n136 vss 0.0349f
C2772 vdd.n137 vss 0.0555f
C2773 vdd.n138 vss 0.0345f
C2774 vdd.n139 vss 0.00885f
C2775 vdd.n140 vss 0.0163f
C2776 vdd.n141 vss 0.00246f
C2777 vdd.n142 vss 0.00433f
C2778 vdd.n143 vss 0.0289f
C2779 vdd.n144 vss 0.0298f
C2780 vdd.n145 vss 0.388f
C2781 vdd.n146 vss 0.387f
C2782 vdd.n147 vss 0.0158f
C2783 vdd.n148 vss 0.00885f
C2784 vdd.t36 vss 0.0064f
C2785 vdd.t107 vss 0.00608f
C2786 vdd.n149 vss 0.0131f
C2787 vdd.n150 vss 0.0424f
C2788 vdd.t106 vss 0.12f
C2789 vdd.n151 vss 0.138f
C2790 vdd.n152 vss 0.0216f
C2791 vdd.n153 vss 0.0231f
C2792 vdd.n154 vss 0.0691f
C2793 vdd.n155 vss 0.156f
C2794 vdd.n156 vss 0.0215f
C2795 vdd.n157 vss 0.0347f
C2796 vdd.n158 vss 0.0691f
C2797 vdd.t98 vss 0.118f
C2798 vdd.n159 vss 0.109f
C2799 vdd.n160 vss 0.0213f
C2800 vdd.n161 vss 0.0233f
C2801 vdd.n162 vss 0.0231f
C2802 vdd.n163 vss 0.0379f
C2803 vdd.t6 vss 0.0156f
C2804 vdd.t129 vss 0.0416f
C2805 vdd.n164 vss 0.0599f
C2806 vdd.t5 vss 0.117f
C2807 vdd.n165 vss 0.0234f
C2808 vdd.n166 vss 0.0231f
C2809 vdd.n167 vss 0.0213f
C2810 vdd.n168 vss 0.165f
C2811 vdd.n169 vss 0.0793f
C2812 vdd.n170 vss 0.0217f
C2813 vdd.n171 vss 0.0231f
C2814 vdd.n172 vss 0.0401f
C2815 vdd.n173 vss 0.0409f
C2816 vdd.t70 vss 0.118f
C2817 vdd.t128 vss 0.065f
C2818 vdd.n174 vss 0.0624f
C2819 vdd.n175 vss 0.0218f
C2820 vdd.n176 vss 0.0234f
C2821 vdd.n177 vss 0.013f
C2822 vdd.n178 vss 0.0657f
C2823 vdd.n179 vss 0.0345f
C2824 vdd.n180 vss 0.00885f
C2825 vdd.n181 vss 0.0163f
C2826 vdd.n182 vss 0.00246f
C2827 vdd.n183 vss 0.00433f
C2828 vdd.n184 vss 0.0289f
C2829 vdd.n185 vss 0.0298f
C2830 vdd.n186 vss 0.198f
C2831 vdd.n187 vss 0.197f
C2832 vdd.n188 vss 0.116f
C2833 vdd.n189 vss 0.0101f
C2834 vdd.n190 vss 0.00569f
C2835 vdd.n191 vss 0.0175f
C2836 vdd.t43 vss 0.0416f
C2837 vdd.n192 vss 0.00808f
C2838 vdd.n193 vss 0.0102f
C2839 vdd.n194 vss 0.196f
C2840 vdd.n195 vss 0.0114f
C2841 vdd.n196 vss 0.00209f
C2842 vdd.n197 vss 0.00319f
C2843 vdd.n198 vss 0.00713f
C2844 vdd.n199 vss 0.00362f
C2845 vdd.n200 vss 0.0101f
C2846 vdd.n201 vss 0.0139f
C2847 vdd.n202 vss 0.0175f
C2848 vdd.n203 vss 0.0163f
C2849 vdd.n204 vss 0.0216f
C2850 vdd.n205 vss 0.0175f
C2851 vdd.n206 vss 0.00175f
C2852 vdd.n207 vss 0.0213f
C2853 vdd.n208 vss 0.00563f
C2854 vdd.n209 vss 0.00333f
C2855 vdd.n210 vss 0.015f
C2856 vdd.t66 vss 0.0416f
C2857 vdd.n211 vss 0.0458f
C2858 vdd.n212 vss 2.07f
C2859 vdd.n213 vss 1.03f
C2860 vdd.t78 vss 1.43f
C2861 vdd.t110 vss 0.228f
C2862 vdd.n214 vss 0.0102f
C2863 vdd.n215 vss 0.00808f
C2864 vdd.t111 vss 0.0416f
C2865 vdd.n216 vss 0.0175f
C2866 vdd.n217 vss 6.66e-19
C2867 vdd.n218 vss 0.0101f
C2868 vdd.n219 vss 0.0152f
C2869 vdd.n220 vss 0.0101f
C2870 vdd.n221 vss 0.00376f
C2871 vdd.n222 vss 0.00319f
C2872 vdd.n223 vss 0.00209f
C2873 vdd.n224 vss 0.00882f
C2874 vdd.n225 vss 0.00209f
C2875 vdd.n226 vss 0.0256f
C2876 vdd.n227 vss 0.00133f
C2877 vdd.n228 vss 0.116f
C2878 vdd.n229 vss 0.0664f
C2879 vdd.n230 vss 0.00673f
C2880 vdd.n231 vss 0.0163f
C2881 vdd.n232 vss 0.0163f
C2882 vdd.n233 vss 0.0427f
C2883 vdd.n234 vss 0.0313f
C2884 vdd.n235 vss 0.0163f
C2885 vdd.n236 vss 0.00673f
C2886 vdd.n237 vss 0.00518f
C2887 vdd.n238 vss 0.0495f
C2888 vdd.n239 vss 0.0213f
C2889 vdd.n240 vss 0.00362f
C2890 vdd.n241 vss 0.0223f
C2891 vdd.t118 vss 0.0416f
C2892 vdd.n242 vss 0.0224f
C2893 vdd.n243 vss 0.0226f
C2894 vdd.n244 vss 0.00908f
C2895 vdd.n245 vss 0.00994f
C2896 vdd.n246 vss 0.0129f
C2897 vdd.n247 vss 0.251f
C2898 vdd.n248 vss 0.00247f
C2899 vdd.n249 vss 0.00226f
C2900 vdd.n250 vss 2.1f
C2901 vdd.n251 vss 0.0105f
C2902 vdd.n253 vss 0.0105f
C2903 vdd.n257 vss 0.0105f
C2904 vdd.n260 vss 0.00226f
C2905 vdd.n261 vss 0.047f
C2906 vdd.n262 vss 0.008f
C2907 vdd.n263 vss 0.00219f
C2908 vdd.n264 vss 0.00226f
C2909 vdd.n265 vss 0.00219f
C2910 vdd.n266 vss 0.00219f
C2911 vdd.n267 vss 3.87e-19
C2912 vdd.n268 vss 0.00542f
C2913 vdd.n269 vss 0.00271f
C2914 vdd.n270 vss 0.00658f
C2915 vdd.n271 vss 0.00359f
C2916 vdd.n272 vss 0.00638f
C2917 vdd.n273 vss 0.0185f
C2918 vdd.n274 vss -0.173f
C2919 vdd.n275 vss 0.0113f
C2920 vdd.n276 vss 2.66e-19
C2921 vdd.n277 vss 0.0115f
C2922 vdd.n278 vss 0.00359f
C2923 vdd.n279 vss 0.00271f
C2924 vdd.n280 vss 0.00219f
C2925 vdd.n281 vss 3.87e-19
C2926 vdd.n282 vss 0.00219f
C2927 vdd.n283 vss 0.008f
C2928 vdd.n284 vss 0.00851f
C2929 vdd.n285 vss 0.00219f
C2930 vdd.n286 vss 0.00219f
C2931 vdd.n287 vss 3.87e-19
C2932 vdd.n288 vss 0.008f
C2933 vdd.n289 vss 0.00271f
C2934 vdd.n290 vss 0.00542f
C2935 vdd.n291 vss 0.00271f
C2936 vdd.n292 vss 0.00284f
C2937 vdd.n293 vss 0.00658f
C2938 vdd.n294 vss 0.00359f
C2939 vdd.n295 vss 0.00638f
C2940 vdd.n296 vss 0.0182f
C2941 vdd.n297 vss -0.173f
C2942 vdd.n298 vss 0.0111f
C2943 vdd.n299 vss 2.66e-19
C2944 vdd.n300 vss 3.87e-19
C2945 vdd.n301 vss 0.00477f
C2946 vdd.n302 vss 0.00284f
C2947 vdd.n303 vss 0.00219f
C2948 vdd.n304 vss 0.0105f
C2949 vdd.n305 vss 0.008f
C2950 vdd.n306 vss 0.00271f
C2951 vdd.n307 vss 0.00477f
C2952 vdd.n308 vss 0.00284f
C2953 vdd.n309 vss 3.87e-19
C2954 vdd.n310 vss 2.66e-19
C2955 vdd.n311 vss 0.00399f
C2956 vdd.n312 vss 0.0186f
C2957 vdd.n313 vss 0.00359f
C2958 vdd.n314 vss 0.00335f
C2959 vdd.n315 vss 0.00284f
C2960 vdd.n316 vss 0.00748f
C2961 vdd.n317 vss 0.00219f
C2962 vdd.n318 vss 0.008f
C2963 vdd.n319 vss 0.008f
C2964 vdd.n320 vss 0.00219f
C2965 vdd.n322 vss 0.00226f
C2966 vdd.n323 vss 0.00219f
C2967 vdd.n324 vss 0.0105f
C2968 vdd.n325 vss 0.00219f
C2969 vdd.n326 vss 0.00219f
C2970 vdd.n327 vss 0.00284f
C2971 vdd.n328 vss 0.00638f
C2972 vdd.n329 vss 0.0115f
C2973 vdd.n330 vss -0.0615f
C2974 vdd.n331 vss 0.00335f
C2975 vdd.n332 vss 0.00748f
C2976 vdd.n333 vss 0.00219f
C2977 vdd.n334 vss 0.00219f
C2978 vdd.n335 vss 0.00284f
C2979 vdd.n336 vss 0.0233f
C2980 vdd.n337 vss 0.0115f
C2981 vdd.n338 vss 2.66e-19
C2982 vdd.n339 vss 0.00271f
C2983 vdd.n340 vss 0.00284f
C2984 vdd.n341 vss 0.00748f
C2985 vdd.n342 vss 0.00219f
C2986 vdd.n343 vss 0.00219f
C2987 vdd.n344 vss 0.024f
C2988 vdd.n345 vss 0.00271f
C2989 vdd.n346 vss 0.0213f
C2990 vdd.n347 vss 0.0234f
C2991 vdd.n348 vss 0.0234f
C2992 vdd.n349 vss 0.0213f
C2993 vdd.n350 vss 0.00271f
C2994 vdd.n351 vss 0.024f
C2995 vdd.n352 vss 0.00219f
C2996 vdd.n353 vss 0.00851f
C2997 vdd.n354 vss 0.00219f
C2998 vdd.n355 vss 0.00219f
C2999 vdd.n356 vss 0.00284f
C3000 vdd.n357 vss 0.00335f
C3001 vdd.n358 vss 0.00306f
C3002 vdd.n359 vss 0.0115f
C3003 vdd.n360 vss 2.66e-19
C3004 vdd.n361 vss 0.00271f
C3005 vdd.n362 vss 0.00748f
C3006 vdd.n363 vss 0.008f
C3007 vdd.n364 vss 0.00226f
C3008 vdd.n365 vss 0.00219f
C3009 vdd.n366 vss 0.00219f
C3010 vdd.n367 vss 0.00748f
C3011 vdd.n368 vss 3.87e-19
C3012 vdd.n369 vss 0.008f
C3013 vdd.n370 vss 0.00271f
C3014 vdd.n371 vss 0.00335f
C3015 vdd.n372 vss 0.00306f
C3016 vdd.n373 vss -0.069f
C3017 vdd.n374 vss 0.00385f
C3018 vdd.n375 vss 0.0111f
C3019 vdd.n376 vss 0.00284f
C3020 vdd.n377 vss 0.00219f
C3021 vdd.n378 vss 0.00219f
C3022 vdd.n379 vss 2.58e-19
C3023 vdd.n380 vss 0.0105f
C3024 vdd.n381 vss 0.00219f
C3025 vdd.n382 vss 0.00219f
C3026 vdd.n383 vss 0.00748f
C3027 vdd.n384 vss 0.00284f
C3028 vdd.n385 vss 0.00335f
C3029 vdd.n386 vss 0.00306f
C3030 vdd.n387 vss 2.66e-19
C3031 vdd.n388 vss 0.0115f
C3032 vdd.n389 vss 2.66e-19
C3033 vdd.n390 vss 0.00271f
C3034 vdd.n391 vss 0.00748f
C3035 vdd.n392 vss 0.00219f
C3036 vdd.n393 vss 0.00851f
C3037 vdd.n394 vss 0.00219f
C3038 vdd.n395 vss 0.00219f
C3039 vdd.n396 vss 0.00284f
C3040 vdd.n397 vss 0.00335f
C3041 vdd.n398 vss 0.00306f
C3042 vdd.n399 vss -0.069f
C3043 vdd.n400 vss 2.66e-19
C3044 vdd.n401 vss 0.00271f
C3045 vdd.n402 vss 0.0241f
C3046 vdd.n403 vss 0.00219f
C3047 vdd.n404 vss 0.0105f
C3048 vdd.n405 vss 0.00219f
C3049 vdd.n406 vss 0.00219f
C3050 vdd.n407 vss 3.87e-19
C3051 vdd.n408 vss 0.00271f
C3052 vdd.n409 vss 0.00335f
C3053 vdd.n410 vss 0.0205f
C3054 vdd.n411 vss 0.00359f
C3055 vdd.n412 vss 0.0197f
C3056 vdd.n413 vss -0.148f
C3057 vdd.n414 vss 0.00399f
C3058 vdd.n415 vss 0.0111f
C3059 vdd.n416 vss 2.66e-19
C3060 vdd.n417 vss 3.87e-19
C3061 vdd.n418 vss 0.00477f
C3062 vdd.n419 vss 0.00284f
C3063 vdd.n420 vss 2.58e-19
C3064 vdd.n421 vss 0.00226f
C3065 vdd.n422 vss 0.00219f
C3066 vdd.n423 vss 0.00219f
C3067 vdd.n424 vss 0.00542f
C3068 vdd.n425 vss 0.00335f
C3069 vdd.n426 vss -0.0615f
C3070 vdd.n427 vss 0.00385f
C3071 vdd.n428 vss 0.00638f
C3072 vdd.n429 vss 0.0182f
C3073 vdd.n430 vss 0.00638f
C3074 vdd.n431 vss 0.00284f
C3075 vdd.n432 vss 0.00271f
C3076 vdd.n433 vss 0.00219f
C3077 vdd.n434 vss 0.00748f
C3078 vdd.n435 vss 0.00219f
C3079 vdd.n436 vss 0.008f
C3080 vdd.n437 vss 0.00851f
C3081 vdd.n438 vss 0.00219f
C3082 vdd.n439 vss 0.00219f
C3083 vdd.n440 vss 3.87e-19
C3084 vdd.n441 vss 0.008f
C3085 vdd.n442 vss 0.00271f
C3086 vdd.n443 vss 0.00542f
C3087 vdd.n444 vss 0.00271f
C3088 vdd.n445 vss 0.00658f
C3089 vdd.n446 vss 0.00359f
C3090 vdd.n447 vss -0.148f
C3091 vdd.n448 vss 0.00399f
C3092 vdd.n449 vss 0.0111f
C3093 vdd.n450 vss 2.66e-19
C3094 vdd.n451 vss 3.87e-19
C3095 vdd.n452 vss 0.00477f
C3096 vdd.n453 vss 0.00284f
C3097 vdd.n454 vss 0.00219f
C3098 vdd.n455 vss 0.0105f
C3099 vdd.n456 vss 0.008f
C3100 vdd.n457 vss 0.00271f
C3101 vdd.n458 vss 0.00477f
C3102 vdd.n459 vss 0.00284f
C3103 vdd.n460 vss 3.87e-19
C3104 vdd.n461 vss 2.66e-19
C3105 vdd.n462 vss -0.173f
C3106 vdd.n463 vss 0.0657f
C3107 vdd.n464 vss 2.66e-19
C3108 vdd.n465 vss 0.00271f
C3109 vdd.n466 vss 0.00284f
C3110 vdd.n467 vss 0.00748f
C3111 vdd.n468 vss 0.00219f
C3112 vdd.n469 vss 0.00219f
C3113 vdd.n470 vss 0.024f
C3114 vdd.n471 vss 0.0213f
C3115 vdd.n472 vss 0.00271f
C3116 vdd.n473 vss 0.008f
C3117 vdd.n474 vss 0.00219f
C3118 vdd.n476 vss 0.00226f
C3119 vdd.n477 vss 0.0193f
C3120 vdd.n478 vss 2.58e-19
C3121 vdd.n479 vss 0.00219f
C3122 vdd.n480 vss 0.00219f
C3123 vdd.n481 vss 0.00284f
C3124 vdd.n482 vss 0.0234f
C3125 vdd.n483 vss 0.0234f
C3126 vdd.n484 vss 0.0213f
C3127 vdd.n485 vss 0.00271f
C3128 vdd.n486 vss 0.024f
C3129 vdd.n487 vss 0.00219f
C3130 vdd.n488 vss 0.00851f
C3131 vdd.n489 vss 0.00219f
C3132 vdd.n490 vss 0.00219f
C3133 vdd.n491 vss 0.00284f
C3134 vdd.n492 vss 0.00335f
C3135 vdd.n493 vss 0.00306f
C3136 vdd.n494 vss 0.0115f
C3137 vdd.n495 vss 2.66e-19
C3138 vdd.n496 vss 0.00271f
C3139 vdd.n497 vss 0.00748f
C3140 vdd.n498 vss 0.008f
C3141 vdd.n499 vss 0.00226f
C3142 vdd.n500 vss 0.00219f
C3143 vdd.n501 vss 0.00219f
C3144 vdd.n502 vss 0.00748f
C3145 vdd.n503 vss 3.87e-19
C3146 vdd.n504 vss 0.008f
C3147 vdd.n505 vss 0.00271f
C3148 vdd.n506 vss 0.00335f
C3149 vdd.n507 vss 0.00306f
C3150 vdd.n508 vss -0.069f
C3151 vdd.n509 vss 0.00385f
C3152 vdd.n510 vss 0.0111f
C3153 vdd.n511 vss 0.00284f
C3154 vdd.n512 vss 0.00219f
C3155 vdd.n513 vss 0.00219f
C3156 vdd.n514 vss 2.58e-19
C3157 vdd.n515 vss 0.0105f
C3158 vdd.n516 vss 0.00219f
C3159 vdd.n517 vss 0.00219f
C3160 vdd.n518 vss 0.00748f
C3161 vdd.n519 vss 0.00284f
C3162 vdd.n520 vss 0.00335f
C3163 vdd.n521 vss 0.00306f
C3164 vdd.n522 vss 2.66e-19
C3165 vdd.n523 vss 0.0115f
C3166 vdd.n524 vss 2.66e-19
C3167 vdd.n525 vss 0.00271f
C3168 vdd.n526 vss 0.00748f
C3169 vdd.n527 vss 0.00219f
C3170 vdd.n528 vss 0.00851f
C3171 vdd.n529 vss 0.00219f
C3172 vdd.n530 vss 0.00219f
C3173 vdd.n531 vss 0.00284f
C3174 vdd.n532 vss 0.00335f
C3175 vdd.n533 vss 0.00306f
C3176 vdd.n534 vss -0.069f
C3177 vdd.n535 vss 2.66e-19
C3178 vdd.n536 vss 0.00271f
C3179 vdd.n537 vss 0.0241f
C3180 vdd.n538 vss 0.00219f
C3181 vdd.n539 vss 0.0105f
C3182 vdd.n540 vss 0.00219f
C3183 vdd.n541 vss 0.00219f
C3184 vdd.n542 vss 3.87e-19
C3185 vdd.n543 vss 0.00271f
C3186 vdd.n544 vss 0.00335f
C3187 vdd.n545 vss 0.0205f
C3188 vdd.n546 vss 0.00359f
C3189 vdd.n547 vss 0.0197f
C3190 vdd.n548 vss -0.148f
C3191 vdd.n549 vss 0.00399f
C3192 vdd.n550 vss 0.0111f
C3193 vdd.n551 vss 2.66e-19
C3194 vdd.n552 vss 3.87e-19
C3195 vdd.n553 vss 0.00477f
C3196 vdd.n554 vss 0.00284f
C3197 vdd.n555 vss 2.58e-19
C3198 vdd.n556 vss 0.00226f
C3199 vdd.n557 vss 0.00219f
C3200 vdd.n558 vss 0.00219f
C3201 vdd.n559 vss 0.00542f
C3202 vdd.n560 vss 0.00335f
C3203 vdd.n561 vss -0.0615f
C3204 vdd.n562 vss 0.00385f
C3205 vdd.n563 vss 0.00638f
C3206 vdd.n564 vss 0.0182f
C3207 vdd.n565 vss 0.00638f
C3208 vdd.n566 vss 0.00284f
C3209 vdd.n567 vss 0.00271f
C3210 vdd.n568 vss 0.00219f
C3211 vdd.n569 vss 0.00748f
C3212 vdd.n570 vss 0.00219f
C3213 vdd.n571 vss 0.008f
C3214 vdd.n572 vss 0.00851f
C3215 vdd.n573 vss 0.00219f
C3216 vdd.n574 vss 0.00219f
C3217 vdd.n575 vss 3.87e-19
C3218 vdd.n576 vss 0.008f
C3219 vdd.n577 vss 0.00271f
C3220 vdd.n578 vss 0.00542f
C3221 vdd.n579 vss 0.00271f
C3222 vdd.n580 vss 0.00658f
C3223 vdd.n581 vss 0.00359f
C3224 vdd.n582 vss -0.148f
C3225 vdd.n583 vss 0.00399f
C3226 vdd.n584 vss 0.0111f
C3227 vdd.n585 vss 2.66e-19
C3228 vdd.n586 vss 3.87e-19
C3229 vdd.n587 vss 0.00477f
C3230 vdd.n588 vss 0.00284f
C3231 vdd.n589 vss 0.00219f
C3232 vdd.n590 vss 0.0105f
C3233 vdd.n591 vss 0.008f
C3234 vdd.n592 vss 0.00271f
C3235 vdd.n593 vss 0.00477f
C3236 vdd.n594 vss 0.00284f
C3237 vdd.n595 vss 3.87e-19
C3238 vdd.n596 vss 2.66e-19
C3239 vdd.n597 vss -0.173f
C3240 vdd.n598 vss 0.0657f
C3241 vdd.n599 vss 2.66e-19
C3242 vdd.n600 vss 0.00271f
C3243 vdd.n601 vss 0.00284f
C3244 vdd.n602 vss 0.00748f
C3245 vdd.n603 vss 0.00219f
C3246 vdd.n604 vss 0.00219f
C3247 vdd.n605 vss 0.024f
C3248 vdd.n606 vss 0.0213f
C3249 vdd.n607 vss 0.00271f
C3250 vdd.n608 vss 0.008f
C3251 vdd.n609 vss 0.00219f
C3252 vdd.n611 vss 0.00226f
C3253 vdd.n612 vss 0.0193f
C3254 vdd.n613 vss 2.58e-19
C3255 vdd.n614 vss 0.00219f
C3256 vdd.n615 vss 0.00219f
C3257 vdd.n616 vss 0.00284f
C3258 vdd.n617 vss 0.0234f
C3259 vdd.n618 vss 0.0234f
C3260 vdd.n619 vss 0.0213f
C3261 vdd.n620 vss 0.00271f
C3262 vdd.n621 vss 0.024f
C3263 vdd.n622 vss 0.00219f
C3264 vdd.n623 vss 0.00851f
C3265 vdd.n624 vss 0.00219f
C3266 vdd.n625 vss 0.00219f
C3267 vdd.n626 vss 0.00284f
C3268 vdd.n627 vss 0.00335f
C3269 vdd.n628 vss 0.00306f
C3270 vdd.n629 vss 0.0115f
C3271 vdd.n630 vss 2.66e-19
C3272 vdd.n631 vss 0.00271f
C3273 vdd.n632 vss 0.00748f
C3274 vdd.n633 vss 0.008f
C3275 vdd.n634 vss 0.00226f
C3276 vdd.n635 vss 0.00219f
C3277 vdd.n636 vss 0.00219f
C3278 vdd.n637 vss 0.00748f
C3279 vdd.n638 vss 3.87e-19
C3280 vdd.n639 vss 0.008f
C3281 vdd.n640 vss 0.00271f
C3282 vdd.n641 vss 0.00335f
C3283 vdd.n642 vss 0.00306f
C3284 vdd.n643 vss -0.069f
C3285 vdd.n644 vss 0.00385f
C3286 vdd.n645 vss 0.0111f
C3287 vdd.n646 vss 0.00284f
C3288 vdd.n647 vss 0.00219f
C3289 vdd.n648 vss 0.00219f
C3290 vdd.n649 vss 2.58e-19
C3291 vdd.n650 vss 0.0105f
C3292 vdd.n651 vss 0.00219f
C3293 vdd.n652 vss 0.00219f
C3294 vdd.n653 vss 0.00748f
C3295 vdd.n654 vss 0.00284f
C3296 vdd.n655 vss 0.00335f
C3297 vdd.n656 vss 0.00306f
C3298 vdd.n657 vss 2.66e-19
C3299 vdd.n658 vss 0.0115f
C3300 vdd.n659 vss 2.66e-19
C3301 vdd.n660 vss 0.00271f
C3302 vdd.n661 vss 0.00748f
C3303 vdd.n662 vss 0.00219f
C3304 vdd.n663 vss 0.00851f
C3305 vdd.n664 vss 0.00219f
C3306 vdd.n665 vss 0.00219f
C3307 vdd.n666 vss 0.00284f
C3308 vdd.n667 vss 0.00335f
C3309 vdd.n668 vss 0.00306f
C3310 vdd.n669 vss -0.069f
C3311 vdd.n670 vss 2.66e-19
C3312 vdd.n671 vss 0.00271f
C3313 vdd.n672 vss 0.0241f
C3314 vdd.n673 vss 0.00219f
C3315 vdd.n674 vss 0.0105f
C3316 vdd.n675 vss 0.00219f
C3317 vdd.n676 vss 0.00219f
C3318 vdd.n677 vss 3.87e-19
C3319 vdd.n678 vss 0.00271f
C3320 vdd.n679 vss 0.00335f
C3321 vdd.n680 vss 0.0205f
C3322 vdd.n681 vss 0.00359f
C3323 vdd.n682 vss 0.0197f
C3324 vdd.n683 vss -0.148f
C3325 vdd.n684 vss 0.00399f
C3326 vdd.n685 vss 0.0111f
C3327 vdd.n686 vss 2.66e-19
C3328 vdd.n687 vss 3.87e-19
C3329 vdd.n688 vss 0.00477f
C3330 vdd.n689 vss 0.00284f
C3331 vdd.n690 vss 2.58e-19
C3332 vdd.n691 vss 0.00226f
C3333 vdd.n692 vss 0.00219f
C3334 vdd.n693 vss 0.00219f
C3335 vdd.n694 vss 0.00542f
C3336 vdd.n695 vss 0.00335f
C3337 vdd.n696 vss -0.0615f
C3338 vdd.n697 vss 0.00385f
C3339 vdd.n698 vss 0.00638f
C3340 vdd.n699 vss 0.0182f
C3341 vdd.n700 vss 0.00638f
C3342 vdd.n701 vss 0.00284f
C3343 vdd.n702 vss 0.00271f
C3344 vdd.n703 vss 0.00219f
C3345 vdd.n704 vss 0.00748f
C3346 vdd.n705 vss 0.00219f
C3347 vdd.n706 vss 0.008f
C3348 vdd.n707 vss 0.00851f
C3349 vdd.n708 vss 0.00219f
C3350 vdd.n709 vss 0.00219f
C3351 vdd.n710 vss 3.87e-19
C3352 vdd.n711 vss 0.008f
C3353 vdd.n712 vss 0.00271f
C3354 vdd.n713 vss 0.00542f
C3355 vdd.n714 vss 0.00271f
C3356 vdd.n715 vss 0.00658f
C3357 vdd.n716 vss 0.00359f
C3358 vdd.n717 vss -0.148f
C3359 vdd.n718 vss 0.00399f
C3360 vdd.n719 vss 0.0111f
C3361 vdd.n720 vss 2.66e-19
C3362 vdd.n721 vss 3.87e-19
C3363 vdd.n722 vss 0.00477f
C3364 vdd.n723 vss 0.00284f
C3365 vdd.n724 vss 0.00219f
C3366 vdd.n725 vss 0.0105f
C3367 vdd.n726 vss 0.008f
C3368 vdd.n727 vss 0.00271f
C3369 vdd.n728 vss 0.00477f
C3370 vdd.n729 vss 0.00284f
C3371 vdd.n730 vss 3.87e-19
C3372 vdd.n731 vss 2.66e-19
C3373 vdd.n732 vss -0.173f
C3374 vdd.n733 vss 0.0657f
C3375 vdd.n734 vss 2.66e-19
C3376 vdd.n735 vss 0.00271f
C3377 vdd.n736 vss 0.00284f
C3378 vdd.n737 vss 0.00748f
C3379 vdd.n738 vss 0.00219f
C3380 vdd.n739 vss 0.00219f
C3381 vdd.n740 vss 0.024f
C3382 vdd.n741 vss 0.0213f
C3383 vdd.n742 vss 0.00271f
C3384 vdd.n743 vss 0.008f
C3385 vdd.n744 vss 0.00219f
C3386 vdd.n746 vss 0.00226f
C3387 vdd.n747 vss 0.0193f
C3388 vdd.n748 vss 2.58e-19
C3389 vdd.n749 vss 0.00219f
C3390 vdd.n750 vss 0.00219f
C3391 vdd.n751 vss 0.00284f
C3392 vdd.n752 vss 0.0234f
C3393 vdd.n753 vss 0.0234f
C3394 vdd.n754 vss 0.0213f
C3395 vdd.n755 vss 0.00271f
C3396 vdd.n756 vss 0.024f
C3397 vdd.n757 vss 0.00219f
C3398 vdd.n758 vss 0.00851f
C3399 vdd.n759 vss 0.00219f
C3400 vdd.n760 vss 0.00219f
C3401 vdd.n761 vss 0.00284f
C3402 vdd.n762 vss 0.00335f
C3403 vdd.n763 vss 0.00306f
C3404 vdd.n764 vss 0.0115f
C3405 vdd.n765 vss 2.66e-19
C3406 vdd.n766 vss 0.00271f
C3407 vdd.n767 vss 0.00748f
C3408 vdd.n768 vss 0.008f
C3409 vdd.n769 vss 0.00226f
C3410 vdd.n770 vss 0.00219f
C3411 vdd.n771 vss 0.00219f
C3412 vdd.n772 vss 0.00748f
C3413 vdd.n773 vss 3.87e-19
C3414 vdd.n774 vss 0.008f
C3415 vdd.n775 vss 0.00271f
C3416 vdd.n776 vss 0.00335f
C3417 vdd.n777 vss 0.00306f
C3418 vdd.n778 vss -0.069f
C3419 vdd.n779 vss 0.00385f
C3420 vdd.n780 vss 0.0111f
C3421 vdd.n781 vss 0.00284f
C3422 vdd.n782 vss 0.00219f
C3423 vdd.n783 vss 0.00219f
C3424 vdd.n784 vss 2.58e-19
C3425 vdd.n785 vss 0.0105f
C3426 vdd.n786 vss 0.00219f
C3427 vdd.n787 vss 0.00219f
C3428 vdd.n788 vss 0.00748f
C3429 vdd.n789 vss 0.00284f
C3430 vdd.n790 vss 0.00335f
C3431 vdd.n791 vss 0.00306f
C3432 vdd.n792 vss 2.66e-19
C3433 vdd.n793 vss 0.0115f
C3434 vdd.n794 vss 2.66e-19
C3435 vdd.n795 vss 0.00271f
C3436 vdd.n796 vss 0.00748f
C3437 vdd.n797 vss 0.00219f
C3438 vdd.n798 vss 0.0226f
C3439 vdd.n799 vss 0.00219f
C3440 vdd.n800 vss 0.00219f
C3441 vdd.n801 vss 0.00284f
C3442 vdd.n802 vss 0.00335f
C3443 vdd.n803 vss 0.00306f
C3444 vdd.n804 vss -0.069f
C3445 vdd.n805 vss 2.66e-19
C3446 vdd.n806 vss 0.00271f
C3447 vdd.n807 vss 0.131f
C3448 vdd.n808 vss 0.00887f
C3449 vdd.n809 vss 0.0131f
C3450 vdd.n810 vss 0.00887f
C3451 vdd.n811 vss 0.00518f
C3452 vdd.t86 vss 0.206f
C3453 vdd.t85 vss 1.36f
C3454 vdd.n812 vss 0.385f
C3455 vdd.n813 vss 0.0131f
C3456 vdd.n814 vss 0.0131f
C3457 vdd.n815 vss 0.00887f
C3458 vdd.n816 vss 0.0163f
C3459 vdd.n817 vss 0.00518f
C3460 vdd.n818 vss 0.0635f
C3461 vdd.n819 vss 0.0547f
C3462 vdd.n820 vss 0.00673f
C3463 vdd.n821 vss 0.0163f
C3464 vdd.n822 vss 0.0163f
C3465 vdd.n823 vss 0.00887f
C3466 vdd.n824 vss 0.00518f
C3467 vdd.n825 vss 0.00668f
C3468 vdd.n826 vss 0.0664f
C3469 vdd.n827 vss 1.65f
C3470 vdd.t90 vss 1.84f
C3471 vdd.n828 vss 0.0157f
C3472 vdd.n829 vss 0.014f
C3473 vdd.n830 vss 0.00642f
C3474 vdd.n831 vss 0.0137f
C3475 vdd.n832 vss 0.00541f
C3476 vdd.t38 vss 0.00542f
C3477 vdd.t41 vss 0.00542f
C3478 vdd.n833 vss 0.0133f
C3479 vdd.n834 vss 0.0394f
C3480 vdd.n835 vss 0.00658f
C3481 vdd.n836 vss 0.0134f
C3482 vdd.n837 vss 0.0818f
C3483 vdd.n838 vss 0.0927f
C3484 vdd.n839 vss 0.00327f
C3485 vdd.n840 vss 0.0101f
C3486 vdd.n841 vss 0.013f
C3487 vdd.n842 vss 0.0189f
C3488 vdd.n843 vss 0.0158f
C3489 vdd.t121 vss 0.0416f
C3490 vdd.n844 vss 0.0454f
C3491 vdd.n845 vss 0.00651f
C3492 vdd.n846 vss 0.00209f
C3493 vdd.n847 vss 0.0166f
C3494 vdd.n848 vss 0.00133f
C3495 vdd.n849 vss 0.0517f
C3496 vdd.t120 vss 0.0847f
C3497 vdd.t126 vss 0.101f
C3498 vdd.n850 vss 0.0522f
C3499 vdd.n851 vss 0.043f
C3500 vdd.n852 vss 0.00226f
C3501 vdd.n853 vss 0.00219f
C3502 vdd.n854 vss 0.00284f
C3503 vdd.n855 vss 0.0105f
C3504 vdd.n856 vss 0.162f
C3505 vdd.n857 vss 0.00851f
C3506 vdd.n858 vss 0.008f
C3507 vdd.n859 vss 0.00219f
C3508 vdd.n860 vss 0.00748f
C3509 vdd.n861 vss 3.87e-19
C3510 vdd.n862 vss 0.00271f
C3511 vdd.n863 vss 0.00477f
C3512 vdd.n864 vss 0.00284f
C3513 vdd.n865 vss 3.87e-19
C3514 vdd.n866 vss -0.173f
C3515 vdd.n867 vss 2.66e-19
C3516 vdd.n868 vss 0.0191f
C3517 vdd.n869 vss 0.00359f
C3518 vdd.n870 vss -0.142f
C3519 vdd.n871 vss 0.00651f
C3520 vdd.n872 vss 0.00271f
C3521 vdd.n873 vss 0.00359f
C3522 vdd.n874 vss 0.00686f
C3523 vdd.n875 vss 0.00994f
C3524 vdd.t40 vss 0.00477f
C3525 vdd.n876 vss 0.0469f
C3526 vdd.n877 vss 0.00504f
C3527 vdd.n878 vss 0.0248f
C3528 vdd.n879 vss 0.0229f
C3529 vdd.n880 vss 0.00908f
C3530 vdd.n881 vss 8.67e-19
C3531 vdd.n882 vss 0.0142f
C3532 vdd.n883 vss 0.0295f
C3533 vdd.n884 vss 0.0129f
C3534 vdd.n885 vss 0.00335f
C3535 vdd.n886 vss 0.00637f
C3536 vdd.n887 vss 0.00385f
C3537 vdd.n888 vss 0.0062f
C3538 vdd.n889 vss 0.0118f
C3539 vdd.n890 vss 0.0114f
C3540 vdd.n891 vss -0.0687f
C3541 vdd.n892 vss 2.66e-19
C3542 vdd.n893 vss 0.00399f
C3543 vdd.n894 vss 3.87e-19
C3544 vdd.n895 vss 0.00284f
C3545 vdd.n896 vss 0.00219f
C3546 vdd.n897 vss 0.008f
C3547 vdd.n898 vss 0.00271f
C3548 vdd.n899 vss 0.00542f
C3549 vdd.n900 vss 0.00658f
C3550 vdd.n901 vss 0.00271f
C3551 vdd.n902 vss 0.00335f
C3552 vdd.n903 vss 0.00477f
C3553 vdd.n904 vss 0.00385f
C3554 vdd.n905 vss 0.00306f
C3555 vdd.n906 vss 0.0187f
C3556 vdd.n907 vss 0.0114f
C3557 vdd.n908 vss 0.0118f
C3558 vdd.n909 vss 2.66e-19
C3559 vdd.n910 vss 0.00399f
C3560 vdd.n911 vss 0.00651f
C3561 vdd.n912 vss 0.00306f
C3562 vdd.n913 vss 0.0187f
C3563 vdd.n914 vss 0.0187f
C3564 vdd.n915 vss 0.00399f
C3565 vdd.n916 vss 0.00359f
C3566 vdd.n917 vss 0.00658f
C3567 vdd.n918 vss 0.00271f
C3568 vdd.n919 vss 0.00542f
C3569 vdd.n920 vss 3.87e-19
C3570 vdd.n921 vss 0.00219f
C3571 vdd.n922 vss 0.00219f
C3572 vdd.n923 vss 0.00219f
C3573 vdd.n924 vss 0.00226f
C3574 vdd.n925 vss 0.0105f
C3575 vdd.n926 vss 0.162f
C3576 vdd.n927 vss 0.00851f
C3577 vdd.n928 vss 0.008f
C3578 vdd.n929 vss 0.008f
C3579 vdd.n930 vss 0.0105f
C3580 vdd.n931 vss 0.2f
C3581 vdd.n932 vss 0.043f
C3582 vdd.n933 vss 0.00226f
C3583 vdd.n934 vss 0.00219f
C3584 vdd.n935 vss 2.58e-19
C3585 vdd.n936 vss 0.00219f
C3586 vdd.n937 vss 0.00284f
C3587 vdd.n938 vss 0.00219f
C3588 vdd.n939 vss 0.00271f
C3589 vdd.n940 vss 0.008f
C3590 vdd.n941 vss 0.008f
C3591 vdd.n942 vss 0.0105f
C3592 vdd.n943 vss 0.2f
C3593 vdd.n944 vss 0.043f
C3594 vdd.n945 vss 0.162f
C3595 vdd.n946 vss 0.00851f
C3596 vdd.n947 vss 0.008f
C3597 vdd.n948 vss 0.00219f
C3598 vdd.n949 vss 0.00748f
C3599 vdd.n950 vss 3.87e-19
C3600 vdd.n951 vss 0.00271f
C3601 vdd.n952 vss 0.00477f
C3602 vdd.n953 vss 0.0471f
C3603 vdd.n954 vss 0.0354f
C3604 vdd.n955 vss -0.173f
C3605 vdd.n956 vss 2.66e-19
C3606 vdd.n957 vss 0.0191f
C3607 vdd.n958 vss 0.00359f
C3608 vdd.n959 vss -0.142f
C3609 vdd.n960 vss 0.0114f
C3610 vdd.n961 vss -0.0687f
C3611 vdd.n962 vss 2.66e-19
C3612 vdd.n963 vss 0.00399f
C3613 vdd.n964 vss 0.00651f
C3614 vdd.n965 vss 0.00284f
C3615 vdd.n966 vss 0.008f
C3616 vdd.n967 vss 0.00271f
C3617 vdd.n968 vss 0.00542f
C3618 vdd.n969 vss 0.00658f
C3619 vdd.n970 vss 0.00271f
C3620 vdd.n971 vss 0.00335f
C3621 vdd.n972 vss 0.00477f
C3622 vdd.n973 vss 0.00385f
C3623 vdd.n974 vss 0.00306f
C3624 vdd.n975 vss 0.0187f
C3625 vdd.n976 vss 0.0114f
C3626 vdd.n977 vss 0.0118f
C3627 vdd.n978 vss 2.66e-19
C3628 vdd.n979 vss 0.00399f
C3629 vdd.n980 vss 0.00651f
C3630 vdd.n981 vss 0.00306f
C3631 vdd.n982 vss 0.0187f
C3632 vdd.n983 vss 0.0113f
C3633 vdd.n984 vss 0.00359f
C3634 vdd.n985 vss 0.00271f
C3635 vdd.n986 vss 3.87e-19
C3636 vdd.n987 vss 0.00219f
C3637 vdd.n988 vss 0.0147f
C3638 vdd.n989 vss 0.00219f
C3639 vdd.n990 vss 0.00226f
C3640 vdd.n991 vss 0.0105f
C3641 vdd.n992 vss 0.043f
C3642 vdd.n993 vss 0.00226f
C3643 vdd.n994 vss 0.008f
C3644 vdd.n995 vss 0.2f
C3645 vdd.n996 vss 0.0105f
C3646 vdd.n997 vss 0.008f
C3647 vdd.n998 vss 0.00219f
C3648 vdd.n999 vss 0.0257f
C3649 vdd.n1000 vss 0.0193f
C3650 vdd.n1001 vss 0.101f
C3651 vdd.t103 vss 0.4f
C3652 vdd.n1002 vss 0.494f
C3653 vdd.n1003 vss 0.043f
C3654 vdd.n1004 vss 0.162f
C3655 vdd.n1005 vss 0.00851f
C3656 vdd.n1006 vss 0.008f
C3657 vdd.n1007 vss 0.00219f
C3658 vdd.n1008 vss 0.00748f
C3659 vdd.n1009 vss 3.87e-19
C3660 vdd.n1010 vss 0.00271f
C3661 vdd.n1011 vss 0.00477f
C3662 vdd.n1012 vss 0.00284f
C3663 vdd.n1013 vss 3.87e-19
C3664 vdd.n1014 vss -0.173f
C3665 vdd.n1015 vss 2.66e-19
C3666 vdd.n1016 vss 0.0188f
C3667 vdd.n1017 vss 0.00359f
C3668 vdd.n1018 vss -0.142f
C3669 vdd.n1019 vss -0.0689f
C3670 vdd.n1020 vss 2.66e-19
C3671 vdd.n1021 vss 0.00399f
C3672 vdd.n1022 vss 0.00651f
C3673 vdd.n1023 vss 0.00284f
C3674 vdd.n1024 vss 0.008f
C3675 vdd.n1025 vss 0.00271f
C3676 vdd.n1026 vss 0.00542f
C3677 vdd.n1027 vss 0.00658f
C3678 vdd.n1028 vss 0.00271f
C3679 vdd.n1029 vss 0.00335f
C3680 vdd.n1030 vss 0.00477f
C3681 vdd.n1031 vss 0.00385f
C3682 vdd.n1032 vss 0.00306f
C3683 vdd.n1033 vss 0.0184f
C3684 vdd.n1034 vss 0.0113f
C3685 vdd.n1035 vss 0.0116f
C3686 vdd.n1036 vss 2.66e-19
C3687 vdd.n1037 vss 0.00399f
C3688 vdd.n1038 vss 0.00651f
C3689 vdd.n1039 vss 0.00306f
C3690 vdd.n1040 vss 0.0184f
C3691 vdd.n1041 vss 0.0184f
C3692 vdd.n1042 vss 0.00399f
C3693 vdd.n1043 vss 0.00359f
C3694 vdd.n1044 vss 0.00658f
C3695 vdd.n1045 vss 0.00271f
C3696 vdd.n1046 vss 0.00542f
C3697 vdd.n1047 vss 3.87e-19
C3698 vdd.n1048 vss 0.00219f
C3699 vdd.n1049 vss 0.00219f
C3700 vdd.n1050 vss 0.00219f
C3701 vdd.n1051 vss 0.00226f
C3702 vdd.n1052 vss 0.0105f
C3703 vdd.n1053 vss 0.162f
C3704 vdd.n1054 vss 0.00851f
C3705 vdd.n1055 vss 0.008f
C3706 vdd.n1056 vss 0.008f
C3707 vdd.n1057 vss 0.0105f
C3708 vdd.n1058 vss 0.2f
C3709 vdd.n1059 vss 0.043f
C3710 vdd.n1060 vss 0.00226f
C3711 vdd.n1061 vss 0.00219f
C3712 vdd.n1062 vss 2.58e-19
C3713 vdd.n1063 vss 0.00219f
C3714 vdd.n1064 vss 0.00284f
C3715 vdd.n1065 vss 0.00219f
C3716 vdd.n1066 vss 0.00271f
C3717 vdd.n1067 vss 0.008f
C3718 vdd.n1068 vss 0.008f
C3719 vdd.n1069 vss 0.0105f
C3720 vdd.n1070 vss 0.2f
C3721 vdd.n1071 vss 0.043f
C3722 vdd.n1072 vss 0.162f
C3723 vdd.n1073 vss 0.00851f
C3724 vdd.n1074 vss 0.008f
C3725 vdd.n1075 vss 0.00219f
C3726 vdd.n1076 vss 0.00748f
C3727 vdd.n1077 vss 3.87e-19
C3728 vdd.n1078 vss 0.00271f
C3729 vdd.n1079 vss 0.00477f
C3730 vdd.n1080 vss 0.00284f
C3731 vdd.n1081 vss 3.87e-19
C3732 vdd.n1082 vss -0.173f
C3733 vdd.n1083 vss 2.66e-19
C3734 vdd.n1084 vss 0.0188f
C3735 vdd.n1085 vss 0.00359f
C3736 vdd.n1086 vss -0.142f
C3737 vdd.n1087 vss 0.0113f
C3738 vdd.n1088 vss -0.0689f
C3739 vdd.n1089 vss 2.66e-19
C3740 vdd.n1090 vss 0.00399f
C3741 vdd.n1091 vss 0.00651f
C3742 vdd.n1092 vss 0.00284f
C3743 vdd.n1093 vss 0.008f
C3744 vdd.n1094 vss 0.00271f
C3745 vdd.n1095 vss 0.00542f
C3746 vdd.n1096 vss 0.00658f
C3747 vdd.n1097 vss 0.00271f
C3748 vdd.n1098 vss 0.00335f
C3749 vdd.n1099 vss 0.00477f
C3750 vdd.n1100 vss 0.00385f
C3751 vdd.n1101 vss 0.00306f
C3752 vdd.n1102 vss 0.0184f
C3753 vdd.n1103 vss 0.0113f
C3754 vdd.n1104 vss 0.0116f
C3755 vdd.n1105 vss 2.66e-19
C3756 vdd.n1106 vss 0.00399f
C3757 vdd.n1107 vss 0.00651f
C3758 vdd.n1108 vss 0.00306f
C3759 vdd.n1109 vss 0.0184f
C3760 vdd.n1110 vss 0.0661f
C3761 vdd.n1111 vss 0.00399f
C3762 vdd.n1112 vss 2.66e-19
C3763 vdd.n1113 vss 0.00284f
C3764 vdd.n1114 vss 0.00271f
C3765 vdd.n1115 vss 0.00219f
C3766 vdd.n1116 vss 0.00748f
C3767 vdd.n1117 vss 0.00219f
C3768 vdd.n1118 vss 0.00219f
C3769 vdd.n1119 vss 0.00226f
C3770 vdd.n1120 vss 0.043f
C3771 vdd.n1121 vss 0.00226f
C3772 vdd.n1122 vss 0.008f
C3773 vdd.n1123 vss 0.2f
C3774 vdd.n1124 vss 0.0105f
C3775 vdd.n1125 vss 0.008f
C3776 vdd.n1126 vss 0.00219f
C3777 vdd.n1127 vss 0.024f
C3778 vdd.n1128 vss 0.00271f
C3779 vdd.n1129 vss 0.0234f
C3780 vdd.n1130 vss 0.024f
C3781 vdd.n1131 vss 0.00271f
C3782 vdd.n1132 vss 0.0213f
C3783 vdd.n1133 vss 0.0213f
C3784 vdd.n1134 vss 0.0234f
C3785 vdd.n1135 vss 0.00284f
C3786 vdd.n1136 vss 0.00219f
C3787 vdd.n1137 vss 0.00219f
C3788 vdd.n1138 vss 2.58e-19
C3789 vdd.n1139 vss 0.0193f
C3790 vdd.n1140 vss 0.101f
C3791 vdd.t63 vss 0.384f
C3792 vdd.n1141 vss 0.169f
C3793 vdd.t74 vss 0.207f
C3794 vdd.n1142 vss 0.162f
C3795 vdd.n1143 vss 0.00851f
C3796 vdd.n1144 vss 0.00219f
C3797 vdd.n1145 vss 0.00542f
C3798 vdd.n1146 vss 0.00284f
C3799 vdd.n1147 vss 0.00658f
C3800 vdd.n1148 vss 0.00271f
C3801 vdd.n1149 vss 0.00638f
C3802 vdd.n1150 vss 0.00359f
C3803 vdd.n1151 vss 0.0113f
C3804 vdd.n1152 vss 0.0116f
C3805 vdd.n1153 vss -0.0615f
C3806 vdd.n1154 vss 0.00335f
C3807 vdd.n1155 vss 0.00477f
C3808 vdd.n1156 vss -0.173f
C3809 vdd.n1157 vss 0.00319f
C3810 vdd.n1158 vss 0.0188f
C3811 vdd.n1159 vss 0.0184f
C3812 vdd.n1160 vss -0.148f
C3813 vdd.n1161 vss 0.00399f
C3814 vdd.n1162 vss 2.66e-19
C3815 vdd.n1163 vss 0.00284f
C3816 vdd.n1164 vss 0.00271f
C3817 vdd.n1165 vss 0.00219f
C3818 vdd.n1166 vss 0.00748f
C3819 vdd.n1167 vss 0.00219f
C3820 vdd.n1168 vss 0.00219f
C3821 vdd.n1169 vss 0.0105f
C3822 vdd.n1170 vss 0.00226f
C3823 vdd.n1171 vss 2.58e-19
C3824 vdd.n1172 vss 0.00748f
C3825 vdd.n1173 vss 0.00335f
C3826 vdd.n1174 vss 0.00477f
C3827 vdd.n1175 vss 0.00658f
C3828 vdd.n1176 vss 0.00542f
C3829 vdd.n1177 vss 0.00271f
C3830 vdd.n1178 vss 0.008f
C3831 vdd.n1179 vss 0.008f
C3832 vdd.n1180 vss 0.00219f
C3833 vdd.n1181 vss 0.00226f
C3834 vdd.n1182 vss 0.043f
C3835 vdd.n1183 vss 0.2f
C3836 vdd.n1184 vss 0.162f
C3837 vdd.n1185 vss 0.00851f
C3838 vdd.n1186 vss 0.00219f
C3839 vdd.n1187 vss 0.00542f
C3840 vdd.n1188 vss 0.00284f
C3841 vdd.n1189 vss 0.00658f
C3842 vdd.n1190 vss 0.00271f
C3843 vdd.n1191 vss 0.00638f
C3844 vdd.n1192 vss -0.0615f
C3845 vdd.n1193 vss -0.0637f
C3846 vdd.n1194 vss 0.0116f
C3847 vdd.n1195 vss 0.00359f
C3848 vdd.n1196 vss 0.00335f
C3849 vdd.n1197 vss 0.00477f
C3850 vdd.n1198 vss 0.00399f
C3851 vdd.n1199 vss 0.00319f
C3852 vdd.n1200 vss 0.0188f
C3853 vdd.n1201 vss 0.0184f
C3854 vdd.n1202 vss 0.0184f
C3855 vdd.n1203 vss -0.173f
C3856 vdd.n1204 vss 2.66e-19
C3857 vdd.n1205 vss 0.00284f
C3858 vdd.n1206 vss 0.00271f
C3859 vdd.n1207 vss 0.00219f
C3860 vdd.n1208 vss 0.00748f
C3861 vdd.n1209 vss 0.00219f
C3862 vdd.n1210 vss 0.00219f
C3863 vdd.n1211 vss 0.0105f
C3864 vdd.n1212 vss 0.00226f
C3865 vdd.n1213 vss 2.58e-19
C3866 vdd.n1214 vss 0.00748f
C3867 vdd.n1215 vss 0.00335f
C3868 vdd.n1216 vss 0.00477f
C3869 vdd.n1217 vss 0.00658f
C3870 vdd.n1218 vss 0.00542f
C3871 vdd.n1219 vss 0.00271f
C3872 vdd.n1220 vss 0.008f
C3873 vdd.n1221 vss 0.008f
C3874 vdd.n1222 vss 0.00219f
C3875 vdd.n1223 vss 0.00226f
C3876 vdd.n1224 vss 0.043f
C3877 vdd.n1225 vss 0.2f
C3878 vdd.n1226 vss 0.162f
C3879 vdd.n1227 vss 0.00851f
C3880 vdd.n1228 vss 0.00219f
C3881 vdd.n1229 vss 0.00542f
C3882 vdd.n1230 vss 0.00284f
C3883 vdd.n1231 vss 0.00658f
C3884 vdd.n1232 vss 0.00271f
C3885 vdd.n1233 vss 0.00638f
C3886 vdd.n1234 vss 0.00359f
C3887 vdd.n1235 vss 0.0113f
C3888 vdd.n1236 vss 0.0116f
C3889 vdd.n1237 vss 0.00359f
C3890 vdd.n1238 vss 0.00335f
C3891 vdd.n1239 vss 0.00477f
C3892 vdd.n1240 vss 0.00399f
C3893 vdd.n1241 vss 0.00319f
C3894 vdd.n1242 vss 0.0188f
C3895 vdd.n1243 vss -0.148f
C3896 vdd.n1244 vss 0.00399f
C3897 vdd.n1245 vss 0.00385f
C3898 vdd.n1246 vss -0.0689f
C3899 vdd.n1247 vss 2.66e-19
C3900 vdd.n1248 vss 0.00335f
C3901 vdd.n1249 vss 0.00284f
C3902 vdd.n1250 vss 0.00399f
C3903 vdd.n1251 vss 0.0205f
C3904 vdd.n1252 vss 0.0205f
C3905 vdd.n1253 vss 0.00335f
C3906 vdd.n1254 vss 0.0241f
C3907 vdd.n1255 vss 0.0241f
C3908 vdd.n1256 vss 0.00219f
C3909 vdd.n1257 vss 0.00219f
C3910 vdd.n1258 vss 0.00219f
C3911 vdd.n1259 vss 0.00226f
C3912 vdd.n1260 vss 0.0105f
C3913 vdd.n1261 vss 2.58e-19
C3914 vdd.n1262 vss 0.00219f
C3915 vdd.n1263 vss 0.00226f
C3916 vdd.n1264 vss 0.043f
C3917 vdd.n1265 vss 0.336f
C3918 vdd.n1266 vss 0.0152f
C3919 vdd.n1267 vss 0.0245f
C3920 vdd.n1268 vss 0.0245f
C3921 vdd.n1269 vss 0.0152f
C3922 vdd.n1270 vss 0.185f
C3923 vdd.n1271 vss 0.043f
C3924 vdd.n1272 vss 0.162f
C3925 vdd.n1273 vss 0.00851f
C3926 vdd.n1274 vss 0.008f
C3927 vdd.n1275 vss 0.00219f
C3928 vdd.n1276 vss 0.00748f
C3929 vdd.n1277 vss 3.87e-19
C3930 vdd.n1278 vss 0.00271f
C3931 vdd.n1279 vss 0.00477f
C3932 vdd.n1280 vss 0.00284f
C3933 vdd.n1281 vss 3.87e-19
C3934 vdd.n1282 vss -0.173f
C3935 vdd.n1283 vss 2.66e-19
C3936 vdd.n1284 vss 0.0188f
C3937 vdd.n1285 vss 0.00359f
C3938 vdd.n1286 vss -0.142f
C3939 vdd.n1287 vss 0.00651f
C3940 vdd.n1288 vss 0.008f
C3941 vdd.n1289 vss 0.00271f
C3942 vdd.n1290 vss 0.00542f
C3943 vdd.n1291 vss 0.00658f
C3944 vdd.n1292 vss 0.00271f
C3945 vdd.n1293 vss 0.00335f
C3946 vdd.n1294 vss 0.00477f
C3947 vdd.n1295 vss 0.00385f
C3948 vdd.n1296 vss 0.00306f
C3949 vdd.n1297 vss 0.0184f
C3950 vdd.n1298 vss 0.0113f
C3951 vdd.n1299 vss 0.0116f
C3952 vdd.n1300 vss 2.66e-19
C3953 vdd.n1301 vss 0.00399f
C3954 vdd.n1302 vss 0.00651f
C3955 vdd.n1303 vss 0.00306f
C3956 vdd.n1304 vss 0.0184f
C3957 vdd.n1305 vss 0.0184f
C3958 vdd.n1306 vss 0.00399f
C3959 vdd.n1307 vss 0.00359f
C3960 vdd.n1308 vss 0.00658f
C3961 vdd.n1309 vss 0.00271f
C3962 vdd.n1310 vss 0.00542f
C3963 vdd.n1311 vss 3.87e-19
C3964 vdd.n1312 vss 0.00219f
C3965 vdd.n1313 vss 0.00219f
C3966 vdd.n1314 vss 0.00219f
C3967 vdd.n1315 vss 0.00226f
C3968 vdd.n1316 vss 0.0105f
C3969 vdd.n1317 vss 0.162f
C3970 vdd.n1318 vss 0.00851f
C3971 vdd.n1319 vss 0.008f
C3972 vdd.n1320 vss 0.008f
C3973 vdd.n1321 vss 0.0105f
C3974 vdd.n1322 vss 0.2f
C3975 vdd.n1323 vss 0.043f
C3976 vdd.n1324 vss 0.00226f
C3977 vdd.n1325 vss 0.00219f
C3978 vdd.n1326 vss 2.58e-19
C3979 vdd.n1327 vss 0.00219f
C3980 vdd.n1328 vss 0.00284f
C3981 vdd.n1329 vss 0.00219f
C3982 vdd.n1330 vss 0.00271f
C3983 vdd.n1331 vss 0.008f
C3984 vdd.n1332 vss 0.008f
C3985 vdd.n1333 vss 0.0105f
C3986 vdd.n1334 vss 0.2f
C3987 vdd.n1335 vss 0.043f
C3988 vdd.n1336 vss 0.162f
C3989 vdd.n1337 vss 0.00851f
C3990 vdd.n1338 vss 0.008f
C3991 vdd.n1339 vss 0.00219f
C3992 vdd.n1340 vss 0.00748f
C3993 vdd.n1341 vss 3.87e-19
C3994 vdd.n1342 vss 0.00271f
C3995 vdd.n1343 vss 0.00477f
C3996 vdd.n1344 vss 0.00284f
C3997 vdd.n1345 vss 3.87e-19
C3998 vdd.n1346 vss -0.173f
C3999 vdd.n1347 vss 2.66e-19
C4000 vdd.n1348 vss 0.0188f
C4001 vdd.n1349 vss 0.00359f
C4002 vdd.n1350 vss -0.142f
C4003 vdd.n1351 vss 0.0113f
C4004 vdd.n1352 vss -0.0689f
C4005 vdd.n1353 vss 2.66e-19
C4006 vdd.n1354 vss 0.00399f
C4007 vdd.n1355 vss 0.00651f
C4008 vdd.n1356 vss 0.00284f
C4009 vdd.n1357 vss 0.008f
C4010 vdd.n1358 vss 0.00271f
C4011 vdd.n1359 vss 0.00542f
C4012 vdd.n1360 vss 0.00658f
C4013 vdd.n1361 vss 0.00271f
C4014 vdd.n1362 vss 0.00335f
C4015 vdd.n1363 vss 0.00477f
C4016 vdd.n1364 vss 0.00385f
C4017 vdd.n1365 vss 0.00306f
C4018 vdd.n1366 vss 0.0184f
C4019 vdd.n1367 vss 0.0113f
C4020 vdd.n1368 vss 0.0116f
C4021 vdd.n1369 vss 2.66e-19
C4022 vdd.n1370 vss 0.00399f
C4023 vdd.n1371 vss 0.00651f
C4024 vdd.n1372 vss 0.00306f
C4025 vdd.n1373 vss 0.0184f
C4026 vdd.n1374 vss 0.0661f
C4027 vdd.n1375 vss 0.00399f
C4028 vdd.n1376 vss 2.66e-19
C4029 vdd.n1377 vss 0.00284f
C4030 vdd.n1378 vss 0.00271f
C4031 vdd.n1379 vss 0.00219f
C4032 vdd.n1380 vss 0.00748f
C4033 vdd.n1381 vss 0.00219f
C4034 vdd.n1382 vss 0.00219f
C4035 vdd.n1383 vss 0.00226f
C4036 vdd.n1384 vss 0.043f
C4037 vdd.n1385 vss 0.00226f
C4038 vdd.n1386 vss 0.008f
C4039 vdd.n1387 vss 0.2f
C4040 vdd.n1388 vss 0.0105f
C4041 vdd.n1389 vss 0.008f
C4042 vdd.n1390 vss 0.00219f
C4043 vdd.n1391 vss 0.024f
C4044 vdd.n1392 vss 0.00271f
C4045 vdd.n1393 vss 0.0234f
C4046 vdd.n1394 vss 0.024f
C4047 vdd.n1395 vss 0.00271f
C4048 vdd.n1396 vss 0.0213f
C4049 vdd.n1397 vss 0.0213f
C4050 vdd.n1398 vss 0.0234f
C4051 vdd.n1399 vss 0.00284f
C4052 vdd.n1400 vss 0.00219f
C4053 vdd.n1401 vss 0.00219f
C4054 vdd.n1402 vss 2.58e-19
C4055 vdd.n1403 vss 0.0193f
C4056 vdd.n1404 vss 0.101f
C4057 vdd.t94 vss 0.384f
C4058 vdd.n1405 vss 0.169f
C4059 vdd.t125 vss 0.207f
C4060 vdd.n1406 vss 0.162f
C4061 vdd.n1407 vss 0.00851f
C4062 vdd.n1408 vss 0.00219f
C4063 vdd.n1409 vss 0.00542f
C4064 vdd.n1410 vss 0.00284f
C4065 vdd.n1411 vss 0.00658f
C4066 vdd.n1412 vss 0.00271f
C4067 vdd.n1413 vss 0.00638f
C4068 vdd.n1414 vss 0.00359f
C4069 vdd.n1415 vss 0.0113f
C4070 vdd.n1416 vss 0.0116f
C4071 vdd.n1417 vss -0.0615f
C4072 vdd.n1418 vss 0.00335f
C4073 vdd.n1419 vss 0.00477f
C4074 vdd.n1420 vss -0.173f
C4075 vdd.n1421 vss 0.00319f
C4076 vdd.n1422 vss 0.0188f
C4077 vdd.n1423 vss 0.0184f
C4078 vdd.n1424 vss -0.148f
C4079 vdd.n1425 vss 0.00399f
C4080 vdd.n1426 vss 2.66e-19
C4081 vdd.n1427 vss 0.00284f
C4082 vdd.n1428 vss 0.00271f
C4083 vdd.n1429 vss 0.00219f
C4084 vdd.n1430 vss 0.00748f
C4085 vdd.n1431 vss 0.00219f
C4086 vdd.n1432 vss 0.00219f
C4087 vdd.n1433 vss 0.0105f
C4088 vdd.n1434 vss 0.00226f
C4089 vdd.n1435 vss 2.58e-19
C4090 vdd.n1436 vss 0.00748f
C4091 vdd.n1437 vss 0.00335f
C4092 vdd.n1438 vss 0.00477f
C4093 vdd.n1439 vss 0.00658f
C4094 vdd.n1440 vss 0.00542f
C4095 vdd.n1441 vss 0.00271f
C4096 vdd.n1442 vss 0.008f
C4097 vdd.n1443 vss 0.008f
C4098 vdd.n1444 vss 0.00219f
C4099 vdd.n1445 vss 0.00226f
C4100 vdd.n1446 vss 0.043f
C4101 vdd.n1447 vss 0.2f
C4102 vdd.n1448 vss 0.162f
C4103 vdd.n1449 vss 0.00851f
C4104 vdd.n1450 vss 0.00219f
C4105 vdd.n1451 vss 0.00542f
C4106 vdd.n1452 vss 0.00284f
C4107 vdd.n1453 vss 0.00658f
C4108 vdd.n1454 vss 0.00271f
C4109 vdd.n1455 vss 0.00638f
C4110 vdd.n1456 vss -0.0615f
C4111 vdd.n1457 vss -0.0637f
C4112 vdd.n1458 vss 0.0116f
C4113 vdd.n1459 vss 0.00359f
C4114 vdd.n1460 vss 0.00335f
C4115 vdd.n1461 vss 0.00477f
C4116 vdd.n1462 vss 0.00399f
C4117 vdd.n1463 vss 0.00319f
C4118 vdd.n1464 vss 0.0188f
C4119 vdd.n1465 vss 0.0184f
C4120 vdd.n1466 vss 0.0184f
C4121 vdd.n1467 vss -0.173f
C4122 vdd.n1468 vss 2.66e-19
C4123 vdd.n1469 vss 0.00284f
C4124 vdd.n1470 vss 0.00271f
C4125 vdd.n1471 vss 0.00219f
C4126 vdd.n1472 vss 0.00748f
C4127 vdd.n1473 vss 0.00219f
C4128 vdd.n1474 vss 0.00219f
C4129 vdd.n1475 vss 0.0105f
C4130 vdd.n1476 vss 0.00226f
C4131 vdd.n1477 vss 2.58e-19
C4132 vdd.n1478 vss 0.00748f
C4133 vdd.n1479 vss 0.00335f
C4134 vdd.n1480 vss 0.00477f
C4135 vdd.n1481 vss 0.00658f
C4136 vdd.n1482 vss 0.00542f
C4137 vdd.n1483 vss 0.00271f
C4138 vdd.n1484 vss 0.008f
C4139 vdd.n1485 vss 0.008f
C4140 vdd.n1486 vss 0.00219f
C4141 vdd.n1487 vss 0.00226f
C4142 vdd.n1488 vss 0.043f
C4143 vdd.n1489 vss 0.2f
C4144 vdd.n1490 vss 0.162f
C4145 vdd.n1491 vss 0.00851f
C4146 vdd.n1492 vss 0.00219f
C4147 vdd.n1493 vss 0.00542f
C4148 vdd.n1494 vss 0.00284f
C4149 vdd.n1495 vss 0.00658f
C4150 vdd.n1496 vss 0.00271f
C4151 vdd.n1497 vss 0.00638f
C4152 vdd.n1498 vss 0.00359f
C4153 vdd.n1499 vss 0.0113f
C4154 vdd.n1500 vss 0.0116f
C4155 vdd.n1501 vss 0.00359f
C4156 vdd.n1502 vss 0.00335f
C4157 vdd.n1503 vss 0.00477f
C4158 vdd.n1504 vss 0.00399f
C4159 vdd.n1505 vss 0.00319f
C4160 vdd.n1506 vss 0.0188f
C4161 vdd.n1507 vss -0.148f
C4162 vdd.n1508 vss 0.00399f
C4163 vdd.n1509 vss 0.00385f
C4164 vdd.n1510 vss -0.0689f
C4165 vdd.n1511 vss 2.66e-19
C4166 vdd.n1512 vss 0.00335f
C4167 vdd.n1513 vss 0.00284f
C4168 vdd.n1514 vss 0.00399f
C4169 vdd.n1515 vss 0.0205f
C4170 vdd.n1516 vss 0.0205f
C4171 vdd.n1517 vss 0.00335f
C4172 vdd.n1518 vss 0.0241f
C4173 vdd.n1519 vss 0.0241f
C4174 vdd.n1520 vss 0.00219f
C4175 vdd.n1521 vss 0.00219f
C4176 vdd.n1522 vss 0.00219f
C4177 vdd.n1523 vss 0.00226f
C4178 vdd.n1524 vss 0.0105f
C4179 vdd.n1525 vss 2.58e-19
C4180 vdd.n1526 vss 0.00219f
C4181 vdd.n1527 vss 0.00226f
C4182 vdd.n1528 vss 0.043f
C4183 vdd.n1529 vss 0.336f
C4184 vdd.n1530 vss 0.0152f
C4185 vdd.n1531 vss 0.0245f
C4186 vdd.n1532 vss 0.0245f
C4187 vdd.n1533 vss 0.0152f
C4188 vdd.n1534 vss 0.185f
C4189 vdd.n1535 vss 0.043f
C4190 vdd.n1536 vss 0.162f
C4191 vdd.n1537 vss 0.00851f
C4192 vdd.n1538 vss 0.008f
C4193 vdd.n1539 vss 0.00219f
C4194 vdd.n1540 vss 0.00748f
C4195 vdd.n1541 vss 3.87e-19
C4196 vdd.n1542 vss 0.00271f
C4197 vdd.n1543 vss 0.00477f
C4198 vdd.n1544 vss 0.00284f
C4199 vdd.n1545 vss 3.87e-19
C4200 vdd.n1546 vss -0.173f
C4201 vdd.n1547 vss 2.66e-19
C4202 vdd.n1548 vss 0.0188f
C4203 vdd.n1549 vss 0.00359f
C4204 vdd.n1550 vss -0.142f
C4205 vdd.n1551 vss 0.00651f
C4206 vdd.n1552 vss 0.008f
C4207 vdd.n1553 vss 0.00271f
C4208 vdd.n1554 vss 0.00542f
C4209 vdd.n1555 vss 0.00658f
C4210 vdd.n1556 vss 0.00271f
C4211 vdd.n1557 vss 0.00335f
C4212 vdd.n1558 vss 0.00477f
C4213 vdd.n1559 vss 0.00385f
C4214 vdd.n1560 vss 0.00306f
C4215 vdd.n1561 vss 0.0184f
C4216 vdd.n1562 vss 0.0113f
C4217 vdd.n1563 vss 0.0116f
C4218 vdd.n1564 vss 2.66e-19
C4219 vdd.n1565 vss 0.00399f
C4220 vdd.n1566 vss 0.00651f
C4221 vdd.n1567 vss 0.00306f
C4222 vdd.n1568 vss 0.0184f
C4223 vdd.n1569 vss 0.0184f
C4224 vdd.n1570 vss 0.00399f
C4225 vdd.n1571 vss 0.00359f
C4226 vdd.n1572 vss 0.00658f
C4227 vdd.n1573 vss 0.00271f
C4228 vdd.n1574 vss 0.00542f
C4229 vdd.n1575 vss 3.87e-19
C4230 vdd.n1576 vss 0.00219f
C4231 vdd.n1577 vss 0.00219f
C4232 vdd.n1578 vss 0.00219f
C4233 vdd.n1579 vss 0.00226f
C4234 vdd.n1580 vss 0.0105f
C4235 vdd.n1581 vss 0.162f
C4236 vdd.n1582 vss 0.00851f
C4237 vdd.n1583 vss 0.008f
C4238 vdd.n1584 vss 0.008f
C4239 vdd.n1585 vss 0.0105f
C4240 vdd.n1586 vss 0.2f
C4241 vdd.n1587 vss 0.043f
C4242 vdd.n1588 vss 0.00226f
C4243 vdd.n1589 vss 0.00219f
C4244 vdd.n1590 vss 2.58e-19
C4245 vdd.n1591 vss 0.00219f
C4246 vdd.n1592 vss 0.00284f
C4247 vdd.n1593 vss 0.00219f
C4248 vdd.n1594 vss 0.00271f
C4249 vdd.n1595 vss 0.008f
C4250 vdd.n1596 vss 0.008f
C4251 vdd.n1597 vss 0.0105f
C4252 vdd.n1598 vss 0.2f
C4253 vdd.n1599 vss 0.043f
C4254 vdd.n1600 vss 0.162f
C4255 vdd.n1601 vss 0.00851f
C4256 vdd.n1602 vss 0.008f
C4257 vdd.n1603 vss 0.00219f
C4258 vdd.n1604 vss 0.00748f
C4259 vdd.n1605 vss 3.87e-19
C4260 vdd.n1606 vss 0.00271f
C4261 vdd.n1607 vss 0.00477f
C4262 vdd.n1608 vss 0.00284f
C4263 vdd.n1609 vss 3.87e-19
C4264 vdd.n1610 vss -0.173f
C4265 vdd.n1611 vss 2.66e-19
C4266 vdd.n1612 vss 0.0188f
C4267 vdd.n1613 vss 0.00359f
C4268 vdd.n1614 vss -0.142f
C4269 vdd.n1615 vss 0.0113f
C4270 vdd.n1616 vss -0.0689f
C4271 vdd.n1617 vss 2.66e-19
C4272 vdd.n1618 vss 0.00399f
C4273 vdd.n1619 vss 0.00651f
C4274 vdd.n1620 vss 0.00284f
C4275 vdd.n1621 vss 0.008f
C4276 vdd.n1622 vss 0.00271f
C4277 vdd.n1623 vss 0.00542f
C4278 vdd.n1624 vss 0.00658f
C4279 vdd.n1625 vss 0.00271f
C4280 vdd.n1626 vss 0.00335f
C4281 vdd.n1627 vss 0.00477f
C4282 vdd.n1628 vss 0.00385f
C4283 vdd.n1629 vss 0.00306f
C4284 vdd.n1630 vss 0.0184f
C4285 vdd.n1631 vss 0.0113f
C4286 vdd.n1632 vss 0.0116f
C4287 vdd.n1633 vss 2.66e-19
C4288 vdd.n1634 vss 0.00399f
C4289 vdd.n1635 vss 0.00651f
C4290 vdd.n1636 vss 0.00306f
C4291 vdd.n1637 vss 0.0184f
C4292 vdd.n1638 vss 0.0661f
C4293 vdd.n1639 vss 0.00399f
C4294 vdd.n1640 vss 2.66e-19
C4295 vdd.n1641 vss 0.00284f
C4296 vdd.n1642 vss 0.00271f
C4297 vdd.n1643 vss 0.00219f
C4298 vdd.n1644 vss 0.00748f
C4299 vdd.n1645 vss 0.00219f
C4300 vdd.n1646 vss 0.00219f
C4301 vdd.n1647 vss 0.00226f
C4302 vdd.n1648 vss 0.043f
C4303 vdd.n1649 vss 0.00226f
C4304 vdd.n1650 vss 0.008f
C4305 vdd.n1651 vss 0.2f
C4306 vdd.n1652 vss 0.0105f
C4307 vdd.n1653 vss 0.008f
C4308 vdd.n1654 vss 0.00219f
C4309 vdd.n1655 vss 0.024f
C4310 vdd.n1656 vss 0.00271f
C4311 vdd.n1657 vss 0.0234f
C4312 vdd.n1658 vss 0.024f
C4313 vdd.n1659 vss 0.00271f
C4314 vdd.n1660 vss 0.0213f
C4315 vdd.n1661 vss 0.0213f
C4316 vdd.n1662 vss 0.0234f
C4317 vdd.n1663 vss 0.00284f
C4318 vdd.n1664 vss 0.00219f
C4319 vdd.n1665 vss 0.00219f
C4320 vdd.n1666 vss 2.58e-19
C4321 vdd.n1667 vss 0.0193f
C4322 vdd.n1668 vss 0.101f
C4323 vdd.t124 vss 0.384f
C4324 vdd.n1669 vss 0.169f
C4325 vdd.t112 vss 0.207f
C4326 vdd.n1670 vss 0.162f
C4327 vdd.n1671 vss 0.00851f
C4328 vdd.n1672 vss 0.00219f
C4329 vdd.n1673 vss 0.00542f
C4330 vdd.n1674 vss 0.00284f
C4331 vdd.n1675 vss 0.00658f
C4332 vdd.n1676 vss 0.00271f
C4333 vdd.n1677 vss 0.00638f
C4334 vdd.n1678 vss 0.00359f
C4335 vdd.n1679 vss 0.0113f
C4336 vdd.n1680 vss 0.0116f
C4337 vdd.n1681 vss -0.0615f
C4338 vdd.n1682 vss 0.00335f
C4339 vdd.n1683 vss 0.00477f
C4340 vdd.n1684 vss -0.173f
C4341 vdd.n1685 vss 0.00319f
C4342 vdd.n1686 vss 0.0188f
C4343 vdd.n1687 vss 0.0184f
C4344 vdd.n1688 vss -0.148f
C4345 vdd.n1689 vss 0.00399f
C4346 vdd.n1690 vss 2.66e-19
C4347 vdd.n1691 vss 0.00284f
C4348 vdd.n1692 vss 0.00271f
C4349 vdd.n1693 vss 0.00219f
C4350 vdd.n1694 vss 0.00748f
C4351 vdd.n1695 vss 0.00219f
C4352 vdd.n1696 vss 0.00219f
C4353 vdd.n1697 vss 0.0105f
C4354 vdd.n1698 vss 0.00226f
C4355 vdd.n1699 vss 2.58e-19
C4356 vdd.n1700 vss 0.00748f
C4357 vdd.n1701 vss 0.00335f
C4358 vdd.n1702 vss 0.00477f
C4359 vdd.n1703 vss 0.00658f
C4360 vdd.n1704 vss 0.00542f
C4361 vdd.n1705 vss 0.00271f
C4362 vdd.n1706 vss 0.008f
C4363 vdd.n1707 vss 0.008f
C4364 vdd.n1708 vss 0.00219f
C4365 vdd.n1709 vss 0.00226f
C4366 vdd.n1710 vss 0.043f
C4367 vdd.n1711 vss 0.2f
C4368 vdd.n1712 vss 0.162f
C4369 vdd.n1713 vss 0.00851f
C4370 vdd.n1714 vss 0.00219f
C4371 vdd.n1715 vss 0.00542f
C4372 vdd.n1716 vss 0.00284f
C4373 vdd.n1717 vss 0.00658f
C4374 vdd.n1718 vss 0.00271f
C4375 vdd.n1719 vss 0.00638f
C4376 vdd.n1720 vss -0.0615f
C4377 vdd.n1721 vss -0.0637f
C4378 vdd.n1722 vss 0.0116f
C4379 vdd.n1723 vss 0.00359f
C4380 vdd.n1724 vss 0.00335f
C4381 vdd.n1725 vss 0.00477f
C4382 vdd.n1726 vss 0.00399f
C4383 vdd.n1727 vss 0.00319f
C4384 vdd.n1728 vss 0.0188f
C4385 vdd.n1729 vss 0.0184f
C4386 vdd.n1730 vss 0.0184f
C4387 vdd.n1731 vss -0.173f
C4388 vdd.n1732 vss 2.66e-19
C4389 vdd.n1733 vss 0.00284f
C4390 vdd.n1734 vss 0.00271f
C4391 vdd.n1735 vss 0.00219f
C4392 vdd.n1736 vss 0.00748f
C4393 vdd.n1737 vss 0.00219f
C4394 vdd.n1738 vss 0.00219f
C4395 vdd.n1739 vss 0.0105f
C4396 vdd.n1740 vss 0.00226f
C4397 vdd.n1741 vss 2.58e-19
C4398 vdd.n1742 vss 0.00748f
C4399 vdd.n1743 vss 0.00335f
C4400 vdd.n1744 vss 0.00477f
C4401 vdd.n1745 vss 0.00658f
C4402 vdd.n1746 vss 0.00542f
C4403 vdd.n1747 vss 0.00271f
C4404 vdd.n1748 vss 0.008f
C4405 vdd.n1749 vss 0.008f
C4406 vdd.n1750 vss 0.00219f
C4407 vdd.n1751 vss 0.00226f
C4408 vdd.n1752 vss 0.043f
C4409 vdd.n1753 vss 0.2f
C4410 vdd.n1754 vss 0.162f
C4411 vdd.n1755 vss 0.00851f
C4412 vdd.n1756 vss 0.00219f
C4413 vdd.n1757 vss 0.00542f
C4414 vdd.n1758 vss 0.00284f
C4415 vdd.n1759 vss 0.00658f
C4416 vdd.n1760 vss 0.00271f
C4417 vdd.n1761 vss 0.00638f
C4418 vdd.n1762 vss 0.00359f
C4419 vdd.n1763 vss 0.0113f
C4420 vdd.n1764 vss 0.0116f
C4421 vdd.n1765 vss 0.00359f
C4422 vdd.n1766 vss 0.00335f
C4423 vdd.n1767 vss 0.00477f
C4424 vdd.n1768 vss 0.00399f
C4425 vdd.n1769 vss 0.00319f
C4426 vdd.n1770 vss 0.0188f
C4427 vdd.n1771 vss -0.148f
C4428 vdd.n1772 vss 0.00399f
C4429 vdd.n1773 vss 0.00385f
C4430 vdd.n1774 vss -0.0689f
C4431 vdd.n1775 vss 2.66e-19
C4432 vdd.n1776 vss 0.00335f
C4433 vdd.n1777 vss 0.00284f
C4434 vdd.n1778 vss 0.00399f
C4435 vdd.n1779 vss 0.0205f
C4436 vdd.n1780 vss 0.0205f
C4437 vdd.n1781 vss 0.00335f
C4438 vdd.n1782 vss 0.0241f
C4439 vdd.n1783 vss 0.0241f
C4440 vdd.n1784 vss 0.00219f
C4441 vdd.n1785 vss 0.00219f
C4442 vdd.n1786 vss 0.00219f
C4443 vdd.n1787 vss 0.00226f
C4444 vdd.n1788 vss 0.0105f
C4445 vdd.n1789 vss 2.58e-19
C4446 vdd.n1790 vss 0.00219f
C4447 vdd.n1791 vss 0.00226f
C4448 vdd.n1792 vss 0.043f
C4449 vdd.n1793 vss 0.336f
C4450 vdd.n1794 vss 0.0152f
C4451 vdd.n1795 vss 0.0245f
C4452 vdd.n1796 vss 0.0245f
C4453 vdd.n1797 vss 0.0152f
C4454 vdd.n1798 vss 0.185f
C4455 vdd.n1799 vss 0.043f
C4456 vdd.n1800 vss 0.162f
C4457 vdd.n1801 vss 0.00851f
C4458 vdd.n1802 vss 0.008f
C4459 vdd.n1803 vss 0.00219f
C4460 vdd.n1804 vss 0.00748f
C4461 vdd.n1805 vss 3.87e-19
C4462 vdd.n1806 vss 0.00271f
C4463 vdd.n1807 vss 0.00477f
C4464 vdd.n1808 vss 0.00284f
C4465 vdd.n1809 vss 3.87e-19
C4466 vdd.n1810 vss -0.173f
C4467 vdd.n1811 vss 2.66e-19
C4468 vdd.n1812 vss 0.0188f
C4469 vdd.n1813 vss 0.00359f
C4470 vdd.n1814 vss -0.142f
C4471 vdd.n1815 vss 0.00651f
C4472 vdd.n1816 vss 0.008f
C4473 vdd.n1817 vss 0.00271f
C4474 vdd.n1818 vss 0.00542f
C4475 vdd.n1819 vss 0.00658f
C4476 vdd.n1820 vss 0.00271f
C4477 vdd.n1821 vss 0.00335f
C4478 vdd.n1822 vss 0.00477f
C4479 vdd.n1823 vss 0.00385f
C4480 vdd.n1824 vss 0.00306f
C4481 vdd.n1825 vss 0.0184f
C4482 vdd.n1826 vss 0.0113f
C4483 vdd.n1827 vss 0.0116f
C4484 vdd.n1828 vss 2.66e-19
C4485 vdd.n1829 vss 0.00399f
C4486 vdd.n1830 vss 0.00651f
C4487 vdd.n1831 vss 0.00306f
C4488 vdd.n1832 vss 0.0184f
C4489 vdd.n1833 vss 0.0184f
C4490 vdd.n1834 vss 0.00399f
C4491 vdd.n1835 vss 0.00359f
C4492 vdd.n1836 vss 0.00658f
C4493 vdd.n1837 vss 0.00271f
C4494 vdd.n1838 vss 0.00542f
C4495 vdd.n1839 vss 3.87e-19
C4496 vdd.n1840 vss 0.00219f
C4497 vdd.n1841 vss 0.00219f
C4498 vdd.n1842 vss 0.00219f
C4499 vdd.n1843 vss 0.00226f
C4500 vdd.n1844 vss 0.0105f
C4501 vdd.n1845 vss 0.162f
C4502 vdd.n1846 vss 0.00851f
C4503 vdd.n1847 vss 0.008f
C4504 vdd.n1848 vss 0.008f
C4505 vdd.n1849 vss 0.0105f
C4506 vdd.n1850 vss 0.2f
C4507 vdd.n1851 vss 0.043f
C4508 vdd.n1852 vss 0.00226f
C4509 vdd.n1853 vss 0.00219f
C4510 vdd.n1854 vss 2.58e-19
C4511 vdd.n1855 vss 0.00219f
C4512 vdd.n1856 vss 0.00284f
C4513 vdd.n1857 vss 0.00219f
C4514 vdd.n1858 vss 0.00271f
C4515 vdd.n1859 vss 0.008f
C4516 vdd.n1860 vss 0.008f
C4517 vdd.n1861 vss 0.0105f
C4518 vdd.n1862 vss 0.2f
C4519 vdd.n1863 vss 0.043f
C4520 vdd.n1864 vss 0.162f
C4521 vdd.n1865 vss 0.00851f
C4522 vdd.n1866 vss 0.008f
C4523 vdd.n1867 vss 0.00219f
C4524 vdd.n1868 vss 0.00748f
C4525 vdd.n1869 vss 3.87e-19
C4526 vdd.n1870 vss 0.00271f
C4527 vdd.n1871 vss 0.00477f
C4528 vdd.n1872 vss 0.00284f
C4529 vdd.n1873 vss 3.87e-19
C4530 vdd.n1874 vss -0.173f
C4531 vdd.n1875 vss 2.66e-19
C4532 vdd.n1876 vss 0.0188f
C4533 vdd.n1877 vss 0.00359f
C4534 vdd.n1878 vss -0.142f
C4535 vdd.n1879 vss 0.0113f
C4536 vdd.n1880 vss -0.0689f
C4537 vdd.n1881 vss 2.66e-19
C4538 vdd.n1882 vss 0.00399f
C4539 vdd.n1883 vss 0.00651f
C4540 vdd.n1884 vss 0.00284f
C4541 vdd.n1885 vss 0.008f
C4542 vdd.n1886 vss 0.00271f
C4543 vdd.n1887 vss 0.00542f
C4544 vdd.n1888 vss 0.00658f
C4545 vdd.n1889 vss 0.00271f
C4546 vdd.n1890 vss 0.00335f
C4547 vdd.n1891 vss 0.00477f
C4548 vdd.n1892 vss 0.00385f
C4549 vdd.n1893 vss 0.00306f
C4550 vdd.n1894 vss 0.0184f
C4551 vdd.n1895 vss 0.0113f
C4552 vdd.n1896 vss 0.0116f
C4553 vdd.n1897 vss 2.66e-19
C4554 vdd.n1898 vss 0.00399f
C4555 vdd.n1899 vss 0.00651f
C4556 vdd.n1900 vss 0.00306f
C4557 vdd.n1901 vss 0.0184f
C4558 vdd.n1902 vss 0.0661f
C4559 vdd.n1903 vss 0.00399f
C4560 vdd.n1904 vss 2.66e-19
C4561 vdd.n1905 vss 0.00284f
C4562 vdd.n1906 vss 0.00271f
C4563 vdd.n1907 vss 0.00219f
C4564 vdd.n1908 vss 0.00748f
C4565 vdd.n1909 vss 0.00219f
C4566 vdd.n1910 vss 0.00219f
C4567 vdd.n1911 vss 0.00226f
C4568 vdd.n1912 vss 0.043f
C4569 vdd.n1913 vss 0.00226f
C4570 vdd.n1914 vss 0.008f
C4571 vdd.n1915 vss 0.2f
C4572 vdd.n1916 vss 0.0105f
C4573 vdd.n1917 vss 0.008f
C4574 vdd.n1918 vss 0.00219f
C4575 vdd.n1919 vss 0.024f
C4576 vdd.n1920 vss 0.00271f
C4577 vdd.n1921 vss 0.0234f
C4578 vdd.n1922 vss 0.024f
C4579 vdd.n1923 vss 0.00271f
C4580 vdd.n1924 vss 0.0213f
C4581 vdd.n1925 vss 0.0213f
C4582 vdd.n1926 vss 0.0234f
C4583 vdd.n1927 vss 0.00284f
C4584 vdd.n1928 vss 0.00219f
C4585 vdd.n1929 vss 0.00219f
C4586 vdd.n1930 vss 2.58e-19
C4587 vdd.n1931 vss 0.0193f
C4588 vdd.n1932 vss 0.101f
C4589 vdd.t62 vss 0.384f
C4590 vdd.n1933 vss 0.169f
C4591 vdd.t2 vss 0.207f
C4592 vdd.n1934 vss 0.162f
C4593 vdd.n1935 vss 0.00851f
C4594 vdd.n1936 vss 0.00219f
C4595 vdd.n1937 vss 0.00542f
C4596 vdd.n1938 vss 0.00284f
C4597 vdd.n1939 vss 0.00658f
C4598 vdd.n1940 vss 0.00271f
C4599 vdd.n1941 vss 0.00638f
C4600 vdd.n1942 vss 0.00359f
C4601 vdd.n1943 vss 0.0113f
C4602 vdd.n1944 vss 0.0116f
C4603 vdd.n1945 vss -0.0615f
C4604 vdd.n1946 vss 0.00335f
C4605 vdd.n1947 vss 0.00477f
C4606 vdd.n1948 vss -0.173f
C4607 vdd.n1949 vss 0.00319f
C4608 vdd.n1950 vss 0.0188f
C4609 vdd.n1951 vss 0.0184f
C4610 vdd.n1952 vss -0.148f
C4611 vdd.n1953 vss 0.00399f
C4612 vdd.n1954 vss 2.66e-19
C4613 vdd.n1955 vss 0.00284f
C4614 vdd.n1956 vss 0.00271f
C4615 vdd.n1957 vss 0.00219f
C4616 vdd.n1958 vss 0.00748f
C4617 vdd.n1959 vss 0.00219f
C4618 vdd.n1960 vss 0.00219f
C4619 vdd.n1961 vss 0.0105f
C4620 vdd.n1962 vss 0.00226f
C4621 vdd.n1963 vss 2.58e-19
C4622 vdd.n1964 vss 0.00748f
C4623 vdd.n1965 vss 0.00335f
C4624 vdd.n1966 vss 0.00477f
C4625 vdd.n1967 vss 0.00658f
C4626 vdd.n1968 vss 0.00542f
C4627 vdd.n1969 vss 0.00271f
C4628 vdd.n1970 vss 0.008f
C4629 vdd.n1971 vss 0.008f
C4630 vdd.n1972 vss 0.00219f
C4631 vdd.n1973 vss 0.00226f
C4632 vdd.n1974 vss 0.043f
C4633 vdd.n1975 vss 0.2f
C4634 vdd.n1976 vss 0.162f
C4635 vdd.n1977 vss 0.00851f
C4636 vdd.n1978 vss 0.00219f
C4637 vdd.n1979 vss 0.00542f
C4638 vdd.n1980 vss 0.00284f
C4639 vdd.n1981 vss 0.00658f
C4640 vdd.n1982 vss 0.00271f
C4641 vdd.n1983 vss 0.00638f
C4642 vdd.n1984 vss -0.0615f
C4643 vdd.n1985 vss -0.0637f
C4644 vdd.n1986 vss 0.0116f
C4645 vdd.n1987 vss 0.00359f
C4646 vdd.n1988 vss 0.00335f
C4647 vdd.n1989 vss 0.00477f
C4648 vdd.n1990 vss 0.00399f
C4649 vdd.n1991 vss 0.00319f
C4650 vdd.n1992 vss 0.0188f
C4651 vdd.n1993 vss 0.0184f
C4652 vdd.n1994 vss 0.0184f
C4653 vdd.n1995 vss -0.173f
C4654 vdd.n1996 vss 2.66e-19
C4655 vdd.n1997 vss 0.00284f
C4656 vdd.n1998 vss 0.00271f
C4657 vdd.n1999 vss 0.00219f
C4658 vdd.n2000 vss 0.00748f
C4659 vdd.n2001 vss 0.00219f
C4660 vdd.n2002 vss 0.00219f
C4661 vdd.n2003 vss 0.0105f
C4662 vdd.n2004 vss 0.00226f
C4663 vdd.n2005 vss 2.58e-19
C4664 vdd.n2006 vss 0.00748f
C4665 vdd.n2007 vss 0.00335f
C4666 vdd.n2008 vss 0.00477f
C4667 vdd.n2009 vss 0.00658f
C4668 vdd.n2010 vss 0.00542f
C4669 vdd.n2011 vss 0.00271f
C4670 vdd.n2012 vss 0.008f
C4671 vdd.n2013 vss 0.008f
C4672 vdd.n2014 vss 0.00219f
C4673 vdd.n2015 vss 0.00226f
C4674 vdd.n2016 vss 0.043f
C4675 vdd.n2017 vss 0.2f
C4676 vdd.n2018 vss 0.162f
C4677 vdd.n2019 vss 0.00851f
C4678 vdd.n2020 vss 0.00219f
C4679 vdd.n2021 vss 0.00542f
C4680 vdd.n2022 vss 0.0344f
C4681 vdd.n2023 vss 0.00658f
C4682 vdd.n2024 vss 0.00271f
C4683 vdd.n2025 vss 0.00638f
C4684 vdd.n2026 vss 0.00359f
C4685 vdd.n2027 vss 0.0113f
C4686 vdd.n2028 vss 0.0116f
C4687 vdd.n2029 vss 0.00359f
C4688 vdd.n2030 vss 0.00335f
C4689 vdd.n2031 vss 0.00477f
C4690 vdd.n2032 vss 0.00399f
C4691 vdd.n2033 vss 0.00319f
C4692 vdd.n2034 vss 0.0188f
C4693 vdd.n2035 vss -0.148f
C4694 vdd.n2036 vss 0.0727f
C4695 vdd.n2037 vss 0.0229f
C4696 vdd.n2038 vss 0.0142f
C4697 vdd.n2039 vss 0.00686f
C4698 vdd.n2040 vss 0.00335f
C4699 vdd.n2041 vss 0.0062f
C4700 vdd.n2042 vss 2.66e-19
C4701 vdd.n2043 vss 0.00271f
C4702 vdd.n2044 vss 0.0248f
C4703 vdd.n2045 vss 0.0118f
C4704 vdd.n2046 vss 0.0187f
C4705 vdd.n2047 vss 0.00399f
C4706 vdd.n2048 vss 0.00359f
C4707 vdd.n2049 vss 0.00658f
C4708 vdd.n2050 vss 0.00271f
C4709 vdd.n2051 vss 0.00542f
C4710 vdd.n2052 vss 3.87e-19
C4711 vdd.n2053 vss 0.00219f
C4712 vdd.n2054 vss 0.00219f
C4713 vdd.n2055 vss 0.00219f
C4714 vdd.n2056 vss 0.00226f
C4715 vdd.n2057 vss 0.0105f
C4716 vdd.n2064 vss 0.0193f
C4717 vdd.n2065 vss 0.355f
C4718 vdd.n2066 vss 0.00851f
C4719 vdd.n2067 vss 0.00226f
C4720 vdd.t26 vss 2.19f
C4721 vdd.n2068 vss 0.0527f
C4722 vdd.n2069 vss 0.29f
C4723 vdd.n2070 vss 0.00685f
C4724 vdd.n2071 vss 0.00518f
C4725 vdd.n2072 vss 0.00887f
C4726 vdd.n2073 vss 0.0641f
C4727 vdd.n2074 vss 0.0303f
C4728 vdd.n2075 vss 0.0163f
C4729 vdd.n2076 vss 0.0615f
C4730 vdd.n2077 vss 0.00518f
C4731 vdd.n2078 vss 0.00685f
C4732 vdd.n2079 vss 0.0261f
C4733 vdd.n2080 vss 0.0664f
C4734 vdd.n2081 vss 0.00685f
C4735 vdd.n2082 vss 0.00518f
C4736 vdd.n2083 vss 0.00887f
C4737 vdd.n2084 vss 0.114f
C4738 vdd.n2085 vss 0.0361f
C4739 vdd.n2086 vss 0.0163f
C4740 vdd.n2087 vss 0.114f
C4741 vdd.n2088 vss 0.00685f
C4742 vdd.n2089 vss 0.00518f
C4743 vdd.n2090 vss 0.00661f
C4744 vdd.n2091 vss 0.0163f
C4745 vdd.n2092 vss 0.00887f
C4746 vdd.n2093 vss 0.0512f
C4747 vdd.n2094 vss 0.00433f
C4748 vdd.n2095 vss 0.0253f
C4749 vdd.n2096 vss 0.0158f
C4750 vdd.n2097 vss 0.00246f
C4751 vdd.n2098 vss 0.00885f
C4752 vdd.n2099 vss 0.0159f
C4753 vdd.n2100 vss 0.0842f
C4754 vdd.t45 vss 0.0428f
C4755 vdd.n2101 vss 0.0451f
C4756 vdd.t64 vss 0.043f
C4757 vdd.n2102 vss 0.0378f
C4758 vdd.n2103 vss 0.00113f
C4759 vdd.n2104 vss 0.0445f
C4760 vdd.t132 vss 0.00929f
C4761 vdd.n2105 vss 0.0556f
C4762 vdd.n2106 vss 0.00607f
C4763 vdd.t77 vss 0.043f
C4764 vdd.n2107 vss 0.0329f
C4765 vdd.n2108 vss 0.0411f
C4766 vdd.n2109 vss 0.00885f
C4767 vdd.n2110 vss 0.00246f
C4768 vdd.n2111 vss 0.0307f
C4769 vdd.n2112 vss 0.00449f
C4770 vdd.n2113 vss 0.0157f
C4771 vdd.n2114 vss 0.0297f
C4772 vdd.n2115 vss 0.00885f
C4773 vdd.n2116 vss 0.00433f
C4774 vdd.n2117 vss 0.0158f
C4775 vdd.n2118 vss 0.00885f
C4776 vdd.n2119 vss 0.00433f
C4777 vdd.n2120 vss 0.0157f
C4778 vdd.n2121 vss 0.0137f
C4779 vdd.n2122 vss 0.00642f
C4780 vdd.n2123 vss 0.014f
C4781 vdd.n2124 vss 0.00538f
C4782 vdd.t48 vss 0.00542f
C4783 vdd.t47 vss 0.00542f
C4784 vdd.n2125 vss 0.0133f
C4785 vdd.n2126 vss 0.0394f
C4786 vdd.n2127 vss 0.00658f
C4787 vdd.n2128 vss 0.0134f
C4788 vdd.n2129 vss 0.125f
C4789 vdd.n2130 vss 0.371f
C4790 vdd.n2131 vss 0.0157f
C4791 vdd.n2132 vss 0.014f
C4792 vdd.n2133 vss 0.00449f
C4793 vdd.n2134 vss 0.00642f
C4794 vdd.n2135 vss 0.00804f
C4795 vdd.n2136 vss 0.0789f
C4796 vdd.n2137 vss 0.0128f
C4797 vdd.n2138 vss 8.33e-19
C4798 vdd.n2139 vss 0.0025f
C4799 vdd.n2140 vss 3.21e-19
C4800 vdd.n2141 vss 0.0516f
C4801 vdd.n2142 vss 0.0873f
C4802 vdd.n2143 vss 0.0227f
C4803 vdd.n2144 vss 0.126f
C4804 vdd.n2145 vss 0.0287f
C4805 vdd.n2146 vss 0.0168f
C4806 vdd.n2147 vss 0.00246f
C4807 vdd.n2148 vss 0.0163f
C4808 vdd.n2149 vss 0.0288f
C4809 vdd.n2150 vss 0.0158f
C4810 vdd.n2151 vss 0.00433f
C4811 vdd.n2152 vss 3.21e-19
C4812 vdd.n2153 vss 0.00286f
C4813 vdd.n2154 vss 0.00305f
C4814 vdd.n2155 vss 4.73e-19
C4815 vdd.n2156 vss 0.00839f
C4816 vdd.n2157 vss 0.014f
C4817 vdd.n2158 vss 0.107f
C4818 vdd.n2159 vss 0.106f
C4819 vdd.n2160 vss 0.0158f
C4820 vdd.n2161 vss 0.00433f
C4821 vdd.n2162 vss 0.0297f
C4822 vdd.n2163 vss 0.0307f
C4823 vdd.n2164 vss 0.0297f
C4824 vdd.n2165 vss 0.00433f
C4825 vdd.n2166 vss 0.00274f
C4826 vdd.t51 vss 0.106f
C4827 vdd.t61 vss 0.101f
C4828 vdd.n2167 vss 0.0155f
C4829 vdd.n2168 vss 0.0243f
C4830 vdd.n2169 vss 0.013f
C4831 vdd.t50 vss 0.393f
C4832 vdd.t52 vss 0.12f
C4833 vdd.t60 vss 0.393f
C4834 vdd.t9 vss 0.371f
C4835 vdd.t44 vss 0.493f
C4836 vdd.t122 vss 0.197f
C4837 vdd.t46 vss 0.244f
C4838 vdd.t56 vss 0.148f
C4839 vdd.t119 vss 0.705f
C4840 vdd.t0 vss 4.13f
C4841 vdd.t28 vss 3.12f
C4842 vdd.t19 vss 2.87f
C4843 vdd.n2170 vss 5.38f
C4844 vdd.n2171 vss 0.841f
C4845 vdd.n2172 vss 0.184f
C4846 vdd.n2174 vss 0.334f
C4847 vdd.n2175 vss 0.0163f
C4848 vdd.n2176 vss 0.0141f
C4849 vdd.n2177 vss 0.0156f
C4850 vdd.t123 vss 0.0159f
C4851 vdd.n2178 vss 0.108f
C4852 vdd.n2179 vss 0.0637f
C4853 vdd.n2180 vss 0.0732f
C4854 vdd.n2181 vss 0.0621f
C4855 vdd.n2182 vss 0.0482f
C4856 vdd.n2183 vss 0.0146f
C4857 vdd.n2184 vss 0.00286f
C4858 vdd.n2185 vss 0.00449f
C4859 vdd.n2186 vss 3.21e-19
C4860 vdd.n2187 vss 0.925f
C4861 vdd.n2188 vss 0.0147f
C4862 vdd.n2189 vss 0.00607f
C4863 vdd.t55 vss 0.0997f
C4864 vdd.t11 vss 0.0997f
C4865 vdd.t54 vss 0.0163f
C4866 vdd.t53 vss 0.0163f
C4867 vdd.n2190 vss 0.106f
C4868 vdd.t10 vss 0.0163f
C4869 vdd.t12 vss 0.0163f
C4870 vdd.n2191 vss 0.106f
C4871 vdd.n2192 vss 0.0554f
C4872 vdd.n2193 vss 0.133f
C4873 vdd.n2194 vss 0.022f
C4874 vdd.n2195 vss 0.0229f
C4875 vdd.n2196 vss 0.00683f
C4876 vdd.n2197 vss 0.0212f
C4877 vdd.n2198 vss 0.00619f
C4878 vdd.n2199 vss 0.0157f
C4879 vdd.n2200 vss 0.322f
C4880 vdd.n2201 vss 0.324f
C4881 vdd.n2202 vss 0.0163f
C4882 vdd.n2203 vss 0.00885f
C4883 vdd.n2204 vss 0.061f
C4884 vdd.n2205 vss 0.0592f
C4885 vdd.n2206 vss 0.0524f
C4886 vdd.n2207 vss 0.00459f
C4887 vdd.n2208 vss 0.022f
C4888 vdd.n2209 vss 0.0104f
C4889 vdd.n2210 vss 0.00488f
C4890 vdd.n2211 vss 0.00432f
C4891 vdd.n2212 vss 0.0633f
C4892 vdd.n2213 vss 0.0103f
C4893 vdd.n2214 vss 0.00798f
C4894 vdd.n2215 vss 0.0768f
C4895 vdd.n2216 vss 0.0329f
C4896 vdd.n2217 vss 0.0113f
C4897 vdd.n2218 vss 0.0139f
C4898 vdd.n2219 vss 0.0316f
C4899 vdd.n2220 vss 0.0659f
C4900 vdd.n2221 vss 0.0596f
C4901 vdd.n2222 vss 0.0162f
C4902 vdd.t57 vss 0.0077f
C4903 vdd.n2223 vss 0.111f
C4904 vdd.n2224 vss 0.0163f
C4905 vdd.n2225 vss 0.00891f
C4906 vdd.n2226 vss 0.0924f
C4907 vdd.n2227 vss 0.0303f
C4908 vdd.n2228 vss 0.0163f
C4909 vdd.n2229 vss 0.0641f
C4910 vdd.n2230 vss 0.00518f
C4911 vdd.n2231 vss 0.00685f
C4912 vdd.n2232 vss 0.0664f
C4913 vdd.n2233 vss 0.00661f
C4914 vdd.n2234 vss 0.0163f
C4915 vdd.n2235 vss 0.00887f
C4916 vdd.n2236 vss 0.0202f
C4917 vdd.n2237 vss 0.392f
C4918 vdd.n2238 vss 0.286f
C4919 vdd.n2239 vss 0.0303f
C4920 vdd.n2240 vss 0.0163f
C4921 vdd.n2241 vss 0.00518f
C4922 vdd.n2242 vss 0.00685f
C4923 vdd.n2243 vss 0.0664f
C4924 vdd.n2244 vss 0.00661f
C4925 vdd.n2245 vss 0.0163f
C4926 vdd.n2246 vss 0.0615f
C4927 vdd.n2247 vss 0.00887f
C4928 vdd.n2248 vss 0.0212f
C4929 vdd.n2249 vss 0.00887f
C4930 vdd.n2250 vss 0.0163f
C4931 vdd.n2251 vss 0.0116f
C4932 vdd.n2252 vss 0.00359f
C4933 vdd.n2253 vss 0.00271f
C4934 vdd.n2254 vss 0.00219f
C4935 vdd.n2255 vss 3.87e-19
C4936 vdd.n2256 vss 0.00219f
C4937 vdd.n2257 vss 0.008f
C4938 vdd.n2258 vss 0.00851f
C4939 vdd.n2259 vss 0.00219f
C4940 vdd.n2260 vss 0.00219f
C4941 vdd.n2261 vss 3.87e-19
C4942 vdd.n2262 vss 0.008f
C4943 vdd.n2263 vss 0.00271f
C4944 vdd.n2264 vss 0.00542f
C4945 vdd.n2265 vss 0.00271f
C4946 vdd.n2266 vss 0.00284f
C4947 vdd.n2267 vss 0.00658f
C4948 vdd.n2268 vss 0.00359f
C4949 vdd.n2269 vss 0.00638f
C4950 vdd.n2270 vss 0.0184f
C4951 vdd.n2271 vss -0.173f
C4952 vdd.n2272 vss 0.0113f
C4953 vdd.n2273 vss 2.66e-19
C4954 vdd.n2274 vss 3.87e-19
C4955 vdd.n2275 vss 0.00477f
C4956 vdd.n2276 vss 0.00284f
C4957 vdd.n2277 vss 0.00219f
C4958 vdd.n2278 vss 0.0105f
C4959 vdd.n2279 vss 0.008f
C4960 vdd.n2280 vss 0.00271f
C4961 vdd.n2281 vss 0.00477f
C4962 vdd.n2282 vss 0.00284f
C4963 vdd.n2283 vss 3.87e-19
C4964 vdd.n2284 vss 2.66e-19
C4965 vdd.n2285 vss 0.00399f
C4966 vdd.n2286 vss 0.0188f
C4967 vdd.n2287 vss 0.00359f
C4968 vdd.n2288 vss 0.00335f
C4969 vdd.n2289 vss 0.00284f
C4970 vdd.n2290 vss 0.00748f
C4971 vdd.n2291 vss 0.00219f
C4972 vdd.n2292 vss 0.008f
C4973 vdd.n2293 vss 0.008f
C4974 vdd.n2294 vss 0.00219f
C4975 vdd.n2296 vss 0.00226f
C4976 vdd.n2297 vss 0.00219f
C4977 vdd.n2298 vss 0.0105f
C4978 vdd.n2299 vss 0.00219f
C4979 vdd.n2300 vss 0.00219f
C4980 vdd.n2301 vss 0.00284f
C4981 vdd.n2302 vss 0.00271f
C4982 vdd.n2303 vss 0.00638f
C4983 vdd.n2304 vss 0.0116f
C4984 vdd.n2305 vss -0.0615f
C4985 vdd.n2306 vss 0.00335f
C4986 vdd.n2307 vss 0.00748f
C4987 vdd.n2308 vss 0.00219f
C4988 vdd.n2309 vss 0.00219f
C4989 vdd.n2310 vss 0.00284f
C4990 vdd.n2311 vss 0.00271f
C4991 vdd.n2312 vss 0.0233f
C4992 vdd.n2313 vss 0.0116f
C4993 vdd.n2314 vss 2.66e-19
C4994 vdd.n2315 vss 0.00271f
C4995 vdd.n2316 vss 0.00284f
C4996 vdd.n2317 vss 0.00748f
C4997 vdd.n2318 vss 0.00219f
C4998 vdd.n2319 vss 0.00219f
C4999 vdd.n2320 vss 0.024f
C5000 vdd.n2321 vss 0.00271f
C5001 vdd.n2322 vss 0.0213f
C5002 vdd.n2323 vss 0.0234f
C5003 vdd.n2324 vss 0.0234f
C5004 vdd.n2325 vss 0.0213f
C5005 vdd.n2326 vss 0.00271f
C5006 vdd.n2327 vss 0.024f
C5007 vdd.n2328 vss 0.00219f
C5008 vdd.n2329 vss 0.00851f
C5009 vdd.n2330 vss 0.00219f
C5010 vdd.n2331 vss 0.00219f
C5011 vdd.n2332 vss 0.00284f
C5012 vdd.n2333 vss 0.00335f
C5013 vdd.n2334 vss 0.00306f
C5014 vdd.n2335 vss 0.0116f
C5015 vdd.n2336 vss 2.66e-19
C5016 vdd.n2337 vss 0.00271f
C5017 vdd.n2338 vss 0.00748f
C5018 vdd.n2339 vss 0.008f
C5019 vdd.n2340 vss 0.00226f
C5020 vdd.n2341 vss 0.00219f
C5021 vdd.n2342 vss 0.00219f
C5022 vdd.n2343 vss 0.00748f
C5023 vdd.n2344 vss 3.87e-19
C5024 vdd.n2345 vss 0.008f
C5025 vdd.n2346 vss 0.00271f
C5026 vdd.n2347 vss 0.00335f
C5027 vdd.n2348 vss 0.00306f
C5028 vdd.n2349 vss -0.0689f
C5029 vdd.n2350 vss 0.00385f
C5030 vdd.n2351 vss 0.0113f
C5031 vdd.n2352 vss 0.00284f
C5032 vdd.n2353 vss 0.00219f
C5033 vdd.n2354 vss 0.00219f
C5034 vdd.n2355 vss 2.58e-19
C5035 vdd.n2356 vss 0.0105f
C5036 vdd.n2357 vss 0.00219f
C5037 vdd.n2358 vss 0.00219f
C5038 vdd.n2359 vss 0.00748f
C5039 vdd.n2360 vss 0.00284f
C5040 vdd.n2361 vss 0.00335f
C5041 vdd.n2362 vss 0.00306f
C5042 vdd.n2363 vss 2.66e-19
C5043 vdd.n2364 vss 0.0116f
C5044 vdd.n2365 vss 2.66e-19
C5045 vdd.n2366 vss 0.00271f
C5046 vdd.n2367 vss 0.00748f
C5047 vdd.n2368 vss 0.00219f
C5048 vdd.n2369 vss 0.00851f
C5049 vdd.n2370 vss 0.00219f
C5050 vdd.n2371 vss 0.00219f
C5051 vdd.n2372 vss 0.00284f
C5052 vdd.n2373 vss 0.00335f
C5053 vdd.n2374 vss 0.00306f
C5054 vdd.n2375 vss -0.0689f
C5055 vdd.n2376 vss 2.66e-19
C5056 vdd.n2377 vss 0.00271f
C5057 vdd.n2378 vss 0.0241f
C5058 vdd.n2379 vss 0.00219f
C5059 vdd.n2380 vss 0.0105f
C5060 vdd.n2381 vss 0.00219f
C5061 vdd.n2382 vss 0.00219f
C5062 vdd.n2383 vss 3.87e-19
C5063 vdd.n2384 vss 0.00271f
C5064 vdd.n2385 vss 0.00335f
C5065 vdd.n2386 vss 0.0205f
C5066 vdd.n2387 vss 0.00359f
C5067 vdd.n2388 vss 0.0197f
C5068 vdd.n2389 vss -0.148f
C5069 vdd.n2390 vss 0.00399f
C5070 vdd.n2391 vss 0.0113f
C5071 vdd.n2392 vss 2.66e-19
C5072 vdd.n2393 vss 3.87e-19
C5073 vdd.n2394 vss 0.00477f
C5074 vdd.n2395 vss 0.00284f
C5075 vdd.n2396 vss 2.58e-19
C5076 vdd.n2397 vss 0.00226f
C5077 vdd.n2398 vss 0.00219f
C5078 vdd.n2399 vss 0.00219f
C5079 vdd.n2400 vss 0.00542f
C5080 vdd.n2401 vss 0.00335f
C5081 vdd.n2402 vss -0.0615f
C5082 vdd.n2403 vss 0.00385f
C5083 vdd.n2404 vss 0.00638f
C5084 vdd.n2405 vss 0.0184f
C5085 vdd.n2406 vss 0.00638f
C5086 vdd.n2407 vss 0.00284f
C5087 vdd.n2408 vss 0.00271f
C5088 vdd.n2409 vss 0.00219f
C5089 vdd.n2410 vss 0.00748f
C5090 vdd.n2411 vss 0.00219f
C5091 vdd.n2412 vss 0.008f
C5092 vdd.n2413 vss 0.00851f
C5093 vdd.n2414 vss 0.00219f
C5094 vdd.n2415 vss 0.00219f
C5095 vdd.n2416 vss 3.87e-19
C5096 vdd.n2417 vss 0.008f
C5097 vdd.n2418 vss 0.00271f
C5098 vdd.n2419 vss 0.00542f
C5099 vdd.n2420 vss 0.00271f
C5100 vdd.n2421 vss 0.00658f
C5101 vdd.n2422 vss 0.00359f
C5102 vdd.n2423 vss -0.148f
C5103 vdd.n2424 vss 0.00399f
C5104 vdd.n2425 vss 0.0113f
C5105 vdd.n2426 vss 2.66e-19
C5106 vdd.n2427 vss 3.87e-19
C5107 vdd.n2428 vss 0.00477f
C5108 vdd.n2429 vss 0.00284f
C5109 vdd.n2430 vss 0.00219f
C5110 vdd.n2431 vss 0.0105f
C5111 vdd.n2432 vss 0.008f
C5112 vdd.n2433 vss 0.00271f
C5113 vdd.n2434 vss 0.00477f
C5114 vdd.n2435 vss 0.00284f
C5115 vdd.n2436 vss 3.87e-19
C5116 vdd.n2437 vss 2.66e-19
C5117 vdd.n2438 vss -0.173f
C5118 vdd.n2439 vss 0.0664f
C5119 vdd.n2440 vss 2.66e-19
C5120 vdd.n2441 vss 0.00271f
C5121 vdd.n2442 vss 0.00284f
C5122 vdd.n2443 vss 0.00748f
C5123 vdd.n2444 vss 0.00219f
C5124 vdd.n2445 vss 0.00219f
C5125 vdd.n2446 vss 0.024f
C5126 vdd.n2447 vss 0.0213f
C5127 vdd.n2448 vss 0.00271f
C5128 vdd.n2449 vss 0.008f
C5129 vdd.n2450 vss 0.00219f
C5130 vdd.n2452 vss 0.00226f
C5131 vdd.n2453 vss 0.0193f
C5132 vdd.n2454 vss 2.58e-19
C5133 vdd.n2455 vss 0.00219f
C5134 vdd.n2456 vss 0.00219f
C5135 vdd.n2457 vss 0.00284f
C5136 vdd.n2458 vss 0.0234f
C5137 vdd.n2459 vss 0.0234f
C5138 vdd.n2460 vss 0.0213f
C5139 vdd.n2461 vss 0.00271f
C5140 vdd.n2462 vss 0.024f
C5141 vdd.n2463 vss 0.00219f
C5142 vdd.n2464 vss 0.00851f
C5143 vdd.n2465 vss 0.00219f
C5144 vdd.n2466 vss 0.00219f
C5145 vdd.n2467 vss 0.00284f
C5146 vdd.n2468 vss 0.00335f
C5147 vdd.n2469 vss 0.00306f
C5148 vdd.n2470 vss 0.0116f
C5149 vdd.n2471 vss 2.66e-19
C5150 vdd.n2472 vss 0.00271f
C5151 vdd.n2473 vss 0.00748f
C5152 vdd.n2474 vss 0.008f
C5153 vdd.n2475 vss 0.00226f
C5154 vdd.n2476 vss 0.00219f
C5155 vdd.n2477 vss 0.00219f
C5156 vdd.n2478 vss 0.00748f
C5157 vdd.n2479 vss 3.87e-19
C5158 vdd.n2480 vss 0.008f
C5159 vdd.n2481 vss 0.00271f
C5160 vdd.n2482 vss 0.00335f
C5161 vdd.n2483 vss 0.00306f
C5162 vdd.n2484 vss -0.0689f
C5163 vdd.n2485 vss 0.00385f
C5164 vdd.n2486 vss 0.0113f
C5165 vdd.n2487 vss 0.00284f
C5166 vdd.n2488 vss 0.00219f
C5167 vdd.n2489 vss 0.00219f
C5168 vdd.n2490 vss 2.58e-19
C5169 vdd.n2491 vss 0.0105f
C5170 vdd.n2492 vss 0.00219f
C5171 vdd.n2493 vss 0.00219f
C5172 vdd.n2494 vss 0.00748f
C5173 vdd.n2495 vss 0.00284f
C5174 vdd.n2496 vss 0.00335f
C5175 vdd.n2497 vss 0.00306f
C5176 vdd.n2498 vss 2.66e-19
C5177 vdd.n2499 vss 0.0116f
C5178 vdd.n2500 vss 2.66e-19
C5179 vdd.n2501 vss 0.00271f
C5180 vdd.n2502 vss 0.00748f
C5181 vdd.n2503 vss 0.00219f
C5182 vdd.n2504 vss 0.00851f
C5183 vdd.n2505 vss 0.00219f
C5184 vdd.n2506 vss 0.00219f
C5185 vdd.n2507 vss 0.00284f
C5186 vdd.n2508 vss 0.00335f
C5187 vdd.n2509 vss 0.00306f
C5188 vdd.n2510 vss -0.0689f
C5189 vdd.n2511 vss 2.66e-19
C5190 vdd.n2512 vss 0.00271f
C5191 vdd.n2513 vss 0.0241f
C5192 vdd.n2514 vss 0.00219f
C5193 vdd.n2515 vss 0.0105f
C5194 vdd.n2516 vss 0.00219f
C5195 vdd.n2517 vss 0.00219f
C5196 vdd.n2518 vss 3.87e-19
C5197 vdd.n2519 vss 0.00271f
C5198 vdd.n2520 vss 0.00335f
C5199 vdd.n2521 vss 0.0205f
C5200 vdd.n2522 vss 0.00359f
C5201 vdd.n2523 vss 0.0197f
C5202 vdd.n2524 vss -0.148f
C5203 vdd.n2525 vss 0.00399f
C5204 vdd.n2526 vss 0.0113f
C5205 vdd.n2527 vss 2.66e-19
C5206 vdd.n2528 vss 3.87e-19
C5207 vdd.n2529 vss 0.00477f
C5208 vdd.n2530 vss 0.00284f
C5209 vdd.n2531 vss 2.58e-19
C5210 vdd.n2532 vss 0.00226f
C5211 vdd.n2533 vss 0.00219f
C5212 vdd.n2534 vss 0.00219f
C5213 vdd.n2535 vss 0.00542f
C5214 vdd.n2536 vss 0.00335f
C5215 vdd.n2537 vss -0.0615f
C5216 vdd.n2538 vss 0.00385f
C5217 vdd.n2539 vss 0.00638f
C5218 vdd.n2540 vss 0.0184f
C5219 vdd.n2541 vss 0.00638f
C5220 vdd.n2542 vss 0.00284f
C5221 vdd.n2543 vss 0.00271f
C5222 vdd.n2544 vss 0.00219f
C5223 vdd.n2545 vss 0.00748f
C5224 vdd.n2546 vss 0.00219f
C5225 vdd.n2547 vss 0.008f
C5226 vdd.n2548 vss 0.00851f
C5227 vdd.n2549 vss 0.00219f
C5228 vdd.n2550 vss 0.00219f
C5229 vdd.n2551 vss 3.87e-19
C5230 vdd.n2552 vss 0.008f
C5231 vdd.n2553 vss 0.00271f
C5232 vdd.n2554 vss 0.00542f
C5233 vdd.n2555 vss 0.00271f
C5234 vdd.n2556 vss 0.00658f
C5235 vdd.n2557 vss 0.00359f
C5236 vdd.n2558 vss -0.148f
C5237 vdd.n2559 vss 0.00399f
C5238 vdd.n2560 vss 0.0113f
C5239 vdd.n2561 vss 2.66e-19
C5240 vdd.n2562 vss 3.87e-19
C5241 vdd.n2563 vss 0.00477f
C5242 vdd.n2564 vss 0.00284f
C5243 vdd.n2565 vss 0.00219f
C5244 vdd.n2566 vss 0.0105f
C5245 vdd.n2567 vss 0.008f
C5246 vdd.n2568 vss 0.00271f
C5247 vdd.n2569 vss 0.00477f
C5248 vdd.n2570 vss 0.00284f
C5249 vdd.n2571 vss 3.87e-19
C5250 vdd.n2572 vss 2.66e-19
C5251 vdd.n2573 vss -0.173f
C5252 vdd.n2574 vss 0.0664f
C5253 vdd.n2575 vss 2.66e-19
C5254 vdd.n2576 vss 0.00271f
C5255 vdd.n2577 vss 0.00284f
C5256 vdd.n2578 vss 0.00748f
C5257 vdd.n2579 vss 0.00219f
C5258 vdd.n2580 vss 0.00219f
C5259 vdd.n2581 vss 0.024f
C5260 vdd.n2582 vss 0.0213f
C5261 vdd.n2583 vss 0.00271f
C5262 vdd.n2584 vss 0.008f
C5263 vdd.n2585 vss 0.00219f
C5264 vdd.n2587 vss 0.00226f
C5265 vdd.n2588 vss 0.0193f
C5266 vdd.n2589 vss 2.58e-19
C5267 vdd.n2590 vss 0.00219f
C5268 vdd.n2591 vss 0.00219f
C5269 vdd.n2592 vss 0.00284f
C5270 vdd.n2593 vss 0.0234f
C5271 vdd.n2594 vss 0.0234f
C5272 vdd.n2595 vss 0.0213f
C5273 vdd.n2596 vss 0.00271f
C5274 vdd.n2597 vss 0.024f
C5275 vdd.n2598 vss 0.00219f
C5276 vdd.n2599 vss 0.00851f
C5277 vdd.n2600 vss 0.00219f
C5278 vdd.n2601 vss 0.00219f
C5279 vdd.n2602 vss 0.00284f
C5280 vdd.n2603 vss 0.00335f
C5281 vdd.n2604 vss 0.00306f
C5282 vdd.n2605 vss 0.0116f
C5283 vdd.n2606 vss 2.66e-19
C5284 vdd.n2607 vss 0.00271f
C5285 vdd.n2608 vss 0.00748f
C5286 vdd.n2609 vss 0.008f
C5287 vdd.n2610 vss 0.00226f
C5288 vdd.n2611 vss 0.00219f
C5289 vdd.n2612 vss 0.00219f
C5290 vdd.n2613 vss 0.00748f
C5291 vdd.n2614 vss 3.87e-19
C5292 vdd.n2615 vss 0.008f
C5293 vdd.n2616 vss 0.00271f
C5294 vdd.n2617 vss 0.00335f
C5295 vdd.n2618 vss 0.00306f
C5296 vdd.n2619 vss -0.0689f
C5297 vdd.n2620 vss 0.00385f
C5298 vdd.n2621 vss 0.0113f
C5299 vdd.n2622 vss 0.00284f
C5300 vdd.n2623 vss 0.00219f
C5301 vdd.n2624 vss 0.00219f
C5302 vdd.n2625 vss 2.58e-19
C5303 vdd.n2626 vss 0.0105f
C5304 vdd.n2627 vss 0.00219f
C5305 vdd.n2628 vss 0.00219f
C5306 vdd.n2629 vss 0.00748f
C5307 vdd.n2630 vss 0.00284f
C5308 vdd.n2631 vss 0.00335f
C5309 vdd.n2632 vss 0.00306f
C5310 vdd.n2633 vss 2.66e-19
C5311 vdd.n2634 vss 0.0116f
C5312 vdd.n2635 vss 2.66e-19
C5313 vdd.n2636 vss 0.00271f
C5314 vdd.n2637 vss 0.00748f
C5315 vdd.n2638 vss 0.00219f
C5316 vdd.n2639 vss 0.00851f
C5317 vdd.n2640 vss 0.00219f
C5318 vdd.n2641 vss 0.00219f
C5319 vdd.n2642 vss 0.00284f
C5320 vdd.n2643 vss 0.00335f
C5321 vdd.n2644 vss 0.00306f
C5322 vdd.n2645 vss -0.0689f
C5323 vdd.n2646 vss 2.66e-19
C5324 vdd.n2647 vss 0.00271f
C5325 vdd.n2648 vss 0.0241f
C5326 vdd.n2649 vss 0.00219f
C5327 vdd.n2650 vss 0.0105f
C5328 vdd.n2651 vss 0.00219f
C5329 vdd.n2652 vss 0.00219f
C5330 vdd.n2653 vss 3.87e-19
C5331 vdd.n2654 vss 0.00271f
C5332 vdd.n2655 vss 0.00335f
C5333 vdd.n2656 vss 0.0205f
C5334 vdd.n2657 vss 0.00359f
C5335 vdd.n2658 vss 0.0197f
C5336 vdd.n2659 vss -0.148f
C5337 vdd.n2660 vss 0.00399f
C5338 vdd.n2661 vss 0.0113f
C5339 vdd.n2662 vss 2.66e-19
C5340 vdd.n2663 vss 3.87e-19
C5341 vdd.n2664 vss 0.00477f
C5342 vdd.n2665 vss 0.00284f
C5343 vdd.n2666 vss 2.58e-19
C5344 vdd.n2667 vss 0.00226f
C5345 vdd.n2668 vss 0.00219f
C5346 vdd.n2669 vss 0.00219f
C5347 vdd.n2670 vss 0.00542f
C5348 vdd.n2671 vss 0.00335f
C5349 vdd.n2672 vss -0.0615f
C5350 vdd.n2673 vss 0.00385f
C5351 vdd.n2674 vss 0.00638f
C5352 vdd.n2675 vss 0.0184f
C5353 vdd.n2676 vss 0.00638f
C5354 vdd.n2677 vss 0.00284f
C5355 vdd.n2678 vss 0.00271f
C5356 vdd.n2679 vss 0.00219f
C5357 vdd.n2680 vss 0.00748f
C5358 vdd.n2681 vss 0.00219f
C5359 vdd.n2682 vss 0.008f
C5360 vdd.n2683 vss 0.00851f
C5361 vdd.n2684 vss 0.00219f
C5362 vdd.n2685 vss 0.00219f
C5363 vdd.n2686 vss 3.87e-19
C5364 vdd.n2687 vss 0.008f
C5365 vdd.n2688 vss 0.00271f
C5366 vdd.n2689 vss 0.00542f
C5367 vdd.n2690 vss 0.00271f
C5368 vdd.n2691 vss 0.00658f
C5369 vdd.n2692 vss 0.00359f
C5370 vdd.n2693 vss -0.148f
C5371 vdd.n2694 vss 0.00399f
C5372 vdd.n2695 vss 0.0113f
C5373 vdd.n2696 vss 2.66e-19
C5374 vdd.n2697 vss 3.87e-19
C5375 vdd.n2698 vss 0.00477f
C5376 vdd.n2699 vss 0.00284f
C5377 vdd.n2700 vss 0.00219f
C5378 vdd.n2701 vss 0.0105f
C5379 vdd.n2702 vss 0.008f
C5380 vdd.n2703 vss 0.00271f
C5381 vdd.n2704 vss 0.00477f
C5382 vdd.n2705 vss 0.00284f
C5383 vdd.n2706 vss 3.87e-19
C5384 vdd.n2707 vss 2.66e-19
C5385 vdd.n2708 vss -0.173f
C5386 vdd.n2709 vss 0.0664f
C5387 vdd.n2710 vss 2.66e-19
C5388 vdd.n2711 vss 0.00271f
C5389 vdd.n2712 vss 0.00284f
C5390 vdd.n2713 vss 0.00748f
C5391 vdd.n2714 vss 0.00219f
C5392 vdd.n2715 vss 0.00219f
C5393 vdd.n2716 vss 0.024f
C5394 vdd.n2717 vss 0.0213f
C5395 vdd.n2718 vss 0.00271f
C5396 vdd.n2719 vss 0.008f
C5397 vdd.n2720 vss 0.00219f
C5398 vdd.n2722 vss 0.00226f
C5399 vdd.n2723 vss 0.0193f
C5400 vdd.n2724 vss 2.58e-19
C5401 vdd.n2725 vss 0.00219f
C5402 vdd.n2726 vss 0.00219f
C5403 vdd.n2727 vss 0.00284f
C5404 vdd.n2728 vss 0.0234f
C5405 vdd.n2729 vss 0.0234f
C5406 vdd.n2730 vss 0.0213f
C5407 vdd.n2731 vss 0.00271f
C5408 vdd.n2732 vss 0.024f
C5409 vdd.n2733 vss 0.00219f
C5410 vdd.n2734 vss 0.00851f
C5411 vdd.n2735 vss 0.00219f
C5412 vdd.n2736 vss 0.00219f
C5413 vdd.n2737 vss 0.00284f
C5414 vdd.n2738 vss 0.00335f
C5415 vdd.n2739 vss 0.00306f
C5416 vdd.n2740 vss 0.0116f
C5417 vdd.n2741 vss 2.66e-19
C5418 vdd.n2742 vss 0.00271f
C5419 vdd.n2743 vss 0.00748f
C5420 vdd.n2744 vss 0.008f
C5421 vdd.n2745 vss 0.00226f
C5422 vdd.n2746 vss 0.00219f
C5423 vdd.n2747 vss 0.00219f
C5424 vdd.n2748 vss 0.00748f
C5425 vdd.n2749 vss 3.87e-19
C5426 vdd.n2750 vss 0.008f
C5427 vdd.n2751 vss 0.00271f
C5428 vdd.n2752 vss 0.00335f
C5429 vdd.n2753 vss 0.00306f
C5430 vdd.n2754 vss -0.0689f
C5431 vdd.n2755 vss 0.00385f
C5432 vdd.n2756 vss 0.0113f
C5433 vdd.n2757 vss 0.00284f
C5434 vdd.n2758 vss 0.00219f
C5435 vdd.n2759 vss 0.00219f
C5436 vdd.n2760 vss 2.58e-19
C5437 vdd.n2761 vss 0.0105f
C5438 vdd.n2762 vss 0.00219f
C5439 vdd.n2763 vss 0.00219f
C5440 vdd.n2764 vss 0.00748f
C5441 vdd.n2765 vss 0.00284f
C5442 vdd.n2766 vss 0.00335f
C5443 vdd.n2767 vss 0.00306f
C5444 vdd.n2768 vss 2.66e-19
C5445 vdd.n2769 vss 0.0116f
C5446 vdd.n2770 vss 2.66e-19
C5447 vdd.n2771 vss 0.00271f
C5448 vdd.n2772 vss 0.00748f
C5449 vdd.n2773 vss 0.00219f
C5450 vdd.n2774 vss 0.0226f
C5451 vdd.n2775 vss 0.00219f
C5452 vdd.n2776 vss 0.00219f
C5453 vdd.n2777 vss 0.00284f
C5454 vdd.n2778 vss 0.00335f
C5455 vdd.n2779 vss 0.00306f
C5456 vdd.n2780 vss -0.0689f
C5457 vdd.n2781 vss 2.66e-19
C5458 vdd.n2782 vss 0.00271f
C5459 vdd.n2783 vss 0.0118f
C5460 vdd.n2784 vss 2.66e-19
C5461 vdd.n2785 vss 0.00271f
C5462 vdd.n2786 vss 0.0257f
C5463 vdd.n2787 vss 0.00542f
C5464 vdd.n2788 vss 0.00658f
C5465 vdd.n2789 vss 0.00306f
C5466 vdd.n2790 vss 0.0118f
C5467 vdd.n2791 vss 2.66e-19
C5468 vdd.n2792 vss 0.00271f
C5469 vdd.n2793 vss 0.00284f
C5470 vdd.n2794 vss 0.00748f
C5471 vdd.n2795 vss 0.00219f
C5472 vdd.n2796 vss 0.00219f
C5473 vdd.n2797 vss 0.00219f
C5474 vdd.n2798 vss 0.00284f
C5475 vdd.n2799 vss 0.00335f
C5476 vdd.n2800 vss 0.00306f
C5477 vdd.n2801 vss -0.0687f
C5478 vdd.n2802 vss 2.66e-19
C5479 vdd.n2803 vss 0.00271f
C5480 vdd.n2804 vss 0.00748f
C5481 vdd.n2805 vss 0.008f
C5482 vdd.n2806 vss 0.00226f
C5483 vdd.n2807 vss 0.00219f
C5484 vdd.n2808 vss 0.00219f
C5485 vdd.n2809 vss 0.00748f
C5486 vdd.n2810 vss 3.87e-19
C5487 vdd.n2811 vss 0.00271f
C5488 vdd.n2812 vss 0.00335f
C5489 vdd.n2813 vss 0.00306f
C5490 vdd.n2814 vss 0.0118f
C5491 vdd.n2815 vss -0.173f
C5492 vdd.n2816 vss 0.0191f
C5493 vdd.n2817 vss 0.0114f
C5494 vdd.n2818 vss 0.0118f
C5495 vdd.n2819 vss 2.66e-19
C5496 vdd.n2820 vss 0.00399f
C5497 vdd.n2821 vss 0.00651f
C5498 vdd.n2822 vss 0.00306f
C5499 vdd.n2823 vss 0.0187f
C5500 vdd.n2824 vss 0.0114f
C5501 vdd.n2825 vss 0.00284f
C5502 vdd.n2826 vss 0.008f
C5503 vdd.n2827 vss 0.008f
C5504 vdd.n2828 vss 0.00271f
C5505 vdd.n2829 vss 0.00542f
C5506 vdd.n2830 vss 0.00658f
C5507 vdd.n2831 vss 0.00477f
C5508 vdd.n2832 vss 0.00335f
C5509 vdd.n2833 vss 0.00271f
C5510 vdd.n2834 vss -0.0615f
C5511 vdd.n2835 vss 2.66e-19
C5512 vdd.n2836 vss 0.00399f
C5513 vdd.n2837 vss 0.00651f
C5514 vdd.n2838 vss 0.0191f
C5515 vdd.n2839 vss 0.0187f
C5516 vdd.n2840 vss 0.0114f
C5517 vdd.n2841 vss 0.00359f
C5518 vdd.n2842 vss 0.00385f
C5519 vdd.n2843 vss 0.00477f
C5520 vdd.n2844 vss 0.00542f
C5521 vdd.n2845 vss 0.00658f
C5522 vdd.n2846 vss 0.00284f
C5523 vdd.n2847 vss 0.00219f
C5524 vdd.n2848 vss 0.00284f
C5525 vdd.n2849 vss 2.58e-19
C5526 vdd.n2850 vss 0.00851f
C5527 vdd.n2851 vss 0.0105f
C5528 vdd.n2852 vss 0.008f
C5529 vdd.n2853 vss 0.00219f
C5530 vdd.n2854 vss 0.00226f
C5531 vdd.n2855 vss 0.00851f
C5532 vdd.n2856 vss 2.58e-19
C5533 vdd.n2857 vss 0.00284f
C5534 vdd.n2858 vss 3.87e-19
C5535 vdd.n2859 vss 0.00399f
C5536 vdd.n2860 vss 0.00651f
C5537 vdd.n2861 vss -0.142f
C5538 vdd.n2862 vss 0.0187f
C5539 vdd.n2863 vss 0.0114f
C5540 vdd.n2864 vss 0.00359f
C5541 vdd.n2865 vss 0.00385f
C5542 vdd.n2866 vss 0.00477f
C5543 vdd.n2867 vss 0.00658f
C5544 vdd.n2868 vss 0.00542f
C5545 vdd.n2869 vss 0.00271f
C5546 vdd.n2870 vss 0.008f
C5547 vdd.n2871 vss 0.008f
C5548 vdd.n2872 vss 0.0105f
C5549 vdd.n2873 vss 0.00226f
C5550 vdd.n2874 vss 0.00219f
C5551 vdd.n2875 vss 0.00219f
C5552 vdd.n2876 vss 0.00271f
C5553 vdd.n2877 vss 0.008f
C5554 vdd.n2878 vss 0.00226f
C5555 vdd.n2879 vss 0.00219f
C5556 vdd.n2880 vss 0.008f
C5557 vdd.n2881 vss 0.0105f
C5558 vdd.n2882 vss 0.00851f
C5559 vdd.n2883 vss 2.58e-19
C5560 vdd.n2884 vss 0.00284f
C5561 vdd.n2885 vss 3.87e-19
C5562 vdd.n2886 vss 0.00399f
C5563 vdd.n2887 vss 0.00651f
C5564 vdd.n2888 vss 0.0191f
C5565 vdd.n2889 vss 0.0187f
C5566 vdd.n2890 vss 0.0114f
C5567 vdd.n2891 vss -0.0615f
C5568 vdd.n2892 vss -0.173f
C5569 vdd.n2893 vss 0.00477f
C5570 vdd.n2894 vss 0.00335f
C5571 vdd.n2895 vss 0.00776f
C5572 vdd.n2896 vss 0.0471f
C5573 vdd.n2897 vss 0.0354f
C5574 vdd.n2898 vss 0.0358f
C5575 vdd.n2899 vss 0.114f
C5576 vdd.n2900 vss 0.0117f
C5577 vdd.n2901 vss 0.0113f
C5578 vdd.n2902 vss 0.00359f
C5579 vdd.n2903 vss 0.0325f
C5580 vdd.n2904 vss 0.0318f
C5581 vdd.n2905 vss 0.0361f
C5582 vdd.n2906 vss 0.0344f
C5583 vdd.n2907 vss 3.87e-19
C5584 vdd.n2908 vss 0.00399f
C5585 vdd.n2909 vss 0.00651f
C5586 vdd.n2910 vss -0.142f
C5587 vdd.n2911 vss 0.0184f
C5588 vdd.n2912 vss 0.0113f
C5589 vdd.n2913 vss 0.00359f
C5590 vdd.n2914 vss 0.00385f
C5591 vdd.n2915 vss 0.00477f
C5592 vdd.n2916 vss 0.00658f
C5593 vdd.n2917 vss 0.00542f
C5594 vdd.n2918 vss 0.00271f
C5595 vdd.n2919 vss 0.008f
C5596 vdd.n2920 vss 0.008f
C5597 vdd.n2921 vss 0.0105f
C5598 vdd.n2923 vss 0.00226f
C5599 vdd.n2925 vss 0.00851f
C5600 vdd.n2926 vss 2.58e-19
C5601 vdd.n2927 vss 0.00284f
C5602 vdd.n2928 vss 3.87e-19
C5603 vdd.n2929 vss 0.00399f
C5604 vdd.n2930 vss 0.00651f
C5605 vdd.n2931 vss 0.0188f
C5606 vdd.n2932 vss 0.0184f
C5607 vdd.n2933 vss 0.0113f
C5608 vdd.n2934 vss 0.00306f
C5609 vdd.n2935 vss 0.0116f
C5610 vdd.n2936 vss 0.0184f
C5611 vdd.n2937 vss 0.0188f
C5612 vdd.n2938 vss 0.00651f
C5613 vdd.n2939 vss 0.00399f
C5614 vdd.n2940 vss 0.00284f
C5615 vdd.n2941 vss 3.87e-19
C5616 vdd.n2942 vss 0.00271f
C5617 vdd.n2943 vss -0.0615f
C5618 vdd.n2944 vss -0.173f
C5619 vdd.n2945 vss 0.00477f
C5620 vdd.n2946 vss 0.00658f
C5621 vdd.n2947 vss 0.00542f
C5622 vdd.n2948 vss 0.00271f
C5623 vdd.n2949 vss 0.008f
C5624 vdd.n2950 vss 0.008f
C5625 vdd.n2951 vss 0.00219f
C5626 vdd.n2952 vss 0.00226f
C5627 vdd.n2954 vss 0.00851f
C5628 vdd.n2956 vss 0.0105f
C5629 vdd.n2957 vss 0.008f
C5630 vdd.n2958 vss 0.008f
C5631 vdd.n2959 vss 0.00271f
C5632 vdd.n2960 vss 0.00542f
C5633 vdd.n2961 vss 0.00658f
C5634 vdd.n2962 vss 0.00477f
C5635 vdd.n2963 vss 0.00335f
C5636 vdd.n2964 vss 0.00271f
C5637 vdd.n2965 vss 0.00359f
C5638 vdd.n2966 vss 2.66e-19
C5639 vdd.n2967 vss 0.00399f
C5640 vdd.n2968 vss 0.00651f
C5641 vdd.n2969 vss -0.142f
C5642 vdd.n2970 vss 0.0184f
C5643 vdd.n2971 vss 0.0113f
C5644 vdd.n2972 vss 0.00359f
C5645 vdd.n2973 vss 0.00385f
C5646 vdd.n2974 vss 0.00477f
C5647 vdd.n2975 vss 0.00542f
C5648 vdd.n2976 vss 0.00658f
C5649 vdd.n2977 vss 0.00284f
C5650 vdd.n2978 vss 0.00219f
C5651 vdd.n2979 vss 0.00284f
C5652 vdd.n2980 vss 2.58e-19
C5653 vdd.n2981 vss 0.00851f
C5654 vdd.n2983 vss 0.0105f
C5655 vdd.n2985 vss 0.00226f
C5656 vdd.n2986 vss 0.00219f
C5657 vdd.n2987 vss 2.58e-19
C5658 vdd.n2988 vss 0.00284f
C5659 vdd.n2989 vss 3.87e-19
C5660 vdd.n2990 vss 0.00399f
C5661 vdd.n2991 vss 0.00651f
C5662 vdd.n2992 vss 0.0188f
C5663 vdd.n2993 vss 0.0184f
C5664 vdd.n2994 vss 0.0116f
C5665 vdd.n2995 vss 0.0113f
C5666 vdd.n2996 vss -0.0615f
C5667 vdd.n2997 vss -0.173f
C5668 vdd.n2998 vss 0.00477f
C5669 vdd.n2999 vss 0.00658f
C5670 vdd.n3000 vss 0.00542f
C5671 vdd.n3001 vss 0.00271f
C5672 vdd.n3002 vss 0.008f
C5673 vdd.n3003 vss 0.008f
C5674 vdd.n3004 vss 0.0105f
C5675 vdd.n3006 vss 0.00226f
C5676 vdd.n3007 vss 0.0193f
C5677 vdd.n3008 vss 2.58e-19
C5678 vdd.n3009 vss 0.00284f
C5679 vdd.n3010 vss 3.87e-19
C5680 vdd.n3011 vss 0.00399f
C5681 vdd.n3012 vss 0.0234f
C5682 vdd.n3013 vss 0.00385f
C5683 vdd.n3014 vss 0.0233f
C5684 vdd.n3015 vss 0.0661f
C5685 vdd.n3016 vss 0.0113f
C5686 vdd.n3017 vss 0.0184f
C5687 vdd.n3018 vss 0.00385f
C5688 vdd.n3019 vss 0.00638f
C5689 vdd.n3020 vss 0.00319f
C5690 vdd.n3021 vss 0.0188f
C5691 vdd.n3022 vss 0.0116f
C5692 vdd.n3023 vss -0.0615f
C5693 vdd.n3024 vss 0.00271f
C5694 vdd.n3025 vss 0.00335f
C5695 vdd.n3026 vss 0.00748f
C5696 vdd.n3027 vss 0.00542f
C5697 vdd.n3028 vss 0.00658f
C5698 vdd.n3029 vss 0.00284f
C5699 vdd.n3030 vss 0.00219f
C5700 vdd.n3031 vss 0.00219f
C5701 vdd.n3032 vss 2.58e-19
C5702 vdd.n3033 vss 0.00851f
C5703 vdd.n3035 vss 0.00226f
C5704 vdd.n3037 vss 0.0105f
C5705 vdd.n3038 vss 0.008f
C5706 vdd.n3039 vss 0.008f
C5707 vdd.n3040 vss 0.00271f
C5708 vdd.n3041 vss 0.00284f
C5709 vdd.n3042 vss 0.00658f
C5710 vdd.n3043 vss 0.00542f
C5711 vdd.n3044 vss 0.00748f
C5712 vdd.n3045 vss 0.00335f
C5713 vdd.n3046 vss 0.00271f
C5714 vdd.n3047 vss 0.00359f
C5715 vdd.n3048 vss 0.0116f
C5716 vdd.n3049 vss 0.0188f
C5717 vdd.n3050 vss 0.00319f
C5718 vdd.n3051 vss 0.00638f
C5719 vdd.n3052 vss 0.00385f
C5720 vdd.n3053 vss 2.66e-19
C5721 vdd.n3054 vss -0.0637f
C5722 vdd.n3055 vss 0.0116f
C5723 vdd.n3056 vss 0.0188f
C5724 vdd.n3057 vss 0.00319f
C5725 vdd.n3058 vss 0.00399f
C5726 vdd.n3059 vss 0.00477f
C5727 vdd.n3060 vss 0.00335f
C5728 vdd.n3061 vss 0.00748f
C5729 vdd.n3062 vss 0.00284f
C5730 vdd.n3063 vss 2.58e-19
C5731 vdd.n3064 vss 0.00219f
C5732 vdd.n3065 vss 0.00226f
C5733 vdd.n3067 vss 0.0105f
C5734 vdd.n3069 vss 0.00851f
C5735 vdd.n3070 vss 2.58e-19
C5736 vdd.n3071 vss 0.00284f
C5737 vdd.n3072 vss 3.87e-19
C5738 vdd.n3073 vss 0.00385f
C5739 vdd.n3074 vss 2.66e-19
C5740 vdd.n3075 vss 0.0113f
C5741 vdd.n3076 vss 0.0116f
C5742 vdd.n3077 vss 0.0184f
C5743 vdd.n3078 vss 0.0188f
C5744 vdd.n3079 vss 0.00319f
C5745 vdd.n3080 vss -0.173f
C5746 vdd.n3081 vss 0.00477f
C5747 vdd.n3082 vss 0.00658f
C5748 vdd.n3083 vss 0.00284f
C5749 vdd.n3084 vss 0.00219f
C5750 vdd.n3085 vss 0.00271f
C5751 vdd.n3086 vss 0.008f
C5752 vdd.n3087 vss 0.008f
C5753 vdd.n3088 vss 0.0105f
C5754 vdd.n3090 vss 0.00851f
C5755 vdd.n3092 vss 0.00226f
C5756 vdd.n3093 vss 0.00219f
C5757 vdd.n3094 vss 0.008f
C5758 vdd.n3095 vss 0.008f
C5759 vdd.n3096 vss 0.00271f
C5760 vdd.n3097 vss 0.00284f
C5761 vdd.n3098 vss 0.00658f
C5762 vdd.n3099 vss 0.00542f
C5763 vdd.n3100 vss 0.00748f
C5764 vdd.n3101 vss 0.00335f
C5765 vdd.n3102 vss 0.00271f
C5766 vdd.n3103 vss 0.00359f
C5767 vdd.n3104 vss 0.0116f
C5768 vdd.n3105 vss 0.0188f
C5769 vdd.n3106 vss 0.00319f
C5770 vdd.n3107 vss 0.00638f
C5771 vdd.n3108 vss 0.00385f
C5772 vdd.n3109 vss 2.66e-19
C5773 vdd.n3110 vss -0.0637f
C5774 vdd.n3111 vss 0.0116f
C5775 vdd.n3112 vss 0.00385f
C5776 vdd.n3113 vss 0.00359f
C5777 vdd.n3114 vss 0.0113f
C5778 vdd.n3115 vss 0.0116f
C5779 vdd.n3116 vss 0.0495f
C5780 vdd.n3117 vss 0.0198f
C5781 vdd.n3118 vss 0.00399f
C5782 vdd.n3119 vss 0.0205f
C5783 vdd.n3120 vss 0.00335f
C5784 vdd.n3121 vss 0.0241f
C5785 vdd.n3122 vss 0.00284f
C5786 vdd.n3123 vss 2.58e-19
C5787 vdd.n3124 vss 0.00851f
C5788 vdd.n3126 vss 0.00226f
C5789 vdd.n3127 vss 0.0152f
C5790 vdd.n3128 vss 0.0245f
C5791 vdd.n3129 vss 0.0255f
C5792 vdd.n3130 vss 0.0142f
C5793 vdd.n3131 vss 0.00226f
C5794 vdd.n3132 vss 0.00219f
C5795 vdd.n3133 vss 2.58e-19
C5796 vdd.n3134 vss 0.00284f
C5797 vdd.n3135 vss 3.87e-19
C5798 vdd.n3136 vss 0.00399f
C5799 vdd.n3137 vss 0.00651f
C5800 vdd.n3138 vss -0.142f
C5801 vdd.n3139 vss 0.0184f
C5802 vdd.n3140 vss 0.0113f
C5803 vdd.n3141 vss 0.00359f
C5804 vdd.n3142 vss 0.00385f
C5805 vdd.n3143 vss 0.00477f
C5806 vdd.n3144 vss 0.00658f
C5807 vdd.n3145 vss 0.00542f
C5808 vdd.n3146 vss 0.00271f
C5809 vdd.n3147 vss 0.008f
C5810 vdd.n3148 vss 0.008f
C5811 vdd.n3149 vss 0.0105f
C5812 vdd.n3151 vss 0.00226f
C5813 vdd.n3153 vss 0.00851f
C5814 vdd.n3154 vss 2.58e-19
C5815 vdd.n3155 vss 0.00284f
C5816 vdd.n3156 vss 3.87e-19
C5817 vdd.n3157 vss 0.00399f
C5818 vdd.n3158 vss 0.00651f
C5819 vdd.n3159 vss 0.0188f
C5820 vdd.n3160 vss 0.0184f
C5821 vdd.n3161 vss 0.0113f
C5822 vdd.n3162 vss 0.00306f
C5823 vdd.n3163 vss 0.0116f
C5824 vdd.n3164 vss 0.0184f
C5825 vdd.n3165 vss 0.0188f
C5826 vdd.n3166 vss 0.00651f
C5827 vdd.n3167 vss 0.00399f
C5828 vdd.n3168 vss 0.00284f
C5829 vdd.n3169 vss 3.87e-19
C5830 vdd.n3170 vss 0.00271f
C5831 vdd.n3171 vss -0.0615f
C5832 vdd.n3172 vss -0.173f
C5833 vdd.n3173 vss 0.00477f
C5834 vdd.n3174 vss 0.00658f
C5835 vdd.n3175 vss 0.00542f
C5836 vdd.n3176 vss 0.00271f
C5837 vdd.n3177 vss 0.008f
C5838 vdd.n3178 vss 0.008f
C5839 vdd.n3179 vss 0.00219f
C5840 vdd.n3180 vss 0.00226f
C5841 vdd.n3182 vss 0.00851f
C5842 vdd.n3184 vss 0.0105f
C5843 vdd.n3185 vss 0.008f
C5844 vdd.n3186 vss 0.008f
C5845 vdd.n3187 vss 0.00271f
C5846 vdd.n3188 vss 0.00542f
C5847 vdd.n3189 vss 0.00658f
C5848 vdd.n3190 vss 0.00477f
C5849 vdd.n3191 vss 0.00335f
C5850 vdd.n3192 vss 0.00271f
C5851 vdd.n3193 vss 0.00359f
C5852 vdd.n3194 vss 2.66e-19
C5853 vdd.n3195 vss 0.00399f
C5854 vdd.n3196 vss 0.00651f
C5855 vdd.n3197 vss -0.142f
C5856 vdd.n3198 vss 0.0184f
C5857 vdd.n3199 vss 0.0113f
C5858 vdd.n3200 vss 0.00359f
C5859 vdd.n3201 vss 0.00385f
C5860 vdd.n3202 vss 0.00477f
C5861 vdd.n3203 vss 0.00542f
C5862 vdd.n3204 vss 0.00658f
C5863 vdd.n3205 vss 0.00284f
C5864 vdd.n3206 vss 0.00219f
C5865 vdd.n3207 vss 0.00284f
C5866 vdd.n3208 vss 2.58e-19
C5867 vdd.n3209 vss 0.00851f
C5868 vdd.n3211 vss 0.0105f
C5869 vdd.n3213 vss 0.00226f
C5870 vdd.n3214 vss 0.00219f
C5871 vdd.n3215 vss 2.58e-19
C5872 vdd.n3216 vss 0.00284f
C5873 vdd.n3217 vss 3.87e-19
C5874 vdd.n3218 vss 0.00399f
C5875 vdd.n3219 vss 0.00651f
C5876 vdd.n3220 vss 0.0188f
C5877 vdd.n3221 vss 0.0184f
C5878 vdd.n3222 vss 0.0116f
C5879 vdd.n3223 vss 0.0113f
C5880 vdd.n3224 vss -0.0615f
C5881 vdd.n3225 vss -0.173f
C5882 vdd.n3226 vss 0.00477f
C5883 vdd.n3227 vss 0.00658f
C5884 vdd.n3228 vss 0.00542f
C5885 vdd.n3229 vss 0.00271f
C5886 vdd.n3230 vss 0.008f
C5887 vdd.n3231 vss 0.008f
C5888 vdd.n3232 vss 0.0105f
C5889 vdd.n3234 vss 0.00226f
C5890 vdd.n3235 vss 0.0193f
C5891 vdd.n3236 vss 2.58e-19
C5892 vdd.n3237 vss 0.00284f
C5893 vdd.n3238 vss 3.87e-19
C5894 vdd.n3239 vss 0.00399f
C5895 vdd.n3240 vss 0.0234f
C5896 vdd.n3241 vss 0.00385f
C5897 vdd.n3242 vss 0.0233f
C5898 vdd.n3243 vss 0.0661f
C5899 vdd.n3244 vss 0.0113f
C5900 vdd.n3245 vss 0.0184f
C5901 vdd.n3246 vss 0.00385f
C5902 vdd.n3247 vss 0.00638f
C5903 vdd.n3248 vss 0.00319f
C5904 vdd.n3249 vss 0.0188f
C5905 vdd.n3250 vss 0.0116f
C5906 vdd.n3251 vss -0.0615f
C5907 vdd.n3252 vss 0.00271f
C5908 vdd.n3253 vss 0.00335f
C5909 vdd.n3254 vss 0.00748f
C5910 vdd.n3255 vss 0.00542f
C5911 vdd.n3256 vss 0.00658f
C5912 vdd.n3257 vss 0.00284f
C5913 vdd.n3258 vss 0.00219f
C5914 vdd.n3259 vss 0.00219f
C5915 vdd.n3260 vss 2.58e-19
C5916 vdd.n3261 vss 0.00851f
C5917 vdd.n3263 vss 0.00226f
C5918 vdd.n3265 vss 0.0105f
C5919 vdd.n3266 vss 0.008f
C5920 vdd.n3267 vss 0.008f
C5921 vdd.n3268 vss 0.00271f
C5922 vdd.n3269 vss 0.00284f
C5923 vdd.n3270 vss 0.00658f
C5924 vdd.n3271 vss 0.00542f
C5925 vdd.n3272 vss 0.00748f
C5926 vdd.n3273 vss 0.00335f
C5927 vdd.n3274 vss 0.00271f
C5928 vdd.n3275 vss 0.00359f
C5929 vdd.n3276 vss 0.0116f
C5930 vdd.n3277 vss 0.0188f
C5931 vdd.n3278 vss 0.00319f
C5932 vdd.n3279 vss 0.00638f
C5933 vdd.n3280 vss 0.00385f
C5934 vdd.n3281 vss 2.66e-19
C5935 vdd.n3282 vss -0.0637f
C5936 vdd.n3283 vss 0.0116f
C5937 vdd.n3284 vss 0.0188f
C5938 vdd.n3285 vss 0.00319f
C5939 vdd.n3286 vss 0.00399f
C5940 vdd.n3287 vss 0.00477f
C5941 vdd.n3288 vss 0.00335f
C5942 vdd.n3289 vss 0.00748f
C5943 vdd.n3290 vss 0.00284f
C5944 vdd.n3291 vss 2.58e-19
C5945 vdd.n3292 vss 0.00219f
C5946 vdd.n3293 vss 0.00226f
C5947 vdd.n3295 vss 0.0105f
C5948 vdd.n3297 vss 0.00851f
C5949 vdd.n3298 vss 2.58e-19
C5950 vdd.n3299 vss 0.00284f
C5951 vdd.n3300 vss 3.87e-19
C5952 vdd.n3301 vss 0.00385f
C5953 vdd.n3302 vss 2.66e-19
C5954 vdd.n3303 vss 0.0113f
C5955 vdd.n3304 vss 0.0116f
C5956 vdd.n3305 vss 0.0184f
C5957 vdd.n3306 vss 0.0188f
C5958 vdd.n3307 vss 0.00319f
C5959 vdd.n3308 vss -0.173f
C5960 vdd.n3309 vss 0.00477f
C5961 vdd.n3310 vss 0.00658f
C5962 vdd.n3311 vss 0.00284f
C5963 vdd.n3312 vss 0.00219f
C5964 vdd.n3313 vss 0.00271f
C5965 vdd.n3314 vss 0.008f
C5966 vdd.n3315 vss 0.008f
C5967 vdd.n3316 vss 0.0105f
C5968 vdd.n3318 vss 0.00851f
C5969 vdd.n3320 vss 0.00226f
C5970 vdd.n3321 vss 0.00219f
C5971 vdd.n3322 vss 0.008f
C5972 vdd.n3323 vss 0.008f
C5973 vdd.n3324 vss 0.00271f
C5974 vdd.n3325 vss 0.00284f
C5975 vdd.n3326 vss 0.00658f
C5976 vdd.n3327 vss 0.00542f
C5977 vdd.n3328 vss 0.00748f
C5978 vdd.n3329 vss 0.00335f
C5979 vdd.n3330 vss 0.00271f
C5980 vdd.n3331 vss 0.00359f
C5981 vdd.n3332 vss 0.0116f
C5982 vdd.n3333 vss 0.0188f
C5983 vdd.n3334 vss 0.00319f
C5984 vdd.n3335 vss 0.00638f
C5985 vdd.n3336 vss 0.00385f
C5986 vdd.n3337 vss 2.66e-19
C5987 vdd.n3338 vss -0.0637f
C5988 vdd.n3339 vss 0.0116f
C5989 vdd.n3340 vss 0.00385f
C5990 vdd.n3341 vss 0.00359f
C5991 vdd.n3342 vss 0.0113f
C5992 vdd.n3343 vss 0.0116f
C5993 vdd.n3344 vss 0.0495f
C5994 vdd.n3345 vss 0.0198f
C5995 vdd.n3346 vss 0.00399f
C5996 vdd.n3347 vss 0.0205f
C5997 vdd.n3348 vss 0.00335f
C5998 vdd.n3349 vss 0.0241f
C5999 vdd.n3350 vss 0.00284f
C6000 vdd.n3351 vss 2.58e-19
C6001 vdd.n3352 vss 0.00851f
C6002 vdd.n3354 vss 0.00226f
C6003 vdd.n3355 vss 0.0152f
C6004 vdd.n3356 vss 0.0245f
C6005 vdd.n3357 vss 0.0255f
C6006 vdd.n3358 vss 0.0142f
C6007 vdd.n3359 vss 0.00226f
C6008 vdd.n3360 vss 0.00219f
C6009 vdd.n3361 vss 2.58e-19
C6010 vdd.n3362 vss 0.00284f
C6011 vdd.n3363 vss 3.87e-19
C6012 vdd.n3364 vss 0.00399f
C6013 vdd.n3365 vss 0.00651f
C6014 vdd.n3366 vss -0.142f
C6015 vdd.n3367 vss 0.0184f
C6016 vdd.n3368 vss 0.0113f
C6017 vdd.n3369 vss 0.00359f
C6018 vdd.n3370 vss 0.00385f
C6019 vdd.n3371 vss 0.00477f
C6020 vdd.n3372 vss 0.00658f
C6021 vdd.n3373 vss 0.00542f
C6022 vdd.n3374 vss 0.00271f
C6023 vdd.n3375 vss 0.008f
C6024 vdd.n3376 vss 0.008f
C6025 vdd.n3377 vss 0.0105f
C6026 vdd.n3379 vss 0.00226f
C6027 vdd.n3381 vss 0.00851f
C6028 vdd.n3382 vss 2.58e-19
C6029 vdd.n3383 vss 0.00284f
C6030 vdd.n3384 vss 3.87e-19
C6031 vdd.n3385 vss 0.00399f
C6032 vdd.n3386 vss 0.00651f
C6033 vdd.n3387 vss 0.0188f
C6034 vdd.n3388 vss 0.0184f
C6035 vdd.n3389 vss 0.0113f
C6036 vdd.n3390 vss 0.00306f
C6037 vdd.n3391 vss 0.0116f
C6038 vdd.n3392 vss 0.0184f
C6039 vdd.n3393 vss 0.0188f
C6040 vdd.n3394 vss 0.00651f
C6041 vdd.n3395 vss 0.00399f
C6042 vdd.n3396 vss 0.00284f
C6043 vdd.n3397 vss 3.87e-19
C6044 vdd.n3398 vss 0.00271f
C6045 vdd.n3399 vss -0.0615f
C6046 vdd.n3400 vss -0.173f
C6047 vdd.n3401 vss 0.00477f
C6048 vdd.n3402 vss 0.00658f
C6049 vdd.n3403 vss 0.00542f
C6050 vdd.n3404 vss 0.00271f
C6051 vdd.n3405 vss 0.008f
C6052 vdd.n3406 vss 0.008f
C6053 vdd.n3407 vss 0.00219f
C6054 vdd.n3408 vss 0.00226f
C6055 vdd.n3410 vss 0.00851f
C6056 vdd.n3412 vss 0.0105f
C6057 vdd.n3413 vss 0.008f
C6058 vdd.n3414 vss 0.008f
C6059 vdd.n3415 vss 0.00271f
C6060 vdd.n3416 vss 0.00542f
C6061 vdd.n3417 vss 0.00658f
C6062 vdd.n3418 vss 0.00477f
C6063 vdd.n3419 vss 0.00335f
C6064 vdd.n3420 vss 0.00271f
C6065 vdd.n3421 vss 0.00359f
C6066 vdd.n3422 vss 2.66e-19
C6067 vdd.n3423 vss 0.00399f
C6068 vdd.n3424 vss 0.00651f
C6069 vdd.n3425 vss -0.142f
C6070 vdd.n3426 vss 0.0184f
C6071 vdd.n3427 vss 0.0113f
C6072 vdd.n3428 vss 0.00359f
C6073 vdd.n3429 vss 0.00385f
C6074 vdd.n3430 vss 0.00477f
C6075 vdd.n3431 vss 0.00542f
C6076 vdd.n3432 vss 0.00658f
C6077 vdd.n3433 vss 0.00284f
C6078 vdd.n3434 vss 0.00219f
C6079 vdd.n3435 vss 0.00284f
C6080 vdd.n3436 vss 2.58e-19
C6081 vdd.n3437 vss 0.00851f
C6082 vdd.n3439 vss 0.0105f
C6083 vdd.n3441 vss 0.00226f
C6084 vdd.n3442 vss 0.00219f
C6085 vdd.n3443 vss 2.58e-19
C6086 vdd.n3444 vss 0.00284f
C6087 vdd.n3445 vss 3.87e-19
C6088 vdd.n3446 vss 0.00399f
C6089 vdd.n3447 vss 0.00651f
C6090 vdd.n3448 vss 0.0188f
C6091 vdd.n3449 vss 0.0184f
C6092 vdd.n3450 vss 0.0116f
C6093 vdd.n3451 vss 0.0113f
C6094 vdd.n3452 vss -0.0615f
C6095 vdd.n3453 vss -0.173f
C6096 vdd.n3454 vss 0.00477f
C6097 vdd.n3455 vss 0.00658f
C6098 vdd.n3456 vss 0.00542f
C6099 vdd.n3457 vss 0.00271f
C6100 vdd.n3458 vss 0.008f
C6101 vdd.n3459 vss 0.008f
C6102 vdd.n3460 vss 0.0105f
C6103 vdd.n3462 vss 0.00226f
C6104 vdd.n3463 vss 0.0193f
C6105 vdd.n3464 vss 2.58e-19
C6106 vdd.n3465 vss 0.00284f
C6107 vdd.n3466 vss 3.87e-19
C6108 vdd.n3467 vss 0.00399f
C6109 vdd.n3468 vss 0.0234f
C6110 vdd.n3469 vss 0.00385f
C6111 vdd.n3470 vss 0.0233f
C6112 vdd.n3471 vss 0.0661f
C6113 vdd.n3472 vss 0.0113f
C6114 vdd.n3473 vss 0.0184f
C6115 vdd.n3474 vss 0.00385f
C6116 vdd.n3475 vss 0.00638f
C6117 vdd.n3476 vss 0.00319f
C6118 vdd.n3477 vss 0.0188f
C6119 vdd.n3478 vss 0.0116f
C6120 vdd.n3479 vss -0.0615f
C6121 vdd.n3480 vss 0.00271f
C6122 vdd.n3481 vss 0.00335f
C6123 vdd.n3482 vss 0.00748f
C6124 vdd.n3483 vss 0.00542f
C6125 vdd.n3484 vss 0.00658f
C6126 vdd.n3485 vss 0.00284f
C6127 vdd.n3486 vss 0.00219f
C6128 vdd.n3487 vss 0.00219f
C6129 vdd.n3488 vss 2.58e-19
C6130 vdd.n3489 vss 0.00851f
C6131 vdd.n3491 vss 0.00226f
C6132 vdd.n3493 vss 0.0105f
C6133 vdd.n3494 vss 0.008f
C6134 vdd.n3495 vss 0.008f
C6135 vdd.n3496 vss 0.00271f
C6136 vdd.n3497 vss 0.00284f
C6137 vdd.n3498 vss 0.00658f
C6138 vdd.n3499 vss 0.00542f
C6139 vdd.n3500 vss 0.00748f
C6140 vdd.n3501 vss 0.00335f
C6141 vdd.n3502 vss 0.00271f
C6142 vdd.n3503 vss 0.00359f
C6143 vdd.n3504 vss 0.0116f
C6144 vdd.n3505 vss 0.0188f
C6145 vdd.n3506 vss 0.00319f
C6146 vdd.n3507 vss 0.00638f
C6147 vdd.n3508 vss 0.00385f
C6148 vdd.n3509 vss 2.66e-19
C6149 vdd.n3510 vss -0.0637f
C6150 vdd.n3511 vss 0.0116f
C6151 vdd.n3512 vss 0.0188f
C6152 vdd.n3513 vss 0.00319f
C6153 vdd.n3514 vss 0.00399f
C6154 vdd.n3515 vss 0.00477f
C6155 vdd.n3516 vss 0.00335f
C6156 vdd.n3517 vss 0.00748f
C6157 vdd.n3518 vss 0.00284f
C6158 vdd.n3519 vss 2.58e-19
C6159 vdd.n3520 vss 0.00219f
C6160 vdd.n3521 vss 0.00226f
C6161 vdd.n3523 vss 0.0105f
C6162 vdd.n3525 vss 0.00851f
C6163 vdd.n3526 vss 2.58e-19
C6164 vdd.n3527 vss 0.00284f
C6165 vdd.n3528 vss 3.87e-19
C6166 vdd.n3529 vss 0.00385f
C6167 vdd.n3530 vss 2.66e-19
C6168 vdd.n3531 vss 0.0113f
C6169 vdd.n3532 vss 0.0116f
C6170 vdd.n3533 vss 0.0184f
C6171 vdd.n3534 vss 0.0188f
C6172 vdd.n3535 vss 0.00319f
C6173 vdd.n3536 vss -0.173f
C6174 vdd.n3537 vss 0.00477f
C6175 vdd.n3538 vss 0.00658f
C6176 vdd.n3539 vss 0.00284f
C6177 vdd.n3540 vss 0.00219f
C6178 vdd.n3541 vss 0.00271f
C6179 vdd.n3542 vss 0.008f
C6180 vdd.n3543 vss 0.008f
C6181 vdd.n3544 vss 0.0105f
C6182 vdd.n3546 vss 0.00851f
C6183 vdd.n3548 vss 0.00226f
C6184 vdd.n3549 vss 0.00219f
C6185 vdd.n3550 vss 0.008f
C6186 vdd.n3551 vss 0.008f
C6187 vdd.n3552 vss 0.00271f
C6188 vdd.n3553 vss 0.00284f
C6189 vdd.n3554 vss 0.00658f
C6190 vdd.n3555 vss 0.00542f
C6191 vdd.n3556 vss 0.00748f
C6192 vdd.n3557 vss 0.00335f
C6193 vdd.n3558 vss 0.00271f
C6194 vdd.n3559 vss 0.00359f
C6195 vdd.n3560 vss 0.0116f
C6196 vdd.n3561 vss 0.0188f
C6197 vdd.n3562 vss 0.00319f
C6198 vdd.n3563 vss 0.00638f
C6199 vdd.n3564 vss 0.00385f
C6200 vdd.n3565 vss 2.66e-19
C6201 vdd.n3566 vss -0.0637f
C6202 vdd.n3567 vss 0.0116f
C6203 vdd.n3568 vss 0.00385f
C6204 vdd.n3569 vss 0.00359f
C6205 vdd.n3570 vss 0.0113f
C6206 vdd.n3571 vss 0.0116f
C6207 vdd.n3572 vss 0.0495f
C6208 vdd.n3573 vss 0.0198f
C6209 vdd.n3574 vss 0.00399f
C6210 vdd.n3575 vss 0.0205f
C6211 vdd.n3576 vss 0.00335f
C6212 vdd.n3577 vss 0.0241f
C6213 vdd.n3578 vss 0.00284f
C6214 vdd.n3579 vss 2.58e-19
C6215 vdd.n3580 vss 0.00851f
C6216 vdd.n3582 vss 0.00226f
C6217 vdd.n3583 vss 0.0152f
C6218 vdd.n3584 vss 0.0245f
C6219 vdd.n3585 vss 0.0255f
C6220 vdd.n3586 vss 0.0142f
C6221 vdd.n3587 vss 0.00226f
C6222 vdd.n3588 vss 0.00219f
C6223 vdd.n3589 vss 2.58e-19
C6224 vdd.n3590 vss 0.00284f
C6225 vdd.n3591 vss 3.87e-19
C6226 vdd.n3592 vss 0.00399f
C6227 vdd.n3593 vss 0.00651f
C6228 vdd.n3594 vss -0.142f
C6229 vdd.n3595 vss 0.0184f
C6230 vdd.n3596 vss 0.0113f
C6231 vdd.n3597 vss 0.00359f
C6232 vdd.n3598 vss 0.00385f
C6233 vdd.n3599 vss 0.00477f
C6234 vdd.n3600 vss 0.00658f
C6235 vdd.n3601 vss 0.00542f
C6236 vdd.n3602 vss 0.00271f
C6237 vdd.n3603 vss 0.008f
C6238 vdd.n3604 vss 0.008f
C6239 vdd.n3605 vss 0.0105f
C6240 vdd.n3607 vss 0.00226f
C6241 vdd.n3609 vss 0.00851f
C6242 vdd.n3610 vss 2.58e-19
C6243 vdd.n3611 vss 0.00284f
C6244 vdd.n3612 vss 3.87e-19
C6245 vdd.n3613 vss 0.00399f
C6246 vdd.n3614 vss 0.00651f
C6247 vdd.n3615 vss 0.0188f
C6248 vdd.n3616 vss 0.0184f
C6249 vdd.n3617 vss 0.0113f
C6250 vdd.n3618 vss 0.00306f
C6251 vdd.n3619 vss 0.0116f
C6252 vdd.n3620 vss 0.0184f
C6253 vdd.n3621 vss 0.0188f
C6254 vdd.n3622 vss 0.00651f
C6255 vdd.n3623 vss 0.00399f
C6256 vdd.n3624 vss 0.00284f
C6257 vdd.n3625 vss 3.87e-19
C6258 vdd.n3626 vss 0.00271f
C6259 vdd.n3627 vss -0.0615f
C6260 vdd.n3628 vss -0.173f
C6261 vdd.n3629 vss 0.00477f
C6262 vdd.n3630 vss 0.00658f
C6263 vdd.n3631 vss 0.00542f
C6264 vdd.n3632 vss 0.00271f
C6265 vdd.n3633 vss 0.008f
C6266 vdd.n3634 vss 0.008f
C6267 vdd.n3635 vss 0.00219f
C6268 vdd.n3636 vss 0.00226f
C6269 vdd.n3638 vss 0.00851f
C6270 vdd.n3640 vss 0.0105f
C6271 vdd.n3641 vss 0.008f
C6272 vdd.n3642 vss 0.008f
C6273 vdd.n3643 vss 0.00271f
C6274 vdd.n3644 vss 0.00542f
C6275 vdd.n3645 vss 0.00658f
C6276 vdd.n3646 vss 0.00477f
C6277 vdd.n3647 vss 0.00335f
C6278 vdd.n3648 vss 0.00271f
C6279 vdd.n3649 vss 0.00359f
C6280 vdd.n3650 vss 2.66e-19
C6281 vdd.n3651 vss 0.00399f
C6282 vdd.n3652 vss 0.00651f
C6283 vdd.n3653 vss -0.142f
C6284 vdd.n3654 vss 0.0184f
C6285 vdd.n3655 vss 0.0113f
C6286 vdd.n3656 vss 0.00359f
C6287 vdd.n3657 vss 0.00385f
C6288 vdd.n3658 vss 0.00477f
C6289 vdd.n3659 vss 0.00542f
C6290 vdd.n3660 vss 0.00658f
C6291 vdd.n3661 vss 0.00284f
C6292 vdd.n3662 vss 0.00219f
C6293 vdd.n3663 vss 0.00284f
C6294 vdd.n3664 vss 2.58e-19
C6295 vdd.n3665 vss 0.00851f
C6296 vdd.n3667 vss 0.0105f
C6297 vdd.n3669 vss 0.00226f
C6298 vdd.n3670 vss 0.00219f
C6299 vdd.n3671 vss 2.58e-19
C6300 vdd.n3672 vss 0.00284f
C6301 vdd.n3673 vss 3.87e-19
C6302 vdd.n3674 vss 0.00399f
C6303 vdd.n3675 vss 0.00651f
C6304 vdd.n3676 vss 0.0188f
C6305 vdd.n3677 vss 0.0184f
C6306 vdd.n3678 vss 0.0113f
C6307 vdd.n3679 vss -0.0615f
C6308 vdd.n3680 vss -0.173f
C6309 vdd.n3681 vss 0.00477f
C6310 vdd.n3682 vss 0.00658f
C6311 vdd.n3683 vss 0.00542f
C6312 vdd.n3684 vss 0.00271f
C6313 vdd.n3685 vss 0.008f
C6314 vdd.n3686 vss 0.008f
C6315 vdd.n3687 vss 0.0105f
C6316 vdd.n3689 vss 0.00226f
C6317 vdd.n3690 vss 0.0193f
C6318 vdd.n3691 vss 2.58e-19
C6319 vdd.n3692 vss 0.00284f
C6320 vdd.n3693 vss 3.87e-19
C6321 vdd.n3694 vss 0.00399f
C6322 vdd.n3695 vss 0.0234f
C6323 vdd.n3696 vss 0.0664f
C6324 vdd.n3697 vss 0.0661f
C6325 vdd.n3698 vss 0.0113f
C6326 vdd.n3699 vss 2.66e-19
C6327 vdd.n3700 vss 0.00385f
C6328 vdd.n3701 vss 3.87e-19
C6329 vdd.n3702 vss 0.00284f
C6330 vdd.n3703 vss 2.58e-19
C6331 vdd.n3704 vss 0.0193f
C6332 vdd.n3706 vss 0.00226f
C6333 vdd.n3707 vss 0.00219f
C6334 vdd.n3708 vss 0.008f
C6335 vdd.n3709 vss 0.008f
C6336 vdd.n3710 vss 0.00271f
C6337 vdd.n3711 vss 0.00542f
C6338 vdd.n3712 vss 0.00658f
C6339 vdd.n3713 vss 0.00477f
C6340 vdd.n3714 vss -0.173f
C6341 vdd.n3715 vss 0.00319f
C6342 vdd.n3716 vss 0.0188f
C6343 vdd.n3717 vss 0.0184f
C6344 vdd.n3718 vss 0.0116f
C6345 vdd.n3719 vss 0.0113f
C6346 vdd.n3720 vss 2.66e-19
C6347 vdd.n3721 vss 0.00385f
C6348 vdd.n3722 vss 3.87e-19
C6349 vdd.n3723 vss 0.00284f
C6350 vdd.n3724 vss 2.58e-19
C6351 vdd.n3725 vss 0.00851f
C6352 vdd.n3727 vss 0.00226f
C6353 vdd.n3728 vss 0.0105f
C6354 vdd.n3730 vss 0.00851f
C6355 vdd.n3731 vss 2.58e-19
C6356 vdd.n3732 vss 0.00219f
C6357 vdd.n3733 vss 0.008f
C6358 vdd.n3734 vss 0.00271f
C6359 vdd.n3735 vss 0.00542f
C6360 vdd.n3736 vss 0.00658f
C6361 vdd.n3737 vss 0.00477f
C6362 vdd.n3738 vss 0.00399f
C6363 vdd.n3739 vss 0.00319f
C6364 vdd.n3740 vss 0.00385f
C6365 vdd.n3741 vss 0.00638f
C6366 vdd.n3742 vss -0.148f
C6367 vdd.n3743 vss -0.0637f
C6368 vdd.n3744 vss 0.0184f
C6369 vdd.n3745 vss 0.00385f
C6370 vdd.n3746 vss 0.00638f
C6371 vdd.n3747 vss 0.00319f
C6372 vdd.n3748 vss 0.0188f
C6373 vdd.n3749 vss 0.0116f
C6374 vdd.n3750 vss 0.00359f
C6375 vdd.n3751 vss 0.00271f
C6376 vdd.n3752 vss 0.00335f
C6377 vdd.n3753 vss 0.00748f
C6378 vdd.n3754 vss 0.00542f
C6379 vdd.n3755 vss 0.00658f
C6380 vdd.n3756 vss 0.00284f
C6381 vdd.n3757 vss 0.00219f
C6382 vdd.n3758 vss 0.00219f
C6383 vdd.n3759 vss 2.58e-19
C6384 vdd.n3760 vss 0.00851f
C6385 vdd.n3762 vss 0.00226f
C6386 vdd.n3764 vss 0.0105f
C6387 vdd.n3765 vss 0.008f
C6388 vdd.n3766 vss 0.008f
C6389 vdd.n3767 vss 0.00271f
C6390 vdd.n3768 vss 0.00284f
C6391 vdd.n3769 vss 0.00658f
C6392 vdd.n3770 vss 0.00542f
C6393 vdd.n3771 vss 0.00748f
C6394 vdd.n3772 vss 0.00335f
C6395 vdd.n3773 vss 0.00271f
C6396 vdd.n3774 vss -0.0615f
C6397 vdd.n3775 vss 0.0116f
C6398 vdd.n3776 vss 0.0188f
C6399 vdd.n3777 vss 0.00319f
C6400 vdd.n3778 vss 0.00638f
C6401 vdd.n3779 vss 0.00385f
C6402 vdd.n3780 vss 2.66e-19
C6403 vdd.n3781 vss 0.0113f
C6404 vdd.n3782 vss 0.0116f
C6405 vdd.n3783 vss 0.00385f
C6406 vdd.n3784 vss 2.66e-19
C6407 vdd.n3785 vss -0.0637f
C6408 vdd.n3786 vss -0.148f
C6409 vdd.n3787 vss 0.0188f
C6410 vdd.n3788 vss 0.00319f
C6411 vdd.n3789 vss 0.00399f
C6412 vdd.n3790 vss 0.00477f
C6413 vdd.n3791 vss 0.00335f
C6414 vdd.n3792 vss 0.00748f
C6415 vdd.n3793 vss 0.00284f
C6416 vdd.n3794 vss 2.58e-19
C6417 vdd.n3795 vss 0.00219f
C6418 vdd.n3796 vss 0.00226f
C6419 vdd.n3798 vss 0.0105f
C6420 vdd.n3799 vss 0.0226f
C6421 vdd.n3800 vss 0.0361f
C6422 vdd.n3801 vss 0.0344f
C6423 vdd.n3802 vss 0.0318f
C6424 vdd.n3803 vss 0.0325f
C6425 vdd.n3804 vss 0.0496f
C6426 vdd.n3805 vss 0.14f
C6427 vdd.n3806 vss 0.00518f
C6428 vdd.n3807 vss 0.00661f
C6429 vdd.n3808 vss 0.0664f
C6430 vdd.n3809 vss 0.0068f
C6431 vdd.n3810 vss 0.0163f
C6432 vdd.n3811 vss 0.0303f
C6433 vdd.n3812 vss 0.0391f
C6434 vdd.n3813 vss 0.173f
C6435 vdd.n3814 vss 0.428f
C6436 vdd.n3815 vss 0.0163f
C6437 vdd.n3816 vss 0.0361f
C6438 vdd.n3817 vss 0.0163f
C6439 vdd.n3818 vss 0.00661f
C6440 vdd.n3819 vss 0.0664f
C6441 vdd.t3 vss 0.367f
C6442 vdd.n3820 vss 0.199f
C6443 vdd.n3821 vss 0.397f
C6444 vdd.n3822 vss 0.391f
C6445 vdd.n3823 vss 0.0664f
C6446 vdd.n3824 vss 0.00661f
C6447 vdd.n3825 vss 0.0163f
C6448 vdd.n3826 vss 0.00887f
C6449 vdd.n3827 vss 0.0706f
C6450 vdd.n3828 vss 0.0706f
C6451 vdd.n3829 vss 0.0163f
C6452 vdd.n3830 vss 0.0303f
C6453 vdd.n3831 vss 0.0163f
C6454 vdd.n3832 vss 0.00661f
C6455 vdd.n3833 vss 0.0664f
C6456 vdd.n3834 vss 0.178f
C6457 vdd.n3835 vss 0.342f
C6458 vdd.n3836 vss 0.392f
C6459 vdd.t108 vss 0.244f
C6460 vdd.n3837 vss 0.0114f
C6461 vdd.n3838 vss 0.00864f
C6462 vdd.t109 vss 0.0416f
C6463 vdd.n3839 vss 0.0169f
C6464 vdd.n3840 vss 6.66e-19
C6465 vdd.n3841 vss 0.0101f
C6466 vdd.n3842 vss 0.0151f
C6467 vdd.n3843 vss 0.00563f
C6468 vdd.n3844 vss 0.0152f
C6469 vdd.n3845 vss 0.00564f
C6470 vdd.n3846 vss 0.00362f
C6471 vdd.n3847 vss 0.0972f
C6472 vdd.n3848 vss 0.013f
C6473 vdd.n3849 vss 0.0139f
C6474 vdd.n3850 vss 0.0334f
C6475 vdd.n3851 vss 0.0189f
C6476 vdd.n3852 vss 0.00563f
C6477 vdd.n3853 vss 0.0158f
C6478 vdd.t131 vss 0.0416f
C6479 vdd.n3854 vss 0.0454f
C6480 vdd.n3855 vss 0.00651f
C6481 vdd.n3856 vss 0.00209f
C6482 vdd.n3857 vss 0.00394f
C6483 vdd.n3858 vss 0.00886f
C6484 vdd.n3859 vss 0.00338f
C6485 vdd.n3860 vss 0.00619f
C6486 vdd.n3861 vss 0.00318f
C6487 vdd.n3862 vss 0.00376f
C6488 vdd.n3863 vss 0.00319f
C6489 vdd.n3864 vss 0.0015f
C6490 vdd.n3865 vss 0.00111f
C6491 vdd.n3866 vss 0.00209f
C6492 vdd.n3867 vss 0.0166f
C6493 vdd.n3868 vss 0.00133f
C6494 vdd.t130 vss 0.224f
C6495 vdd.t20 vss 0.392f
C6496 vdd.n3869 vss 0.0568f
C6497 vdd.n3870 vss 0.0664f
C6498 vdd.n3871 vss 0.00685f
C6499 vdd.n3872 vss 0.00518f
C6500 vdd.n3873 vss 0.00887f
C6501 vdd.n3874 vss 0.0373f
C6502 vdd.n3875 vss 0.0163f
C6503 vdd.n3876 vss 0.00685f
C6504 vdd.n3877 vss 0.00518f
C6505 vdd.n3878 vss 0.00661f
C6506 vdd.n3879 vss 0.0163f
C6507 vdd.n3880 vss 0.0373f
C6508 vdd.n3881 vss 0.0163f
C6509 vdd.n3882 vss 0.00518f
C6510 vdd.n3883 vss 0.00685f
C6511 vdd.n3884 vss 0.0664f
C6512 vdd.n3885 vss 0.00661f
C6513 vdd.n3886 vss 0.0163f
C6514 vdd.n3887 vss 0.0374f
C6515 vdd.n3888 vss 0.0162f
C6516 vdd.t101 vss 0.0077f
C6517 vdd.n3889 vss 0.111f
C6518 vdd.n3890 vss 0.0163f
C6519 vdd.n3891 vss 0.0157f
C6520 vdd.n3892 vss 0.0137f
C6521 vdd.n3893 vss 0.00642f
C6522 vdd.n3894 vss 0.014f
C6523 vdd.n3895 vss 0.00538f
C6524 vdd.t27 vss 0.00542f
C6525 vdd.t21 vss 0.00542f
C6526 vdd.n3896 vss 0.0133f
C6527 vdd.n3897 vss 0.0394f
C6528 vdd.n3898 vss 0.00658f
C6529 vdd.n3899 vss 0.0134f
C6530 vdd.n3900 vss 0.0793f
C6531 vdd.n3901 vss 0.0947f
C6532 vdd.n3902 vss 0.00887f
C6533 vdd.n3903 vss 0.132f
C6534 vdd.n3904 vss 0.132f
C6535 vdd.n3905 vss 0.00887f
C6536 vdd.n3906 vss 0.0789f
C6537 vdd.n3907 vss 0.0789f
C6538 vdd.n3908 vss 0.00887f
C6539 vdd.n3909 vss 0.087f
C6540 vdd.n3910 vss 0.087f
C6541 vdd.n3911 vss 0.0373f
C6542 vdd.n3912 vss 0.0163f
C6543 vdd.n3913 vss 0.0373f
C6544 vdd.n3914 vss 0.0163f
C6545 vdd.n3915 vss 0.00518f
C6546 vdd.n3916 vss 0.00685f
C6547 vdd.n3917 vss 0.043f
C6548 vdd.n3918 vss 0.00226f
C6549 vdd.n3919 vss 0.0341f
C6550 vdd.n3920 vss 0.0147f
C6551 vdd.n3921 vss 0.337f
C6552 vdd.t100 vss 0.453f
C6553 vdd.t25 vss 0.252f
C6554 vdd.n3922 vss 0.108f
C6555 vdd.n3923 vss 0.122f
C6556 vdd.n3924 vss 0.0664f
C6557 vdd.n3925 vss 0.00661f
C6558 vdd.n3926 vss 0.0163f
C6559 vdd.n3927 vss 0.00887f
C6560 vdd.n3928 vss 0.0709f
C6561 vdd.n3929 vss 0.0709f
C6562 vdd.n3930 vss 0.00518f
C6563 vdd.n3931 vss 0.00685f
C6564 vdd.n3932 vss 0.0664f
C6565 vdd.n3933 vss 0.00661f
C6566 vdd.n3934 vss 0.0163f
C6567 vdd.n3935 vss 0.00887f
C6568 vdd.n3936 vss 0.0758f
C6569 vdd.n3937 vss 0.0758f
C6570 vdd.n3938 vss 0.0163f
C6571 vdd.n3939 vss 0.0373f
C6572 vdd.n3940 vss 0.0163f
C6573 vdd.n3941 vss 0.00661f
C6574 vdd.n3942 vss 0.0664f
C6575 vdd.n3943 vss 0.176f
C6576 vdd.n3944 vss 0.0769f
C6577 vdd.n3945 vss 0.136f
C6578 vdd.n3946 vss 0.452f
C6579 vdd.n3947 vss 0.0664f
C6580 vdd.n3948 vss 0.0664f
C6581 vdd.n3949 vss 0.00685f
C6582 vdd.n3950 vss 0.00518f
C6583 vdd.n3951 vss 0.00887f
C6584 vdd.n3952 vss 0.049f
C6585 vdd.n3953 vss 0.0163f
C6586 vdd.n3954 vss 0.00685f
C6587 vdd.n3955 vss 0.00518f
C6588 vdd.n3956 vss 0.00661f
C6589 vdd.n3957 vss 0.0163f
C6590 vdd.n3958 vss 0.049f
C6591 vdd.n3959 vss 0.0163f
C6592 vdd.n3960 vss 0.00685f
C6593 vdd.n3961 vss 0.00518f
C6594 vdd.n3962 vss 0.00661f
C6595 vdd.n3963 vss 0.0163f
C6596 vdd.n3964 vss 0.00887f
C6597 vdd.n3965 vss 0.136f
C6598 vdd.n3966 vss 0.136f
C6599 vdd.n3967 vss 0.00887f
C6600 vdd.n3968 vss 0.118f
C6601 vdd.n3969 vss 0.118f
C6602 vdd.n3970 vss 0.0997f
C6603 vdd.n3971 vss 0.0163f
C6604 vdd.n3972 vss 0.049f
C6605 vdd.n3973 vss 0.0163f
C6606 vdd.n3974 vss 0.00661f
C6607 vdd.n3975 vss 0.0664f
C6608 vdd.n3976 vss 0.242f
C6609 vdd.n3977 vss 0.027f
C6610 vdd.n3978 vss 0.017f
C6611 vdd.n3979 vss 0.0322f
C6612 vdd.n3980 vss 0.163f
C6613 vdd.n3981 vss 0.0102f
C6614 vdd.n3982 vss 0.00888f
C6615 vdd.n3983 vss 0.00814f
C6616 vdd.n3984 vss 0.0214f
C6617 vdd.n3985 vss 0.0141f
C6618 vdd.n3986 vss 0.0161f
C6619 vdd.n3987 vss 6.66e-19
C6620 vdd.n3988 vss 0.0101f
C6621 vdd.n3989 vss 0.0735f
C6622 vdd.n3990 vss 0.00327f
C6623 vdd.n3991 vss 0.0101f
C6624 vdd.n3992 vss 0.00903f
C6625 vdd.n3993 vss 0.00466f
C6626 vdd.n3994 vss 0.0163f
C6627 vdd.n3995 vss 0.0213f
C6628 vdd.n3996 vss 0.0493f
C6629 vdd.n3997 vss 0.0224f
C6630 vdd.n3998 vss 0.0162f
C6631 vdd.n3999 vss 0.0173f
C6632 vdd.n4000 vss 0.019f
C6633 vdd.n4001 vss 0.0458f
C6634 vdd.n4002 vss 0.00651f
C6635 vdd.n4003 vss 0.0256f
C6636 vdd.n4004 vss 0.201f
C6637 vdd.n4005 vss 1.68f
C6638 vdd.t22 vss 1.62f
C6639 vdd.n4006 vss 1.56f
C6640 vdd.t23 vss 1.9f
C6641 vdd.t29 vss 1.6f
C6642 vdd.n4007 vss 0.916f
C6643 vdd.n4008 vss 0.0522f
C6644 vdd.n4009 vss 0.00219f
C6645 vdd.t24 vss 0.00477f
C6646 vdd.n4010 vss 0.0469f
C6647 vdd.n4011 vss 0.0295f
C6648 vdd.n4012 vss 0.0129f
C6649 vdd.n4013 vss 3.87e-19
C6650 vdd.n4014 vss 0.0105f
C6651 vdd.n4015 vss 0.008f
C6652 vdd.n4016 vss 0.008f
C6653 vdd.n4017 vss 0.00271f
C6654 vdd.n4018 vss 0.00284f
C6655 vdd.n4019 vss 0.00219f
C6656 vdd.n4020 vss 0.00284f
C6657 vdd.n4021 vss 2.58e-19
C6658 vdd.n4022 vss 0.00247f
C6659 vdd.n4023 vss 0.00811f
C6660 vdd.n4024 vss 0.0142f
C6661 vdd.n4025 vss 0.113f
C6662 vdd.n4027 vss 0.00851f
C6663 vdd.n4028 vss 2.58e-19
C6664 vdd.n4029 vss 0.00284f
C6665 vdd.n4030 vss 0.00748f
C6666 vdd.n4031 vss 0.00335f
C6667 vdd.n4032 vss 0.00477f
C6668 vdd.n4033 vss 0.00385f
C6669 vdd.n4034 vss 0.00306f
C6670 vdd.n4035 vss 0.00651f
C6671 vdd.n4036 vss -0.142f
C6672 vdd.n4037 vss -0.0687f
C6673 vdd.n4038 vss 0.0114f
C6674 vdd.n4039 vss 0.00359f
C6675 vdd.n4040 vss 0.00385f
C6676 vdd.n4041 vss 0.00637f
C6677 vdd.n4042 vss 0.00994f
C6678 vdd.n4043 vss 0.00504f
C6679 vdd.n4044 vss 0.00908f
C6680 vdd.n4045 vss 8.67e-19
C6681 vdd.n4046 vss 0.0927f
C6682 vdd.n4047 vss 0.27f
C6683 vdd.n4048 vss 0.213f
C6684 vdd.n4049 vss 0.0318f
C6685 vdd.n4050 vss 0.0325f
C6686 vdd.n4051 vss 0.0496f
C6687 vdd.n4052 vss 0.0116f
C6688 vdd.n4053 vss -0.0637f
C6689 vdd.n4054 vss 2.66e-19
C6690 vdd.n4055 vss 0.00385f
C6691 vdd.n4056 vss 3.87e-19
C6692 vdd.n4057 vss 0.00284f
C6693 vdd.n4058 vss 0.00219f
C6694 vdd.n4059 vss 0.00271f
C6695 vdd.n4060 vss 0.008f
C6696 vdd.n4061 vss 0.008f
C6697 vdd.n4062 vss 0.0105f
C6698 vdd.n4063 vss 0.2f
C6699 vdd.n4064 vss 0.043f
C6700 vdd.n4065 vss 0.162f
C6701 vdd.n4066 vss 0.00851f
C6702 vdd.n4067 vss 2.58e-19
C6703 vdd.n4068 vss 0.00284f
C6704 vdd.n4069 vss 3.87e-19
C6705 vdd.n4070 vss 0.00385f
C6706 vdd.n4071 vss 0.00638f
C6707 vdd.n4072 vss 0.00319f
C6708 vdd.n4073 vss 0.0188f
C6709 vdd.n4074 vss 0.0116f
C6710 vdd.n4075 vss 0.0113f
C6711 vdd.n4076 vss 2.66e-19
C6712 vdd.n4077 vss 0.00385f
C6713 vdd.n4078 vss 3.87e-19
C6714 vdd.n4079 vss 0.00284f
C6715 vdd.n4080 vss 0.00219f
C6716 vdd.n4081 vss 0.00271f
C6717 vdd.n4082 vss 0.008f
C6718 vdd.n4083 vss 0.008f
C6719 vdd.n4084 vss 0.0105f
C6720 vdd.n4085 vss 0.2f
C6721 vdd.n4086 vss 0.043f
C6722 vdd.n4087 vss 0.162f
C6723 vdd.n4088 vss 0.00851f
C6724 vdd.n4089 vss 2.58e-19
C6725 vdd.n4090 vss 0.00284f
C6726 vdd.n4091 vss 3.87e-19
C6727 vdd.n4092 vss 0.00385f
C6728 vdd.n4093 vss 0.00638f
C6729 vdd.n4094 vss 0.00319f
C6730 vdd.n4095 vss 0.0188f
C6731 vdd.n4096 vss 0.0116f
C6732 vdd.n4097 vss 0.0113f
C6733 vdd.n4098 vss 2.66e-19
C6734 vdd.n4099 vss 0.00385f
C6735 vdd.n4100 vss 3.87e-19
C6736 vdd.n4101 vss 0.00284f
C6737 vdd.n4102 vss 0.00219f
C6738 vdd.n4103 vss 0.00271f
C6739 vdd.n4104 vss 0.008f
C6740 vdd.n4105 vss 0.008f
C6741 vdd.n4106 vss 0.0105f
C6742 vdd.n4107 vss 0.2f
C6743 vdd.n4108 vss 0.043f
C6744 vdd.n4109 vss 0.101f
C6745 vdd.n4110 vss 0.0193f
C6746 vdd.n4111 vss 2.58e-19
C6747 vdd.n4112 vss 0.00284f
C6748 vdd.n4113 vss 3.87e-19
C6749 vdd.n4114 vss 0.00385f
C6750 vdd.n4115 vss 0.0233f
C6751 vdd.n4116 vss 0.0234f
C6752 vdd.n4117 vss 0.0664f
C6753 vdd.n4118 vss 0.0116f
C6754 vdd.n4119 vss 0.0113f
C6755 vdd.n4120 vss -0.0615f
C6756 vdd.n4121 vss 0.00271f
C6757 vdd.n4122 vss 0.00335f
C6758 vdd.n4123 vss 0.00748f
C6759 vdd.n4124 vss 0.00542f
C6760 vdd.n4125 vss 0.00658f
C6761 vdd.n4126 vss 0.00284f
C6762 vdd.n4127 vss 0.00219f
C6763 vdd.n4128 vss 0.00284f
C6764 vdd.n4129 vss 2.58e-19
C6765 vdd.n4130 vss 0.00219f
C6766 vdd.n4131 vss 0.00226f
C6767 vdd.n4132 vss 0.043f
C6768 vdd.n4133 vss 0.2f
C6769 vdd.n4134 vss 0.162f
C6770 vdd.n4135 vss 0.00851f
C6771 vdd.n4136 vss 2.58e-19
C6772 vdd.n4137 vss 0.00284f
C6773 vdd.n4138 vss 0.00748f
C6774 vdd.n4139 vss 0.00335f
C6775 vdd.n4140 vss 0.00477f
C6776 vdd.n4141 vss 0.00385f
C6777 vdd.n4142 vss 0.00306f
C6778 vdd.n4143 vss 0.00651f
C6779 vdd.n4144 vss 0.0188f
C6780 vdd.n4145 vss 0.0116f
C6781 vdd.n4146 vss 0.0113f
C6782 vdd.n4147 vss -0.0615f
C6783 vdd.n4148 vss 0.00271f
C6784 vdd.n4149 vss 0.00335f
C6785 vdd.n4150 vss 0.00748f
C6786 vdd.n4151 vss 0.00542f
C6787 vdd.n4152 vss 0.00658f
C6788 vdd.n4153 vss 0.00284f
C6789 vdd.n4154 vss 0.00219f
C6790 vdd.n4155 vss 0.00284f
C6791 vdd.n4156 vss 2.58e-19
C6792 vdd.n4157 vss 0.00219f
C6793 vdd.n4158 vss 0.00226f
C6794 vdd.n4159 vss 0.043f
C6795 vdd.n4160 vss 0.2f
C6796 vdd.n4161 vss 0.162f
C6797 vdd.n4162 vss 0.00851f
C6798 vdd.n4163 vss 2.58e-19
C6799 vdd.n4164 vss 0.00284f
C6800 vdd.n4165 vss 3.87e-19
C6801 vdd.n4166 vss 0.00271f
C6802 vdd.n4167 vss 0.00359f
C6803 vdd.n4168 vss 0.0113f
C6804 vdd.n4169 vss 0.0116f
C6805 vdd.n4170 vss 0.0197f
C6806 vdd.n4171 vss 0.0198f
C6807 vdd.n4172 vss 0.0495f
C6808 vdd.n4173 vss 0.0116f
C6809 vdd.n4174 vss -0.0637f
C6810 vdd.n4175 vss 2.66e-19
C6811 vdd.n4176 vss 0.00385f
C6812 vdd.n4177 vss 3.87e-19
C6813 vdd.n4178 vss 0.00284f
C6814 vdd.n4179 vss 0.00219f
C6815 vdd.n4180 vss 0.00271f
C6816 vdd.n4181 vss 0.008f
C6817 vdd.n4182 vss 0.008f
C6818 vdd.n4183 vss 0.0105f
C6819 vdd.n4184 vss 0.2f
C6820 vdd.n4185 vss 0.043f
C6821 vdd.n4186 vss 0.162f
C6822 vdd.n4187 vss 0.00851f
C6823 vdd.n4188 vss 2.58e-19
C6824 vdd.n4189 vss 0.00284f
C6825 vdd.n4190 vss 3.87e-19
C6826 vdd.n4191 vss 0.00385f
C6827 vdd.n4192 vss 0.00638f
C6828 vdd.n4193 vss 0.00319f
C6829 vdd.n4194 vss 0.0188f
C6830 vdd.n4195 vss 0.0116f
C6831 vdd.n4196 vss 0.0113f
C6832 vdd.n4197 vss 2.66e-19
C6833 vdd.n4198 vss 0.00385f
C6834 vdd.n4199 vss 3.87e-19
C6835 vdd.n4200 vss 0.00284f
C6836 vdd.n4201 vss 0.00219f
C6837 vdd.n4202 vss 0.00271f
C6838 vdd.n4203 vss 0.008f
C6839 vdd.n4204 vss 0.008f
C6840 vdd.n4205 vss 0.0105f
C6841 vdd.n4206 vss 0.2f
C6842 vdd.n4207 vss 0.043f
C6843 vdd.n4208 vss 0.162f
C6844 vdd.n4209 vss 0.00851f
C6845 vdd.n4210 vss 2.58e-19
C6846 vdd.n4211 vss 0.00284f
C6847 vdd.n4212 vss 3.87e-19
C6848 vdd.n4213 vss 0.00385f
C6849 vdd.n4214 vss 0.00638f
C6850 vdd.n4215 vss 0.00319f
C6851 vdd.n4216 vss 0.0188f
C6852 vdd.n4217 vss 0.0116f
C6853 vdd.n4218 vss 0.0113f
C6854 vdd.n4219 vss 2.66e-19
C6855 vdd.n4220 vss 0.00385f
C6856 vdd.n4221 vss 3.87e-19
C6857 vdd.n4222 vss 0.00284f
C6858 vdd.n4223 vss 0.00219f
C6859 vdd.n4224 vss 0.00271f
C6860 vdd.n4225 vss 0.008f
C6861 vdd.n4226 vss 0.008f
C6862 vdd.n4227 vss 0.0105f
C6863 vdd.n4228 vss 0.2f
C6864 vdd.n4229 vss 0.043f
C6865 vdd.n4230 vss 0.101f
C6866 vdd.n4231 vss 0.0193f
C6867 vdd.n4232 vss 2.58e-19
C6868 vdd.n4233 vss 0.00284f
C6869 vdd.n4234 vss 3.87e-19
C6870 vdd.n4235 vss 0.00385f
C6871 vdd.n4236 vss 0.0233f
C6872 vdd.n4237 vss 0.0234f
C6873 vdd.n4238 vss 0.0664f
C6874 vdd.n4239 vss 0.0116f
C6875 vdd.n4240 vss 0.0113f
C6876 vdd.n4241 vss -0.0615f
C6877 vdd.n4242 vss 0.00271f
C6878 vdd.n4243 vss 0.00335f
C6879 vdd.n4244 vss 0.00748f
C6880 vdd.n4245 vss 0.00542f
C6881 vdd.n4246 vss 0.00658f
C6882 vdd.n4247 vss 0.00284f
C6883 vdd.n4248 vss 0.00219f
C6884 vdd.n4249 vss 0.00284f
C6885 vdd.n4250 vss 2.58e-19
C6886 vdd.n4251 vss 0.00219f
C6887 vdd.n4252 vss 0.00226f
C6888 vdd.n4253 vss 0.043f
C6889 vdd.n4254 vss 0.2f
C6890 vdd.n4255 vss 0.162f
C6891 vdd.n4256 vss 0.00851f
C6892 vdd.n4257 vss 2.58e-19
C6893 vdd.n4258 vss 0.00284f
C6894 vdd.n4259 vss 0.00748f
C6895 vdd.n4260 vss 0.00335f
C6896 vdd.n4261 vss 0.00477f
C6897 vdd.n4262 vss 0.00385f
C6898 vdd.n4263 vss 0.00306f
C6899 vdd.n4264 vss 0.00651f
C6900 vdd.n4265 vss 0.0188f
C6901 vdd.n4266 vss 0.0116f
C6902 vdd.n4267 vss 0.0113f
C6903 vdd.n4268 vss -0.0615f
C6904 vdd.n4269 vss 0.00271f
C6905 vdd.n4270 vss 0.00335f
C6906 vdd.n4271 vss 0.00748f
C6907 vdd.n4272 vss 0.00542f
C6908 vdd.n4273 vss 0.00658f
C6909 vdd.n4274 vss 0.00284f
C6910 vdd.n4275 vss 0.00219f
C6911 vdd.n4276 vss 0.00284f
C6912 vdd.n4277 vss 2.58e-19
C6913 vdd.n4278 vss 0.00219f
C6914 vdd.n4279 vss 0.00226f
C6915 vdd.n4280 vss 0.043f
C6916 vdd.n4281 vss 0.2f
C6917 vdd.n4282 vss 0.162f
C6918 vdd.n4283 vss 0.00851f
C6919 vdd.n4284 vss 2.58e-19
C6920 vdd.n4285 vss 0.00284f
C6921 vdd.n4286 vss 3.87e-19
C6922 vdd.n4287 vss 0.00271f
C6923 vdd.n4288 vss 0.00359f
C6924 vdd.n4289 vss 0.0113f
C6925 vdd.n4290 vss 0.0116f
C6926 vdd.n4291 vss 0.0197f
C6927 vdd.n4292 vss 0.0198f
C6928 vdd.n4293 vss 0.0495f
C6929 vdd.n4294 vss 0.0116f
C6930 vdd.n4295 vss -0.0637f
C6931 vdd.n4296 vss 2.66e-19
C6932 vdd.n4297 vss 0.00385f
C6933 vdd.n4298 vss 3.87e-19
C6934 vdd.n4299 vss 0.00284f
C6935 vdd.n4300 vss 0.00219f
C6936 vdd.n4301 vss 0.00271f
C6937 vdd.n4302 vss 0.008f
C6938 vdd.n4303 vss 0.008f
C6939 vdd.n4304 vss 0.0105f
C6940 vdd.n4305 vss 0.2f
C6941 vdd.n4306 vss 0.043f
C6942 vdd.n4307 vss 0.162f
C6943 vdd.n4308 vss 0.00851f
C6944 vdd.n4309 vss 2.58e-19
C6945 vdd.n4310 vss 0.00284f
C6946 vdd.n4311 vss 3.87e-19
C6947 vdd.n4312 vss 0.00385f
C6948 vdd.n4313 vss 0.00638f
C6949 vdd.n4314 vss 0.00319f
C6950 vdd.n4315 vss 0.0188f
C6951 vdd.n4316 vss 0.0116f
C6952 vdd.n4317 vss 0.0113f
C6953 vdd.n4318 vss 2.66e-19
C6954 vdd.n4319 vss 0.00385f
C6955 vdd.n4320 vss 3.87e-19
C6956 vdd.n4321 vss 0.00284f
C6957 vdd.n4322 vss 0.00219f
C6958 vdd.n4323 vss 0.00271f
C6959 vdd.n4324 vss 0.008f
C6960 vdd.n4325 vss 0.008f
C6961 vdd.n4326 vss 0.0105f
C6962 vdd.n4327 vss 0.2f
C6963 vdd.n4328 vss 0.043f
C6964 vdd.n4329 vss 0.162f
C6965 vdd.n4330 vss 0.00851f
C6966 vdd.n4331 vss 2.58e-19
C6967 vdd.n4332 vss 0.00284f
C6968 vdd.n4333 vss 3.87e-19
C6969 vdd.n4334 vss 0.00385f
C6970 vdd.n4335 vss 0.00638f
C6971 vdd.n4336 vss 0.00319f
C6972 vdd.n4337 vss 0.0188f
C6973 vdd.n4338 vss 0.0116f
C6974 vdd.n4339 vss 0.0113f
C6975 vdd.n4340 vss 2.66e-19
C6976 vdd.n4341 vss 0.00385f
C6977 vdd.n4342 vss 3.87e-19
C6978 vdd.n4343 vss 0.00284f
C6979 vdd.n4344 vss 0.00219f
C6980 vdd.n4345 vss 0.00271f
C6981 vdd.n4346 vss 0.008f
C6982 vdd.n4347 vss 0.008f
C6983 vdd.n4348 vss 0.0105f
C6984 vdd.n4349 vss 0.2f
C6985 vdd.n4350 vss 0.043f
C6986 vdd.n4351 vss 0.101f
C6987 vdd.n4352 vss 0.0193f
C6988 vdd.n4353 vss 2.58e-19
C6989 vdd.n4354 vss 0.00284f
C6990 vdd.n4355 vss 3.87e-19
C6991 vdd.n4356 vss 0.00385f
C6992 vdd.n4357 vss 0.0233f
C6993 vdd.n4358 vss 0.0234f
C6994 vdd.n4359 vss 0.0664f
C6995 vdd.n4360 vss 0.0116f
C6996 vdd.n4361 vss 0.0113f
C6997 vdd.n4362 vss -0.0615f
C6998 vdd.n4363 vss 0.00271f
C6999 vdd.n4364 vss 0.00335f
C7000 vdd.n4365 vss 0.00748f
C7001 vdd.n4366 vss 0.00542f
C7002 vdd.n4367 vss 0.00658f
C7003 vdd.n4368 vss 0.00284f
C7004 vdd.n4369 vss 0.00219f
C7005 vdd.n4370 vss 0.00284f
C7006 vdd.n4371 vss 2.58e-19
C7007 vdd.n4372 vss 0.00219f
C7008 vdd.n4373 vss 0.00226f
C7009 vdd.n4374 vss 0.043f
C7010 vdd.n4375 vss 0.2f
C7011 vdd.n4376 vss 0.162f
C7012 vdd.n4377 vss 0.00851f
C7013 vdd.n4378 vss 2.58e-19
C7014 vdd.n4379 vss 0.00284f
C7015 vdd.n4380 vss 0.00748f
C7016 vdd.n4381 vss 0.00335f
C7017 vdd.n4382 vss 0.00477f
C7018 vdd.n4383 vss 0.00385f
C7019 vdd.n4384 vss 0.00306f
C7020 vdd.n4385 vss 0.00651f
C7021 vdd.n4386 vss 0.0188f
C7022 vdd.n4387 vss 0.0116f
C7023 vdd.n4388 vss 0.0113f
C7024 vdd.n4389 vss -0.0615f
C7025 vdd.n4390 vss 0.00271f
C7026 vdd.n4391 vss 0.00335f
C7027 vdd.n4392 vss 0.00748f
C7028 vdd.n4393 vss 0.00542f
C7029 vdd.n4394 vss 0.00658f
C7030 vdd.n4395 vss 0.00284f
C7031 vdd.n4396 vss 0.00219f
C7032 vdd.n4397 vss 0.00284f
C7033 vdd.n4398 vss 2.58e-19
C7034 vdd.n4399 vss 0.00219f
C7035 vdd.n4400 vss 0.00226f
C7036 vdd.n4401 vss 0.043f
C7037 vdd.n4402 vss 0.2f
C7038 vdd.n4403 vss 0.162f
C7039 vdd.n4404 vss 0.00851f
C7040 vdd.n4405 vss 2.58e-19
C7041 vdd.n4406 vss 0.00284f
C7042 vdd.n4407 vss 3.87e-19
C7043 vdd.n4408 vss 0.00271f
C7044 vdd.n4409 vss 0.00359f
C7045 vdd.n4410 vss 0.0113f
C7046 vdd.n4411 vss 0.0116f
C7047 vdd.n4412 vss 0.0197f
C7048 vdd.n4413 vss 0.0198f
C7049 vdd.n4414 vss 0.0495f
C7050 vdd.n4415 vss 0.0116f
C7051 vdd.n4416 vss -0.0637f
C7052 vdd.n4417 vss 2.66e-19
C7053 vdd.n4418 vss 0.00385f
C7054 vdd.n4419 vss 3.87e-19
C7055 vdd.n4420 vss 0.00284f
C7056 vdd.n4421 vss 0.00219f
C7057 vdd.n4422 vss 0.00271f
C7058 vdd.n4423 vss 0.008f
C7059 vdd.n4424 vss 0.008f
C7060 vdd.n4425 vss 0.0105f
C7061 vdd.n4426 vss 0.2f
C7062 vdd.n4427 vss 0.043f
C7063 vdd.n4428 vss 0.162f
C7064 vdd.n4429 vss 0.00851f
C7065 vdd.n4430 vss 2.58e-19
C7066 vdd.n4431 vss 0.00284f
C7067 vdd.n4432 vss 3.87e-19
C7068 vdd.n4433 vss 0.00385f
C7069 vdd.n4434 vss 0.00638f
C7070 vdd.n4435 vss 0.00319f
C7071 vdd.n4436 vss 0.0188f
C7072 vdd.n4437 vss 0.0116f
C7073 vdd.n4438 vss 0.0113f
C7074 vdd.n4439 vss 2.66e-19
C7075 vdd.n4440 vss 0.00385f
C7076 vdd.n4441 vss 3.87e-19
C7077 vdd.n4442 vss 0.00284f
C7078 vdd.n4443 vss 0.00219f
C7079 vdd.n4444 vss 0.00271f
C7080 vdd.n4445 vss 0.008f
C7081 vdd.n4446 vss 0.008f
C7082 vdd.n4447 vss 0.0105f
C7083 vdd.n4448 vss 0.2f
C7084 vdd.n4449 vss 0.043f
C7085 vdd.n4450 vss 0.162f
C7086 vdd.n4451 vss 0.00851f
C7087 vdd.n4452 vss 2.58e-19
C7088 vdd.n4453 vss 0.00284f
C7089 vdd.n4454 vss 3.87e-19
C7090 vdd.n4455 vss 0.00385f
C7091 vdd.n4456 vss 0.00638f
C7092 vdd.n4457 vss 0.00319f
C7093 vdd.n4458 vss 0.0188f
C7094 vdd.n4459 vss 0.0116f
C7095 vdd.n4460 vss 0.0113f
C7096 vdd.n4461 vss 2.66e-19
C7097 vdd.n4462 vss 0.00385f
C7098 vdd.n4463 vss 3.87e-19
C7099 vdd.n4464 vss 0.00284f
C7100 vdd.n4465 vss 0.00219f
C7101 vdd.n4466 vss 0.00271f
C7102 vdd.n4467 vss 0.008f
C7103 vdd.n4468 vss 0.008f
C7104 vdd.n4469 vss 0.0105f
C7105 vdd.n4470 vss 0.2f
C7106 vdd.n4471 vss 0.043f
C7107 vdd.n4472 vss 0.101f
C7108 vdd.n4473 vss 0.0193f
C7109 vdd.n4474 vss 2.58e-19
C7110 vdd.n4475 vss 0.00284f
C7111 vdd.n4476 vss 3.87e-19
C7112 vdd.n4477 vss 0.00385f
C7113 vdd.n4478 vss 0.0233f
C7114 vdd.n4479 vss 0.0234f
C7115 vdd.n4480 vss 0.0664f
C7116 vdd.n4481 vss 0.0116f
C7117 vdd.n4482 vss 0.0113f
C7118 vdd.n4483 vss -0.0615f
C7119 vdd.n4484 vss 0.00271f
C7120 vdd.n4485 vss 0.00335f
C7121 vdd.n4486 vss 0.00748f
C7122 vdd.n4487 vss 0.00542f
C7123 vdd.n4488 vss 0.00658f
C7124 vdd.n4489 vss 0.00284f
C7125 vdd.n4490 vss 0.00219f
C7126 vdd.n4491 vss 0.00284f
C7127 vdd.n4492 vss 2.58e-19
C7128 vdd.n4493 vss 0.00219f
C7129 vdd.n4494 vss 0.00226f
C7130 vdd.n4495 vss 0.043f
C7131 vdd.n4496 vss 0.2f
C7132 vdd.n4497 vss 0.162f
C7133 vdd.n4498 vss 0.00851f
C7134 vdd.n4499 vss 2.58e-19
C7135 vdd.n4500 vss 0.00284f
C7136 vdd.n4501 vss 0.00748f
C7137 vdd.n4502 vss 0.00335f
C7138 vdd.n4503 vss 0.00477f
C7139 vdd.n4504 vss 0.00385f
C7140 vdd.n4505 vss 0.00306f
C7141 vdd.n4506 vss 0.00651f
C7142 vdd.n4507 vss 0.0188f
C7143 vdd.n4508 vss 0.0116f
C7144 vdd.n4509 vss 0.0113f
C7145 vdd.n4510 vss -0.0615f
C7146 vdd.n4511 vss 0.00271f
C7147 vdd.n4512 vss 0.00335f
C7148 vdd.n4513 vss 0.00748f
C7149 vdd.n4514 vss 0.00542f
C7150 vdd.n4515 vss 0.00658f
C7151 vdd.n4516 vss 0.00284f
C7152 vdd.n4517 vss 0.00219f
C7153 vdd.n4518 vss 0.00284f
C7154 vdd.n4519 vss 2.58e-19
C7155 vdd.n4520 vss 0.00219f
C7156 vdd.n4521 vss 0.00226f
C7157 vdd.n4522 vss 0.043f
C7158 vdd.n4523 vss 0.2f
C7159 vdd.n4524 vss 0.162f
C7160 vdd.n4525 vss 0.00851f
C7161 vdd.n4526 vss 0.0341f
C7162 vdd.n4527 vss 0.0344f
C7163 vdd.n4528 vss 0.0318f
C7164 vdd.n4529 vss 0.0325f
C7165 vdd.n4530 vss 0.0117f
C7166 vdd.n4531 vss 0.0358f
C7167 vdd.n4532 vss 0.114f
C7168 vdd.n4533 vss 0.0118f
C7169 vdd.n4534 vss 0.0114f
C7170 vdd.n4535 vss -0.0615f
C7171 vdd.n4536 vss 0.00271f
C7172 vdd.n4537 vss 0.00335f
C7173 vdd.n4538 vss 0.00776f
C7174 vdd.n4539 vss 0.00542f
C7175 vdd.n4540 vss 0.00658f
C7176 vdd.n4541 vss 0.00284f
C7177 vdd.n4542 vss 0.00219f
C7178 vdd.n4543 vss 0.00284f
C7179 vdd.n4544 vss 2.58e-19
C7180 vdd.n4545 vss 0.00219f
C7181 vdd.n4546 vss 0.00226f
C7182 vdd.n4547 vss 0.043f
C7183 vdd.n4548 vss 0.2f
C7184 vdd.n4549 vss 0.162f
C7185 vdd.n4550 vss 0.00851f
C7186 vdd.n4551 vss 2.58e-19
C7187 vdd.n4552 vss 0.00284f
C7188 vdd.n4553 vss 0.00748f
C7189 vdd.n4554 vss 0.00335f
C7190 vdd.n4555 vss 0.00477f
C7191 vdd.n4556 vss 0.00385f
C7192 vdd.n4557 vss 0.00306f
C7193 vdd.n4558 vss 0.00651f
C7194 vdd.n4559 vss 0.0191f
C7195 vdd.n4560 vss 0.0118f
C7196 vdd.n4561 vss 0.0114f
C7197 vdd.n4562 vss -0.0615f
C7198 vdd.n4563 vss 0.00271f
C7199 vdd.n4564 vss 0.00335f
C7200 vdd.n4565 vss 0.00748f
C7201 vdd.n4566 vss 0.00542f
C7202 vdd.n4567 vss 0.00658f
C7203 vdd.n4568 vss 0.00284f
C7204 vdd.n4569 vss 0.00219f
C7205 vdd.n4570 vss 0.00284f
C7206 vdd.n4571 vss 2.58e-19
C7207 vdd.n4572 vss 0.00219f
C7208 vdd.n4573 vss 0.00226f
C7209 vdd.n4574 vss 0.043f
C7210 vdd.n4575 vss 0.2f
C7211 vdd.n4576 vss 0.162f
C7212 vdd.n4577 vss 0.00851f
C7213 vdd.n4578 vss 2.58e-19
C7214 vdd.n4579 vss 0.00247f
C7215 vdd.n4580 vss 0.0071f
C7216 vdd.n4581 vss 0.0152f
C7217 vdd.n4582 vss 0.0835f
C7218 vdd.n4583 vss 0.361f
C7219 vdd.t37 vss 0.651f
C7220 vdd.n4584 vss 0.076f
C7221 vdd.n4585 vss 0.0256f
C7222 vdd.n4586 vss 0.00209f
C7223 vdd.n4587 vss 0.00394f
C7224 vdd.n4588 vss 0.00338f
C7225 vdd.n4589 vss 0.00362f
C7226 vdd.n4590 vss 0.00563f
C7227 vdd.n4591 vss 6.66e-19
C7228 vdd.n4592 vss 0.0151f
C7229 vdd.n4593 vss 0.0334f
C7230 vdd.n4594 vss 0.0152f
C7231 vdd.n4595 vss 0.0139f
C7232 vdd.n4596 vss 0.00563f
C7233 vdd.n4597 vss 0.00564f
C7234 vdd.n4598 vss 0.0101f
C7235 vdd.n4599 vss 0.00903f
C7236 vdd.n4600 vss 0.00466f
C7237 vdd.n4601 vss 0.0163f
C7238 vdd.n4602 vss 0.0213f
C7239 vdd.n4603 vss 0.0493f
C7240 vdd.n4604 vss 0.0224f
C7241 vdd.n4605 vss 0.0162f
C7242 vdd.n4606 vss 0.0173f
C7243 vdd.n4607 vss 0.00886f
C7244 vdd.t127 vss 0.0416f
C7245 vdd.n4608 vss 0.019f
C7246 vdd.n4609 vss 0.0458f
C7247 vdd.n4610 vss 0.00651f
C7248 vdd.n4611 vss 0.00864f
C7249 vdd.n4612 vss 0.0169f
C7250 vdd.n4613 vss 0.00619f
C7251 vdd.n4614 vss 0.00318f
C7252 vdd.n4615 vss 0.00376f
C7253 vdd.n4616 vss 0.00319f
C7254 vdd.n4617 vss 0.0015f
C7255 vdd.n4618 vss 0.00111f
C7256 vdd.n4619 vss 0.0114f
C7257 vdd.n4620 vss 0.0746f
C7258 vdd.n4621 vss 0.0122f
C7259 vdd.n4622 vss 0.0617f
C7260 vdd.n4623 vss 0.0102f
C7261 vdd.n4624 vss 0.00888f
C7262 vdd.n4625 vss 0.00814f
C7263 vdd.n4626 vss 0.0214f
C7264 vdd.n4627 vss 0.0141f
C7265 vdd.n4628 vss 0.0161f
C7266 vdd.n4629 vss 6.66e-19
C7267 vdd.n4630 vss 0.0101f
C7268 vdd.n4631 vss 0.501f
C7269 vdd.n4632 vss 3.96f
C7270 vdd.n4633 vss 7.21f
C7271 vdd.n4634 vss 0.363f
C7272 vdd.n4635 vss 0.243f
C7273 vdd.n4636 vss 0.0163f
C7274 vdd.n4637 vss 0.00673f
C7275 vdd.n4638 vss 0.0163f
C7276 vdd.n4639 vss 0.00518f
C7277 vdd.n4640 vss 0.00668f
C7278 vdd.n4641 vss 0.0664f
C7279 vdd.n4642 vss 1.03f
C7280 vdd.t117 vss 0.156f
C7281 vdd.n4643 vss 0.14f
C7282 vdd.n4644 vss 1.49f
C7283 vdd.t88 vss 1.43f
C7284 vdd.n4645 vss 0.00673f
C7285 vdd.n4646 vss 0.0163f
C7286 vdd.n4647 vss 0.0163f
C7287 vdd.n4648 vss 0.00887f
C7288 vdd.n4649 vss 0.00518f
C7289 vdd.n4650 vss 0.00668f
C7290 vdd.n4651 vss 0.0664f
C7291 vdd.t4 vss 0.35f
C7292 vdd.t99 vss 0.732f
C7293 vdd.n4652 vss 0.0127f
C7294 vdd.t39 vss 1.8f
C7295 vdd.t71 vss 5.45f
C7296 vdd.t89 vss 4.45f
C7297 vdd.n4653 vss 1.69f
C7298 vdd.t93 vss 1.9f
C7299 vdd.n4654 vss 1.69f
C7300 vdd.n4655 vss 0.00673f
C7301 vdd.n4656 vss 0.0664f
C7302 vdd.n4657 vss 0.00668f
C7303 vdd.n4658 vss 0.0163f
C7304 vdd.n4659 vss 0.00887f
C7305 vdd.n4660 vss 0.0547f
C7306 vdd.n4661 vss 0.0635f
C7307 vdd.n4662 vss 0.0163f
C7308 vdd.n4663 vss 0.00673f
C7309 vdd.n4664 vss 0.0664f
C7310 vdd.n4665 vss 0.00668f
C7311 vdd.n4666 vss 0.0163f
C7312 vdd.n4667 vss 0.0482f
C7313 vdd.n4668 vss 0.103f
C7314 vdd.n4669 vss 0.0163f
C7315 vdd.t72 vss 0.0077f
C7316 vdd.n4670 vss 0.111f
C7317 vdd.n4671 vss 0.0163f
C7318 vdd.n4672 vss 0.142f
C7319 vdd.n4673 vss 28.7f
C7320 vdd.n4674 vss 0.0115f
C7321 vdd.n4675 vss 0.0111f
C7322 vdd.n4676 vss 0.00359f
C7323 vdd.n4677 vss 0.0325f
C7324 vdd.n4678 vss 0.0318f
C7325 vdd.n4679 vss 0.0361f
C7326 vdd.n4680 vss 0.0344f
C7327 vdd.n4681 vss 3.87e-19
C7328 vdd.n4682 vss 0.00399f
C7329 vdd.n4683 vss 0.00651f
C7330 vdd.n4684 vss -0.143f
C7331 vdd.n4685 vss 0.0182f
C7332 vdd.n4686 vss 0.0111f
C7333 vdd.n4687 vss 0.00359f
C7334 vdd.n4688 vss 0.00385f
C7335 vdd.n4689 vss 0.00477f
C7336 vdd.n4690 vss 0.00658f
C7337 vdd.n4691 vss 0.00542f
C7338 vdd.n4692 vss 0.00271f
C7339 vdd.n4693 vss 0.008f
C7340 vdd.n4694 vss 0.008f
C7341 vdd.n4695 vss 0.0105f
C7342 vdd.n4697 vss 0.00226f
C7343 vdd.n4699 vss 0.00851f
C7344 vdd.n4700 vss 2.58e-19
C7345 vdd.n4701 vss 0.00284f
C7346 vdd.n4702 vss 3.87e-19
C7347 vdd.n4703 vss 0.00399f
C7348 vdd.n4704 vss 0.00651f
C7349 vdd.n4705 vss 0.0186f
C7350 vdd.n4706 vss 0.0182f
C7351 vdd.n4707 vss 0.0111f
C7352 vdd.n4708 vss 0.00306f
C7353 vdd.n4709 vss 0.0115f
C7354 vdd.n4710 vss 0.0182f
C7355 vdd.n4711 vss 0.0186f
C7356 vdd.n4712 vss 0.00651f
C7357 vdd.n4713 vss 0.00399f
C7358 vdd.n4714 vss 0.00284f
C7359 vdd.n4715 vss 3.87e-19
C7360 vdd.n4716 vss 0.00271f
C7361 vdd.n4717 vss -0.0615f
C7362 vdd.n4718 vss -0.173f
C7363 vdd.n4719 vss 0.00477f
C7364 vdd.n4720 vss 0.00658f
C7365 vdd.n4721 vss 0.00542f
C7366 vdd.n4722 vss 0.00271f
C7367 vdd.n4723 vss 0.008f
C7368 vdd.n4724 vss 0.008f
C7369 vdd.n4725 vss 0.00219f
C7370 vdd.n4726 vss 0.00226f
C7371 vdd.n4728 vss 0.00851f
C7372 vdd.n4730 vss 0.0105f
C7373 vdd.n4731 vss 0.008f
C7374 vdd.n4732 vss 0.008f
C7375 vdd.n4733 vss 0.00271f
C7376 vdd.n4734 vss 0.00542f
C7377 vdd.n4735 vss 0.00658f
C7378 vdd.n4736 vss 0.00477f
C7379 vdd.n4737 vss 0.00335f
C7380 vdd.n4738 vss 0.00271f
C7381 vdd.n4739 vss 0.00359f
C7382 vdd.n4740 vss 2.66e-19
C7383 vdd.n4741 vss 0.00399f
C7384 vdd.n4742 vss 0.00651f
C7385 vdd.n4743 vss -0.143f
C7386 vdd.n4744 vss 0.0182f
C7387 vdd.n4745 vss 0.0111f
C7388 vdd.n4746 vss 0.00359f
C7389 vdd.n4747 vss 0.00385f
C7390 vdd.n4748 vss 0.00477f
C7391 vdd.n4749 vss 0.00542f
C7392 vdd.n4750 vss 0.00658f
C7393 vdd.n4751 vss 0.00284f
C7394 vdd.n4752 vss 0.00219f
C7395 vdd.n4753 vss 0.00284f
C7396 vdd.n4754 vss 2.58e-19
C7397 vdd.n4755 vss 0.00851f
C7398 vdd.n4757 vss 0.0105f
C7399 vdd.n4759 vss 0.00226f
C7400 vdd.n4760 vss 0.00219f
C7401 vdd.n4761 vss 2.58e-19
C7402 vdd.n4762 vss 0.00284f
C7403 vdd.n4763 vss 3.87e-19
C7404 vdd.n4764 vss 0.00399f
C7405 vdd.n4765 vss 0.00651f
C7406 vdd.n4766 vss 0.0186f
C7407 vdd.n4767 vss 0.0182f
C7408 vdd.n4768 vss 0.0115f
C7409 vdd.n4769 vss 0.0111f
C7410 vdd.n4770 vss -0.0615f
C7411 vdd.n4771 vss -0.173f
C7412 vdd.n4772 vss 0.00477f
C7413 vdd.n4773 vss 0.00658f
C7414 vdd.n4774 vss 0.00542f
C7415 vdd.n4775 vss 0.00271f
C7416 vdd.n4776 vss 0.008f
C7417 vdd.n4777 vss 0.008f
C7418 vdd.n4778 vss 0.0105f
C7419 vdd.n4780 vss 0.00226f
C7420 vdd.n4781 vss 0.0193f
C7421 vdd.n4782 vss 2.58e-19
C7422 vdd.n4783 vss 0.00284f
C7423 vdd.n4784 vss 3.87e-19
C7424 vdd.n4785 vss 0.00399f
C7425 vdd.n4786 vss 0.0234f
C7426 vdd.n4787 vss 0.00385f
C7427 vdd.n4788 vss 0.0233f
C7428 vdd.n4789 vss 0.0654f
C7429 vdd.n4790 vss 0.0111f
C7430 vdd.n4791 vss 0.0182f
C7431 vdd.n4792 vss 0.00385f
C7432 vdd.n4793 vss 0.00638f
C7433 vdd.n4794 vss 0.00319f
C7434 vdd.n4795 vss 0.0186f
C7435 vdd.n4796 vss 0.0115f
C7436 vdd.n4797 vss -0.0615f
C7437 vdd.n4798 vss 0.00271f
C7438 vdd.n4799 vss 0.00335f
C7439 vdd.n4800 vss 0.00748f
C7440 vdd.n4801 vss 0.00542f
C7441 vdd.n4802 vss 0.00658f
C7442 vdd.n4803 vss 0.00284f
C7443 vdd.n4804 vss 0.00219f
C7444 vdd.n4805 vss 0.00219f
C7445 vdd.n4806 vss 2.58e-19
C7446 vdd.n4807 vss 0.00851f
C7447 vdd.n4809 vss 0.00226f
C7448 vdd.n4811 vss 0.0105f
C7449 vdd.n4812 vss 0.008f
C7450 vdd.n4813 vss 0.008f
C7451 vdd.n4814 vss 0.00271f
C7452 vdd.n4815 vss 0.00284f
C7453 vdd.n4816 vss 0.00658f
C7454 vdd.n4817 vss 0.00542f
C7455 vdd.n4818 vss 0.00748f
C7456 vdd.n4819 vss 0.00335f
C7457 vdd.n4820 vss 0.00271f
C7458 vdd.n4821 vss 0.00359f
C7459 vdd.n4822 vss 0.0115f
C7460 vdd.n4823 vss 0.0186f
C7461 vdd.n4824 vss 0.00319f
C7462 vdd.n4825 vss 0.00638f
C7463 vdd.n4826 vss 0.00385f
C7464 vdd.n4827 vss 2.66e-19
C7465 vdd.n4828 vss -0.0638f
C7466 vdd.n4829 vss 0.0115f
C7467 vdd.n4830 vss 0.0186f
C7468 vdd.n4831 vss 0.00319f
C7469 vdd.n4832 vss 0.00399f
C7470 vdd.n4833 vss 0.00477f
C7471 vdd.n4834 vss 0.00335f
C7472 vdd.n4835 vss 0.00748f
C7473 vdd.n4836 vss 0.00284f
C7474 vdd.n4837 vss 2.58e-19
C7475 vdd.n4838 vss 0.00219f
C7476 vdd.n4839 vss 0.00226f
C7477 vdd.n4841 vss 0.0105f
C7478 vdd.n4843 vss 0.00851f
C7479 vdd.n4844 vss 2.58e-19
C7480 vdd.n4845 vss 0.00284f
C7481 vdd.n4846 vss 3.87e-19
C7482 vdd.n4847 vss 0.00385f
C7483 vdd.n4848 vss 2.66e-19
C7484 vdd.n4849 vss 0.0111f
C7485 vdd.n4850 vss 0.0115f
C7486 vdd.n4851 vss 0.0182f
C7487 vdd.n4852 vss 0.0186f
C7488 vdd.n4853 vss 0.00319f
C7489 vdd.n4854 vss -0.173f
C7490 vdd.n4855 vss 0.00477f
C7491 vdd.n4856 vss 0.00658f
C7492 vdd.n4857 vss 0.00284f
C7493 vdd.n4858 vss 0.00219f
C7494 vdd.n4859 vss 0.00271f
C7495 vdd.n4860 vss 0.008f
C7496 vdd.n4861 vss 0.008f
C7497 vdd.n4862 vss 0.0105f
C7498 vdd.n4864 vss 0.00851f
C7499 vdd.n4866 vss 0.00226f
C7500 vdd.n4867 vss 0.00219f
C7501 vdd.n4868 vss 0.008f
C7502 vdd.n4869 vss 0.008f
C7503 vdd.n4870 vss 0.00271f
C7504 vdd.n4871 vss 0.00284f
C7505 vdd.n4872 vss 0.00658f
C7506 vdd.n4873 vss 0.00542f
C7507 vdd.n4874 vss 0.00748f
C7508 vdd.n4875 vss 0.00335f
C7509 vdd.n4876 vss 0.00271f
C7510 vdd.n4877 vss 0.00359f
C7511 vdd.n4878 vss 0.0115f
C7512 vdd.n4879 vss 0.0186f
C7513 vdd.n4880 vss 0.00319f
C7514 vdd.n4881 vss 0.00638f
C7515 vdd.n4882 vss 0.00385f
C7516 vdd.n4883 vss 2.66e-19
C7517 vdd.n4884 vss -0.0638f
C7518 vdd.n4885 vss 0.0115f
C7519 vdd.n4886 vss 0.00385f
C7520 vdd.n4887 vss 0.00359f
C7521 vdd.n4888 vss 0.0111f
C7522 vdd.n4889 vss 0.0115f
C7523 vdd.n4890 vss 0.049f
C7524 vdd.n4891 vss 0.0198f
C7525 vdd.n4892 vss 0.00399f
C7526 vdd.n4893 vss 0.0205f
C7527 vdd.n4894 vss 0.00335f
C7528 vdd.n4895 vss 0.0241f
C7529 vdd.n4896 vss 0.00284f
C7530 vdd.n4897 vss 2.58e-19
C7531 vdd.n4898 vss 0.00851f
C7532 vdd.n4900 vss 0.00226f
C7533 vdd.n4901 vss 0.0152f
C7534 vdd.n4902 vss 0.0245f
C7535 vdd.n4903 vss 0.0255f
C7536 vdd.n4904 vss 0.0142f
C7537 vdd.n4905 vss 0.00226f
C7538 vdd.n4906 vss 0.00219f
C7539 vdd.n4907 vss 2.58e-19
C7540 vdd.n4908 vss 0.00284f
C7541 vdd.n4909 vss 3.87e-19
C7542 vdd.n4910 vss 0.00399f
C7543 vdd.n4911 vss 0.00651f
C7544 vdd.n4912 vss -0.143f
C7545 vdd.n4913 vss 0.0182f
C7546 vdd.n4914 vss 0.0111f
C7547 vdd.n4915 vss 0.00359f
C7548 vdd.n4916 vss 0.00385f
C7549 vdd.n4917 vss 0.00477f
C7550 vdd.n4918 vss 0.00658f
C7551 vdd.n4919 vss 0.00542f
C7552 vdd.n4920 vss 0.00271f
C7553 vdd.n4921 vss 0.008f
C7554 vdd.n4922 vss 0.008f
C7555 vdd.n4923 vss 0.0105f
C7556 vdd.n4925 vss 0.00226f
C7557 vdd.n4927 vss 0.00851f
C7558 vdd.n4928 vss 2.58e-19
C7559 vdd.n4929 vss 0.00284f
C7560 vdd.n4930 vss 3.87e-19
C7561 vdd.n4931 vss 0.00399f
C7562 vdd.n4932 vss 0.00651f
C7563 vdd.n4933 vss 0.0186f
C7564 vdd.n4934 vss 0.0182f
C7565 vdd.n4935 vss 0.0111f
C7566 vdd.n4936 vss 0.00306f
C7567 vdd.n4937 vss 0.0115f
C7568 vdd.n4938 vss 0.0182f
C7569 vdd.n4939 vss 0.0186f
C7570 vdd.n4940 vss 0.00651f
C7571 vdd.n4941 vss 0.00399f
C7572 vdd.n4942 vss 0.00284f
C7573 vdd.n4943 vss 3.87e-19
C7574 vdd.n4944 vss 0.00271f
C7575 vdd.n4945 vss -0.0615f
C7576 vdd.n4946 vss -0.173f
C7577 vdd.n4947 vss 0.00477f
C7578 vdd.n4948 vss 0.00658f
C7579 vdd.n4949 vss 0.00542f
C7580 vdd.n4950 vss 0.00271f
C7581 vdd.n4951 vss 0.008f
C7582 vdd.n4952 vss 0.008f
C7583 vdd.n4953 vss 0.00219f
C7584 vdd.n4954 vss 0.00226f
C7585 vdd.n4956 vss 0.00851f
C7586 vdd.n4958 vss 0.0105f
C7587 vdd.n4959 vss 0.008f
C7588 vdd.n4960 vss 0.008f
C7589 vdd.n4961 vss 0.00271f
C7590 vdd.n4962 vss 0.00542f
C7591 vdd.n4963 vss 0.00658f
C7592 vdd.n4964 vss 0.00477f
C7593 vdd.n4965 vss 0.00335f
C7594 vdd.n4966 vss 0.00271f
C7595 vdd.n4967 vss 0.00359f
C7596 vdd.n4968 vss 2.66e-19
C7597 vdd.n4969 vss 0.00399f
C7598 vdd.n4970 vss 0.00651f
C7599 vdd.n4971 vss -0.143f
C7600 vdd.n4972 vss 0.0182f
C7601 vdd.n4973 vss 0.0111f
C7602 vdd.n4974 vss 0.00359f
C7603 vdd.n4975 vss 0.00385f
C7604 vdd.n4976 vss 0.00477f
C7605 vdd.n4977 vss 0.00542f
C7606 vdd.n4978 vss 0.00658f
C7607 vdd.n4979 vss 0.00284f
C7608 vdd.n4980 vss 0.00219f
C7609 vdd.n4981 vss 0.00284f
C7610 vdd.n4982 vss 2.58e-19
C7611 vdd.n4983 vss 0.00851f
C7612 vdd.n4985 vss 0.0105f
C7613 vdd.n4987 vss 0.00226f
C7614 vdd.n4988 vss 0.00219f
C7615 vdd.n4989 vss 2.58e-19
C7616 vdd.n4990 vss 0.00284f
C7617 vdd.n4991 vss 3.87e-19
C7618 vdd.n4992 vss 0.00399f
C7619 vdd.n4993 vss 0.00651f
C7620 vdd.n4994 vss 0.0186f
C7621 vdd.n4995 vss 0.0182f
C7622 vdd.n4996 vss 0.0115f
C7623 vdd.n4997 vss 0.0111f
C7624 vdd.n4998 vss -0.0615f
C7625 vdd.n4999 vss -0.173f
C7626 vdd.n5000 vss 0.00477f
C7627 vdd.n5001 vss 0.00658f
C7628 vdd.n5002 vss 0.00542f
C7629 vdd.n5003 vss 0.00271f
C7630 vdd.n5004 vss 0.008f
C7631 vdd.n5005 vss 0.008f
C7632 vdd.n5006 vss 0.0105f
C7633 vdd.n5008 vss 0.00226f
C7634 vdd.n5009 vss 0.0193f
C7635 vdd.n5010 vss 2.58e-19
C7636 vdd.n5011 vss 0.00284f
C7637 vdd.n5012 vss 3.87e-19
C7638 vdd.n5013 vss 0.00399f
C7639 vdd.n5014 vss 0.0234f
C7640 vdd.n5015 vss 0.00385f
C7641 vdd.n5016 vss 0.0233f
C7642 vdd.n5017 vss 0.0654f
C7643 vdd.n5018 vss 0.0111f
C7644 vdd.n5019 vss 0.0182f
C7645 vdd.n5020 vss 0.00385f
C7646 vdd.n5021 vss 0.00638f
C7647 vdd.n5022 vss 0.00319f
C7648 vdd.n5023 vss 0.0186f
C7649 vdd.n5024 vss 0.0115f
C7650 vdd.n5025 vss -0.0615f
C7651 vdd.n5026 vss 0.00271f
C7652 vdd.n5027 vss 0.00335f
C7653 vdd.n5028 vss 0.00748f
C7654 vdd.n5029 vss 0.00542f
C7655 vdd.n5030 vss 0.00658f
C7656 vdd.n5031 vss 0.00284f
C7657 vdd.n5032 vss 0.00219f
C7658 vdd.n5033 vss 0.00219f
C7659 vdd.n5034 vss 2.58e-19
C7660 vdd.n5035 vss 0.00851f
C7661 vdd.n5037 vss 0.00226f
C7662 vdd.n5039 vss 0.0105f
C7663 vdd.n5040 vss 0.008f
C7664 vdd.n5041 vss 0.008f
C7665 vdd.n5042 vss 0.00271f
C7666 vdd.n5043 vss 0.00284f
C7667 vdd.n5044 vss 0.00658f
C7668 vdd.n5045 vss 0.00542f
C7669 vdd.n5046 vss 0.00748f
C7670 vdd.n5047 vss 0.00335f
C7671 vdd.n5048 vss 0.00271f
C7672 vdd.n5049 vss 0.00359f
C7673 vdd.n5050 vss 0.0115f
C7674 vdd.n5051 vss 0.0186f
C7675 vdd.n5052 vss 0.00319f
C7676 vdd.n5053 vss 0.00638f
C7677 vdd.n5054 vss 0.00385f
C7678 vdd.n5055 vss 2.66e-19
C7679 vdd.n5056 vss -0.0638f
C7680 vdd.n5057 vss 0.0115f
C7681 vdd.n5058 vss 0.0186f
C7682 vdd.n5059 vss 0.00319f
C7683 vdd.n5060 vss 0.00399f
C7684 vdd.n5061 vss 0.00477f
C7685 vdd.n5062 vss 0.00335f
C7686 vdd.n5063 vss 0.00748f
C7687 vdd.n5064 vss 0.00284f
C7688 vdd.n5065 vss 2.58e-19
C7689 vdd.n5066 vss 0.00219f
C7690 vdd.n5067 vss 0.00226f
C7691 vdd.n5069 vss 0.0105f
C7692 vdd.n5071 vss 0.00851f
C7693 vdd.n5072 vss 2.58e-19
C7694 vdd.n5073 vss 0.00284f
C7695 vdd.n5074 vss 3.87e-19
C7696 vdd.n5075 vss 0.00385f
C7697 vdd.n5076 vss 2.66e-19
C7698 vdd.n5077 vss 0.0111f
C7699 vdd.n5078 vss 0.0115f
C7700 vdd.n5079 vss 0.0182f
C7701 vdd.n5080 vss 0.0186f
C7702 vdd.n5081 vss 0.00319f
C7703 vdd.n5082 vss -0.173f
C7704 vdd.n5083 vss 0.00477f
C7705 vdd.n5084 vss 0.00658f
C7706 vdd.n5085 vss 0.00284f
C7707 vdd.n5086 vss 0.00219f
C7708 vdd.n5087 vss 0.00271f
C7709 vdd.n5088 vss 0.008f
C7710 vdd.n5089 vss 0.008f
C7711 vdd.n5090 vss 0.0105f
C7712 vdd.n5092 vss 0.00851f
C7713 vdd.n5094 vss 0.00226f
C7714 vdd.n5095 vss 0.00219f
C7715 vdd.n5096 vss 0.008f
C7716 vdd.n5097 vss 0.008f
C7717 vdd.n5098 vss 0.00271f
C7718 vdd.n5099 vss 0.00284f
C7719 vdd.n5100 vss 0.00658f
C7720 vdd.n5101 vss 0.00542f
C7721 vdd.n5102 vss 0.00748f
C7722 vdd.n5103 vss 0.00335f
C7723 vdd.n5104 vss 0.00271f
C7724 vdd.n5105 vss 0.00359f
C7725 vdd.n5106 vss 0.0115f
C7726 vdd.n5107 vss 0.0186f
C7727 vdd.n5108 vss 0.00319f
C7728 vdd.n5109 vss 0.00638f
C7729 vdd.n5110 vss 0.00385f
C7730 vdd.n5111 vss 2.66e-19
C7731 vdd.n5112 vss -0.0638f
C7732 vdd.n5113 vss 0.0115f
C7733 vdd.n5114 vss 0.00385f
C7734 vdd.n5115 vss 0.00359f
C7735 vdd.n5116 vss 0.0111f
C7736 vdd.n5117 vss 0.0115f
C7737 vdd.n5118 vss 0.049f
C7738 vdd.n5119 vss 0.0198f
C7739 vdd.n5120 vss 0.00399f
C7740 vdd.n5121 vss 0.0205f
C7741 vdd.n5122 vss 0.00335f
C7742 vdd.n5123 vss 0.0241f
C7743 vdd.n5124 vss 0.00284f
C7744 vdd.n5125 vss 2.58e-19
C7745 vdd.n5126 vss 0.00851f
C7746 vdd.n5128 vss 0.00226f
C7747 vdd.n5129 vss 0.0152f
C7748 vdd.n5130 vss 0.0245f
C7749 vdd.n5131 vss 0.0255f
C7750 vdd.n5132 vss 0.0142f
C7751 vdd.n5133 vss 0.00226f
C7752 vdd.n5134 vss 0.00219f
C7753 vdd.n5135 vss 2.58e-19
C7754 vdd.n5136 vss 0.00284f
C7755 vdd.n5137 vss 3.87e-19
C7756 vdd.n5138 vss 0.00399f
C7757 vdd.n5139 vss 0.00651f
C7758 vdd.n5140 vss -0.143f
C7759 vdd.n5141 vss 0.0182f
C7760 vdd.n5142 vss 0.0111f
C7761 vdd.n5143 vss 0.00359f
C7762 vdd.n5144 vss 0.00385f
C7763 vdd.n5145 vss 0.00477f
C7764 vdd.n5146 vss 0.00658f
C7765 vdd.n5147 vss 0.00542f
C7766 vdd.n5148 vss 0.00271f
C7767 vdd.n5149 vss 0.008f
C7768 vdd.n5150 vss 0.008f
C7769 vdd.n5151 vss 0.0105f
C7770 vdd.n5153 vss 0.00226f
C7771 vdd.n5155 vss 0.00851f
C7772 vdd.n5156 vss 2.58e-19
C7773 vdd.n5157 vss 0.00284f
C7774 vdd.n5158 vss 3.87e-19
C7775 vdd.n5159 vss 0.00399f
C7776 vdd.n5160 vss 0.00651f
C7777 vdd.n5161 vss 0.0186f
C7778 vdd.n5162 vss 0.0182f
C7779 vdd.n5163 vss 0.0111f
C7780 vdd.n5164 vss 0.00306f
C7781 vdd.n5165 vss 0.0115f
C7782 vdd.n5166 vss 0.0182f
C7783 vdd.n5167 vss 0.0186f
C7784 vdd.n5168 vss 0.00651f
C7785 vdd.n5169 vss 0.00399f
C7786 vdd.n5170 vss 0.00284f
C7787 vdd.n5171 vss 3.87e-19
C7788 vdd.n5172 vss 0.00271f
C7789 vdd.n5173 vss -0.0615f
C7790 vdd.n5174 vss -0.173f
C7791 vdd.n5175 vss 0.00477f
C7792 vdd.n5176 vss 0.00658f
C7793 vdd.n5177 vss 0.00542f
C7794 vdd.n5178 vss 0.00271f
C7795 vdd.n5179 vss 0.008f
C7796 vdd.n5180 vss 0.008f
C7797 vdd.n5181 vss 0.00219f
C7798 vdd.n5182 vss 0.00226f
C7799 vdd.n5184 vss 0.00851f
C7800 vdd.n5186 vss 0.0105f
C7801 vdd.n5187 vss 0.008f
C7802 vdd.n5188 vss 0.008f
C7803 vdd.n5189 vss 0.00271f
C7804 vdd.n5190 vss 0.00542f
C7805 vdd.n5191 vss 0.00658f
C7806 vdd.n5192 vss 0.00477f
C7807 vdd.n5193 vss 0.00335f
C7808 vdd.n5194 vss 0.00271f
C7809 vdd.n5195 vss 0.00359f
C7810 vdd.n5196 vss 2.66e-19
C7811 vdd.n5197 vss 0.00399f
C7812 vdd.n5198 vss 0.00651f
C7813 vdd.n5199 vss -0.143f
C7814 vdd.n5200 vss 0.0182f
C7815 vdd.n5201 vss 0.0111f
C7816 vdd.n5202 vss 0.00359f
C7817 vdd.n5203 vss 0.00385f
C7818 vdd.n5204 vss 0.00477f
C7819 vdd.n5205 vss 0.00542f
C7820 vdd.n5206 vss 0.00658f
C7821 vdd.n5207 vss 0.00284f
C7822 vdd.n5208 vss 0.00219f
C7823 vdd.n5209 vss 0.00284f
C7824 vdd.n5210 vss 2.58e-19
C7825 vdd.n5211 vss 0.00851f
C7826 vdd.n5213 vss 0.0105f
C7827 vdd.n5215 vss 0.00226f
C7828 vdd.n5216 vss 0.00219f
C7829 vdd.n5217 vss 2.58e-19
C7830 vdd.n5218 vss 0.00284f
C7831 vdd.n5219 vss 3.87e-19
C7832 vdd.n5220 vss 0.00399f
C7833 vdd.n5221 vss 0.00651f
C7834 vdd.n5222 vss 0.0186f
C7835 vdd.n5223 vss 0.0182f
C7836 vdd.n5224 vss 0.0115f
C7837 vdd.n5225 vss 0.0111f
C7838 vdd.n5226 vss -0.0615f
C7839 vdd.n5227 vss -0.173f
C7840 vdd.n5228 vss 0.00477f
C7841 vdd.n5229 vss 0.00658f
C7842 vdd.n5230 vss 0.00542f
C7843 vdd.n5231 vss 0.00271f
C7844 vdd.n5232 vss 0.008f
C7845 vdd.n5233 vss 0.008f
C7846 vdd.n5234 vss 0.0105f
C7847 vdd.n5236 vss 0.00226f
C7848 vdd.n5237 vss 0.0193f
C7849 vdd.n5238 vss 2.58e-19
C7850 vdd.n5239 vss 0.00284f
C7851 vdd.n5240 vss 3.87e-19
C7852 vdd.n5241 vss 0.00399f
C7853 vdd.n5242 vss 0.0234f
C7854 vdd.n5243 vss 0.00385f
C7855 vdd.n5244 vss 0.0233f
C7856 vdd.n5245 vss 0.0654f
C7857 vdd.n5246 vss 0.0111f
C7858 vdd.n5247 vss 0.0182f
C7859 vdd.n5248 vss 0.00385f
C7860 vdd.n5249 vss 0.00638f
C7861 vdd.n5250 vss 0.00319f
C7862 vdd.n5251 vss 0.0186f
C7863 vdd.n5252 vss 0.0115f
C7864 vdd.n5253 vss -0.0615f
C7865 vdd.n5254 vss 0.00271f
C7866 vdd.n5255 vss 0.00335f
C7867 vdd.n5256 vss 0.00748f
C7868 vdd.n5257 vss 0.00542f
C7869 vdd.n5258 vss 0.00658f
C7870 vdd.n5259 vss 0.00284f
C7871 vdd.n5260 vss 0.00219f
C7872 vdd.n5261 vss 0.00219f
C7873 vdd.n5262 vss 2.58e-19
C7874 vdd.n5263 vss 0.00851f
C7875 vdd.n5265 vss 0.00226f
C7876 vdd.n5267 vss 0.0105f
C7877 vdd.n5268 vss 0.008f
C7878 vdd.n5269 vss 0.008f
C7879 vdd.n5270 vss 0.00271f
C7880 vdd.n5271 vss 0.00284f
C7881 vdd.n5272 vss 0.00658f
C7882 vdd.n5273 vss 0.00542f
C7883 vdd.n5274 vss 0.00748f
C7884 vdd.n5275 vss 0.00335f
C7885 vdd.n5276 vss 0.00271f
C7886 vdd.n5277 vss 0.00359f
C7887 vdd.n5278 vss 0.0115f
C7888 vdd.n5279 vss 0.0186f
C7889 vdd.n5280 vss 0.00319f
C7890 vdd.n5281 vss 0.00638f
C7891 vdd.n5282 vss 0.00385f
C7892 vdd.n5283 vss 2.66e-19
C7893 vdd.n5284 vss -0.0638f
C7894 vdd.n5285 vss 0.0115f
C7895 vdd.n5286 vss 0.0186f
C7896 vdd.n5287 vss 0.00319f
C7897 vdd.n5288 vss 0.00399f
C7898 vdd.n5289 vss 0.00477f
C7899 vdd.n5290 vss 0.00335f
C7900 vdd.n5291 vss 0.00748f
C7901 vdd.n5292 vss 0.00284f
C7902 vdd.n5293 vss 2.58e-19
C7903 vdd.n5294 vss 0.00219f
C7904 vdd.n5295 vss 0.00226f
C7905 vdd.n5297 vss 0.0105f
C7906 vdd.n5299 vss 0.00851f
C7907 vdd.n5300 vss 2.58e-19
C7908 vdd.n5301 vss 0.00284f
C7909 vdd.n5302 vss 3.87e-19
C7910 vdd.n5303 vss 0.00385f
C7911 vdd.n5304 vss 2.66e-19
C7912 vdd.n5305 vss 0.0111f
C7913 vdd.n5306 vss 0.0115f
C7914 vdd.n5307 vss 0.0182f
C7915 vdd.n5308 vss 0.0186f
C7916 vdd.n5309 vss 0.00319f
C7917 vdd.n5310 vss -0.173f
C7918 vdd.n5311 vss 0.00477f
C7919 vdd.n5312 vss 0.00658f
C7920 vdd.n5313 vss 0.00284f
C7921 vdd.n5314 vss 0.00219f
C7922 vdd.n5315 vss 0.00271f
C7923 vdd.n5316 vss 0.008f
C7924 vdd.n5317 vss 0.008f
C7925 vdd.n5318 vss 0.0105f
C7926 vdd.n5320 vss 0.00851f
C7927 vdd.n5322 vss 0.00226f
C7928 vdd.n5323 vss 0.00219f
C7929 vdd.n5324 vss 0.008f
C7930 vdd.n5325 vss 0.008f
C7931 vdd.n5326 vss 0.00271f
C7932 vdd.n5327 vss 0.00284f
C7933 vdd.n5328 vss 0.00658f
C7934 vdd.n5329 vss 0.00542f
C7935 vdd.n5330 vss 0.00748f
C7936 vdd.n5331 vss 0.00335f
C7937 vdd.n5332 vss 0.00271f
C7938 vdd.n5333 vss 0.00359f
C7939 vdd.n5334 vss 0.0115f
C7940 vdd.n5335 vss 0.0186f
C7941 vdd.n5336 vss 0.00319f
C7942 vdd.n5337 vss 0.00638f
C7943 vdd.n5338 vss 0.00385f
C7944 vdd.n5339 vss 2.66e-19
C7945 vdd.n5340 vss -0.0638f
C7946 vdd.n5341 vss 0.0115f
C7947 vdd.n5342 vss 0.00385f
C7948 vdd.n5343 vss 0.00359f
C7949 vdd.n5344 vss 0.0111f
C7950 vdd.n5345 vss 0.0115f
C7951 vdd.n5346 vss 0.049f
C7952 vdd.n5347 vss 0.0198f
C7953 vdd.n5348 vss 0.00399f
C7954 vdd.n5349 vss 0.0205f
C7955 vdd.n5350 vss 0.00335f
C7956 vdd.n5351 vss 0.0241f
C7957 vdd.n5352 vss 0.00284f
C7958 vdd.n5353 vss 2.58e-19
C7959 vdd.n5354 vss 0.00851f
C7960 vdd.n5356 vss 0.00226f
C7961 vdd.n5357 vss 0.0152f
C7962 vdd.n5358 vss 0.0245f
C7963 vdd.n5359 vss 0.0255f
C7964 vdd.n5360 vss 0.0142f
C7965 vdd.n5361 vss 0.00226f
C7966 vdd.n5362 vss 0.00219f
C7967 vdd.n5363 vss 2.58e-19
C7968 vdd.n5364 vss 0.00284f
C7969 vdd.n5365 vss 3.87e-19
C7970 vdd.n5366 vss 0.00399f
C7971 vdd.n5367 vss 0.00651f
C7972 vdd.n5368 vss -0.143f
C7973 vdd.n5369 vss 0.0182f
C7974 vdd.n5370 vss 0.0111f
C7975 vdd.n5371 vss 0.00359f
C7976 vdd.n5372 vss 0.00385f
C7977 vdd.n5373 vss 0.00477f
C7978 vdd.n5374 vss 0.00658f
C7979 vdd.n5375 vss 0.00542f
C7980 vdd.n5376 vss 0.00271f
C7981 vdd.n5377 vss 0.008f
C7982 vdd.n5378 vss 0.008f
C7983 vdd.n5379 vss 0.0105f
C7984 vdd.n5381 vss 0.00226f
C7985 vdd.n5383 vss 0.00851f
C7986 vdd.n5384 vss 2.58e-19
C7987 vdd.n5385 vss 0.00284f
C7988 vdd.n5386 vss 3.87e-19
C7989 vdd.n5387 vss 0.00399f
C7990 vdd.n5388 vss 0.00651f
C7991 vdd.n5389 vss 0.0186f
C7992 vdd.n5390 vss 0.0182f
C7993 vdd.n5391 vss 0.0111f
C7994 vdd.n5392 vss 0.00306f
C7995 vdd.n5393 vss 0.0115f
C7996 vdd.n5394 vss 0.0182f
C7997 vdd.n5395 vss 0.0186f
C7998 vdd.n5396 vss 0.00651f
C7999 vdd.n5397 vss 0.00399f
C8000 vdd.n5398 vss 0.00284f
C8001 vdd.n5399 vss 3.87e-19
C8002 vdd.n5400 vss 0.00271f
C8003 vdd.n5401 vss -0.0615f
C8004 vdd.n5402 vss -0.173f
C8005 vdd.n5403 vss 0.00477f
C8006 vdd.n5404 vss 0.00658f
C8007 vdd.n5405 vss 0.00542f
C8008 vdd.n5406 vss 0.00271f
C8009 vdd.n5407 vss 0.008f
C8010 vdd.n5408 vss 0.008f
C8011 vdd.n5409 vss 0.00219f
C8012 vdd.n5410 vss 0.00226f
C8013 vdd.n5412 vss 0.00851f
C8014 vdd.n5414 vss 0.0105f
C8015 vdd.n5415 vss 0.008f
C8016 vdd.n5416 vss 0.008f
C8017 vdd.n5417 vss 0.00271f
C8018 vdd.n5418 vss 0.00542f
C8019 vdd.n5419 vss 0.00658f
C8020 vdd.n5420 vss 0.00477f
C8021 vdd.n5421 vss 0.00335f
C8022 vdd.n5422 vss 0.00271f
C8023 vdd.n5423 vss 0.00359f
C8024 vdd.n5424 vss 2.66e-19
C8025 vdd.n5425 vss 0.00399f
C8026 vdd.n5426 vss 0.00651f
C8027 vdd.n5427 vss -0.143f
C8028 vdd.n5428 vss 0.0182f
C8029 vdd.n5429 vss 0.0111f
C8030 vdd.n5430 vss 0.00359f
C8031 vdd.n5431 vss 0.00385f
C8032 vdd.n5432 vss 0.00477f
C8033 vdd.n5433 vss 0.00542f
C8034 vdd.n5434 vss 0.00658f
C8035 vdd.n5435 vss 0.00284f
C8036 vdd.n5436 vss 0.00219f
C8037 vdd.n5437 vss 0.00284f
C8038 vdd.n5438 vss 2.58e-19
C8039 vdd.n5439 vss 0.00851f
C8040 vdd.n5441 vss 0.0105f
C8041 vdd.n5443 vss 0.00226f
C8042 vdd.n5444 vss 0.00219f
C8043 vdd.n5445 vss 2.58e-19
C8044 vdd.n5446 vss 0.00284f
C8045 vdd.n5447 vss 3.87e-19
C8046 vdd.n5448 vss 0.00399f
C8047 vdd.n5449 vss 0.00651f
C8048 vdd.n5450 vss 0.0186f
C8049 vdd.n5451 vss 0.0182f
C8050 vdd.n5452 vss 0.0111f
C8051 vdd.n5453 vss -0.0615f
C8052 vdd.n5454 vss -0.173f
C8053 vdd.n5455 vss 0.00477f
C8054 vdd.n5456 vss 0.00658f
C8055 vdd.n5457 vss 0.00542f
C8056 vdd.n5458 vss 0.00271f
C8057 vdd.n5459 vss 0.008f
C8058 vdd.n5460 vss 0.008f
C8059 vdd.n5461 vss 0.0105f
C8060 vdd.n5463 vss 0.00226f
C8061 vdd.n5464 vss 0.0193f
C8062 vdd.n5465 vss 2.58e-19
C8063 vdd.n5466 vss 0.00284f
C8064 vdd.n5467 vss 3.87e-19
C8065 vdd.n5468 vss 0.00399f
C8066 vdd.n5469 vss 0.0234f
C8067 vdd.n5470 vss 0.0657f
C8068 vdd.n5471 vss 0.0654f
C8069 vdd.n5472 vss 0.0111f
C8070 vdd.n5473 vss 2.66e-19
C8071 vdd.n5474 vss 0.00385f
C8072 vdd.n5475 vss 0.00271f
C8073 vdd.n5476 vss 3.87e-19
C8074 vdd.n5477 vss 0.00284f
C8075 vdd.n5478 vss 2.58e-19
C8076 vdd.n5479 vss 0.0193f
C8077 vdd.n5481 vss 0.00226f
C8078 vdd.n5482 vss 0.00219f
C8079 vdd.n5483 vss 0.008f
C8080 vdd.n5484 vss 0.008f
C8081 vdd.n5485 vss 0.00271f
C8082 vdd.n5486 vss 0.00542f
C8083 vdd.n5487 vss 0.00658f
C8084 vdd.n5488 vss 0.00477f
C8085 vdd.n5489 vss -0.173f
C8086 vdd.n5490 vss 0.00319f
C8087 vdd.n5491 vss 0.0186f
C8088 vdd.n5492 vss 0.0182f
C8089 vdd.n5493 vss 0.0115f
C8090 vdd.n5494 vss 0.0111f
C8091 vdd.n5495 vss 2.66e-19
C8092 vdd.n5496 vss 0.00385f
C8093 vdd.n5497 vss 0.00271f
C8094 vdd.n5498 vss 3.87e-19
C8095 vdd.n5499 vss 0.00284f
C8096 vdd.n5500 vss 2.58e-19
C8097 vdd.n5501 vss 0.00851f
C8098 vdd.n5503 vss 0.00226f
C8099 vdd.n5504 vss 0.0105f
C8100 vdd.n5506 vss 0.00851f
C8101 vdd.n5507 vss 2.58e-19
C8102 vdd.n5508 vss 0.00219f
C8103 vdd.n5509 vss 0.008f
C8104 vdd.n5510 vss 0.00271f
C8105 vdd.n5511 vss 0.00542f
C8106 vdd.n5512 vss 0.00658f
C8107 vdd.n5513 vss 0.00477f
C8108 vdd.n5514 vss 0.00399f
C8109 vdd.n5515 vss 0.00319f
C8110 vdd.n5516 vss 0.00385f
C8111 vdd.n5517 vss 0.00638f
C8112 vdd.n5518 vss -0.148f
C8113 vdd.n5519 vss -0.0638f
C8114 vdd.n5520 vss 0.0182f
C8115 vdd.n5521 vss 0.00385f
C8116 vdd.n5522 vss 0.00638f
C8117 vdd.n5523 vss 0.00319f
C8118 vdd.n5524 vss 0.0186f
C8119 vdd.n5525 vss 0.0115f
C8120 vdd.n5526 vss 0.00359f
C8121 vdd.n5527 vss 0.00271f
C8122 vdd.n5528 vss 0.00335f
C8123 vdd.n5529 vss 0.00748f
C8124 vdd.n5530 vss 0.00542f
C8125 vdd.n5531 vss 0.00658f
C8126 vdd.n5532 vss 0.00284f
C8127 vdd.n5533 vss 0.00219f
C8128 vdd.n5534 vss 0.00219f
C8129 vdd.n5535 vss 2.58e-19
C8130 vdd.n5536 vss 0.00851f
C8131 vdd.n5538 vss 0.00226f
C8132 vdd.n5540 vss 0.0105f
C8133 vdd.n5541 vss 0.008f
C8134 vdd.n5542 vss 0.008f
C8135 vdd.n5543 vss 0.00271f
C8136 vdd.n5544 vss 0.00284f
C8137 vdd.n5545 vss 0.00658f
C8138 vdd.n5546 vss 0.00542f
C8139 vdd.n5547 vss 0.00748f
C8140 vdd.n5548 vss 0.00335f
C8141 vdd.n5549 vss 0.00271f
C8142 vdd.n5550 vss -0.0615f
C8143 vdd.n5551 vss 0.0115f
C8144 vdd.n5552 vss 0.0186f
C8145 vdd.n5553 vss 0.00319f
C8146 vdd.n5554 vss 0.00638f
C8147 vdd.n5555 vss 0.00385f
C8148 vdd.n5556 vss 2.66e-19
C8149 vdd.n5557 vss 0.0111f
C8150 vdd.n5558 vss 0.0115f
C8151 vdd.n5559 vss 0.00385f
C8152 vdd.n5560 vss 2.66e-19
C8153 vdd.n5561 vss -0.0638f
C8154 vdd.n5562 vss -0.148f
C8155 vdd.n5563 vss 0.0186f
C8156 vdd.n5564 vss 0.00319f
C8157 vdd.n5565 vss 0.00399f
C8158 vdd.n5566 vss 0.00477f
C8159 vdd.n5567 vss 0.00335f
C8160 vdd.n5568 vss 0.00748f
C8161 vdd.n5569 vss 0.00284f
C8162 vdd.n5570 vss 2.58e-19
C8163 vdd.n5571 vss 0.00219f
C8164 vdd.n5572 vss 0.00226f
C8165 vdd.n5574 vss 0.0105f
C8166 vdd.n5575 vss 0.0226f
C8167 vdd.n5576 vss 0.0361f
C8168 vdd.n5577 vss 0.0344f
C8169 vdd.n5578 vss 0.0318f
C8170 vdd.n5579 vss 0.0325f
C8171 vdd.n5580 vss 0.0491f
C8172 vdd.n5581 vss 3f
C8173 vdd.n5582 vss 3.05f
C8174 vdd.n5583 vss 0.0515f
C8175 vdd.n5584 vss 0.0358f
C8176 vdd.n5585 vss 0.0354f
C8177 vdd.n5586 vss 0.00477f
C8178 vdd.n5587 vss 0.00271f
C8179 vdd.n5588 vss 0.00284f
C8180 vdd.n5589 vss 0.00658f
C8181 vdd.n5590 vss 0.00542f
C8182 vdd.n5591 vss 0.00781f
C8183 vdd.n5592 vss 0.00335f
C8184 vdd.n5593 vss 0.00271f
C8185 vdd.n5594 vss -0.0615f
C8186 vdd.n5595 vss 0.0117f
C8187 vdd.n5596 vss 0.0189f
C8188 vdd.n5597 vss 0.00319f
C8189 vdd.n5598 vss 0.00638f
C8190 vdd.n5599 vss 0.00385f
C8191 vdd.n5600 vss 2.66e-19
C8192 vdd.n5601 vss 0.0113f
C8193 vdd.n5602 vss 0.0117f
C8194 vdd.n5603 vss 0.0117f
C8195 vdd.n5604 vss 0.00385f
C8196 vdd.n5605 vss 0.00399f
C8197 vdd.n5606 vss 3.87e-19
C8198 vdd.n5607 vss 0.00477f
C8199 vdd.n5608 vss 0.00284f
C8200 vdd.n5609 vss 0.00271f
C8201 vdd.n5610 vss 3.87e-19
C8202 vdd.n5611 vss 0.00284f
C8203 vdd.n5612 vss 0.008f
C8204 vdd.n5613 vss 0.008f
C8205 vdd.n5614 vss 0.00271f
C8206 vdd.n5615 vss 0.00284f
C8207 vdd.n5616 vss 0.00219f
C8208 vdd.n5617 vss 0.00219f
C8209 vdd.n5618 vss 0.00851f
C8210 vdd.n5619 vss 2.58e-19
C8211 vdd.n5620 vss 0.00226f
C8212 vdd.n5621 vss 0.00219f
C8213 vdd.n5622 vss 0.008f
C8214 vdd.n5623 vss 0.008f
C8215 vdd.n5624 vss 0.00219f
C8216 vdd.n5625 vss 0.00542f
C8217 vdd.n5626 vss 0.00284f
C8218 vdd.n5627 vss 0.00658f
C8219 vdd.n5628 vss 0.00271f
C8220 vdd.n5629 vss 0.00638f
C8221 vdd.n5630 vss 0.00359f
C8222 vdd.n5631 vss 0.0117f
C8223 vdd.n5632 vss 0.00385f
C8224 vdd.n5633 vss 0.0189f
C8225 vdd.n5634 vss 0.00319f
C8226 vdd.n5635 vss 0.00638f
C8227 vdd.n5636 vss 0.0185f
C8228 vdd.n5637 vss 0.0113f
C8229 vdd.n5638 vss 2.66e-19
C8230 vdd.n5639 vss -0.0615f
C8231 vdd.n5640 vss 0.00271f
C8232 vdd.n5641 vss 0.00748f
C8233 vdd.n5642 vss 0.00335f
C8234 vdd.n5643 vss 0.00477f
C8235 vdd.n5644 vss -0.173f
C8236 vdd.n5645 vss 0.00319f
C8237 vdd.n5646 vss 0.0189f
C8238 vdd.n5647 vss 0.0185f
C8239 vdd.n5648 vss -0.148f
C8240 vdd.n5649 vss 0.00399f
C8241 vdd.n5650 vss 2.66e-19
C8242 vdd.n5651 vss 0.00284f
C8243 vdd.n5652 vss 0.00335f
C8244 vdd.n5653 vss 0.00637f
C8245 vdd.n5654 vss 0.00399f
C8246 vdd.n5655 vss -0.0637f
C8247 vdd.n5656 vss 0.0249f
C8248 vdd.n5657 vss 0.00504f
C8249 vdd.n5658 vss 0.00667f
C8250 vdd.n5659 vss 0.00626f
C8251 vdd.n5660 vss 0.0249f
C8252 vdd.n5661 vss 0.0117f
C8253 vdd.n5662 vss 0.00359f
C8254 vdd.n5663 vss 0.00271f
C8255 vdd.n5664 vss 0.00219f
C8256 vdd.n5665 vss 0.00851f
C8257 vdd.n5666 vss 2.58e-19
C8258 vdd.n5667 vss 0.00219f
C8259 vdd.n5668 vss 0.00226f
C8260 vdd.n5669 vss 0.0105f
C8261 vdd.n5670 vss 0.008f
C8262 vdd.n5671 vss 0.00748f
C8263 vdd.n5672 vss 0.00335f
C8264 vdd.n5673 vss 0.00477f
C8265 vdd.n5674 vss 0.00658f
C8266 vdd.n5675 vss 0.00542f
C8267 vdd.n5676 vss 0.00271f
C8268 vdd.n5677 vss 0.008f
C8269 vdd.n5678 vss 0.00219f
C8270 vdd.n5679 vss 0.00851f
C8271 vdd.n5680 vss 2.58e-19
C8272 vdd.n5681 vss 0.00284f
C8273 vdd.n5682 vss 3.87e-19
C8274 vdd.n5683 vss 0.00385f
C8275 vdd.n5684 vss 0.00638f
C8276 vdd.n5685 vss 0.00319f
C8277 vdd.n5686 vss 0.0189f
C8278 vdd.n5687 vss 0.0117f
C8279 vdd.n5688 vss 0.0113f
C8280 vdd.n5689 vss 2.66e-19
C8281 vdd.n5690 vss 0.00385f
C8282 vdd.n5691 vss 3.87e-19
C8283 vdd.n5692 vss 0.00284f
C8284 vdd.n5693 vss 0.00219f
C8285 vdd.n5694 vss 0.00271f
C8286 vdd.n5695 vss 0.008f
C8287 vdd.n5696 vss 0.008f
C8288 vdd.n5697 vss 0.00226f
C8289 vdd.n5698 vss 0.00219f
C8290 vdd.n5699 vss 0.00851f
C8291 vdd.n5700 vss 2.58e-19
C8292 vdd.n5701 vss 0.00219f
C8293 vdd.n5702 vss 0.00219f
C8294 vdd.n5703 vss 0.00284f
C8295 vdd.n5704 vss 0.00658f
C8296 vdd.n5705 vss 0.00542f
C8297 vdd.n5706 vss 0.00748f
C8298 vdd.n5707 vss 0.00335f
C8299 vdd.n5708 vss 0.00271f
C8300 vdd.n5709 vss 0.00359f
C8301 vdd.n5710 vss 2.66e-19
C8302 vdd.n5711 vss -0.0637f
C8303 vdd.n5712 vss -0.148f
C8304 vdd.n5713 vss 0.0189f
C8305 vdd.n5714 vss 0.00319f
C8306 vdd.n5715 vss 0.00399f
C8307 vdd.n5716 vss 0.00477f
C8308 vdd.n5717 vss 0.00335f
C8309 vdd.n5718 vss 0.00748f
C8310 vdd.n5719 vss 0.00284f
C8311 vdd.n5720 vss 2.58e-19
C8312 vdd.n5721 vss 0.00851f
C8313 vdd.n5722 vss 0.0105f
C8314 vdd.n5723 vss 0.008f
C8315 vdd.n5724 vss 0.00219f
C8316 vdd.n5725 vss 0.0257f
C8317 vdd.n5726 vss 0.0193f
C8318 vdd.n5727 vss 0.376f
C8319 vdd.n5728 vss 0.0142f
C8320 vdd.n5729 vss 0.00832f
C8321 vdd.n5730 vss 0.0517f
C8322 vdd.t87 vss 0.00477f
C8323 vdd.n5731 vss 0.0473f
C8324 vdd.n5732 vss 0.0295f
C8325 vdd.n5733 vss 0.0142f
C8326 vdd.n5734 vss 8.67e-19
C8327 vdd.n5735 vss 0.0136f
C8328 vdd.n5736 vss 2.85f
C8329 vdd.n5737 vss 2.86f
C8330 vdd.n5738 vss 0.0427f
C8331 vdd.n5739 vss 0.00887f
C8332 vdd.n5740 vss 0.00518f
C8333 vdd.n5741 vss 0.0163f
C8334 vdd.n5742 vss 0.00668f
C8335 vdd.n5743 vss 0.0664f
C8336 vdd.n5744 vss 0.00673f
C8337 vdd.n5745 vss 0.0163f
C8338 vdd.n5746 vss 0.0882f
C8339 vdd.n5747 vss 0.209f
C8340 vdd.n5748 vss 0.0101f
C8341 vdd.n5749 vss 6.66e-19
C8342 vdd.n5750 vss 0.0162f
C8343 vdd.n5751 vss 0.0141f
C8344 vdd.n5752 vss 0.0458f
C8345 vdd.n5753 vss 0.00651f
C8346 vdd.n5754 vss 0.00869f
C8347 vdd.n5755 vss 0.00893f
C8348 vdd.n5756 vss 0.00319f
C8349 vdd.n5757 vss 0.015f
C8350 vdd.n5758 vss 0.00333f
C8351 vdd.n5759 vss 0.00563f
C8352 vdd.n5760 vss 0.0163f
C8353 vdd.n5761 vss 0.00903f
C8354 vdd.n5762 vss 0.0328f
C8355 vdd.n5763 vss 0.0157f
C8356 vdd.n5764 vss 0.014f
C8357 vdd.n5765 vss 0.00642f
C8358 vdd.n5766 vss 0.0137f
C8359 vdd.n5767 vss 0.00541f
C8360 vdd.t92 vss 0.00542f
C8361 vdd.t91 vss 0.00542f
C8362 vdd.n5768 vss 0.0133f
C8363 vdd.n5769 vss 0.0394f
C8364 vdd.n5770 vss 0.00658f
C8365 vdd.n5771 vss 0.0134f
C8366 vdd.n5772 vss 0.0818f
C8367 vdd.n5773 vss 0.0163f
C8368 vdd.n5774 vss 0.0131f
C8369 vdd.n5775 vss 0.00887f
C8370 vdd.n5776 vss 0.00518f
C8371 vdd.n5777 vss 1.69f
C8372 vdd.n5778 vss 0.0635f
C8373 vdd.n5779 vss 0.0163f
C8374 vdd.n5780 vss 0.0163f
C8375 vdd.n5781 vss 0.0482f
C8376 vdd.n5782 vss 0.00673f
C8377 vdd.n5783 vss 0.0664f
C8378 vdd.n5784 vss 0.00668f
C8379 vdd.n5785 vss 0.00518f
C8380 vdd.n5786 vss 0.00887f
C8381 vdd.n5787 vss 0.0547f
C8382 vdd.n5788 vss 0.0163f
C8383 vdd.n5789 vss 0.00673f
C8384 vdd.t82 vss 1.36f
C8385 vdd.n5790 vss 0.00832f
C8386 vdd.t76 vss 0.00477f
C8387 vdd.n5791 vss 0.0129f
C8388 vdd.n5792 vss 0.00994f
C8389 vdd.n5793 vss 0.00908f
C8390 vdd.n5794 vss 0.0249f
C8391 vdd.n5795 vss 0.00359f
C8392 vdd.n5796 vss 0.00284f
C8393 vdd.n5797 vss 0.00385f
C8394 vdd.n5798 vss 0.00219f
C8395 vdd.n5799 vss 0.00219f
C8396 vdd.n5800 vss 0.00247f
C8397 vdd.n5801 vss 0.00226f
C8398 vdd.n5802 vss 0.0142f
C8399 vdd.n5803 vss 0.00673f
C8400 vdd.n5804 vss 0.0163f
C8401 vdd.n5805 vss 0.0635f
C8402 vdd.n5806 vss 0.0163f
C8403 vdd.n5807 vss 0.00887f
C8404 vdd.n5808 vss 0.00518f
C8405 vdd.n5809 vss 0.00668f
C8406 vdd.n5810 vss 0.0664f
C8407 vdd.n5811 vss 0.385f
C8408 vdd.t75 vss 0.206f
C8409 vdd.n5812 vss 0.376f
C8410 vdd.n5813 vss 0.00226f
C8411 vdd.n5814 vss 0.00219f
C8412 vdd.n5815 vss 0.00748f
C8413 vdd.n5816 vss 0.00335f
C8414 vdd.n5817 vss 0.00359f
C8415 vdd.n5818 vss 0.00638f
C8416 vdd.n5819 vss 0.0185f
C8417 vdd.n5820 vss 0.00638f
C8418 vdd.n5821 vss 0.00284f
C8419 vdd.n5822 vss 0.00271f
C8420 vdd.n5823 vss 0.00219f
C8421 vdd.n5824 vss 0.00219f
C8422 vdd.n5825 vss 0.00226f
C8423 vdd.n5826 vss 0.00219f
C8424 vdd.n5827 vss 0.00748f
C8425 vdd.n5828 vss 0.00335f
C8426 vdd.n5829 vss -0.0615f
C8427 vdd.n5830 vss 0.0185f
C8428 vdd.n5831 vss 0.00638f
C8429 vdd.n5832 vss 0.00284f
C8430 vdd.n5833 vss 0.00271f
C8431 vdd.n5834 vss 0.00219f
C8432 vdd.n5835 vss 0.00219f
C8433 vdd.n5836 vss 0.00226f
C8434 vdd.n5837 vss 0.00219f
C8435 vdd.n5838 vss 0.00748f
C8436 vdd.n5839 vss 0.00335f
C8437 vdd.n5840 vss 0.00359f
C8438 vdd.n5841 vss -0.148f
C8439 vdd.n5842 vss 0.00638f
C8440 vdd.n5843 vss 0.00284f
C8441 vdd.n5844 vss 0.00271f
C8442 vdd.n5845 vss 0.00219f
C8443 vdd.n5846 vss 0.00219f
C8444 vdd.n5847 vss 0.00226f
C8445 vdd.n5848 vss 0.00219f
C8446 vdd.n5849 vss 0.00748f
C8447 vdd.n5850 vss 0.00335f
C8448 vdd.n5851 vss 0.00359f
C8449 vdd.n5852 vss 0.0185f
C8450 vdd.n5853 vss 0.00638f
C8451 vdd.n5854 vss 0.00284f
C8452 vdd.n5855 vss 0.00271f
C8453 vdd.n5856 vss 0.00219f
C8454 vdd.n5857 vss 0.00219f
C8455 vdd.n5859 vss 0.00219f
C8456 vdd.n5860 vss 0.00776f
C8457 vdd.n5861 vss 0.00335f
C8458 vdd.n5862 vss -0.0615f
C8459 vdd.n5863 vss 0.0115f
C8460 vdd.n5864 vss 0.00359f
C8461 vdd.n5865 vss 0.00271f
C8462 vdd.n5866 vss 0.00219f
C8463 vdd.n5867 vss 3.87e-19
C8464 vdd.n5868 vss 0.00219f
C8465 vdd.n5869 vss 0.00226f
C8466 vdd.n5870 vss 0.00219f
C8467 vdd.n5871 vss 0.00748f
C8468 vdd.n5872 vss 0.00335f
C8469 vdd.n5873 vss 0.00359f
C8470 vdd.n5874 vss 0.00638f
C8471 vdd.n5875 vss 0.0182f
C8472 vdd.n5876 vss 0.00638f
C8473 vdd.n5877 vss 0.00284f
C8474 vdd.n5878 vss 0.00271f
C8475 vdd.n5879 vss 0.00219f
C8476 vdd.n5880 vss 0.00219f
C8477 vdd.n5881 vss 0.008f
C8478 vdd.n5882 vss 0.00851f
C8479 vdd.n5883 vss 0.00219f
C8480 vdd.n5884 vss 0.00219f
C8481 vdd.n5885 vss 3.87e-19
C8482 vdd.n5886 vss 0.008f
C8483 vdd.n5887 vss 0.00271f
C8484 vdd.n5888 vss 0.00542f
C8485 vdd.n5889 vss 0.00271f
C8486 vdd.n5890 vss 0.00658f
C8487 vdd.n5891 vss -0.0615f
C8488 vdd.n5892 vss 0.0182f
C8489 vdd.n5893 vss 0.00399f
C8490 vdd.n5894 vss -0.0638f
C8491 vdd.n5895 vss 2.66e-19
C8492 vdd.n5896 vss 3.87e-19
C8493 vdd.n5897 vss 0.00477f
C8494 vdd.n5898 vss 0.00284f
C8495 vdd.n5899 vss 0.00219f
C8496 vdd.n5900 vss 0.0105f
C8497 vdd.n5901 vss 0.008f
C8498 vdd.n5902 vss 0.00271f
C8499 vdd.n5903 vss 0.00477f
C8500 vdd.n5904 vss 0.00284f
C8501 vdd.n5905 vss 3.87e-19
C8502 vdd.n5906 vss 2.66e-19
C8503 vdd.n5907 vss 0.00399f
C8504 vdd.n5908 vss 0.0186f
C8505 vdd.n5909 vss -0.0615f
C8506 vdd.n5910 vss 0.00335f
C8507 vdd.n5911 vss 0.00284f
C8508 vdd.n5912 vss 0.00748f
C8509 vdd.n5913 vss 0.00219f
C8510 vdd.n5914 vss 0.008f
C8511 vdd.n5915 vss 0.008f
C8512 vdd.n5916 vss 0.00219f
C8513 vdd.n5917 vss 0.00219f
C8514 vdd.n5918 vss 0.00219f
C8515 vdd.n5919 vss 0.00219f
C8516 vdd.n5920 vss 0.00284f
C8517 vdd.n5921 vss 0.0233f
C8518 vdd.n5922 vss 0.0115f
C8519 vdd.n5923 vss 2.66e-19
C8520 vdd.n5924 vss 0.00271f
C8521 vdd.n5925 vss 0.00284f
C8522 vdd.n5926 vss 0.00748f
C8523 vdd.n5927 vss 0.00219f
C8524 vdd.n5928 vss 0.00219f
C8525 vdd.n5929 vss 0.024f
C8526 vdd.n5930 vss 0.00271f
C8527 vdd.n5931 vss 0.0213f
C8528 vdd.n5932 vss 0.0234f
C8529 vdd.n5933 vss 0.0234f
C8530 vdd.n5934 vss 0.0213f
C8531 vdd.n5935 vss 0.00271f
C8532 vdd.n5936 vss 0.024f
C8533 vdd.n5937 vss 0.00219f
C8534 vdd.n5939 vss 0.00219f
C8535 vdd.n5940 vss 0.00219f
C8536 vdd.n5941 vss 0.00284f
C8537 vdd.n5942 vss 0.00335f
C8538 vdd.n5943 vss 0.00306f
C8539 vdd.n5944 vss 0.0115f
C8540 vdd.n5945 vss 2.66e-19
C8541 vdd.n5946 vss 0.00271f
C8542 vdd.n5947 vss 0.00748f
C8543 vdd.n5948 vss 0.00219f
C8544 vdd.n5949 vss 0.00851f
C8545 vdd.n5950 vss 0.00219f
C8546 vdd.n5951 vss 0.00219f
C8547 vdd.n5952 vss 0.00284f
C8548 vdd.n5953 vss 0.00335f
C8549 vdd.n5954 vss 0.00306f
C8550 vdd.n5955 vss -0.069f
C8551 vdd.n5956 vss 2.66e-19
C8552 vdd.n5957 vss 0.00271f
C8553 vdd.n5958 vss 0.00748f
C8554 vdd.n5959 vss 0.008f
C8555 vdd.n5960 vss 0.00226f
C8556 vdd.n5961 vss 0.00219f
C8557 vdd.n5962 vss 0.00219f
C8558 vdd.n5963 vss 0.00748f
C8559 vdd.n5964 vss 3.87e-19
C8560 vdd.n5965 vss 0.008f
C8561 vdd.n5966 vss 0.00271f
C8562 vdd.n5967 vss 0.00335f
C8563 vdd.n5968 vss 0.00306f
C8564 vdd.n5969 vss 0.0115f
C8565 vdd.n5970 vss -0.173f
C8566 vdd.n5971 vss 0.0111f
C8567 vdd.n5972 vss 0.00284f
C8568 vdd.n5973 vss 0.00219f
C8569 vdd.n5974 vss 0.00219f
C8570 vdd.n5975 vss 0.00226f
C8571 vdd.n5976 vss 0.00219f
C8572 vdd.n5977 vss 0.00748f
C8573 vdd.n5978 vss 0.00271f
C8574 vdd.n5979 vss 2.66e-19
C8575 vdd.n5980 vss 0.00306f
C8576 vdd.n5981 vss 0.0182f
C8577 vdd.n5982 vss 0.00306f
C8578 vdd.n5983 vss 0.00284f
C8579 vdd.n5984 vss 0.00219f
C8580 vdd.n5985 vss 0.00219f
C8581 vdd.n5986 vss 0.00226f
C8582 vdd.n5987 vss 0.00219f
C8583 vdd.n5988 vss 0.0241f
C8584 vdd.n5989 vss 0.00271f
C8585 vdd.n5990 vss 2.66e-19
C8586 vdd.n5991 vss 0.0115f
C8587 vdd.n5992 vss 0.0197f
C8588 vdd.n5993 vss 0.00335f
C8589 vdd.n5994 vss 0.00359f
C8590 vdd.n5995 vss -0.148f
C8591 vdd.n5996 vss 0.00638f
C8592 vdd.n5997 vss 0.00284f
C8593 vdd.n5998 vss 0.00271f
C8594 vdd.n5999 vss 0.00219f
C8595 vdd.n6000 vss 0.0241f
C8596 vdd.n6001 vss 0.00219f
C8597 vdd.n6002 vss 0.00219f
C8598 vdd.n6003 vss 0.00226f
C8599 vdd.n6004 vss 0.00219f
C8600 vdd.n6005 vss 0.00748f
C8601 vdd.n6006 vss 0.00335f
C8602 vdd.n6007 vss 0.00359f
C8603 vdd.n6008 vss 0.0182f
C8604 vdd.n6009 vss 0.00638f
C8605 vdd.n6010 vss 0.00284f
C8606 vdd.n6011 vss 0.00271f
C8607 vdd.n6012 vss 0.00219f
C8608 vdd.n6013 vss 0.00219f
C8609 vdd.n6014 vss 0.008f
C8610 vdd.n6015 vss 0.00851f
C8611 vdd.n6016 vss 0.00219f
C8612 vdd.n6017 vss 0.00219f
C8613 vdd.n6018 vss 3.87e-19
C8614 vdd.n6019 vss 0.008f
C8615 vdd.n6020 vss 0.00271f
C8616 vdd.n6021 vss 0.00542f
C8617 vdd.n6022 vss 0.00271f
C8618 vdd.n6023 vss 0.00658f
C8619 vdd.n6024 vss -0.0615f
C8620 vdd.n6025 vss 0.0182f
C8621 vdd.n6026 vss 0.00399f
C8622 vdd.n6027 vss -0.0638f
C8623 vdd.n6028 vss 2.66e-19
C8624 vdd.n6029 vss 3.87e-19
C8625 vdd.n6030 vss 0.00477f
C8626 vdd.n6031 vss 0.00284f
C8627 vdd.n6032 vss 0.00219f
C8628 vdd.n6033 vss 0.0105f
C8629 vdd.n6034 vss 0.008f
C8630 vdd.n6035 vss 0.00271f
C8631 vdd.n6036 vss 0.00477f
C8632 vdd.n6037 vss 0.00284f
C8633 vdd.n6038 vss 3.87e-19
C8634 vdd.n6039 vss 2.66e-19
C8635 vdd.n6040 vss 0.00399f
C8636 vdd.n6041 vss 0.0186f
C8637 vdd.n6042 vss -0.0615f
C8638 vdd.n6043 vss 0.00335f
C8639 vdd.n6044 vss 0.00284f
C8640 vdd.n6045 vss 0.00748f
C8641 vdd.n6046 vss 0.00219f
C8642 vdd.n6047 vss 0.008f
C8643 vdd.n6048 vss 0.008f
C8644 vdd.n6049 vss 0.00219f
C8645 vdd.n6050 vss 0.00219f
C8646 vdd.n6051 vss 0.00219f
C8647 vdd.n6052 vss 0.00219f
C8648 vdd.n6053 vss 0.00284f
C8649 vdd.n6054 vss 0.0233f
C8650 vdd.n6055 vss 0.0115f
C8651 vdd.n6056 vss 2.66e-19
C8652 vdd.n6057 vss 0.00271f
C8653 vdd.n6058 vss 0.00284f
C8654 vdd.n6059 vss 0.00748f
C8655 vdd.n6060 vss 0.00219f
C8656 vdd.n6061 vss 0.00219f
C8657 vdd.n6062 vss 0.024f
C8658 vdd.n6063 vss 0.00271f
C8659 vdd.n6064 vss 0.0213f
C8660 vdd.n6065 vss 0.0234f
C8661 vdd.n6066 vss 0.0234f
C8662 vdd.n6067 vss 0.0213f
C8663 vdd.n6068 vss 0.00271f
C8664 vdd.n6069 vss 0.024f
C8665 vdd.n6070 vss 0.00219f
C8666 vdd.n6072 vss 0.00219f
C8667 vdd.n6073 vss 0.00219f
C8668 vdd.n6074 vss 0.00284f
C8669 vdd.n6075 vss 0.00335f
C8670 vdd.n6076 vss 0.00306f
C8671 vdd.n6077 vss 0.0115f
C8672 vdd.n6078 vss 2.66e-19
C8673 vdd.n6079 vss 0.00271f
C8674 vdd.n6080 vss 0.00748f
C8675 vdd.n6081 vss 0.00219f
C8676 vdd.n6082 vss 0.00851f
C8677 vdd.n6083 vss 0.00219f
C8678 vdd.n6084 vss 0.00219f
C8679 vdd.n6085 vss 0.00284f
C8680 vdd.n6086 vss 0.00335f
C8681 vdd.n6087 vss 0.00306f
C8682 vdd.n6088 vss -0.069f
C8683 vdd.n6089 vss 2.66e-19
C8684 vdd.n6090 vss 0.00271f
C8685 vdd.n6091 vss 0.00748f
C8686 vdd.n6092 vss 0.008f
C8687 vdd.n6093 vss 0.00226f
C8688 vdd.n6094 vss 0.00219f
C8689 vdd.n6095 vss 0.00219f
C8690 vdd.n6096 vss 0.00748f
C8691 vdd.n6097 vss 3.87e-19
C8692 vdd.n6098 vss 0.008f
C8693 vdd.n6099 vss 0.00271f
C8694 vdd.n6100 vss 0.00335f
C8695 vdd.n6101 vss 0.00306f
C8696 vdd.n6102 vss 0.0115f
C8697 vdd.n6103 vss -0.173f
C8698 vdd.n6104 vss 0.0111f
C8699 vdd.n6105 vss 0.00284f
C8700 vdd.n6106 vss 0.00219f
C8701 vdd.n6107 vss 0.00219f
C8702 vdd.n6108 vss 0.00226f
C8703 vdd.n6109 vss 0.00219f
C8704 vdd.n6110 vss 0.00748f
C8705 vdd.n6111 vss 0.00271f
C8706 vdd.n6112 vss 2.66e-19
C8707 vdd.n6113 vss 0.00306f
C8708 vdd.n6114 vss 0.0182f
C8709 vdd.n6115 vss 0.00306f
C8710 vdd.n6116 vss 0.00284f
C8711 vdd.n6117 vss 0.00219f
C8712 vdd.n6118 vss 0.00219f
C8713 vdd.n6119 vss 0.00226f
C8714 vdd.n6120 vss 0.00219f
C8715 vdd.n6121 vss 0.0241f
C8716 vdd.n6122 vss 0.00271f
C8717 vdd.n6123 vss 2.66e-19
C8718 vdd.n6124 vss 0.0115f
C8719 vdd.n6125 vss 0.0197f
C8720 vdd.n6126 vss 0.00335f
C8721 vdd.n6127 vss 0.00359f
C8722 vdd.n6128 vss -0.148f
C8723 vdd.n6129 vss 0.00638f
C8724 vdd.n6130 vss 0.00284f
C8725 vdd.n6131 vss 0.00271f
C8726 vdd.n6132 vss 0.00219f
C8727 vdd.n6133 vss 0.0241f
C8728 vdd.n6134 vss 0.00219f
C8729 vdd.n6135 vss 0.00219f
C8730 vdd.n6136 vss 0.00226f
C8731 vdd.n6137 vss 0.00219f
C8732 vdd.n6138 vss 0.00748f
C8733 vdd.n6139 vss 0.00335f
C8734 vdd.n6140 vss 0.00359f
C8735 vdd.n6141 vss 0.0182f
C8736 vdd.n6142 vss 0.00638f
C8737 vdd.n6143 vss 0.00284f
C8738 vdd.n6144 vss 0.00271f
C8739 vdd.n6145 vss 0.00219f
C8740 vdd.n6146 vss 0.00219f
C8741 vdd.n6147 vss 0.008f
C8742 vdd.n6148 vss 0.00851f
C8743 vdd.n6149 vss 0.00219f
C8744 vdd.n6150 vss 0.00219f
C8745 vdd.n6151 vss 3.87e-19
C8746 vdd.n6152 vss 0.008f
C8747 vdd.n6153 vss 0.00271f
C8748 vdd.n6154 vss 0.00542f
C8749 vdd.n6155 vss 0.00271f
C8750 vdd.n6156 vss 0.00658f
C8751 vdd.n6157 vss -0.0615f
C8752 vdd.n6158 vss 0.0182f
C8753 vdd.n6159 vss 0.00399f
C8754 vdd.n6160 vss -0.0638f
C8755 vdd.n6161 vss 2.66e-19
C8756 vdd.n6162 vss 3.87e-19
C8757 vdd.n6163 vss 0.00477f
C8758 vdd.n6164 vss 0.00284f
C8759 vdd.n6165 vss 0.00219f
C8760 vdd.n6166 vss 0.0105f
C8761 vdd.n6167 vss 0.008f
C8762 vdd.n6168 vss 0.00271f
C8763 vdd.n6169 vss 0.00477f
C8764 vdd.n6170 vss 0.00284f
C8765 vdd.n6171 vss 3.87e-19
C8766 vdd.n6172 vss 2.66e-19
C8767 vdd.n6173 vss 0.00399f
C8768 vdd.n6174 vss 0.0186f
C8769 vdd.n6175 vss -0.0615f
C8770 vdd.n6176 vss 0.00335f
C8771 vdd.n6177 vss 0.00284f
C8772 vdd.n6178 vss 0.00748f
C8773 vdd.n6179 vss 0.00219f
C8774 vdd.n6180 vss 0.008f
C8775 vdd.n6181 vss 0.008f
C8776 vdd.n6182 vss 0.00219f
C8777 vdd.n6183 vss 0.00219f
C8778 vdd.n6184 vss 0.00219f
C8779 vdd.n6185 vss 0.00219f
C8780 vdd.n6186 vss 0.00284f
C8781 vdd.n6187 vss 0.0233f
C8782 vdd.n6188 vss 0.0115f
C8783 vdd.n6189 vss 2.66e-19
C8784 vdd.n6190 vss 0.00271f
C8785 vdd.n6191 vss 0.00284f
C8786 vdd.n6192 vss 0.00748f
C8787 vdd.n6193 vss 0.00219f
C8788 vdd.n6194 vss 0.00219f
C8789 vdd.n6195 vss 0.024f
C8790 vdd.n6196 vss 0.00271f
C8791 vdd.n6197 vss 0.0213f
C8792 vdd.n6198 vss 0.0234f
C8793 vdd.n6199 vss 0.0234f
C8794 vdd.n6200 vss 0.0213f
C8795 vdd.n6201 vss 0.00271f
C8796 vdd.n6202 vss 0.024f
C8797 vdd.n6203 vss 0.00219f
C8798 vdd.n6205 vss 0.00219f
C8799 vdd.n6206 vss 0.00219f
C8800 vdd.n6207 vss 0.00284f
C8801 vdd.n6208 vss 0.00335f
C8802 vdd.n6209 vss 0.00306f
C8803 vdd.n6210 vss 0.0115f
C8804 vdd.n6211 vss 2.66e-19
C8805 vdd.n6212 vss 0.00271f
C8806 vdd.n6213 vss 0.00748f
C8807 vdd.n6214 vss 0.00219f
C8808 vdd.n6215 vss 0.00851f
C8809 vdd.n6216 vss 0.00219f
C8810 vdd.n6217 vss 0.00219f
C8811 vdd.n6218 vss 0.00284f
C8812 vdd.n6219 vss 0.00335f
C8813 vdd.n6220 vss 0.00306f
C8814 vdd.n6221 vss -0.069f
C8815 vdd.n6222 vss 2.66e-19
C8816 vdd.n6223 vss 0.00271f
C8817 vdd.n6224 vss 0.00748f
C8818 vdd.n6225 vss 0.008f
C8819 vdd.n6226 vss 0.00226f
C8820 vdd.n6227 vss 0.00219f
C8821 vdd.n6228 vss 0.00219f
C8822 vdd.n6229 vss 0.00748f
C8823 vdd.n6230 vss 3.87e-19
C8824 vdd.n6231 vss 0.008f
C8825 vdd.n6232 vss 0.00271f
C8826 vdd.n6233 vss 0.00335f
C8827 vdd.n6234 vss 0.00306f
C8828 vdd.n6235 vss 0.0115f
C8829 vdd.n6236 vss -0.173f
C8830 vdd.n6237 vss 0.0111f
C8831 vdd.n6238 vss 0.00284f
C8832 vdd.n6239 vss 0.00219f
C8833 vdd.n6240 vss 0.00219f
C8834 vdd.n6241 vss 0.00226f
C8835 vdd.n6242 vss 0.00219f
C8836 vdd.n6243 vss 0.00748f
C8837 vdd.n6244 vss 0.00271f
C8838 vdd.n6245 vss 2.66e-19
C8839 vdd.n6246 vss 0.00306f
C8840 vdd.n6247 vss 0.0182f
C8841 vdd.n6248 vss 0.00306f
C8842 vdd.n6249 vss 0.00284f
C8843 vdd.n6250 vss 0.00219f
C8844 vdd.n6251 vss 0.00219f
C8845 vdd.n6252 vss 0.00226f
C8846 vdd.n6253 vss 0.00219f
C8847 vdd.n6254 vss 0.0241f
C8848 vdd.n6255 vss 0.00271f
C8849 vdd.n6256 vss 2.66e-19
C8850 vdd.n6257 vss 0.0115f
C8851 vdd.n6258 vss 0.0197f
C8852 vdd.n6259 vss 0.00335f
C8853 vdd.n6260 vss 0.00359f
C8854 vdd.n6261 vss -0.148f
C8855 vdd.n6262 vss 0.00638f
C8856 vdd.n6263 vss 0.00284f
C8857 vdd.n6264 vss 0.00271f
C8858 vdd.n6265 vss 0.00219f
C8859 vdd.n6266 vss 0.0241f
C8860 vdd.n6267 vss 0.00219f
C8861 vdd.n6268 vss 0.00219f
C8862 vdd.n6269 vss 0.00226f
C8863 vdd.n6270 vss 0.00219f
C8864 vdd.n6271 vss 0.00748f
C8865 vdd.n6272 vss 0.00335f
C8866 vdd.n6273 vss 0.00359f
C8867 vdd.n6274 vss 0.0182f
C8868 vdd.n6275 vss 0.00638f
C8869 vdd.n6276 vss 0.00284f
C8870 vdd.n6277 vss 0.00271f
C8871 vdd.n6278 vss 0.00219f
C8872 vdd.n6279 vss 0.00219f
C8873 vdd.n6280 vss 0.008f
C8874 vdd.n6281 vss 0.00851f
C8875 vdd.n6282 vss 0.00219f
C8876 vdd.n6283 vss 0.00219f
C8877 vdd.n6284 vss 3.87e-19
C8878 vdd.n6285 vss 0.008f
C8879 vdd.n6286 vss 0.00271f
C8880 vdd.n6287 vss 0.00542f
C8881 vdd.n6288 vss 0.00271f
C8882 vdd.n6289 vss 0.00658f
C8883 vdd.n6290 vss -0.0615f
C8884 vdd.n6291 vss 0.0182f
C8885 vdd.n6292 vss 0.00399f
C8886 vdd.n6293 vss -0.0638f
C8887 vdd.n6294 vss 2.66e-19
C8888 vdd.n6295 vss 3.87e-19
C8889 vdd.n6296 vss 0.00477f
C8890 vdd.n6297 vss 0.00284f
C8891 vdd.n6298 vss 0.00219f
C8892 vdd.n6299 vss 0.0105f
C8893 vdd.n6300 vss 0.008f
C8894 vdd.n6301 vss 0.00271f
C8895 vdd.n6302 vss 0.00477f
C8896 vdd.n6303 vss 0.00284f
C8897 vdd.n6304 vss 3.87e-19
C8898 vdd.n6305 vss 2.66e-19
C8899 vdd.n6306 vss 0.00399f
C8900 vdd.n6307 vss 0.0186f
C8901 vdd.n6308 vss -0.0615f
C8902 vdd.n6309 vss 0.00335f
C8903 vdd.n6310 vss 0.00284f
C8904 vdd.n6311 vss 0.00748f
C8905 vdd.n6312 vss 0.00219f
C8906 vdd.n6313 vss 0.008f
C8907 vdd.n6314 vss 0.008f
C8908 vdd.n6315 vss 0.00219f
C8909 vdd.n6316 vss 0.00219f
C8910 vdd.n6317 vss 0.00219f
C8911 vdd.n6318 vss 0.00219f
C8912 vdd.n6319 vss 0.00284f
C8913 vdd.n6320 vss 0.0233f
C8914 vdd.n6321 vss 0.0115f
C8915 vdd.n6322 vss 2.66e-19
C8916 vdd.n6323 vss 0.00271f
C8917 vdd.n6324 vss 0.00284f
C8918 vdd.n6325 vss 0.00748f
C8919 vdd.n6326 vss 0.00219f
C8920 vdd.n6327 vss 0.00219f
C8921 vdd.n6328 vss 0.024f
C8922 vdd.n6329 vss 0.00271f
C8923 vdd.n6330 vss 0.0213f
C8924 vdd.n6331 vss 0.0234f
C8925 vdd.n6332 vss 0.0234f
C8926 vdd.n6333 vss 0.0213f
C8927 vdd.n6334 vss 0.00271f
C8928 vdd.n6335 vss 0.024f
C8929 vdd.n6336 vss 0.00219f
C8930 vdd.n6338 vss 0.00219f
C8931 vdd.n6339 vss 0.00219f
C8932 vdd.n6340 vss 0.00284f
C8933 vdd.n6341 vss 0.00335f
C8934 vdd.n6342 vss 0.00306f
C8935 vdd.n6343 vss 0.0115f
C8936 vdd.n6344 vss 2.66e-19
C8937 vdd.n6345 vss 0.00271f
C8938 vdd.n6346 vss 0.00748f
C8939 vdd.n6347 vss 0.00219f
C8940 vdd.n6348 vss 0.00851f
C8941 vdd.n6349 vss 0.00219f
C8942 vdd.n6350 vss 0.00219f
C8943 vdd.n6351 vss 0.00284f
C8944 vdd.n6352 vss 0.00335f
C8945 vdd.n6353 vss 0.00306f
C8946 vdd.n6354 vss -0.069f
C8947 vdd.n6355 vss 2.66e-19
C8948 vdd.n6356 vss 0.00271f
C8949 vdd.n6357 vss 0.00748f
C8950 vdd.n6358 vss 0.008f
C8951 vdd.n6359 vss 0.00226f
C8952 vdd.n6360 vss 0.00219f
C8953 vdd.n6361 vss 0.00219f
C8954 vdd.n6362 vss 0.00748f
C8955 vdd.n6363 vss 3.87e-19
C8956 vdd.n6364 vss 0.008f
C8957 vdd.n6365 vss 0.00271f
C8958 vdd.n6366 vss 0.00335f
C8959 vdd.n6367 vss 0.00306f
C8960 vdd.n6368 vss 0.0115f
C8961 vdd.n6369 vss -0.173f
C8962 vdd.n6370 vss 0.0111f
C8963 vdd.n6371 vss 0.00284f
C8964 vdd.n6372 vss 0.00219f
C8965 vdd.n6373 vss 0.00219f
C8966 vdd.n6375 vss 0.00219f
C8967 vdd.n6376 vss 0.00748f
C8968 vdd.n6377 vss 0.00271f
C8969 vdd.n6378 vss 2.66e-19
C8970 vdd.n6379 vss 0.00306f
C8971 vdd.n6380 vss 0.0182f
C8972 vdd.n6381 vss 0.00306f
C8973 vdd.n6382 vss 0.00284f
C8974 vdd.n6383 vss 0.00219f
C8975 vdd.n6384 vss 0.00219f
C8976 vdd.n6385 vss 0.0318f
C8977 vdd.n6386 vss 0.00271f
C8978 vdd.n6387 vss 2.66e-19
C8979 vdd.n6388 vss 0.131f
C8980 vdd.n6389 vss 0.00887f
C8981 vdd.n6390 vss 0.103f
C8982 vdd.n6391 vss 0.0163f
C8983 vdd.t31 vss 0.0077f
C8984 vdd.n6392 vss 0.111f
C8985 vdd.n6393 vss 0.0163f
C8986 vdd.n6394 vss 0.142f
C8987 vdd.n6395 vss 14f
C8988 vdd.n6396 vss 0.0115f
C8989 vdd.n6397 vss 0.0325f
C8990 vdd.n6398 vss 0.00359f
C8991 vdd.n6399 vss 0.0111f
C8992 vdd.n6400 vss -0.069f
C8993 vdd.n6401 vss -0.143f
C8994 vdd.n6402 vss 0.00651f
C8995 vdd.n6403 vss 0.00399f
C8996 vdd.n6404 vss 3.87e-19
C8997 vdd.n6405 vss 0.0344f
C8998 vdd.n6406 vss 0.0421f
C8999 vdd.n6407 vss 0.0165f
C9000 vdd.n6408 vss 0.00226f
C9001 vdd.n6409 vss 0.0105f
C9002 vdd.n6410 vss 0.008f
C9003 vdd.n6411 vss 0.008f
C9004 vdd.n6412 vss 0.00271f
C9005 vdd.n6413 vss 0.00542f
C9006 vdd.n6414 vss 0.00658f
C9007 vdd.n6415 vss 0.00335f
C9008 vdd.n6416 vss 0.00477f
C9009 vdd.n6417 vss 0.00385f
C9010 vdd.n6418 vss 0.00359f
C9011 vdd.n6419 vss 0.0111f
C9012 vdd.n6420 vss 0.0115f
C9013 vdd.n6421 vss 0.0182f
C9014 vdd.n6422 vss 0.0186f
C9015 vdd.n6423 vss 0.00651f
C9016 vdd.n6424 vss 0.00399f
C9017 vdd.n6425 vss 3.87e-19
C9018 vdd.n6426 vss 0.00284f
C9019 vdd.n6427 vss 2.58e-19
C9020 vdd.n6428 vss 0.00851f
C9021 vdd.n6430 vss 0.0105f
C9022 vdd.n6431 vss 0.008f
C9023 vdd.n6432 vss 0.008f
C9024 vdd.n6433 vss 0.00271f
C9025 vdd.n6434 vss 0.00542f
C9026 vdd.n6435 vss 0.00658f
C9027 vdd.n6436 vss 0.00477f
C9028 vdd.n6437 vss 0.00335f
C9029 vdd.n6438 vss 0.00271f
C9030 vdd.n6439 vss -0.0615f
C9031 vdd.n6440 vss 2.66e-19
C9032 vdd.n6441 vss 0.00399f
C9033 vdd.n6442 vss 0.00651f
C9034 vdd.n6443 vss 0.0186f
C9035 vdd.n6444 vss 0.0182f
C9036 vdd.n6445 vss 0.0111f
C9037 vdd.n6446 vss 0.00359f
C9038 vdd.n6447 vss 0.00385f
C9039 vdd.n6448 vss 0.00477f
C9040 vdd.n6449 vss 0.00542f
C9041 vdd.n6450 vss 0.00658f
C9042 vdd.n6451 vss 0.00284f
C9043 vdd.n6452 vss 0.00219f
C9044 vdd.n6453 vss 0.00284f
C9045 vdd.n6454 vss 2.58e-19
C9046 vdd.n6455 vss 0.00851f
C9047 vdd.n6456 vss 0.0105f
C9048 vdd.n6458 vss 0.00226f
C9049 vdd.n6459 vss 0.00219f
C9050 vdd.n6460 vss 2.58e-19
C9051 vdd.n6461 vss 0.00284f
C9052 vdd.n6462 vss 3.87e-19
C9053 vdd.n6463 vss 0.00399f
C9054 vdd.n6464 vss 0.00651f
C9055 vdd.n6465 vss -0.143f
C9056 vdd.n6466 vss 0.0182f
C9057 vdd.n6467 vss 0.0111f
C9058 vdd.n6468 vss 0.00359f
C9059 vdd.n6469 vss 0.00385f
C9060 vdd.n6470 vss 0.00477f
C9061 vdd.n6471 vss 0.00658f
C9062 vdd.n6472 vss 0.00542f
C9063 vdd.n6473 vss 0.00271f
C9064 vdd.n6474 vss 0.008f
C9065 vdd.n6475 vss 0.008f
C9066 vdd.n6476 vss 0.0105f
C9067 vdd.n6478 vss 0.00226f
C9068 vdd.n6479 vss 0.00851f
C9069 vdd.n6480 vss 2.58e-19
C9070 vdd.n6481 vss 0.00284f
C9071 vdd.n6482 vss 3.87e-19
C9072 vdd.n6483 vss 0.00399f
C9073 vdd.n6484 vss 0.00651f
C9074 vdd.n6485 vss 0.0186f
C9075 vdd.n6486 vss 0.0182f
C9076 vdd.n6487 vss 0.0111f
C9077 vdd.n6488 vss -0.0615f
C9078 vdd.n6489 vss -0.173f
C9079 vdd.n6490 vss 0.00477f
C9080 vdd.n6491 vss 0.00658f
C9081 vdd.n6492 vss 0.00542f
C9082 vdd.n6493 vss 0.00271f
C9083 vdd.n6494 vss 0.008f
C9084 vdd.n6495 vss 0.008f
C9085 vdd.n6496 vss 0.0105f
C9086 vdd.n6497 vss 0.00226f
C9087 vdd.n6498 vss 0.0191f
C9088 vdd.n6499 vss 4.31e-19
C9089 vdd.n6500 vss 0.00284f
C9090 vdd.n6501 vss 3.87e-19
C9091 vdd.n6502 vss 0.00399f
C9092 vdd.n6503 vss 0.0234f
C9093 vdd.n6504 vss 0.0657f
C9094 vdd.n6505 vss 0.0654f
C9095 vdd.n6506 vss 0.0115f
C9096 vdd.n6507 vss 0.0111f
C9097 vdd.n6508 vss 2.66e-19
C9098 vdd.n6509 vss 0.00385f
C9099 vdd.n6510 vss 0.00271f
C9100 vdd.n6511 vss 3.87e-19
C9101 vdd.n6512 vss 0.00284f
C9102 vdd.n6513 vss 4.31e-19
C9103 vdd.n6514 vss 0.0191f
C9104 vdd.n6515 vss 0.00226f
C9105 vdd.n6516 vss 0.0105f
C9106 vdd.n6519 vss 0.00226f
C9107 vdd.n6520 vss 0.00851f
C9108 vdd.n6521 vss 2.58e-19
C9109 vdd.n6522 vss 0.00219f
C9110 vdd.n6523 vss 0.008f
C9111 vdd.n6524 vss 0.00271f
C9112 vdd.n6525 vss 0.00542f
C9113 vdd.n6526 vss 0.00658f
C9114 vdd.n6527 vss 0.00477f
C9115 vdd.n6528 vss -0.173f
C9116 vdd.n6529 vss 0.00319f
C9117 vdd.n6530 vss 0.00385f
C9118 vdd.n6531 vss 0.00638f
C9119 vdd.n6532 vss 0.0182f
C9120 vdd.n6533 vss 0.0111f
C9121 vdd.n6534 vss -0.148f
C9122 vdd.n6535 vss 0.00385f
C9123 vdd.n6536 vss 0.00638f
C9124 vdd.n6537 vss 0.00319f
C9125 vdd.n6538 vss 0.0186f
C9126 vdd.n6539 vss 0.0115f
C9127 vdd.n6540 vss 0.00359f
C9128 vdd.n6541 vss 0.00271f
C9129 vdd.n6542 vss 0.00335f
C9130 vdd.n6543 vss 0.00748f
C9131 vdd.n6544 vss 0.00542f
C9132 vdd.n6545 vss 0.00658f
C9133 vdd.n6546 vss 0.00284f
C9134 vdd.n6547 vss 0.00219f
C9135 vdd.n6548 vss 0.00219f
C9136 vdd.n6549 vss 2.58e-19
C9137 vdd.n6550 vss 0.00851f
C9138 vdd.n6552 vss 0.00226f
C9139 vdd.n6554 vss 0.0105f
C9140 vdd.n6555 vss 0.008f
C9141 vdd.n6556 vss 0.008f
C9142 vdd.n6557 vss 0.00271f
C9143 vdd.n6558 vss 0.00284f
C9144 vdd.n6559 vss 0.00658f
C9145 vdd.n6560 vss 0.00542f
C9146 vdd.n6561 vss 0.00748f
C9147 vdd.n6562 vss 0.00335f
C9148 vdd.n6563 vss 0.00271f
C9149 vdd.n6564 vss 0.00359f
C9150 vdd.n6565 vss 0.0115f
C9151 vdd.n6566 vss 0.0186f
C9152 vdd.n6567 vss 0.00319f
C9153 vdd.n6568 vss 0.00638f
C9154 vdd.n6569 vss 0.00385f
C9155 vdd.n6570 vss 2.66e-19
C9156 vdd.n6571 vss 0.0111f
C9157 vdd.n6572 vss 0.0115f
C9158 vdd.n6573 vss 0.0186f
C9159 vdd.n6574 vss 0.00319f
C9160 vdd.n6575 vss -0.173f
C9161 vdd.n6576 vss 0.00477f
C9162 vdd.n6577 vss 0.00335f
C9163 vdd.n6578 vss 0.00748f
C9164 vdd.n6579 vss 0.00284f
C9165 vdd.n6580 vss 2.58e-19
C9166 vdd.n6581 vss 0.00219f
C9167 vdd.n6582 vss 0.00226f
C9168 vdd.n6584 vss 0.0105f
C9169 vdd.n6586 vss 0.00851f
C9170 vdd.n6587 vss 2.58e-19
C9171 vdd.n6588 vss 0.00284f
C9172 vdd.n6589 vss 3.87e-19
C9173 vdd.n6590 vss 0.00385f
C9174 vdd.n6591 vss 2.66e-19
C9175 vdd.n6592 vss 0.0111f
C9176 vdd.n6593 vss 0.0115f
C9177 vdd.n6594 vss 0.0186f
C9178 vdd.n6595 vss 0.00319f
C9179 vdd.n6596 vss 0.00399f
C9180 vdd.n6597 vss 0.00477f
C9181 vdd.n6598 vss 0.00658f
C9182 vdd.n6599 vss 0.00542f
C9183 vdd.n6600 vss 0.00271f
C9184 vdd.n6601 vss 0.008f
C9185 vdd.n6602 vss 0.008f
C9186 vdd.n6603 vss 0.0105f
C9187 vdd.n6605 vss 0.0142f
C9188 vdd.n6606 vss 0.0255f
C9189 vdd.n6607 vss 0.0255f
C9190 vdd.n6608 vss 0.0142f
C9191 vdd.n6609 vss 0.00226f
C9192 vdd.n6610 vss 0.00851f
C9193 vdd.n6611 vss 2.58e-19
C9194 vdd.n6612 vss 0.00284f
C9195 vdd.n6613 vss 3.87e-19
C9196 vdd.n6614 vss 0.00385f
C9197 vdd.n6615 vss 2.66e-19
C9198 vdd.n6616 vss -0.0638f
C9199 vdd.n6617 vss 0.0115f
C9200 vdd.n6618 vss 0.049f
C9201 vdd.n6619 vss 0.0198f
C9202 vdd.n6620 vss 0.00399f
C9203 vdd.n6621 vss 0.0205f
C9204 vdd.n6622 vss 0.00335f
C9205 vdd.n6623 vss 0.0205f
C9206 vdd.n6624 vss 0.00385f
C9207 vdd.n6625 vss 0.00359f
C9208 vdd.n6626 vss 0.0111f
C9209 vdd.n6627 vss -0.069f
C9210 vdd.n6628 vss -0.143f
C9211 vdd.n6629 vss 0.00651f
C9212 vdd.n6630 vss 0.00399f
C9213 vdd.n6631 vss 3.87e-19
C9214 vdd.n6632 vss 0.00284f
C9215 vdd.n6633 vss 2.58e-19
C9216 vdd.n6634 vss 0.00851f
C9217 vdd.n6636 vss 0.0105f
C9218 vdd.n6637 vss 0.008f
C9219 vdd.n6638 vss 0.008f
C9220 vdd.n6639 vss 0.00271f
C9221 vdd.n6640 vss 0.00542f
C9222 vdd.n6641 vss 0.00658f
C9223 vdd.n6642 vss 0.00335f
C9224 vdd.n6643 vss 0.00477f
C9225 vdd.n6644 vss 0.00385f
C9226 vdd.n6645 vss 0.00359f
C9227 vdd.n6646 vss 0.0111f
C9228 vdd.n6647 vss 0.0115f
C9229 vdd.n6648 vss 0.0182f
C9230 vdd.n6649 vss 0.0186f
C9231 vdd.n6650 vss 0.00651f
C9232 vdd.n6651 vss 0.00399f
C9233 vdd.n6652 vss 3.87e-19
C9234 vdd.n6653 vss 0.00284f
C9235 vdd.n6654 vss 2.58e-19
C9236 vdd.n6655 vss 0.00851f
C9237 vdd.n6657 vss 0.0105f
C9238 vdd.n6658 vss 0.008f
C9239 vdd.n6659 vss 0.008f
C9240 vdd.n6660 vss 0.00271f
C9241 vdd.n6661 vss 0.00542f
C9242 vdd.n6662 vss 0.00658f
C9243 vdd.n6663 vss 0.00477f
C9244 vdd.n6664 vss 0.00335f
C9245 vdd.n6665 vss 0.00271f
C9246 vdd.n6666 vss -0.0615f
C9247 vdd.n6667 vss 2.66e-19
C9248 vdd.n6668 vss 0.00399f
C9249 vdd.n6669 vss 0.00651f
C9250 vdd.n6670 vss 0.0186f
C9251 vdd.n6671 vss 0.0182f
C9252 vdd.n6672 vss 0.0111f
C9253 vdd.n6673 vss 0.00359f
C9254 vdd.n6674 vss 0.00385f
C9255 vdd.n6675 vss 0.00477f
C9256 vdd.n6676 vss 0.00542f
C9257 vdd.n6677 vss 0.00658f
C9258 vdd.n6678 vss 0.00284f
C9259 vdd.n6679 vss 0.00219f
C9260 vdd.n6680 vss 0.00284f
C9261 vdd.n6681 vss 2.58e-19
C9262 vdd.n6682 vss 0.00851f
C9263 vdd.n6683 vss 0.0105f
C9264 vdd.n6685 vss 0.00226f
C9265 vdd.n6686 vss 0.00219f
C9266 vdd.n6687 vss 2.58e-19
C9267 vdd.n6688 vss 0.00284f
C9268 vdd.n6689 vss 3.87e-19
C9269 vdd.n6690 vss 0.00399f
C9270 vdd.n6691 vss 0.00651f
C9271 vdd.n6692 vss -0.143f
C9272 vdd.n6693 vss 0.0182f
C9273 vdd.n6694 vss 0.0111f
C9274 vdd.n6695 vss 0.00359f
C9275 vdd.n6696 vss 0.00385f
C9276 vdd.n6697 vss 0.00477f
C9277 vdd.n6698 vss 0.00658f
C9278 vdd.n6699 vss 0.00542f
C9279 vdd.n6700 vss 0.00271f
C9280 vdd.n6701 vss 0.008f
C9281 vdd.n6702 vss 0.008f
C9282 vdd.n6703 vss 0.0105f
C9283 vdd.n6705 vss 0.00226f
C9284 vdd.n6706 vss 0.00851f
C9285 vdd.n6707 vss 2.58e-19
C9286 vdd.n6708 vss 0.00284f
C9287 vdd.n6709 vss 3.87e-19
C9288 vdd.n6710 vss 0.00399f
C9289 vdd.n6711 vss 0.00651f
C9290 vdd.n6712 vss 0.0186f
C9291 vdd.n6713 vss 0.0182f
C9292 vdd.n6714 vss 0.0111f
C9293 vdd.n6715 vss -0.0615f
C9294 vdd.n6716 vss -0.173f
C9295 vdd.n6717 vss 0.00477f
C9296 vdd.n6718 vss 0.00658f
C9297 vdd.n6719 vss 0.00542f
C9298 vdd.n6720 vss 0.00271f
C9299 vdd.n6721 vss 0.008f
C9300 vdd.n6722 vss 0.008f
C9301 vdd.n6723 vss 0.0105f
C9302 vdd.n6724 vss 0.00226f
C9303 vdd.n6725 vss 0.0191f
C9304 vdd.n6726 vss 4.31e-19
C9305 vdd.n6727 vss 0.00284f
C9306 vdd.n6728 vss 3.87e-19
C9307 vdd.n6729 vss 0.00399f
C9308 vdd.n6730 vss 0.0234f
C9309 vdd.n6731 vss 0.0657f
C9310 vdd.n6732 vss 0.0654f
C9311 vdd.n6733 vss 0.0115f
C9312 vdd.n6734 vss 0.0111f
C9313 vdd.n6735 vss 2.66e-19
C9314 vdd.n6736 vss 0.00385f
C9315 vdd.n6737 vss 0.00271f
C9316 vdd.n6738 vss 3.87e-19
C9317 vdd.n6739 vss 0.00284f
C9318 vdd.n6740 vss 4.31e-19
C9319 vdd.n6741 vss 0.0191f
C9320 vdd.n6742 vss 0.00226f
C9321 vdd.n6743 vss 0.0105f
C9322 vdd.n6746 vss 0.00226f
C9323 vdd.n6747 vss 0.00851f
C9324 vdd.n6748 vss 2.58e-19
C9325 vdd.n6749 vss 0.00219f
C9326 vdd.n6750 vss 0.008f
C9327 vdd.n6751 vss 0.00271f
C9328 vdd.n6752 vss 0.00542f
C9329 vdd.n6753 vss 0.00658f
C9330 vdd.n6754 vss 0.00477f
C9331 vdd.n6755 vss -0.173f
C9332 vdd.n6756 vss 0.00319f
C9333 vdd.n6757 vss 0.00385f
C9334 vdd.n6758 vss 0.00638f
C9335 vdd.n6759 vss 0.0182f
C9336 vdd.n6760 vss 0.0111f
C9337 vdd.n6761 vss -0.148f
C9338 vdd.n6762 vss 0.00385f
C9339 vdd.n6763 vss 0.00638f
C9340 vdd.n6764 vss 0.00319f
C9341 vdd.n6765 vss 0.0186f
C9342 vdd.n6766 vss 0.0115f
C9343 vdd.n6767 vss 0.00359f
C9344 vdd.n6768 vss 0.00271f
C9345 vdd.n6769 vss 0.00335f
C9346 vdd.n6770 vss 0.00748f
C9347 vdd.n6771 vss 0.00542f
C9348 vdd.n6772 vss 0.00658f
C9349 vdd.n6773 vss 0.00284f
C9350 vdd.n6774 vss 0.00219f
C9351 vdd.n6775 vss 0.00219f
C9352 vdd.n6776 vss 2.58e-19
C9353 vdd.n6777 vss 0.00851f
C9354 vdd.n6779 vss 0.00226f
C9355 vdd.n6781 vss 0.0105f
C9356 vdd.n6782 vss 0.008f
C9357 vdd.n6783 vss 0.008f
C9358 vdd.n6784 vss 0.00271f
C9359 vdd.n6785 vss 0.00284f
C9360 vdd.n6786 vss 0.00658f
C9361 vdd.n6787 vss 0.00542f
C9362 vdd.n6788 vss 0.00748f
C9363 vdd.n6789 vss 0.00335f
C9364 vdd.n6790 vss 0.00271f
C9365 vdd.n6791 vss 0.00359f
C9366 vdd.n6792 vss 0.0115f
C9367 vdd.n6793 vss 0.0186f
C9368 vdd.n6794 vss 0.00319f
C9369 vdd.n6795 vss 0.00638f
C9370 vdd.n6796 vss 0.00385f
C9371 vdd.n6797 vss 2.66e-19
C9372 vdd.n6798 vss 0.0111f
C9373 vdd.n6799 vss 0.0115f
C9374 vdd.n6800 vss 0.0186f
C9375 vdd.n6801 vss 0.00319f
C9376 vdd.n6802 vss -0.173f
C9377 vdd.n6803 vss 0.00477f
C9378 vdd.n6804 vss 0.00335f
C9379 vdd.n6805 vss 0.00748f
C9380 vdd.n6806 vss 0.00284f
C9381 vdd.n6807 vss 2.58e-19
C9382 vdd.n6808 vss 0.00219f
C9383 vdd.n6809 vss 0.00226f
C9384 vdd.n6811 vss 0.0105f
C9385 vdd.n6813 vss 0.00851f
C9386 vdd.n6814 vss 2.58e-19
C9387 vdd.n6815 vss 0.00284f
C9388 vdd.n6816 vss 3.87e-19
C9389 vdd.n6817 vss 0.00385f
C9390 vdd.n6818 vss 2.66e-19
C9391 vdd.n6819 vss 0.0111f
C9392 vdd.n6820 vss 0.0115f
C9393 vdd.n6821 vss 0.0186f
C9394 vdd.n6822 vss 0.00319f
C9395 vdd.n6823 vss 0.00399f
C9396 vdd.n6824 vss 0.00477f
C9397 vdd.n6825 vss 0.00658f
C9398 vdd.n6826 vss 0.00542f
C9399 vdd.n6827 vss 0.00271f
C9400 vdd.n6828 vss 0.008f
C9401 vdd.n6829 vss 0.008f
C9402 vdd.n6830 vss 0.0105f
C9403 vdd.n6832 vss 0.0142f
C9404 vdd.n6833 vss 0.0255f
C9405 vdd.n6834 vss 0.0255f
C9406 vdd.n6835 vss 0.0142f
C9407 vdd.n6836 vss 0.00226f
C9408 vdd.n6837 vss 0.00851f
C9409 vdd.n6838 vss 2.58e-19
C9410 vdd.n6839 vss 0.00284f
C9411 vdd.n6840 vss 3.87e-19
C9412 vdd.n6841 vss 0.00385f
C9413 vdd.n6842 vss 2.66e-19
C9414 vdd.n6843 vss -0.0638f
C9415 vdd.n6844 vss 0.0115f
C9416 vdd.n6845 vss 0.049f
C9417 vdd.n6846 vss 0.0198f
C9418 vdd.n6847 vss 0.00399f
C9419 vdd.n6848 vss 0.0205f
C9420 vdd.n6849 vss 0.00335f
C9421 vdd.n6850 vss 0.0205f
C9422 vdd.n6851 vss 0.00385f
C9423 vdd.n6852 vss 0.00359f
C9424 vdd.n6853 vss 0.0111f
C9425 vdd.n6854 vss -0.069f
C9426 vdd.n6855 vss -0.143f
C9427 vdd.n6856 vss 0.00651f
C9428 vdd.n6857 vss 0.00399f
C9429 vdd.n6858 vss 3.87e-19
C9430 vdd.n6859 vss 0.00284f
C9431 vdd.n6860 vss 2.58e-19
C9432 vdd.n6861 vss 0.00851f
C9433 vdd.n6863 vss 0.0105f
C9434 vdd.n6864 vss 0.008f
C9435 vdd.n6865 vss 0.008f
C9436 vdd.n6866 vss 0.00271f
C9437 vdd.n6867 vss 0.00542f
C9438 vdd.n6868 vss 0.00658f
C9439 vdd.n6869 vss 0.00335f
C9440 vdd.n6870 vss 0.00477f
C9441 vdd.n6871 vss 0.00385f
C9442 vdd.n6872 vss 0.00359f
C9443 vdd.n6873 vss 0.0111f
C9444 vdd.n6874 vss 0.0115f
C9445 vdd.n6875 vss 0.0182f
C9446 vdd.n6876 vss 0.0186f
C9447 vdd.n6877 vss 0.00651f
C9448 vdd.n6878 vss 0.00399f
C9449 vdd.n6879 vss 3.87e-19
C9450 vdd.n6880 vss 0.00284f
C9451 vdd.n6881 vss 2.58e-19
C9452 vdd.n6882 vss 0.00851f
C9453 vdd.n6884 vss 0.0105f
C9454 vdd.n6885 vss 0.008f
C9455 vdd.n6886 vss 0.008f
C9456 vdd.n6887 vss 0.00271f
C9457 vdd.n6888 vss 0.00542f
C9458 vdd.n6889 vss 0.00658f
C9459 vdd.n6890 vss 0.00477f
C9460 vdd.n6891 vss 0.00335f
C9461 vdd.n6892 vss 0.00271f
C9462 vdd.n6893 vss -0.0615f
C9463 vdd.n6894 vss 2.66e-19
C9464 vdd.n6895 vss 0.00399f
C9465 vdd.n6896 vss 0.00651f
C9466 vdd.n6897 vss 0.0186f
C9467 vdd.n6898 vss 0.0182f
C9468 vdd.n6899 vss 0.0111f
C9469 vdd.n6900 vss 0.00359f
C9470 vdd.n6901 vss 0.00385f
C9471 vdd.n6902 vss 0.00477f
C9472 vdd.n6903 vss 0.00542f
C9473 vdd.n6904 vss 0.00658f
C9474 vdd.n6905 vss 0.00284f
C9475 vdd.n6906 vss 0.00219f
C9476 vdd.n6907 vss 0.00284f
C9477 vdd.n6908 vss 2.58e-19
C9478 vdd.n6909 vss 0.00851f
C9479 vdd.n6910 vss 0.0105f
C9480 vdd.n6912 vss 0.00226f
C9481 vdd.n6913 vss 0.00219f
C9482 vdd.n6914 vss 2.58e-19
C9483 vdd.n6915 vss 0.00284f
C9484 vdd.n6916 vss 3.87e-19
C9485 vdd.n6917 vss 0.00399f
C9486 vdd.n6918 vss 0.00651f
C9487 vdd.n6919 vss -0.143f
C9488 vdd.n6920 vss 0.0182f
C9489 vdd.n6921 vss 0.0111f
C9490 vdd.n6922 vss 0.00359f
C9491 vdd.n6923 vss 0.00385f
C9492 vdd.n6924 vss 0.00477f
C9493 vdd.n6925 vss 0.00658f
C9494 vdd.n6926 vss 0.00542f
C9495 vdd.n6927 vss 0.00271f
C9496 vdd.n6928 vss 0.008f
C9497 vdd.n6929 vss 0.008f
C9498 vdd.n6930 vss 0.0105f
C9499 vdd.n6932 vss 0.00226f
C9500 vdd.n6933 vss 0.00851f
C9501 vdd.n6934 vss 2.58e-19
C9502 vdd.n6935 vss 0.00284f
C9503 vdd.n6936 vss 3.87e-19
C9504 vdd.n6937 vss 0.00399f
C9505 vdd.n6938 vss 0.00651f
C9506 vdd.n6939 vss 0.0186f
C9507 vdd.n6940 vss 0.0182f
C9508 vdd.n6941 vss 0.0111f
C9509 vdd.n6942 vss -0.0615f
C9510 vdd.n6943 vss -0.173f
C9511 vdd.n6944 vss 0.00477f
C9512 vdd.n6945 vss 0.00658f
C9513 vdd.n6946 vss 0.00542f
C9514 vdd.n6947 vss 0.00271f
C9515 vdd.n6948 vss 0.008f
C9516 vdd.n6949 vss 0.008f
C9517 vdd.n6950 vss 0.0105f
C9518 vdd.n6951 vss 0.00226f
C9519 vdd.n6952 vss 0.0191f
C9520 vdd.n6953 vss 4.31e-19
C9521 vdd.n6954 vss 0.00284f
C9522 vdd.n6955 vss 3.87e-19
C9523 vdd.n6956 vss 0.00399f
C9524 vdd.n6957 vss 0.0234f
C9525 vdd.n6958 vss 0.0657f
C9526 vdd.n6959 vss 0.0654f
C9527 vdd.n6960 vss 0.0115f
C9528 vdd.n6961 vss 0.0111f
C9529 vdd.n6962 vss 2.66e-19
C9530 vdd.n6963 vss 0.00385f
C9531 vdd.n6964 vss 0.00271f
C9532 vdd.n6965 vss 3.87e-19
C9533 vdd.n6966 vss 0.00284f
C9534 vdd.n6967 vss 4.31e-19
C9535 vdd.n6968 vss 0.0191f
C9536 vdd.n6969 vss 0.00226f
C9537 vdd.n6970 vss 0.0105f
C9538 vdd.n6973 vss 0.00226f
C9539 vdd.n6974 vss 0.00851f
C9540 vdd.n6975 vss 2.58e-19
C9541 vdd.n6976 vss 0.00219f
C9542 vdd.n6977 vss 0.008f
C9543 vdd.n6978 vss 0.00271f
C9544 vdd.n6979 vss 0.00542f
C9545 vdd.n6980 vss 0.00658f
C9546 vdd.n6981 vss 0.00477f
C9547 vdd.n6982 vss -0.173f
C9548 vdd.n6983 vss 0.00319f
C9549 vdd.n6984 vss 0.00385f
C9550 vdd.n6985 vss 0.00638f
C9551 vdd.n6986 vss 0.0182f
C9552 vdd.n6987 vss 0.0111f
C9553 vdd.n6988 vss -0.148f
C9554 vdd.n6989 vss 0.00385f
C9555 vdd.n6990 vss 0.00638f
C9556 vdd.n6991 vss 0.00319f
C9557 vdd.n6992 vss 0.0186f
C9558 vdd.n6993 vss 0.0115f
C9559 vdd.n6994 vss 0.00359f
C9560 vdd.n6995 vss 0.00271f
C9561 vdd.n6996 vss 0.00335f
C9562 vdd.n6997 vss 0.00748f
C9563 vdd.n6998 vss 0.00542f
C9564 vdd.n6999 vss 0.00658f
C9565 vdd.n7000 vss 0.00284f
C9566 vdd.n7001 vss 0.00219f
C9567 vdd.n7002 vss 0.00219f
C9568 vdd.n7003 vss 2.58e-19
C9569 vdd.n7004 vss 0.00851f
C9570 vdd.n7006 vss 0.00226f
C9571 vdd.n7008 vss 0.0105f
C9572 vdd.n7009 vss 0.008f
C9573 vdd.n7010 vss 0.008f
C9574 vdd.n7011 vss 0.00271f
C9575 vdd.n7012 vss 0.00284f
C9576 vdd.n7013 vss 0.00658f
C9577 vdd.n7014 vss 0.00542f
C9578 vdd.n7015 vss 0.00748f
C9579 vdd.n7016 vss 0.00335f
C9580 vdd.n7017 vss 0.00271f
C9581 vdd.n7018 vss 0.00359f
C9582 vdd.n7019 vss 0.0115f
C9583 vdd.n7020 vss 0.0186f
C9584 vdd.n7021 vss 0.00319f
C9585 vdd.n7022 vss 0.00638f
C9586 vdd.n7023 vss 0.00385f
C9587 vdd.n7024 vss 2.66e-19
C9588 vdd.n7025 vss 0.0111f
C9589 vdd.n7026 vss 0.0115f
C9590 vdd.n7027 vss 0.0186f
C9591 vdd.n7028 vss 0.00319f
C9592 vdd.n7029 vss -0.173f
C9593 vdd.n7030 vss 0.00477f
C9594 vdd.n7031 vss 0.00335f
C9595 vdd.n7032 vss 0.00748f
C9596 vdd.n7033 vss 0.00284f
C9597 vdd.n7034 vss 2.58e-19
C9598 vdd.n7035 vss 0.00219f
C9599 vdd.n7036 vss 0.00226f
C9600 vdd.n7038 vss 0.0105f
C9601 vdd.n7040 vss 0.00851f
C9602 vdd.n7041 vss 2.58e-19
C9603 vdd.n7042 vss 0.00284f
C9604 vdd.n7043 vss 3.87e-19
C9605 vdd.n7044 vss 0.00385f
C9606 vdd.n7045 vss 2.66e-19
C9607 vdd.n7046 vss 0.0111f
C9608 vdd.n7047 vss 0.0115f
C9609 vdd.n7048 vss 0.0186f
C9610 vdd.n7049 vss 0.00319f
C9611 vdd.n7050 vss 0.00399f
C9612 vdd.n7051 vss 0.00477f
C9613 vdd.n7052 vss 0.00658f
C9614 vdd.n7053 vss 0.00542f
C9615 vdd.n7054 vss 0.00271f
C9616 vdd.n7055 vss 0.008f
C9617 vdd.n7056 vss 0.008f
C9618 vdd.n7057 vss 0.0105f
C9619 vdd.n7059 vss 0.0142f
C9620 vdd.n7060 vss 0.0255f
C9621 vdd.n7061 vss 0.0255f
C9622 vdd.n7062 vss 0.0142f
C9623 vdd.n7063 vss 0.00226f
C9624 vdd.n7064 vss 0.00851f
C9625 vdd.n7065 vss 2.58e-19
C9626 vdd.n7066 vss 0.00284f
C9627 vdd.n7067 vss 3.87e-19
C9628 vdd.n7068 vss 0.00385f
C9629 vdd.n7069 vss 2.66e-19
C9630 vdd.n7070 vss -0.0638f
C9631 vdd.n7071 vss 0.0115f
C9632 vdd.n7072 vss 0.049f
C9633 vdd.n7073 vss 0.0198f
C9634 vdd.n7074 vss 0.00399f
C9635 vdd.n7075 vss 0.0205f
C9636 vdd.n7076 vss 0.00335f
C9637 vdd.n7077 vss 0.0205f
C9638 vdd.n7078 vss 0.00385f
C9639 vdd.n7079 vss 0.00359f
C9640 vdd.n7080 vss 0.0111f
C9641 vdd.n7081 vss -0.069f
C9642 vdd.n7082 vss -0.143f
C9643 vdd.n7083 vss 0.00651f
C9644 vdd.n7084 vss 0.00399f
C9645 vdd.n7085 vss 3.87e-19
C9646 vdd.n7086 vss 0.00284f
C9647 vdd.n7087 vss 2.58e-19
C9648 vdd.n7088 vss 0.00851f
C9649 vdd.n7090 vss 0.0105f
C9650 vdd.n7091 vss 0.008f
C9651 vdd.n7092 vss 0.008f
C9652 vdd.n7093 vss 0.00271f
C9653 vdd.n7094 vss 0.00542f
C9654 vdd.n7095 vss 0.00658f
C9655 vdd.n7096 vss 0.00335f
C9656 vdd.n7097 vss 0.00477f
C9657 vdd.n7098 vss 0.00385f
C9658 vdd.n7099 vss 0.00359f
C9659 vdd.n7100 vss 0.0111f
C9660 vdd.n7101 vss 0.0115f
C9661 vdd.n7102 vss 0.0182f
C9662 vdd.n7103 vss 0.0186f
C9663 vdd.n7104 vss 0.00651f
C9664 vdd.n7105 vss 0.00399f
C9665 vdd.n7106 vss 3.87e-19
C9666 vdd.n7107 vss 0.00284f
C9667 vdd.n7108 vss 2.58e-19
C9668 vdd.n7109 vss 0.00851f
C9669 vdd.n7111 vss 0.0105f
C9670 vdd.n7112 vss 0.008f
C9671 vdd.n7113 vss 0.008f
C9672 vdd.n7114 vss 0.00271f
C9673 vdd.n7115 vss 0.00542f
C9674 vdd.n7116 vss 0.00658f
C9675 vdd.n7117 vss 0.00477f
C9676 vdd.n7118 vss 0.00335f
C9677 vdd.n7119 vss 0.00271f
C9678 vdd.n7120 vss -0.0615f
C9679 vdd.n7121 vss 2.66e-19
C9680 vdd.n7122 vss 0.00399f
C9681 vdd.n7123 vss 0.00651f
C9682 vdd.n7124 vss 0.0186f
C9683 vdd.n7125 vss 0.0182f
C9684 vdd.n7126 vss 0.0111f
C9685 vdd.n7127 vss 0.00359f
C9686 vdd.n7128 vss 0.00385f
C9687 vdd.n7129 vss 0.00477f
C9688 vdd.n7130 vss 0.00542f
C9689 vdd.n7131 vss 0.00658f
C9690 vdd.n7132 vss 0.00284f
C9691 vdd.n7133 vss 0.00219f
C9692 vdd.n7134 vss 0.00284f
C9693 vdd.n7135 vss 2.58e-19
C9694 vdd.n7136 vss 0.00851f
C9695 vdd.n7137 vss 0.0105f
C9696 vdd.n7139 vss 0.00226f
C9697 vdd.n7140 vss 0.00219f
C9698 vdd.n7141 vss 2.58e-19
C9699 vdd.n7142 vss 0.00284f
C9700 vdd.n7143 vss 3.87e-19
C9701 vdd.n7144 vss 0.00399f
C9702 vdd.n7145 vss 0.00651f
C9703 vdd.n7146 vss -0.143f
C9704 vdd.n7147 vss 0.0182f
C9705 vdd.n7148 vss 0.0111f
C9706 vdd.n7149 vss 0.00359f
C9707 vdd.n7150 vss 0.00385f
C9708 vdd.n7151 vss 0.00477f
C9709 vdd.n7152 vss 0.00658f
C9710 vdd.n7153 vss 0.00542f
C9711 vdd.n7154 vss 0.00271f
C9712 vdd.n7155 vss 0.008f
C9713 vdd.n7156 vss 0.008f
C9714 vdd.n7157 vss 0.0105f
C9715 vdd.n7159 vss 0.00226f
C9716 vdd.n7160 vss 0.00851f
C9717 vdd.n7161 vss 2.58e-19
C9718 vdd.n7162 vss 0.00284f
C9719 vdd.n7163 vss 3.87e-19
C9720 vdd.n7164 vss 0.00399f
C9721 vdd.n7165 vss 0.00651f
C9722 vdd.n7166 vss 0.0186f
C9723 vdd.n7167 vss 0.0182f
C9724 vdd.n7168 vss 0.0111f
C9725 vdd.n7169 vss -0.0615f
C9726 vdd.n7170 vss -0.173f
C9727 vdd.n7171 vss 0.00477f
C9728 vdd.n7172 vss 0.00658f
C9729 vdd.n7173 vss 0.00542f
C9730 vdd.n7174 vss 0.00271f
C9731 vdd.n7175 vss 0.008f
C9732 vdd.n7176 vss 0.008f
C9733 vdd.n7177 vss 0.0105f
C9734 vdd.n7178 vss 0.00226f
C9735 vdd.n7179 vss 0.0191f
C9736 vdd.n7180 vss 4.31e-19
C9737 vdd.n7181 vss 0.00284f
C9738 vdd.n7182 vss 3.87e-19
C9739 vdd.n7183 vss 0.00399f
C9740 vdd.n7184 vss 0.0234f
C9741 vdd.n7185 vss 0.0657f
C9742 vdd.n7186 vss 0.0654f
C9743 vdd.n7187 vss 0.0115f
C9744 vdd.n7188 vss 0.0111f
C9745 vdd.n7189 vss 2.66e-19
C9746 vdd.n7190 vss 0.00385f
C9747 vdd.n7191 vss 0.00271f
C9748 vdd.n7192 vss 3.87e-19
C9749 vdd.n7193 vss 0.00284f
C9750 vdd.n7194 vss 4.31e-19
C9751 vdd.n7195 vss 0.0191f
C9752 vdd.n7196 vss 0.00226f
C9753 vdd.n7197 vss 0.0105f
C9754 vdd.n7200 vss 0.00226f
C9755 vdd.n7201 vss 0.00851f
C9756 vdd.n7202 vss 2.58e-19
C9757 vdd.n7203 vss 0.00219f
C9758 vdd.n7204 vss 0.008f
C9759 vdd.n7205 vss 0.00271f
C9760 vdd.n7206 vss 0.00542f
C9761 vdd.n7207 vss 0.00658f
C9762 vdd.n7208 vss 0.00477f
C9763 vdd.n7209 vss -0.173f
C9764 vdd.n7210 vss 0.00319f
C9765 vdd.n7211 vss 0.00385f
C9766 vdd.n7212 vss 0.00638f
C9767 vdd.n7213 vss 0.0182f
C9768 vdd.n7214 vss 0.0111f
C9769 vdd.n7215 vss -0.148f
C9770 vdd.n7216 vss 0.00385f
C9771 vdd.n7217 vss 0.00638f
C9772 vdd.n7218 vss 0.00319f
C9773 vdd.n7219 vss 0.0186f
C9774 vdd.n7220 vss 0.0115f
C9775 vdd.n7221 vss 0.00359f
C9776 vdd.n7222 vss 0.00271f
C9777 vdd.n7223 vss 0.00335f
C9778 vdd.n7224 vss 0.00748f
C9779 vdd.n7225 vss 0.00542f
C9780 vdd.n7226 vss 0.00658f
C9781 vdd.n7227 vss 0.00284f
C9782 vdd.n7228 vss 0.00219f
C9783 vdd.n7229 vss 0.00219f
C9784 vdd.n7230 vss 2.58e-19
C9785 vdd.n7231 vss 0.00851f
C9786 vdd.n7233 vss 0.00226f
C9787 vdd.n7235 vss 0.0105f
C9788 vdd.n7236 vss 0.008f
C9789 vdd.n7237 vss 0.008f
C9790 vdd.n7238 vss 0.00271f
C9791 vdd.n7239 vss 0.00284f
C9792 vdd.n7240 vss 0.00658f
C9793 vdd.n7241 vss 0.00542f
C9794 vdd.n7242 vss 0.00748f
C9795 vdd.n7243 vss 0.00335f
C9796 vdd.n7244 vss 0.00271f
C9797 vdd.n7245 vss 0.00359f
C9798 vdd.n7246 vss 0.0115f
C9799 vdd.n7247 vss 0.0186f
C9800 vdd.n7248 vss 0.00319f
C9801 vdd.n7249 vss 0.00638f
C9802 vdd.n7250 vss 0.00385f
C9803 vdd.n7251 vss 2.66e-19
C9804 vdd.n7252 vss 0.0111f
C9805 vdd.n7253 vss 0.0115f
C9806 vdd.n7254 vss 0.0186f
C9807 vdd.n7255 vss 0.00319f
C9808 vdd.n7256 vss -0.173f
C9809 vdd.n7257 vss 0.00477f
C9810 vdd.n7258 vss 0.00335f
C9811 vdd.n7259 vss 0.00748f
C9812 vdd.n7260 vss 0.00284f
C9813 vdd.n7261 vss 2.58e-19
C9814 vdd.n7262 vss 0.00219f
C9815 vdd.n7263 vss 0.00226f
C9816 vdd.n7265 vss 0.0105f
C9817 vdd.n7267 vss 0.00851f
C9818 vdd.n7268 vss 2.58e-19
C9819 vdd.n7269 vss 0.00284f
C9820 vdd.n7270 vss 3.87e-19
C9821 vdd.n7271 vss 0.00385f
C9822 vdd.n7272 vss 2.66e-19
C9823 vdd.n7273 vss 0.0111f
C9824 vdd.n7274 vss 0.0115f
C9825 vdd.n7275 vss 0.00385f
C9826 vdd.n7276 vss 2.66e-19
C9827 vdd.n7277 vss -0.0638f
C9828 vdd.n7278 vss -0.148f
C9829 vdd.n7279 vss 0.0186f
C9830 vdd.n7280 vss 0.00319f
C9831 vdd.n7281 vss 0.00399f
C9832 vdd.n7282 vss 0.00477f
C9833 vdd.n7283 vss 0.00284f
C9834 vdd.n7284 vss 0.00658f
C9835 vdd.n7285 vss 0.00542f
C9836 vdd.n7286 vss 0.00271f
C9837 vdd.n7287 vss 0.008f
C9838 vdd.n7288 vss 0.008f
C9839 vdd.n7289 vss 0.0105f
C9840 vdd.n7290 vss 0.0165f
C9841 vdd.n7291 vss 0.0421f
C9842 vdd.n7292 vss 0.0344f
C9843 vdd.n7293 vss 0.0318f
C9844 vdd.n7294 vss 0.0325f
C9845 vdd.n7295 vss 0.0491f
C9846 vdd.n7296 vss 0.506f
C9847 vdd.n7297 vss 0.528f
C9848 vdd.n7298 vss 0.0515f
C9849 vdd.n7299 vss 0.00226f
C9850 vdd.n7300 vss 0.0193f
C9851 vdd.n7301 vss 0.0256f
C9852 vdd.n7302 vss 0.0471f
C9853 vdd.n7303 vss 0.00271f
C9854 vdd.n7304 vss 0.0354f
C9855 vdd.n7305 vss 0.0358f
C9856 vdd.n7306 vss 2.66e-19
C9857 vdd.n7307 vss 0.0113f
C9858 vdd.n7308 vss 0.0117f
C9859 vdd.n7309 vss 0.0189f
C9860 vdd.n7310 vss 0.00319f
C9861 vdd.n7311 vss -0.173f
C9862 vdd.n7312 vss 0.00477f
C9863 vdd.n7313 vss 0.00658f
C9864 vdd.n7314 vss 0.00542f
C9865 vdd.n7315 vss 0.00271f
C9866 vdd.n7316 vss 0.008f
C9867 vdd.n7317 vss 0.008f
C9868 vdd.n7318 vss 0.0105f
C9869 vdd.n7320 vss 0.00851f
C9870 vdd.n7321 vss 2.58e-19
C9871 vdd.n7322 vss 0.00284f
C9872 vdd.n7323 vss 3.87e-19
C9873 vdd.n7324 vss 0.00385f
C9874 vdd.n7325 vss 2.66e-19
C9875 vdd.n7326 vss 0.0113f
C9876 vdd.n7327 vss 0.0117f
C9877 vdd.n7328 vss 0.0189f
C9878 vdd.n7329 vss 0.00319f
C9879 vdd.n7330 vss 0.00399f
C9880 vdd.n7331 vss 0.00477f
C9881 vdd.n7332 vss 0.00658f
C9882 vdd.n7333 vss 0.00542f
C9883 vdd.n7334 vss 0.00271f
C9884 vdd.n7335 vss 0.008f
C9885 vdd.n7336 vss 0.008f
C9886 vdd.n7337 vss 0.0105f
C9887 vdd.n7339 vss 0.00851f
C9888 vdd.n7340 vss 2.58e-19
C9889 vdd.n7341 vss 0.00284f
C9890 vdd.n7342 vss 3.87e-19
C9891 vdd.n7343 vss 0.00385f
C9892 vdd.n7344 vss 2.66e-19
C9893 vdd.n7345 vss -0.0637f
C9894 vdd.n7346 vss 0.0117f
C9895 vdd.n7347 vss 0.0189f
C9896 vdd.n7348 vss 0.00319f
C9897 vdd.n7349 vss 0.00399f
C9898 vdd.n7350 vss 0.00477f
C9899 vdd.n7351 vss 0.00658f
C9900 vdd.n7352 vss 0.00542f
C9901 vdd.n7353 vss 0.00271f
C9902 vdd.n7354 vss 0.008f
C9903 vdd.n7355 vss 0.008f
C9904 vdd.n7356 vss 0.0105f
C9905 vdd.n7358 vss 0.00851f
C9906 vdd.n7359 vss 2.58e-19
C9907 vdd.n7360 vss 0.00284f
C9908 vdd.n7361 vss 3.87e-19
C9909 vdd.n7362 vss 0.00385f
C9910 vdd.n7363 vss 2.66e-19
C9911 vdd.n7364 vss 0.0113f
C9912 vdd.n7365 vss 0.0117f
C9913 vdd.n7366 vss 0.0189f
C9914 vdd.n7367 vss 0.00319f
C9915 vdd.n7368 vss -0.173f
C9916 vdd.n7369 vss 0.00477f
C9917 vdd.n7370 vss 0.00658f
C9918 vdd.n7371 vss 0.00542f
C9919 vdd.n7372 vss 0.00271f
C9920 vdd.n7373 vss 0.008f
C9921 vdd.n7374 vss 0.008f
C9922 vdd.n7375 vss 0.0105f
C9923 vdd.n7377 vss 0.00851f
C9924 vdd.n7378 vss 2.58e-19
C9925 vdd.n7379 vss 0.00284f
C9926 vdd.n7380 vss 3.87e-19
C9927 vdd.n7381 vss 0.00385f
C9928 vdd.n7382 vss 2.66e-19
C9929 vdd.n7383 vss 0.0113f
C9930 vdd.n7384 vss 0.0117f
C9931 vdd.n7385 vss 0.0117f
C9932 vdd.n7386 vss 2.66e-19
C9933 vdd.n7387 vss -0.0637f
C9934 vdd.n7388 vss -0.148f
C9935 vdd.n7389 vss 0.0189f
C9936 vdd.n7390 vss 0.00319f
C9937 vdd.n7391 vss 0.00399f
C9938 vdd.n7392 vss 0.00477f
C9939 vdd.n7393 vss 0.00658f
C9940 vdd.n7394 vss 0.00542f
C9941 vdd.n7395 vss 0.00271f
C9942 vdd.n7396 vss 0.008f
C9943 vdd.n7397 vss 0.008f
C9944 vdd.n7398 vss 0.0105f
C9945 vdd.n7400 vss 0.00851f
C9946 vdd.n7401 vss 2.58e-19
C9947 vdd.n7402 vss 0.00284f
C9948 vdd.n7403 vss 3.87e-19
C9949 vdd.n7404 vss 0.00271f
C9950 vdd.n7405 vss 0.00335f
C9951 vdd.n7406 vss 0.00637f
C9952 vdd.n7407 vss 0.00399f
C9953 vdd.n7408 vss 0.00626f
C9954 vdd.n7409 vss 0.00504f
C9955 vdd.n7410 vss 0.00667f
C9956 vdd.n7411 vss 0.0249f
C9957 vdd.n7412 vss 0.0226f
C9958 vdd.n7413 vss 0.139f
C9959 vdd.n7414 vss 0.29f
C9960 vdd.n7415 vss 0.164f
C9961 vdd.n7416 vss 0.233f
C9962 vdd.n7417 vss 0.314f
C9963 vdd.n7418 vss 0.0136f
C9964 vdd.n7419 vss 8.67e-19
C9965 vdd.n7420 vss 0.0142f
C9966 vdd.n7421 vss 0.0295f
C9967 vdd.n7422 vss 0.0473f
C9968 vdd.n7423 vss 0.0517f
C9969 vdd.n7424 vss 0.251f
C9970 vdd.t80 vss 1.84f
C9971 vdd.n7425 vss 1.65f
C9972 vdd.n7426 vss 0.0664f
C9973 vdd.n7427 vss 0.00668f
C9974 vdd.n7428 vss 0.00518f
C9975 vdd.n7429 vss 0.00887f
C9976 vdd.n7430 vss 0.0131f
C9977 vdd.n7431 vss 0.00887f
C9978 vdd.n7432 vss 0.00518f
C9979 vdd.n7433 vss 0.0163f
C9980 vdd.n7434 vss 0.00673f
C9981 vdd.t81 vss 1.9f
C9982 vdd.t1 vss 0.35f
C9983 vdd.t102 vss 0.732f
C9984 vdd.n7435 vss 0.0127f
C9985 vdd.t32 vss 1.8f
C9986 vdd.t30 vss 5.45f
C9987 vdd.t79 vss 4.45f
C9988 vdd.n7436 vss 1.69f
C9989 vdd.n7437 vss 0.0664f
C9990 vdd.n7438 vss 0.00668f
C9991 vdd.n7439 vss 0.0163f
C9992 vdd.n7440 vss 0.0131f
C9993 vdd.n7441 vss 0.0547f
C9994 vdd.n7442 vss 0.0163f
C9995 vdd.n7443 vss 0.00668f
C9996 vdd.n7444 vss 0.0664f
C9997 vdd.n7445 vss 0.00673f
C9998 vdd.n7446 vss 0.0163f
C9999 vdd.n7447 vss 0.243f
C10000 vdd.n7448 vss 0.363f
C10001 vdd.n7449 vss 1.68f
C10002 vdd.n7450 vss 0.253f
C10003 vdd.n7451 vss 0.218f
C10004 vdd.n7452 vss 0.0427f
C10005 vdd.n7453 vss 0.00668f
C10006 vdd.n7454 vss 0.0163f
C10007 vdd.n7455 vss 0.00887f
C10008 vdd.n7456 vss 0.0427f
C10009 vdd.n7457 vss 0.00887f
C10010 vdd.n7458 vss 0.00518f
C10011 vdd.n7459 vss 0.00668f
C10012 vdd.n7460 vss 0.0664f
C10013 vdd.n7461 vss 0.162f
C10014 vdd.n7462 vss 0.167f
C10015 vdd.n7463 vss 0.0331f
C10016 vdd.n7464 vss 0.107f
C10017 vdd.n7465 vss 0.0114f
C10018 vdd.n7466 vss 0.00111f
C10019 vdd.n7467 vss 0.0015f
C10020 vdd.n7468 vss 0.00394f
C10021 vdd.n7469 vss 0.00713f
C10022 vdd.n7470 vss 0.00549f
C10023 vdd.n7471 vss 0.00564f
C10024 vdd.n7472 vss 0.0139f
C10025 vdd.n7473 vss 0.0189f
C10026 vdd.n7474 vss 0.0334f
C10027 vdd.n7475 vss 0.013f
C10028 vdd.n7476 vss 0.0161f
C10029 vdd.n7477 vss 0.0173f
C10030 vdd.n7478 vss 0.0183f
C10031 vdd.n7479 vss 0.0454f
C10032 vdd.n7480 vss 0.00651f
C10033 vdd.n7481 vss 0.0165f
C10034 vdd.n7482 vss 0.206f
C10035 vdd.n7483 vss 1.57f
C10036 vdd.t65 vss 0.268f
C10037 vdd.n7484 vss 0.136f
C10038 vdd.n7485 vss 0.0256f
C10039 vdd.n7486 vss 0.00651f
C10040 vdd.n7487 vss 0.00319f
C10041 vdd.n7488 vss 0.00893f
C10042 vdd.n7489 vss 0.00869f
C10043 vdd.n7490 vss 0.0223f
C10044 vdd.n7491 vss 0.0141f
C10045 vdd.n7492 vss 0.0162f
C10046 vdd.n7493 vss 6.66e-19
C10047 vdd.n7494 vss 0.0102f
C10048 vdd.n7495 vss 0.0413f
C10049 vdd.n7496 vss 0.0175f
C10050 vdd.n7497 vss 0.0139f
C10051 vdd.n7498 vss 0.00564f
C10052 vdd.n7499 vss 0.00549f
C10053 vdd.n7500 vss 0.00376f
C10054 vdd.n7501 vss 0.00394f
C10055 vdd.n7502 vss 0.0015f
C10056 vdd.n7503 vss 0.00111f
C10057 vdd.n7504 vss 0.00882f
C10058 vdd.n7505 vss 0.00209f
C10059 vdd.n7506 vss 0.00133f
C10060 vdd.n7507 vss 0.032f
C10061 vdd.n7508 vss 0.162f
C10062 vdd.t42 vss 0.22f
C10063 vdd.n7509 vss 0.2f
C10064 vdd.n7510 vss 0.0165f
C10065 vdd.n7511 vss 0.00651f
C10066 vdd.n7512 vss 0.0454f
C10067 vdd.n7513 vss 0.0183f
C10068 vdd.n7514 vss 0.0173f
C10069 vdd.n7515 vss 0.0161f
C10070 vdd.n7516 vss 0.0126f
C10071 vdd.n7517 vss 0.0909f
C10072 vdd.n7518 vss 5.43f
C10073 vdd.n7519 vss 0.721f
C10074 vdd.n7520 vss 0.0298f
C10075 vdd.n7521 vss 0.0289f
C10076 vdd.n7522 vss 0.163f
C10077 vdd.n7523 vss 0.164f
C10078 vdd.n7524 vss 0.0298f
C10079 vdd.n7525 vss 0.0289f
C10080 vdd.n7526 vss 0.00433f
C10081 vdd.n7527 vss 0.00246f
C10082 vdd.n7528 vss 0.0163f
C10083 vdd.n7529 vss 0.00885f
C10084 vdd.n7530 vss 0.0173f
C10085 CAP_CTRL_CODE0[0].t0 vss 0.0571f
C10086 CAP_CTRL_CODE0[0].n0 vss 12.1f
.ends

