magic
tech sky130A
magscale 1 2
timestamp 1698575955
<< error_s >>
rect 666 2102 724 2108
rect 666 2068 678 2102
rect 666 2062 724 2068
rect 666 1908 724 1914
rect 666 1874 678 1908
rect 666 1868 724 1874
use hgu_cdac_unit  x2
timestamp 1698474146
transform 1 0 -317 0 1 -51
box 686 598 1358 1826
use sky130_fd_pr__nfet_01v8_L7T3GD  XM14
timestamp 1698474146
transform 1 0 695 0 1 1988
box -211 -252 211 252
<< end >>
