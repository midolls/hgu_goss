magic
tech sky130A
magscale 1 2
timestamp 1698913543
<< nwell >>
rect -38 1236 666 1250
rect -38 1058 668 1236
rect -38 861 666 1058
<< pwell >>
rect 42 621 228 803
rect 394 621 580 803
rect 42 617 63 621
rect 394 617 415 621
rect 29 583 63 617
rect 381 583 415 617
<< scnmos >>
rect 120 647 150 777
rect 472 647 502 777
<< scpmoshvt >>
rect 120 897 150 1097
rect 472 897 502 1097
<< ndiff >>
rect 68 765 120 777
rect 68 731 76 765
rect 110 731 120 765
rect 68 697 120 731
rect 68 663 76 697
rect 110 663 120 697
rect 68 647 120 663
rect 150 765 202 777
rect 150 731 160 765
rect 194 731 202 765
rect 150 697 202 731
rect 150 663 160 697
rect 194 663 202 697
rect 150 647 202 663
rect 420 765 472 777
rect 420 731 428 765
rect 462 731 472 765
rect 420 697 472 731
rect 420 663 428 697
rect 462 663 472 697
rect 420 647 472 663
rect 502 765 554 777
rect 502 731 512 765
rect 546 731 554 765
rect 502 697 554 731
rect 502 663 512 697
rect 546 663 554 697
rect 502 647 554 663
<< pdiff >>
rect 68 1085 120 1097
rect 68 1051 76 1085
rect 110 1051 120 1085
rect 68 1017 120 1051
rect 68 983 76 1017
rect 110 983 120 1017
rect 68 949 120 983
rect 68 915 76 949
rect 110 915 120 949
rect 68 897 120 915
rect 150 1085 202 1097
rect 150 1051 160 1085
rect 194 1051 202 1085
rect 150 1017 202 1051
rect 150 983 160 1017
rect 194 983 202 1017
rect 150 949 202 983
rect 150 915 160 949
rect 194 915 202 949
rect 150 897 202 915
rect 420 1085 472 1097
rect 420 1051 428 1085
rect 462 1051 472 1085
rect 420 1017 472 1051
rect 420 983 428 1017
rect 462 983 472 1017
rect 420 949 472 983
rect 420 915 428 949
rect 462 915 472 949
rect 420 897 472 915
rect 502 1085 554 1097
rect 502 1051 512 1085
rect 546 1051 554 1085
rect 502 1017 554 1051
rect 502 983 512 1017
rect 546 983 554 1017
rect 502 949 554 983
rect 502 915 512 949
rect 546 915 554 949
rect 502 897 554 915
<< ndiffc >>
rect 76 731 110 765
rect 76 663 110 697
rect 160 731 194 765
rect 160 663 194 697
rect 428 731 462 765
rect 428 663 462 697
rect 512 731 546 765
rect 512 663 546 697
<< pdiffc >>
rect 76 1051 110 1085
rect 76 983 110 1017
rect 76 915 110 949
rect 160 1051 194 1085
rect 160 983 194 1017
rect 160 915 194 949
rect 428 1051 462 1085
rect 428 983 462 1017
rect 428 915 462 949
rect 512 1051 546 1085
rect 512 983 546 1017
rect 512 915 546 949
<< psubdiff >>
rect 2 586 630 590
rect 2 552 156 586
rect 190 552 630 586
<< nsubdiff >>
rect 0 1188 628 1190
rect 0 1154 121 1188
rect 155 1154 628 1188
rect 0 1152 628 1154
<< psubdiffcont >>
rect 156 552 190 586
<< nsubdiffcont >>
rect 121 1154 155 1188
<< poly >>
rect 120 1097 150 1123
rect 472 1097 502 1123
rect 120 865 150 897
rect 472 865 502 897
rect 64 849 150 865
rect 64 815 80 849
rect 114 815 150 849
rect 64 799 150 815
rect 416 849 502 865
rect 416 815 432 849
rect 466 815 502 849
rect 416 799 502 815
rect 120 777 150 799
rect 472 777 502 799
rect 120 621 150 647
rect 472 621 502 647
<< polycont >>
rect 80 815 114 849
rect 432 815 466 849
<< locali >>
rect 104 1188 172 1190
rect 104 1161 121 1188
rect 155 1161 172 1188
rect 0 1127 29 1161
rect 63 1127 121 1161
rect 155 1127 213 1161
rect 247 1127 276 1161
rect 352 1127 381 1161
rect 415 1127 473 1161
rect 507 1127 565 1161
rect 599 1127 628 1161
rect 68 1085 110 1127
rect 68 1051 76 1085
rect 68 1017 110 1051
rect 68 983 76 1017
rect 68 949 110 983
rect 68 915 76 949
rect 68 899 110 915
rect 144 1085 210 1093
rect 144 1051 160 1085
rect 194 1051 210 1085
rect 144 1017 210 1051
rect 144 983 160 1017
rect 194 983 210 1017
rect 144 949 210 983
rect 144 915 160 949
rect 194 915 210 949
rect 144 897 210 915
rect 420 1085 462 1127
rect 420 1051 428 1085
rect 420 1017 462 1051
rect 420 983 428 1017
rect 420 949 462 983
rect 420 915 428 949
rect 420 899 462 915
rect 496 1085 562 1093
rect 496 1051 512 1085
rect 546 1051 562 1085
rect 496 1017 562 1051
rect 496 983 512 1017
rect 546 983 562 1017
rect 496 949 562 983
rect 496 915 512 949
rect 546 915 562 949
rect 496 897 562 915
rect 64 852 130 863
rect 64 818 74 852
rect 108 849 130 852
rect 64 815 80 818
rect 114 815 130 849
rect 164 854 210 897
rect 416 854 482 863
rect 164 849 482 854
rect 164 820 432 849
rect 64 765 110 781
rect 164 777 210 820
rect 416 815 432 820
rect 466 815 482 849
rect 516 858 562 897
rect 516 824 526 858
rect 560 824 562 858
rect 64 731 76 765
rect 64 697 110 731
rect 64 663 76 697
rect 64 617 110 663
rect 144 765 210 777
rect 144 731 160 765
rect 194 731 210 765
rect 144 697 210 731
rect 144 663 160 697
rect 194 663 210 697
rect 144 651 210 663
rect 416 765 462 781
rect 516 777 562 824
rect 416 731 428 765
rect 416 697 462 731
rect 416 663 428 697
rect 416 617 462 663
rect 496 765 562 777
rect 496 731 512 765
rect 546 731 562 765
rect 496 697 562 731
rect 496 663 512 697
rect 546 663 562 697
rect 496 651 562 663
rect 0 583 29 617
rect 63 583 121 617
rect 155 586 213 617
rect 155 583 156 586
rect 138 552 156 583
rect 190 583 213 586
rect 247 583 276 617
rect 352 583 381 617
rect 415 583 473 617
rect 507 583 565 617
rect 599 583 628 617
rect 190 552 206 583
<< viali >>
rect 29 1127 63 1161
rect 121 1154 155 1161
rect 121 1127 155 1154
rect 213 1127 247 1161
rect 381 1127 415 1161
rect 473 1127 507 1161
rect 565 1127 599 1161
rect 74 849 108 852
rect 74 818 80 849
rect 80 818 108 849
rect 526 824 560 858
rect 29 583 63 617
rect 121 583 155 617
rect 213 583 247 617
rect 381 583 415 617
rect 473 583 507 617
rect 565 583 599 617
<< metal1 >>
rect 0 1192 626 1206
rect 0 1161 628 1192
rect 0 1127 29 1161
rect 63 1127 121 1161
rect 155 1127 213 1161
rect 247 1127 381 1161
rect 415 1127 473 1161
rect 507 1127 565 1161
rect 599 1127 628 1161
rect 0 1108 628 1127
rect 0 1096 276 1108
rect 352 1096 628 1108
rect 514 858 684 866
rect -54 852 124 858
rect -54 818 74 852
rect 108 818 124 852
rect -54 810 124 818
rect 514 824 526 858
rect 560 824 684 858
rect 514 816 684 824
rect -54 808 106 810
rect 0 628 276 648
rect 352 628 628 648
rect 0 617 628 628
rect 0 583 29 617
rect 63 583 121 617
rect 155 583 213 617
rect 247 583 381 617
rect 415 583 473 617
rect 507 583 565 617
rect 599 583 628 617
rect 0 552 628 583
rect 0 530 626 552
<< labels >>
flabel metal1 0 1108 550 1206 0 FreeSans 320 0 0 0 VDD
port 0 nsew
flabel metal1 0 530 550 628 0 FreeSans 320 0 0 0 VSS
port 1 nsew
flabel metal1 -54 808 106 858 0 FreeSans 320 0 0 0 in
port 2 nsew
flabel metal1 524 816 684 866 0 FreeSans 320 0 0 0 out
port 4 nsew
flabel locali 516 889 550 923 0 FreeSans 340 0 0 0 x2.Y
flabel locali 516 821 550 855 0 FreeSans 340 0 0 0 x2.Y
flabel locali 424 821 458 855 0 FreeSans 340 0 0 0 x2.A
flabel metal1 381 583 415 617 0 FreeSans 200 0 0 0 x2.VGND
flabel metal1 381 1127 415 1161 0 FreeSans 200 0 0 0 x2.VPWR
rlabel comment 352 600 352 600 4 x2.inv_1
rlabel metal1 352 552 628 648 1 x2.VGND
rlabel metal1 352 1096 628 1192 1 x2.VPWR
flabel pwell 381 583 415 617 0 FreeSans 200 0 0 0 x2.VNB
flabel nwell 381 1127 415 1161 0 FreeSans 200 0 0 0 x2.VPB
flabel locali 164 889 198 923 0 FreeSans 340 0 0 0 x1.Y
flabel locali 164 821 198 855 0 FreeSans 340 0 0 0 x1.Y
flabel locali 72 821 106 855 0 FreeSans 340 0 0 0 x1.A
flabel metal1 29 583 63 617 0 FreeSans 200 0 0 0 x1.VGND
flabel metal1 29 1127 63 1161 0 FreeSans 200 0 0 0 x1.VPWR
rlabel comment 0 600 0 600 4 x1.inv_1
rlabel metal1 0 552 276 648 1 x1.VGND
rlabel metal1 0 1096 276 1192 1 x1.VPWR
flabel pwell 29 583 63 617 0 FreeSans 200 0 0 0 x1.VNB
flabel nwell 29 1127 63 1161 0 FreeSans 200 0 0 0 x1.VPB
<< end >>
