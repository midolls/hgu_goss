magic
tech sky130A
magscale 1 2
timestamp 1701698102
<< nwell >>
rect -2452 8582 -2345 8954
rect -2557 7301 -2294 7964
<< psubdiff >>
rect -49900 6691 -49891 6739
<< poly >>
rect -49498 1455 -49380 1465
rect -49498 1421 -49482 1455
rect -49448 1421 -49380 1455
rect -49498 1411 -49380 1421
rect -48256 1402 -48122 1421
rect -46737 1405 -46590 1432
rect -48256 1392 -48080 1402
rect -48256 1391 -48133 1392
rect -48152 1376 -48133 1391
rect -48149 1358 -48133 1376
rect -48099 1358 -48080 1392
rect -46737 1392 -46554 1405
rect -46737 1387 -46604 1392
rect -48149 1348 -48080 1358
rect -46620 1358 -46604 1387
rect -46570 1358 -46554 1392
rect -44613 1396 -44412 1429
rect -41148 1411 -40990 1430
rect -41191 1398 -40990 1411
rect -44613 1388 -44383 1396
rect -46620 1348 -46554 1358
rect -44449 1383 -44383 1388
rect -44449 1349 -44433 1383
rect -44399 1349 -44383 1383
rect -41191 1364 -41175 1398
rect -41141 1386 -40990 1398
rect -33422 1429 -33241 1442
rect -33422 1395 -33406 1429
rect -33372 1395 -33241 1429
rect -19968 1439 -19697 1452
rect -19968 1405 -19952 1439
rect -19918 1405 -19697 1439
rect -19968 1395 -19697 1405
rect -33422 1386 -33241 1395
rect -41141 1379 -41122 1386
rect -33422 1385 -33353 1386
rect -41141 1364 -41125 1379
rect -41191 1354 -41125 1364
rect -44449 1339 -44383 1349
rect -47255 773 -47123 779
rect -49411 749 -49342 759
rect -49957 714 -49891 727
rect -49957 680 -49941 714
rect -49907 680 -49891 714
rect -49411 715 -49395 749
rect -49361 715 -49342 749
rect -49411 705 -49342 715
rect -48385 749 -48295 762
rect -48385 715 -48345 749
rect -48311 715 -48295 749
rect -48385 705 -48295 715
rect -47255 760 -47075 773
rect -47255 726 -47125 760
rect -47091 726 -47075 760
rect -47255 716 -47075 726
rect -34465 745 -34345 758
rect -47255 710 -47123 716
rect -45117 685 -44972 718
rect -41603 686 -41388 724
rect -34465 711 -34395 745
rect -34361 711 -34345 745
rect -34465 701 -34345 711
rect -20531 725 -20317 735
rect -20531 691 -20367 725
rect -20333 691 -20317 725
rect -20531 686 -20317 691
rect -45117 683 -44971 685
rect -45117 680 -44937 683
rect -41603 680 -41360 686
rect -49957 670 -49891 680
rect -45004 674 -44937 680
rect -41429 678 -41360 680
rect -20386 678 -20317 686
rect -45003 670 -44937 674
rect -45003 636 -44987 670
rect -44953 636 -44937 670
rect -45003 626 -44937 636
rect -41426 673 -41360 678
rect -41426 639 -41410 673
rect -41376 639 -41360 673
rect -41426 629 -41360 639
<< polycont >>
rect -49482 1421 -49448 1455
rect -48133 1358 -48099 1392
rect -46604 1358 -46570 1392
rect -44433 1349 -44399 1383
rect -41175 1364 -41141 1398
rect -33406 1395 -33372 1429
rect -19952 1405 -19918 1439
rect -49941 680 -49907 714
rect -49395 715 -49361 749
rect -48345 715 -48311 749
rect -47125 726 -47091 760
rect -34395 711 -34361 745
rect -20367 691 -20333 725
rect -44987 636 -44953 670
rect -41410 639 -41376 673
<< locali >>
rect -49693 19027 -185 19358
rect -49635 16048 102 16379
rect -49900 6691 -49891 6739
rect -49498 1417 -49487 1460
rect -49442 1417 -49432 1460
rect -48149 1354 -48138 1397
rect -48093 1354 -48083 1397
rect -46620 1354 -46609 1397
rect -46564 1354 -46554 1397
rect -44449 1345 -44438 1388
rect -44393 1345 -44383 1388
rect -41191 1360 -41180 1403
rect -41135 1360 -41125 1403
rect -33422 1391 -33411 1434
rect -33366 1391 -33356 1434
rect -19968 1401 -19957 1444
rect -19912 1401 -19902 1444
rect -49957 676 -49946 719
rect -49901 676 -49891 719
rect -49411 711 -49400 754
rect -49355 711 -49345 754
rect -48361 711 -48350 754
rect -48305 711 -48295 754
rect -47141 722 -47130 765
rect -47085 722 -47075 765
rect -34411 707 -34400 750
rect -34355 707 -34345 750
rect -20383 686 -20373 729
rect -20328 686 -20317 729
rect -45003 632 -44992 675
rect -44947 632 -44937 675
rect -41426 635 -41415 678
rect -41370 635 -41360 678
<< viali >>
rect -49487 1455 -49442 1460
rect -49487 1421 -49482 1455
rect -49482 1421 -49448 1455
rect -49448 1421 -49442 1455
rect -49487 1417 -49442 1421
rect -48138 1392 -48093 1397
rect -48138 1358 -48133 1392
rect -48133 1358 -48099 1392
rect -48099 1358 -48093 1392
rect -48138 1354 -48093 1358
rect -46609 1392 -46564 1397
rect -46609 1358 -46604 1392
rect -46604 1358 -46570 1392
rect -46570 1358 -46564 1392
rect -46609 1354 -46564 1358
rect -44438 1383 -44393 1388
rect -44438 1349 -44433 1383
rect -44433 1349 -44399 1383
rect -44399 1349 -44393 1383
rect -44438 1345 -44393 1349
rect -41180 1398 -41135 1403
rect -41180 1364 -41175 1398
rect -41175 1364 -41141 1398
rect -41141 1364 -41135 1398
rect -41180 1360 -41135 1364
rect -33411 1429 -33366 1434
rect -33411 1395 -33406 1429
rect -33406 1395 -33372 1429
rect -33372 1395 -33366 1429
rect -33411 1391 -33366 1395
rect -19957 1439 -19912 1444
rect -19957 1405 -19952 1439
rect -19952 1405 -19918 1439
rect -19918 1405 -19912 1439
rect -19957 1401 -19912 1405
rect -49946 714 -49901 719
rect -49946 680 -49941 714
rect -49941 680 -49907 714
rect -49907 680 -49901 714
rect -49946 676 -49901 680
rect -49400 749 -49355 754
rect -49400 715 -49395 749
rect -49395 715 -49361 749
rect -49361 715 -49355 749
rect -49400 711 -49355 715
rect -48350 749 -48305 754
rect -48350 715 -48345 749
rect -48345 715 -48311 749
rect -48311 715 -48305 749
rect -48350 711 -48305 715
rect -47130 760 -47085 765
rect -47130 726 -47125 760
rect -47125 726 -47091 760
rect -47091 726 -47085 760
rect -47130 722 -47085 726
rect -34400 745 -34355 750
rect -34400 711 -34395 745
rect -34395 711 -34361 745
rect -34361 711 -34355 745
rect -34400 707 -34355 711
rect -20373 725 -20328 729
rect -20373 691 -20367 725
rect -20367 691 -20333 725
rect -20333 691 -20328 725
rect -20373 686 -20328 691
rect -44992 670 -44947 675
rect -44992 636 -44987 670
rect -44987 636 -44953 670
rect -44953 636 -44947 670
rect -44992 632 -44947 636
rect -41415 673 -41370 678
rect -41415 639 -41410 673
rect -41410 639 -41376 673
rect -41376 639 -41370 673
rect -41415 635 -41370 639
<< metal1 >>
rect -1294 20649 -1264 27894
rect -7726 14613 -7720 14665
rect -7668 14663 -7662 14665
rect -7668 14616 -7607 14663
rect -7668 14613 -7662 14616
rect -46 13742 18 13748
rect -46 13690 -40 13742
rect 12 13734 18 13742
rect 1886 13742 1950 13748
rect 1886 13734 1892 13742
rect 12 13697 1892 13734
rect 12 13690 18 13697
rect -46 13684 18 13690
rect 1886 13690 1892 13697
rect 1944 13690 1950 13742
rect 1886 13684 1950 13690
rect -155 12709 -91 12715
rect -155 12657 -149 12709
rect -97 12702 -91 12709
rect 1775 12711 1839 12717
rect 1775 12702 1781 12711
rect -97 12665 1781 12702
rect -97 12657 -91 12665
rect -155 12651 -91 12657
rect 1775 12659 1781 12665
rect 1833 12659 1839 12711
rect 1775 12653 1839 12659
rect 1883 11866 1947 11872
rect 1883 11814 1889 11866
rect 1941 11814 1947 11866
rect 1883 11808 1947 11814
rect 1786 10836 1850 10842
rect -50095 10792 -49983 10799
rect -50095 10690 -50089 10792
rect -49990 10690 -49983 10792
rect 1786 10784 1792 10836
rect 1844 10831 1850 10836
rect 1844 10794 1889 10831
rect 1844 10784 1850 10794
rect 1786 10778 1850 10784
rect -50095 10685 -49983 10690
rect -50079 9932 -49998 10685
rect -5518 10156 -5512 10208
rect -5460 10156 -5454 10208
rect -110 9906 -104 9916
rect -7939 9876 -104 9906
rect -110 9864 -104 9876
rect -52 9906 -46 9916
rect -52 9876 -37 9906
rect -52 9864 -46 9876
rect -203 9836 -197 9846
rect -7936 9806 -197 9836
rect -203 9794 -197 9806
rect -145 9836 -139 9846
rect -145 9806 -37 9836
rect -145 9794 -139 9806
rect -665 9766 -659 9778
rect -7945 9736 -659 9766
rect -665 9726 -659 9736
rect -607 9766 -601 9778
rect -607 9736 -37 9766
rect -607 9726 -601 9736
rect -943 9697 -937 9708
rect -1537 9696 -937 9697
rect -7939 9666 -937 9696
rect -943 9656 -937 9666
rect -885 9697 -879 9708
rect -885 9696 -247 9697
rect -885 9666 -37 9696
rect -885 9656 -879 9666
rect -793 9627 -787 9638
rect -7943 9597 -787 9627
rect -793 9586 -787 9597
rect -735 9627 -729 9638
rect -735 9597 -37 9627
rect -735 9586 -729 9597
rect -1457 9557 -1451 9568
rect -7944 9527 -1451 9557
rect -1457 9516 -1451 9527
rect -1399 9557 -1393 9568
rect -1399 9527 -37 9557
rect -1399 9516 -1393 9527
rect -385 9488 -379 9498
rect -7945 9458 -379 9488
rect -385 9446 -379 9458
rect -327 9488 -321 9498
rect -327 9458 -37 9488
rect -327 9446 -321 9458
rect -2394 9418 -2388 9429
rect -7941 9388 -2388 9418
rect -2394 9377 -2388 9388
rect -2336 9418 -2330 9429
rect -2336 9388 -37 9418
rect -2336 9377 -2330 9388
rect -2481 9348 -2475 9358
rect -7940 9318 -2475 9348
rect -2481 9306 -2475 9318
rect -2423 9348 -2417 9358
rect -2423 9318 -37 9348
rect -2423 9306 -2417 9318
rect -2843 9278 -2837 9290
rect -7943 9248 -2837 9278
rect -2843 9238 -2837 9248
rect -2785 9278 -2779 9290
rect -2785 9248 -37 9278
rect -2785 9238 -2779 9248
rect -3121 9209 -3115 9220
rect -7945 9179 -3115 9209
rect -3121 9168 -3115 9179
rect -3063 9209 -3057 9220
rect -3063 9179 -37 9209
rect -3063 9168 -3057 9179
rect -2971 9139 -2965 9150
rect -7945 9109 -2965 9139
rect -2971 9098 -2965 9109
rect -2913 9139 -2907 9150
rect -2913 9109 -37 9139
rect -2913 9098 -2907 9109
rect -3635 9069 -3629 9080
rect -7940 9039 -3629 9069
rect -3635 9028 -3629 9039
rect -3577 9069 -3571 9080
rect -3577 9039 -37 9069
rect -3577 9028 -3571 9039
rect -2568 9000 -2562 9010
rect -9006 8970 -2562 9000
rect -2568 8958 -2562 8970
rect -2510 9000 -2504 9010
rect -2510 8970 -37 9000
rect -2510 8958 -2504 8970
rect -7725 8776 -7719 8828
rect -7667 8814 -7661 8828
rect -2494 8816 -2318 8912
rect -7667 8786 -5130 8814
rect -7667 8776 -7661 8786
rect -5158 6724 -5130 8786
rect -2607 8337 -2310 8368
rect -4166 8303 -4162 8337
rect -2603 8303 -2545 8337
rect -2511 8303 -2310 8337
rect -2607 8176 -2310 8303
rect -2603 7536 -2306 7728
rect -2581 6992 -2320 7088
rect -4557 6783 -4551 6799
rect -4582 6748 -4551 6783
rect -4557 6747 -4551 6748
rect -4499 6783 -4493 6799
rect -4499 6748 1004 6783
rect -4499 6747 -4493 6748
rect -5171 6672 -5165 6724
rect -5113 6672 -5107 6724
rect -474 6590 -468 6642
rect -416 6631 -410 6642
rect -288 6631 -282 6641
rect -416 6601 -282 6631
rect -416 6590 -410 6601
rect -288 6589 -282 6601
rect -230 6589 -224 6641
rect -749 6521 -743 6573
rect -691 6561 -685 6573
rect -374 6561 -368 6571
rect -691 6531 -368 6561
rect -691 6521 -685 6531
rect -374 6519 -368 6531
rect -316 6519 -310 6571
rect -1024 6451 -1018 6503
rect -966 6491 -960 6503
rect -461 6491 -455 6502
rect -966 6461 -455 6491
rect -966 6451 -960 6461
rect -461 6450 -455 6461
rect -403 6450 -397 6502
rect -1566 6381 -1560 6433
rect -1508 6422 -1502 6433
rect -547 6422 -541 6432
rect -1508 6392 -541 6422
rect -1508 6381 -1502 6392
rect -547 6380 -541 6392
rect -489 6380 -483 6432
rect -2131 6312 -2125 6364
rect -2073 6352 -2067 6364
rect -634 6352 -628 6363
rect -2073 6322 -628 6352
rect -2073 6312 -2067 6322
rect -634 6311 -628 6322
rect -576 6311 -570 6363
rect -2395 6242 -2389 6294
rect -2337 6283 -2331 6294
rect -720 6283 -714 6293
rect -2337 6253 -714 6283
rect -2337 6242 -2331 6253
rect -720 6241 -714 6253
rect -662 6241 -656 6293
rect -2483 6172 -2477 6224
rect -2425 6213 -2419 6224
rect -806 6213 -800 6223
rect -2425 6183 -800 6213
rect -2425 6172 -2419 6183
rect -806 6171 -800 6183
rect -748 6171 -742 6223
rect -2657 6102 -2651 6154
rect -2599 6143 -2593 6154
rect -892 6143 -886 6153
rect -2599 6113 -886 6143
rect -2599 6102 -2593 6113
rect -892 6101 -886 6113
rect -834 6101 -828 6153
rect -2930 6033 -2924 6085
rect -2872 6073 -2866 6085
rect -979 6073 -973 6084
rect -2872 6043 -973 6073
rect -2872 6033 -2866 6043
rect -979 6032 -973 6043
rect -921 6032 -915 6084
rect -3209 5963 -3203 6015
rect -3151 6004 -3145 6015
rect -1065 6004 -1059 6014
rect -3151 5974 -1059 6004
rect -3151 5963 -3145 5974
rect -1065 5962 -1059 5974
rect -1007 5962 -1001 6014
rect -3756 5894 -3750 5946
rect -3698 5934 -3692 5946
rect -1151 5934 -1145 5944
rect -3698 5904 -1145 5934
rect -3698 5894 -3692 5904
rect -1151 5892 -1145 5904
rect -1093 5892 -1087 5944
rect -4307 5824 -4301 5876
rect -4249 5864 -4243 5876
rect -1238 5864 -1232 5875
rect -4249 5834 -1232 5864
rect -4249 5824 -4243 5834
rect -1238 5823 -1232 5834
rect -1180 5823 -1174 5875
rect -50079 4516 -49998 5205
rect -50094 4511 -49982 4516
rect -50094 4409 -50087 4511
rect -49988 4409 -49982 4511
rect -50094 4402 -49982 4409
rect -49501 1468 -49429 1474
rect -49501 1411 -49495 1468
rect -49435 1411 -49429 1468
rect -19971 1452 -19899 1458
rect -33425 1442 -33353 1448
rect -41194 1411 -41122 1417
rect -49501 1405 -49429 1411
rect -48152 1405 -48080 1411
rect -48152 1348 -48146 1405
rect -48086 1348 -48080 1405
rect -48152 1342 -48080 1348
rect -46623 1405 -46551 1411
rect -46623 1348 -46617 1405
rect -46557 1348 -46551 1405
rect -46623 1342 -46551 1348
rect -44452 1396 -44380 1402
rect -44452 1339 -44446 1396
rect -44386 1339 -44380 1396
rect -41194 1354 -41188 1411
rect -41128 1354 -41122 1411
rect -33425 1385 -33419 1442
rect -33359 1385 -33353 1442
rect -19971 1395 -19965 1452
rect -19905 1395 -19899 1452
rect -19971 1389 -19899 1395
rect -33425 1379 -33353 1385
rect -41194 1348 -41122 1354
rect -44452 1333 -44380 1339
rect -512 972 -506 1024
rect -454 1014 -448 1024
rect -454 984 15324 1014
rect -454 972 -448 984
rect 36 902 42 954
rect 94 944 100 954
rect 94 914 15324 944
rect 94 902 100 914
rect 303 833 309 885
rect 361 874 367 885
rect 361 844 15324 874
rect 361 833 367 844
rect -47144 773 -47072 779
rect -49414 762 -49342 767
rect -49960 727 -49888 733
rect -49960 670 -49954 727
rect -49894 670 -49888 727
rect -49414 705 -49408 762
rect -49348 705 -49342 762
rect -49414 699 -49342 705
rect -48364 762 -48292 768
rect -48364 705 -48358 762
rect -48298 705 -48292 762
rect -47144 716 -47138 773
rect -47078 716 -47072 773
rect -47144 710 -47072 716
rect -34414 758 -34342 764
rect 589 763 595 815
rect 647 805 653 815
rect 647 775 15324 805
rect 647 763 653 775
rect -48364 699 -48292 705
rect -34414 701 -34408 758
rect -34348 701 -34342 758
rect -34414 695 -34342 701
rect -20386 735 -20314 741
rect -49960 664 -49888 670
rect -45006 683 -44934 689
rect -45006 626 -45000 683
rect -44940 626 -44934 683
rect -45006 620 -44934 626
rect -41429 686 -41357 692
rect -41429 629 -41423 686
rect -41363 629 -41357 686
rect -20386 678 -20380 735
rect -20320 678 -20314 735
rect 816 694 822 746
rect 874 735 880 746
rect 874 705 15324 735
rect 874 694 880 705
rect -20386 672 -20314 678
rect -41429 623 -41357 629
rect 952 624 958 676
rect 1010 666 1016 676
rect 1010 636 15324 666
rect 1010 624 1016 636
rect 1288 554 1294 606
rect 1346 596 1352 606
rect 1346 566 15324 596
rect 1346 554 1352 566
rect 1834 484 1840 536
rect 1892 526 1898 536
rect 1892 496 15324 526
rect 1892 484 1898 496
rect 2381 415 2387 467
rect 2439 456 2445 467
rect 2439 426 15324 456
rect 2439 415 2445 426
rect 2667 345 2673 397
rect 2725 387 2731 397
rect 2725 357 15324 387
rect 2725 345 2731 357
rect 2933 275 2939 327
rect 2991 317 2997 327
rect 2991 287 15324 317
rect 2991 275 2997 287
rect 3178 206 3184 258
rect 3236 247 3242 258
rect 3236 217 15324 247
rect 3236 206 3242 217
rect 3316 137 3322 189
rect 3374 178 3380 189
rect 3374 148 15324 178
rect 3374 137 3380 148
rect -19963 -1898 -19899 -1892
rect -19963 -1950 -19957 -1898
rect -19905 -1922 -19899 -1898
rect 676 -1922 682 -1910
rect -19905 -1950 682 -1922
rect -19963 -1952 682 -1950
rect -19963 -1957 -19899 -1952
rect 676 -1962 682 -1952
rect 734 -1922 740 -1910
rect 734 -1952 3482 -1922
rect 734 -1962 740 -1952
rect -33422 -1973 -33358 -1967
rect -33422 -2025 -33416 -1973
rect -33364 -1991 -33358 -1973
rect -396 -1991 -390 -1980
rect -33364 -2021 -390 -1991
rect -33364 -2025 -33358 -2021
rect -33422 -2032 -33358 -2025
rect -396 -2032 -390 -2021
rect -338 -1991 -332 -1980
rect -338 -2021 3482 -1991
rect -338 -2032 -332 -2021
rect -41201 -2042 -41137 -2036
rect -41201 -2094 -41195 -2042
rect -41143 -2061 -41137 -2042
rect 268 -2061 274 -2050
rect -41143 -2091 274 -2061
rect -41143 -2094 -41137 -2091
rect -44447 -2106 -44383 -2100
rect -41201 -2101 -41137 -2094
rect 268 -2102 274 -2091
rect 326 -2061 332 -2050
rect 326 -2091 3482 -2061
rect 326 -2102 332 -2091
rect -44447 -2158 -44441 -2106
rect -44389 -2131 -44383 -2106
rect 118 -2131 124 -2120
rect -44389 -2158 124 -2131
rect -44447 -2161 124 -2158
rect -44447 -2165 -44383 -2161
rect 118 -2172 124 -2161
rect 176 -2131 182 -2120
rect 176 -2161 3482 -2131
rect 176 -2172 182 -2161
rect -46618 -2183 -46554 -2177
rect -46618 -2235 -46612 -2183
rect -46560 -2200 -46554 -2183
rect 396 -2200 402 -2190
rect -46560 -2230 402 -2200
rect -46560 -2235 -46554 -2230
rect -46618 -2242 -46554 -2235
rect 396 -2242 402 -2230
rect 454 -2200 460 -2190
rect 454 -2230 3482 -2200
rect 454 -2242 460 -2230
rect -48148 -2252 -48084 -2246
rect -48148 -2304 -48142 -2252
rect -48090 -2270 -48084 -2252
rect 818 -2270 824 -2258
rect -48090 -2300 824 -2270
rect -48090 -2304 -48084 -2300
rect -48148 -2311 -48084 -2304
rect 818 -2310 824 -2300
rect 876 -2270 882 -2258
rect 876 -2300 3482 -2270
rect 876 -2310 882 -2300
rect -49498 -2330 -49434 -2324
rect -49498 -2382 -49492 -2330
rect -49440 -2340 -49434 -2330
rect 952 -2340 958 -2328
rect -49440 -2370 958 -2340
rect -49440 -2382 -49434 -2370
rect 952 -2380 958 -2370
rect 1010 -2340 1016 -2328
rect 1010 -2370 3482 -2340
rect 1010 -2380 1016 -2370
rect -49498 -2389 -49434 -2382
rect -20387 -2451 -20381 -2399
rect -20329 -2410 -20323 -2399
rect 3030 -2410 3036 -2398
rect -20329 -2440 3036 -2410
rect -20329 -2451 -20323 -2440
rect 3030 -2450 3036 -2440
rect 3088 -2410 3094 -2398
rect 3088 -2440 3482 -2410
rect 3088 -2450 3094 -2440
rect -34410 -2459 -34346 -2453
rect -34410 -2511 -34404 -2459
rect -34352 -2479 -34346 -2459
rect 1958 -2479 1964 -2468
rect -34352 -2509 1964 -2479
rect -34352 -2511 -34346 -2509
rect -34410 -2518 -34346 -2511
rect 1958 -2520 1964 -2509
rect 2016 -2479 2022 -2468
rect 2016 -2509 3482 -2479
rect 2016 -2520 2022 -2509
rect -41424 -2530 -41360 -2524
rect -41424 -2582 -41418 -2530
rect -41366 -2549 -41360 -2530
rect 2622 -2549 2628 -2538
rect -41366 -2579 2628 -2549
rect -41366 -2582 -41360 -2579
rect -41424 -2589 -41360 -2582
rect 2622 -2590 2628 -2579
rect 2680 -2549 2686 -2538
rect 2680 -2579 3482 -2549
rect 2680 -2590 2686 -2579
rect -45001 -2600 -44937 -2594
rect -45001 -2652 -44995 -2600
rect -44943 -2618 -44937 -2600
rect 2472 -2618 2478 -2608
rect -44943 -2648 2478 -2618
rect -44943 -2652 -44937 -2648
rect 1878 -2649 2478 -2648
rect -45001 -2659 -44937 -2652
rect 2472 -2660 2478 -2649
rect 2530 -2618 2536 -2608
rect 2530 -2648 3482 -2618
rect 2530 -2649 3168 -2648
rect 2530 -2660 2536 -2649
rect -47141 -2671 -47077 -2665
rect -47141 -2723 -47135 -2671
rect -47083 -2688 -47077 -2671
rect 2750 -2688 2756 -2678
rect -47083 -2718 2756 -2688
rect -47083 -2723 -47077 -2718
rect -47141 -2730 -47077 -2723
rect 2750 -2730 2756 -2718
rect 2808 -2688 2814 -2678
rect 2808 -2718 3482 -2688
rect 2808 -2730 2814 -2718
rect -48360 -2739 -48296 -2733
rect -48360 -2791 -48354 -2739
rect -48302 -2758 -48296 -2739
rect 3177 -2758 3183 -2746
rect -48302 -2788 3183 -2758
rect -48302 -2791 -48296 -2788
rect -48360 -2798 -48296 -2791
rect 3177 -2798 3183 -2788
rect 3235 -2758 3241 -2746
rect 3235 -2788 3482 -2758
rect 3235 -2798 3241 -2788
rect -49356 -2818 -49292 -2812
rect -49356 -2870 -49350 -2818
rect -49298 -2828 -49292 -2818
rect 3321 -2828 3327 -2816
rect -49298 -2858 3327 -2828
rect -49298 -2870 -49292 -2858
rect 3321 -2868 3327 -2858
rect 3379 -2828 3385 -2816
rect 3379 -2858 3481 -2828
rect 3379 -2868 3385 -2858
rect -49356 -2877 -49292 -2870
<< via1 >>
rect -7720 14613 -7668 14665
rect -40 13690 12 13742
rect 1892 13690 1944 13742
rect -149 12657 -97 12709
rect 1781 12659 1833 12711
rect 1889 11814 1941 11866
rect -50089 10690 -49990 10792
rect 1792 10784 1844 10836
rect -5512 10156 -5460 10208
rect -104 9864 -52 9916
rect -197 9794 -145 9846
rect -659 9726 -607 9778
rect -937 9656 -885 9708
rect -787 9586 -735 9638
rect -1451 9516 -1399 9568
rect -379 9446 -327 9498
rect -2388 9377 -2336 9429
rect -2475 9306 -2423 9358
rect -2837 9238 -2785 9290
rect -3115 9168 -3063 9220
rect -2965 9098 -2913 9150
rect -3629 9028 -3577 9080
rect -2562 8958 -2510 9010
rect -7719 8776 -7667 8828
rect -4551 6747 -4499 6799
rect -5165 6672 -5113 6724
rect -468 6590 -416 6642
rect -282 6589 -230 6641
rect -743 6521 -691 6573
rect -368 6519 -316 6571
rect -1018 6451 -966 6503
rect -455 6450 -403 6502
rect -1560 6381 -1508 6433
rect -541 6380 -489 6432
rect -2125 6312 -2073 6364
rect -628 6311 -576 6363
rect -2389 6242 -2337 6294
rect -714 6241 -662 6293
rect -2477 6172 -2425 6224
rect -800 6171 -748 6223
rect -2651 6102 -2599 6154
rect -886 6101 -834 6153
rect -2924 6033 -2872 6085
rect -973 6032 -921 6084
rect -3203 5963 -3151 6015
rect -1059 5962 -1007 6014
rect -3750 5894 -3698 5946
rect -1145 5892 -1093 5944
rect -4301 5824 -4249 5876
rect -1232 5823 -1180 5875
rect -50087 4409 -49988 4511
rect -49495 1460 -49435 1468
rect -49495 1417 -49487 1460
rect -49487 1417 -49442 1460
rect -49442 1417 -49435 1460
rect -49495 1411 -49435 1417
rect -48146 1397 -48086 1405
rect -48146 1354 -48138 1397
rect -48138 1354 -48093 1397
rect -48093 1354 -48086 1397
rect -48146 1348 -48086 1354
rect -46617 1397 -46557 1405
rect -46617 1354 -46609 1397
rect -46609 1354 -46564 1397
rect -46564 1354 -46557 1397
rect -46617 1348 -46557 1354
rect -44446 1388 -44386 1396
rect -44446 1345 -44438 1388
rect -44438 1345 -44393 1388
rect -44393 1345 -44386 1388
rect -44446 1339 -44386 1345
rect -41188 1403 -41128 1411
rect -41188 1360 -41180 1403
rect -41180 1360 -41135 1403
rect -41135 1360 -41128 1403
rect -41188 1354 -41128 1360
rect -33419 1434 -33359 1442
rect -33419 1391 -33411 1434
rect -33411 1391 -33366 1434
rect -33366 1391 -33359 1434
rect -33419 1385 -33359 1391
rect -19965 1444 -19905 1452
rect -19965 1401 -19957 1444
rect -19957 1401 -19912 1444
rect -19912 1401 -19905 1444
rect -19965 1395 -19905 1401
rect -506 972 -454 1024
rect 42 902 94 954
rect 309 833 361 885
rect -49954 719 -49894 727
rect -49954 676 -49946 719
rect -49946 676 -49901 719
rect -49901 676 -49894 719
rect -49954 670 -49894 676
rect -49408 754 -49348 762
rect -49408 711 -49400 754
rect -49400 711 -49355 754
rect -49355 711 -49348 754
rect -49408 705 -49348 711
rect -48358 754 -48298 762
rect -48358 711 -48350 754
rect -48350 711 -48305 754
rect -48305 711 -48298 754
rect -48358 705 -48298 711
rect -47138 765 -47078 773
rect -47138 722 -47130 765
rect -47130 722 -47085 765
rect -47085 722 -47078 765
rect -47138 716 -47078 722
rect 595 763 647 815
rect -34408 750 -34348 758
rect -34408 707 -34400 750
rect -34400 707 -34355 750
rect -34355 707 -34348 750
rect -34408 701 -34348 707
rect -45000 675 -44940 683
rect -45000 632 -44992 675
rect -44992 632 -44947 675
rect -44947 632 -44940 675
rect -45000 626 -44940 632
rect -41423 678 -41363 686
rect -41423 635 -41415 678
rect -41415 635 -41370 678
rect -41370 635 -41363 678
rect -41423 629 -41363 635
rect -20380 729 -20320 735
rect -20380 686 -20373 729
rect -20373 686 -20328 729
rect -20328 686 -20320 729
rect -20380 678 -20320 686
rect 822 694 874 746
rect 958 624 1010 676
rect 1294 554 1346 606
rect 1840 484 1892 536
rect 2387 415 2439 467
rect 2673 345 2725 397
rect 2939 275 2991 327
rect 3184 206 3236 258
rect 3322 137 3374 189
rect -19957 -1950 -19905 -1898
rect 682 -1962 734 -1910
rect -33416 -2025 -33364 -1973
rect -390 -2032 -338 -1980
rect -41195 -2094 -41143 -2042
rect 274 -2102 326 -2050
rect -44441 -2158 -44389 -2106
rect 124 -2172 176 -2120
rect -46612 -2235 -46560 -2183
rect 402 -2242 454 -2190
rect -48142 -2304 -48090 -2252
rect 824 -2310 876 -2258
rect -49492 -2382 -49440 -2330
rect 958 -2380 1010 -2328
rect -20381 -2451 -20329 -2399
rect 3036 -2450 3088 -2398
rect -34404 -2511 -34352 -2459
rect 1964 -2520 2016 -2468
rect -41418 -2582 -41366 -2530
rect 2628 -2590 2680 -2538
rect -44995 -2652 -44943 -2600
rect 2478 -2660 2530 -2608
rect -47135 -2723 -47083 -2671
rect 2756 -2730 2808 -2678
rect -48354 -2791 -48302 -2739
rect 3183 -2798 3235 -2746
rect -49350 -2870 -49298 -2818
rect 3327 -2868 3379 -2816
<< metal2 >>
rect -316 18304 -119 18313
rect -49826 18264 -49660 18273
rect -49826 18120 -49817 18264
rect -49669 18120 -49660 18264
rect -49826 18110 -49660 18120
rect -316 18119 -308 18304
rect -128 18224 -119 18304
rect -128 18191 6 18224
rect -128 18119 -119 18191
rect -316 18110 -119 18119
rect -49767 18093 -49722 18110
rect -49984 17276 -49818 17285
rect -49984 17132 -49975 17276
rect -49827 17132 -49818 17276
rect -49984 17122 -49818 17132
rect -49917 17105 -49844 17122
rect -49877 14572 -49844 17105
rect -50109 10801 -49970 10811
rect -50109 10680 -50099 10801
rect -49979 10680 -49970 10801
rect -50109 10670 -49970 10680
rect -49877 8497 -49843 14572
rect -49767 8637 -49733 18093
rect -427 17304 -230 17313
rect -427 17119 -419 17304
rect -239 17224 -230 17304
rect -239 17191 -105 17224
rect -239 17119 -230 17191
rect -427 17110 -230 17119
rect -7726 14613 -7720 14665
rect -7668 14613 -7662 14665
rect -7712 8828 -7684 14613
rect -142 12715 -105 17191
rect -31 13748 6 18191
rect -46 13742 18 13748
rect -46 13690 -40 13742
rect 12 13690 18 13742
rect -46 13684 18 13690
rect 1886 13742 1950 13748
rect 1886 13690 1892 13742
rect 1944 13690 1950 13742
rect 1886 13684 1950 13690
rect -155 12709 -91 12715
rect -155 12657 -149 12709
rect -97 12657 -91 12709
rect -155 12651 -91 12657
rect 1775 12711 1839 12717
rect 1775 12659 1781 12711
rect 1833 12659 1839 12711
rect 1775 12653 1839 12659
rect 1789 10842 1826 12653
rect 1900 11872 1937 13684
rect 1883 11866 1947 11872
rect 1883 11814 1889 11866
rect 1941 11814 1947 11866
rect 1883 11808 1947 11814
rect 1786 10836 1850 10842
rect 1786 10784 1792 10836
rect 1844 10784 1850 10836
rect 1786 10778 1850 10784
rect -5518 10156 -5512 10208
rect -5460 10156 -5454 10208
rect -7725 8776 -7719 8828
rect -7667 8776 -7661 8828
rect -5498 8739 -5470 10156
rect -110 9864 -104 9916
rect -52 9864 -46 9916
rect -203 9794 -197 9846
rect -145 9794 -139 9846
rect -665 9726 -659 9778
rect -607 9726 -601 9778
rect -943 9656 -937 9708
rect -885 9656 -879 9708
rect -1457 9516 -1451 9568
rect -1399 9516 -1393 9568
rect -2394 9377 -2388 9429
rect -2336 9377 -2330 9429
rect -2481 9306 -2475 9358
rect -2423 9306 -2417 9358
rect -2843 9238 -2837 9290
rect -2785 9238 -2779 9290
rect -3121 9168 -3115 9220
rect -3063 9168 -3057 9220
rect -3635 9028 -3629 9080
rect -3577 9028 -3571 9080
rect -3624 8944 -3583 9028
rect -3105 8944 -3064 9168
rect -2971 9098 -2965 9150
rect -2913 9098 -2907 9150
rect -2961 8944 -2920 9098
rect -2829 8944 -2788 9238
rect -2568 8958 -2562 9010
rect -2510 8958 -2504 9010
rect -2551 8944 -2510 8958
rect -49791 8628 -49717 8637
rect -49791 8572 -49782 8628
rect -49726 8572 -49717 8628
rect -49791 8563 -49717 8572
rect -49894 8488 -49819 8497
rect -49894 8432 -49884 8488
rect -49828 8432 -49819 8488
rect -49894 8423 -49819 8432
rect -49876 6739 -49842 8423
rect -49900 6730 -49818 6739
rect -49900 6674 -49891 6730
rect -49828 6674 -49818 6730
rect -49900 6665 -49818 6674
rect -49767 6605 -49733 8563
rect -4557 6747 -4551 6799
rect -4499 6747 -4493 6799
rect -5171 6672 -5165 6724
rect -5113 6672 -5107 6724
rect -49800 6596 -49726 6605
rect -49800 6540 -49791 6596
rect -49735 6540 -49726 6596
rect -49800 6531 -49726 6540
rect -4295 5876 -4253 6958
rect -3746 5946 -3704 6953
rect -3198 6015 -3156 6955
rect -2918 6085 -2876 6956
rect -2646 6154 -2604 6952
rect -2472 6224 -2430 9306
rect -2383 6294 -2341 9377
rect -1446 8944 -1405 9516
rect -927 8944 -886 9656
rect -793 9586 -787 9638
rect -735 9586 -729 9638
rect -783 8944 -742 9586
rect -651 8944 -610 9726
rect -385 9446 -379 9498
rect -327 9446 -321 9498
rect -373 8944 -332 9446
rect -2119 6364 -2077 6949
rect -1555 6433 -1513 6954
rect -1012 6503 -970 6957
rect -738 6573 -696 6957
rect -463 6642 -421 6965
rect -474 6590 -468 6642
rect -416 6590 -410 6642
rect -288 6589 -282 6641
rect -230 6589 -224 6641
rect -749 6521 -743 6573
rect -691 6521 -685 6573
rect -374 6519 -368 6571
rect -316 6519 -310 6571
rect -1024 6451 -1018 6503
rect -966 6451 -960 6503
rect -461 6450 -455 6502
rect -403 6450 -397 6502
rect -1566 6381 -1560 6433
rect -1508 6381 -1502 6433
rect -547 6380 -541 6432
rect -489 6380 -483 6432
rect -2131 6312 -2125 6364
rect -2073 6312 -2067 6364
rect -634 6311 -628 6363
rect -576 6311 -570 6363
rect -2395 6242 -2389 6294
rect -2337 6242 -2331 6294
rect -720 6241 -714 6293
rect -662 6241 -656 6293
rect -2483 6172 -2477 6224
rect -2425 6172 -2419 6224
rect -806 6171 -800 6223
rect -748 6171 -742 6223
rect -2657 6102 -2651 6154
rect -2599 6102 -2593 6154
rect -892 6101 -886 6153
rect -834 6101 -828 6153
rect -2930 6033 -2924 6085
rect -2872 6033 -2866 6085
rect -979 6032 -973 6084
rect -921 6032 -915 6084
rect -3209 5963 -3203 6015
rect -3151 5963 -3145 6015
rect -1065 5962 -1059 6014
rect -1007 5962 -1001 6014
rect -3756 5894 -3750 5946
rect -3698 5894 -3692 5946
rect -1151 5892 -1145 5944
rect -1093 5892 -1087 5944
rect -4307 5824 -4301 5876
rect -4249 5824 -4243 5876
rect -1238 5823 -1232 5875
rect -1180 5823 -1174 5875
rect -1222 5715 -1180 5823
rect -1140 5715 -1098 5892
rect -1056 5715 -1014 5962
rect -968 5715 -926 6032
rect -881 5715 -839 6101
rect -795 5715 -753 6171
rect -709 5715 -667 6241
rect -622 5715 -580 6311
rect -536 5715 -494 6380
rect -450 5715 -408 6450
rect -363 5715 -321 6519
rect -278 5715 -236 6589
rect -191 5716 -149 9794
rect -104 5716 -62 9864
rect -50107 4521 -49968 4531
rect -50107 4400 -50098 4521
rect -49978 4400 -49968 4521
rect -50107 4390 -49968 4400
rect -49501 1468 -49429 1474
rect -49501 1411 -49495 1468
rect -49435 1411 -49429 1468
rect -19971 1452 -19899 1458
rect -33425 1442 -33353 1448
rect -41194 1411 -41122 1417
rect -49501 1405 -49429 1411
rect -48152 1405 -48080 1411
rect -49960 727 -49888 733
rect -49960 670 -49954 727
rect -49894 670 -49888 727
rect -49960 664 -49888 670
rect -49490 -2324 -49442 1405
rect -48152 1348 -48146 1405
rect -48086 1348 -48080 1405
rect -48152 1342 -48080 1348
rect -46623 1405 -46551 1411
rect -46623 1348 -46617 1405
rect -46557 1348 -46551 1405
rect -46623 1342 -46551 1348
rect -44452 1396 -44380 1402
rect -49342 767 -49300 769
rect -49414 762 -49300 767
rect -49414 705 -49408 762
rect -49348 705 -49300 762
rect -49414 699 -49300 705
rect -48364 762 -48292 768
rect -48364 705 -48358 762
rect -48298 705 -48292 762
rect -48364 699 -48292 705
rect -49498 -2330 -49434 -2324
rect -49498 -2382 -49492 -2330
rect -49440 -2382 -49434 -2330
rect -49498 -2389 -49434 -2382
rect -49348 -2812 -49300 699
rect -48352 -2733 -48304 699
rect -48140 -2246 -48092 1342
rect -47144 773 -47072 779
rect -47144 716 -47138 773
rect -47078 716 -47072 773
rect -47144 710 -47072 716
rect -48148 -2252 -48084 -2246
rect -48148 -2304 -48142 -2252
rect -48090 -2304 -48084 -2252
rect -48148 -2311 -48084 -2304
rect -47132 -2665 -47084 710
rect -46610 -2177 -46562 1342
rect -44452 1339 -44446 1396
rect -44386 1339 -44380 1396
rect -41194 1354 -41188 1411
rect -41128 1354 -41122 1411
rect -33425 1385 -33419 1442
rect -33359 1385 -33353 1442
rect -19971 1395 -19965 1452
rect -19905 1395 -19899 1452
rect -19971 1389 -19899 1395
rect -33425 1379 -33353 1385
rect -41194 1348 -41122 1354
rect -44452 1333 -44380 1339
rect -45006 683 -44934 689
rect -45006 626 -45000 683
rect -44940 626 -44934 683
rect -45006 620 -44934 626
rect -46618 -2183 -46554 -2177
rect -46618 -2235 -46612 -2183
rect -46560 -2235 -46554 -2183
rect -46618 -2242 -46554 -2235
rect -44994 -2594 -44946 620
rect -44439 -2100 -44391 1333
rect -41429 686 -41357 692
rect -41429 629 -41423 686
rect -41363 629 -41357 686
rect -41429 623 -41357 629
rect -44447 -2106 -44383 -2100
rect -44447 -2158 -44441 -2106
rect -44389 -2158 -44383 -2106
rect -44447 -2165 -44383 -2158
rect -41416 -2524 -41368 623
rect -41192 -2036 -41144 1348
rect -34414 758 -34342 764
rect -34414 701 -34408 758
rect -34348 701 -34342 758
rect -34414 695 -34342 701
rect -41201 -2042 -41137 -2036
rect -41201 -2094 -41195 -2042
rect -41143 -2094 -41137 -2042
rect -41201 -2101 -41137 -2094
rect -34401 -2453 -34353 695
rect -33413 -1967 -33365 1379
rect -20386 735 -20314 741
rect -20386 678 -20380 735
rect -20320 678 -20314 735
rect -20386 672 -20314 678
rect -33422 -1973 -33358 -1967
rect -33422 -2025 -33416 -1973
rect -33364 -2025 -33358 -1973
rect -33422 -2032 -33358 -2025
rect -20377 -2399 -20329 672
rect -19958 -1892 -19910 1389
rect -512 972 -506 1024
rect -454 972 -448 1024
rect -1062 138 -1020 906
rect -500 93 -458 972
rect 36 902 42 954
rect 94 902 100 954
rect 46 93 88 902
rect 303 833 309 885
rect 361 833 367 885
rect 314 93 356 833
rect 589 763 595 815
rect 647 763 653 815
rect 601 93 643 763
rect 816 694 822 746
rect 874 694 880 746
rect -19963 -1898 -19899 -1892
rect -19963 -1950 -19957 -1898
rect -19905 -1950 -19899 -1898
rect -19963 -1957 -19899 -1950
rect -385 -1980 -344 -1718
rect -396 -2032 -390 -1980
rect -338 -2032 -332 -1980
rect 134 -2120 175 -1838
rect 278 -2050 319 -1791
rect 268 -2102 274 -2050
rect 326 -2102 332 -2050
rect 118 -2172 124 -2120
rect 176 -2172 182 -2120
rect 410 -2190 451 -1903
rect 676 -1962 682 -1910
rect 734 -1962 740 -1910
rect 396 -2242 402 -2190
rect 454 -2242 460 -2190
rect 827 -2258 869 694
rect 952 624 958 676
rect 1010 624 1016 676
rect 818 -2310 824 -2258
rect 876 -2310 882 -2258
rect 963 -2328 1005 624
rect 1288 554 1294 606
rect 1346 554 1352 606
rect 1300 93 1342 554
rect 1834 484 1840 536
rect 1892 484 1898 536
rect 1846 93 1888 484
rect 2381 415 2387 467
rect 2439 415 2445 467
rect 2392 93 2434 415
rect 2667 345 2673 397
rect 2725 345 2731 397
rect 2679 93 2721 345
rect 2933 275 2939 327
rect 2991 275 2997 327
rect 2944 93 2986 275
rect 3178 206 3184 258
rect 3236 206 3242 258
rect 952 -2380 958 -2328
rect 1010 -2380 1016 -2328
rect -20387 -2451 -20381 -2399
rect -20329 -2451 -20323 -2399
rect -34410 -2459 -34346 -2453
rect -34410 -2511 -34404 -2459
rect -34352 -2511 -34346 -2459
rect 1969 -2468 2010 -1625
rect -34410 -2518 -34346 -2511
rect 1958 -2520 1964 -2468
rect 2016 -2520 2022 -2468
rect -41424 -2530 -41360 -2524
rect -41424 -2582 -41418 -2530
rect -41366 -2582 -41360 -2530
rect -41424 -2589 -41360 -2582
rect -45001 -2600 -44937 -2594
rect -45001 -2652 -44995 -2600
rect -44943 -2652 -44937 -2600
rect 2488 -2608 2529 -1766
rect 2632 -2538 2673 -1680
rect 2622 -2590 2628 -2538
rect 2680 -2590 2686 -2538
rect -45001 -2659 -44937 -2652
rect 2472 -2660 2478 -2608
rect 2530 -2660 2536 -2608
rect -47141 -2671 -47077 -2665
rect -47141 -2723 -47135 -2671
rect -47083 -2723 -47077 -2671
rect 2764 -2678 2805 -1820
rect 3042 -2398 3083 -1892
rect 3030 -2450 3036 -2398
rect 3088 -2450 3094 -2398
rect -47141 -2730 -47077 -2723
rect 2750 -2730 2756 -2678
rect 2808 -2730 2814 -2678
rect -48360 -2739 -48296 -2733
rect -48360 -2791 -48354 -2739
rect -48302 -2791 -48296 -2739
rect 3189 -2746 3231 206
rect 3316 137 3322 189
rect 3374 137 3380 189
rect -48360 -2798 -48296 -2791
rect 3177 -2798 3183 -2746
rect 3235 -2798 3241 -2746
rect -49356 -2818 -49292 -2812
rect 3327 -2816 3369 137
rect -49356 -2870 -49350 -2818
rect -49298 -2870 -49292 -2818
rect 3321 -2868 3327 -2816
rect 3379 -2868 3385 -2816
rect -49356 -2877 -49292 -2870
<< via2 >>
rect -49817 18120 -49669 18264
rect -308 18119 -128 18304
rect -49975 17132 -49827 17276
rect -50099 10792 -49979 10801
rect -50099 10690 -50089 10792
rect -50089 10690 -49990 10792
rect -49990 10690 -49979 10792
rect -50099 10680 -49979 10690
rect -419 17119 -239 17304
rect -49782 8572 -49726 8628
rect -49884 8432 -49828 8488
rect -49891 6674 -49828 6730
rect -49791 6540 -49735 6596
rect -50098 4511 -49978 4521
rect -50098 4409 -50087 4511
rect -50087 4409 -49988 4511
rect -49988 4409 -49978 4511
rect -50098 4400 -49978 4409
<< metal3 >>
rect -338 18318 -102 18319
rect -49845 18290 -49640 18296
rect -49845 18093 -49839 18290
rect -49646 18093 -49640 18290
rect -338 18105 -325 18318
rect -114 18105 -102 18318
rect -49845 18087 -49640 18093
rect -449 17318 -213 17319
rect -50003 17302 -49798 17308
rect -50003 17105 -49997 17302
rect -49804 17105 -49798 17302
rect -449 17105 -436 17318
rect -225 17105 -213 17318
rect -50003 17099 -49798 17105
rect -50133 10828 -49945 10835
rect -50133 10652 -50127 10828
rect -49950 10652 -49945 10828
rect -50133 10646 -49945 10652
rect -49791 8628 -49717 8637
rect -49791 8623 -49782 8628
rect -49977 8572 -49782 8623
rect -49726 8572 -49717 8628
rect -49977 8563 -49717 8572
rect -50070 8488 -49819 8497
rect -50070 8437 -49884 8488
rect -49894 8432 -49884 8437
rect -49828 8432 -49819 8488
rect -49894 8423 -49819 8432
rect -9304 7723 -9294 7791
rect -9230 7787 -9220 7791
rect -9230 7727 -8803 7787
rect -7941 7727 -7904 7787
rect -9230 7723 -9220 7727
rect -9304 7405 -9294 7473
rect -9230 7469 -9220 7473
rect -9230 7409 -8803 7469
rect -7941 7409 -7904 7469
rect -9230 7405 -9220 7409
rect -49900 6730 -49818 6739
rect -49900 6726 -49891 6730
rect -50066 6674 -49891 6726
rect -49828 6674 -49818 6730
rect -50066 6666 -49818 6674
rect -49900 6665 -49818 6666
rect -49977 6596 -49726 6605
rect -49977 6545 -49791 6596
rect -49800 6540 -49791 6545
rect -49735 6540 -49726 6596
rect -49800 6531 -49726 6540
rect -50132 4549 -49944 4555
rect -50132 4373 -50127 4549
rect -49950 4373 -49944 4549
rect -50132 4366 -49944 4373
<< via3 >>
rect -49839 18264 -49646 18290
rect -49839 18120 -49817 18264
rect -49817 18120 -49669 18264
rect -49669 18120 -49646 18264
rect -49839 18093 -49646 18120
rect -325 18304 -114 18318
rect -325 18119 -308 18304
rect -308 18119 -128 18304
rect -128 18119 -114 18304
rect -325 18105 -114 18119
rect -49997 17276 -49804 17302
rect -49997 17132 -49975 17276
rect -49975 17132 -49827 17276
rect -49827 17132 -49804 17276
rect -49997 17105 -49804 17132
rect -436 17304 -225 17318
rect -436 17119 -419 17304
rect -419 17119 -239 17304
rect -239 17119 -225 17304
rect -436 17105 -225 17119
rect -50127 10801 -49950 10828
rect -50127 10680 -50099 10801
rect -50099 10680 -49979 10801
rect -49979 10680 -49950 10801
rect -50127 10652 -49950 10680
rect -9294 7723 -9230 7791
rect -9294 7405 -9230 7473
rect -50127 4521 -49950 4549
rect -50127 4400 -50098 4521
rect -50098 4400 -49978 4521
rect -49978 4400 -49950 4521
rect -50127 4373 -49950 4400
<< metal4 >>
rect -462 17329 -201 17330
rect -462 17093 -449 17329
rect -213 17093 -201 17329
rect 1775 12653 1839 12717
rect -50084 12269 -49569 12337
rect -50084 10859 -50006 12269
rect -9312 10856 -9208 10902
rect -9312 7791 -9209 10620
rect -6065 10334 -6010 10340
rect -9312 7723 -9294 7791
rect -9230 7723 -9209 7791
rect -9312 7712 -9209 7723
rect -4916 10302 -4835 10334
rect -4771 10302 -4755 10334
rect -4691 10302 -4675 10334
rect -4611 10302 -4595 10334
rect -4531 10302 -4515 10334
rect -4451 10302 -4435 10340
rect -4371 10302 -4229 10340
rect -4165 10302 -4149 10340
rect -4085 10302 -4069 10340
rect -4005 10302 -3989 10340
rect -3925 10302 -3909 10340
rect -3845 10302 -3829 10340
rect -3765 10302 -3623 10340
rect -3559 10302 -3543 10340
rect -4916 10155 -3542 10302
rect -4916 10063 -4728 10155
rect -4538 10153 -3542 10155
rect -4538 10063 -4334 10153
rect -4916 10061 -4334 10063
rect -4144 10151 -3542 10153
rect -4144 10061 -3927 10151
rect -4916 10059 -3927 10061
rect -3737 10059 -3542 10151
rect -4916 8900 -3542 10059
rect -4916 8899 -4147 8900
rect -4916 8889 -4371 8899
rect -4307 8889 -4147 8899
rect -4083 8897 -3542 8900
rect -4083 8895 -3947 8897
rect -3883 8896 -3542 8897
rect -3883 8895 -3746 8896
rect -3682 8895 -3542 8896
rect -2331 10143 -1367 10302
rect -2331 10051 -2202 10143
rect -2012 10139 -1367 10143
rect -2012 10051 -1776 10139
rect -2331 10047 -1776 10051
rect -1586 10047 -1367 10139
rect -2331 8901 -1367 10047
rect -2331 8900 -1969 8901
rect -4083 8889 -3952 8895
rect -4916 8645 -4504 8889
rect -2331 8858 -2193 8900
rect -2129 8858 -1969 8900
rect -1905 8898 -1367 8901
rect -1905 8858 -1769 8898
rect -1705 8897 -1367 8898
rect -1705 8858 -1568 8897
rect -1504 8858 -1367 8897
rect -4916 8535 -4906 8645
rect -4640 8535 -4504 8645
rect -9312 7473 -9209 7483
rect -9312 7405 -9294 7473
rect -9230 7405 -9209 7473
rect -9312 4676 -9209 7405
rect -4916 6995 -4504 8535
rect -3460 7071 -2483 7099
rect -3460 7067 -2783 7071
rect -3460 7003 -3347 7067
rect -3283 7003 -3042 7067
rect -2978 7007 -2783 7067
rect -2719 7007 -2483 7071
rect -2978 7003 -2483 7007
rect -5304 5674 -5022 6314
rect -3460 5674 -2483 7003
rect -331 6988 141 8917
rect -5304 5380 -1745 5674
rect -5304 5376 -5022 5380
rect -9312 4580 -9208 4676
rect -50084 2927 -50006 4342
rect -50084 2859 -49569 2927
<< via4 >>
rect -338 18318 -102 18329
rect -49868 18290 -49614 18314
rect -49868 18093 -49839 18290
rect -49839 18093 -49646 18290
rect -49646 18093 -49614 18290
rect -338 18105 -325 18318
rect -325 18105 -114 18318
rect -114 18105 -102 18318
rect -338 18093 -102 18105
rect -49868 18065 -49614 18093
rect -50026 17302 -49772 17326
rect -50026 17105 -49997 17302
rect -49997 17105 -49804 17302
rect -49804 17105 -49772 17302
rect -50026 17077 -49772 17105
rect -449 17318 -213 17329
rect -449 17105 -436 17318
rect -436 17105 -225 17318
rect -225 17105 -213 17318
rect -449 17093 -213 17105
rect -50157 10828 -49920 10859
rect -50157 10652 -50127 10828
rect -50127 10652 -49950 10828
rect -49950 10652 -49920 10828
rect -50157 10623 -49920 10652
rect -9380 10620 -9144 10856
rect -50157 4549 -49920 4578
rect -50157 4373 -50127 4549
rect -50127 4373 -49950 4549
rect -49950 4373 -49920 4549
rect -50157 4342 -49920 4373
rect -9380 4344 -9144 4580
<< metal5 >>
rect -49894 18329 -76 18365
rect -49894 18314 -338 18329
rect -49894 18065 -49868 18314
rect -49614 18093 -338 18314
rect -102 18093 -76 18329
rect -49614 18065 -76 18093
rect -49894 18034 -76 18065
rect -50051 17329 -187 17372
rect -50051 17326 -449 17329
rect -50051 17077 -50026 17326
rect -49772 17093 -449 17326
rect -213 17093 -187 17329
rect -49772 17077 -187 17093
rect -50051 17041 -187 17077
rect -50203 10903 -49852 10904
rect -50203 10902 -49437 10903
rect -50203 10859 -9105 10902
rect -50203 10623 -50157 10859
rect -49920 10856 -9105 10859
rect -49920 10623 -9380 10856
rect -50203 10620 -9380 10623
rect -9144 10620 -9105 10856
rect -50203 10570 -9105 10620
rect -50137 10569 -49437 10570
rect -50202 4580 -9105 4626
rect -50202 4578 -9380 4580
rect -50202 4342 -50157 4578
rect -49920 4344 -9380 4578
rect -9144 4344 -9105 4580
rect -49920 4342 -9105 4344
rect -50202 4294 -9105 4342
rect -50202 4292 -49508 4294
use hgu_cdac_half  hgu_cdac_half_0
timestamp 1701696200
transform 1 0 -49110 0 -1 6793
box -459 -645 39606 6322
use hgu_cdac_half  hgu_cdac_half_1
timestamp 1701696200
transform 1 0 -49110 0 1 8403
box -459 -645 39606 6322
use hgu_cdac_sw_buffer  hgu_cdac_sw_buffer_0
timestamp 1699539897
transform -1 0 525 0 -1 -2647
box -270 -2798 1830 -714
use hgu_cdac_sw_buffer  hgu_cdac_sw_buffer_1
timestamp 1699539897
transform -1 0 2879 0 -1 -2643
box -270 -2798 1830 -714
use hgu_cdac_sw_buffer  hgu_cdac_sw_buffer_2
timestamp 1699539897
transform -1 0 -536 0 1 9721
box -270 -2798 1830 -714
use hgu_cdac_sw_buffer  hgu_cdac_sw_buffer_3
timestamp 1699539897
transform -1 0 -2714 0 1 9720
box -270 -2798 1830 -714
use hgu_comp_flat  hgu_comp_flat_0
timestamp 1698719859
transform 1 0 -8242 0 1 8167
box 338 -1940 3788 618
use hgu_sarlogic_flat  hgu_sarlogic_flat_0
timestamp 1700302578
transform 1 0 -9938 0 1 2806
box 2064 -1908 31250 13749
use hgu_tah  hgu_tah_0
timestamp 1701281041
transform 1 0 -51706 0 1 4757
box 339 297 1858 5355
use hgu_vgen_vref  hgu_vgen_vref_0
timestamp 1701018915
transform -1 0 -51162 0 1 -30367
box 0 0 22370 76000
<< end >>
