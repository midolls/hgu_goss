magic
tech sky130A
magscale 1 2
timestamp 1699356299
<< error_s >>
rect -148 2906 -144 2934
rect -120 2904 -116 2906
<< nwell >>
rect -36 2961 2892 3031
rect -13 2937 2892 2961
rect 4348 2950 7276 3031
rect -13 2933 2 2937
rect -42 1819 16670 1890
rect -42 1795 3158 1819
rect 3192 1818 6245 1819
rect 6279 1818 9374 1819
rect 3192 1795 9374 1818
rect 9408 1795 16670 1819
rect -42 1526 16670 1795
rect -38 1107 16782 1201
rect -38 463 16782 513
rect 557 460 3056 463
rect 6353 442 6518 463
rect 7606 460 7761 463
rect 8745 418 8749 463
rect 11116 442 11315 463
rect 12322 462 12601 463
rect 12322 442 12589 462
rect 13510 442 13639 463
rect 14786 462 14911 463
rect 15921 442 16102 463
rect 16736 453 16782 463
rect 15943 419 16009 442
<< pwell >>
rect 10592 710 10646 713
<< psubdiff >>
rect 2 2369 31 2403
rect 65 2369 123 2403
rect 157 2369 215 2403
rect 249 2369 307 2403
rect 341 2369 399 2403
rect 433 2369 491 2403
rect 525 2369 583 2403
rect 617 2369 675 2403
rect 709 2369 767 2403
rect 801 2369 859 2403
rect 893 2369 951 2403
rect 985 2369 1043 2403
rect 1077 2369 1135 2403
rect 1169 2369 1227 2403
rect 1261 2369 1319 2403
rect 1353 2369 1411 2403
rect 1445 2369 1503 2403
rect 1537 2369 1595 2403
rect 1629 2369 1687 2403
rect 1721 2369 1779 2403
rect 1813 2369 1871 2403
rect 1905 2369 1963 2403
rect 1997 2369 2055 2403
rect 2089 2369 2147 2403
rect 2181 2369 2239 2403
rect 2273 2369 2331 2403
rect 2365 2369 2423 2403
rect 2457 2369 2515 2403
rect 2549 2369 2607 2403
rect 2641 2369 2699 2403
rect 2733 2369 2791 2403
rect 2825 2369 2854 2403
rect 4386 2369 4415 2403
rect 4449 2369 4507 2403
rect 4541 2369 4599 2403
rect 4633 2369 4691 2403
rect 4725 2369 4783 2403
rect 4817 2369 4875 2403
rect 4909 2369 4967 2403
rect 5001 2369 5059 2403
rect 5093 2369 5151 2403
rect 5185 2369 5243 2403
rect 5277 2369 5335 2403
rect 5369 2369 5427 2403
rect 5461 2369 5519 2403
rect 5553 2369 5611 2403
rect 5645 2369 5703 2403
rect 5737 2369 5795 2403
rect 5829 2369 5887 2403
rect 5921 2369 5979 2403
rect 6013 2369 6071 2403
rect 6105 2369 6163 2403
rect 6197 2369 6255 2403
rect 6289 2369 6347 2403
rect 6381 2369 6439 2403
rect 6473 2369 6531 2403
rect 6565 2369 6623 2403
rect 6657 2369 6715 2403
rect 6749 2369 6807 2403
rect 6841 2369 6899 2403
rect 6933 2369 6991 2403
rect 7025 2369 7083 2403
rect 7117 2369 7175 2403
rect 7209 2369 7238 2403
rect 0 1227 29 1261
rect 63 1227 121 1261
rect 155 1227 213 1261
rect 247 1227 305 1261
rect 339 1227 397 1261
rect 431 1227 489 1261
rect 523 1227 581 1261
rect 615 1227 673 1261
rect 707 1227 765 1261
rect 799 1227 857 1261
rect 891 1227 949 1261
rect 983 1227 1041 1261
rect 1075 1227 1133 1261
rect 1167 1227 1225 1261
rect 1259 1227 1317 1261
rect 1351 1227 1409 1261
rect 1443 1227 1501 1261
rect 1535 1227 1593 1261
rect 1627 1227 1685 1261
rect 1719 1227 1777 1261
rect 1811 1227 1869 1261
rect 1903 1227 1961 1261
rect 1995 1227 2053 1261
rect 2087 1227 2145 1261
rect 2179 1227 2237 1261
rect 2271 1227 2329 1261
rect 2363 1227 2421 1261
rect 2455 1227 2513 1261
rect 2547 1227 2605 1261
rect 2639 1227 2697 1261
rect 2731 1227 2789 1261
rect 2823 1227 2881 1261
rect 2915 1227 2973 1261
rect 3007 1227 3065 1261
rect 3099 1227 3157 1261
rect 3191 1227 3249 1261
rect 3283 1227 3341 1261
rect 3375 1227 3433 1261
rect 3467 1227 3525 1261
rect 3559 1227 3617 1261
rect 3651 1227 3709 1261
rect 3743 1227 3801 1261
rect 3835 1227 3893 1261
rect 3927 1227 3985 1261
rect 4019 1227 4077 1261
rect 4111 1227 4169 1261
rect 4203 1227 4261 1261
rect 4295 1227 4353 1261
rect 4387 1227 4445 1261
rect 4479 1227 4537 1261
rect 4571 1227 4629 1261
rect 4663 1227 4721 1261
rect 4755 1227 4813 1261
rect 4847 1227 4905 1261
rect 4939 1227 4997 1261
rect 5031 1227 5089 1261
rect 5123 1227 5181 1261
rect 5215 1227 5273 1261
rect 5307 1227 5365 1261
rect 5399 1227 5457 1261
rect 5491 1227 5549 1261
rect 5583 1227 5641 1261
rect 5675 1231 6245 1261
rect 5675 1227 5704 1231
rect 6216 1227 6245 1231
rect 6279 1227 6337 1261
rect 6371 1227 6429 1261
rect 6463 1227 6521 1261
rect 6555 1227 6613 1261
rect 6647 1227 6705 1261
rect 6739 1227 6797 1261
rect 6831 1227 6889 1261
rect 6923 1227 6981 1261
rect 7015 1227 7073 1261
rect 7107 1227 7165 1261
rect 7199 1227 7257 1261
rect 7291 1227 7349 1261
rect 7383 1227 7441 1261
rect 7475 1227 7533 1261
rect 7567 1227 7625 1261
rect 7659 1227 7717 1261
rect 7751 1227 7809 1261
rect 7843 1227 7901 1261
rect 7935 1227 7993 1261
rect 8027 1227 8085 1261
rect 8119 1227 8177 1261
rect 8211 1227 8269 1261
rect 8303 1227 8361 1261
rect 8395 1227 8453 1261
rect 8487 1227 8545 1261
rect 8579 1227 8637 1261
rect 8671 1227 8729 1261
rect 8763 1227 8821 1261
rect 8855 1227 8913 1261
rect 8947 1227 9005 1261
rect 9039 1227 9097 1261
rect 9131 1227 9189 1261
rect 9223 1227 9281 1261
rect 9315 1227 9373 1261
rect 9407 1227 9465 1261
rect 9499 1227 9557 1261
rect 9591 1227 9649 1261
rect 9683 1227 9741 1261
rect 9775 1227 9833 1261
rect 9867 1227 9925 1261
rect 9959 1227 10017 1261
rect 10051 1227 10109 1261
rect 10143 1227 10201 1261
rect 10235 1227 10293 1261
rect 10327 1227 10385 1261
rect 10419 1227 10477 1261
rect 10511 1227 10569 1261
rect 10603 1227 10661 1261
rect 10695 1227 10753 1261
rect 10787 1227 10845 1261
rect 10879 1227 10937 1261
rect 10971 1227 11029 1261
rect 11063 1227 11121 1261
rect 11155 1227 11213 1261
rect 11247 1227 11305 1261
rect 11339 1227 11397 1261
rect 11431 1227 11489 1261
rect 11523 1227 11581 1261
rect 11615 1227 11673 1261
rect 11707 1227 11765 1261
rect 11799 1227 11857 1261
rect 11891 1231 12011 1261
rect 11891 1227 11920 1231
rect 11982 1227 12011 1231
rect 12045 1227 12103 1261
rect 12137 1227 12195 1261
rect 12229 1227 12287 1261
rect 12321 1227 12379 1261
rect 12413 1227 12471 1261
rect 12505 1227 12563 1261
rect 12597 1227 12655 1261
rect 12689 1227 12747 1261
rect 12781 1227 12839 1261
rect 12873 1227 12931 1261
rect 12965 1227 13023 1261
rect 13057 1227 13115 1261
rect 13149 1227 13207 1261
rect 13241 1227 13299 1261
rect 13333 1227 13391 1261
rect 13425 1227 13483 1261
rect 13517 1227 13575 1261
rect 13609 1227 13667 1261
rect 13701 1227 13759 1261
rect 13793 1227 13851 1261
rect 13885 1227 13943 1261
rect 13977 1227 14035 1261
rect 14069 1227 14127 1261
rect 14161 1227 14219 1261
rect 14253 1227 14311 1261
rect 14345 1227 14403 1261
rect 14437 1227 14495 1261
rect 14529 1227 14587 1261
rect 14621 1227 14679 1261
rect 14713 1227 14771 1261
rect 14805 1227 14863 1261
rect 14897 1227 14955 1261
rect 14989 1227 15047 1261
rect 15081 1227 15139 1261
rect 15173 1227 15231 1261
rect 15265 1227 15323 1261
rect 15357 1227 15415 1261
rect 15449 1227 15507 1261
rect 15541 1227 15599 1261
rect 15633 1227 15691 1261
rect 15725 1227 15783 1261
rect 15817 1227 15875 1261
rect 15909 1227 15967 1261
rect 16001 1227 16059 1261
rect 16093 1227 16151 1261
rect 16185 1227 16243 1261
rect 16277 1227 16335 1261
rect 16369 1227 16427 1261
rect 16461 1227 16519 1261
rect 16553 1231 16614 1261
rect 16553 1227 16582 1231
rect -1 543 29 573
rect 0 539 29 543
rect 63 539 121 573
rect 155 539 213 573
rect 247 539 305 573
rect 339 539 397 573
rect 431 539 489 573
rect 523 539 581 573
rect 615 539 673 573
rect 707 539 765 573
rect 799 539 857 573
rect 891 539 949 573
rect 983 539 1041 573
rect 1075 539 1133 573
rect 1167 539 1225 573
rect 1259 539 1317 573
rect 1351 539 1409 573
rect 1443 539 1501 573
rect 1535 539 1593 573
rect 1627 539 1685 573
rect 1719 539 1777 573
rect 1811 539 1869 573
rect 1903 539 1961 573
rect 1995 539 2053 573
rect 2087 539 2145 573
rect 2179 539 2237 573
rect 2271 539 2329 573
rect 2363 539 2421 573
rect 2455 539 2513 573
rect 2547 539 2605 573
rect 2639 539 2697 573
rect 2731 539 2789 573
rect 2823 539 2881 573
rect 2915 539 2973 573
rect 3007 539 3065 573
rect 3099 539 3157 573
rect 3191 539 3249 573
rect 3283 539 3341 573
rect 3375 539 3433 573
rect 3467 539 3525 573
rect 3559 539 3617 573
rect 3651 539 3709 573
rect 3743 539 3801 573
rect 3835 539 3893 573
rect 3927 539 3985 573
rect 4019 539 4077 573
rect 4111 539 4169 573
rect 4203 539 4261 573
rect 4295 539 4353 573
rect 4387 539 4445 573
rect 4479 539 4537 573
rect 4571 539 4629 573
rect 4663 539 4721 573
rect 4755 539 4813 573
rect 4847 539 4905 573
rect 4939 539 4997 573
rect 5031 539 5089 573
rect 5123 539 5181 573
rect 5215 539 5273 573
rect 5307 539 5365 573
rect 5399 539 5457 573
rect 5491 539 5549 573
rect 5583 539 5641 573
rect 5675 539 5733 573
rect 5767 539 5825 573
rect 5859 539 5917 573
rect 5951 539 6009 573
rect 6043 539 6101 573
rect 6135 539 6193 573
rect 6227 539 6285 573
rect 6319 539 6377 573
rect 6411 539 6469 573
rect 6503 539 6561 573
rect 6595 539 6653 573
rect 6687 539 6745 573
rect 6779 539 6837 573
rect 6871 539 6929 573
rect 6963 539 7021 573
rect 7055 539 7113 573
rect 7147 539 7205 573
rect 7239 539 7297 573
rect 7331 539 7389 573
rect 7423 539 7481 573
rect 7515 539 7573 573
rect 7607 539 7665 573
rect 7699 539 7757 573
rect 7791 539 7849 573
rect 7883 539 7941 573
rect 7975 539 8033 573
rect 8067 539 8125 573
rect 8159 539 8217 573
rect 8251 539 8309 573
rect 8343 539 8401 573
rect 8435 539 8493 573
rect 8527 539 8585 573
rect 8619 539 8677 573
rect 8711 539 8769 573
rect 8803 539 8861 573
rect 8895 539 8953 573
rect 8987 539 9045 573
rect 9079 539 9137 573
rect 9171 539 9229 573
rect 9263 539 9321 573
rect 9355 539 9413 573
rect 9447 539 9505 573
rect 9539 539 9597 573
rect 9631 539 9689 573
rect 9723 539 9781 573
rect 9815 539 9873 573
rect 9907 539 9965 573
rect 9999 539 10057 573
rect 10091 539 10149 573
rect 10183 539 10241 573
rect 10275 539 10333 573
rect 10367 539 10425 573
rect 10459 539 10517 573
rect 10551 539 10609 573
rect 10643 539 10701 573
rect 10735 539 10793 573
rect 10827 539 10885 573
rect 10919 539 10977 573
rect 11011 539 11069 573
rect 11103 539 11161 573
rect 11195 539 11253 573
rect 11287 539 11345 573
rect 11379 539 11437 573
rect 11471 539 11529 573
rect 11563 539 11621 573
rect 11655 539 11713 573
rect 11747 539 11805 573
rect 11839 539 11897 573
rect 11931 539 11989 573
rect 12023 539 12081 573
rect 12115 539 12173 573
rect 12207 539 12265 573
rect 12299 539 12357 573
rect 12391 539 12449 573
rect 12483 539 12541 573
rect 12575 539 12633 573
rect 12667 539 12725 573
rect 12759 539 12817 573
rect 12851 539 12909 573
rect 12943 539 13001 573
rect 13035 539 13093 573
rect 13127 539 13185 573
rect 13219 539 13277 573
rect 13311 539 13369 573
rect 13403 539 13461 573
rect 13495 539 13553 573
rect 13587 539 13645 573
rect 13679 539 13737 573
rect 13771 539 13829 573
rect 13863 539 13921 573
rect 13955 539 14013 573
rect 14047 539 14105 573
rect 14139 539 14197 573
rect 14231 539 14289 573
rect 14323 539 14381 573
rect 14415 539 14473 573
rect 14507 539 14565 573
rect 14599 539 14657 573
rect 14691 539 14749 573
rect 14783 539 14841 573
rect 14875 539 14933 573
rect 14967 539 15025 573
rect 15059 539 15117 573
rect 15151 539 15209 573
rect 15243 539 15301 573
rect 15335 539 15393 573
rect 15427 539 15485 573
rect 15519 539 15577 573
rect 15611 539 15669 573
rect 15703 539 15761 573
rect 15795 539 15853 573
rect 15887 539 15945 573
rect 15979 539 16037 573
rect 16071 539 16129 573
rect 16163 539 16221 573
rect 16255 539 16313 573
rect 16347 539 16405 573
rect 16439 539 16497 573
rect 16531 539 16589 573
rect 16623 539 16681 573
rect 16715 539 16744 573
rect 0 -150 29 -116
rect 63 -150 121 -116
rect 155 -150 213 -116
rect 247 -150 305 -116
rect 339 -150 397 -116
rect 431 -150 489 -116
rect 523 -150 581 -116
rect 615 -150 673 -116
rect 707 -150 765 -116
rect 799 -150 857 -116
rect 891 -150 949 -116
rect 983 -150 1041 -116
rect 1075 -150 1133 -116
rect 1167 -150 1225 -116
rect 1259 -150 1317 -116
rect 1351 -150 1409 -116
rect 1443 -150 1501 -116
rect 1535 -150 1593 -116
rect 1627 -150 1685 -116
rect 1719 -150 1777 -116
rect 1811 -150 1869 -116
rect 1903 -150 1961 -116
rect 1995 -150 2053 -116
rect 2087 -150 2145 -116
rect 2179 -150 2237 -116
rect 2271 -150 2329 -116
rect 2363 -150 2421 -116
rect 2455 -150 2513 -116
rect 2547 -150 2605 -116
rect 2639 -150 2697 -116
rect 2731 -150 2789 -116
rect 2823 -150 2881 -116
rect 2915 -150 2973 -116
rect 3007 -150 3065 -116
rect 3099 -150 3157 -116
rect 3191 -150 3249 -116
rect 3283 -150 3341 -116
rect 3375 -150 3433 -116
rect 3467 -150 3525 -116
rect 3559 -150 3617 -116
rect 3651 -150 3709 -116
rect 3743 -150 3801 -116
rect 3835 -150 3893 -116
rect 3927 -150 3985 -116
rect 4019 -150 4077 -116
rect 4111 -150 4169 -116
rect 4203 -150 4261 -116
rect 4295 -150 4353 -116
rect 4387 -150 4445 -116
rect 4479 -150 4537 -116
rect 4571 -150 4629 -116
rect 4663 -150 4721 -116
rect 4755 -150 4813 -116
rect 4847 -150 4905 -116
rect 4939 -150 4997 -116
rect 5031 -150 5089 -116
rect 5123 -150 5181 -116
rect 5215 -150 5273 -116
rect 5307 -150 5365 -116
rect 5399 -150 5457 -116
rect 5491 -150 5549 -116
rect 5583 -150 5641 -116
rect 5675 -150 5733 -116
rect 5767 -150 5825 -116
rect 5859 -150 5917 -116
rect 5951 -150 6009 -116
rect 6043 -150 6101 -116
rect 6135 -150 6193 -116
rect 6227 -150 6285 -116
rect 6319 -150 6377 -116
rect 6411 -150 6469 -116
rect 6503 -150 6561 -116
rect 6595 -150 6653 -116
rect 6687 -150 6745 -116
rect 6779 -150 6837 -116
rect 6871 -150 6929 -116
rect 6963 -150 7021 -116
rect 7055 -150 7113 -116
rect 7147 -150 7205 -116
rect 7239 -150 7297 -116
rect 7331 -150 7389 -116
rect 7423 -150 7481 -116
rect 7515 -150 7573 -116
rect 7607 -150 7665 -116
rect 7699 -150 7757 -116
rect 7791 -150 7849 -116
rect 7883 -150 7941 -116
rect 7975 -150 8033 -116
rect 8067 -150 8125 -116
rect 8159 -150 8217 -116
rect 8251 -150 8309 -116
rect 8343 -150 8401 -116
rect 8435 -150 8493 -116
rect 8527 -150 8585 -116
rect 8619 -150 8677 -116
rect 8711 -150 8769 -116
rect 8803 -150 8861 -116
rect 8895 -150 8953 -116
rect 8987 -150 9045 -116
rect 9079 -150 9137 -116
rect 9171 -150 9229 -116
rect 9263 -150 9321 -116
rect 9355 -150 9413 -116
rect 9447 -150 9505 -116
rect 9539 -150 9597 -116
rect 9631 -150 9689 -116
rect 9723 -150 9781 -116
rect 9815 -150 9873 -116
rect 9907 -150 9965 -116
rect 9999 -150 10057 -116
rect 10091 -150 10149 -116
rect 10183 -150 10241 -116
rect 10275 -150 10333 -116
rect 10367 -150 10425 -116
rect 10459 -150 10517 -116
rect 10551 -150 10609 -116
rect 10643 -150 10701 -116
rect 10735 -150 10793 -116
rect 10827 -150 10885 -116
rect 10919 -150 10977 -116
rect 11011 -150 11069 -116
rect 11103 -150 11161 -116
rect 11195 -150 11253 -116
rect 11287 -150 11345 -116
rect 11379 -150 11437 -116
rect 11471 -150 11529 -116
rect 11563 -150 11621 -116
rect 11655 -150 11713 -116
rect 11747 -150 11805 -116
rect 11839 -150 11897 -116
rect 11931 -150 11989 -116
rect 12023 -150 12081 -116
rect 12115 -150 12173 -116
rect 12207 -150 12265 -116
rect 12299 -150 12357 -116
rect 12391 -150 12449 -116
rect 12483 -150 12541 -116
rect 12575 -150 12633 -116
rect 12667 -150 12725 -116
rect 12759 -150 12817 -116
rect 12851 -150 12909 -116
rect 12943 -150 13001 -116
rect 13035 -150 13093 -116
rect 13127 -150 13185 -116
rect 13219 -150 13277 -116
rect 13311 -150 13369 -116
rect 13403 -150 13461 -116
rect 13495 -150 13553 -116
rect 13587 -150 13645 -116
rect 13679 -150 13737 -116
rect 13771 -150 13829 -116
rect 13863 -150 13921 -116
rect 13955 -150 14013 -116
rect 14047 -150 14105 -116
rect 14139 -150 14197 -116
rect 14231 -150 14289 -116
rect 14323 -150 14381 -116
rect 14415 -150 14473 -116
rect 14507 -150 14565 -116
rect 14599 -150 14657 -116
rect 14691 -150 14749 -116
rect 14783 -150 14841 -116
rect 14875 -150 14933 -116
rect 14967 -150 15025 -116
rect 15059 -150 15117 -116
rect 15151 -150 15209 -116
rect 15243 -150 15301 -116
rect 15335 -150 15393 -116
rect 15427 -150 15485 -116
rect 15519 -150 15577 -116
rect 15611 -150 15669 -116
rect 15703 -150 15761 -116
rect 15795 -150 15853 -116
rect 15887 -150 15945 -116
rect 15979 -150 16037 -116
rect 16071 -150 16129 -116
rect 16163 -150 16221 -116
rect 16255 -150 16313 -116
rect 16347 -150 16405 -116
rect 16439 -150 16497 -116
rect 16531 -150 16589 -116
rect 16623 -150 16681 -116
rect 16715 -150 16744 -116
<< nsubdiff >>
rect 2 2961 31 2995
rect 65 2961 123 2995
rect 157 2961 215 2995
rect 249 2961 307 2995
rect 341 2961 399 2995
rect 433 2961 491 2995
rect 525 2961 583 2995
rect 617 2961 675 2995
rect 709 2961 767 2995
rect 801 2961 859 2995
rect 893 2961 951 2995
rect 985 2961 1043 2995
rect 1077 2961 1135 2995
rect 1169 2961 1227 2995
rect 1261 2961 1319 2995
rect 1353 2961 1411 2995
rect 1445 2961 1503 2995
rect 1537 2961 1595 2995
rect 1629 2961 1687 2995
rect 1721 2961 1779 2995
rect 1813 2961 1871 2995
rect 1905 2961 1963 2995
rect 1997 2961 2055 2995
rect 2089 2961 2147 2995
rect 2181 2961 2239 2995
rect 2273 2961 2331 2995
rect 2365 2961 2423 2995
rect 2457 2961 2515 2995
rect 2549 2961 2607 2995
rect 2641 2961 2699 2995
rect 2733 2961 2791 2995
rect 2825 2961 2854 2995
rect 4386 2961 4415 2995
rect 4449 2961 4507 2995
rect 4541 2961 4599 2995
rect 4633 2961 4691 2995
rect 4725 2961 4783 2995
rect 4817 2961 4875 2995
rect 4909 2961 4967 2995
rect 5001 2961 5059 2995
rect 5093 2961 5151 2995
rect 5185 2961 5243 2995
rect 5277 2961 5335 2995
rect 5369 2961 5427 2995
rect 5461 2961 5519 2995
rect 5553 2961 5611 2995
rect 5645 2961 5703 2995
rect 5737 2961 5795 2995
rect 5829 2961 5887 2995
rect 5921 2961 5979 2995
rect 6013 2961 6071 2995
rect 6105 2961 6163 2995
rect 6197 2961 6255 2995
rect 6289 2961 6347 2995
rect 6381 2961 6439 2995
rect 6473 2961 6531 2995
rect 6565 2961 6623 2995
rect 6657 2961 6715 2995
rect 6749 2961 6807 2995
rect 6841 2961 6899 2995
rect 6933 2961 6991 2995
rect 7025 2961 7083 2995
rect 7117 2961 7175 2995
rect 7209 2961 7238 2995
rect 0 1819 29 1853
rect 63 1819 121 1853
rect 155 1819 213 1853
rect 247 1819 305 1853
rect 339 1819 397 1853
rect 431 1819 489 1853
rect 523 1819 581 1853
rect 615 1819 673 1853
rect 707 1819 765 1853
rect 799 1819 857 1853
rect 891 1819 949 1853
rect 983 1819 1041 1853
rect 1075 1819 1133 1853
rect 1167 1819 1225 1853
rect 1259 1819 1317 1853
rect 1351 1819 1409 1853
rect 1443 1819 1501 1853
rect 1535 1819 1593 1853
rect 1627 1819 1685 1853
rect 1719 1819 1777 1853
rect 1811 1819 1869 1853
rect 1903 1819 1961 1853
rect 1995 1819 2053 1853
rect 2087 1819 2145 1853
rect 2179 1819 2237 1853
rect 2271 1819 2329 1853
rect 2363 1819 2421 1853
rect 2455 1819 2513 1853
rect 2547 1819 2605 1853
rect 2639 1819 2697 1853
rect 2731 1819 2789 1853
rect 2823 1819 2881 1853
rect 2915 1819 2973 1853
rect 3007 1819 3065 1853
rect 3099 1819 3157 1853
rect 3191 1819 3249 1853
rect 3283 1819 3341 1853
rect 3375 1819 3433 1853
rect 3467 1819 3525 1853
rect 3559 1819 3617 1853
rect 3651 1819 3709 1853
rect 3743 1819 3801 1853
rect 3835 1819 3893 1853
rect 3927 1819 3985 1853
rect 4019 1819 4077 1853
rect 4111 1819 4169 1853
rect 4203 1819 4261 1853
rect 4295 1819 4353 1853
rect 4387 1819 4445 1853
rect 4479 1819 4537 1853
rect 4571 1819 4629 1853
rect 4663 1819 4721 1853
rect 4755 1819 4813 1853
rect 4847 1819 4905 1853
rect 4939 1819 4997 1853
rect 5031 1819 5089 1853
rect 5123 1819 5181 1853
rect 5215 1819 5273 1853
rect 5307 1819 5365 1853
rect 5399 1819 5457 1853
rect 5491 1819 5549 1853
rect 5583 1819 5641 1853
rect 5675 1849 5704 1853
rect 6216 1849 6245 1853
rect 5675 1819 6245 1849
rect 6279 1819 6337 1853
rect 6371 1819 6429 1853
rect 6463 1819 6521 1853
rect 6555 1819 6613 1853
rect 6647 1819 6705 1853
rect 6739 1819 6797 1853
rect 6831 1819 6889 1853
rect 6923 1819 6981 1853
rect 7015 1819 7073 1853
rect 7107 1819 7165 1853
rect 7199 1819 7257 1853
rect 7291 1819 7349 1853
rect 7383 1819 7441 1853
rect 7475 1819 7533 1853
rect 7567 1819 7625 1853
rect 7659 1819 7717 1853
rect 7751 1819 7809 1853
rect 7843 1819 7901 1853
rect 7935 1819 7993 1853
rect 8027 1819 8085 1853
rect 8119 1819 8177 1853
rect 8211 1819 8269 1853
rect 8303 1819 8361 1853
rect 8395 1819 8453 1853
rect 8487 1819 8545 1853
rect 8579 1819 8637 1853
rect 8671 1819 8729 1853
rect 8763 1819 8821 1853
rect 8855 1819 8913 1853
rect 8947 1819 9005 1853
rect 9039 1819 9097 1853
rect 9131 1819 9189 1853
rect 9223 1819 9281 1853
rect 9315 1819 9373 1853
rect 9407 1819 9465 1853
rect 9499 1819 9557 1853
rect 9591 1819 9649 1853
rect 9683 1819 9741 1853
rect 9775 1819 9833 1853
rect 9867 1819 9925 1853
rect 9959 1819 10017 1853
rect 10051 1819 10109 1853
rect 10143 1819 10201 1853
rect 10235 1819 10293 1853
rect 10327 1819 10385 1853
rect 10419 1819 10477 1853
rect 10511 1819 10569 1853
rect 10603 1819 10661 1853
rect 10695 1819 10753 1853
rect 10787 1819 10845 1853
rect 10879 1819 10937 1853
rect 10971 1819 11029 1853
rect 11063 1819 11121 1853
rect 11155 1819 11213 1853
rect 11247 1819 11305 1853
rect 11339 1819 11397 1853
rect 11431 1819 11489 1853
rect 11523 1819 11581 1853
rect 11615 1819 11673 1853
rect 11707 1819 11765 1853
rect 11799 1819 11857 1853
rect 11891 1849 11920 1853
rect 11982 1849 12011 1853
rect 11891 1819 12011 1849
rect 12045 1819 12103 1853
rect 12137 1819 12195 1853
rect 12229 1819 12287 1853
rect 12321 1819 12379 1853
rect 12413 1819 12471 1853
rect 12505 1819 12563 1853
rect 12597 1819 12655 1853
rect 12689 1819 12747 1853
rect 12781 1819 12839 1853
rect 12873 1819 12931 1853
rect 12965 1819 13023 1853
rect 13057 1819 13115 1853
rect 13149 1819 13207 1853
rect 13241 1819 13299 1853
rect 13333 1819 13391 1853
rect 13425 1819 13483 1853
rect 13517 1819 13575 1853
rect 13609 1819 13667 1853
rect 13701 1819 13759 1853
rect 13793 1819 13851 1853
rect 13885 1819 13943 1853
rect 13977 1819 14035 1853
rect 14069 1819 14127 1853
rect 14161 1819 14219 1853
rect 14253 1819 14311 1853
rect 14345 1819 14403 1853
rect 14437 1819 14495 1853
rect 14529 1819 14587 1853
rect 14621 1819 14679 1853
rect 14713 1819 14771 1853
rect 14805 1819 14863 1853
rect 14897 1819 14955 1853
rect 14989 1819 15047 1853
rect 15081 1819 15139 1853
rect 15173 1819 15231 1853
rect 15265 1819 15323 1853
rect 15357 1819 15415 1853
rect 15449 1819 15507 1853
rect 15541 1819 15599 1853
rect 15633 1819 15691 1853
rect 15725 1819 15783 1853
rect 15817 1819 15875 1853
rect 15909 1819 15967 1853
rect 16001 1819 16059 1853
rect 16093 1819 16151 1853
rect 16185 1819 16243 1853
rect 16277 1819 16335 1853
rect 16369 1819 16427 1853
rect 16461 1819 16519 1853
rect 16553 1849 16582 1853
rect 16553 1819 16614 1849
rect 3704 1804 3757 1819
rect 1 1161 29 1165
rect -1 1131 29 1161
rect 63 1131 121 1165
rect 155 1131 213 1165
rect 247 1131 305 1165
rect 339 1131 397 1165
rect 431 1131 489 1165
rect 523 1131 581 1165
rect 615 1131 673 1165
rect 707 1131 765 1165
rect 799 1131 857 1165
rect 891 1131 949 1165
rect 983 1131 1041 1165
rect 1075 1131 1133 1165
rect 1167 1131 1225 1165
rect 1259 1131 1317 1165
rect 1351 1131 1409 1165
rect 1443 1131 1501 1165
rect 1535 1131 1593 1165
rect 1627 1131 1685 1165
rect 1719 1131 1777 1165
rect 1811 1161 1835 1165
rect 1811 1131 1843 1161
rect 2029 1161 2053 1165
rect 1995 1131 2053 1161
rect 2087 1131 2145 1165
rect 2179 1131 2237 1165
rect 2271 1131 2329 1165
rect 2363 1131 2421 1165
rect 2455 1131 2513 1165
rect 2547 1131 2605 1165
rect 2639 1131 2697 1165
rect 2731 1131 2789 1165
rect 2823 1131 2881 1165
rect 2915 1131 2973 1165
rect 3007 1131 3065 1165
rect 3099 1131 3157 1165
rect 3191 1131 3249 1165
rect 3283 1131 3341 1165
rect 3375 1131 3433 1165
rect 3467 1131 3525 1165
rect 3559 1131 3617 1165
rect 3651 1131 3709 1165
rect 3743 1131 3801 1165
rect 3835 1131 3893 1165
rect 3927 1131 3985 1165
rect 4019 1131 4077 1165
rect 4111 1131 4169 1165
rect 4203 1161 4227 1165
rect 4203 1131 4254 1161
rect 4421 1161 4445 1165
rect 4387 1131 4445 1161
rect 4479 1131 4537 1165
rect 4571 1131 4629 1165
rect 4663 1131 4721 1165
rect 4755 1131 4813 1165
rect 4847 1131 4905 1165
rect 4939 1131 4997 1165
rect 5031 1131 5089 1165
rect 5123 1131 5181 1165
rect 5215 1131 5273 1165
rect 5307 1131 5365 1165
rect 5399 1131 5457 1165
rect 5491 1131 5549 1165
rect 5583 1131 5641 1165
rect 5675 1131 5733 1165
rect 5767 1131 5825 1165
rect 5859 1131 5917 1165
rect 5951 1131 6009 1165
rect 6043 1131 6101 1165
rect 6135 1131 6193 1165
rect 6227 1131 6285 1165
rect 6319 1131 6377 1165
rect 6411 1131 6469 1165
rect 6503 1131 6561 1165
rect 6595 1161 6619 1165
rect 6595 1131 6643 1161
rect 6813 1161 6837 1165
rect 6779 1131 6837 1161
rect 6871 1131 6929 1165
rect 6963 1131 7021 1165
rect 7055 1131 7113 1165
rect 7147 1131 7205 1165
rect 7239 1131 7297 1165
rect 7331 1131 7389 1165
rect 7423 1131 7481 1165
rect 7515 1131 7573 1165
rect 7607 1131 7665 1165
rect 7699 1131 7757 1165
rect 7791 1131 7849 1165
rect 7883 1131 7941 1165
rect 7975 1131 8033 1165
rect 8067 1131 8125 1165
rect 8159 1131 8217 1165
rect 8251 1131 8309 1165
rect 8343 1131 8401 1165
rect 8435 1131 8493 1165
rect 8527 1131 8585 1165
rect 8619 1131 8677 1165
rect 8711 1131 8769 1165
rect 8803 1131 8861 1165
rect 8895 1131 8953 1165
rect 8987 1161 9011 1165
rect 8987 1131 9037 1161
rect 9205 1161 9229 1165
rect 9171 1131 9229 1161
rect 9263 1131 9321 1165
rect 9355 1131 9413 1165
rect 9447 1131 9505 1165
rect 9539 1131 9597 1165
rect 9631 1131 9689 1165
rect 9723 1131 9781 1165
rect 9815 1131 9873 1165
rect 9907 1131 9965 1165
rect 9999 1131 10057 1165
rect 10091 1131 10149 1165
rect 10183 1131 10241 1165
rect 10275 1131 10333 1165
rect 10367 1131 10425 1165
rect 10459 1131 10517 1165
rect 10551 1131 10609 1165
rect 10643 1131 10701 1165
rect 10735 1131 10793 1165
rect 10827 1131 10885 1165
rect 10919 1131 10977 1165
rect 11011 1131 11069 1165
rect 11103 1131 11161 1165
rect 11195 1131 11253 1165
rect 11287 1131 11345 1165
rect 11379 1161 11403 1165
rect 11379 1131 11427 1161
rect 11597 1161 11621 1165
rect 11563 1131 11621 1161
rect 11655 1131 11713 1165
rect 11747 1131 11805 1165
rect 11839 1131 11897 1165
rect 11931 1131 11989 1165
rect 12023 1131 12081 1165
rect 12115 1131 12173 1165
rect 12207 1131 12265 1165
rect 12299 1131 12357 1165
rect 12391 1131 12449 1165
rect 12483 1131 12541 1165
rect 12575 1131 12633 1165
rect 12667 1131 12725 1165
rect 12759 1131 12817 1165
rect 12851 1131 12909 1165
rect 12943 1131 13001 1165
rect 13035 1131 13093 1165
rect 13127 1131 13185 1165
rect 13219 1131 13277 1165
rect 13311 1131 13369 1165
rect 13403 1131 13461 1165
rect 13495 1131 13553 1165
rect 13587 1131 13645 1165
rect 13679 1131 13737 1165
rect 13771 1161 13795 1165
rect 13771 1131 13819 1161
rect 13989 1161 14013 1165
rect 13955 1131 14013 1161
rect 14047 1131 14105 1165
rect 14139 1131 14197 1165
rect 14231 1131 14289 1165
rect 14323 1131 14381 1165
rect 14415 1131 14473 1165
rect 14507 1131 14565 1165
rect 14599 1131 14657 1165
rect 14691 1131 14749 1165
rect 14783 1131 14841 1165
rect 14875 1131 14933 1165
rect 14967 1131 15025 1165
rect 15059 1131 15117 1165
rect 15151 1131 15209 1165
rect 15243 1131 15301 1165
rect 15335 1131 15393 1165
rect 15427 1131 15485 1165
rect 15519 1131 15577 1165
rect 15611 1131 15669 1165
rect 15703 1131 15761 1165
rect 15795 1131 15853 1165
rect 15887 1131 15945 1165
rect 15979 1131 16037 1165
rect 16071 1131 16129 1165
rect 16163 1161 16187 1165
rect 16163 1131 16211 1161
rect 16381 1161 16405 1165
rect 16347 1131 16405 1161
rect 16439 1131 16497 1165
rect 16531 1131 16589 1165
rect 16623 1131 16681 1165
rect 16715 1131 16744 1165
rect 0 476 571 477
rect 0 442 29 476
rect 63 442 121 476
rect 155 442 213 476
rect 247 442 305 476
rect 339 442 394 476
rect 428 442 496 476
rect 530 442 581 476
rect 615 442 673 476
rect 707 442 765 476
rect 799 442 857 476
rect 891 442 949 476
rect 983 442 1041 476
rect 1075 442 1133 476
rect 1167 442 1225 476
rect 1259 442 1317 476
rect 1351 442 1409 476
rect 1443 442 1501 476
rect 1535 442 1559 476
rect 1753 442 1777 476
rect 1811 442 1869 476
rect 1903 442 1961 476
rect 1995 442 2053 476
rect 2087 442 2145 476
rect 2179 442 2237 476
rect 2271 442 2329 476
rect 2363 442 2421 476
rect 2455 442 2513 476
rect 2547 442 2605 476
rect 2639 442 2697 476
rect 2731 442 2791 476
rect 2825 442 2882 476
rect 2916 442 2973 476
rect 3007 442 3065 476
rect 3099 442 3157 476
rect 3191 442 3249 476
rect 3283 442 3341 476
rect 3375 442 3433 476
rect 3467 442 3525 476
rect 3559 442 3617 476
rect 3651 442 3709 476
rect 3743 442 3801 476
rect 3835 442 3893 476
rect 3927 442 3955 476
rect 4145 442 4169 476
rect 4203 442 4261 476
rect 4295 442 4353 476
rect 4387 442 4445 476
rect 4479 442 4537 476
rect 4571 442 4629 476
rect 4663 442 4721 476
rect 4755 442 4813 476
rect 4847 442 4905 476
rect 4939 442 4997 476
rect 5031 442 5089 476
rect 5123 442 5179 476
rect 5213 442 5273 476
rect 5307 442 5365 476
rect 5399 442 5457 476
rect 5491 442 5549 476
rect 5583 442 5641 476
rect 5675 442 5733 476
rect 5767 442 5825 476
rect 5859 442 5917 476
rect 5951 442 6009 476
rect 6043 442 6101 476
rect 6135 442 6193 476
rect 6227 442 6285 476
rect 6319 442 6353 476
rect 6518 442 6561 476
rect 6595 442 6653 476
rect 6687 442 6745 476
rect 6779 442 6837 476
rect 6871 442 6929 476
rect 6963 442 7021 476
rect 7055 442 7113 476
rect 7147 442 7205 476
rect 7239 442 7297 476
rect 7331 442 7389 476
rect 7423 442 7481 476
rect 7515 442 7574 476
rect 7608 442 7665 476
rect 7699 442 7757 476
rect 7791 442 7849 476
rect 7883 442 7941 476
rect 7975 442 8033 476
rect 8067 442 8125 476
rect 8159 442 8217 476
rect 8251 442 8309 476
rect 8343 442 8401 476
rect 8435 442 8493 476
rect 8527 442 8585 476
rect 8619 442 8677 476
rect 8711 442 8745 476
rect 8929 442 8953 476
rect 8987 442 9045 476
rect 9079 442 9137 476
rect 9171 442 9229 476
rect 9263 442 9321 476
rect 9355 442 9413 476
rect 9447 442 9505 476
rect 9539 442 9597 476
rect 9631 442 9689 476
rect 9723 442 9781 476
rect 9815 442 9873 476
rect 9907 442 9963 476
rect 9997 442 10058 476
rect 10092 442 10149 476
rect 10183 442 10241 476
rect 10275 442 10333 476
rect 10367 442 10425 476
rect 10459 442 10517 476
rect 10551 442 10609 476
rect 10643 442 10701 476
rect 10735 442 10793 476
rect 10827 442 10885 476
rect 10919 442 10977 476
rect 11011 442 11069 476
rect 11103 442 11127 476
rect 11315 442 11345 476
rect 11379 442 11437 476
rect 11471 442 11529 476
rect 11563 442 11621 476
rect 11655 442 11713 476
rect 11747 442 11805 476
rect 11839 442 11897 476
rect 11931 442 11989 476
rect 12023 442 12081 476
rect 12115 442 12173 476
rect 12207 442 12265 476
rect 12299 442 12357 476
rect 12391 442 12448 476
rect 12482 442 12541 476
rect 12575 442 12633 476
rect 12667 442 12725 476
rect 12759 442 12817 476
rect 12851 442 12909 476
rect 12943 442 13001 476
rect 13035 442 13093 476
rect 13127 442 13185 476
rect 13219 442 13277 476
rect 13311 442 13369 476
rect 13403 442 13461 476
rect 13495 442 13519 476
rect 13639 442 13737 476
rect 13771 442 13829 476
rect 13863 442 13921 476
rect 13955 442 14013 476
rect 14047 442 14105 476
rect 14139 442 14197 476
rect 14231 442 14289 476
rect 14323 442 14381 476
rect 14415 442 14473 476
rect 14507 442 14565 476
rect 14599 442 14657 476
rect 14691 442 14748 476
rect 14782 442 14842 476
rect 14876 442 14933 476
rect 14967 442 15025 476
rect 15059 442 15117 476
rect 15151 442 15209 476
rect 15243 442 15301 476
rect 15335 442 15393 476
rect 15427 442 15485 476
rect 15519 442 15577 476
rect 15611 442 15669 476
rect 15703 442 15761 476
rect 15795 442 15853 476
rect 15887 442 15921 476
rect 16031 442 16129 476
rect 16163 442 16221 476
rect 16255 442 16313 476
rect 16347 442 16405 476
rect 16439 442 16497 476
rect 16531 442 16589 476
rect 16623 442 16681 476
rect 16715 442 16744 476
<< psubdiffcont >>
rect 31 2369 65 2403
rect 123 2369 157 2403
rect 215 2369 249 2403
rect 307 2369 341 2403
rect 399 2369 433 2403
rect 491 2369 525 2403
rect 583 2369 617 2403
rect 675 2369 709 2403
rect 767 2369 801 2403
rect 859 2369 893 2403
rect 951 2369 985 2403
rect 1043 2369 1077 2403
rect 1135 2369 1169 2403
rect 1227 2369 1261 2403
rect 1319 2369 1353 2403
rect 1411 2369 1445 2403
rect 1503 2369 1537 2403
rect 1595 2369 1629 2403
rect 1687 2369 1721 2403
rect 1779 2369 1813 2403
rect 1871 2369 1905 2403
rect 1963 2369 1997 2403
rect 2055 2369 2089 2403
rect 2147 2369 2181 2403
rect 2239 2369 2273 2403
rect 2331 2369 2365 2403
rect 2423 2369 2457 2403
rect 2515 2369 2549 2403
rect 2607 2369 2641 2403
rect 2699 2369 2733 2403
rect 2791 2369 2825 2403
rect 4415 2369 4449 2403
rect 4507 2369 4541 2403
rect 4599 2369 4633 2403
rect 4691 2369 4725 2403
rect 4783 2369 4817 2403
rect 4875 2369 4909 2403
rect 4967 2369 5001 2403
rect 5059 2369 5093 2403
rect 5151 2369 5185 2403
rect 5243 2369 5277 2403
rect 5335 2369 5369 2403
rect 5427 2369 5461 2403
rect 5519 2369 5553 2403
rect 5611 2369 5645 2403
rect 5703 2369 5737 2403
rect 5795 2369 5829 2403
rect 5887 2369 5921 2403
rect 5979 2369 6013 2403
rect 6071 2369 6105 2403
rect 6163 2369 6197 2403
rect 6255 2369 6289 2403
rect 6347 2369 6381 2403
rect 6439 2369 6473 2403
rect 6531 2369 6565 2403
rect 6623 2369 6657 2403
rect 6715 2369 6749 2403
rect 6807 2369 6841 2403
rect 6899 2369 6933 2403
rect 6991 2369 7025 2403
rect 7083 2369 7117 2403
rect 7175 2369 7209 2403
rect 29 1227 63 1261
rect 121 1227 155 1261
rect 213 1227 247 1261
rect 305 1227 339 1261
rect 397 1227 431 1261
rect 489 1227 523 1261
rect 581 1227 615 1261
rect 673 1227 707 1261
rect 765 1227 799 1261
rect 857 1227 891 1261
rect 949 1227 983 1261
rect 1041 1227 1075 1261
rect 1133 1227 1167 1261
rect 1225 1227 1259 1261
rect 1317 1227 1351 1261
rect 1409 1227 1443 1261
rect 1501 1227 1535 1261
rect 1593 1227 1627 1261
rect 1685 1227 1719 1261
rect 1777 1227 1811 1261
rect 1869 1227 1903 1261
rect 1961 1227 1995 1261
rect 2053 1227 2087 1261
rect 2145 1227 2179 1261
rect 2237 1227 2271 1261
rect 2329 1227 2363 1261
rect 2421 1227 2455 1261
rect 2513 1227 2547 1261
rect 2605 1227 2639 1261
rect 2697 1227 2731 1261
rect 2789 1227 2823 1261
rect 2881 1227 2915 1261
rect 2973 1227 3007 1261
rect 3065 1227 3099 1261
rect 3157 1227 3191 1261
rect 3249 1227 3283 1261
rect 3341 1227 3375 1261
rect 3433 1227 3467 1261
rect 3525 1227 3559 1261
rect 3617 1227 3651 1261
rect 3709 1227 3743 1261
rect 3801 1227 3835 1261
rect 3893 1227 3927 1261
rect 3985 1227 4019 1261
rect 4077 1227 4111 1261
rect 4169 1227 4203 1261
rect 4261 1227 4295 1261
rect 4353 1227 4387 1261
rect 4445 1227 4479 1261
rect 4537 1227 4571 1261
rect 4629 1227 4663 1261
rect 4721 1227 4755 1261
rect 4813 1227 4847 1261
rect 4905 1227 4939 1261
rect 4997 1227 5031 1261
rect 5089 1227 5123 1261
rect 5181 1227 5215 1261
rect 5273 1227 5307 1261
rect 5365 1227 5399 1261
rect 5457 1227 5491 1261
rect 5549 1227 5583 1261
rect 5641 1227 5675 1261
rect 6245 1227 6279 1261
rect 6337 1227 6371 1261
rect 6429 1227 6463 1261
rect 6521 1227 6555 1261
rect 6613 1227 6647 1261
rect 6705 1227 6739 1261
rect 6797 1227 6831 1261
rect 6889 1227 6923 1261
rect 6981 1227 7015 1261
rect 7073 1227 7107 1261
rect 7165 1227 7199 1261
rect 7257 1227 7291 1261
rect 7349 1227 7383 1261
rect 7441 1227 7475 1261
rect 7533 1227 7567 1261
rect 7625 1227 7659 1261
rect 7717 1227 7751 1261
rect 7809 1227 7843 1261
rect 7901 1227 7935 1261
rect 7993 1227 8027 1261
rect 8085 1227 8119 1261
rect 8177 1227 8211 1261
rect 8269 1227 8303 1261
rect 8361 1227 8395 1261
rect 8453 1227 8487 1261
rect 8545 1227 8579 1261
rect 8637 1227 8671 1261
rect 8729 1227 8763 1261
rect 8821 1227 8855 1261
rect 8913 1227 8947 1261
rect 9005 1227 9039 1261
rect 9097 1227 9131 1261
rect 9189 1227 9223 1261
rect 9281 1227 9315 1261
rect 9373 1227 9407 1261
rect 9465 1227 9499 1261
rect 9557 1227 9591 1261
rect 9649 1227 9683 1261
rect 9741 1227 9775 1261
rect 9833 1227 9867 1261
rect 9925 1227 9959 1261
rect 10017 1227 10051 1261
rect 10109 1227 10143 1261
rect 10201 1227 10235 1261
rect 10293 1227 10327 1261
rect 10385 1227 10419 1261
rect 10477 1227 10511 1261
rect 10569 1227 10603 1261
rect 10661 1227 10695 1261
rect 10753 1227 10787 1261
rect 10845 1227 10879 1261
rect 10937 1227 10971 1261
rect 11029 1227 11063 1261
rect 11121 1227 11155 1261
rect 11213 1227 11247 1261
rect 11305 1227 11339 1261
rect 11397 1227 11431 1261
rect 11489 1227 11523 1261
rect 11581 1227 11615 1261
rect 11673 1227 11707 1261
rect 11765 1227 11799 1261
rect 11857 1227 11891 1261
rect 12011 1227 12045 1261
rect 12103 1227 12137 1261
rect 12195 1227 12229 1261
rect 12287 1227 12321 1261
rect 12379 1227 12413 1261
rect 12471 1227 12505 1261
rect 12563 1227 12597 1261
rect 12655 1227 12689 1261
rect 12747 1227 12781 1261
rect 12839 1227 12873 1261
rect 12931 1227 12965 1261
rect 13023 1227 13057 1261
rect 13115 1227 13149 1261
rect 13207 1227 13241 1261
rect 13299 1227 13333 1261
rect 13391 1227 13425 1261
rect 13483 1227 13517 1261
rect 13575 1227 13609 1261
rect 13667 1227 13701 1261
rect 13759 1227 13793 1261
rect 13851 1227 13885 1261
rect 13943 1227 13977 1261
rect 14035 1227 14069 1261
rect 14127 1227 14161 1261
rect 14219 1227 14253 1261
rect 14311 1227 14345 1261
rect 14403 1227 14437 1261
rect 14495 1227 14529 1261
rect 14587 1227 14621 1261
rect 14679 1227 14713 1261
rect 14771 1227 14805 1261
rect 14863 1227 14897 1261
rect 14955 1227 14989 1261
rect 15047 1227 15081 1261
rect 15139 1227 15173 1261
rect 15231 1227 15265 1261
rect 15323 1227 15357 1261
rect 15415 1227 15449 1261
rect 15507 1227 15541 1261
rect 15599 1227 15633 1261
rect 15691 1227 15725 1261
rect 15783 1227 15817 1261
rect 15875 1227 15909 1261
rect 15967 1227 16001 1261
rect 16059 1227 16093 1261
rect 16151 1227 16185 1261
rect 16243 1227 16277 1261
rect 16335 1227 16369 1261
rect 16427 1227 16461 1261
rect 16519 1227 16553 1261
rect 29 539 63 573
rect 121 539 155 573
rect 213 539 247 573
rect 305 539 339 573
rect 397 539 431 573
rect 489 539 523 573
rect 581 539 615 573
rect 673 539 707 573
rect 765 539 799 573
rect 857 539 891 573
rect 949 539 983 573
rect 1041 539 1075 573
rect 1133 539 1167 573
rect 1225 539 1259 573
rect 1317 539 1351 573
rect 1409 539 1443 573
rect 1501 539 1535 573
rect 1593 539 1627 573
rect 1685 539 1719 573
rect 1777 539 1811 573
rect 1869 539 1903 573
rect 1961 539 1995 573
rect 2053 539 2087 573
rect 2145 539 2179 573
rect 2237 539 2271 573
rect 2329 539 2363 573
rect 2421 539 2455 573
rect 2513 539 2547 573
rect 2605 539 2639 573
rect 2697 539 2731 573
rect 2789 539 2823 573
rect 2881 539 2915 573
rect 2973 539 3007 573
rect 3065 539 3099 573
rect 3157 539 3191 573
rect 3249 539 3283 573
rect 3341 539 3375 573
rect 3433 539 3467 573
rect 3525 539 3559 573
rect 3617 539 3651 573
rect 3709 539 3743 573
rect 3801 539 3835 573
rect 3893 539 3927 573
rect 3985 539 4019 573
rect 4077 539 4111 573
rect 4169 539 4203 573
rect 4261 539 4295 573
rect 4353 539 4387 573
rect 4445 539 4479 573
rect 4537 539 4571 573
rect 4629 539 4663 573
rect 4721 539 4755 573
rect 4813 539 4847 573
rect 4905 539 4939 573
rect 4997 539 5031 573
rect 5089 539 5123 573
rect 5181 539 5215 573
rect 5273 539 5307 573
rect 5365 539 5399 573
rect 5457 539 5491 573
rect 5549 539 5583 573
rect 5641 539 5675 573
rect 5733 539 5767 573
rect 5825 539 5859 573
rect 5917 539 5951 573
rect 6009 539 6043 573
rect 6101 539 6135 573
rect 6193 539 6227 573
rect 6285 539 6319 573
rect 6377 539 6411 573
rect 6469 539 6503 573
rect 6561 539 6595 573
rect 6653 539 6687 573
rect 6745 539 6779 573
rect 6837 539 6871 573
rect 6929 539 6963 573
rect 7021 539 7055 573
rect 7113 539 7147 573
rect 7205 539 7239 573
rect 7297 539 7331 573
rect 7389 539 7423 573
rect 7481 539 7515 573
rect 7573 539 7607 573
rect 7665 539 7699 573
rect 7757 539 7791 573
rect 7849 539 7883 573
rect 7941 539 7975 573
rect 8033 539 8067 573
rect 8125 539 8159 573
rect 8217 539 8251 573
rect 8309 539 8343 573
rect 8401 539 8435 573
rect 8493 539 8527 573
rect 8585 539 8619 573
rect 8677 539 8711 573
rect 8769 539 8803 573
rect 8861 539 8895 573
rect 8953 539 8987 573
rect 9045 539 9079 573
rect 9137 539 9171 573
rect 9229 539 9263 573
rect 9321 539 9355 573
rect 9413 539 9447 573
rect 9505 539 9539 573
rect 9597 539 9631 573
rect 9689 539 9723 573
rect 9781 539 9815 573
rect 9873 539 9907 573
rect 9965 539 9999 573
rect 10057 539 10091 573
rect 10149 539 10183 573
rect 10241 539 10275 573
rect 10333 539 10367 573
rect 10425 539 10459 573
rect 10517 539 10551 573
rect 10609 539 10643 573
rect 10701 539 10735 573
rect 10793 539 10827 573
rect 10885 539 10919 573
rect 10977 539 11011 573
rect 11069 539 11103 573
rect 11161 539 11195 573
rect 11253 539 11287 573
rect 11345 539 11379 573
rect 11437 539 11471 573
rect 11529 539 11563 573
rect 11621 539 11655 573
rect 11713 539 11747 573
rect 11805 539 11839 573
rect 11897 539 11931 573
rect 11989 539 12023 573
rect 12081 539 12115 573
rect 12173 539 12207 573
rect 12265 539 12299 573
rect 12357 539 12391 573
rect 12449 539 12483 573
rect 12541 539 12575 573
rect 12633 539 12667 573
rect 12725 539 12759 573
rect 12817 539 12851 573
rect 12909 539 12943 573
rect 13001 539 13035 573
rect 13093 539 13127 573
rect 13185 539 13219 573
rect 13277 539 13311 573
rect 13369 539 13403 573
rect 13461 539 13495 573
rect 13553 539 13587 573
rect 13645 539 13679 573
rect 13737 539 13771 573
rect 13829 539 13863 573
rect 13921 539 13955 573
rect 14013 539 14047 573
rect 14105 539 14139 573
rect 14197 539 14231 573
rect 14289 539 14323 573
rect 14381 539 14415 573
rect 14473 539 14507 573
rect 14565 539 14599 573
rect 14657 539 14691 573
rect 14749 539 14783 573
rect 14841 539 14875 573
rect 14933 539 14967 573
rect 15025 539 15059 573
rect 15117 539 15151 573
rect 15209 539 15243 573
rect 15301 539 15335 573
rect 15393 539 15427 573
rect 15485 539 15519 573
rect 15577 539 15611 573
rect 15669 539 15703 573
rect 15761 539 15795 573
rect 15853 539 15887 573
rect 15945 539 15979 573
rect 16037 539 16071 573
rect 16129 539 16163 573
rect 16221 539 16255 573
rect 16313 539 16347 573
rect 16405 539 16439 573
rect 16497 539 16531 573
rect 16589 539 16623 573
rect 16681 539 16715 573
rect 29 -150 63 -116
rect 121 -150 155 -116
rect 213 -150 247 -116
rect 305 -150 339 -116
rect 397 -150 431 -116
rect 489 -150 523 -116
rect 581 -150 615 -116
rect 673 -150 707 -116
rect 765 -150 799 -116
rect 857 -150 891 -116
rect 949 -150 983 -116
rect 1041 -150 1075 -116
rect 1133 -150 1167 -116
rect 1225 -150 1259 -116
rect 1317 -150 1351 -116
rect 1409 -150 1443 -116
rect 1501 -150 1535 -116
rect 1593 -150 1627 -116
rect 1685 -150 1719 -116
rect 1777 -150 1811 -116
rect 1869 -150 1903 -116
rect 1961 -150 1995 -116
rect 2053 -150 2087 -116
rect 2145 -150 2179 -116
rect 2237 -150 2271 -116
rect 2329 -150 2363 -116
rect 2421 -150 2455 -116
rect 2513 -150 2547 -116
rect 2605 -150 2639 -116
rect 2697 -150 2731 -116
rect 2789 -150 2823 -116
rect 2881 -150 2915 -116
rect 2973 -150 3007 -116
rect 3065 -150 3099 -116
rect 3157 -150 3191 -116
rect 3249 -150 3283 -116
rect 3341 -150 3375 -116
rect 3433 -150 3467 -116
rect 3525 -150 3559 -116
rect 3617 -150 3651 -116
rect 3709 -150 3743 -116
rect 3801 -150 3835 -116
rect 3893 -150 3927 -116
rect 3985 -150 4019 -116
rect 4077 -150 4111 -116
rect 4169 -150 4203 -116
rect 4261 -150 4295 -116
rect 4353 -150 4387 -116
rect 4445 -150 4479 -116
rect 4537 -150 4571 -116
rect 4629 -150 4663 -116
rect 4721 -150 4755 -116
rect 4813 -150 4847 -116
rect 4905 -150 4939 -116
rect 4997 -150 5031 -116
rect 5089 -150 5123 -116
rect 5181 -150 5215 -116
rect 5273 -150 5307 -116
rect 5365 -150 5399 -116
rect 5457 -150 5491 -116
rect 5549 -150 5583 -116
rect 5641 -150 5675 -116
rect 5733 -150 5767 -116
rect 5825 -150 5859 -116
rect 5917 -150 5951 -116
rect 6009 -150 6043 -116
rect 6101 -150 6135 -116
rect 6193 -150 6227 -116
rect 6285 -150 6319 -116
rect 6377 -150 6411 -116
rect 6469 -150 6503 -116
rect 6561 -150 6595 -116
rect 6653 -150 6687 -116
rect 6745 -150 6779 -116
rect 6837 -150 6871 -116
rect 6929 -150 6963 -116
rect 7021 -150 7055 -116
rect 7113 -150 7147 -116
rect 7205 -150 7239 -116
rect 7297 -150 7331 -116
rect 7389 -150 7423 -116
rect 7481 -150 7515 -116
rect 7573 -150 7607 -116
rect 7665 -150 7699 -116
rect 7757 -150 7791 -116
rect 7849 -150 7883 -116
rect 7941 -150 7975 -116
rect 8033 -150 8067 -116
rect 8125 -150 8159 -116
rect 8217 -150 8251 -116
rect 8309 -150 8343 -116
rect 8401 -150 8435 -116
rect 8493 -150 8527 -116
rect 8585 -150 8619 -116
rect 8677 -150 8711 -116
rect 8769 -150 8803 -116
rect 8861 -150 8895 -116
rect 8953 -150 8987 -116
rect 9045 -150 9079 -116
rect 9137 -150 9171 -116
rect 9229 -150 9263 -116
rect 9321 -150 9355 -116
rect 9413 -150 9447 -116
rect 9505 -150 9539 -116
rect 9597 -150 9631 -116
rect 9689 -150 9723 -116
rect 9781 -150 9815 -116
rect 9873 -150 9907 -116
rect 9965 -150 9999 -116
rect 10057 -150 10091 -116
rect 10149 -150 10183 -116
rect 10241 -150 10275 -116
rect 10333 -150 10367 -116
rect 10425 -150 10459 -116
rect 10517 -150 10551 -116
rect 10609 -150 10643 -116
rect 10701 -150 10735 -116
rect 10793 -150 10827 -116
rect 10885 -150 10919 -116
rect 10977 -150 11011 -116
rect 11069 -150 11103 -116
rect 11161 -150 11195 -116
rect 11253 -150 11287 -116
rect 11345 -150 11379 -116
rect 11437 -150 11471 -116
rect 11529 -150 11563 -116
rect 11621 -150 11655 -116
rect 11713 -150 11747 -116
rect 11805 -150 11839 -116
rect 11897 -150 11931 -116
rect 11989 -150 12023 -116
rect 12081 -150 12115 -116
rect 12173 -150 12207 -116
rect 12265 -150 12299 -116
rect 12357 -150 12391 -116
rect 12449 -150 12483 -116
rect 12541 -150 12575 -116
rect 12633 -150 12667 -116
rect 12725 -150 12759 -116
rect 12817 -150 12851 -116
rect 12909 -150 12943 -116
rect 13001 -150 13035 -116
rect 13093 -150 13127 -116
rect 13185 -150 13219 -116
rect 13277 -150 13311 -116
rect 13369 -150 13403 -116
rect 13461 -150 13495 -116
rect 13553 -150 13587 -116
rect 13645 -150 13679 -116
rect 13737 -150 13771 -116
rect 13829 -150 13863 -116
rect 13921 -150 13955 -116
rect 14013 -150 14047 -116
rect 14105 -150 14139 -116
rect 14197 -150 14231 -116
rect 14289 -150 14323 -116
rect 14381 -150 14415 -116
rect 14473 -150 14507 -116
rect 14565 -150 14599 -116
rect 14657 -150 14691 -116
rect 14749 -150 14783 -116
rect 14841 -150 14875 -116
rect 14933 -150 14967 -116
rect 15025 -150 15059 -116
rect 15117 -150 15151 -116
rect 15209 -150 15243 -116
rect 15301 -150 15335 -116
rect 15393 -150 15427 -116
rect 15485 -150 15519 -116
rect 15577 -150 15611 -116
rect 15669 -150 15703 -116
rect 15761 -150 15795 -116
rect 15853 -150 15887 -116
rect 15945 -150 15979 -116
rect 16037 -150 16071 -116
rect 16129 -150 16163 -116
rect 16221 -150 16255 -116
rect 16313 -150 16347 -116
rect 16405 -150 16439 -116
rect 16497 -150 16531 -116
rect 16589 -150 16623 -116
rect 16681 -150 16715 -116
<< nsubdiffcont >>
rect 31 2961 65 2995
rect 123 2961 157 2995
rect 215 2961 249 2995
rect 307 2961 341 2995
rect 399 2961 433 2995
rect 491 2961 525 2995
rect 583 2961 617 2995
rect 675 2961 709 2995
rect 767 2961 801 2995
rect 859 2961 893 2995
rect 951 2961 985 2995
rect 1043 2961 1077 2995
rect 1135 2961 1169 2995
rect 1227 2961 1261 2995
rect 1319 2961 1353 2995
rect 1411 2961 1445 2995
rect 1503 2961 1537 2995
rect 1595 2961 1629 2995
rect 1687 2961 1721 2995
rect 1779 2961 1813 2995
rect 1871 2961 1905 2995
rect 1963 2961 1997 2995
rect 2055 2961 2089 2995
rect 2147 2961 2181 2995
rect 2239 2961 2273 2995
rect 2331 2961 2365 2995
rect 2423 2961 2457 2995
rect 2515 2961 2549 2995
rect 2607 2961 2641 2995
rect 2699 2961 2733 2995
rect 2791 2961 2825 2995
rect 4415 2961 4449 2995
rect 4507 2961 4541 2995
rect 4599 2961 4633 2995
rect 4691 2961 4725 2995
rect 4783 2961 4817 2995
rect 4875 2961 4909 2995
rect 4967 2961 5001 2995
rect 5059 2961 5093 2995
rect 5151 2961 5185 2995
rect 5243 2961 5277 2995
rect 5335 2961 5369 2995
rect 5427 2961 5461 2995
rect 5519 2961 5553 2995
rect 5611 2961 5645 2995
rect 5703 2961 5737 2995
rect 5795 2961 5829 2995
rect 5887 2961 5921 2995
rect 5979 2961 6013 2995
rect 6071 2961 6105 2995
rect 6163 2961 6197 2995
rect 6255 2961 6289 2995
rect 6347 2961 6381 2995
rect 6439 2961 6473 2995
rect 6531 2961 6565 2995
rect 6623 2961 6657 2995
rect 6715 2961 6749 2995
rect 6807 2961 6841 2995
rect 6899 2961 6933 2995
rect 6991 2961 7025 2995
rect 7083 2961 7117 2995
rect 7175 2961 7209 2995
rect 29 1819 63 1853
rect 121 1819 155 1853
rect 213 1819 247 1853
rect 305 1819 339 1853
rect 397 1819 431 1853
rect 489 1819 523 1853
rect 581 1819 615 1853
rect 673 1819 707 1853
rect 765 1819 799 1853
rect 857 1819 891 1853
rect 949 1819 983 1853
rect 1041 1819 1075 1853
rect 1133 1819 1167 1853
rect 1225 1819 1259 1853
rect 1317 1819 1351 1853
rect 1409 1819 1443 1853
rect 1501 1819 1535 1853
rect 1593 1819 1627 1853
rect 1685 1819 1719 1853
rect 1777 1819 1811 1853
rect 1869 1819 1903 1853
rect 1961 1819 1995 1853
rect 2053 1819 2087 1853
rect 2145 1819 2179 1853
rect 2237 1819 2271 1853
rect 2329 1819 2363 1853
rect 2421 1819 2455 1853
rect 2513 1819 2547 1853
rect 2605 1819 2639 1853
rect 2697 1819 2731 1853
rect 2789 1819 2823 1853
rect 2881 1819 2915 1853
rect 2973 1819 3007 1853
rect 3065 1819 3099 1853
rect 3157 1819 3191 1853
rect 3249 1819 3283 1853
rect 3341 1819 3375 1853
rect 3433 1819 3467 1853
rect 3525 1819 3559 1853
rect 3617 1819 3651 1853
rect 3709 1819 3743 1853
rect 3801 1819 3835 1853
rect 3893 1819 3927 1853
rect 3985 1819 4019 1853
rect 4077 1819 4111 1853
rect 4169 1819 4203 1853
rect 4261 1819 4295 1853
rect 4353 1819 4387 1853
rect 4445 1819 4479 1853
rect 4537 1819 4571 1853
rect 4629 1819 4663 1853
rect 4721 1819 4755 1853
rect 4813 1819 4847 1853
rect 4905 1819 4939 1853
rect 4997 1819 5031 1853
rect 5089 1819 5123 1853
rect 5181 1819 5215 1853
rect 5273 1819 5307 1853
rect 5365 1819 5399 1853
rect 5457 1819 5491 1853
rect 5549 1819 5583 1853
rect 5641 1819 5675 1853
rect 6245 1819 6279 1853
rect 6337 1819 6371 1853
rect 6429 1819 6463 1853
rect 6521 1819 6555 1853
rect 6613 1819 6647 1853
rect 6705 1819 6739 1853
rect 6797 1819 6831 1853
rect 6889 1819 6923 1853
rect 6981 1819 7015 1853
rect 7073 1819 7107 1853
rect 7165 1819 7199 1853
rect 7257 1819 7291 1853
rect 7349 1819 7383 1853
rect 7441 1819 7475 1853
rect 7533 1819 7567 1853
rect 7625 1819 7659 1853
rect 7717 1819 7751 1853
rect 7809 1819 7843 1853
rect 7901 1819 7935 1853
rect 7993 1819 8027 1853
rect 8085 1819 8119 1853
rect 8177 1819 8211 1853
rect 8269 1819 8303 1853
rect 8361 1819 8395 1853
rect 8453 1819 8487 1853
rect 8545 1819 8579 1853
rect 8637 1819 8671 1853
rect 8729 1819 8763 1853
rect 8821 1819 8855 1853
rect 8913 1819 8947 1853
rect 9005 1819 9039 1853
rect 9097 1819 9131 1853
rect 9189 1819 9223 1853
rect 9281 1819 9315 1853
rect 9373 1819 9407 1853
rect 9465 1819 9499 1853
rect 9557 1819 9591 1853
rect 9649 1819 9683 1853
rect 9741 1819 9775 1853
rect 9833 1819 9867 1853
rect 9925 1819 9959 1853
rect 10017 1819 10051 1853
rect 10109 1819 10143 1853
rect 10201 1819 10235 1853
rect 10293 1819 10327 1853
rect 10385 1819 10419 1853
rect 10477 1819 10511 1853
rect 10569 1819 10603 1853
rect 10661 1819 10695 1853
rect 10753 1819 10787 1853
rect 10845 1819 10879 1853
rect 10937 1819 10971 1853
rect 11029 1819 11063 1853
rect 11121 1819 11155 1853
rect 11213 1819 11247 1853
rect 11305 1819 11339 1853
rect 11397 1819 11431 1853
rect 11489 1819 11523 1853
rect 11581 1819 11615 1853
rect 11673 1819 11707 1853
rect 11765 1819 11799 1853
rect 11857 1819 11891 1853
rect 12011 1819 12045 1853
rect 12103 1819 12137 1853
rect 12195 1819 12229 1853
rect 12287 1819 12321 1853
rect 12379 1819 12413 1853
rect 12471 1819 12505 1853
rect 12563 1819 12597 1853
rect 12655 1819 12689 1853
rect 12747 1819 12781 1853
rect 12839 1819 12873 1853
rect 12931 1819 12965 1853
rect 13023 1819 13057 1853
rect 13115 1819 13149 1853
rect 13207 1819 13241 1853
rect 13299 1819 13333 1853
rect 13391 1819 13425 1853
rect 13483 1819 13517 1853
rect 13575 1819 13609 1853
rect 13667 1819 13701 1853
rect 13759 1819 13793 1853
rect 13851 1819 13885 1853
rect 13943 1819 13977 1853
rect 14035 1819 14069 1853
rect 14127 1819 14161 1853
rect 14219 1819 14253 1853
rect 14311 1819 14345 1853
rect 14403 1819 14437 1853
rect 14495 1819 14529 1853
rect 14587 1819 14621 1853
rect 14679 1819 14713 1853
rect 14771 1819 14805 1853
rect 14863 1819 14897 1853
rect 14955 1819 14989 1853
rect 15047 1819 15081 1853
rect 15139 1819 15173 1853
rect 15231 1819 15265 1853
rect 15323 1819 15357 1853
rect 15415 1819 15449 1853
rect 15507 1819 15541 1853
rect 15599 1819 15633 1853
rect 15691 1819 15725 1853
rect 15783 1819 15817 1853
rect 15875 1819 15909 1853
rect 15967 1819 16001 1853
rect 16059 1819 16093 1853
rect 16151 1819 16185 1853
rect 16243 1819 16277 1853
rect 16335 1819 16369 1853
rect 16427 1819 16461 1853
rect 16519 1819 16553 1853
rect 29 1131 63 1165
rect 121 1131 155 1165
rect 213 1131 247 1165
rect 305 1131 339 1165
rect 397 1131 431 1165
rect 489 1131 523 1165
rect 581 1131 615 1165
rect 673 1131 707 1165
rect 765 1131 799 1165
rect 857 1131 891 1165
rect 949 1131 983 1165
rect 1041 1131 1075 1165
rect 1133 1131 1167 1165
rect 1225 1131 1259 1165
rect 1317 1131 1351 1165
rect 1409 1131 1443 1165
rect 1501 1131 1535 1165
rect 1593 1131 1627 1165
rect 1685 1131 1719 1165
rect 1777 1131 1811 1165
rect 2053 1131 2087 1165
rect 2145 1131 2179 1165
rect 2237 1131 2271 1165
rect 2329 1131 2363 1165
rect 2421 1131 2455 1165
rect 2513 1131 2547 1165
rect 2605 1131 2639 1165
rect 2697 1131 2731 1165
rect 2789 1131 2823 1165
rect 2881 1131 2915 1165
rect 2973 1131 3007 1165
rect 3065 1131 3099 1165
rect 3157 1131 3191 1165
rect 3249 1131 3283 1165
rect 3341 1131 3375 1165
rect 3433 1131 3467 1165
rect 3525 1131 3559 1165
rect 3617 1131 3651 1165
rect 3709 1131 3743 1165
rect 3801 1131 3835 1165
rect 3893 1131 3927 1165
rect 3985 1131 4019 1165
rect 4077 1131 4111 1165
rect 4169 1131 4203 1165
rect 4445 1131 4479 1165
rect 4537 1131 4571 1165
rect 4629 1131 4663 1165
rect 4721 1131 4755 1165
rect 4813 1131 4847 1165
rect 4905 1131 4939 1165
rect 4997 1131 5031 1165
rect 5089 1131 5123 1165
rect 5181 1131 5215 1165
rect 5273 1131 5307 1165
rect 5365 1131 5399 1165
rect 5457 1131 5491 1165
rect 5549 1131 5583 1165
rect 5641 1131 5675 1165
rect 5733 1131 5767 1165
rect 5825 1131 5859 1165
rect 5917 1131 5951 1165
rect 6009 1131 6043 1165
rect 6101 1131 6135 1165
rect 6193 1131 6227 1165
rect 6285 1131 6319 1165
rect 6377 1131 6411 1165
rect 6469 1131 6503 1165
rect 6561 1131 6595 1165
rect 6837 1131 6871 1165
rect 6929 1131 6963 1165
rect 7021 1131 7055 1165
rect 7113 1131 7147 1165
rect 7205 1131 7239 1165
rect 7297 1131 7331 1165
rect 7389 1131 7423 1165
rect 7481 1131 7515 1165
rect 7573 1131 7607 1165
rect 7665 1131 7699 1165
rect 7757 1131 7791 1165
rect 7849 1131 7883 1165
rect 7941 1131 7975 1165
rect 8033 1131 8067 1165
rect 8125 1131 8159 1165
rect 8217 1131 8251 1165
rect 8309 1131 8343 1165
rect 8401 1131 8435 1165
rect 8493 1131 8527 1165
rect 8585 1131 8619 1165
rect 8677 1131 8711 1165
rect 8769 1131 8803 1165
rect 8861 1131 8895 1165
rect 8953 1131 8987 1165
rect 9229 1131 9263 1165
rect 9321 1131 9355 1165
rect 9413 1131 9447 1165
rect 9505 1131 9539 1165
rect 9597 1131 9631 1165
rect 9689 1131 9723 1165
rect 9781 1131 9815 1165
rect 9873 1131 9907 1165
rect 9965 1131 9999 1165
rect 10057 1131 10091 1165
rect 10149 1131 10183 1165
rect 10241 1131 10275 1165
rect 10333 1131 10367 1165
rect 10425 1131 10459 1165
rect 10517 1131 10551 1165
rect 10609 1131 10643 1165
rect 10701 1131 10735 1165
rect 10793 1131 10827 1165
rect 10885 1131 10919 1165
rect 10977 1131 11011 1165
rect 11069 1131 11103 1165
rect 11161 1131 11195 1165
rect 11253 1131 11287 1165
rect 11345 1131 11379 1165
rect 11621 1131 11655 1165
rect 11713 1131 11747 1165
rect 11805 1131 11839 1165
rect 11897 1131 11931 1165
rect 11989 1131 12023 1165
rect 12081 1131 12115 1165
rect 12173 1131 12207 1165
rect 12265 1131 12299 1165
rect 12357 1131 12391 1165
rect 12449 1131 12483 1165
rect 12541 1131 12575 1165
rect 12633 1131 12667 1165
rect 12725 1131 12759 1165
rect 12817 1131 12851 1165
rect 12909 1131 12943 1165
rect 13001 1131 13035 1165
rect 13093 1131 13127 1165
rect 13185 1131 13219 1165
rect 13277 1131 13311 1165
rect 13369 1131 13403 1165
rect 13461 1131 13495 1165
rect 13553 1131 13587 1165
rect 13645 1131 13679 1165
rect 13737 1131 13771 1165
rect 14013 1131 14047 1165
rect 14105 1131 14139 1165
rect 14197 1131 14231 1165
rect 14289 1131 14323 1165
rect 14381 1131 14415 1165
rect 14473 1131 14507 1165
rect 14565 1131 14599 1165
rect 14657 1131 14691 1165
rect 14749 1131 14783 1165
rect 14841 1131 14875 1165
rect 14933 1131 14967 1165
rect 15025 1131 15059 1165
rect 15117 1131 15151 1165
rect 15209 1131 15243 1165
rect 15301 1131 15335 1165
rect 15393 1131 15427 1165
rect 15485 1131 15519 1165
rect 15577 1131 15611 1165
rect 15669 1131 15703 1165
rect 15761 1131 15795 1165
rect 15853 1131 15887 1165
rect 15945 1131 15979 1165
rect 16037 1131 16071 1165
rect 16129 1131 16163 1165
rect 16405 1131 16439 1165
rect 16497 1131 16531 1165
rect 16589 1131 16623 1165
rect 16681 1131 16715 1165
rect 29 442 63 476
rect 121 442 155 476
rect 213 442 247 476
rect 305 442 339 476
rect 394 442 428 476
rect 496 442 530 476
rect 581 442 615 476
rect 673 442 707 476
rect 765 442 799 476
rect 857 442 891 476
rect 949 442 983 476
rect 1041 442 1075 476
rect 1133 442 1167 476
rect 1225 442 1259 476
rect 1317 442 1351 476
rect 1409 442 1443 476
rect 1501 442 1535 476
rect 1777 442 1811 476
rect 1869 442 1903 476
rect 1961 442 1995 476
rect 2053 442 2087 476
rect 2145 442 2179 476
rect 2237 442 2271 476
rect 2329 442 2363 476
rect 2421 442 2455 476
rect 2513 442 2547 476
rect 2605 442 2639 476
rect 2697 442 2731 476
rect 2791 442 2825 476
rect 2882 442 2916 476
rect 2973 442 3007 476
rect 3065 442 3099 476
rect 3157 442 3191 476
rect 3249 442 3283 476
rect 3341 442 3375 476
rect 3433 442 3467 476
rect 3525 442 3559 476
rect 3617 442 3651 476
rect 3709 442 3743 476
rect 3801 442 3835 476
rect 3893 442 3927 476
rect 4169 442 4203 476
rect 4261 442 4295 476
rect 4353 442 4387 476
rect 4445 442 4479 476
rect 4537 442 4571 476
rect 4629 442 4663 476
rect 4721 442 4755 476
rect 4813 442 4847 476
rect 4905 442 4939 476
rect 4997 442 5031 476
rect 5089 442 5123 476
rect 5179 442 5213 476
rect 5273 442 5307 476
rect 5365 442 5399 476
rect 5457 442 5491 476
rect 5549 442 5583 476
rect 5641 442 5675 476
rect 5733 442 5767 476
rect 5825 442 5859 476
rect 5917 442 5951 476
rect 6009 442 6043 476
rect 6101 442 6135 476
rect 6193 442 6227 476
rect 6285 442 6319 476
rect 6561 442 6595 476
rect 6653 442 6687 476
rect 6745 442 6779 476
rect 6837 442 6871 476
rect 6929 442 6963 476
rect 7021 442 7055 476
rect 7113 442 7147 476
rect 7205 442 7239 476
rect 7297 442 7331 476
rect 7389 442 7423 476
rect 7481 442 7515 476
rect 7574 442 7608 476
rect 7665 442 7699 476
rect 7757 442 7791 476
rect 7849 442 7883 476
rect 7941 442 7975 476
rect 8033 442 8067 476
rect 8125 442 8159 476
rect 8217 442 8251 476
rect 8309 442 8343 476
rect 8401 442 8435 476
rect 8493 442 8527 476
rect 8585 442 8619 476
rect 8677 442 8711 476
rect 8953 442 8987 476
rect 9045 442 9079 476
rect 9137 442 9171 476
rect 9229 442 9263 476
rect 9321 442 9355 476
rect 9413 442 9447 476
rect 9505 442 9539 476
rect 9597 442 9631 476
rect 9689 442 9723 476
rect 9781 442 9815 476
rect 9873 442 9907 476
rect 9963 442 9997 476
rect 10058 442 10092 476
rect 10149 442 10183 476
rect 10241 442 10275 476
rect 10333 442 10367 476
rect 10425 442 10459 476
rect 10517 442 10551 476
rect 10609 442 10643 476
rect 10701 442 10735 476
rect 10793 442 10827 476
rect 10885 442 10919 476
rect 10977 442 11011 476
rect 11069 442 11103 476
rect 11345 442 11379 476
rect 11437 442 11471 476
rect 11529 442 11563 476
rect 11621 442 11655 476
rect 11713 442 11747 476
rect 11805 442 11839 476
rect 11897 442 11931 476
rect 11989 442 12023 476
rect 12081 442 12115 476
rect 12173 442 12207 476
rect 12265 442 12299 476
rect 12357 442 12391 476
rect 12448 442 12482 476
rect 12541 442 12575 476
rect 12633 442 12667 476
rect 12725 442 12759 476
rect 12817 442 12851 476
rect 12909 442 12943 476
rect 13001 442 13035 476
rect 13093 442 13127 476
rect 13185 442 13219 476
rect 13277 442 13311 476
rect 13369 442 13403 476
rect 13461 442 13495 476
rect 13737 442 13771 476
rect 13829 442 13863 476
rect 13921 442 13955 476
rect 14013 442 14047 476
rect 14105 442 14139 476
rect 14197 442 14231 476
rect 14289 442 14323 476
rect 14381 442 14415 476
rect 14473 442 14507 476
rect 14565 442 14599 476
rect 14657 442 14691 476
rect 14748 442 14782 476
rect 14842 442 14876 476
rect 14933 442 14967 476
rect 15025 442 15059 476
rect 15117 442 15151 476
rect 15209 442 15243 476
rect 15301 442 15335 476
rect 15393 442 15427 476
rect 15485 442 15519 476
rect 15577 442 15611 476
rect 15669 442 15703 476
rect 15761 442 15795 476
rect 15853 442 15887 476
rect 16129 442 16163 476
rect 16221 442 16255 476
rect 16313 442 16347 476
rect 16405 442 16439 476
rect 16497 442 16531 476
rect 16589 442 16623 476
rect 16681 442 16715 476
<< poly >>
rect 1885 1158 1951 1174
rect 1885 1124 1901 1158
rect 1935 1124 1951 1158
rect 4277 1157 4343 1173
rect 1885 1108 1951 1124
rect 4277 1123 4293 1157
rect 4327 1123 4343 1157
rect 6669 1157 6735 1173
rect 1903 1030 1933 1108
rect 4277 1107 4343 1123
rect 6669 1123 6685 1157
rect 6719 1123 6735 1157
rect 9061 1158 9127 1174
rect 6669 1107 6735 1123
rect 9061 1124 9077 1158
rect 9111 1124 9127 1158
rect 11453 1158 11519 1174
rect 9061 1108 9127 1124
rect 11453 1124 11469 1158
rect 11503 1124 11519 1158
rect 13845 1157 13911 1173
rect 11453 1108 11519 1124
rect 13845 1123 13861 1157
rect 13895 1123 13911 1157
rect 16237 1157 16303 1173
rect 4295 1029 4325 1107
rect 6687 1029 6717 1107
rect 9079 1030 9109 1108
rect 11471 1030 11501 1108
rect 13845 1107 13911 1123
rect 16237 1123 16253 1157
rect 16287 1123 16303 1157
rect 16237 1107 16303 1123
rect 13863 1029 13893 1107
rect 16255 1029 16285 1107
rect 1591 472 1657 488
rect 1591 438 1607 472
rect 1641 438 1657 472
rect 3983 472 4049 488
rect 1591 422 1657 438
rect 3983 438 3999 472
rect 4033 438 4049 472
rect 6375 472 6441 488
rect 3983 422 4049 438
rect 6375 438 6391 472
rect 6425 438 6441 472
rect 8767 472 8833 488
rect 6375 422 6441 438
rect 8767 438 8783 472
rect 8817 438 8833 472
rect 11159 472 11225 488
rect 8767 422 8833 438
rect 11159 438 11175 472
rect 11209 438 11225 472
rect 13551 472 13617 488
rect 11159 422 11225 438
rect 13551 438 13567 472
rect 13601 438 13617 472
rect 15943 469 16009 485
rect 13551 422 13617 438
rect 15943 435 15959 469
rect 15993 435 16009 469
rect 1609 390 1639 422
rect 4001 390 4031 422
rect 6393 390 6423 422
rect 8785 390 8815 422
rect 11177 390 11207 422
rect 13569 390 13599 422
rect 15943 419 16009 435
rect 15961 388 15991 419
<< polycont >>
rect 1901 1124 1935 1158
rect 4293 1123 4327 1157
rect 6685 1123 6719 1157
rect 9077 1124 9111 1158
rect 11469 1124 11503 1158
rect 13861 1123 13895 1157
rect 16253 1123 16287 1157
rect 1607 438 1641 472
rect 3999 438 4033 472
rect 6391 438 6425 472
rect 8783 438 8817 472
rect 11175 438 11209 472
rect 13567 438 13601 472
rect 15959 435 15993 469
<< locali >>
rect 2 2961 31 2995
rect 65 2961 123 2995
rect 157 2961 215 2995
rect 249 2961 307 2995
rect 341 2961 399 2995
rect 433 2961 491 2995
rect 525 2961 583 2995
rect 617 2961 675 2995
rect 709 2961 767 2995
rect 801 2961 859 2995
rect 893 2961 951 2995
rect 985 2961 1043 2995
rect 1077 2961 1135 2995
rect 1169 2961 1227 2995
rect 1261 2961 1319 2995
rect 1353 2961 1411 2995
rect 1445 2961 1503 2995
rect 1537 2961 1595 2995
rect 1629 2961 1687 2995
rect 1721 2961 1779 2995
rect 1813 2961 1871 2995
rect 1905 2961 1963 2995
rect 1997 2961 2055 2995
rect 2089 2961 2147 2995
rect 2181 2961 2239 2995
rect 2273 2961 2331 2995
rect 2365 2961 2423 2995
rect 2457 2961 2515 2995
rect 2549 2961 2607 2995
rect 2641 2961 2699 2995
rect 2733 2961 2791 2995
rect 2825 2961 2854 2995
rect 2 2954 2854 2961
rect 4386 2961 4415 2995
rect 4449 2961 4507 2995
rect 4541 2961 4599 2995
rect 4633 2961 4691 2995
rect 4725 2961 4783 2995
rect 4817 2961 4875 2995
rect 4909 2961 4967 2995
rect 5001 2961 5059 2995
rect 5093 2961 5151 2995
rect 5185 2961 5243 2995
rect 5277 2961 5335 2995
rect 5369 2961 5427 2995
rect 5461 2961 5519 2995
rect 5553 2961 5611 2995
rect 5645 2961 5703 2995
rect 5737 2961 5795 2995
rect 5829 2961 5887 2995
rect 5921 2961 5979 2995
rect 6013 2961 6071 2995
rect 6105 2961 6163 2995
rect 6197 2961 6255 2995
rect 6289 2961 6347 2995
rect 6381 2961 6439 2995
rect 6473 2961 6531 2995
rect 6565 2961 6623 2995
rect 6657 2961 6715 2995
rect 6749 2961 6807 2995
rect 6841 2961 6899 2995
rect 6933 2961 6991 2995
rect 7025 2961 7083 2995
rect 7117 2961 7175 2995
rect 7209 2961 7238 2995
rect 4386 2955 7238 2961
rect 232 2626 350 2670
rect 2810 2664 2915 2665
rect 666 2626 874 2664
rect 2810 2630 2876 2664
rect 2910 2630 2915 2664
rect 2810 2629 2915 2630
rect 4630 2626 4692 2672
rect 5032 2626 5238 2666
rect 3 2403 2854 2410
rect 2 2369 31 2403
rect 65 2369 123 2403
rect 157 2369 215 2403
rect 249 2369 307 2403
rect 341 2369 399 2403
rect 433 2369 491 2403
rect 525 2369 583 2403
rect 617 2369 675 2403
rect 709 2369 767 2403
rect 801 2369 859 2403
rect 893 2369 951 2403
rect 985 2369 1043 2403
rect 1077 2369 1135 2403
rect 1169 2369 1227 2403
rect 1261 2369 1319 2403
rect 1353 2369 1411 2403
rect 1445 2369 1503 2403
rect 1537 2369 1595 2403
rect 1629 2369 1687 2403
rect 1721 2369 1779 2403
rect 1813 2369 1871 2403
rect 1905 2369 1963 2403
rect 1997 2369 2055 2403
rect 2089 2369 2147 2403
rect 2181 2369 2239 2403
rect 2273 2369 2331 2403
rect 2365 2369 2423 2403
rect 2457 2369 2515 2403
rect 2549 2369 2607 2403
rect 2641 2369 2699 2403
rect 2733 2369 2791 2403
rect 2825 2369 2854 2403
rect 4386 2403 7238 2410
rect 4386 2369 4415 2403
rect 4449 2369 4507 2403
rect 4541 2369 4599 2403
rect 4633 2369 4691 2403
rect 4725 2369 4783 2403
rect 4817 2369 4875 2403
rect 4909 2369 4967 2403
rect 5001 2369 5059 2403
rect 5093 2369 5151 2403
rect 5185 2369 5243 2403
rect 5277 2369 5335 2403
rect 5369 2369 5427 2403
rect 5461 2369 5519 2403
rect 5553 2369 5611 2403
rect 5645 2369 5703 2403
rect 5737 2369 5795 2403
rect 5829 2369 5887 2403
rect 5921 2369 5979 2403
rect 6013 2369 6071 2403
rect 6105 2369 6163 2403
rect 6197 2369 6255 2403
rect 6289 2369 6347 2403
rect 6381 2369 6439 2403
rect 6473 2369 6531 2403
rect 6565 2369 6623 2403
rect 6657 2369 6715 2403
rect 6749 2369 6807 2403
rect 6841 2369 6899 2403
rect 6933 2369 6991 2403
rect 7025 2369 7083 2403
rect 7117 2369 7175 2403
rect 7209 2369 7238 2403
rect 0 1819 29 1853
rect 63 1819 121 1853
rect 155 1819 213 1853
rect 247 1819 305 1853
rect 339 1819 397 1853
rect 431 1819 489 1853
rect 523 1819 581 1853
rect 615 1819 673 1853
rect 707 1819 765 1853
rect 799 1819 857 1853
rect 891 1819 949 1853
rect 983 1819 1041 1853
rect 1075 1819 1133 1853
rect 1167 1819 1225 1853
rect 1259 1819 1317 1853
rect 1351 1819 1409 1853
rect 1443 1819 1501 1853
rect 1535 1819 1593 1853
rect 1627 1819 1685 1853
rect 1719 1819 1777 1853
rect 1811 1819 1869 1853
rect 1903 1819 1961 1853
rect 1995 1819 2053 1853
rect 2087 1819 2145 1853
rect 2179 1819 2237 1853
rect 2271 1819 2329 1853
rect 2363 1819 2421 1853
rect 2455 1819 2513 1853
rect 2547 1819 2605 1853
rect 2639 1819 2697 1853
rect 2731 1819 2789 1853
rect 2823 1819 2881 1853
rect 2915 1819 2973 1853
rect 3007 1819 3065 1853
rect 3099 1819 3157 1853
rect 3191 1819 3249 1853
rect 3283 1819 3341 1853
rect 3375 1819 3433 1853
rect 3467 1819 3525 1853
rect 3559 1819 3617 1853
rect 3651 1819 3709 1853
rect 3743 1819 3801 1853
rect 3835 1819 3893 1853
rect 3927 1819 3985 1853
rect 4019 1819 4077 1853
rect 4111 1819 4169 1853
rect 4203 1819 4261 1853
rect 4295 1819 4353 1853
rect 4387 1819 4445 1853
rect 4479 1819 4537 1853
rect 4571 1819 4629 1853
rect 4663 1819 4721 1853
rect 4755 1819 4813 1853
rect 4847 1819 4905 1853
rect 4939 1819 4997 1853
rect 5031 1819 5089 1853
rect 5123 1819 5181 1853
rect 5215 1819 5273 1853
rect 5307 1819 5365 1853
rect 5399 1819 5457 1853
rect 5491 1819 5549 1853
rect 5583 1819 5641 1853
rect 5675 1819 6245 1853
rect 6279 1819 6337 1853
rect 6371 1819 6429 1853
rect 6463 1819 6521 1853
rect 6555 1819 6613 1853
rect 6647 1819 6705 1853
rect 6739 1819 6797 1853
rect 6831 1819 6889 1853
rect 6923 1819 6981 1853
rect 7015 1819 7073 1853
rect 7107 1819 7165 1853
rect 7199 1819 7257 1853
rect 7291 1819 7349 1853
rect 7383 1819 7441 1853
rect 7475 1819 7533 1853
rect 7567 1819 7625 1853
rect 7659 1819 7717 1853
rect 7751 1819 7809 1853
rect 7843 1819 7901 1853
rect 7935 1819 7993 1853
rect 8027 1819 8085 1853
rect 8119 1819 8177 1853
rect 8211 1819 8269 1853
rect 8303 1819 8361 1853
rect 8395 1819 8453 1853
rect 8487 1819 8545 1853
rect 8579 1819 8637 1853
rect 8671 1819 8729 1853
rect 8763 1819 8821 1853
rect 8855 1819 8913 1853
rect 8947 1819 9005 1853
rect 9039 1819 9097 1853
rect 9131 1819 9189 1853
rect 9223 1819 9281 1853
rect 9315 1819 9373 1853
rect 9407 1819 9465 1853
rect 9499 1819 9557 1853
rect 9591 1819 9649 1853
rect 9683 1819 9741 1853
rect 9775 1819 9833 1853
rect 9867 1819 9925 1853
rect 9959 1819 10017 1853
rect 10051 1819 10109 1853
rect 10143 1819 10201 1853
rect 10235 1819 10293 1853
rect 10327 1819 10385 1853
rect 10419 1819 10477 1853
rect 10511 1819 10569 1853
rect 10603 1819 10661 1853
rect 10695 1819 10753 1853
rect 10787 1819 10845 1853
rect 10879 1819 10937 1853
rect 10971 1819 11029 1853
rect 11063 1819 11121 1853
rect 11155 1819 11213 1853
rect 11247 1819 11305 1853
rect 11339 1819 11397 1853
rect 11431 1819 11489 1853
rect 11523 1819 11581 1853
rect 11615 1819 11673 1853
rect 11707 1819 11765 1853
rect 11799 1819 11857 1853
rect 11891 1819 12011 1853
rect 12045 1819 12103 1853
rect 12137 1819 12195 1853
rect 12229 1819 12287 1853
rect 12321 1819 12379 1853
rect 12413 1819 12471 1853
rect 12505 1819 12563 1853
rect 12597 1819 12655 1853
rect 12689 1819 12747 1853
rect 12781 1819 12839 1853
rect 12873 1819 12931 1853
rect 12965 1819 13023 1853
rect 13057 1819 13115 1853
rect 13149 1819 13207 1853
rect 13241 1819 13299 1853
rect 13333 1819 13391 1853
rect 13425 1819 13483 1853
rect 13517 1819 13575 1853
rect 13609 1819 13667 1853
rect 13701 1819 13759 1853
rect 13793 1819 13851 1853
rect 13885 1819 13943 1853
rect 13977 1819 14035 1853
rect 14069 1819 14127 1853
rect 14161 1819 14219 1853
rect 14253 1819 14311 1853
rect 14345 1819 14403 1853
rect 14437 1819 14495 1853
rect 14529 1819 14587 1853
rect 14621 1819 14679 1853
rect 14713 1819 14771 1853
rect 14805 1819 14863 1853
rect 14897 1819 14955 1853
rect 14989 1819 15047 1853
rect 15081 1819 15139 1853
rect 15173 1819 15231 1853
rect 15265 1819 15323 1853
rect 15357 1819 15415 1853
rect 15449 1819 15507 1853
rect 15541 1819 15599 1853
rect 15633 1819 15691 1853
rect 15725 1819 15783 1853
rect 15817 1819 15875 1853
rect 15909 1819 15967 1853
rect 16001 1819 16059 1853
rect 16093 1819 16151 1853
rect 16185 1819 16243 1853
rect 16277 1819 16335 1853
rect 16369 1819 16427 1853
rect 16461 1819 16519 1853
rect 16553 1819 16614 1853
rect 0 1818 6245 1819
rect 6279 1818 16614 1819
rect 0 1804 16614 1818
rect 29 1795 63 1804
rect 306 1795 340 1804
rect 3158 1795 3192 1804
rect 6522 1795 6556 1804
rect 9374 1795 9408 1804
rect 398 1276 453 1322
rect 1809 1278 1864 1325
rect 2790 1279 2845 1326
rect 4201 1276 4256 1323
rect 5182 1279 5237 1326
rect 6591 1276 6646 1323
rect 7574 1277 7629 1324
rect 8985 1277 9040 1324
rect 9966 1278 10021 1325
rect 11377 1279 11432 1326
rect 12358 1276 12413 1323
rect 13767 1280 13822 1327
rect 14750 1276 14805 1321
rect 16161 1278 16216 1325
rect 0 1261 16614 1276
rect 0 1227 29 1261
rect 63 1227 121 1261
rect 155 1227 213 1261
rect 247 1227 305 1261
rect 339 1227 397 1261
rect 431 1227 489 1261
rect 523 1227 581 1261
rect 615 1227 673 1261
rect 707 1227 765 1261
rect 799 1227 857 1261
rect 891 1227 949 1261
rect 983 1227 1041 1261
rect 1075 1227 1133 1261
rect 1167 1227 1225 1261
rect 1259 1227 1317 1261
rect 1351 1227 1409 1261
rect 1443 1227 1501 1261
rect 1535 1227 1593 1261
rect 1627 1227 1685 1261
rect 1719 1227 1777 1261
rect 1811 1227 1869 1261
rect 1903 1227 1961 1261
rect 1995 1227 2053 1261
rect 2087 1227 2145 1261
rect 2179 1227 2237 1261
rect 2271 1227 2329 1261
rect 2363 1227 2421 1261
rect 2455 1227 2513 1261
rect 2547 1227 2605 1261
rect 2639 1227 2697 1261
rect 2731 1227 2789 1261
rect 2823 1227 2881 1261
rect 2915 1227 2973 1261
rect 3007 1227 3065 1261
rect 3099 1227 3157 1261
rect 3191 1227 3249 1261
rect 3283 1227 3341 1261
rect 3375 1227 3433 1261
rect 3467 1227 3525 1261
rect 3559 1227 3617 1261
rect 3651 1227 3709 1261
rect 3743 1227 3801 1261
rect 3835 1227 3893 1261
rect 3927 1227 3985 1261
rect 4019 1227 4077 1261
rect 4111 1227 4169 1261
rect 4203 1227 4261 1261
rect 4295 1227 4353 1261
rect 4387 1227 4445 1261
rect 4479 1227 4537 1261
rect 4571 1227 4629 1261
rect 4663 1227 4721 1261
rect 4755 1227 4813 1261
rect 4847 1227 4905 1261
rect 4939 1227 4997 1261
rect 5031 1227 5089 1261
rect 5123 1227 5181 1261
rect 5215 1227 5273 1261
rect 5307 1227 5365 1261
rect 5399 1227 5457 1261
rect 5491 1227 5549 1261
rect 5583 1227 5641 1261
rect 5675 1227 6245 1261
rect 6279 1227 6337 1261
rect 6371 1227 6429 1261
rect 6463 1227 6521 1261
rect 6555 1227 6613 1261
rect 6647 1227 6705 1261
rect 6739 1227 6797 1261
rect 6831 1227 6889 1261
rect 6923 1227 6981 1261
rect 7015 1227 7073 1261
rect 7107 1227 7165 1261
rect 7199 1227 7257 1261
rect 7291 1227 7349 1261
rect 7383 1227 7441 1261
rect 7475 1227 7533 1261
rect 7567 1227 7625 1261
rect 7659 1227 7717 1261
rect 7751 1227 7809 1261
rect 7843 1227 7901 1261
rect 7935 1227 7993 1261
rect 8027 1227 8085 1261
rect 8119 1227 8177 1261
rect 8211 1227 8269 1261
rect 8303 1227 8361 1261
rect 8395 1227 8453 1261
rect 8487 1227 8545 1261
rect 8579 1227 8637 1261
rect 8671 1227 8729 1261
rect 8763 1227 8821 1261
rect 8855 1227 8913 1261
rect 8947 1227 9005 1261
rect 9039 1227 9097 1261
rect 9131 1227 9189 1261
rect 9223 1227 9281 1261
rect 9315 1227 9373 1261
rect 9407 1227 9465 1261
rect 9499 1227 9557 1261
rect 9591 1227 9649 1261
rect 9683 1227 9741 1261
rect 9775 1227 9833 1261
rect 9867 1227 9925 1261
rect 9959 1227 10017 1261
rect 10051 1227 10109 1261
rect 10143 1227 10201 1261
rect 10235 1227 10293 1261
rect 10327 1227 10385 1261
rect 10419 1227 10477 1261
rect 10511 1227 10569 1261
rect 10603 1227 10661 1261
rect 10695 1227 10753 1261
rect 10787 1227 10845 1261
rect 10879 1227 10937 1261
rect 10971 1227 11029 1261
rect 11063 1227 11121 1261
rect 11155 1227 11213 1261
rect 11247 1227 11305 1261
rect 11339 1227 11397 1261
rect 11431 1227 11489 1261
rect 11523 1227 11581 1261
rect 11615 1227 11673 1261
rect 11707 1227 11765 1261
rect 11799 1227 11857 1261
rect 11891 1227 12011 1261
rect 12045 1227 12103 1261
rect 12137 1227 12195 1261
rect 12229 1227 12287 1261
rect 12321 1227 12379 1261
rect 12413 1227 12471 1261
rect 12505 1227 12563 1261
rect 12597 1227 12655 1261
rect 12689 1227 12747 1261
rect 12781 1227 12839 1261
rect 12873 1227 12931 1261
rect 12965 1227 13023 1261
rect 13057 1227 13115 1261
rect 13149 1227 13207 1261
rect 13241 1227 13299 1261
rect 13333 1227 13391 1261
rect 13425 1227 13483 1261
rect 13517 1227 13575 1261
rect 13609 1227 13667 1261
rect 13701 1227 13759 1261
rect 13793 1227 13851 1261
rect 13885 1227 13943 1261
rect 13977 1227 14035 1261
rect 14069 1227 14127 1261
rect 14161 1227 14219 1261
rect 14253 1227 14311 1261
rect 14345 1227 14403 1261
rect 14437 1227 14495 1261
rect 14529 1227 14587 1261
rect 14621 1227 14679 1261
rect 14713 1227 14771 1261
rect 14805 1227 14863 1261
rect 14897 1227 14955 1261
rect 14989 1227 15047 1261
rect 15081 1227 15139 1261
rect 15173 1227 15231 1261
rect 15265 1227 15323 1261
rect 15357 1227 15415 1261
rect 15449 1227 15507 1261
rect 15541 1227 15599 1261
rect 15633 1227 15691 1261
rect 15725 1227 15783 1261
rect 15817 1227 15875 1261
rect 15909 1227 15967 1261
rect 16001 1227 16059 1261
rect 16093 1227 16151 1261
rect 16185 1227 16243 1261
rect 16277 1227 16335 1261
rect 16369 1227 16427 1261
rect 16461 1227 16519 1261
rect 16553 1227 16614 1261
rect 16237 1165 16303 1173
rect 0 1131 29 1165
rect 63 1131 121 1165
rect 155 1131 213 1165
rect 247 1131 305 1165
rect 339 1131 397 1165
rect 431 1131 489 1165
rect 523 1131 581 1165
rect 615 1131 673 1165
rect 707 1131 765 1165
rect 799 1131 857 1165
rect 891 1131 949 1165
rect 983 1131 1041 1165
rect 1075 1131 1133 1165
rect 1167 1131 1225 1165
rect 1259 1131 1317 1165
rect 1351 1131 1409 1165
rect 1443 1131 1501 1165
rect 1535 1131 1593 1165
rect 1627 1131 1685 1165
rect 1719 1131 1777 1165
rect 1811 1158 2053 1165
rect 1811 1132 1901 1158
rect 1811 1131 1869 1132
rect 0 1126 1901 1131
rect 1885 1124 1901 1126
rect 1935 1138 2053 1158
rect 1935 1131 1961 1138
rect 1995 1131 2053 1138
rect 2087 1131 2145 1165
rect 2179 1131 2237 1165
rect 2271 1131 2329 1165
rect 2363 1131 2421 1165
rect 2455 1131 2513 1165
rect 2547 1131 2605 1165
rect 2639 1131 2697 1165
rect 2731 1131 2789 1165
rect 2823 1131 2881 1165
rect 2915 1131 2973 1165
rect 3007 1131 3065 1165
rect 3099 1131 3157 1165
rect 3191 1131 3249 1165
rect 3283 1131 3341 1165
rect 3375 1131 3433 1165
rect 3467 1131 3525 1165
rect 3559 1131 3617 1165
rect 3651 1131 3709 1165
rect 3743 1131 3801 1165
rect 3835 1131 3893 1165
rect 3927 1131 3985 1165
rect 4019 1131 4077 1165
rect 4111 1131 4169 1165
rect 4203 1157 4445 1165
rect 4203 1131 4293 1157
rect 1935 1126 4293 1131
rect 1935 1124 1951 1126
rect 4261 1123 4293 1126
rect 4327 1134 4445 1157
rect 4327 1131 4353 1134
rect 4387 1131 4445 1134
rect 4479 1131 4537 1165
rect 4571 1131 4629 1165
rect 4663 1131 4721 1165
rect 4755 1131 4813 1165
rect 4847 1131 4905 1165
rect 4939 1131 4997 1165
rect 5031 1131 5089 1165
rect 5123 1131 5181 1165
rect 5215 1131 5273 1165
rect 5307 1131 5365 1165
rect 5399 1131 5457 1165
rect 5491 1131 5549 1165
rect 5583 1131 5641 1165
rect 5675 1131 5733 1165
rect 5767 1131 5825 1165
rect 5859 1131 5917 1165
rect 5951 1131 6009 1165
rect 6043 1131 6101 1165
rect 6135 1131 6193 1165
rect 6227 1131 6285 1165
rect 6319 1131 6377 1165
rect 6411 1131 6469 1165
rect 6503 1131 6561 1165
rect 6595 1157 6837 1165
rect 6595 1135 6685 1157
rect 6595 1131 6653 1135
rect 4327 1126 6685 1131
rect 4327 1123 4343 1126
rect 6669 1123 6685 1126
rect 6719 1135 6837 1157
rect 6719 1131 6745 1135
rect 6779 1131 6837 1135
rect 6871 1131 6929 1165
rect 6963 1131 7021 1165
rect 7055 1131 7113 1165
rect 7147 1131 7205 1165
rect 7239 1131 7297 1165
rect 7331 1131 7389 1165
rect 7423 1131 7481 1165
rect 7515 1131 7573 1165
rect 7607 1131 7665 1165
rect 7699 1131 7757 1165
rect 7791 1131 7849 1165
rect 7883 1131 7941 1165
rect 7975 1131 8033 1165
rect 8067 1131 8125 1165
rect 8159 1131 8217 1165
rect 8251 1131 8309 1165
rect 8343 1131 8401 1165
rect 8435 1131 8493 1165
rect 8527 1131 8585 1165
rect 8619 1131 8677 1165
rect 8711 1131 8769 1165
rect 8803 1131 8861 1165
rect 8895 1131 8953 1165
rect 8987 1158 9229 1165
rect 8987 1131 9077 1158
rect 6719 1126 9077 1131
rect 6719 1123 6735 1126
rect 9061 1124 9077 1126
rect 9111 1131 9229 1158
rect 9263 1131 9321 1165
rect 9355 1131 9413 1165
rect 9447 1131 9505 1165
rect 9539 1131 9597 1165
rect 9631 1131 9689 1165
rect 9723 1131 9781 1165
rect 9815 1131 9873 1165
rect 9907 1131 9965 1165
rect 9999 1131 10057 1165
rect 10091 1131 10149 1165
rect 10183 1131 10241 1165
rect 10275 1131 10333 1165
rect 10367 1131 10425 1165
rect 10459 1131 10517 1165
rect 10551 1131 10609 1165
rect 10643 1131 10701 1165
rect 10735 1131 10793 1165
rect 10827 1131 10885 1165
rect 10919 1131 10977 1165
rect 11011 1131 11069 1165
rect 11103 1131 11161 1165
rect 11195 1131 11253 1165
rect 11287 1131 11345 1165
rect 11379 1158 11621 1165
rect 11379 1135 11469 1158
rect 11379 1131 11437 1135
rect 9111 1126 11469 1131
rect 9111 1124 9127 1126
rect 11453 1124 11469 1126
rect 11503 1135 11621 1158
rect 11503 1131 11529 1135
rect 11563 1131 11621 1135
rect 11655 1131 11713 1165
rect 11747 1131 11805 1165
rect 11839 1131 11897 1165
rect 11931 1131 11989 1165
rect 12023 1131 12081 1165
rect 12115 1131 12173 1165
rect 12207 1131 12265 1165
rect 12299 1131 12357 1165
rect 12391 1131 12449 1165
rect 12483 1131 12541 1165
rect 12575 1131 12633 1165
rect 12667 1131 12725 1165
rect 12759 1131 12817 1165
rect 12851 1131 12909 1165
rect 12943 1131 13001 1165
rect 13035 1131 13093 1165
rect 13127 1131 13185 1165
rect 13219 1131 13277 1165
rect 13311 1131 13369 1165
rect 13403 1131 13461 1165
rect 13495 1131 13553 1165
rect 13587 1131 13645 1165
rect 13679 1131 13737 1165
rect 13771 1157 14013 1165
rect 13771 1131 13861 1157
rect 11503 1126 13861 1131
rect 11503 1124 11519 1126
rect 13828 1123 13861 1126
rect 13895 1131 14013 1157
rect 14047 1131 14105 1165
rect 14139 1131 14197 1165
rect 14231 1131 14289 1165
rect 14323 1131 14381 1165
rect 14415 1131 14473 1165
rect 14507 1131 14565 1165
rect 14599 1131 14657 1165
rect 14691 1131 14749 1165
rect 14783 1131 14841 1165
rect 14875 1131 14933 1165
rect 14967 1131 15025 1165
rect 15059 1131 15117 1165
rect 15151 1131 15209 1165
rect 15243 1131 15301 1165
rect 15335 1131 15393 1165
rect 15427 1131 15485 1165
rect 15519 1131 15577 1165
rect 15611 1131 15669 1165
rect 15703 1131 15761 1165
rect 15795 1131 15853 1165
rect 15887 1131 15945 1165
rect 15979 1131 16037 1165
rect 16071 1131 16129 1165
rect 16163 1157 16405 1165
rect 16163 1131 16253 1157
rect 13895 1126 16253 1131
rect 13895 1123 13976 1126
rect 4261 1121 4336 1123
rect 13828 1121 13976 1123
rect 16237 1123 16253 1126
rect 16287 1135 16405 1157
rect 16287 1131 16313 1135
rect 16347 1131 16405 1135
rect 16439 1131 16497 1165
rect 16531 1131 16589 1165
rect 16623 1131 16681 1165
rect 16715 1131 16744 1165
rect 16287 1126 16744 1131
rect 16287 1123 16303 1126
rect 16583 1125 16744 1126
rect 16237 1107 16303 1123
rect 0 573 16614 578
rect 0 539 29 573
rect 63 539 121 573
rect 155 539 213 573
rect 247 539 305 573
rect 339 539 397 573
rect 431 539 489 573
rect 523 539 581 573
rect 615 539 673 573
rect 707 539 765 573
rect 799 539 857 573
rect 891 539 949 573
rect 983 539 1041 573
rect 1075 539 1133 573
rect 1167 539 1225 573
rect 1259 539 1317 573
rect 1351 539 1409 573
rect 1443 539 1501 573
rect 1535 539 1593 573
rect 1627 539 1685 573
rect 1719 539 1777 573
rect 1811 539 1869 573
rect 1903 539 1961 573
rect 1995 539 2053 573
rect 2087 539 2145 573
rect 2179 539 2237 573
rect 2271 539 2329 573
rect 2363 539 2421 573
rect 2455 539 2513 573
rect 2547 539 2605 573
rect 2639 539 2697 573
rect 2731 539 2789 573
rect 2823 539 2881 573
rect 2915 539 2973 573
rect 3007 539 3065 573
rect 3099 539 3157 573
rect 3191 539 3249 573
rect 3283 539 3341 573
rect 3375 539 3433 573
rect 3467 539 3525 573
rect 3559 539 3617 573
rect 3651 539 3709 573
rect 3743 539 3801 573
rect 3835 539 3893 573
rect 3927 539 3985 573
rect 4019 539 4077 573
rect 4111 539 4169 573
rect 4203 539 4261 573
rect 4295 539 4353 573
rect 4387 539 4445 573
rect 4479 539 4537 573
rect 4571 539 4629 573
rect 4663 539 4721 573
rect 4755 539 4813 573
rect 4847 539 4905 573
rect 4939 539 4997 573
rect 5031 539 5089 573
rect 5123 539 5181 573
rect 5215 539 5273 573
rect 5307 539 5365 573
rect 5399 539 5457 573
rect 5491 539 5549 573
rect 5583 539 5641 573
rect 5675 539 5733 573
rect 5767 539 5825 573
rect 5859 539 5917 573
rect 5951 539 6009 573
rect 6043 539 6101 573
rect 6135 539 6193 573
rect 6227 539 6285 573
rect 6319 539 6377 573
rect 6411 539 6469 573
rect 6503 539 6561 573
rect 6595 539 6653 573
rect 6687 539 6745 573
rect 6779 539 6837 573
rect 6871 539 6929 573
rect 6963 539 7021 573
rect 7055 539 7113 573
rect 7147 539 7205 573
rect 7239 539 7297 573
rect 7331 539 7389 573
rect 7423 539 7481 573
rect 7515 539 7573 573
rect 7607 539 7665 573
rect 7699 539 7757 573
rect 7791 539 7849 573
rect 7883 539 7941 573
rect 7975 539 8033 573
rect 8067 539 8125 573
rect 8159 539 8217 573
rect 8251 539 8309 573
rect 8343 539 8401 573
rect 8435 539 8493 573
rect 8527 539 8585 573
rect 8619 539 8677 573
rect 8711 539 8769 573
rect 8803 539 8861 573
rect 8895 539 8953 573
rect 8987 539 9045 573
rect 9079 539 9137 573
rect 9171 539 9229 573
rect 9263 539 9321 573
rect 9355 539 9413 573
rect 9447 539 9505 573
rect 9539 539 9597 573
rect 9631 539 9689 573
rect 9723 539 9781 573
rect 9815 539 9873 573
rect 9907 539 9965 573
rect 9999 539 10057 573
rect 10091 539 10149 573
rect 10183 539 10241 573
rect 10275 539 10333 573
rect 10367 539 10425 573
rect 10459 539 10517 573
rect 10551 539 10609 573
rect 10643 539 10701 573
rect 10735 539 10793 573
rect 10827 539 10885 573
rect 10919 539 10977 573
rect 11011 539 11069 573
rect 11103 539 11161 573
rect 11195 539 11253 573
rect 11287 539 11345 573
rect 11379 539 11437 573
rect 11471 539 11529 573
rect 11563 539 11621 573
rect 11655 539 11713 573
rect 11747 539 11805 573
rect 11839 539 11897 573
rect 11931 539 11989 573
rect 12023 539 12081 573
rect 12115 539 12173 573
rect 12207 539 12265 573
rect 12299 539 12357 573
rect 12391 539 12449 573
rect 12483 539 12541 573
rect 12575 539 12633 573
rect 12667 539 12725 573
rect 12759 539 12817 573
rect 12851 539 12909 573
rect 12943 539 13001 573
rect 13035 539 13093 573
rect 13127 539 13185 573
rect 13219 539 13277 573
rect 13311 539 13369 573
rect 13403 539 13461 573
rect 13495 539 13553 573
rect 13587 539 13645 573
rect 13679 539 13737 573
rect 13771 539 13829 573
rect 13863 539 13921 573
rect 13955 539 14013 573
rect 14047 539 14105 573
rect 14139 539 14197 573
rect 14231 539 14289 573
rect 14323 539 14381 573
rect 14415 539 14473 573
rect 14507 539 14565 573
rect 14599 539 14657 573
rect 14691 539 14749 573
rect 14783 539 14841 573
rect 14875 539 14933 573
rect 14967 539 15025 573
rect 15059 539 15117 573
rect 15151 539 15209 573
rect 15243 539 15301 573
rect 15335 539 15393 573
rect 15427 539 15485 573
rect 15519 539 15577 573
rect 15611 539 15669 573
rect 15703 539 15761 573
rect 15795 539 15853 573
rect 15887 539 15945 573
rect 15979 539 16037 573
rect 16071 539 16129 573
rect 16163 539 16221 573
rect 16255 539 16313 573
rect 16347 539 16405 573
rect 16439 539 16497 573
rect 16531 539 16589 573
rect 16623 539 16681 573
rect 16715 539 16744 573
rect 0 476 571 477
rect 0 442 29 476
rect 63 442 121 476
rect 155 442 213 476
rect 247 442 305 476
rect 339 442 394 476
rect 428 442 496 476
rect 530 442 581 476
rect 615 442 673 476
rect 707 442 765 476
rect 799 442 857 476
rect 891 442 949 476
rect 983 442 1041 476
rect 1075 442 1133 476
rect 1167 442 1225 476
rect 1259 442 1317 476
rect 1351 442 1409 476
rect 1443 442 1501 476
rect 1535 472 1777 476
rect 1535 442 1607 472
rect 0 438 1607 442
rect 1641 442 1777 472
rect 1811 442 1869 476
rect 1903 442 1961 476
rect 1995 442 2053 476
rect 2087 442 2145 476
rect 2179 442 2237 476
rect 2271 442 2329 476
rect 2363 442 2421 476
rect 2455 442 2513 476
rect 2547 442 2605 476
rect 2639 442 2697 476
rect 2731 442 2791 476
rect 2825 442 2882 476
rect 2916 442 2973 476
rect 3007 442 3065 476
rect 3099 442 3157 476
rect 3191 442 3249 476
rect 3283 442 3341 476
rect 3375 442 3433 476
rect 3467 442 3525 476
rect 3559 442 3617 476
rect 3651 442 3709 476
rect 3743 442 3801 476
rect 3835 442 3893 476
rect 3927 472 4169 476
rect 3927 442 3999 472
rect 1641 438 3999 442
rect 4033 442 4169 472
rect 4203 442 4261 476
rect 4295 442 4353 476
rect 4387 442 4445 476
rect 4479 442 4537 476
rect 4571 442 4629 476
rect 4663 442 4721 476
rect 4755 442 4813 476
rect 4847 442 4905 476
rect 4939 442 4997 476
rect 5031 442 5089 476
rect 5123 442 5179 476
rect 5213 442 5273 476
rect 5307 442 5365 476
rect 5399 442 5457 476
rect 5491 442 5549 476
rect 5583 442 5641 476
rect 5675 442 5733 476
rect 5767 442 5825 476
rect 5859 442 5917 476
rect 5951 442 6009 476
rect 6043 442 6101 476
rect 6135 442 6193 476
rect 6227 442 6285 476
rect 6319 472 6561 476
rect 6319 442 6391 472
rect 4033 438 6391 442
rect 6425 442 6561 472
rect 6595 442 6653 476
rect 6687 442 6745 476
rect 6779 442 6837 476
rect 6871 442 6929 476
rect 6963 442 7021 476
rect 7055 442 7113 476
rect 7147 442 7205 476
rect 7239 442 7297 476
rect 7331 442 7389 476
rect 7423 442 7481 476
rect 7515 442 7574 476
rect 7608 442 7665 476
rect 7699 442 7757 476
rect 7791 442 7849 476
rect 7883 442 7941 476
rect 7975 442 8033 476
rect 8067 442 8125 476
rect 8159 442 8217 476
rect 8251 442 8309 476
rect 8343 442 8401 476
rect 8435 442 8493 476
rect 8527 442 8585 476
rect 8619 442 8677 476
rect 8711 472 8953 476
rect 8711 442 8783 472
rect 6425 438 8783 442
rect 8817 442 8953 472
rect 8987 442 9045 476
rect 9079 442 9137 476
rect 9171 442 9229 476
rect 9263 442 9321 476
rect 9355 442 9413 476
rect 9447 442 9505 476
rect 9539 442 9597 476
rect 9631 442 9689 476
rect 9723 442 9781 476
rect 9815 442 9873 476
rect 9907 442 9963 476
rect 9997 442 10058 476
rect 10092 442 10149 476
rect 10183 442 10241 476
rect 10275 442 10333 476
rect 10367 442 10425 476
rect 10459 442 10517 476
rect 10551 442 10609 476
rect 10643 442 10701 476
rect 10735 442 10793 476
rect 10827 442 10885 476
rect 10919 442 10977 476
rect 11011 442 11069 476
rect 11103 472 11345 476
rect 11103 442 11175 472
rect 8817 438 11175 442
rect 11209 442 11345 472
rect 11379 442 11437 476
rect 11471 442 11529 476
rect 11563 442 11621 476
rect 11655 442 11713 476
rect 11747 442 11805 476
rect 11839 442 11897 476
rect 11931 442 11989 476
rect 12023 442 12081 476
rect 12115 442 12173 476
rect 12207 442 12265 476
rect 12299 442 12357 476
rect 12391 442 12448 476
rect 12482 442 12541 476
rect 12575 442 12633 476
rect 12667 442 12725 476
rect 12759 442 12817 476
rect 12851 442 12909 476
rect 12943 442 13001 476
rect 13035 442 13093 476
rect 13127 442 13185 476
rect 13219 442 13277 476
rect 13311 442 13369 476
rect 13403 442 13461 476
rect 13495 472 13737 476
rect 13495 442 13567 472
rect 11209 438 13567 442
rect 13601 442 13737 472
rect 13771 442 13829 476
rect 13863 442 13921 476
rect 13955 442 14013 476
rect 14047 442 14105 476
rect 14139 442 14197 476
rect 14231 442 14289 476
rect 14323 442 14381 476
rect 14415 442 14473 476
rect 14507 442 14565 476
rect 14599 442 14657 476
rect 14691 442 14748 476
rect 14782 442 14842 476
rect 14876 442 14933 476
rect 14967 442 15025 476
rect 15059 442 15117 476
rect 15151 442 15209 476
rect 15243 442 15301 476
rect 15335 442 15393 476
rect 15427 442 15485 476
rect 15519 442 15577 476
rect 15611 442 15669 476
rect 15703 442 15761 476
rect 15795 442 15853 476
rect 15887 469 16129 476
rect 15887 442 15959 469
rect 13601 438 15959 442
rect 0 437 1591 438
rect 1657 437 8767 438
rect 8833 437 11159 438
rect 11225 437 15959 438
rect 7683 436 7727 437
rect 8745 418 8749 437
rect 15943 435 15959 437
rect 15993 442 16129 469
rect 16163 442 16221 476
rect 16255 442 16313 476
rect 16347 442 16405 476
rect 16439 442 16497 476
rect 16531 442 16589 476
rect 16623 448 16681 476
rect 16715 448 16744 476
rect 15993 437 16614 442
rect 15993 435 16009 437
rect 15943 419 16009 435
rect 16561 -111 16744 -104
rect 0 -116 16744 -111
rect 0 -150 29 -116
rect 63 -150 121 -116
rect 155 -150 213 -116
rect 247 -150 305 -116
rect 339 -150 397 -116
rect 431 -150 489 -116
rect 523 -150 581 -116
rect 615 -150 673 -116
rect 707 -150 765 -116
rect 799 -150 857 -116
rect 891 -150 949 -116
rect 983 -150 1041 -116
rect 1075 -150 1133 -116
rect 1167 -150 1225 -116
rect 1259 -150 1317 -116
rect 1351 -150 1409 -116
rect 1443 -150 1501 -116
rect 1535 -150 1593 -116
rect 1627 -150 1685 -116
rect 1719 -150 1777 -116
rect 1811 -150 1869 -116
rect 1903 -150 1961 -116
rect 1995 -150 2053 -116
rect 2087 -150 2145 -116
rect 2179 -150 2237 -116
rect 2271 -150 2329 -116
rect 2363 -150 2421 -116
rect 2455 -150 2513 -116
rect 2547 -150 2605 -116
rect 2639 -150 2697 -116
rect 2731 -150 2789 -116
rect 2823 -150 2881 -116
rect 2915 -150 2973 -116
rect 3007 -150 3065 -116
rect 3099 -150 3157 -116
rect 3191 -150 3249 -116
rect 3283 -150 3341 -116
rect 3375 -150 3433 -116
rect 3467 -150 3525 -116
rect 3559 -150 3617 -116
rect 3651 -150 3709 -116
rect 3743 -150 3801 -116
rect 3835 -150 3893 -116
rect 3927 -150 3985 -116
rect 4019 -150 4077 -116
rect 4111 -150 4169 -116
rect 4203 -150 4261 -116
rect 4295 -150 4353 -116
rect 4387 -150 4445 -116
rect 4479 -150 4537 -116
rect 4571 -150 4629 -116
rect 4663 -150 4721 -116
rect 4755 -150 4813 -116
rect 4847 -150 4905 -116
rect 4939 -150 4997 -116
rect 5031 -150 5089 -116
rect 5123 -150 5181 -116
rect 5215 -150 5273 -116
rect 5307 -150 5365 -116
rect 5399 -150 5457 -116
rect 5491 -150 5549 -116
rect 5583 -150 5641 -116
rect 5675 -150 5733 -116
rect 5767 -150 5825 -116
rect 5859 -150 5917 -116
rect 5951 -150 6009 -116
rect 6043 -150 6101 -116
rect 6135 -150 6193 -116
rect 6227 -150 6285 -116
rect 6319 -150 6377 -116
rect 6411 -150 6469 -116
rect 6503 -150 6561 -116
rect 6595 -150 6653 -116
rect 6687 -150 6745 -116
rect 6779 -150 6837 -116
rect 6871 -150 6929 -116
rect 6963 -150 7021 -116
rect 7055 -150 7113 -116
rect 7147 -150 7205 -116
rect 7239 -150 7297 -116
rect 7331 -150 7389 -116
rect 7423 -150 7481 -116
rect 7515 -150 7573 -116
rect 7607 -150 7665 -116
rect 7699 -150 7757 -116
rect 7791 -150 7849 -116
rect 7883 -150 7941 -116
rect 7975 -150 8033 -116
rect 8067 -150 8125 -116
rect 8159 -150 8217 -116
rect 8251 -150 8309 -116
rect 8343 -150 8401 -116
rect 8435 -150 8493 -116
rect 8527 -150 8585 -116
rect 8619 -150 8677 -116
rect 8711 -150 8769 -116
rect 8803 -150 8861 -116
rect 8895 -150 8953 -116
rect 8987 -150 9045 -116
rect 9079 -150 9137 -116
rect 9171 -150 9229 -116
rect 9263 -150 9321 -116
rect 9355 -150 9413 -116
rect 9447 -150 9505 -116
rect 9539 -150 9597 -116
rect 9631 -150 9689 -116
rect 9723 -150 9781 -116
rect 9815 -150 9873 -116
rect 9907 -150 9965 -116
rect 9999 -150 10057 -116
rect 10091 -150 10149 -116
rect 10183 -150 10241 -116
rect 10275 -150 10333 -116
rect 10367 -150 10425 -116
rect 10459 -150 10517 -116
rect 10551 -150 10609 -116
rect 10643 -150 10701 -116
rect 10735 -150 10793 -116
rect 10827 -150 10885 -116
rect 10919 -150 10977 -116
rect 11011 -150 11069 -116
rect 11103 -150 11161 -116
rect 11195 -150 11253 -116
rect 11287 -150 11345 -116
rect 11379 -150 11437 -116
rect 11471 -150 11529 -116
rect 11563 -150 11621 -116
rect 11655 -150 11713 -116
rect 11747 -150 11805 -116
rect 11839 -150 11897 -116
rect 11931 -150 11989 -116
rect 12023 -150 12081 -116
rect 12115 -150 12173 -116
rect 12207 -150 12265 -116
rect 12299 -150 12357 -116
rect 12391 -150 12449 -116
rect 12483 -150 12541 -116
rect 12575 -150 12633 -116
rect 12667 -150 12725 -116
rect 12759 -150 12817 -116
rect 12851 -150 12909 -116
rect 12943 -150 13001 -116
rect 13035 -150 13093 -116
rect 13127 -150 13185 -116
rect 13219 -150 13277 -116
rect 13311 -150 13369 -116
rect 13403 -150 13461 -116
rect 13495 -150 13553 -116
rect 13587 -150 13645 -116
rect 13679 -150 13737 -116
rect 13771 -150 13829 -116
rect 13863 -150 13921 -116
rect 13955 -150 14013 -116
rect 14047 -150 14105 -116
rect 14139 -150 14197 -116
rect 14231 -150 14289 -116
rect 14323 -150 14381 -116
rect 14415 -150 14473 -116
rect 14507 -150 14565 -116
rect 14599 -150 14657 -116
rect 14691 -150 14749 -116
rect 14783 -150 14841 -116
rect 14875 -150 14933 -116
rect 14967 -150 15025 -116
rect 15059 -150 15117 -116
rect 15151 -150 15209 -116
rect 15243 -150 15301 -116
rect 15335 -150 15393 -116
rect 15427 -150 15485 -116
rect 15519 -150 15577 -116
rect 15611 -150 15669 -116
rect 15703 -150 15761 -116
rect 15795 -150 15853 -116
rect 15887 -150 15945 -116
rect 15979 -150 16037 -116
rect 16071 -150 16129 -116
rect 16163 -150 16221 -116
rect 16255 -150 16313 -116
rect 16347 -150 16405 -116
rect 16439 -150 16497 -116
rect 16531 -150 16589 -116
rect 16623 -150 16681 -116
rect 16715 -150 16744 -116
<< viali >>
rect 39 2641 73 2675
rect 2876 2630 2910 2664
rect 4423 2624 4457 2658
rect 7176 2632 7210 2666
rect 484 1573 518 1607
rect 656 1557 690 1591
rect 1566 1558 1600 1592
rect 1746 1573 1780 1607
rect 2877 1572 2911 1606
rect 3048 1556 3082 1590
rect 3958 1557 3992 1591
rect 4138 1573 4172 1607
rect 5269 1572 5303 1606
rect 5439 1557 5473 1591
rect 6348 1557 6382 1591
rect 6529 1574 6563 1608
rect 7661 1573 7695 1607
rect 7832 1557 7866 1591
rect 8742 1558 8776 1592
rect 8922 1574 8956 1608
rect 10052 1572 10086 1606
rect 10223 1558 10257 1592
rect 11134 1557 11168 1591
rect 11315 1574 11349 1608
rect 12444 1571 12478 1605
rect 12615 1558 12649 1592
rect 13523 1557 13557 1591
rect 13704 1574 13738 1608
rect 14836 1572 14870 1606
rect 15008 1558 15042 1592
rect 15918 1558 15952 1592
rect 16099 1574 16133 1608
rect 28 1372 62 1406
rect 2204 1370 2238 1404
rect 2420 1372 2454 1406
rect 4598 1370 4632 1404
rect 4812 1372 4846 1406
rect 6988 1372 7022 1406
rect 7204 1372 7238 1406
rect 9380 1370 9414 1404
rect 9595 1373 9629 1407
rect 11772 1372 11806 1406
rect 11987 1372 12021 1406
rect 14164 1370 14198 1404
rect 14380 1373 14414 1407
rect 16556 1372 16590 1406
rect 2334 1000 2368 1034
rect 4726 1000 4760 1034
rect 7118 1000 7152 1034
rect 9510 1000 9544 1034
rect 11902 1000 11936 1034
rect 14294 1000 14328 1034
rect 16686 1000 16720 1034
rect 2051 921 2085 955
rect 4443 922 4477 956
rect 6834 922 6868 956
rect 9227 923 9261 957
rect 11618 922 11652 956
rect 14011 921 14045 955
rect 16404 923 16438 957
rect 26 825 60 859
rect 366 849 400 883
rect 2418 825 2452 859
rect 2758 849 2792 883
rect 4810 825 4844 859
rect 5150 850 5184 884
rect 7202 825 7236 859
rect 7542 850 7576 884
rect 9593 826 9627 860
rect 9934 849 9968 883
rect 11985 825 12019 859
rect 12326 850 12360 884
rect 14378 826 14412 860
rect 14719 849 14753 883
rect 26 308 60 342
rect 2418 308 2452 342
rect 4811 308 4845 342
rect 7202 308 7236 342
rect 9594 307 9628 341
rect 11987 309 12021 343
rect 14378 309 14412 343
rect 306 242 340 276
rect 2698 242 2732 276
rect 5089 242 5123 276
rect 7482 242 7516 276
rect 9874 242 9908 276
rect 12265 243 12299 277
rect 14658 242 14692 276
rect 2314 171 2348 205
rect 4708 171 4742 205
rect 7098 173 7132 207
rect 9490 171 9524 205
rect 11882 173 11916 207
rect 14274 171 14308 205
rect 16666 173 16700 207
rect 502 114 536 148
rect 1968 115 2002 149
rect 2891 116 2925 150
rect 4360 115 4394 149
rect 5284 116 5318 150
rect 6751 116 6785 150
rect 7677 116 7711 150
rect 9144 115 9178 149
rect 10068 116 10102 150
rect 11535 115 11569 149
rect 12461 116 12495 150
rect 13928 115 13962 149
rect 14852 116 14886 150
rect 16321 115 16355 149
<< metal1 >>
rect 723 3435 775 3441
rect 723 3377 775 3383
rect -126 2990 16861 3002
rect -144 2980 16861 2990
rect -144 2978 1265 2980
rect -144 2976 255 2978
rect -144 2924 53 2976
rect 105 2926 255 2976
rect 307 2976 864 2978
rect 307 2926 466 2976
rect 105 2924 466 2926
rect 518 2924 656 2976
rect 708 2926 864 2976
rect 916 2926 1066 2978
rect 1118 2928 1265 2978
rect 1317 2979 2152 2980
rect 1317 2977 1661 2979
rect 1317 2928 1460 2977
rect 1118 2926 1460 2928
rect 708 2925 1460 2926
rect 1512 2927 1661 2977
rect 1713 2977 2152 2979
rect 1713 2927 1878 2977
rect 1512 2925 1878 2927
rect 1930 2928 2152 2977
rect 2204 2976 16861 2980
rect 2204 2973 2652 2976
rect 2204 2928 2429 2973
rect 1930 2925 2429 2928
rect 708 2924 2429 2925
rect -144 2921 2429 2924
rect 2481 2924 2652 2973
rect 2704 2975 16861 2976
rect 2704 2924 2884 2975
rect 2481 2923 2884 2924
rect 2936 2974 5903 2975
rect 2936 2973 5028 2974
rect 2936 2972 4828 2973
rect 2936 2923 4520 2972
rect 2481 2921 4520 2923
rect -144 2920 4520 2921
rect 4572 2921 4828 2972
rect 4880 2922 5028 2973
rect 5080 2973 5701 2974
rect 5080 2922 5247 2973
rect 4880 2921 5247 2922
rect 5299 2972 5701 2973
rect 5299 2921 5493 2972
rect 4572 2920 5493 2921
rect 5545 2922 5701 2972
rect 5753 2923 5903 2974
rect 5955 2974 16861 2975
rect 5955 2923 6096 2974
rect 5753 2922 6096 2923
rect 6148 2973 16861 2974
rect 6148 2922 6468 2973
rect 5545 2921 6468 2922
rect 6520 2971 7220 2973
rect 6520 2921 6657 2971
rect 5545 2920 6657 2921
rect -144 2919 6657 2920
rect 6709 2919 6947 2971
rect 6999 2921 7220 2971
rect 7272 2921 16861 2973
rect 6999 2919 16861 2921
rect -144 2906 16861 2919
rect -144 2904 -120 2906
rect -126 2722 -34 2756
rect -68 2681 -34 2722
rect 27 2681 85 2687
rect -68 2675 85 2681
rect -68 2647 39 2675
rect 26 2641 39 2647
rect 73 2641 85 2675
rect 26 2631 85 2641
rect 2860 2622 2866 2674
rect 2918 2622 2924 2674
rect 7164 2668 7216 2674
rect 7421 2668 7427 2674
rect 7164 2666 7427 2668
rect 4411 2658 4469 2664
rect 4411 2656 4423 2658
rect 4270 2624 4423 2656
rect 4457 2624 4469 2658
rect 4270 2560 4302 2624
rect 4411 2618 4469 2624
rect 7164 2632 7176 2666
rect 7210 2632 7427 2666
rect 7164 2626 7427 2632
rect 7164 2620 7216 2626
rect 7421 2622 7427 2626
rect 7479 2622 7485 2674
rect -126 2526 4302 2560
rect -126 2448 16861 2458
rect -126 2441 16876 2448
rect -126 2437 1390 2441
rect -126 2385 1171 2437
rect 1223 2389 1390 2437
rect 1442 2389 1673 2441
rect 1725 2389 1882 2441
rect 1934 2440 16876 2441
rect 1934 2439 4477 2440
rect 1934 2389 2153 2439
rect 1223 2387 2153 2389
rect 2205 2437 4477 2439
rect 2205 2387 4228 2437
rect 1223 2385 4228 2387
rect 4280 2388 4477 2437
rect 4529 2439 16876 2440
rect 4529 2437 7226 2439
rect 4529 2432 7022 2437
rect 4529 2426 5075 2432
rect 4529 2388 4821 2426
rect 4280 2385 4821 2388
rect -126 2374 4821 2385
rect 4873 2380 5075 2426
rect 5127 2380 5304 2432
rect 5356 2385 7022 2432
rect 7074 2387 7226 2437
rect 7278 2437 16876 2439
rect 7278 2387 7549 2437
rect 7074 2385 7549 2387
rect 7601 2385 16876 2437
rect 5356 2380 16876 2385
rect 4873 2374 16876 2380
rect -126 2362 16876 2374
rect 1018 2294 1024 2303
rect 95 2260 1024 2294
rect 1018 2250 1024 2260
rect 1077 2294 1083 2303
rect 2860 2294 2866 2302
rect 1077 2260 2866 2294
rect 1077 2250 1083 2260
rect 2860 2250 2866 2260
rect 2918 2294 2924 2302
rect 3412 2294 3418 2309
rect 2918 2260 3418 2294
rect 2918 2250 2924 2260
rect 3412 2256 3418 2260
rect 3471 2294 3477 2309
rect 5803 2294 5809 2309
rect 3471 2260 5809 2294
rect 3471 2256 3477 2260
rect 3412 2255 3477 2256
rect 5803 2256 5809 2260
rect 5862 2294 5868 2309
rect 8194 2294 8200 2309
rect 5862 2260 8200 2294
rect 5862 2256 5868 2260
rect 7416 2259 7533 2260
rect 5803 2255 5868 2256
rect 8194 2256 8200 2260
rect 8253 2294 8259 2309
rect 10586 2294 10592 2309
rect 8253 2260 10592 2294
rect 8253 2256 8259 2260
rect 8194 2255 8259 2256
rect 10586 2256 10592 2260
rect 10645 2294 10651 2309
rect 12977 2294 12983 2309
rect 10645 2260 12983 2294
rect 10645 2256 10651 2260
rect 10586 2255 10651 2256
rect 12977 2256 12983 2260
rect 13036 2294 13042 2309
rect 15370 2294 15376 2309
rect 13036 2260 15376 2294
rect 13036 2256 13042 2260
rect 12977 2255 13042 2256
rect 15370 2256 15376 2260
rect 15429 2294 15435 2309
rect 15429 2260 16861 2294
rect 15429 2256 15435 2260
rect 15370 2255 15435 2256
rect 1018 2249 1083 2250
rect 95 2186 16861 2188
rect 95 2154 16876 2186
rect 7419 2153 7528 2154
rect 467 2082 474 2091
rect 95 2048 474 2082
rect 467 2039 474 2048
rect 526 2082 533 2091
rect 1729 2082 1736 2091
rect 526 2048 1736 2082
rect 526 2039 533 2048
rect 1729 2039 1736 2048
rect 1788 2082 1795 2091
rect 2860 2082 2867 2090
rect 1788 2048 2867 2082
rect 1788 2039 1795 2048
rect 2860 2038 2867 2048
rect 2919 2082 2926 2090
rect 4121 2082 4128 2091
rect 2919 2048 4128 2082
rect 2919 2038 2926 2048
rect 4121 2039 4128 2048
rect 4180 2082 4187 2091
rect 5252 2082 5259 2090
rect 4180 2048 5259 2082
rect 4180 2039 4187 2048
rect 5252 2038 5259 2048
rect 5311 2082 5318 2090
rect 6512 2082 6519 2092
rect 5311 2048 6519 2082
rect 5311 2038 5318 2048
rect 6512 2040 6519 2048
rect 6571 2082 6578 2092
rect 7421 2082 7427 2090
rect 6571 2048 7427 2082
rect 6571 2040 6578 2048
rect 7421 2038 7427 2048
rect 7479 2082 7485 2090
rect 7644 2082 7651 2091
rect 7479 2048 7651 2082
rect 7479 2038 7485 2048
rect 7644 2039 7651 2048
rect 7703 2082 7710 2091
rect 8905 2082 8912 2092
rect 7703 2048 8912 2082
rect 7703 2039 7710 2048
rect 8905 2040 8912 2048
rect 8964 2082 8971 2092
rect 10035 2082 10042 2090
rect 8964 2048 10042 2082
rect 8964 2040 8971 2048
rect 10035 2038 10042 2048
rect 10094 2082 10101 2090
rect 11298 2082 11305 2092
rect 10094 2048 11305 2082
rect 10094 2038 10101 2048
rect 11298 2040 11305 2048
rect 11357 2082 11364 2092
rect 12427 2082 12434 2089
rect 11357 2048 12434 2082
rect 11357 2040 11364 2048
rect 12427 2037 12434 2048
rect 12486 2082 12493 2089
rect 13687 2082 13694 2092
rect 12486 2048 13694 2082
rect 12486 2037 12493 2048
rect 13687 2040 13694 2048
rect 13746 2082 13753 2092
rect 14819 2082 14826 2090
rect 13746 2048 14826 2082
rect 13746 2040 13753 2048
rect 14819 2038 14826 2048
rect 14878 2082 14885 2090
rect 16082 2082 16089 2092
rect 14878 2048 16089 2082
rect 14878 2038 14885 2048
rect 16082 2040 16089 2048
rect 16141 2082 16148 2092
rect 16141 2048 16861 2082
rect 16141 2040 16148 2048
rect 95 1944 16876 1976
rect 95 1942 16861 1944
rect -126 1856 16861 1860
rect -144 1840 16861 1856
rect -144 1837 5962 1840
rect -144 1836 5596 1837
rect -144 1834 3028 1836
rect -144 1832 2703 1834
rect -144 1780 19 1832
rect 71 1830 2703 1832
rect 71 1780 259 1830
rect -144 1778 259 1780
rect 311 1829 799 1830
rect 311 1778 581 1829
rect -144 1777 581 1778
rect 633 1778 799 1829
rect 851 1782 2703 1830
rect 2755 1784 3028 1834
rect 3080 1819 3296 1836
rect 3080 1795 3158 1819
rect 3192 1795 3296 1819
rect 3080 1784 3296 1795
rect 3348 1784 3562 1836
rect 3614 1834 5596 1836
rect 3614 1784 3802 1834
rect 2755 1782 3802 1784
rect 3854 1785 5596 1834
rect 5648 1788 5962 1837
rect 6014 1788 6206 1840
rect 6258 1838 16861 1840
rect 6258 1833 9030 1838
rect 6258 1831 8572 1833
rect 6258 1819 6629 1831
rect 6279 1818 6629 1819
rect 6258 1788 6629 1818
rect 5648 1785 6629 1788
rect 3854 1782 6629 1785
rect 851 1779 6629 1782
rect 6681 1781 8572 1831
rect 8624 1830 9030 1833
rect 8624 1781 8824 1830
rect 6681 1779 8824 1781
rect 851 1778 8824 1779
rect 8876 1786 9030 1830
rect 9082 1836 16861 1838
rect 9082 1834 11653 1836
rect 9082 1833 11443 1834
rect 9082 1832 9611 1833
rect 9082 1786 9313 1832
rect 8876 1780 9313 1786
rect 9365 1819 9611 1832
rect 9365 1795 9374 1819
rect 9408 1795 9611 1819
rect 9365 1781 9611 1795
rect 9663 1782 11443 1833
rect 11495 1784 11653 1834
rect 11705 1834 16861 1836
rect 11705 1784 12004 1834
rect 11495 1782 12004 1784
rect 12056 1782 12284 1834
rect 12336 1833 15547 1834
rect 12336 1782 12601 1833
rect 9663 1781 12601 1782
rect 12653 1831 15547 1833
rect 12653 1781 14391 1831
rect 9365 1780 14391 1781
rect 8876 1779 14391 1780
rect 14443 1779 14686 1831
rect 14738 1779 14973 1831
rect 15025 1779 15263 1831
rect 15315 1782 15547 1831
rect 15599 1782 16861 1834
rect 15315 1779 16861 1782
rect 8876 1778 16861 1779
rect 633 1777 16861 1778
rect -144 1770 16861 1777
rect -126 1764 16861 1770
rect 468 1565 475 1617
rect 527 1565 534 1617
rect 641 1591 710 1608
rect 1551 1591 1557 1603
rect 641 1557 656 1591
rect 690 1557 1557 1591
rect 641 1542 710 1557
rect 1551 1550 1557 1557
rect 1609 1550 1616 1603
rect 1730 1565 1737 1617
rect 1789 1565 1796 1617
rect 2861 1564 2868 1616
rect 2920 1564 2927 1616
rect 3033 1590 3103 1611
rect 3943 1590 3949 1602
rect 1551 1549 1616 1550
rect 3033 1556 3048 1590
rect 3082 1556 3949 1590
rect 3033 1541 3103 1556
rect 3943 1549 3949 1556
rect 4001 1549 4008 1602
rect 4122 1565 4129 1617
rect 4181 1565 4188 1617
rect 5253 1564 5260 1616
rect 5312 1564 5319 1616
rect 5424 1602 5488 1605
rect 5424 1591 5489 1602
rect 3943 1548 4008 1549
rect 5424 1557 5439 1591
rect 5473 1590 5489 1591
rect 6333 1590 6339 1602
rect 5473 1559 6339 1590
rect 5473 1557 5489 1559
rect 5424 1548 5489 1557
rect 6333 1549 6339 1559
rect 6391 1549 6398 1602
rect 6513 1566 6520 1618
rect 6572 1566 6579 1618
rect 7645 1565 7652 1617
rect 7704 1565 7711 1617
rect 7817 1591 7884 1604
rect 8727 1591 8733 1603
rect 6333 1548 6398 1549
rect 7817 1557 7832 1591
rect 7866 1558 8733 1591
rect 7866 1557 7884 1558
rect 5424 1546 5488 1548
rect 7817 1543 7884 1557
rect 8727 1550 8733 1558
rect 8785 1550 8792 1603
rect 8906 1566 8913 1618
rect 8965 1566 8972 1618
rect 10036 1564 10043 1616
rect 10095 1564 10102 1616
rect 10208 1592 10270 1607
rect 8727 1549 8792 1550
rect 10208 1558 10223 1592
rect 10257 1591 10270 1592
rect 11119 1591 11125 1602
rect 10257 1559 11125 1591
rect 10257 1558 10270 1559
rect 10208 1544 10270 1558
rect 11119 1549 11125 1559
rect 11177 1549 11184 1602
rect 11299 1566 11306 1618
rect 11358 1566 11365 1618
rect 12428 1563 12435 1615
rect 12487 1563 12494 1615
rect 12600 1593 12658 1604
rect 13508 1593 13514 1602
rect 12600 1592 13514 1593
rect 11119 1548 11184 1549
rect 12600 1558 12615 1592
rect 12649 1559 13514 1592
rect 12649 1558 12658 1559
rect 12600 1546 12658 1558
rect 13508 1549 13514 1559
rect 13566 1549 13573 1602
rect 13688 1566 13695 1618
rect 13747 1566 13754 1618
rect 14820 1564 14827 1616
rect 14879 1564 14886 1616
rect 14996 1592 15048 1598
rect 15903 1592 15909 1603
rect 14996 1558 15008 1592
rect 15042 1558 15909 1592
rect 14996 1552 15048 1558
rect 15903 1550 15909 1558
rect 15961 1550 15968 1603
rect 16083 1566 16090 1618
rect 16142 1566 16149 1618
rect 15903 1549 15968 1550
rect 13508 1548 13573 1549
rect 17 1414 71 1420
rect 17 1362 18 1414
rect 70 1362 71 1414
rect 349 1400 356 1452
rect 408 1448 414 1452
rect 1950 1448 1957 1453
rect 408 1406 1957 1448
rect 408 1400 414 1406
rect 1950 1401 1957 1406
rect 2009 1401 2015 1453
rect 2409 1414 2463 1420
rect 2188 1362 2194 1414
rect 2246 1362 2254 1414
rect 2409 1362 2410 1414
rect 2462 1362 2463 1414
rect 2741 1400 2748 1452
rect 2800 1448 2806 1452
rect 4342 1448 4349 1453
rect 2800 1406 4349 1448
rect 2800 1400 2806 1406
rect 4342 1401 4349 1406
rect 4401 1401 4407 1453
rect 4801 1414 4855 1420
rect 4582 1362 4588 1414
rect 4640 1362 4648 1414
rect 4801 1362 4802 1414
rect 4854 1362 4855 1414
rect 5132 1401 5139 1453
rect 5191 1449 5197 1453
rect 6733 1449 6740 1454
rect 5191 1407 6740 1449
rect 5191 1401 5197 1407
rect 6733 1402 6740 1407
rect 6792 1402 6798 1454
rect 6972 1364 6978 1416
rect 7030 1364 7038 1416
rect 7193 1414 7247 1420
rect 17 1356 71 1362
rect 2409 1356 2463 1362
rect 4801 1356 4855 1362
rect 7193 1362 7194 1414
rect 7246 1362 7247 1414
rect 7525 1400 7532 1452
rect 7584 1448 7590 1452
rect 9126 1448 9133 1453
rect 7584 1406 9133 1448
rect 7584 1400 7590 1406
rect 9126 1401 9133 1406
rect 9185 1401 9191 1453
rect 9584 1415 9638 1421
rect 9364 1362 9370 1414
rect 9422 1362 9430 1414
rect 9584 1363 9585 1415
rect 9637 1363 9638 1415
rect 9917 1401 9924 1453
rect 9976 1449 9982 1453
rect 11518 1449 11525 1454
rect 9976 1407 11525 1449
rect 9976 1401 9982 1407
rect 11518 1402 11525 1407
rect 11577 1402 11583 1454
rect 11756 1364 11762 1416
rect 11814 1364 11822 1416
rect 11976 1414 12030 1420
rect 7193 1356 7247 1362
rect 9584 1357 9638 1363
rect 11976 1362 11977 1414
rect 12029 1362 12030 1414
rect 12309 1401 12316 1453
rect 12368 1449 12374 1453
rect 13910 1449 13917 1454
rect 12368 1407 13917 1449
rect 12368 1401 12374 1407
rect 13910 1402 13917 1407
rect 13969 1402 13975 1454
rect 14369 1415 14423 1421
rect 14148 1362 14154 1414
rect 14206 1362 14214 1414
rect 14369 1363 14370 1415
rect 14422 1363 14423 1415
rect 14704 1401 14711 1453
rect 14763 1449 14769 1453
rect 16305 1449 16312 1454
rect 14763 1407 16312 1449
rect 14763 1401 14769 1407
rect 16305 1402 16312 1407
rect 16364 1402 16370 1454
rect 16540 1364 16546 1416
rect 16598 1364 16606 1416
rect 11976 1356 12030 1362
rect 14369 1357 14423 1363
rect 16175 1316 16205 1362
rect -126 1314 16861 1316
rect -126 1301 16876 1314
rect -126 1299 10510 1301
rect -126 1297 7858 1299
rect -126 1294 7668 1297
rect -126 1242 1210 1294
rect 1262 1242 1427 1294
rect 1479 1242 1646 1294
rect 1698 1290 5044 1294
rect 1698 1242 1859 1290
rect -126 1238 1859 1242
rect 1911 1238 2070 1290
rect 2122 1238 4194 1290
rect 4246 1289 5044 1290
rect 4246 1238 4472 1289
rect -126 1237 4472 1238
rect 4524 1242 5044 1289
rect 5096 1242 5283 1294
rect 5335 1292 7668 1294
rect 5335 1242 7441 1292
rect 4524 1240 7441 1242
rect 7493 1245 7668 1292
rect 7720 1247 7858 1297
rect 7910 1296 10510 1299
rect 7910 1293 10284 1296
rect 7910 1290 10055 1293
rect 7910 1247 8074 1290
rect 7720 1245 8074 1247
rect 7493 1240 8074 1245
rect 4524 1238 8074 1240
rect 8126 1241 10055 1290
rect 10107 1244 10284 1293
rect 10336 1249 10510 1296
rect 10562 1299 16876 1301
rect 10562 1293 10974 1299
rect 10562 1249 10738 1293
rect 10336 1244 10738 1249
rect 10107 1241 10738 1244
rect 10790 1247 10974 1293
rect 11026 1298 16876 1299
rect 11026 1295 16022 1298
rect 11026 1290 13105 1295
rect 11026 1247 11166 1290
rect 10790 1241 11166 1247
rect 8126 1238 11166 1241
rect 11218 1238 12901 1290
rect 12953 1243 13105 1290
rect 13157 1294 16022 1295
rect 13157 1290 15828 1294
rect 13157 1243 13296 1290
rect 12953 1238 13296 1243
rect 13348 1289 13788 1290
rect 13348 1238 13498 1289
rect 4524 1237 13498 1238
rect 13550 1238 13788 1289
rect 13840 1289 15828 1290
rect 13840 1238 14073 1289
rect 13550 1237 14073 1238
rect 14125 1242 15828 1289
rect 15880 1246 16022 1294
rect 16074 1297 16876 1298
rect 16074 1295 16434 1297
rect 16074 1246 16211 1295
rect 15880 1243 16211 1246
rect 16263 1245 16434 1295
rect 16486 1245 16876 1297
rect 16263 1243 16876 1245
rect 15880 1242 16876 1243
rect 14125 1237 16876 1242
rect -126 1228 16876 1237
rect -126 1220 16861 1228
rect 16237 1172 16303 1173
rect -126 1164 16782 1172
rect -144 1151 16782 1164
rect -144 1150 8753 1151
rect -144 1149 3262 1150
rect -144 1097 265 1149
rect 317 1146 3262 1149
rect 317 1145 2654 1146
rect 317 1097 467 1145
rect -144 1093 467 1097
rect 519 1143 2654 1145
rect 519 1142 885 1143
rect 519 1093 656 1142
rect -144 1090 656 1093
rect 708 1091 885 1142
rect 937 1094 2654 1143
rect 2706 1143 3262 1146
rect 2706 1094 2869 1143
rect 937 1091 2869 1094
rect 2921 1140 3262 1143
rect 2921 1091 3067 1140
rect 708 1090 3067 1091
rect -144 1088 3067 1090
rect 3119 1098 3262 1140
rect 3314 1149 8753 1150
rect 3314 1148 8563 1149
rect 3314 1098 3542 1148
rect 3119 1096 3542 1098
rect 3594 1147 8563 1148
rect 3594 1146 6518 1147
rect 3594 1096 3761 1146
rect 3119 1094 3761 1096
rect 3813 1145 6518 1146
rect 3813 1143 6327 1145
rect 3813 1094 5582 1143
rect 3119 1091 5582 1094
rect 5634 1140 6327 1143
rect 5634 1091 5933 1140
rect 3119 1088 5933 1091
rect 5985 1138 6327 1140
rect 5985 1088 6122 1138
rect -144 1086 6122 1088
rect 6174 1093 6327 1138
rect 6379 1095 6518 1145
rect 6570 1097 8563 1147
rect 8615 1099 8753 1149
rect 8805 1150 16782 1151
rect 8805 1149 14613 1150
rect 8805 1099 8947 1149
rect 8615 1097 8947 1099
rect 8999 1145 14613 1149
rect 8999 1097 9258 1145
rect 6570 1095 9258 1097
rect 6379 1093 9258 1095
rect 9310 1144 14613 1145
rect 9310 1093 11441 1144
rect 6174 1092 11441 1093
rect 11493 1092 11645 1144
rect 11697 1142 14613 1144
rect 11697 1140 12449 1142
rect 11697 1092 12210 1140
rect 6174 1088 12210 1092
rect 12262 1090 12449 1140
rect 12501 1090 12653 1142
rect 12705 1098 14613 1142
rect 14665 1148 15542 1150
rect 14665 1098 14846 1148
rect 12705 1096 14846 1098
rect 14898 1146 15262 1148
rect 14898 1096 15053 1146
rect 12705 1094 15053 1096
rect 15105 1096 15262 1146
rect 15314 1098 15542 1148
rect 15594 1098 16782 1150
rect 15314 1096 16782 1098
rect 15105 1094 16782 1096
rect 12705 1090 16782 1094
rect 12262 1088 16782 1090
rect 6174 1086 16782 1088
rect -144 1078 16782 1086
rect -126 1076 16782 1078
rect 2324 1042 2376 1048
rect 2324 984 2376 990
rect 4716 1042 4768 1048
rect 4716 984 4768 990
rect 7108 1042 7160 1048
rect 7108 984 7160 990
rect 9500 1042 9552 1048
rect 9500 984 9552 990
rect 11892 1042 11944 1048
rect 11892 984 11944 990
rect 14284 1042 14336 1048
rect 14284 984 14336 990
rect 16676 1042 16728 1048
rect 16676 984 16728 990
rect 2042 965 2094 971
rect 2042 907 2094 913
rect 4434 966 4486 972
rect 4434 908 4486 914
rect 6825 966 6877 972
rect 6825 908 6877 914
rect 9218 967 9270 973
rect 9218 909 9270 915
rect 11609 966 11661 972
rect 11609 908 11661 914
rect 14002 965 14054 971
rect 14002 907 14054 913
rect 16395 967 16447 973
rect 16395 909 16447 915
rect 17 869 71 875
rect 17 817 18 869
rect 70 817 71 869
rect 351 841 357 894
rect 409 841 416 894
rect 351 840 416 841
rect 2409 869 2463 875
rect 17 811 71 817
rect 2409 817 2410 869
rect 2462 817 2463 869
rect 2743 841 2749 894
rect 2801 841 2808 894
rect 2743 840 2808 841
rect 4801 869 4855 875
rect 2409 811 2463 817
rect 4801 817 4802 869
rect 4854 817 4855 869
rect 5135 842 5141 895
rect 5193 842 5200 895
rect 5135 841 5200 842
rect 7193 869 7247 875
rect 4801 811 4855 817
rect 7193 817 7194 869
rect 7246 817 7247 869
rect 7527 842 7533 895
rect 7585 842 7592 895
rect 7527 841 7592 842
rect 9584 870 9638 876
rect 7193 811 7247 817
rect 9584 818 9585 870
rect 9637 818 9638 870
rect 9919 841 9925 894
rect 9977 841 9984 894
rect 9919 840 9984 841
rect 11976 869 12030 875
rect 9584 812 9638 818
rect 11976 817 11977 869
rect 12029 817 12030 869
rect 12311 842 12317 895
rect 12369 842 12376 895
rect 12311 841 12376 842
rect 14369 870 14423 876
rect 11976 811 12030 817
rect 14369 818 14370 870
rect 14422 818 14423 870
rect 14704 841 14710 894
rect 14762 841 14769 894
rect 14704 840 14769 841
rect 14369 812 14423 818
rect 1024 770 1078 776
rect 1024 718 1025 770
rect 1077 718 1078 770
rect 1024 712 1078 718
rect 3417 770 3471 776
rect 3417 718 3418 770
rect 3470 718 3471 770
rect 3417 712 3471 718
rect 5809 770 5863 776
rect 5809 718 5810 770
rect 5862 718 5863 770
rect 5809 712 5863 718
rect 8201 770 8255 776
rect 8201 718 8202 770
rect 8254 718 8255 770
rect 8201 712 8255 718
rect 10592 770 10646 776
rect 10592 718 10593 770
rect 10645 718 10646 770
rect 10592 710 10646 718
rect 12984 770 13038 776
rect 12984 718 12985 770
rect 13037 718 13038 770
rect 12984 712 13038 718
rect 15376 770 15430 776
rect 15376 718 15377 770
rect 15429 718 15430 770
rect 15376 712 15430 718
rect 16816 628 16861 632
rect -126 612 16876 628
rect -126 600 1421 612
rect -126 548 1192 600
rect 1244 560 1421 600
rect 1473 611 16876 612
rect 1473 609 5038 611
rect 1473 606 4708 609
rect 1473 602 1832 606
rect 1473 560 1640 602
rect 1244 550 1640 560
rect 1692 554 1832 602
rect 1884 604 4708 606
rect 1884 554 2326 604
rect 1692 552 2326 554
rect 2378 603 4708 604
rect 2378 552 4118 603
rect 1692 551 4118 552
rect 4170 601 4708 603
rect 4170 551 4511 601
rect 1692 550 4511 551
rect 1244 549 4511 550
rect 4563 557 4708 601
rect 4760 559 5038 609
rect 5090 559 5234 611
rect 5286 609 8069 611
rect 5286 608 7648 609
rect 5286 604 7442 608
rect 5286 559 7141 604
rect 4760 557 7141 559
rect 4563 552 7141 557
rect 7193 556 7442 604
rect 7494 557 7648 608
rect 7700 605 8069 609
rect 7700 557 7858 605
rect 7494 556 7858 557
rect 7193 553 7858 556
rect 7910 559 8069 605
rect 8121 608 10968 611
rect 8121 607 10727 608
rect 8121 600 10206 607
rect 8121 559 9949 600
rect 7910 553 9949 559
rect 7193 552 9949 553
rect 4563 549 9949 552
rect 1244 548 9949 549
rect 10001 555 10206 600
rect 10258 603 10727 607
rect 10258 555 10456 603
rect 10001 551 10456 555
rect 10508 556 10727 603
rect 10779 559 10968 608
rect 11020 610 16876 611
rect 11020 608 16216 610
rect 11020 607 16021 608
rect 11020 559 11193 607
rect 10779 556 11193 559
rect 10508 555 11193 556
rect 11245 606 16021 607
rect 11245 605 13101 606
rect 11245 555 12900 605
rect 10508 553 12900 555
rect 12952 554 13101 605
rect 13153 602 13526 606
rect 13153 554 13319 602
rect 12952 553 13319 554
rect 10508 551 13319 553
rect 10001 550 13319 551
rect 13371 554 13526 602
rect 13578 605 16021 606
rect 13578 554 13731 605
rect 13371 553 13731 554
rect 13783 601 15830 605
rect 13783 553 14078 601
rect 13371 550 14078 553
rect 10001 549 14078 550
rect 14130 553 15830 601
rect 15882 556 16021 605
rect 16073 558 16216 608
rect 16268 605 16876 610
rect 16268 558 16663 605
rect 16073 556 16663 558
rect 15882 553 16663 556
rect 16715 553 16876 605
rect 14130 549 16876 553
rect 10001 548 16876 549
rect -126 542 16876 548
rect -126 536 16861 542
rect -126 532 16816 536
rect 1591 483 1657 487
rect 3983 483 4049 487
rect 6375 483 6441 487
rect 8767 483 8833 487
rect 11159 483 11225 487
rect 13551 483 13617 487
rect 15943 483 16009 485
rect 16816 483 16861 487
rect -126 476 16861 483
rect -144 464 16861 476
rect -144 461 15022 464
rect -144 459 3786 461
rect -144 456 495 459
rect -144 404 47 456
rect 99 452 495 456
rect 99 404 280 452
rect -144 400 280 404
rect 332 407 495 452
rect 547 457 3786 459
rect 547 456 929 457
rect 547 407 713 456
rect 332 404 713 407
rect 765 405 929 456
rect 981 456 3786 457
rect 981 453 3050 456
rect 981 405 2650 453
rect 765 404 2650 405
rect 332 401 2650 404
rect 2702 401 2840 453
rect 2892 404 3050 453
rect 3102 453 3562 456
rect 3102 404 3267 453
rect 2892 401 3267 404
rect 3319 404 3562 453
rect 3614 409 3786 456
rect 3838 456 6433 461
rect 3838 454 6216 456
rect 3838 409 5664 454
rect 3614 404 5664 409
rect 3319 402 5664 404
rect 5716 452 6216 454
rect 5716 402 5964 452
rect 3319 401 5964 402
rect 332 400 5964 401
rect 6016 404 6216 452
rect 6268 409 6433 456
rect 6485 458 14390 461
rect 6485 409 6634 458
rect 6268 406 6634 409
rect 6686 457 14390 458
rect 6686 449 9529 457
rect 6686 406 8519 449
rect 6268 404 8519 406
rect 6016 400 8519 404
rect -144 397 8519 400
rect 8571 397 8711 449
rect 8763 397 8911 449
rect 8963 405 9529 449
rect 9581 455 14390 457
rect 9581 453 12210 455
rect 9581 405 11430 453
rect 8963 401 11430 405
rect 11482 401 11686 453
rect 11738 401 11921 453
rect 11973 403 12210 453
rect 12262 453 12604 455
rect 12262 403 12400 453
rect 11973 401 12400 403
rect 12452 403 12604 453
rect 12656 409 14390 455
rect 14442 457 15022 461
rect 14442 409 14632 457
rect 12656 405 14632 409
rect 14684 456 15022 457
rect 14684 405 14832 456
rect 12656 404 14832 405
rect 14884 412 15022 456
rect 15074 462 16861 464
rect 15074 412 15243 462
rect 14884 410 15243 412
rect 15295 457 16861 462
rect 15295 410 15539 457
rect 14884 405 15539 410
rect 15591 405 16861 457
rect 14884 404 16861 405
rect 12656 403 16861 404
rect 12452 401 16861 403
rect 8963 397 16861 401
rect -144 391 16861 397
rect -144 390 1591 391
rect -126 387 1591 390
rect 1657 387 16816 391
rect 12384 386 12481 387
rect 17 350 69 356
rect 2409 350 2461 356
rect 1019 302 1025 314
rect 17 292 69 298
rect 297 286 349 292
rect 297 228 349 234
rect 508 271 1025 302
rect 508 154 537 271
rect 1019 262 1025 271
rect 1077 262 1083 314
rect 4802 350 4854 356
rect 3411 303 3417 315
rect 2409 292 2461 298
rect 2689 286 2741 292
rect 2689 228 2741 234
rect 2900 272 3417 303
rect 2298 163 2304 215
rect 2358 163 2364 215
rect 490 148 548 154
rect 490 114 502 148
rect 536 114 548 148
rect 490 108 548 114
rect 508 107 537 108
rect 1953 107 1959 160
rect 2011 107 2018 160
rect 2900 156 2929 272
rect 3411 263 3417 272
rect 3469 263 3475 315
rect 7193 350 7245 356
rect 5803 302 5809 314
rect 4802 292 4854 298
rect 5080 286 5132 292
rect 5080 228 5132 234
rect 5292 271 5809 302
rect 4692 163 4698 215
rect 4752 163 4758 215
rect 2879 150 2937 156
rect 2879 116 2891 150
rect 2925 116 2937 150
rect 2879 110 2937 116
rect 2900 108 2929 110
rect 1953 106 2018 107
rect 4345 107 4351 160
rect 4403 107 4410 160
rect 5292 156 5321 271
rect 5803 262 5809 271
rect 5861 262 5867 314
rect 9585 349 9637 355
rect 8195 302 8201 314
rect 7193 292 7245 298
rect 7473 286 7525 292
rect 7473 228 7525 234
rect 7684 271 8201 302
rect 7082 165 7088 217
rect 7142 165 7148 217
rect 6736 160 6801 161
rect 5272 150 5330 156
rect 5272 116 5284 150
rect 5318 116 5330 150
rect 5272 110 5330 116
rect 5292 107 5321 110
rect 6736 108 6742 160
rect 6794 108 6801 160
rect 7684 156 7713 271
rect 8195 262 8201 271
rect 8253 262 8259 314
rect 11978 351 12030 357
rect 10587 302 10593 314
rect 9585 291 9637 297
rect 9865 286 9917 292
rect 9865 228 9917 234
rect 10076 271 10593 302
rect 9474 163 9480 215
rect 9534 163 9540 215
rect 7665 150 7723 156
rect 7665 116 7677 150
rect 7711 116 7723 150
rect 7665 110 7723 116
rect 6736 107 6801 108
rect 7684 107 7713 110
rect 9129 107 9135 160
rect 9187 107 9194 160
rect 10076 156 10105 271
rect 10587 262 10593 271
rect 10645 262 10651 314
rect 14369 351 14421 357
rect 12979 303 12985 315
rect 11978 293 12030 299
rect 12256 287 12308 293
rect 12256 229 12308 235
rect 12468 272 12985 303
rect 11866 165 11872 217
rect 11926 165 11932 217
rect 10056 150 10114 156
rect 10056 116 10068 150
rect 10102 116 10114 150
rect 10056 110 10114 116
rect 10076 107 10105 110
rect 11520 107 11526 160
rect 11578 107 11585 160
rect 12468 156 12497 272
rect 12979 263 12985 272
rect 13037 263 13043 315
rect 15371 303 15377 315
rect 14369 293 14421 299
rect 14649 286 14701 292
rect 14649 228 14701 234
rect 14860 272 15377 303
rect 14258 163 14264 215
rect 14318 163 14324 215
rect 12449 150 12507 156
rect 12449 116 12461 150
rect 12495 116 12507 150
rect 12449 110 12507 116
rect 12468 108 12497 110
rect 4345 106 4410 107
rect 9129 106 9194 107
rect 11520 106 11585 107
rect 13913 107 13919 160
rect 13971 107 13978 160
rect 14860 156 14889 272
rect 15371 263 15377 272
rect 15429 263 15435 315
rect 16650 165 16656 217
rect 16710 165 16716 217
rect 14840 150 14898 156
rect 14840 116 14852 150
rect 14886 116 14898 150
rect 14840 110 14898 116
rect 14860 108 14889 110
rect 13913 106 13978 107
rect 16306 107 16312 160
rect 16364 107 16371 160
rect 16306 106 16371 107
rect 16816 -61 16861 -57
rect -126 -64 16861 -61
rect -126 -74 16876 -64
rect -126 -76 2163 -74
rect -126 -128 421 -76
rect 473 -79 2163 -76
rect 473 -128 620 -79
rect -126 -131 620 -128
rect 672 -131 831 -79
rect 883 -131 1037 -79
rect 1089 -81 1739 -79
rect 1089 -131 1265 -81
rect -126 -133 1265 -131
rect 1317 -133 1509 -81
rect 1561 -131 1739 -81
rect 1791 -131 1945 -79
rect 1997 -126 2163 -79
rect 2215 -77 16876 -74
rect 2215 -80 2574 -77
rect 2215 -126 2366 -80
rect 1997 -131 2366 -126
rect 1561 -132 2366 -131
rect 2418 -129 2574 -80
rect 2626 -80 3455 -77
rect 2626 -81 3045 -80
rect 2626 -129 2837 -81
rect 2418 -132 2837 -129
rect 1561 -133 2837 -132
rect 2889 -132 3045 -81
rect 3097 -83 3455 -80
rect 3097 -132 3255 -83
rect 2889 -133 3255 -132
rect -126 -135 3255 -133
rect 3307 -129 3455 -83
rect 3507 -78 7335 -77
rect 3507 -79 4285 -78
rect 3507 -80 4069 -79
rect 3507 -129 3658 -80
rect 3307 -132 3658 -129
rect 3710 -132 3868 -80
rect 3920 -131 4069 -80
rect 4121 -130 4285 -79
rect 4337 -80 5212 -78
rect 4337 -130 4566 -80
rect 4121 -131 4566 -130
rect 3920 -132 4566 -131
rect 4618 -84 5212 -80
rect 4618 -85 4991 -84
rect 4618 -132 4786 -85
rect 3307 -135 4786 -132
rect -126 -137 4786 -135
rect 4838 -136 4991 -85
rect 5043 -130 5212 -84
rect 5264 -79 7335 -78
rect 5264 -84 6057 -79
rect 5264 -85 5626 -84
rect 5264 -130 5417 -85
rect 5043 -136 5417 -130
rect 4838 -137 5417 -136
rect 5469 -136 5626 -85
rect 5678 -136 5843 -84
rect 5895 -131 6057 -84
rect 6109 -80 7132 -79
rect 6109 -81 6933 -80
rect 6109 -131 6252 -81
rect 5895 -133 6252 -131
rect 6304 -84 6649 -81
rect 6304 -133 6447 -84
rect 5895 -136 6447 -133
rect 6499 -133 6649 -84
rect 6701 -132 6933 -81
rect 6985 -131 7132 -80
rect 7184 -129 7335 -79
rect 7387 -78 10817 -77
rect 7387 -79 9034 -78
rect 7387 -80 7987 -79
rect 7387 -129 7600 -80
rect 7184 -131 7600 -129
rect 6985 -132 7600 -131
rect 7652 -81 7987 -80
rect 7652 -132 7798 -81
rect 6701 -133 7798 -132
rect 7850 -131 7987 -81
rect 8039 -131 8199 -79
rect 8251 -131 8416 -79
rect 8468 -83 9034 -79
rect 8468 -131 8621 -83
rect 7850 -133 8621 -131
rect 6499 -135 8621 -133
rect 8673 -135 8826 -83
rect 8878 -130 9034 -83
rect 9086 -79 10817 -78
rect 9086 -130 9317 -79
rect 8878 -131 9317 -130
rect 9369 -81 10195 -79
rect 9369 -131 9510 -81
rect 8878 -133 9510 -131
rect 9562 -83 10195 -81
rect 9562 -133 9736 -83
rect 8878 -135 9736 -133
rect 9788 -135 10001 -83
rect 10053 -131 10195 -83
rect 10247 -80 10817 -79
rect 10247 -88 10597 -80
rect 10247 -131 10393 -88
rect 10053 -135 10393 -131
rect 6499 -136 10393 -135
rect 5469 -137 10393 -136
rect -126 -140 10393 -137
rect 10445 -132 10597 -88
rect 10649 -129 10817 -80
rect 10869 -78 16876 -77
rect 10869 -81 11260 -78
rect 10869 -129 11032 -81
rect 10649 -132 11032 -129
rect 10445 -133 11032 -132
rect 11084 -130 11260 -81
rect 11312 -79 11895 -78
rect 11312 -81 11702 -79
rect 11312 -130 11464 -81
rect 11084 -133 11464 -130
rect 11516 -131 11702 -81
rect 11754 -130 11895 -79
rect 11947 -80 16876 -78
rect 11947 -83 12348 -80
rect 11947 -130 12092 -83
rect 11754 -131 12092 -130
rect 11516 -133 12092 -131
rect 10445 -135 12092 -133
rect 12144 -132 12348 -83
rect 12400 -81 16876 -80
rect 12400 -83 13460 -81
rect 12400 -84 13041 -83
rect 12400 -132 12587 -84
rect 12144 -135 12587 -132
rect 10445 -136 12587 -135
rect 12639 -88 13041 -84
rect 12639 -136 12820 -88
rect 10445 -140 12820 -136
rect 12872 -135 13041 -88
rect 13093 -135 13232 -83
rect 13284 -133 13460 -83
rect 13512 -82 14511 -81
rect 13512 -83 14285 -82
rect 13512 -86 14096 -83
rect 13512 -133 13657 -86
rect 13284 -135 13657 -133
rect 12872 -138 13657 -135
rect 13709 -138 13869 -86
rect 13921 -135 14096 -86
rect 14148 -134 14285 -83
rect 14337 -133 14511 -82
rect 14563 -133 14765 -81
rect 14817 -82 16497 -81
rect 14817 -84 15497 -82
rect 14817 -133 15009 -84
rect 14337 -134 15009 -133
rect 14148 -135 15009 -134
rect 13921 -136 15009 -135
rect 15061 -85 15497 -84
rect 15061 -136 15239 -85
rect 13921 -137 15239 -136
rect 15291 -134 15497 -85
rect 15549 -134 15707 -82
rect 15759 -134 15932 -82
rect 15984 -85 16497 -82
rect 15984 -134 16151 -85
rect 15291 -137 16151 -134
rect 16203 -133 16497 -85
rect 16549 -84 16876 -81
rect 16549 -133 16696 -84
rect 16203 -136 16696 -133
rect 16748 -136 16876 -84
rect 16203 -137 16876 -136
rect 13921 -138 16876 -137
rect 12872 -140 16876 -138
rect -126 -150 16876 -140
rect -126 -153 16861 -150
rect -126 -157 16816 -153
<< via1 >>
rect 723 3383 775 3435
rect 53 2924 105 2976
rect 255 2926 307 2978
rect 466 2924 518 2976
rect 656 2924 708 2976
rect 864 2926 916 2978
rect 1066 2926 1118 2978
rect 1265 2928 1317 2980
rect 1460 2925 1512 2977
rect 1661 2927 1713 2979
rect 1878 2925 1930 2977
rect 2152 2928 2204 2980
rect 2429 2921 2481 2973
rect 2652 2924 2704 2976
rect 2884 2923 2936 2975
rect 4520 2920 4572 2972
rect 4828 2921 4880 2973
rect 5028 2922 5080 2974
rect 5247 2921 5299 2973
rect 5493 2920 5545 2972
rect 5701 2922 5753 2974
rect 5903 2923 5955 2975
rect 6096 2922 6148 2974
rect 6468 2921 6520 2973
rect 6657 2919 6709 2971
rect 6947 2919 6999 2971
rect 7220 2921 7272 2973
rect 2866 2664 2918 2674
rect 2866 2630 2876 2664
rect 2876 2630 2910 2664
rect 2910 2630 2918 2664
rect 2866 2622 2918 2630
rect 7427 2622 7479 2674
rect 1171 2385 1223 2437
rect 1390 2389 1442 2441
rect 1673 2389 1725 2441
rect 1882 2389 1934 2441
rect 2153 2387 2205 2439
rect 4228 2385 4280 2437
rect 4477 2388 4529 2440
rect 4821 2374 4873 2426
rect 5075 2380 5127 2432
rect 5304 2380 5356 2432
rect 7022 2385 7074 2437
rect 7226 2387 7278 2439
rect 7549 2385 7601 2437
rect 1024 2250 1077 2303
rect 2866 2250 2918 2302
rect 3418 2256 3471 2309
rect 5809 2256 5862 2309
rect 8200 2256 8253 2309
rect 10592 2256 10645 2309
rect 12983 2256 13036 2309
rect 15376 2256 15429 2309
rect 474 2039 526 2091
rect 1736 2039 1788 2091
rect 2867 2038 2919 2090
rect 4128 2039 4180 2091
rect 5259 2038 5311 2090
rect 6519 2040 6571 2092
rect 7427 2038 7479 2090
rect 7651 2039 7703 2091
rect 8912 2040 8964 2092
rect 10042 2038 10094 2090
rect 11305 2040 11357 2092
rect 12434 2037 12486 2089
rect 13694 2040 13746 2092
rect 14826 2038 14878 2090
rect 16089 2040 16141 2092
rect 19 1780 71 1832
rect 259 1778 311 1830
rect 581 1777 633 1829
rect 799 1778 851 1830
rect 2703 1782 2755 1834
rect 3028 1784 3080 1836
rect 3296 1784 3348 1836
rect 3562 1784 3614 1836
rect 3802 1782 3854 1834
rect 5596 1785 5648 1837
rect 5962 1788 6014 1840
rect 6206 1788 6258 1840
rect 6629 1779 6681 1831
rect 8572 1781 8624 1833
rect 8824 1778 8876 1830
rect 9030 1786 9082 1838
rect 9313 1780 9365 1832
rect 9611 1781 9663 1833
rect 11443 1782 11495 1834
rect 11653 1784 11705 1836
rect 12004 1782 12056 1834
rect 12284 1782 12336 1834
rect 12601 1781 12653 1833
rect 14391 1779 14443 1831
rect 14686 1779 14738 1831
rect 14973 1779 15025 1831
rect 15263 1779 15315 1831
rect 15547 1782 15599 1834
rect 475 1607 527 1617
rect 475 1573 484 1607
rect 484 1573 518 1607
rect 518 1573 527 1607
rect 475 1565 527 1573
rect 1557 1592 1609 1603
rect 1557 1558 1566 1592
rect 1566 1558 1600 1592
rect 1600 1558 1609 1592
rect 1557 1550 1609 1558
rect 1737 1607 1789 1617
rect 1737 1573 1746 1607
rect 1746 1573 1780 1607
rect 1780 1573 1789 1607
rect 1737 1565 1789 1573
rect 2868 1606 2920 1616
rect 2868 1572 2877 1606
rect 2877 1572 2911 1606
rect 2911 1572 2920 1606
rect 2868 1564 2920 1572
rect 3949 1591 4001 1602
rect 3949 1557 3958 1591
rect 3958 1557 3992 1591
rect 3992 1557 4001 1591
rect 3949 1549 4001 1557
rect 4129 1607 4181 1617
rect 4129 1573 4138 1607
rect 4138 1573 4172 1607
rect 4172 1573 4181 1607
rect 4129 1565 4181 1573
rect 5260 1606 5312 1616
rect 5260 1572 5269 1606
rect 5269 1572 5303 1606
rect 5303 1572 5312 1606
rect 5260 1564 5312 1572
rect 6339 1591 6391 1602
rect 6339 1557 6348 1591
rect 6348 1557 6382 1591
rect 6382 1557 6391 1591
rect 6339 1549 6391 1557
rect 6520 1608 6572 1618
rect 6520 1574 6529 1608
rect 6529 1574 6563 1608
rect 6563 1574 6572 1608
rect 6520 1566 6572 1574
rect 7652 1607 7704 1617
rect 7652 1573 7661 1607
rect 7661 1573 7695 1607
rect 7695 1573 7704 1607
rect 7652 1565 7704 1573
rect 8733 1592 8785 1603
rect 8733 1558 8742 1592
rect 8742 1558 8776 1592
rect 8776 1558 8785 1592
rect 8733 1550 8785 1558
rect 8913 1608 8965 1618
rect 8913 1574 8922 1608
rect 8922 1574 8956 1608
rect 8956 1574 8965 1608
rect 8913 1566 8965 1574
rect 10043 1606 10095 1616
rect 10043 1572 10052 1606
rect 10052 1572 10086 1606
rect 10086 1572 10095 1606
rect 10043 1564 10095 1572
rect 11125 1591 11177 1602
rect 11125 1557 11134 1591
rect 11134 1557 11168 1591
rect 11168 1557 11177 1591
rect 11125 1549 11177 1557
rect 11306 1608 11358 1618
rect 11306 1574 11315 1608
rect 11315 1574 11349 1608
rect 11349 1574 11358 1608
rect 11306 1566 11358 1574
rect 12435 1605 12487 1615
rect 12435 1571 12444 1605
rect 12444 1571 12478 1605
rect 12478 1571 12487 1605
rect 12435 1563 12487 1571
rect 13514 1591 13566 1602
rect 13514 1557 13523 1591
rect 13523 1557 13557 1591
rect 13557 1557 13566 1591
rect 13514 1549 13566 1557
rect 13695 1608 13747 1618
rect 13695 1574 13704 1608
rect 13704 1574 13738 1608
rect 13738 1574 13747 1608
rect 13695 1566 13747 1574
rect 14827 1606 14879 1616
rect 14827 1572 14836 1606
rect 14836 1572 14870 1606
rect 14870 1572 14879 1606
rect 14827 1564 14879 1572
rect 15909 1592 15961 1603
rect 15909 1558 15918 1592
rect 15918 1558 15952 1592
rect 15952 1558 15961 1592
rect 15909 1550 15961 1558
rect 16090 1608 16142 1618
rect 16090 1574 16099 1608
rect 16099 1574 16133 1608
rect 16133 1574 16142 1608
rect 16090 1566 16142 1574
rect 18 1406 70 1414
rect 18 1372 28 1406
rect 28 1372 62 1406
rect 62 1372 70 1406
rect 18 1362 70 1372
rect 356 1400 408 1452
rect 1957 1401 2009 1453
rect 2194 1404 2246 1414
rect 2194 1370 2204 1404
rect 2204 1370 2238 1404
rect 2238 1370 2246 1404
rect 2194 1362 2246 1370
rect 2410 1406 2462 1414
rect 2410 1372 2420 1406
rect 2420 1372 2454 1406
rect 2454 1372 2462 1406
rect 2410 1362 2462 1372
rect 2748 1400 2800 1452
rect 4349 1401 4401 1453
rect 4588 1404 4640 1414
rect 4588 1370 4598 1404
rect 4598 1370 4632 1404
rect 4632 1370 4640 1404
rect 4588 1362 4640 1370
rect 4802 1406 4854 1414
rect 4802 1372 4812 1406
rect 4812 1372 4846 1406
rect 4846 1372 4854 1406
rect 4802 1362 4854 1372
rect 5139 1401 5191 1453
rect 6740 1402 6792 1454
rect 6978 1406 7030 1416
rect 6978 1372 6988 1406
rect 6988 1372 7022 1406
rect 7022 1372 7030 1406
rect 6978 1364 7030 1372
rect 7194 1406 7246 1414
rect 7194 1372 7204 1406
rect 7204 1372 7238 1406
rect 7238 1372 7246 1406
rect 7194 1362 7246 1372
rect 7532 1400 7584 1452
rect 9133 1401 9185 1453
rect 9370 1404 9422 1414
rect 9370 1370 9380 1404
rect 9380 1370 9414 1404
rect 9414 1370 9422 1404
rect 9370 1362 9422 1370
rect 9585 1407 9637 1415
rect 9585 1373 9595 1407
rect 9595 1373 9629 1407
rect 9629 1373 9637 1407
rect 9585 1363 9637 1373
rect 9924 1401 9976 1453
rect 11525 1402 11577 1454
rect 11762 1406 11814 1416
rect 11762 1372 11772 1406
rect 11772 1372 11806 1406
rect 11806 1372 11814 1406
rect 11762 1364 11814 1372
rect 11977 1406 12029 1414
rect 11977 1372 11987 1406
rect 11987 1372 12021 1406
rect 12021 1372 12029 1406
rect 11977 1362 12029 1372
rect 12316 1401 12368 1453
rect 13917 1402 13969 1454
rect 14154 1404 14206 1414
rect 14154 1370 14164 1404
rect 14164 1370 14198 1404
rect 14198 1370 14206 1404
rect 14154 1362 14206 1370
rect 14370 1407 14422 1415
rect 14370 1373 14380 1407
rect 14380 1373 14414 1407
rect 14414 1373 14422 1407
rect 14370 1363 14422 1373
rect 14711 1401 14763 1453
rect 16312 1402 16364 1454
rect 16546 1406 16598 1416
rect 16546 1372 16556 1406
rect 16556 1372 16590 1406
rect 16590 1372 16598 1406
rect 16546 1364 16598 1372
rect 1210 1242 1262 1294
rect 1427 1242 1479 1294
rect 1646 1242 1698 1294
rect 1859 1238 1911 1290
rect 2070 1238 2122 1290
rect 4194 1238 4246 1290
rect 4472 1237 4524 1289
rect 5044 1242 5096 1294
rect 5283 1242 5335 1294
rect 7441 1240 7493 1292
rect 7668 1245 7720 1297
rect 7858 1247 7910 1299
rect 8074 1238 8126 1290
rect 10055 1241 10107 1293
rect 10284 1244 10336 1296
rect 10510 1249 10562 1301
rect 10738 1241 10790 1293
rect 10974 1247 11026 1299
rect 11166 1238 11218 1290
rect 12901 1238 12953 1290
rect 13105 1243 13157 1295
rect 13296 1238 13348 1290
rect 13498 1237 13550 1289
rect 13788 1238 13840 1290
rect 14073 1237 14125 1289
rect 15828 1242 15880 1294
rect 16022 1246 16074 1298
rect 16211 1243 16263 1295
rect 16434 1245 16486 1297
rect 265 1097 317 1149
rect 467 1093 519 1145
rect 656 1090 708 1142
rect 885 1091 937 1143
rect 2654 1094 2706 1146
rect 2869 1091 2921 1143
rect 3067 1088 3119 1140
rect 3262 1098 3314 1150
rect 3542 1096 3594 1148
rect 3761 1094 3813 1146
rect 5582 1091 5634 1143
rect 5933 1088 5985 1140
rect 6122 1086 6174 1138
rect 6327 1093 6379 1145
rect 6518 1095 6570 1147
rect 8563 1097 8615 1149
rect 8753 1099 8805 1151
rect 8947 1097 8999 1149
rect 9258 1093 9310 1145
rect 11441 1092 11493 1144
rect 11645 1092 11697 1144
rect 12210 1088 12262 1140
rect 12449 1090 12501 1142
rect 12653 1090 12705 1142
rect 14613 1098 14665 1150
rect 14846 1096 14898 1148
rect 15053 1094 15105 1146
rect 15262 1096 15314 1148
rect 15542 1098 15594 1150
rect 2324 1034 2376 1042
rect 2324 1000 2334 1034
rect 2334 1000 2368 1034
rect 2368 1000 2376 1034
rect 2324 990 2376 1000
rect 4716 1034 4768 1042
rect 4716 1000 4726 1034
rect 4726 1000 4760 1034
rect 4760 1000 4768 1034
rect 4716 990 4768 1000
rect 7108 1034 7160 1042
rect 7108 1000 7118 1034
rect 7118 1000 7152 1034
rect 7152 1000 7160 1034
rect 7108 990 7160 1000
rect 9500 1034 9552 1042
rect 9500 1000 9510 1034
rect 9510 1000 9544 1034
rect 9544 1000 9552 1034
rect 9500 990 9552 1000
rect 11892 1034 11944 1042
rect 11892 1000 11902 1034
rect 11902 1000 11936 1034
rect 11936 1000 11944 1034
rect 11892 990 11944 1000
rect 14284 1034 14336 1042
rect 14284 1000 14294 1034
rect 14294 1000 14328 1034
rect 14328 1000 14336 1034
rect 14284 990 14336 1000
rect 16676 1034 16728 1042
rect 16676 1000 16686 1034
rect 16686 1000 16720 1034
rect 16720 1000 16728 1034
rect 16676 990 16728 1000
rect 2042 955 2094 965
rect 2042 921 2051 955
rect 2051 921 2085 955
rect 2085 921 2094 955
rect 2042 913 2094 921
rect 4434 956 4486 966
rect 4434 922 4443 956
rect 4443 922 4477 956
rect 4477 922 4486 956
rect 4434 914 4486 922
rect 6825 956 6877 966
rect 6825 922 6834 956
rect 6834 922 6868 956
rect 6868 922 6877 956
rect 6825 914 6877 922
rect 9218 957 9270 967
rect 9218 923 9227 957
rect 9227 923 9261 957
rect 9261 923 9270 957
rect 9218 915 9270 923
rect 11609 956 11661 966
rect 11609 922 11618 956
rect 11618 922 11652 956
rect 11652 922 11661 956
rect 11609 914 11661 922
rect 14002 955 14054 965
rect 14002 921 14011 955
rect 14011 921 14045 955
rect 14045 921 14054 955
rect 14002 913 14054 921
rect 16395 957 16447 967
rect 16395 923 16404 957
rect 16404 923 16438 957
rect 16438 923 16447 957
rect 16395 915 16447 923
rect 18 859 70 869
rect 18 825 26 859
rect 26 825 60 859
rect 60 825 70 859
rect 18 817 70 825
rect 357 883 409 894
rect 357 849 366 883
rect 366 849 400 883
rect 400 849 409 883
rect 357 841 409 849
rect 2410 859 2462 869
rect 2410 825 2418 859
rect 2418 825 2452 859
rect 2452 825 2462 859
rect 2410 817 2462 825
rect 2749 883 2801 894
rect 2749 849 2758 883
rect 2758 849 2792 883
rect 2792 849 2801 883
rect 2749 841 2801 849
rect 4802 859 4854 869
rect 4802 825 4810 859
rect 4810 825 4844 859
rect 4844 825 4854 859
rect 4802 817 4854 825
rect 5141 884 5193 895
rect 5141 850 5150 884
rect 5150 850 5184 884
rect 5184 850 5193 884
rect 5141 842 5193 850
rect 7194 859 7246 869
rect 7194 825 7202 859
rect 7202 825 7236 859
rect 7236 825 7246 859
rect 7194 817 7246 825
rect 7533 884 7585 895
rect 7533 850 7542 884
rect 7542 850 7576 884
rect 7576 850 7585 884
rect 7533 842 7585 850
rect 9585 860 9637 870
rect 9585 826 9593 860
rect 9593 826 9627 860
rect 9627 826 9637 860
rect 9585 818 9637 826
rect 9925 883 9977 894
rect 9925 849 9934 883
rect 9934 849 9968 883
rect 9968 849 9977 883
rect 9925 841 9977 849
rect 11977 859 12029 869
rect 11977 825 11985 859
rect 11985 825 12019 859
rect 12019 825 12029 859
rect 11977 817 12029 825
rect 12317 884 12369 895
rect 12317 850 12326 884
rect 12326 850 12360 884
rect 12360 850 12369 884
rect 12317 842 12369 850
rect 14370 860 14422 870
rect 14370 826 14378 860
rect 14378 826 14412 860
rect 14412 826 14422 860
rect 14370 818 14422 826
rect 14710 883 14762 894
rect 14710 849 14719 883
rect 14719 849 14753 883
rect 14753 849 14762 883
rect 14710 841 14762 849
rect 1025 718 1077 770
rect 3418 718 3470 770
rect 5810 718 5862 770
rect 8202 718 8254 770
rect 10593 718 10645 770
rect 12985 718 13037 770
rect 15377 718 15429 770
rect 1192 548 1244 600
rect 1421 560 1473 612
rect 1640 550 1692 602
rect 1832 554 1884 606
rect 2326 552 2378 604
rect 4118 551 4170 603
rect 4511 549 4563 601
rect 4708 557 4760 609
rect 5038 559 5090 611
rect 5234 559 5286 611
rect 7141 552 7193 604
rect 7442 556 7494 608
rect 7648 557 7700 609
rect 7858 553 7910 605
rect 8069 559 8121 611
rect 9949 548 10001 600
rect 10206 555 10258 607
rect 10456 551 10508 603
rect 10727 556 10779 608
rect 10968 559 11020 611
rect 11193 555 11245 607
rect 12900 553 12952 605
rect 13101 554 13153 606
rect 13319 550 13371 602
rect 13526 554 13578 606
rect 13731 553 13783 605
rect 14078 549 14130 601
rect 15830 553 15882 605
rect 16021 556 16073 608
rect 16216 558 16268 610
rect 16663 553 16715 605
rect 47 404 99 456
rect 280 400 332 452
rect 495 407 547 459
rect 713 404 765 456
rect 929 405 981 457
rect 2650 401 2702 453
rect 2840 401 2892 453
rect 3050 404 3102 456
rect 3267 401 3319 453
rect 3562 404 3614 456
rect 3786 409 3838 461
rect 5664 402 5716 454
rect 5964 400 6016 452
rect 6216 404 6268 456
rect 6433 409 6485 461
rect 6634 406 6686 458
rect 8519 397 8571 449
rect 8711 397 8763 449
rect 8911 397 8963 449
rect 9529 405 9581 457
rect 11430 401 11482 453
rect 11686 401 11738 453
rect 11921 401 11973 453
rect 12210 403 12262 455
rect 12400 401 12452 453
rect 12604 403 12656 455
rect 14390 409 14442 461
rect 14632 405 14684 457
rect 14832 404 14884 456
rect 15022 412 15074 464
rect 15243 410 15295 462
rect 15539 405 15591 457
rect 17 342 69 350
rect 17 308 26 342
rect 26 308 60 342
rect 60 308 69 342
rect 2409 342 2461 350
rect 17 298 69 308
rect 297 276 349 286
rect 297 242 306 276
rect 306 242 340 276
rect 340 242 349 276
rect 297 234 349 242
rect 1025 262 1077 314
rect 2409 308 2418 342
rect 2418 308 2452 342
rect 2452 308 2461 342
rect 4802 342 4854 350
rect 2409 298 2461 308
rect 2689 276 2741 286
rect 2689 242 2698 276
rect 2698 242 2732 276
rect 2732 242 2741 276
rect 2689 234 2741 242
rect 2304 205 2358 215
rect 2304 171 2314 205
rect 2314 171 2348 205
rect 2348 171 2358 205
rect 2304 163 2358 171
rect 1959 149 2011 160
rect 1959 115 1968 149
rect 1968 115 2002 149
rect 2002 115 2011 149
rect 1959 107 2011 115
rect 3417 263 3469 315
rect 4802 308 4811 342
rect 4811 308 4845 342
rect 4845 308 4854 342
rect 7193 342 7245 350
rect 4802 298 4854 308
rect 5080 276 5132 286
rect 5080 242 5089 276
rect 5089 242 5123 276
rect 5123 242 5132 276
rect 5080 234 5132 242
rect 4698 205 4752 215
rect 4698 171 4708 205
rect 4708 171 4742 205
rect 4742 171 4752 205
rect 4698 163 4752 171
rect 4351 149 4403 160
rect 4351 115 4360 149
rect 4360 115 4394 149
rect 4394 115 4403 149
rect 4351 107 4403 115
rect 5809 262 5861 314
rect 7193 308 7202 342
rect 7202 308 7236 342
rect 7236 308 7245 342
rect 9585 341 9637 349
rect 7193 298 7245 308
rect 7473 276 7525 286
rect 7473 242 7482 276
rect 7482 242 7516 276
rect 7516 242 7525 276
rect 7473 234 7525 242
rect 7088 207 7142 217
rect 7088 173 7098 207
rect 7098 173 7132 207
rect 7132 173 7142 207
rect 7088 165 7142 173
rect 6742 150 6794 160
rect 6742 116 6751 150
rect 6751 116 6785 150
rect 6785 116 6794 150
rect 6742 108 6794 116
rect 8201 262 8253 314
rect 9585 307 9594 341
rect 9594 307 9628 341
rect 9628 307 9637 341
rect 11978 343 12030 351
rect 9585 297 9637 307
rect 9865 276 9917 286
rect 9865 242 9874 276
rect 9874 242 9908 276
rect 9908 242 9917 276
rect 9865 234 9917 242
rect 9480 205 9534 215
rect 9480 171 9490 205
rect 9490 171 9524 205
rect 9524 171 9534 205
rect 9480 163 9534 171
rect 9135 149 9187 160
rect 9135 115 9144 149
rect 9144 115 9178 149
rect 9178 115 9187 149
rect 9135 107 9187 115
rect 10593 262 10645 314
rect 11978 309 11987 343
rect 11987 309 12021 343
rect 12021 309 12030 343
rect 14369 343 14421 351
rect 11978 299 12030 309
rect 12256 277 12308 287
rect 12256 243 12265 277
rect 12265 243 12299 277
rect 12299 243 12308 277
rect 12256 235 12308 243
rect 11872 207 11926 217
rect 11872 173 11882 207
rect 11882 173 11916 207
rect 11916 173 11926 207
rect 11872 165 11926 173
rect 11526 149 11578 160
rect 11526 115 11535 149
rect 11535 115 11569 149
rect 11569 115 11578 149
rect 11526 107 11578 115
rect 12985 263 13037 315
rect 14369 309 14378 343
rect 14378 309 14412 343
rect 14412 309 14421 343
rect 14369 299 14421 309
rect 14649 276 14701 286
rect 14649 242 14658 276
rect 14658 242 14692 276
rect 14692 242 14701 276
rect 14649 234 14701 242
rect 14264 205 14318 215
rect 14264 171 14274 205
rect 14274 171 14308 205
rect 14308 171 14318 205
rect 14264 163 14318 171
rect 13919 149 13971 160
rect 13919 115 13928 149
rect 13928 115 13962 149
rect 13962 115 13971 149
rect 13919 107 13971 115
rect 15377 263 15429 315
rect 16656 207 16710 217
rect 16656 173 16666 207
rect 16666 173 16700 207
rect 16700 173 16710 207
rect 16656 165 16710 173
rect 16312 149 16364 160
rect 16312 115 16321 149
rect 16321 115 16355 149
rect 16355 115 16364 149
rect 16312 107 16364 115
rect 421 -128 473 -76
rect 620 -131 672 -79
rect 831 -131 883 -79
rect 1037 -131 1089 -79
rect 1265 -133 1317 -81
rect 1509 -133 1561 -81
rect 1739 -131 1791 -79
rect 1945 -131 1997 -79
rect 2163 -126 2215 -74
rect 2366 -132 2418 -80
rect 2574 -129 2626 -77
rect 2837 -133 2889 -81
rect 3045 -132 3097 -80
rect 3255 -135 3307 -83
rect 3455 -129 3507 -77
rect 3658 -132 3710 -80
rect 3868 -132 3920 -80
rect 4069 -131 4121 -79
rect 4285 -130 4337 -78
rect 4566 -132 4618 -80
rect 4786 -137 4838 -85
rect 4991 -136 5043 -84
rect 5212 -130 5264 -78
rect 5417 -137 5469 -85
rect 5626 -136 5678 -84
rect 5843 -136 5895 -84
rect 6057 -131 6109 -79
rect 6252 -133 6304 -81
rect 6447 -136 6499 -84
rect 6649 -133 6701 -81
rect 6933 -132 6985 -80
rect 7132 -131 7184 -79
rect 7335 -129 7387 -77
rect 7600 -132 7652 -80
rect 7798 -133 7850 -81
rect 7987 -131 8039 -79
rect 8199 -131 8251 -79
rect 8416 -131 8468 -79
rect 8621 -135 8673 -83
rect 8826 -135 8878 -83
rect 9034 -130 9086 -78
rect 9317 -131 9369 -79
rect 9510 -133 9562 -81
rect 9736 -135 9788 -83
rect 10001 -135 10053 -83
rect 10195 -131 10247 -79
rect 10393 -140 10445 -88
rect 10597 -132 10649 -80
rect 10817 -129 10869 -77
rect 11032 -133 11084 -81
rect 11260 -130 11312 -78
rect 11464 -133 11516 -81
rect 11702 -131 11754 -79
rect 11895 -130 11947 -78
rect 12092 -135 12144 -83
rect 12348 -132 12400 -80
rect 12587 -136 12639 -84
rect 12820 -140 12872 -88
rect 13041 -135 13093 -83
rect 13232 -135 13284 -83
rect 13460 -133 13512 -81
rect 13657 -138 13709 -86
rect 13869 -138 13921 -86
rect 14096 -135 14148 -83
rect 14285 -134 14337 -82
rect 14511 -133 14563 -81
rect 14765 -133 14817 -81
rect 15009 -136 15061 -84
rect 15239 -137 15291 -85
rect 15497 -134 15549 -82
rect 15707 -134 15759 -82
rect 15932 -134 15984 -82
rect 16151 -137 16203 -85
rect 16497 -133 16549 -81
rect 16696 -136 16748 -84
<< metal2 >>
rect 721 3437 777 3446
rect 721 3372 777 3381
rect 51 2978 107 2987
rect 51 2913 107 2922
rect 17 1834 73 1843
rect 17 1769 73 1778
rect 17 1414 71 1420
rect 17 1362 18 1414
rect 70 1362 71 1414
rect 17 1356 71 1362
rect 23 875 65 1356
rect 17 869 71 875
rect 17 817 18 869
rect 70 817 71 869
rect 17 811 71 817
rect 45 458 101 467
rect 45 393 101 402
rect 17 350 69 356
rect 141 346 183 3300
rect 253 2980 309 2989
rect 253 2915 309 2924
rect 464 2978 520 2987
rect 464 2913 520 2922
rect 654 2978 710 2987
rect 654 2913 710 2922
rect 862 2980 918 2989
rect 862 2915 918 2924
rect 1064 2980 1120 2989
rect 1064 2915 1120 2924
rect 1263 2982 1319 2991
rect 1263 2917 1319 2926
rect 1458 2979 1514 2988
rect 1458 2914 1514 2923
rect 1169 2439 1225 2448
rect 1169 2374 1225 2383
rect 1388 2443 1444 2452
rect 1388 2378 1444 2387
rect 1018 2250 1024 2303
rect 1077 2250 1083 2303
rect 1018 2249 1083 2250
rect 467 2039 474 2091
rect 526 2039 533 2091
rect 257 1832 313 1841
rect 257 1767 313 1776
rect 482 1617 519 2039
rect 579 1831 635 1840
rect 579 1766 635 1775
rect 797 1832 853 1841
rect 797 1767 853 1776
rect 468 1565 475 1617
rect 527 1565 534 1617
rect 349 1400 356 1452
rect 408 1400 414 1452
rect 263 1151 319 1160
rect 263 1086 319 1095
rect 362 894 404 1400
rect 465 1147 521 1156
rect 465 1082 521 1091
rect 654 1144 710 1153
rect 654 1079 710 1088
rect 883 1145 939 1154
rect 883 1080 939 1089
rect 351 841 357 894
rect 409 841 416 894
rect 351 840 416 841
rect 1030 776 1072 2249
rect 1562 1603 1604 3300
rect 1659 2981 1715 2990
rect 1659 2916 1715 2925
rect 1876 2979 1932 2988
rect 1876 2914 1932 2923
rect 1671 2443 1727 2452
rect 1671 2378 1727 2387
rect 1880 2443 1936 2452
rect 1880 2378 1936 2387
rect 1729 2039 1736 2091
rect 1788 2039 1795 2091
rect 1744 1617 1781 2039
rect 1551 1550 1557 1603
rect 1609 1550 1616 1603
rect 1730 1565 1737 1617
rect 1789 1565 1796 1617
rect 1551 1549 1616 1550
rect 1964 1453 2006 3300
rect 2150 2982 2206 2991
rect 2150 2917 2206 2926
rect 2151 2441 2207 2450
rect 2151 2376 2207 2385
rect 1950 1401 1957 1453
rect 2009 1401 2015 1453
rect 1208 1296 1264 1305
rect 1208 1231 1264 1240
rect 1425 1296 1481 1305
rect 1425 1231 1481 1240
rect 1644 1296 1700 1305
rect 1644 1231 1700 1240
rect 1857 1292 1913 1301
rect 1857 1227 1913 1236
rect 1024 770 1078 776
rect 1024 718 1025 770
rect 1077 718 1078 770
rect 1024 712 1078 718
rect 278 454 334 463
rect 278 389 334 398
rect 493 461 549 470
rect 493 396 549 405
rect 711 458 767 467
rect 711 393 767 402
rect 927 459 983 468
rect 927 394 983 403
rect 69 304 183 346
rect 1030 314 1072 712
rect 1419 614 1475 623
rect 1190 602 1246 611
rect 1419 549 1475 558
rect 1638 604 1694 613
rect 1190 537 1246 546
rect 1638 539 1694 548
rect 1830 608 1886 617
rect 1830 543 1886 552
rect 17 292 69 298
rect 297 286 349 292
rect 1019 262 1025 314
rect 1077 262 1083 314
rect 297 228 349 234
rect 301 -343 343 228
rect 1964 160 2006 1401
rect 2188 1362 2194 1414
rect 2246 1362 2254 1414
rect 2068 1292 2124 1301
rect 2068 1227 2124 1236
rect 2042 965 2094 971
rect 2042 907 2094 913
rect 1953 107 1959 160
rect 2011 107 2018 160
rect 1953 106 2018 107
rect 419 -74 475 -65
rect 419 -139 475 -130
rect 618 -77 674 -68
rect 618 -142 674 -133
rect 829 -77 885 -68
rect 829 -142 885 -133
rect 1035 -77 1091 -68
rect 1035 -142 1091 -133
rect 1263 -79 1319 -70
rect 1263 -144 1319 -135
rect 1507 -79 1563 -70
rect 1507 -144 1563 -135
rect 1737 -77 1793 -68
rect 1737 -142 1793 -133
rect 1943 -77 1999 -68
rect 1943 -142 1999 -133
rect 2046 -343 2088 907
rect 2200 215 2242 1362
rect 2330 1048 2372 3300
rect 2427 2975 2483 2984
rect 2427 2910 2483 2919
rect 2409 1414 2463 1420
rect 2409 1362 2410 1414
rect 2462 1362 2463 1414
rect 2409 1356 2463 1362
rect 2324 1042 2376 1048
rect 2324 984 2376 990
rect 2415 875 2457 1356
rect 2409 869 2463 875
rect 2409 817 2410 869
rect 2462 817 2463 869
rect 2409 811 2463 817
rect 2324 606 2380 615
rect 2324 541 2380 550
rect 2409 350 2461 356
rect 2533 346 2575 3300
rect 2650 2978 2706 2987
rect 2650 2913 2706 2922
rect 2882 2977 2938 2986
rect 2882 2912 2938 2921
rect 2860 2622 2866 2674
rect 2918 2622 2924 2674
rect 2866 2302 2918 2622
rect 2860 2250 2866 2302
rect 2918 2250 2924 2302
rect 3412 2256 3418 2309
rect 3471 2256 3477 2309
rect 3412 2255 3477 2256
rect 2860 2038 2867 2090
rect 2919 2038 2926 2090
rect 2701 1836 2757 1845
rect 2701 1771 2757 1780
rect 2875 1616 2912 2038
rect 3026 1838 3082 1847
rect 3026 1773 3082 1782
rect 3294 1838 3350 1847
rect 3294 1773 3350 1782
rect 2861 1564 2868 1616
rect 2920 1564 2927 1616
rect 2741 1400 2748 1452
rect 2800 1400 2806 1452
rect 2652 1148 2708 1157
rect 2652 1083 2708 1092
rect 2754 894 2796 1400
rect 2867 1145 2923 1154
rect 3260 1152 3316 1161
rect 2867 1080 2923 1089
rect 3065 1142 3121 1151
rect 3260 1087 3316 1096
rect 3065 1077 3121 1086
rect 2743 841 2749 894
rect 2801 841 2808 894
rect 2743 840 2808 841
rect 3424 776 3466 2255
rect 3560 1838 3616 1847
rect 3560 1773 3616 1782
rect 3800 1836 3856 1845
rect 3800 1771 3856 1780
rect 3954 1602 3996 3300
rect 4226 2439 4282 2448
rect 4226 2374 4282 2383
rect 4121 2039 4128 2091
rect 4180 2039 4187 2091
rect 4136 1617 4173 2039
rect 3943 1549 3949 1602
rect 4001 1549 4008 1602
rect 4122 1565 4129 1617
rect 4181 1565 4188 1617
rect 3943 1548 4008 1549
rect 4356 1453 4398 3300
rect 4518 2974 4574 2983
rect 4518 2909 4574 2918
rect 4475 2442 4531 2451
rect 4475 2377 4531 2386
rect 4342 1401 4349 1453
rect 4401 1401 4407 1453
rect 4192 1292 4248 1301
rect 4192 1227 4248 1236
rect 3540 1150 3596 1159
rect 3540 1085 3596 1094
rect 3759 1148 3815 1157
rect 3759 1083 3815 1092
rect 3417 770 3471 776
rect 3417 718 3418 770
rect 3470 718 3471 770
rect 3417 712 3471 718
rect 2648 455 2704 464
rect 2648 390 2704 399
rect 2838 455 2894 464
rect 2838 390 2894 399
rect 3048 458 3104 467
rect 3048 393 3104 402
rect 3265 455 3321 464
rect 3265 390 3321 399
rect 2461 304 2575 346
rect 3422 315 3464 712
rect 4116 605 4172 614
rect 4116 540 4172 549
rect 3560 458 3616 467
rect 3560 393 3616 402
rect 3784 463 3840 472
rect 3784 398 3840 407
rect 2409 292 2461 298
rect 2689 286 2741 292
rect 3411 263 3417 315
rect 3469 263 3475 315
rect 2689 228 2741 234
rect 2200 175 2304 215
rect 2298 163 2304 175
rect 2358 163 2364 215
rect 2161 -72 2217 -63
rect 2161 -137 2217 -128
rect 2364 -78 2420 -69
rect 2364 -143 2420 -134
rect 2572 -75 2628 -66
rect 2572 -140 2628 -131
rect 2693 -343 2735 228
rect 4356 160 4398 1401
rect 4582 1362 4588 1414
rect 4640 1362 4648 1414
rect 4470 1291 4526 1300
rect 4470 1226 4526 1235
rect 4434 966 4486 972
rect 4434 908 4486 914
rect 4345 107 4351 160
rect 4403 107 4410 160
rect 4345 106 4410 107
rect 2835 -79 2891 -70
rect 2835 -144 2891 -135
rect 3043 -78 3099 -69
rect 3043 -143 3099 -134
rect 3253 -81 3309 -72
rect 3253 -146 3309 -137
rect 3453 -75 3509 -66
rect 3453 -140 3509 -131
rect 3656 -78 3712 -69
rect 3656 -143 3712 -134
rect 3866 -78 3922 -69
rect 3866 -143 3922 -134
rect 4067 -77 4123 -68
rect 4067 -142 4123 -133
rect 4283 -76 4339 -67
rect 4283 -141 4339 -132
rect 4438 -343 4480 908
rect 4509 603 4565 612
rect 4509 538 4565 547
rect 4594 215 4636 1362
rect 4722 1048 4764 3300
rect 4826 2975 4882 2984
rect 4826 2910 4882 2919
rect 4819 2428 4875 2437
rect 4819 2363 4875 2372
rect 4801 1414 4855 1420
rect 4801 1362 4802 1414
rect 4854 1362 4855 1414
rect 4801 1356 4855 1362
rect 4716 1042 4768 1048
rect 4716 984 4768 990
rect 4807 875 4849 1356
rect 4801 869 4855 875
rect 4801 817 4802 869
rect 4854 817 4855 869
rect 4801 811 4855 817
rect 4706 611 4762 620
rect 4706 546 4762 555
rect 4802 350 4854 356
rect 4926 346 4968 3300
rect 5026 2976 5082 2985
rect 5026 2911 5082 2920
rect 5245 2975 5301 2984
rect 5245 2910 5301 2919
rect 5491 2974 5547 2983
rect 5491 2909 5547 2918
rect 5699 2976 5755 2985
rect 5699 2911 5755 2920
rect 5901 2977 5957 2986
rect 5901 2912 5957 2921
rect 6094 2976 6150 2985
rect 6094 2911 6150 2920
rect 5073 2434 5129 2443
rect 5073 2369 5129 2378
rect 5302 2434 5358 2443
rect 5302 2369 5358 2378
rect 5803 2256 5809 2309
rect 5862 2256 5868 2309
rect 5803 2255 5868 2256
rect 5252 2038 5259 2090
rect 5311 2038 5318 2090
rect 5267 1616 5304 2038
rect 5594 1839 5650 1848
rect 5594 1774 5650 1783
rect 5253 1564 5260 1616
rect 5312 1564 5319 1616
rect 5132 1401 5139 1453
rect 5191 1401 5197 1453
rect 5042 1296 5098 1305
rect 5042 1231 5098 1240
rect 5146 895 5188 1401
rect 5281 1296 5337 1305
rect 5281 1231 5337 1240
rect 5580 1145 5636 1154
rect 5580 1080 5636 1089
rect 5135 842 5141 895
rect 5193 842 5200 895
rect 5135 841 5200 842
rect 5815 776 5857 2255
rect 5960 1842 6016 1851
rect 5960 1777 6016 1786
rect 6204 1842 6260 1851
rect 6204 1777 6260 1786
rect 6344 1602 6386 3300
rect 6466 2975 6522 2984
rect 6466 2910 6522 2919
rect 6655 2973 6711 2982
rect 6655 2908 6711 2917
rect 6512 2040 6519 2092
rect 6571 2040 6578 2092
rect 6527 1853 6564 2040
rect 6521 1819 6564 1853
rect 6527 1618 6564 1819
rect 6627 1833 6683 1842
rect 6627 1768 6683 1777
rect 6333 1549 6339 1602
rect 6391 1549 6398 1602
rect 6513 1566 6520 1618
rect 6572 1566 6579 1618
rect 6333 1548 6398 1549
rect 6747 1454 6789 3300
rect 6945 2973 7001 2982
rect 6945 2908 7001 2917
rect 7020 2439 7076 2448
rect 7020 2374 7076 2383
rect 6733 1402 6740 1454
rect 6792 1402 6798 1454
rect 5931 1142 5987 1151
rect 5931 1077 5987 1086
rect 6120 1140 6176 1149
rect 6120 1075 6176 1084
rect 6325 1147 6381 1156
rect 6325 1082 6381 1091
rect 6516 1149 6572 1158
rect 6516 1084 6572 1093
rect 5809 770 5863 776
rect 5809 718 5810 770
rect 5862 718 5863 770
rect 5809 712 5863 718
rect 5036 613 5092 622
rect 5036 548 5092 557
rect 5232 613 5288 622
rect 5232 548 5288 557
rect 5662 456 5718 465
rect 5662 391 5718 400
rect 4854 304 4968 346
rect 5814 314 5856 712
rect 5962 454 6018 463
rect 5962 389 6018 398
rect 6214 458 6270 467
rect 6214 393 6270 402
rect 6431 463 6487 472
rect 6431 398 6487 407
rect 6632 460 6688 469
rect 6632 395 6688 404
rect 4802 292 4854 298
rect 5080 286 5132 292
rect 5803 262 5809 314
rect 5861 262 5867 314
rect 5080 228 5132 234
rect 4594 175 4698 215
rect 4692 163 4698 175
rect 4752 163 4758 215
rect 4564 -78 4620 -69
rect 4564 -143 4620 -134
rect 4784 -83 4840 -74
rect 4784 -148 4840 -139
rect 4989 -82 5045 -73
rect 4989 -147 5045 -138
rect 5084 -343 5126 228
rect 6747 161 6789 1402
rect 6972 1364 6978 1416
rect 7030 1364 7038 1416
rect 6825 966 6877 972
rect 6825 908 6877 914
rect 6736 160 6801 161
rect 6736 108 6742 160
rect 6794 108 6801 160
rect 6736 107 6801 108
rect 5210 -76 5266 -67
rect 5210 -141 5266 -132
rect 5415 -83 5471 -74
rect 5415 -148 5471 -139
rect 5624 -82 5680 -73
rect 5624 -147 5680 -138
rect 5841 -82 5897 -73
rect 5841 -147 5897 -138
rect 6055 -77 6111 -68
rect 6055 -142 6111 -133
rect 6250 -79 6306 -70
rect 6250 -144 6306 -135
rect 6445 -82 6501 -73
rect 6445 -147 6501 -138
rect 6647 -79 6703 -70
rect 6647 -144 6703 -135
rect 6829 -343 6871 908
rect 6984 217 7026 1364
rect 7114 1048 7156 3300
rect 7218 2975 7274 2984
rect 7218 2910 7274 2919
rect 7224 2441 7280 2450
rect 7224 2376 7280 2385
rect 7193 1414 7247 1420
rect 7193 1362 7194 1414
rect 7246 1362 7247 1414
rect 7193 1356 7247 1362
rect 7108 1042 7160 1048
rect 7108 984 7160 990
rect 7199 875 7241 1356
rect 7193 869 7247 875
rect 7193 817 7194 869
rect 7246 817 7247 869
rect 7193 811 7247 817
rect 7139 606 7195 615
rect 7139 541 7195 550
rect 7193 350 7245 356
rect 7317 346 7359 3300
rect 7421 2622 7427 2674
rect 7479 2622 7485 2674
rect 7427 2090 7479 2622
rect 7547 2439 7603 2448
rect 7547 2374 7603 2383
rect 8194 2256 8200 2309
rect 8253 2256 8259 2309
rect 8194 2255 8259 2256
rect 7421 2038 7427 2090
rect 7479 2038 7485 2090
rect 7644 2039 7651 2091
rect 7703 2039 7710 2091
rect 7659 1617 7696 2039
rect 7645 1565 7652 1617
rect 7704 1565 7711 1617
rect 7525 1400 7532 1452
rect 7584 1400 7590 1452
rect 7439 1294 7495 1303
rect 7439 1229 7495 1238
rect 7538 895 7580 1400
rect 7666 1299 7722 1308
rect 7666 1234 7722 1243
rect 7856 1301 7912 1310
rect 7856 1236 7912 1245
rect 8072 1292 8128 1301
rect 8072 1227 8128 1236
rect 7527 842 7533 895
rect 7585 842 7592 895
rect 7527 841 7592 842
rect 8206 776 8248 2255
rect 8570 1835 8626 1844
rect 8570 1770 8626 1779
rect 8738 1603 8780 3300
rect 8905 2040 8912 2092
rect 8964 2040 8971 2092
rect 8822 1832 8878 1841
rect 8822 1767 8878 1776
rect 8920 1618 8957 2040
rect 9028 1840 9084 1849
rect 9028 1775 9084 1784
rect 8727 1550 8733 1603
rect 8785 1550 8792 1603
rect 8906 1566 8913 1618
rect 8965 1566 8972 1618
rect 8727 1549 8792 1550
rect 9140 1453 9182 3300
rect 9311 1834 9367 1843
rect 9311 1769 9367 1778
rect 9126 1401 9133 1453
rect 9185 1401 9191 1453
rect 8561 1151 8617 1160
rect 8561 1086 8617 1095
rect 8751 1153 8807 1162
rect 8751 1088 8807 1097
rect 8945 1151 9001 1160
rect 8945 1086 9001 1095
rect 8201 770 8255 776
rect 8201 718 8202 770
rect 8254 718 8255 770
rect 8201 712 8255 718
rect 7440 610 7496 619
rect 7440 545 7496 554
rect 7646 611 7702 620
rect 7646 546 7702 555
rect 7856 607 7912 616
rect 7856 542 7912 551
rect 8067 613 8123 622
rect 8067 548 8123 557
rect 7245 304 7359 346
rect 8206 314 8248 712
rect 8517 451 8573 460
rect 8517 386 8573 395
rect 8709 451 8765 460
rect 8709 386 8765 395
rect 8909 451 8965 460
rect 8909 386 8965 395
rect 7193 292 7245 298
rect 7473 286 7525 292
rect 8195 262 8201 314
rect 8253 262 8259 314
rect 7473 228 7525 234
rect 6984 177 7088 217
rect 7082 165 7088 177
rect 7142 165 7148 217
rect 6931 -78 6987 -69
rect 6931 -143 6987 -134
rect 7130 -77 7186 -68
rect 7130 -142 7186 -133
rect 7333 -75 7389 -66
rect 7333 -140 7389 -131
rect 7477 -343 7519 228
rect 9140 160 9182 1401
rect 9364 1362 9370 1414
rect 9422 1362 9430 1414
rect 9256 1147 9312 1156
rect 9256 1082 9312 1091
rect 9218 967 9270 973
rect 9218 909 9270 915
rect 9129 107 9135 160
rect 9187 107 9194 160
rect 9129 106 9194 107
rect 7598 -78 7654 -69
rect 7598 -143 7654 -134
rect 7796 -79 7852 -70
rect 7796 -144 7852 -135
rect 7985 -77 8041 -68
rect 7985 -142 8041 -133
rect 8197 -77 8253 -68
rect 8197 -142 8253 -133
rect 8414 -77 8470 -68
rect 8414 -142 8470 -133
rect 8619 -81 8675 -72
rect 8619 -146 8675 -137
rect 8824 -81 8880 -72
rect 8824 -146 8880 -137
rect 9032 -76 9088 -67
rect 9032 -141 9088 -132
rect 9222 -343 9264 909
rect 9376 215 9418 1362
rect 9506 1048 9548 3300
rect 9609 1835 9665 1844
rect 9609 1770 9665 1779
rect 9584 1415 9638 1421
rect 9584 1363 9585 1415
rect 9637 1363 9638 1415
rect 9584 1357 9638 1363
rect 9500 1042 9552 1048
rect 9500 984 9552 990
rect 9590 876 9632 1357
rect 9584 870 9638 876
rect 9584 818 9585 870
rect 9637 818 9638 870
rect 9584 812 9638 818
rect 9527 459 9583 468
rect 9527 394 9583 403
rect 9585 349 9637 355
rect 9709 345 9751 3300
rect 10586 2256 10592 2309
rect 10645 2256 10651 2309
rect 10586 2255 10651 2256
rect 10035 2038 10042 2090
rect 10094 2038 10101 2090
rect 10050 1616 10087 2038
rect 10036 1564 10043 1616
rect 10095 1564 10102 1616
rect 9917 1401 9924 1453
rect 9976 1401 9982 1453
rect 9930 894 9972 1401
rect 10053 1295 10109 1304
rect 10053 1230 10109 1239
rect 10282 1298 10338 1307
rect 10282 1233 10338 1242
rect 10508 1303 10564 1312
rect 10508 1238 10564 1247
rect 9919 841 9925 894
rect 9977 841 9984 894
rect 9919 840 9984 841
rect 10598 776 10640 2255
rect 11130 1602 11172 3300
rect 11298 2040 11305 2092
rect 11357 2040 11364 2092
rect 11313 1618 11350 2040
rect 11441 1836 11497 1845
rect 11441 1771 11497 1780
rect 11119 1549 11125 1602
rect 11177 1549 11184 1602
rect 11299 1566 11306 1618
rect 11358 1566 11365 1618
rect 11119 1548 11184 1549
rect 11531 1454 11573 3300
rect 11651 1838 11707 1847
rect 11651 1773 11707 1782
rect 11518 1402 11525 1454
rect 11577 1402 11583 1454
rect 10736 1295 10792 1304
rect 10736 1230 10792 1239
rect 10972 1301 11028 1310
rect 10972 1236 11028 1245
rect 11164 1292 11220 1301
rect 11164 1227 11220 1236
rect 11439 1146 11495 1155
rect 11439 1081 11495 1090
rect 10592 770 10646 776
rect 10592 718 10593 770
rect 10645 718 10646 770
rect 10592 710 10646 718
rect 9947 602 10003 611
rect 9947 537 10003 546
rect 10204 609 10260 618
rect 10204 544 10260 553
rect 10454 605 10510 614
rect 10454 540 10510 549
rect 9637 303 9751 345
rect 10598 314 10640 710
rect 10725 610 10781 619
rect 10725 545 10781 554
rect 10966 613 11022 622
rect 10966 548 11022 557
rect 11191 609 11247 618
rect 11191 544 11247 553
rect 11428 455 11484 464
rect 11428 390 11484 399
rect 9585 291 9637 297
rect 9865 286 9917 292
rect 10587 262 10593 314
rect 10645 262 10651 314
rect 9865 228 9917 234
rect 9376 175 9480 215
rect 9474 163 9480 175
rect 9534 163 9540 215
rect 9315 -77 9371 -68
rect 9315 -142 9371 -133
rect 9508 -79 9564 -70
rect 9508 -144 9564 -135
rect 9734 -81 9790 -72
rect 9734 -146 9790 -137
rect 9869 -343 9911 228
rect 11531 160 11573 1402
rect 11756 1364 11762 1416
rect 11814 1364 11822 1416
rect 11643 1146 11699 1155
rect 11643 1081 11699 1090
rect 11609 966 11661 972
rect 11609 908 11661 914
rect 11520 107 11526 160
rect 11578 107 11585 160
rect 11520 106 11585 107
rect 9999 -81 10055 -72
rect 9999 -146 10055 -137
rect 10193 -77 10249 -68
rect 10193 -142 10249 -133
rect 10391 -86 10447 -77
rect 10391 -151 10447 -142
rect 10595 -78 10651 -69
rect 10595 -143 10651 -134
rect 10815 -75 10871 -66
rect 10815 -140 10871 -131
rect 11030 -79 11086 -70
rect 11030 -144 11086 -135
rect 11258 -76 11314 -67
rect 11258 -141 11314 -132
rect 11462 -79 11518 -70
rect 11462 -144 11518 -135
rect 11613 -343 11655 908
rect 11684 455 11740 464
rect 11684 390 11740 399
rect 11768 217 11810 1364
rect 11898 1048 11940 3300
rect 12002 1836 12058 1845
rect 12002 1771 12058 1780
rect 11976 1414 12030 1420
rect 11976 1362 11977 1414
rect 12029 1362 12030 1414
rect 11976 1356 12030 1362
rect 11892 1042 11944 1048
rect 11892 984 11944 990
rect 11982 875 12024 1356
rect 11976 869 12030 875
rect 11976 817 11977 869
rect 12029 817 12030 869
rect 11976 811 12030 817
rect 11919 455 11975 464
rect 11919 390 11975 399
rect 11978 351 12030 357
rect 12102 347 12144 3300
rect 12977 2256 12983 2309
rect 13036 2256 13042 2309
rect 12977 2255 13042 2256
rect 12427 2037 12434 2089
rect 12486 2037 12493 2089
rect 12282 1836 12338 1845
rect 12282 1771 12338 1780
rect 12442 1615 12479 2037
rect 12599 1835 12655 1844
rect 12599 1770 12655 1779
rect 12428 1563 12435 1615
rect 12487 1563 12494 1615
rect 12309 1401 12316 1453
rect 12368 1401 12374 1453
rect 12208 1142 12264 1151
rect 12208 1077 12264 1086
rect 12322 895 12364 1401
rect 12899 1292 12955 1301
rect 12899 1227 12955 1236
rect 12447 1144 12503 1153
rect 12447 1079 12503 1088
rect 12651 1144 12707 1153
rect 12651 1079 12707 1088
rect 12311 842 12317 895
rect 12369 842 12376 895
rect 12311 841 12376 842
rect 12989 776 13031 2255
rect 13519 1602 13561 3300
rect 13687 2040 13694 2092
rect 13746 2040 13753 2092
rect 13702 1618 13739 2040
rect 13508 1549 13514 1602
rect 13566 1549 13573 1602
rect 13688 1566 13695 1618
rect 13747 1566 13754 1618
rect 13508 1548 13573 1549
rect 13924 1454 13966 3300
rect 13910 1402 13917 1454
rect 13969 1402 13975 1454
rect 13103 1297 13159 1306
rect 13103 1232 13159 1241
rect 13294 1292 13350 1301
rect 13294 1227 13350 1236
rect 13496 1291 13552 1300
rect 13496 1226 13552 1235
rect 13786 1292 13842 1301
rect 13786 1227 13842 1236
rect 12984 770 13038 776
rect 12984 718 12985 770
rect 13037 718 13038 770
rect 12984 712 13038 718
rect 12898 607 12954 616
rect 12898 542 12954 551
rect 12208 457 12264 466
rect 12208 392 12264 401
rect 12398 455 12454 464
rect 12398 390 12454 399
rect 12602 457 12658 466
rect 12602 392 12658 401
rect 12030 305 12144 347
rect 12990 315 13032 712
rect 13099 608 13155 617
rect 13099 543 13155 552
rect 13317 604 13373 613
rect 13317 539 13373 548
rect 13524 608 13580 617
rect 13524 543 13580 552
rect 13729 607 13785 616
rect 13729 542 13785 551
rect 11978 293 12030 299
rect 12256 287 12308 293
rect 12979 263 12985 315
rect 13037 263 13043 315
rect 12256 229 12308 235
rect 11768 177 11872 217
rect 11866 165 11872 177
rect 11926 165 11932 217
rect 11700 -77 11756 -68
rect 11700 -142 11756 -133
rect 11893 -76 11949 -67
rect 11893 -141 11949 -132
rect 12090 -81 12146 -72
rect 12090 -146 12146 -137
rect 12260 -343 12302 229
rect 13924 160 13966 1402
rect 14148 1362 14154 1414
rect 14206 1362 14214 1414
rect 14071 1291 14127 1300
rect 14071 1226 14127 1235
rect 14002 965 14054 971
rect 14002 907 14054 913
rect 13913 107 13919 160
rect 13971 107 13978 160
rect 13913 106 13978 107
rect 12346 -78 12402 -69
rect 12346 -143 12402 -134
rect 12585 -82 12641 -73
rect 12585 -147 12641 -138
rect 12818 -86 12874 -77
rect 12818 -151 12874 -142
rect 13039 -81 13095 -72
rect 13039 -146 13095 -137
rect 13230 -81 13286 -72
rect 13230 -146 13286 -137
rect 13458 -79 13514 -70
rect 13458 -144 13514 -135
rect 13655 -84 13711 -75
rect 13655 -149 13711 -140
rect 13867 -84 13923 -75
rect 13867 -149 13923 -140
rect 14006 -343 14048 907
rect 14076 603 14132 612
rect 14076 538 14132 547
rect 14160 215 14202 1362
rect 14290 1048 14332 3300
rect 14389 1833 14445 1842
rect 14389 1768 14445 1777
rect 14369 1415 14423 1421
rect 14369 1363 14370 1415
rect 14422 1363 14423 1415
rect 14369 1357 14423 1363
rect 14284 1042 14336 1048
rect 14284 984 14336 990
rect 14375 876 14417 1357
rect 14369 870 14423 876
rect 14369 818 14370 870
rect 14422 818 14423 870
rect 14369 812 14423 818
rect 14388 463 14444 472
rect 14388 398 14444 407
rect 14369 351 14421 357
rect 14493 347 14535 3300
rect 15370 2256 15376 2309
rect 15429 2256 15435 2309
rect 15370 2255 15435 2256
rect 14819 2038 14826 2090
rect 14878 2038 14885 2090
rect 14684 1833 14740 1842
rect 14684 1768 14740 1777
rect 14834 1616 14871 2038
rect 14971 1833 15027 1842
rect 14971 1768 15027 1777
rect 15261 1833 15317 1842
rect 15261 1768 15317 1777
rect 14820 1564 14827 1616
rect 14879 1564 14886 1616
rect 14704 1401 14711 1453
rect 14763 1401 14769 1453
rect 14611 1152 14667 1161
rect 14611 1087 14667 1096
rect 14715 894 14757 1401
rect 14844 1150 14900 1159
rect 14844 1085 14900 1094
rect 15051 1148 15107 1157
rect 15051 1083 15107 1092
rect 15260 1150 15316 1159
rect 15260 1085 15316 1094
rect 14704 841 14710 894
rect 14762 841 14769 894
rect 14704 840 14769 841
rect 15382 776 15424 2255
rect 15545 1836 15601 1845
rect 15545 1771 15601 1780
rect 15914 1603 15956 3300
rect 16082 2040 16089 2092
rect 16141 2040 16148 2092
rect 16097 1618 16134 2040
rect 15903 1550 15909 1603
rect 15961 1550 15968 1603
rect 16083 1566 16090 1618
rect 16142 1566 16149 1618
rect 15903 1549 15968 1550
rect 16317 1454 16359 3300
rect 16305 1402 16312 1454
rect 16364 1402 16370 1454
rect 15826 1296 15882 1305
rect 15826 1231 15882 1240
rect 16020 1300 16076 1309
rect 16020 1235 16076 1244
rect 16209 1297 16265 1306
rect 16209 1232 16265 1241
rect 15540 1152 15596 1161
rect 15540 1087 15596 1096
rect 15376 770 15430 776
rect 15376 718 15377 770
rect 15429 718 15430 770
rect 15376 712 15430 718
rect 14630 459 14686 468
rect 14630 394 14686 403
rect 14830 458 14886 467
rect 14830 393 14886 402
rect 15020 466 15076 475
rect 15020 401 15076 410
rect 15241 464 15297 473
rect 15241 399 15297 408
rect 14421 305 14535 347
rect 15382 315 15424 712
rect 15828 607 15884 616
rect 15828 542 15884 551
rect 16019 610 16075 619
rect 16019 545 16075 554
rect 16214 612 16270 621
rect 16214 547 16270 556
rect 15537 459 15593 468
rect 15537 394 15593 403
rect 14369 293 14421 299
rect 14649 286 14701 292
rect 15371 263 15377 315
rect 15429 263 15435 315
rect 14649 228 14701 234
rect 14160 175 14264 215
rect 14258 163 14264 175
rect 14318 163 14324 215
rect 14094 -81 14150 -72
rect 14094 -146 14150 -137
rect 14283 -80 14339 -71
rect 14283 -145 14339 -136
rect 14509 -79 14565 -70
rect 14509 -144 14565 -135
rect 14653 -343 14695 228
rect 16317 160 16359 1402
rect 16540 1364 16546 1416
rect 16598 1364 16606 1416
rect 16432 1299 16488 1308
rect 16432 1234 16488 1243
rect 16395 967 16447 973
rect 16395 909 16447 915
rect 16306 107 16312 160
rect 16364 107 16371 160
rect 16306 106 16371 107
rect 14763 -79 14819 -70
rect 14763 -144 14819 -135
rect 15007 -82 15063 -73
rect 15007 -147 15063 -138
rect 15237 -83 15293 -74
rect 15237 -148 15293 -139
rect 15495 -80 15551 -71
rect 15495 -145 15551 -136
rect 15705 -80 15761 -71
rect 15705 -145 15761 -136
rect 15930 -80 15986 -71
rect 15930 -145 15986 -136
rect 16149 -83 16205 -74
rect 16149 -148 16205 -139
rect 16399 -343 16441 909
rect 16552 217 16594 1364
rect 16682 1048 16724 3300
rect 16676 1042 16728 1048
rect 16676 984 16728 990
rect 16661 607 16717 616
rect 16661 542 16717 551
rect 16552 177 16656 217
rect 16650 165 16656 177
rect 16710 165 16716 217
rect 16495 -79 16551 -70
rect 16495 -144 16551 -135
rect 16694 -82 16750 -73
rect 16694 -147 16750 -138
<< via2 >>
rect 721 3435 777 3437
rect 721 3383 723 3435
rect 723 3383 775 3435
rect 775 3383 777 3435
rect 721 3381 777 3383
rect 51 2976 107 2978
rect 51 2924 53 2976
rect 53 2924 105 2976
rect 105 2924 107 2976
rect 51 2922 107 2924
rect 17 1832 73 1834
rect 17 1780 19 1832
rect 19 1780 71 1832
rect 71 1780 73 1832
rect 17 1778 73 1780
rect 45 456 101 458
rect 45 404 47 456
rect 47 404 99 456
rect 99 404 101 456
rect 45 402 101 404
rect 253 2978 309 2980
rect 253 2926 255 2978
rect 255 2926 307 2978
rect 307 2926 309 2978
rect 253 2924 309 2926
rect 464 2976 520 2978
rect 464 2924 466 2976
rect 466 2924 518 2976
rect 518 2924 520 2976
rect 464 2922 520 2924
rect 654 2976 710 2978
rect 654 2924 656 2976
rect 656 2924 708 2976
rect 708 2924 710 2976
rect 654 2922 710 2924
rect 862 2978 918 2980
rect 862 2926 864 2978
rect 864 2926 916 2978
rect 916 2926 918 2978
rect 862 2924 918 2926
rect 1064 2978 1120 2980
rect 1064 2926 1066 2978
rect 1066 2926 1118 2978
rect 1118 2926 1120 2978
rect 1064 2924 1120 2926
rect 1263 2980 1319 2982
rect 1263 2928 1265 2980
rect 1265 2928 1317 2980
rect 1317 2928 1319 2980
rect 1263 2926 1319 2928
rect 1458 2977 1514 2979
rect 1458 2925 1460 2977
rect 1460 2925 1512 2977
rect 1512 2925 1514 2977
rect 1458 2923 1514 2925
rect 1169 2437 1225 2439
rect 1169 2385 1171 2437
rect 1171 2385 1223 2437
rect 1223 2385 1225 2437
rect 1169 2383 1225 2385
rect 1388 2441 1444 2443
rect 1388 2389 1390 2441
rect 1390 2389 1442 2441
rect 1442 2389 1444 2441
rect 1388 2387 1444 2389
rect 257 1830 313 1832
rect 257 1778 259 1830
rect 259 1778 311 1830
rect 311 1778 313 1830
rect 257 1776 313 1778
rect 579 1829 635 1831
rect 579 1777 581 1829
rect 581 1777 633 1829
rect 633 1777 635 1829
rect 579 1775 635 1777
rect 797 1830 853 1832
rect 797 1778 799 1830
rect 799 1778 851 1830
rect 851 1778 853 1830
rect 797 1776 853 1778
rect 263 1149 319 1151
rect 263 1097 265 1149
rect 265 1097 317 1149
rect 317 1097 319 1149
rect 263 1095 319 1097
rect 465 1145 521 1147
rect 465 1093 467 1145
rect 467 1093 519 1145
rect 519 1093 521 1145
rect 465 1091 521 1093
rect 654 1142 710 1144
rect 654 1090 656 1142
rect 656 1090 708 1142
rect 708 1090 710 1142
rect 654 1088 710 1090
rect 883 1143 939 1145
rect 883 1091 885 1143
rect 885 1091 937 1143
rect 937 1091 939 1143
rect 883 1089 939 1091
rect 1659 2979 1715 2981
rect 1659 2927 1661 2979
rect 1661 2927 1713 2979
rect 1713 2927 1715 2979
rect 1659 2925 1715 2927
rect 1876 2977 1932 2979
rect 1876 2925 1878 2977
rect 1878 2925 1930 2977
rect 1930 2925 1932 2977
rect 1876 2923 1932 2925
rect 1671 2441 1727 2443
rect 1671 2389 1673 2441
rect 1673 2389 1725 2441
rect 1725 2389 1727 2441
rect 1671 2387 1727 2389
rect 1880 2441 1936 2443
rect 1880 2389 1882 2441
rect 1882 2389 1934 2441
rect 1934 2389 1936 2441
rect 1880 2387 1936 2389
rect 2150 2980 2206 2982
rect 2150 2928 2152 2980
rect 2152 2928 2204 2980
rect 2204 2928 2206 2980
rect 2150 2926 2206 2928
rect 2151 2439 2207 2441
rect 2151 2387 2153 2439
rect 2153 2387 2205 2439
rect 2205 2387 2207 2439
rect 2151 2385 2207 2387
rect 1208 1294 1264 1296
rect 1208 1242 1210 1294
rect 1210 1242 1262 1294
rect 1262 1242 1264 1294
rect 1208 1240 1264 1242
rect 1425 1294 1481 1296
rect 1425 1242 1427 1294
rect 1427 1242 1479 1294
rect 1479 1242 1481 1294
rect 1425 1240 1481 1242
rect 1644 1294 1700 1296
rect 1644 1242 1646 1294
rect 1646 1242 1698 1294
rect 1698 1242 1700 1294
rect 1644 1240 1700 1242
rect 1857 1290 1913 1292
rect 1857 1238 1859 1290
rect 1859 1238 1911 1290
rect 1911 1238 1913 1290
rect 1857 1236 1913 1238
rect 278 452 334 454
rect 278 400 280 452
rect 280 400 332 452
rect 332 400 334 452
rect 278 398 334 400
rect 493 459 549 461
rect 493 407 495 459
rect 495 407 547 459
rect 547 407 549 459
rect 493 405 549 407
rect 711 456 767 458
rect 711 404 713 456
rect 713 404 765 456
rect 765 404 767 456
rect 711 402 767 404
rect 927 457 983 459
rect 927 405 929 457
rect 929 405 981 457
rect 981 405 983 457
rect 927 403 983 405
rect 1419 612 1475 614
rect 1190 600 1246 602
rect 1190 548 1192 600
rect 1192 548 1244 600
rect 1244 548 1246 600
rect 1419 560 1421 612
rect 1421 560 1473 612
rect 1473 560 1475 612
rect 1419 558 1475 560
rect 1638 602 1694 604
rect 1638 550 1640 602
rect 1640 550 1692 602
rect 1692 550 1694 602
rect 1190 546 1246 548
rect 1638 548 1694 550
rect 1830 606 1886 608
rect 1830 554 1832 606
rect 1832 554 1884 606
rect 1884 554 1886 606
rect 1830 552 1886 554
rect 2068 1290 2124 1292
rect 2068 1238 2070 1290
rect 2070 1238 2122 1290
rect 2122 1238 2124 1290
rect 2068 1236 2124 1238
rect 419 -76 475 -74
rect 419 -128 421 -76
rect 421 -128 473 -76
rect 473 -128 475 -76
rect 419 -130 475 -128
rect 618 -79 674 -77
rect 618 -131 620 -79
rect 620 -131 672 -79
rect 672 -131 674 -79
rect 618 -133 674 -131
rect 829 -79 885 -77
rect 829 -131 831 -79
rect 831 -131 883 -79
rect 883 -131 885 -79
rect 829 -133 885 -131
rect 1035 -79 1091 -77
rect 1035 -131 1037 -79
rect 1037 -131 1089 -79
rect 1089 -131 1091 -79
rect 1035 -133 1091 -131
rect 1263 -81 1319 -79
rect 1263 -133 1265 -81
rect 1265 -133 1317 -81
rect 1317 -133 1319 -81
rect 1263 -135 1319 -133
rect 1507 -81 1563 -79
rect 1507 -133 1509 -81
rect 1509 -133 1561 -81
rect 1561 -133 1563 -81
rect 1507 -135 1563 -133
rect 1737 -79 1793 -77
rect 1737 -131 1739 -79
rect 1739 -131 1791 -79
rect 1791 -131 1793 -79
rect 1737 -133 1793 -131
rect 1943 -79 1999 -77
rect 1943 -131 1945 -79
rect 1945 -131 1997 -79
rect 1997 -131 1999 -79
rect 1943 -133 1999 -131
rect 2427 2973 2483 2975
rect 2427 2921 2429 2973
rect 2429 2921 2481 2973
rect 2481 2921 2483 2973
rect 2427 2919 2483 2921
rect 2324 604 2380 606
rect 2324 552 2326 604
rect 2326 552 2378 604
rect 2378 552 2380 604
rect 2324 550 2380 552
rect 2650 2976 2706 2978
rect 2650 2924 2652 2976
rect 2652 2924 2704 2976
rect 2704 2924 2706 2976
rect 2650 2922 2706 2924
rect 2882 2975 2938 2977
rect 2882 2923 2884 2975
rect 2884 2923 2936 2975
rect 2936 2923 2938 2975
rect 2882 2921 2938 2923
rect 2701 1834 2757 1836
rect 2701 1782 2703 1834
rect 2703 1782 2755 1834
rect 2755 1782 2757 1834
rect 2701 1780 2757 1782
rect 3026 1836 3082 1838
rect 3026 1784 3028 1836
rect 3028 1784 3080 1836
rect 3080 1784 3082 1836
rect 3026 1782 3082 1784
rect 3294 1836 3350 1838
rect 3294 1784 3296 1836
rect 3296 1784 3348 1836
rect 3348 1784 3350 1836
rect 3294 1782 3350 1784
rect 2652 1146 2708 1148
rect 2652 1094 2654 1146
rect 2654 1094 2706 1146
rect 2706 1094 2708 1146
rect 2652 1092 2708 1094
rect 2867 1143 2923 1145
rect 2867 1091 2869 1143
rect 2869 1091 2921 1143
rect 2921 1091 2923 1143
rect 2867 1089 2923 1091
rect 3065 1140 3121 1142
rect 3065 1088 3067 1140
rect 3067 1088 3119 1140
rect 3119 1088 3121 1140
rect 3065 1086 3121 1088
rect 3260 1150 3316 1152
rect 3260 1098 3262 1150
rect 3262 1098 3314 1150
rect 3314 1098 3316 1150
rect 3260 1096 3316 1098
rect 3560 1836 3616 1838
rect 3560 1784 3562 1836
rect 3562 1784 3614 1836
rect 3614 1784 3616 1836
rect 3560 1782 3616 1784
rect 3800 1834 3856 1836
rect 3800 1782 3802 1834
rect 3802 1782 3854 1834
rect 3854 1782 3856 1834
rect 3800 1780 3856 1782
rect 4226 2437 4282 2439
rect 4226 2385 4228 2437
rect 4228 2385 4280 2437
rect 4280 2385 4282 2437
rect 4226 2383 4282 2385
rect 4518 2972 4574 2974
rect 4518 2920 4520 2972
rect 4520 2920 4572 2972
rect 4572 2920 4574 2972
rect 4518 2918 4574 2920
rect 4475 2440 4531 2442
rect 4475 2388 4477 2440
rect 4477 2388 4529 2440
rect 4529 2388 4531 2440
rect 4475 2386 4531 2388
rect 4192 1290 4248 1292
rect 4192 1238 4194 1290
rect 4194 1238 4246 1290
rect 4246 1238 4248 1290
rect 4192 1236 4248 1238
rect 3540 1148 3596 1150
rect 3540 1096 3542 1148
rect 3542 1096 3594 1148
rect 3594 1096 3596 1148
rect 3540 1094 3596 1096
rect 3759 1146 3815 1148
rect 3759 1094 3761 1146
rect 3761 1094 3813 1146
rect 3813 1094 3815 1146
rect 3759 1092 3815 1094
rect 2648 453 2704 455
rect 2648 401 2650 453
rect 2650 401 2702 453
rect 2702 401 2704 453
rect 2648 399 2704 401
rect 2838 453 2894 455
rect 2838 401 2840 453
rect 2840 401 2892 453
rect 2892 401 2894 453
rect 2838 399 2894 401
rect 3048 456 3104 458
rect 3048 404 3050 456
rect 3050 404 3102 456
rect 3102 404 3104 456
rect 3048 402 3104 404
rect 3265 453 3321 455
rect 3265 401 3267 453
rect 3267 401 3319 453
rect 3319 401 3321 453
rect 3265 399 3321 401
rect 4116 603 4172 605
rect 4116 551 4118 603
rect 4118 551 4170 603
rect 4170 551 4172 603
rect 4116 549 4172 551
rect 3560 456 3616 458
rect 3560 404 3562 456
rect 3562 404 3614 456
rect 3614 404 3616 456
rect 3560 402 3616 404
rect 3784 461 3840 463
rect 3784 409 3786 461
rect 3786 409 3838 461
rect 3838 409 3840 461
rect 3784 407 3840 409
rect 2161 -74 2217 -72
rect 2161 -126 2163 -74
rect 2163 -126 2215 -74
rect 2215 -126 2217 -74
rect 2161 -128 2217 -126
rect 2364 -80 2420 -78
rect 2364 -132 2366 -80
rect 2366 -132 2418 -80
rect 2418 -132 2420 -80
rect 2364 -134 2420 -132
rect 2572 -77 2628 -75
rect 2572 -129 2574 -77
rect 2574 -129 2626 -77
rect 2626 -129 2628 -77
rect 2572 -131 2628 -129
rect 4470 1289 4526 1291
rect 4470 1237 4472 1289
rect 4472 1237 4524 1289
rect 4524 1237 4526 1289
rect 4470 1235 4526 1237
rect 2835 -81 2891 -79
rect 2835 -133 2837 -81
rect 2837 -133 2889 -81
rect 2889 -133 2891 -81
rect 2835 -135 2891 -133
rect 3043 -80 3099 -78
rect 3043 -132 3045 -80
rect 3045 -132 3097 -80
rect 3097 -132 3099 -80
rect 3043 -134 3099 -132
rect 3253 -83 3309 -81
rect 3253 -135 3255 -83
rect 3255 -135 3307 -83
rect 3307 -135 3309 -83
rect 3253 -137 3309 -135
rect 3453 -77 3509 -75
rect 3453 -129 3455 -77
rect 3455 -129 3507 -77
rect 3507 -129 3509 -77
rect 3453 -131 3509 -129
rect 3656 -80 3712 -78
rect 3656 -132 3658 -80
rect 3658 -132 3710 -80
rect 3710 -132 3712 -80
rect 3656 -134 3712 -132
rect 3866 -80 3922 -78
rect 3866 -132 3868 -80
rect 3868 -132 3920 -80
rect 3920 -132 3922 -80
rect 3866 -134 3922 -132
rect 4067 -79 4123 -77
rect 4067 -131 4069 -79
rect 4069 -131 4121 -79
rect 4121 -131 4123 -79
rect 4067 -133 4123 -131
rect 4283 -78 4339 -76
rect 4283 -130 4285 -78
rect 4285 -130 4337 -78
rect 4337 -130 4339 -78
rect 4283 -132 4339 -130
rect 4509 601 4565 603
rect 4509 549 4511 601
rect 4511 549 4563 601
rect 4563 549 4565 601
rect 4509 547 4565 549
rect 4826 2973 4882 2975
rect 4826 2921 4828 2973
rect 4828 2921 4880 2973
rect 4880 2921 4882 2973
rect 4826 2919 4882 2921
rect 4819 2426 4875 2428
rect 4819 2374 4821 2426
rect 4821 2374 4873 2426
rect 4873 2374 4875 2426
rect 4819 2372 4875 2374
rect 4706 609 4762 611
rect 4706 557 4708 609
rect 4708 557 4760 609
rect 4760 557 4762 609
rect 4706 555 4762 557
rect 5026 2974 5082 2976
rect 5026 2922 5028 2974
rect 5028 2922 5080 2974
rect 5080 2922 5082 2974
rect 5026 2920 5082 2922
rect 5245 2973 5301 2975
rect 5245 2921 5247 2973
rect 5247 2921 5299 2973
rect 5299 2921 5301 2973
rect 5245 2919 5301 2921
rect 5491 2972 5547 2974
rect 5491 2920 5493 2972
rect 5493 2920 5545 2972
rect 5545 2920 5547 2972
rect 5491 2918 5547 2920
rect 5699 2974 5755 2976
rect 5699 2922 5701 2974
rect 5701 2922 5753 2974
rect 5753 2922 5755 2974
rect 5699 2920 5755 2922
rect 5901 2975 5957 2977
rect 5901 2923 5903 2975
rect 5903 2923 5955 2975
rect 5955 2923 5957 2975
rect 5901 2921 5957 2923
rect 6094 2974 6150 2976
rect 6094 2922 6096 2974
rect 6096 2922 6148 2974
rect 6148 2922 6150 2974
rect 6094 2920 6150 2922
rect 5073 2432 5129 2434
rect 5073 2380 5075 2432
rect 5075 2380 5127 2432
rect 5127 2380 5129 2432
rect 5073 2378 5129 2380
rect 5302 2432 5358 2434
rect 5302 2380 5304 2432
rect 5304 2380 5356 2432
rect 5356 2380 5358 2432
rect 5302 2378 5358 2380
rect 5594 1837 5650 1839
rect 5594 1785 5596 1837
rect 5596 1785 5648 1837
rect 5648 1785 5650 1837
rect 5594 1783 5650 1785
rect 5042 1294 5098 1296
rect 5042 1242 5044 1294
rect 5044 1242 5096 1294
rect 5096 1242 5098 1294
rect 5042 1240 5098 1242
rect 5281 1294 5337 1296
rect 5281 1242 5283 1294
rect 5283 1242 5335 1294
rect 5335 1242 5337 1294
rect 5281 1240 5337 1242
rect 5580 1143 5636 1145
rect 5580 1091 5582 1143
rect 5582 1091 5634 1143
rect 5634 1091 5636 1143
rect 5580 1089 5636 1091
rect 5960 1840 6016 1842
rect 5960 1788 5962 1840
rect 5962 1788 6014 1840
rect 6014 1788 6016 1840
rect 5960 1786 6016 1788
rect 6204 1840 6260 1842
rect 6204 1788 6206 1840
rect 6206 1788 6258 1840
rect 6258 1788 6260 1840
rect 6204 1786 6260 1788
rect 6466 2973 6522 2975
rect 6466 2921 6468 2973
rect 6468 2921 6520 2973
rect 6520 2921 6522 2973
rect 6466 2919 6522 2921
rect 6655 2971 6711 2973
rect 6655 2919 6657 2971
rect 6657 2919 6709 2971
rect 6709 2919 6711 2971
rect 6655 2917 6711 2919
rect 6627 1831 6683 1833
rect 6627 1779 6629 1831
rect 6629 1779 6681 1831
rect 6681 1779 6683 1831
rect 6627 1777 6683 1779
rect 6945 2971 7001 2973
rect 6945 2919 6947 2971
rect 6947 2919 6999 2971
rect 6999 2919 7001 2971
rect 6945 2917 7001 2919
rect 7020 2437 7076 2439
rect 7020 2385 7022 2437
rect 7022 2385 7074 2437
rect 7074 2385 7076 2437
rect 7020 2383 7076 2385
rect 5931 1140 5987 1142
rect 5931 1088 5933 1140
rect 5933 1088 5985 1140
rect 5985 1088 5987 1140
rect 5931 1086 5987 1088
rect 6120 1138 6176 1140
rect 6120 1086 6122 1138
rect 6122 1086 6174 1138
rect 6174 1086 6176 1138
rect 6120 1084 6176 1086
rect 6325 1145 6381 1147
rect 6325 1093 6327 1145
rect 6327 1093 6379 1145
rect 6379 1093 6381 1145
rect 6325 1091 6381 1093
rect 6516 1147 6572 1149
rect 6516 1095 6518 1147
rect 6518 1095 6570 1147
rect 6570 1095 6572 1147
rect 6516 1093 6572 1095
rect 5036 611 5092 613
rect 5036 559 5038 611
rect 5038 559 5090 611
rect 5090 559 5092 611
rect 5036 557 5092 559
rect 5232 611 5288 613
rect 5232 559 5234 611
rect 5234 559 5286 611
rect 5286 559 5288 611
rect 5232 557 5288 559
rect 5662 454 5718 456
rect 5662 402 5664 454
rect 5664 402 5716 454
rect 5716 402 5718 454
rect 5662 400 5718 402
rect 5962 452 6018 454
rect 5962 400 5964 452
rect 5964 400 6016 452
rect 6016 400 6018 452
rect 5962 398 6018 400
rect 6214 456 6270 458
rect 6214 404 6216 456
rect 6216 404 6268 456
rect 6268 404 6270 456
rect 6214 402 6270 404
rect 6431 461 6487 463
rect 6431 409 6433 461
rect 6433 409 6485 461
rect 6485 409 6487 461
rect 6431 407 6487 409
rect 6632 458 6688 460
rect 6632 406 6634 458
rect 6634 406 6686 458
rect 6686 406 6688 458
rect 6632 404 6688 406
rect 4564 -80 4620 -78
rect 4564 -132 4566 -80
rect 4566 -132 4618 -80
rect 4618 -132 4620 -80
rect 4564 -134 4620 -132
rect 4784 -85 4840 -83
rect 4784 -137 4786 -85
rect 4786 -137 4838 -85
rect 4838 -137 4840 -85
rect 4784 -139 4840 -137
rect 4989 -84 5045 -82
rect 4989 -136 4991 -84
rect 4991 -136 5043 -84
rect 5043 -136 5045 -84
rect 4989 -138 5045 -136
rect 5210 -78 5266 -76
rect 5210 -130 5212 -78
rect 5212 -130 5264 -78
rect 5264 -130 5266 -78
rect 5210 -132 5266 -130
rect 5415 -85 5471 -83
rect 5415 -137 5417 -85
rect 5417 -137 5469 -85
rect 5469 -137 5471 -85
rect 5415 -139 5471 -137
rect 5624 -84 5680 -82
rect 5624 -136 5626 -84
rect 5626 -136 5678 -84
rect 5678 -136 5680 -84
rect 5624 -138 5680 -136
rect 5841 -84 5897 -82
rect 5841 -136 5843 -84
rect 5843 -136 5895 -84
rect 5895 -136 5897 -84
rect 5841 -138 5897 -136
rect 6055 -79 6111 -77
rect 6055 -131 6057 -79
rect 6057 -131 6109 -79
rect 6109 -131 6111 -79
rect 6055 -133 6111 -131
rect 6250 -81 6306 -79
rect 6250 -133 6252 -81
rect 6252 -133 6304 -81
rect 6304 -133 6306 -81
rect 6250 -135 6306 -133
rect 6445 -84 6501 -82
rect 6445 -136 6447 -84
rect 6447 -136 6499 -84
rect 6499 -136 6501 -84
rect 6445 -138 6501 -136
rect 6647 -81 6703 -79
rect 6647 -133 6649 -81
rect 6649 -133 6701 -81
rect 6701 -133 6703 -81
rect 6647 -135 6703 -133
rect 7218 2973 7274 2975
rect 7218 2921 7220 2973
rect 7220 2921 7272 2973
rect 7272 2921 7274 2973
rect 7218 2919 7274 2921
rect 7224 2439 7280 2441
rect 7224 2387 7226 2439
rect 7226 2387 7278 2439
rect 7278 2387 7280 2439
rect 7224 2385 7280 2387
rect 7139 604 7195 606
rect 7139 552 7141 604
rect 7141 552 7193 604
rect 7193 552 7195 604
rect 7139 550 7195 552
rect 7547 2437 7603 2439
rect 7547 2385 7549 2437
rect 7549 2385 7601 2437
rect 7601 2385 7603 2437
rect 7547 2383 7603 2385
rect 7439 1292 7495 1294
rect 7439 1240 7441 1292
rect 7441 1240 7493 1292
rect 7493 1240 7495 1292
rect 7439 1238 7495 1240
rect 7666 1297 7722 1299
rect 7666 1245 7668 1297
rect 7668 1245 7720 1297
rect 7720 1245 7722 1297
rect 7666 1243 7722 1245
rect 7856 1299 7912 1301
rect 7856 1247 7858 1299
rect 7858 1247 7910 1299
rect 7910 1247 7912 1299
rect 7856 1245 7912 1247
rect 8072 1290 8128 1292
rect 8072 1238 8074 1290
rect 8074 1238 8126 1290
rect 8126 1238 8128 1290
rect 8072 1236 8128 1238
rect 8570 1833 8626 1835
rect 8570 1781 8572 1833
rect 8572 1781 8624 1833
rect 8624 1781 8626 1833
rect 8570 1779 8626 1781
rect 8822 1830 8878 1832
rect 8822 1778 8824 1830
rect 8824 1778 8876 1830
rect 8876 1778 8878 1830
rect 8822 1776 8878 1778
rect 9028 1838 9084 1840
rect 9028 1786 9030 1838
rect 9030 1786 9082 1838
rect 9082 1786 9084 1838
rect 9028 1784 9084 1786
rect 9311 1832 9367 1834
rect 9311 1780 9313 1832
rect 9313 1780 9365 1832
rect 9365 1780 9367 1832
rect 9311 1778 9367 1780
rect 8561 1149 8617 1151
rect 8561 1097 8563 1149
rect 8563 1097 8615 1149
rect 8615 1097 8617 1149
rect 8561 1095 8617 1097
rect 8751 1151 8807 1153
rect 8751 1099 8753 1151
rect 8753 1099 8805 1151
rect 8805 1099 8807 1151
rect 8751 1097 8807 1099
rect 8945 1149 9001 1151
rect 8945 1097 8947 1149
rect 8947 1097 8999 1149
rect 8999 1097 9001 1149
rect 8945 1095 9001 1097
rect 7440 608 7496 610
rect 7440 556 7442 608
rect 7442 556 7494 608
rect 7494 556 7496 608
rect 7440 554 7496 556
rect 7646 609 7702 611
rect 7646 557 7648 609
rect 7648 557 7700 609
rect 7700 557 7702 609
rect 7646 555 7702 557
rect 7856 605 7912 607
rect 7856 553 7858 605
rect 7858 553 7910 605
rect 7910 553 7912 605
rect 7856 551 7912 553
rect 8067 611 8123 613
rect 8067 559 8069 611
rect 8069 559 8121 611
rect 8121 559 8123 611
rect 8067 557 8123 559
rect 8517 449 8573 451
rect 8517 397 8519 449
rect 8519 397 8571 449
rect 8571 397 8573 449
rect 8517 395 8573 397
rect 8709 449 8765 451
rect 8709 397 8711 449
rect 8711 397 8763 449
rect 8763 397 8765 449
rect 8709 395 8765 397
rect 8909 449 8965 451
rect 8909 397 8911 449
rect 8911 397 8963 449
rect 8963 397 8965 449
rect 8909 395 8965 397
rect 6931 -80 6987 -78
rect 6931 -132 6933 -80
rect 6933 -132 6985 -80
rect 6985 -132 6987 -80
rect 6931 -134 6987 -132
rect 7130 -79 7186 -77
rect 7130 -131 7132 -79
rect 7132 -131 7184 -79
rect 7184 -131 7186 -79
rect 7130 -133 7186 -131
rect 7333 -77 7389 -75
rect 7333 -129 7335 -77
rect 7335 -129 7387 -77
rect 7387 -129 7389 -77
rect 7333 -131 7389 -129
rect 9256 1145 9312 1147
rect 9256 1093 9258 1145
rect 9258 1093 9310 1145
rect 9310 1093 9312 1145
rect 9256 1091 9312 1093
rect 7598 -80 7654 -78
rect 7598 -132 7600 -80
rect 7600 -132 7652 -80
rect 7652 -132 7654 -80
rect 7598 -134 7654 -132
rect 7796 -81 7852 -79
rect 7796 -133 7798 -81
rect 7798 -133 7850 -81
rect 7850 -133 7852 -81
rect 7796 -135 7852 -133
rect 7985 -79 8041 -77
rect 7985 -131 7987 -79
rect 7987 -131 8039 -79
rect 8039 -131 8041 -79
rect 7985 -133 8041 -131
rect 8197 -79 8253 -77
rect 8197 -131 8199 -79
rect 8199 -131 8251 -79
rect 8251 -131 8253 -79
rect 8197 -133 8253 -131
rect 8414 -79 8470 -77
rect 8414 -131 8416 -79
rect 8416 -131 8468 -79
rect 8468 -131 8470 -79
rect 8414 -133 8470 -131
rect 8619 -83 8675 -81
rect 8619 -135 8621 -83
rect 8621 -135 8673 -83
rect 8673 -135 8675 -83
rect 8619 -137 8675 -135
rect 8824 -83 8880 -81
rect 8824 -135 8826 -83
rect 8826 -135 8878 -83
rect 8878 -135 8880 -83
rect 8824 -137 8880 -135
rect 9032 -78 9088 -76
rect 9032 -130 9034 -78
rect 9034 -130 9086 -78
rect 9086 -130 9088 -78
rect 9032 -132 9088 -130
rect 9609 1833 9665 1835
rect 9609 1781 9611 1833
rect 9611 1781 9663 1833
rect 9663 1781 9665 1833
rect 9609 1779 9665 1781
rect 9527 457 9583 459
rect 9527 405 9529 457
rect 9529 405 9581 457
rect 9581 405 9583 457
rect 9527 403 9583 405
rect 10053 1293 10109 1295
rect 10053 1241 10055 1293
rect 10055 1241 10107 1293
rect 10107 1241 10109 1293
rect 10053 1239 10109 1241
rect 10282 1296 10338 1298
rect 10282 1244 10284 1296
rect 10284 1244 10336 1296
rect 10336 1244 10338 1296
rect 10282 1242 10338 1244
rect 10508 1301 10564 1303
rect 10508 1249 10510 1301
rect 10510 1249 10562 1301
rect 10562 1249 10564 1301
rect 10508 1247 10564 1249
rect 11441 1834 11497 1836
rect 11441 1782 11443 1834
rect 11443 1782 11495 1834
rect 11495 1782 11497 1834
rect 11441 1780 11497 1782
rect 11651 1836 11707 1838
rect 11651 1784 11653 1836
rect 11653 1784 11705 1836
rect 11705 1784 11707 1836
rect 11651 1782 11707 1784
rect 10736 1293 10792 1295
rect 10736 1241 10738 1293
rect 10738 1241 10790 1293
rect 10790 1241 10792 1293
rect 10736 1239 10792 1241
rect 10972 1299 11028 1301
rect 10972 1247 10974 1299
rect 10974 1247 11026 1299
rect 11026 1247 11028 1299
rect 10972 1245 11028 1247
rect 11164 1290 11220 1292
rect 11164 1238 11166 1290
rect 11166 1238 11218 1290
rect 11218 1238 11220 1290
rect 11164 1236 11220 1238
rect 11439 1144 11495 1146
rect 11439 1092 11441 1144
rect 11441 1092 11493 1144
rect 11493 1092 11495 1144
rect 11439 1090 11495 1092
rect 9947 600 10003 602
rect 9947 548 9949 600
rect 9949 548 10001 600
rect 10001 548 10003 600
rect 9947 546 10003 548
rect 10204 607 10260 609
rect 10204 555 10206 607
rect 10206 555 10258 607
rect 10258 555 10260 607
rect 10204 553 10260 555
rect 10454 603 10510 605
rect 10454 551 10456 603
rect 10456 551 10508 603
rect 10508 551 10510 603
rect 10454 549 10510 551
rect 10725 608 10781 610
rect 10725 556 10727 608
rect 10727 556 10779 608
rect 10779 556 10781 608
rect 10725 554 10781 556
rect 10966 611 11022 613
rect 10966 559 10968 611
rect 10968 559 11020 611
rect 11020 559 11022 611
rect 10966 557 11022 559
rect 11191 607 11247 609
rect 11191 555 11193 607
rect 11193 555 11245 607
rect 11245 555 11247 607
rect 11191 553 11247 555
rect 11428 453 11484 455
rect 11428 401 11430 453
rect 11430 401 11482 453
rect 11482 401 11484 453
rect 11428 399 11484 401
rect 9315 -79 9371 -77
rect 9315 -131 9317 -79
rect 9317 -131 9369 -79
rect 9369 -131 9371 -79
rect 9315 -133 9371 -131
rect 9508 -81 9564 -79
rect 9508 -133 9510 -81
rect 9510 -133 9562 -81
rect 9562 -133 9564 -81
rect 9508 -135 9564 -133
rect 9734 -83 9790 -81
rect 9734 -135 9736 -83
rect 9736 -135 9788 -83
rect 9788 -135 9790 -83
rect 9734 -137 9790 -135
rect 11643 1144 11699 1146
rect 11643 1092 11645 1144
rect 11645 1092 11697 1144
rect 11697 1092 11699 1144
rect 11643 1090 11699 1092
rect 9999 -83 10055 -81
rect 9999 -135 10001 -83
rect 10001 -135 10053 -83
rect 10053 -135 10055 -83
rect 9999 -137 10055 -135
rect 10193 -79 10249 -77
rect 10193 -131 10195 -79
rect 10195 -131 10247 -79
rect 10247 -131 10249 -79
rect 10193 -133 10249 -131
rect 10391 -88 10447 -86
rect 10391 -140 10393 -88
rect 10393 -140 10445 -88
rect 10445 -140 10447 -88
rect 10391 -142 10447 -140
rect 10595 -80 10651 -78
rect 10595 -132 10597 -80
rect 10597 -132 10649 -80
rect 10649 -132 10651 -80
rect 10595 -134 10651 -132
rect 10815 -77 10871 -75
rect 10815 -129 10817 -77
rect 10817 -129 10869 -77
rect 10869 -129 10871 -77
rect 10815 -131 10871 -129
rect 11030 -81 11086 -79
rect 11030 -133 11032 -81
rect 11032 -133 11084 -81
rect 11084 -133 11086 -81
rect 11030 -135 11086 -133
rect 11258 -78 11314 -76
rect 11258 -130 11260 -78
rect 11260 -130 11312 -78
rect 11312 -130 11314 -78
rect 11258 -132 11314 -130
rect 11462 -81 11518 -79
rect 11462 -133 11464 -81
rect 11464 -133 11516 -81
rect 11516 -133 11518 -81
rect 11462 -135 11518 -133
rect 11684 453 11740 455
rect 11684 401 11686 453
rect 11686 401 11738 453
rect 11738 401 11740 453
rect 11684 399 11740 401
rect 12002 1834 12058 1836
rect 12002 1782 12004 1834
rect 12004 1782 12056 1834
rect 12056 1782 12058 1834
rect 12002 1780 12058 1782
rect 11919 453 11975 455
rect 11919 401 11921 453
rect 11921 401 11973 453
rect 11973 401 11975 453
rect 11919 399 11975 401
rect 12282 1834 12338 1836
rect 12282 1782 12284 1834
rect 12284 1782 12336 1834
rect 12336 1782 12338 1834
rect 12282 1780 12338 1782
rect 12599 1833 12655 1835
rect 12599 1781 12601 1833
rect 12601 1781 12653 1833
rect 12653 1781 12655 1833
rect 12599 1779 12655 1781
rect 12208 1140 12264 1142
rect 12208 1088 12210 1140
rect 12210 1088 12262 1140
rect 12262 1088 12264 1140
rect 12208 1086 12264 1088
rect 12899 1290 12955 1292
rect 12899 1238 12901 1290
rect 12901 1238 12953 1290
rect 12953 1238 12955 1290
rect 12899 1236 12955 1238
rect 12447 1142 12503 1144
rect 12447 1090 12449 1142
rect 12449 1090 12501 1142
rect 12501 1090 12503 1142
rect 12447 1088 12503 1090
rect 12651 1142 12707 1144
rect 12651 1090 12653 1142
rect 12653 1090 12705 1142
rect 12705 1090 12707 1142
rect 12651 1088 12707 1090
rect 13103 1295 13159 1297
rect 13103 1243 13105 1295
rect 13105 1243 13157 1295
rect 13157 1243 13159 1295
rect 13103 1241 13159 1243
rect 13294 1290 13350 1292
rect 13294 1238 13296 1290
rect 13296 1238 13348 1290
rect 13348 1238 13350 1290
rect 13294 1236 13350 1238
rect 13496 1289 13552 1291
rect 13496 1237 13498 1289
rect 13498 1237 13550 1289
rect 13550 1237 13552 1289
rect 13496 1235 13552 1237
rect 13786 1290 13842 1292
rect 13786 1238 13788 1290
rect 13788 1238 13840 1290
rect 13840 1238 13842 1290
rect 13786 1236 13842 1238
rect 12898 605 12954 607
rect 12898 553 12900 605
rect 12900 553 12952 605
rect 12952 553 12954 605
rect 12898 551 12954 553
rect 12208 455 12264 457
rect 12208 403 12210 455
rect 12210 403 12262 455
rect 12262 403 12264 455
rect 12208 401 12264 403
rect 12398 453 12454 455
rect 12398 401 12400 453
rect 12400 401 12452 453
rect 12452 401 12454 453
rect 12398 399 12454 401
rect 12602 455 12658 457
rect 12602 403 12604 455
rect 12604 403 12656 455
rect 12656 403 12658 455
rect 12602 401 12658 403
rect 13099 606 13155 608
rect 13099 554 13101 606
rect 13101 554 13153 606
rect 13153 554 13155 606
rect 13099 552 13155 554
rect 13317 602 13373 604
rect 13317 550 13319 602
rect 13319 550 13371 602
rect 13371 550 13373 602
rect 13317 548 13373 550
rect 13524 606 13580 608
rect 13524 554 13526 606
rect 13526 554 13578 606
rect 13578 554 13580 606
rect 13524 552 13580 554
rect 13729 605 13785 607
rect 13729 553 13731 605
rect 13731 553 13783 605
rect 13783 553 13785 605
rect 13729 551 13785 553
rect 11700 -79 11756 -77
rect 11700 -131 11702 -79
rect 11702 -131 11754 -79
rect 11754 -131 11756 -79
rect 11700 -133 11756 -131
rect 11893 -78 11949 -76
rect 11893 -130 11895 -78
rect 11895 -130 11947 -78
rect 11947 -130 11949 -78
rect 11893 -132 11949 -130
rect 12090 -83 12146 -81
rect 12090 -135 12092 -83
rect 12092 -135 12144 -83
rect 12144 -135 12146 -83
rect 12090 -137 12146 -135
rect 14071 1289 14127 1291
rect 14071 1237 14073 1289
rect 14073 1237 14125 1289
rect 14125 1237 14127 1289
rect 14071 1235 14127 1237
rect 12346 -80 12402 -78
rect 12346 -132 12348 -80
rect 12348 -132 12400 -80
rect 12400 -132 12402 -80
rect 12346 -134 12402 -132
rect 12585 -84 12641 -82
rect 12585 -136 12587 -84
rect 12587 -136 12639 -84
rect 12639 -136 12641 -84
rect 12585 -138 12641 -136
rect 12818 -88 12874 -86
rect 12818 -140 12820 -88
rect 12820 -140 12872 -88
rect 12872 -140 12874 -88
rect 12818 -142 12874 -140
rect 13039 -83 13095 -81
rect 13039 -135 13041 -83
rect 13041 -135 13093 -83
rect 13093 -135 13095 -83
rect 13039 -137 13095 -135
rect 13230 -83 13286 -81
rect 13230 -135 13232 -83
rect 13232 -135 13284 -83
rect 13284 -135 13286 -83
rect 13230 -137 13286 -135
rect 13458 -81 13514 -79
rect 13458 -133 13460 -81
rect 13460 -133 13512 -81
rect 13512 -133 13514 -81
rect 13458 -135 13514 -133
rect 13655 -86 13711 -84
rect 13655 -138 13657 -86
rect 13657 -138 13709 -86
rect 13709 -138 13711 -86
rect 13655 -140 13711 -138
rect 13867 -86 13923 -84
rect 13867 -138 13869 -86
rect 13869 -138 13921 -86
rect 13921 -138 13923 -86
rect 13867 -140 13923 -138
rect 14076 601 14132 603
rect 14076 549 14078 601
rect 14078 549 14130 601
rect 14130 549 14132 601
rect 14076 547 14132 549
rect 14389 1831 14445 1833
rect 14389 1779 14391 1831
rect 14391 1779 14443 1831
rect 14443 1779 14445 1831
rect 14389 1777 14445 1779
rect 14388 461 14444 463
rect 14388 409 14390 461
rect 14390 409 14442 461
rect 14442 409 14444 461
rect 14388 407 14444 409
rect 14684 1831 14740 1833
rect 14684 1779 14686 1831
rect 14686 1779 14738 1831
rect 14738 1779 14740 1831
rect 14684 1777 14740 1779
rect 14971 1831 15027 1833
rect 14971 1779 14973 1831
rect 14973 1779 15025 1831
rect 15025 1779 15027 1831
rect 14971 1777 15027 1779
rect 15261 1831 15317 1833
rect 15261 1779 15263 1831
rect 15263 1779 15315 1831
rect 15315 1779 15317 1831
rect 15261 1777 15317 1779
rect 14611 1150 14667 1152
rect 14611 1098 14613 1150
rect 14613 1098 14665 1150
rect 14665 1098 14667 1150
rect 14611 1096 14667 1098
rect 14844 1148 14900 1150
rect 14844 1096 14846 1148
rect 14846 1096 14898 1148
rect 14898 1096 14900 1148
rect 14844 1094 14900 1096
rect 15051 1146 15107 1148
rect 15051 1094 15053 1146
rect 15053 1094 15105 1146
rect 15105 1094 15107 1146
rect 15051 1092 15107 1094
rect 15260 1148 15316 1150
rect 15260 1096 15262 1148
rect 15262 1096 15314 1148
rect 15314 1096 15316 1148
rect 15260 1094 15316 1096
rect 15545 1834 15601 1836
rect 15545 1782 15547 1834
rect 15547 1782 15599 1834
rect 15599 1782 15601 1834
rect 15545 1780 15601 1782
rect 15826 1294 15882 1296
rect 15826 1242 15828 1294
rect 15828 1242 15880 1294
rect 15880 1242 15882 1294
rect 15826 1240 15882 1242
rect 16020 1298 16076 1300
rect 16020 1246 16022 1298
rect 16022 1246 16074 1298
rect 16074 1246 16076 1298
rect 16020 1244 16076 1246
rect 16209 1295 16265 1297
rect 16209 1243 16211 1295
rect 16211 1243 16263 1295
rect 16263 1243 16265 1295
rect 16209 1241 16265 1243
rect 15540 1150 15596 1152
rect 15540 1098 15542 1150
rect 15542 1098 15594 1150
rect 15594 1098 15596 1150
rect 15540 1096 15596 1098
rect 14630 457 14686 459
rect 14630 405 14632 457
rect 14632 405 14684 457
rect 14684 405 14686 457
rect 14630 403 14686 405
rect 14830 456 14886 458
rect 14830 404 14832 456
rect 14832 404 14884 456
rect 14884 404 14886 456
rect 14830 402 14886 404
rect 15020 464 15076 466
rect 15020 412 15022 464
rect 15022 412 15074 464
rect 15074 412 15076 464
rect 15020 410 15076 412
rect 15241 462 15297 464
rect 15241 410 15243 462
rect 15243 410 15295 462
rect 15295 410 15297 462
rect 15241 408 15297 410
rect 15828 605 15884 607
rect 15828 553 15830 605
rect 15830 553 15882 605
rect 15882 553 15884 605
rect 15828 551 15884 553
rect 16019 608 16075 610
rect 16019 556 16021 608
rect 16021 556 16073 608
rect 16073 556 16075 608
rect 16019 554 16075 556
rect 16214 610 16270 612
rect 16214 558 16216 610
rect 16216 558 16268 610
rect 16268 558 16270 610
rect 16214 556 16270 558
rect 15537 457 15593 459
rect 15537 405 15539 457
rect 15539 405 15591 457
rect 15591 405 15593 457
rect 15537 403 15593 405
rect 14094 -83 14150 -81
rect 14094 -135 14096 -83
rect 14096 -135 14148 -83
rect 14148 -135 14150 -83
rect 14094 -137 14150 -135
rect 14283 -82 14339 -80
rect 14283 -134 14285 -82
rect 14285 -134 14337 -82
rect 14337 -134 14339 -82
rect 14283 -136 14339 -134
rect 14509 -81 14565 -79
rect 14509 -133 14511 -81
rect 14511 -133 14563 -81
rect 14563 -133 14565 -81
rect 14509 -135 14565 -133
rect 16432 1297 16488 1299
rect 16432 1245 16434 1297
rect 16434 1245 16486 1297
rect 16486 1245 16488 1297
rect 16432 1243 16488 1245
rect 14763 -81 14819 -79
rect 14763 -133 14765 -81
rect 14765 -133 14817 -81
rect 14817 -133 14819 -81
rect 14763 -135 14819 -133
rect 15007 -84 15063 -82
rect 15007 -136 15009 -84
rect 15009 -136 15061 -84
rect 15061 -136 15063 -84
rect 15007 -138 15063 -136
rect 15237 -85 15293 -83
rect 15237 -137 15239 -85
rect 15239 -137 15291 -85
rect 15291 -137 15293 -85
rect 15237 -139 15293 -137
rect 15495 -82 15551 -80
rect 15495 -134 15497 -82
rect 15497 -134 15549 -82
rect 15549 -134 15551 -82
rect 15495 -136 15551 -134
rect 15705 -82 15761 -80
rect 15705 -134 15707 -82
rect 15707 -134 15759 -82
rect 15759 -134 15761 -82
rect 15705 -136 15761 -134
rect 15930 -82 15986 -80
rect 15930 -134 15932 -82
rect 15932 -134 15984 -82
rect 15984 -134 15986 -82
rect 15930 -136 15986 -134
rect 16149 -85 16205 -83
rect 16149 -137 16151 -85
rect 16151 -137 16203 -85
rect 16203 -137 16205 -85
rect 16149 -139 16205 -137
rect 16661 605 16717 607
rect 16661 553 16663 605
rect 16663 553 16715 605
rect 16715 553 16717 605
rect 16661 551 16717 553
rect 16495 -81 16551 -79
rect 16495 -133 16497 -81
rect 16497 -133 16549 -81
rect 16549 -133 16551 -81
rect 16495 -135 16551 -133
rect 16694 -84 16750 -82
rect 16694 -136 16696 -84
rect 16696 -136 16748 -84
rect 16748 -136 16750 -84
rect 16694 -138 16750 -136
<< metal3 >>
rect 686 3441 815 3452
rect 686 3377 717 3441
rect 781 3377 815 3441
rect 686 3366 815 3377
rect 16 2982 145 2993
rect 16 2918 47 2982
rect 111 2918 145 2982
rect 16 2907 145 2918
rect 218 2984 347 2995
rect 218 2920 249 2984
rect 313 2920 347 2984
rect 218 2909 347 2920
rect 429 2982 558 2993
rect 429 2918 460 2982
rect 524 2918 558 2982
rect 429 2907 558 2918
rect 619 2982 748 2993
rect 619 2918 650 2982
rect 714 2918 748 2982
rect 619 2907 748 2918
rect 827 2984 956 2995
rect 827 2920 858 2984
rect 922 2920 956 2984
rect 827 2909 956 2920
rect 1029 2984 1158 2995
rect 1029 2920 1060 2984
rect 1124 2920 1158 2984
rect 1029 2909 1158 2920
rect 1228 2986 1357 2997
rect 1228 2922 1259 2986
rect 1323 2922 1357 2986
rect 1228 2911 1357 2922
rect 1423 2983 1552 2994
rect 1423 2919 1454 2983
rect 1518 2919 1552 2983
rect 1423 2908 1552 2919
rect 1624 2985 1753 2996
rect 1624 2921 1655 2985
rect 1719 2921 1753 2985
rect 1624 2910 1753 2921
rect 1841 2983 1970 2994
rect 1841 2919 1872 2983
rect 1936 2919 1970 2983
rect 1841 2908 1970 2919
rect 2115 2986 2244 2997
rect 2115 2922 2146 2986
rect 2210 2922 2244 2986
rect 2115 2911 2244 2922
rect 2392 2979 2521 2990
rect 2392 2915 2423 2979
rect 2487 2915 2521 2979
rect 2392 2904 2521 2915
rect 2615 2982 2744 2993
rect 2615 2918 2646 2982
rect 2710 2918 2744 2982
rect 2615 2907 2744 2918
rect 2847 2981 2976 2992
rect 2847 2917 2878 2981
rect 2942 2917 2976 2981
rect 2847 2906 2976 2917
rect 4483 2978 4612 2989
rect 4483 2914 4514 2978
rect 4578 2914 4612 2978
rect 4483 2903 4612 2914
rect 4791 2979 4920 2990
rect 4791 2915 4822 2979
rect 4886 2915 4920 2979
rect 4791 2904 4920 2915
rect 4991 2980 5120 2991
rect 4991 2916 5022 2980
rect 5086 2916 5120 2980
rect 4991 2905 5120 2916
rect 5210 2979 5339 2990
rect 5210 2915 5241 2979
rect 5305 2915 5339 2979
rect 5210 2904 5339 2915
rect 5456 2978 5585 2989
rect 5456 2914 5487 2978
rect 5551 2914 5585 2978
rect 5456 2903 5585 2914
rect 5664 2980 5793 2991
rect 5664 2916 5695 2980
rect 5759 2916 5793 2980
rect 5664 2905 5793 2916
rect 5866 2981 5995 2992
rect 5866 2917 5897 2981
rect 5961 2917 5995 2981
rect 5866 2906 5995 2917
rect 6059 2980 6188 2991
rect 6059 2916 6090 2980
rect 6154 2916 6188 2980
rect 6059 2905 6188 2916
rect 6431 2979 6560 2990
rect 6431 2915 6462 2979
rect 6526 2915 6560 2979
rect 6431 2904 6560 2915
rect 6620 2977 6749 2988
rect 6620 2913 6651 2977
rect 6715 2913 6749 2977
rect 6620 2902 6749 2913
rect 6910 2977 7039 2988
rect 6910 2913 6941 2977
rect 7005 2913 7039 2977
rect 6910 2902 7039 2913
rect 7183 2979 7312 2990
rect 7183 2915 7214 2979
rect 7278 2915 7312 2979
rect 7183 2904 7312 2915
rect 1134 2443 1263 2454
rect 1134 2379 1165 2443
rect 1229 2379 1263 2443
rect 1134 2368 1263 2379
rect 1353 2447 1482 2458
rect 1353 2383 1384 2447
rect 1448 2383 1482 2447
rect 1353 2372 1482 2383
rect 1636 2447 1765 2458
rect 1636 2383 1667 2447
rect 1731 2383 1765 2447
rect 1636 2372 1765 2383
rect 1845 2447 1974 2458
rect 1845 2383 1876 2447
rect 1940 2383 1974 2447
rect 1845 2372 1974 2383
rect 2116 2445 2245 2456
rect 2116 2381 2147 2445
rect 2211 2381 2245 2445
rect 2116 2370 2245 2381
rect 4191 2443 4320 2454
rect 4191 2379 4222 2443
rect 4286 2379 4320 2443
rect 4191 2368 4320 2379
rect 4440 2446 4569 2457
rect 4440 2382 4471 2446
rect 4535 2382 4569 2446
rect 4440 2371 4569 2382
rect 4784 2432 4913 2443
rect 4784 2368 4815 2432
rect 4879 2368 4913 2432
rect 4784 2357 4913 2368
rect 5038 2438 5167 2449
rect 5038 2374 5069 2438
rect 5133 2374 5167 2438
rect 5038 2363 5167 2374
rect 5267 2438 5396 2449
rect 5267 2374 5298 2438
rect 5362 2374 5396 2438
rect 5267 2363 5396 2374
rect 6985 2443 7114 2454
rect 6985 2379 7016 2443
rect 7080 2379 7114 2443
rect 6985 2368 7114 2379
rect 7189 2445 7318 2456
rect 7189 2381 7220 2445
rect 7284 2381 7318 2445
rect 7189 2370 7318 2381
rect 7512 2443 7641 2454
rect 7512 2379 7543 2443
rect 7607 2379 7641 2443
rect 7512 2368 7641 2379
rect -18 1838 111 1849
rect -18 1774 13 1838
rect 77 1774 111 1838
rect -18 1763 111 1774
rect 222 1836 351 1847
rect 222 1772 253 1836
rect 317 1772 351 1836
rect 222 1761 351 1772
rect 544 1835 673 1846
rect 544 1771 575 1835
rect 639 1771 673 1835
rect 544 1760 673 1771
rect 762 1836 891 1847
rect 762 1772 793 1836
rect 857 1772 891 1836
rect 762 1761 891 1772
rect 2666 1840 2795 1851
rect 2666 1776 2697 1840
rect 2761 1776 2795 1840
rect 2666 1765 2795 1776
rect 2991 1842 3120 1853
rect 2991 1778 3022 1842
rect 3086 1778 3120 1842
rect 2991 1767 3120 1778
rect 3259 1842 3388 1853
rect 3259 1778 3290 1842
rect 3354 1778 3388 1842
rect 3259 1767 3388 1778
rect 3525 1842 3654 1853
rect 3525 1778 3556 1842
rect 3620 1778 3654 1842
rect 3525 1767 3654 1778
rect 3765 1840 3894 1851
rect 3765 1776 3796 1840
rect 3860 1776 3894 1840
rect 3765 1765 3894 1776
rect 5559 1843 5688 1854
rect 5559 1779 5590 1843
rect 5654 1779 5688 1843
rect 5559 1768 5688 1779
rect 5925 1846 6054 1857
rect 5925 1782 5956 1846
rect 6020 1782 6054 1846
rect 5925 1771 6054 1782
rect 6169 1846 6298 1857
rect 6169 1782 6200 1846
rect 6264 1782 6298 1846
rect 6169 1771 6298 1782
rect 6592 1837 6721 1848
rect 6592 1773 6623 1837
rect 6687 1773 6721 1837
rect 6592 1762 6721 1773
rect 8535 1839 8664 1850
rect 8535 1775 8566 1839
rect 8630 1775 8664 1839
rect 8535 1764 8664 1775
rect 8787 1836 8916 1847
rect 8787 1772 8818 1836
rect 8882 1772 8916 1836
rect 8787 1761 8916 1772
rect 8993 1844 9122 1855
rect 8993 1780 9024 1844
rect 9088 1780 9122 1844
rect 8993 1769 9122 1780
rect 9276 1838 9405 1849
rect 9276 1774 9307 1838
rect 9371 1774 9405 1838
rect 9276 1763 9405 1774
rect 9574 1839 9703 1850
rect 9574 1775 9605 1839
rect 9669 1775 9703 1839
rect 9574 1764 9703 1775
rect 11406 1840 11535 1851
rect 11406 1776 11437 1840
rect 11501 1776 11535 1840
rect 11406 1765 11535 1776
rect 11616 1842 11745 1853
rect 11616 1778 11647 1842
rect 11711 1778 11745 1842
rect 11616 1767 11745 1778
rect 11967 1840 12096 1851
rect 11967 1776 11998 1840
rect 12062 1776 12096 1840
rect 11967 1765 12096 1776
rect 12247 1840 12376 1851
rect 12247 1776 12278 1840
rect 12342 1776 12376 1840
rect 12247 1765 12376 1776
rect 12564 1839 12693 1850
rect 12564 1775 12595 1839
rect 12659 1775 12693 1839
rect 12564 1764 12693 1775
rect 14354 1837 14483 1848
rect 14354 1773 14385 1837
rect 14449 1773 14483 1837
rect 14354 1762 14483 1773
rect 14649 1837 14778 1848
rect 14649 1773 14680 1837
rect 14744 1773 14778 1837
rect 14649 1762 14778 1773
rect 14936 1837 15065 1848
rect 14936 1773 14967 1837
rect 15031 1773 15065 1837
rect 14936 1762 15065 1773
rect 15226 1837 15355 1848
rect 15226 1773 15257 1837
rect 15321 1773 15355 1837
rect 15226 1762 15355 1773
rect 15510 1840 15639 1851
rect 15510 1776 15541 1840
rect 15605 1776 15639 1840
rect 15510 1765 15639 1776
rect 1173 1300 1302 1311
rect 1173 1236 1204 1300
rect 1268 1236 1302 1300
rect 1173 1225 1302 1236
rect 1390 1300 1519 1311
rect 1390 1236 1421 1300
rect 1485 1236 1519 1300
rect 1390 1225 1519 1236
rect 1609 1300 1738 1311
rect 1609 1236 1640 1300
rect 1704 1236 1738 1300
rect 1609 1225 1738 1236
rect 1822 1296 1951 1307
rect 1822 1232 1853 1296
rect 1917 1232 1951 1296
rect 1822 1221 1951 1232
rect 2033 1296 2162 1307
rect 2033 1232 2064 1296
rect 2128 1232 2162 1296
rect 2033 1221 2162 1232
rect 4157 1296 4286 1307
rect 4157 1232 4188 1296
rect 4252 1232 4286 1296
rect 4157 1221 4286 1232
rect 4435 1295 4564 1306
rect 4435 1231 4466 1295
rect 4530 1231 4564 1295
rect 4435 1220 4564 1231
rect 5007 1300 5136 1311
rect 5007 1236 5038 1300
rect 5102 1236 5136 1300
rect 5007 1225 5136 1236
rect 5246 1300 5375 1311
rect 5246 1236 5277 1300
rect 5341 1236 5375 1300
rect 5246 1225 5375 1236
rect 7404 1298 7533 1309
rect 7404 1234 7435 1298
rect 7499 1234 7533 1298
rect 7404 1223 7533 1234
rect 7631 1303 7760 1314
rect 7631 1239 7662 1303
rect 7726 1239 7760 1303
rect 7631 1228 7760 1239
rect 7821 1305 7950 1316
rect 7821 1241 7852 1305
rect 7916 1241 7950 1305
rect 7821 1230 7950 1241
rect 8037 1296 8166 1307
rect 8037 1232 8068 1296
rect 8132 1232 8166 1296
rect 8037 1221 8166 1232
rect 10018 1299 10147 1310
rect 10018 1235 10049 1299
rect 10113 1235 10147 1299
rect 10018 1224 10147 1235
rect 10247 1302 10376 1313
rect 10247 1238 10278 1302
rect 10342 1238 10376 1302
rect 10247 1227 10376 1238
rect 10473 1307 10602 1318
rect 10473 1243 10504 1307
rect 10568 1243 10602 1307
rect 10473 1232 10602 1243
rect 10701 1299 10830 1310
rect 10701 1235 10732 1299
rect 10796 1235 10830 1299
rect 10701 1224 10830 1235
rect 10937 1305 11066 1316
rect 10937 1241 10968 1305
rect 11032 1241 11066 1305
rect 10937 1230 11066 1241
rect 11129 1296 11258 1307
rect 11129 1232 11160 1296
rect 11224 1232 11258 1296
rect 11129 1221 11258 1232
rect 12864 1296 12993 1307
rect 12864 1232 12895 1296
rect 12959 1232 12993 1296
rect 12864 1221 12993 1232
rect 13068 1301 13197 1312
rect 13068 1237 13099 1301
rect 13163 1237 13197 1301
rect 13068 1226 13197 1237
rect 13259 1296 13388 1307
rect 13259 1232 13290 1296
rect 13354 1232 13388 1296
rect 13259 1221 13388 1232
rect 13461 1295 13590 1306
rect 13461 1231 13492 1295
rect 13556 1231 13590 1295
rect 13461 1220 13590 1231
rect 13751 1296 13880 1307
rect 13751 1232 13782 1296
rect 13846 1232 13880 1296
rect 13751 1221 13880 1232
rect 14036 1295 14165 1306
rect 14036 1231 14067 1295
rect 14131 1231 14165 1295
rect 14036 1220 14165 1231
rect 15791 1300 15920 1311
rect 15791 1236 15822 1300
rect 15886 1236 15920 1300
rect 15791 1225 15920 1236
rect 15985 1304 16114 1315
rect 15985 1240 16016 1304
rect 16080 1240 16114 1304
rect 15985 1229 16114 1240
rect 16174 1301 16303 1312
rect 16174 1237 16205 1301
rect 16269 1237 16303 1301
rect 16174 1226 16303 1237
rect 16397 1303 16526 1314
rect 16397 1239 16428 1303
rect 16492 1239 16526 1303
rect 16397 1228 16526 1239
rect 228 1155 357 1166
rect 228 1091 259 1155
rect 323 1091 357 1155
rect 228 1080 357 1091
rect 430 1151 559 1162
rect 430 1087 461 1151
rect 525 1087 559 1151
rect 430 1076 559 1087
rect 619 1148 748 1159
rect 619 1084 650 1148
rect 714 1084 748 1148
rect 619 1073 748 1084
rect 848 1149 977 1160
rect 848 1085 879 1149
rect 943 1085 977 1149
rect 848 1074 977 1085
rect 2617 1152 2746 1163
rect 2617 1088 2648 1152
rect 2712 1088 2746 1152
rect 2617 1077 2746 1088
rect 2832 1149 2961 1160
rect 2832 1085 2863 1149
rect 2927 1085 2961 1149
rect 2832 1074 2961 1085
rect 3030 1146 3159 1157
rect 3030 1082 3061 1146
rect 3125 1082 3159 1146
rect 3030 1071 3159 1082
rect 3225 1156 3354 1167
rect 3225 1092 3256 1156
rect 3320 1092 3354 1156
rect 3225 1081 3354 1092
rect 3505 1154 3634 1165
rect 3505 1090 3536 1154
rect 3600 1090 3634 1154
rect 3505 1079 3634 1090
rect 3724 1152 3853 1163
rect 3724 1088 3755 1152
rect 3819 1088 3853 1152
rect 3724 1077 3853 1088
rect 5545 1149 5674 1160
rect 5545 1085 5576 1149
rect 5640 1085 5674 1149
rect 5545 1074 5674 1085
rect 5896 1146 6025 1157
rect 5896 1082 5927 1146
rect 5991 1082 6025 1146
rect 5896 1071 6025 1082
rect 6085 1144 6214 1155
rect 6085 1080 6116 1144
rect 6180 1080 6214 1144
rect 6085 1069 6214 1080
rect 6290 1151 6419 1162
rect 6290 1087 6321 1151
rect 6385 1087 6419 1151
rect 6290 1076 6419 1087
rect 6481 1153 6610 1164
rect 6481 1089 6512 1153
rect 6576 1089 6610 1153
rect 6481 1078 6610 1089
rect 8526 1155 8655 1166
rect 8526 1091 8557 1155
rect 8621 1091 8655 1155
rect 8526 1080 8655 1091
rect 8716 1157 8845 1168
rect 8716 1093 8747 1157
rect 8811 1093 8845 1157
rect 8716 1082 8845 1093
rect 8910 1155 9039 1166
rect 8910 1091 8941 1155
rect 9005 1091 9039 1155
rect 8910 1080 9039 1091
rect 9221 1151 9350 1162
rect 9221 1087 9252 1151
rect 9316 1087 9350 1151
rect 9221 1076 9350 1087
rect 11404 1150 11533 1161
rect 11404 1086 11435 1150
rect 11499 1086 11533 1150
rect 11404 1075 11533 1086
rect 11608 1150 11737 1161
rect 11608 1086 11639 1150
rect 11703 1086 11737 1150
rect 11608 1075 11737 1086
rect 12173 1146 12302 1157
rect 12173 1082 12204 1146
rect 12268 1082 12302 1146
rect 12173 1071 12302 1082
rect 12412 1148 12541 1159
rect 12412 1084 12443 1148
rect 12507 1084 12541 1148
rect 12412 1073 12541 1084
rect 12616 1148 12745 1159
rect 12616 1084 12647 1148
rect 12711 1084 12745 1148
rect 12616 1073 12745 1084
rect 14576 1156 14705 1167
rect 14576 1092 14607 1156
rect 14671 1092 14705 1156
rect 14576 1081 14705 1092
rect 14809 1154 14938 1165
rect 14809 1090 14840 1154
rect 14904 1090 14938 1154
rect 14809 1079 14938 1090
rect 15016 1152 15145 1163
rect 15016 1088 15047 1152
rect 15111 1088 15145 1152
rect 15016 1077 15145 1088
rect 15225 1154 15354 1165
rect 15225 1090 15256 1154
rect 15320 1090 15354 1154
rect 15225 1079 15354 1090
rect 15505 1156 15634 1167
rect 15505 1092 15536 1156
rect 15600 1092 15634 1156
rect 15505 1081 15634 1092
rect 1384 618 1513 629
rect 1155 606 1284 617
rect 1155 542 1186 606
rect 1250 542 1284 606
rect 1384 554 1415 618
rect 1479 554 1513 618
rect 1384 543 1513 554
rect 1603 608 1732 619
rect 1603 544 1634 608
rect 1698 544 1732 608
rect 1155 531 1284 542
rect 1603 533 1732 544
rect 1795 612 1924 623
rect 1795 548 1826 612
rect 1890 548 1924 612
rect 1795 537 1924 548
rect 2289 610 2418 621
rect 2289 546 2320 610
rect 2384 546 2418 610
rect 2289 535 2418 546
rect 4081 609 4210 620
rect 4081 545 4112 609
rect 4176 545 4210 609
rect 4081 534 4210 545
rect 4474 607 4603 618
rect 4474 543 4505 607
rect 4569 543 4603 607
rect 4474 532 4603 543
rect 4671 615 4800 626
rect 4671 551 4702 615
rect 4766 551 4800 615
rect 4671 540 4800 551
rect 5001 617 5130 628
rect 5001 553 5032 617
rect 5096 553 5130 617
rect 5001 542 5130 553
rect 5197 617 5326 628
rect 5197 553 5228 617
rect 5292 553 5326 617
rect 5197 542 5326 553
rect 7104 610 7233 621
rect 7104 546 7135 610
rect 7199 546 7233 610
rect 7104 535 7233 546
rect 7405 614 7534 625
rect 7405 550 7436 614
rect 7500 550 7534 614
rect 7405 539 7534 550
rect 7611 615 7740 626
rect 7611 551 7642 615
rect 7706 551 7740 615
rect 7611 540 7740 551
rect 7821 611 7950 622
rect 7821 547 7852 611
rect 7916 547 7950 611
rect 7821 536 7950 547
rect 8032 617 8161 628
rect 8032 553 8063 617
rect 8127 553 8161 617
rect 8032 542 8161 553
rect 9912 606 10041 617
rect 9912 542 9943 606
rect 10007 542 10041 606
rect 9912 531 10041 542
rect 10169 613 10298 624
rect 10169 549 10200 613
rect 10264 549 10298 613
rect 10169 538 10298 549
rect 10419 609 10548 620
rect 10419 545 10450 609
rect 10514 545 10548 609
rect 10419 534 10548 545
rect 10690 614 10819 625
rect 10690 550 10721 614
rect 10785 550 10819 614
rect 10690 539 10819 550
rect 10931 617 11060 628
rect 10931 553 10962 617
rect 11026 553 11060 617
rect 10931 542 11060 553
rect 11156 613 11285 624
rect 11156 549 11187 613
rect 11251 549 11285 613
rect 11156 538 11285 549
rect 12863 611 12992 622
rect 12863 547 12894 611
rect 12958 547 12992 611
rect 12863 536 12992 547
rect 13064 612 13193 623
rect 13064 548 13095 612
rect 13159 548 13193 612
rect 13064 537 13193 548
rect 13282 608 13411 619
rect 13282 544 13313 608
rect 13377 544 13411 608
rect 13282 533 13411 544
rect 13489 612 13618 623
rect 13489 548 13520 612
rect 13584 548 13618 612
rect 13489 537 13618 548
rect 13694 611 13823 622
rect 13694 547 13725 611
rect 13789 547 13823 611
rect 13694 536 13823 547
rect 14041 607 14170 618
rect 14041 543 14072 607
rect 14136 543 14170 607
rect 14041 532 14170 543
rect 15793 611 15922 622
rect 15793 547 15824 611
rect 15888 547 15922 611
rect 15793 536 15922 547
rect 15984 614 16113 625
rect 15984 550 16015 614
rect 16079 550 16113 614
rect 15984 539 16113 550
rect 16179 616 16308 627
rect 16179 552 16210 616
rect 16274 552 16308 616
rect 16179 541 16308 552
rect 16626 611 16755 622
rect 16626 547 16657 611
rect 16721 547 16755 611
rect 16626 536 16755 547
rect 10 462 139 473
rect 10 398 41 462
rect 105 398 139 462
rect 10 387 139 398
rect 243 458 372 469
rect 243 394 274 458
rect 338 394 372 458
rect 243 383 372 394
rect 458 465 587 476
rect 458 401 489 465
rect 553 401 587 465
rect 458 390 587 401
rect 676 462 805 473
rect 676 398 707 462
rect 771 398 805 462
rect 676 387 805 398
rect 892 463 1021 474
rect 892 399 923 463
rect 987 399 1021 463
rect 892 388 1021 399
rect 2613 459 2742 470
rect 2613 395 2644 459
rect 2708 395 2742 459
rect 2613 384 2742 395
rect 2803 459 2932 470
rect 2803 395 2834 459
rect 2898 395 2932 459
rect 2803 384 2932 395
rect 3013 462 3142 473
rect 3013 398 3044 462
rect 3108 398 3142 462
rect 3013 387 3142 398
rect 3230 459 3359 470
rect 3230 395 3261 459
rect 3325 395 3359 459
rect 3230 384 3359 395
rect 3525 462 3654 473
rect 3525 398 3556 462
rect 3620 398 3654 462
rect 3525 387 3654 398
rect 3749 467 3878 478
rect 3749 403 3780 467
rect 3844 403 3878 467
rect 3749 392 3878 403
rect 5627 460 5756 471
rect 5627 396 5658 460
rect 5722 396 5756 460
rect 5627 385 5756 396
rect 5927 458 6056 469
rect 5927 394 5958 458
rect 6022 394 6056 458
rect 5927 383 6056 394
rect 6179 462 6308 473
rect 6179 398 6210 462
rect 6274 398 6308 462
rect 6179 387 6308 398
rect 6396 467 6525 478
rect 6396 403 6427 467
rect 6491 403 6525 467
rect 6396 392 6525 403
rect 6597 464 6726 475
rect 6597 400 6628 464
rect 6692 400 6726 464
rect 6597 389 6726 400
rect 8482 455 8611 466
rect 8482 391 8513 455
rect 8577 391 8611 455
rect 8482 380 8611 391
rect 8674 455 8803 466
rect 8674 391 8705 455
rect 8769 391 8803 455
rect 8674 380 8803 391
rect 8874 455 9003 466
rect 8874 391 8905 455
rect 8969 391 9003 455
rect 8874 380 9003 391
rect 9492 463 9621 474
rect 9492 399 9523 463
rect 9587 399 9621 463
rect 9492 388 9621 399
rect 11393 459 11522 470
rect 11393 395 11424 459
rect 11488 395 11522 459
rect 11393 384 11522 395
rect 11649 459 11778 470
rect 11649 395 11680 459
rect 11744 395 11778 459
rect 11649 384 11778 395
rect 11884 459 12013 470
rect 11884 395 11915 459
rect 11979 395 12013 459
rect 11884 384 12013 395
rect 12173 461 12302 472
rect 12173 397 12204 461
rect 12268 397 12302 461
rect 12173 386 12302 397
rect 12363 459 12492 470
rect 12363 395 12394 459
rect 12458 395 12492 459
rect 12363 384 12492 395
rect 12567 461 12696 472
rect 12567 397 12598 461
rect 12662 397 12696 461
rect 12567 386 12696 397
rect 14353 467 14482 478
rect 14353 403 14384 467
rect 14448 403 14482 467
rect 14353 392 14482 403
rect 14595 463 14724 474
rect 14595 399 14626 463
rect 14690 399 14724 463
rect 14595 388 14724 399
rect 14795 462 14924 473
rect 14795 398 14826 462
rect 14890 398 14924 462
rect 14795 387 14924 398
rect 14985 470 15114 481
rect 14985 406 15016 470
rect 15080 406 15114 470
rect 14985 395 15114 406
rect 15206 468 15335 479
rect 15206 404 15237 468
rect 15301 404 15335 468
rect 15206 393 15335 404
rect 15502 463 15631 474
rect 15502 399 15533 463
rect 15597 399 15631 463
rect 15502 388 15631 399
rect 384 -70 513 -59
rect 384 -134 415 -70
rect 479 -134 513 -70
rect 384 -145 513 -134
rect 583 -73 712 -62
rect 583 -137 614 -73
rect 678 -137 712 -73
rect 583 -148 712 -137
rect 794 -73 923 -62
rect 794 -137 825 -73
rect 889 -137 923 -73
rect 794 -148 923 -137
rect 1000 -73 1129 -62
rect 1000 -137 1031 -73
rect 1095 -137 1129 -73
rect 1000 -148 1129 -137
rect 1228 -75 1357 -64
rect 1228 -139 1259 -75
rect 1323 -139 1357 -75
rect 1228 -150 1357 -139
rect 1472 -75 1601 -64
rect 1472 -139 1503 -75
rect 1567 -139 1601 -75
rect 1472 -150 1601 -139
rect 1702 -73 1831 -62
rect 1702 -137 1733 -73
rect 1797 -137 1831 -73
rect 1702 -148 1831 -137
rect 1908 -73 2037 -62
rect 1908 -137 1939 -73
rect 2003 -137 2037 -73
rect 1908 -148 2037 -137
rect 2126 -68 2255 -57
rect 2126 -132 2157 -68
rect 2221 -132 2255 -68
rect 2126 -143 2255 -132
rect 2329 -74 2458 -63
rect 2329 -138 2360 -74
rect 2424 -138 2458 -74
rect 2329 -149 2458 -138
rect 2537 -71 2666 -60
rect 2537 -135 2568 -71
rect 2632 -135 2666 -71
rect 2537 -146 2666 -135
rect 2800 -75 2929 -64
rect 2800 -139 2831 -75
rect 2895 -139 2929 -75
rect 2800 -150 2929 -139
rect 3008 -74 3137 -63
rect 3008 -138 3039 -74
rect 3103 -138 3137 -74
rect 3008 -149 3137 -138
rect 3218 -77 3347 -66
rect 3218 -141 3249 -77
rect 3313 -141 3347 -77
rect 3218 -152 3347 -141
rect 3418 -71 3547 -60
rect 3418 -135 3449 -71
rect 3513 -135 3547 -71
rect 3418 -146 3547 -135
rect 3621 -74 3750 -63
rect 3621 -138 3652 -74
rect 3716 -138 3750 -74
rect 3621 -149 3750 -138
rect 3831 -74 3960 -63
rect 3831 -138 3862 -74
rect 3926 -138 3960 -74
rect 3831 -149 3960 -138
rect 4032 -73 4161 -62
rect 4032 -137 4063 -73
rect 4127 -137 4161 -73
rect 4032 -148 4161 -137
rect 4248 -72 4377 -61
rect 4248 -136 4279 -72
rect 4343 -136 4377 -72
rect 4248 -147 4377 -136
rect 4529 -74 4658 -63
rect 4529 -138 4560 -74
rect 4624 -138 4658 -74
rect 4529 -149 4658 -138
rect 4749 -79 4878 -68
rect 4749 -143 4780 -79
rect 4844 -143 4878 -79
rect 4749 -154 4878 -143
rect 4954 -78 5083 -67
rect 4954 -142 4985 -78
rect 5049 -142 5083 -78
rect 4954 -153 5083 -142
rect 5175 -72 5304 -61
rect 5175 -136 5206 -72
rect 5270 -136 5304 -72
rect 5175 -147 5304 -136
rect 5380 -79 5509 -68
rect 5380 -143 5411 -79
rect 5475 -143 5509 -79
rect 5380 -154 5509 -143
rect 5589 -78 5718 -67
rect 5589 -142 5620 -78
rect 5684 -142 5718 -78
rect 5589 -153 5718 -142
rect 5806 -78 5935 -67
rect 5806 -142 5837 -78
rect 5901 -142 5935 -78
rect 5806 -153 5935 -142
rect 6020 -73 6149 -62
rect 6020 -137 6051 -73
rect 6115 -137 6149 -73
rect 6020 -148 6149 -137
rect 6215 -75 6344 -64
rect 6215 -139 6246 -75
rect 6310 -139 6344 -75
rect 6215 -150 6344 -139
rect 6410 -78 6539 -67
rect 6410 -142 6441 -78
rect 6505 -142 6539 -78
rect 6410 -153 6539 -142
rect 6612 -75 6741 -64
rect 6612 -139 6643 -75
rect 6707 -139 6741 -75
rect 6612 -150 6741 -139
rect 6896 -74 7025 -63
rect 6896 -138 6927 -74
rect 6991 -138 7025 -74
rect 6896 -149 7025 -138
rect 7095 -73 7224 -62
rect 7095 -137 7126 -73
rect 7190 -137 7224 -73
rect 7095 -148 7224 -137
rect 7298 -71 7427 -60
rect 7298 -135 7329 -71
rect 7393 -135 7427 -71
rect 7298 -146 7427 -135
rect 7563 -74 7692 -63
rect 7563 -138 7594 -74
rect 7658 -138 7692 -74
rect 7563 -149 7692 -138
rect 7761 -75 7890 -64
rect 7761 -139 7792 -75
rect 7856 -139 7890 -75
rect 7761 -150 7890 -139
rect 7950 -73 8079 -62
rect 7950 -137 7981 -73
rect 8045 -137 8079 -73
rect 7950 -148 8079 -137
rect 8162 -73 8291 -62
rect 8162 -137 8193 -73
rect 8257 -137 8291 -73
rect 8162 -148 8291 -137
rect 8379 -73 8508 -62
rect 8379 -137 8410 -73
rect 8474 -137 8508 -73
rect 8379 -148 8508 -137
rect 8584 -77 8713 -66
rect 8584 -141 8615 -77
rect 8679 -141 8713 -77
rect 8584 -152 8713 -141
rect 8789 -77 8918 -66
rect 8789 -141 8820 -77
rect 8884 -141 8918 -77
rect 8789 -152 8918 -141
rect 8997 -72 9126 -61
rect 8997 -136 9028 -72
rect 9092 -136 9126 -72
rect 8997 -147 9126 -136
rect 9280 -73 9409 -62
rect 9280 -137 9311 -73
rect 9375 -137 9409 -73
rect 9280 -148 9409 -137
rect 9473 -75 9602 -64
rect 9473 -139 9504 -75
rect 9568 -139 9602 -75
rect 9473 -150 9602 -139
rect 9699 -77 9828 -66
rect 9699 -141 9730 -77
rect 9794 -141 9828 -77
rect 9699 -152 9828 -141
rect 9964 -77 10093 -66
rect 9964 -141 9995 -77
rect 10059 -141 10093 -77
rect 9964 -152 10093 -141
rect 10158 -73 10287 -62
rect 10158 -137 10189 -73
rect 10253 -137 10287 -73
rect 10158 -148 10287 -137
rect 10356 -82 10485 -71
rect 10356 -146 10387 -82
rect 10451 -146 10485 -82
rect 10356 -157 10485 -146
rect 10560 -74 10689 -63
rect 10560 -138 10591 -74
rect 10655 -138 10689 -74
rect 10560 -149 10689 -138
rect 10780 -71 10909 -60
rect 10780 -135 10811 -71
rect 10875 -135 10909 -71
rect 10780 -146 10909 -135
rect 10995 -75 11124 -64
rect 10995 -139 11026 -75
rect 11090 -139 11124 -75
rect 10995 -150 11124 -139
rect 11223 -72 11352 -61
rect 11223 -136 11254 -72
rect 11318 -136 11352 -72
rect 11223 -147 11352 -136
rect 11427 -75 11556 -64
rect 11427 -139 11458 -75
rect 11522 -139 11556 -75
rect 11427 -150 11556 -139
rect 11665 -73 11794 -62
rect 11665 -137 11696 -73
rect 11760 -137 11794 -73
rect 11665 -148 11794 -137
rect 11858 -72 11987 -61
rect 11858 -136 11889 -72
rect 11953 -136 11987 -72
rect 11858 -147 11987 -136
rect 12055 -77 12184 -66
rect 12055 -141 12086 -77
rect 12150 -141 12184 -77
rect 12055 -152 12184 -141
rect 12311 -74 12440 -63
rect 12311 -138 12342 -74
rect 12406 -138 12440 -74
rect 12311 -149 12440 -138
rect 12550 -78 12679 -67
rect 12550 -142 12581 -78
rect 12645 -142 12679 -78
rect 12550 -153 12679 -142
rect 12783 -82 12912 -71
rect 12783 -146 12814 -82
rect 12878 -146 12912 -82
rect 12783 -157 12912 -146
rect 13004 -77 13133 -66
rect 13004 -141 13035 -77
rect 13099 -141 13133 -77
rect 13004 -152 13133 -141
rect 13195 -77 13324 -66
rect 13195 -141 13226 -77
rect 13290 -141 13324 -77
rect 13195 -152 13324 -141
rect 13423 -75 13552 -64
rect 13423 -139 13454 -75
rect 13518 -139 13552 -75
rect 13423 -150 13552 -139
rect 13620 -80 13749 -69
rect 13620 -144 13651 -80
rect 13715 -144 13749 -80
rect 13620 -155 13749 -144
rect 13832 -80 13961 -69
rect 13832 -144 13863 -80
rect 13927 -144 13961 -80
rect 13832 -155 13961 -144
rect 14059 -77 14188 -66
rect 14059 -141 14090 -77
rect 14154 -141 14188 -77
rect 14059 -152 14188 -141
rect 14248 -76 14377 -65
rect 14248 -140 14279 -76
rect 14343 -140 14377 -76
rect 14248 -151 14377 -140
rect 14474 -75 14603 -64
rect 14474 -139 14505 -75
rect 14569 -139 14603 -75
rect 14474 -150 14603 -139
rect 14728 -75 14857 -64
rect 14728 -139 14759 -75
rect 14823 -139 14857 -75
rect 14728 -150 14857 -139
rect 14972 -78 15101 -67
rect 14972 -142 15003 -78
rect 15067 -142 15101 -78
rect 14972 -153 15101 -142
rect 15202 -79 15331 -68
rect 15202 -143 15233 -79
rect 15297 -143 15331 -79
rect 15202 -154 15331 -143
rect 15460 -76 15589 -65
rect 15460 -140 15491 -76
rect 15555 -140 15589 -76
rect 15460 -151 15589 -140
rect 15670 -76 15799 -65
rect 15670 -140 15701 -76
rect 15765 -140 15799 -76
rect 15670 -151 15799 -140
rect 15895 -76 16024 -65
rect 15895 -140 15926 -76
rect 15990 -140 16024 -76
rect 15895 -151 16024 -140
rect 16114 -79 16243 -68
rect 16114 -143 16145 -79
rect 16209 -143 16243 -79
rect 16114 -154 16243 -143
rect 16460 -75 16589 -64
rect 16460 -139 16491 -75
rect 16555 -139 16589 -75
rect 16460 -150 16589 -139
rect 16659 -78 16788 -67
rect 16659 -142 16690 -78
rect 16754 -142 16788 -78
rect 16659 -153 16788 -142
<< via3 >>
rect 717 3437 781 3441
rect 717 3381 721 3437
rect 721 3381 777 3437
rect 777 3381 781 3437
rect 717 3377 781 3381
rect 47 2978 111 2982
rect 47 2922 51 2978
rect 51 2922 107 2978
rect 107 2922 111 2978
rect 47 2918 111 2922
rect 249 2980 313 2984
rect 249 2924 253 2980
rect 253 2924 309 2980
rect 309 2924 313 2980
rect 249 2920 313 2924
rect 460 2978 524 2982
rect 460 2922 464 2978
rect 464 2922 520 2978
rect 520 2922 524 2978
rect 460 2918 524 2922
rect 650 2978 714 2982
rect 650 2922 654 2978
rect 654 2922 710 2978
rect 710 2922 714 2978
rect 650 2918 714 2922
rect 858 2980 922 2984
rect 858 2924 862 2980
rect 862 2924 918 2980
rect 918 2924 922 2980
rect 858 2920 922 2924
rect 1060 2980 1124 2984
rect 1060 2924 1064 2980
rect 1064 2924 1120 2980
rect 1120 2924 1124 2980
rect 1060 2920 1124 2924
rect 1259 2982 1323 2986
rect 1259 2926 1263 2982
rect 1263 2926 1319 2982
rect 1319 2926 1323 2982
rect 1259 2922 1323 2926
rect 1454 2979 1518 2983
rect 1454 2923 1458 2979
rect 1458 2923 1514 2979
rect 1514 2923 1518 2979
rect 1454 2919 1518 2923
rect 1655 2981 1719 2985
rect 1655 2925 1659 2981
rect 1659 2925 1715 2981
rect 1715 2925 1719 2981
rect 1655 2921 1719 2925
rect 1872 2979 1936 2983
rect 1872 2923 1876 2979
rect 1876 2923 1932 2979
rect 1932 2923 1936 2979
rect 1872 2919 1936 2923
rect 2146 2982 2210 2986
rect 2146 2926 2150 2982
rect 2150 2926 2206 2982
rect 2206 2926 2210 2982
rect 2146 2922 2210 2926
rect 2423 2975 2487 2979
rect 2423 2919 2427 2975
rect 2427 2919 2483 2975
rect 2483 2919 2487 2975
rect 2423 2915 2487 2919
rect 2646 2978 2710 2982
rect 2646 2922 2650 2978
rect 2650 2922 2706 2978
rect 2706 2922 2710 2978
rect 2646 2918 2710 2922
rect 2878 2977 2942 2981
rect 2878 2921 2882 2977
rect 2882 2921 2938 2977
rect 2938 2921 2942 2977
rect 2878 2917 2942 2921
rect 4514 2974 4578 2978
rect 4514 2918 4518 2974
rect 4518 2918 4574 2974
rect 4574 2918 4578 2974
rect 4514 2914 4578 2918
rect 4822 2975 4886 2979
rect 4822 2919 4826 2975
rect 4826 2919 4882 2975
rect 4882 2919 4886 2975
rect 4822 2915 4886 2919
rect 5022 2976 5086 2980
rect 5022 2920 5026 2976
rect 5026 2920 5082 2976
rect 5082 2920 5086 2976
rect 5022 2916 5086 2920
rect 5241 2975 5305 2979
rect 5241 2919 5245 2975
rect 5245 2919 5301 2975
rect 5301 2919 5305 2975
rect 5241 2915 5305 2919
rect 5487 2974 5551 2978
rect 5487 2918 5491 2974
rect 5491 2918 5547 2974
rect 5547 2918 5551 2974
rect 5487 2914 5551 2918
rect 5695 2976 5759 2980
rect 5695 2920 5699 2976
rect 5699 2920 5755 2976
rect 5755 2920 5759 2976
rect 5695 2916 5759 2920
rect 5897 2977 5961 2981
rect 5897 2921 5901 2977
rect 5901 2921 5957 2977
rect 5957 2921 5961 2977
rect 5897 2917 5961 2921
rect 6090 2976 6154 2980
rect 6090 2920 6094 2976
rect 6094 2920 6150 2976
rect 6150 2920 6154 2976
rect 6090 2916 6154 2920
rect 6462 2975 6526 2979
rect 6462 2919 6466 2975
rect 6466 2919 6522 2975
rect 6522 2919 6526 2975
rect 6462 2915 6526 2919
rect 6651 2973 6715 2977
rect 6651 2917 6655 2973
rect 6655 2917 6711 2973
rect 6711 2917 6715 2973
rect 6651 2913 6715 2917
rect 6941 2973 7005 2977
rect 6941 2917 6945 2973
rect 6945 2917 7001 2973
rect 7001 2917 7005 2973
rect 6941 2913 7005 2917
rect 7214 2975 7278 2979
rect 7214 2919 7218 2975
rect 7218 2919 7274 2975
rect 7274 2919 7278 2975
rect 7214 2915 7278 2919
rect 1165 2439 1229 2443
rect 1165 2383 1169 2439
rect 1169 2383 1225 2439
rect 1225 2383 1229 2439
rect 1165 2379 1229 2383
rect 1384 2443 1448 2447
rect 1384 2387 1388 2443
rect 1388 2387 1444 2443
rect 1444 2387 1448 2443
rect 1384 2383 1448 2387
rect 1667 2443 1731 2447
rect 1667 2387 1671 2443
rect 1671 2387 1727 2443
rect 1727 2387 1731 2443
rect 1667 2383 1731 2387
rect 1876 2443 1940 2447
rect 1876 2387 1880 2443
rect 1880 2387 1936 2443
rect 1936 2387 1940 2443
rect 1876 2383 1940 2387
rect 2147 2441 2211 2445
rect 2147 2385 2151 2441
rect 2151 2385 2207 2441
rect 2207 2385 2211 2441
rect 2147 2381 2211 2385
rect 4222 2439 4286 2443
rect 4222 2383 4226 2439
rect 4226 2383 4282 2439
rect 4282 2383 4286 2439
rect 4222 2379 4286 2383
rect 4471 2442 4535 2446
rect 4471 2386 4475 2442
rect 4475 2386 4531 2442
rect 4531 2386 4535 2442
rect 4471 2382 4535 2386
rect 4815 2428 4879 2432
rect 4815 2372 4819 2428
rect 4819 2372 4875 2428
rect 4875 2372 4879 2428
rect 4815 2368 4879 2372
rect 5069 2434 5133 2438
rect 5069 2378 5073 2434
rect 5073 2378 5129 2434
rect 5129 2378 5133 2434
rect 5069 2374 5133 2378
rect 5298 2434 5362 2438
rect 5298 2378 5302 2434
rect 5302 2378 5358 2434
rect 5358 2378 5362 2434
rect 5298 2374 5362 2378
rect 7016 2439 7080 2443
rect 7016 2383 7020 2439
rect 7020 2383 7076 2439
rect 7076 2383 7080 2439
rect 7016 2379 7080 2383
rect 7220 2441 7284 2445
rect 7220 2385 7224 2441
rect 7224 2385 7280 2441
rect 7280 2385 7284 2441
rect 7220 2381 7284 2385
rect 7543 2439 7607 2443
rect 7543 2383 7547 2439
rect 7547 2383 7603 2439
rect 7603 2383 7607 2439
rect 7543 2379 7607 2383
rect 13 1834 77 1838
rect 13 1778 17 1834
rect 17 1778 73 1834
rect 73 1778 77 1834
rect 13 1774 77 1778
rect 253 1832 317 1836
rect 253 1776 257 1832
rect 257 1776 313 1832
rect 313 1776 317 1832
rect 253 1772 317 1776
rect 575 1831 639 1835
rect 575 1775 579 1831
rect 579 1775 635 1831
rect 635 1775 639 1831
rect 575 1771 639 1775
rect 793 1832 857 1836
rect 793 1776 797 1832
rect 797 1776 853 1832
rect 853 1776 857 1832
rect 793 1772 857 1776
rect 2697 1836 2761 1840
rect 2697 1780 2701 1836
rect 2701 1780 2757 1836
rect 2757 1780 2761 1836
rect 2697 1776 2761 1780
rect 3022 1838 3086 1842
rect 3022 1782 3026 1838
rect 3026 1782 3082 1838
rect 3082 1782 3086 1838
rect 3022 1778 3086 1782
rect 3290 1838 3354 1842
rect 3290 1782 3294 1838
rect 3294 1782 3350 1838
rect 3350 1782 3354 1838
rect 3290 1778 3354 1782
rect 3556 1838 3620 1842
rect 3556 1782 3560 1838
rect 3560 1782 3616 1838
rect 3616 1782 3620 1838
rect 3556 1778 3620 1782
rect 3796 1836 3860 1840
rect 3796 1780 3800 1836
rect 3800 1780 3856 1836
rect 3856 1780 3860 1836
rect 3796 1776 3860 1780
rect 5590 1839 5654 1843
rect 5590 1783 5594 1839
rect 5594 1783 5650 1839
rect 5650 1783 5654 1839
rect 5590 1779 5654 1783
rect 5956 1842 6020 1846
rect 5956 1786 5960 1842
rect 5960 1786 6016 1842
rect 6016 1786 6020 1842
rect 5956 1782 6020 1786
rect 6200 1842 6264 1846
rect 6200 1786 6204 1842
rect 6204 1786 6260 1842
rect 6260 1786 6264 1842
rect 6200 1782 6264 1786
rect 6623 1833 6687 1837
rect 6623 1777 6627 1833
rect 6627 1777 6683 1833
rect 6683 1777 6687 1833
rect 6623 1773 6687 1777
rect 8566 1835 8630 1839
rect 8566 1779 8570 1835
rect 8570 1779 8626 1835
rect 8626 1779 8630 1835
rect 8566 1775 8630 1779
rect 8818 1832 8882 1836
rect 8818 1776 8822 1832
rect 8822 1776 8878 1832
rect 8878 1776 8882 1832
rect 8818 1772 8882 1776
rect 9024 1840 9088 1844
rect 9024 1784 9028 1840
rect 9028 1784 9084 1840
rect 9084 1784 9088 1840
rect 9024 1780 9088 1784
rect 9307 1834 9371 1838
rect 9307 1778 9311 1834
rect 9311 1778 9367 1834
rect 9367 1778 9371 1834
rect 9307 1774 9371 1778
rect 9605 1835 9669 1839
rect 9605 1779 9609 1835
rect 9609 1779 9665 1835
rect 9665 1779 9669 1835
rect 9605 1775 9669 1779
rect 11437 1836 11501 1840
rect 11437 1780 11441 1836
rect 11441 1780 11497 1836
rect 11497 1780 11501 1836
rect 11437 1776 11501 1780
rect 11647 1838 11711 1842
rect 11647 1782 11651 1838
rect 11651 1782 11707 1838
rect 11707 1782 11711 1838
rect 11647 1778 11711 1782
rect 11998 1836 12062 1840
rect 11998 1780 12002 1836
rect 12002 1780 12058 1836
rect 12058 1780 12062 1836
rect 11998 1776 12062 1780
rect 12278 1836 12342 1840
rect 12278 1780 12282 1836
rect 12282 1780 12338 1836
rect 12338 1780 12342 1836
rect 12278 1776 12342 1780
rect 12595 1835 12659 1839
rect 12595 1779 12599 1835
rect 12599 1779 12655 1835
rect 12655 1779 12659 1835
rect 12595 1775 12659 1779
rect 14385 1833 14449 1837
rect 14385 1777 14389 1833
rect 14389 1777 14445 1833
rect 14445 1777 14449 1833
rect 14385 1773 14449 1777
rect 14680 1833 14744 1837
rect 14680 1777 14684 1833
rect 14684 1777 14740 1833
rect 14740 1777 14744 1833
rect 14680 1773 14744 1777
rect 14967 1833 15031 1837
rect 14967 1777 14971 1833
rect 14971 1777 15027 1833
rect 15027 1777 15031 1833
rect 14967 1773 15031 1777
rect 15257 1833 15321 1837
rect 15257 1777 15261 1833
rect 15261 1777 15317 1833
rect 15317 1777 15321 1833
rect 15257 1773 15321 1777
rect 15541 1836 15605 1840
rect 15541 1780 15545 1836
rect 15545 1780 15601 1836
rect 15601 1780 15605 1836
rect 15541 1776 15605 1780
rect 1204 1296 1268 1300
rect 1204 1240 1208 1296
rect 1208 1240 1264 1296
rect 1264 1240 1268 1296
rect 1204 1236 1268 1240
rect 1421 1296 1485 1300
rect 1421 1240 1425 1296
rect 1425 1240 1481 1296
rect 1481 1240 1485 1296
rect 1421 1236 1485 1240
rect 1640 1296 1704 1300
rect 1640 1240 1644 1296
rect 1644 1240 1700 1296
rect 1700 1240 1704 1296
rect 1640 1236 1704 1240
rect 1853 1292 1917 1296
rect 1853 1236 1857 1292
rect 1857 1236 1913 1292
rect 1913 1236 1917 1292
rect 1853 1232 1917 1236
rect 2064 1292 2128 1296
rect 2064 1236 2068 1292
rect 2068 1236 2124 1292
rect 2124 1236 2128 1292
rect 2064 1232 2128 1236
rect 4188 1292 4252 1296
rect 4188 1236 4192 1292
rect 4192 1236 4248 1292
rect 4248 1236 4252 1292
rect 4188 1232 4252 1236
rect 4466 1291 4530 1295
rect 4466 1235 4470 1291
rect 4470 1235 4526 1291
rect 4526 1235 4530 1291
rect 4466 1231 4530 1235
rect 5038 1296 5102 1300
rect 5038 1240 5042 1296
rect 5042 1240 5098 1296
rect 5098 1240 5102 1296
rect 5038 1236 5102 1240
rect 5277 1296 5341 1300
rect 5277 1240 5281 1296
rect 5281 1240 5337 1296
rect 5337 1240 5341 1296
rect 5277 1236 5341 1240
rect 7435 1294 7499 1298
rect 7435 1238 7439 1294
rect 7439 1238 7495 1294
rect 7495 1238 7499 1294
rect 7435 1234 7499 1238
rect 7662 1299 7726 1303
rect 7662 1243 7666 1299
rect 7666 1243 7722 1299
rect 7722 1243 7726 1299
rect 7662 1239 7726 1243
rect 7852 1301 7916 1305
rect 7852 1245 7856 1301
rect 7856 1245 7912 1301
rect 7912 1245 7916 1301
rect 7852 1241 7916 1245
rect 8068 1292 8132 1296
rect 8068 1236 8072 1292
rect 8072 1236 8128 1292
rect 8128 1236 8132 1292
rect 8068 1232 8132 1236
rect 10049 1295 10113 1299
rect 10049 1239 10053 1295
rect 10053 1239 10109 1295
rect 10109 1239 10113 1295
rect 10049 1235 10113 1239
rect 10278 1298 10342 1302
rect 10278 1242 10282 1298
rect 10282 1242 10338 1298
rect 10338 1242 10342 1298
rect 10278 1238 10342 1242
rect 10504 1303 10568 1307
rect 10504 1247 10508 1303
rect 10508 1247 10564 1303
rect 10564 1247 10568 1303
rect 10504 1243 10568 1247
rect 10732 1295 10796 1299
rect 10732 1239 10736 1295
rect 10736 1239 10792 1295
rect 10792 1239 10796 1295
rect 10732 1235 10796 1239
rect 10968 1301 11032 1305
rect 10968 1245 10972 1301
rect 10972 1245 11028 1301
rect 11028 1245 11032 1301
rect 10968 1241 11032 1245
rect 11160 1292 11224 1296
rect 11160 1236 11164 1292
rect 11164 1236 11220 1292
rect 11220 1236 11224 1292
rect 11160 1232 11224 1236
rect 12895 1292 12959 1296
rect 12895 1236 12899 1292
rect 12899 1236 12955 1292
rect 12955 1236 12959 1292
rect 12895 1232 12959 1236
rect 13099 1297 13163 1301
rect 13099 1241 13103 1297
rect 13103 1241 13159 1297
rect 13159 1241 13163 1297
rect 13099 1237 13163 1241
rect 13290 1292 13354 1296
rect 13290 1236 13294 1292
rect 13294 1236 13350 1292
rect 13350 1236 13354 1292
rect 13290 1232 13354 1236
rect 13492 1291 13556 1295
rect 13492 1235 13496 1291
rect 13496 1235 13552 1291
rect 13552 1235 13556 1291
rect 13492 1231 13556 1235
rect 13782 1292 13846 1296
rect 13782 1236 13786 1292
rect 13786 1236 13842 1292
rect 13842 1236 13846 1292
rect 13782 1232 13846 1236
rect 14067 1291 14131 1295
rect 14067 1235 14071 1291
rect 14071 1235 14127 1291
rect 14127 1235 14131 1291
rect 14067 1231 14131 1235
rect 15822 1296 15886 1300
rect 15822 1240 15826 1296
rect 15826 1240 15882 1296
rect 15882 1240 15886 1296
rect 15822 1236 15886 1240
rect 16016 1300 16080 1304
rect 16016 1244 16020 1300
rect 16020 1244 16076 1300
rect 16076 1244 16080 1300
rect 16016 1240 16080 1244
rect 16205 1297 16269 1301
rect 16205 1241 16209 1297
rect 16209 1241 16265 1297
rect 16265 1241 16269 1297
rect 16205 1237 16269 1241
rect 16428 1299 16492 1303
rect 16428 1243 16432 1299
rect 16432 1243 16488 1299
rect 16488 1243 16492 1299
rect 16428 1239 16492 1243
rect 259 1151 323 1155
rect 259 1095 263 1151
rect 263 1095 319 1151
rect 319 1095 323 1151
rect 259 1091 323 1095
rect 461 1147 525 1151
rect 461 1091 465 1147
rect 465 1091 521 1147
rect 521 1091 525 1147
rect 461 1087 525 1091
rect 650 1144 714 1148
rect 650 1088 654 1144
rect 654 1088 710 1144
rect 710 1088 714 1144
rect 650 1084 714 1088
rect 879 1145 943 1149
rect 879 1089 883 1145
rect 883 1089 939 1145
rect 939 1089 943 1145
rect 879 1085 943 1089
rect 2648 1148 2712 1152
rect 2648 1092 2652 1148
rect 2652 1092 2708 1148
rect 2708 1092 2712 1148
rect 2648 1088 2712 1092
rect 2863 1145 2927 1149
rect 2863 1089 2867 1145
rect 2867 1089 2923 1145
rect 2923 1089 2927 1145
rect 2863 1085 2927 1089
rect 3061 1142 3125 1146
rect 3061 1086 3065 1142
rect 3065 1086 3121 1142
rect 3121 1086 3125 1142
rect 3061 1082 3125 1086
rect 3256 1152 3320 1156
rect 3256 1096 3260 1152
rect 3260 1096 3316 1152
rect 3316 1096 3320 1152
rect 3256 1092 3320 1096
rect 3536 1150 3600 1154
rect 3536 1094 3540 1150
rect 3540 1094 3596 1150
rect 3596 1094 3600 1150
rect 3536 1090 3600 1094
rect 3755 1148 3819 1152
rect 3755 1092 3759 1148
rect 3759 1092 3815 1148
rect 3815 1092 3819 1148
rect 3755 1088 3819 1092
rect 5576 1145 5640 1149
rect 5576 1089 5580 1145
rect 5580 1089 5636 1145
rect 5636 1089 5640 1145
rect 5576 1085 5640 1089
rect 5927 1142 5991 1146
rect 5927 1086 5931 1142
rect 5931 1086 5987 1142
rect 5987 1086 5991 1142
rect 5927 1082 5991 1086
rect 6116 1140 6180 1144
rect 6116 1084 6120 1140
rect 6120 1084 6176 1140
rect 6176 1084 6180 1140
rect 6116 1080 6180 1084
rect 6321 1147 6385 1151
rect 6321 1091 6325 1147
rect 6325 1091 6381 1147
rect 6381 1091 6385 1147
rect 6321 1087 6385 1091
rect 6512 1149 6576 1153
rect 6512 1093 6516 1149
rect 6516 1093 6572 1149
rect 6572 1093 6576 1149
rect 6512 1089 6576 1093
rect 8557 1151 8621 1155
rect 8557 1095 8561 1151
rect 8561 1095 8617 1151
rect 8617 1095 8621 1151
rect 8557 1091 8621 1095
rect 8747 1153 8811 1157
rect 8747 1097 8751 1153
rect 8751 1097 8807 1153
rect 8807 1097 8811 1153
rect 8747 1093 8811 1097
rect 8941 1151 9005 1155
rect 8941 1095 8945 1151
rect 8945 1095 9001 1151
rect 9001 1095 9005 1151
rect 8941 1091 9005 1095
rect 9252 1147 9316 1151
rect 9252 1091 9256 1147
rect 9256 1091 9312 1147
rect 9312 1091 9316 1147
rect 9252 1087 9316 1091
rect 11435 1146 11499 1150
rect 11435 1090 11439 1146
rect 11439 1090 11495 1146
rect 11495 1090 11499 1146
rect 11435 1086 11499 1090
rect 11639 1146 11703 1150
rect 11639 1090 11643 1146
rect 11643 1090 11699 1146
rect 11699 1090 11703 1146
rect 11639 1086 11703 1090
rect 12204 1142 12268 1146
rect 12204 1086 12208 1142
rect 12208 1086 12264 1142
rect 12264 1086 12268 1142
rect 12204 1082 12268 1086
rect 12443 1144 12507 1148
rect 12443 1088 12447 1144
rect 12447 1088 12503 1144
rect 12503 1088 12507 1144
rect 12443 1084 12507 1088
rect 12647 1144 12711 1148
rect 12647 1088 12651 1144
rect 12651 1088 12707 1144
rect 12707 1088 12711 1144
rect 12647 1084 12711 1088
rect 14607 1152 14671 1156
rect 14607 1096 14611 1152
rect 14611 1096 14667 1152
rect 14667 1096 14671 1152
rect 14607 1092 14671 1096
rect 14840 1150 14904 1154
rect 14840 1094 14844 1150
rect 14844 1094 14900 1150
rect 14900 1094 14904 1150
rect 14840 1090 14904 1094
rect 15047 1148 15111 1152
rect 15047 1092 15051 1148
rect 15051 1092 15107 1148
rect 15107 1092 15111 1148
rect 15047 1088 15111 1092
rect 15256 1150 15320 1154
rect 15256 1094 15260 1150
rect 15260 1094 15316 1150
rect 15316 1094 15320 1150
rect 15256 1090 15320 1094
rect 15536 1152 15600 1156
rect 15536 1096 15540 1152
rect 15540 1096 15596 1152
rect 15596 1096 15600 1152
rect 15536 1092 15600 1096
rect 1186 602 1250 606
rect 1186 546 1190 602
rect 1190 546 1246 602
rect 1246 546 1250 602
rect 1186 542 1250 546
rect 1415 614 1479 618
rect 1415 558 1419 614
rect 1419 558 1475 614
rect 1475 558 1479 614
rect 1415 554 1479 558
rect 1634 604 1698 608
rect 1634 548 1638 604
rect 1638 548 1694 604
rect 1694 548 1698 604
rect 1634 544 1698 548
rect 1826 608 1890 612
rect 1826 552 1830 608
rect 1830 552 1886 608
rect 1886 552 1890 608
rect 1826 548 1890 552
rect 2320 606 2384 610
rect 2320 550 2324 606
rect 2324 550 2380 606
rect 2380 550 2384 606
rect 2320 546 2384 550
rect 4112 605 4176 609
rect 4112 549 4116 605
rect 4116 549 4172 605
rect 4172 549 4176 605
rect 4112 545 4176 549
rect 4505 603 4569 607
rect 4505 547 4509 603
rect 4509 547 4565 603
rect 4565 547 4569 603
rect 4505 543 4569 547
rect 4702 611 4766 615
rect 4702 555 4706 611
rect 4706 555 4762 611
rect 4762 555 4766 611
rect 4702 551 4766 555
rect 5032 613 5096 617
rect 5032 557 5036 613
rect 5036 557 5092 613
rect 5092 557 5096 613
rect 5032 553 5096 557
rect 5228 613 5292 617
rect 5228 557 5232 613
rect 5232 557 5288 613
rect 5288 557 5292 613
rect 5228 553 5292 557
rect 7135 606 7199 610
rect 7135 550 7139 606
rect 7139 550 7195 606
rect 7195 550 7199 606
rect 7135 546 7199 550
rect 7436 610 7500 614
rect 7436 554 7440 610
rect 7440 554 7496 610
rect 7496 554 7500 610
rect 7436 550 7500 554
rect 7642 611 7706 615
rect 7642 555 7646 611
rect 7646 555 7702 611
rect 7702 555 7706 611
rect 7642 551 7706 555
rect 7852 607 7916 611
rect 7852 551 7856 607
rect 7856 551 7912 607
rect 7912 551 7916 607
rect 7852 547 7916 551
rect 8063 613 8127 617
rect 8063 557 8067 613
rect 8067 557 8123 613
rect 8123 557 8127 613
rect 8063 553 8127 557
rect 9943 602 10007 606
rect 9943 546 9947 602
rect 9947 546 10003 602
rect 10003 546 10007 602
rect 9943 542 10007 546
rect 10200 609 10264 613
rect 10200 553 10204 609
rect 10204 553 10260 609
rect 10260 553 10264 609
rect 10200 549 10264 553
rect 10450 605 10514 609
rect 10450 549 10454 605
rect 10454 549 10510 605
rect 10510 549 10514 605
rect 10450 545 10514 549
rect 10721 610 10785 614
rect 10721 554 10725 610
rect 10725 554 10781 610
rect 10781 554 10785 610
rect 10721 550 10785 554
rect 10962 613 11026 617
rect 10962 557 10966 613
rect 10966 557 11022 613
rect 11022 557 11026 613
rect 10962 553 11026 557
rect 11187 609 11251 613
rect 11187 553 11191 609
rect 11191 553 11247 609
rect 11247 553 11251 609
rect 11187 549 11251 553
rect 12894 607 12958 611
rect 12894 551 12898 607
rect 12898 551 12954 607
rect 12954 551 12958 607
rect 12894 547 12958 551
rect 13095 608 13159 612
rect 13095 552 13099 608
rect 13099 552 13155 608
rect 13155 552 13159 608
rect 13095 548 13159 552
rect 13313 604 13377 608
rect 13313 548 13317 604
rect 13317 548 13373 604
rect 13373 548 13377 604
rect 13313 544 13377 548
rect 13520 608 13584 612
rect 13520 552 13524 608
rect 13524 552 13580 608
rect 13580 552 13584 608
rect 13520 548 13584 552
rect 13725 607 13789 611
rect 13725 551 13729 607
rect 13729 551 13785 607
rect 13785 551 13789 607
rect 13725 547 13789 551
rect 14072 603 14136 607
rect 14072 547 14076 603
rect 14076 547 14132 603
rect 14132 547 14136 603
rect 14072 543 14136 547
rect 15824 607 15888 611
rect 15824 551 15828 607
rect 15828 551 15884 607
rect 15884 551 15888 607
rect 15824 547 15888 551
rect 16015 610 16079 614
rect 16015 554 16019 610
rect 16019 554 16075 610
rect 16075 554 16079 610
rect 16015 550 16079 554
rect 16210 612 16274 616
rect 16210 556 16214 612
rect 16214 556 16270 612
rect 16270 556 16274 612
rect 16210 552 16274 556
rect 16657 607 16721 611
rect 16657 551 16661 607
rect 16661 551 16717 607
rect 16717 551 16721 607
rect 16657 547 16721 551
rect 41 458 105 462
rect 41 402 45 458
rect 45 402 101 458
rect 101 402 105 458
rect 41 398 105 402
rect 274 454 338 458
rect 274 398 278 454
rect 278 398 334 454
rect 334 398 338 454
rect 274 394 338 398
rect 489 461 553 465
rect 489 405 493 461
rect 493 405 549 461
rect 549 405 553 461
rect 489 401 553 405
rect 707 458 771 462
rect 707 402 711 458
rect 711 402 767 458
rect 767 402 771 458
rect 707 398 771 402
rect 923 459 987 463
rect 923 403 927 459
rect 927 403 983 459
rect 983 403 987 459
rect 923 399 987 403
rect 2644 455 2708 459
rect 2644 399 2648 455
rect 2648 399 2704 455
rect 2704 399 2708 455
rect 2644 395 2708 399
rect 2834 455 2898 459
rect 2834 399 2838 455
rect 2838 399 2894 455
rect 2894 399 2898 455
rect 2834 395 2898 399
rect 3044 458 3108 462
rect 3044 402 3048 458
rect 3048 402 3104 458
rect 3104 402 3108 458
rect 3044 398 3108 402
rect 3261 455 3325 459
rect 3261 399 3265 455
rect 3265 399 3321 455
rect 3321 399 3325 455
rect 3261 395 3325 399
rect 3556 458 3620 462
rect 3556 402 3560 458
rect 3560 402 3616 458
rect 3616 402 3620 458
rect 3556 398 3620 402
rect 3780 463 3844 467
rect 3780 407 3784 463
rect 3784 407 3840 463
rect 3840 407 3844 463
rect 3780 403 3844 407
rect 5658 456 5722 460
rect 5658 400 5662 456
rect 5662 400 5718 456
rect 5718 400 5722 456
rect 5658 396 5722 400
rect 5958 454 6022 458
rect 5958 398 5962 454
rect 5962 398 6018 454
rect 6018 398 6022 454
rect 5958 394 6022 398
rect 6210 458 6274 462
rect 6210 402 6214 458
rect 6214 402 6270 458
rect 6270 402 6274 458
rect 6210 398 6274 402
rect 6427 463 6491 467
rect 6427 407 6431 463
rect 6431 407 6487 463
rect 6487 407 6491 463
rect 6427 403 6491 407
rect 6628 460 6692 464
rect 6628 404 6632 460
rect 6632 404 6688 460
rect 6688 404 6692 460
rect 6628 400 6692 404
rect 8513 451 8577 455
rect 8513 395 8517 451
rect 8517 395 8573 451
rect 8573 395 8577 451
rect 8513 391 8577 395
rect 8705 451 8769 455
rect 8705 395 8709 451
rect 8709 395 8765 451
rect 8765 395 8769 451
rect 8705 391 8769 395
rect 8905 451 8969 455
rect 8905 395 8909 451
rect 8909 395 8965 451
rect 8965 395 8969 451
rect 8905 391 8969 395
rect 9523 459 9587 463
rect 9523 403 9527 459
rect 9527 403 9583 459
rect 9583 403 9587 459
rect 9523 399 9587 403
rect 11424 455 11488 459
rect 11424 399 11428 455
rect 11428 399 11484 455
rect 11484 399 11488 455
rect 11424 395 11488 399
rect 11680 455 11744 459
rect 11680 399 11684 455
rect 11684 399 11740 455
rect 11740 399 11744 455
rect 11680 395 11744 399
rect 11915 455 11979 459
rect 11915 399 11919 455
rect 11919 399 11975 455
rect 11975 399 11979 455
rect 11915 395 11979 399
rect 12204 457 12268 461
rect 12204 401 12208 457
rect 12208 401 12264 457
rect 12264 401 12268 457
rect 12204 397 12268 401
rect 12394 455 12458 459
rect 12394 399 12398 455
rect 12398 399 12454 455
rect 12454 399 12458 455
rect 12394 395 12458 399
rect 12598 457 12662 461
rect 12598 401 12602 457
rect 12602 401 12658 457
rect 12658 401 12662 457
rect 12598 397 12662 401
rect 14384 463 14448 467
rect 14384 407 14388 463
rect 14388 407 14444 463
rect 14444 407 14448 463
rect 14384 403 14448 407
rect 14626 459 14690 463
rect 14626 403 14630 459
rect 14630 403 14686 459
rect 14686 403 14690 459
rect 14626 399 14690 403
rect 14826 458 14890 462
rect 14826 402 14830 458
rect 14830 402 14886 458
rect 14886 402 14890 458
rect 14826 398 14890 402
rect 15016 466 15080 470
rect 15016 410 15020 466
rect 15020 410 15076 466
rect 15076 410 15080 466
rect 15016 406 15080 410
rect 15237 464 15301 468
rect 15237 408 15241 464
rect 15241 408 15297 464
rect 15297 408 15301 464
rect 15237 404 15301 408
rect 15533 459 15597 463
rect 15533 403 15537 459
rect 15537 403 15593 459
rect 15593 403 15597 459
rect 15533 399 15597 403
rect 415 -74 479 -70
rect 415 -130 419 -74
rect 419 -130 475 -74
rect 475 -130 479 -74
rect 415 -134 479 -130
rect 614 -77 678 -73
rect 614 -133 618 -77
rect 618 -133 674 -77
rect 674 -133 678 -77
rect 614 -137 678 -133
rect 825 -77 889 -73
rect 825 -133 829 -77
rect 829 -133 885 -77
rect 885 -133 889 -77
rect 825 -137 889 -133
rect 1031 -77 1095 -73
rect 1031 -133 1035 -77
rect 1035 -133 1091 -77
rect 1091 -133 1095 -77
rect 1031 -137 1095 -133
rect 1259 -79 1323 -75
rect 1259 -135 1263 -79
rect 1263 -135 1319 -79
rect 1319 -135 1323 -79
rect 1259 -139 1323 -135
rect 1503 -79 1567 -75
rect 1503 -135 1507 -79
rect 1507 -135 1563 -79
rect 1563 -135 1567 -79
rect 1503 -139 1567 -135
rect 1733 -77 1797 -73
rect 1733 -133 1737 -77
rect 1737 -133 1793 -77
rect 1793 -133 1797 -77
rect 1733 -137 1797 -133
rect 1939 -77 2003 -73
rect 1939 -133 1943 -77
rect 1943 -133 1999 -77
rect 1999 -133 2003 -77
rect 1939 -137 2003 -133
rect 2157 -72 2221 -68
rect 2157 -128 2161 -72
rect 2161 -128 2217 -72
rect 2217 -128 2221 -72
rect 2157 -132 2221 -128
rect 2360 -78 2424 -74
rect 2360 -134 2364 -78
rect 2364 -134 2420 -78
rect 2420 -134 2424 -78
rect 2360 -138 2424 -134
rect 2568 -75 2632 -71
rect 2568 -131 2572 -75
rect 2572 -131 2628 -75
rect 2628 -131 2632 -75
rect 2568 -135 2632 -131
rect 2831 -79 2895 -75
rect 2831 -135 2835 -79
rect 2835 -135 2891 -79
rect 2891 -135 2895 -79
rect 2831 -139 2895 -135
rect 3039 -78 3103 -74
rect 3039 -134 3043 -78
rect 3043 -134 3099 -78
rect 3099 -134 3103 -78
rect 3039 -138 3103 -134
rect 3249 -81 3313 -77
rect 3249 -137 3253 -81
rect 3253 -137 3309 -81
rect 3309 -137 3313 -81
rect 3249 -141 3313 -137
rect 3449 -75 3513 -71
rect 3449 -131 3453 -75
rect 3453 -131 3509 -75
rect 3509 -131 3513 -75
rect 3449 -135 3513 -131
rect 3652 -78 3716 -74
rect 3652 -134 3656 -78
rect 3656 -134 3712 -78
rect 3712 -134 3716 -78
rect 3652 -138 3716 -134
rect 3862 -78 3926 -74
rect 3862 -134 3866 -78
rect 3866 -134 3922 -78
rect 3922 -134 3926 -78
rect 3862 -138 3926 -134
rect 4063 -77 4127 -73
rect 4063 -133 4067 -77
rect 4067 -133 4123 -77
rect 4123 -133 4127 -77
rect 4063 -137 4127 -133
rect 4279 -76 4343 -72
rect 4279 -132 4283 -76
rect 4283 -132 4339 -76
rect 4339 -132 4343 -76
rect 4279 -136 4343 -132
rect 4560 -78 4624 -74
rect 4560 -134 4564 -78
rect 4564 -134 4620 -78
rect 4620 -134 4624 -78
rect 4560 -138 4624 -134
rect 4780 -83 4844 -79
rect 4780 -139 4784 -83
rect 4784 -139 4840 -83
rect 4840 -139 4844 -83
rect 4780 -143 4844 -139
rect 4985 -82 5049 -78
rect 4985 -138 4989 -82
rect 4989 -138 5045 -82
rect 5045 -138 5049 -82
rect 4985 -142 5049 -138
rect 5206 -76 5270 -72
rect 5206 -132 5210 -76
rect 5210 -132 5266 -76
rect 5266 -132 5270 -76
rect 5206 -136 5270 -132
rect 5411 -83 5475 -79
rect 5411 -139 5415 -83
rect 5415 -139 5471 -83
rect 5471 -139 5475 -83
rect 5411 -143 5475 -139
rect 5620 -82 5684 -78
rect 5620 -138 5624 -82
rect 5624 -138 5680 -82
rect 5680 -138 5684 -82
rect 5620 -142 5684 -138
rect 5837 -82 5901 -78
rect 5837 -138 5841 -82
rect 5841 -138 5897 -82
rect 5897 -138 5901 -82
rect 5837 -142 5901 -138
rect 6051 -77 6115 -73
rect 6051 -133 6055 -77
rect 6055 -133 6111 -77
rect 6111 -133 6115 -77
rect 6051 -137 6115 -133
rect 6246 -79 6310 -75
rect 6246 -135 6250 -79
rect 6250 -135 6306 -79
rect 6306 -135 6310 -79
rect 6246 -139 6310 -135
rect 6441 -82 6505 -78
rect 6441 -138 6445 -82
rect 6445 -138 6501 -82
rect 6501 -138 6505 -82
rect 6441 -142 6505 -138
rect 6643 -79 6707 -75
rect 6643 -135 6647 -79
rect 6647 -135 6703 -79
rect 6703 -135 6707 -79
rect 6643 -139 6707 -135
rect 6927 -78 6991 -74
rect 6927 -134 6931 -78
rect 6931 -134 6987 -78
rect 6987 -134 6991 -78
rect 6927 -138 6991 -134
rect 7126 -77 7190 -73
rect 7126 -133 7130 -77
rect 7130 -133 7186 -77
rect 7186 -133 7190 -77
rect 7126 -137 7190 -133
rect 7329 -75 7393 -71
rect 7329 -131 7333 -75
rect 7333 -131 7389 -75
rect 7389 -131 7393 -75
rect 7329 -135 7393 -131
rect 7594 -78 7658 -74
rect 7594 -134 7598 -78
rect 7598 -134 7654 -78
rect 7654 -134 7658 -78
rect 7594 -138 7658 -134
rect 7792 -79 7856 -75
rect 7792 -135 7796 -79
rect 7796 -135 7852 -79
rect 7852 -135 7856 -79
rect 7792 -139 7856 -135
rect 7981 -77 8045 -73
rect 7981 -133 7985 -77
rect 7985 -133 8041 -77
rect 8041 -133 8045 -77
rect 7981 -137 8045 -133
rect 8193 -77 8257 -73
rect 8193 -133 8197 -77
rect 8197 -133 8253 -77
rect 8253 -133 8257 -77
rect 8193 -137 8257 -133
rect 8410 -77 8474 -73
rect 8410 -133 8414 -77
rect 8414 -133 8470 -77
rect 8470 -133 8474 -77
rect 8410 -137 8474 -133
rect 8615 -81 8679 -77
rect 8615 -137 8619 -81
rect 8619 -137 8675 -81
rect 8675 -137 8679 -81
rect 8615 -141 8679 -137
rect 8820 -81 8884 -77
rect 8820 -137 8824 -81
rect 8824 -137 8880 -81
rect 8880 -137 8884 -81
rect 8820 -141 8884 -137
rect 9028 -76 9092 -72
rect 9028 -132 9032 -76
rect 9032 -132 9088 -76
rect 9088 -132 9092 -76
rect 9028 -136 9092 -132
rect 9311 -77 9375 -73
rect 9311 -133 9315 -77
rect 9315 -133 9371 -77
rect 9371 -133 9375 -77
rect 9311 -137 9375 -133
rect 9504 -79 9568 -75
rect 9504 -135 9508 -79
rect 9508 -135 9564 -79
rect 9564 -135 9568 -79
rect 9504 -139 9568 -135
rect 9730 -81 9794 -77
rect 9730 -137 9734 -81
rect 9734 -137 9790 -81
rect 9790 -137 9794 -81
rect 9730 -141 9794 -137
rect 9995 -81 10059 -77
rect 9995 -137 9999 -81
rect 9999 -137 10055 -81
rect 10055 -137 10059 -81
rect 9995 -141 10059 -137
rect 10189 -77 10253 -73
rect 10189 -133 10193 -77
rect 10193 -133 10249 -77
rect 10249 -133 10253 -77
rect 10189 -137 10253 -133
rect 10387 -86 10451 -82
rect 10387 -142 10391 -86
rect 10391 -142 10447 -86
rect 10447 -142 10451 -86
rect 10387 -146 10451 -142
rect 10591 -78 10655 -74
rect 10591 -134 10595 -78
rect 10595 -134 10651 -78
rect 10651 -134 10655 -78
rect 10591 -138 10655 -134
rect 10811 -75 10875 -71
rect 10811 -131 10815 -75
rect 10815 -131 10871 -75
rect 10871 -131 10875 -75
rect 10811 -135 10875 -131
rect 11026 -79 11090 -75
rect 11026 -135 11030 -79
rect 11030 -135 11086 -79
rect 11086 -135 11090 -79
rect 11026 -139 11090 -135
rect 11254 -76 11318 -72
rect 11254 -132 11258 -76
rect 11258 -132 11314 -76
rect 11314 -132 11318 -76
rect 11254 -136 11318 -132
rect 11458 -79 11522 -75
rect 11458 -135 11462 -79
rect 11462 -135 11518 -79
rect 11518 -135 11522 -79
rect 11458 -139 11522 -135
rect 11696 -77 11760 -73
rect 11696 -133 11700 -77
rect 11700 -133 11756 -77
rect 11756 -133 11760 -77
rect 11696 -137 11760 -133
rect 11889 -76 11953 -72
rect 11889 -132 11893 -76
rect 11893 -132 11949 -76
rect 11949 -132 11953 -76
rect 11889 -136 11953 -132
rect 12086 -81 12150 -77
rect 12086 -137 12090 -81
rect 12090 -137 12146 -81
rect 12146 -137 12150 -81
rect 12086 -141 12150 -137
rect 12342 -78 12406 -74
rect 12342 -134 12346 -78
rect 12346 -134 12402 -78
rect 12402 -134 12406 -78
rect 12342 -138 12406 -134
rect 12581 -82 12645 -78
rect 12581 -138 12585 -82
rect 12585 -138 12641 -82
rect 12641 -138 12645 -82
rect 12581 -142 12645 -138
rect 12814 -86 12878 -82
rect 12814 -142 12818 -86
rect 12818 -142 12874 -86
rect 12874 -142 12878 -86
rect 12814 -146 12878 -142
rect 13035 -81 13099 -77
rect 13035 -137 13039 -81
rect 13039 -137 13095 -81
rect 13095 -137 13099 -81
rect 13035 -141 13099 -137
rect 13226 -81 13290 -77
rect 13226 -137 13230 -81
rect 13230 -137 13286 -81
rect 13286 -137 13290 -81
rect 13226 -141 13290 -137
rect 13454 -79 13518 -75
rect 13454 -135 13458 -79
rect 13458 -135 13514 -79
rect 13514 -135 13518 -79
rect 13454 -139 13518 -135
rect 13651 -84 13715 -80
rect 13651 -140 13655 -84
rect 13655 -140 13711 -84
rect 13711 -140 13715 -84
rect 13651 -144 13715 -140
rect 13863 -84 13927 -80
rect 13863 -140 13867 -84
rect 13867 -140 13923 -84
rect 13923 -140 13927 -84
rect 13863 -144 13927 -140
rect 14090 -81 14154 -77
rect 14090 -137 14094 -81
rect 14094 -137 14150 -81
rect 14150 -137 14154 -81
rect 14090 -141 14154 -137
rect 14279 -80 14343 -76
rect 14279 -136 14283 -80
rect 14283 -136 14339 -80
rect 14339 -136 14343 -80
rect 14279 -140 14343 -136
rect 14505 -79 14569 -75
rect 14505 -135 14509 -79
rect 14509 -135 14565 -79
rect 14565 -135 14569 -79
rect 14505 -139 14569 -135
rect 14759 -79 14823 -75
rect 14759 -135 14763 -79
rect 14763 -135 14819 -79
rect 14819 -135 14823 -79
rect 14759 -139 14823 -135
rect 15003 -82 15067 -78
rect 15003 -138 15007 -82
rect 15007 -138 15063 -82
rect 15063 -138 15067 -82
rect 15003 -142 15067 -138
rect 15233 -83 15297 -79
rect 15233 -139 15237 -83
rect 15237 -139 15293 -83
rect 15293 -139 15297 -83
rect 15233 -143 15297 -139
rect 15491 -80 15555 -76
rect 15491 -136 15495 -80
rect 15495 -136 15551 -80
rect 15551 -136 15555 -80
rect 15491 -140 15555 -136
rect 15701 -80 15765 -76
rect 15701 -136 15705 -80
rect 15705 -136 15761 -80
rect 15761 -136 15765 -80
rect 15701 -140 15765 -136
rect 15926 -80 15990 -76
rect 15926 -136 15930 -80
rect 15930 -136 15986 -80
rect 15986 -136 15990 -80
rect 15926 -140 15990 -136
rect 16145 -83 16209 -79
rect 16145 -139 16149 -83
rect 16149 -139 16205 -83
rect 16205 -139 16209 -83
rect 16145 -143 16209 -139
rect 16491 -79 16555 -75
rect 16491 -135 16495 -79
rect 16495 -135 16551 -79
rect 16551 -135 16555 -79
rect 16491 -139 16555 -135
rect 16690 -82 16754 -78
rect 16690 -138 16694 -82
rect 16694 -138 16750 -82
rect 16750 -138 16754 -82
rect 16690 -142 16754 -138
<< metal4 >>
rect 686 3441 815 3452
rect 686 3377 717 3441
rect 781 3377 815 3441
rect 686 3366 815 3377
rect -144 2986 16604 3041
rect -144 2984 1259 2986
rect -144 2982 249 2984
rect -144 2918 47 2982
rect 111 2920 249 2982
rect 313 2982 858 2984
rect 313 2920 460 2982
rect 111 2918 460 2920
rect 524 2918 650 2982
rect 714 2920 858 2982
rect 922 2920 1060 2984
rect 1124 2922 1259 2984
rect 1323 2985 2146 2986
rect 1323 2983 1655 2985
rect 1323 2922 1454 2983
rect 1124 2920 1454 2922
rect 714 2919 1454 2920
rect 1518 2921 1655 2983
rect 1719 2983 2146 2985
rect 1719 2921 1872 2983
rect 1518 2919 1872 2921
rect 1936 2922 2146 2983
rect 2210 2982 16604 2986
rect 2210 2979 2646 2982
rect 2210 2922 2423 2979
rect 1936 2919 2423 2922
rect 714 2918 2423 2919
rect -144 2915 2423 2918
rect 2487 2918 2646 2979
rect 2710 2981 16604 2982
rect 2710 2918 2878 2981
rect 2487 2917 2878 2918
rect 2942 2980 5897 2981
rect 2942 2979 5022 2980
rect 2942 2978 4822 2979
rect 2942 2917 4514 2978
rect 2487 2915 4514 2917
rect -144 2914 4514 2915
rect 4578 2915 4822 2978
rect 4886 2916 5022 2979
rect 5086 2979 5695 2980
rect 5086 2916 5241 2979
rect 4886 2915 5241 2916
rect 5305 2978 5695 2979
rect 5305 2915 5487 2978
rect 4578 2914 5487 2915
rect 5551 2916 5695 2978
rect 5759 2917 5897 2980
rect 5961 2980 16604 2981
rect 5961 2917 6090 2980
rect 5759 2916 6090 2917
rect 6154 2979 16604 2980
rect 6154 2916 6462 2979
rect 5551 2915 6462 2916
rect 6526 2977 7214 2979
rect 6526 2915 6651 2977
rect 5551 2914 6651 2915
rect -144 2913 6651 2914
rect 6715 2913 6941 2977
rect 7005 2915 7214 2977
rect 7278 2915 16604 2979
rect 7005 2913 16604 2915
rect -144 2721 16604 2913
rect -144 1838 1030 2721
rect -144 1774 13 1838
rect 77 1836 1030 1838
rect 77 1774 253 1836
rect -144 1772 253 1774
rect 317 1835 793 1836
rect 317 1772 575 1835
rect -144 1771 575 1772
rect 639 1772 793 1835
rect 857 1772 1030 1836
rect 639 1771 1030 1772
rect -144 1155 1030 1771
rect -144 1091 259 1155
rect 323 1151 1030 1155
rect 323 1091 461 1151
rect -144 1087 461 1091
rect 525 1149 1030 1151
rect 525 1148 879 1149
rect 525 1087 650 1148
rect -144 1084 650 1087
rect 714 1085 879 1148
rect 943 1085 1030 1149
rect 714 1084 1030 1085
rect -144 465 1030 1084
rect -144 462 489 465
rect -144 398 41 462
rect 105 458 489 462
rect 105 398 274 458
rect -144 394 274 398
rect 338 401 489 458
rect 553 463 1030 465
rect 553 462 923 463
rect 553 401 707 462
rect 338 398 707 401
rect 771 399 923 462
rect 987 399 1030 463
rect 771 398 1030 399
rect 338 394 1030 398
rect -144 195 1030 394
rect 1110 2447 2496 2640
rect 1110 2443 1384 2447
rect 1110 2379 1165 2443
rect 1229 2383 1384 2443
rect 1448 2383 1667 2447
rect 1731 2383 1876 2447
rect 1940 2445 2496 2447
rect 1940 2383 2147 2445
rect 1229 2381 2147 2383
rect 2211 2381 2496 2445
rect 1229 2379 2496 2381
rect 1110 1300 2496 2379
rect 1110 1236 1204 1300
rect 1268 1236 1421 1300
rect 1485 1236 1640 1300
rect 1704 1296 2496 1300
rect 1704 1236 1853 1296
rect 1110 1232 1853 1236
rect 1917 1232 2064 1296
rect 2128 1232 2496 1296
rect 1110 618 2496 1232
rect 1110 606 1415 618
rect 1110 542 1186 606
rect 1250 554 1415 606
rect 1479 612 2496 618
rect 1479 608 1826 612
rect 1479 554 1634 608
rect 1250 544 1634 554
rect 1698 548 1826 608
rect 1890 610 2496 612
rect 1890 548 2320 610
rect 1698 546 2320 548
rect 2384 546 2496 610
rect 1698 544 2496 546
rect 1250 542 2496 544
rect 1110 114 2496 542
rect 2576 1842 3962 2721
rect 2576 1840 3022 1842
rect 2576 1776 2697 1840
rect 2761 1778 3022 1840
rect 3086 1778 3290 1842
rect 3354 1778 3556 1842
rect 3620 1840 3962 1842
rect 3620 1778 3796 1840
rect 2761 1776 3796 1778
rect 3860 1776 3962 1840
rect 2576 1156 3962 1776
rect 2576 1152 3256 1156
rect 2576 1088 2648 1152
rect 2712 1149 3256 1152
rect 2712 1088 2863 1149
rect 2576 1085 2863 1088
rect 2927 1146 3256 1149
rect 2927 1085 3061 1146
rect 2576 1082 3061 1085
rect 3125 1092 3256 1146
rect 3320 1154 3962 1156
rect 3320 1092 3536 1154
rect 3125 1090 3536 1092
rect 3600 1152 3962 1154
rect 3600 1090 3755 1152
rect 3125 1088 3755 1090
rect 3819 1088 3962 1152
rect 3125 1082 3962 1088
rect 2576 467 3962 1082
rect 2576 462 3780 467
rect 2576 459 3044 462
rect 2576 395 2644 459
rect 2708 395 2834 459
rect 2898 398 3044 459
rect 3108 459 3556 462
rect 3108 398 3261 459
rect 2898 395 3261 398
rect 3325 398 3556 459
rect 3620 403 3780 462
rect 3844 403 3962 467
rect 3620 398 3962 403
rect 3325 395 3962 398
rect 2576 195 3962 395
rect 4042 2446 5428 2640
rect 4042 2443 4471 2446
rect 4042 2379 4222 2443
rect 4286 2382 4471 2443
rect 4535 2438 5428 2446
rect 4535 2432 5069 2438
rect 4535 2382 4815 2432
rect 4286 2379 4815 2382
rect 4042 2368 4815 2379
rect 4879 2374 5069 2432
rect 5133 2374 5298 2438
rect 5362 2374 5428 2438
rect 4879 2368 5428 2374
rect 4042 1300 5428 2368
rect 4042 1296 5038 1300
rect 4042 1232 4188 1296
rect 4252 1295 5038 1296
rect 4252 1232 4466 1295
rect 4042 1231 4466 1232
rect 4530 1236 5038 1295
rect 5102 1236 5277 1300
rect 5341 1236 5428 1300
rect 4530 1231 5428 1236
rect 4042 617 5428 1231
rect 4042 615 5032 617
rect 4042 609 4702 615
rect 4042 545 4112 609
rect 4176 607 4702 609
rect 4176 545 4505 607
rect 4042 543 4505 545
rect 4569 551 4702 607
rect 4766 553 5032 615
rect 5096 553 5228 617
rect 5292 553 5428 617
rect 4766 551 5428 553
rect 4569 543 5428 551
rect 4042 114 5428 543
rect 5508 1846 6894 2721
rect 5508 1843 5956 1846
rect 5508 1779 5590 1843
rect 5654 1782 5956 1843
rect 6020 1782 6200 1846
rect 6264 1837 6894 1846
rect 6264 1782 6623 1837
rect 5654 1779 6623 1782
rect 5508 1773 6623 1779
rect 6687 1773 6894 1837
rect 5508 1153 6894 1773
rect 5508 1151 6512 1153
rect 5508 1149 6321 1151
rect 5508 1085 5576 1149
rect 5640 1146 6321 1149
rect 5640 1085 5927 1146
rect 5508 1082 5927 1085
rect 5991 1144 6321 1146
rect 5991 1082 6116 1144
rect 5508 1080 6116 1082
rect 6180 1087 6321 1144
rect 6385 1089 6512 1151
rect 6576 1089 6894 1153
rect 6385 1087 6894 1089
rect 6180 1080 6894 1087
rect 5508 467 6894 1080
rect 5508 462 6427 467
rect 5508 460 6210 462
rect 5508 396 5658 460
rect 5722 458 6210 460
rect 5722 396 5958 458
rect 5508 394 5958 396
rect 6022 398 6210 458
rect 6274 403 6427 462
rect 6491 464 6894 467
rect 6491 403 6628 464
rect 6274 400 6628 403
rect 6692 400 6894 464
rect 6274 398 6894 400
rect 6022 394 6894 398
rect 5508 194 6894 394
rect 6974 2445 8360 2640
rect 6974 2443 7220 2445
rect 6974 2379 7016 2443
rect 7080 2381 7220 2443
rect 7284 2443 8360 2445
rect 7284 2381 7543 2443
rect 7080 2379 7543 2381
rect 7607 2379 8360 2443
rect 6974 1305 8360 2379
rect 6974 1303 7852 1305
rect 6974 1298 7662 1303
rect 6974 1234 7435 1298
rect 7499 1239 7662 1298
rect 7726 1241 7852 1303
rect 7916 1296 8360 1305
rect 7916 1241 8068 1296
rect 7726 1239 8068 1241
rect 7499 1234 8068 1239
rect 6974 1232 8068 1234
rect 8132 1232 8360 1296
rect 6974 617 8360 1232
rect 6974 615 8063 617
rect 6974 614 7642 615
rect 6974 610 7436 614
rect 6974 546 7135 610
rect 7199 550 7436 610
rect 7500 551 7642 614
rect 7706 611 8063 615
rect 7706 551 7852 611
rect 7500 550 7852 551
rect 7199 547 7852 550
rect 7916 553 8063 611
rect 8127 553 8360 617
rect 7916 547 8360 553
rect 7199 546 8360 547
rect 6974 114 8360 546
rect 8440 1844 9826 2721
rect 8440 1839 9024 1844
rect 8440 1775 8566 1839
rect 8630 1836 9024 1839
rect 8630 1775 8818 1836
rect 8440 1772 8818 1775
rect 8882 1780 9024 1836
rect 9088 1839 9826 1844
rect 9088 1838 9605 1839
rect 9088 1780 9307 1838
rect 8882 1774 9307 1780
rect 9371 1775 9605 1838
rect 9669 1775 9826 1839
rect 9371 1774 9826 1775
rect 8882 1772 9826 1774
rect 8440 1157 9826 1772
rect 8440 1155 8747 1157
rect 8440 1091 8557 1155
rect 8621 1093 8747 1155
rect 8811 1155 9826 1157
rect 8811 1093 8941 1155
rect 8621 1091 8941 1093
rect 9005 1151 9826 1155
rect 9005 1091 9252 1151
rect 8440 1087 9252 1091
rect 9316 1087 9826 1151
rect 8440 463 9826 1087
rect 8440 455 9523 463
rect 8440 391 8513 455
rect 8577 391 8705 455
rect 8769 391 8905 455
rect 8969 399 9523 455
rect 9587 399 9826 463
rect 8969 391 9826 399
rect 8440 195 9826 391
rect 9906 1307 11292 2641
rect 9906 1302 10504 1307
rect 9906 1299 10278 1302
rect 9906 1235 10049 1299
rect 10113 1238 10278 1299
rect 10342 1243 10504 1302
rect 10568 1305 11292 1307
rect 10568 1299 10968 1305
rect 10568 1243 10732 1299
rect 10342 1238 10732 1243
rect 10113 1235 10732 1238
rect 10796 1241 10968 1299
rect 11032 1296 11292 1305
rect 11032 1241 11160 1296
rect 10796 1235 11160 1241
rect 9906 1232 11160 1235
rect 11224 1232 11292 1296
rect 9906 617 11292 1232
rect 9906 614 10962 617
rect 9906 613 10721 614
rect 9906 606 10200 613
rect 9906 542 9943 606
rect 10007 549 10200 606
rect 10264 609 10721 613
rect 10264 549 10450 609
rect 10007 545 10450 549
rect 10514 550 10721 609
rect 10785 553 10962 614
rect 11026 613 11292 617
rect 11026 553 11187 613
rect 10785 550 11187 553
rect 10514 549 11187 550
rect 11251 549 11292 613
rect 10514 545 11292 549
rect 10007 542 11292 545
rect 9906 114 11292 542
rect 11372 1842 12758 2721
rect 11372 1840 11647 1842
rect 11372 1776 11437 1840
rect 11501 1778 11647 1840
rect 11711 1840 12758 1842
rect 11711 1778 11998 1840
rect 11501 1776 11998 1778
rect 12062 1776 12278 1840
rect 12342 1839 12758 1840
rect 12342 1776 12595 1839
rect 11372 1775 12595 1776
rect 12659 1775 12758 1839
rect 11372 1150 12758 1775
rect 11372 1086 11435 1150
rect 11499 1086 11639 1150
rect 11703 1148 12758 1150
rect 11703 1146 12443 1148
rect 11703 1086 12204 1146
rect 11372 1082 12204 1086
rect 12268 1084 12443 1146
rect 12507 1084 12647 1148
rect 12711 1084 12758 1148
rect 12268 1082 12758 1084
rect 11372 461 12758 1082
rect 11372 459 12204 461
rect 11372 395 11424 459
rect 11488 395 11680 459
rect 11744 395 11915 459
rect 11979 397 12204 459
rect 12268 459 12598 461
rect 12268 397 12394 459
rect 11979 395 12394 397
rect 12458 397 12598 459
rect 12662 397 12758 461
rect 12458 395 12758 397
rect 11372 195 12758 395
rect 12838 1301 14224 2640
rect 12838 1296 13099 1301
rect 12838 1232 12895 1296
rect 12959 1237 13099 1296
rect 13163 1296 14224 1301
rect 13163 1237 13290 1296
rect 12959 1232 13290 1237
rect 13354 1295 13782 1296
rect 13354 1232 13492 1295
rect 12838 1231 13492 1232
rect 13556 1232 13782 1295
rect 13846 1295 14224 1296
rect 13846 1232 14067 1295
rect 13556 1231 14067 1232
rect 14131 1231 14224 1295
rect 12838 612 14224 1231
rect 12838 611 13095 612
rect 12838 547 12894 611
rect 12958 548 13095 611
rect 13159 608 13520 612
rect 13159 548 13313 608
rect 12958 547 13313 548
rect 12838 544 13313 547
rect 13377 548 13520 608
rect 13584 611 14224 612
rect 13584 548 13725 611
rect 13377 547 13725 548
rect 13789 607 14224 611
rect 13789 547 14072 607
rect 13377 544 14072 547
rect 12838 543 14072 544
rect 14136 543 14224 607
rect 12838 114 14224 543
rect 14304 1840 15690 2721
rect 14304 1837 15541 1840
rect 14304 1773 14385 1837
rect 14449 1773 14680 1837
rect 14744 1773 14967 1837
rect 15031 1773 15257 1837
rect 15321 1776 15541 1837
rect 15605 1776 15690 1840
rect 15321 1773 15690 1776
rect 14304 1156 15690 1773
rect 14304 1092 14607 1156
rect 14671 1154 15536 1156
rect 14671 1092 14840 1154
rect 14304 1090 14840 1092
rect 14904 1152 15256 1154
rect 14904 1090 15047 1152
rect 14304 1088 15047 1090
rect 15111 1090 15256 1152
rect 15320 1092 15536 1154
rect 15600 1092 15690 1156
rect 15320 1090 15690 1092
rect 15111 1088 15690 1090
rect 14304 470 15690 1088
rect 14304 467 15016 470
rect 14304 403 14384 467
rect 14448 463 15016 467
rect 14448 403 14626 463
rect 14304 399 14626 403
rect 14690 462 15016 463
rect 14690 399 14826 462
rect 14304 398 14826 399
rect 14890 406 15016 462
rect 15080 468 15690 470
rect 15080 406 15237 468
rect 14890 404 15237 406
rect 15301 463 15690 468
rect 15301 404 15533 463
rect 14890 399 15533 404
rect 15597 399 15690 463
rect 14890 398 15690 399
rect 14304 195 15690 398
rect 15770 1304 16876 2640
rect 15770 1300 16016 1304
rect 15770 1236 15822 1300
rect 15886 1240 16016 1300
rect 16080 1303 16876 1304
rect 16080 1301 16428 1303
rect 16080 1240 16205 1301
rect 15886 1237 16205 1240
rect 16269 1239 16428 1301
rect 16492 1239 16876 1303
rect 16269 1237 16876 1239
rect 15886 1236 16876 1237
rect 15770 616 16876 1236
rect 15770 614 16210 616
rect 15770 611 16015 614
rect 15770 547 15824 611
rect 15888 550 16015 611
rect 16079 552 16210 614
rect 16274 611 16876 616
rect 16274 552 16657 611
rect 16079 550 16657 552
rect 15888 547 16657 550
rect 16721 547 16876 611
rect 15770 114 16876 547
rect 196 -68 16876 114
rect 196 -70 2157 -68
rect 196 -134 415 -70
rect 479 -73 2157 -70
rect 479 -134 614 -73
rect 196 -137 614 -134
rect 678 -137 825 -73
rect 889 -137 1031 -73
rect 1095 -75 1733 -73
rect 1095 -137 1259 -75
rect 196 -139 1259 -137
rect 1323 -139 1503 -75
rect 1567 -137 1733 -75
rect 1797 -137 1939 -73
rect 2003 -132 2157 -73
rect 2221 -71 16876 -68
rect 2221 -74 2568 -71
rect 2221 -132 2360 -74
rect 2003 -137 2360 -132
rect 1567 -138 2360 -137
rect 2424 -135 2568 -74
rect 2632 -74 3449 -71
rect 2632 -75 3039 -74
rect 2632 -135 2831 -75
rect 2424 -138 2831 -135
rect 1567 -139 2831 -138
rect 2895 -138 3039 -75
rect 3103 -77 3449 -74
rect 3103 -138 3249 -77
rect 2895 -139 3249 -138
rect 196 -141 3249 -139
rect 3313 -135 3449 -77
rect 3513 -72 7329 -71
rect 3513 -73 4279 -72
rect 3513 -74 4063 -73
rect 3513 -135 3652 -74
rect 3313 -138 3652 -135
rect 3716 -138 3862 -74
rect 3926 -137 4063 -74
rect 4127 -136 4279 -73
rect 4343 -74 5206 -72
rect 4343 -136 4560 -74
rect 4127 -137 4560 -136
rect 3926 -138 4560 -137
rect 4624 -78 5206 -74
rect 4624 -79 4985 -78
rect 4624 -138 4780 -79
rect 3313 -141 4780 -138
rect 196 -143 4780 -141
rect 4844 -142 4985 -79
rect 5049 -136 5206 -78
rect 5270 -73 7329 -72
rect 5270 -78 6051 -73
rect 5270 -79 5620 -78
rect 5270 -136 5411 -79
rect 5049 -142 5411 -136
rect 4844 -143 5411 -142
rect 5475 -142 5620 -79
rect 5684 -142 5837 -78
rect 5901 -137 6051 -78
rect 6115 -74 7126 -73
rect 6115 -75 6927 -74
rect 6115 -137 6246 -75
rect 5901 -139 6246 -137
rect 6310 -78 6643 -75
rect 6310 -139 6441 -78
rect 5901 -142 6441 -139
rect 6505 -139 6643 -78
rect 6707 -138 6927 -75
rect 6991 -137 7126 -74
rect 7190 -135 7329 -73
rect 7393 -72 10811 -71
rect 7393 -73 9028 -72
rect 7393 -74 7981 -73
rect 7393 -135 7594 -74
rect 7190 -137 7594 -135
rect 6991 -138 7594 -137
rect 7658 -75 7981 -74
rect 7658 -138 7792 -75
rect 6707 -139 7792 -138
rect 7856 -137 7981 -75
rect 8045 -137 8193 -73
rect 8257 -137 8410 -73
rect 8474 -77 9028 -73
rect 8474 -137 8615 -77
rect 7856 -139 8615 -137
rect 6505 -141 8615 -139
rect 8679 -141 8820 -77
rect 8884 -136 9028 -77
rect 9092 -73 10811 -72
rect 9092 -136 9311 -73
rect 8884 -137 9311 -136
rect 9375 -75 10189 -73
rect 9375 -137 9504 -75
rect 8884 -139 9504 -137
rect 9568 -77 10189 -75
rect 9568 -139 9730 -77
rect 8884 -141 9730 -139
rect 9794 -141 9995 -77
rect 10059 -137 10189 -77
rect 10253 -74 10811 -73
rect 10253 -82 10591 -74
rect 10253 -137 10387 -82
rect 10059 -141 10387 -137
rect 6505 -142 10387 -141
rect 5475 -143 10387 -142
rect 196 -146 10387 -143
rect 10451 -138 10591 -82
rect 10655 -135 10811 -74
rect 10875 -72 16876 -71
rect 10875 -75 11254 -72
rect 10875 -135 11026 -75
rect 10655 -138 11026 -135
rect 10451 -139 11026 -138
rect 11090 -136 11254 -75
rect 11318 -73 11889 -72
rect 11318 -75 11696 -73
rect 11318 -136 11458 -75
rect 11090 -139 11458 -136
rect 11522 -137 11696 -75
rect 11760 -136 11889 -73
rect 11953 -74 16876 -72
rect 11953 -77 12342 -74
rect 11953 -136 12086 -77
rect 11760 -137 12086 -136
rect 11522 -139 12086 -137
rect 10451 -141 12086 -139
rect 12150 -138 12342 -77
rect 12406 -75 16876 -74
rect 12406 -77 13454 -75
rect 12406 -78 13035 -77
rect 12406 -138 12581 -78
rect 12150 -141 12581 -138
rect 10451 -142 12581 -141
rect 12645 -82 13035 -78
rect 12645 -142 12814 -82
rect 10451 -146 12814 -142
rect 12878 -141 13035 -82
rect 13099 -141 13226 -77
rect 13290 -139 13454 -77
rect 13518 -76 14505 -75
rect 13518 -77 14279 -76
rect 13518 -80 14090 -77
rect 13518 -139 13651 -80
rect 13290 -141 13651 -139
rect 12878 -144 13651 -141
rect 13715 -144 13863 -80
rect 13927 -141 14090 -80
rect 14154 -140 14279 -77
rect 14343 -139 14505 -76
rect 14569 -139 14759 -75
rect 14823 -76 16491 -75
rect 14823 -78 15491 -76
rect 14823 -139 15003 -78
rect 14343 -140 15003 -139
rect 14154 -141 15003 -140
rect 13927 -142 15003 -141
rect 15067 -79 15491 -78
rect 15067 -142 15233 -79
rect 13927 -143 15233 -142
rect 15297 -140 15491 -79
rect 15555 -140 15701 -76
rect 15765 -140 15926 -76
rect 15990 -79 16491 -76
rect 15990 -140 16145 -79
rect 15297 -143 16145 -140
rect 16209 -139 16491 -79
rect 16555 -78 16876 -75
rect 16555 -139 16690 -78
rect 16209 -142 16690 -139
rect 16754 -142 16876 -78
rect 16209 -143 16876 -142
rect 13927 -144 16876 -143
rect 12878 -146 16876 -144
rect 196 -206 16876 -146
use sky130_fd_sc_hd__dfbbn_1  sky130_fd_sc_hd__dfbbn_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1699356299
transform 1 0 0 0 1 580
box -38 -48 2430 592
use sky130_fd_sc_hd__buf_1  x1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698323353
transform 1 0 2 0 1 2410
box -38 -48 314 592
use sky130_fd_sc_hd__buf_16  x2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698323353
transform 1 0 830 0 1 2410
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_4  x3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698323353
transform 1 0 278 0 1 2410
box -38 -48 590 592
use sky130_fd_sc_hd__dfbbn_1  x5
timestamp 1699356299
transform -1 0 2392 0 1 -109
box -38 -48 2430 592
use sky130_fd_sc_hd__mux2_1  x6 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 0 0 1 1268
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  x7
timestamp 1683767628
transform -1 0 2262 0 1 1268
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  x8
timestamp 1683767628
transform 1 0 2392 0 1 1268
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  x9
timestamp 1683767628
transform -1 0 4654 0 1 1268
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  x10
timestamp 1683767628
transform 1 0 4784 0 1 1268
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  x11
timestamp 1683767628
transform -1 0 7044 0 1 1268
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  x12
timestamp 1683767628
transform 1 0 7176 0 1 1268
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  x13
timestamp 1683767628
transform -1 0 9438 0 1 1268
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  x14
timestamp 1683767628
transform 1 0 9568 0 1 1268
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  x15
timestamp 1683767628
transform -1 0 11830 0 1 1268
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  x16
timestamp 1683767628
transform 1 0 11960 0 1 1268
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  x17
timestamp 1683767628
transform -1 0 14220 0 1 1268
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  x18
timestamp 1683767628
transform 1 0 14352 0 1 1268
box -38 -48 866 592
use sky130_fd_sc_hd__dfbbn_1  x19
timestamp 1699356299
transform 1 0 2392 0 1 580
box -38 -48 2430 592
use sky130_fd_sc_hd__mux2_1  x20
timestamp 1683767628
transform -1 0 16614 0 1 1268
box -38 -48 866 592
use sky130_fd_sc_hd__dfbbn_1  x21
timestamp 1699356299
transform -1 0 4784 0 1 -109
box -38 -48 2430 592
use sky130_fd_sc_hd__buf_1  x22
timestamp 1698323353
transform 1 0 4386 0 1 2410
box -38 -48 314 592
use sky130_fd_sc_hd__dfbbn_1  x23
timestamp 1699356299
transform 1 0 4784 0 1 580
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbn_1  x24
timestamp 1699356299
transform -1 0 7176 0 1 -109
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbn_1  x25
timestamp 1699356299
transform 1 0 7176 0 1 580
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbn_1  x26
timestamp 1699356299
transform -1 0 9568 0 1 -109
box -38 -48 2430 592
use sky130_fd_sc_hd__buf_4  x27
timestamp 1698323353
transform 1 0 4662 0 1 2410
box -38 -48 590 592
use sky130_fd_sc_hd__dfbbn_1  x28
timestamp 1699356299
transform 1 0 9568 0 1 580
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbn_1  x29
timestamp 1699356299
transform -1 0 11960 0 1 -109
box -38 -48 2430 592
use sky130_fd_sc_hd__buf_16  x30
timestamp 1698323353
transform 1 0 5214 0 1 2410
box -38 -48 2062 592
use sky130_fd_sc_hd__dfbbn_1  x31
timestamp 1699356299
transform 1 0 11960 0 1 580
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbn_1  x32
timestamp 1699356299
transform -1 0 14352 0 1 -109
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbn_1  x34
timestamp 1699356299
transform 1 0 14352 0 1 580
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbn_1  x35
timestamp 1699356299
transform -1 0 16744 0 1 -109
box -38 -48 2430 592
<< labels >>
flabel metal2 9709 344 9751 3300 0 FreeSans 320 0 0 0 VSS_SW[3]
port 6 nsew
flabel metal2 7317 345 7359 3300 0 FreeSans 320 0 0 0 VSS_SW[4]
port 7 nsew
flabel metal2 4926 345 4968 3300 0 FreeSans 320 0 0 0 VSS_SW[5]
port 8 nsew
flabel metal2 14290 1062 14332 3300 0 FreeSans 320 0 0 0 VDD_SW[2]
port 11 nsew
flabel metal2 11898 1062 11940 3300 0 FreeSans 320 0 0 0 VDD_SW[3]
port 12 nsew
flabel metal2 9506 1062 9548 3300 0 FreeSans 320 0 0 0 VDD_SW[4]
port 13 nsew
flabel metal2 7114 1062 7156 3300 0 FreeSans 320 0 0 0 VDD_SW[5]
port 14 nsew
flabel metal2 4722 1062 4764 3300 0 FreeSans 320 0 0 0 VDD_SW[6]
port 15 nsew
flabel metal2 13924 1454 13966 3300 0 FreeSans 320 0 0 0 D[2]
port 17 nsew
flabel metal2 11531 1454 11573 3300 0 FreeSans 320 0 0 0 D[3]
port 18 nsew
flabel metal2 9140 1453 9182 3300 0 FreeSans 320 0 0 0 D[4]
port 19 nsew
flabel metal2 6747 1454 6789 3300 0 FreeSans 320 0 0 0 D[5]
port 20 nsew
flabel metal2 4356 1453 4398 3300 0 FreeSans 320 0 0 0 D[6]
port 21 nsew
flabel metal2 15914 1603 15956 3300 0 FreeSans 320 0 0 0 check[0]
port 23 nsew
flabel metal2 13519 1602 13561 3300 0 FreeSans 320 0 0 0 check[1]
port 24 nsew
flabel metal2 11130 1602 11172 3300 0 FreeSans 320 0 0 0 check[2]
port 25 nsew
flabel metal2 8738 1603 8780 3300 0 FreeSans 320 0 0 0 check[3]
port 26 nsew
flabel metal2 6344 1602 6386 3300 0 FreeSans 320 0 0 0 check[4]
port 27 nsew
flabel metal2 3954 1602 3996 3300 0 FreeSans 320 0 0 0 check[5]
port 28 nsew
flabel metal2 16317 1454 16359 3300 0 FreeSans 320 0 0 0 D[1]
port 46 nsew
flabel metal2 16682 1062 16724 3300 0 FreeSans 320 0 0 0 VDD_SW[1]
port 49 nsew
flabel metal2 1562 1603 1604 3300 0 FreeSans 320 0 0 0 check[6]
port 29 nsew
flabel metal2 1964 1453 2006 3300 0 FreeSans 320 0 0 0 D[7]
port 22 nsew
flabel metal2 2330 1062 2372 3300 0 FreeSans 320 0 0 0 VDD_SW[7]
port 16 nsew
flabel metal2 2533 345 2575 3300 0 FreeSans 320 0 0 0 VSS_SW[6]
port 9 nsew
flabel metal2 141 345 183 3300 0 FreeSans 320 0 0 0 VSS_SW[7]
port 10 nsew
rlabel comment s 4386 2410 4386 2410 4 buf_1
rlabel comment s 5214 2410 5214 2410 4 buf_16
rlabel comment s 4662 2410 4662 2410 4 buf_4
rlabel comment s 276 1268 276 1268 4 buf_4
rlabel comment s 828 1268 828 1268 4 buf_16
rlabel comment s 0 1268 0 1268 4 buf_1
rlabel comment s 3128 1268 3128 1268 4 buf_4
rlabel comment s 3680 1268 3680 1268 4 buf_16
rlabel comment s 2852 1268 2852 1268 4 buf_1
rlabel comment s 6216 1268 6216 1268 4 buf_1
rlabel comment s 7044 1268 7044 1268 4 buf_16
rlabel comment s 6492 1268 6492 1268 4 buf_4
rlabel comment s 9068 1268 9068 1268 4 buf_1
rlabel comment s 9896 1268 9896 1268 4 buf_16
rlabel comment s 9344 1268 9344 1268 4 buf_4
rlabel comment s 11982 1268 11982 1268 4 buf_1
rlabel comment s 12810 1268 12810 1268 4 buf_16
rlabel comment s 12258 1268 12258 1268 4 buf_4
rlabel comment s 13730 1268 13730 1268 4 buf_1
rlabel comment s 14558 1268 14558 1268 4 buf_16
rlabel comment s 14006 1268 14006 1268 4 buf_4
flabel metal2 16399 -322 16441 915 0 FreeSans 320 0 0 0 VDD_SW_b[1]
port 30 nsew
flabel metal2 14006 -322 14048 913 0 FreeSans 320 0 0 0 VDD_SW_b[2]
port 31 nsew
flabel metal2 11613 -322 11655 914 0 FreeSans 320 0 0 0 VDD_SW_b[3]
port 32 nsew
flabel metal2 9222 -322 9264 915 0 FreeSans 320 0 0 0 VDD_SW_b[4]
port 33 nsew
flabel metal2 4438 -322 4480 914 0 FreeSans 320 0 0 0 VDD_SW_b[6]
port 35 nsew
flabel metal2 2046 -322 2088 913 0 FreeSans 320 0 0 0 VDD_SW_b[7]
port 36 nsew
rlabel comment s 276 580 276 580 4 buf_4
rlabel comment s 828 580 828 580 4 buf_16
rlabel comment s 0 580 0 580 4 buf_1
rlabel comment s 2852 580 2852 580 4 buf_1
rlabel comment s 3680 580 3680 580 4 buf_16
rlabel comment s 3128 580 3128 580 4 buf_4
rlabel comment s 5980 580 5980 580 4 buf_4
rlabel comment s 6532 580 6532 580 4 buf_16
rlabel comment s 5704 580 5704 580 4 buf_1
rlabel comment s 8556 580 8556 580 4 buf_1
rlabel comment s 9384 580 9384 580 4 buf_16
rlabel comment s 8832 580 8832 580 4 buf_4
rlabel comment s 11408 580 11408 580 4 buf_1
rlabel comment s 12236 580 12236 580 4 buf_16
rlabel comment s 11684 580 11684 580 4 buf_4
rlabel comment s 14260 580 14260 580 4 buf_1
rlabel comment s 15088 580 15088 580 4 buf_16
rlabel comment s 14536 580 14536 580 4 buf_4
flabel metal2 14653 -343 14695 234 0 FreeSans 320 0 0 0 VSS_SW_b[1]
port 37 nsew
flabel metal2 12260 -343 12302 235 0 FreeSans 320 0 0 0 VSS_SW_b[2]
port 38 nsew
flabel metal2 9869 -343 9911 234 0 FreeSans 320 0 0 0 VSS_SW_b[3]
port 39 nsew
flabel metal2 7477 -343 7519 234 0 FreeSans 320 0 0 0 VSS_SW_b[4]
port 40 nsew
flabel metal2 5084 -343 5126 234 0 FreeSans 320 0 0 0 VSS_SW_b[5]
port 41 nsew
flabel metal2 2693 -343 2735 234 0 FreeSans 320 0 0 0 VSS_SW_b[6]
port 42 nsew
flabel metal2 301 -343 343 234 0 FreeSans 320 0 0 0 VSS_SW_b[7]
port 44 nsew
flabel metal2 14493 346 14535 3300 0 FreeSans 320 0 0 0 VSS_SW[1]
port 4 nsew
flabel metal2 12102 346 12144 3300 0 FreeSans 320 0 0 0 VSS_SW[2]
port 5 nsew
flabel metal1 -126 2526 4302 2560 0 FreeSans 320 0 0 0 ready
port 51 nsew
flabel metal1 -126 2722 -34 2756 0 FreeSans 320 0 0 0 reset
port 52 nsew
flabel metal2 6829 -322 6871 914 0 FreeSans 320 0 0 0 VDD_SW_b[5]
port 34 nsew
flabel metal4 8673 2721 16604 3041 0 FreeSans 1600 0 0 0 VDD
port 58 nsew
flabel metal4 12406 -75 16876 114 0 FreeSans 1600 0 0 0 VSS
port 59 nsew
<< end >>
