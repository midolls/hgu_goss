magic
tech sky130A
timestamp 1699890160
<< psubdiff >>
rect 9808 -899 9830 -853
<< metal4 >>
rect 9593 -797 9615 -751
rect 9837 -799 9859 -753
rect 9776 -1059 9798 -1013
use hgu_cdac_unit  x1[0]
timestamp 1699890160
transform 1 0 7245 0 1 -1822
box 343 299 679 913
use hgu_cdac_unit  x1[1]
timestamp 1699890160
transform -1 0 8267 0 -1 -30
box 343 299 679 913
use hgu_cdac_unit  x1[2]
timestamp 1699890160
transform 1 0 7548 0 1 -1822
box 343 299 679 913
use hgu_cdac_unit  x1[3]
timestamp 1699890160
transform -1 0 8570 0 -1 -30
box 343 299 679 913
use hgu_cdac_unit  x1[4]
timestamp 1699890160
transform 1 0 7851 0 1 -1822
box 343 299 679 913
use hgu_cdac_unit  x1[5]
timestamp 1699890160
transform -1 0 8873 0 -1 -30
box 343 299 679 913
use hgu_cdac_unit  x1[6]
timestamp 1699890160
transform 1 0 8154 0 1 -1822
box 343 299 679 913
use hgu_cdac_unit  x1[7]
timestamp 1699890160
transform -1 0 9176 0 -1 -30
box 343 299 679 913
use hgu_cdac_unit  x1[8]
timestamp 1699890160
transform 1 0 8457 0 1 -1822
box 343 299 679 913
use hgu_cdac_unit  x1[9]
timestamp 1699890160
transform -1 0 9479 0 -1 -30
box 343 299 679 913
use hgu_cdac_unit  x1[10]
timestamp 1699890160
transform 1 0 8760 0 1 -1822
box 343 299 679 913
use hgu_cdac_unit  x1[11]
timestamp 1699890160
transform -1 0 9782 0 -1 -30
box 343 299 679 913
use hgu_cdac_unit  x1[12]
timestamp 1699890160
transform 1 0 9063 0 1 -1822
box 343 299 679 913
use hgu_cdac_unit  x1[13]
timestamp 1699890160
transform -1 0 10085 0 -1 -30
box 343 299 679 913
use hgu_cdac_unit  x1[14]
timestamp 1699890160
transform 1 0 9366 0 1 -1822
box 343 299 679 913
use hgu_cdac_unit  x1[15]
timestamp 1699890160
transform -1 0 10388 0 -1 -30
box 343 299 679 913
use hgu_cdac_unit  x1[16]
timestamp 1699890160
transform 1 0 9669 0 1 -1822
box 343 299 679 913
use hgu_cdac_unit  x1[17]
timestamp 1699890160
transform -1 0 10691 0 -1 -30
box 343 299 679 913
use hgu_cdac_unit  x1[18]
timestamp 1699890160
transform 1 0 9972 0 1 -1822
box 343 299 679 913
use hgu_cdac_unit  x1[19]
timestamp 1699890160
transform -1 0 10994 0 -1 -30
box 343 299 679 913
use hgu_cdac_unit  x1[20]
timestamp 1699890160
transform 1 0 10275 0 1 -1822
box 343 299 679 913
use hgu_cdac_unit  x1[21]
timestamp 1699890160
transform -1 0 11297 0 -1 -30
box 343 299 679 913
use hgu_cdac_unit  x1[22]
timestamp 1699890160
transform 1 0 10578 0 1 -1822
box 343 299 679 913
use hgu_cdac_unit  x1[23]
timestamp 1699890160
transform -1 0 11600 0 -1 -30
box 343 299 679 913
use hgu_cdac_unit  x1[24]
timestamp 1699890160
transform 1 0 10881 0 1 -1822
box 343 299 679 913
use hgu_cdac_unit  x1[25]
timestamp 1699890160
transform -1 0 11903 0 -1 -30
box 343 299 679 913
use hgu_cdac_unit  x1[26]
timestamp 1699890160
transform 1 0 11184 0 1 -1822
box 343 299 679 913
use hgu_cdac_unit  x1[27]
timestamp 1699890160
transform -1 0 12206 0 -1 -30
box 343 299 679 913
use hgu_cdac_unit  x1[28]
timestamp 1699890160
transform 1 0 11487 0 1 -1822
box 343 299 679 913
use hgu_cdac_unit  x1[29]
timestamp 1699890160
transform -1 0 12509 0 -1 -30
box 343 299 679 913
use hgu_cdac_unit  x1[30]
timestamp 1699890160
transform 1 0 11790 0 1 -1822
box 343 299 679 913
use hgu_cdac_unit  x1[31]
timestamp 1699890160
transform -1 0 12812 0 -1 -30
box 343 299 679 913
<< labels >>
flabel psubdiff 9808 -899 9830 -853 0 FreeSans 160 0 0 0 SUB
port 2 nsew
flabel metal4 9593 -797 9615 -751 0 FreeSans 160 0 0 0 CBOT
port 4 nsew
flabel metal4 9837 -799 9859 -753 0 FreeSans 160 0 0 0 CTOP
port 6 nsew
flabel metal4 9776 -1059 9798 -1013 0 FreeSans 160 0 0 0 CTOP
port 8 nsew
<< end >>
