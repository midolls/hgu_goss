* NGSPICE file created from hgu_sarlogic_8bit_logic_flat.ext - technology: sky130A

.subckt hgu_sarlogic_8bit_logic_RC sel_bit[0] sel_bit[1] eob clk_sar D[0] D[1] D[2] D[3] D[4] D[5] D[6] D[7] comparator_out check[0] check[1] check[2] check[3] check[4] check[5] check[6] reset VDD VSS
X0 VDD.t263 a_10680_2340# D[3].t0 VDD.t262 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X1 VDD.t266 a_8289_4086# check[1].t0 VDD.t265 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X2 VDD.t333 D[0].t2 a_8236_3239# VDD.t332 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3 VDD.t585 a_2389_5648# eob.t3 VDD.t584 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.135 ps=1.27 w=1 l=0.15
X4 a_12030_3213# a_11856_3239# a_12146_3239# VSS.t550 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X5 a_4971_4801# VDD.t725 VSS.t246 VSS.t245 sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X6 a_2147_5083# a_1682_4775# VDD.t542 VDD.t541 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X7 a_1822_4801# x4.X.t32 VSS.t543 VSS.t542 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X8 a_11330_2340# a_11628_2640# a_11564_2732# VDD.t261 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0924 ps=0.86 w=0.42 l=0.15
X9 VSS.t586 a_12030_3213# a_12737_3239# VSS.t585 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X10 a_4213_3239# a_4367_3213# a_4073_3213# VSS.t533 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X11 a_8591_4801# check[5].t2 VSS.t150 VSS.t149 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X12 a_9710_4296# a_9238_4086# a_9954_4478# VDD.t609 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X13 VSS.t605 x30.Q_N a_7185_2366# VSS.t604 sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.101 ps=0.99 w=0.42 l=0.15
X14 VDD.t156 a_11250_4775# a_11160_5167# VDD.t155 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X15 VSS.t570 a_5992_4086# x45.Q_N VSS.t569 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X16 a_3599_2340# a_3912_2366# a_4018_2366# VSS.t600 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X17 x72.Q_N a_7246_3213# VSS.t144 VSS.t143 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X18 VSS.t521 x27.Q_N a_4018_2366# VSS.t520 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.12 ps=1.08 w=0.42 l=0.15
X19 a_4854_3213# x77.Y VDD.t7 VDD.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X20 a_7072_3239# a_5844_3239# a_6930_3521# VDD.t637 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X21 a_9442_4086# a_8697_4112# a_9578_4112# VSS.t116 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X22 VSS.t263 x4.X.t33 a_9151_3213# VSS.t262 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X23 VDD.t137 a_7246_3213# a_7158_3605# VDD.t136 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X24 VDD.t180 a_5897_4086# check[0].t1 VDD.t179 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X25 a_11089_4112# x4.X.t34 VDD.t276 VDD.t275 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.154 ps=1.34 w=0.64 l=0.15
X26 a_4793_2366# a_4925_2550# a_4657_2340# VSS.t410 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0864 ps=0.91 w=0.64 l=0.15
X27 VDD.t170 x75.Q a_5844_3239# VDD.t169 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X28 a_6978_4801# a_6466_4775# VSS.t529 VSS.t528 sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X29 a_4388_2732# a_3599_2340# VDD.t712 VDD.t711 sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0819 ps=0.81 w=0.42 l=0.15
X30 a_2788_5674# check[2].t2 VSS.t136 VSS.t135 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.107 ps=1 w=0.42 l=0.15
X31 a_10794_3239# a_10628_3239# VDD.t337 VDD.t336 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X32 VSS.t45 D[0].t3 a_8236_3239# VSS.t44 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X33 VDD.t325 x4.X.t35 a_4368_4775# VDD.t324 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X34 a_9465_4801# a_8403_4801# a_9370_4801# VSS.t592 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X35 VSS.t484 a_1511_4112# x4.X.t15 VSS.t483 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X36 a_12048_4394# a_11089_4112# VDD.t3 VDD.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X37 a_9101_3521# a_8683_3605# a_8857_3213# VDD.t533 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X38 a_7247_4775# VDD.t257 VDD.t259 VDD.t258 sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X39 VDD.t107 a_6846_4086# a_6845_4386# VDD.t106 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X40 VSS.t541 x20.Q_N a_1626_2366# VSS.t540 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.12 ps=1.08 w=0.42 l=0.15
X41 D[2].t0 a_12737_3239# VSS.t580 VSS.t579 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X42 a_11250_4775# a_11076_5167# a_11390_4801# VSS.t28 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X43 a_4680_3239# a_3452_3239# a_4538_3521# VDD.t200 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X44 a_2479_2648# a_1520_2366# VDD.t694 VDD.t693 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X45 VDD.t349 a_4854_3213# a_4766_3605# VDD.t348 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X46 a_11184_4801# a_10795_4801# a_11076_5167# VSS.t91 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X47 VSS.t609 a_1338_5674# x5.X.t1 VSS.t608 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X48 a_2784_5996# check[2].t3 VDD.t129 VDD.t128 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=0.995 as=0.154 ps=1.34 w=0.64 l=0.15
X49 a_4593_4112# a_4453_4386# a_4155_4086# VSS.t138 sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.0711 ps=0.755 w=0.36 l=0.15
X50 a_1996_2732# a_1207_2340# VDD.t331 VDD.t330 sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0819 ps=0.81 w=0.42 l=0.15
X51 a_7181_3239# a_5844_3239# a_7072_3239# VSS.t598 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X52 a_6198_3239# comparator_out.t0 VSS.t353 VSS.t352 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X53 x4.X.t31 a_1511_4112# VDD.t511 VDD.t510 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X54 a_2265_2340# a_1520_2366# a_2401_2366# VSS.t643 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X55 a_12031_4775# a_11857_4801# a_12147_4801# VSS.t662 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X56 VSS.t178 x75.Q a_5844_3239# VSS.t177 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X57 VDD.t256 VDD.t254 a_1976_4775# VDD.t255 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X58 VSS.t549 a_7050_4086# a_6985_4112# VSS.t548 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0935 ps=0.965 w=0.64 l=0.15
X59 a_1762_2340# a_2060_2640# a_1996_2732# VDD.t164 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0924 ps=0.86 w=0.42 l=0.15
X60 VDD.t447 check[1].t2 a_2969_6040# VDD.t446 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.138 ps=1.16 w=0.64 l=0.15
X61 a_2883_5674# a_2853_5648# a_2788_5674# VSS.t407 sky130_fd_pr__nfet_01v8 ad=0.072 pd=0.76 as=0.066 ps=0.745 w=0.36 l=0.15
X62 a_7562_4478# a_7050_4086# VDD.t576 VDD.t575 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X63 a_10775_2340# a_11088_2366# a_11194_2366# VSS.t397 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X64 a_6504_2648# a_6304_2366# VDD.t322 VDD.t321 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X65 a_4214_4801# a_4368_4775# a_4074_4775# VSS.t210 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X66 VSS.t261 x36.Q_N a_11194_2366# VSS.t260 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.12 ps=1.08 w=0.42 l=0.15
X67 a_10794_3239# a_10628_3239# VSS.t314 VSS.t313 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X68 a_1511_4112# x4.A VSS.t286 VSS.t285 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X69 a_4855_4775# VDD.t251 VDD.t253 VDD.t252 sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X70 a_7073_4801# a_5845_4801# a_6931_5083# VDD.t392 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X71 VDD.t519 a_4454_4086# a_4453_4386# VDD.t518 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X72 VDD.t366 a_7247_4775# a_7159_5167# VDD.t365 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X73 x4.A a_897_4112# VDD.t386 VDD.t385 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X74 x30.Q_N a_7247_4775# VSS.t343 VSS.t342 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X75 x4.X.t30 a_1511_4112# VDD.t509 VDD.t508 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X76 a_12345_2732# a_11833_2340# VDD.t360 VDD.t359 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X77 VSS.t412 check[0].t2 a_5372_4112# VSS.t411 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X78 a_8803_4112# a_8939_4086# a_8384_4086# VSS.t189 sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0864 ps=0.91 w=0.64 l=0.15
X79 VSS.t304 x4.X.t36 a_9152_4775# VSS.t303 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X80 a_3806_3239# VSS.t68 VSS.t70 VSS.t69 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X81 VDD.t570 x20.Q_N a_1207_2340# VDD.t569 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.123 ps=1.17 w=0.42 l=0.15
X82 VSS.t133 check[1].t3 a_2993_5674# VSS.t132 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0786 ps=0.805 w=0.42 l=0.15
X83 VSS.t244 VDD.t726 a_8803_4112# VSS.t243 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.12 ps=1.08 w=0.42 l=0.15
X84 VSS.t80 a_10776_4086# x39.Q_N VSS.t79 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X85 a_6291_3605# a_5844_3239# a_6198_3239# VSS.t597 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X86 x75.Q_N a_4854_3213# VDD.t347 VDD.t346 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X87 VSS.t7 x5.X.t4 a_8237_4801# VSS.t6 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X88 VSS.t507 a_6465_3213# a_6399_3239# VSS.t506 sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X89 a_1822_4801# a_1976_4775# a_1682_4775# VSS.t442 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X90 VDD.t162 a_10775_2340# x63.Q_N VDD.t161 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X91 a_9102_5083# a_8684_5167# a_8858_4775# VDD.t78 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X92 a_11856_3239# a_10628_3239# a_11714_3521# VDD.t335 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X93 a_4681_4801# a_3453_4801# a_4539_5083# VDD.t523 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X94 VDD.t686 a_4855_4775# a_4767_5167# VDD.t685 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X95 a_9953_2366# a_9441_2340# VSS.t154 VSS.t153 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.084 ps=0.82 w=0.42 l=0.15
X96 check[3].t0 a_12738_4801# VSS.t333 VSS.t332 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X97 a_1112_2340# a_1207_2340# VSS.t310 VSS.t309 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X98 a_11769_4112# a_11629_4386# a_11331_4086# VSS.t269 sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.0711 ps=0.755 w=0.36 l=0.15
X99 a_2579_4801# x4.X.t37 VSS.t432 VSS.t431 sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X100 a_4155_4086# a_4453_4386# a_4389_4478# VDD.t131 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0924 ps=0.86 w=0.42 l=0.15
X101 a_7480_3521# a_7072_3239# a_7246_3213# VDD.t182 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X102 VSS.t242 VDD.t727 a_9578_4112# VSS.t241 sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.101 ps=0.99 w=0.42 l=0.15
X103 a_5992_4086# a_6305_4112# a_6411_4112# VSS.t379 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X104 VDD.t376 comparator_out.t1 a_12547_2366# VDD.t375 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0662 ps=0.735 w=0.42 l=0.15
X105 a_6199_4801# check[6].t2 VSS.t625 VSS.t624 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X106 a_7182_4801# a_5845_4801# a_7073_4801# VSS.t369 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X107 VSS.t240 VDD.t728 a_6411_4112# VSS.t239 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.12 ps=1.08 w=0.42 l=0.15
X108 VDD.t455 x4.X.t38 a_6759_3213# VDD.t454 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X109 x33.Q_N a_9639_4775# VSS.t97 VSS.t96 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X110 VSS.t519 x27.Q_N a_4793_2366# VSS.t518 sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.101 ps=0.99 w=0.42 l=0.15
X111 a_3899_3605# a_3452_3239# a_3806_3239# VSS.t206 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X112 VSS.t420 x5.X.t5 a_5845_4801# VSS.t419 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X113 D[1].t1 a_10345_3239# VDD.t459 VDD.t458 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X114 a_6710_5083# a_6292_5167# a_6466_4775# VDD.t538 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X115 a_11195_4112# a_11331_4086# a_10776_4086# VSS.t327 sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0864 ps=0.91 w=0.64 l=0.15
X116 a_6375_3605# a_5844_3239# a_6291_3605# VDD.t636 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X117 a_2969_6040# a_2853_5648# a_2883_5674# VDD.t434 sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.16 as=0.0567 ps=0.69 w=0.42 l=0.15
X118 a_8288_2340# a_8383_2340# VDD.t400 VDD.t399 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X119 a_10795_4801# a_10629_4801# VSS.t267 VSS.t266 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X120 a_7050_4086# a_6305_4112# a_7186_4112# VSS.t378 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X121 a_11965_3239# a_10628_3239# a_11856_3239# VSS.t312 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X122 a_12102_4296# a_11629_4386# a_12346_4112# VSS.t268 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0671 ps=0.75 w=0.36 l=0.15
X123 VSS.t202 a_2463_4775# a_3170_4801# VSS.t201 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X124 a_11970_4112# a_12102_4296# a_11834_4086# VSS.t29 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0864 ps=0.91 w=0.64 l=0.15
X125 VDD.t120 a_3505_4086# x48.Q VDD.t119 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X126 a_8590_3239# comparator_out.t2 VDD.t116 VDD.t115 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X127 VDD.t152 VSS.t674 a_3452_3239# VDD.t151 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X128 x4.X.t29 a_1511_4112# VDD.t507 VDD.t506 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X129 a_4113_4394# a_3913_4112# VDD.t141 VDD.t140 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X130 VSS.t347 a_11834_4086# a_11769_4112# VSS.t346 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0935 ps=0.965 w=0.64 l=0.15
X131 a_3807_4801# x27.D VSS.t371 VSS.t370 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X132 a_4790_4801# a_3453_4801# a_4681_4801# VSS.t494 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X133 VSS.t539 x20.Q_N a_2401_2366# VSS.t538 sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.101 ps=0.99 w=0.42 l=0.15
X134 a_1511_4112# x4.A VSS.t284 VSS.t283 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X135 a_11564_2366# a_10775_2340# VSS.t168 VSS.t167 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0588 ps=0.7 w=0.42 l=0.15
X136 a_7763_2366# a_6844_2640# a_7317_2550# VDD.t633 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X137 a_11714_3521# a_11249_3213# VDD.t188 VDD.t187 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X138 a_11857_4801# a_10629_4801# a_11715_5083# VDD.t280 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X139 x4.A a_897_4112# VDD.t384 VDD.t383 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X140 a_6292_5167# a_5845_4801# a_6199_4801# VSS.t368 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X141 VDD.t329 a_1207_2340# x51.Q_N VDD.t328 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X142 a_3983_3605# a_3452_3239# a_3899_3605# VDD.t199 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X143 a_2389_5648# a_3258_5648# a_2883_5674# VSS.t46 sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X144 a_5896_2340# a_5991_2340# VDD.t58 VDD.t57 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X145 VSS.t527 a_6466_4775# a_6400_4801# VSS.t526 sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X146 a_4658_4086# a_3913_4112# a_4794_4112# VSS.t146 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X147 VDD.t194 a_2463_4775# a_3170_4801# VDD.t193 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X148 a_7481_5083# a_7073_4801# a_7247_4775# VDD.t289 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X149 a_9237_2340# D[3].t2 VDD.t619 VDD.t618 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X150 VDD.t49 reset.t0 a_621_4112# VDD.t48 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X151 a_9173_4112# a_8384_4086# VSS.t185 VSS.t184 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0588 ps=0.7 w=0.42 l=0.15
X152 VDD.t118 comparator_out.t3 a_2979_2366# VDD.t117 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0662 ps=0.735 w=0.42 l=0.15
X153 VDD.t358 a_11833_2340# a_11766_2732# VDD.t357 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X154 VSS.t67 VSS.t65 a_3452_3239# VSS.t66 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X155 VDD.t168 a_9442_4086# a_9375_4478# VDD.t167 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X156 VDD.t650 x30.Q_N a_7049_2340# VDD.t649 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X157 a_4317_3521# a_3899_3605# a_4073_3213# VDD.t114 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X158 a_6376_5167# a_5845_4801# a_6292_5167# VDD.t391 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X159 a_3900_5167# a_3453_4801# a_3807_4801# VSS.t493 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X160 VSS.t377 a_8383_2340# x60.Q_N VSS.t376 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X161 a_11249_3213# x39.Q_N VDD.t343 VDD.t342 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X162 a_1227_4801# a_1061_4801# VSS.t25 VSS.t24 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X163 a_4074_4775# VDD.t248 VDD.t250 VDD.t249 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X164 a_8997_3239# x42.Q_N VSS.t574 VSS.t573 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X165 x5.X.t3 a_1338_5674# VDD.t654 VDD.t653 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X166 a_8591_4801# check[5].t3 VDD.t305 VDD.t304 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X167 a_11289_4394# a_11089_4112# VDD.t1 VDD.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X168 a_1511_4112# x4.A VDD.t303 VDD.t302 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X169 x4.X.t14 a_1511_4112# VSS.t482 VSS.t481 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X170 x75.Q a_5561_3239# VDD.t123 VDD.t122 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X171 a_11966_4801# a_10629_4801# a_11857_4801# VSS.t265 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X172 a_9376_2366# a_9236_2640# a_8938_2340# VSS.t647 sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.0711 ps=0.755 w=0.36 l=0.15
X173 eob.t4 a_2389_5648# VSS.t558 VSS.t557 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X174 a_6781_4112# a_5992_4086# VSS.t568 VSS.t567 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0588 ps=0.7 w=0.42 l=0.15
X175 x77.Y eob.t8 VDD.t196 VDD.t195 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X176 a_9237_2340# D[3].t3 VSS.t588 VSS.t587 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X177 a_11715_5083# a_11250_4775# VDD.t154 VDD.t153 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X178 x27.Q_N a_4855_4775# VDD.t684 VDD.t683 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X179 a_3984_5167# a_3453_4801# a_3900_5167# VDD.t522 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X180 a_8791_3239# a_8402_3239# a_8683_3605# VSS.t43 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X181 a_11089_4112# x4.X.t39 VSS.t502 VSS.t501 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X182 a_5991_2340# a_6546_2340# a_6504_2648# VDD.t716 sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0882 ps=1.05 w=0.84 l=0.15
X183 a_11075_3605# a_10794_3239# a_10982_3239# VDD.t39 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X184 VDD.t439 check[0].t3 a_5372_4112# VDD.t438 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0662 ps=0.735 w=0.42 l=0.15
X185 VDD.t463 a_11629_2340# a_11628_2640# VDD.t462 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X186 a_9638_3213# a_9464_3239# a_9754_3239# VSS.t87 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X187 a_5088_3521# a_4680_3239# a_4854_3213# VDD.t178 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X188 x4.X.t28 a_1511_4112# VDD.t505 VDD.t504 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X189 VDD.t247 VDD.t245 a_9442_4086# VDD.t246 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X190 a_6984_2366# a_6844_2640# a_6546_2340# VSS.t594 sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.0711 ps=0.755 w=0.36 l=0.15
X191 VDD.t527 x4.X.t40 a_4367_3213# VDD.t526 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X192 a_7318_4296# a_6846_4086# a_7562_4478# VDD.t105 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X193 VSS.t152 a_9441_2340# a_9376_2366# VSS.t151 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0935 ps=0.965 w=0.64 l=0.15
X194 a_4318_5083# a_3900_5167# a_4074_4775# VDD.t264 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X195 check[4].t1 a_10346_4801# VDD.t291 VDD.t290 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X196 VDD.t503 a_1511_4112# x4.X.t27 VDD.t502 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X197 a_12101_2550# a_11629_2340# a_12345_2732# VDD.t461 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X198 a_12548_4112# a_11629_4386# a_12102_4296# VDD.t282 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X199 VSS.t422 x5.X.t6 a_3453_4801# VSS.t421 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X200 a_11250_4775# VDD.t230 VDD.t232 VDD.t231 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X201 a_4453_2340# D[5].t2 VDD.t676 VDD.t675 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X202 a_3373_5674# a_3258_5648# a_2389_5648# VDD.t52 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.6 as=0.0729 ps=0.81 w=0.54 l=0.15
X203 VSS.t444 x4.X.t41 a_6759_3213# VSS.t443 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X204 VSS.t172 reset.t1 a_621_4112# VSS.t171 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X205 a_1762_2340# a_2061_2340# a_1996_2366# VSS.t673 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.066 ps=0.745 w=0.36 l=0.15
X206 a_9550_3605# a_8402_3239# a_9464_3239# VDD.t51 sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X207 a_8998_4801# VDD.t729 VSS.t238 VSS.t237 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X208 x4.X.t13 a_1511_4112# VSS.t480 VSS.t479 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X209 a_7049_2340# a_7317_2550# a_7263_2648# VDD.t201 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X210 a_6198_3239# comparator_out.t4 VDD.t451 VDD.t450 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X211 VSS.t428 comparator_out.t5 a_7763_2366# VSS.t427 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X212 a_2398_4801# a_1061_4801# a_2289_4801# VSS.t23 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X213 VSS.t440 a_11629_2340# a_11628_2640# VSS.t439 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X214 VDD.t288 a_6759_3213# a_7480_3521# VDD.t287 sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X215 a_3877_5674# a_2853_5648# a_3373_5674# VSS.t406 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.072 ps=0.76 w=0.36 l=0.15
X216 a_9656_4394# a_8697_4112# VDD.t113 VDD.t112 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X217 a_7185_2366# a_7317_2550# a_7049_2340# VSS.t207 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0864 ps=0.91 w=0.64 l=0.15
X218 a_10155_2366# a_9237_2340# a_9709_2550# VSS.t15 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X219 a_1926_5083# a_1508_5167# a_1682_4775# VDD.t124 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X220 a_9370_4801# a_8858_4775# VSS.t401 VSS.t400 sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X221 a_3504_2340# a_3599_2340# VDD.t710 VDD.t709 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X222 VDD.t244 VDD.t242 a_11834_4086# VDD.t243 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X223 a_11076_5167# a_10795_4801# a_10983_4801# VDD.t88 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X224 a_8792_4801# a_8403_4801# a_8684_5167# VSS.t591 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X225 a_5089_5083# a_4681_4801# a_4855_4775# VDD.t127 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X226 x4.X.t12 a_1511_4112# VSS.t478 VSS.t477 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X227 VDD.t724 a_2061_2340# a_2060_2640# VDD.t723 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X228 a_3671_5674# x48.Q VSS.t89 VSS.t88 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0819 ps=0.81 w=0.42 l=0.15
X229 a_4453_2340# D[5].t3 VSS.t627 VSS.t626 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X230 a_4657_2340# a_4925_2550# a_4871_2648# VDD.t437 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X231 a_3806_3239# VSS.t675 VDD.t284 VDD.t283 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X232 a_9639_4775# a_9465_4801# a_9755_4801# VSS.t655 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X233 VDD.t617 a_12030_3213# a_12737_3239# VDD.t616 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X234 a_4970_3239# a_4367_3213# a_4854_3213# VSS.t532 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X235 a_8857_3213# a_8683_3605# a_8997_3239# VSS.t508 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X236 a_3600_4086# a_4155_4086# a_4113_4394# VDD.t171 sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0882 ps=1.05 w=0.84 l=0.15
X237 a_8383_2340# a_8696_2366# a_8802_2366# VSS.t31 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X238 VDD.t532 a_6465_3213# a_6375_3605# VDD.t531 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X239 VSS.t58 check[0].t4 a_3877_5674# VSS.t57 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.066 ps=0.745 w=0.42 l=0.15
X240 VSS.t200 a_2463_4775# a_2398_4801# VSS.t199 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X241 VSS.t253 a_8289_4086# check[1].t1 VSS.t252 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X242 x5.A a_1062_5674# VDD.t21 VDD.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X243 VDD.t60 check[0].t5 a_3876_6040# VDD.t59 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.0974 ps=0.97 w=0.64 l=0.15
X244 a_11390_4801# VDD.t730 VSS.t236 VSS.t235 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X245 VSS.t52 a_5991_2340# x57.Q_N VSS.t51 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X246 a_4590_2732# a_4453_2340# a_4154_2340# VDD.t432 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X247 VDD.t566 a_8288_2340# D[4].t1 VDD.t565 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X248 VSS.t125 comparator_out.t6 a_10155_2366# VSS.t124 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X249 a_9953_2732# a_9441_2340# VDD.t146 VDD.t145 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X250 a_8289_4086# a_8384_4086# VDD.t177 VDD.t176 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X251 a_2697_5083# a_2289_4801# a_2463_4775# VDD.t705 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X252 a_9551_5167# a_8403_4801# a_9465_4801# VDD.t631 sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X253 a_9441_2340# a_8696_2366# a_9577_2366# VSS.t30 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X254 a_6199_4801# check[6].t3 VDD.t674 VDD.t673 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X255 a_11630_4086# x5.X.t7 VSS.t590 VSS.t589 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X256 VSS.t446 x4.X.t42 a_6760_4775# VSS.t445 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X257 a_5170_4112# a_4658_4086# VSS.t395 VSS.t394 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.084 ps=0.82 w=0.42 l=0.15
X258 a_10680_2340# a_10775_2340# VSS.t166 VSS.t165 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X259 VSS.t60 sel_bit[1].t0 a_3258_5648# VSS.t59 sky130_fd_pr__nfet_01v8 ad=0.0819 pd=0.81 as=0.113 ps=1.38 w=0.42 l=0.15
X260 a_9173_4478# a_8384_4086# VDD.t175 VDD.t174 sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0819 ps=0.81 w=0.42 l=0.15
X261 VDD.t658 sel_bit[1].t1 a_3258_5648# VDD.t657 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X262 check[6].t1 a_5562_4801# VDD.t97 VDD.t96 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X263 VDD.t101 a_6760_4775# a_7481_5083# VDD.t100 sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X264 a_4389_4112# a_3600_4086# VSS.t292 VSS.t291 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0588 ps=0.7 w=0.42 l=0.15
X265 a_5372_4112# a_4454_4086# a_4926_4296# VSS.t490 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X266 a_9375_4478# a_9238_4086# a_8939_4086# VDD.t608 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X267 VSS.t672 a_2061_2340# a_2060_2640# VSS.t671 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X268 a_6465_3213# a_6291_3605# a_6605_3239# VSS.t295 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X269 VSS.t188 a_5897_4086# check[0].t0 VSS.t187 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X270 a_6399_3239# a_6010_3239# a_6291_3605# VSS.t17 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X271 VSS.t661 a_3599_2340# x54.Q_N VSS.t660 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X272 eob.t2 a_2389_5648# VDD.t583 VDD.t582 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.335 ps=2.67 w=1 l=0.15
X273 VDD.t621 x5.X.t8 a_1061_4801# VDD.t620 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X274 VDD.t378 a_5896_2340# D[5].t1 VDD.t377 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X275 VDD.t546 x27.Q_N a_3599_2340# VDD.t545 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.123 ps=1.17 w=0.42 l=0.15
X276 a_11389_3239# a_11543_3213# a_11249_3213# VSS.t619 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X277 VDD.t420 a_4658_4086# a_4591_4478# VDD.t419 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X278 VDD.t15 a_9237_2340# a_9236_2640# VDD.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X279 a_5897_4086# a_5992_4086# VDD.t601 VDD.t600 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X280 a_8289_4086# a_8384_4086# VSS.t183 VSS.t182 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X281 a_6304_2366# x4.X.t43 VSS.t424 VSS.t423 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X282 a_3807_4801# x27.D VDD.t394 VDD.t393 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X283 a_12146_3239# x39.Q_N VSS.t320 VSS.t319 sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X284 VSS.t615 a_12031_4775# a_12738_4801# VSS.t614 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X285 a_6781_4478# a_5992_4086# VDD.t599 VDD.t598 sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0819 ps=0.81 w=0.42 l=0.15
X286 VSS.t564 a_1112_2340# D[7].t0 VSS.t563 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X287 a_12146_3239# a_11543_3213# a_12030_3213# VSS.t618 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X288 a_6983_4478# a_6846_4086# a_6547_4086# VDD.t104 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X289 VDD.t241 VDD.t239 a_8384_4086# VDD.t240 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.123 ps=1.17 w=0.42 l=0.15
X290 a_9238_4086# x5.X.t9 VDD.t67 VDD.t66 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X291 a_12047_2648# a_11088_2366# VDD.t424 VDD.t423 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X292 a_6546_2340# a_6844_2640# a_6780_2732# VDD.t632 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0924 ps=0.86 w=0.42 l=0.15
X293 a_1520_2366# x4.X.t44 VDD.t443 VDD.t442 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.154 ps=1.34 w=0.64 l=0.15
X294 a_4585_3239# a_4073_3213# VSS.t641 VSS.t640 sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X295 VDD.t554 a_6466_4775# a_6376_5167# VDD.t553 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X296 VSS.t651 a_7049_2340# a_6984_2366# VSS.t650 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0935 ps=0.965 w=0.64 l=0.15
X297 a_11564_2732# a_10775_2340# VDD.t160 VDD.t159 sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0819 ps=0.81 w=0.42 l=0.15
X298 x4.X.t26 a_1511_4112# VDD.t501 VDD.t500 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X299 a_11766_2732# a_11629_2340# a_11330_2340# VDD.t460 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X300 a_11833_2340# a_11088_2366# a_11969_2366# VSS.t396 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X301 a_4971_4801# a_4368_4775# a_4855_4775# VSS.t209 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X302 a_4155_4086# a_4454_4086# a_4389_4112# VSS.t489 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.066 ps=0.745 w=0.36 l=0.15
X303 a_10156_4112# a_9237_4386# a_9710_4296# VDD.t372 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X304 a_7072_3239# a_6010_3239# a_6977_3239# VSS.t16 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X305 a_4007_3239# a_3618_3239# a_3899_3605# VSS.t114 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X306 a_8858_4775# a_8684_5167# a_8998_4801# VSS.t81 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X307 x4.X.t11 a_1511_4112# VSS.t476 VSS.t475 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X308 VDD.t644 x4.X.t45 a_11544_4775# VDD.t643 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X309 a_6305_4112# x4.X.t46 VDD.t646 VDD.t645 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.154 ps=1.34 w=0.64 l=0.15
X310 a_4018_2366# a_4154_2340# a_3599_2340# VSS.t98 sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0864 ps=0.91 w=0.64 l=0.15
X311 a_5897_4086# a_5992_4086# VSS.t566 VSS.t565 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X312 VDD.t664 a_12031_4775# a_12738_4801# VDD.t663 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X313 a_3912_2366# x4.X.t47 VSS.t531 VSS.t530 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X314 a_7158_3605# a_6010_3239# a_7072_3239# VDD.t17 sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X315 a_12346_4112# a_11834_4086# VSS.t345 VSS.t344 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.084 ps=0.82 w=0.42 l=0.15
X316 a_9578_4112# a_9710_4296# a_9442_4086# VSS.t433 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0864 ps=0.91 w=0.64 l=0.15
X317 a_12548_4112# a_11630_4086# a_12102_4296# VSS.t450 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X318 VDD.t173 a_8384_4086# x42.Q_N VDD.t172 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X319 VSS.t14 a_9237_2340# a_9236_2640# VSS.t13 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X320 a_4925_2550# a_4452_2640# a_5169_2366# VSS.t108 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0671 ps=0.75 w=0.36 l=0.15
X321 VDD.t238 VDD.t236 a_5992_4086# VDD.t237 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.123 ps=1.17 w=0.42 l=0.15
X322 x4.A a_897_4112# VSS.t363 VSS.t362 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X323 VSS.t11 a_4657_2340# a_4592_2366# VSS.t10 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0935 ps=0.965 w=0.64 l=0.15
X324 x5.A a_1062_5674# VSS.t21 VSS.t20 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X325 x4.X.t10 a_1511_4112# VSS.t474 VSS.t473 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X326 a_2579_4801# a_1976_4775# a_2463_4775# VSS.t441 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X327 VDD.t274 x36.Q_N a_10775_2340# VDD.t273 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.123 ps=1.17 w=0.42 l=0.15
X328 a_4680_3239# a_3618_3239# a_4585_3239# VSS.t113 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X329 a_6466_4775# a_6292_5167# a_6606_4801# VSS.t513 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X330 VDD.t301 x4.A a_1511_4112# VDD.t300 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X331 a_3913_4112# x4.X.t48 VDD.t556 VDD.t555 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.154 ps=1.34 w=0.64 l=0.15
X332 a_1626_2366# a_1762_2340# a_1207_2340# VSS.t364 sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0864 ps=0.91 w=0.64 l=0.15
X333 VSS.t41 a_9638_3213# a_10345_3239# VSS.t40 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X334 VDD.t564 a_9151_3213# a_9101_3521# VDD.t563 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X335 a_1112_2340# a_1207_2340# VDD.t327 VDD.t326 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X336 a_11390_4801# a_11544_4775# a_11250_4775# VSS.t486 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X337 VSS.t112 a_6846_4086# a_6845_4386# VSS.t111 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X338 a_4766_3605# a_3618_3239# a_4680_3239# VDD.t109 sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X339 x75.Q_N a_4854_3213# VSS.t326 VSS.t325 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X340 VDD.t471 a_11630_4086# a_11629_4386# VDD.t470 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X341 a_2533_2550# a_2060_2640# a_2777_2366# VSS.t170 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0671 ps=0.75 w=0.36 l=0.15
X342 a_2401_2366# a_2533_2550# a_2265_2340# VSS.t120 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0864 ps=0.91 w=0.64 l=0.15
X343 a_12147_4801# VDD.t731 VSS.t234 VSS.t233 sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X344 VSS.t294 check[3].t2 a_12548_4112# VSS.t293 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X345 a_12147_4801# a_11544_4775# a_12031_4775# VSS.t485 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X346 a_10982_3239# comparator_out.t7 VSS.t127 VSS.t126 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X347 a_4586_4801# a_4074_4775# VSS.t64 VSS.t63 sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X348 a_2198_2732# a_2061_2340# a_1762_2340# VDD.t722 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X349 a_8857_3213# x42.Q_N VDD.t605 VDD.t604 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X350 a_8403_4801# a_8237_4801# VDD.t537 VDD.t536 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X351 a_4008_4801# a_3619_4801# a_3900_5167# VSS.t500 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X352 a_7073_4801# a_6011_4801# a_6978_4801# VSS.t560 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X353 x66.Q_N a_12030_3213# VDD.t615 VDD.t614 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X354 VDD.t286 a_6759_3213# a_6709_3521# VDD.t285 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X355 a_7159_5167# a_6011_4801# a_7073_4801# VDD.t589 sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X356 a_4454_4086# x5.X.t10 VDD.t69 VDD.t68 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X357 VSS.t488 a_4454_4086# a_4453_4386# VSS.t487 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X358 a_8897_4394# a_8697_4112# VDD.t111 VDD.t110 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X359 a_12030_3213# x39.Q_N VDD.t341 VDD.t340 sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X360 D[1].t0 a_10345_3239# VSS.t436 VSS.t435 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X361 a_3373_5674# a_2853_5648# a_3648_5972# VDD.t433 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.164 ps=1.33 w=0.42 l=0.15
X362 a_11331_4086# a_11629_4386# a_11565_4478# VDD.t281 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0924 ps=0.86 w=0.42 l=0.15
X363 a_11856_3239# a_10794_3239# a_11761_3239# VSS.t33 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X364 a_8697_4112# x4.X.t49 VSS.t426 VSS.t425 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X365 a_8683_3605# a_8402_3239# a_8590_3239# VDD.t50 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X366 D[0].t0 a_7953_3239# VDD.t670 VDD.t669 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X367 a_6011_4801# a_5845_4801# VDD.t390 VDD.t389 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X368 VSS.t259 x36.Q_N a_11969_2366# VSS.t258 sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.101 ps=0.99 w=0.42 l=0.15
X369 a_4681_4801# a_3619_4801# a_4586_4801# VSS.t499 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X370 VDD.t479 a_9152_4775# a_9102_5083# VDD.t478 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X371 VSS.t119 a_3505_4086# x48.Q VSS.t118 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X372 a_4767_5167# a_3619_4801# a_4681_4801# VDD.t525 sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X373 x4.X.t9 a_1511_4112# VSS.t472 VSS.t471 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X374 VSS.t232 VDD.t732 a_1976_4775# VSS.t231 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X375 a_5170_4478# a_4658_4086# VDD.t418 VDD.t417 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X376 a_4112_2648# a_3912_2366# VDD.t641 VDD.t640 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X377 VDD.t126 a_3504_2340# D[6].t1 VDD.t125 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X378 VSS.t95 a_9639_4775# a_10346_4801# VSS.t94 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X379 a_2463_4775# x4.X.t50 VDD.t449 VDD.t448 sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X380 a_3505_4086# a_3600_4086# VDD.t311 VDD.t310 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X381 a_4389_4478# a_3600_4086# VDD.t309 VDD.t308 sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0819 ps=0.81 w=0.42 l=0.15
X382 VDD.t678 comparator_out.t8 a_7763_2366# VDD.t677 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0662 ps=0.735 w=0.42 l=0.15
X383 VSS.t556 a_2389_5648# eob.t7 VSS.t555 sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X384 VDD.t467 a_1976_4775# a_2697_5083# VDD.t466 sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X385 x4.A a_897_4112# VSS.t361 VSS.t360 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X386 x27.Q_N a_4855_4775# VSS.t637 VSS.t636 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X387 a_6411_4112# a_6547_4086# a_5992_4086# VSS.t302 sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0864 ps=0.91 w=0.64 l=0.15
X388 VDD.t299 x4.A a_1511_4112# VDD.t298 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X389 a_8858_4775# VDD.t233 VDD.t235 VDD.t234 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X390 a_10983_4801# check[4].t2 VSS.t391 VSS.t390 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X391 VDD.t99 a_6760_4775# a_6710_5083# VDD.t98 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X392 a_7318_4296# a_6845_4386# a_7562_4112# VSS.t545 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0671 ps=0.75 w=0.36 l=0.15
X393 VDD.t94 a_9639_4775# a_10346_4801# VDD.t93 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X394 a_12031_4775# VDD.t227 VDD.t229 VDD.t228 sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X395 a_1720_2648# a_1520_2366# VDD.t692 VDD.t691 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X396 VSS.t639 a_4073_3213# a_4007_3239# VSS.t638 sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X397 a_3505_4086# a_3600_4086# VSS.t290 VSS.t289 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X398 VSS.t39 a_9638_3213# a_9573_3239# VSS.t38 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X399 a_2289_4801# a_1061_4801# a_2147_5083# VDD.t25 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X400 a_6845_2340# D[4].t2 VDD.t412 VDD.t411 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X401 VDD.t192 a_2463_4775# a_2375_5167# VDD.t191 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X402 a_7561_2366# a_7049_2340# VSS.t649 VSS.t648 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.084 ps=0.82 w=0.42 l=0.15
X403 a_7763_2366# a_6845_2340# a_7317_2550# VSS.t331 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X404 check[4].t0 a_10346_4801# VSS.t274 VSS.t273 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X405 VDD.t499 a_1511_4112# x4.X.t25 VDD.t498 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X406 VDD.t144 a_9441_2340# a_9374_2732# VDD.t143 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X407 VSS.t230 VDD.t733 a_7186_4112# VSS.t229 sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.101 ps=0.99 w=0.42 l=0.15
X408 a_8684_5167# a_8403_4801# a_8591_4801# VDD.t630 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X409 a_11857_4801# a_10795_4801# a_11762_4801# VSS.t90 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X410 VDD.t680 comparator_out.t9 a_10155_2366# VDD.t679 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0662 ps=0.735 w=0.42 l=0.15
X411 a_8938_2340# a_9237_2340# a_9172_2366# VSS.t12 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.066 ps=0.745 w=0.36 l=0.15
X412 a_6930_3521# a_6465_3213# VDD.t530 VDD.t529 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X413 VDD.t382 a_897_4112# x4.A VDD.t381 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X414 a_3600_4086# a_3913_4112# a_4019_4112# VSS.t145 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X415 a_1511_4112# x4.A VSS.t282 VSS.t281 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X416 VSS.t228 VDD.t734 a_4019_4112# VSS.t227 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.12 ps=1.08 w=0.42 l=0.15
X417 a_11288_2648# a_11088_2366# VDD.t422 VDD.t421 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X418 x75.Q a_5561_3239# VSS.t122 VSS.t121 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X419 a_12346_4478# a_11834_4086# VDD.t370 VDD.t369 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X420 x77.Y eob.t9 VSS.t498 VSS.t497 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X421 VDD.t607 a_9238_4086# a_9237_4386# VDD.t606 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X422 a_11493_3521# a_11075_3605# a_11249_3213# VDD.t83 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X423 a_3373_5674# sel_bit[1].t2 a_2389_5648# VSS.t147 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X424 VDD.t307 a_3600_4086# x48.Q_N VDD.t306 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X425 a_9710_4296# a_9237_4386# a_9954_4112# VSS.t349 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0671 ps=0.75 w=0.36 l=0.15
X426 a_6845_2340# D[4].t3 VSS.t387 VSS.t386 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X427 x4.X.t8 a_1511_4112# VSS.t470 VSS.t469 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X428 a_6546_2340# a_6845_2340# a_6780_2366# VSS.t330 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.066 ps=0.745 w=0.36 l=0.15
X429 VSS.t584 a_12030_3213# a_11965_3239# VSS.t583 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X430 a_11075_3605# a_10628_3239# a_10982_3239# VSS.t311 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X431 x69.Q_N a_9638_3213# VDD.t47 VDD.t46 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X432 a_1415_4801# eob.t10 VSS.t496 VSS.t495 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X433 VSS.t196 a_11249_3213# a_11183_3239# VSS.t195 sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X434 VDD.t453 x5.X.t11 a_10629_4801# VDD.t452 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X435 x36.Q_N a_12031_4775# VDD.t662 VDD.t661 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X436 a_5371_2366# a_4452_2640# a_4925_2550# VDD.t103 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X437 VDD.t652 a_1338_5674# x5.X.t2 VDD.t651 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X438 VSS.t62 a_4074_4775# a_4008_4801# VSS.t61 sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X439 a_2993_5674# sel_bit[0].t0 a_2883_5674# VSS.t622 sky130_fd_pr__nfet_01v8 ad=0.0786 pd=0.805 as=0.072 ps=0.76 w=0.36 l=0.15
X440 VSS.t250 a_10680_2340# D[3].t1 VSS.t249 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X441 VDD.t313 check[3].t3 a_12548_4112# VDD.t312 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0662 ps=0.735 w=0.42 l=0.15
X442 VDD.t297 x4.A a_1511_4112# VDD.t296 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X443 VSS.t468 a_1511_4112# x4.X.t7 VSS.t467 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X444 a_12264_3521# a_11856_3239# a_12030_3213# VDD.t577 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X445 VSS.t93 a_9639_4775# a_9574_4801# VSS.t92 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X446 VSS.t554 a_2389_5648# eob.t5 VSS.t553 sky130_fd_pr__nfet_01v8 ad=0.107 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X447 a_6931_5083# a_6466_4775# VDD.t552 VDD.t551 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X448 a_10776_4086# a_11089_4112# a_11195_4112# VSS.t1 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X449 VDD.t35 x4.X.t51 a_11543_3213# VDD.t34 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X450 a_3619_4801# a_3453_4801# VDD.t521 VDD.t520 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X451 VSS.t226 VDD.t735 a_11195_4112# VSS.t225 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.12 ps=1.08 w=0.42 l=0.15
X452 a_2289_4801# a_1227_4801# a_2194_4801# VSS.t664 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X453 check[5].t1 a_7954_4801# VDD.t591 VDD.t590 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X454 a_11494_5083# a_11076_5167# a_11250_4775# VDD.t28 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X455 VDD.t544 x27.Q_N a_4657_2340# VDD.t543 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X456 a_2979_2366# a_2060_2640# a_2533_2550# VDD.t163 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X457 a_11159_3605# a_10628_3239# a_11075_3605# VDD.t334 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X458 check[6].t0 a_5562_4801# VSS.t100 VSS.t99 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X459 VDD.t574 a_7050_4086# a_6983_4478# VDD.t573 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X460 a_9754_3239# x42.Q_N VSS.t572 VSS.t571 sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X461 a_1508_5167# a_1061_4801# a_1415_4801# VSS.t22 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X462 a_9754_3239# a_9151_3213# a_9638_3213# VSS.t535 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X463 VSS.t517 a_1682_4775# a_1616_4801# VSS.t516 sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X464 a_9655_2648# a_8696_2366# VDD.t33 VDD.t32 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X465 VDD.t497 a_1511_4112# x4.X.t24 VDD.t496 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X466 a_8384_4086# a_8939_4086# a_8897_4394# VDD.t181 sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0882 ps=1.05 w=0.84 l=0.15
X467 a_6605_3239# x45.Q_N VSS.t85 VSS.t84 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X468 a_7764_4112# a_6845_4386# a_7318_4296# VDD.t572 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X469 a_3899_3605# a_3618_3239# a_3806_3239# VDD.t108 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X470 a_8938_2340# a_9236_2640# a_9172_2732# VDD.t698 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0924 ps=0.86 w=0.42 l=0.15
X471 a_12547_2366# a_11628_2640# a_12101_2550# VDD.t260 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X472 a_9954_4112# a_9442_4086# VSS.t176 VSS.t175 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.084 ps=0.82 w=0.42 l=0.15
X473 x20.Q_N a_2463_4775# VDD.t190 VDD.t189 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X474 a_11076_5167# a_10629_4801# a_10983_4801# VSS.t264 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X475 VSS.t613 a_12031_4775# a_11966_4801# VSS.t612 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X476 VDD.t495 a_1511_4112# x4.X.t23 VDD.t494 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X477 VDD.t568 x20.Q_N a_2265_2340# VDD.t567 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X478 a_1592_5167# a_1061_4801# a_1508_5167# VDD.t24 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X479 a_8696_2366# x4.X.t52 VDD.t37 VDD.t36 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.154 ps=1.34 w=0.64 l=0.15
X480 a_10680_2340# a_10775_2340# VDD.t158 VDD.t157 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X481 a_5169_2366# a_4657_2340# VSS.t9 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.084 ps=0.82 w=0.42 l=0.15
X482 a_3599_2340# a_4154_2340# a_4112_2648# VDD.t95 sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0882 ps=1.05 w=0.84 l=0.15
X483 a_12265_5083# a_11857_4801# a_12031_4775# VDD.t713 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X484 a_10982_3239# comparator_out.t10 VDD.t184 VDD.t183 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X485 a_7246_3213# a_7072_3239# a_7362_3239# VSS.t190 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X486 VDD.t374 x3.A a_897_4112# VDD.t373 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X487 VDD.t226 VDD.t224 a_7050_4086# VDD.t225 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X488 a_4592_2366# a_4452_2640# a_4154_2340# VSS.t107 sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.0711 ps=0.755 w=0.36 l=0.15
X489 a_8402_3239# a_8236_3239# VDD.t270 VDD.t269 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X490 a_4538_3521# a_4073_3213# VDD.t690 VDD.t689 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X491 a_4926_4296# a_4454_4086# a_5170_4478# VDD.t517 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X492 a_10776_4086# a_11331_4086# a_11289_4394# VDD.t350 sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0882 ps=1.05 w=0.84 l=0.15
X493 VDD.t272 x36.Q_N a_11833_2340# VDD.t271 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X494 a_9709_2550# a_9237_2340# a_9953_2732# VDD.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X495 a_2061_2340# D[6].t2 VDD.t41 VDD.t40 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X496 VSS.t430 x5.X.t12 a_1061_4801# VSS.t429 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X497 a_2777_2366# a_2265_2340# VSS.t669 VSS.t668 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.084 ps=0.82 w=0.42 l=0.15
X498 a_1207_2340# a_1762_2340# a_1720_2648# VDD.t387 sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0882 ps=1.05 w=0.84 l=0.15
X499 a_9755_4801# VDD.t736 VSS.t224 VSS.t223 sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X500 a_2979_2366# a_2061_2340# a_2533_2550# VSS.t670 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X501 VSS.t297 x4.X.t53 a_4367_3213# VSS.t296 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X502 a_9755_4801# a_9152_4775# a_9639_4775# VSS.t452 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X503 a_6606_4801# VDD.t737 VSS.t222 VSS.t221 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X504 a_8802_2366# a_8938_2340# a_8383_2340# VSS.t434 sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0864 ps=0.91 w=0.64 l=0.15
X505 a_11088_2366# x4.X.t54 VDD.t316 VDD.t315 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.154 ps=1.34 w=0.64 l=0.15
X506 VSS.t192 comparator_out.t11 a_5371_2366# VSS.t191 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X507 VDD.t11 a_4657_2340# a_4590_2732# VDD.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X508 a_6010_3239# a_5844_3239# VDD.t635 VDD.t634 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X509 a_11565_4112# a_10776_4086# VSS.t78 VSS.t77 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0588 ps=0.7 w=0.42 l=0.15
X510 VDD.t560 a_4367_3213# a_5088_3521# VDD.t559 sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X511 a_7264_4394# a_6305_4112# VDD.t404 VDD.t403 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X512 a_8402_3239# a_8236_3239# VSS.t257 VSS.t256 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X513 VSS.t158 x33.Q_N a_8802_2366# VSS.t157 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.12 ps=1.08 w=0.42 l=0.15
X514 a_9638_3213# x42.Q_N VDD.t603 VDD.t602 sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X515 VDD.t493 a_1511_4112# x4.X.t22 VDD.t492 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X516 VSS.t164 a_10775_2340# x63.Q_N VSS.t163 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X517 x4.X.t6 a_1511_4112# VSS.t466 VSS.t465 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X518 a_11834_4086# a_12102_4296# a_12048_4394# VDD.t29 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X519 a_3648_5972# x48.Q VDD.t86 VDD.t85 sky130_fd_pr__pfet_01v8_hvt ad=0.164 pd=1.33 as=0.0864 ps=0.91 w=0.64 l=0.15
X520 a_6400_4801# a_6011_4801# a_6292_5167# VSS.t559 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X521 a_10983_4801# check[4].t3 VDD.t416 VDD.t415 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X522 a_6846_4086# x5.X.t13 VDD.t71 VDD.t70 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X523 a_11768_2366# a_11628_2640# a_11330_2340# VSS.t248 sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.0711 ps=0.755 w=0.36 l=0.15
X524 a_2061_2340# D[6].t3 VSS.t35 VSS.t34 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X525 a_4539_5083# a_4074_4775# VDD.t65 VDD.t64 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X526 a_2265_2340# a_2533_2550# a_2479_2648# VDD.t121 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X527 a_6605_3239# a_6759_3213# a_6465_3213# VSS.t271 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X528 a_7247_4775# a_7073_4801# a_7363_4801# VSS.t272 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X529 a_11761_3239# a_11249_3213# VSS.t194 VSS.t193 sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X530 a_12102_4296# a_11630_4086# a_12346_4478# VDD.t469 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X531 VSS.t156 x33.Q_N a_9577_2366# VSS.t155 sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.101 ps=0.99 w=0.42 l=0.15
X532 VDD.t45 a_9638_3213# a_10345_3239# VDD.t44 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X533 VDD.t491 a_1511_4112# x4.X.t21 VDD.t490 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X534 a_4872_4394# a_3913_4112# VDD.t139 VDD.t138 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X535 VSS.t181 a_8384_4086# x42.Q_N VSS.t180 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X536 VDD.t398 a_8383_2340# x60.Q_N VDD.t397 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X537 a_5991_2340# a_6304_2366# a_6410_2366# VSS.t301 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X538 a_6010_3239# a_5844_3239# VSS.t596 VSS.t595 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X539 VDD.t688 a_4073_3213# a_3983_3605# VDD.t687 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X540 a_11331_4086# a_11630_4086# a_11565_4112# VSS.t449 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.066 ps=0.745 w=0.36 l=0.15
X541 VSS.t603 x30.Q_N a_6410_2366# VSS.t602 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.12 ps=1.08 w=0.42 l=0.15
X542 a_9464_3239# a_8236_3239# a_9322_3521# VDD.t268 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X543 VDD.t43 a_9638_3213# a_9550_3605# VDD.t42 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X544 VDD.t380 a_897_4112# x4.A VDD.t379 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X545 VSS.t54 x4.X.t55 a_11543_3213# VSS.t53 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X546 a_11194_2366# a_11330_2340# a_10775_2340# VSS.t148 sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0864 ps=0.91 w=0.64 l=0.15
X547 a_7561_2732# a_7049_2340# VDD.t702 VDD.t701 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X548 a_9377_4112# a_9237_4386# a_8939_4086# VSS.t348 sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.0711 ps=0.755 w=0.36 l=0.15
X549 VSS.t280 x4.A a_1511_4112# VSS.t279 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X550 a_7049_2340# a_6304_2366# a_7185_2366# VSS.t300 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X551 VSS.t56 x4.X.t56 a_4368_4775# VSS.t55 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X552 a_9238_4086# x5.X.t14 VSS.t74 VSS.t73 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X553 a_12101_2550# a_11628_2640# a_12345_2366# VSS.t247 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0671 ps=0.75 w=0.36 l=0.15
X554 eob.t1 a_2389_5648# VDD.t581 VDD.t580 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.175 ps=1.35 w=1 l=0.15
X555 VDD.t668 a_11543_3213# a_12264_3521# VDD.t667 sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X556 x27.D a_3170_4801# VDD.t208 VDD.t207 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X557 VDD.t206 a_4368_4775# a_5089_5083# VDD.t205 sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X558 VDD.t489 a_1511_4112# x4.X.t20 VDD.t488 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X559 a_11969_2366# a_12101_2550# a_11833_2340# VSS.t208 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0864 ps=0.91 w=0.64 l=0.15
X560 VSS.t337 a_11833_2340# a_11768_2366# VSS.t336 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0935 ps=0.965 w=0.64 l=0.15
X561 a_4073_3213# a_3899_3605# a_4213_3239# VSS.t117 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X562 a_9639_4775# VDD.t221 VDD.t223 VDD.t222 sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X563 VSS.t142 a_7246_3213# a_7953_3239# VSS.t141 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X564 VSS.t308 a_1207_2340# x51.Q_N VSS.t307 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X565 a_8403_4801# a_8237_4801# VSS.t512 VSS.t511 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X566 a_6985_4112# a_6845_4386# a_6547_4086# VSS.t544 sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.0711 ps=0.755 w=0.36 l=0.15
X567 a_9573_3239# a_8236_3239# a_9464_3239# VSS.t255 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X568 a_11942_3605# a_10794_3239# a_11856_3239# VDD.t38 sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X569 a_4854_3213# a_4680_3239# a_4970_3239# VSS.t186 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X570 a_4657_2340# a_3912_2366# a_4793_2366# VSS.t599 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X571 x66.Q_N a_12030_3213# VSS.t582 VSS.t581 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X572 a_1415_4801# eob.t11 VDD.t595 VDD.t594 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X573 VSS.t174 a_9442_4086# a_9377_4112# VSS.t173 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0935 ps=0.965 w=0.64 l=0.15
X574 VDD.t613 a_12030_3213# a_11942_3605# VDD.t612 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X575 a_4591_4478# a_4454_4086# a_4155_4086# VDD.t516 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X576 a_4154_2340# a_4452_2640# a_4388_2732# VDD.t102 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0924 ps=0.86 w=0.42 l=0.15
X577 VDD.t339 D[1].t2 a_10628_3239# VDD.t338 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X578 a_9954_4478# a_9442_4086# VDD.t166 VDD.t165 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X579 VDD.t27 a_10681_4086# check[2].t1 VDD.t26 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X580 a_8896_2648# a_8696_2366# VDD.t31 VDD.t30 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X581 VDD.t186 a_11249_3213# a_11159_3605# VDD.t185 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X582 VDD.t63 a_4074_4775# a_3984_5167# VDD.t62 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X583 a_11762_4801# a_11250_4775# VSS.t162 VSS.t161 sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X584 a_9322_3521# a_8857_3213# VDD.t550 VDD.t549 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X585 a_9172_2366# a_8383_2340# VSS.t375 VSS.t374 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0588 ps=0.7 w=0.42 l=0.15
X586 a_9465_4801# a_8237_4801# a_9323_5083# VDD.t535 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X587 VSS.t324 a_4854_3213# a_5561_3239# VSS.t323 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X588 VDD.t92 a_9639_4775# a_9551_5167# VDD.t91 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X589 a_6011_4801# a_5845_4801# VSS.t367 VSS.t366 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X590 VDD.t414 x4.X.t57 a_9152_4775# VDD.t413 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X591 VSS.t131 check[1].t4 a_7764_4112# VSS.t130 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X592 D[0].t1 a_7953_3239# VSS.t621 VSS.t620 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X593 VSS.t389 x4.X.t58 a_11544_4775# VSS.t388 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X594 VSS.t448 a_11630_4086# a_11629_4386# VSS.t447 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X595 a_1520_2366# x4.X.t59 VSS.t629 VSS.t628 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X596 VDD.t656 clk_sar.t0 a_1062_5674# VDD.t655 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X597 x5.X.t0 a_1338_5674# VSS.t607 VSS.t606 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X598 a_7186_4112# a_7318_4296# a_7050_4086# VSS.t365 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0864 ps=0.91 w=0.64 l=0.15
X599 a_10156_4112# a_9238_4086# a_9710_4296# VSS.t578 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X600 VDD.t515 a_11544_4775# a_12265_5083# VDD.t514 sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X601 a_3618_3239# a_3452_3239# VDD.t198 VDD.t197 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X602 VDD.t597 a_5992_4086# x45.Q_N VDD.t596 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X603 a_8683_3605# a_8236_3239# a_8590_3239# VSS.t254 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X604 VDD.t220 VDD.t218 a_3600_4086# VDD.t219 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.123 ps=1.17 w=0.42 l=0.15
X605 a_11249_3213# a_11075_3605# a_11389_3239# VSS.t86 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X606 x72.Q_N a_7246_3213# VDD.t135 VDD.t134 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X607 VSS.t525 a_8857_3213# a_8791_3239# VSS.t524 sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X608 VDD.t540 a_1682_4775# a_1592_5167# VDD.t539 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X609 x3.A a_621_4112# VDD.t696 VDD.t695 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X610 a_6780_2366# a_5991_2340# VSS.t50 VSS.t49 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0588 ps=0.7 w=0.42 l=0.15
X611 VSS.t667 a_2265_2340# a_2200_2366# VSS.t666 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0935 ps=0.965 w=0.64 l=0.15
X612 a_4074_4775# a_3900_5167# a_4214_4801# VSS.t251 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X613 VSS.t316 D[1].t3 a_10628_3239# VSS.t315 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X614 VSS.t278 x4.A a_1511_4112# VSS.t277 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X615 a_4454_4086# x5.X.t15 VSS.t416 VSS.t415 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X616 VSS.t341 a_7247_4775# a_7954_4801# VSS.t340 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X617 a_6547_4086# a_6845_4386# a_6781_4478# VDD.t571 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0924 ps=0.86 w=0.42 l=0.15
X618 a_10681_4086# a_10776_4086# VDD.t77 VDD.t76 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X619 a_11943_5167# a_10795_4801# a_11857_4801# VDD.t87 sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X620 a_11088_2366# x4.X.t60 VSS.t631 VSS.t630 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X621 a_9872_3521# a_9464_3239# a_9638_3213# VDD.t84 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X622 a_3876_6040# sel_bit[0].t1 a_3373_5674# VDD.t671 sky130_fd_pr__pfet_01v8_hvt ad=0.0974 pd=0.97 as=0.0567 ps=0.69 w=0.42 l=0.15
X623 a_11565_4478# a_10776_4086# VDD.t75 VDD.t74 sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0819 ps=0.81 w=0.42 l=0.15
X624 VDD.t487 a_1511_4112# x4.X.t19 VDD.t486 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X625 a_4794_4112# a_4926_4296# a_4658_4086# VSS.t601 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0864 ps=0.91 w=0.64 l=0.15
X626 a_4855_4775# a_4681_4801# a_4971_4801# VSS.t134 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X627 a_9574_4801# a_8237_4801# a_9465_4801# VSS.t510 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X628 a_8384_4086# a_8697_4112# a_8803_4112# VSS.t115 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X629 a_11767_4478# a_11630_4086# a_11331_4086# VDD.t468 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X630 VDD.t660 a_12031_4775# a_11943_5167# VDD.t659 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X631 x36.Q_N a_12031_4775# VSS.t611 VSS.t610 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X632 D[2].t1 a_12737_3239# VDD.t611 VDD.t610 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X633 a_9323_5083# a_8858_4775# VDD.t428 VDD.t427 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X634 VSS.t299 check[2].t4 a_10156_4112# VSS.t298 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X635 VDD.t56 a_5991_2340# x57.Q_N VDD.t55 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X636 a_8767_3605# a_8236_3239# a_8683_3605# VDD.t267 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X637 a_3618_3239# a_3452_3239# VSS.t205 VSS.t204 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X638 a_2194_4801# a_1682_4775# VSS.t515 VSS.t514 sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X639 a_1682_4775# a_1508_5167# a_1822_4801# VSS.t123 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X640 VDD.t364 a_7247_4775# a_7954_4801# VDD.t363 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X641 VSS.t464 a_1511_4112# x4.X.t5 VSS.t463 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X642 a_5169_2732# a_4657_2340# VDD.t9 VDD.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X643 a_6465_3213# x45.Q_N VDD.t82 VDD.t81 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X644 VSS.t635 a_4855_4775# a_5562_4801# VSS.t634 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X645 a_10681_4086# a_10776_4086# VSS.t76 VSS.t75 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X646 a_1616_4801# a_1227_4801# a_1508_5167# VSS.t663 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X647 VDD.t558 a_4367_3213# a_4317_3521# VDD.t557 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X648 VSS.t359 a_897_4112# x4.A VSS.t358 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X649 a_6505_4394# a_6305_4112# VDD.t402 VDD.t401 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X650 a_9709_2550# a_9236_2640# a_9953_2366# VSS.t646 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0671 ps=0.75 w=0.36 l=0.15
X651 a_2463_4775# a_2289_4801# a_2579_4801# VSS.t654 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X652 check[5].t0 a_7954_4801# VSS.t562 VSS.t561 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X653 VDD.t217 VDD.t215 a_10776_4086# VDD.t216 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.123 ps=1.17 w=0.42 l=0.15
X654 a_1511_4112# x4.A VDD.t295 VDD.t294 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X655 VSS.t288 a_3600_4086# x48.Q_N VSS.t287 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X656 VDD.t708 a_3599_2340# x54.Q_N VDD.t707 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X657 a_1207_2340# a_1520_2366# a_1626_2366# VSS.t642 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X658 a_8684_5167# a_8237_4801# a_8591_4801# VSS.t509 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X659 VSS.t399 a_8858_4775# a_8792_4801# VSS.t398 sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X660 VDD.t682 a_4855_4775# a_5562_4801# VDD.t681 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X661 a_6305_4112# x4.X.t61 VSS.t104 VSS.t103 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X662 a_3373_5674# sel_bit[0].t2 a_3671_5674# VSS.t623 sky130_fd_pr__nfet_01v8 ad=0.072 pd=0.76 as=0.0671 ps=0.75 w=0.36 l=0.15
X663 a_2777_2732# a_2265_2340# VDD.t720 VDD.t719 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X664 a_6291_3605# a_6010_3239# a_6198_3239# VDD.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X665 a_2883_5674# sel_bit[0].t3 a_2784_5996# VDD.t672 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.105 ps=0.995 w=0.42 l=0.15
X666 a_9873_5083# a_9465_4801# a_9639_4775# VDD.t706 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X667 VSS.t418 x5.X.t16 a_10629_4801# VSS.t417 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X668 a_11629_2340# D[2].t2 VDD.t19 VDD.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X669 VSS.t617 clk_sar.t1 a_1062_5674# VSS.t616 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X670 a_2375_5167# a_1227_4801# a_2289_4801# VDD.t715 sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X671 VDD.t593 a_1112_2340# D[7].t1 VDD.t592 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X672 x69.Q_N a_9638_3213# VSS.t37 VSS.t36 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X673 VDD.t73 a_10776_4086# x39.Q_N VDD.t72 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X674 VDD.t436 comparator_out.t12 a_5371_2366# VDD.t435 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0662 ps=0.735 w=0.42 l=0.15
X675 a_11834_4086# a_11089_4112# a_11970_4112# VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X676 x20.Q_N a_2463_4775# VSS.t198 VSS.t197 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X677 VDD.t406 x5.X.t17 a_8237_4801# VDD.t405 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X678 x3.A a_621_4112# VSS.t645 VSS.t644 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X679 VDD.t150 x33.Q_N a_9441_2340# VDD.t149 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X680 a_8768_5167# a_8237_4801# a_8684_5167# VDD.t534 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X681 a_6709_3521# a_6291_3605# a_6465_3213# VDD.t314 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X682 a_4019_4112# a_4155_4086# a_3600_4086# VSS.t179 sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0864 ps=0.91 w=0.64 l=0.15
X683 VSS.t276 x4.A a_1511_4112# VSS.t275 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X684 a_7317_2550# a_6845_2340# a_7561_2732# VDD.t354 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X685 a_6466_4775# VDD.t212 VDD.t214 VDD.t213 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X686 a_3913_4112# x4.X.t62 VSS.t106 VSS.t105 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X687 a_3619_4801# a_3453_4801# VSS.t492 VSS.t491 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X688 VSS.t537 a_8288_2340# D[4].t0 VSS.t536 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X689 VDD.t666 a_11543_3213# a_11493_3521# VDD.t665 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X690 a_4926_4296# a_4453_4386# a_5170_4112# VSS.t137 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0671 ps=0.75 w=0.36 l=0.15
X691 VSS.t577 a_9238_4086# a_9237_4386# VSS.t576 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X692 a_4789_3239# a_3452_3239# a_4680_3239# VSS.t203 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X693 VDD.t204 a_4368_4775# a_4318_5083# VDD.t203 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X694 VSS.t160 a_11250_4775# a_11184_4801# VSS.t159 sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X695 VSS.t393 a_4658_4086# a_4593_4112# VSS.t392 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0935 ps=0.965 w=0.64 l=0.15
X696 a_11629_2340# D[2].t3 VSS.t19 VSS.t18 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X697 VSS.t140 a_7246_3213# a_7181_3239# VSS.t139 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X698 VDD.t408 x5.X.t18 a_5845_4801# VDD.t407 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X699 x30.Q_N a_7247_4775# VDD.t362 VDD.t361 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X700 VDD.t700 a_7049_2340# a_6982_2732# VDD.t699 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X701 a_5371_2366# a_4453_2340# a_4925_2550# VSS.t405 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X702 a_4388_2366# a_3599_2340# VSS.t659 VSS.t658 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0588 ps=0.7 w=0.42 l=0.15
X703 VSS.t462 a_1511_4112# x4.X.t4 VSS.t461 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X704 VSS.t220 VDD.t738 a_4794_4112# VSS.t219 sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.101 ps=0.99 w=0.42 l=0.15
X705 a_8383_2340# a_8938_2340# a_8896_2648# VDD.t457 sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0882 ps=1.05 w=0.84 l=0.15
X706 a_10795_4801# a_10629_4801# VDD.t279 VDD.t278 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X707 VDD.t445 check[1].t5 a_7764_4112# VDD.t444 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0662 ps=0.735 w=0.42 l=0.15
X708 a_9442_4086# a_9710_4296# a_9656_4394# VDD.t456 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X709 a_6292_5167# a_6011_4801# a_6199_4801# VDD.t588 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X710 VSS.t355 a_5896_2340# D[5].t0 VSS.t354 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X711 eob.t6 a_2389_5648# VSS.t552 VSS.t551 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.218 ps=1.97 w=0.65 l=0.15
X712 VDD.t465 a_1976_4775# a_1926_5083# VDD.t464 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X713 a_11160_5167# a_10629_4801# a_11076_5167# VDD.t277 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X714 a_1511_4112# x4.A VDD.t293 VDD.t292 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X715 a_8288_2340# a_8383_2340# VSS.t373 VSS.t372 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X716 VSS.t322 a_4854_3213# a_4789_3239# VSS.t321 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X717 VSS.t456 a_1511_4112# x4.X.t3 VSS.t455 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X718 a_1996_2366# a_1207_2340# VSS.t306 VSS.t305 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0588 ps=0.7 w=0.42 l=0.15
X719 check[3].t1 a_12738_4801# VDD.t356 VDD.t355 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X720 a_4073_3213# x77.Y VDD.t5 VDD.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X721 a_8997_3239# a_9151_3213# a_8857_3213# VSS.t534 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X722 a_3900_5167# a_3619_4801# a_3807_4801# VDD.t524 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X723 VDD.t513 a_11544_4775# a_11494_5083# VDD.t512 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X724 a_4154_2340# a_4453_2340# a_4388_2366# VSS.t404 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.066 ps=0.745 w=0.36 l=0.15
X725 VSS.t351 x3.A a_897_4112# VSS.t350 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X726 VDD.t353 a_6845_2340# a_6844_2640# VDD.t352 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X727 x33.Q_N a_9639_4775# VDD.t90 VDD.t89 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X728 a_9441_2340# a_9709_2550# a_9655_2648# VDD.t528 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X729 VDD.t368 a_11834_4086# a_11767_4478# VDD.t367 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X730 a_5896_2340# a_5991_2340# VSS.t48 VSS.t47 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X731 VDD.t562 a_9151_3213# a_9872_3521# VDD.t561 sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X732 a_10775_2340# a_11330_2340# a_11288_2648# VDD.t142 sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0882 ps=1.05 w=0.84 l=0.15
X733 a_12345_2366# a_11833_2340# VSS.t335 VSS.t334 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.084 ps=0.82 w=0.42 l=0.15
X734 VDD.t318 check[2].t5 a_10156_4112# VDD.t317 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0662 ps=0.735 w=0.42 l=0.15
X735 a_9577_2366# a_9709_2550# a_9441_2340# VSS.t503 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0864 ps=0.91 w=0.64 l=0.15
X736 a_12547_2366# a_11629_2340# a_12101_2550# VSS.t438 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X737 VSS.t339 a_7247_4775# a_7182_4801# VSS.t338 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X738 a_9172_2732# a_8383_2340# VDD.t396 VDD.t395 sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0819 ps=0.81 w=0.42 l=0.15
X739 VSS.t218 VDD.t739 a_11970_4112# VSS.t217 sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.101 ps=0.99 w=0.42 l=0.15
X740 a_9374_2732# a_9237_2340# a_8938_2340# VDD.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X741 VDD.t473 x4.X.t63 a_9151_3213# VDD.t472 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X742 a_1227_4801# a_1061_4801# VDD.t23 VDD.t22 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X743 x4.X.t18 a_1511_4112# VDD.t485 VDD.t484 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X744 VDD.t431 a_4453_2340# a_4452_2640# VDD.t430 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X745 a_2389_5648# sel_bit[1].t3 a_2883_5674# VDD.t61 sky130_fd_pr__pfet_01v8_hvt ad=0.0729 pd=0.81 as=0.14 ps=1.6 w=0.54 l=0.15
X746 VDD.t579 a_2389_5648# eob.t0 VDD.t578 sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X747 x27.D a_3170_4801# VSS.t212 VSS.t211 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X748 VSS.t329 a_6845_2340# a_6844_2640# VSS.t328 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X749 a_7362_3239# x45.Q_N VSS.t83 VSS.t82 sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X750 a_7263_2648# a_6304_2366# VDD.t320 VDD.t319 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X751 a_7362_3239# a_6759_3213# a_7246_3213# VSS.t270 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X752 VSS.t460 a_1511_4112# x4.X.t2 VSS.t459 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X753 a_5992_4086# a_6547_4086# a_6505_4394# VDD.t323 sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0882 ps=1.05 w=0.84 l=0.15
X754 VDD.t548 a_8857_3213# a_8767_3605# VDD.t547 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X755 a_4213_3239# x77.Y VSS.t5 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X756 VSS.t633 a_4855_4775# a_4790_4801# VSS.t632 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X757 a_6780_2732# a_5991_2340# VDD.t54 VDD.t53 sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0819 ps=0.81 w=0.42 l=0.15
X758 a_5372_4112# a_4453_4386# a_4926_4296# VDD.t130 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X759 VDD.t148 x33.Q_N a_8383_2340# VDD.t147 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.123 ps=1.17 w=0.42 l=0.15
X760 a_11833_2340# a_12101_2550# a_12047_2648# VDD.t202 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X761 a_6982_2732# a_6845_2340# a_6546_2340# VDD.t351 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X762 a_4925_2550# a_4453_2340# a_5169_2732# VDD.t429 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X763 a_11330_2340# a_11629_2340# a_11564_2366# VSS.t437 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.066 ps=0.745 w=0.36 l=0.15
X764 VSS.t409 comparator_out.t13 a_12547_2366# VSS.t408 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X765 VDD.t410 x5.A a_1338_5674# VDD.t409 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X766 VDD.t475 x4.X.t64 a_6760_4775# VDD.t474 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X767 a_8998_4801# a_9152_4775# a_8858_4775# VSS.t451 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X768 a_10155_2366# a_9236_2640# a_9709_2550# VDD.t697 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X769 a_7562_4112# a_7050_4086# VSS.t547 VSS.t546 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.084 ps=0.82 w=0.42 l=0.15
X770 VDD.t477 a_9152_4775# a_9873_5083# VDD.t476 sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X771 VSS.t458 a_1511_4112# x4.X.t1 VSS.t457 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X772 a_7764_4112# a_6846_4086# a_7318_4296# VSS.t110 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X773 VSS.t403 a_4453_2340# a_4452_2640# VSS.t402 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X774 a_6304_2366# x4.X.t65 VDD.t627 VDD.t626 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.154 ps=1.34 w=0.64 l=0.15
X775 a_9369_3239# a_8857_3213# VSS.t523 VSS.t522 sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X776 a_4970_3239# x77.Y VSS.t3 VSS.t2 sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X777 a_4871_2648# a_3912_2366# VDD.t639 VDD.t638 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X778 VSS.t385 x5.A a_1338_5674# VSS.t384 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X779 VSS.t357 a_897_4112# x4.A VSS.t356 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X780 a_8939_4086# a_9238_4086# a_9173_4112# VSS.t575 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.066 ps=0.745 w=0.36 l=0.15
X781 a_8590_3239# comparator_out.t14 VSS.t381 VSS.t380 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X782 VDD.t133 a_7246_3213# a_7953_3239# VDD.t132 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X783 VDD.t648 x30.Q_N a_5991_2340# VDD.t647 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.123 ps=1.17 w=0.42 l=0.15
X784 a_2533_2550# a_2061_2340# a_2777_2732# VDD.t721 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X785 a_1682_4775# x4.X.t66 VDD.t629 VDD.t628 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X786 VDD.t623 x5.X.t19 a_3453_4801# VDD.t622 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X787 VDD.t211 VDD.t209 a_4658_4086# VDD.t210 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X788 a_7050_4086# a_7318_4296# a_7264_4394# VDD.t388 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X789 x4.X.t17 a_1511_4112# VDD.t483 VDD.t482 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X790 a_2200_2366# a_2060_2640# a_1762_2340# VSS.t169 sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.0711 ps=0.755 w=0.36 l=0.15
X791 a_2853_5648# sel_bit[0].t4 VDD.t704 VDD.t703 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X792 a_2853_5648# sel_bit[0].t5 VSS.t653 VSS.t652 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X793 a_8696_2366# x4.X.t67 VSS.t414 VSS.t413 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X794 a_6606_4801# a_6760_4775# a_6466_4775# VSS.t102 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X795 VSS.t454 a_1511_4112# x4.X.t0 VSS.t453 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X796 VSS.t129 a_3504_2340# D[6].t0 VSS.t128 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X797 a_11630_4086# x5.X.t20 VDD.t625 VDD.t624 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X798 a_3912_2366# x4.X.t68 VDD.t441 VDD.t440 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.154 ps=1.34 w=0.64 l=0.15
X799 a_6977_3239# a_6465_3213# VSS.t505 VSS.t504 sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X800 a_6846_4086# x5.X.t21 VSS.t72 VSS.t71 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X801 a_11389_3239# x39.Q_N VSS.t318 VSS.t317 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X802 VDD.t426 a_8858_4775# a_8768_5167# VDD.t425 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X803 a_7363_4801# VDD.t740 VSS.t216 VSS.t215 sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X804 a_8939_4086# a_9237_4386# a_9173_4478# VDD.t371 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0924 ps=0.86 w=0.42 l=0.15
X805 a_7363_4801# a_6760_4775# a_7247_4775# VSS.t101 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X806 a_6547_4086# a_6846_4086# a_6781_4112# VSS.t109 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.066 ps=0.745 w=0.36 l=0.15
X807 a_9464_3239# a_8402_3239# a_9369_3239# VSS.t42 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X808 VDD.t345 a_4854_3213# a_5561_3239# VDD.t344 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X809 a_4214_4801# VDD.t741 VSS.t214 VSS.t213 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X810 x4.X.t16 a_1511_4112# VDD.t481 VDD.t480 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X811 a_4658_4086# a_4926_4296# a_4872_4394# VDD.t642 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X812 a_8697_4112# x4.X.t69 VDD.t587 VDD.t586 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.154 ps=1.34 w=0.64 l=0.15
X813 VSS.t383 comparator_out.t15 a_2979_2366# VSS.t382 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X814 VDD.t718 a_2265_2340# a_2198_2732# VDD.t717 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X815 a_1508_5167# a_1227_4801# a_1415_4801# VDD.t714 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X816 a_6410_2366# a_6546_2340# a_5991_2340# VSS.t665 sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0864 ps=0.91 w=0.64 l=0.15
X817 VSS.t27 a_10681_4086# check[2].t0 VSS.t26 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X818 a_7317_2550# a_6844_2640# a_7561_2366# VSS.t593 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0671 ps=0.75 w=0.36 l=0.15
X819 a_3504_2340# a_3599_2340# VSS.t657 VSS.t656 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X820 a_11183_3239# a_10794_3239# a_11075_3605# VSS.t32 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X821 a_7246_3213# x45.Q_N VDD.t80 VDD.t79 sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
R0 D[3].n8 D[3].t2 269.921
R1 D[3].n8 D[3].t3 234.573
R2 D[3].n7 D[3].t0 207.373
R3 D[3].n9 D[3].n8 76.0005
R4 D[3].n14 D[3].t1 34.8148
R5 D[3].n11 D[3] 26.5622
R6 D[3].n12 D[3].n11 19.8539
R7 D[3].n11 D[3].n10 14.6672
R8 D[3] D[3].n7 9.01934
R9 D[3] D[3].n14 8.8299
R10 D[3].n9 D[3] 7.57233
R11 D[3].n7 D[3] 7.45876
R12 D[3].n13 D[3].n12 3.14374
R13 D[3].n12 D[3].n6 2.74043
R14 D[3].n10 D[3].n9 2.70473
R15 D[3].n3 D[3] 2.62982
R16 D[3].n5 D[3].n1 2.26284
R17 D[3].n4 D[3].n3 2.23869
R18 D[3].n10 D[3] 1.9836
R19 D[3].n14 D[3].n13 0.412636
R20 D[3].n6 D[3].n0 0.0232273
R21 D[3].n4 D[3].n2 0.00807576
R22 D[3].n5 D[3].n4 0.00195195
R23 D[3].n6 D[3].n5 0.00194159
R24 VDD.n2087 VDD.n1996 1858.01
R25 VDD.n1416 VDD.t692 500.865
R26 VDD.n1454 VDD.t641 500.865
R27 VDD.n1497 VDD.t322 500.865
R28 VDD.n1535 VDD.t31 500.865
R29 VDD.n1578 VDD.t422 500.865
R30 VDD.n856 VDD.t560 500.865
R31 VDD.n1152 VDD.t288 500.865
R32 VDD.n932 VDD.t562 500.865
R33 VDD.n994 VDD.t668 500.865
R34 VDD.n220 VDD.t1 500.865
R35 VDD.n185 VDD.t111 500.865
R36 VDD.n150 VDD.t402 500.865
R37 VDD.n115 VDD.t141 500.865
R38 VDD.n2193 VDD.t467 500.865
R39 VDD.n2327 VDD.t206 500.865
R40 VDD.n2451 VDD.t101 500.865
R41 VDD.n2575 VDD.t477 500.865
R42 VDD.n2631 VDD.t515 500.865
R43 VDD.n1413 VDD.n1412 440.25
R44 VDD.n1452 VDD.n1451 440.25
R45 VDD.n1494 VDD.n1493 440.25
R46 VDD.n1533 VDD.n1532 440.25
R47 VDD.n1575 VDD.n1574 440.25
R48 VDD.n1227 VDD.n1226 440.25
R49 VDD.n895 VDD.n894 440.25
R50 VDD.n1069 VDD.n1068 440.25
R51 VDD.n971 VDD.n970 440.25
R52 VDD.n218 VDD.n217 440.25
R53 VDD.n183 VDD.n182 440.25
R54 VDD.n148 VDD.n147 440.25
R55 VDD.n113 VDD.n112 440.25
R56 VDD.n2205 VDD.n2204 440.25
R57 VDD.n2337 VDD.n2336 440.25
R58 VDD.n2461 VDD.n2460 440.25
R59 VDD.n2585 VDD.n2584 440.25
R60 VDD.n2622 VDD.n2621 440.25
R61 VDD.n288 VDD.t242 397.163
R62 VDD.n377 VDD.t245 397.163
R63 VDD.n466 VDD.t224 397.163
R64 VDD.n555 VDD.t209 397.163
R65 VDD.t230 VDD.n2688 397.144
R66 VDD.t233 VDD.n2524 397.144
R67 VDD.t212 VDD.n2400 397.144
R68 VDD.t248 VDD.n2276 397.144
R69 VDD.n2679 VDD.t227 394.462
R70 VDD.n2515 VDD.t221 394.462
R71 VDD.n2391 VDD.t257 394.462
R72 VDD.n2267 VDD.t251 394.462
R73 VDD.t215 VDD.n296 385.733
R74 VDD.t239 VDD.n385 385.733
R75 VDD.t236 VDD.n474 385.733
R76 VDD.t218 VDD.n563 385.733
R77 VDD.n1614 VDD.t376 374.342
R78 VDD.n1693 VDD.t680 374.342
R79 VDD.n1767 VDD.t678 374.342
R80 VDD.n1846 VDD.t436 374.342
R81 VDD.n1920 VDD.t118 374.342
R82 VDD.n1042 VDD.t184 374.342
R83 VDD.n1121 VDD.t116 374.342
R84 VDD.n1200 VDD.t451 374.342
R85 VDD.n520 VDD.t439 374.342
R86 VDD.n431 VDD.t445 374.342
R87 VDD.n342 VDD.t318 374.342
R88 VDD.n253 VDD.t313 374.342
R89 VDD.n2124 VDD.t595 374.342
R90 VDD.n2247 VDD.t394 374.342
R91 VDD.n2371 VDD.t674 374.342
R92 VDD.n2495 VDD.t305 374.342
R93 VDD.n2713 VDD.t416 374.342
R94 VDD.n1365 VDD.t284 373.63
R95 VDD.n2058 VDD.t447 354.697
R96 VDD.n2191 VDD.t255 326.317
R97 VDD.n2031 VDD.n2029 324.707
R98 VDD.n2035 VDD.n2029 324.707
R99 VDD.n2035 VDD.n2022 324.707
R100 VDD.n2041 VDD.n2022 324.707
R101 VDD.n2041 VDD.n2021 324.707
R102 VDD.n2046 VDD.n2021 324.707
R103 VDD.n2046 VDD.n2016 324.707
R104 VDD.n2052 VDD.n2016 324.707
R105 VDD.n2052 VDD.n2015 324.707
R106 VDD.n2056 VDD.n2015 324.707
R107 VDD.n2056 VDD.n2011 324.707
R108 VDD.n2063 VDD.n2011 324.707
R109 VDD.n2063 VDD.n2009 324.707
R110 VDD.n2068 VDD.n2009 324.707
R111 VDD.n2068 VDD.n2000 324.707
R112 VDD.n2075 VDD.n2000 324.707
R113 VDD.n2075 VDD.n1999 324.707
R114 VDD.n2079 VDD.n1999 324.707
R115 VDD.n2080 VDD.n2079 324.707
R116 VDD.n2086 VDD.n1995 324.707
R117 VDD.n2091 VDD.n1995 324.707
R118 VDD.n2091 VDD.n1992 324.707
R119 VDD.n2099 VDD.n1992 324.707
R120 VDD.n2099 VDD.n1991 324.707
R121 VDD.n2103 VDD.n1991 324.707
R122 VDD.n1607 VDD.n1605 324.707
R123 VDD.n1605 VDD.n1602 324.707
R124 VDD.n1616 VDD.n1602 324.707
R125 VDD.n1616 VDD.n1600 324.707
R126 VDD.n1621 VDD.n1600 324.707
R127 VDD.n1621 VDD.n1596 324.707
R128 VDD.n1630 VDD.n1596 324.707
R129 VDD.n1630 VDD.n1595 324.707
R130 VDD.n1634 VDD.n1595 324.707
R131 VDD.n1634 VDD.n1590 324.707
R132 VDD.n1640 VDD.n1590 324.707
R133 VDD.n1640 VDD.n1588 324.707
R134 VDD.n1643 VDD.n1588 324.707
R135 VDD.n1643 VDD.n1584 324.707
R136 VDD.n1652 VDD.n1584 324.707
R137 VDD.n1652 VDD.n1582 324.707
R138 VDD.n1657 VDD.n1582 324.707
R139 VDD.n1657 VDD.n1577 324.707
R140 VDD.n1663 VDD.n1577 324.707
R141 VDD.n1663 VDD.n1576 324.707
R142 VDD.n1667 VDD.n1576 324.707
R143 VDD.n1667 VDD.n1571 324.707
R144 VDD.n1673 VDD.n1571 324.707
R145 VDD.n1673 VDD.n1569 324.707
R146 VDD.n1678 VDD.n1569 324.707
R147 VDD.n1678 VDD.n1563 324.707
R148 VDD.n1686 VDD.n1563 324.707
R149 VDD.n1686 VDD.n1562 324.707
R150 VDD.n1691 VDD.n1562 324.707
R151 VDD.n1691 VDD.n1558 324.707
R152 VDD.n1698 VDD.n1558 324.707
R153 VDD.n1698 VDD.n1557 324.707
R154 VDD.n1702 VDD.n1557 324.707
R155 VDD.n1702 VDD.n1551 324.707
R156 VDD.n1709 VDD.n1551 324.707
R157 VDD.n1709 VDD.n1549 324.707
R158 VDD.n1713 VDD.n1549 324.707
R159 VDD.n1713 VDD.n1544 324.707
R160 VDD.n1719 VDD.n1544 324.707
R161 VDD.n1719 VDD.n1542 324.707
R162 VDD.n1723 VDD.n1542 324.707
R163 VDD.n1723 VDD.n1537 324.707
R164 VDD.n1732 VDD.n1537 324.707
R165 VDD.n1732 VDD.n1536 324.707
R166 VDD.n1737 VDD.n1536 324.707
R167 VDD.n1737 VDD.n1531 324.707
R168 VDD.n1743 VDD.n1531 324.707
R169 VDD.n1743 VDD.n1530 324.707
R170 VDD.n1748 VDD.n1530 324.707
R171 VDD.n1748 VDD.n1526 324.707
R172 VDD.n1757 VDD.n1526 324.707
R173 VDD.n1757 VDD.n1525 324.707
R174 VDD.n1761 VDD.n1525 324.707
R175 VDD.n1761 VDD.n1521 324.707
R176 VDD.n1769 VDD.n1521 324.707
R177 VDD.n1769 VDD.n1519 324.707
R178 VDD.n1774 VDD.n1519 324.707
R179 VDD.n1774 VDD.n1515 324.707
R180 VDD.n1783 VDD.n1515 324.707
R181 VDD.n1783 VDD.n1514 324.707
R182 VDD.n1787 VDD.n1514 324.707
R183 VDD.n1787 VDD.n1509 324.707
R184 VDD.n1793 VDD.n1509 324.707
R185 VDD.n1793 VDD.n1507 324.707
R186 VDD.n1796 VDD.n1507 324.707
R187 VDD.n1796 VDD.n1503 324.707
R188 VDD.n1805 VDD.n1503 324.707
R189 VDD.n1805 VDD.n1501 324.707
R190 VDD.n1810 VDD.n1501 324.707
R191 VDD.n1810 VDD.n1496 324.707
R192 VDD.n1816 VDD.n1496 324.707
R193 VDD.n1816 VDD.n1495 324.707
R194 VDD.n1820 VDD.n1495 324.707
R195 VDD.n1820 VDD.n1490 324.707
R196 VDD.n1826 VDD.n1490 324.707
R197 VDD.n1826 VDD.n1488 324.707
R198 VDD.n1831 VDD.n1488 324.707
R199 VDD.n1831 VDD.n1482 324.707
R200 VDD.n1839 VDD.n1482 324.707
R201 VDD.n1839 VDD.n1481 324.707
R202 VDD.n1844 VDD.n1481 324.707
R203 VDD.n1844 VDD.n1477 324.707
R204 VDD.n1851 VDD.n1477 324.707
R205 VDD.n1851 VDD.n1476 324.707
R206 VDD.n1855 VDD.n1476 324.707
R207 VDD.n1855 VDD.n1470 324.707
R208 VDD.n1862 VDD.n1470 324.707
R209 VDD.n1862 VDD.n1468 324.707
R210 VDD.n1866 VDD.n1468 324.707
R211 VDD.n1866 VDD.n1463 324.707
R212 VDD.n1872 VDD.n1463 324.707
R213 VDD.n1872 VDD.n1461 324.707
R214 VDD.n1876 VDD.n1461 324.707
R215 VDD.n1876 VDD.n1456 324.707
R216 VDD.n1885 VDD.n1456 324.707
R217 VDD.n1885 VDD.n1455 324.707
R218 VDD.n1890 VDD.n1455 324.707
R219 VDD.n1890 VDD.n1450 324.707
R220 VDD.n1896 VDD.n1450 324.707
R221 VDD.n1896 VDD.n1449 324.707
R222 VDD.n1901 VDD.n1449 324.707
R223 VDD.n1901 VDD.n1445 324.707
R224 VDD.n1910 VDD.n1445 324.707
R225 VDD.n1910 VDD.n1444 324.707
R226 VDD.n1914 VDD.n1444 324.707
R227 VDD.n1914 VDD.n1440 324.707
R228 VDD.n1922 VDD.n1440 324.707
R229 VDD.n1922 VDD.n1438 324.707
R230 VDD.n1927 VDD.n1438 324.707
R231 VDD.n1927 VDD.n1434 324.707
R232 VDD.n1936 VDD.n1434 324.707
R233 VDD.n1936 VDD.n1433 324.707
R234 VDD.n1940 VDD.n1433 324.707
R235 VDD.n1940 VDD.n1428 324.707
R236 VDD.n1946 VDD.n1428 324.707
R237 VDD.n1946 VDD.n1426 324.707
R238 VDD.n1949 VDD.n1426 324.707
R239 VDD.n1949 VDD.n1422 324.707
R240 VDD.n1958 VDD.n1422 324.707
R241 VDD.n1958 VDD.n1420 324.707
R242 VDD.n1963 VDD.n1420 324.707
R243 VDD.n1963 VDD.n1415 324.707
R244 VDD.n1969 VDD.n1415 324.707
R245 VDD.n1969 VDD.n1414 324.707
R246 VDD.n1973 VDD.n1414 324.707
R247 VDD.n1973 VDD.n1409 324.707
R248 VDD.n1979 VDD.n1409 324.707
R249 VDD.n1979 VDD.n1407 324.707
R250 VDD.n1982 VDD.n1407 324.707
R251 VDD.n978 VDD.n976 324.707
R252 VDD.n982 VDD.n976 324.707
R253 VDD.n982 VDD.n968 324.707
R254 VDD.n988 VDD.n968 324.707
R255 VDD.n988 VDD.n967 324.707
R256 VDD.n993 VDD.n967 324.707
R257 VDD.n993 VDD.n963 324.707
R258 VDD.n1000 VDD.n963 324.707
R259 VDD.n1000 VDD.n962 324.707
R260 VDD.n1005 VDD.n962 324.707
R261 VDD.n1005 VDD.n956 324.707
R262 VDD.n1011 VDD.n956 324.707
R263 VDD.n1011 VDD.n955 324.707
R264 VDD.n1015 VDD.n955 324.707
R265 VDD.n1015 VDD.n951 324.707
R266 VDD.n1023 VDD.n951 324.707
R267 VDD.n1023 VDD.n950 324.707
R268 VDD.n1028 VDD.n950 324.707
R269 VDD.n1028 VDD.n945 324.707
R270 VDD.n1035 VDD.n945 324.707
R271 VDD.n1035 VDD.n944 324.707
R272 VDD.n1040 VDD.n944 324.707
R273 VDD.n1040 VDD.n940 324.707
R274 VDD.n1050 VDD.n940 324.707
R275 VDD.n1050 VDD.n939 324.707
R276 VDD.n1055 VDD.n939 324.707
R277 VDD.n1055 VDD.n936 324.707
R278 VDD.n1063 VDD.n936 324.707
R279 VDD.n1063 VDD.n935 324.707
R280 VDD.n1067 VDD.n935 324.707
R281 VDD.n1067 VDD.n930 324.707
R282 VDD.n1075 VDD.n930 324.707
R283 VDD.n1075 VDD.n928 324.707
R284 VDD.n1080 VDD.n928 324.707
R285 VDD.n1080 VDD.n924 324.707
R286 VDD.n1088 VDD.n924 324.707
R287 VDD.n1088 VDD.n923 324.707
R288 VDD.n1092 VDD.n923 324.707
R289 VDD.n1092 VDD.n917 324.707
R290 VDD.n1098 VDD.n917 324.707
R291 VDD.n1098 VDD.n916 324.707
R292 VDD.n1103 VDD.n916 324.707
R293 VDD.n1103 VDD.n912 324.707
R294 VDD.n1111 VDD.n912 324.707
R295 VDD.n1111 VDD.n911 324.707
R296 VDD.n1116 VDD.n911 324.707
R297 VDD.n1116 VDD.n907 324.707
R298 VDD.n1123 VDD.n907 324.707
R299 VDD.n1123 VDD.n906 324.707
R300 VDD.n1128 VDD.n906 324.707
R301 VDD.n1128 VDD.n901 324.707
R302 VDD.n1135 VDD.n901 324.707
R303 VDD.n1135 VDD.n900 324.707
R304 VDD.n1140 VDD.n900 324.707
R305 VDD.n1140 VDD.n892 324.707
R306 VDD.n1146 VDD.n892 324.707
R307 VDD.n1146 VDD.n891 324.707
R308 VDD.n1151 VDD.n891 324.707
R309 VDD.n1151 VDD.n887 324.707
R310 VDD.n1158 VDD.n887 324.707
R311 VDD.n1158 VDD.n886 324.707
R312 VDD.n1163 VDD.n886 324.707
R313 VDD.n1163 VDD.n880 324.707
R314 VDD.n1169 VDD.n880 324.707
R315 VDD.n1169 VDD.n879 324.707
R316 VDD.n1173 VDD.n879 324.707
R317 VDD.n1173 VDD.n875 324.707
R318 VDD.n1181 VDD.n875 324.707
R319 VDD.n1181 VDD.n874 324.707
R320 VDD.n1186 VDD.n874 324.707
R321 VDD.n1186 VDD.n869 324.707
R322 VDD.n1193 VDD.n869 324.707
R323 VDD.n1193 VDD.n868 324.707
R324 VDD.n1198 VDD.n868 324.707
R325 VDD.n1198 VDD.n864 324.707
R326 VDD.n1208 VDD.n864 324.707
R327 VDD.n1208 VDD.n863 324.707
R328 VDD.n1213 VDD.n863 324.707
R329 VDD.n1213 VDD.n860 324.707
R330 VDD.n1221 VDD.n860 324.707
R331 VDD.n1221 VDD.n859 324.707
R332 VDD.n1225 VDD.n859 324.707
R333 VDD.n1225 VDD.n854 324.707
R334 VDD.n1233 VDD.n854 324.707
R335 VDD.n1233 VDD.n851 324.707
R336 VDD.n1242 VDD.n851 324.707
R337 VDD.n1396 VDD.n767 324.707
R338 VDD.n1400 VDD.n767 324.707
R339 VDD.n579 VDD.n116 324.707
R340 VDD.n579 VDD.n111 324.707
R341 VDD.n586 VDD.n111 324.707
R342 VDD.n586 VDD.n110 324.707
R343 VDD.n591 VDD.n110 324.707
R344 VDD.n591 VDD.n108 324.707
R345 VDD.n108 VDD.n103 324.707
R346 VDD.n599 VDD.n103 324.707
R347 VDD.n599 VDD.n101 324.707
R348 VDD.n604 VDD.n101 324.707
R349 VDD.n604 VDD.n95 324.707
R350 VDD.n612 VDD.n95 324.707
R351 VDD.n612 VDD.n93 324.707
R352 VDD.n618 VDD.n93 324.707
R353 VDD.n618 VDD.n94 324.707
R354 VDD.n94 VDD.n88 324.707
R355 VDD.n628 VDD.n88 324.707
R356 VDD.n628 VDD.n86 324.707
R357 VDD.n738 VDD.n22 324.707
R358 VDD.n747 VDD.n22 324.707
R359 VDD.n747 VDD.n21 324.707
R360 VDD.n752 VDD.n21 324.707
R361 VDD.n752 VDD.n17 324.707
R362 VDD.n758 VDD.n17 324.707
R363 VDD.n758 VDD.n16 324.707
R364 VDD.n762 VDD.n16 324.707
R365 VDD.n490 VDD.n151 324.707
R366 VDD.n490 VDD.n146 324.707
R367 VDD.n496 VDD.n146 324.707
R368 VDD.n496 VDD.n145 324.707
R369 VDD.n501 VDD.n145 324.707
R370 VDD.n501 VDD.n141 324.707
R371 VDD.n510 VDD.n141 324.707
R372 VDD.n510 VDD.n140 324.707
R373 VDD.n514 VDD.n140 324.707
R374 VDD.n514 VDD.n136 324.707
R375 VDD.n522 VDD.n136 324.707
R376 VDD.n522 VDD.n134 324.707
R377 VDD.n527 VDD.n134 324.707
R378 VDD.n527 VDD.n130 324.707
R379 VDD.n536 VDD.n130 324.707
R380 VDD.n536 VDD.n129 324.707
R381 VDD.n540 VDD.n129 324.707
R382 VDD.n540 VDD.n124 324.707
R383 VDD.n546 VDD.n124 324.707
R384 VDD.n546 VDD.n122 324.707
R385 VDD.n549 VDD.n122 324.707
R386 VDD.n549 VDD.n118 324.707
R387 VDD.n574 VDD.n118 324.707
R388 VDD.n401 VDD.n186 324.707
R389 VDD.n401 VDD.n181 324.707
R390 VDD.n407 VDD.n181 324.707
R391 VDD.n407 VDD.n180 324.707
R392 VDD.n412 VDD.n180 324.707
R393 VDD.n412 VDD.n176 324.707
R394 VDD.n421 VDD.n176 324.707
R395 VDD.n421 VDD.n175 324.707
R396 VDD.n425 VDD.n175 324.707
R397 VDD.n425 VDD.n171 324.707
R398 VDD.n433 VDD.n171 324.707
R399 VDD.n433 VDD.n169 324.707
R400 VDD.n438 VDD.n169 324.707
R401 VDD.n438 VDD.n165 324.707
R402 VDD.n447 VDD.n165 324.707
R403 VDD.n447 VDD.n164 324.707
R404 VDD.n451 VDD.n164 324.707
R405 VDD.n451 VDD.n159 324.707
R406 VDD.n457 VDD.n159 324.707
R407 VDD.n457 VDD.n157 324.707
R408 VDD.n460 VDD.n157 324.707
R409 VDD.n460 VDD.n153 324.707
R410 VDD.n485 VDD.n153 324.707
R411 VDD.n312 VDD.n221 324.707
R412 VDD.n312 VDD.n216 324.707
R413 VDD.n318 VDD.n216 324.707
R414 VDD.n318 VDD.n215 324.707
R415 VDD.n323 VDD.n215 324.707
R416 VDD.n323 VDD.n211 324.707
R417 VDD.n332 VDD.n211 324.707
R418 VDD.n332 VDD.n210 324.707
R419 VDD.n336 VDD.n210 324.707
R420 VDD.n336 VDD.n206 324.707
R421 VDD.n344 VDD.n206 324.707
R422 VDD.n344 VDD.n204 324.707
R423 VDD.n349 VDD.n204 324.707
R424 VDD.n349 VDD.n200 324.707
R425 VDD.n358 VDD.n200 324.707
R426 VDD.n358 VDD.n199 324.707
R427 VDD.n362 VDD.n199 324.707
R428 VDD.n362 VDD.n194 324.707
R429 VDD.n368 VDD.n194 324.707
R430 VDD.n368 VDD.n192 324.707
R431 VDD.n371 VDD.n192 324.707
R432 VDD.n371 VDD.n188 324.707
R433 VDD.n396 VDD.n188 324.707
R434 VDD.n246 VDD.n244 324.707
R435 VDD.n244 VDD.n241 324.707
R436 VDD.n255 VDD.n241 324.707
R437 VDD.n255 VDD.n239 324.707
R438 VDD.n260 VDD.n239 324.707
R439 VDD.n260 VDD.n235 324.707
R440 VDD.n269 VDD.n235 324.707
R441 VDD.n269 VDD.n234 324.707
R442 VDD.n273 VDD.n234 324.707
R443 VDD.n273 VDD.n229 324.707
R444 VDD.n279 VDD.n229 324.707
R445 VDD.n279 VDD.n227 324.707
R446 VDD.n282 VDD.n227 324.707
R447 VDD.n282 VDD.n223 324.707
R448 VDD.n307 VDD.n223 324.707
R449 VDD.n2020 VDD.n2019 315.596
R450 VDD.n1684 VDD.n1683 312.132
R451 VDD.n1763 VDD.n1523 312.132
R452 VDD.n1837 VDD.n1836 312.132
R453 VDD.n1916 VDD.n1442 312.132
R454 VDD.n1610 VDD.n1604 312.132
R455 VDD.n1048 VDD.n1047 312.132
R456 VDD.n1130 VDD.n904 312.132
R457 VDD.n1206 VDD.n1205 312.132
R458 VDD.n516 VDD.n138 312.132
R459 VDD.n427 VDD.n173 312.132
R460 VDD.n338 VDD.n208 312.132
R461 VDD.n249 VDD.n243 312.132
R462 VDD.n2115 VDD.n2108 312.132
R463 VDD.n2230 VDD.n9 312.132
R464 VDD.n2362 VDD.n5 312.132
R465 VDD.n2486 VDD.n1 312.132
R466 VDD.n2722 VDD.n2721 312.132
R467 VDD.n1380 VDD.n1378 311.387
R468 VDD.n2027 VDD.n2026 307.478
R469 VDD.n1628 VDD.n1627 307.212
R470 VDD.n1704 VDD.n1555 307.212
R471 VDD.n1781 VDD.n1780 307.212
R472 VDD.n1857 VDD.n1474 307.212
R473 VDD.n1934 VDD.n1933 307.212
R474 VDD.n1030 VDD.n948 307.212
R475 VDD.n1109 VDD.n1108 307.212
R476 VDD.n1188 VDD.n872 307.212
R477 VDD.n534 VDD.n533 307.212
R478 VDD.n445 VDD.n444 307.212
R479 VDD.n356 VDD.n355 307.212
R480 VDD.n267 VDD.n266 307.212
R481 VDD.n2142 VDD.n2138 307.212
R482 VDD.n2263 VDD.n2262 306.985
R483 VDD.n2387 VDD.n2386 306.985
R484 VDD.n2511 VDD.n2510 306.985
R485 VDD.n2696 VDD.n2695 306.985
R486 VDD.n1327 VDD.n1325 306.546
R487 VDD.n1648 VDD.n1647 305.529
R488 VDD.n1727 VDD.n1726 305.529
R489 VDD.n1801 VDD.n1800 305.529
R490 VDD.n1880 VDD.n1879 305.529
R491 VDD.n1954 VDD.n1953 305.529
R492 VDD.n960 VDD.n959 305.529
R493 VDD.n1084 VDD.n1083 305.529
R494 VDD.n884 VDD.n883 305.529
R495 VDD.n2181 VDD.n2177 305.529
R496 VDD.n2315 VDD.n2311 305.529
R497 VDD.n2439 VDD.n2435 305.529
R498 VDD.n2563 VDD.n2559 305.529
R499 VDD.n2646 VDD.n2642 305.529
R500 VDD.n571 VDD.n565 305.3
R501 VDD.n482 VDD.n476 305.3
R502 VDD.n393 VDD.n387 305.3
R503 VDD.n304 VDD.n298 305.3
R504 VDD.n1247 VDD.n1246 304.861
R505 VDD.n2198 VDD.t254 289.93
R506 VDD.n1396 VDD.n768 289.413
R507 VDD.n738 VDD.n27 289.413
R508 VDD.t216 VDD.t74 281.096
R509 VDD.t240 VDD.t174 281.096
R510 VDD.t237 VDD.t598 281.096
R511 VDD.t219 VDD.t308 281.096
R512 VDD.n2673 VDD.t231 276.317
R513 VDD.n2530 VDD.t234 276.317
R514 VDD.n2406 VDD.t213 276.317
R515 VDD.n2282 VDD.t249 276.317
R516 VDD.n1236 VDD.n844 264.707
R517 VDD.n1257 VDD.n842 264.707
R518 VDD.n1264 VDD.n834 264.707
R519 VDD.n1277 VDD.n830 264.707
R520 VDD.n1281 VDD.n823 264.707
R521 VDD.n1296 VDD.n821 264.707
R522 VDD.n1306 VDD.n816 264.707
R523 VDD.n1310 VDD.n809 264.707
R524 VDD.n1324 VDD.n807 264.707
R525 VDD.n1330 VDD.n802 264.707
R526 VDD.n1343 VDD.n798 264.707
R527 VDD.n1347 VDD.n791 264.707
R528 VDD.n1364 VDD.n788 264.707
R529 VDD.n1360 VDD.n781 264.707
R530 VDD.n1377 VDD.n779 264.707
R531 VDD.n1383 VDD.n773 264.707
R532 VDD.n646 VDD.n74 264.707
R533 VDD.n658 VDD.n72 264.707
R534 VDD.n666 VDD.n63 264.707
R535 VDD.n680 VDD.n58 264.707
R536 VDD.n684 VDD.n52 264.707
R537 VDD.n696 VDD.n50 264.707
R538 VDD.n704 VDD.n41 264.707
R539 VDD.n718 VDD.n36 264.707
R540 VDD.n722 VDD.n29 264.707
R541 VDD.t350 VDD.t216 249.863
R542 VDD.t181 VDD.t240 249.863
R543 VDD.t323 VDD.t237 249.863
R544 VDD.t171 VDD.t219 249.863
R545 VDD.n1617 VDD.n1601 242.779
R546 VDD.n1633 VDD.n1632 242.779
R547 VDD.n1641 VDD.n1589 242.779
R548 VDD.t460 VDD.n1642 242.779
R549 VDD.n1653 VDD.n1583 242.779
R550 VDD.n1665 VDD.n1664 242.779
R551 VDD.n1674 VDD.n1570 242.779
R552 VDD.n1677 VDD.n1676 242.779
R553 VDD.n1690 VDD.n1688 242.779
R554 VDD.n1710 VDD.n1550 242.779
R555 VDD.n1712 VDD.n1711 242.779
R556 VDD.t12 VDD.n1543 242.779
R557 VDD.n1722 VDD.n1720 242.779
R558 VDD.n1736 VDD.n1735 242.779
R559 VDD.n1747 VDD.n1745 242.779
R560 VDD.n1759 VDD.n1758 242.779
R561 VDD.n1770 VDD.n1520 242.779
R562 VDD.n1786 VDD.n1785 242.779
R563 VDD.n1794 VDD.n1508 242.779
R564 VDD.t351 VDD.n1795 242.779
R565 VDD.n1806 VDD.n1502 242.779
R566 VDD.n1818 VDD.n1817 242.779
R567 VDD.n1827 VDD.n1489 242.779
R568 VDD.n1830 VDD.n1829 242.779
R569 VDD.n1843 VDD.n1841 242.779
R570 VDD.n1863 VDD.n1469 242.779
R571 VDD.n1865 VDD.n1864 242.779
R572 VDD.t432 VDD.n1462 242.779
R573 VDD.n1875 VDD.n1873 242.779
R574 VDD.n1889 VDD.n1888 242.779
R575 VDD.n1900 VDD.n1898 242.779
R576 VDD.n1912 VDD.n1911 242.779
R577 VDD.n1923 VDD.n1439 242.779
R578 VDD.n1939 VDD.n1938 242.779
R579 VDD.n1947 VDD.n1427 242.779
R580 VDD.t722 VDD.n1948 242.779
R581 VDD.n1959 VDD.n1421 242.779
R582 VDD.n1971 VDD.n1970 242.779
R583 VDD.n1980 VDD.n1408 242.779
R584 VDD.n2045 VDD.n2044 241.436
R585 VDD.n2055 VDD.n2054 241.436
R586 VDD.n2064 VDD.n2010 241.436
R587 VDD.n256 VDD.n240 239.452
R588 VDD.n272 VDD.n271 239.452
R589 VDD.n280 VDD.n228 239.452
R590 VDD.t468 VDD.n281 239.452
R591 VDD.n308 VDD.n222 239.452
R592 VDD.n311 VDD.n310 239.452
R593 VDD.n322 VDD.n320 239.452
R594 VDD.n334 VDD.n333 239.452
R595 VDD.n345 VDD.n205 239.452
R596 VDD.n361 VDD.n360 239.452
R597 VDD.n369 VDD.n193 239.452
R598 VDD.t608 VDD.n370 239.452
R599 VDD.n397 VDD.n187 239.452
R600 VDD.n400 VDD.n399 239.452
R601 VDD.n411 VDD.n409 239.452
R602 VDD.n423 VDD.n422 239.452
R603 VDD.n434 VDD.n170 239.452
R604 VDD.n450 VDD.n449 239.452
R605 VDD.n458 VDD.n158 239.452
R606 VDD.t104 VDD.n459 239.452
R607 VDD.n486 VDD.n152 239.452
R608 VDD.n489 VDD.n488 239.452
R609 VDD.n500 VDD.n498 239.452
R610 VDD.n512 VDD.n511 239.452
R611 VDD.n523 VDD.n135 239.452
R612 VDD.n539 VDD.n538 239.452
R613 VDD.n547 VDD.n123 239.452
R614 VDD.t516 VDD.n548 239.452
R615 VDD.n575 VDD.n117 239.452
R616 VDD.n578 VDD.n577 239.452
R617 VDD.n590 VDD.n588 239.452
R618 VDD.n600 VDD.n102 239.452
R619 VDD.n601 VDD.n600 239.452
R620 VDD.n981 VDD.n980 237.5
R621 VDD.n992 VDD.n990 237.5
R622 VDD.n1004 VDD.n1003 237.5
R623 VDD.n1012 VDD.t335 237.5
R624 VDD.n1014 VDD.n1013 237.5
R625 VDD.n1025 VDD.n1024 237.5
R626 VDD.n1039 VDD.n1038 237.5
R627 VDD.n1065 VDD.n1064 237.5
R628 VDD.n1076 VDD.n929 237.5
R629 VDD.n1090 VDD.n1089 237.5
R630 VDD.t268 VDD.n1091 237.5
R631 VDD.n1100 VDD.n1099 237.5
R632 VDD.n1102 VDD.n1101 237.5
R633 VDD.n1125 VDD.n1124 237.5
R634 VDD.n1139 VDD.n1138 237.5
R635 VDD.n1150 VDD.n1148 237.5
R636 VDD.n1162 VDD.n1161 237.5
R637 VDD.n1170 VDD.t637 237.5
R638 VDD.n1172 VDD.n1171 237.5
R639 VDD.n1183 VDD.n1182 237.5
R640 VDD.n1197 VDD.n1196 237.5
R641 VDD.n1223 VDD.n1222 237.5
R642 VDD.n1234 VDD.n853 237.5
R643 VDD.n1398 VDD.n1397 237.5
R644 VDD.n1242 VDD.n852 232.941
R645 VDD.t85 VDD.n2042 230.94
R646 VDD.n1399 VDD.t195 229.756
R647 VDD.n634 VDD.n86 229.412
R648 VDD.n642 VDD.n81 229.412
R649 VDD.n297 VDD.t215 229.072
R650 VDD.n386 VDD.t239 229.072
R651 VDD.n475 VDD.t236 229.072
R652 VDD.n564 VDD.t218 229.072
R653 VDD.t202 VDD.t423 221.667
R654 VDD.t460 VDD.t261 221.667
R655 VDD.t32 VDD.t528 221.667
R656 VDD.t698 VDD.t12 221.667
R657 VDD.t201 VDD.t319 221.667
R658 VDD.t351 VDD.t632 221.667
R659 VDD.t638 VDD.t437 221.667
R660 VDD.t102 VDD.t432 221.667
R661 VDD.t121 VDD.t693 221.667
R662 VDD.t722 VDD.t164 221.667
R663 VDD.n2044 VDD.t52 220.442
R664 VDD.t29 VDD.t2 218.631
R665 VDD.t468 VDD.t281 218.631
R666 VDD.t456 VDD.t112 218.631
R667 VDD.t608 VDD.t371 218.631
R668 VDD.t388 VDD.t403 218.631
R669 VDD.t104 VDD.t571 218.631
R670 VDD.t642 VDD.t138 218.631
R671 VDD.t516 VDD.t131 218.631
R672 VDD.t502 VDD.t508 218.631
R673 VDD.t335 VDD.t38 216.849
R674 VDD.t665 VDD.t83 216.849
R675 VDD.t268 VDD.t51 216.849
R676 VDD.t533 VDD.t563 216.849
R677 VDD.t637 VDD.t17 216.849
R678 VDD.t285 VDD.t314 216.849
R679 VDD.t657 VDD.n2043 209.946
R680 VDD.n2055 VDD.t446 209.946
R681 VDD.t271 VDD.n1631 208.472
R682 VDD.n1701 VDD.t149 208.472
R683 VDD.t649 VDD.n1784 208.472
R684 VDD.n1854 VDD.t543 208.472
R685 VDD.t567 VDD.n1937 208.472
R686 VDD.n613 VDD.t486 208.22
R687 VDD.t484 VDD.n614 208.22
R688 VDD.n2197 VDD.t732 208.013
R689 VDD.t243 VDD.n270 205.617
R690 VDD.t246 VDD.n359 205.617
R691 VDD.t225 VDD.n448 205.617
R692 VDD.t210 VDD.n537 205.617
R693 VDD.n1027 VDD.t342 203.94
R694 VDD.n1112 VDD.t604 203.94
R695 VDD.n1185 VDD.t81 203.94
R696 VDD.n105 VDD.t489 201.19
R697 VDD.n2728 VDD 200
R698 VDD.n2 VDD 200
R699 VDD.n6 VDD 200
R700 VDD.n10 VDD 200
R701 VDD.t61 VDD.n2053 199.448
R702 VDD.n737 VDD.t379 197.809
R703 VDD.n759 VDD 197.809
R704 VDD.n2100 VDD 196.823
R705 VDD.n1054 VDD 196.196
R706 VDD.n1136 VDD 196.196
R707 VDD.n1212 VDD 196.196
R708 VDD.n1654 VDD.t159 195.279
R709 VDD.n1664 VDD.t421 195.279
R710 VDD.t395 VDD.n1721 195.279
R711 VDD.n1736 VDD.t30 195.279
R712 VDD.n1807 VDD.t53 195.279
R713 VDD.n1817 VDD.t321 195.279
R714 VDD.t711 VDD.n1874 195.279
R715 VDD.n1889 VDD.t640 195.279
R716 VDD.n1960 VDD.t330 195.279
R717 VDD.n1970 VDD.t691 195.279
R718 VDD.n695 VDD.n694 195.206
R719 VDD.n1237 VDD.n843 193.614
R720 VDD.n1256 VDD.n1255 193.614
R721 VDD.n1295 VDD.n1292 193.614
R722 VDD.n1361 VDD.n780 193.614
R723 VDD.n311 VDD.t0 192.603
R724 VDD.n400 VDD.t110 192.603
R725 VDD.n489 VDD.t401 192.603
R726 VDD.n578 VDD.t140 192.603
R727 VDD.n992 VDD.t667 191.034
R728 VDD.t612 VDD.n1002 191.034
R729 VDD.t561 VDD.n1076 191.034
R730 VDD.n1078 VDD.t42 191.034
R731 VDD.n1150 VDD.t287 191.034
R732 VDD.t136 VDD.n1160 191.034
R733 VDD.t559 VDD.n1234 191.034
R734 VDD.t300 VDD.n51 190
R735 VDD.t500 VDD.n602 187.398
R736 VDD.n617 VDD.t494 187.398
R737 VDD.n773 VDD.n772 185
R738 VDD.n1385 VDD.n773 185
R739 VDD.n1381 VDD.n1377 185
R740 VDD.n1377 VDD.n1376 185
R741 VDD.n782 VDD.n781 185
R742 VDD.n781 VDD.n780 185
R743 VDD.n1366 VDD.n1364 185
R744 VDD.n1364 VDD.n1363 185
R745 VDD.n792 VDD.n791 185
R746 VDD.n791 VDD.n790 185
R747 VDD.n1343 VDD.n1342 185
R748 VDD.n1344 VDD.n1343 185
R749 VDD.n802 VDD.n801 185
R750 VDD.n1332 VDD.n802 185
R751 VDD.n1328 VDD.n1324 185
R752 VDD.n1324 VDD.n1323 185
R753 VDD.n810 VDD.n809 185
R754 VDD.n809 VDD.n808 185
R755 VDD.n1306 VDD.n1305 185
R756 VDD.n1307 VDD.n1306 185
R757 VDD.n1296 VDD.n1295 185
R758 VDD.n824 VDD.n823 185
R759 VDD.n823 VDD.n822 185
R760 VDD.n1277 VDD.n1276 185
R761 VDD.n1278 VDD.n1277 185
R762 VDD.n834 VDD.n833 185
R763 VDD.n1266 VDD.n834 185
R764 VDD.n1258 VDD.n1257 185
R765 VDD.n1257 VDD.n1256 185
R766 VDD.n845 VDD.n844 185
R767 VDD.n844 VDD.n843 185
R768 VDD.n852 VDD.n847 185
R769 VDD.n1240 VDD.n852 185
R770 VDD.n30 VDD.n29 185
R771 VDD.n29 VDD.n28 185
R772 VDD.n718 VDD.n717 185
R773 VDD.n719 VDD.n718 185
R774 VDD.n41 VDD.n40 185
R775 VDD.n706 VDD.n41 185
R776 VDD.n697 VDD.n696 185
R777 VDD.n696 VDD.n695 185
R778 VDD.n53 VDD.n52 185
R779 VDD.n52 VDD.n51 185
R780 VDD.n680 VDD.n679 185
R781 VDD.n681 VDD.n680 185
R782 VDD.n63 VDD.n62 185
R783 VDD.n668 VDD.n63 185
R784 VDD.n659 VDD.n658 185
R785 VDD.n658 VDD.n657 185
R786 VDD.n75 VDD.n74 185
R787 VDD.n74 VDD.n73 185
R788 VDD.n642 VDD.n641 185
R789 VDD.n643 VDD.n642 185
R790 VDD.n635 VDD.n634 185
R791 VDD.n634 VDD.n633 185
R792 VDD.t292 VDD.n705 182.192
R793 VDD.n2067 VDD.t672 181.077
R794 VDD.t254 VDD.n2197 179.094
R795 VDD.t114 VDD.n808 178.125
R796 VDD.n736 VDD.t385 176.987
R797 VDD.n2008 VDD.n2007 174.595
R798 VDD.n716 VDD.n37 174.595
R799 VDD.n698 VDD.n49 174.595
R800 VDD.n678 VDD.n59 174.595
R801 VDD.n660 VDD.n71 174.595
R802 VDD.n78 VDD.n77 174.595
R803 VDD.n85 VDD.n84 174.595
R804 VDD.n626 VDD.n89 174.595
R805 VDD.n620 VDD.n619 174.595
R806 VDD.n98 VDD.n97 174.595
R807 VDD.n606 VDD.n605 174.595
R808 VDD.n1619 VDD.t359 171.529
R809 VDD.t145 VDD.n1700 171.529
R810 VDD.n1772 VDD.t701 171.529
R811 VDD.t8 VDD.n1853 171.529
R812 VDD.n1925 VDD.t719 171.529
R813 VDD.n2698 VDD.t155 171.054
R814 VDD.n2505 VDD.t425 171.054
R815 VDD.n2381 VDD.t553 171.054
R816 VDD.n2257 VDD.t62 171.054
R817 VDD.n1278 VDD.t200 170.381
R818 VDD.n1567 VDD.n1566 169.184
R819 VDD.n1752 VDD.n1751 169.184
R820 VDD.n1486 VDD.n1485 169.184
R821 VDD.n1905 VDD.n1904 169.184
R822 VDD.n1405 VDD.n1404 169.184
R823 VDD.n1059 VDD.n1058 169.184
R824 VDD.n898 VDD.n897 169.184
R825 VDD.n1217 VDD.n1216 169.184
R826 VDD.n974 VDD.n973 169.184
R827 VDD.n594 VDD.n107 169.184
R828 VDD.n505 VDD.n504 169.184
R829 VDD.n416 VDD.n415 169.184
R830 VDD.n327 VDD.n326 169.184
R831 VDD.n2220 VDD.n2216 169.184
R832 VDD.n2352 VDD.n2348 169.184
R833 VDD.n2476 VDD.n2472 169.184
R834 VDD.n2600 VDD.n2596 169.184
R835 VDD.n2609 VDD.n2605 169.184
R836 VDD.n258 VDD.t369 169.179
R837 VDD.n347 VDD.t165 169.179
R838 VDD.n436 VDD.t575 169.179
R839 VDD.n525 VDD.t417 169.179
R840 VDD.n681 VDD.t482 169.179
R841 VDD.t185 VDD.n1026 167.799
R842 VDD.n1113 VDD.t547 167.799
R843 VDD.t531 VDD.n1184 167.799
R844 VDD.n603 VDD.t488 166.576
R845 VDD.n616 VDD.t480 166.576
R846 VDD.n1592 VDD.n1591 166.542
R847 VDD.n1548 VDD.n1547 166.542
R848 VDD.n1511 VDD.n1510 166.542
R849 VDD.n1467 VDD.n1466 166.542
R850 VDD.n1430 VDD.n1429 166.542
R851 VDD.n1017 VDD.n1016 166.542
R852 VDD.n920 VDD.n919 166.542
R853 VDD.n1175 VDD.n1174 166.542
R854 VDD.n1299 VDD.n1298 166.542
R855 VDD.n126 VDD.n125 166.542
R856 VDD.n161 VDD.n160 166.542
R857 VDD.n196 VDD.n195 166.542
R858 VDD.n231 VDD.n230 166.542
R859 VDD.n2153 VDD.n2152 166.542
R860 VDD.n2287 VDD.n2286 166.542
R861 VDD.n2411 VDD.n2410 166.542
R862 VDD.n2535 VDD.n2534 166.542
R863 VDD.n2668 VDD.n2667 166.542
R864 VDD.n20 VDD.n19 166.381
R865 VDD.n2093 VDD.n2092 166.006
R866 VDD.n1989 VDD.n1988 166.006
R867 VDD.n14 VDD.n13 166.006
R868 VDD.n2077 VDD.t580 165.332
R869 VDD.t582 VDD.n1996 165.332
R870 VDD.n1333 VDD.t199 165.218
R871 VDD.n25 VDD.n24 164.453
R872 VDD.n2081 VDD.t583 163.582
R873 VDD.n707 VDD.t296 161.37
R874 VDD.n2065 VDD.t434 160.083
R875 VDD.n31 VDD.t303 159.46
R876 VDD.n1666 VDD.t315 158.333
R877 VDD.n1744 VDD.t36 158.333
R878 VDD.n1819 VDD.t626 158.333
R879 VDD.n1897 VDD.t440 158.333
R880 VDD.n1972 VDD.t442 158.333
R881 VDD.n1280 VDD.t689 157.474
R882 VDD.n1307 VDD.t557 157.474
R883 VDD.t197 VDD.n1375 157.474
R884 VDD.t128 VDD.n2066 157.459
R885 VDD.n319 VDD.t275 156.165
R886 VDD.n408 VDD.t586 156.165
R887 VDD.n497 VDD.t645 156.165
R888 VDD.n587 VDD.t555 156.165
R889 VDD.t381 VDD.n748 156.165
R890 VDD.t34 VDD.n989 154.892
R891 VDD.n1066 VDD.t472 154.892
R892 VDD.t454 VDD.n1147 154.892
R893 VDD.n1224 VDD.t526 154.892
R894 VDD.n1656 VDD.t273 153.056
R895 VDD.n1733 VDD.t147 153.056
R896 VDD.n1809 VDD.t647 153.056
R897 VDD.n1886 VDD.t545 153.056
R898 VDD.n1962 VDD.t569 153.056
R899 VDD.n766 VDD.t196 152.88
R900 VDD.n2689 VDD.t230 152.694
R901 VDD.n295 VDD.n294 152
R902 VDD.n384 VDD.n383 152
R903 VDD.n473 VDD.n472 152
R904 VDD.n562 VDD.n561 152
R905 VDD.n2525 VDD.t233 151.811
R906 VDD.n2401 VDD.t212 151.811
R907 VDD.t340 VDD.n1001 149.728
R908 VDD.n1079 VDD.t602 149.728
R909 VDD.t79 VDD.n1159 149.728
R910 VDD.n1241 VDD.t6 149.728
R911 VDD.n1266 VDD.t109 149.728
R912 VDD.n2277 VDD.t248 149.322
R913 VDD.n668 VDD.t492 148.357
R914 VDD.n739 VDD.t380 148.195
R915 VDD.n2085 VDD.t652 147.891
R916 VDD.t283 VDD.n1359 147.148
R917 VDD.n1397 VDD 147.148
R918 VDD.n2042 VDD.t433 146.962
R919 VDD.n615 VDD.t490 145.754
R920 VDD.n737 VDD 145.754
R921 VDD.t461 VDD.n1619 145.139
R922 VDD.t161 VDD.n1570 145.139
R923 VDD.n1700 VDD.t13 145.139
R924 VDD.n1745 VDD.t397 145.139
R925 VDD.t354 VDD.n1772 145.139
R926 VDD.t55 VDD.n1489 145.139
R927 VDD.n1853 VDD.t429 145.139
R928 VDD.n1898 VDD.t707 145.139
R929 VDD.t721 VDD.n1925 145.139
R930 VDD.t328 VDD.n1408 145.139
R931 VDD.n2208 VDD.t189 144.738
R932 VDD.n1346 VDD.t108 144.565
R933 VDD.n2076 VDD.t584 144.338
R934 VDD.n2078 VDD.t578 144.338
R935 VDD.t469 VDD.n258 143.151
R936 VDD.n320 VDD.t72 143.151
R937 VDD.t609 VDD.n347 143.151
R938 VDD.n409 VDD.t172 143.151
R939 VDD.t105 VDD.n436 143.151
R940 VDD.n498 VDD.t596 143.151
R941 VDD.t517 VDD.n525 143.151
R942 VDD.n588 VDD.t306 143.151
R943 VDD.t142 VDD.n1655 142.5
R944 VDD.n1734 VDD.t457 142.5
R945 VDD.t716 VDD.n1808 142.5
R946 VDD.n1887 VDD.t95 142.5
R947 VDD.t387 VDD.n1961 142.5
R948 VDD.n980 VDD.t614 141.984
R949 VDD.n1026 VDD.t334 141.984
R950 VDD.t46 VDD.n1065 141.984
R951 VDD.t267 VDD.n1113 141.984
R952 VDD.n1138 VDD.t134 141.984
R953 VDD.n1184 VDD.t636 141.984
R954 VDD.t346 VDD.n1223 141.984
R955 VDD.n309 VDD.t350 140.548
R956 VDD.n398 VDD.t181 140.548
R957 VDD.n487 VDD.t323 140.548
R958 VDD.n576 VDD.t171 140.548
R959 VDD.n721 VDD.t302 140.548
R960 VDD.n991 VDD.t577 139.403
R961 VDD.t84 VDD.n1077 139.403
R962 VDD.n1149 VDD.t182 139.403
R963 VDD.t178 VDD.n1235 139.403
R964 VDD.t462 VDD.n1601 137.222
R965 VDD.n1642 VDD.t357 137.222
R966 VDD.n1688 VDD.t14 137.222
R967 VDD.t143 VDD.n1543 137.222
R968 VDD.t352 VDD.n1520 137.222
R969 VDD.n1795 VDD.t699 137.222
R970 VDD.n1841 VDD.t430 137.222
R971 VDD.t10 VDD.n1462 137.222
R972 VDD.t723 VDD.n1439 137.222
R973 VDD.n1948 VDD.t717 137.222
R974 VDD.n1323 VDD.t4 136.821
R975 VDD.t151 VDD.n1384 136.821
R976 VDD.n2034 VDD.t59 136.464
R977 VDD.t470 VDD.n240 135.343
R978 VDD.n281 VDD.t367 135.343
R979 VDD.t606 VDD.n205 135.343
R980 VDD.n370 VDD.t167 135.343
R981 VDD.t106 VDD.n170 135.343
R982 VDD.n459 VDD.t573 135.343
R983 VDD.t518 VDD.n135 135.343
R984 VDD.n548 VDD.t419 135.343
R985 VDD.t383 VDD.n749 135.343
R986 VDD.n1982 VDD.t592 135.118
R987 VDD.n2688 VDD.t730 134.986
R988 VDD.n2524 VDD.t729 134.986
R989 VDD.n2400 VDD.t737 134.986
R990 VDD.n2276 VDD.t741 134.986
R991 VDD.n288 VDD.t739 134.966
R992 VDD.n377 VDD.t727 134.966
R993 VDD.n466 VDD.t733 134.966
R994 VDD.n555 VDD.t738 134.966
R995 VDD.n1675 VDD.t157 134.583
R996 VDD.t399 VDD.n1746 134.583
R997 VDD.n1828 VDD.t57 134.583
R998 VDD.t709 VDD.n1899 134.583
R999 VDD.n1981 VDD.t326 134.583
R1000 VDD.n2679 VDD.t731 134.484
R1001 VDD.n2515 VDD.t736 134.484
R1002 VDD.n2391 VDD.t740 134.484
R1003 VDD.n2267 VDD.t725 134.484
R1004 VDD.t187 VDD.n1012 134.239
R1005 VDD.n1038 VDD.t336 134.239
R1006 VDD.n1091 VDD.t549 134.239
R1007 VDD.t269 VDD.n1125 134.239
R1008 VDD.t529 VDD.n1170 134.239
R1009 VDD.n1196 VDD.t634 134.239
R1010 VDD.n2090 VDD.t653 133.84
R1011 VDD.n295 VDD.t735 133.5
R1012 VDD.n384 VDD.t726 133.5
R1013 VDD.n473 VDD.t728 133.5
R1014 VDD.n562 VDD.t734 133.5
R1015 VDD.t76 VDD.n321 132.74
R1016 VDD.t176 VDD.n410 132.74
R1017 VDD.t600 VDD.n499 132.74
R1018 VDD.t310 VDD.n589 132.74
R1019 VDD.t610 VDD.n978 132.363
R1020 VDD.t616 VDD.n979 131.659
R1021 VDD.n1053 VDD.t44 131.659
R1022 VDD.t132 VDD.n1137 131.659
R1023 VDD.n1211 VDD.t344 131.659
R1024 VDD.t651 VDD.n2087 128.591
R1025 VDD.n657 VDD.t504 127.534
R1026 VDD.n1618 VDD.t375 126.668
R1027 VDD.n1677 VDD.t262 126.668
R1028 VDD.t679 VDD.n1689 126.668
R1029 VDD.n1758 VDD.t565 126.668
R1030 VDD.n1771 VDD.t677 126.668
R1031 VDD.n1830 VDD.t377 126.668
R1032 VDD.t435 VDD.n1842 126.668
R1033 VDD.n1911 VDD.t125 126.668
R1034 VDD.n1924 VDD.t117 126.668
R1035 VDD.t671 VDD.n2033 125.968
R1036 VDD.t409 VDD.n2089 125.968
R1037 VDD.t20 VDD.n2100 125.968
R1038 VDD.n2102 VDD.t655 125.968
R1039 VDD.n257 VDD.t312 124.933
R1040 VDD.n333 VDD.t26 124.933
R1041 VDD.n346 VDD.t317 124.933
R1042 VDD.n422 VDD.t265 124.933
R1043 VDD.n435 VDD.t444 124.933
R1044 VDD.n511 VDD.t179 124.933
R1045 VDD.n524 VDD.t438 124.933
R1046 VDD.t119 VDD.n102 124.933
R1047 VDD.t510 VDD.n629 124.933
R1048 VDD.t373 VDD.n750 124.933
R1049 VDD.t695 VDD.n759 124.933
R1050 VDD.n761 VDD.t48 124.933
R1051 VDD.n1620 VDD.t260 124.028
R1052 VDD.n1699 VDD.t697 124.028
R1053 VDD.n1773 VDD.t633 124.028
R1054 VDD.n1852 VDD.t103 124.028
R1055 VDD.n1926 VDD.t163 124.028
R1056 VDD.t183 VDD.n1037 123.913
R1057 VDD.n1054 VDD.t458 123.913
R1058 VDD.n1114 VDD.t115 123.913
R1059 VDD.t669 VDD.n1136 123.913
R1060 VDD.t450 VDD.n1195 123.913
R1061 VDD.n1212 VDD.t122 123.913
R1062 VDD VDD.t452 123.684
R1063 VDD.t405 VDD 123.684
R1064 VDD.t407 VDD 123.684
R1065 VDD.t622 VDD 123.684
R1066 VDD.t620 VDD 123.684
R1067 VDD.n259 VDD.t282 122.329
R1068 VDD.n348 VDD.t372 122.329
R1069 VDD.n437 VDD.t572 122.329
R1070 VDD.n526 VDD.t130 122.329
R1071 VDD.n2003 VDD.n2002 121.769
R1072 VDD.t39 VDD.n1036 121.332
R1073 VDD VDD.t338 121.332
R1074 VDD.n1115 VDD.t50 121.332
R1075 VDD.t332 VDD 121.332
R1076 VDD.t16 VDD.n1194 121.332
R1077 VDD VDD.t169 121.332
R1078 VDD.t260 VDD.n1618 118.751
R1079 VDD.n1689 VDD.t697 118.751
R1080 VDD.t633 VDD.n1771 118.751
R1081 VDD.n1842 VDD.t103 118.751
R1082 VDD.t163 VDD.n1924 118.751
R1083 VDD.n2706 VDD.t88 118.421
R1084 VDD.n2497 VDD.t630 118.421
R1085 VDD.n2373 VDD.t588 118.421
R1086 VDD.n2249 VDD.t524 118.421
R1087 VDD.n2126 VDD.t714 118.421
R1088 VDD.t282 VDD.n257 117.124
R1089 VDD.t372 VDD.n346 117.124
R1090 VDD.t572 VDD.n435 117.124
R1091 VDD.t130 VDD.n524 117.124
R1092 VDD.n1037 VDD.t39 116.168
R1093 VDD.t50 VDD.n1114 116.168
R1094 VDD.n1195 VDD.t16 116.168
R1095 VDD.t18 VDD.n1606 116.112
R1096 VDD.t375 VDD.n1617 116.112
R1097 VDD.t262 VDD.n1675 116.112
R1098 VDD.n1687 VDD.t618 116.112
R1099 VDD.n1690 VDD.t679 116.112
R1100 VDD.n1746 VDD.t565 116.112
R1101 VDD.n1760 VDD.t411 116.112
R1102 VDD.t677 VDD.n1770 116.112
R1103 VDD.t377 VDD.n1828 116.112
R1104 VDD.n1840 VDD.t675 116.112
R1105 VDD.n1843 VDD.t435 116.112
R1106 VDD.n1899 VDD.t125 116.112
R1107 VDD.n1913 VDD.t40 116.112
R1108 VDD.t117 VDD.n1923 116.112
R1109 VDD.t592 VDD.n1981 116.112
R1110 VDD.n2606 VDD.t355 115.79
R1111 VDD.n2710 VDD.t415 115.79
R1112 VDD.t452 VDD.n2725 115.79
R1113 VDD.n2597 VDD.t290 115.79
R1114 VDD.n2492 VDD.t304 115.79
R1115 VDD.n2483 VDD.t405 115.79
R1116 VDD.n2473 VDD.t590 115.79
R1117 VDD.n2368 VDD.t673 115.79
R1118 VDD.n2359 VDD.t407 115.79
R1119 VDD.n2349 VDD.t96 115.79
R1120 VDD.n2244 VDD.t393 115.79
R1121 VDD.n2227 VDD.t622 115.79
R1122 VDD.n2217 VDD.t207 115.79
R1123 VDD.n2121 VDD.t594 115.79
R1124 VDD.n2112 VDD.t620 115.79
R1125 VDD.n2032 VDD.t703 115.471
R1126 VDD.n2034 VDD.t671 115.471
R1127 VDD.n2090 VDD.t409 115.471
R1128 VDD.n2101 VDD.t20 115.471
R1129 VDD.t655 VDD.n2101 115.471
R1130 VDD.t624 VDD.n245 114.522
R1131 VDD.t312 VDD.n256 114.522
R1132 VDD.n321 VDD.t26 114.522
R1133 VDD.n335 VDD.t66 114.522
R1134 VDD.t317 VDD.n345 114.522
R1135 VDD.n410 VDD.t265 114.522
R1136 VDD.n424 VDD.t70 114.522
R1137 VDD.t444 VDD.n434 114.522
R1138 VDD.n499 VDD.t179 114.522
R1139 VDD.n513 VDD.t68 114.522
R1140 VDD.t438 VDD.n523 114.522
R1141 VDD.n589 VDD.t119 114.522
R1142 VDD.n630 VDD.t510 114.522
R1143 VDD.n751 VDD.t373 114.522
R1144 VDD.n760 VDD.t695 114.522
R1145 VDD.t48 VDD.n760 114.522
R1146 VDD.n979 VDD.t610 113.588
R1147 VDD.n1039 VDD.t183 113.588
R1148 VDD.t338 VDD.n1051 113.588
R1149 VDD.t458 VDD.n1053 113.588
R1150 VDD.n1124 VDD.t115 113.588
R1151 VDD.n1127 VDD.t332 113.588
R1152 VDD.n1137 VDD.t669 113.588
R1153 VDD.n1197 VDD.t450 113.588
R1154 VDD.t169 VDD.n1209 113.588
R1155 VDD.t122 VDD.n1211 113.588
R1156 VDD.n2088 VDD.t651 112.846
R1157 VDD.t157 VDD.n1674 108.195
R1158 VDD.n1747 VDD.t399 108.195
R1159 VDD.t57 VDD.n1827 108.195
R1160 VDD.n1900 VDD.t709 108.195
R1161 VDD.t326 VDD.n1980 108.195
R1162 VDD.n2611 VDD.t663 107.895
R1163 VDD.n2592 VDD.t93 107.895
R1164 VDD.n2468 VDD.t363 107.895
R1165 VDD.n2344 VDD.t681 107.895
R1166 VDD.n2212 VDD.t193 107.895
R1167 VDD.t653 VDD.n2088 107.597
R1168 VDD.n322 VDD.t76 106.713
R1169 VDD.n411 VDD.t176 106.713
R1170 VDD.n500 VDD.t600 106.713
R1171 VDD.n590 VDD.t310 106.713
R1172 VDD.t496 VDD.n73 106.713
R1173 VDD.n981 VDD.t616 105.843
R1174 VDD.n1064 VDD.t44 105.843
R1175 VDD.n1139 VDD.t132 105.843
R1176 VDD.n1222 VDD.t344 105.843
R1177 VDD.n1606 VDD.t462 105.556
R1178 VDD.t357 VDD.n1641 105.556
R1179 VDD.t14 VDD.n1687 105.556
R1180 VDD.n1712 VDD.t143 105.556
R1181 VDD.n1760 VDD.t352 105.556
R1182 VDD.t699 VDD.n1794 105.556
R1183 VDD.t430 VDD.n1840 105.556
R1184 VDD.n1865 VDD.t10 105.556
R1185 VDD.n1913 VDD.t723 105.556
R1186 VDD.t717 VDD.n1947 105.556
R1187 VDD.n2663 VDD.t153 105.263
R1188 VDD.n2725 VDD.t278 105.263
R1189 VDD.n2540 VDD.t427 105.263
R1190 VDD.n2483 VDD.t536 105.263
R1191 VDD.n2416 VDD.t551 105.263
R1192 VDD.n2359 VDD.t389 105.263
R1193 VDD.n2292 VDD.t64 105.263
R1194 VDD.n2227 VDD.t520 105.263
R1195 VDD.n2158 VDD.t541 105.263
R1196 VDD.n2112 VDD.t22 105.263
R1197 VDD.t59 VDD.n2032 104.972
R1198 VDD.n245 VDD.t470 104.111
R1199 VDD.t367 VDD.n280 104.111
R1200 VDD.n335 VDD.t606 104.111
R1201 VDD.t167 VDD.n369 104.111
R1202 VDD.n424 VDD.t106 104.111
R1203 VDD.t573 VDD.n458 104.111
R1204 VDD.n513 VDD.t518 104.111
R1205 VDD.t419 VDD.n547 104.111
R1206 VDD.t498 VDD.n630 104.111
R1207 VDD.n751 VDD.t383 104.111
R1208 VDD.n1014 VDD.t187 103.261
R1209 VDD.n1051 VDD.t336 103.261
R1210 VDD.n1099 VDD.t549 103.261
R1211 VDD.n1127 VDD.t269 103.261
R1212 VDD.n1172 VDD.t529 103.261
R1213 VDD.n1209 VDD.t634 103.261
R1214 VDD.n1332 VDD.t687 100.68
R1215 VDD.n1656 VDD.t142 100.278
R1216 VDD.t457 VDD.n1733 100.278
R1217 VDD.n1809 VDD.t716 100.278
R1218 VDD.t95 VDD.n1886 100.278
R1219 VDD.n1962 VDD.t387 100.278
R1220 VDD.n2638 VDD.t713 100.001
R1221 VDD.n2565 VDD.t706 100.001
R1222 VDD.n2441 VDD.t289 100.001
R1223 VDD.n2317 VDD.t127 100.001
R1224 VDD.n2183 VDD.t705 100.001
R1225 VDD.n1001 VDD.t577 98.0983
R1226 VDD.n1079 VDD.t84 98.0983
R1227 VDD.n1159 VDD.t182 98.0983
R1228 VDD.n1241 VDD.t178 98.0983
R1229 VDD.n1620 VDD.t461 97.6394
R1230 VDD.n1666 VDD.t161 97.6394
R1231 VDD.t13 VDD.n1699 97.6394
R1232 VDD.t397 VDD.n1744 97.6394
R1233 VDD.n1773 VDD.t354 97.6394
R1234 VDD.n1819 VDD.t55 97.6394
R1235 VDD.t429 VDD.n1852 97.6394
R1236 VDD.t707 VDD.n1897 97.6394
R1237 VDD.n1926 VDD.t721 97.6394
R1238 VDD.n1972 VDD.t328 97.6394
R1239 VDD.n2619 VDD.t661 97.3689
R1240 VDD.n2702 VDD.t277 97.3689
R1241 VDD.n2582 VDD.t89 97.3689
R1242 VDD.n2501 VDD.t534 97.3689
R1243 VDD.n2458 VDD.t361 97.3689
R1244 VDD.n2377 VDD.t391 97.3689
R1245 VDD.n2334 VDD.t683 97.3689
R1246 VDD.n2253 VDD.t522 97.3689
R1247 VDD.n2130 VDD.t24 97.3689
R1248 VDD.n2066 VDD.t584 97.0999
R1249 VDD.t578 VDD.n2077 97.0999
R1250 VDD.n259 VDD.t469 96.3019
R1251 VDD.t72 VDD.n319 96.3019
R1252 VDD.n348 VDD.t609 96.3019
R1253 VDD.t172 VDD.n408 96.3019
R1254 VDD.n437 VDD.t105 96.3019
R1255 VDD.t596 VDD.n497 96.3019
R1256 VDD.n526 VDD.t517 96.3019
R1257 VDD.t306 VDD.n587 96.3019
R1258 VDD.n989 VDD.t614 95.5168
R1259 VDD.n1036 VDD.t334 95.5168
R1260 VDD.n1066 VDD.t46 95.5168
R1261 VDD.n1115 VDD.t267 95.5168
R1262 VDD.n1147 VDD.t134 95.5168
R1263 VDD.n1194 VDD.t636 95.5168
R1264 VDD.n1224 VDD.t346 95.5168
R1265 VDD.n2033 VDD.t433 94.4756
R1266 VDD.n629 VDD.t490 93.6991
R1267 VDD.t687 VDD.n1331 92.9353
R1268 VDD.n1388 VDD.n1387 92.5005
R1269 VDD.n775 VDD.n774 92.5005
R1270 VDD.n1374 VDD.n1373 92.5005
R1271 VDD.n1362 VDD.n789 92.5005
R1272 VDD.n1358 VDD.n1357 92.5005
R1273 VDD.n1345 VDD.n797 92.5005
R1274 VDD.n1335 VDD.n1334 92.5005
R1275 VDD.n804 VDD.n803 92.5005
R1276 VDD.n1321 VDD.n1320 92.5005
R1277 VDD.n1308 VDD.n815 92.5005
R1278 VDD.n1294 VDD.n820 92.5005
R1279 VDD.n1291 VDD.n1290 92.5005
R1280 VDD.n1279 VDD.n829 92.5005
R1281 VDD.n1269 VDD.n1268 92.5005
R1282 VDD.n836 VDD.n835 92.5005
R1283 VDD.n1254 VDD.n1253 92.5005
R1284 VDD.n1239 VDD.n1238 92.5005
R1285 VDD.n1389 VDD.n1388 92.5005
R1286 VDD.n1373 VDD.n1372 92.5005
R1287 VDD.n1357 VDD.n1356 92.5005
R1288 VDD.n797 VDD.n795 92.5005
R1289 VDD.n1336 VDD.n1335 92.5005
R1290 VDD.n1320 VDD.n1319 92.5005
R1291 VDD.n815 VDD.n813 92.5005
R1292 VDD.n1290 VDD.n1289 92.5005
R1293 VDD.n829 VDD.n827 92.5005
R1294 VDD.n1270 VDD.n1269 92.5005
R1295 VDD.n837 VDD.n836 92.5005
R1296 VDD.n1253 VDD.n1252 92.5005
R1297 VDD.n734 VDD.n733 92.5005
R1298 VDD.n720 VDD.n35 92.5005
R1299 VDD.n709 VDD.n708 92.5005
R1300 VDD.n43 VDD.n42 92.5005
R1301 VDD.n693 VDD.n692 92.5005
R1302 VDD.n682 VDD.n57 92.5005
R1303 VDD.n671 VDD.n670 92.5005
R1304 VDD.n65 VDD.n64 92.5005
R1305 VDD.n655 VDD.n654 92.5005
R1306 VDD.n644 VDD.n80 92.5005
R1307 VDD.n733 VDD.n732 92.5005
R1308 VDD.n35 VDD.n33 92.5005
R1309 VDD.n710 VDD.n709 92.5005
R1310 VDD.n44 VDD.n43 92.5005
R1311 VDD.n692 VDD.n691 92.5005
R1312 VDD.n57 VDD.n55 92.5005
R1313 VDD.n672 VDD.n671 92.5005
R1314 VDD.n66 VDD.n65 92.5005
R1315 VDD.n654 VDD.n653 92.5005
R1316 VDD.n640 VDD.n80 92.5005
R1317 VDD.n1627 VDD.t272 91.4648
R1318 VDD.n1647 VDD.t160 91.4648
R1319 VDD.n1647 VDD.t274 91.4648
R1320 VDD.n1555 VDD.t150 91.4648
R1321 VDD.n1726 VDD.t396 91.4648
R1322 VDD.n1726 VDD.t148 91.4648
R1323 VDD.n1780 VDD.t650 91.4648
R1324 VDD.n1800 VDD.t54 91.4648
R1325 VDD.n1800 VDD.t648 91.4648
R1326 VDD.n1474 VDD.t544 91.4648
R1327 VDD.n1879 VDD.t712 91.4648
R1328 VDD.n1879 VDD.t546 91.4648
R1329 VDD.n1933 VDD.t568 91.4648
R1330 VDD.n1953 VDD.t331 91.4648
R1331 VDD.n1953 VDD.t570 91.4648
R1332 VDD.n959 VDD.t341 91.4648
R1333 VDD.n959 VDD.t613 91.4648
R1334 VDD.n948 VDD.t343 91.4648
R1335 VDD.n1083 VDD.t603 91.4648
R1336 VDD.n1083 VDD.t43 91.4648
R1337 VDD.n1108 VDD.t605 91.4648
R1338 VDD.n883 VDD.t80 91.4648
R1339 VDD.n883 VDD.t137 91.4648
R1340 VDD.n872 VDD.t82 91.4648
R1341 VDD.n1246 VDD.t7 91.4648
R1342 VDD.n1246 VDD.t349 91.4648
R1343 VDD.n1325 VDD.t5 91.4648
R1344 VDD.n565 VDD.t309 91.4648
R1345 VDD.n565 VDD.t220 91.4648
R1346 VDD.n533 VDD.t211 91.4648
R1347 VDD.n476 VDD.t599 91.4648
R1348 VDD.n476 VDD.t238 91.4648
R1349 VDD.n444 VDD.t226 91.4648
R1350 VDD.n387 VDD.t175 91.4648
R1351 VDD.n387 VDD.t241 91.4648
R1352 VDD.n355 VDD.t247 91.4648
R1353 VDD.n298 VDD.t75 91.4648
R1354 VDD.n298 VDD.t217 91.4648
R1355 VDD.n266 VDD.t244 91.4648
R1356 VDD.n2138 VDD.t629 91.4648
R1357 VDD.n2177 VDD.t449 91.4648
R1358 VDD.n2177 VDD.t192 91.4648
R1359 VDD.n2262 VDD.t250 91.4648
R1360 VDD.n2311 VDD.t253 91.4648
R1361 VDD.n2311 VDD.t686 91.4648
R1362 VDD.n2386 VDD.t214 91.4648
R1363 VDD.n2435 VDD.t259 91.4648
R1364 VDD.n2435 VDD.t366 91.4648
R1365 VDD.n2510 VDD.t235 91.4648
R1366 VDD.n2559 VDD.t223 91.4648
R1367 VDD.n2559 VDD.t92 91.4648
R1368 VDD.n2695 VDD.t232 91.4648
R1369 VDD.n2642 VDD.t229 91.4648
R1370 VDD.n2642 VDD.t660 91.4648
R1371 VDD.t273 VDD.n1654 89.7227
R1372 VDD.n1721 VDD.t147 89.7227
R1373 VDD.t647 VDD.n1807 89.7227
R1374 VDD.n1874 VDD.t545 89.7227
R1375 VDD.t569 VDD.n1960 89.7227
R1376 VDD.n2643 VDD.t228 89.4742
R1377 VDD.n2560 VDD.t222 89.4742
R1378 VDD.n2436 VDD.t258 89.4742
R1379 VDD.n2312 VDD.t252 89.4742
R1380 VDD.n2178 VDD.t448 89.4742
R1381 VDD.n645 VDD.t496 88.4936
R1382 VDD.n1002 VDD.t340 87.7722
R1383 VDD.t602 VDD.n1078 87.7722
R1384 VDD.n1160 VDD.t79 87.7722
R1385 VDD.n2197 VDD 87.6875
R1386 VDD.n1627 VDD.t360 86.7743
R1387 VDD.n1591 VDD.t358 86.7743
R1388 VDD.n1555 VDD.t146 86.7743
R1389 VDD.n1547 VDD.t144 86.7743
R1390 VDD.n1780 VDD.t702 86.7743
R1391 VDD.n1510 VDD.t700 86.7743
R1392 VDD.n1474 VDD.t9 86.7743
R1393 VDD.n1466 VDD.t11 86.7743
R1394 VDD.n1933 VDD.t720 86.7743
R1395 VDD.n1429 VDD.t718 86.7743
R1396 VDD.n1016 VDD.t188 86.7743
R1397 VDD.n948 VDD.t186 86.7743
R1398 VDD.n919 VDD.t550 86.7743
R1399 VDD.n1108 VDD.t548 86.7743
R1400 VDD.n1174 VDD.t530 86.7743
R1401 VDD.n872 VDD.t532 86.7743
R1402 VDD.n1298 VDD.t690 86.7743
R1403 VDD.n1325 VDD.t688 86.7743
R1404 VDD.n533 VDD.t418 86.7743
R1405 VDD.n125 VDD.t420 86.7743
R1406 VDD.n444 VDD.t576 86.7743
R1407 VDD.n160 VDD.t574 86.7743
R1408 VDD.n355 VDD.t166 86.7743
R1409 VDD.n195 VDD.t168 86.7743
R1410 VDD.n266 VDD.t370 86.7743
R1411 VDD.n230 VDD.t368 86.7743
R1412 VDD.n2152 VDD.t542 86.7743
R1413 VDD.n2138 VDD.t540 86.7743
R1414 VDD.n2262 VDD.t63 86.7743
R1415 VDD.n2286 VDD.t65 86.7743
R1416 VDD.n2386 VDD.t554 86.7743
R1417 VDD.n2410 VDD.t552 86.7743
R1418 VDD.n2510 VDD.t426 86.7743
R1419 VDD.n2534 VDD.t428 86.7743
R1420 VDD.n2695 VDD.t156 86.7743
R1421 VDD.n2667 VDD.t154 86.7743
R1422 VDD.n643 VDD.t506 85.8909
R1423 VDD.t315 VDD.n1665 84.4449
R1424 VDD.n1735 VDD.t36 84.4449
R1425 VDD.t626 VDD.n1818 84.4449
R1426 VDD.n1888 VDD.t440 84.4449
R1427 VDD.t442 VDD.n1971 84.4449
R1428 VDD.n2625 VDD.t643 84.211
R1429 VDD.n2578 VDD.t413 84.211
R1430 VDD.n2454 VDD.t474 84.211
R1431 VDD.n2330 VDD.t324 84.211
R1432 VDD.n2067 VDD.t128 83.9784
R1433 VDD.n310 VDD.t275 83.2882
R1434 VDD.n399 VDD.t586 83.2882
R1435 VDD.n488 VDD.t645 83.2882
R1436 VDD.n577 VDD.t555 83.2882
R1437 VDD.n631 VDD.t506 83.2882
R1438 VDD.n749 VDD.t381 83.2882
R1439 VDD.n990 VDD.t34 82.6092
R1440 VDD.t472 VDD.n929 82.6092
R1441 VDD.n1148 VDD.t454 82.6092
R1442 VDD.t526 VDD.n853 82.6092
R1443 VDD.t434 VDD.n2064 81.3541
R1444 VDD VDD.t18 79.1672
R1445 VDD VDD.t618 79.1672
R1446 VDD.t411 VDD 79.1672
R1447 VDD VDD.t675 79.1672
R1448 VDD.t40 VDD 79.1672
R1449 VDD.t703 VDD 78.7298
R1450 VDD VDD.t624 78.0827
R1451 VDD.t66 VDD 78.0827
R1452 VDD.t70 VDD 78.0827
R1453 VDD.t68 VDD 78.0827
R1454 VDD.t580 VDD.n2076 76.1055
R1455 VDD.n2078 VDD.t582 76.1055
R1456 VDD.n296 VDD.n287 75.2776
R1457 VDD.n385 VDD.n376 75.2776
R1458 VDD.n474 VDD.n465 75.2776
R1459 VDD.n563 VDD.n554 75.2776
R1460 VDD.t488 VDD.n601 72.8772
R1461 VDD.t480 VDD.n615 72.8772
R1462 VDD.n1631 VDD.t359 71.2505
R1463 VDD.n1701 VDD.t145 71.2505
R1464 VDD.n1784 VDD.t701 71.2505
R1465 VDD.n1854 VDD.t8 71.2505
R1466 VDD.n1937 VDD.t719 71.2505
R1467 VDD.n2139 VDD.t539 71.0531
R1468 VDD.n270 VDD.t369 70.2745
R1469 VDD.n359 VDD.t165 70.2745
R1470 VDD.n448 VDD.t575 70.2745
R1471 VDD.n537 VDD.t417 70.2745
R1472 VDD.n1027 VDD.t185 69.7016
R1473 VDD.t547 VDD.n1112 69.7016
R1474 VDD.n1185 VDD.t531 69.7016
R1475 VDD.t504 VDD.n656 67.6717
R1476 VDD VDD.n735 67.6717
R1477 VDD.n633 VDD.t498 65.069
R1478 VDD.n1412 VDD.t443 63.1021
R1479 VDD.n1451 VDD.t441 63.1021
R1480 VDD.n1493 VDD.t627 63.1021
R1481 VDD.n1532 VDD.t37 63.1021
R1482 VDD.n1574 VDD.t316 63.1021
R1483 VDD.n1226 VDD.t527 63.1021
R1484 VDD.n894 VDD.t455 63.1021
R1485 VDD.n1068 VDD.t473 63.1021
R1486 VDD.n970 VDD.t35 63.1021
R1487 VDD.n217 VDD.t276 63.1021
R1488 VDD.n182 VDD.t587 63.1021
R1489 VDD.n147 VDD.t646 63.1021
R1490 VDD.n112 VDD.t556 63.1021
R1491 VDD.n2204 VDD.t256 63.1021
R1492 VDD.n2336 VDD.t325 63.1021
R1493 VDD.n2460 VDD.t475 63.1021
R1494 VDD.n2584 VDD.t414 63.1021
R1495 VDD.n2621 VDD.t644 63.1021
R1496 VDD.n748 VDD.t385 62.4663
R1497 VDD.n2007 VDD.t129 61.563
R1498 VDD.t672 VDD.n2065 60.3596
R1499 VDD.n634 VDD.n87 60.0005
R1500 VDD.n1566 VDD.t158 58.4849
R1501 VDD.n1751 VDD.t400 58.4849
R1502 VDD.n1485 VDD.t58 58.4849
R1503 VDD.n1904 VDD.t710 58.4849
R1504 VDD.n1404 VDD.t327 58.4849
R1505 VDD.n1058 VDD.t45 58.4849
R1506 VDD.n897 VDD.t133 58.4849
R1507 VDD.n1216 VDD.t345 58.4849
R1508 VDD.n973 VDD.t617 58.4849
R1509 VDD.n107 VDD.t311 58.4849
R1510 VDD.n504 VDD.t601 58.4849
R1511 VDD.n415 VDD.t177 58.4849
R1512 VDD.n326 VDD.t77 58.4849
R1513 VDD.n2216 VDD.t194 58.4849
R1514 VDD.n2348 VDD.t682 58.4849
R1515 VDD.n2472 VDD.t364 58.4849
R1516 VDD.n2596 VDD.t94 58.4849
R1517 VDD.n2605 VDD.t664 58.4849
R1518 VDD.n1299 VDD.n1297 57.7084
R1519 VDD.t4 VDD.n1322 56.794
R1520 VDD.n1385 VDD.t151 56.794
R1521 VDD.n2236 VDD.n2235 56.4711
R1522 VDD VDD.n2031 55.6885
R1523 VDD.n2092 VDD.t410 55.4067
R1524 VDD.t302 VDD.n28 54.658
R1525 VDD.n603 VDD.t500 52.0553
R1526 VDD.t494 VDD.n616 52.0553
R1527 VDD.t108 VDD.n790 49.0494
R1528 VDD.t159 VDD.n1653 47.5005
R1529 VDD.n1655 VDD.t421 47.5005
R1530 VDD.n1722 VDD.t395 47.5005
R1531 VDD.t30 VDD.n1734 47.5005
R1532 VDD.t53 VDD.n1806 47.5005
R1533 VDD.n1808 VDD.t321 47.5005
R1534 VDD.n1875 VDD.t711 47.5005
R1535 VDD.t640 VDD.n1887 47.5005
R1536 VDD.t330 VDD.n1959 47.5005
R1537 VDD.n1961 VDD.t691 47.5005
R1538 VDD.n2634 VDD.t514 47.3689
R1539 VDD.n2648 VDD.t659 47.3689
R1540 VDD.n2569 VDD.t476 47.3689
R1541 VDD.n2555 VDD.t91 47.3689
R1542 VDD.n2445 VDD.t100 47.3689
R1543 VDD.n2431 VDD.t365 47.3689
R1544 VDD.n2321 VDD.t205 47.3689
R1545 VDD.n2307 VDD.t685 47.3689
R1546 VDD.n2187 VDD.t466 47.3689
R1547 VDD.n2173 VDD.t191 47.3689
R1548 VDD.t74 VDD.n308 46.8498
R1549 VDD.t0 VDD.n309 46.8498
R1550 VDD.t174 VDD.n397 46.8498
R1551 VDD.t110 VDD.n398 46.8498
R1552 VDD.t598 VDD.n486 46.8498
R1553 VDD.t401 VDD.n487 46.8498
R1554 VDD.t308 VDD.n575 46.8498
R1555 VDD.t140 VDD.n576 46.8498
R1556 VDD.t492 VDD.n667 46.8498
R1557 VDD.t667 VDD.n991 46.4679
R1558 VDD.n1004 VDD.t612 46.4679
R1559 VDD.n1077 VDD.t561 46.4679
R1560 VDD.n1089 VDD.t42 46.4679
R1561 VDD.t287 VDD.n1149 46.4679
R1562 VDD.n1162 VDD.t136 46.4679
R1563 VDD.n1235 VDD.t559 46.4679
R1564 VDD.n1363 VDD.t283 46.4679
R1565 VDD.n2089 VDD 44.6138
R1566 VDD.n2102 VDD 44.6138
R1567 VDD.n633 VDD.n632 44.2471
R1568 VDD.n761 VDD 44.2471
R1569 VDD.t109 VDD.n1265 43.8864
R1570 VDD.n1399 VDD 43.8864
R1571 VDD.n2002 VDD.t581 42.3555
R1572 VDD VDD.n2727 42.1058
R1573 VDD.n2482 VDD 42.1058
R1574 VDD.n2358 VDD 42.1058
R1575 VDD.n2238 VDD.n2237 42.1058
R1576 VDD.n2226 VDD 42.1058
R1577 VDD.n2111 VDD 42.1058
R1578 VDD.n2054 VDD.t61 41.9894
R1579 VDD.t379 VDD.n736 41.6443
R1580 VDD.n750 VDD 41.6443
R1581 VDD.n2026 VDD.t704 41.5552
R1582 VDD.n2026 VDD.t60 41.5552
R1583 VDD.n2019 VDD.t86 41.5552
R1584 VDD.n2019 VDD.t658 41.5552
R1585 VDD.n1683 VDD.t619 41.5552
R1586 VDD.n1683 VDD.t15 41.5552
R1587 VDD.n1523 VDD.t412 41.5552
R1588 VDD.n1523 VDD.t353 41.5552
R1589 VDD.n1836 VDD.t676 41.5552
R1590 VDD.n1836 VDD.t431 41.5552
R1591 VDD.n1442 VDD.t41 41.5552
R1592 VDD.n1442 VDD.t724 41.5552
R1593 VDD.n1604 VDD.t19 41.5552
R1594 VDD.n1604 VDD.t463 41.5552
R1595 VDD.n1047 VDD.t337 41.5552
R1596 VDD.n1047 VDD.t339 41.5552
R1597 VDD.n904 VDD.t270 41.5552
R1598 VDD.n904 VDD.t333 41.5552
R1599 VDD.n1205 VDD.t635 41.5552
R1600 VDD.n1205 VDD.t170 41.5552
R1601 VDD.n1378 VDD.t198 41.5552
R1602 VDD.n1378 VDD.t152 41.5552
R1603 VDD.n138 VDD.t69 41.5552
R1604 VDD.n138 VDD.t519 41.5552
R1605 VDD.n173 VDD.t71 41.5552
R1606 VDD.n173 VDD.t107 41.5552
R1607 VDD.n208 VDD.t67 41.5552
R1608 VDD.n208 VDD.t607 41.5552
R1609 VDD.n243 VDD.t625 41.5552
R1610 VDD.n243 VDD.t471 41.5552
R1611 VDD.n2108 VDD.t23 41.5552
R1612 VDD.n2108 VDD.t621 41.5552
R1613 VDD.n9 VDD.t521 41.5552
R1614 VDD.n9 VDD.t623 41.5552
R1615 VDD.n5 VDD.t390 41.5552
R1616 VDD.n5 VDD.t408 41.5552
R1617 VDD.n1 VDD.t537 41.5552
R1618 VDD.n1 VDD.t406 41.5552
R1619 VDD.n2721 VDD.t279 41.5552
R1620 VDD.n2721 VDD.t453 41.5552
R1621 VDD VDD.n1052 41.3048
R1622 VDD.n1126 VDD 41.3048
R1623 VDD VDD.n1210 41.3048
R1624 VDD.n1591 VDD.t424 38.6969
R1625 VDD.n1547 VDD.t33 38.6969
R1626 VDD.n1510 VDD.t320 38.6969
R1627 VDD.n1466 VDD.t639 38.6969
R1628 VDD.n1429 VDD.t694 38.6969
R1629 VDD.n1016 VDD.t666 38.6969
R1630 VDD.n919 VDD.t564 38.6969
R1631 VDD.n1174 VDD.t286 38.6969
R1632 VDD.n1298 VDD.t558 38.6969
R1633 VDD.n125 VDD.t139 38.6969
R1634 VDD.n160 VDD.t404 38.6969
R1635 VDD.n195 VDD.t113 38.6969
R1636 VDD.n230 VDD.t3 38.6969
R1637 VDD.n2152 VDD.t465 38.6969
R1638 VDD.n2286 VDD.t204 38.6969
R1639 VDD.n2410 VDD.t99 38.6969
R1640 VDD.n2534 VDD.t479 38.6969
R1641 VDD.n2667 VDD.t513 38.6969
R1642 VDD.n1988 VDD.t21 36.1587
R1643 VDD.n1988 VDD.t656 36.1587
R1644 VDD.n13 VDD.t696 36.1587
R1645 VDD.n13 VDD.t49 36.1587
R1646 VDD.t689 VDD.n822 36.1418
R1647 VDD.n1293 VDD.t557 36.1418
R1648 VDD.n1376 VDD.t197 36.1418
R1649 VDD.n1253 VDD.n842 35.2946
R1650 VDD.n1264 VDD.n836 35.2946
R1651 VDD.n1269 VDD.n830 35.2946
R1652 VDD.n1281 VDD.n829 35.2946
R1653 VDD.n1290 VDD.n821 35.2946
R1654 VDD.n820 VDD.n816 35.2946
R1655 VDD.n1310 VDD.n815 35.2946
R1656 VDD.n1320 VDD.n807 35.2946
R1657 VDD.n1335 VDD.n798 35.2946
R1658 VDD.n1347 VDD.n797 35.2946
R1659 VDD.n1357 VDD.n788 35.2946
R1660 VDD.n1373 VDD.n779 35.2946
R1661 VDD.n1388 VDD.n768 35.2946
R1662 VDD.n87 VDD.n81 35.2946
R1663 VDD.n646 VDD.n80 35.2946
R1664 VDD.n654 VDD.n72 35.2946
R1665 VDD.n666 VDD.n65 35.2946
R1666 VDD.n671 VDD.n58 35.2946
R1667 VDD.n684 VDD.n57 35.2946
R1668 VDD.n692 VDD.n50 35.2946
R1669 VDD.n704 VDD.n43 35.2946
R1670 VDD.n709 VDD.n36 35.2946
R1671 VDD.n722 VDD.n35 35.2946
R1672 VDD.n733 VDD.n27 35.2946
R1673 VDD.n1632 VDD.t271 34.3061
R1674 VDD.t149 VDD.n1550 34.3061
R1675 VDD.n1785 VDD.t649 34.3061
R1676 VDD.t543 VDD.n1469 34.3061
R1677 VDD.n1938 VDD.t567 34.3061
R1678 VDD.n2144 VDD.t628 34.211
R1679 VDD.n2092 VDD.t654 34.0906
R1680 VDD.n271 VDD.t243 33.8361
R1681 VDD.n360 VDD.t246 33.8361
R1682 VDD.n449 VDD.t225 33.8361
R1683 VDD.n538 VDD.t210 33.8361
R1684 VDD.n719 VDD.t296 33.8361
R1685 VDD.t342 VDD.n1025 33.5603
R1686 VDD.n1101 VDD.t604 33.5603
R1687 VDD.t81 VDD.n1183 33.5603
R1688 VDD.n1566 VDD.t263 31.831
R1689 VDD.n1751 VDD.t566 31.831
R1690 VDD.n1485 VDD.t378 31.831
R1691 VDD.n1904 VDD.t126 31.831
R1692 VDD.n1404 VDD.t593 31.831
R1693 VDD.n1058 VDD.t459 31.831
R1694 VDD.n897 VDD.t670 31.831
R1695 VDD.n1216 VDD.t123 31.831
R1696 VDD.n973 VDD.t611 31.831
R1697 VDD.n107 VDD.t120 31.831
R1698 VDD.n504 VDD.t180 31.831
R1699 VDD.n415 VDD.t266 31.831
R1700 VDD.n326 VDD.t27 31.831
R1701 VDD.n2216 VDD.t208 31.831
R1702 VDD.n2348 VDD.t97 31.831
R1703 VDD.n2472 VDD.t591 31.831
R1704 VDD.n2596 VDD.t291 31.831
R1705 VDD.n2605 VDD.t356 31.831
R1706 VDD.n2045 VDD.t657 31.4922
R1707 VDD.t446 VDD.n2010 31.4922
R1708 VDD.n602 VDD.t486 31.2334
R1709 VDD.n617 VDD.t484 31.2334
R1710 VDD.n2007 VDD.t585 30.5947
R1711 VDD.n1344 VDD.t199 28.3972
R1712 VDD.n1412 VDD.t329 28.0332
R1713 VDD.n1451 VDD.t708 28.0332
R1714 VDD.n1493 VDD.t56 28.0332
R1715 VDD.n1532 VDD.t398 28.0332
R1716 VDD.n1574 VDD.t162 28.0332
R1717 VDD.n1226 VDD.t347 28.0332
R1718 VDD.n894 VDD.t135 28.0332
R1719 VDD.n1068 VDD.t47 28.0332
R1720 VDD.n970 VDD.t615 28.0332
R1721 VDD.n217 VDD.t73 28.0332
R1722 VDD.n182 VDD.t173 28.0332
R1723 VDD.n147 VDD.t597 28.0332
R1724 VDD.n112 VDD.t307 28.0332
R1725 VDD.n2204 VDD.t190 28.0332
R1726 VDD.n2336 VDD.t684 28.0332
R1727 VDD.n2460 VDD.t362 28.0332
R1728 VDD.n2584 VDD.t90 28.0332
R1729 VDD.n2621 VDD.t662 28.0332
R1730 VDD.n2002 VDD.t579 26.5955
R1731 VDD.n37 VDD.t293 26.5955
R1732 VDD.n37 VDD.t297 26.5955
R1733 VDD.n49 VDD.t295 26.5955
R1734 VDD.n49 VDD.t299 26.5955
R1735 VDD.n59 VDD.t483 26.5955
R1736 VDD.n59 VDD.t301 26.5955
R1737 VDD.n71 VDD.t505 26.5955
R1738 VDD.n71 VDD.t493 26.5955
R1739 VDD.n77 VDD.t507 26.5955
R1740 VDD.n77 VDD.t497 26.5955
R1741 VDD.n84 VDD.t511 26.5955
R1742 VDD.n84 VDD.t499 26.5955
R1743 VDD.n89 VDD.t481 26.5955
R1744 VDD.n89 VDD.t491 26.5955
R1745 VDD.n619 VDD.t485 26.5955
R1746 VDD.n619 VDD.t495 26.5955
R1747 VDD.n97 VDD.t509 26.5955
R1748 VDD.n97 VDD.t503 26.5955
R1749 VDD.n605 VDD.t501 26.5955
R1750 VDD.n605 VDD.t487 26.5955
R1751 VDD.n24 VDD.t386 26.5955
R1752 VDD.n24 VDD.t382 26.5955
R1753 VDD.n19 VDD.t384 26.5955
R1754 VDD.n19 VDD.t374 26.5955
R1755 VDD.n632 VDD.n631 26.0279
R1756 VDD.n645 VDD.n644 26.0279
R1757 VDD.n656 VDD.n655 26.0279
R1758 VDD.n667 VDD.n64 26.0279
R1759 VDD.n670 VDD.n669 26.0279
R1760 VDD.n669 VDD.t482 26.0279
R1761 VDD.n683 VDD.n682 26.0279
R1762 VDD.n705 VDD.n42 26.0279
R1763 VDD.n708 VDD.n707 26.0279
R1764 VDD.n721 VDD.n720 26.0279
R1765 VDD.n735 VDD.n734 26.0279
R1766 VDD.n1239 VDD.n1237 25.8157
R1767 VDD.n1265 VDD.n835 25.8157
R1768 VDD.n1268 VDD.n1267 25.8157
R1769 VDD.n1280 VDD.n1279 25.8157
R1770 VDD.n1292 VDD.n1291 25.8157
R1771 VDD.n1294 VDD.n1293 25.8157
R1772 VDD.n1309 VDD.n1308 25.8157
R1773 VDD.n1322 VDD.n1321 25.8157
R1774 VDD.n1331 VDD.n803 25.8157
R1775 VDD.n1334 VDD.n1333 25.8157
R1776 VDD.n1346 VDD.n1345 25.8157
R1777 VDD.n1359 VDD.n1358 25.8157
R1778 VDD.n1362 VDD.n1361 25.8157
R1779 VDD.n1375 VDD.n1374 25.8157
R1780 VDD.n1384 VDD.n774 25.8157
R1781 VDD.n1387 VDD.n1386 25.8157
R1782 VDD.n1238 VDD.n852 24.7064
R1783 VDD.n1253 VDD.n844 24.7064
R1784 VDD.n1257 VDD.n836 24.7064
R1785 VDD.n1269 VDD.n834 24.7064
R1786 VDD.n1277 VDD.n829 24.7064
R1787 VDD.n1290 VDD.n823 24.7064
R1788 VDD.n1306 VDD.n815 24.7064
R1789 VDD.n1320 VDD.n809 24.7064
R1790 VDD.n1324 VDD.n804 24.7064
R1791 VDD.n1335 VDD.n802 24.7064
R1792 VDD.n1343 VDD.n797 24.7064
R1793 VDD.n1357 VDD.n791 24.7064
R1794 VDD.n1364 VDD.n789 24.7064
R1795 VDD.n1373 VDD.n781 24.7064
R1796 VDD.n1377 VDD.n775 24.7064
R1797 VDD.n1388 VDD.n773 24.7064
R1798 VDD.n642 VDD.n80 24.7064
R1799 VDD.n654 VDD.n74 24.7064
R1800 VDD.n658 VDD.n65 24.7064
R1801 VDD.n671 VDD.n63 24.7064
R1802 VDD.n680 VDD.n57 24.7064
R1803 VDD.n692 VDD.n52 24.7064
R1804 VDD.n696 VDD.n43 24.7064
R1805 VDD.n709 VDD.n41 24.7064
R1806 VDD.n718 VDD.n35 24.7064
R1807 VDD.n733 VDD.n29 24.7064
R1808 VDD.n1382 VDD.n775 24.0258
R1809 VDD.n789 VDD.n786 24.0139
R1810 VDD.n1238 VDD.n848 23.9985
R1811 VDD.n1329 VDD.n804 23.9985
R1812 VDD.n1255 VDD.t348 23.2342
R1813 VDD.n1267 VDD.t200 23.2342
R1814 VDD.t261 VDD.n1583 21.1116
R1815 VDD.n1720 VDD.t698 21.1116
R1816 VDD.t632 VDD.n1502 21.1116
R1817 VDD.n1873 VDD.t102 21.1116
R1818 VDD.t164 VDD.n1421 21.1116
R1819 VDD.n2652 VDD.t87 21.0531
R1820 VDD.n2551 VDD.t631 21.0531
R1821 VDD.n2427 VDD.t589 21.0531
R1822 VDD.n2303 VDD.t525 21.0531
R1823 VDD.n2169 VDD.t715 21.0531
R1824 VDD.n2053 VDD.t52 20.995
R1825 VDD.t281 VDD.n222 20.8224
R1826 VDD.t371 VDD.n187 20.8224
R1827 VDD.t571 VDD.n152 20.8224
R1828 VDD.t131 VDD.n117 20.8224
R1829 VDD.n1003 VDD.t38 20.6527
R1830 VDD.t51 VDD.n1090 20.6527
R1831 VDD.n1161 VDD.t17 20.6527
R1832 VDD.t6 VDD.n1240 20.6527
R1833 VDD.n1386 VDD 20.6527
R1834 VDD.n2036 VDD.n2023 20.3039
R1835 VDD.n2040 VDD.n2023 20.3039
R1836 VDD.n2040 VDD.n2024 20.3039
R1837 VDD.n2047 VDD.n2017 20.3039
R1838 VDD.n2051 VDD.n2017 20.3039
R1839 VDD.n2051 VDD.n2014 20.3039
R1840 VDD.n2062 VDD.n2012 20.3039
R1841 VDD.n2062 VDD.n2006 20.3039
R1842 VDD.n2069 VDD.n2006 20.3039
R1843 VDD.n2074 VDD.n2001 20.3039
R1844 VDD.n2074 VDD.n2004 20.3039
R1845 VDD.n2081 VDD.n1998 20.3039
R1846 VDD.n2085 VDD.n1994 20.3039
R1847 VDD.n1622 VDD.n1599 20.3039
R1848 VDD.n1622 VDD.n1597 20.3039
R1849 VDD.n1635 VDD.n1594 20.3039
R1850 VDD.n1636 VDD.n1635 20.3039
R1851 VDD.n1639 VDD.n1587 20.3039
R1852 VDD.n1644 VDD.n1587 20.3039
R1853 VDD.n1644 VDD.n1585 20.3039
R1854 VDD.n1651 VDD.n1585 20.3039
R1855 VDD.n1659 VDD.n1658 20.3039
R1856 VDD.n1672 VDD.n1572 20.3039
R1857 VDD.n1679 VDD.n1564 20.3039
R1858 VDD.n1697 VDD.n1559 20.3039
R1859 VDD.n1697 VDD.n1556 20.3039
R1860 VDD.n1708 VDD.n1552 20.3039
R1861 VDD.n1708 VDD.n1553 20.3039
R1862 VDD.n1714 VDD.n1545 20.3039
R1863 VDD.n1718 VDD.n1545 20.3039
R1864 VDD.n1718 VDD.n1541 20.3039
R1865 VDD.n1724 VDD.n1541 20.3039
R1866 VDD.n1731 VDD.n1539 20.3039
R1867 VDD.n1749 VDD.n1529 20.3039
R1868 VDD.n1756 VDD.n1524 20.3039
R1869 VDD.n1775 VDD.n1518 20.3039
R1870 VDD.n1775 VDD.n1516 20.3039
R1871 VDD.n1788 VDD.n1513 20.3039
R1872 VDD.n1789 VDD.n1788 20.3039
R1873 VDD.n1792 VDD.n1506 20.3039
R1874 VDD.n1797 VDD.n1506 20.3039
R1875 VDD.n1797 VDD.n1504 20.3039
R1876 VDD.n1804 VDD.n1504 20.3039
R1877 VDD.n1812 VDD.n1811 20.3039
R1878 VDD.n1825 VDD.n1491 20.3039
R1879 VDD.n1832 VDD.n1483 20.3039
R1880 VDD.n1850 VDD.n1478 20.3039
R1881 VDD.n1850 VDD.n1475 20.3039
R1882 VDD.n1861 VDD.n1471 20.3039
R1883 VDD.n1861 VDD.n1472 20.3039
R1884 VDD.n1867 VDD.n1464 20.3039
R1885 VDD.n1871 VDD.n1464 20.3039
R1886 VDD.n1871 VDD.n1460 20.3039
R1887 VDD.n1877 VDD.n1460 20.3039
R1888 VDD.n1884 VDD.n1458 20.3039
R1889 VDD.n1902 VDD.n1448 20.3039
R1890 VDD.n1909 VDD.n1443 20.3039
R1891 VDD.n1928 VDD.n1437 20.3039
R1892 VDD.n1928 VDD.n1435 20.3039
R1893 VDD.n1941 VDD.n1432 20.3039
R1894 VDD.n1942 VDD.n1941 20.3039
R1895 VDD.n1945 VDD.n1425 20.3039
R1896 VDD.n1950 VDD.n1425 20.3039
R1897 VDD.n1950 VDD.n1423 20.3039
R1898 VDD.n1957 VDD.n1423 20.3039
R1899 VDD.n1965 VDD.n1964 20.3039
R1900 VDD.n1978 VDD.n1410 20.3039
R1901 VDD.n983 VDD.n969 20.3039
R1902 VDD.n999 VDD.n964 20.3039
R1903 VDD.n1006 VDD.n957 20.3039
R1904 VDD.n1010 VDD.n957 20.3039
R1905 VDD.n1010 VDD.n954 20.3039
R1906 VDD.n1018 VDD.n954 20.3039
R1907 VDD.n1022 VDD.n952 20.3039
R1908 VDD.n1022 VDD.n949 20.3039
R1909 VDD.n1034 VDD.n946 20.3039
R1910 VDD.n1034 VDD.n943 20.3039
R1911 VDD.n1056 VDD.n938 20.3039
R1912 VDD.n1062 VDD.n934 20.3039
R1913 VDD.n1081 VDD.n927 20.3039
R1914 VDD.n1087 VDD.n922 20.3039
R1915 VDD.n1093 VDD.n922 20.3039
R1916 VDD.n1093 VDD.n918 20.3039
R1917 VDD.n1097 VDD.n918 20.3039
R1918 VDD.n1104 VDD.n915 20.3039
R1919 VDD.n1104 VDD.n913 20.3039
R1920 VDD.n1117 VDD.n910 20.3039
R1921 VDD.n1117 VDD.n908 20.3039
R1922 VDD.n1134 VDD.n902 20.3039
R1923 VDD.n1141 VDD.n893 20.3039
R1924 VDD.n1157 VDD.n888 20.3039
R1925 VDD.n1164 VDD.n881 20.3039
R1926 VDD.n1168 VDD.n881 20.3039
R1927 VDD.n1168 VDD.n878 20.3039
R1928 VDD.n1176 VDD.n878 20.3039
R1929 VDD.n1180 VDD.n876 20.3039
R1930 VDD.n1180 VDD.n873 20.3039
R1931 VDD.n1192 VDD.n870 20.3039
R1932 VDD.n1192 VDD.n867 20.3039
R1933 VDD.n1214 VDD.n862 20.3039
R1934 VDD.n1220 VDD.n858 20.3039
R1935 VDD.n1243 VDD.n850 20.3039
R1936 VDD.n1395 VDD.n770 20.3039
R1937 VDD.n598 VDD.n104 20.3039
R1938 VDD.n607 VDD.n100 20.3039
R1939 VDD.n611 VDD.n96 20.3039
R1940 VDD.n621 VDD.n92 20.3039
R1941 VDD.n625 VDD.n90 20.3039
R1942 VDD.n754 VDD.n753 20.3039
R1943 VDD.n592 VDD.n109 20.3039
R1944 VDD.n568 VDD.n567 20.3039
R1945 VDD.n509 VDD.n139 20.3039
R1946 VDD.n528 VDD.n133 20.3039
R1947 VDD.n528 VDD.n131 20.3039
R1948 VDD.n541 VDD.n128 20.3039
R1949 VDD.n542 VDD.n541 20.3039
R1950 VDD.n545 VDD.n121 20.3039
R1951 VDD.n550 VDD.n121 20.3039
R1952 VDD.n550 VDD.n119 20.3039
R1953 VDD.n573 VDD.n119 20.3039
R1954 VDD.n502 VDD.n144 20.3039
R1955 VDD.n479 VDD.n478 20.3039
R1956 VDD.n420 VDD.n174 20.3039
R1957 VDD.n439 VDD.n168 20.3039
R1958 VDD.n439 VDD.n166 20.3039
R1959 VDD.n452 VDD.n163 20.3039
R1960 VDD.n453 VDD.n452 20.3039
R1961 VDD.n456 VDD.n156 20.3039
R1962 VDD.n461 VDD.n156 20.3039
R1963 VDD.n461 VDD.n154 20.3039
R1964 VDD.n484 VDD.n154 20.3039
R1965 VDD.n413 VDD.n179 20.3039
R1966 VDD.n390 VDD.n389 20.3039
R1967 VDD.n331 VDD.n209 20.3039
R1968 VDD.n350 VDD.n203 20.3039
R1969 VDD.n350 VDD.n201 20.3039
R1970 VDD.n363 VDD.n198 20.3039
R1971 VDD.n364 VDD.n363 20.3039
R1972 VDD.n367 VDD.n191 20.3039
R1973 VDD.n372 VDD.n191 20.3039
R1974 VDD.n372 VDD.n189 20.3039
R1975 VDD.n395 VDD.n189 20.3039
R1976 VDD.n324 VDD.n214 20.3039
R1977 VDD.n301 VDD.n300 20.3039
R1978 VDD.n261 VDD.n238 20.3039
R1979 VDD.n261 VDD.n236 20.3039
R1980 VDD.n274 VDD.n233 20.3039
R1981 VDD.n275 VDD.n274 20.3039
R1982 VDD.n278 VDD.n226 20.3039
R1983 VDD.n283 VDD.n226 20.3039
R1984 VDD.n283 VDD.n224 20.3039
R1985 VDD.n306 VDD.n224 20.3039
R1986 VDD.n2224 VDD.n2223 20.3039
R1987 VDD.n2356 VDD.n2355 20.3039
R1988 VDD.n2480 VDD.n2479 20.3039
R1989 VDD.n2730 VDD.n2602 20.3039
R1990 VDD.n627 VDD.n85 19.8626
R1991 VDD.n2003 VDD.n1998 19.6419
R1992 VDD.n2069 VDD.n2008 19.2005
R1993 VDD.n745 VDD.n20 19.2005
R1994 VDD.n1629 VDD.n1597 18.5384
R1995 VDD.n1703 VDD.n1556 18.5384
R1996 VDD.n1782 VDD.n1516 18.5384
R1997 VDD.n1856 VDD.n1475 18.5384
R1998 VDD.n1935 VDD.n1435 18.5384
R1999 VDD.n1029 VDD.n946 18.5384
R2000 VDD.n1110 VDD.n910 18.5384
R2001 VDD.n1187 VDD.n870 18.5384
R2002 VDD.n535 VDD.n131 18.5384
R2003 VDD.n446 VDD.n166 18.5384
R2004 VDD.n357 VDD.n201 18.5384
R2005 VDD.n268 VDD.n236 18.5384
R2006 VDD.n644 VDD.n643 18.2197
R2007 VDD.n655 VDD.n73 18.2197
R2008 VDD.n657 VDD.n64 18.2197
R2009 VDD.n670 VDD.n668 18.2197
R2010 VDD.n682 VDD.n681 18.2197
R2011 VDD.n693 VDD.n51 18.2197
R2012 VDD.n708 VDD.n706 18.2197
R2013 VDD.n720 VDD.n719 18.2197
R2014 VDD.n734 VDD.n28 18.2197
R2015 VDD.n1240 VDD.n1239 18.0712
R2016 VDD.n1254 VDD.n843 18.0712
R2017 VDD.n1256 VDD.n835 18.0712
R2018 VDD.n1268 VDD.n1266 18.0712
R2019 VDD.n1279 VDD.n1278 18.0712
R2020 VDD.n1291 VDD.n822 18.0712
R2021 VDD.n1295 VDD.n1294 18.0712
R2022 VDD.n1308 VDD.n1307 18.0712
R2023 VDD.n1321 VDD.n808 18.0712
R2024 VDD.n1323 VDD.n803 18.0712
R2025 VDD.n1334 VDD.n1332 18.0712
R2026 VDD.n1345 VDD.n1344 18.0712
R2027 VDD.n1358 VDD.n790 18.0712
R2028 VDD.n1363 VDD.n1362 18.0712
R2029 VDD.n1374 VDD.n780 18.0712
R2030 VDD.n1376 VDD.n774 18.0712
R2031 VDD.n1387 VDD.n1385 18.0712
R2032 VDD.n2057 VDD.n2014 17.2143
R2033 VDD.n598 VDD.n105 17.2143
R2034 VDD.n627 VDD.n626 17.2143
R2035 VDD.n746 VDD.n23 16.9936
R2036 VDD.n1668 VDD.n1572 16.7993
R2037 VDD.n1742 VDD.n1529 16.7993
R2038 VDD.n1821 VDD.n1491 16.7993
R2039 VDD.n1895 VDD.n1448 16.7993
R2040 VDD.n1974 VDD.n1410 16.7993
R2041 VDD.n987 VDD.n969 16.7993
R2042 VDD.n1070 VDD.n934 16.7993
R2043 VDD.n1145 VDD.n893 16.7993
R2044 VDD.n1228 VDD.n858 16.7993
R2045 VDD.n585 VDD.n109 16.7993
R2046 VDD.n495 VDD.n144 16.7993
R2047 VDD.n406 VDD.n179 16.7993
R2048 VDD.n317 VDD.n214 16.7993
R2049 VDD.n757 VDD 16.7729
R2050 VDD.n2098 VDD 16.5522
R2051 VDD.n694 VDD.t294 15.6169
R2052 VDD.n1309 VDD.t114 15.4896
R2053 VDD.n1658 VDD.n1581 15.2281
R2054 VDD.n1731 VDD.n1538 15.2281
R2055 VDD.n1811 VDD.n1500 15.2281
R2056 VDD.n1884 VDD.n1457 15.2281
R2057 VDD.n1964 VDD.n1419 15.2281
R2058 VDD.n999 VDD.n961 15.2281
R2059 VDD.n1081 VDD.n925 15.2281
R2060 VDD.n1157 VDD.n885 15.2281
R2061 VDD.n1672 VDD.n1568 15.0074
R2062 VDD.n1749 VDD.n1527 15.0074
R2063 VDD.n1825 VDD.n1487 15.0074
R2064 VDD.n1902 VDD.n1446 15.0074
R2065 VDD.n1978 VDD.n1406 15.0074
R2066 VDD.n983 VDD.n975 15.0074
R2067 VDD.n1062 VDD.n937 15.0074
R2068 VDD.n1141 VDD.n899 15.0074
R2069 VDD.n1220 VDD.n861 15.0074
R2070 VDD.n593 VDD.n592 15.0074
R2071 VDD.n502 VDD.n142 15.0074
R2072 VDD.n413 VDD.n177 15.0074
R2073 VDD.n324 VDD.n212 15.0074
R2074 VDD.n1297 VDD.n1296 14.9976
R2075 VDD.n2095 VDD.n2094 14.566
R2076 VDD.n1243 VDD.n847 14.566
R2077 VDD.n1395 VDD.n769 14.3453
R2078 VDD.n636 VDD.n635 14.3453
R2079 VDD.n641 VDD.n639 14.3453
R2080 VDD.n740 VDD.n26 14.3453
R2081 VDD.n607 VDD.n606 13.6833
R2082 VDD.n620 VDD.n90 13.6833
R2083 VDD.n289 VDD 13.6005
R2084 VDD.n378 VDD 13.6005
R2085 VDD.n467 VDD 13.6005
R2086 VDD.n556 VDD 13.6005
R2087 VDD.n2686 VDD 13.6005
R2088 VDD.n2522 VDD 13.6005
R2089 VDD.n2398 VDD 13.6005
R2090 VDD.n2274 VDD 13.6005
R2091 VDD.n2036 VDD.n2028 13.4626
R2092 VDD.n1609 VDD.n1603 13.4626
R2093 VDD.n1685 VDD.n1561 13.4626
R2094 VDD.n1762 VDD.n1522 13.4626
R2095 VDD.n1838 VDD.n1480 13.4626
R2096 VDD.n1915 VDD.n1441 13.4626
R2097 VDD.n1049 VDD.n941 13.4626
R2098 VDD.n1129 VDD.n905 13.4626
R2099 VDD.n1207 VDD.n865 13.4626
R2100 VDD.n515 VDD.n137 13.4626
R2101 VDD.n426 VDD.n172 13.4626
R2102 VDD.n337 VDD.n207 13.4626
R2103 VDD.n248 VDD.n242 13.4626
R2104 VDD.t423 VDD.n1589 13.1949
R2105 VDD.n1711 VDD.t32 13.1949
R2106 VDD.t319 VDD.n1508 13.1949
R2107 VDD.n1864 VDD.t638 13.1949
R2108 VDD.t693 VDD.n1427 13.1949
R2109 VDD.n2669 VDD.t512 13.1584
R2110 VDD.n2536 VDD.t478 13.1584
R2111 VDD.n2412 VDD.t98 13.1584
R2112 VDD.n2288 VDD.t203 13.1584
R2113 VDD.n2154 VDD.t464 13.1584
R2114 VDD.n2098 VDD.n1990 13.0212
R2115 VDD.n2104 VDD.n1990 13.0212
R2116 VDD.n757 VDD.n15 13.0212
R2117 VDD.n763 VDD.n15 13.0212
R2118 VDD.t2 VDD.n228 13.0142
R2119 VDD.t112 VDD.n193 13.0142
R2120 VDD.t403 VDD.n158 13.0142
R2121 VDD.t138 VDD.n123 13.0142
R2122 VDD.n706 VDD.t292 13.0142
R2123 VDD.n1013 VDD.t665 12.9081
R2124 VDD.t563 VDD.n1100 12.9081
R2125 VDD.n1171 VDD.t285 12.9081
R2126 VDD.n1259 VDD.n1258 12.8005
R2127 VDD.n838 VDD.n833 12.8005
R2128 VDD.n1276 VDD.n1275 12.8005
R2129 VDD.n1284 VDD.n824 12.8005
R2130 VDD.n1305 VDD.n1304 12.8005
R2131 VDD.n1313 VDD.n810 12.8005
R2132 VDD.n1328 VDD.n801 12.8005
R2133 VDD.n1342 VDD.n1341 12.8005
R2134 VDD.n1350 VDD.n792 12.8005
R2135 VDD.n649 VDD.n75 12.8005
R2136 VDD.n67 VDD.n62 12.8005
R2137 VDD.n687 VDD.n53 12.8005
R2138 VDD.n45 VDD.n40 12.8005
R2139 VDD.n725 VDD.n30 12.8005
R2140 VDD.n2030 VDD.n2028 12.5798
R2141 VDD.n1615 VDD.n1603 12.5798
R2142 VDD.n1615 VDD.n1599 12.5798
R2143 VDD.n1679 VDD.n1568 12.5798
R2144 VDD.n1685 VDD.n1564 12.5798
R2145 VDD.n1692 VDD.n1561 12.5798
R2146 VDD.n1692 VDD.n1559 12.5798
R2147 VDD.n1756 VDD.n1527 12.5798
R2148 VDD.n1762 VDD.n1524 12.5798
R2149 VDD.n1768 VDD.n1522 12.5798
R2150 VDD.n1768 VDD.n1518 12.5798
R2151 VDD.n1832 VDD.n1487 12.5798
R2152 VDD.n1838 VDD.n1483 12.5798
R2153 VDD.n1845 VDD.n1480 12.5798
R2154 VDD.n1845 VDD.n1478 12.5798
R2155 VDD.n1909 VDD.n1446 12.5798
R2156 VDD.n1915 VDD.n1443 12.5798
R2157 VDD.n1921 VDD.n1441 12.5798
R2158 VDD.n1921 VDD.n1437 12.5798
R2159 VDD.n1983 VDD.n1406 12.5798
R2160 VDD.n1609 VDD.n1608 12.5798
R2161 VDD.n1041 VDD.n943 12.5798
R2162 VDD.n1041 VDD.n941 12.5798
R2163 VDD.n1049 VDD.n938 12.5798
R2164 VDD.n1056 VDD.n937 12.5798
R2165 VDD.n1122 VDD.n908 12.5798
R2166 VDD.n1122 VDD.n905 12.5798
R2167 VDD.n1129 VDD.n902 12.5798
R2168 VDD.n1134 VDD.n899 12.5798
R2169 VDD.n1199 VDD.n867 12.5798
R2170 VDD.n1199 VDD.n865 12.5798
R2171 VDD.n1207 VDD.n862 12.5798
R2172 VDD.n1214 VDD.n861 12.5798
R2173 VDD.n977 VDD.n975 12.5798
R2174 VDD.n593 VDD.n104 12.5798
R2175 VDD.n568 VDD.n564 12.5798
R2176 VDD.n509 VDD.n142 12.5798
R2177 VDD.n515 VDD.n139 12.5798
R2178 VDD.n521 VDD.n137 12.5798
R2179 VDD.n521 VDD.n133 12.5798
R2180 VDD.n479 VDD.n475 12.5798
R2181 VDD.n420 VDD.n177 12.5798
R2182 VDD.n426 VDD.n174 12.5798
R2183 VDD.n432 VDD.n172 12.5798
R2184 VDD.n432 VDD.n168 12.5798
R2185 VDD.n390 VDD.n386 12.5798
R2186 VDD.n331 VDD.n212 12.5798
R2187 VDD.n337 VDD.n209 12.5798
R2188 VDD.n343 VDD.n207 12.5798
R2189 VDD.n343 VDD.n203 12.5798
R2190 VDD.n301 VDD.n297 12.5798
R2191 VDD.n254 VDD.n242 12.5798
R2192 VDD.n254 VDD.n238 12.5798
R2193 VDD.n248 VDD.n247 12.5798
R2194 VDD.n2047 VDD.n2020 12.1384
R2195 VDD.n717 VDD.n716 12.1384
R2196 VDD.n1381 VDD.n776 11.6971
R2197 VDD.n2094 VDD.n1994 11.4764
R2198 VDD.n661 VDD.n660 11.2557
R2199 VDD.n1607 VDD 11.0898
R2200 VDD.n246 VDD 11.0536
R2201 VDD.n296 VDD.n295 10.9416
R2202 VDD.n385 VDD.n384 10.9416
R2203 VDD.n474 VDD.n473 10.9416
R2204 VDD.n563 VDD.n562 10.9416
R2205 VDD.n1366 VDD.n785 10.8143
R2206 VDD.n770 VDD.n766 10.8143
R2207 VDD.n2043 VDD.t85 10.4977
R2208 VDD.t508 VDD.n613 10.4115
R2209 VDD.n614 VDD.t502 10.4115
R2210 VDD.t294 VDD.n693 10.4115
R2211 VDD.t298 VDD.n42 10.4115
R2212 VDD.n611 VDD.n98 10.1522
R2213 VDD.n98 VDD.n92 10.1522
R2214 VDD.n1401 VDD.n766 9.49016
R2215 VDD.n1393 VDD.n769 9.3005
R2216 VDD.n1390 VDD.n771 9.3005
R2217 VDD.n1390 VDD.n768 9.3005
R2218 VDD.n1386 VDD.n768 9.3005
R2219 VDD.n1381 VDD.n778 9.3005
R2220 VDD.n1384 VDD.n1383 9.3005
R2221 VDD.n1381 VDD.n777 9.3005
R2222 VDD.n1371 VDD.n1370 9.3005
R2223 VDD.n1371 VDD.n779 9.3005
R2224 VDD.n1375 VDD.n779 9.3005
R2225 VDD.n1368 VDD.n776 9.3005
R2226 VDD.n1366 VDD.n787 9.3005
R2227 VDD.n1361 VDD.n1360 9.3005
R2228 VDD.n1367 VDD.n1366 9.3005
R2229 VDD.n1355 VDD.n1354 9.3005
R2230 VDD.n1355 VDD.n788 9.3005
R2231 VDD.n1359 VDD.n788 9.3005
R2232 VDD.n1352 VDD.n785 9.3005
R2233 VDD.n1348 VDD.n796 9.3005
R2234 VDD.n1348 VDD.n1347 9.3005
R2235 VDD.n1347 VDD.n1346 9.3005
R2236 VDD.n1351 VDD.n1350 9.3005
R2237 VDD.n1338 VDD.n1337 9.3005
R2238 VDD.n1337 VDD.n798 9.3005
R2239 VDD.n1333 VDD.n798 9.3005
R2240 VDD.n1341 VDD.n1340 9.3005
R2241 VDD.n1328 VDD.n806 9.3005
R2242 VDD.n1331 VDD.n1330 9.3005
R2243 VDD.n1328 VDD.n800 9.3005
R2244 VDD.n1318 VDD.n1317 9.3005
R2245 VDD.n1318 VDD.n807 9.3005
R2246 VDD.n1322 VDD.n807 9.3005
R2247 VDD.n1315 VDD.n805 9.3005
R2248 VDD.n1311 VDD.n814 9.3005
R2249 VDD.n1311 VDD.n1310 9.3005
R2250 VDD.n1310 VDD.n1309 9.3005
R2251 VDD.n1314 VDD.n1313 9.3005
R2252 VDD.n1301 VDD.n1300 9.3005
R2253 VDD.n1300 VDD.n816 9.3005
R2254 VDD.n1293 VDD.n816 9.3005
R2255 VDD.n1304 VDD.n1303 9.3005
R2256 VDD.n1288 VDD.n1287 9.3005
R2257 VDD.n1288 VDD.n821 9.3005
R2258 VDD.n1292 VDD.n821 9.3005
R2259 VDD.n819 VDD.n818 9.3005
R2260 VDD.n1282 VDD.n828 9.3005
R2261 VDD.n1282 VDD.n1281 9.3005
R2262 VDD.n1281 VDD.n1280 9.3005
R2263 VDD.n1285 VDD.n1284 9.3005
R2264 VDD.n1272 VDD.n1271 9.3005
R2265 VDD.n1271 VDD.n830 9.3005
R2266 VDD.n1267 VDD.n830 9.3005
R2267 VDD.n1275 VDD.n1274 9.3005
R2268 VDD.n1263 VDD.n1262 9.3005
R2269 VDD.n1264 VDD.n1263 9.3005
R2270 VDD.n1265 VDD.n1264 9.3005
R2271 VDD.n838 VDD.n832 9.3005
R2272 VDD.n1251 VDD.n1250 9.3005
R2273 VDD.n1251 VDD.n842 9.3005
R2274 VDD.n1255 VDD.n842 9.3005
R2275 VDD.n1260 VDD.n1259 9.3005
R2276 VDD.n1248 VDD.n1245 9.3005
R2277 VDD.n1237 VDD.n1236 9.3005
R2278 VDD.n1249 VDD.n1248 9.3005
R2279 VDD.n295 VDD.n293 9.3005
R2280 VDD.n384 VDD.n382 9.3005
R2281 VDD.n473 VDD.n471 9.3005
R2282 VDD.n562 VDD.n560 9.3005
R2283 VDD.n727 VDD.n26 9.3005
R2284 VDD.n731 VDD.n730 9.3005
R2285 VDD.n731 VDD.n27 9.3005
R2286 VDD.n735 VDD.n27 9.3005
R2287 VDD.n723 VDD.n34 9.3005
R2288 VDD.n723 VDD.n722 9.3005
R2289 VDD.n722 VDD.n721 9.3005
R2290 VDD.n726 VDD.n725 9.3005
R2291 VDD.n712 VDD.n711 9.3005
R2292 VDD.n711 VDD.n36 9.3005
R2293 VDD.n707 VDD.n36 9.3005
R2294 VDD.n715 VDD.n714 9.3005
R2295 VDD.n703 VDD.n702 9.3005
R2296 VDD.n704 VDD.n703 9.3005
R2297 VDD.n705 VDD.n704 9.3005
R2298 VDD.n45 VDD.n39 9.3005
R2299 VDD.n690 VDD.n689 9.3005
R2300 VDD.n690 VDD.n50 9.3005
R2301 VDD.n694 VDD.n50 9.3005
R2302 VDD.n700 VDD.n699 9.3005
R2303 VDD.n685 VDD.n56 9.3005
R2304 VDD.n685 VDD.n684 9.3005
R2305 VDD.n684 VDD.n683 9.3005
R2306 VDD.n688 VDD.n687 9.3005
R2307 VDD.n674 VDD.n673 9.3005
R2308 VDD.n673 VDD.n58 9.3005
R2309 VDD.n669 VDD.n58 9.3005
R2310 VDD.n677 VDD.n676 9.3005
R2311 VDD.n665 VDD.n664 9.3005
R2312 VDD.n666 VDD.n665 9.3005
R2313 VDD.n667 VDD.n666 9.3005
R2314 VDD.n67 VDD.n61 9.3005
R2315 VDD.n652 VDD.n651 9.3005
R2316 VDD.n652 VDD.n72 9.3005
R2317 VDD.n656 VDD.n72 9.3005
R2318 VDD.n662 VDD.n661 9.3005
R2319 VDD.n647 VDD.n79 9.3005
R2320 VDD.n647 VDD.n646 9.3005
R2321 VDD.n646 VDD.n645 9.3005
R2322 VDD.n650 VDD.n649 9.3005
R2323 VDD.n639 VDD.n81 9.3005
R2324 VDD.n631 VDD.n81 9.3005
R2325 VDD.n2242 VDD.n2240 9.3005
R2326 VDD.n2240 VDD.n2239 9.3005
R2327 VDD.n1659 VDD.n1578 9.11136
R2328 VDD.n1539 VDD.n1535 9.11136
R2329 VDD.n1812 VDD.n1497 9.11136
R2330 VDD.n1458 VDD.n1454 9.11136
R2331 VDD.n1965 VDD.n1416 9.11136
R2332 VDD.n994 VDD.n964 9.11136
R2333 VDD.n932 VDD.n927 9.11136
R2334 VDD.n1152 VDD.n888 9.11136
R2335 VDD.n856 VDD.n850 9.11136
R2336 VDD.n567 VDD.n115 9.11136
R2337 VDD.n478 VDD.n150 9.11136
R2338 VDD.n389 VDD.n185 9.11136
R2339 VDD.n300 VDD.n220 9.11136
R2340 VDD.n746 VDD.n745 9.04877
R2341 VDD.n290 VDD.n288 8.91563
R2342 VDD.n379 VDD.n377 8.91563
R2343 VDD.n468 VDD.n466 8.91563
R2344 VDD.n557 VDD.n555 8.91563
R2345 VDD.n1662 VDD.n1579 8.78856
R2346 VDD.n1739 VDD.n1738 8.78856
R2347 VDD.n1815 VDD.n1498 8.78856
R2348 VDD.n1892 VDD.n1891 8.78856
R2349 VDD.n1968 VDD.n1417 8.78856
R2350 VDD.n995 VDD.n966 8.78856
R2351 VDD.n1074 VDD.n931 8.78856
R2352 VDD.n1153 VDD.n890 8.78856
R2353 VDD.n1232 VDD.n855 8.78856
R2354 VDD.n581 VDD.n580 8.78856
R2355 VDD.n492 VDD.n491 8.78856
R2356 VDD.n403 VDD.n402 8.78856
R2357 VDD.n314 VDD.n313 8.78856
R2358 VDD.n1651 VDD.n1581 8.6074
R2359 VDD.n1724 VDD.n1538 8.6074
R2360 VDD.n1804 VDD.n1500 8.6074
R2361 VDD.n1877 VDD.n1457 8.6074
R2362 VDD.n1957 VDD.n1419 8.6074
R2363 VDD.n1006 VDD.n961 8.6074
R2364 VDD.n1087 VDD.n925 8.6074
R2365 VDD.n1164 VDD.n885 8.6074
R2366 VDD.n698 VDD.n697 8.6074
R2367 VDD.n573 VDD.n572 8.6074
R2368 VDD.n484 VDD.n483 8.6074
R2369 VDD.n395 VDD.n394 8.6074
R2370 VDD.n306 VDD.n305 8.6074
R2371 VDD.n976 VDD.n975 8.47522
R2372 VDD.n593 VDD.n108 8.47522
R2373 VDD.n142 VDD.n141 8.47522
R2374 VDD.n177 VDD.n176 8.47522
R2375 VDD.n212 VDD.n211 8.47522
R2376 VDD.n2608 VDD.n2607 8.47522
R2377 VDD.n1407 VDD.n1406 8.47518
R2378 VDD.n1446 VDD.n1445 8.47518
R2379 VDD.n1488 VDD.n1487 8.47518
R2380 VDD.n1527 VDD.n1526 8.47518
R2381 VDD.n1569 VDD.n1568 8.47518
R2382 VDD.n861 VDD.n860 8.47518
R2383 VDD.n900 VDD.n899 8.47518
R2384 VDD.n937 VDD.n936 8.47518
R2385 VDD.n2219 VDD.n2218 8.47518
R2386 VDD.n2351 VDD.n2350 8.47518
R2387 VDD.n2475 VDD.n2474 8.47518
R2388 VDD.n2599 VDD.n2598 8.47518
R2389 VDD.n1991 VDD.n1990 8.47281
R2390 VDD.n1609 VDD.n1605 8.47281
R2391 VDD.n248 VDD.n244 8.47281
R2392 VDD.n2094 VDD.n2091 8.47276
R2393 VDD.n1915 VDD.n1914 8.47276
R2394 VDD.n1839 VDD.n1838 8.47276
R2395 VDD.n1762 VDD.n1761 8.47276
R2396 VDD.n1686 VDD.n1685 8.47276
R2397 VDD.n1208 VDD.n1207 8.47276
R2398 VDD.n1129 VDD.n1128 8.47276
R2399 VDD.n1050 VDD.n1049 8.47276
R2400 VDD.n16 VDD.n15 8.47276
R2401 VDD.n747 VDD.n746 8.47276
R2402 VDD.n515 VDD.n514 8.47276
R2403 VDD.n426 VDD.n425 8.47276
R2404 VDD.n337 VDD.n336 8.47276
R2405 VDD.n2114 VDD.n2113 8.47276
R2406 VDD.n2229 VDD.n2228 8.47276
R2407 VDD.n2361 VDD.n2360 8.47276
R2408 VDD.n2485 VDD.n2484 8.47276
R2409 VDD.n2724 VDD.n2723 8.47276
R2410 VDD.n2029 VDD.n2028 8.47181
R2411 VDD.n2246 VDD.n2245 8.47164
R2412 VDD.n2370 VDD.n2369 8.47164
R2413 VDD.n2494 VDD.n2493 8.47164
R2414 VDD.n2712 VDD.n2711 8.47164
R2415 VDD.n1922 VDD.n1921 8.4716
R2416 VDD.n1845 VDD.n1844 8.4716
R2417 VDD.n1769 VDD.n1768 8.4716
R2418 VDD.n1692 VDD.n1691 8.4716
R2419 VDD.n1616 VDD.n1615 8.4716
R2420 VDD.n1199 VDD.n1198 8.4716
R2421 VDD.n1123 VDD.n1122 8.4716
R2422 VDD.n1041 VDD.n1040 8.4716
R2423 VDD.n522 VDD.n521 8.4716
R2424 VDD.n433 VDD.n432 8.4716
R2425 VDD.n344 VDD.n343 8.4716
R2426 VDD.n255 VDD.n254 8.4716
R2427 VDD.n2123 VDD.n2122 8.4716
R2428 VDD.n2057 VDD.n2056 8.47092
R2429 VDD.n2180 VDD.n2179 8.47011
R2430 VDD.n1420 VDD.n1419 8.47007
R2431 VDD.n1936 VDD.n1935 8.47007
R2432 VDD.n1457 VDD.n1456 8.47007
R2433 VDD.n1856 VDD.n1855 8.47007
R2434 VDD.n1501 VDD.n1500 8.47007
R2435 VDD.n1783 VDD.n1782 8.47007
R2436 VDD.n1538 VDD.n1537 8.47007
R2437 VDD.n1703 VDD.n1702 8.47007
R2438 VDD.n1582 VDD.n1581 8.47007
R2439 VDD.n1630 VDD.n1629 8.47007
R2440 VDD.n1187 VDD.n1186 8.47007
R2441 VDD.n886 VDD.n885 8.47007
R2442 VDD.n1111 VDD.n1110 8.47007
R2443 VDD.n925 VDD.n924 8.47007
R2444 VDD.n1029 VDD.n1028 8.47007
R2445 VDD.n962 VDD.n961 8.47007
R2446 VDD.n536 VDD.n535 8.47007
R2447 VDD.n447 VDD.n446 8.47007
R2448 VDD.n358 VDD.n357 8.47007
R2449 VDD.n269 VDD.n268 8.47007
R2450 VDD.n2141 VDD.n2140 8.47007
R2451 VDD.n2314 VDD.n2313 8.47007
R2452 VDD.n2438 VDD.n2437 8.47007
R2453 VDD.n2562 VDD.n2561 8.47007
R2454 VDD.n2645 VDD.n2644 8.47007
R2455 VDD.n2081 VDD.n2080 8.45089
R2456 VDD.n2080 VDD.n1996 8.45089
R2457 VDD.n2079 VDD.n2078 8.45089
R2458 VDD.n2077 VDD.n1999 8.45089
R2459 VDD.n2076 VDD.n2075 8.45089
R2460 VDD.n2066 VDD.n2000 8.45089
R2461 VDD.n2068 VDD.n2067 8.45089
R2462 VDD.n2065 VDD.n2009 8.45089
R2463 VDD.n2064 VDD.n2063 8.45089
R2464 VDD.n2011 VDD.n2010 8.45089
R2465 VDD.n2056 VDD.n2055 8.45089
R2466 VDD.n2054 VDD.n2015 8.45089
R2467 VDD.n2053 VDD.n2052 8.45089
R2468 VDD.n2044 VDD.n2016 8.45089
R2469 VDD.n2046 VDD.n2045 8.45089
R2470 VDD.n2043 VDD.n2021 8.45089
R2471 VDD.n2042 VDD.n2041 8.45089
R2472 VDD.n2033 VDD.n2022 8.45089
R2473 VDD.n2035 VDD.n2034 8.45089
R2474 VDD.n2032 VDD.n2029 8.45089
R2475 VDD.n2099 VDD.n2098 8.45089
R2476 VDD.n2100 VDD.n2099 8.45089
R2477 VDD.n2089 VDD.n1992 8.45089
R2478 VDD.n2091 VDD.n2090 8.45089
R2479 VDD.n2088 VDD.n1995 8.45089
R2480 VDD.n2087 VDD.n2086 8.45089
R2481 VDD.n2101 VDD.n1991 8.45089
R2482 VDD.n2104 VDD.n2103 8.45089
R2483 VDD.n2103 VDD.n2102 8.45089
R2484 VDD.n1983 VDD.n1982 8.45089
R2485 VDD.n1981 VDD.n1407 8.45089
R2486 VDD.n1980 VDD.n1979 8.45089
R2487 VDD.n1409 VDD.n1408 8.45089
R2488 VDD.n1973 VDD.n1972 8.45089
R2489 VDD.n1971 VDD.n1414 8.45089
R2490 VDD.n1970 VDD.n1969 8.45089
R2491 VDD.n1961 VDD.n1415 8.45089
R2492 VDD.n1963 VDD.n1962 8.45089
R2493 VDD.n1960 VDD.n1420 8.45089
R2494 VDD.n1959 VDD.n1958 8.45089
R2495 VDD.n1422 VDD.n1421 8.45089
R2496 VDD.n1949 VDD.t722 8.45089
R2497 VDD.n1948 VDD.n1426 8.45089
R2498 VDD.n1947 VDD.n1946 8.45089
R2499 VDD.n1428 VDD.n1427 8.45089
R2500 VDD.n1940 VDD.n1939 8.45089
R2501 VDD.n1938 VDD.n1433 8.45089
R2502 VDD.n1937 VDD.n1936 8.45089
R2503 VDD.n1925 VDD.n1434 8.45089
R2504 VDD.n1927 VDD.n1926 8.45089
R2505 VDD.n1924 VDD.n1438 8.45089
R2506 VDD.n1923 VDD.n1922 8.45089
R2507 VDD.n1440 VDD.n1439 8.45089
R2508 VDD.n1914 VDD.n1913 8.45089
R2509 VDD.n1912 VDD.n1444 8.45089
R2510 VDD.n1911 VDD.n1910 8.45089
R2511 VDD.n1899 VDD.n1445 8.45089
R2512 VDD.n1901 VDD.n1900 8.45089
R2513 VDD.n1898 VDD.n1449 8.45089
R2514 VDD.n1897 VDD.n1896 8.45089
R2515 VDD.n1888 VDD.n1450 8.45089
R2516 VDD.n1890 VDD.n1889 8.45089
R2517 VDD.n1887 VDD.n1455 8.45089
R2518 VDD.n1886 VDD.n1885 8.45089
R2519 VDD.n1874 VDD.n1456 8.45089
R2520 VDD.n1876 VDD.n1875 8.45089
R2521 VDD.n1873 VDD.n1461 8.45089
R2522 VDD.t432 VDD.n1872 8.45089
R2523 VDD.n1463 VDD.n1462 8.45089
R2524 VDD.n1866 VDD.n1865 8.45089
R2525 VDD.n1864 VDD.n1468 8.45089
R2526 VDD.n1863 VDD.n1862 8.45089
R2527 VDD.n1470 VDD.n1469 8.45089
R2528 VDD.n1855 VDD.n1854 8.45089
R2529 VDD.n1853 VDD.n1476 8.45089
R2530 VDD.n1852 VDD.n1851 8.45089
R2531 VDD.n1842 VDD.n1477 8.45089
R2532 VDD.n1844 VDD.n1843 8.45089
R2533 VDD.n1841 VDD.n1481 8.45089
R2534 VDD.n1840 VDD.n1839 8.45089
R2535 VDD.n1829 VDD.n1482 8.45089
R2536 VDD.n1831 VDD.n1830 8.45089
R2537 VDD.n1828 VDD.n1488 8.45089
R2538 VDD.n1827 VDD.n1826 8.45089
R2539 VDD.n1490 VDD.n1489 8.45089
R2540 VDD.n1820 VDD.n1819 8.45089
R2541 VDD.n1818 VDD.n1495 8.45089
R2542 VDD.n1817 VDD.n1816 8.45089
R2543 VDD.n1808 VDD.n1496 8.45089
R2544 VDD.n1810 VDD.n1809 8.45089
R2545 VDD.n1807 VDD.n1501 8.45089
R2546 VDD.n1806 VDD.n1805 8.45089
R2547 VDD.n1503 VDD.n1502 8.45089
R2548 VDD.n1796 VDD.t351 8.45089
R2549 VDD.n1795 VDD.n1507 8.45089
R2550 VDD.n1794 VDD.n1793 8.45089
R2551 VDD.n1509 VDD.n1508 8.45089
R2552 VDD.n1787 VDD.n1786 8.45089
R2553 VDD.n1785 VDD.n1514 8.45089
R2554 VDD.n1784 VDD.n1783 8.45089
R2555 VDD.n1772 VDD.n1515 8.45089
R2556 VDD.n1774 VDD.n1773 8.45089
R2557 VDD.n1771 VDD.n1519 8.45089
R2558 VDD.n1770 VDD.n1769 8.45089
R2559 VDD.n1521 VDD.n1520 8.45089
R2560 VDD.n1761 VDD.n1760 8.45089
R2561 VDD.n1759 VDD.n1525 8.45089
R2562 VDD.n1758 VDD.n1757 8.45089
R2563 VDD.n1746 VDD.n1526 8.45089
R2564 VDD.n1748 VDD.n1747 8.45089
R2565 VDD.n1745 VDD.n1530 8.45089
R2566 VDD.n1744 VDD.n1743 8.45089
R2567 VDD.n1735 VDD.n1531 8.45089
R2568 VDD.n1737 VDD.n1736 8.45089
R2569 VDD.n1734 VDD.n1536 8.45089
R2570 VDD.n1733 VDD.n1732 8.45089
R2571 VDD.n1721 VDD.n1537 8.45089
R2572 VDD.n1723 VDD.n1722 8.45089
R2573 VDD.n1720 VDD.n1542 8.45089
R2574 VDD.t12 VDD.n1719 8.45089
R2575 VDD.n1544 VDD.n1543 8.45089
R2576 VDD.n1713 VDD.n1712 8.45089
R2577 VDD.n1711 VDD.n1549 8.45089
R2578 VDD.n1710 VDD.n1709 8.45089
R2579 VDD.n1551 VDD.n1550 8.45089
R2580 VDD.n1702 VDD.n1701 8.45089
R2581 VDD.n1700 VDD.n1557 8.45089
R2582 VDD.n1699 VDD.n1698 8.45089
R2583 VDD.n1689 VDD.n1558 8.45089
R2584 VDD.n1691 VDD.n1690 8.45089
R2585 VDD.n1688 VDD.n1562 8.45089
R2586 VDD.n1687 VDD.n1686 8.45089
R2587 VDD.n1676 VDD.n1563 8.45089
R2588 VDD.n1678 VDD.n1677 8.45089
R2589 VDD.n1675 VDD.n1569 8.45089
R2590 VDD.n1674 VDD.n1673 8.45089
R2591 VDD.n1571 VDD.n1570 8.45089
R2592 VDD.n1667 VDD.n1666 8.45089
R2593 VDD.n1665 VDD.n1576 8.45089
R2594 VDD.n1664 VDD.n1663 8.45089
R2595 VDD.n1655 VDD.n1577 8.45089
R2596 VDD.n1657 VDD.n1656 8.45089
R2597 VDD.n1654 VDD.n1582 8.45089
R2598 VDD.n1653 VDD.n1652 8.45089
R2599 VDD.n1584 VDD.n1583 8.45089
R2600 VDD.n1643 VDD.t460 8.45089
R2601 VDD.n1642 VDD.n1588 8.45089
R2602 VDD.n1641 VDD.n1640 8.45089
R2603 VDD.n1590 VDD.n1589 8.45089
R2604 VDD.n1634 VDD.n1633 8.45089
R2605 VDD.n1632 VDD.n1595 8.45089
R2606 VDD.n1631 VDD.n1630 8.45089
R2607 VDD.n1619 VDD.n1596 8.45089
R2608 VDD.n1621 VDD.n1620 8.45089
R2609 VDD.n1618 VDD.n1600 8.45089
R2610 VDD.n1617 VDD.n1616 8.45089
R2611 VDD.n1602 VDD.n1601 8.45089
R2612 VDD.n1606 VDD.n1605 8.45089
R2613 VDD.n1608 VDD.n1607 8.45089
R2614 VDD.n1401 VDD.n1400 8.45089
R2615 VDD.n1400 VDD.n1399 8.45089
R2616 VDD.n1398 VDD.n767 8.45089
R2617 VDD.n1397 VDD.n1396 8.45089
R2618 VDD.n1242 VDD.n1241 8.45089
R2619 VDD.n1235 VDD.n851 8.45089
R2620 VDD.n1234 VDD.n1233 8.45089
R2621 VDD.n854 VDD.n853 8.45089
R2622 VDD.n1225 VDD.n1224 8.45089
R2623 VDD.n1223 VDD.n859 8.45089
R2624 VDD.n1222 VDD.n1221 8.45089
R2625 VDD.n1211 VDD.n860 8.45089
R2626 VDD.n1213 VDD.n1212 8.45089
R2627 VDD.n1210 VDD.n863 8.45089
R2628 VDD.n1209 VDD.n1208 8.45089
R2629 VDD.n1196 VDD.n864 8.45089
R2630 VDD.n1198 VDD.n1197 8.45089
R2631 VDD.n1195 VDD.n868 8.45089
R2632 VDD.n1194 VDD.n1193 8.45089
R2633 VDD.n1184 VDD.n869 8.45089
R2634 VDD.n1186 VDD.n1185 8.45089
R2635 VDD.n1183 VDD.n874 8.45089
R2636 VDD.n1182 VDD.n1181 8.45089
R2637 VDD.n1171 VDD.n875 8.45089
R2638 VDD.n1173 VDD.n1172 8.45089
R2639 VDD.n1170 VDD.n879 8.45089
R2640 VDD.t637 VDD.n1169 8.45089
R2641 VDD.n1161 VDD.n880 8.45089
R2642 VDD.n1163 VDD.n1162 8.45089
R2643 VDD.n1160 VDD.n886 8.45089
R2644 VDD.n1159 VDD.n1158 8.45089
R2645 VDD.n1149 VDD.n887 8.45089
R2646 VDD.n1151 VDD.n1150 8.45089
R2647 VDD.n1148 VDD.n891 8.45089
R2648 VDD.n1147 VDD.n1146 8.45089
R2649 VDD.n1138 VDD.n892 8.45089
R2650 VDD.n1140 VDD.n1139 8.45089
R2651 VDD.n1137 VDD.n900 8.45089
R2652 VDD.n1136 VDD.n1135 8.45089
R2653 VDD.n1126 VDD.n901 8.45089
R2654 VDD.n1128 VDD.n1127 8.45089
R2655 VDD.n1125 VDD.n906 8.45089
R2656 VDD.n1124 VDD.n1123 8.45089
R2657 VDD.n1114 VDD.n907 8.45089
R2658 VDD.n1116 VDD.n1115 8.45089
R2659 VDD.n1113 VDD.n911 8.45089
R2660 VDD.n1112 VDD.n1111 8.45089
R2661 VDD.n1101 VDD.n912 8.45089
R2662 VDD.n1103 VDD.n1102 8.45089
R2663 VDD.n1100 VDD.n916 8.45089
R2664 VDD.n1099 VDD.n1098 8.45089
R2665 VDD.n1091 VDD.n917 8.45089
R2666 VDD.n1092 VDD.t268 8.45089
R2667 VDD.n1090 VDD.n923 8.45089
R2668 VDD.n1089 VDD.n1088 8.45089
R2669 VDD.n1078 VDD.n924 8.45089
R2670 VDD.n1080 VDD.n1079 8.45089
R2671 VDD.n1077 VDD.n928 8.45089
R2672 VDD.n1076 VDD.n1075 8.45089
R2673 VDD.n930 VDD.n929 8.45089
R2674 VDD.n1067 VDD.n1066 8.45089
R2675 VDD.n1065 VDD.n935 8.45089
R2676 VDD.n1064 VDD.n1063 8.45089
R2677 VDD.n1053 VDD.n936 8.45089
R2678 VDD.n1055 VDD.n1054 8.45089
R2679 VDD.n1052 VDD.n939 8.45089
R2680 VDD.n1051 VDD.n1050 8.45089
R2681 VDD.n1038 VDD.n940 8.45089
R2682 VDD.n1040 VDD.n1039 8.45089
R2683 VDD.n1037 VDD.n944 8.45089
R2684 VDD.n1036 VDD.n1035 8.45089
R2685 VDD.n1026 VDD.n945 8.45089
R2686 VDD.n1028 VDD.n1027 8.45089
R2687 VDD.n1025 VDD.n950 8.45089
R2688 VDD.n1024 VDD.n1023 8.45089
R2689 VDD.n1013 VDD.n951 8.45089
R2690 VDD.n1015 VDD.n1014 8.45089
R2691 VDD.n1012 VDD.n955 8.45089
R2692 VDD.t335 VDD.n1011 8.45089
R2693 VDD.n1003 VDD.n956 8.45089
R2694 VDD.n1005 VDD.n1004 8.45089
R2695 VDD.n1002 VDD.n962 8.45089
R2696 VDD.n1001 VDD.n1000 8.45089
R2697 VDD.n991 VDD.n963 8.45089
R2698 VDD.n993 VDD.n992 8.45089
R2699 VDD.n990 VDD.n967 8.45089
R2700 VDD.n989 VDD.n988 8.45089
R2701 VDD.n980 VDD.n968 8.45089
R2702 VDD.n982 VDD.n981 8.45089
R2703 VDD.n979 VDD.n976 8.45089
R2704 VDD.n978 VDD.n977 8.45089
R2705 VDD.n763 VDD.n762 8.45089
R2706 VDD.n762 VDD.n761 8.45089
R2707 VDD.n760 VDD.n16 8.45089
R2708 VDD.n759 VDD.n758 8.45089
R2709 VDD.n750 VDD.n17 8.45089
R2710 VDD.n752 VDD.n751 8.45089
R2711 VDD.n749 VDD.n21 8.45089
R2712 VDD.n748 VDD.n747 8.45089
R2713 VDD.n736 VDD.n22 8.45089
R2714 VDD.n738 VDD.n737 8.45089
R2715 VDD.n630 VDD.n86 8.45089
R2716 VDD.n629 VDD.n628 8.45089
R2717 VDD.n615 VDD.n88 8.45089
R2718 VDD.n616 VDD.n94 8.45089
R2719 VDD.n618 VDD.n617 8.45089
R2720 VDD.n614 VDD.n93 8.45089
R2721 VDD.n613 VDD.n612 8.45089
R2722 VDD.n602 VDD.n95 8.45089
R2723 VDD.n604 VDD.n603 8.45089
R2724 VDD.n601 VDD.n101 8.45089
R2725 VDD.n600 VDD.n599 8.45089
R2726 VDD.n103 VDD.n102 8.45089
R2727 VDD.n589 VDD.n108 8.45089
R2728 VDD.n591 VDD.n590 8.45089
R2729 VDD.n588 VDD.n110 8.45089
R2730 VDD.n587 VDD.n586 8.45089
R2731 VDD.n577 VDD.n111 8.45089
R2732 VDD.n579 VDD.n578 8.45089
R2733 VDD.n576 VDD.n116 8.45089
R2734 VDD.n574 VDD.n573 8.45089
R2735 VDD.n575 VDD.n574 8.45089
R2736 VDD.n118 VDD.n117 8.45089
R2737 VDD.n549 VDD.t516 8.45089
R2738 VDD.n548 VDD.n122 8.45089
R2739 VDD.n547 VDD.n546 8.45089
R2740 VDD.n124 VDD.n123 8.45089
R2741 VDD.n540 VDD.n539 8.45089
R2742 VDD.n538 VDD.n129 8.45089
R2743 VDD.n537 VDD.n536 8.45089
R2744 VDD.n525 VDD.n130 8.45089
R2745 VDD.n527 VDD.n526 8.45089
R2746 VDD.n524 VDD.n134 8.45089
R2747 VDD.n523 VDD.n522 8.45089
R2748 VDD.n136 VDD.n135 8.45089
R2749 VDD.n514 VDD.n513 8.45089
R2750 VDD.n512 VDD.n140 8.45089
R2751 VDD.n511 VDD.n510 8.45089
R2752 VDD.n499 VDD.n141 8.45089
R2753 VDD.n501 VDD.n500 8.45089
R2754 VDD.n498 VDD.n145 8.45089
R2755 VDD.n497 VDD.n496 8.45089
R2756 VDD.n488 VDD.n146 8.45089
R2757 VDD.n490 VDD.n489 8.45089
R2758 VDD.n487 VDD.n151 8.45089
R2759 VDD.n485 VDD.n484 8.45089
R2760 VDD.n486 VDD.n485 8.45089
R2761 VDD.n153 VDD.n152 8.45089
R2762 VDD.n460 VDD.t104 8.45089
R2763 VDD.n459 VDD.n157 8.45089
R2764 VDD.n458 VDD.n457 8.45089
R2765 VDD.n159 VDD.n158 8.45089
R2766 VDD.n451 VDD.n450 8.45089
R2767 VDD.n449 VDD.n164 8.45089
R2768 VDD.n448 VDD.n447 8.45089
R2769 VDD.n436 VDD.n165 8.45089
R2770 VDD.n438 VDD.n437 8.45089
R2771 VDD.n435 VDD.n169 8.45089
R2772 VDD.n434 VDD.n433 8.45089
R2773 VDD.n171 VDD.n170 8.45089
R2774 VDD.n425 VDD.n424 8.45089
R2775 VDD.n423 VDD.n175 8.45089
R2776 VDD.n422 VDD.n421 8.45089
R2777 VDD.n410 VDD.n176 8.45089
R2778 VDD.n412 VDD.n411 8.45089
R2779 VDD.n409 VDD.n180 8.45089
R2780 VDD.n408 VDD.n407 8.45089
R2781 VDD.n399 VDD.n181 8.45089
R2782 VDD.n401 VDD.n400 8.45089
R2783 VDD.n398 VDD.n186 8.45089
R2784 VDD.n396 VDD.n395 8.45089
R2785 VDD.n397 VDD.n396 8.45089
R2786 VDD.n188 VDD.n187 8.45089
R2787 VDD.n371 VDD.t608 8.45089
R2788 VDD.n370 VDD.n192 8.45089
R2789 VDD.n369 VDD.n368 8.45089
R2790 VDD.n194 VDD.n193 8.45089
R2791 VDD.n362 VDD.n361 8.45089
R2792 VDD.n360 VDD.n199 8.45089
R2793 VDD.n359 VDD.n358 8.45089
R2794 VDD.n347 VDD.n200 8.45089
R2795 VDD.n349 VDD.n348 8.45089
R2796 VDD.n346 VDD.n204 8.45089
R2797 VDD.n345 VDD.n344 8.45089
R2798 VDD.n206 VDD.n205 8.45089
R2799 VDD.n336 VDD.n335 8.45089
R2800 VDD.n334 VDD.n210 8.45089
R2801 VDD.n333 VDD.n332 8.45089
R2802 VDD.n321 VDD.n211 8.45089
R2803 VDD.n323 VDD.n322 8.45089
R2804 VDD.n320 VDD.n215 8.45089
R2805 VDD.n319 VDD.n318 8.45089
R2806 VDD.n310 VDD.n216 8.45089
R2807 VDD.n312 VDD.n311 8.45089
R2808 VDD.n309 VDD.n221 8.45089
R2809 VDD.n307 VDD.n306 8.45089
R2810 VDD.n308 VDD.n307 8.45089
R2811 VDD.n223 VDD.n222 8.45089
R2812 VDD.n282 VDD.t468 8.45089
R2813 VDD.n281 VDD.n227 8.45089
R2814 VDD.n280 VDD.n279 8.45089
R2815 VDD.n229 VDD.n228 8.45089
R2816 VDD.n273 VDD.n272 8.45089
R2817 VDD.n271 VDD.n234 8.45089
R2818 VDD.n270 VDD.n269 8.45089
R2819 VDD.n258 VDD.n235 8.45089
R2820 VDD.n260 VDD.n259 8.45089
R2821 VDD.n257 VDD.n239 8.45089
R2822 VDD.n256 VDD.n255 8.45089
R2823 VDD.n241 VDD.n240 8.45089
R2824 VDD.n245 VDD.n244 8.45089
R2825 VDD.n247 VDD.n246 8.45089
R2826 VDD.n2110 VDD.n2109 8.45089
R2827 VDD.n2111 VDD.n2110 8.45089
R2828 VDD.n2113 VDD.n2112 8.45089
R2829 VDD.n2118 VDD.n2117 8.45089
R2830 VDD.n2122 VDD.n2121 8.45089
R2831 VDD.n2127 VDD.n2126 8.45089
R2832 VDD.n2131 VDD.n2130 8.45089
R2833 VDD.n2135 VDD.n2134 8.45089
R2834 VDD.n2140 VDD.n2139 8.45089
R2835 VDD.n2145 VDD.n2144 8.45089
R2836 VDD.n2149 VDD.n2148 8.45089
R2837 VDD.n2155 VDD.n2154 8.45089
R2838 VDD.n2159 VDD.n2158 8.45089
R2839 VDD.n2163 VDD.n2162 8.45089
R2840 VDD.n2166 VDD.t25 8.45089
R2841 VDD.n2170 VDD.n2169 8.45089
R2842 VDD.n2174 VDD.n2173 8.45089
R2843 VDD.n2179 VDD.n2178 8.45089
R2844 VDD.n2184 VDD.n2183 8.45089
R2845 VDD.n2188 VDD.n2187 8.45089
R2846 VDD.n2192 VDD.n2191 8.45089
R2847 VDD.n2210 VDD.n2209 8.45089
R2848 VDD.n2209 VDD.n2208 8.45089
R2849 VDD.n2213 VDD.n2212 8.45089
R2850 VDD.n2218 VDD.n2217 8.45089
R2851 VDD.n11 VDD.n10 8.45089
R2852 VDD.n2226 VDD.n2225 8.45089
R2853 VDD.n2228 VDD.n2227 8.45089
R2854 VDD.n2245 VDD.n2244 8.45089
R2855 VDD.n2250 VDD.n2249 8.45089
R2856 VDD.n2254 VDD.n2253 8.45089
R2857 VDD.n2258 VDD.n2257 8.45089
R2858 VDD.n2284 VDD.n2283 8.45089
R2859 VDD.n2283 VDD.n2282 8.45089
R2860 VDD.n2289 VDD.n2288 8.45089
R2861 VDD.n2293 VDD.n2292 8.45089
R2862 VDD.n2297 VDD.n2296 8.45089
R2863 VDD.n2300 VDD.t523 8.45089
R2864 VDD.n2304 VDD.n2303 8.45089
R2865 VDD.n2308 VDD.n2307 8.45089
R2866 VDD.n2313 VDD.n2312 8.45089
R2867 VDD.n2318 VDD.n2317 8.45089
R2868 VDD.n2322 VDD.n2321 8.45089
R2869 VDD.n2326 VDD.n2325 8.45089
R2870 VDD.n2331 VDD.n2330 8.45089
R2871 VDD.n2335 VDD.n2334 8.45089
R2872 VDD.n2341 VDD.n2340 8.45089
R2873 VDD.n2345 VDD.n2344 8.45089
R2874 VDD.n2350 VDD.n2349 8.45089
R2875 VDD.n7 VDD.n6 8.45089
R2876 VDD.n2358 VDD.n2357 8.45089
R2877 VDD.n2360 VDD.n2359 8.45089
R2878 VDD.n2365 VDD.n2364 8.45089
R2879 VDD.n2369 VDD.n2368 8.45089
R2880 VDD.n2374 VDD.n2373 8.45089
R2881 VDD.n2378 VDD.n2377 8.45089
R2882 VDD.n2382 VDD.n2381 8.45089
R2883 VDD.n2408 VDD.n2407 8.45089
R2884 VDD.n2407 VDD.n2406 8.45089
R2885 VDD.n2413 VDD.n2412 8.45089
R2886 VDD.n2417 VDD.n2416 8.45089
R2887 VDD.n2421 VDD.n2420 8.45089
R2888 VDD.n2424 VDD.t392 8.45089
R2889 VDD.n2428 VDD.n2427 8.45089
R2890 VDD.n2432 VDD.n2431 8.45089
R2891 VDD.n2437 VDD.n2436 8.45089
R2892 VDD.n2442 VDD.n2441 8.45089
R2893 VDD.n2446 VDD.n2445 8.45089
R2894 VDD.n2450 VDD.n2449 8.45089
R2895 VDD.n2455 VDD.n2454 8.45089
R2896 VDD.n2459 VDD.n2458 8.45089
R2897 VDD.n2465 VDD.n2464 8.45089
R2898 VDD.n2469 VDD.n2468 8.45089
R2899 VDD.n2474 VDD.n2473 8.45089
R2900 VDD.n3 VDD.n2 8.45089
R2901 VDD.n2482 VDD.n2481 8.45089
R2902 VDD.n2484 VDD.n2483 8.45089
R2903 VDD.n2489 VDD.n2488 8.45089
R2904 VDD.n2493 VDD.n2492 8.45089
R2905 VDD.n2498 VDD.n2497 8.45089
R2906 VDD.n2502 VDD.n2501 8.45089
R2907 VDD.n2506 VDD.n2505 8.45089
R2908 VDD.n2532 VDD.n2531 8.45089
R2909 VDD.n2531 VDD.n2530 8.45089
R2910 VDD.n2537 VDD.n2536 8.45089
R2911 VDD.n2541 VDD.n2540 8.45089
R2912 VDD.n2545 VDD.n2544 8.45089
R2913 VDD.n2548 VDD.t535 8.45089
R2914 VDD.n2552 VDD.n2551 8.45089
R2915 VDD.n2556 VDD.n2555 8.45089
R2916 VDD.n2561 VDD.n2560 8.45089
R2917 VDD.n2566 VDD.n2565 8.45089
R2918 VDD.n2570 VDD.n2569 8.45089
R2919 VDD.n2574 VDD.n2573 8.45089
R2920 VDD.n2579 VDD.n2578 8.45089
R2921 VDD.n2583 VDD.n2582 8.45089
R2922 VDD.n2589 VDD.n2588 8.45089
R2923 VDD.n2593 VDD.n2592 8.45089
R2924 VDD.n2598 VDD.n2597 8.45089
R2925 VDD.n2729 VDD.n2728 8.45089
R2926 VDD.n2727 VDD.n2726 8.45089
R2927 VDD.n2725 VDD.n2724 8.45089
R2928 VDD.n2716 VDD.n2715 8.45089
R2929 VDD.n2711 VDD.n2710 8.45089
R2930 VDD.n2707 VDD.n2706 8.45089
R2931 VDD.n2703 VDD.n2702 8.45089
R2932 VDD.n2699 VDD.n2698 8.45089
R2933 VDD.n2675 VDD.n2674 8.45089
R2934 VDD.n2674 VDD.n2673 8.45089
R2935 VDD.n2670 VDD.n2669 8.45089
R2936 VDD.n2664 VDD.n2663 8.45089
R2937 VDD.n2660 VDD.n2659 8.45089
R2938 VDD.n2656 VDD.t280 8.45089
R2939 VDD.n2653 VDD.n2652 8.45089
R2940 VDD.n2649 VDD.n2648 8.45089
R2941 VDD.n2644 VDD.n2643 8.45089
R2942 VDD.n2639 VDD.n2638 8.45089
R2943 VDD.n2635 VDD.n2634 8.45089
R2944 VDD.n2630 VDD.n2629 8.45089
R2945 VDD.n2626 VDD.n2625 8.45089
R2946 VDD.n2620 VDD.n2619 8.45089
R2947 VDD.n2616 VDD.n2615 8.45089
R2948 VDD.n2612 VDD.n2611 8.45089
R2949 VDD.n2607 VDD.n2606 8.45089
R2950 VDD.n2604 VDD.n2603 8.45089
R2951 VDD.n2095 VDD.n1992 8.45089
R2952 VDD.n1995 VDD.n1994 8.45089
R2953 VDD.n2086 VDD.n2085 8.45089
R2954 VDD.n2079 VDD.n1998 8.45089
R2955 VDD.n2004 VDD.n1999 8.45089
R2956 VDD.n2075 VDD.n2074 8.45089
R2957 VDD.n2001 VDD.n2000 8.45089
R2958 VDD.n2069 VDD.n2068 8.45089
R2959 VDD.n2009 VDD.n2006 8.45089
R2960 VDD.n2063 VDD.n2062 8.45089
R2961 VDD.n2012 VDD.n2011 8.45089
R2962 VDD.n2015 VDD.n2014 8.45089
R2963 VDD.n2052 VDD.n2051 8.45089
R2964 VDD.n2017 VDD.n2016 8.45089
R2965 VDD.n2047 VDD.n2046 8.45089
R2966 VDD.n2024 VDD.n2021 8.45089
R2967 VDD.n2041 VDD.n2040 8.45089
R2968 VDD.n2023 VDD.n2022 8.45089
R2969 VDD.n2036 VDD.n2035 8.45089
R2970 VDD.n2031 VDD.n2030 8.45089
R2971 VDD.n1979 VDD.n1978 8.45089
R2972 VDD.n1410 VDD.n1409 8.45089
R2973 VDD.n1974 VDD.n1973 8.45089
R2974 VDD.n1417 VDD.n1414 8.45089
R2975 VDD.n1969 VDD.n1968 8.45089
R2976 VDD.n1965 VDD.n1415 8.45089
R2977 VDD.n1964 VDD.n1963 8.45089
R2978 VDD.n1958 VDD.n1957 8.45089
R2979 VDD.n1423 VDD.n1422 8.45089
R2980 VDD.n1950 VDD.n1949 8.45089
R2981 VDD.n1426 VDD.n1425 8.45089
R2982 VDD.n1946 VDD.n1945 8.45089
R2983 VDD.n1942 VDD.n1428 8.45089
R2984 VDD.n1941 VDD.n1940 8.45089
R2985 VDD.n1433 VDD.n1432 8.45089
R2986 VDD.n1435 VDD.n1434 8.45089
R2987 VDD.n1928 VDD.n1927 8.45089
R2988 VDD.n1438 VDD.n1437 8.45089
R2989 VDD.n1441 VDD.n1440 8.45089
R2990 VDD.n1444 VDD.n1443 8.45089
R2991 VDD.n1910 VDD.n1909 8.45089
R2992 VDD.n1902 VDD.n1901 8.45089
R2993 VDD.n1449 VDD.n1448 8.45089
R2994 VDD.n1896 VDD.n1895 8.45089
R2995 VDD.n1892 VDD.n1450 8.45089
R2996 VDD.n1891 VDD.n1890 8.45089
R2997 VDD.n1458 VDD.n1455 8.45089
R2998 VDD.n1885 VDD.n1884 8.45089
R2999 VDD.n1877 VDD.n1876 8.45089
R3000 VDD.n1461 VDD.n1460 8.45089
R3001 VDD.n1872 VDD.n1871 8.45089
R3002 VDD.n1464 VDD.n1463 8.45089
R3003 VDD.n1867 VDD.n1866 8.45089
R3004 VDD.n1472 VDD.n1468 8.45089
R3005 VDD.n1862 VDD.n1861 8.45089
R3006 VDD.n1471 VDD.n1470 8.45089
R3007 VDD.n1476 VDD.n1475 8.45089
R3008 VDD.n1851 VDD.n1850 8.45089
R3009 VDD.n1478 VDD.n1477 8.45089
R3010 VDD.n1481 VDD.n1480 8.45089
R3011 VDD.n1483 VDD.n1482 8.45089
R3012 VDD.n1832 VDD.n1831 8.45089
R3013 VDD.n1826 VDD.n1825 8.45089
R3014 VDD.n1491 VDD.n1490 8.45089
R3015 VDD.n1821 VDD.n1820 8.45089
R3016 VDD.n1498 VDD.n1495 8.45089
R3017 VDD.n1816 VDD.n1815 8.45089
R3018 VDD.n1812 VDD.n1496 8.45089
R3019 VDD.n1811 VDD.n1810 8.45089
R3020 VDD.n1805 VDD.n1804 8.45089
R3021 VDD.n1504 VDD.n1503 8.45089
R3022 VDD.n1797 VDD.n1796 8.45089
R3023 VDD.n1507 VDD.n1506 8.45089
R3024 VDD.n1793 VDD.n1792 8.45089
R3025 VDD.n1789 VDD.n1509 8.45089
R3026 VDD.n1788 VDD.n1787 8.45089
R3027 VDD.n1514 VDD.n1513 8.45089
R3028 VDD.n1516 VDD.n1515 8.45089
R3029 VDD.n1775 VDD.n1774 8.45089
R3030 VDD.n1519 VDD.n1518 8.45089
R3031 VDD.n1522 VDD.n1521 8.45089
R3032 VDD.n1525 VDD.n1524 8.45089
R3033 VDD.n1757 VDD.n1756 8.45089
R3034 VDD.n1749 VDD.n1748 8.45089
R3035 VDD.n1530 VDD.n1529 8.45089
R3036 VDD.n1743 VDD.n1742 8.45089
R3037 VDD.n1739 VDD.n1531 8.45089
R3038 VDD.n1738 VDD.n1737 8.45089
R3039 VDD.n1539 VDD.n1536 8.45089
R3040 VDD.n1732 VDD.n1731 8.45089
R3041 VDD.n1724 VDD.n1723 8.45089
R3042 VDD.n1542 VDD.n1541 8.45089
R3043 VDD.n1719 VDD.n1718 8.45089
R3044 VDD.n1545 VDD.n1544 8.45089
R3045 VDD.n1714 VDD.n1713 8.45089
R3046 VDD.n1553 VDD.n1549 8.45089
R3047 VDD.n1709 VDD.n1708 8.45089
R3048 VDD.n1552 VDD.n1551 8.45089
R3049 VDD.n1557 VDD.n1556 8.45089
R3050 VDD.n1698 VDD.n1697 8.45089
R3051 VDD.n1559 VDD.n1558 8.45089
R3052 VDD.n1562 VDD.n1561 8.45089
R3053 VDD.n1564 VDD.n1563 8.45089
R3054 VDD.n1679 VDD.n1678 8.45089
R3055 VDD.n1673 VDD.n1672 8.45089
R3056 VDD.n1572 VDD.n1571 8.45089
R3057 VDD.n1668 VDD.n1667 8.45089
R3058 VDD.n1579 VDD.n1576 8.45089
R3059 VDD.n1663 VDD.n1662 8.45089
R3060 VDD.n1659 VDD.n1577 8.45089
R3061 VDD.n1658 VDD.n1657 8.45089
R3062 VDD.n1652 VDD.n1651 8.45089
R3063 VDD.n1585 VDD.n1584 8.45089
R3064 VDD.n1644 VDD.n1643 8.45089
R3065 VDD.n1588 VDD.n1587 8.45089
R3066 VDD.n1640 VDD.n1639 8.45089
R3067 VDD.n1636 VDD.n1590 8.45089
R3068 VDD.n1635 VDD.n1634 8.45089
R3069 VDD.n1595 VDD.n1594 8.45089
R3070 VDD.n1597 VDD.n1596 8.45089
R3071 VDD.n1622 VDD.n1621 8.45089
R3072 VDD.n1600 VDD.n1599 8.45089
R3073 VDD.n1603 VDD.n1602 8.45089
R3074 VDD.n770 VDD.n767 8.45089
R3075 VDD.n1396 VDD.n1395 8.45089
R3076 VDD.n1243 VDD.n1242 8.45089
R3077 VDD.n851 VDD.n850 8.45089
R3078 VDD.n1233 VDD.n1232 8.45089
R3079 VDD.n855 VDD.n854 8.45089
R3080 VDD.n1228 VDD.n1225 8.45089
R3081 VDD.n859 VDD.n858 8.45089
R3082 VDD.n1221 VDD.n1220 8.45089
R3083 VDD.n1214 VDD.n1213 8.45089
R3084 VDD.n863 VDD.n862 8.45089
R3085 VDD.n865 VDD.n864 8.45089
R3086 VDD.n868 VDD.n867 8.45089
R3087 VDD.n1193 VDD.n1192 8.45089
R3088 VDD.n870 VDD.n869 8.45089
R3089 VDD.n874 VDD.n873 8.45089
R3090 VDD.n1181 VDD.n1180 8.45089
R3091 VDD.n876 VDD.n875 8.45089
R3092 VDD.n1176 VDD.n1173 8.45089
R3093 VDD.n879 VDD.n878 8.45089
R3094 VDD.n1169 VDD.n1168 8.45089
R3095 VDD.n881 VDD.n880 8.45089
R3096 VDD.n1164 VDD.n1163 8.45089
R3097 VDD.n1158 VDD.n1157 8.45089
R3098 VDD.n888 VDD.n887 8.45089
R3099 VDD.n1153 VDD.n1151 8.45089
R3100 VDD.n891 VDD.n890 8.45089
R3101 VDD.n1146 VDD.n1145 8.45089
R3102 VDD.n893 VDD.n892 8.45089
R3103 VDD.n1141 VDD.n1140 8.45089
R3104 VDD.n1135 VDD.n1134 8.45089
R3105 VDD.n902 VDD.n901 8.45089
R3106 VDD.n906 VDD.n905 8.45089
R3107 VDD.n908 VDD.n907 8.45089
R3108 VDD.n1117 VDD.n1116 8.45089
R3109 VDD.n911 VDD.n910 8.45089
R3110 VDD.n913 VDD.n912 8.45089
R3111 VDD.n1104 VDD.n1103 8.45089
R3112 VDD.n916 VDD.n915 8.45089
R3113 VDD.n1098 VDD.n1097 8.45089
R3114 VDD.n918 VDD.n917 8.45089
R3115 VDD.n1093 VDD.n1092 8.45089
R3116 VDD.n923 VDD.n922 8.45089
R3117 VDD.n1088 VDD.n1087 8.45089
R3118 VDD.n1081 VDD.n1080 8.45089
R3119 VDD.n928 VDD.n927 8.45089
R3120 VDD.n1075 VDD.n1074 8.45089
R3121 VDD.n931 VDD.n930 8.45089
R3122 VDD.n1070 VDD.n1067 8.45089
R3123 VDD.n935 VDD.n934 8.45089
R3124 VDD.n1063 VDD.n1062 8.45089
R3125 VDD.n1056 VDD.n1055 8.45089
R3126 VDD.n939 VDD.n938 8.45089
R3127 VDD.n941 VDD.n940 8.45089
R3128 VDD.n944 VDD.n943 8.45089
R3129 VDD.n1035 VDD.n1034 8.45089
R3130 VDD.n946 VDD.n945 8.45089
R3131 VDD.n950 VDD.n949 8.45089
R3132 VDD.n1023 VDD.n1022 8.45089
R3133 VDD.n952 VDD.n951 8.45089
R3134 VDD.n1018 VDD.n1015 8.45089
R3135 VDD.n955 VDD.n954 8.45089
R3136 VDD.n1011 VDD.n1010 8.45089
R3137 VDD.n957 VDD.n956 8.45089
R3138 VDD.n1006 VDD.n1005 8.45089
R3139 VDD.n1000 VDD.n999 8.45089
R3140 VDD.n964 VDD.n963 8.45089
R3141 VDD.n995 VDD.n993 8.45089
R3142 VDD.n967 VDD.n966 8.45089
R3143 VDD.n988 VDD.n987 8.45089
R3144 VDD.n969 VDD.n968 8.45089
R3145 VDD.n983 VDD.n982 8.45089
R3146 VDD.n758 VDD.n757 8.45089
R3147 VDD.n754 VDD.n17 8.45089
R3148 VDD.n753 VDD.n752 8.45089
R3149 VDD.n745 VDD.n21 8.45089
R3150 VDD.n23 VDD.n22 8.45089
R3151 VDD.n740 VDD.n738 8.45089
R3152 VDD.n636 VDD.n86 8.45089
R3153 VDD.n628 VDD.n627 8.45089
R3154 VDD.n625 VDD.n88 8.45089
R3155 VDD.n94 VDD.n90 8.45089
R3156 VDD.n621 VDD.n618 8.45089
R3157 VDD.n93 VDD.n92 8.45089
R3158 VDD.n612 VDD.n611 8.45089
R3159 VDD.n96 VDD.n95 8.45089
R3160 VDD.n607 VDD.n604 8.45089
R3161 VDD.n101 VDD.n100 8.45089
R3162 VDD.n599 VDD.n598 8.45089
R3163 VDD.n104 VDD.n103 8.45089
R3164 VDD.n592 VDD.n591 8.45089
R3165 VDD.n110 VDD.n109 8.45089
R3166 VDD.n586 VDD.n585 8.45089
R3167 VDD.n581 VDD.n111 8.45089
R3168 VDD.n580 VDD.n579 8.45089
R3169 VDD.n567 VDD.n116 8.45089
R3170 VDD.n119 VDD.n118 8.45089
R3171 VDD.n550 VDD.n549 8.45089
R3172 VDD.n122 VDD.n121 8.45089
R3173 VDD.n546 VDD.n545 8.45089
R3174 VDD.n542 VDD.n124 8.45089
R3175 VDD.n541 VDD.n540 8.45089
R3176 VDD.n129 VDD.n128 8.45089
R3177 VDD.n131 VDD.n130 8.45089
R3178 VDD.n528 VDD.n527 8.45089
R3179 VDD.n134 VDD.n133 8.45089
R3180 VDD.n137 VDD.n136 8.45089
R3181 VDD.n140 VDD.n139 8.45089
R3182 VDD.n510 VDD.n509 8.45089
R3183 VDD.n502 VDD.n501 8.45089
R3184 VDD.n145 VDD.n144 8.45089
R3185 VDD.n496 VDD.n495 8.45089
R3186 VDD.n492 VDD.n146 8.45089
R3187 VDD.n491 VDD.n490 8.45089
R3188 VDD.n478 VDD.n151 8.45089
R3189 VDD.n154 VDD.n153 8.45089
R3190 VDD.n461 VDD.n460 8.45089
R3191 VDD.n157 VDD.n156 8.45089
R3192 VDD.n457 VDD.n456 8.45089
R3193 VDD.n453 VDD.n159 8.45089
R3194 VDD.n452 VDD.n451 8.45089
R3195 VDD.n164 VDD.n163 8.45089
R3196 VDD.n166 VDD.n165 8.45089
R3197 VDD.n439 VDD.n438 8.45089
R3198 VDD.n169 VDD.n168 8.45089
R3199 VDD.n172 VDD.n171 8.45089
R3200 VDD.n175 VDD.n174 8.45089
R3201 VDD.n421 VDD.n420 8.45089
R3202 VDD.n413 VDD.n412 8.45089
R3203 VDD.n180 VDD.n179 8.45089
R3204 VDD.n407 VDD.n406 8.45089
R3205 VDD.n403 VDD.n181 8.45089
R3206 VDD.n402 VDD.n401 8.45089
R3207 VDD.n389 VDD.n186 8.45089
R3208 VDD.n189 VDD.n188 8.45089
R3209 VDD.n372 VDD.n371 8.45089
R3210 VDD.n192 VDD.n191 8.45089
R3211 VDD.n368 VDD.n367 8.45089
R3212 VDD.n364 VDD.n194 8.45089
R3213 VDD.n363 VDD.n362 8.45089
R3214 VDD.n199 VDD.n198 8.45089
R3215 VDD.n201 VDD.n200 8.45089
R3216 VDD.n350 VDD.n349 8.45089
R3217 VDD.n204 VDD.n203 8.45089
R3218 VDD.n207 VDD.n206 8.45089
R3219 VDD.n210 VDD.n209 8.45089
R3220 VDD.n332 VDD.n331 8.45089
R3221 VDD.n324 VDD.n323 8.45089
R3222 VDD.n215 VDD.n214 8.45089
R3223 VDD.n318 VDD.n317 8.45089
R3224 VDD.n314 VDD.n216 8.45089
R3225 VDD.n313 VDD.n312 8.45089
R3226 VDD.n300 VDD.n221 8.45089
R3227 VDD.n224 VDD.n223 8.45089
R3228 VDD.n283 VDD.n282 8.45089
R3229 VDD.n227 VDD.n226 8.45089
R3230 VDD.n279 VDD.n278 8.45089
R3231 VDD.n275 VDD.n229 8.45089
R3232 VDD.n274 VDD.n273 8.45089
R3233 VDD.n234 VDD.n233 8.45089
R3234 VDD.n236 VDD.n235 8.45089
R3235 VDD.n261 VDD.n260 8.45089
R3236 VDD.n239 VDD.n238 8.45089
R3237 VDD.n242 VDD.n241 8.45089
R3238 VDD.n2119 VDD.n2118 8.45089
R3239 VDD.n2128 VDD.n2127 8.45089
R3240 VDD.n2132 VDD.n2131 8.45089
R3241 VDD.n2136 VDD.n2135 8.45089
R3242 VDD.n2146 VDD.n2145 8.45089
R3243 VDD.n2150 VDD.n2149 8.45089
R3244 VDD.n2156 VDD.n2155 8.45089
R3245 VDD.n2160 VDD.n2159 8.45089
R3246 VDD.n2164 VDD.n2163 8.45089
R3247 VDD.n2167 VDD.n2166 8.45089
R3248 VDD.n2171 VDD.n2170 8.45089
R3249 VDD.n2175 VDD.n2174 8.45089
R3250 VDD.n2185 VDD.n2184 8.45089
R3251 VDD.n2189 VDD.n2188 8.45089
R3252 VDD.n2194 VDD.n2192 8.45089
R3253 VDD.n2214 VDD.n2213 8.45089
R3254 VDD.n2223 VDD.n11 8.45089
R3255 VDD.n2225 VDD.n2224 8.45089
R3256 VDD.n2251 VDD.n2250 8.45089
R3257 VDD.n2255 VDD.n2254 8.45089
R3258 VDD.n2259 VDD.n2258 8.45089
R3259 VDD.n2290 VDD.n2289 8.45089
R3260 VDD.n2294 VDD.n2293 8.45089
R3261 VDD.n2298 VDD.n2297 8.45089
R3262 VDD.n2301 VDD.n2300 8.45089
R3263 VDD.n2305 VDD.n2304 8.45089
R3264 VDD.n2309 VDD.n2308 8.45089
R3265 VDD.n2319 VDD.n2318 8.45089
R3266 VDD.n2323 VDD.n2322 8.45089
R3267 VDD.n2328 VDD.n2326 8.45089
R3268 VDD.n2332 VDD.n2331 8.45089
R3269 VDD.n2338 VDD.n2335 8.45089
R3270 VDD.n2342 VDD.n2341 8.45089
R3271 VDD.n2346 VDD.n2345 8.45089
R3272 VDD.n2355 VDD.n7 8.45089
R3273 VDD.n2357 VDD.n2356 8.45089
R3274 VDD.n2366 VDD.n2365 8.45089
R3275 VDD.n2375 VDD.n2374 8.45089
R3276 VDD.n2379 VDD.n2378 8.45089
R3277 VDD.n2383 VDD.n2382 8.45089
R3278 VDD.n2414 VDD.n2413 8.45089
R3279 VDD.n2418 VDD.n2417 8.45089
R3280 VDD.n2422 VDD.n2421 8.45089
R3281 VDD.n2425 VDD.n2424 8.45089
R3282 VDD.n2429 VDD.n2428 8.45089
R3283 VDD.n2433 VDD.n2432 8.45089
R3284 VDD.n2443 VDD.n2442 8.45089
R3285 VDD.n2447 VDD.n2446 8.45089
R3286 VDD.n2452 VDD.n2450 8.45089
R3287 VDD.n2456 VDD.n2455 8.45089
R3288 VDD.n2462 VDD.n2459 8.45089
R3289 VDD.n2466 VDD.n2465 8.45089
R3290 VDD.n2470 VDD.n2469 8.45089
R3291 VDD.n2479 VDD.n3 8.45089
R3292 VDD.n2481 VDD.n2480 8.45089
R3293 VDD.n2490 VDD.n2489 8.45089
R3294 VDD.n2499 VDD.n2498 8.45089
R3295 VDD.n2503 VDD.n2502 8.45089
R3296 VDD.n2507 VDD.n2506 8.45089
R3297 VDD.n2538 VDD.n2537 8.45089
R3298 VDD.n2542 VDD.n2541 8.45089
R3299 VDD.n2546 VDD.n2545 8.45089
R3300 VDD.n2549 VDD.n2548 8.45089
R3301 VDD.n2553 VDD.n2552 8.45089
R3302 VDD.n2557 VDD.n2556 8.45089
R3303 VDD.n2567 VDD.n2566 8.45089
R3304 VDD.n2571 VDD.n2570 8.45089
R3305 VDD.n2576 VDD.n2574 8.45089
R3306 VDD.n2580 VDD.n2579 8.45089
R3307 VDD.n2586 VDD.n2583 8.45089
R3308 VDD.n2590 VDD.n2589 8.45089
R3309 VDD.n2594 VDD.n2593 8.45089
R3310 VDD.n2730 VDD.n2729 8.45089
R3311 VDD.n2726 VDD.n2602 8.45089
R3312 VDD.n2717 VDD.n2716 8.45089
R3313 VDD.n2708 VDD.n2707 8.45089
R3314 VDD.n2704 VDD.n2703 8.45089
R3315 VDD.n2700 VDD.n2699 8.45089
R3316 VDD.n2671 VDD.n2670 8.45089
R3317 VDD.n2665 VDD.n2664 8.45089
R3318 VDD.n2661 VDD.n2660 8.45089
R3319 VDD.n2657 VDD.n2656 8.45089
R3320 VDD.n2654 VDD.n2653 8.45089
R3321 VDD.n2650 VDD.n2649 8.45089
R3322 VDD.n2640 VDD.n2639 8.45089
R3323 VDD.n2636 VDD.n2635 8.45089
R3324 VDD.n2632 VDD.n2630 8.45089
R3325 VDD.n2627 VDD.n2626 8.45089
R3326 VDD.n2623 VDD.n2620 8.45089
R3327 VDD.n2617 VDD.n2616 8.45089
R3328 VDD.n2613 VDD.n2612 8.45089
R3329 VDD.n1579 VDD.n1575 8.31095
R3330 VDD.n1739 VDD.n1533 8.31095
R3331 VDD.n1498 VDD.n1494 8.31095
R3332 VDD.n1892 VDD.n1452 8.31095
R3333 VDD.n1417 VDD.n1413 8.31095
R3334 VDD.n971 VDD.n966 8.31095
R3335 VDD.n1069 VDD.n931 8.31095
R3336 VDD.n895 VDD.n890 8.31095
R3337 VDD.n1227 VDD.n855 8.31095
R3338 VDD.n581 VDD.n113 8.31095
R3339 VDD.n492 VDD.n148 8.31095
R3340 VDD.n403 VDD.n183 8.31095
R3341 VDD.n314 VDD.n218 8.31095
R3342 VDD.n2024 VDD.n2020 8.16602
R3343 VDD.n2057 VDD.n2012 8.16602
R3344 VDD.n2680 VDD.n2679 8.00414
R3345 VDD.n2516 VDD.n2515 8.00414
R3346 VDD.n2392 VDD.n2391 8.00414
R3347 VDD.n2268 VDD.n2267 8.00414
R3348 VDD.n1633 VDD.t202 7.91717
R3349 VDD.t528 VDD.n1710 7.91717
R3350 VDD.n1786 VDD.t201 7.91717
R3351 VDD.t437 VDD.n1863 7.91717
R3352 VDD.n1939 VDD.t121 7.91717
R3353 VDD.n2673 VDD.t28 7.89524
R3354 VDD.n2530 VDD.t78 7.89524
R3355 VDD.n2406 VDD.t538 7.89524
R3356 VDD.n2282 VDD.t264 7.89524
R3357 VDD.n2148 VDD.t124 7.89524
R3358 VDD.n272 VDD.t29 7.80872
R3359 VDD.n361 VDD.t456 7.80872
R3360 VDD.n450 VDD.t388 7.80872
R3361 VDD.n539 VDD.t642 7.80872
R3362 VDD.n695 VDD.t298 7.80872
R3363 VDD.n1024 VDD.t83 7.74507
R3364 VDD.n1102 VDD.t533 7.74507
R3365 VDD.n1182 VDD.t314 7.74507
R3366 VDD.t195 VDD.n1398 7.74507
R3367 VDD.n678 VDD.n677 7.72464
R3368 VDD.n1297 VDD.n820 7.70756
R3369 VDD.n2688 VDD.n2687 6.95412
R3370 VDD.n2524 VDD.n2523 6.95412
R3371 VDD.n2400 VDD.n2399 6.95412
R3372 VDD.n2276 VDD.n2275 6.95412
R3373 VDD.n1366 VDD.n782 6.84188
R3374 VDD.n1381 VDD.n772 6.84188
R3375 VDD.n606 VDD.n96 6.62119
R3376 VDD.n621 VDD.n620 6.62119
R3377 VDD.n1382 VDD.n1381 6.33153
R3378 VDD.n1366 VDD.n786 6.32841
R3379 VDD.n1248 VDD.n848 6.32433
R3380 VDD.n1329 VDD.n1328 6.32433
R3381 VDD.n739 VDD.n23 5.51774
R3382 VDD.n1629 VDD.n1594 5.29705
R3383 VDD.n1703 VDD.n1552 5.29705
R3384 VDD.n1782 VDD.n1513 5.29705
R3385 VDD.n1856 VDD.n1471 5.29705
R3386 VDD.n1935 VDD.n1432 5.29705
R3387 VDD.n1029 VDD.n949 5.29705
R3388 VDD.n1110 VDD.n913 5.29705
R3389 VDD.n1187 VDD.n873 5.29705
R3390 VDD.n535 VDD.n128 5.29705
R3391 VDD.n446 VDD.n163 5.29705
R3392 VDD.n357 VDD.n198 5.29705
R3393 VDD.n268 VDD.n233 5.29705
R3394 VDD.n683 VDD.t300 5.20598
R3395 VDD.n679 VDD.n678 5.07636
R3396 VDD.n294 VDD 5.04292
R3397 VDD.n383 VDD 5.04292
R3398 VDD.n472 VDD 5.04292
R3399 VDD.n561 VDD 5.04292
R3400 VDD.n841 VDD.n840 4.6505
R3401 VDD.n1261 VDD.n839 4.6505
R3402 VDD.n1273 VDD.n831 4.6505
R3403 VDD.n1283 VDD.n826 4.6505
R3404 VDD.n1286 VDD.n825 4.6505
R3405 VDD.n1302 VDD.n817 4.6505
R3406 VDD.n1312 VDD.n812 4.6505
R3407 VDD.n1316 VDD.n811 4.6505
R3408 VDD.n1339 VDD.n799 4.6505
R3409 VDD.n1349 VDD.n794 4.6505
R3410 VDD.n1353 VDD.n793 4.6505
R3411 VDD.n1369 VDD.n783 4.6505
R3412 VDD.n1392 VDD.n1391 4.6505
R3413 VDD.n304 VDD.n303 4.6505
R3414 VDD.n302 VDD.n301 4.6505
R3415 VDD.n393 VDD.n392 4.6505
R3416 VDD.n391 VDD.n390 4.6505
R3417 VDD.n482 VDD.n481 4.6505
R3418 VDD.n480 VDD.n479 4.6505
R3419 VDD.n571 VDD.n570 4.6505
R3420 VDD.n569 VDD.n568 4.6505
R3421 VDD.n648 VDD.n76 4.6505
R3422 VDD.n70 VDD.n69 4.6505
R3423 VDD.n663 VDD.n68 4.6505
R3424 VDD.n675 VDD.n60 4.6505
R3425 VDD.n686 VDD.n54 4.6505
R3426 VDD.n48 VDD.n47 4.6505
R3427 VDD.n701 VDD.n46 4.6505
R3428 VDD.n713 VDD.n38 4.6505
R3429 VDD.n724 VDD.n32 4.6505
R3430 VDD.n729 VDD.n728 4.6505
R3431 VDD.n2692 VDD.n2691 4.6505
R3432 VDD.n2697 VDD.n2696 4.6505
R3433 VDD.n2528 VDD.n2527 4.6505
R3434 VDD.n2512 VDD.n2511 4.6505
R3435 VDD.n2404 VDD.n2403 4.6505
R3436 VDD.n2388 VDD.n2387 4.6505
R3437 VDD.n2280 VDD.n2279 4.6505
R3438 VDD.n2264 VDD.n2263 4.6505
R3439 VDD.n2207 VDD.n2206 4.6505
R3440 VDD.n2202 VDD.n2201 4.6505
R3441 VDD.n2680 VDD 4.55532
R3442 VDD.n2516 VDD 4.55532
R3443 VDD.n2392 VDD 4.55532
R3444 VDD.n2268 VDD 4.55532
R3445 VDD.n2685 VDD.n2684 4.46483
R3446 VDD.n2521 VDD.n2520 4.46483
R3447 VDD.n2397 VDD.n2396 4.46483
R3448 VDD.n2273 VDD.n2272 4.46483
R3449 VDD.n1247 VDD.n846 4.44959
R3450 VDD.n1327 VDD.n1326 4.44959
R3451 VDD.n1365 VDD.n784 4.43314
R3452 VDD.n1380 VDD.n1379 4.42059
R3453 VDD.n699 VDD.n698 4.1936
R3454 VDD.n2095 VDD 3.75222
R3455 VDD.n635 VDD.n82 3.75222
R3456 VDD.n763 VDD 3.75222
R3457 VDD.n2242 VDD.n2241 3.75222
R3458 VDD.n1639 VDD.n1592 3.53153
R3459 VDD.n1714 VDD.n1548 3.53153
R3460 VDD.n1792 VDD.n1511 3.53153
R3461 VDD.n1867 VDD.n1467 3.53153
R3462 VDD.n1945 VDD.n1430 3.53153
R3463 VDD.n1018 VDD.n1017 3.53153
R3464 VDD.n1097 VDD.n920 3.53153
R3465 VDD.n1176 VDD.n1175 3.53153
R3466 VDD.n1328 VDD.n805 3.53153
R3467 VDD.n754 VDD 3.53153
R3468 VDD.n545 VDD.n126 3.53153
R3469 VDD.n456 VDD.n161 3.53153
R3470 VDD.n367 VDD.n196 3.53153
R3471 VDD.n278 VDD.n231 3.53153
R3472 VDD.n2234 VDD.n2233 3.53153
R3473 VDD.n2240 VDD.n2236 3.52991
R3474 VDD.n977 VDD.n972 3.22029
R3475 VDD.n2610 VDD.n2604 3.22029
R3476 VDD.n2030 VDD 3.12394
R3477 VDD.n1608 VDD 3.12394
R3478 VDD.n247 VDD 3.12394
R3479 VDD.n289 VDD 3.10353
R3480 VDD.n378 VDD 3.10353
R3481 VDD.n467 VDD 3.10353
R3482 VDD.n556 VDD 3.10353
R3483 VDD.n2105 VDD.n2104 3.1005
R3484 VDD.n2098 VDD.n2097 3.1005
R3485 VDD.n2082 VDD.n2081 3.1005
R3486 VDD.n2037 VDD.n2036 3.1005
R3487 VDD.n2038 VDD.n2023 3.1005
R3488 VDD.n2040 VDD.n2039 3.1005
R3489 VDD.n2024 VDD.n2018 3.1005
R3490 VDD.n2048 VDD.n2047 3.1005
R3491 VDD.n2049 VDD.n2017 3.1005
R3492 VDD.n2051 VDD.n2050 3.1005
R3493 VDD.n2014 VDD.n2013 3.1005
R3494 VDD.n2060 VDD.n2012 3.1005
R3495 VDD.n2062 VDD.n2061 3.1005
R3496 VDD.n2006 VDD.n2005 3.1005
R3497 VDD.n2070 VDD.n2069 3.1005
R3498 VDD.n2071 VDD.n2001 3.1005
R3499 VDD.n2074 VDD.n2073 3.1005
R3500 VDD.n2072 VDD.n2004 3.1005
R3501 VDD.n1998 VDD.n1997 3.1005
R3502 VDD.n2085 VDD.n2084 3.1005
R3503 VDD.n2083 VDD.n1994 3.1005
R3504 VDD.n2096 VDD.n2095 3.1005
R3505 VDD.n1984 VDD.n1983 3.1005
R3506 VDD.n1612 VDD.n1603 3.1005
R3507 VDD.n1599 VDD.n1598 3.1005
R3508 VDD.n1623 VDD.n1622 3.1005
R3509 VDD.n1624 VDD.n1597 3.1005
R3510 VDD.n1625 VDD.n1594 3.1005
R3511 VDD.n1635 VDD.n1593 3.1005
R3512 VDD.n1637 VDD.n1636 3.1005
R3513 VDD.n1639 VDD.n1638 3.1005
R3514 VDD.n1587 VDD.n1586 3.1005
R3515 VDD.n1645 VDD.n1644 3.1005
R3516 VDD.n1646 VDD.n1585 3.1005
R3517 VDD.n1651 VDD.n1650 3.1005
R3518 VDD.n1658 VDD.n1580 3.1005
R3519 VDD.n1660 VDD.n1659 3.1005
R3520 VDD.n1662 VDD.n1661 3.1005
R3521 VDD.n1579 VDD.n1573 3.1005
R3522 VDD.n1669 VDD.n1668 3.1005
R3523 VDD.n1670 VDD.n1572 3.1005
R3524 VDD.n1672 VDD.n1671 3.1005
R3525 VDD.n1680 VDD.n1679 3.1005
R3526 VDD.n1681 VDD.n1564 3.1005
R3527 VDD.n1561 VDD.n1560 3.1005
R3528 VDD.n1695 VDD.n1559 3.1005
R3529 VDD.n1697 VDD.n1696 3.1005
R3530 VDD.n1556 VDD.n1554 3.1005
R3531 VDD.n1706 VDD.n1552 3.1005
R3532 VDD.n1708 VDD.n1707 3.1005
R3533 VDD.n1553 VDD.n1546 3.1005
R3534 VDD.n1715 VDD.n1714 3.1005
R3535 VDD.n1716 VDD.n1545 3.1005
R3536 VDD.n1718 VDD.n1717 3.1005
R3537 VDD.n1541 VDD.n1540 3.1005
R3538 VDD.n1725 VDD.n1724 3.1005
R3539 VDD.n1731 VDD.n1730 3.1005
R3540 VDD.n1729 VDD.n1539 3.1005
R3541 VDD.n1738 VDD.n1534 3.1005
R3542 VDD.n1740 VDD.n1739 3.1005
R3543 VDD.n1742 VDD.n1741 3.1005
R3544 VDD.n1529 VDD.n1528 3.1005
R3545 VDD.n1750 VDD.n1749 3.1005
R3546 VDD.n1756 VDD.n1755 3.1005
R3547 VDD.n1754 VDD.n1524 3.1005
R3548 VDD.n1765 VDD.n1522 3.1005
R3549 VDD.n1518 VDD.n1517 3.1005
R3550 VDD.n1776 VDD.n1775 3.1005
R3551 VDD.n1777 VDD.n1516 3.1005
R3552 VDD.n1778 VDD.n1513 3.1005
R3553 VDD.n1788 VDD.n1512 3.1005
R3554 VDD.n1790 VDD.n1789 3.1005
R3555 VDD.n1792 VDD.n1791 3.1005
R3556 VDD.n1506 VDD.n1505 3.1005
R3557 VDD.n1798 VDD.n1797 3.1005
R3558 VDD.n1799 VDD.n1504 3.1005
R3559 VDD.n1804 VDD.n1803 3.1005
R3560 VDD.n1811 VDD.n1499 3.1005
R3561 VDD.n1813 VDD.n1812 3.1005
R3562 VDD.n1815 VDD.n1814 3.1005
R3563 VDD.n1498 VDD.n1492 3.1005
R3564 VDD.n1822 VDD.n1821 3.1005
R3565 VDD.n1823 VDD.n1491 3.1005
R3566 VDD.n1825 VDD.n1824 3.1005
R3567 VDD.n1833 VDD.n1832 3.1005
R3568 VDD.n1834 VDD.n1483 3.1005
R3569 VDD.n1480 VDD.n1479 3.1005
R3570 VDD.n1848 VDD.n1478 3.1005
R3571 VDD.n1850 VDD.n1849 3.1005
R3572 VDD.n1475 VDD.n1473 3.1005
R3573 VDD.n1859 VDD.n1471 3.1005
R3574 VDD.n1861 VDD.n1860 3.1005
R3575 VDD.n1472 VDD.n1465 3.1005
R3576 VDD.n1868 VDD.n1867 3.1005
R3577 VDD.n1869 VDD.n1464 3.1005
R3578 VDD.n1871 VDD.n1870 3.1005
R3579 VDD.n1460 VDD.n1459 3.1005
R3580 VDD.n1878 VDD.n1877 3.1005
R3581 VDD.n1884 VDD.n1883 3.1005
R3582 VDD.n1882 VDD.n1458 3.1005
R3583 VDD.n1891 VDD.n1453 3.1005
R3584 VDD.n1893 VDD.n1892 3.1005
R3585 VDD.n1895 VDD.n1894 3.1005
R3586 VDD.n1448 VDD.n1447 3.1005
R3587 VDD.n1903 VDD.n1902 3.1005
R3588 VDD.n1909 VDD.n1908 3.1005
R3589 VDD.n1907 VDD.n1443 3.1005
R3590 VDD.n1918 VDD.n1441 3.1005
R3591 VDD.n1437 VDD.n1436 3.1005
R3592 VDD.n1929 VDD.n1928 3.1005
R3593 VDD.n1930 VDD.n1435 3.1005
R3594 VDD.n1931 VDD.n1432 3.1005
R3595 VDD.n1941 VDD.n1431 3.1005
R3596 VDD.n1943 VDD.n1942 3.1005
R3597 VDD.n1945 VDD.n1944 3.1005
R3598 VDD.n1425 VDD.n1424 3.1005
R3599 VDD.n1951 VDD.n1950 3.1005
R3600 VDD.n1952 VDD.n1423 3.1005
R3601 VDD.n1957 VDD.n1956 3.1005
R3602 VDD.n1964 VDD.n1418 3.1005
R3603 VDD.n1966 VDD.n1965 3.1005
R3604 VDD.n1968 VDD.n1967 3.1005
R3605 VDD.n1417 VDD.n1411 3.1005
R3606 VDD.n1975 VDD.n1974 3.1005
R3607 VDD.n1976 VDD.n1410 3.1005
R3608 VDD.n1978 VDD.n1977 3.1005
R3609 VDD.n1402 VDD.n1401 3.1005
R3610 VDD.n984 VDD.n983 3.1005
R3611 VDD.n985 VDD.n969 3.1005
R3612 VDD.n987 VDD.n986 3.1005
R3613 VDD.n966 VDD.n965 3.1005
R3614 VDD.n996 VDD.n995 3.1005
R3615 VDD.n997 VDD.n964 3.1005
R3616 VDD.n999 VDD.n998 3.1005
R3617 VDD.n1007 VDD.n1006 3.1005
R3618 VDD.n1008 VDD.n957 3.1005
R3619 VDD.n1010 VDD.n1009 3.1005
R3620 VDD.n954 VDD.n953 3.1005
R3621 VDD.n1019 VDD.n1018 3.1005
R3622 VDD.n1020 VDD.n952 3.1005
R3623 VDD.n1022 VDD.n1021 3.1005
R3624 VDD.n949 VDD.n947 3.1005
R3625 VDD.n1032 VDD.n946 3.1005
R3626 VDD.n1034 VDD.n1033 3.1005
R3627 VDD.n943 VDD.n942 3.1005
R3628 VDD.n1044 VDD.n941 3.1005
R3629 VDD.n1045 VDD.n938 3.1005
R3630 VDD.n1057 VDD.n1056 3.1005
R3631 VDD.n1062 VDD.n1061 3.1005
R3632 VDD.n934 VDD.n933 3.1005
R3633 VDD.n1071 VDD.n1070 3.1005
R3634 VDD.n1072 VDD.n931 3.1005
R3635 VDD.n1074 VDD.n1073 3.1005
R3636 VDD.n927 VDD.n926 3.1005
R3637 VDD.n1082 VDD.n1081 3.1005
R3638 VDD.n1087 VDD.n1086 3.1005
R3639 VDD.n922 VDD.n921 3.1005
R3640 VDD.n1094 VDD.n1093 3.1005
R3641 VDD.n1095 VDD.n918 3.1005
R3642 VDD.n1097 VDD.n1096 3.1005
R3643 VDD.n915 VDD.n914 3.1005
R3644 VDD.n1105 VDD.n1104 3.1005
R3645 VDD.n1106 VDD.n913 3.1005
R3646 VDD.n910 VDD.n909 3.1005
R3647 VDD.n1118 VDD.n1117 3.1005
R3648 VDD.n1119 VDD.n908 3.1005
R3649 VDD.n905 VDD.n903 3.1005
R3650 VDD.n1132 VDD.n902 3.1005
R3651 VDD.n1134 VDD.n1133 3.1005
R3652 VDD.n1142 VDD.n1141 3.1005
R3653 VDD.n1143 VDD.n893 3.1005
R3654 VDD.n1145 VDD.n1144 3.1005
R3655 VDD.n890 VDD.n889 3.1005
R3656 VDD.n1154 VDD.n1153 3.1005
R3657 VDD.n1155 VDD.n888 3.1005
R3658 VDD.n1157 VDD.n1156 3.1005
R3659 VDD.n1165 VDD.n1164 3.1005
R3660 VDD.n1166 VDD.n881 3.1005
R3661 VDD.n1168 VDD.n1167 3.1005
R3662 VDD.n878 VDD.n877 3.1005
R3663 VDD.n1177 VDD.n1176 3.1005
R3664 VDD.n1178 VDD.n876 3.1005
R3665 VDD.n1180 VDD.n1179 3.1005
R3666 VDD.n873 VDD.n871 3.1005
R3667 VDD.n1190 VDD.n870 3.1005
R3668 VDD.n1192 VDD.n1191 3.1005
R3669 VDD.n867 VDD.n866 3.1005
R3670 VDD.n1202 VDD.n865 3.1005
R3671 VDD.n1203 VDD.n862 3.1005
R3672 VDD.n1215 VDD.n1214 3.1005
R3673 VDD.n1220 VDD.n1219 3.1005
R3674 VDD.n858 VDD.n857 3.1005
R3675 VDD.n1229 VDD.n1228 3.1005
R3676 VDD.n1230 VDD.n855 3.1005
R3677 VDD.n1232 VDD.n1231 3.1005
R3678 VDD.n850 VDD.n849 3.1005
R3679 VDD.n1244 VDD.n1243 3.1005
R3680 VDD.n1395 VDD.n1394 3.1005
R3681 VDD.n770 VDD.n765 3.1005
R3682 VDD.n306 VDD.n286 3.1005
R3683 VDD.n395 VDD.n375 3.1005
R3684 VDD.n484 VDD.n464 3.1005
R3685 VDD.n573 VDD.n553 3.1005
R3686 VDD.n764 VDD.n763 3.1005
R3687 VDD.n251 VDD.n242 3.1005
R3688 VDD.n238 VDD.n237 3.1005
R3689 VDD.n262 VDD.n261 3.1005
R3690 VDD.n263 VDD.n236 3.1005
R3691 VDD.n264 VDD.n233 3.1005
R3692 VDD.n274 VDD.n232 3.1005
R3693 VDD.n276 VDD.n275 3.1005
R3694 VDD.n278 VDD.n277 3.1005
R3695 VDD.n226 VDD.n225 3.1005
R3696 VDD.n284 VDD.n283 3.1005
R3697 VDD.n285 VDD.n224 3.1005
R3698 VDD.n300 VDD.n299 3.1005
R3699 VDD.n313 VDD.n219 3.1005
R3700 VDD.n315 VDD.n314 3.1005
R3701 VDD.n317 VDD.n316 3.1005
R3702 VDD.n214 VDD.n213 3.1005
R3703 VDD.n325 VDD.n324 3.1005
R3704 VDD.n331 VDD.n330 3.1005
R3705 VDD.n329 VDD.n209 3.1005
R3706 VDD.n340 VDD.n207 3.1005
R3707 VDD.n203 VDD.n202 3.1005
R3708 VDD.n351 VDD.n350 3.1005
R3709 VDD.n352 VDD.n201 3.1005
R3710 VDD.n353 VDD.n198 3.1005
R3711 VDD.n363 VDD.n197 3.1005
R3712 VDD.n365 VDD.n364 3.1005
R3713 VDD.n367 VDD.n366 3.1005
R3714 VDD.n191 VDD.n190 3.1005
R3715 VDD.n373 VDD.n372 3.1005
R3716 VDD.n374 VDD.n189 3.1005
R3717 VDD.n389 VDD.n388 3.1005
R3718 VDD.n402 VDD.n184 3.1005
R3719 VDD.n404 VDD.n403 3.1005
R3720 VDD.n406 VDD.n405 3.1005
R3721 VDD.n179 VDD.n178 3.1005
R3722 VDD.n414 VDD.n413 3.1005
R3723 VDD.n420 VDD.n419 3.1005
R3724 VDD.n418 VDD.n174 3.1005
R3725 VDD.n429 VDD.n172 3.1005
R3726 VDD.n168 VDD.n167 3.1005
R3727 VDD.n440 VDD.n439 3.1005
R3728 VDD.n441 VDD.n166 3.1005
R3729 VDD.n442 VDD.n163 3.1005
R3730 VDD.n452 VDD.n162 3.1005
R3731 VDD.n454 VDD.n453 3.1005
R3732 VDD.n456 VDD.n455 3.1005
R3733 VDD.n156 VDD.n155 3.1005
R3734 VDD.n462 VDD.n461 3.1005
R3735 VDD.n463 VDD.n154 3.1005
R3736 VDD.n478 VDD.n477 3.1005
R3737 VDD.n491 VDD.n149 3.1005
R3738 VDD.n493 VDD.n492 3.1005
R3739 VDD.n495 VDD.n494 3.1005
R3740 VDD.n144 VDD.n143 3.1005
R3741 VDD.n503 VDD.n502 3.1005
R3742 VDD.n509 VDD.n508 3.1005
R3743 VDD.n507 VDD.n139 3.1005
R3744 VDD.n518 VDD.n137 3.1005
R3745 VDD.n133 VDD.n132 3.1005
R3746 VDD.n529 VDD.n528 3.1005
R3747 VDD.n530 VDD.n131 3.1005
R3748 VDD.n531 VDD.n128 3.1005
R3749 VDD.n541 VDD.n127 3.1005
R3750 VDD.n543 VDD.n542 3.1005
R3751 VDD.n545 VDD.n544 3.1005
R3752 VDD.n121 VDD.n120 3.1005
R3753 VDD.n551 VDD.n550 3.1005
R3754 VDD.n552 VDD.n119 3.1005
R3755 VDD.n567 VDD.n566 3.1005
R3756 VDD.n580 VDD.n114 3.1005
R3757 VDD.n582 VDD.n581 3.1005
R3758 VDD.n585 VDD.n584 3.1005
R3759 VDD.n583 VDD.n109 3.1005
R3760 VDD.n592 VDD.n106 3.1005
R3761 VDD.n596 VDD.n104 3.1005
R3762 VDD.n598 VDD.n597 3.1005
R3763 VDD.n100 VDD.n99 3.1005
R3764 VDD.n608 VDD.n607 3.1005
R3765 VDD.n609 VDD.n96 3.1005
R3766 VDD.n611 VDD.n610 3.1005
R3767 VDD.n92 VDD.n91 3.1005
R3768 VDD.n622 VDD.n621 3.1005
R3769 VDD.n623 VDD.n90 3.1005
R3770 VDD.n625 VDD.n624 3.1005
R3771 VDD.n627 VDD.n83 3.1005
R3772 VDD.n637 VDD.n636 3.1005
R3773 VDD.n639 VDD.n638 3.1005
R3774 VDD.n741 VDD.n740 3.1005
R3775 VDD.n742 VDD.n23 3.1005
R3776 VDD.n745 VDD.n744 3.1005
R3777 VDD.n753 VDD.n18 3.1005
R3778 VDD.n755 VDD.n754 3.1005
R3779 VDD.n757 VDD.n756 3.1005
R3780 VDD.n2676 VDD.n2675 3.1005
R3781 VDD.n2533 VDD.n2532 3.1005
R3782 VDD.n2409 VDD.n2408 3.1005
R3783 VDD.n2285 VDD.n2284 3.1005
R3784 VDD.n2211 VDD.n2210 3.1005
R3785 VDD.n2109 VDD.n2107 3.1005
R3786 VDD.n2614 VDD.n2613 3.1005
R3787 VDD.n2618 VDD.n2617 3.1005
R3788 VDD.n2624 VDD.n2623 3.1005
R3789 VDD.n2628 VDD.n2627 3.1005
R3790 VDD.n2633 VDD.n2632 3.1005
R3791 VDD.n2637 VDD.n2636 3.1005
R3792 VDD.n2641 VDD.n2640 3.1005
R3793 VDD.n2651 VDD.n2650 3.1005
R3794 VDD.n2655 VDD.n2654 3.1005
R3795 VDD.n2658 VDD.n2657 3.1005
R3796 VDD.n2662 VDD.n2661 3.1005
R3797 VDD.n2666 VDD.n2665 3.1005
R3798 VDD.n2672 VDD.n2671 3.1005
R3799 VDD.n2701 VDD.n2700 3.1005
R3800 VDD.n2705 VDD.n2704 3.1005
R3801 VDD.n2709 VDD.n2708 3.1005
R3802 VDD.n2718 VDD.n2717 3.1005
R3803 VDD.n2719 VDD.n2602 3.1005
R3804 VDD.n2731 VDD.n2730 3.1005
R3805 VDD.n2595 VDD.n2594 3.1005
R3806 VDD.n2591 VDD.n2590 3.1005
R3807 VDD.n2587 VDD.n2586 3.1005
R3808 VDD.n2581 VDD.n2580 3.1005
R3809 VDD.n2577 VDD.n2576 3.1005
R3810 VDD.n2572 VDD.n2571 3.1005
R3811 VDD.n2568 VDD.n2567 3.1005
R3812 VDD.n2558 VDD.n2557 3.1005
R3813 VDD.n2554 VDD.n2553 3.1005
R3814 VDD.n2550 VDD.n2549 3.1005
R3815 VDD.n2547 VDD.n2546 3.1005
R3816 VDD.n2543 VDD.n2542 3.1005
R3817 VDD.n2539 VDD.n2538 3.1005
R3818 VDD.n2508 VDD.n2507 3.1005
R3819 VDD.n2504 VDD.n2503 3.1005
R3820 VDD.n2500 VDD.n2499 3.1005
R3821 VDD.n2491 VDD.n2490 3.1005
R3822 VDD.n2480 VDD.n0 3.1005
R3823 VDD.n2479 VDD.n2478 3.1005
R3824 VDD.n2471 VDD.n2470 3.1005
R3825 VDD.n2467 VDD.n2466 3.1005
R3826 VDD.n2463 VDD.n2462 3.1005
R3827 VDD.n2457 VDD.n2456 3.1005
R3828 VDD.n2453 VDD.n2452 3.1005
R3829 VDD.n2448 VDD.n2447 3.1005
R3830 VDD.n2444 VDD.n2443 3.1005
R3831 VDD.n2434 VDD.n2433 3.1005
R3832 VDD.n2430 VDD.n2429 3.1005
R3833 VDD.n2426 VDD.n2425 3.1005
R3834 VDD.n2423 VDD.n2422 3.1005
R3835 VDD.n2419 VDD.n2418 3.1005
R3836 VDD.n2415 VDD.n2414 3.1005
R3837 VDD.n2384 VDD.n2383 3.1005
R3838 VDD.n2380 VDD.n2379 3.1005
R3839 VDD.n2376 VDD.n2375 3.1005
R3840 VDD.n2367 VDD.n2366 3.1005
R3841 VDD.n2356 VDD.n4 3.1005
R3842 VDD.n2355 VDD.n2354 3.1005
R3843 VDD.n2347 VDD.n2346 3.1005
R3844 VDD.n2343 VDD.n2342 3.1005
R3845 VDD.n2339 VDD.n2338 3.1005
R3846 VDD.n2333 VDD.n2332 3.1005
R3847 VDD.n2329 VDD.n2328 3.1005
R3848 VDD.n2324 VDD.n2323 3.1005
R3849 VDD.n2320 VDD.n2319 3.1005
R3850 VDD.n2310 VDD.n2309 3.1005
R3851 VDD.n2306 VDD.n2305 3.1005
R3852 VDD.n2302 VDD.n2301 3.1005
R3853 VDD.n2299 VDD.n2298 3.1005
R3854 VDD.n2295 VDD.n2294 3.1005
R3855 VDD.n2291 VDD.n2290 3.1005
R3856 VDD.n2260 VDD.n2259 3.1005
R3857 VDD.n2256 VDD.n2255 3.1005
R3858 VDD.n2252 VDD.n2251 3.1005
R3859 VDD.n2243 VDD.n2242 3.1005
R3860 VDD.n2224 VDD.n8 3.1005
R3861 VDD.n2223 VDD.n2222 3.1005
R3862 VDD.n2215 VDD.n2214 3.1005
R3863 VDD.n2195 VDD.n2194 3.1005
R3864 VDD.n2190 VDD.n2189 3.1005
R3865 VDD.n2186 VDD.n2185 3.1005
R3866 VDD.n2176 VDD.n2175 3.1005
R3867 VDD.n2172 VDD.n2171 3.1005
R3868 VDD.n2168 VDD.n2167 3.1005
R3869 VDD.n2165 VDD.n2164 3.1005
R3870 VDD.n2161 VDD.n2160 3.1005
R3871 VDD.n2157 VDD.n2156 3.1005
R3872 VDD.n2151 VDD.n2150 3.1005
R3873 VDD.n2147 VDD.n2146 3.1005
R3874 VDD.n2137 VDD.n2136 3.1005
R3875 VDD.n2133 VDD.n2132 3.1005
R3876 VDD.n2129 VDD.n2128 3.1005
R3877 VDD.n2120 VDD.n2119 3.1005
R3878 VDD.n105 VDD.n100 3.09016
R3879 VDD.n626 VDD.n625 3.09016
R3880 VDD.n1662 VDD.n1578 3.05722
R3881 VDD.n1738 VDD.n1535 3.05722
R3882 VDD.n1815 VDD.n1497 3.05722
R3883 VDD.n1891 VDD.n1454 3.05722
R3884 VDD.n1968 VDD.n1416 3.05722
R3885 VDD.n995 VDD.n994 3.05722
R3886 VDD.n1074 VDD.n932 3.05722
R3887 VDD.n1153 VDD.n1152 3.05722
R3888 VDD.n1232 VDD.n856 3.05722
R3889 VDD.n580 VDD.n115 3.05722
R3890 VDD.n491 VDD.n150 3.05722
R3891 VDD.n402 VDD.n185 3.05722
R3892 VDD.n313 VDD.n220 3.05722
R3893 VDD.n2194 VDD.n2193 3.05722
R3894 VDD.n2328 VDD.n2327 3.05722
R3895 VDD.n2452 VDD.n2451 3.05722
R3896 VDD.n2576 VDD.n2575 3.05722
R3897 VDD.n2632 VDD.n2631 3.05722
R3898 VDD.n291 VDD 3.02729
R3899 VDD.n380 VDD 3.02729
R3900 VDD.n469 VDD 3.02729
R3901 VDD.n558 VDD 3.02729
R3902 VDD.n2681 VDD 3.02729
R3903 VDD.n2517 VDD 3.02729
R3904 VDD.n2393 VDD 3.02729
R3905 VDD.n2269 VDD 3.02729
R3906 VDD.n293 VDD.n292 2.92946
R3907 VDD.n382 VDD.n381 2.92946
R3908 VDD.n471 VDD.n470 2.92946
R3909 VDD.n560 VDD.n559 2.92946
R3910 VDD.n2685 VDD 2.89456
R3911 VDD.n2521 VDD 2.89456
R3912 VDD.n2397 VDD 2.89456
R3913 VDD.n2273 VDD 2.89456
R3914 VDD.n1248 VDD.n845 2.86947
R3915 VDD.n1381 VDD.n1380 2.7891
R3916 VDD.n572 VDD.n564 2.64878
R3917 VDD.n483 VDD.n475 2.64878
R3918 VDD.n394 VDD.n386 2.64878
R3919 VDD.n305 VDD.n297 2.64878
R3920 VDD.n1676 VDD 2.63939
R3921 VDD VDD.n1759 2.63939
R3922 VDD.n1829 VDD 2.63939
R3923 VDD VDD.n1912 2.63939
R3924 VDD.n2727 VDD 2.63208
R3925 VDD VDD.n2482 2.63208
R3926 VDD VDD.n2358 2.63208
R3927 VDD.n2239 VDD.n2238 2.63208
R3928 VDD VDD.n2226 2.63208
R3929 VDD VDD.n2111 2.63208
R3930 VDD.n1366 VDD.n1365 2.63101
R3931 VDD VDD.n334 2.60324
R3932 VDD VDD.n423 2.60324
R3933 VDD VDD.n512 2.60324
R3934 VDD.n1052 VDD 2.58202
R3935 VDD VDD.n1126 2.58202
R3936 VDD.n1210 VDD 2.58202
R3937 VDD.t348 VDD.n1254 2.58202
R3938 VDD.n1628 VDD.n1626 2.55931
R3939 VDD.n1649 VDD.n1648 2.55931
R3940 VDD.n1705 VDD.n1704 2.55931
R3941 VDD.n1728 VDD.n1727 2.55931
R3942 VDD.n1781 VDD.n1779 2.55931
R3943 VDD.n1802 VDD.n1801 2.55931
R3944 VDD.n1858 VDD.n1857 2.55931
R3945 VDD.n1881 VDD.n1880 2.55931
R3946 VDD.n1934 VDD.n1932 2.55931
R3947 VDD.n1955 VDD.n1954 2.55931
R3948 VDD.n960 VDD.n958 2.55931
R3949 VDD.n1031 VDD.n1030 2.55931
R3950 VDD.n1085 VDD.n1084 2.55931
R3951 VDD.n1109 VDD.n1107 2.55931
R3952 VDD.n884 VDD.n882 2.55931
R3953 VDD.n1189 VDD.n1188 2.55931
R3954 VDD.n267 VDD.n265 2.55931
R3955 VDD.n356 VDD.n354 2.55931
R3956 VDD.n445 VDD.n443 2.55931
R3957 VDD.n534 VDD.n532 2.55931
R3958 VDD.n2647 VDD.n2646 2.55931
R3959 VDD.n2564 VDD.n2563 2.55931
R3960 VDD.n2440 VDD.n2439 2.55931
R3961 VDD.n2316 VDD.n2315 2.55931
R3962 VDD.n2182 VDD.n2181 2.55931
R3963 VDD.n2143 VDD.n2142 2.55931
R3964 VDD.n294 VDD.n287 2.52171
R3965 VDD.n383 VDD.n376 2.52171
R3966 VDD.n472 VDD.n465 2.52171
R3967 VDD.n561 VDD.n554 2.52171
R3968 VDD.n2687 VDD.n2686 2.52171
R3969 VDD.n2523 VDD.n2522 2.52171
R3970 VDD.n2399 VDD.n2398 2.52171
R3971 VDD.n2275 VDD.n2274 2.52171
R3972 VDD.n1614 VDD.n1613 2.5203
R3973 VDD.n1694 VDD.n1693 2.5203
R3974 VDD.n1767 VDD.n1766 2.5203
R3975 VDD.n1847 VDD.n1846 2.5203
R3976 VDD.n1920 VDD.n1919 2.5203
R3977 VDD.n1043 VDD.n1042 2.5203
R3978 VDD.n1121 VDD.n1120 2.5203
R3979 VDD.n1201 VDD.n1200 2.5203
R3980 VDD.n253 VDD.n252 2.5203
R3981 VDD.n342 VDD.n341 2.5203
R3982 VDD.n431 VDD.n430 2.5203
R3983 VDD.n520 VDD.n519 2.5203
R3984 VDD.n2714 VDD.n2713 2.5203
R3985 VDD.n2496 VDD.n2495 2.5203
R3986 VDD.n2372 VDD.n2371 2.5203
R3987 VDD.n2248 VDD.n2247 2.5203
R3988 VDD.n2125 VDD.n2124 2.5203
R3989 VDD.n2059 VDD.n2058 2.51325
R3990 VDD.n2027 VDD.n2025 2.49102
R3991 VDD.n2093 VDD.n1993 2.49102
R3992 VDD.n1989 VDD.n1987 2.49102
R3993 VDD.n1611 VDD.n1610 2.49102
R3994 VDD.n1684 VDD.n1682 2.49102
R3995 VDD.n1764 VDD.n1763 2.49102
R3996 VDD.n1837 VDD.n1835 2.49102
R3997 VDD.n1917 VDD.n1916 2.49102
R3998 VDD.n1048 VDD.n1046 2.49102
R3999 VDD.n1131 VDD.n1130 2.49102
R4000 VDD.n1206 VDD.n1204 2.49102
R4001 VDD.n250 VDD.n249 2.49102
R4002 VDD.n339 VDD.n338 2.49102
R4003 VDD.n428 VDD.n427 2.49102
R4004 VDD.n517 VDD.n516 2.49102
R4005 VDD.n743 VDD.n25 2.49102
R4006 VDD.n14 VDD.n12 2.49102
R4007 VDD.n2722 VDD.n2720 2.49102
R4008 VDD.n2487 VDD.n2486 2.49102
R4009 VDD.n2363 VDD.n2362 2.49102
R4010 VDD.n2231 VDD.n2230 2.49102
R4011 VDD.n2116 VDD.n2115 2.49102
R4012 VDD.n1567 VDD.n1565 2.43201
R4013 VDD.n1753 VDD.n1752 2.43201
R4014 VDD.n1486 VDD.n1484 2.43201
R4015 VDD.n1906 VDD.n1905 2.43201
R4016 VDD.n1405 VDD.n1403 2.43201
R4017 VDD.n974 VDD.n972 2.43201
R4018 VDD.n1060 VDD.n1059 2.43201
R4019 VDD.n898 VDD.n896 2.43201
R4020 VDD.n1218 VDD.n1217 2.43201
R4021 VDD.n328 VDD.n327 2.43201
R4022 VDD.n417 VDD.n416 2.43201
R4023 VDD.n506 VDD.n505 2.43201
R4024 VDD.n595 VDD.n594 2.43201
R4025 VDD.n2610 VDD.n2609 2.43201
R4026 VDD.n2601 VDD.n2600 2.43201
R4027 VDD.n2477 VDD.n2476 2.43201
R4028 VDD.n2353 VDD.n2352 2.43201
R4029 VDD.n2221 VDD.n2220 2.43201
R4030 VDD.n1248 VDD.n1247 2.42487
R4031 VDD.n1328 VDD.n1327 2.42487
R4032 VDD.n1330 VDD.n1329 2.35689
R4033 VDD.n1236 VDD.n848 2.35689
R4034 VDD.n1360 VDD.n786 2.35366
R4035 VDD.n1383 VDD.n1382 2.35119
R4036 VDD.n1636 VDD.n1592 2.2074
R4037 VDD.n1553 VDD.n1548 2.2074
R4038 VDD.n1789 VDD.n1511 2.2074
R4039 VDD.n1472 VDD.n1467 2.2074
R4040 VDD.n1942 VDD.n1430 2.2074
R4041 VDD.n1017 VDD.n952 2.2074
R4042 VDD.n920 VDD.n915 2.2074
R4043 VDD.n1175 VDD.n876 2.2074
R4044 VDD.n1252 VDD.n1251 2.2074
R4045 VDD.n1263 VDD.n837 2.2074
R4046 VDD.n1271 VDD.n1270 2.2074
R4047 VDD.n1282 VDD.n827 2.2074
R4048 VDD.n1289 VDD.n1288 2.2074
R4049 VDD.n1311 VDD.n813 2.2074
R4050 VDD.n1319 VDD.n1318 2.2074
R4051 VDD.n1337 VDD.n1336 2.2074
R4052 VDD.n1348 VDD.n795 2.2074
R4053 VDD.n1356 VDD.n1355 2.2074
R4054 VDD.n1372 VDD.n1371 2.2074
R4055 VDD.n1390 VDD.n1389 2.2074
R4056 VDD.n639 VDD.n82 2.2074
R4057 VDD.n648 VDD.n647 2.2074
R4058 VDD.n653 VDD.n652 2.2074
R4059 VDD.n652 VDD.n70 2.2074
R4060 VDD.n665 VDD.n66 2.2074
R4061 VDD.n665 VDD.n68 2.2074
R4062 VDD.n673 VDD.n672 2.2074
R4063 VDD.n673 VDD.n60 2.2074
R4064 VDD.n685 VDD.n55 2.2074
R4065 VDD.n686 VDD.n685 2.2074
R4066 VDD.n691 VDD.n690 2.2074
R4067 VDD.n690 VDD.n48 2.2074
R4068 VDD.n703 VDD.n44 2.2074
R4069 VDD.n703 VDD.n46 2.2074
R4070 VDD.n711 VDD.n710 2.2074
R4071 VDD.n711 VDD.n38 2.2074
R4072 VDD.n723 VDD.n33 2.2074
R4073 VDD.n724 VDD.n723 2.2074
R4074 VDD.n732 VDD.n731 2.2074
R4075 VDD.n542 VDD.n126 2.2074
R4076 VDD.n453 VDD.n161 2.2074
R4077 VDD.n364 VDD.n196 2.2074
R4078 VDD.n275 VDD.n231 2.2074
R4079 VDD.n2156 VDD.n2153 2.2074
R4080 VDD.n2290 VDD.n2287 2.2074
R4081 VDD.n2279 VDD.n2266 2.2074
R4082 VDD.n2414 VDD.n2411 2.2074
R4083 VDD.n2403 VDD.n2390 2.2074
R4084 VDD.n2538 VDD.n2535 2.2074
R4085 VDD.n2527 VDD.n2514 2.2074
R4086 VDD.n2671 VDD.n2668 2.2074
R4087 VDD.n2691 VDD.n2678 2.2074
R4088 VDD.n572 VDD.n571 2.02155
R4089 VDD.n483 VDD.n482 2.02155
R4090 VDD.n394 VDD.n393 2.02155
R4091 VDD.n305 VDD.n304 2.02155
R4092 VDD.n2263 VDD.n2261 2.02155
R4093 VDD.n2387 VDD.n2385 2.02155
R4094 VDD.n2511 VDD.n2509 2.02155
R4095 VDD.n2696 VDD.n2694 2.02155
R4096 VDD.n1251 VDD.n841 1.98671
R4097 VDD.n1263 VDD.n839 1.98671
R4098 VDD.n1271 VDD.n831 1.98671
R4099 VDD.n1283 VDD.n1282 1.98671
R4100 VDD.n1288 VDD.n825 1.98671
R4101 VDD.n1300 VDD.n817 1.98671
R4102 VDD.n1312 VDD.n1311 1.98671
R4103 VDD.n1318 VDD.n811 1.98671
R4104 VDD.n1337 VDD.n799 1.98671
R4105 VDD.n1349 VDD.n1348 1.98671
R4106 VDD.n1355 VDD.n793 1.98671
R4107 VDD.n1371 VDD.n783 1.98671
R4108 VDD.n1391 VDD.n1390 1.98671
R4109 VDD VDD.n290 1.91393
R4110 VDD VDD.n379 1.91393
R4111 VDD VDD.n468 1.91393
R4112 VDD VDD.n557 1.91393
R4113 VDD VDD.n2680 1.85046
R4114 VDD VDD.n2516 1.85046
R4115 VDD VDD.n2392 1.85046
R4116 VDD VDD.n2268 1.85046
R4117 VDD.n1259 VDD.n841 1.76602
R4118 VDD.n839 VDD.n838 1.76602
R4119 VDD.n1275 VDD.n831 1.76602
R4120 VDD.n1284 VDD.n1283 1.76602
R4121 VDD.n825 VDD.n819 1.76602
R4122 VDD.n1299 VDD.n819 1.76602
R4123 VDD.n1304 VDD.n817 1.76602
R4124 VDD.n1313 VDD.n1312 1.76602
R4125 VDD.n811 VDD.n805 1.76602
R4126 VDD.n1341 VDD.n799 1.76602
R4127 VDD.n1350 VDD.n1349 1.76602
R4128 VDD.n793 VDD.n785 1.76602
R4129 VDD.n783 VDD.n776 1.76602
R4130 VDD.n1391 VDD.n769 1.76602
R4131 VDD.n647 VDD.n78 1.76602
R4132 VDD.n1568 VDD.n1567 1.72554
R4133 VDD.n1752 VDD.n1527 1.72554
R4134 VDD.n1487 VDD.n1486 1.72554
R4135 VDD.n1905 VDD.n1446 1.72554
R4136 VDD.n1406 VDD.n1405 1.72554
R4137 VDD.n975 VDD.n974 1.72554
R4138 VDD.n1059 VDD.n937 1.72554
R4139 VDD.n899 VDD.n898 1.72554
R4140 VDD.n1217 VDD.n861 1.72554
R4141 VDD.n327 VDD.n212 1.72554
R4142 VDD.n416 VDD.n177 1.72554
R4143 VDD.n505 VDD.n142 1.72554
R4144 VDD.n594 VDD.n593 1.72554
R4145 VDD.n2609 VDD.n2608 1.72554
R4146 VDD.n2600 VDD.n2599 1.72554
R4147 VDD.n2476 VDD.n2475 1.72554
R4148 VDD.n2352 VDD.n2351 1.72554
R4149 VDD.n2220 VDD.n2219 1.72554
R4150 VDD.n2028 VDD.n2027 1.57241
R4151 VDD.n2094 VDD.n2093 1.57241
R4152 VDD.n1990 VDD.n1989 1.57241
R4153 VDD.n1610 VDD.n1609 1.57241
R4154 VDD.n1685 VDD.n1684 1.57241
R4155 VDD.n1763 VDD.n1762 1.57241
R4156 VDD.n1838 VDD.n1837 1.57241
R4157 VDD.n1916 VDD.n1915 1.57241
R4158 VDD.n1049 VDD.n1048 1.57241
R4159 VDD.n1130 VDD.n1129 1.57241
R4160 VDD.n1207 VDD.n1206 1.57241
R4161 VDD.n249 VDD.n248 1.57241
R4162 VDD.n338 VDD.n337 1.57241
R4163 VDD.n427 VDD.n426 1.57241
R4164 VDD.n516 VDD.n515 1.57241
R4165 VDD.n746 VDD.n25 1.57241
R4166 VDD.n15 VDD.n14 1.57241
R4167 VDD.n2723 VDD.n2722 1.57241
R4168 VDD.n2486 VDD.n2485 1.57241
R4169 VDD.n2362 VDD.n2361 1.57241
R4170 VDD.n2230 VDD.n2229 1.57241
R4171 VDD.n2115 VDD.n2114 1.57241
R4172 VDD.n1252 VDD.n845 1.54533
R4173 VDD.n1258 VDD.n837 1.54533
R4174 VDD.n1270 VDD.n833 1.54533
R4175 VDD.n1276 VDD.n827 1.54533
R4176 VDD.n1289 VDD.n824 1.54533
R4177 VDD.n1305 VDD.n813 1.54533
R4178 VDD.n1319 VDD.n810 1.54533
R4179 VDD.n1336 VDD.n801 1.54533
R4180 VDD.n1342 VDD.n795 1.54533
R4181 VDD.n1356 VDD.n792 1.54533
R4182 VDD.n1372 VDD.n782 1.54533
R4183 VDD.n1389 VDD.n772 1.54533
R4184 VDD.n641 VDD.n640 1.54533
R4185 VDD.n649 VDD.n648 1.54533
R4186 VDD.n653 VDD.n75 1.54533
R4187 VDD.n661 VDD.n70 1.54533
R4188 VDD.n660 VDD.n659 1.54533
R4189 VDD.n659 VDD.n66 1.54533
R4190 VDD.n68 VDD.n67 1.54533
R4191 VDD.n672 VDD.n62 1.54533
R4192 VDD.n677 VDD.n60 1.54533
R4193 VDD.n679 VDD.n55 1.54533
R4194 VDD.n687 VDD.n686 1.54533
R4195 VDD.n691 VDD.n53 1.54533
R4196 VDD.n699 VDD.n48 1.54533
R4197 VDD.n697 VDD.n44 1.54533
R4198 VDD.n46 VDD.n45 1.54533
R4199 VDD.n710 VDD.n40 1.54533
R4200 VDD.n715 VDD.n38 1.54533
R4201 VDD.n717 VDD.n33 1.54533
R4202 VDD.n725 VDD.n724 1.54533
R4203 VDD.n732 VDD.n30 1.54533
R4204 VDD.n728 VDD.n26 1.54533
R4205 VDD.n2279 VDD.n2278 1.54533
R4206 VDD.n2403 VDD.n2402 1.54533
R4207 VDD.n2527 VDD.n2526 1.54533
R4208 VDD.n2691 VDD.n2690 1.54533
R4209 VDD.n2058 VDD.n2057 1.5148
R4210 VDD.n1615 VDD.n1614 1.49652
R4211 VDD.n1693 VDD.n1692 1.49652
R4212 VDD.n1768 VDD.n1767 1.49652
R4213 VDD.n1846 VDD.n1845 1.49652
R4214 VDD.n1921 VDD.n1920 1.49652
R4215 VDD.n1042 VDD.n1041 1.49652
R4216 VDD.n1122 VDD.n1121 1.49652
R4217 VDD.n1200 VDD.n1199 1.49652
R4218 VDD.n254 VDD.n253 1.49652
R4219 VDD.n343 VDD.n342 1.49652
R4220 VDD.n432 VDD.n431 1.49652
R4221 VDD.n521 VDD.n520 1.49652
R4222 VDD.n2713 VDD.n2712 1.49652
R4223 VDD.n2495 VDD.n2494 1.49652
R4224 VDD.n2371 VDD.n2370 1.49652
R4225 VDD.n2247 VDD.n2246 1.49652
R4226 VDD.n2124 VDD.n2123 1.49652
R4227 VDD.n2201 VDD.n2199 1.43334
R4228 VDD.n1629 VDD.n1628 1.39551
R4229 VDD.n1648 VDD.n1581 1.39551
R4230 VDD.n1704 VDD.n1703 1.39551
R4231 VDD.n1727 VDD.n1538 1.39551
R4232 VDD.n1782 VDD.n1781 1.39551
R4233 VDD.n1801 VDD.n1500 1.39551
R4234 VDD.n1857 VDD.n1856 1.39551
R4235 VDD.n1880 VDD.n1457 1.39551
R4236 VDD.n1935 VDD.n1934 1.39551
R4237 VDD.n1954 VDD.n1419 1.39551
R4238 VDD.n961 VDD.n960 1.39551
R4239 VDD.n1030 VDD.n1029 1.39551
R4240 VDD.n1084 VDD.n925 1.39551
R4241 VDD.n1110 VDD.n1109 1.39551
R4242 VDD.n885 VDD.n884 1.39551
R4243 VDD.n1188 VDD.n1187 1.39551
R4244 VDD.n268 VDD.n267 1.39551
R4245 VDD.n357 VDD.n356 1.39551
R4246 VDD.n446 VDD.n445 1.39551
R4247 VDD.n535 VDD.n534 1.39551
R4248 VDD.n2646 VDD.n2645 1.39551
R4249 VDD.n2563 VDD.n2562 1.39551
R4250 VDD.n2439 VDD.n2438 1.39551
R4251 VDD.n2315 VDD.n2314 1.39551
R4252 VDD.n2181 VDD.n2180 1.39551
R4253 VDD.n2142 VDD.n2141 1.39551
R4254 VDD.n728 VDD.n31 1.32464
R4255 VDD.n2008 VDD.n2001 1.10395
R4256 VDD.n753 VDD.n20 1.10395
R4257 VDD.n731 VDD.n31 0.883259
R4258 VDD.n2084 VDD 0.862479
R4259 VDD.n293 VDD.n287 0.776258
R4260 VDD.n382 VDD.n376 0.776258
R4261 VDD.n471 VDD.n465 0.776258
R4262 VDD.n560 VDD.n554 0.776258
R4263 VDD.n290 VDD.n289 0.750619
R4264 VDD.n379 VDD.n378 0.750619
R4265 VDD.n468 VDD.n467 0.750619
R4266 VDD.n557 VDD.n556 0.750619
R4267 VDD.n2004 VDD.n2003 0.662569
R4268 VDD.n1248 VDD.n847 0.662569
R4269 VDD.n716 VDD.n715 0.662569
R4270 VDD.n1668 VDD.n1575 0.478112
R4271 VDD.n1742 VDD.n1533 0.478112
R4272 VDD.n1821 VDD.n1494 0.478112
R4273 VDD.n1895 VDD.n1452 0.478112
R4274 VDD.n1974 VDD.n1413 0.478112
R4275 VDD.n987 VDD.n971 0.478112
R4276 VDD.n1070 VDD.n1069 0.478112
R4277 VDD.n1145 VDD.n895 0.478112
R4278 VDD.n1228 VDD.n1227 0.478112
R4279 VDD.n585 VDD.n113 0.478112
R4280 VDD.n495 VDD.n148 0.478112
R4281 VDD.n406 VDD.n183 0.478112
R4282 VDD.n317 VDD.n218 0.478112
R4283 VDD.n2206 VDD.n2205 0.478112
R4284 VDD.n2338 VDD.n2337 0.478112
R4285 VDD.n2462 VDD.n2461 0.478112
R4286 VDD.n2586 VDD.n2585 0.478112
R4287 VDD.n2623 VDD.n2622 0.478112
R4288 VDD.n636 VDD.n85 0.441879
R4289 VDD.n640 VDD.n78 0.441879
R4290 VDD.n632 VDD.n87 0.426767
R4291 VDD.n87 VDD.n82 0.426767
R4292 VDD.n2686 VDD.n2685 0.373349
R4293 VDD.n2522 VDD.n2521 0.373349
R4294 VDD.n2398 VDD.n2397 0.373349
R4295 VDD.n2274 VDD.n2273 0.373349
R4296 VDD.n2278 VDD.n2277 0.332764
R4297 VDD.n2402 VDD.n2401 0.332063
R4298 VDD.n2526 VDD.n2525 0.332063
R4299 VDD.n2690 VDD.n2689 0.331371
R4300 VDD.n1985 VDD 0.28318
R4301 VDD.n291 VDD 0.259429
R4302 VDD.n380 VDD 0.259429
R4303 VDD.n469 VDD 0.259429
R4304 VDD.n558 VDD 0.259429
R4305 VDD.n2681 VDD 0.259429
R4306 VDD.n2517 VDD 0.259429
R4307 VDD.n2393 VDD 0.259429
R4308 VDD.n2269 VDD 0.259429
R4309 VDD.n2199 VDD.n2198 0.225571
R4310 VDD.n1300 VDD.n1299 0.22119
R4311 VDD.n740 VDD.n739 0.22119
R4312 VDD.n2242 VDD.n2234 0.22119
R4313 VDD.n2201 VDD.n2200 0.191545
R4314 VDD.n1986 VDD 0.151171
R4315 VDD.n2037 VDD.n2025 0.120292
R4316 VDD.n2038 VDD.n2037 0.120292
R4317 VDD.n2039 VDD.n2038 0.120292
R4318 VDD.n2039 VDD.n2018 0.120292
R4319 VDD.n2048 VDD.n2018 0.120292
R4320 VDD.n2049 VDD.n2048 0.120292
R4321 VDD.n2050 VDD.n2049 0.120292
R4322 VDD.n2050 VDD.n2013 0.120292
R4323 VDD.n2059 VDD.n2013 0.120292
R4324 VDD.n2060 VDD.n2059 0.120292
R4325 VDD.n2061 VDD.n2060 0.120292
R4326 VDD.n2061 VDD.n2005 0.120292
R4327 VDD.n2070 VDD.n2005 0.120292
R4328 VDD.n2071 VDD.n2070 0.120292
R4329 VDD.n2073 VDD.n2071 0.120292
R4330 VDD.n2073 VDD.n2072 0.120292
R4331 VDD.n2072 VDD.n1997 0.120292
R4332 VDD.n2082 VDD.n1997 0.120292
R4333 VDD.n2084 VDD.n2083 0.120292
R4334 VDD.n2083 VDD.n1993 0.120292
R4335 VDD.n2096 VDD.n1993 0.120292
R4336 VDD.n2097 VDD.n1987 0.120292
R4337 VDD.n2105 VDD.n1987 0.120292
R4338 VDD.n1612 VDD.n1611 0.120292
R4339 VDD.n1613 VDD.n1612 0.120292
R4340 VDD.n1613 VDD.n1598 0.120292
R4341 VDD.n1623 VDD.n1598 0.120292
R4342 VDD.n1624 VDD.n1623 0.120292
R4343 VDD.n1626 VDD.n1624 0.120292
R4344 VDD.n1626 VDD.n1625 0.120292
R4345 VDD.n1625 VDD.n1593 0.120292
R4346 VDD.n1637 VDD.n1593 0.120292
R4347 VDD.n1638 VDD.n1637 0.120292
R4348 VDD.n1638 VDD.n1586 0.120292
R4349 VDD.n1645 VDD.n1586 0.120292
R4350 VDD.n1646 VDD.n1645 0.120292
R4351 VDD.n1650 VDD.n1646 0.120292
R4352 VDD.n1650 VDD.n1649 0.120292
R4353 VDD.n1649 VDD.n1580 0.120292
R4354 VDD.n1660 VDD.n1580 0.120292
R4355 VDD.n1661 VDD.n1660 0.120292
R4356 VDD.n1661 VDD.n1573 0.120292
R4357 VDD.n1669 VDD.n1573 0.120292
R4358 VDD.n1670 VDD.n1669 0.120292
R4359 VDD.n1671 VDD.n1670 0.120292
R4360 VDD.n1671 VDD.n1565 0.120292
R4361 VDD.n1680 VDD.n1565 0.120292
R4362 VDD.n1682 VDD.n1560 0.120292
R4363 VDD.n1694 VDD.n1560 0.120292
R4364 VDD.n1695 VDD.n1694 0.120292
R4365 VDD.n1696 VDD.n1695 0.120292
R4366 VDD.n1696 VDD.n1554 0.120292
R4367 VDD.n1705 VDD.n1554 0.120292
R4368 VDD.n1706 VDD.n1705 0.120292
R4369 VDD.n1707 VDD.n1706 0.120292
R4370 VDD.n1707 VDD.n1546 0.120292
R4371 VDD.n1715 VDD.n1546 0.120292
R4372 VDD.n1716 VDD.n1715 0.120292
R4373 VDD.n1717 VDD.n1716 0.120292
R4374 VDD.n1717 VDD.n1540 0.120292
R4375 VDD.n1725 VDD.n1540 0.120292
R4376 VDD.n1728 VDD.n1725 0.120292
R4377 VDD.n1730 VDD.n1728 0.120292
R4378 VDD.n1730 VDD.n1729 0.120292
R4379 VDD.n1729 VDD.n1534 0.120292
R4380 VDD.n1740 VDD.n1534 0.120292
R4381 VDD.n1741 VDD.n1740 0.120292
R4382 VDD.n1741 VDD.n1528 0.120292
R4383 VDD.n1750 VDD.n1528 0.120292
R4384 VDD.n1753 VDD.n1750 0.120292
R4385 VDD.n1755 VDD.n1753 0.120292
R4386 VDD.n1765 VDD.n1764 0.120292
R4387 VDD.n1766 VDD.n1765 0.120292
R4388 VDD.n1766 VDD.n1517 0.120292
R4389 VDD.n1776 VDD.n1517 0.120292
R4390 VDD.n1777 VDD.n1776 0.120292
R4391 VDD.n1779 VDD.n1777 0.120292
R4392 VDD.n1779 VDD.n1778 0.120292
R4393 VDD.n1778 VDD.n1512 0.120292
R4394 VDD.n1790 VDD.n1512 0.120292
R4395 VDD.n1791 VDD.n1790 0.120292
R4396 VDD.n1791 VDD.n1505 0.120292
R4397 VDD.n1798 VDD.n1505 0.120292
R4398 VDD.n1799 VDD.n1798 0.120292
R4399 VDD.n1803 VDD.n1799 0.120292
R4400 VDD.n1803 VDD.n1802 0.120292
R4401 VDD.n1802 VDD.n1499 0.120292
R4402 VDD.n1813 VDD.n1499 0.120292
R4403 VDD.n1814 VDD.n1813 0.120292
R4404 VDD.n1814 VDD.n1492 0.120292
R4405 VDD.n1822 VDD.n1492 0.120292
R4406 VDD.n1823 VDD.n1822 0.120292
R4407 VDD.n1824 VDD.n1823 0.120292
R4408 VDD.n1824 VDD.n1484 0.120292
R4409 VDD.n1833 VDD.n1484 0.120292
R4410 VDD.n1835 VDD.n1479 0.120292
R4411 VDD.n1847 VDD.n1479 0.120292
R4412 VDD.n1848 VDD.n1847 0.120292
R4413 VDD.n1849 VDD.n1848 0.120292
R4414 VDD.n1849 VDD.n1473 0.120292
R4415 VDD.n1858 VDD.n1473 0.120292
R4416 VDD.n1859 VDD.n1858 0.120292
R4417 VDD.n1860 VDD.n1859 0.120292
R4418 VDD.n1860 VDD.n1465 0.120292
R4419 VDD.n1868 VDD.n1465 0.120292
R4420 VDD.n1869 VDD.n1868 0.120292
R4421 VDD.n1870 VDD.n1869 0.120292
R4422 VDD.n1870 VDD.n1459 0.120292
R4423 VDD.n1878 VDD.n1459 0.120292
R4424 VDD.n1881 VDD.n1878 0.120292
R4425 VDD.n1883 VDD.n1881 0.120292
R4426 VDD.n1883 VDD.n1882 0.120292
R4427 VDD.n1882 VDD.n1453 0.120292
R4428 VDD.n1893 VDD.n1453 0.120292
R4429 VDD.n1894 VDD.n1893 0.120292
R4430 VDD.n1894 VDD.n1447 0.120292
R4431 VDD.n1903 VDD.n1447 0.120292
R4432 VDD.n1906 VDD.n1903 0.120292
R4433 VDD.n1908 VDD.n1906 0.120292
R4434 VDD.n1918 VDD.n1917 0.120292
R4435 VDD.n1919 VDD.n1918 0.120292
R4436 VDD.n1919 VDD.n1436 0.120292
R4437 VDD.n1929 VDD.n1436 0.120292
R4438 VDD.n1930 VDD.n1929 0.120292
R4439 VDD.n1932 VDD.n1930 0.120292
R4440 VDD.n1932 VDD.n1931 0.120292
R4441 VDD.n1931 VDD.n1431 0.120292
R4442 VDD.n1943 VDD.n1431 0.120292
R4443 VDD.n1944 VDD.n1943 0.120292
R4444 VDD.n1944 VDD.n1424 0.120292
R4445 VDD.n1951 VDD.n1424 0.120292
R4446 VDD.n1952 VDD.n1951 0.120292
R4447 VDD.n1956 VDD.n1952 0.120292
R4448 VDD.n1956 VDD.n1955 0.120292
R4449 VDD.n1955 VDD.n1418 0.120292
R4450 VDD.n1966 VDD.n1418 0.120292
R4451 VDD.n1967 VDD.n1966 0.120292
R4452 VDD.n1967 VDD.n1411 0.120292
R4453 VDD.n1975 VDD.n1411 0.120292
R4454 VDD.n1976 VDD.n1975 0.120292
R4455 VDD.n1977 VDD.n1976 0.120292
R4456 VDD.n1977 VDD.n1403 0.120292
R4457 VDD.n1984 VDD.n1403 0.120292
R4458 VDD.n984 VDD.n972 0.120292
R4459 VDD.n985 VDD.n984 0.120292
R4460 VDD.n986 VDD.n985 0.120292
R4461 VDD.n986 VDD.n965 0.120292
R4462 VDD.n996 VDD.n965 0.120292
R4463 VDD.n997 VDD.n996 0.120292
R4464 VDD.n998 VDD.n997 0.120292
R4465 VDD.n998 VDD.n958 0.120292
R4466 VDD.n1007 VDD.n958 0.120292
R4467 VDD.n1008 VDD.n1007 0.120292
R4468 VDD.n1009 VDD.n1008 0.120292
R4469 VDD.n1009 VDD.n953 0.120292
R4470 VDD.n1019 VDD.n953 0.120292
R4471 VDD.n1020 VDD.n1019 0.120292
R4472 VDD.n1021 VDD.n1020 0.120292
R4473 VDD.n1021 VDD.n947 0.120292
R4474 VDD.n1031 VDD.n947 0.120292
R4475 VDD.n1032 VDD.n1031 0.120292
R4476 VDD.n1033 VDD.n1032 0.120292
R4477 VDD.n1033 VDD.n942 0.120292
R4478 VDD.n1043 VDD.n942 0.120292
R4479 VDD.n1044 VDD.n1043 0.120292
R4480 VDD.n1046 VDD.n1044 0.120292
R4481 VDD.n1046 VDD.n1045 0.120292
R4482 VDD.n1060 VDD.n1057 0.120292
R4483 VDD.n1061 VDD.n1060 0.120292
R4484 VDD.n1061 VDD.n933 0.120292
R4485 VDD.n1071 VDD.n933 0.120292
R4486 VDD.n1072 VDD.n1071 0.120292
R4487 VDD.n1073 VDD.n1072 0.120292
R4488 VDD.n1073 VDD.n926 0.120292
R4489 VDD.n1082 VDD.n926 0.120292
R4490 VDD.n1085 VDD.n1082 0.120292
R4491 VDD.n1086 VDD.n1085 0.120292
R4492 VDD.n1086 VDD.n921 0.120292
R4493 VDD.n1094 VDD.n921 0.120292
R4494 VDD.n1095 VDD.n1094 0.120292
R4495 VDD.n1096 VDD.n1095 0.120292
R4496 VDD.n1096 VDD.n914 0.120292
R4497 VDD.n1105 VDD.n914 0.120292
R4498 VDD.n1106 VDD.n1105 0.120292
R4499 VDD.n1107 VDD.n1106 0.120292
R4500 VDD.n1107 VDD.n909 0.120292
R4501 VDD.n1118 VDD.n909 0.120292
R4502 VDD.n1119 VDD.n1118 0.120292
R4503 VDD.n1120 VDD.n1119 0.120292
R4504 VDD.n1120 VDD.n903 0.120292
R4505 VDD.n1131 VDD.n903 0.120292
R4506 VDD.n1132 VDD.n1131 0.120292
R4507 VDD.n1133 VDD.n896 0.120292
R4508 VDD.n1142 VDD.n896 0.120292
R4509 VDD.n1143 VDD.n1142 0.120292
R4510 VDD.n1144 VDD.n1143 0.120292
R4511 VDD.n1144 VDD.n889 0.120292
R4512 VDD.n1154 VDD.n889 0.120292
R4513 VDD.n1155 VDD.n1154 0.120292
R4514 VDD.n1156 VDD.n1155 0.120292
R4515 VDD.n1156 VDD.n882 0.120292
R4516 VDD.n1165 VDD.n882 0.120292
R4517 VDD.n1166 VDD.n1165 0.120292
R4518 VDD.n1167 VDD.n1166 0.120292
R4519 VDD.n1167 VDD.n877 0.120292
R4520 VDD.n1177 VDD.n877 0.120292
R4521 VDD.n1178 VDD.n1177 0.120292
R4522 VDD.n1179 VDD.n1178 0.120292
R4523 VDD.n1179 VDD.n871 0.120292
R4524 VDD.n1189 VDD.n871 0.120292
R4525 VDD.n1190 VDD.n1189 0.120292
R4526 VDD.n1191 VDD.n1190 0.120292
R4527 VDD.n1191 VDD.n866 0.120292
R4528 VDD.n1201 VDD.n866 0.120292
R4529 VDD.n1202 VDD.n1201 0.120292
R4530 VDD.n1204 VDD.n1202 0.120292
R4531 VDD.n1204 VDD.n1203 0.120292
R4532 VDD.n1218 VDD.n1215 0.120292
R4533 VDD.n1219 VDD.n1218 0.120292
R4534 VDD.n1219 VDD.n857 0.120292
R4535 VDD.n1229 VDD.n857 0.120292
R4536 VDD.n1230 VDD.n1229 0.120292
R4537 VDD.n1231 VDD.n1230 0.120292
R4538 VDD.n1231 VDD.n849 0.120292
R4539 VDD.n1244 VDD.n849 0.120292
R4540 VDD.n1394 VDD.n765 0.120292
R4541 VDD.n1402 VDD.n765 0.120292
R4542 VDD.n251 VDD.n250 0.120292
R4543 VDD.n252 VDD.n251 0.120292
R4544 VDD.n252 VDD.n237 0.120292
R4545 VDD.n262 VDD.n237 0.120292
R4546 VDD.n263 VDD.n262 0.120292
R4547 VDD.n265 VDD.n263 0.120292
R4548 VDD.n265 VDD.n264 0.120292
R4549 VDD.n264 VDD.n232 0.120292
R4550 VDD.n276 VDD.n232 0.120292
R4551 VDD.n277 VDD.n276 0.120292
R4552 VDD.n277 VDD.n225 0.120292
R4553 VDD.n284 VDD.n225 0.120292
R4554 VDD.n285 VDD.n284 0.120292
R4555 VDD.n286 VDD.n285 0.120292
R4556 VDD.n303 VDD.n286 0.120292
R4557 VDD.n303 VDD.n302 0.120292
R4558 VDD.n302 VDD.n299 0.120292
R4559 VDD.n299 VDD.n219 0.120292
R4560 VDD.n315 VDD.n219 0.120292
R4561 VDD.n316 VDD.n315 0.120292
R4562 VDD.n316 VDD.n213 0.120292
R4563 VDD.n325 VDD.n213 0.120292
R4564 VDD.n328 VDD.n325 0.120292
R4565 VDD.n330 VDD.n328 0.120292
R4566 VDD.n340 VDD.n339 0.120292
R4567 VDD.n341 VDD.n340 0.120292
R4568 VDD.n341 VDD.n202 0.120292
R4569 VDD.n351 VDD.n202 0.120292
R4570 VDD.n352 VDD.n351 0.120292
R4571 VDD.n354 VDD.n352 0.120292
R4572 VDD.n354 VDD.n353 0.120292
R4573 VDD.n353 VDD.n197 0.120292
R4574 VDD.n365 VDD.n197 0.120292
R4575 VDD.n366 VDD.n365 0.120292
R4576 VDD.n366 VDD.n190 0.120292
R4577 VDD.n373 VDD.n190 0.120292
R4578 VDD.n374 VDD.n373 0.120292
R4579 VDD.n375 VDD.n374 0.120292
R4580 VDD.n392 VDD.n375 0.120292
R4581 VDD.n392 VDD.n391 0.120292
R4582 VDD.n391 VDD.n388 0.120292
R4583 VDD.n388 VDD.n184 0.120292
R4584 VDD.n404 VDD.n184 0.120292
R4585 VDD.n405 VDD.n404 0.120292
R4586 VDD.n405 VDD.n178 0.120292
R4587 VDD.n414 VDD.n178 0.120292
R4588 VDD.n417 VDD.n414 0.120292
R4589 VDD.n419 VDD.n417 0.120292
R4590 VDD.n429 VDD.n428 0.120292
R4591 VDD.n430 VDD.n429 0.120292
R4592 VDD.n430 VDD.n167 0.120292
R4593 VDD.n440 VDD.n167 0.120292
R4594 VDD.n441 VDD.n440 0.120292
R4595 VDD.n443 VDD.n441 0.120292
R4596 VDD.n443 VDD.n442 0.120292
R4597 VDD.n442 VDD.n162 0.120292
R4598 VDD.n454 VDD.n162 0.120292
R4599 VDD.n455 VDD.n454 0.120292
R4600 VDD.n455 VDD.n155 0.120292
R4601 VDD.n462 VDD.n155 0.120292
R4602 VDD.n463 VDD.n462 0.120292
R4603 VDD.n464 VDD.n463 0.120292
R4604 VDD.n481 VDD.n464 0.120292
R4605 VDD.n481 VDD.n480 0.120292
R4606 VDD.n480 VDD.n477 0.120292
R4607 VDD.n477 VDD.n149 0.120292
R4608 VDD.n493 VDD.n149 0.120292
R4609 VDD.n494 VDD.n493 0.120292
R4610 VDD.n494 VDD.n143 0.120292
R4611 VDD.n503 VDD.n143 0.120292
R4612 VDD.n506 VDD.n503 0.120292
R4613 VDD.n508 VDD.n506 0.120292
R4614 VDD.n518 VDD.n517 0.120292
R4615 VDD.n519 VDD.n518 0.120292
R4616 VDD.n519 VDD.n132 0.120292
R4617 VDD.n529 VDD.n132 0.120292
R4618 VDD.n530 VDD.n529 0.120292
R4619 VDD.n532 VDD.n530 0.120292
R4620 VDD.n532 VDD.n531 0.120292
R4621 VDD.n531 VDD.n127 0.120292
R4622 VDD.n543 VDD.n127 0.120292
R4623 VDD.n544 VDD.n543 0.120292
R4624 VDD.n544 VDD.n120 0.120292
R4625 VDD.n551 VDD.n120 0.120292
R4626 VDD.n552 VDD.n551 0.120292
R4627 VDD.n553 VDD.n552 0.120292
R4628 VDD.n570 VDD.n553 0.120292
R4629 VDD.n570 VDD.n569 0.120292
R4630 VDD.n569 VDD.n566 0.120292
R4631 VDD.n566 VDD.n114 0.120292
R4632 VDD.n582 VDD.n114 0.120292
R4633 VDD.n584 VDD.n582 0.120292
R4634 VDD.n584 VDD.n583 0.120292
R4635 VDD.n583 VDD.n106 0.120292
R4636 VDD.n595 VDD.n106 0.120292
R4637 VDD.n596 VDD.n595 0.120292
R4638 VDD.n597 VDD.n99 0.120292
R4639 VDD.n608 VDD.n99 0.120292
R4640 VDD.n609 VDD.n608 0.120292
R4641 VDD.n610 VDD.n609 0.120292
R4642 VDD.n610 VDD.n91 0.120292
R4643 VDD.n622 VDD.n91 0.120292
R4644 VDD.n623 VDD.n622 0.120292
R4645 VDD.n624 VDD.n623 0.120292
R4646 VDD.n624 VDD.n83 0.120292
R4647 VDD.n637 VDD.n83 0.120292
R4648 VDD.n638 VDD.n637 0.120292
R4649 VDD.n742 VDD.n741 0.120292
R4650 VDD.n743 VDD.n742 0.120292
R4651 VDD.n744 VDD.n743 0.120292
R4652 VDD.n744 VDD.n18 0.120292
R4653 VDD.n755 VDD.n18 0.120292
R4654 VDD.n756 VDD.n12 0.120292
R4655 VDD.n764 VDD.n12 0.120292
R4656 VDD.n2614 VDD.n2610 0.120292
R4657 VDD.n2618 VDD.n2614 0.120292
R4658 VDD.n2624 VDD.n2618 0.120292
R4659 VDD.n2628 VDD.n2624 0.120292
R4660 VDD.n2633 VDD.n2628 0.120292
R4661 VDD.n2637 VDD.n2633 0.120292
R4662 VDD.n2641 VDD.n2637 0.120292
R4663 VDD.n2647 VDD.n2641 0.120292
R4664 VDD.n2651 VDD.n2647 0.120292
R4665 VDD.n2655 VDD.n2651 0.120292
R4666 VDD.n2658 VDD.n2655 0.120292
R4667 VDD.n2662 VDD.n2658 0.120292
R4668 VDD.n2666 VDD.n2662 0.120292
R4669 VDD.n2672 VDD.n2666 0.120292
R4670 VDD.n2676 VDD.n2672 0.120292
R4671 VDD.n2701 VDD.n2697 0.120292
R4672 VDD.n2705 VDD.n2701 0.120292
R4673 VDD.n2709 VDD.n2705 0.120292
R4674 VDD.n2714 VDD.n2709 0.120292
R4675 VDD.n2718 VDD.n2714 0.120292
R4676 VDD.n2720 VDD.n2718 0.120292
R4677 VDD.n2720 VDD.n2719 0.120292
R4678 VDD.n2731 VDD.n2601 0.120292
R4679 VDD.n2601 VDD.n2595 0.120292
R4680 VDD.n2595 VDD.n2591 0.120292
R4681 VDD.n2591 VDD.n2587 0.120292
R4682 VDD.n2587 VDD.n2581 0.120292
R4683 VDD.n2581 VDD.n2577 0.120292
R4684 VDD.n2577 VDD.n2572 0.120292
R4685 VDD.n2572 VDD.n2568 0.120292
R4686 VDD.n2568 VDD.n2564 0.120292
R4687 VDD.n2564 VDD.n2558 0.120292
R4688 VDD.n2558 VDD.n2554 0.120292
R4689 VDD.n2554 VDD.n2550 0.120292
R4690 VDD.n2550 VDD.n2547 0.120292
R4691 VDD.n2547 VDD.n2543 0.120292
R4692 VDD.n2543 VDD.n2539 0.120292
R4693 VDD.n2539 VDD.n2533 0.120292
R4694 VDD.n2512 VDD.n2508 0.120292
R4695 VDD.n2508 VDD.n2504 0.120292
R4696 VDD.n2504 VDD.n2500 0.120292
R4697 VDD.n2500 VDD.n2496 0.120292
R4698 VDD.n2496 VDD.n2491 0.120292
R4699 VDD.n2491 VDD.n2487 0.120292
R4700 VDD.n2487 VDD.n0 0.120292
R4701 VDD.n2478 VDD.n2477 0.120292
R4702 VDD.n2477 VDD.n2471 0.120292
R4703 VDD.n2471 VDD.n2467 0.120292
R4704 VDD.n2467 VDD.n2463 0.120292
R4705 VDD.n2463 VDD.n2457 0.120292
R4706 VDD.n2457 VDD.n2453 0.120292
R4707 VDD.n2453 VDD.n2448 0.120292
R4708 VDD.n2448 VDD.n2444 0.120292
R4709 VDD.n2444 VDD.n2440 0.120292
R4710 VDD.n2440 VDD.n2434 0.120292
R4711 VDD.n2434 VDD.n2430 0.120292
R4712 VDD.n2430 VDD.n2426 0.120292
R4713 VDD.n2426 VDD.n2423 0.120292
R4714 VDD.n2423 VDD.n2419 0.120292
R4715 VDD.n2419 VDD.n2415 0.120292
R4716 VDD.n2415 VDD.n2409 0.120292
R4717 VDD.n2388 VDD.n2384 0.120292
R4718 VDD.n2384 VDD.n2380 0.120292
R4719 VDD.n2380 VDD.n2376 0.120292
R4720 VDD.n2376 VDD.n2372 0.120292
R4721 VDD.n2372 VDD.n2367 0.120292
R4722 VDD.n2367 VDD.n2363 0.120292
R4723 VDD.n2363 VDD.n4 0.120292
R4724 VDD.n2354 VDD.n2353 0.120292
R4725 VDD.n2353 VDD.n2347 0.120292
R4726 VDD.n2347 VDD.n2343 0.120292
R4727 VDD.n2343 VDD.n2339 0.120292
R4728 VDD.n2339 VDD.n2333 0.120292
R4729 VDD.n2333 VDD.n2329 0.120292
R4730 VDD.n2329 VDD.n2324 0.120292
R4731 VDD.n2324 VDD.n2320 0.120292
R4732 VDD.n2320 VDD.n2316 0.120292
R4733 VDD.n2316 VDD.n2310 0.120292
R4734 VDD.n2310 VDD.n2306 0.120292
R4735 VDD.n2306 VDD.n2302 0.120292
R4736 VDD.n2302 VDD.n2299 0.120292
R4737 VDD.n2299 VDD.n2295 0.120292
R4738 VDD.n2295 VDD.n2291 0.120292
R4739 VDD.n2291 VDD.n2285 0.120292
R4740 VDD.n2264 VDD.n2260 0.120292
R4741 VDD.n2260 VDD.n2256 0.120292
R4742 VDD.n2256 VDD.n2252 0.120292
R4743 VDD.n2252 VDD.n2248 0.120292
R4744 VDD.n2248 VDD.n2243 0.120292
R4745 VDD.n2231 VDD.n8 0.120292
R4746 VDD.n2222 VDD.n2221 0.120292
R4747 VDD.n2221 VDD.n2215 0.120292
R4748 VDD.n2215 VDD.n2211 0.120292
R4749 VDD.n2211 VDD.n2207 0.120292
R4750 VDD.n2195 VDD.n2190 0.120292
R4751 VDD.n2190 VDD.n2186 0.120292
R4752 VDD.n2186 VDD.n2182 0.120292
R4753 VDD.n2182 VDD.n2176 0.120292
R4754 VDD.n2176 VDD.n2172 0.120292
R4755 VDD.n2172 VDD.n2168 0.120292
R4756 VDD.n2168 VDD.n2165 0.120292
R4757 VDD.n2165 VDD.n2161 0.120292
R4758 VDD.n2161 VDD.n2157 0.120292
R4759 VDD.n2157 VDD.n2151 0.120292
R4760 VDD.n2151 VDD.n2147 0.120292
R4761 VDD.n2147 VDD.n2143 0.120292
R4762 VDD.n2143 VDD.n2137 0.120292
R4763 VDD.n2137 VDD.n2133 0.120292
R4764 VDD.n2133 VDD.n2129 0.120292
R4765 VDD.n2129 VDD.n2125 0.120292
R4766 VDD.n2125 VDD.n2120 0.120292
R4767 VDD.n2120 VDD.n2116 0.120292
R4768 VDD.n2116 VDD.n2107 0.120292
R4769 VDD.n1985 VDD 0.119803
R4770 VDD VDD.n2106 0.119505
R4771 VDD.n2196 VDD.n2195 0.117688
R4772 VDD.n2697 VDD.n2693 0.111177
R4773 VDD.n2513 VDD.n2512 0.111177
R4774 VDD.n2389 VDD.n2388 0.111177
R4775 VDD.n2265 VDD.n2264 0.111177
R4776 VDD.n1245 VDD.n1244 0.108573
R4777 VDD.n638 VDD.n79 0.107271
R4778 VDD.n2677 VDD.n2676 0.107271
R4779 VDD.n2533 VDD.n2529 0.107271
R4780 VDD.n2409 VDD.n2405 0.107271
R4781 VDD.n2285 VDD.n2281 0.107271
R4782 VDD.n2207 VDD.n2203 0.10076
R4783 VDD.n1250 VDD.n1249 0.0981562
R4784 VDD.n1262 VDD.n1260 0.0981562
R4785 VDD.n1272 VDD.n832 0.0981562
R4786 VDD.n1274 VDD.n828 0.0981562
R4787 VDD.n1287 VDD.n1285 0.0981562
R4788 VDD.n1301 VDD.n818 0.0981562
R4789 VDD.n1303 VDD.n814 0.0981562
R4790 VDD.n1317 VDD.n1314 0.0981562
R4791 VDD.n1315 VDD.n806 0.0981562
R4792 VDD.n1338 VDD.n800 0.0981562
R4793 VDD.n1340 VDD.n796 0.0981562
R4794 VDD.n1354 VDD.n1351 0.0981562
R4795 VDD.n1352 VDD.n787 0.0981562
R4796 VDD.n1370 VDD.n1367 0.0981562
R4797 VDD.n1368 VDD.n778 0.0981562
R4798 VDD.n777 VDD.n771 0.0981562
R4799 VDD.n651 VDD.n650 0.0981562
R4800 VDD.n664 VDD.n662 0.0981562
R4801 VDD.n674 VDD.n61 0.0981562
R4802 VDD.n676 VDD.n56 0.0981562
R4803 VDD.n689 VDD.n688 0.0981562
R4804 VDD.n702 VDD.n700 0.0981562
R4805 VDD.n712 VDD.n39 0.0981562
R4806 VDD.n714 VDD.n34 0.0981562
R4807 VDD.n730 VDD.n726 0.0981562
R4808 VDD.n2232 VDD.n2231 0.0981562
R4809 VDD VDD.n2025 0.0968542
R4810 VDD.n1611 VDD 0.0968542
R4811 VDD.n1682 VDD 0.0968542
R4812 VDD.n1764 VDD 0.0968542
R4813 VDD.n1835 VDD 0.0968542
R4814 VDD.n1917 VDD 0.0968542
R4815 VDD.n250 VDD 0.0968542
R4816 VDD.n339 VDD 0.0968542
R4817 VDD.n428 VDD 0.0968542
R4818 VDD.n517 VDD 0.0968542
R4819 VDD.n292 VDD 0.0821977
R4820 VDD.n381 VDD 0.0821977
R4821 VDD.n470 VDD 0.0821977
R4822 VDD.n559 VDD 0.0821977
R4823 VDD.n292 VDD.n291 0.0783056
R4824 VDD.n381 VDD.n380 0.0783056
R4825 VDD.n470 VDD.n469 0.0783056
R4826 VDD.n559 VDD.n558 0.0783056
R4827 VDD.n2682 VDD.n2681 0.076587
R4828 VDD.n2518 VDD.n2517 0.076587
R4829 VDD.n2394 VDD.n2393 0.076587
R4830 VDD.n2270 VDD.n2269 0.076587
R4831 VDD VDD.n2082 0.0603958
R4832 VDD VDD.n2096 0.0603958
R4833 VDD.n2097 VDD 0.0603958
R4834 VDD VDD.n1680 0.0603958
R4835 VDD.n1681 VDD 0.0603958
R4836 VDD.n1755 VDD 0.0603958
R4837 VDD VDD.n1754 0.0603958
R4838 VDD VDD.n1833 0.0603958
R4839 VDD.n1834 VDD 0.0603958
R4840 VDD.n1908 VDD 0.0603958
R4841 VDD VDD.n1907 0.0603958
R4842 VDD VDD.n1984 0.0603958
R4843 VDD.n1057 VDD 0.0603958
R4844 VDD.n1133 VDD 0.0603958
R4845 VDD.n1215 VDD 0.0603958
R4846 VDD.n330 VDD 0.0603958
R4847 VDD VDD.n329 0.0603958
R4848 VDD.n419 VDD 0.0603958
R4849 VDD VDD.n418 0.0603958
R4850 VDD.n508 VDD 0.0603958
R4851 VDD VDD.n507 0.0603958
R4852 VDD VDD.n596 0.0603958
R4853 VDD.n597 VDD 0.0603958
R4854 VDD VDD.n755 0.0603958
R4855 VDD.n756 VDD 0.0603958
R4856 VDD VDD.n764 0.0603958
R4857 VDD VDD.n2731 0.0603958
R4858 VDD.n2478 VDD 0.0603958
R4859 VDD.n2354 VDD 0.0603958
R4860 VDD.n2222 VDD 0.0603958
R4861 VDD.n2684 VDD.n2683 0.0439783
R4862 VDD.n2520 VDD.n2519 0.0439783
R4863 VDD.n2396 VDD.n2395 0.0439783
R4864 VDD.n2272 VDD.n2271 0.0439783
R4865 VDD.n2683 VDD 0.0358261
R4866 VDD.n2519 VDD 0.0358261
R4867 VDD.n2395 VDD 0.0358261
R4868 VDD.n2271 VDD 0.0358261
R4869 VDD.n1394 VDD 0.0356562
R4870 VDD.n741 VDD 0.0343542
R4871 VDD VDD.n1681 0.0239375
R4872 VDD.n1754 VDD 0.0239375
R4873 VDD VDD.n1834 0.0239375
R4874 VDD.n1907 VDD 0.0239375
R4875 VDD.n329 VDD 0.0239375
R4876 VDD.n418 VDD 0.0239375
R4877 VDD.n507 VDD 0.0239375
R4878 VDD VDD.n2105 0.0226354
R4879 VDD VDD.n1402 0.0226354
R4880 VDD.n2243 VDD.n2232 0.0226354
R4881 VDD.n1045 VDD 0.0213333
R4882 VDD VDD.n1132 0.0213333
R4883 VDD.n1203 VDD 0.0213333
R4884 VDD.n2719 VDD 0.0213333
R4885 VDD VDD.n0 0.0213333
R4886 VDD VDD.n4 0.0213333
R4887 VDD VDD.n8 0.0213333
R4888 VDD.n2107 VDD 0.0213333
R4889 VDD.n2203 VDD.n2202 0.0200312
R4890 VDD.n1986 VDD.n1985 0.0141161
R4891 VDD.n79 VDD.n76 0.0135208
R4892 VDD.n651 VDD.n69 0.0135208
R4893 VDD.n664 VDD.n663 0.0135208
R4894 VDD.n675 VDD.n674 0.0135208
R4895 VDD.n56 VDD.n54 0.0135208
R4896 VDD.n689 VDD.n47 0.0135208
R4897 VDD.n702 VDD.n701 0.0135208
R4898 VDD.n713 VDD.n712 0.0135208
R4899 VDD.n34 VDD.n32 0.0135208
R4900 VDD.n730 VDD.n729 0.0135208
R4901 VDD.n2692 VDD.n2677 0.0135208
R4902 VDD.n2529 VDD.n2528 0.0135208
R4903 VDD.n2405 VDD.n2404 0.0135208
R4904 VDD.n2281 VDD.n2280 0.0135208
R4905 VDD.n1245 VDD.n846 0.0122188
R4906 VDD.n1250 VDD.n840 0.0122188
R4907 VDD.n1262 VDD.n1261 0.0122188
R4908 VDD.n1273 VDD.n1272 0.0122188
R4909 VDD.n828 VDD.n826 0.0122188
R4910 VDD.n1287 VDD.n1286 0.0122188
R4911 VDD.n1302 VDD.n1301 0.0122188
R4912 VDD.n814 VDD.n812 0.0122188
R4913 VDD.n1317 VDD.n1316 0.0122188
R4914 VDD.n1326 VDD.n806 0.0122188
R4915 VDD.n1339 VDD.n1338 0.0122188
R4916 VDD.n796 VDD.n794 0.0122188
R4917 VDD.n1354 VDD.n1353 0.0122188
R4918 VDD.n787 VDD.n784 0.0122188
R4919 VDD.n1370 VDD.n1369 0.0122188
R4920 VDD.n1379 VDD.n778 0.0122188
R4921 VDD.n1392 VDD.n771 0.0122188
R4922 VDD.n727 VDD 0.0122188
R4923 VDD.n1249 VDD.n846 0.0109167
R4924 VDD.n1260 VDD.n840 0.0109167
R4925 VDD.n1261 VDD.n832 0.0109167
R4926 VDD.n1274 VDD.n1273 0.0109167
R4927 VDD.n1285 VDD.n826 0.0109167
R4928 VDD.n1286 VDD.n818 0.0109167
R4929 VDD.n1303 VDD.n1302 0.0109167
R4930 VDD.n1314 VDD.n812 0.0109167
R4931 VDD.n1316 VDD.n1315 0.0109167
R4932 VDD.n1326 VDD.n800 0.0109167
R4933 VDD.n1340 VDD.n1339 0.0109167
R4934 VDD.n1351 VDD.n794 0.0109167
R4935 VDD.n1353 VDD.n1352 0.0109167
R4936 VDD.n1367 VDD.n784 0.0109167
R4937 VDD.n1369 VDD.n1368 0.0109167
R4938 VDD.n1379 VDD.n777 0.0109167
R4939 VDD.n1393 VDD.n1392 0.0109167
R4940 VDD VDD.n1393 0.0109167
R4941 VDD.n650 VDD.n76 0.00961458
R4942 VDD.n662 VDD.n69 0.00961458
R4943 VDD.n663 VDD.n61 0.00961458
R4944 VDD.n676 VDD.n675 0.00961458
R4945 VDD.n688 VDD.n54 0.00961458
R4946 VDD.n700 VDD.n47 0.00961458
R4947 VDD.n701 VDD.n39 0.00961458
R4948 VDD.n714 VDD.n713 0.00961458
R4949 VDD.n726 VDD.n32 0.00961458
R4950 VDD.n729 VDD.n727 0.00961458
R4951 VDD.n2693 VDD.n2692 0.00961458
R4952 VDD.n2528 VDD.n2513 0.00961458
R4953 VDD.n2404 VDD.n2389 0.00961458
R4954 VDD.n2280 VDD.n2265 0.00961458
R4955 VDD.n2106 VDD.n1986 0.0093414
R4956 VDD.n2684 VDD.n2682 0.00321739
R4957 VDD.n2520 VDD.n2518 0.00321739
R4958 VDD.n2396 VDD.n2394 0.00321739
R4959 VDD.n2272 VDD.n2270 0.00321739
R4960 VDD.n2202 VDD.n2196 0.00310417
R4961 VDD.n2106 VDD 0.00195147
R4962 check[1].n3 check[1].t5 331.51
R4963 check[1].n1 check[1].t2 280.899
R4964 check[1].n1 check[1].t3 216.238
R4965 check[1].n3 check[1].t4 209.403
R4966 check[1].n0 check[1].t0 207.373
R4967 check[1].n4 check[1].n3 76.0005
R4968 check[1].n7 check[1].n6 50.467
R4969 check[1].n2 check[1].n1 35.7166
R4970 check[1].n8 check[1].t1 33.1309
R4971 check[1].n5 check[1].n2 32.9012
R4972 check[1].n7 check[1] 15.9389
R4973 check[1].n6 check[1] 12.062
R4974 check[1] check[1].n0 9.01934
R4975 check[1].n5 check[1] 8.68932
R4976 check[1] check[1].n4 8.58587
R4977 check[1] check[1].n8 8.00801
R4978 check[1].n0 check[1] 7.45876
R4979 check[1].n6 check[1].n5 3.04357
R4980 check[1].n2 check[1] 2.56973
R4981 check[1].n4 check[1] 2.02977
R4982 check[1].n8 check[1].n7 1.94232
R4983 D[0].n8 D[0].t2 269.921
R4984 D[0].n8 D[0].t3 234.573
R4985 D[0].n7 D[0].t0 207.373
R4986 D[0].n9 D[0].n8 76.0005
R4987 D[0].n14 D[0].t1 33.3405
R4988 D[0].n12 D[0].n11 26.2261
R4989 D[0].n11 D[0] 19.418
R4990 D[0].n11 D[0].n10 14.9338
R4991 D[0] D[0].n14 9.32876
R4992 D[0] D[0].n7 9.01934
R4993 D[0].n7 D[0] 7.45876
R4994 D[0].n3 D[0] 6.42
R4995 D[0].n10 D[0] 5.9498
R4996 D[0].n9 D[0] 4.68782
R4997 D[0].n13 D[0].n12 3.50069
R4998 D[0].n12 D[0].n6 2.83165
R4999 D[0].n5 D[0].n1 2.26284
R5000 D[0].n4 D[0].n3 2.23869
R5001 D[0].n10 D[0].n9 1.62304
R5002 D[0].n14 D[0].n13 0.391757
R5003 D[0].n4 D[0].n2 0.0213333
R5004 D[0].n6 D[0].n0 0.0099697
R5005 D[0].n5 D[0].n4 0.00195195
R5006 D[0].n6 D[0].n5 0.00194159
R5007 eob.n10 eob.t11 331.51
R5008 eob.n4 eob 298.998
R5009 eob.n5 eob.n4 292.5
R5010 eob.n0 eob.t8 230.576
R5011 eob.n10 eob.t10 209.403
R5012 eob.n3 eob.n1 180.082
R5013 eob.n0 eob.t9 158.275
R5014 eob.n3 eob.n2 124.501
R5015 eob.n8 eob.n7 92.5005
R5016 eob eob.n0 82.6672
R5017 eob.n11 eob.n10 76.0005
R5018 eob.n6 eob.n3 36.0005
R5019 eob.n4 eob.t0 26.5955
R5020 eob.n4 eob.t2 26.5955
R5021 eob.n1 eob.t3 26.5955
R5022 eob.n1 eob.t1 26.5955
R5023 eob eob.n13 25.8571
R5024 eob.n7 eob.t7 24.9236
R5025 eob.n7 eob.t6 24.9236
R5026 eob.n2 eob.t5 24.9236
R5027 eob.n2 eob.t4 24.9236
R5028 eob.n12 eob.n9 11.9351
R5029 eob.n12 eob 11.6575
R5030 eob.n6 eob 10.2405
R5031 eob.n13 eob.n12 9.41338
R5032 eob eob.n11 8.58587
R5033 eob eob.n5 8.46819
R5034 eob eob.n8 8.07435
R5035 eob.n13 eob 6.9444
R5036 eob.n8 eob 5.31742
R5037 eob.n5 eob 4.92358
R5038 eob.n9 eob 2.95435
R5039 eob.n11 eob 2.02977
R5040 eob.n9 eob.n6 0.197423
R5041 VSS.n4120 VSS 52235.6
R5042 VSS.n3839 VSS 8025.31
R5043 VSS VSS.n3839 5751.89
R5044 VSS.n1246 VSS.n1240 2560.8
R5045 VSS.n1833 VSS.n1832 2487.33
R5046 VSS.n4121 VSS.n4120 1234.15
R5047 VSS.n3839 VSS 1073.17
R5048 VSS.n4235 VSS 1019.51
R5049 VSS.n3495 VSS 1019.51
R5050 VSS.n3609 VSS 1019.51
R5051 VSS.n3723 VSS 1019.51
R5052 VSS VSS.n3853 643.275
R5053 VSS VSS.t417 630.489
R5054 VSS VSS.t6 630.489
R5055 VSS VSS.t419 630.489
R5056 VSS VSS.t421 630.489
R5057 VSS.t429 VSS 630.489
R5058 VSS.n4210 VSS.t264 603.659
R5059 VSS.n3470 VSS.t509 603.659
R5060 VSS.n3584 VSS.t368 603.659
R5061 VSS.n3698 VSS.t493 603.659
R5062 VSS.n3812 VSS.t22 603.659
R5063 VSS.n4125 VSS.t332 590.245
R5064 VSS.n4218 VSS.t390 590.245
R5065 VSS.t417 VSS.n4231 590.245
R5066 VSS.n1 VSS.t273 590.245
R5067 VSS.n3478 VSS.t149 590.245
R5068 VSS.t6 VSS.n3493 590.245
R5069 VSS.n3499 VSS.t561 590.245
R5070 VSS.n3592 VSS.t624 590.245
R5071 VSS.t419 VSS.n3607 590.245
R5072 VSS.n3613 VSS.t99 590.245
R5073 VSS.n3706 VSS.t370 590.245
R5074 VSS.t421 VSS.n3721 590.245
R5075 VSS.n3727 VSS.t211 590.245
R5076 VSS.n3820 VSS.t495 590.245
R5077 VSS.n3829 VSS.t429 590.245
R5078 VSS.n3074 VSS 574.659
R5079 VSS.n4131 VSS.t614 550
R5080 VSS.n3391 VSS.t94 550
R5081 VSS.n3505 VSS.t340 550
R5082 VSS.n3619 VSS.t634 550
R5083 VSS.n3733 VSS.t201 550
R5084 VSS.n4231 VSS.t266 536.586
R5085 VSS.n3493 VSS.t511 536.586
R5086 VSS.n3607 VSS.t366 536.586
R5087 VSS.n3721 VSS.t491 536.586
R5088 VSS.n3829 VSS.t24 536.586
R5089 VSS.n3372 VSS.n3369 533.059
R5090 VSS.n3855 VSS.n3852 533.059
R5091 VSS.n3496 VSS.n3389 533.059
R5092 VSS.n3610 VSS.n3387 533.059
R5093 VSS.n3724 VSS.n3385 533.059
R5094 VSS.n4157 VSS.t662 509.757
R5095 VSS.n3417 VSS.t655 509.757
R5096 VSS.n3531 VSS.t272 509.757
R5097 VSS.n3645 VSS.t134 509.757
R5098 VSS.n3759 VSS.t654 509.757
R5099 VSS.n4139 VSS.t610 496.341
R5100 VSS.n3399 VSS.t96 496.341
R5101 VSS.n3513 VSS.t342 496.341
R5102 VSS.n3627 VSS.t636 496.341
R5103 VSS.n3741 VSS.t197 496.341
R5104 VSS.n3062 VSS 488.889
R5105 VSS.n3063 VSS.n3058 475.118
R5106 VSS.n4145 VSS.t388 456.099
R5107 VSS.n3405 VSS.t303 456.099
R5108 VSS.n3519 VSS.t445 456.099
R5109 VSS.n3633 VSS.t55 456.099
R5110 VSS.n3747 VSS.t231 456.099
R5111 VSS.n2354 VSS.n110 434.56
R5112 VSS.n2705 VSS.n98 434.56
R5113 VSS.n2030 VSS 428.851
R5114 VSS.n2356 VSS 428.851
R5115 VSS.n2707 VSS 428.851
R5116 VSS.n4206 VSS.t91 415.854
R5117 VSS.n3466 VSS.t591 415.854
R5118 VSS.n3580 VSS.t559 415.854
R5119 VSS.n3694 VSS.t500 415.854
R5120 VSS.n3808 VSS.t663 415.854
R5121 VSS.n4153 VSS.t485 402.44
R5122 VSS.n3413 VSS.t452 402.44
R5123 VSS.n3527 VSS.t101 402.44
R5124 VSS.n3641 VSS.t209 402.44
R5125 VSS.n3755 VSS.t441 402.44
R5126 VSS.n1226 VSS.t450 396
R5127 VSS.n1125 VSS.t578 396
R5128 VSS.t589 VSS.n1245 387.2
R5129 VSS.n123 VSS.t293 387.2
R5130 VSS.n132 VSS.t26 387.2
R5131 VSS.t73 VSS.n1143 387.2
R5132 VSS.n138 VSS.t298 387.2
R5133 VSS.n987 VSS.t425 387.2
R5134 VSS.n678 VSS.t103 387.2
R5135 VSS.n369 VSS.t105 387.2
R5136 VSS.n2028 VSS.n116 382.413
R5137 VSS.n3858 VSS.t384 377.389
R5138 VSS.n3844 VSS.t20 377.389
R5139 VSS.n3844 VSS.t616 377.389
R5140 VSS.n1837 VSS.t579 377.389
R5141 VSS.n3935 VSS.t557 368.812
R5142 VSS.n3906 VSS.t551 368.812
R5143 VSS.n3864 VSS.t608 368.812
R5144 VSS.n4202 VSS.t159 362.195
R5145 VSS.n3462 VSS.t398 362.195
R5146 VSS.n3576 VSS.t526 362.195
R5147 VSS.n3690 VSS.t61 362.195
R5148 VSS.n3804 VSS.t516 362.195
R5149 VSS.n1152 VSS.t75 360.8
R5150 VSS.n3964 VSS.t135 360.235
R5151 VSS.n1245 VSS.t447 352
R5152 VSS.n1143 VSS.t576 352
R5153 VSS.n1015 VSS.t115 352
R5154 VSS.n706 VSS.t379 352
R5155 VSS.n397 VSS.t145 352
R5156 VSS.n3864 VSS.t606 351.658
R5157 VSS.n1843 VSS.t585 351.658
R5158 VSS.n2275 VSS.t43 343.08
R5159 VSS.n2626 VSS.t17 343.08
R5160 VSS.n2977 VSS.t114 343.08
R5161 VSS.n3978 VSS.t407 334.503
R5162 VSS.n1173 VSS.t327 334.401
R5163 VSS.n305 VSS.t453 334.401
R5164 VSS.n86 VSS.t675 327.046
R5165 VSS.n1869 VSS.t550 325.926
R5166 VSS.n127 VSS.t79 325.601
R5167 VSS.n1851 VSS.t581 317.349
R5168 VSS.n2261 VSS.t524 308.772
R5169 VSS.n2612 VSS.t506 308.772
R5170 VSS.n2963 VSS.t638 308.772
R5171 VSS.n1161 VSS.t501 299.2
R5172 VSS.n3893 VSS.n3892 292.5
R5173 VSS.n3892 VSS.n3891 292.5
R5174 VSS.n3890 VSS.n3889 292.5
R5175 VSS.n3889 VSS.n3888 292.5
R5176 VSS.n3887 VSS.n3886 292.5
R5177 VSS.n3886 VSS.n3885 292.5
R5178 VSS.n3884 VSS.n3883 292.5
R5179 VSS.n3883 VSS.n3882 292.5
R5180 VSS.n3881 VSS.n3880 292.5
R5181 VSS.n3880 VSS.n3879 292.5
R5182 VSS.n3878 VSS.n3877 292.5
R5183 VSS.n3877 VSS.n3876 292.5
R5184 VSS.n3875 VSS.n3874 292.5
R5185 VSS.n3874 VSS.n3873 292.5
R5186 VSS.n1857 VSS.t53 291.618
R5187 VSS.n1222 VSS.t268 272.8
R5188 VSS.n1121 VSS.t349 272.8
R5189 VSS.n1971 VSS.t32 265.887
R5190 VSS VSS.t589 264
R5191 VSS.n1169 VSS.t1 264
R5192 VSS VSS.t73 264
R5193 VSS VSS.t71 264
R5194 VSS VSS.t415 264
R5195 VSS.n291 VSS.t465 264
R5196 VSS.n79 VSS.t674 260.281
R5197 VSS VSS.t652 257.31
R5198 VSS.n1865 VSS.t618 257.31
R5199 VSS.n1059 VSS.t184 246.4
R5200 VSS.n968 VSS.t180 246.4
R5201 VSS.n750 VSS.t567 246.4
R5202 VSS.n659 VSS.t569 246.4
R5203 VSS.n441 VSS.t291 246.4
R5204 VSS.n350 VSS.t287 246.4
R5205 VSS.n3371 VSS 242.143
R5206 VSS.n4167 VSS.t612 241.464
R5207 VSS.n3427 VSS.t92 241.464
R5208 VSS.n3541 VSS.t338 241.464
R5209 VSS.n3655 VSS.t632 241.464
R5210 VSS.n3769 VSS.t199 241.464
R5211 VSS.n1218 VSS.t344 237.601
R5212 VSS.n1117 VSS.t175 237.601
R5213 VSS.n1013 VSS.t189 237.601
R5214 VSS.n704 VSS.t302 237.601
R5215 VSS.n395 VSS.t179 237.601
R5216 VSS.n1808 VSS.t438 237.126
R5217 VSS.n1707 VSS.t15 237.126
R5218 VSS.n1606 VSS.t331 237.126
R5219 VSS.n1505 VSS.t405 237.126
R5220 VSS.n1404 VSS.t670 237.126
R5221 VSS.t18 VSS.n1826 231.857
R5222 VSS.n1251 VSS.t408 231.857
R5223 VSS.n1260 VSS.t249 231.857
R5224 VSS.t587 VSS.n1725 231.857
R5225 VSS.n1266 VSS.t124 231.857
R5226 VSS.n1275 VSS.t536 231.857
R5227 VSS.t386 VSS.n1624 231.857
R5228 VSS.n1281 VSS.t427 231.857
R5229 VSS.n1290 VSS.t354 231.857
R5230 VSS.t626 VSS.n1523 231.857
R5231 VSS.n1296 VSS.t191 231.857
R5232 VSS.n1305 VSS.t128 231.857
R5233 VSS.t34 VSS.n1422 231.857
R5234 VSS.n1311 VSS.t382 231.857
R5235 VSS.n1320 VSS.t563 231.857
R5236 VSS.n1961 VSS.t195 231.579
R5237 VSS.n81 VSS.t65 229.315
R5238 VSS.n1073 VSS.t575 220
R5239 VSS.n920 VSS.t111 220
R5240 VSS.n764 VSS.t109 220
R5241 VSS.n611 VSS.t487 220
R5242 VSS.n455 VSS.t489 220
R5243 VSS.n1734 VSS.t165 216.048
R5244 VSS.n1633 VSS.t372 216.048
R5245 VSS.n1532 VSS.t47 216.048
R5246 VSS.n1431 VSS.t656 216.048
R5247 VSS.n1330 VSS.t309 216.048
R5248 VSS VSS.n4234 214.635
R5249 VSS VSS.n3494 214.635
R5250 VSS VSS.n3608 214.635
R5251 VSS VSS.n3722 214.635
R5252 VSS VSS.n3838 214.635
R5253 VSS.n154 VSS.t182 211.201
R5254 VSS.n208 VSS.t565 211.201
R5255 VSS.n262 VSS.t289 211.201
R5256 VSS.n1826 VSS.t439 210.779
R5257 VSS.n1725 VSS.t13 210.779
R5258 VSS.n1624 VSS.t328 210.779
R5259 VSS.n1523 VSS.t402 210.779
R5260 VSS.n1422 VSS.t671 210.779
R5261 VSS.n3933 VSS.t553 205.849
R5262 VSS.n3904 VSS.t555 205.849
R5263 VSS.n4171 VSS.t265 201.22
R5264 VSS.n3431 VSS.t510 201.22
R5265 VSS.n3545 VSS.t369 201.22
R5266 VSS.n3659 VSS.t494 201.22
R5267 VSS.n3773 VSS.t23 201.22
R5268 VSS.n1755 VSS.t148 200.24
R5269 VSS.n1654 VSS.t434 200.24
R5270 VSS.n1553 VSS.t665 200.24
R5271 VSS.n1452 VSS.t98 200.24
R5272 VSS.n1351 VSS.t364 200.24
R5273 VSS.n84 VSS.t68 198.691
R5274 VSS.n1255 VSS.t163 194.97
R5275 VSS.n1270 VSS.t376 194.97
R5276 VSS.n1285 VSS.t51 194.97
R5277 VSS.n1300 VSS.t660 194.97
R5278 VSS.n1315 VSS.t307 194.97
R5279 VSS.n1045 VSS.t243 193.601
R5280 VSS.n736 VSS.t239 193.601
R5281 VSS.n427 VSS.t227 193.601
R5282 VSS.n2899 VSS.t641 190.337
R5283 VSS.n2548 VSS.t505 190.337
R5284 VSS.n2197 VSS.t523 190.337
R5285 VSS.n1913 VSS.t194 190.337
R5286 VSS.n1199 VSS.t347 190.337
R5287 VSS.n1098 VSS.t174 190.337
R5288 VSS.n808 VSS.t549 190.337
R5289 VSS.n499 VSS.t393 190.337
R5290 VSS.n1781 VSS.t337 190.337
R5291 VSS.n1680 VSS.t152 190.337
R5292 VSS.n1579 VSS.t651 190.337
R5293 VSS.n1478 VSS.t11 190.337
R5294 VSS.n1377 VSS.t667 190.337
R5295 VSS.n4183 VSS.t162 190.337
R5296 VSS.n3443 VSS.t401 190.337
R5297 VSS.n3557 VSS.t529 190.337
R5298 VSS.n3671 VSS.t64 190.337
R5299 VSS.n3785 VSS.t515 190.337
R5300 VSS.n300 VSS.t454 190.065
R5301 VSS.n119 VSS.t315 188.695
R5302 VSS.n106 VSS.t44 188.695
R5303 VSS.n94 VSS.t177 188.695
R5304 VSS.n3059 VSS.t66 188.695
R5305 VSS.n168 VSS.t252 184.8
R5306 VSS.n903 VSS.t130 184.8
R5307 VSS.n222 VSS.t187 184.8
R5308 VSS.n594 VSS.t411 184.8
R5309 VSS.n276 VSS.t118 184.8
R5310 VSS.n4108 VSS.t57 180.118
R5311 VSS.n3992 VSS.t622 180.118
R5312 VSS.n1987 VSS.t311 180.118
R5313 VSS.n2301 VSS.t254 180.118
R5314 VSS.n2652 VSS.t597 180.118
R5315 VSS.n3003 VSS.t206 180.118
R5316 VSS.n1743 VSS.t630 179.162
R5317 VSS.n1642 VSS.t413 179.162
R5318 VSS.n1541 VSS.t423 179.162
R5319 VSS.n1440 VSS.t530 179.162
R5320 VSS.n1339 VSS.t628 179.162
R5321 VSS.n3346 VSS 178.422
R5322 VSS.n1804 VSS.t247 163.353
R5323 VSS.n1703 VSS.t646 163.353
R5324 VSS.n1602 VSS.t593 163.353
R5325 VSS.n1501 VSS.t108 163.353
R5326 VSS.n1400 VSS.t170 163.353
R5327 VSS.n4163 VSS.t233 160.976
R5328 VSS.n3423 VSS.t223 160.976
R5329 VSS.n3537 VSS.t215 160.976
R5330 VSS.n3651 VSS.t245 160.976
R5331 VSS.n3765 VSS.t431 160.976
R5332 VSS.n1183 VSS.t77 158.4
R5333 VSS.n889 VSS.t110 158.4
R5334 VSS.n580 VSS.t490 158.4
R5335 VSS VSS.t18 158.084
R5336 VSS.n1751 VSS.t397 158.084
R5337 VSS VSS.t587 158.084
R5338 VSS.n1650 VSS.t31 158.084
R5339 VSS VSS.t386 158.084
R5340 VSS.n1549 VSS.t301 158.084
R5341 VSS VSS.t626 158.084
R5342 VSS.n1448 VSS.t600 158.084
R5343 VSS VSS.t34 158.084
R5344 VSS.n1347 VSS.t642 158.084
R5345 VSS.n4089 VSS.t406 154.387
R5346 VSS.n1879 VSS.t583 154.387
R5347 VSS.n1998 VSS.t126 154.387
R5348 VSS.n2039 VSS.t435 154.387
R5349 VSS.n2217 VSS.t534 154.387
R5350 VSS.n2245 VSS.t573 154.387
R5351 VSS.n2311 VSS.t380 154.387
R5352 VSS.n2369 VSS.t620 154.387
R5353 VSS.n2568 VSS.t271 154.387
R5354 VSS.n2596 VSS.t84 154.387
R5355 VSS.n2662 VSS.t352 154.387
R5356 VSS.n2720 VSS.t121 154.387
R5357 VSS.n2919 VSS.t533 154.387
R5358 VSS.n2947 VSS.t4 154.387
R5359 VSS.n3013 VSS.t69 154.387
R5360 VSS.n3371 VSS.t644 152.934
R5361 VSS.t71 VSS.n936 149.601
R5362 VSS.t415 VSS.n627 149.601
R5363 VSS.n3854 VSS 145.81
R5364 VSS.n1896 VSS.n1895 145.81
R5365 VSS.n1906 VSS.n1905 145.81
R5366 VSS.n1916 VSS.n1915 145.81
R5367 VSS.n1926 VSS.n1925 145.81
R5368 VSS.n1936 VSS.n1935 145.81
R5369 VSS.n1946 VSS.n1945 145.81
R5370 VSS.n1958 VSS.n1957 145.81
R5371 VSS.n1968 VSS.n1967 145.81
R5372 VSS.n1978 VSS.n1977 145.81
R5373 VSS.n1988 VSS.n1987 145.81
R5374 VSS.n1999 VSS.n1998 145.81
R5375 VSS.n2008 VSS.n2007 145.81
R5376 VSS.n2019 VSS.n2018 145.81
R5377 VSS.n120 VSS.n119 145.81
R5378 VSS.n2031 VSS.n2030 145.81
R5379 VSS.n2040 VSS.n2039 145.81
R5380 VSS.n2052 VSS.n2051 145.81
R5381 VSS.n2062 VSS.n2061 145.81
R5382 VSS.n2073 VSS.n2072 145.81
R5383 VSS.n2083 VSS.n2082 145.81
R5384 VSS.n2093 VSS.n2092 145.81
R5385 VSS.n2103 VSS.n2102 145.81
R5386 VSS VSS.n3073 145.81
R5387 VSS.n40 VSS.t133 145.303
R5388 VSS.n2003 VSS.t127 145.203
R5389 VSS.n126 VSS.t294 145.203
R5390 VSS.n141 VSS.t299 145.203
R5391 VSS.n1254 VSS.t409 145.203
R5392 VSS.n1269 VSS.t125 145.203
R5393 VSS.n1284 VSS.t428 145.203
R5394 VSS.n1299 VSS.t192 145.203
R5395 VSS.n1314 VSS.t383 145.203
R5396 VSS.n4221 VSS.t391 145.203
R5397 VSS.n3481 VSS.t150 145.203
R5398 VSS.n3595 VSS.t625 145.203
R5399 VSS.n3709 VSS.t371 145.203
R5400 VSS.n3823 VSS.t496 145.203
R5401 VSS.n3021 VSS.t70 144.49
R5402 VSS.n2670 VSS.t353 144.49
R5403 VSS.n2319 VSS.t381 144.49
R5404 VSS.n195 VSS.t131 144.49
R5405 VSS.n249 VSS.t412 144.49
R5406 VSS.n1800 VSS.t334 142.275
R5407 VSS.n1699 VSS.t153 142.275
R5408 VSS.n1598 VSS.t648 142.275
R5409 VSS.n1497 VSS.t8 142.275
R5410 VSS.n1396 VSS.t668 142.275
R5411 VSS.n3363 VSS.t350 140.189
R5412 VSS.n3375 VSS.t171 140.189
R5413 VSS VSS.n2029 137.232
R5414 VSS.n3195 VSS.t471 133.816
R5415 VSS.n1187 VSS.t449 132
R5416 VSS.n3840 VSS 128.655
R5417 VSS.n2051 VSS.t40 128.655
R5418 VSS.n2383 VSS.t141 128.655
R5419 VSS.n2734 VSS.t323 128.655
R5420 VSS.n3363 VSS.t360 127.445
R5421 VSS.n4188 VSS.t486 120.733
R5422 VSS.n4196 VSS.t235 120.733
R5423 VSS.n3448 VSS.t451 120.733
R5424 VSS.n3456 VSS.t237 120.733
R5425 VSS.n3562 VSS.t102 120.733
R5426 VSS.n3570 VSS.t221 120.733
R5427 VSS.n3676 VSS.t210 120.733
R5428 VSS.n3684 VSS.t213 120.733
R5429 VSS.n3790 VSS.t442 120.733
R5430 VSS.n3798 VSS.t542 120.733
R5431 VSS.n4118 VSS.n4117 120.079
R5432 VSS.n4110 VSS.n4109 120.079
R5433 VSS.n4091 VSS.n4090 120.079
R5434 VSS.n4077 VSS.n4076 120.079
R5435 VSS.n4061 VSS.n4060 120.079
R5436 VSS.n4049 VSS.n4048 120.079
R5437 VSS.n4035 VSS.n4034 120.079
R5438 VSS.n4021 VSS.n4020 120.079
R5439 VSS.n34 VSS.n33 120.079
R5440 VSS.n4004 VSS.n4003 120.079
R5441 VSS.n3992 VSS.n3991 120.079
R5442 VSS.n3978 VSS.n3977 120.079
R5443 VSS.n3964 VSS.n3963 120.079
R5444 VSS.n3949 VSS.n3948 120.079
R5445 VSS.n3935 VSS.n3934 120.079
R5446 VSS.n3920 VSS.n3919 120.079
R5447 VSS.n3906 VSS.n3905 120.079
R5448 VSS.n48 VSS.n47 120.079
R5449 VSS.n2018 VSS.t313 120.079
R5450 VSS.n2189 VSS.t522 120.079
R5451 VSS.n2338 VSS.t256 120.079
R5452 VSS.n2540 VSS.t504 120.079
R5453 VSS.n2689 VSS.t595 120.079
R5454 VSS.n2891 VSS.t640 120.079
R5455 VSS.n3040 VSS.t204 120.079
R5456 VSS.n65 VSS.n64 116.219
R5457 VSS.n3094 VSS.n3093 116.219
R5458 VSS.n3124 VSS.n3123 116.219
R5459 VSS.n3153 VSS.n3152 116.219
R5460 VSS.n3183 VSS.n3173 116.219
R5461 VSS.n3206 VSS.n3203 116.219
R5462 VSS.n3234 VSS.n3233 116.219
R5463 VSS.n3259 VSS.n3258 116.219
R5464 VSS.n3289 VSS.n3288 116.219
R5465 VSS.n3319 VSS.n3318 116.219
R5466 VSS.n3342 VSS.t282 114.775
R5467 VSS.n3953 VSS.n3952 114.749
R5468 VSS.n2956 VSS.n2955 113.207
R5469 VSS.n2605 VSS.n2604 113.207
R5470 VSS.n2254 VSS.n2253 113.207
R5471 VSS.n1954 VSS.n1953 113.207
R5472 VSS.n1217 VSS.n1216 113.207
R5473 VSS.n1116 VSS.n1115 113.207
R5474 VSS.n865 VSS.n864 113.207
R5475 VSS.n556 VSS.n555 113.207
R5476 VSS.n1799 VSS.n1798 113.207
R5477 VSS.n1698 VSS.n1697 113.207
R5478 VSS.n1597 VSS.n1596 113.207
R5479 VSS.n1496 VSS.n1495 113.207
R5480 VSS.n1395 VSS.n1394 113.207
R5481 VSS.n4201 VSS.n4200 113.207
R5482 VSS.n3461 VSS.n3460 113.207
R5483 VSS.n3575 VSS.n3574 113.207
R5484 VSS.n3689 VSS.n3688 113.207
R5485 VSS.n3803 VSS.n3802 113.207
R5486 VSS.t652 VSS.n4119 111.501
R5487 VSS.n22 VSS.t88 111.501
R5488 VSS.n3362 VSS.n3361 109.3
R5489 VSS.n2047 VSS.n2046 109.231
R5490 VSS.n1841 VSS.n1840 109.231
R5491 VSS.n136 VSS.n135 109.231
R5492 VSS.n1264 VSS.n1263 109.231
R5493 VSS.n1279 VSS.n1278 109.231
R5494 VSS.n1294 VSS.n1293 109.231
R5495 VSS.n1309 VSS.n1308 109.231
R5496 VSS.n1324 VSS.n1323 109.231
R5497 VSS.n5 VSS.n4 109.231
R5498 VSS.n3503 VSS.n3502 109.231
R5499 VSS.n3617 VSS.n3616 109.231
R5500 VSS.n3731 VSS.n3730 109.231
R5501 VSS.n4129 VSS.n4128 109.231
R5502 VSS.n2726 VSS.n2725 108.416
R5503 VSS.n2375 VSS.n2374 108.416
R5504 VSS.n162 VSS.n152 108.416
R5505 VSS.n216 VSS.n206 108.416
R5506 VSS.n270 VSS.n260 108.416
R5507 VSS.n3211 VSS.t461 108.328
R5508 VSS.n3355 VSS.n3354 108.254
R5509 VSS.n2078 VSS.n2077 107.478
R5510 VSS.n2024 VSS.n2023 107.478
R5511 VSS.n1855 VSS.n1854 107.478
R5512 VSS.n1242 VSS.n1241 107.478
R5513 VSS.n131 VSS.n130 107.478
R5514 VSS.n1140 VSS.n1139 107.478
R5515 VSS.n3379 VSS.n3378 107.478
R5516 VSS.n3862 VSS.n3861 107.478
R5517 VSS.n3848 VSS.n3847 107.478
R5518 VSS.n1259 VSS.n1258 107.478
R5519 VSS.n1722 VSS.n1721 107.478
R5520 VSS.n1274 VSS.n1273 107.478
R5521 VSS.n1621 VSS.n1620 107.478
R5522 VSS.n1289 VSS.n1288 107.478
R5523 VSS.n1520 VSS.n1519 107.478
R5524 VSS.n1304 VSS.n1303 107.478
R5525 VSS.n1419 VSS.n1418 107.478
R5526 VSS.n1319 VSS.n1318 107.478
R5527 VSS.n1823 VSS.n1822 107.478
R5528 VSS.n4143 VSS.n4142 107.478
R5529 VSS.n4228 VSS.n7 107.478
R5530 VSS.n3403 VSS.n3402 107.478
R5531 VSS.n3490 VSS.n3390 107.478
R5532 VSS.n3517 VSS.n3516 107.478
R5533 VSS.n3604 VSS.n3388 107.478
R5534 VSS.n3631 VSS.n3630 107.478
R5535 VSS.n3718 VSS.n3386 107.478
R5536 VSS.n3745 VSS.n3744 107.478
R5537 VSS.n3833 VSS.n3832 107.478
R5538 VSS.n71 VSS.t498 107.195
R5539 VSS.n3048 VSS.n3039 106.731
R5540 VSS.n2767 VSS.n2758 106.731
R5541 VSS.n2697 VSS.n2688 106.731
R5542 VSS.n2416 VSS.n2407 106.731
R5543 VSS.n2346 VSS.n2337 106.731
R5544 VSS.n151 VSS.n142 106.731
R5545 VSS.n931 VSS.n182 106.731
R5546 VSS.n205 VSS.n196 106.731
R5547 VSS.n622 VSS.n236 106.731
R5548 VSS.n259 VSS.n250 106.731
R5549 VSS.n4105 VSS.n13 106.731
R5550 VSS.n27 VSS.n15 106.731
R5551 VSS.n2837 VSS.n2836 106.038
R5552 VSS.n2486 VSS.n2485 106.038
R5553 VSS.n2135 VSS.n2134 106.038
R5554 VSS.n1874 VSS.n1873 106.038
R5555 VSS.n1178 VSS.n1177 106.038
R5556 VSS.n1038 VSS.n1037 106.038
R5557 VSS.n729 VSS.n728 106.038
R5558 VSS.n420 VSS.n419 106.038
R5559 VSS.n1760 VSS.n1759 106.038
R5560 VSS.n1659 VSS.n1658 106.038
R5561 VSS.n1558 VSS.n1557 106.038
R5562 VSS.n1457 VSS.n1456 106.038
R5563 VSS.n1356 VSS.n1355 106.038
R5564 VSS.n4162 VSS.n4161 106.038
R5565 VSS.n3422 VSS.n3421 106.038
R5566 VSS.n3536 VSS.n3535 106.038
R5567 VSS.n3650 VSS.n3649 106.038
R5568 VSS.n3764 VSS.n3763 106.038
R5569 VSS.n56 VSS.t357 105.835
R5570 VSS.n1179 VSS.t225 105.6
R5571 VSS.n3895 VSS.t552 104.103
R5572 VSS.n3872 VSS.t609 103.968
R5573 VSS.n1875 VSS.t319 102.924
R5574 VSS.n2115 VSS.t87 102.924
R5575 VSS.n2466 VSS.t190 102.924
R5576 VSS.n2817 VSS.t186 102.924
R5577 VSS.n3357 VSS.t358 101.956
R5578 VSS.n1887 VSS.n1884 98.5005
R5579 VSS.n1897 VSS.n1894 98.5005
R5580 VSS.n1907 VSS.n1904 98.5005
R5581 VSS.n1917 VSS.n1914 98.5005
R5582 VSS.n1927 VSS.n1924 98.5005
R5583 VSS.n1937 VSS.n1934 98.5005
R5584 VSS.n1947 VSS.n1944 98.5005
R5585 VSS.n1959 VSS.n1956 98.5005
R5586 VSS.n1969 VSS.n1966 98.5005
R5587 VSS.n1979 VSS.n1976 98.5005
R5588 VSS.n1989 VSS.n1986 98.5005
R5589 VSS.n2000 VSS.n1997 98.5005
R5590 VSS.n2009 VSS.n2006 98.5005
R5591 VSS.n2020 VSS.n2017 98.5005
R5592 VSS.n121 VSS.n118 98.5005
R5593 VSS.n2032 VSS.n116 98.5005
R5594 VSS.n2053 VSS.n2050 98.5005
R5595 VSS.n2063 VSS.n2060 98.5005
R5596 VSS.n2074 VSS.n2071 98.5005
R5597 VSS.n2084 VSS.n2081 98.5005
R5598 VSS.n2094 VSS.n2091 98.5005
R5599 VSS.n2104 VSS.n2101 98.5005
R5600 VSS.n937 VSS 96.8005
R5601 VSS.n628 VSS 96.8005
R5602 VSS.n1765 VSS.t167 94.8508
R5603 VSS.n1664 VSS.t374 94.8508
R5604 VSS.n1563 VSS.t49 94.8508
R5605 VSS.n1462 VSS.t658 94.8508
R5606 VSS.n1361 VSS.t305 94.8508
R5607 VSS.t312 VSS.n1885 94.3475
R5608 VSS.n2072 VSS.t36 94.3475
R5609 VSS.n2175 VSS.t42 94.3475
R5610 VSS.n2408 VSS.t143 94.3475
R5611 VSS.n2526 VSS.t16 94.3475
R5612 VSS.n2759 VSS.t325 94.3475
R5613 VSS.n2877 VSS.t113 94.3475
R5614 VSS.n1087 VSS.n1086 88.0005
R5615 VSS.n1073 VSS.n1072 88.0005
R5616 VSS.n1059 VSS.n1058 88.0005
R5617 VSS.n1045 VSS.n1044 88.0005
R5618 VSS.n1029 VSS.n1028 88.0005
R5619 VSS.n1015 VSS.n1014 88.0005
R5620 VSS.n1001 VSS.n1000 88.0005
R5621 VSS.n987 VSS.n986 88.0005
R5622 VSS.n148 VSS.n147 88.0005
R5623 VSS.n970 VSS.n969 88.0005
R5624 VSS.n956 VSS.n955 88.0005
R5625 VSS.n156 VSS.n155 88.0005
R5626 VSS.n170 VSS.n169 88.0005
R5627 VSS.n937 VSS.n177 88.0005
R5628 VSS.n935 VSS.n934 88.0005
R5629 VSS.n922 VSS.n921 88.0005
R5630 VSS.n192 VSS.n191 88.0005
R5631 VSS.n905 VSS.n904 88.0005
R5632 VSS.n891 VSS.n890 88.0005
R5633 VSS.n877 VSS.n876 88.0005
R5634 VSS.n861 VSS.n860 88.0005
R5635 VSS.n848 VSS.n847 88.0005
R5636 VSS.n834 VSS.n833 88.0005
R5637 VSS.n820 VSS.n819 88.0005
R5638 VSS.n805 VSS.n804 88.0005
R5639 VSS.n791 VSS.n790 88.0005
R5640 VSS.n778 VSS.n777 88.0005
R5641 VSS.n764 VSS.n763 88.0005
R5642 VSS.n750 VSS.n749 88.0005
R5643 VSS.n736 VSS.n735 88.0005
R5644 VSS.n720 VSS.n719 88.0005
R5645 VSS.n706 VSS.n705 88.0005
R5646 VSS.n692 VSS.n691 88.0005
R5647 VSS.n678 VSS.n677 88.0005
R5648 VSS.n202 VSS.n201 88.0005
R5649 VSS.n661 VSS.n660 88.0005
R5650 VSS.n647 VSS.n646 88.0005
R5651 VSS.n210 VSS.n209 88.0005
R5652 VSS.n224 VSS.n223 88.0005
R5653 VSS.n628 VSS.n231 88.0005
R5654 VSS.n626 VSS.n625 88.0005
R5655 VSS.n613 VSS.n612 88.0005
R5656 VSS.n246 VSS.n245 88.0005
R5657 VSS.n596 VSS.n595 88.0005
R5658 VSS.n582 VSS.n581 88.0005
R5659 VSS.n568 VSS.n567 88.0005
R5660 VSS.n552 VSS.n551 88.0005
R5661 VSS.n539 VSS.n538 88.0005
R5662 VSS.n525 VSS.n524 88.0005
R5663 VSS.n511 VSS.n510 88.0005
R5664 VSS.n496 VSS.n495 88.0005
R5665 VSS.n482 VSS.n481 88.0005
R5666 VSS.n469 VSS.n468 88.0005
R5667 VSS.n455 VSS.n454 88.0005
R5668 VSS.n441 VSS.n440 88.0005
R5669 VSS.n427 VSS.n426 88.0005
R5670 VSS.n411 VSS.n410 88.0005
R5671 VSS.n397 VSS.n396 88.0005
R5672 VSS.n383 VSS.n382 88.0005
R5673 VSS.n369 VSS.n368 88.0005
R5674 VSS.n256 VSS.n255 88.0005
R5675 VSS.n352 VSS.n351 88.0005
R5676 VSS.n338 VSS.n337 88.0005
R5677 VSS.n264 VSS.n263 88.0005
R5678 VSS.n278 VSS.n277 88.0005
R5679 VSS.n319 VSS.n318 88.0005
R5680 VSS.n305 VSS.n304 88.0005
R5681 VSS.n291 VSS.n290 88.0005
R5682 VSS.n2117 VSS.n2116 85.7705
R5683 VSS.n2175 VSS.n2174 85.7705
R5684 VSS.n2189 VSS.n2188 85.7705
R5685 VSS.n2203 VSS.n2202 85.7705
R5686 VSS.n2217 VSS.n2216 85.7705
R5687 VSS.n2231 VSS.n2230 85.7705
R5688 VSS.n2231 VSS.t508 85.7705
R5689 VSS.n2245 VSS.n2244 85.7705
R5690 VSS.n2261 VSS.n2260 85.7705
R5691 VSS.n2275 VSS.n2274 85.7705
R5692 VSS.n2289 VSS.n2288 85.7705
R5693 VSS.n2303 VSS.n2302 85.7705
R5694 VSS.n2313 VSS.n2312 85.7705
R5695 VSS.n2329 VSS.n2328 85.7705
R5696 VSS.n2340 VSS.n2339 85.7705
R5697 VSS.n2355 VSS.n107 85.7705
R5698 VSS.n2358 VSS.n2357 85.7705
R5699 VSS.n2371 VSS.n2370 85.7705
R5700 VSS.n2385 VSS.n2384 85.7705
R5701 VSS.n2399 VSS.n2398 85.7705
R5702 VSS.n2410 VSS.n2409 85.7705
R5703 VSS.n2426 VSS.n2425 85.7705
R5704 VSS.n2440 VSS.n2439 85.7705
R5705 VSS.n2454 VSS.n2453 85.7705
R5706 VSS.n2468 VSS.n2467 85.7705
R5707 VSS.n2526 VSS.n2525 85.7705
R5708 VSS.n2540 VSS.n2539 85.7705
R5709 VSS.n2554 VSS.n2553 85.7705
R5710 VSS.n2568 VSS.n2567 85.7705
R5711 VSS.n2582 VSS.n2581 85.7705
R5712 VSS.n2582 VSS.t295 85.7705
R5713 VSS.n2596 VSS.n2595 85.7705
R5714 VSS.n2612 VSS.n2611 85.7705
R5715 VSS.n2626 VSS.n2625 85.7705
R5716 VSS.n2640 VSS.n2639 85.7705
R5717 VSS.n2654 VSS.n2653 85.7705
R5718 VSS.n2664 VSS.n2663 85.7705
R5719 VSS.n2680 VSS.n2679 85.7705
R5720 VSS.n2691 VSS.n2690 85.7705
R5721 VSS.n2706 VSS.n95 85.7705
R5722 VSS.n2709 VSS.n2708 85.7705
R5723 VSS.n2722 VSS.n2721 85.7705
R5724 VSS.n2736 VSS.n2735 85.7705
R5725 VSS.n2750 VSS.n2749 85.7705
R5726 VSS.n2761 VSS.n2760 85.7705
R5727 VSS.n2777 VSS.n2776 85.7705
R5728 VSS.n2791 VSS.n2790 85.7705
R5729 VSS.n2805 VSS.n2804 85.7705
R5730 VSS.n2819 VSS.n2818 85.7705
R5731 VSS.n2877 VSS.n2876 85.7705
R5732 VSS.n2891 VSS.n2890 85.7705
R5733 VSS.n2905 VSS.n2904 85.7705
R5734 VSS.n2919 VSS.n2918 85.7705
R5735 VSS.n2933 VSS.n2932 85.7705
R5736 VSS.n2933 VSS.t117 85.7705
R5737 VSS.n2947 VSS.n2946 85.7705
R5738 VSS.n2963 VSS.n2962 85.7705
R5739 VSS.n2977 VSS.n2976 85.7705
R5740 VSS.n2991 VSS.n2990 85.7705
R5741 VSS.n3005 VSS.n3004 85.7705
R5742 VSS.n3015 VSS.n3014 85.7705
R5743 VSS.n3031 VSS.n3030 85.7705
R5744 VSS.n3042 VSS.n3041 85.7705
R5745 VSS.n3061 VSS.n3060 85.7705
R5746 VSS.n2042 VSS.n2038 83.8127
R5747 VSS.n3225 VSS.t469 82.839
R5748 VSS VSS.n3345 82.839
R5749 VSS.n4116 VSS.n10 81.1181
R5750 VSS.n4111 VSS.n4107 81.1181
R5751 VSS.n4092 VSS.n4088 81.1181
R5752 VSS.n4078 VSS.n4075 81.1181
R5753 VSS.n23 VSS.n19 81.1181
R5754 VSS.n4062 VSS.n4058 81.1181
R5755 VSS.n4050 VSS.n4046 81.1181
R5756 VSS.n4036 VSS.n4032 81.1181
R5757 VSS.n4022 VSS.n4018 81.1181
R5758 VSS.n35 VSS.n31 81.1181
R5759 VSS.n4005 VSS.n4001 81.1181
R5760 VSS.n3993 VSS.n3989 81.1181
R5761 VSS.n3979 VSS.n3975 81.1181
R5762 VSS.n3965 VSS.n3961 81.1181
R5763 VSS.n3950 VSS.n3946 81.1181
R5764 VSS.n3936 VSS.n3932 81.1181
R5765 VSS.n3921 VSS.n3917 81.1181
R5766 VSS.n3907 VSS.n3903 81.1181
R5767 VSS.n49 VSS.n45 81.1181
R5768 VSS.n3193 VSS.t463 79.6529
R5769 VSS.n1212 VSS.t217 79.2005
R5770 VSS.n1204 VSS.t0 79.2005
R5771 VSS.n1111 VSS.t241 79.2005
R5772 VSS.n1103 VSS.t116 79.2005
R5773 VSS.n834 VSS.t365 79.2005
R5774 VSS.n525 VSS.t601 79.2005
R5775 VSS.n1769 VSS.t437 79.0424
R5776 VSS.n1668 VSS.t12 79.0424
R5777 VSS.n1567 VSS.t330 79.0424
R5778 VSS.n1466 VSS.t404 79.0424
R5779 VSS.n1365 VSS.t673 79.0424
R5780 VSS.n4035 VSS.t147 77.1935
R5781 VSS.n1929 VSS.t619 77.1935
R5782 VSS.n1949 VSS.t317 77.1935
R5783 VSS.n2147 VSS.t38 77.1935
R5784 VSS.n2498 VSS.t139 77.1935
R5785 VSS.n2849 VSS.t321 77.1935
R5786 VSS.n3351 VSS.t362 76.4668
R5787 VSS.n2955 VSS.t639 75.7148
R5788 VSS.n2604 VSS.t507 75.7148
R5789 VSS.n2253 VSS.t525 75.7148
R5790 VSS.n1953 VSS.t196 75.7148
R5791 VSS.n1216 VSS.t345 75.7148
R5792 VSS.n1115 VSS.t176 75.7148
R5793 VSS.n864 VSS.t547 75.7148
R5794 VSS.n555 VSS.t395 75.7148
R5795 VSS.n1798 VSS.t335 75.7148
R5796 VSS.n1697 VSS.t154 75.7148
R5797 VSS.n1596 VSS.t649 75.7148
R5798 VSS.n1495 VSS.t9 75.7148
R5799 VSS.n1394 VSS.t669 75.7148
R5800 VSS.n4200 VSS.t160 75.7148
R5801 VSS.n3460 VSS.t399 75.7148
R5802 VSS.n3574 VSS.t527 75.7148
R5803 VSS.n3688 VSS.t62 75.7148
R5804 VSS.n3802 VSS.t517 75.7148
R5805 VSS.n1087 VSS.t348 70.4005
R5806 VSS.n778 VSS.t544 70.4005
R5807 VSS.n469 VSS.t138 70.4005
R5808 VSS.n3076 VSS.t483 70.0946
R5809 VSS.n120 VSS 68.6165
R5810 VSS.n2082 VSS.t262 68.6165
R5811 VSS VSS.n2355 68.6165
R5812 VSS.n2424 VSS.t443 68.6165
R5813 VSS VSS.n2706 68.6165
R5814 VSS.n2775 VSS.t296 68.6165
R5815 VSS VSS.n3061 68.6165
R5816 VSS.n4179 VSS.t161 67.0737
R5817 VSS.n3439 VSS.t400 67.0737
R5818 VSS.n3553 VSS.t528 67.0737
R5819 VSS.n3667 VSS.t63 67.0737
R5820 VSS.n3781 VSS.t514 67.0737
R5821 VSS.n57 VSS.t281 66.9085
R5822 VSS.n3924 VSS.n3923 65.3332
R5823 VSS.n1761 VSS.t260 63.234
R5824 VSS.n1660 VSS.t157 63.234
R5825 VSS.n1559 VSS.t602 63.234
R5826 VSS.n1458 VSS.t520 63.234
R5827 VSS.n1357 VSS.t540 63.234
R5828 VSS.n3952 VSS.t136 62.3526
R5829 VSS.n1086 VSS.n1085 61.6005
R5830 VSS.n1072 VSS.n1071 61.6005
R5831 VSS.n1058 VSS.n1057 61.6005
R5832 VSS.n1044 VSS.n1043 61.6005
R5833 VSS.n1028 VSS.n1027 61.6005
R5834 VSS.n1014 VSS.n1013 61.6005
R5835 VSS.n1000 VSS.n999 61.6005
R5836 VSS.n986 VSS.n985 61.6005
R5837 VSS.n147 VSS.n146 61.6005
R5838 VSS.n969 VSS.n968 61.6005
R5839 VSS.n955 VSS.n954 61.6005
R5840 VSS.n155 VSS.n154 61.6005
R5841 VSS.n169 VSS.n168 61.6005
R5842 VSS.n177 VSS.n176 61.6005
R5843 VSS.n936 VSS.n935 61.6005
R5844 VSS.n921 VSS.n920 61.6005
R5845 VSS.n191 VSS.n190 61.6005
R5846 VSS.n904 VSS.n903 61.6005
R5847 VSS.n890 VSS.n889 61.6005
R5848 VSS.n876 VSS.n875 61.6005
R5849 VSS.n860 VSS.t546 61.6005
R5850 VSS.n847 VSS.n846 61.6005
R5851 VSS.n833 VSS.n832 61.6005
R5852 VSS.n819 VSS.n818 61.6005
R5853 VSS.n804 VSS.n803 61.6005
R5854 VSS.n790 VSS.n789 61.6005
R5855 VSS.n777 VSS.n776 61.6005
R5856 VSS.n763 VSS.n762 61.6005
R5857 VSS.n749 VSS.n748 61.6005
R5858 VSS.n735 VSS.n734 61.6005
R5859 VSS.n719 VSS.n718 61.6005
R5860 VSS.n705 VSS.n704 61.6005
R5861 VSS.n691 VSS.n690 61.6005
R5862 VSS.n677 VSS.n676 61.6005
R5863 VSS.n201 VSS.n200 61.6005
R5864 VSS.n660 VSS.n659 61.6005
R5865 VSS.n646 VSS.n645 61.6005
R5866 VSS.n209 VSS.n208 61.6005
R5867 VSS.n223 VSS.n222 61.6005
R5868 VSS.n231 VSS.n230 61.6005
R5869 VSS.n627 VSS.n626 61.6005
R5870 VSS.n612 VSS.n611 61.6005
R5871 VSS.n245 VSS.n244 61.6005
R5872 VSS.n595 VSS.n594 61.6005
R5873 VSS.n581 VSS.n580 61.6005
R5874 VSS.n567 VSS.n566 61.6005
R5875 VSS.n551 VSS.t394 61.6005
R5876 VSS.n538 VSS.n537 61.6005
R5877 VSS.n524 VSS.n523 61.6005
R5878 VSS.n510 VSS.n509 61.6005
R5879 VSS.n495 VSS.n494 61.6005
R5880 VSS.n481 VSS.n480 61.6005
R5881 VSS.n468 VSS.n467 61.6005
R5882 VSS.n454 VSS.n453 61.6005
R5883 VSS.n440 VSS.n439 61.6005
R5884 VSS.n426 VSS.n425 61.6005
R5885 VSS.n410 VSS.n409 61.6005
R5886 VSS.n396 VSS.n395 61.6005
R5887 VSS.n382 VSS.n381 61.6005
R5888 VSS.n368 VSS.n367 61.6005
R5889 VSS.n255 VSS.n254 61.6005
R5890 VSS.n351 VSS.n350 61.6005
R5891 VSS.n337 VSS.n336 61.6005
R5892 VSS.n263 VSS.n262 61.6005
R5893 VSS.n277 VSS.n276 61.6005
R5894 VSS.n318 VSS.n317 61.6005
R5895 VSS.n304 VSS.n303 61.6005
R5896 VSS.n290 VSS.n289 61.6005
R5897 VSS.n2116 VSS.n2115 60.0395
R5898 VSS.n2130 VSS.n2129 60.0395
R5899 VSS.t571 VSS.n2130 60.0395
R5900 VSS.n2146 VSS.n2145 60.0395
R5901 VSS.n2160 VSS.n2159 60.0395
R5902 VSS.n2174 VSS.n2173 60.0395
R5903 VSS.n2188 VSS.n2187 60.0395
R5904 VSS.n2202 VSS.n2201 60.0395
R5905 VSS.n2216 VSS.n2215 60.0395
R5906 VSS.n2230 VSS.n2229 60.0395
R5907 VSS.n2244 VSS.n2243 60.0395
R5908 VSS.n2260 VSS.n2259 60.0395
R5909 VSS.n2274 VSS.n2273 60.0395
R5910 VSS.n2288 VSS.n2287 60.0395
R5911 VSS.n2302 VSS.n2301 60.0395
R5912 VSS.n2312 VSS.n2311 60.0395
R5913 VSS.n2328 VSS.n2327 60.0395
R5914 VSS.n2339 VSS.n2338 60.0395
R5915 VSS.n107 VSS.n106 60.0395
R5916 VSS.n2357 VSS.n2356 60.0395
R5917 VSS.n2370 VSS.n2369 60.0395
R5918 VSS.n2384 VSS.n2383 60.0395
R5919 VSS.n2398 VSS.n2397 60.0395
R5920 VSS.n2409 VSS.n2408 60.0395
R5921 VSS.n2425 VSS.n2424 60.0395
R5922 VSS.n2439 VSS.n2438 60.0395
R5923 VSS.n2453 VSS.n2452 60.0395
R5924 VSS.n2467 VSS.n2466 60.0395
R5925 VSS.n2481 VSS.n2480 60.0395
R5926 VSS.t82 VSS.n2481 60.0395
R5927 VSS.n2497 VSS.n2496 60.0395
R5928 VSS.n2511 VSS.n2510 60.0395
R5929 VSS.n2525 VSS.n2524 60.0395
R5930 VSS.n2539 VSS.n2538 60.0395
R5931 VSS.n2553 VSS.n2552 60.0395
R5932 VSS.n2567 VSS.n2566 60.0395
R5933 VSS.n2581 VSS.n2580 60.0395
R5934 VSS.n2595 VSS.n2594 60.0395
R5935 VSS.n2611 VSS.n2610 60.0395
R5936 VSS.n2625 VSS.n2624 60.0395
R5937 VSS.n2639 VSS.n2638 60.0395
R5938 VSS.n2653 VSS.n2652 60.0395
R5939 VSS.n2663 VSS.n2662 60.0395
R5940 VSS.n2679 VSS.n2678 60.0395
R5941 VSS.n2690 VSS.n2689 60.0395
R5942 VSS.n95 VSS.n94 60.0395
R5943 VSS.n2708 VSS.n2707 60.0395
R5944 VSS.n2721 VSS.n2720 60.0395
R5945 VSS.n2735 VSS.n2734 60.0395
R5946 VSS.n2749 VSS.n2748 60.0395
R5947 VSS.n2760 VSS.n2759 60.0395
R5948 VSS.n2776 VSS.n2775 60.0395
R5949 VSS.n2790 VSS.n2789 60.0395
R5950 VSS.n2804 VSS.n2803 60.0395
R5951 VSS.n2818 VSS.n2817 60.0395
R5952 VSS.n2832 VSS.n2831 60.0395
R5953 VSS.t2 VSS.n2832 60.0395
R5954 VSS.n2848 VSS.n2847 60.0395
R5955 VSS.n2862 VSS.n2861 60.0395
R5956 VSS.n2876 VSS.n2875 60.0395
R5957 VSS.n2890 VSS.n2889 60.0395
R5958 VSS.n2904 VSS.n2903 60.0395
R5959 VSS.n2918 VSS.n2917 60.0395
R5960 VSS.n2932 VSS.n2931 60.0395
R5961 VSS.n2946 VSS.n2945 60.0395
R5962 VSS.n2962 VSS.n2961 60.0395
R5963 VSS.n2976 VSS.n2975 60.0395
R5964 VSS.n2990 VSS.n2989 60.0395
R5965 VSS.n3004 VSS.n3003 60.0395
R5966 VSS.n3014 VSS.n3013 60.0395
R5967 VSS.n3030 VSS.n3029 60.0395
R5968 VSS.n3041 VSS.n3040 60.0395
R5969 VSS.n3060 VSS.n3059 60.0395
R5970 VSS.n2118 VSS.n2114 57.9417
R5971 VSS.n2132 VSS.n2128 57.9417
R5972 VSS.n2148 VSS.n2144 57.9417
R5973 VSS.n2162 VSS.n2158 57.9417
R5974 VSS.n2176 VSS.n2172 57.9417
R5975 VSS.n2190 VSS.n2186 57.9417
R5976 VSS.n2204 VSS.n2200 57.9417
R5977 VSS.n2218 VSS.n2214 57.9417
R5978 VSS.n2232 VSS.n2228 57.9417
R5979 VSS.n2246 VSS.n2242 57.9417
R5980 VSS.n2262 VSS.n2258 57.9417
R5981 VSS.n2276 VSS.n2272 57.9417
R5982 VSS.n2290 VSS.n2286 57.9417
R5983 VSS.n2304 VSS.n2300 57.9417
R5984 VSS.n2330 VSS.n2326 57.9417
R5985 VSS.n2354 VSS.n109 57.9417
R5986 VSS.n2359 VSS.n105 57.9417
R5987 VSS.n2372 VSS.n2368 57.9417
R5988 VSS.n2386 VSS.n2382 57.9417
R5989 VSS.n2400 VSS.n2396 57.9417
R5990 VSS.n2427 VSS.n2423 57.9417
R5991 VSS.n2441 VSS.n2437 57.9417
R5992 VSS.n2455 VSS.n2451 57.9417
R5993 VSS.n2469 VSS.n2465 57.9417
R5994 VSS.n2483 VSS.n2479 57.9417
R5995 VSS.n2499 VSS.n2495 57.9417
R5996 VSS.n2513 VSS.n2509 57.9417
R5997 VSS.n2527 VSS.n2523 57.9417
R5998 VSS.n2541 VSS.n2537 57.9417
R5999 VSS.n2555 VSS.n2551 57.9417
R6000 VSS.n2569 VSS.n2565 57.9417
R6001 VSS.n2583 VSS.n2579 57.9417
R6002 VSS.n2597 VSS.n2593 57.9417
R6003 VSS.n2613 VSS.n2609 57.9417
R6004 VSS.n2627 VSS.n2623 57.9417
R6005 VSS.n2641 VSS.n2637 57.9417
R6006 VSS.n2655 VSS.n2651 57.9417
R6007 VSS.n2681 VSS.n2677 57.9417
R6008 VSS.n2705 VSS.n97 57.9417
R6009 VSS.n2710 VSS.n93 57.9417
R6010 VSS.n2723 VSS.n2719 57.9417
R6011 VSS.n2737 VSS.n2733 57.9417
R6012 VSS.n2751 VSS.n2747 57.9417
R6013 VSS.n2778 VSS.n2774 57.9417
R6014 VSS.n2792 VSS.n2788 57.9417
R6015 VSS.n2806 VSS.n2802 57.9417
R6016 VSS.n2820 VSS.n2816 57.9417
R6017 VSS.n2834 VSS.n2830 57.9417
R6018 VSS.n2850 VSS.n2846 57.9417
R6019 VSS.n2864 VSS.n2860 57.9417
R6020 VSS.n2878 VSS.n2874 57.9417
R6021 VSS.n2892 VSS.n2888 57.9417
R6022 VSS.n2906 VSS.n2902 57.9417
R6023 VSS.n2920 VSS.n2916 57.9417
R6024 VSS.n2934 VSS.n2930 57.9417
R6025 VSS.n2948 VSS.n2944 57.9417
R6026 VSS.n2964 VSS.n2960 57.9417
R6027 VSS.n2978 VSS.n2974 57.9417
R6028 VSS.n2992 VSS.n2988 57.9417
R6029 VSS.n3006 VSS.n3002 57.9417
R6030 VSS.n3032 VSS.n3028 57.9417
R6031 VSS.n3058 VSS.n73 57.9417
R6032 VSS.n1088 VSS.n1084 57.9417
R6033 VSS.n1074 VSS.n1070 57.9417
R6034 VSS.n1060 VSS.n1056 57.9417
R6035 VSS.n1046 VSS.n1042 57.9417
R6036 VSS.n1030 VSS.n1026 57.9417
R6037 VSS.n1016 VSS.n1012 57.9417
R6038 VSS.n1002 VSS.n998 57.9417
R6039 VSS.n988 VSS.n984 57.9417
R6040 VSS.n149 VSS.n145 57.9417
R6041 VSS.n971 VSS.n967 57.9417
R6042 VSS.n957 VSS.n953 57.9417
R6043 VSS.n171 VSS.n167 57.9417
R6044 VSS.n938 VSS.n175 57.9417
R6045 VSS.n933 VSS.n180 57.9417
R6046 VSS.n923 VSS.n919 57.9417
R6047 VSS.n193 VSS.n189 57.9417
R6048 VSS.n906 VSS.n902 57.9417
R6049 VSS.n892 VSS.n888 57.9417
R6050 VSS.n878 VSS.n874 57.9417
R6051 VSS.n862 VSS.n859 57.9417
R6052 VSS.n849 VSS.n845 57.9417
R6053 VSS.n835 VSS.n831 57.9417
R6054 VSS.n821 VSS.n817 57.9417
R6055 VSS.n806 VSS.n802 57.9417
R6056 VSS.n792 VSS.n788 57.9417
R6057 VSS.n779 VSS.n775 57.9417
R6058 VSS.n765 VSS.n761 57.9417
R6059 VSS.n751 VSS.n747 57.9417
R6060 VSS.n737 VSS.n733 57.9417
R6061 VSS.n721 VSS.n717 57.9417
R6062 VSS.n707 VSS.n703 57.9417
R6063 VSS.n693 VSS.n689 57.9417
R6064 VSS.n679 VSS.n675 57.9417
R6065 VSS.n203 VSS.n199 57.9417
R6066 VSS.n662 VSS.n658 57.9417
R6067 VSS.n648 VSS.n644 57.9417
R6068 VSS.n225 VSS.n221 57.9417
R6069 VSS.n629 VSS.n229 57.9417
R6070 VSS.n624 VSS.n234 57.9417
R6071 VSS.n614 VSS.n610 57.9417
R6072 VSS.n247 VSS.n243 57.9417
R6073 VSS.n597 VSS.n593 57.9417
R6074 VSS.n583 VSS.n579 57.9417
R6075 VSS.n569 VSS.n565 57.9417
R6076 VSS.n553 VSS.n550 57.9417
R6077 VSS.n540 VSS.n536 57.9417
R6078 VSS.n526 VSS.n522 57.9417
R6079 VSS.n512 VSS.n508 57.9417
R6080 VSS.n497 VSS.n493 57.9417
R6081 VSS.n483 VSS.n479 57.9417
R6082 VSS.n470 VSS.n466 57.9417
R6083 VSS.n456 VSS.n452 57.9417
R6084 VSS.n442 VSS.n438 57.9417
R6085 VSS.n428 VSS.n424 57.9417
R6086 VSS.n412 VSS.n408 57.9417
R6087 VSS.n398 VSS.n394 57.9417
R6088 VSS.n384 VSS.n380 57.9417
R6089 VSS.n370 VSS.n366 57.9417
R6090 VSS.n257 VSS.n253 57.9417
R6091 VSS.n353 VSS.n349 57.9417
R6092 VSS.n339 VSS.n335 57.9417
R6093 VSS.n279 VSS.n275 57.9417
R6094 VSS.n320 VSS.n316 57.9417
R6095 VSS.n306 VSS.n302 57.9417
R6096 VSS.n292 VSS.n288 57.9417
R6097 VSS.n3077 VSS.n69 57.9417
R6098 VSS.n3091 VSS.n3087 57.9417
R6099 VSS.n3107 VSS.n3103 57.9417
R6100 VSS.n3121 VSS.n3117 57.9417
R6101 VSS.n3136 VSS.n3133 57.9417
R6102 VSS.n3150 VSS.n3146 57.9417
R6103 VSS.n3166 VSS.n3162 57.9417
R6104 VSS.n3181 VSS.n3177 57.9417
R6105 VSS.n3196 VSS.n3192 57.9417
R6106 VSS.n3212 VSS.n3208 57.9417
R6107 VSS.n3226 VSS.n3222 57.9417
R6108 VSS.n3242 VSS.n3238 57.9417
R6109 VSS.n3256 VSS.n3252 57.9417
R6110 VSS.n3272 VSS.n3268 57.9417
R6111 VSS.n3286 VSS.n3282 57.9417
R6112 VSS.n3302 VSS.n3298 57.9417
R6113 VSS.n3316 VSS.n3312 57.9417
R6114 VSS.n3332 VSS.n3328 57.9417
R6115 VSS.n3344 VSS.n60 57.9417
R6116 VSS.n3241 VSS.t459 57.3502
R6117 VSS.n15 VSS.t60 57.1434
R6118 VSS.n2758 VSS.t297 54.2862
R6119 VSS.n2725 VSS.t324 54.2862
R6120 VSS.n2407 VSS.t444 54.2862
R6121 VSS.n2374 VSS.t142 54.2862
R6122 VSS.n2077 VSS.t263 54.2862
R6123 VSS.n2046 VSS.t41 54.2862
R6124 VSS.n1854 VSS.t54 54.2862
R6125 VSS.n1840 VSS.t586 54.2862
R6126 VSS.n130 VSS.t502 54.2862
R6127 VSS.n135 VSS.t76 54.2862
R6128 VSS.n142 VSS.t426 54.2862
R6129 VSS.n152 VSS.t183 54.2862
R6130 VSS.n196 VSS.t104 54.2862
R6131 VSS.n206 VSS.t566 54.2862
R6132 VSS.n250 VSS.t106 54.2862
R6133 VSS.n260 VSS.t290 54.2862
R6134 VSS.n15 VSS.t89 54.2862
R6135 VSS.n1258 VSS.t631 54.2862
R6136 VSS.n1263 VSS.t166 54.2862
R6137 VSS.n1273 VSS.t414 54.2862
R6138 VSS.n1278 VSS.t373 54.2862
R6139 VSS.n1288 VSS.t424 54.2862
R6140 VSS.n1293 VSS.t48 54.2862
R6141 VSS.n1303 VSS.t531 54.2862
R6142 VSS.n1308 VSS.t657 54.2862
R6143 VSS.n1318 VSS.t629 54.2862
R6144 VSS.n1323 VSS.t310 54.2862
R6145 VSS.n4142 VSS.t389 54.2862
R6146 VSS.n4 VSS.t95 54.2862
R6147 VSS.n3402 VSS.t304 54.2862
R6148 VSS.n3502 VSS.t341 54.2862
R6149 VSS.n3516 VSS.t446 54.2862
R6150 VSS.n3616 VSS.t635 54.2862
R6151 VSS.n3630 VSS.t56 54.2862
R6152 VSS.n3730 VSS.t202 54.2862
R6153 VSS.n3744 VSS.t232 54.2862
R6154 VSS.n4128 VSS.t615 54.2862
R6155 VSS.n3178 VSS.t475 54.1641
R6156 VSS.n4004 VSS.t132 51.4625
R6157 VSS.n1886 VSS.t312 51.4625
R6158 VSS.n2161 VSS.t255 51.4625
R6159 VSS.n2512 VSS.t598 51.4625
R6160 VSS.n2863 VSS.t203 51.4625
R6161 VSS.n3861 VSS.t385 51.4291
R6162 VSS.n53 VSS.t356 50.9781
R6163 VSS VSS.n3370 50.9781
R6164 VSS VSS.n3384 47.792
R6165 VSS.n1794 VSS.t258 47.4256
R6166 VSS.n1786 VSS.t396 47.4256
R6167 VSS.n1693 VSS.t155 47.4256
R6168 VSS.n1685 VSS.t30 47.4256
R6169 VSS.n1592 VSS.t604 47.4256
R6170 VSS.n1584 VSS.t300 47.4256
R6171 VSS.n1491 VSS.t518 47.4256
R6172 VSS.n1483 VSS.t599 47.4256
R6173 VSS.n1390 VSS.t538 47.4256
R6174 VSS.n1382 VSS.t643 47.4256
R6175 VSS.n160 VSS.n159 47.1979
R6176 VSS.n214 VSS.n213 47.1979
R6177 VSS.n268 VSS.n267 47.1979
R6178 VSS.n3046 VSS.n3045 47.1889
R6179 VSS.n2765 VSS.n2764 47.1889
R6180 VSS.n2695 VSS.n2694 47.1889
R6181 VSS.n2414 VSS.n2413 47.1889
R6182 VSS.n2344 VSS.n2343 47.1889
R6183 VSS.n3019 VSS.n3018 47.1845
R6184 VSS.n2668 VSS.n2667 47.1845
R6185 VSS.n2317 VSS.n2316 47.1845
R6186 VSS.n3090 VSS.t473 44.6059
R6187 VSS.n1195 VSS.t346 44.0005
R6188 VSS.n1094 VSS.t173 44.0005
R6189 VSS.n791 VSS.t548 44.0005
R6190 VSS.n482 VSS.t392 44.0005
R6191 VSS.n1909 VSS.t193 42.8855
R6192 VSS.n2836 VSS.t322 41.4291
R6193 VSS.n2485 VSS.t140 41.4291
R6194 VSS.n2134 VSS.t39 41.4291
R6195 VSS.n1873 VSS.t584 41.4291
R6196 VSS.n1177 VSS.t78 41.4291
R6197 VSS.n1037 VSS.t185 41.4291
R6198 VSS.n728 VSS.t568 41.4291
R6199 VSS.n419 VSS.t292 41.4291
R6200 VSS.n1759 VSS.t168 41.4291
R6201 VSS.n1658 VSS.t375 41.4291
R6202 VSS.n1557 VSS.t50 41.4291
R6203 VSS.n1456 VSS.t659 41.4291
R6204 VSS.n1355 VSS.t306 41.4291
R6205 VSS.n4161 VSS.t613 41.4291
R6206 VSS.n3421 VSS.t93 41.4291
R6207 VSS.n3535 VSS.t339 41.4291
R6208 VSS.n3649 VSS.t633 41.4291
R6209 VSS.n3763 VSS.t200 41.4291
R6210 VSS.n3329 VSS.t275 41.4198
R6211 VSS.n2114 VSS.n2113 40.5593
R6212 VSS.n2128 VSS.n2127 40.5593
R6213 VSS.n2144 VSS.n2143 40.5593
R6214 VSS.n2158 VSS.n2157 40.5593
R6215 VSS.n2172 VSS.n2171 40.5593
R6216 VSS.n2186 VSS.n2185 40.5593
R6217 VSS.n2214 VSS.n2213 40.5593
R6218 VSS.n2228 VSS.n2227 40.5593
R6219 VSS.n2242 VSS.n2241 40.5593
R6220 VSS.n2258 VSS.n2257 40.5593
R6221 VSS.n2272 VSS.n2271 40.5593
R6222 VSS.n2286 VSS.n2285 40.5593
R6223 VSS.n2300 VSS.n2299 40.5593
R6224 VSS.n2316 VSS.n2315 40.5593
R6225 VSS.n2326 VSS.n2325 40.5593
R6226 VSS.n2343 VSS.n2342 40.5593
R6227 VSS.n109 VSS.n108 40.5593
R6228 VSS.n110 VSS.n105 40.5593
R6229 VSS.n2382 VSS.n2381 40.5593
R6230 VSS.n2396 VSS.n2395 40.5593
R6231 VSS.n2413 VSS.n2412 40.5593
R6232 VSS.n2423 VSS.n2422 40.5593
R6233 VSS.n2437 VSS.n2436 40.5593
R6234 VSS.n2451 VSS.n2450 40.5593
R6235 VSS.n2465 VSS.n2464 40.5593
R6236 VSS.n2479 VSS.n2478 40.5593
R6237 VSS.n2495 VSS.n2494 40.5593
R6238 VSS.n2509 VSS.n2508 40.5593
R6239 VSS.n2523 VSS.n2522 40.5593
R6240 VSS.n2537 VSS.n2536 40.5593
R6241 VSS.n2565 VSS.n2564 40.5593
R6242 VSS.n2579 VSS.n2578 40.5593
R6243 VSS.n2593 VSS.n2592 40.5593
R6244 VSS.n2609 VSS.n2608 40.5593
R6245 VSS.n2623 VSS.n2622 40.5593
R6246 VSS.n2637 VSS.n2636 40.5593
R6247 VSS.n2651 VSS.n2650 40.5593
R6248 VSS.n2667 VSS.n2666 40.5593
R6249 VSS.n2677 VSS.n2676 40.5593
R6250 VSS.n2694 VSS.n2693 40.5593
R6251 VSS.n97 VSS.n96 40.5593
R6252 VSS.n98 VSS.n93 40.5593
R6253 VSS.n2733 VSS.n2732 40.5593
R6254 VSS.n2747 VSS.n2746 40.5593
R6255 VSS.n2764 VSS.n2763 40.5593
R6256 VSS.n2774 VSS.n2773 40.5593
R6257 VSS.n2788 VSS.n2787 40.5593
R6258 VSS.n2802 VSS.n2801 40.5593
R6259 VSS.n2816 VSS.n2815 40.5593
R6260 VSS.n2830 VSS.n2829 40.5593
R6261 VSS.n2846 VSS.n2845 40.5593
R6262 VSS.n2860 VSS.n2859 40.5593
R6263 VSS.n2874 VSS.n2873 40.5593
R6264 VSS.n2888 VSS.n2887 40.5593
R6265 VSS.n2916 VSS.n2915 40.5593
R6266 VSS.n2930 VSS.n2929 40.5593
R6267 VSS.n2944 VSS.n2943 40.5593
R6268 VSS.n2960 VSS.n2959 40.5593
R6269 VSS.n2974 VSS.n2973 40.5593
R6270 VSS.n2988 VSS.n2987 40.5593
R6271 VSS.n3002 VSS.n3001 40.5593
R6272 VSS.n3018 VSS.n3017 40.5593
R6273 VSS.n3028 VSS.n3027 40.5593
R6274 VSS.n3045 VSS.n3044 40.5593
R6275 VSS.n73 VSS.n72 40.5593
R6276 VSS.n1084 VSS.n1083 40.5593
R6277 VSS.n1070 VSS.n1069 40.5593
R6278 VSS.n1056 VSS.n1055 40.5593
R6279 VSS.n1042 VSS.n1041 40.5593
R6280 VSS.n1026 VSS.n1025 40.5593
R6281 VSS.n1012 VSS.n1011 40.5593
R6282 VSS.n998 VSS.n997 40.5593
R6283 VSS.n984 VSS.n983 40.5593
R6284 VSS.n967 VSS.n966 40.5593
R6285 VSS.n953 VSS.n952 40.5593
R6286 VSS.n159 VSS.n158 40.5593
R6287 VSS.n167 VSS.n166 40.5593
R6288 VSS.n175 VSS.n174 40.5593
R6289 VSS.n919 VSS.n918 40.5593
R6290 VSS.n902 VSS.n901 40.5593
R6291 VSS.n888 VSS.n887 40.5593
R6292 VSS.n874 VSS.n873 40.5593
R6293 VSS.n859 VSS.n858 40.5593
R6294 VSS.n845 VSS.n844 40.5593
R6295 VSS.n831 VSS.n830 40.5593
R6296 VSS.n817 VSS.n816 40.5593
R6297 VSS.n802 VSS.n801 40.5593
R6298 VSS.n775 VSS.n774 40.5593
R6299 VSS.n761 VSS.n760 40.5593
R6300 VSS.n747 VSS.n746 40.5593
R6301 VSS.n733 VSS.n732 40.5593
R6302 VSS.n717 VSS.n716 40.5593
R6303 VSS.n703 VSS.n702 40.5593
R6304 VSS.n689 VSS.n688 40.5593
R6305 VSS.n675 VSS.n674 40.5593
R6306 VSS.n658 VSS.n657 40.5593
R6307 VSS.n644 VSS.n643 40.5593
R6308 VSS.n213 VSS.n212 40.5593
R6309 VSS.n221 VSS.n220 40.5593
R6310 VSS.n229 VSS.n228 40.5593
R6311 VSS.n610 VSS.n609 40.5593
R6312 VSS.n593 VSS.n592 40.5593
R6313 VSS.n579 VSS.n578 40.5593
R6314 VSS.n565 VSS.n564 40.5593
R6315 VSS.n550 VSS.n549 40.5593
R6316 VSS.n536 VSS.n535 40.5593
R6317 VSS.n522 VSS.n521 40.5593
R6318 VSS.n508 VSS.n507 40.5593
R6319 VSS.n493 VSS.n492 40.5593
R6320 VSS.n466 VSS.n465 40.5593
R6321 VSS.n452 VSS.n451 40.5593
R6322 VSS.n438 VSS.n437 40.5593
R6323 VSS.n424 VSS.n423 40.5593
R6324 VSS.n408 VSS.n407 40.5593
R6325 VSS.n394 VSS.n393 40.5593
R6326 VSS.n380 VSS.n379 40.5593
R6327 VSS.n366 VSS.n365 40.5593
R6328 VSS.n349 VSS.n348 40.5593
R6329 VSS.n335 VSS.n334 40.5593
R6330 VSS.n267 VSS.n266 40.5593
R6331 VSS.n275 VSS.n274 40.5593
R6332 VSS.n316 VSS.n315 40.5593
R6333 VSS.n302 VSS.n301 40.5593
R6334 VSS.n288 VSS.n287 40.5593
R6335 VSS.n69 VSS.n68 40.5593
R6336 VSS.n3087 VSS.n3086 40.5593
R6337 VSS.n3103 VSS.n3102 40.5593
R6338 VSS.n3117 VSS.n3116 40.5593
R6339 VSS.n3133 VSS.n3132 40.5593
R6340 VSS.n3146 VSS.n3145 40.5593
R6341 VSS.n3162 VSS.n3161 40.5593
R6342 VSS.n3177 VSS.n3176 40.5593
R6343 VSS.n3192 VSS.n3191 40.5593
R6344 VSS.n3208 VSS.n3207 40.5593
R6345 VSS.n3222 VSS.n3221 40.5593
R6346 VSS.n3238 VSS.n3237 40.5593
R6347 VSS.n3252 VSS.n3251 40.5593
R6348 VSS.n3268 VSS.n3267 40.5593
R6349 VSS.n3282 VSS.n3281 40.5593
R6350 VSS.n3298 VSS.n3297 40.5593
R6351 VSS.n3312 VSS.n3311 40.5593
R6352 VSS.n3328 VSS.n3327 40.5593
R6353 VSS.n60 VSS.n59 40.5593
R6354 VSS.n3923 VSS.t558 39.6928
R6355 VSS.n3039 VSS.t205 38.5719
R6356 VSS.n3039 VSS.t67 38.5719
R6357 VSS.n2955 VSS.t5 38.5719
R6358 VSS.n2836 VSS.t3 38.5719
R6359 VSS.n2688 VSS.t596 38.5719
R6360 VSS.n2688 VSS.t178 38.5719
R6361 VSS.n2604 VSS.t85 38.5719
R6362 VSS.n2485 VSS.t83 38.5719
R6363 VSS.n2337 VSS.t257 38.5719
R6364 VSS.n2337 VSS.t45 38.5719
R6365 VSS.n2253 VSS.t574 38.5719
R6366 VSS.n2134 VSS.t572 38.5719
R6367 VSS.n2023 VSS.t314 38.5719
R6368 VSS.n2023 VSS.t316 38.5719
R6369 VSS.n1953 VSS.t318 38.5719
R6370 VSS.n1873 VSS.t320 38.5719
R6371 VSS.n1241 VSS.t590 38.5719
R6372 VSS.n1241 VSS.t448 38.5719
R6373 VSS.n1216 VSS.t218 38.5719
R6374 VSS.n1177 VSS.t226 38.5719
R6375 VSS.n1139 VSS.t74 38.5719
R6376 VSS.n1139 VSS.t577 38.5719
R6377 VSS.n1115 VSS.t242 38.5719
R6378 VSS.n1037 VSS.t244 38.5719
R6379 VSS.n182 VSS.t72 38.5719
R6380 VSS.n182 VSS.t112 38.5719
R6381 VSS.n864 VSS.t230 38.5719
R6382 VSS.n728 VSS.t240 38.5719
R6383 VSS.n236 VSS.t416 38.5719
R6384 VSS.n236 VSS.t488 38.5719
R6385 VSS.n555 VSS.t220 38.5719
R6386 VSS.n419 VSS.t228 38.5719
R6387 VSS.n13 VSS.t653 38.5719
R6388 VSS.n13 VSS.t58 38.5719
R6389 VSS.n1822 VSS.t19 38.5719
R6390 VSS.n1822 VSS.t440 38.5719
R6391 VSS.n1798 VSS.t259 38.5719
R6392 VSS.n1759 VSS.t261 38.5719
R6393 VSS.n1721 VSS.t588 38.5719
R6394 VSS.n1721 VSS.t14 38.5719
R6395 VSS.n1697 VSS.t156 38.5719
R6396 VSS.n1658 VSS.t158 38.5719
R6397 VSS.n1620 VSS.t387 38.5719
R6398 VSS.n1620 VSS.t329 38.5719
R6399 VSS.n1596 VSS.t605 38.5719
R6400 VSS.n1557 VSS.t603 38.5719
R6401 VSS.n1519 VSS.t627 38.5719
R6402 VSS.n1519 VSS.t403 38.5719
R6403 VSS.n1495 VSS.t519 38.5719
R6404 VSS.n1456 VSS.t521 38.5719
R6405 VSS.n1418 VSS.t35 38.5719
R6406 VSS.n1418 VSS.t672 38.5719
R6407 VSS.n1394 VSS.t539 38.5719
R6408 VSS.n1355 VSS.t541 38.5719
R6409 VSS.n4161 VSS.t234 38.5719
R6410 VSS.n4200 VSS.t236 38.5719
R6411 VSS.n7 VSS.t267 38.5719
R6412 VSS.n7 VSS.t418 38.5719
R6413 VSS.n3421 VSS.t224 38.5719
R6414 VSS.n3460 VSS.t238 38.5719
R6415 VSS.n3390 VSS.t512 38.5719
R6416 VSS.n3390 VSS.t7 38.5719
R6417 VSS.n3535 VSS.t216 38.5719
R6418 VSS.n3574 VSS.t222 38.5719
R6419 VSS.n3388 VSS.t367 38.5719
R6420 VSS.n3388 VSS.t420 38.5719
R6421 VSS.n3649 VSS.t246 38.5719
R6422 VSS.n3688 VSS.t214 38.5719
R6423 VSS.n3386 VSS.t492 38.5719
R6424 VSS.n3386 VSS.t422 38.5719
R6425 VSS.n3763 VSS.t432 38.5719
R6426 VSS.n3802 VSS.t543 38.5719
R6427 VSS.n3832 VSS.t25 38.5719
R6428 VSS.n3832 VSS.t430 38.5719
R6429 VSS.n875 VSS.t545 35.2005
R6430 VSS.n566 VSS.t137 35.2005
R6431 VSS.n2102 VSS.t535 34.3085
R6432 VSS.t255 VSS.n2160 34.3085
R6433 VSS.n2452 VSS.t270 34.3085
R6434 VSS.t598 VSS.n2511 34.3085
R6435 VSS.n2803 VSS.t532 34.3085
R6436 VSS.t203 VSS.n2862 34.3085
R6437 VSS.n3378 VSS.t645 33.462
R6438 VSS.n3378 VSS.t172 33.462
R6439 VSS.n3847 VSS.t21 33.462
R6440 VSS.n3847 VSS.t617 33.462
R6441 VSS.n3076 VSS.n3075 31.8615
R6442 VSS.n3090 VSS.n3089 31.8615
R6443 VSS.n3106 VSS.n3105 31.8615
R6444 VSS.n3135 VSS.t455 31.8615
R6445 VSS.n3149 VSS.n3148 31.8615
R6446 VSS.n3165 VSS.n3164 31.8615
R6447 VSS.n3180 VSS.n3179 31.8615
R6448 VSS.n3195 VSS.n3194 31.8615
R6449 VSS.n3211 VSS.n3210 31.8615
R6450 VSS.n3225 VSS.n3224 31.8615
R6451 VSS.n3241 VSS.n3240 31.8615
R6452 VSS.n3255 VSS.n3254 31.8615
R6453 VSS.n3255 VSS.t479 31.8615
R6454 VSS.n3271 VSS.n3270 31.8615
R6455 VSS.n3301 VSS.n3300 31.8615
R6456 VSS.n3315 VSS.n3314 31.8615
R6457 VSS.n3331 VSS.n3330 31.8615
R6458 VSS.n3345 VSS.n58 31.8615
R6459 VSS.n3893 VSS.n3890 30.1954
R6460 VSS.n3890 VSS.n3887 30.1954
R6461 VSS.n3887 VSS.n3884 30.1954
R6462 VSS.n3884 VSS.n3881 30.1954
R6463 VSS.n3881 VSS.n3878 30.1954
R6464 VSS.n3878 VSS.n3875 30.1954
R6465 VSS.n3861 VSS.t607 28.7917
R6466 VSS.n3163 VSS.t457 28.6754
R6467 VSS.n4175 VSS.t90 26.8298
R6468 VSS.n3435 VSS.t592 26.8298
R6469 VSS.n3549 VSS.t560 26.8298
R6470 VSS.n3663 VSS.t499 26.8298
R6471 VSS.n3777 VSS.t664 26.8298
R6472 VSS.n1777 VSS.t336 26.3478
R6473 VSS.n1676 VSS.t151 26.3478
R6474 VSS.n1575 VSS.t650 26.3478
R6475 VSS.n1474 VSS.t10 26.3478
R6476 VSS.n1373 VSS.t666 26.3478
R6477 VSS.n2758 VSS.t326 25.9346
R6478 VSS.n2725 VSS.t122 25.9346
R6479 VSS.n2407 VSS.t144 25.9346
R6480 VSS.n2374 VSS.t621 25.9346
R6481 VSS.n2077 VSS.t37 25.9346
R6482 VSS.n2046 VSS.t436 25.9346
R6483 VSS.n1854 VSS.t582 25.9346
R6484 VSS.n1840 VSS.t580 25.9346
R6485 VSS.n130 VSS.t80 25.9346
R6486 VSS.n135 VSS.t27 25.9346
R6487 VSS.n142 VSS.t181 25.9346
R6488 VSS.n152 VSS.t253 25.9346
R6489 VSS.n196 VSS.t570 25.9346
R6490 VSS.n206 VSS.t188 25.9346
R6491 VSS.n250 VSS.t288 25.9346
R6492 VSS.n260 VSS.t119 25.9346
R6493 VSS.n1258 VSS.t164 25.9346
R6494 VSS.n1263 VSS.t250 25.9346
R6495 VSS.n1273 VSS.t377 25.9346
R6496 VSS.n1278 VSS.t537 25.9346
R6497 VSS.n1288 VSS.t52 25.9346
R6498 VSS.n1293 VSS.t355 25.9346
R6499 VSS.n1303 VSS.t661 25.9346
R6500 VSS.n1308 VSS.t129 25.9346
R6501 VSS.n1318 VSS.t308 25.9346
R6502 VSS.n1323 VSS.t564 25.9346
R6503 VSS.n4142 VSS.t611 25.9346
R6504 VSS.n4 VSS.t274 25.9346
R6505 VSS.n3402 VSS.t97 25.9346
R6506 VSS.n3502 VSS.t562 25.9346
R6507 VSS.n3516 VSS.t343 25.9346
R6508 VSS.n3616 VSS.t100 25.9346
R6509 VSS.n3630 VSS.t637 25.9346
R6510 VSS.n3730 VSS.t212 25.9346
R6511 VSS.n3744 VSS.t198 25.9346
R6512 VSS.n4128 VSS.t333 25.9346
R6513 VSS.n188 VSS.n187 25.7776
R6514 VSS.n242 VSS.n241 25.7776
R6515 VSS.n2199 VSS.n2198 25.7735
R6516 VSS.n2550 VSS.n2549 25.7735
R6517 VSS.n2901 VSS.n2900 25.7735
R6518 VSS.n787 VSS.n786 25.7735
R6519 VSS.n478 VSS.n477 25.7735
R6520 VSS.n144 VSS.n143 25.7735
R6521 VSS.n179 VSS.n178 25.7735
R6522 VSS.n198 VSS.n197 25.7735
R6523 VSS.n233 VSS.n232 25.7735
R6524 VSS.n252 VSS.n251 25.7735
R6525 VSS.n2367 VSS.n2366 25.765
R6526 VSS.n2718 VSS.n2717 25.765
R6527 VSS.n4119 VSS.n4118 25.7315
R6528 VSS.n4109 VSS.n4108 25.7315
R6529 VSS.n4090 VSS.n4089 25.7315
R6530 VSS.n4076 VSS.t623 25.7315
R6531 VSS.n21 VSS.n20 25.7315
R6532 VSS.n4060 VSS.n4059 25.7315
R6533 VSS.n4061 VSS.t59 25.7315
R6534 VSS.n4048 VSS.n4047 25.7315
R6535 VSS.n4034 VSS.n4033 25.7315
R6536 VSS.n4020 VSS.n4019 25.7315
R6537 VSS.n33 VSS.n32 25.7315
R6538 VSS.n4003 VSS.n4002 25.7315
R6539 VSS.n3991 VSS.n3990 25.7315
R6540 VSS.n3977 VSS.n3976 25.7315
R6541 VSS.n3963 VSS.n3962 25.7315
R6542 VSS.n3948 VSS.n3947 25.7315
R6543 VSS.n3934 VSS.n3933 25.7315
R6544 VSS.n3919 VSS.n3918 25.7315
R6545 VSS.n3905 VSS.n3904 25.7315
R6546 VSS.n47 VSS.n46 25.7315
R6547 VSS.n2131 VSS.t571 25.7315
R6548 VSS.n2482 VSS.t82 25.7315
R6549 VSS.n2833 VSS.t2 25.7315
R6550 VSS.n3066 VSS.t497 25.7315
R6551 VSS.t481 VSS.n3119 25.4893
R6552 VSS.n3952 VSS.t554 24.9241
R6553 VSS.n64 VSS.t466 24.9236
R6554 VSS.n64 VSS.t484 24.9236
R6555 VSS.n3093 VSS.t474 24.9236
R6556 VSS.n3093 VSS.t468 24.9236
R6557 VSS.n3123 VSS.t482 24.9236
R6558 VSS.n3123 VSS.t456 24.9236
R6559 VSS.n3152 VSS.t478 24.9236
R6560 VSS.n3152 VSS.t458 24.9236
R6561 VSS.n3173 VSS.t476 24.9236
R6562 VSS.n3173 VSS.t464 24.9236
R6563 VSS.n3203 VSS.t472 24.9236
R6564 VSS.n3203 VSS.t462 24.9236
R6565 VSS.n3233 VSS.t470 24.9236
R6566 VSS.n3233 VSS.t460 24.9236
R6567 VSS.n3258 VSS.t480 24.9236
R6568 VSS.n3258 VSS.t280 24.9236
R6569 VSS.n3288 VSS.t286 24.9236
R6570 VSS.n3288 VSS.t278 24.9236
R6571 VSS.n3318 VSS.t284 24.9236
R6572 VSS.n3318 VSS.t276 24.9236
R6573 VSS.n3354 VSS.t363 24.9236
R6574 VSS.n3354 VSS.t359 24.9236
R6575 VSS.n3361 VSS.t361 24.9236
R6576 VSS.n3361 VSS.t351 24.9236
R6577 VSS.n3923 VSS.t556 24.9236
R6578 VSS.n3875 VSS.n3872 24.8083
R6579 VSS.n3089 VSS.n3088 22.3032
R6580 VSS.n3105 VSS.n3104 22.3032
R6581 VSS.n3119 VSS.n3118 22.3032
R6582 VSS.t455 VSS.n3134 22.3032
R6583 VSS.n3148 VSS.n3147 22.3032
R6584 VSS.n3164 VSS.n3163 22.3032
R6585 VSS.n3179 VSS.n3178 22.3032
R6586 VSS.n3194 VSS.n3193 22.3032
R6587 VSS.n3210 VSS.n3209 22.3032
R6588 VSS.n3224 VSS.n3223 22.3032
R6589 VSS.n3240 VSS.n3239 22.3032
R6590 VSS.n3254 VSS.n3253 22.3032
R6591 VSS.n3270 VSS.n3269 22.3032
R6592 VSS.n3284 VSS.n3283 22.3032
R6593 VSS.n3314 VSS.n3313 22.3032
R6594 VSS.n3330 VSS.n3329 22.3032
R6595 VSS.n58 VSS.n57 22.3032
R6596 VSS.n1149 VSS.n1146 20.3039
R6597 VSS.n1731 VSS.n1728 20.3039
R6598 VSS.n1630 VSS.n1627 20.3039
R6599 VSS.n1529 VSS.n1526 20.3039
R6600 VSS.n1428 VSS.n1425 20.3039
R6601 VSS.n3075 VSS.n3074 19.1171
R6602 VSS.n3106 VSS.t467 19.1171
R6603 VSS.n3285 VSS.t285 19.1171
R6604 VSS.n1191 VSS.t269 17.6005
R6605 VSS.n4107 VSS.n4106 17.3829
R6606 VSS.n4088 VSS.n4087 17.3829
R6607 VSS.n4075 VSS.n4074 17.3829
R6608 VSS.n19 VSS.n18 17.3829
R6609 VSS.n4058 VSS.n4057 17.3829
R6610 VSS.n4046 VSS.n4045 17.3829
R6611 VSS.n4032 VSS.n4031 17.3829
R6612 VSS.n4018 VSS.n4017 17.3829
R6613 VSS.n31 VSS.n30 17.3829
R6614 VSS.n4001 VSS.n4000 17.3829
R6615 VSS.n3989 VSS.n3988 17.3829
R6616 VSS.n3975 VSS.n3974 17.3829
R6617 VSS.n3961 VSS.n3960 17.3829
R6618 VSS.n3946 VSS.n3945 17.3829
R6619 VSS.n3932 VSS.n3931 17.3829
R6620 VSS.n3917 VSS.n3916 17.3829
R6621 VSS.n3903 VSS.n3902 17.3829
R6622 VSS.n45 VSS.n44 17.3829
R6623 VSS.n4115 VSS.n12 17.2298
R6624 VSS.n4021 VSS.t46 17.1545
R6625 VSS.n1899 VSS.t33 17.1545
R6626 VSS.n3373 VSS 16.7729
R6627 VSS.n4237 VSS 16.7729
R6628 VSS.n3497 VSS 16.7729
R6629 VSS.n3611 VSS 16.7729
R6630 VSS.n3725 VSS 16.7729
R6631 VSS.n3851 VSS 16.5522
R6632 VSS.n3313 VSS.t283 15.931
R6633 VSS.n3894 VSS.n3893 15.3978
R6634 VSS.n3348 VSS.n52 14.3453
R6635 VSS.n4192 VSS.t28 13.4151
R6636 VSS.n4234 VSS 13.4151
R6637 VSS.n3452 VSS.t81 13.4151
R6638 VSS.n3494 VSS 13.4151
R6639 VSS.n3566 VSS.t513 13.4151
R6640 VSS.n3608 VSS 13.4151
R6641 VSS.n3680 VSS.t251 13.4151
R6642 VSS.n3722 VSS 13.4151
R6643 VSS.n3794 VSS.t123 13.4151
R6644 VSS.n3838 VSS 13.4151
R6645 VSS.n2368 VSS.n2367 13.0096
R6646 VSS.n2719 VSS.n2718 13.0096
R6647 VSS.n145 VSS.n144 13.0005
R6648 VSS.n180 VSS.n179 13.0005
R6649 VSS.n199 VSS.n198 13.0005
R6650 VSS.n234 VSS.n233 13.0005
R6651 VSS.n253 VSS.n252 13.0005
R6652 VSS.n2902 VSS.n2901 13.0005
R6653 VSS.n2551 VSS.n2550 13.0005
R6654 VSS.n2200 VSS.n2199 13.0005
R6655 VSS.n788 VSS.n787 13.0005
R6656 VSS.n479 VSS.n478 13.0005
R6657 VSS.n189 VSS.n188 12.9961
R6658 VSS.n243 VSS.n242 12.9961
R6659 VSS.n942 VSS.n941 12.8005
R6660 VSS.n633 VSS.n632 12.8005
R6661 VSS.n324 VSS.n323 12.8005
R6662 VSS.n282 VSS.n281 12.8005
R6663 VSS.t285 VSS.n3284 12.7449
R6664 VSS.n3300 VSS.t277 12.7449
R6665 VSS.n3064 VSS 12.5798
R6666 VSS.n1728 VSS.n1723 12.5798
R6667 VSS.n1627 VSS.n1622 12.5798
R6668 VSS.n1526 VSS.n1521 12.5798
R6669 VSS.n1425 VSS.n1420 12.5798
R6670 VSS.n1829 VSS.n1824 12.5798
R6671 VSS.n12 VSS.n11 12.0275
R6672 VSS VSS.n101 11.035
R6673 VSS VSS.n113 11.035
R6674 VSS VSS.n115 11.035
R6675 VSS.n85 VSS.n84 10.7116
R6676 VSS.n1773 VSS.t248 10.5394
R6677 VSS.n1672 VSS.t647 10.5394
R6678 VSS.n1571 VSS.t594 10.5394
R6679 VSS.n1470 VSS.t107 10.5394
R6680 VSS.n1369 VSS.t169 10.5394
R6681 VSS.n80 VSS.n79 9.6405
R6682 VSS.t277 VSS.n3299 9.55879
R6683 VSS.n3384 VSS.n51 9.55879
R6684 VSS.n50 VSS.n49 9.3005
R6685 VSS.n49 VSS.n48 9.3005
R6686 VSS.n3908 VSS.n3907 9.3005
R6687 VSS.n3907 VSS.n3906 9.3005
R6688 VSS.n3922 VSS.n3921 9.3005
R6689 VSS.n3921 VSS.n3920 9.3005
R6690 VSS.n3937 VSS.n3936 9.3005
R6691 VSS.n3936 VSS.n3935 9.3005
R6692 VSS.n3951 VSS.n3950 9.3005
R6693 VSS.n3950 VSS.n3949 9.3005
R6694 VSS.n3966 VSS.n3965 9.3005
R6695 VSS.n3965 VSS.n3964 9.3005
R6696 VSS.n3980 VSS.n3979 9.3005
R6697 VSS.n3979 VSS.n3978 9.3005
R6698 VSS.n3994 VSS.n3993 9.3005
R6699 VSS.n3993 VSS.n3992 9.3005
R6700 VSS.n4006 VSS.n4005 9.3005
R6701 VSS.n4005 VSS.n4004 9.3005
R6702 VSS.n36 VSS.n35 9.3005
R6703 VSS.n35 VSS.n34 9.3005
R6704 VSS.n4023 VSS.n4022 9.3005
R6705 VSS.n4022 VSS.n4021 9.3005
R6706 VSS.n4037 VSS.n4036 9.3005
R6707 VSS.n4036 VSS.n4035 9.3005
R6708 VSS.n4051 VSS.n4050 9.3005
R6709 VSS.n4050 VSS.n4049 9.3005
R6710 VSS.n4063 VSS.n4062 9.3005
R6711 VSS.n4062 VSS.n4061 9.3005
R6712 VSS.n26 VSS.n23 9.3005
R6713 VSS.n23 VSS.n22 9.3005
R6714 VSS.n4079 VSS.n4078 9.3005
R6715 VSS.n4078 VSS.n4077 9.3005
R6716 VSS.n4093 VSS.n4092 9.3005
R6717 VSS.n4092 VSS.n4091 9.3005
R6718 VSS.n4112 VSS.n4111 9.3005
R6719 VSS.n4111 VSS.n4110 9.3005
R6720 VSS.n4116 VSS.n4115 9.3005
R6721 VSS.n4117 VSS.n4116 9.3005
R6722 VSS.n3078 VSS.n3077 9.3005
R6723 VSS.n3077 VSS.n3076 9.3005
R6724 VSS.n3092 VSS.n3091 9.3005
R6725 VSS.n3091 VSS.n3090 9.3005
R6726 VSS.n3108 VSS.n3107 9.3005
R6727 VSS.n3107 VSS.n3106 9.3005
R6728 VSS.n3122 VSS.n3121 9.3005
R6729 VSS.n3121 VSS.n3120 9.3005
R6730 VSS.n3137 VSS.n3136 9.3005
R6731 VSS.n3136 VSS.n3135 9.3005
R6732 VSS.n3151 VSS.n3150 9.3005
R6733 VSS.n3150 VSS.n3149 9.3005
R6734 VSS.n3167 VSS.n3166 9.3005
R6735 VSS.n3166 VSS.n3165 9.3005
R6736 VSS.n3182 VSS.n3181 9.3005
R6737 VSS.n3181 VSS.n3180 9.3005
R6738 VSS.n3197 VSS.n3196 9.3005
R6739 VSS.n3196 VSS.n3195 9.3005
R6740 VSS.n3213 VSS.n3212 9.3005
R6741 VSS.n3212 VSS.n3211 9.3005
R6742 VSS.n3227 VSS.n3226 9.3005
R6743 VSS.n3226 VSS.n3225 9.3005
R6744 VSS.n3243 VSS.n3242 9.3005
R6745 VSS.n3242 VSS.n3241 9.3005
R6746 VSS.n3257 VSS.n3256 9.3005
R6747 VSS.n3256 VSS.n3255 9.3005
R6748 VSS.n3273 VSS.n3272 9.3005
R6749 VSS.n3272 VSS.n3271 9.3005
R6750 VSS.n3287 VSS.n3286 9.3005
R6751 VSS.n3286 VSS.n3285 9.3005
R6752 VSS.n3303 VSS.n3302 9.3005
R6753 VSS.n3302 VSS.n3301 9.3005
R6754 VSS.n3317 VSS.n3316 9.3005
R6755 VSS.n3316 VSS.n3315 9.3005
R6756 VSS.n3333 VSS.n3332 9.3005
R6757 VSS.n3332 VSS.n3331 9.3005
R6758 VSS.n3344 VSS.n3343 9.3005
R6759 VSS.n3345 VSS.n3344 9.3005
R6760 VSS.n1891 VSS.n1890 9.3005
R6761 VSS.n1890 VSS.n1889 9.3005
R6762 VSS.n1901 VSS.n1900 9.3005
R6763 VSS.n1900 VSS.n1899 9.3005
R6764 VSS.n1921 VSS.n1920 9.3005
R6765 VSS.n1920 VSS.n1919 9.3005
R6766 VSS.n1931 VSS.n1930 9.3005
R6767 VSS.n1930 VSS.n1929 9.3005
R6768 VSS.n1941 VSS.n1940 9.3005
R6769 VSS.n1940 VSS.n1939 9.3005
R6770 VSS.n1963 VSS.n1962 9.3005
R6771 VSS.n1962 VSS.n1961 9.3005
R6772 VSS.n1973 VSS.n1972 9.3005
R6773 VSS.n1972 VSS.n1971 9.3005
R6774 VSS.n1983 VSS.n1982 9.3005
R6775 VSS.n1982 VSS.n1981 9.3005
R6776 VSS.n1996 VSS.n1995 9.3005
R6777 VSS.n2013 VSS.n2012 9.3005
R6778 VSS.n2012 VSS.n2011 9.3005
R6779 VSS.n2016 VSS.n2015 9.3005
R6780 VSS.n2036 VSS.n2035 9.3005
R6781 VSS.n2035 VSS.n2034 9.3005
R6782 VSS.n2045 VSS.n2044 9.3005
R6783 VSS.n2044 VSS.n2043 9.3005
R6784 VSS.n2057 VSS.n2056 9.3005
R6785 VSS.n2056 VSS.n2055 9.3005
R6786 VSS.n2070 VSS.n2069 9.3005
R6787 VSS.n2088 VSS.n2087 9.3005
R6788 VSS.n2087 VSS.n2086 9.3005
R6789 VSS.n2098 VSS.n2097 9.3005
R6790 VSS.n2097 VSS.n2096 9.3005
R6791 VSS.n2119 VSS.n2118 9.3005
R6792 VSS.n2118 VSS.n2117 9.3005
R6793 VSS.n2133 VSS.n2132 9.3005
R6794 VSS.n2132 VSS.n2131 9.3005
R6795 VSS.n2149 VSS.n2148 9.3005
R6796 VSS.n2148 VSS.n2147 9.3005
R6797 VSS.n2163 VSS.n2162 9.3005
R6798 VSS.n2162 VSS.n2161 9.3005
R6799 VSS.n2177 VSS.n2176 9.3005
R6800 VSS.n2176 VSS.n2175 9.3005
R6801 VSS.n2191 VSS.n2190 9.3005
R6802 VSS.n2190 VSS.n2189 9.3005
R6803 VSS.n2205 VSS.n2204 9.3005
R6804 VSS.n2204 VSS.n2203 9.3005
R6805 VSS.n2219 VSS.n2218 9.3005
R6806 VSS.n2218 VSS.n2217 9.3005
R6807 VSS.n2233 VSS.n2232 9.3005
R6808 VSS.n2232 VSS.n2231 9.3005
R6809 VSS.n2247 VSS.n2246 9.3005
R6810 VSS.n2246 VSS.n2245 9.3005
R6811 VSS.n2263 VSS.n2262 9.3005
R6812 VSS.n2262 VSS.n2261 9.3005
R6813 VSS.n2277 VSS.n2276 9.3005
R6814 VSS.n2276 VSS.n2275 9.3005
R6815 VSS.n2291 VSS.n2290 9.3005
R6816 VSS.n2290 VSS.n2289 9.3005
R6817 VSS.n2305 VSS.n2304 9.3005
R6818 VSS.n2304 VSS.n2303 9.3005
R6819 VSS.n2314 VSS.n2313 9.3005
R6820 VSS.n2331 VSS.n2330 9.3005
R6821 VSS.n2330 VSS.n2329 9.3005
R6822 VSS.n2341 VSS.n2340 9.3005
R6823 VSS.n2354 VSS.n2353 9.3005
R6824 VSS.n2355 VSS.n2354 9.3005
R6825 VSS.n2360 VSS.n2359 9.3005
R6826 VSS.n2359 VSS.n2358 9.3005
R6827 VSS.n2373 VSS.n2372 9.3005
R6828 VSS.n2372 VSS.n2371 9.3005
R6829 VSS.n2387 VSS.n2386 9.3005
R6830 VSS.n2386 VSS.n2385 9.3005
R6831 VSS.n2401 VSS.n2400 9.3005
R6832 VSS.n2400 VSS.n2399 9.3005
R6833 VSS.n2411 VSS.n2410 9.3005
R6834 VSS.n2428 VSS.n2427 9.3005
R6835 VSS.n2427 VSS.n2426 9.3005
R6836 VSS.n2442 VSS.n2441 9.3005
R6837 VSS.n2441 VSS.n2440 9.3005
R6838 VSS.n2456 VSS.n2455 9.3005
R6839 VSS.n2455 VSS.n2454 9.3005
R6840 VSS.n2470 VSS.n2469 9.3005
R6841 VSS.n2469 VSS.n2468 9.3005
R6842 VSS.n2484 VSS.n2483 9.3005
R6843 VSS.n2483 VSS.n2482 9.3005
R6844 VSS.n2500 VSS.n2499 9.3005
R6845 VSS.n2499 VSS.n2498 9.3005
R6846 VSS.n2514 VSS.n2513 9.3005
R6847 VSS.n2513 VSS.n2512 9.3005
R6848 VSS.n2528 VSS.n2527 9.3005
R6849 VSS.n2527 VSS.n2526 9.3005
R6850 VSS.n2542 VSS.n2541 9.3005
R6851 VSS.n2541 VSS.n2540 9.3005
R6852 VSS.n2556 VSS.n2555 9.3005
R6853 VSS.n2555 VSS.n2554 9.3005
R6854 VSS.n2570 VSS.n2569 9.3005
R6855 VSS.n2569 VSS.n2568 9.3005
R6856 VSS.n2584 VSS.n2583 9.3005
R6857 VSS.n2583 VSS.n2582 9.3005
R6858 VSS.n2598 VSS.n2597 9.3005
R6859 VSS.n2597 VSS.n2596 9.3005
R6860 VSS.n2614 VSS.n2613 9.3005
R6861 VSS.n2613 VSS.n2612 9.3005
R6862 VSS.n2628 VSS.n2627 9.3005
R6863 VSS.n2627 VSS.n2626 9.3005
R6864 VSS.n2642 VSS.n2641 9.3005
R6865 VSS.n2641 VSS.n2640 9.3005
R6866 VSS.n2656 VSS.n2655 9.3005
R6867 VSS.n2655 VSS.n2654 9.3005
R6868 VSS.n2665 VSS.n2664 9.3005
R6869 VSS.n2682 VSS.n2681 9.3005
R6870 VSS.n2681 VSS.n2680 9.3005
R6871 VSS.n2692 VSS.n2691 9.3005
R6872 VSS.n2705 VSS.n2704 9.3005
R6873 VSS.n2706 VSS.n2705 9.3005
R6874 VSS.n2711 VSS.n2710 9.3005
R6875 VSS.n2710 VSS.n2709 9.3005
R6876 VSS.n2724 VSS.n2723 9.3005
R6877 VSS.n2723 VSS.n2722 9.3005
R6878 VSS.n2738 VSS.n2737 9.3005
R6879 VSS.n2737 VSS.n2736 9.3005
R6880 VSS.n2752 VSS.n2751 9.3005
R6881 VSS.n2751 VSS.n2750 9.3005
R6882 VSS.n2762 VSS.n2761 9.3005
R6883 VSS.n2779 VSS.n2778 9.3005
R6884 VSS.n2778 VSS.n2777 9.3005
R6885 VSS.n2793 VSS.n2792 9.3005
R6886 VSS.n2792 VSS.n2791 9.3005
R6887 VSS.n2807 VSS.n2806 9.3005
R6888 VSS.n2806 VSS.n2805 9.3005
R6889 VSS.n2821 VSS.n2820 9.3005
R6890 VSS.n2820 VSS.n2819 9.3005
R6891 VSS.n2835 VSS.n2834 9.3005
R6892 VSS.n2834 VSS.n2833 9.3005
R6893 VSS.n2851 VSS.n2850 9.3005
R6894 VSS.n2850 VSS.n2849 9.3005
R6895 VSS.n2865 VSS.n2864 9.3005
R6896 VSS.n2864 VSS.n2863 9.3005
R6897 VSS.n2879 VSS.n2878 9.3005
R6898 VSS.n2878 VSS.n2877 9.3005
R6899 VSS.n2893 VSS.n2892 9.3005
R6900 VSS.n2892 VSS.n2891 9.3005
R6901 VSS.n2907 VSS.n2906 9.3005
R6902 VSS.n2906 VSS.n2905 9.3005
R6903 VSS.n2921 VSS.n2920 9.3005
R6904 VSS.n2920 VSS.n2919 9.3005
R6905 VSS.n2935 VSS.n2934 9.3005
R6906 VSS.n2934 VSS.n2933 9.3005
R6907 VSS.n2949 VSS.n2948 9.3005
R6908 VSS.n2948 VSS.n2947 9.3005
R6909 VSS.n2965 VSS.n2964 9.3005
R6910 VSS.n2964 VSS.n2963 9.3005
R6911 VSS.n2979 VSS.n2978 9.3005
R6912 VSS.n2978 VSS.n2977 9.3005
R6913 VSS.n2993 VSS.n2992 9.3005
R6914 VSS.n2992 VSS.n2991 9.3005
R6915 VSS.n3007 VSS.n3006 9.3005
R6916 VSS.n3006 VSS.n3005 9.3005
R6917 VSS.n3016 VSS.n3015 9.3005
R6918 VSS.n3033 VSS.n3032 9.3005
R6919 VSS.n3032 VSS.n3031 9.3005
R6920 VSS.n3043 VSS.n3042 9.3005
R6921 VSS.n3058 VSS.n3057 9.3005
R6922 VSS.n3061 VSS.n3058 9.3005
R6923 VSS.n2108 VSS.n2107 9.3005
R6924 VSS.n2107 VSS.n2106 9.3005
R6925 VSS.n2067 VSS.n2066 9.3005
R6926 VSS.n2066 VSS.n2065 9.3005
R6927 VSS.n2028 VSS.n2027 9.3005
R6928 VSS.n2029 VSS.n2028 9.3005
R6929 VSS.n1993 VSS.n1992 9.3005
R6930 VSS.n1992 VSS.n1991 9.3005
R6931 VSS.n1951 VSS.n1950 9.3005
R6932 VSS.n1950 VSS.n1949 9.3005
R6933 VSS.n1911 VSS.n1910 9.3005
R6934 VSS.n1910 VSS.n1909 9.3005
R6935 VSS.n1089 VSS.n1088 9.3005
R6936 VSS.n1088 VSS.n1087 9.3005
R6937 VSS.n1075 VSS.n1074 9.3005
R6938 VSS.n1074 VSS.n1073 9.3005
R6939 VSS.n1061 VSS.n1060 9.3005
R6940 VSS.n1060 VSS.n1059 9.3005
R6941 VSS.n1047 VSS.n1046 9.3005
R6942 VSS.n1046 VSS.n1045 9.3005
R6943 VSS.n1031 VSS.n1030 9.3005
R6944 VSS.n1030 VSS.n1029 9.3005
R6945 VSS.n1017 VSS.n1016 9.3005
R6946 VSS.n1016 VSS.n1015 9.3005
R6947 VSS.n1003 VSS.n1002 9.3005
R6948 VSS.n1002 VSS.n1001 9.3005
R6949 VSS.n989 VSS.n988 9.3005
R6950 VSS.n988 VSS.n987 9.3005
R6951 VSS.n150 VSS.n149 9.3005
R6952 VSS.n149 VSS.n148 9.3005
R6953 VSS.n972 VSS.n971 9.3005
R6954 VSS.n971 VSS.n970 9.3005
R6955 VSS.n958 VSS.n957 9.3005
R6956 VSS.n957 VSS.n956 9.3005
R6957 VSS.n157 VSS.n156 9.3005
R6958 VSS.n172 VSS.n171 9.3005
R6959 VSS.n171 VSS.n170 9.3005
R6960 VSS.n939 VSS.n938 9.3005
R6961 VSS.n938 VSS.n937 9.3005
R6962 VSS.n933 VSS.n932 9.3005
R6963 VSS.n934 VSS.n933 9.3005
R6964 VSS.n924 VSS.n923 9.3005
R6965 VSS.n923 VSS.n922 9.3005
R6966 VSS.n194 VSS.n193 9.3005
R6967 VSS.n193 VSS.n192 9.3005
R6968 VSS.n907 VSS.n906 9.3005
R6969 VSS.n906 VSS.n905 9.3005
R6970 VSS.n893 VSS.n892 9.3005
R6971 VSS.n892 VSS.n891 9.3005
R6972 VSS.n879 VSS.n878 9.3005
R6973 VSS.n878 VSS.n877 9.3005
R6974 VSS.n863 VSS.n862 9.3005
R6975 VSS.n862 VSS.n861 9.3005
R6976 VSS.n850 VSS.n849 9.3005
R6977 VSS.n849 VSS.n848 9.3005
R6978 VSS.n836 VSS.n835 9.3005
R6979 VSS.n835 VSS.n834 9.3005
R6980 VSS.n822 VSS.n821 9.3005
R6981 VSS.n821 VSS.n820 9.3005
R6982 VSS.n807 VSS.n806 9.3005
R6983 VSS.n806 VSS.n805 9.3005
R6984 VSS.n793 VSS.n792 9.3005
R6985 VSS.n792 VSS.n791 9.3005
R6986 VSS.n780 VSS.n779 9.3005
R6987 VSS.n779 VSS.n778 9.3005
R6988 VSS.n766 VSS.n765 9.3005
R6989 VSS.n765 VSS.n764 9.3005
R6990 VSS.n752 VSS.n751 9.3005
R6991 VSS.n751 VSS.n750 9.3005
R6992 VSS.n738 VSS.n737 9.3005
R6993 VSS.n737 VSS.n736 9.3005
R6994 VSS.n722 VSS.n721 9.3005
R6995 VSS.n721 VSS.n720 9.3005
R6996 VSS.n708 VSS.n707 9.3005
R6997 VSS.n707 VSS.n706 9.3005
R6998 VSS.n694 VSS.n693 9.3005
R6999 VSS.n693 VSS.n692 9.3005
R7000 VSS.n680 VSS.n679 9.3005
R7001 VSS.n679 VSS.n678 9.3005
R7002 VSS.n204 VSS.n203 9.3005
R7003 VSS.n203 VSS.n202 9.3005
R7004 VSS.n663 VSS.n662 9.3005
R7005 VSS.n662 VSS.n661 9.3005
R7006 VSS.n649 VSS.n648 9.3005
R7007 VSS.n648 VSS.n647 9.3005
R7008 VSS.n211 VSS.n210 9.3005
R7009 VSS.n226 VSS.n225 9.3005
R7010 VSS.n225 VSS.n224 9.3005
R7011 VSS.n630 VSS.n629 9.3005
R7012 VSS.n629 VSS.n628 9.3005
R7013 VSS.n624 VSS.n623 9.3005
R7014 VSS.n625 VSS.n624 9.3005
R7015 VSS.n615 VSS.n614 9.3005
R7016 VSS.n614 VSS.n613 9.3005
R7017 VSS.n248 VSS.n247 9.3005
R7018 VSS.n247 VSS.n246 9.3005
R7019 VSS.n598 VSS.n597 9.3005
R7020 VSS.n597 VSS.n596 9.3005
R7021 VSS.n584 VSS.n583 9.3005
R7022 VSS.n583 VSS.n582 9.3005
R7023 VSS.n570 VSS.n569 9.3005
R7024 VSS.n569 VSS.n568 9.3005
R7025 VSS.n554 VSS.n553 9.3005
R7026 VSS.n553 VSS.n552 9.3005
R7027 VSS.n541 VSS.n540 9.3005
R7028 VSS.n540 VSS.n539 9.3005
R7029 VSS.n527 VSS.n526 9.3005
R7030 VSS.n526 VSS.n525 9.3005
R7031 VSS.n513 VSS.n512 9.3005
R7032 VSS.n512 VSS.n511 9.3005
R7033 VSS.n498 VSS.n497 9.3005
R7034 VSS.n497 VSS.n496 9.3005
R7035 VSS.n484 VSS.n483 9.3005
R7036 VSS.n483 VSS.n482 9.3005
R7037 VSS.n471 VSS.n470 9.3005
R7038 VSS.n470 VSS.n469 9.3005
R7039 VSS.n457 VSS.n456 9.3005
R7040 VSS.n456 VSS.n455 9.3005
R7041 VSS.n443 VSS.n442 9.3005
R7042 VSS.n442 VSS.n441 9.3005
R7043 VSS.n429 VSS.n428 9.3005
R7044 VSS.n428 VSS.n427 9.3005
R7045 VSS.n413 VSS.n412 9.3005
R7046 VSS.n412 VSS.n411 9.3005
R7047 VSS.n399 VSS.n398 9.3005
R7048 VSS.n398 VSS.n397 9.3005
R7049 VSS.n385 VSS.n384 9.3005
R7050 VSS.n384 VSS.n383 9.3005
R7051 VSS.n371 VSS.n370 9.3005
R7052 VSS.n370 VSS.n369 9.3005
R7053 VSS.n258 VSS.n257 9.3005
R7054 VSS.n257 VSS.n256 9.3005
R7055 VSS.n354 VSS.n353 9.3005
R7056 VSS.n353 VSS.n352 9.3005
R7057 VSS.n340 VSS.n339 9.3005
R7058 VSS.n339 VSS.n338 9.3005
R7059 VSS.n265 VSS.n264 9.3005
R7060 VSS.n280 VSS.n279 9.3005
R7061 VSS.n279 VSS.n278 9.3005
R7062 VSS.n321 VSS.n320 9.3005
R7063 VSS.n320 VSS.n319 9.3005
R7064 VSS.n307 VSS.n306 9.3005
R7065 VSS.n306 VSS.n305 9.3005
R7066 VSS.n293 VSS.n292 9.3005
R7067 VSS.n292 VSS.n291 9.3005
R7068 VSS.n3071 VSS.n71 9.04877
R7069 VSS.n1220 VSS.n1217 9.04877
R7070 VSS.n1119 VSS.n1116 9.04877
R7071 VSS.n1802 VSS.n1799 9.04877
R7072 VSS.n1701 VSS.n1698 9.04877
R7073 VSS.n1600 VSS.n1597 9.04877
R7074 VSS.n1499 VSS.n1496 9.04877
R7075 VSS.n1398 VSS.n1395 9.04877
R7076 VSS.n4204 VSS.n4201 9.04877
R7077 VSS.n3464 VSS.n3461 9.04877
R7078 VSS.n3578 VSS.n3575 9.04877
R7079 VSS.n3692 VSS.n3689 9.04877
R7080 VSS.n3806 VSS.n3803 9.04877
R7081 VSS.n3 VSS.n2 9.01861
R7082 VSS.n3501 VSS.n3500 9.01861
R7083 VSS.n3615 VSS.n3614 9.01861
R7084 VSS.n3729 VSS.n3728 9.01861
R7085 VSS.n3860 VSS.n3859 9.01832
R7086 VSS.n4127 VSS.n4126 9.01761
R7087 VSS.n3846 VSS.n3845 9.01734
R7088 VSS.n4141 VSS.n4140 9.01732
R7089 VSS.n4230 VSS.n4229 9.01732
R7090 VSS.n3401 VSS.n3400 9.01732
R7091 VSS.n3492 VSS.n3491 9.01732
R7092 VSS.n3515 VSS.n3514 9.01732
R7093 VSS.n3606 VSS.n3605 9.01732
R7094 VSS.n3629 VSS.n3628 9.01732
R7095 VSS.n3720 VSS.n3719 9.01732
R7096 VSS.n3743 VSS.n3742 9.01732
R7097 VSS.n3831 VSS.n3830 9.01732
R7098 VSS.n4220 VSS.n4219 9.01719
R7099 VSS.n3480 VSS.n3479 9.01719
R7100 VSS.n3594 VSS.n3593 9.01719
R7101 VSS.n3708 VSS.n3707 9.01719
R7102 VSS.n3822 VSS.n3821 9.01719
R7103 VSS.n1839 VSS.n1838 9.01662
R7104 VSS.n134 VSS.n133 9.01662
R7105 VSS.n1262 VSS.n1261 9.01662
R7106 VSS.n1277 VSS.n1276 9.01662
R7107 VSS.n1292 VSS.n1291 9.01662
R7108 VSS.n1307 VSS.n1306 9.01662
R7109 VSS.n1322 VSS.n1321 9.01662
R7110 VSS.n1853 VSS.n1852 9.01634
R7111 VSS.n1244 VSS.n1243 9.01634
R7112 VSS.n129 VSS.n128 9.01634
R7113 VSS.n1142 VSS.n1141 9.01634
R7114 VSS.n3353 VSS.n3352 9.01634
R7115 VSS.n3377 VSS.n3376 9.01634
R7116 VSS.n1257 VSS.n1256 9.01634
R7117 VSS.n1724 VSS.n1723 9.01634
R7118 VSS.n1272 VSS.n1271 9.01634
R7119 VSS.n1623 VSS.n1622 9.01634
R7120 VSS.n1287 VSS.n1286 9.01634
R7121 VSS.n1522 VSS.n1521 9.01634
R7122 VSS.n1302 VSS.n1301 9.01634
R7123 VSS.n1421 VSS.n1420 9.01634
R7124 VSS.n1317 VSS.n1316 9.01634
R7125 VSS.n1825 VSS.n1824 9.01634
R7126 VSS.n125 VSS.n124 9.0162
R7127 VSS.n140 VSS.n139 9.0162
R7128 VSS.n1253 VSS.n1252 9.0162
R7129 VSS.n1268 VSS.n1267 9.0162
R7130 VSS.n1283 VSS.n1282 9.0162
R7131 VSS.n1298 VSS.n1297 9.0162
R7132 VSS.n1313 VSS.n1312 9.0162
R7133 VSS.n3845 VSS.n3844 9.01392
R7134 VSS.n3871 VSS.n3870 9.01392
R7135 VSS.n3866 VSS.n3865 9.01392
R7136 VSS.n3856 VSS.n3855 9.01392
R7137 VSS.n3852 VSS.n3851 9.01392
R7138 VSS.n1829 VSS.n1828 9.01392
R7139 VSS.n1828 VSS.n1827 9.01392
R7140 VSS.n1819 VSS.n1818 9.01392
R7141 VSS.n1814 VSS.n1813 9.01392
R7142 VSS.n1810 VSS.n1809 9.01392
R7143 VSS.n1806 VSS.n1805 9.01392
R7144 VSS.n1802 VSS.n1801 9.01392
R7145 VSS.n1796 VSS.n1795 9.01392
R7146 VSS.n1792 VSS.n1791 9.01392
R7147 VSS.n1788 VSS.n1787 9.01392
R7148 VSS.n1784 VSS.n1783 9.01392
R7149 VSS.n1779 VSS.n1778 9.01392
R7150 VSS.n1775 VSS.n1774 9.01392
R7151 VSS.n1771 VSS.n1770 9.01392
R7152 VSS.n1767 VSS.n1766 9.01392
R7153 VSS.n1763 VSS.n1762 9.01392
R7154 VSS.n1757 VSS.n1756 9.01392
R7155 VSS.n1753 VSS.n1752 9.01392
R7156 VSS.n1749 VSS.n1748 9.01392
R7157 VSS.n1745 VSS.n1744 9.01392
R7158 VSS.n1740 VSS.n1739 9.01392
R7159 VSS.n1736 VSS.n1735 9.01392
R7160 VSS.n1731 VSS.n1730 9.01392
R7161 VSS.n1728 VSS.n1727 9.01392
R7162 VSS.n1718 VSS.n1717 9.01392
R7163 VSS.n1713 VSS.n1712 9.01392
R7164 VSS.n1709 VSS.n1708 9.01392
R7165 VSS.n1705 VSS.n1704 9.01392
R7166 VSS.n1701 VSS.n1700 9.01392
R7167 VSS.n1695 VSS.n1694 9.01392
R7168 VSS.n1691 VSS.n1690 9.01392
R7169 VSS.n1687 VSS.n1686 9.01392
R7170 VSS.n1683 VSS.n1682 9.01392
R7171 VSS.n1678 VSS.n1677 9.01392
R7172 VSS.n1674 VSS.n1673 9.01392
R7173 VSS.n1670 VSS.n1669 9.01392
R7174 VSS.n1666 VSS.n1665 9.01392
R7175 VSS.n1662 VSS.n1661 9.01392
R7176 VSS.n1656 VSS.n1655 9.01392
R7177 VSS.n1652 VSS.n1651 9.01392
R7178 VSS.n1648 VSS.n1647 9.01392
R7179 VSS.n1644 VSS.n1643 9.01392
R7180 VSS.n1639 VSS.n1638 9.01392
R7181 VSS.n1635 VSS.n1634 9.01392
R7182 VSS.n1630 VSS.n1629 9.01392
R7183 VSS.n1627 VSS.n1626 9.01392
R7184 VSS.n1617 VSS.n1616 9.01392
R7185 VSS.n1612 VSS.n1611 9.01392
R7186 VSS.n1608 VSS.n1607 9.01392
R7187 VSS.n1604 VSS.n1603 9.01392
R7188 VSS.n1600 VSS.n1599 9.01392
R7189 VSS.n1594 VSS.n1593 9.01392
R7190 VSS.n1590 VSS.n1589 9.01392
R7191 VSS.n1586 VSS.n1585 9.01392
R7192 VSS.n1582 VSS.n1581 9.01392
R7193 VSS.n1577 VSS.n1576 9.01392
R7194 VSS.n1573 VSS.n1572 9.01392
R7195 VSS.n1569 VSS.n1568 9.01392
R7196 VSS.n1565 VSS.n1564 9.01392
R7197 VSS.n1561 VSS.n1560 9.01392
R7198 VSS.n1555 VSS.n1554 9.01392
R7199 VSS.n1551 VSS.n1550 9.01392
R7200 VSS.n1547 VSS.n1546 9.01392
R7201 VSS.n1543 VSS.n1542 9.01392
R7202 VSS.n1538 VSS.n1537 9.01392
R7203 VSS.n1534 VSS.n1533 9.01392
R7204 VSS.n1529 VSS.n1528 9.01392
R7205 VSS.n1526 VSS.n1525 9.01392
R7206 VSS.n1516 VSS.n1515 9.01392
R7207 VSS.n1511 VSS.n1510 9.01392
R7208 VSS.n1507 VSS.n1506 9.01392
R7209 VSS.n1503 VSS.n1502 9.01392
R7210 VSS.n1499 VSS.n1498 9.01392
R7211 VSS.n1493 VSS.n1492 9.01392
R7212 VSS.n1489 VSS.n1488 9.01392
R7213 VSS.n1485 VSS.n1484 9.01392
R7214 VSS.n1481 VSS.n1480 9.01392
R7215 VSS.n1476 VSS.n1475 9.01392
R7216 VSS.n1472 VSS.n1471 9.01392
R7217 VSS.n1468 VSS.n1467 9.01392
R7218 VSS.n1464 VSS.n1463 9.01392
R7219 VSS.n1460 VSS.n1459 9.01392
R7220 VSS.n1454 VSS.n1453 9.01392
R7221 VSS.n1450 VSS.n1449 9.01392
R7222 VSS.n1446 VSS.n1445 9.01392
R7223 VSS.n1442 VSS.n1441 9.01392
R7224 VSS.n1437 VSS.n1436 9.01392
R7225 VSS.n1433 VSS.n1432 9.01392
R7226 VSS.n1428 VSS.n1427 9.01392
R7227 VSS.n1425 VSS.n1424 9.01392
R7228 VSS.n1415 VSS.n1414 9.01392
R7229 VSS.n1410 VSS.n1409 9.01392
R7230 VSS.n1406 VSS.n1405 9.01392
R7231 VSS.n1402 VSS.n1401 9.01392
R7232 VSS.n1398 VSS.n1397 9.01392
R7233 VSS.n1392 VSS.n1391 9.01392
R7234 VSS.n1388 VSS.n1387 9.01392
R7235 VSS.n1384 VSS.n1383 9.01392
R7236 VSS.n1380 VSS.n1379 9.01392
R7237 VSS.n1375 VSS.n1374 9.01392
R7238 VSS.n1371 VSS.n1370 9.01392
R7239 VSS.n1367 VSS.n1366 9.01392
R7240 VSS.n1363 VSS.n1362 9.01392
R7241 VSS.n1359 VSS.n1358 9.01392
R7242 VSS.n1353 VSS.n1352 9.01392
R7243 VSS.n1349 VSS.n1348 9.01392
R7244 VSS.n1345 VSS.n1344 9.01392
R7245 VSS.n1341 VSS.n1340 9.01392
R7246 VSS.n1336 VSS.n1335 9.01392
R7247 VSS.n1332 VSS.n1331 9.01392
R7248 VSS.n55 VSS.n54 9.01392
R7249 VSS.n3359 VSS.n3358 9.01392
R7250 VSS.n3365 VSS.n3364 9.01392
R7251 VSS.n3369 VSS.n3368 9.01392
R7252 VSS.n3373 VSS.n3372 9.01392
R7253 VSS.n3348 VSS.n3347 9.01392
R7254 VSS.n1835 VSS.n1834 9.01392
R7255 VSS.n1834 VSS.n1833 9.01392
R7256 VSS.n3068 VSS.n3067 9.01392
R7257 VSS.n3064 VSS.n3063 9.01392
R7258 VSS.n1881 VSS.n1880 9.01392
R7259 VSS.n1871 VSS.n1870 9.01392
R7260 VSS.n1867 VSS.n1866 9.01392
R7261 VSS.n1859 VSS.n1858 9.01392
R7262 VSS.n1845 VSS.n1844 9.01392
R7263 VSS.n1237 VSS.n1236 9.01392
R7264 VSS.n1232 VSS.n1231 9.01392
R7265 VSS.n1228 VSS.n1227 9.01392
R7266 VSS.n1224 VSS.n1223 9.01392
R7267 VSS.n1220 VSS.n1219 9.01392
R7268 VSS.n1214 VSS.n1213 9.01392
R7269 VSS.n1210 VSS.n1209 9.01392
R7270 VSS.n1206 VSS.n1205 9.01392
R7271 VSS.n1202 VSS.n1201 9.01392
R7272 VSS.n1197 VSS.n1196 9.01392
R7273 VSS.n1193 VSS.n1192 9.01392
R7274 VSS.n1189 VSS.n1188 9.01392
R7275 VSS.n1185 VSS.n1184 9.01392
R7276 VSS.n1181 VSS.n1180 9.01392
R7277 VSS.n1175 VSS.n1174 9.01392
R7278 VSS.n1171 VSS.n1170 9.01392
R7279 VSS.n1167 VSS.n1166 9.01392
R7280 VSS.n1163 VSS.n1162 9.01392
R7281 VSS.n1158 VSS.n1157 9.01392
R7282 VSS.n1154 VSS.n1153 9.01392
R7283 VSS.n1149 VSS.n1148 9.01392
R7284 VSS.n1146 VSS.n1145 9.01392
R7285 VSS.n1136 VSS.n1135 9.01392
R7286 VSS.n1131 VSS.n1130 9.01392
R7287 VSS.n1127 VSS.n1126 9.01392
R7288 VSS.n1123 VSS.n1122 9.01392
R7289 VSS.n1119 VSS.n1118 9.01392
R7290 VSS.n1113 VSS.n1112 9.01392
R7291 VSS.n1109 VSS.n1108 9.01392
R7292 VSS.n1105 VSS.n1104 9.01392
R7293 VSS.n1101 VSS.n1100 9.01392
R7294 VSS.n1096 VSS.n1095 9.01392
R7295 VSS.n3837 VSS.n3836 9.01392
R7296 VSS.n3838 VSS.n3837 9.01392
R7297 VSS.n4126 VSS.n4125 9.01392
R7298 VSS.n4123 VSS.n4122 9.01392
R7299 VSS.n3853 VSS.n3852 9.01392
R7300 VSS.n3855 VSS.n3854 9.01392
R7301 VSS.n3859 VSS.n3858 9.01392
R7302 VSS.n3865 VSS.n3864 9.01392
R7303 VSS.n3870 VSS.n3869 9.01392
R7304 VSS.n3842 VSS.n3841 9.01392
R7305 VSS.n3841 VSS.n3840 9.01392
R7306 VSS.n1826 VSS.n1825 9.01392
R7307 VSS.n1818 VSS.n1817 9.01392
R7308 VSS.n1252 VSS.n1251 9.01392
R7309 VSS.n1813 VSS.n1812 9.01392
R7310 VSS.n1809 VSS.n1808 9.01392
R7311 VSS.n1805 VSS.n1804 9.01392
R7312 VSS.n1801 VSS.n1800 9.01392
R7313 VSS.n1795 VSS.n1794 9.01392
R7314 VSS.n1791 VSS.n1790 9.01392
R7315 VSS.n1787 VSS.n1786 9.01392
R7316 VSS.n1783 VSS.n1782 9.01392
R7317 VSS.n1778 VSS.n1777 9.01392
R7318 VSS.n1774 VSS.n1773 9.01392
R7319 VSS.n1770 VSS.n1769 9.01392
R7320 VSS.n1766 VSS.n1765 9.01392
R7321 VSS.n1762 VSS.n1761 9.01392
R7322 VSS.n1756 VSS.n1755 9.01392
R7323 VSS.n1752 VSS.n1751 9.01392
R7324 VSS.n1748 VSS.n1747 9.01392
R7325 VSS.n1744 VSS.n1743 9.01392
R7326 VSS.n1256 VSS.n1255 9.01392
R7327 VSS.n1739 VSS.n1738 9.01392
R7328 VSS.n1735 VSS.n1734 9.01392
R7329 VSS.n1261 VSS.n1260 9.01392
R7330 VSS.n1730 VSS.n1729 9.01392
R7331 VSS.n1727 VSS.n1726 9.01392
R7332 VSS.n1725 VSS.n1724 9.01392
R7333 VSS.n1717 VSS.n1716 9.01392
R7334 VSS.n1267 VSS.n1266 9.01392
R7335 VSS.n1712 VSS.n1711 9.01392
R7336 VSS.n1708 VSS.n1707 9.01392
R7337 VSS.n1704 VSS.n1703 9.01392
R7338 VSS.n1700 VSS.n1699 9.01392
R7339 VSS.n1694 VSS.n1693 9.01392
R7340 VSS.n1690 VSS.n1689 9.01392
R7341 VSS.n1686 VSS.n1685 9.01392
R7342 VSS.n1682 VSS.n1681 9.01392
R7343 VSS.n1677 VSS.n1676 9.01392
R7344 VSS.n1673 VSS.n1672 9.01392
R7345 VSS.n1669 VSS.n1668 9.01392
R7346 VSS.n1665 VSS.n1664 9.01392
R7347 VSS.n1661 VSS.n1660 9.01392
R7348 VSS.n1655 VSS.n1654 9.01392
R7349 VSS.n1651 VSS.n1650 9.01392
R7350 VSS.n1647 VSS.n1646 9.01392
R7351 VSS.n1643 VSS.n1642 9.01392
R7352 VSS.n1271 VSS.n1270 9.01392
R7353 VSS.n1638 VSS.n1637 9.01392
R7354 VSS.n1634 VSS.n1633 9.01392
R7355 VSS.n1276 VSS.n1275 9.01392
R7356 VSS.n1629 VSS.n1628 9.01392
R7357 VSS.n1626 VSS.n1625 9.01392
R7358 VSS.n1624 VSS.n1623 9.01392
R7359 VSS.n1616 VSS.n1615 9.01392
R7360 VSS.n1282 VSS.n1281 9.01392
R7361 VSS.n1611 VSS.n1610 9.01392
R7362 VSS.n1607 VSS.n1606 9.01392
R7363 VSS.n1603 VSS.n1602 9.01392
R7364 VSS.n1599 VSS.n1598 9.01392
R7365 VSS.n1593 VSS.n1592 9.01392
R7366 VSS.n1589 VSS.n1588 9.01392
R7367 VSS.n1585 VSS.n1584 9.01392
R7368 VSS.n1581 VSS.n1580 9.01392
R7369 VSS.n1576 VSS.n1575 9.01392
R7370 VSS.n1572 VSS.n1571 9.01392
R7371 VSS.n1568 VSS.n1567 9.01392
R7372 VSS.n1564 VSS.n1563 9.01392
R7373 VSS.n1560 VSS.n1559 9.01392
R7374 VSS.n1554 VSS.n1553 9.01392
R7375 VSS.n1550 VSS.n1549 9.01392
R7376 VSS.n1546 VSS.n1545 9.01392
R7377 VSS.n1542 VSS.n1541 9.01392
R7378 VSS.n1286 VSS.n1285 9.01392
R7379 VSS.n1537 VSS.n1536 9.01392
R7380 VSS.n1533 VSS.n1532 9.01392
R7381 VSS.n1291 VSS.n1290 9.01392
R7382 VSS.n1528 VSS.n1527 9.01392
R7383 VSS.n1525 VSS.n1524 9.01392
R7384 VSS.n1523 VSS.n1522 9.01392
R7385 VSS.n1515 VSS.n1514 9.01392
R7386 VSS.n1297 VSS.n1296 9.01392
R7387 VSS.n1510 VSS.n1509 9.01392
R7388 VSS.n1506 VSS.n1505 9.01392
R7389 VSS.n1502 VSS.n1501 9.01392
R7390 VSS.n1498 VSS.n1497 9.01392
R7391 VSS.n1492 VSS.n1491 9.01392
R7392 VSS.n1488 VSS.n1487 9.01392
R7393 VSS.n1484 VSS.n1483 9.01392
R7394 VSS.n1480 VSS.n1479 9.01392
R7395 VSS.n1475 VSS.n1474 9.01392
R7396 VSS.n1471 VSS.n1470 9.01392
R7397 VSS.n1467 VSS.n1466 9.01392
R7398 VSS.n1463 VSS.n1462 9.01392
R7399 VSS.n1459 VSS.n1458 9.01392
R7400 VSS.n1453 VSS.n1452 9.01392
R7401 VSS.n1449 VSS.n1448 9.01392
R7402 VSS.n1445 VSS.n1444 9.01392
R7403 VSS.n1441 VSS.n1440 9.01392
R7404 VSS.n1301 VSS.n1300 9.01392
R7405 VSS.n1436 VSS.n1435 9.01392
R7406 VSS.n1432 VSS.n1431 9.01392
R7407 VSS.n1306 VSS.n1305 9.01392
R7408 VSS.n1427 VSS.n1426 9.01392
R7409 VSS.n1424 VSS.n1423 9.01392
R7410 VSS.n1422 VSS.n1421 9.01392
R7411 VSS.n1414 VSS.n1413 9.01392
R7412 VSS.n1312 VSS.n1311 9.01392
R7413 VSS.n1409 VSS.n1408 9.01392
R7414 VSS.n1405 VSS.n1404 9.01392
R7415 VSS.n1401 VSS.n1400 9.01392
R7416 VSS.n1397 VSS.n1396 9.01392
R7417 VSS.n1391 VSS.n1390 9.01392
R7418 VSS.n1387 VSS.n1386 9.01392
R7419 VSS.n1383 VSS.n1382 9.01392
R7420 VSS.n1379 VSS.n1378 9.01392
R7421 VSS.n1374 VSS.n1373 9.01392
R7422 VSS.n1370 VSS.n1369 9.01392
R7423 VSS.n1366 VSS.n1365 9.01392
R7424 VSS.n1362 VSS.n1361 9.01392
R7425 VSS.n1358 VSS.n1357 9.01392
R7426 VSS.n1352 VSS.n1351 9.01392
R7427 VSS.n1348 VSS.n1347 9.01392
R7428 VSS.n1344 VSS.n1343 9.01392
R7429 VSS.n1340 VSS.n1339 9.01392
R7430 VSS.n1316 VSS.n1315 9.01392
R7431 VSS.n1335 VSS.n1334 9.01392
R7432 VSS.n1331 VSS.n1330 9.01392
R7433 VSS.n1321 VSS.n1320 9.01392
R7434 VSS.n1327 VSS.n1326 9.01392
R7435 VSS.n1326 VSS.n1325 9.01392
R7436 VSS.n3347 VSS.n3346 9.01392
R7437 VSS.n54 VSS.n53 9.01392
R7438 VSS.n3352 VSS.n3351 9.01392
R7439 VSS.n3358 VSS.n3357 9.01392
R7440 VSS.n3364 VSS.n3363 9.01392
R7441 VSS.n3370 VSS.n3369 9.01392
R7442 VSS.n3372 VSS.n3371 9.01392
R7443 VSS.n3376 VSS.n3375 9.01392
R7444 VSS.n3383 VSS.n3382 9.01392
R7445 VSS.n3384 VSS.n3383 9.01392
R7446 VSS.n1838 VSS.n1837 9.01392
R7447 VSS.n1844 VSS.n1843 9.01392
R7448 VSS.n1852 VSS.n1851 9.01392
R7449 VSS.n1858 VSS.n1857 9.01392
R7450 VSS.n1866 VSS.n1865 9.01392
R7451 VSS.n1870 VSS.n1869 9.01392
R7452 VSS.n1880 VSS.n1879 9.01392
R7453 VSS.n3063 VSS.n3062 9.01392
R7454 VSS.n3067 VSS.n3066 9.01392
R7455 VSS.n3072 VSS.n3071 9.01392
R7456 VSS.n3073 VSS.n3072 9.01392
R7457 VSS.n1877 VSS.n1876 9.01392
R7458 VSS.n1876 VSS.n1875 9.01392
R7459 VSS.n1863 VSS.n1862 9.01392
R7460 VSS.n1862 VSS.n1861 9.01392
R7461 VSS.n1849 VSS.n1848 9.01392
R7462 VSS.n1848 VSS.n1847 9.01392
R7463 VSS.n1245 VSS.n1244 9.01392
R7464 VSS.n1236 VSS.n1235 9.01392
R7465 VSS.n124 VSS.n123 9.01392
R7466 VSS.n1231 VSS.n1230 9.01392
R7467 VSS.n1227 VSS.n1226 9.01392
R7468 VSS.n1223 VSS.n1222 9.01392
R7469 VSS.n1219 VSS.n1218 9.01392
R7470 VSS.n1213 VSS.n1212 9.01392
R7471 VSS.n1209 VSS.n1208 9.01392
R7472 VSS.n1205 VSS.n1204 9.01392
R7473 VSS.n1201 VSS.n1200 9.01392
R7474 VSS.n1196 VSS.n1195 9.01392
R7475 VSS.n1192 VSS.n1191 9.01392
R7476 VSS.n1188 VSS.n1187 9.01392
R7477 VSS.n1184 VSS.n1183 9.01392
R7478 VSS.n1180 VSS.n1179 9.01392
R7479 VSS.n1174 VSS.n1173 9.01392
R7480 VSS.n1170 VSS.n1169 9.01392
R7481 VSS.n1166 VSS.n1165 9.01392
R7482 VSS.n1162 VSS.n1161 9.01392
R7483 VSS.n128 VSS.n127 9.01392
R7484 VSS.n1157 VSS.n1156 9.01392
R7485 VSS.n1153 VSS.n1152 9.01392
R7486 VSS.n133 VSS.n132 9.01392
R7487 VSS.n1148 VSS.n1147 9.01392
R7488 VSS.n1145 VSS.n1144 9.01392
R7489 VSS.n1143 VSS.n1142 9.01392
R7490 VSS.n1135 VSS.n1134 9.01392
R7491 VSS.n139 VSS.n138 9.01392
R7492 VSS.n1130 VSS.n1129 9.01392
R7493 VSS.n1126 VSS.n1125 9.01392
R7494 VSS.n1122 VSS.n1121 9.01392
R7495 VSS.n1118 VSS.n1117 9.01392
R7496 VSS.n1112 VSS.n1111 9.01392
R7497 VSS.n1108 VSS.n1107 9.01392
R7498 VSS.n1104 VSS.n1103 9.01392
R7499 VSS.n1100 VSS.n1099 9.01392
R7500 VSS.n1095 VSS.n1094 9.01392
R7501 VSS.n1248 VSS.n1247 9.01392
R7502 VSS.n1247 VSS.n1246 9.01392
R7503 VSS.n3830 VSS.n3829 9.01392
R7504 VSS.n3827 VSS.n3826 9.01392
R7505 VSS.n3826 VSS.n3825 9.01392
R7506 VSS.n3821 VSS.n3820 9.01392
R7507 VSS.n3818 VSS.n3817 9.01392
R7508 VSS.n3817 VSS.n3816 9.01392
R7509 VSS.n3814 VSS.n3813 9.01392
R7510 VSS.n3813 VSS.n3812 9.01392
R7511 VSS.n3810 VSS.n3809 9.01392
R7512 VSS.n3809 VSS.n3808 9.01392
R7513 VSS.n3806 VSS.n3805 9.01392
R7514 VSS.n3805 VSS.n3804 9.01392
R7515 VSS.n3800 VSS.n3799 9.01392
R7516 VSS.n3799 VSS.n3798 9.01392
R7517 VSS.n3796 VSS.n3795 9.01392
R7518 VSS.n3795 VSS.n3794 9.01392
R7519 VSS.n3792 VSS.n3791 9.01392
R7520 VSS.n3791 VSS.n3790 9.01392
R7521 VSS.n3788 VSS.n3787 9.01392
R7522 VSS.n3787 VSS.n3786 9.01392
R7523 VSS.n3783 VSS.n3782 9.01392
R7524 VSS.n3782 VSS.n3781 9.01392
R7525 VSS.n3779 VSS.n3778 9.01392
R7526 VSS.n3778 VSS.n3777 9.01392
R7527 VSS.n3775 VSS.n3774 9.01392
R7528 VSS.n3774 VSS.n3773 9.01392
R7529 VSS.n3771 VSS.n3770 9.01392
R7530 VSS.n3770 VSS.n3769 9.01392
R7531 VSS.n3767 VSS.n3766 9.01392
R7532 VSS.n3766 VSS.n3765 9.01392
R7533 VSS.n3761 VSS.n3760 9.01392
R7534 VSS.n3760 VSS.n3759 9.01392
R7535 VSS.n3757 VSS.n3756 9.01392
R7536 VSS.n3756 VSS.n3755 9.01392
R7537 VSS.n3753 VSS.n3752 9.01392
R7538 VSS.n3752 VSS.n3751 9.01392
R7539 VSS.n3749 VSS.n3748 9.01392
R7540 VSS.n3748 VSS.n3747 9.01392
R7541 VSS.n3742 VSS.n3741 9.01392
R7542 VSS.n3739 VSS.n3738 9.01392
R7543 VSS.n3738 VSS.n3737 9.01392
R7544 VSS.n3735 VSS.n3734 9.01392
R7545 VSS.n3734 VSS.n3733 9.01392
R7546 VSS.n3728 VSS.n3727 9.01392
R7547 VSS.n3725 VSS.n3724 9.01392
R7548 VSS.n3724 VSS.n3723 9.01392
R7549 VSS.n3715 VSS.n3385 9.01392
R7550 VSS.n3722 VSS.n3385 9.01392
R7551 VSS.n3721 VSS.n3720 9.01392
R7552 VSS.n3713 VSS.n3712 9.01392
R7553 VSS.n3712 VSS.n3711 9.01392
R7554 VSS.n3707 VSS.n3706 9.01392
R7555 VSS.n3704 VSS.n3703 9.01392
R7556 VSS.n3703 VSS.n3702 9.01392
R7557 VSS.n3700 VSS.n3699 9.01392
R7558 VSS.n3699 VSS.n3698 9.01392
R7559 VSS.n3696 VSS.n3695 9.01392
R7560 VSS.n3695 VSS.n3694 9.01392
R7561 VSS.n3692 VSS.n3691 9.01392
R7562 VSS.n3691 VSS.n3690 9.01392
R7563 VSS.n3686 VSS.n3685 9.01392
R7564 VSS.n3685 VSS.n3684 9.01392
R7565 VSS.n3682 VSS.n3681 9.01392
R7566 VSS.n3681 VSS.n3680 9.01392
R7567 VSS.n3678 VSS.n3677 9.01392
R7568 VSS.n3677 VSS.n3676 9.01392
R7569 VSS.n3674 VSS.n3673 9.01392
R7570 VSS.n3673 VSS.n3672 9.01392
R7571 VSS.n3669 VSS.n3668 9.01392
R7572 VSS.n3668 VSS.n3667 9.01392
R7573 VSS.n3665 VSS.n3664 9.01392
R7574 VSS.n3664 VSS.n3663 9.01392
R7575 VSS.n3661 VSS.n3660 9.01392
R7576 VSS.n3660 VSS.n3659 9.01392
R7577 VSS.n3657 VSS.n3656 9.01392
R7578 VSS.n3656 VSS.n3655 9.01392
R7579 VSS.n3653 VSS.n3652 9.01392
R7580 VSS.n3652 VSS.n3651 9.01392
R7581 VSS.n3647 VSS.n3646 9.01392
R7582 VSS.n3646 VSS.n3645 9.01392
R7583 VSS.n3643 VSS.n3642 9.01392
R7584 VSS.n3642 VSS.n3641 9.01392
R7585 VSS.n3639 VSS.n3638 9.01392
R7586 VSS.n3638 VSS.n3637 9.01392
R7587 VSS.n3635 VSS.n3634 9.01392
R7588 VSS.n3634 VSS.n3633 9.01392
R7589 VSS.n3628 VSS.n3627 9.01392
R7590 VSS.n3625 VSS.n3624 9.01392
R7591 VSS.n3624 VSS.n3623 9.01392
R7592 VSS.n3621 VSS.n3620 9.01392
R7593 VSS.n3620 VSS.n3619 9.01392
R7594 VSS.n3614 VSS.n3613 9.01392
R7595 VSS.n3611 VSS.n3610 9.01392
R7596 VSS.n3610 VSS.n3609 9.01392
R7597 VSS.n3601 VSS.n3387 9.01392
R7598 VSS.n3608 VSS.n3387 9.01392
R7599 VSS.n3607 VSS.n3606 9.01392
R7600 VSS.n3599 VSS.n3598 9.01392
R7601 VSS.n3598 VSS.n3597 9.01392
R7602 VSS.n3593 VSS.n3592 9.01392
R7603 VSS.n3590 VSS.n3589 9.01392
R7604 VSS.n3589 VSS.n3588 9.01392
R7605 VSS.n3586 VSS.n3585 9.01392
R7606 VSS.n3585 VSS.n3584 9.01392
R7607 VSS.n3582 VSS.n3581 9.01392
R7608 VSS.n3581 VSS.n3580 9.01392
R7609 VSS.n3578 VSS.n3577 9.01392
R7610 VSS.n3577 VSS.n3576 9.01392
R7611 VSS.n3572 VSS.n3571 9.01392
R7612 VSS.n3571 VSS.n3570 9.01392
R7613 VSS.n3568 VSS.n3567 9.01392
R7614 VSS.n3567 VSS.n3566 9.01392
R7615 VSS.n3564 VSS.n3563 9.01392
R7616 VSS.n3563 VSS.n3562 9.01392
R7617 VSS.n3560 VSS.n3559 9.01392
R7618 VSS.n3559 VSS.n3558 9.01392
R7619 VSS.n3555 VSS.n3554 9.01392
R7620 VSS.n3554 VSS.n3553 9.01392
R7621 VSS.n3551 VSS.n3550 9.01392
R7622 VSS.n3550 VSS.n3549 9.01392
R7623 VSS.n3547 VSS.n3546 9.01392
R7624 VSS.n3546 VSS.n3545 9.01392
R7625 VSS.n3543 VSS.n3542 9.01392
R7626 VSS.n3542 VSS.n3541 9.01392
R7627 VSS.n3539 VSS.n3538 9.01392
R7628 VSS.n3538 VSS.n3537 9.01392
R7629 VSS.n3533 VSS.n3532 9.01392
R7630 VSS.n3532 VSS.n3531 9.01392
R7631 VSS.n3529 VSS.n3528 9.01392
R7632 VSS.n3528 VSS.n3527 9.01392
R7633 VSS.n3525 VSS.n3524 9.01392
R7634 VSS.n3524 VSS.n3523 9.01392
R7635 VSS.n3521 VSS.n3520 9.01392
R7636 VSS.n3520 VSS.n3519 9.01392
R7637 VSS.n3514 VSS.n3513 9.01392
R7638 VSS.n3511 VSS.n3510 9.01392
R7639 VSS.n3510 VSS.n3509 9.01392
R7640 VSS.n3507 VSS.n3506 9.01392
R7641 VSS.n3506 VSS.n3505 9.01392
R7642 VSS.n3500 VSS.n3499 9.01392
R7643 VSS.n3497 VSS.n3496 9.01392
R7644 VSS.n3496 VSS.n3495 9.01392
R7645 VSS.n3487 VSS.n3389 9.01392
R7646 VSS.n3494 VSS.n3389 9.01392
R7647 VSS.n3493 VSS.n3492 9.01392
R7648 VSS.n3485 VSS.n3484 9.01392
R7649 VSS.n3484 VSS.n3483 9.01392
R7650 VSS.n3479 VSS.n3478 9.01392
R7651 VSS.n3476 VSS.n3475 9.01392
R7652 VSS.n3475 VSS.n3474 9.01392
R7653 VSS.n3472 VSS.n3471 9.01392
R7654 VSS.n3471 VSS.n3470 9.01392
R7655 VSS.n3468 VSS.n3467 9.01392
R7656 VSS.n3467 VSS.n3466 9.01392
R7657 VSS.n3464 VSS.n3463 9.01392
R7658 VSS.n3463 VSS.n3462 9.01392
R7659 VSS.n3458 VSS.n3457 9.01392
R7660 VSS.n3457 VSS.n3456 9.01392
R7661 VSS.n3454 VSS.n3453 9.01392
R7662 VSS.n3453 VSS.n3452 9.01392
R7663 VSS.n3450 VSS.n3449 9.01392
R7664 VSS.n3449 VSS.n3448 9.01392
R7665 VSS.n3446 VSS.n3445 9.01392
R7666 VSS.n3445 VSS.n3444 9.01392
R7667 VSS.n3441 VSS.n3440 9.01392
R7668 VSS.n3440 VSS.n3439 9.01392
R7669 VSS.n3437 VSS.n3436 9.01392
R7670 VSS.n3436 VSS.n3435 9.01392
R7671 VSS.n3433 VSS.n3432 9.01392
R7672 VSS.n3432 VSS.n3431 9.01392
R7673 VSS.n3429 VSS.n3428 9.01392
R7674 VSS.n3428 VSS.n3427 9.01392
R7675 VSS.n3425 VSS.n3424 9.01392
R7676 VSS.n3424 VSS.n3423 9.01392
R7677 VSS.n3419 VSS.n3418 9.01392
R7678 VSS.n3418 VSS.n3417 9.01392
R7679 VSS.n3415 VSS.n3414 9.01392
R7680 VSS.n3414 VSS.n3413 9.01392
R7681 VSS.n3411 VSS.n3410 9.01392
R7682 VSS.n3410 VSS.n3409 9.01392
R7683 VSS.n3407 VSS.n3406 9.01392
R7684 VSS.n3406 VSS.n3405 9.01392
R7685 VSS.n3400 VSS.n3399 9.01392
R7686 VSS.n3397 VSS.n3396 9.01392
R7687 VSS.n3396 VSS.n3395 9.01392
R7688 VSS.n3393 VSS.n3392 9.01392
R7689 VSS.n3392 VSS.n3391 9.01392
R7690 VSS.n2 VSS.n1 9.01392
R7691 VSS.n4237 VSS.n4236 9.01392
R7692 VSS.n4236 VSS.n4235 9.01392
R7693 VSS.n4233 VSS.n4232 9.01392
R7694 VSS.n4234 VSS.n4233 9.01392
R7695 VSS.n4231 VSS.n4230 9.01392
R7696 VSS.n4225 VSS.n4224 9.01392
R7697 VSS.n4224 VSS.n4223 9.01392
R7698 VSS.n4219 VSS.n4218 9.01392
R7699 VSS.n4216 VSS.n4215 9.01392
R7700 VSS.n4215 VSS.n4214 9.01392
R7701 VSS.n4212 VSS.n4211 9.01392
R7702 VSS.n4211 VSS.n4210 9.01392
R7703 VSS.n4208 VSS.n4207 9.01392
R7704 VSS.n4207 VSS.n4206 9.01392
R7705 VSS.n4204 VSS.n4203 9.01392
R7706 VSS.n4203 VSS.n4202 9.01392
R7707 VSS.n4198 VSS.n4197 9.01392
R7708 VSS.n4197 VSS.n4196 9.01392
R7709 VSS.n4194 VSS.n4193 9.01392
R7710 VSS.n4193 VSS.n4192 9.01392
R7711 VSS.n4190 VSS.n4189 9.01392
R7712 VSS.n4189 VSS.n4188 9.01392
R7713 VSS.n4186 VSS.n4185 9.01392
R7714 VSS.n4185 VSS.n4184 9.01392
R7715 VSS.n4181 VSS.n4180 9.01392
R7716 VSS.n4180 VSS.n4179 9.01392
R7717 VSS.n4177 VSS.n4176 9.01392
R7718 VSS.n4176 VSS.n4175 9.01392
R7719 VSS.n4173 VSS.n4172 9.01392
R7720 VSS.n4172 VSS.n4171 9.01392
R7721 VSS.n4169 VSS.n4168 9.01392
R7722 VSS.n4168 VSS.n4167 9.01392
R7723 VSS.n4165 VSS.n4164 9.01392
R7724 VSS.n4164 VSS.n4163 9.01392
R7725 VSS.n4159 VSS.n4158 9.01392
R7726 VSS.n4158 VSS.n4157 9.01392
R7727 VSS.n4155 VSS.n4154 9.01392
R7728 VSS.n4154 VSS.n4153 9.01392
R7729 VSS.n4151 VSS.n4150 9.01392
R7730 VSS.n4150 VSS.n4149 9.01392
R7731 VSS.n4147 VSS.n4146 9.01392
R7732 VSS.n4146 VSS.n4145 9.01392
R7733 VSS.n4140 VSS.n4139 9.01392
R7734 VSS.n4137 VSS.n4136 9.01392
R7735 VSS.n4136 VSS.n4135 9.01392
R7736 VSS.n4133 VSS.n4132 9.01392
R7737 VSS.n4132 VSS.n4131 9.01392
R7738 VSS.n4122 VSS.n4121 9.01392
R7739 VSS.n1246 VSS 8.8005
R7740 VSS.n1208 VSS.t29 8.8005
R7741 VSS.n1144 VSS 8.8005
R7742 VSS.n1107 VSS.t433 8.8005
R7743 VSS.n848 VSS.t229 8.8005
R7744 VSS.n820 VSS.t378 8.8005
R7745 VSS.n539 VSS.t219 8.8005
R7746 VSS.n511 VSS.t146 8.8005
R7747 VSS.n3074 VSS.n70 8.8005
R7748 VSS.n89 VSS.n86 8.76429
R7749 VSS.n82 VSS.n81 8.76429
R7750 VSS.n1877 VSS.n1874 8.6074
R7751 VSS.n1243 VSS 8.6074
R7752 VSS.n1181 VSS.n1178 8.6074
R7753 VSS.n1141 VSS 8.6074
R7754 VSS.n932 VSS 8.6074
R7755 VSS.n623 VSS 8.6074
R7756 VSS.n3095 VSS.n3094 8.6074
R7757 VSS.n1763 VSS.n1760 8.6074
R7758 VSS.n1662 VSS.n1659 8.6074
R7759 VSS.n1561 VSS.n1558 8.6074
R7760 VSS.n1460 VSS.n1457 8.6074
R7761 VSS.n1359 VSS.n1356 8.6074
R7762 VSS.n4165 VSS.n4162 8.6074
R7763 VSS.n3425 VSS.n3422 8.6074
R7764 VSS.n3539 VSS.n3536 8.6074
R7765 VSS.n3653 VSS.n3650 8.6074
R7766 VSS.n3767 VSS.n3764 8.6074
R7767 VSS.t88 VSS.n21 8.5775
R7768 VSS.n1939 VSS.t86 8.5775
R7769 VSS.n2029 VSS 8.5775
R7770 VSS.t38 VSS.n2146 8.5775
R7771 VSS.t139 VSS.n2497 8.5775
R7772 VSS.t321 VSS.n2848 8.5775
R7773 VSS.n3260 VSS.n3259 7.72464
R7774 VSS.n161 VSS.n160 7.57647
R7775 VSS.n215 VSS.n214 7.57647
R7776 VSS.n269 VSS.n268 7.57647
R7777 VSS.n2345 VSS.n2344 7.57501
R7778 VSS.n2415 VSS.n2414 7.57501
R7779 VSS.n2696 VSS.n2695 7.57501
R7780 VSS.n2766 VSS.n2765 7.57501
R7781 VSS.n3047 VSS.n3046 7.57501
R7782 VSS.n2318 VSS.n2317 7.57431
R7783 VSS.n2669 VSS.n2668 7.57431
R7784 VSS.n3020 VSS.n3019 7.57431
R7785 VSS.n866 VSS.n865 7.50395
R7786 VSS.n557 VSS.n556 7.50395
R7787 VSS.n2001 VSS.n1996 7.45502
R7788 VSS.n2021 VSS.n2016 7.43981
R7789 VSS.n2075 VSS.n2070 7.43981
R7790 VSS.n2838 VSS.n2837 6.84188
R7791 VSS.n2487 VSS.n2486 6.84188
R7792 VSS.n2136 VSS.n2135 6.84188
R7793 VSS.n90 VSS 6.66075
R7794 VSS.n4115 VSS.n4114 6.62119
R7795 VSS.n3120 VSS.t481 6.37269
R7796 VSS.n3271 VSS.t279 6.37269
R7797 VSS.n10 VSS.n9 5.71609
R7798 VSS.n77 VSS 5.58923
R7799 VSS.n56 VSS.n55 5.51774
R7800 VSS.n1827 VSS 5.26996
R7801 VSS.n1790 VSS.t208 5.26996
R7802 VSS.n1726 VSS 5.26996
R7803 VSS.n1689 VSS.t503 5.26996
R7804 VSS.n1625 VSS 5.26996
R7805 VSS.n1588 VSS.t207 5.26996
R7806 VSS.n1524 VSS 5.26996
R7807 VSS.n1487 VSS.t410 5.26996
R7808 VSS.n1423 VSS 5.26996
R7809 VSS.n1386 VSS.t120 5.26996
R7810 VSS.n81 VSS.n80 5.25868
R7811 VSS.n3125 VSS.n3124 5.07636
R7812 VSS.n2122 VSS.n2121 4.6505
R7813 VSS.n2138 VSS.n2137 4.6505
R7814 VSS.n2152 VSS.n2151 4.6505
R7815 VSS.n2166 VSS.n2165 4.6505
R7816 VSS.n2180 VSS.n2179 4.6505
R7817 VSS.n2194 VSS.n2193 4.6505
R7818 VSS.n2208 VSS.n2207 4.6505
R7819 VSS.n2222 VSS.n2221 4.6505
R7820 VSS.n2236 VSS.n2235 4.6505
R7821 VSS.n2250 VSS.n2249 4.6505
R7822 VSS.n2266 VSS.n2265 4.6505
R7823 VSS.n2280 VSS.n2279 4.6505
R7824 VSS.n2294 VSS.n2293 4.6505
R7825 VSS.n2308 VSS.n2307 4.6505
R7826 VSS.n2334 VSS.n2333 4.6505
R7827 VSS.n2352 VSS.n2351 4.6505
R7828 VSS.n2363 VSS.n2362 4.6505
R7829 VSS.n2390 VSS.n2389 4.6505
R7830 VSS.n2404 VSS.n2403 4.6505
R7831 VSS.n2431 VSS.n2430 4.6505
R7832 VSS.n2445 VSS.n2444 4.6505
R7833 VSS.n2459 VSS.n2458 4.6505
R7834 VSS.n2473 VSS.n2472 4.6505
R7835 VSS.n2489 VSS.n2488 4.6505
R7836 VSS.n2503 VSS.n2502 4.6505
R7837 VSS.n2517 VSS.n2516 4.6505
R7838 VSS.n2531 VSS.n2530 4.6505
R7839 VSS.n2545 VSS.n2544 4.6505
R7840 VSS.n2559 VSS.n2558 4.6505
R7841 VSS.n2573 VSS.n2572 4.6505
R7842 VSS.n2587 VSS.n2586 4.6505
R7843 VSS.n2601 VSS.n2600 4.6505
R7844 VSS.n2617 VSS.n2616 4.6505
R7845 VSS.n2631 VSS.n2630 4.6505
R7846 VSS.n2645 VSS.n2644 4.6505
R7847 VSS.n2659 VSS.n2658 4.6505
R7848 VSS.n2685 VSS.n2684 4.6505
R7849 VSS.n2703 VSS.n2702 4.6505
R7850 VSS.n2714 VSS.n2713 4.6505
R7851 VSS.n2741 VSS.n2740 4.6505
R7852 VSS.n2755 VSS.n2754 4.6505
R7853 VSS.n2782 VSS.n2781 4.6505
R7854 VSS.n2796 VSS.n2795 4.6505
R7855 VSS.n2810 VSS.n2809 4.6505
R7856 VSS.n2824 VSS.n2823 4.6505
R7857 VSS.n2840 VSS.n2839 4.6505
R7858 VSS.n2854 VSS.n2853 4.6505
R7859 VSS.n2868 VSS.n2867 4.6505
R7860 VSS.n2882 VSS.n2881 4.6505
R7861 VSS.n2896 VSS.n2895 4.6505
R7862 VSS.n2910 VSS.n2909 4.6505
R7863 VSS.n2924 VSS.n2923 4.6505
R7864 VSS.n2938 VSS.n2937 4.6505
R7865 VSS.n2952 VSS.n2951 4.6505
R7866 VSS.n2968 VSS.n2967 4.6505
R7867 VSS.n2982 VSS.n2981 4.6505
R7868 VSS.n2996 VSS.n2995 4.6505
R7869 VSS.n3010 VSS.n3009 4.6505
R7870 VSS.n3036 VSS.n3035 4.6505
R7871 VSS.n3056 VSS.n3055 4.6505
R7872 VSS.n1092 VSS.n1091 4.6505
R7873 VSS.n1078 VSS.n1077 4.6505
R7874 VSS.n1064 VSS.n1063 4.6505
R7875 VSS.n1050 VSS.n1049 4.6505
R7876 VSS.n1034 VSS.n1033 4.6505
R7877 VSS.n1020 VSS.n1019 4.6505
R7878 VSS.n1006 VSS.n1005 4.6505
R7879 VSS.n992 VSS.n991 4.6505
R7880 VSS.n975 VSS.n974 4.6505
R7881 VSS.n961 VSS.n960 4.6505
R7882 VSS.n944 VSS.n943 4.6505
R7883 VSS.n184 VSS.n173 4.6505
R7884 VSS.n927 VSS.n926 4.6505
R7885 VSS.n910 VSS.n909 4.6505
R7886 VSS.n896 VSS.n895 4.6505
R7887 VSS.n882 VSS.n881 4.6505
R7888 VSS.n868 VSS.n867 4.6505
R7889 VSS.n853 VSS.n852 4.6505
R7890 VSS.n839 VSS.n838 4.6505
R7891 VSS.n825 VSS.n824 4.6505
R7892 VSS.n811 VSS.n810 4.6505
R7893 VSS.n796 VSS.n795 4.6505
R7894 VSS.n783 VSS.n782 4.6505
R7895 VSS.n769 VSS.n768 4.6505
R7896 VSS.n755 VSS.n754 4.6505
R7897 VSS.n741 VSS.n740 4.6505
R7898 VSS.n725 VSS.n724 4.6505
R7899 VSS.n711 VSS.n710 4.6505
R7900 VSS.n697 VSS.n696 4.6505
R7901 VSS.n683 VSS.n682 4.6505
R7902 VSS.n666 VSS.n665 4.6505
R7903 VSS.n652 VSS.n651 4.6505
R7904 VSS.n635 VSS.n634 4.6505
R7905 VSS.n238 VSS.n227 4.6505
R7906 VSS.n618 VSS.n617 4.6505
R7907 VSS.n601 VSS.n600 4.6505
R7908 VSS.n587 VSS.n586 4.6505
R7909 VSS.n573 VSS.n572 4.6505
R7910 VSS.n559 VSS.n558 4.6505
R7911 VSS.n544 VSS.n543 4.6505
R7912 VSS.n530 VSS.n529 4.6505
R7913 VSS.n516 VSS.n515 4.6505
R7914 VSS.n502 VSS.n501 4.6505
R7915 VSS.n487 VSS.n486 4.6505
R7916 VSS.n474 VSS.n473 4.6505
R7917 VSS.n460 VSS.n459 4.6505
R7918 VSS.n446 VSS.n445 4.6505
R7919 VSS.n432 VSS.n431 4.6505
R7920 VSS.n416 VSS.n415 4.6505
R7921 VSS.n402 VSS.n401 4.6505
R7922 VSS.n388 VSS.n387 4.6505
R7923 VSS.n374 VSS.n373 4.6505
R7924 VSS.n357 VSS.n356 4.6505
R7925 VSS.n343 VSS.n342 4.6505
R7926 VSS.n326 VSS.n325 4.6505
R7927 VSS.n314 VSS.n313 4.6505
R7928 VSS.n310 VSS.n309 4.6505
R7929 VSS.n296 VSS.n295 4.6505
R7930 VSS.n3081 VSS.n3080 4.6505
R7931 VSS.n3097 VSS.n3096 4.6505
R7932 VSS.n3111 VSS.n3110 4.6505
R7933 VSS.n3127 VSS.n3126 4.6505
R7934 VSS.n3140 VSS.n3139 4.6505
R7935 VSS.n3156 VSS.n3155 4.6505
R7936 VSS.n3170 VSS.n3169 4.6505
R7937 VSS.n3186 VSS.n3185 4.6505
R7938 VSS.n3200 VSS.n3199 4.6505
R7939 VSS.n3216 VSS.n3215 4.6505
R7940 VSS.n3230 VSS.n3229 4.6505
R7941 VSS.n3246 VSS.n3245 4.6505
R7942 VSS.n3262 VSS.n3261 4.6505
R7943 VSS.n3276 VSS.n3275 4.6505
R7944 VSS.n3292 VSS.n3291 4.6505
R7945 VSS.n3306 VSS.n3305 4.6505
R7946 VSS.n3322 VSS.n3321 4.6505
R7947 VSS.n3336 VSS.n3335 4.6505
R7948 VSS.n3341 VSS.n3340 4.6505
R7949 VSS.n4101 VSS.n4100 4.6505
R7950 VSS.n4096 VSS.n4095 4.6505
R7951 VSS.n4082 VSS.n4081 4.6505
R7952 VSS.n4066 VSS.n4065 4.6505
R7953 VSS.n4054 VSS.n4053 4.6505
R7954 VSS.n4040 VSS.n4039 4.6505
R7955 VSS.n4026 VSS.n4025 4.6505
R7956 VSS.n4009 VSS.n4008 4.6505
R7957 VSS.n3997 VSS.n3996 4.6505
R7958 VSS.n3983 VSS.n3982 4.6505
R7959 VSS.n3969 VSS.n3968 4.6505
R7960 VSS.n3955 VSS.n3954 4.6505
R7961 VSS.n3940 VSS.n3939 4.6505
R7962 VSS.n3926 VSS.n3925 4.6505
R7963 VSS.n3911 VSS.n3910 4.6505
R7964 VSS.n3897 VSS.n3896 4.6505
R7965 VSS.n86 VSS.n85 4.46346
R7966 VSS.n2320 VSS.n2319 4.43314
R7967 VSS.n2671 VSS.n2670 4.43314
R7968 VSS.n3022 VSS.n3021 4.43314
R7969 VSS.n604 VSS.n249 4.43314
R7970 VSS.n913 VSS.n195 4.43314
R7971 VSS.n2347 VSS.n2346 4.42059
R7972 VSS.n2417 VSS.n2416 4.42059
R7973 VSS.n2698 VSS.n2697 4.42059
R7974 VSS.n2768 VSS.n2767 4.42059
R7975 VSS.n3049 VSS.n3048 4.42059
R7976 VSS.n360 VSS.n259 4.42059
R7977 VSS.n622 VSS.n621 4.42059
R7978 VSS.n669 VSS.n205 4.42059
R7979 VSS.n931 VSS.n930 4.42059
R7980 VSS.n978 VSS.n151 4.42059
R7981 VSS.n4069 VSS.n27 4.42059
R7982 VSS.n4012 VSS.n40 4.42059
R7983 VSS.n4105 VSS.n4104 4.42059
R7984 VSS.n2376 VSS.n2375 4.39476
R7985 VSS.n2727 VSS.n2726 4.39476
R7986 VSS.n329 VSS.n270 4.39476
R7987 VSS.n638 VSS.n216 4.39476
R7988 VSS.n947 VSS.n162 4.39476
R7989 VSS.n3290 VSS.n3289 4.1936
R7990 VSS.n1248 VSS 3.97291
R7991 VSS.n1146 VSS 3.97291
R7992 VSS.n2085 VSS.n2080 3.75222
R7993 VSS.n2095 VSS.n2090 3.75222
R7994 VSS.n2105 VSS.n2100 3.75222
R7995 VSS.n2054 VSS.n2049 3.75222
R7996 VSS.n2064 VSS.n2059 3.75222
R7997 VSS.n122 VSS.n117 3.75222
R7998 VSS.n2033 VSS.n115 3.75222
R7999 VSS.n2010 VSS.n2005 3.75222
R8000 VSS.n1928 VSS.n1923 3.75222
R8001 VSS.n1938 VSS.n1933 3.75222
R8002 VSS.n1948 VSS.n1943 3.75222
R8003 VSS.n1960 VSS.n1955 3.75222
R8004 VSS.n1970 VSS.n1965 3.75222
R8005 VSS.n1980 VSS.n1975 3.75222
R8006 VSS.n1990 VSS.n1985 3.75222
R8007 VSS.n1888 VSS.n1883 3.75222
R8008 VSS.n1898 VSS.n1893 3.75222
R8009 VSS.n1908 VSS.n1903 3.75222
R8010 VSS.n3856 VSS 3.75222
R8011 VSS.n2027 VSS 3.53153
R8012 VSS.n3368 VSS 3.53153
R8013 VSS.n4232 VSS 3.53153
R8014 VSS.n3487 VSS 3.53153
R8015 VSS.n3601 VSS 3.53153
R8016 VSS.n3715 VSS 3.53153
R8017 VSS.n3836 VSS 3.53153
R8018 VSS.n2045 VSS.n2042 3.42435
R8019 VSS.n2957 VSS.n2956 3.31084
R8020 VSS.n2606 VSS.n2605 3.31084
R8021 VSS.n2255 VSS.n2254 3.31084
R8022 VSS.n1955 VSS.n1954 3.31084
R8023 VSS.n3382 VSS 3.31084
R8024 VSS.n3842 VSS 3.31084
R8025 VSS.n3050 VSS.n90 3.19691
R8026 VSS.n3147 VSS.t477 3.1866
R8027 VSS.n2726 VSS.n2724 3.11687
R8028 VSS.n2375 VSS.n2373 3.11687
R8029 VSS.n162 VSS.n161 3.11687
R8030 VSS.n216 VSS.n215 3.11687
R8031 VSS.n270 VSS.n269 3.11687
R8032 VSS.n1846 VSS.n1845 3.1005
R8033 VSS.n1836 VSS.n1835 3.1005
R8034 VSS.n3382 VSS.n3381 3.1005
R8035 VSS.n3851 VSS.n3850 3.1005
R8036 VSS.n3843 VSS.n3842 3.1005
R8037 VSS.n3857 VSS.n3856 3.1005
R8038 VSS.n3867 VSS.n3866 3.1005
R8039 VSS.n3871 VSS.n3868 3.1005
R8040 VSS.n1328 VSS.n1327 3.1005
R8041 VSS.n1830 VSS.n1829 3.1005
R8042 VSS.n1820 VSS.n1819 3.1005
R8043 VSS.n1815 VSS.n1814 3.1005
R8044 VSS.n1811 VSS.n1810 3.1005
R8045 VSS.n1807 VSS.n1806 3.1005
R8046 VSS.n1803 VSS.n1802 3.1005
R8047 VSS.n1797 VSS.n1796 3.1005
R8048 VSS.n1793 VSS.n1792 3.1005
R8049 VSS.n1789 VSS.n1788 3.1005
R8050 VSS.n1785 VSS.n1784 3.1005
R8051 VSS.n1780 VSS.n1779 3.1005
R8052 VSS.n1776 VSS.n1775 3.1005
R8053 VSS.n1772 VSS.n1771 3.1005
R8054 VSS.n1768 VSS.n1767 3.1005
R8055 VSS.n1764 VSS.n1763 3.1005
R8056 VSS.n1758 VSS.n1757 3.1005
R8057 VSS.n1754 VSS.n1753 3.1005
R8058 VSS.n1750 VSS.n1749 3.1005
R8059 VSS.n1746 VSS.n1745 3.1005
R8060 VSS.n1741 VSS.n1740 3.1005
R8061 VSS.n1737 VSS.n1736 3.1005
R8062 VSS.n1732 VSS.n1731 3.1005
R8063 VSS.n1728 VSS.n1265 3.1005
R8064 VSS.n1719 VSS.n1718 3.1005
R8065 VSS.n1714 VSS.n1713 3.1005
R8066 VSS.n1710 VSS.n1709 3.1005
R8067 VSS.n1706 VSS.n1705 3.1005
R8068 VSS.n1702 VSS.n1701 3.1005
R8069 VSS.n1696 VSS.n1695 3.1005
R8070 VSS.n1692 VSS.n1691 3.1005
R8071 VSS.n1688 VSS.n1687 3.1005
R8072 VSS.n1684 VSS.n1683 3.1005
R8073 VSS.n1679 VSS.n1678 3.1005
R8074 VSS.n1675 VSS.n1674 3.1005
R8075 VSS.n1671 VSS.n1670 3.1005
R8076 VSS.n1667 VSS.n1666 3.1005
R8077 VSS.n1663 VSS.n1662 3.1005
R8078 VSS.n1657 VSS.n1656 3.1005
R8079 VSS.n1653 VSS.n1652 3.1005
R8080 VSS.n1649 VSS.n1648 3.1005
R8081 VSS.n1645 VSS.n1644 3.1005
R8082 VSS.n1640 VSS.n1639 3.1005
R8083 VSS.n1636 VSS.n1635 3.1005
R8084 VSS.n1631 VSS.n1630 3.1005
R8085 VSS.n1627 VSS.n1280 3.1005
R8086 VSS.n1618 VSS.n1617 3.1005
R8087 VSS.n1613 VSS.n1612 3.1005
R8088 VSS.n1609 VSS.n1608 3.1005
R8089 VSS.n1605 VSS.n1604 3.1005
R8090 VSS.n1601 VSS.n1600 3.1005
R8091 VSS.n1595 VSS.n1594 3.1005
R8092 VSS.n1591 VSS.n1590 3.1005
R8093 VSS.n1587 VSS.n1586 3.1005
R8094 VSS.n1583 VSS.n1582 3.1005
R8095 VSS.n1578 VSS.n1577 3.1005
R8096 VSS.n1574 VSS.n1573 3.1005
R8097 VSS.n1570 VSS.n1569 3.1005
R8098 VSS.n1566 VSS.n1565 3.1005
R8099 VSS.n1562 VSS.n1561 3.1005
R8100 VSS.n1556 VSS.n1555 3.1005
R8101 VSS.n1552 VSS.n1551 3.1005
R8102 VSS.n1548 VSS.n1547 3.1005
R8103 VSS.n1544 VSS.n1543 3.1005
R8104 VSS.n1539 VSS.n1538 3.1005
R8105 VSS.n1535 VSS.n1534 3.1005
R8106 VSS.n1530 VSS.n1529 3.1005
R8107 VSS.n1526 VSS.n1295 3.1005
R8108 VSS.n1517 VSS.n1516 3.1005
R8109 VSS.n1512 VSS.n1511 3.1005
R8110 VSS.n1508 VSS.n1507 3.1005
R8111 VSS.n1504 VSS.n1503 3.1005
R8112 VSS.n1500 VSS.n1499 3.1005
R8113 VSS.n1494 VSS.n1493 3.1005
R8114 VSS.n1490 VSS.n1489 3.1005
R8115 VSS.n1486 VSS.n1485 3.1005
R8116 VSS.n1482 VSS.n1481 3.1005
R8117 VSS.n1477 VSS.n1476 3.1005
R8118 VSS.n1473 VSS.n1472 3.1005
R8119 VSS.n1469 VSS.n1468 3.1005
R8120 VSS.n1465 VSS.n1464 3.1005
R8121 VSS.n1461 VSS.n1460 3.1005
R8122 VSS.n1455 VSS.n1454 3.1005
R8123 VSS.n1451 VSS.n1450 3.1005
R8124 VSS.n1447 VSS.n1446 3.1005
R8125 VSS.n1443 VSS.n1442 3.1005
R8126 VSS.n1438 VSS.n1437 3.1005
R8127 VSS.n1434 VSS.n1433 3.1005
R8128 VSS.n1429 VSS.n1428 3.1005
R8129 VSS.n1425 VSS.n1310 3.1005
R8130 VSS.n1416 VSS.n1415 3.1005
R8131 VSS.n1411 VSS.n1410 3.1005
R8132 VSS.n1407 VSS.n1406 3.1005
R8133 VSS.n1403 VSS.n1402 3.1005
R8134 VSS.n1399 VSS.n1398 3.1005
R8135 VSS.n1393 VSS.n1392 3.1005
R8136 VSS.n1389 VSS.n1388 3.1005
R8137 VSS.n1385 VSS.n1384 3.1005
R8138 VSS.n1381 VSS.n1380 3.1005
R8139 VSS.n1376 VSS.n1375 3.1005
R8140 VSS.n1372 VSS.n1371 3.1005
R8141 VSS.n1368 VSS.n1367 3.1005
R8142 VSS.n1364 VSS.n1363 3.1005
R8143 VSS.n1360 VSS.n1359 3.1005
R8144 VSS.n1354 VSS.n1353 3.1005
R8145 VSS.n1350 VSS.n1349 3.1005
R8146 VSS.n1346 VSS.n1345 3.1005
R8147 VSS.n1342 VSS.n1341 3.1005
R8148 VSS.n1337 VSS.n1336 3.1005
R8149 VSS.n1333 VSS.n1332 3.1005
R8150 VSS.n3349 VSS.n3348 3.1005
R8151 VSS.n3360 VSS.n3359 3.1005
R8152 VSS.n3366 VSS.n3365 3.1005
R8153 VSS.n3368 VSS.n3367 3.1005
R8154 VSS.n3374 VSS.n3373 3.1005
R8155 VSS.n1860 VSS.n1859 3.1005
R8156 VSS.n1868 VSS.n1867 3.1005
R8157 VSS.n1872 VSS.n1871 3.1005
R8158 VSS.n1882 VSS.n1881 3.1005
R8159 VSS.n1892 VSS.n1891 3.1005
R8160 VSS.n1902 VSS.n1901 3.1005
R8161 VSS.n1922 VSS.n1921 3.1005
R8162 VSS.n1932 VSS.n1931 3.1005
R8163 VSS.n1942 VSS.n1941 3.1005
R8164 VSS.n1964 VSS.n1963 3.1005
R8165 VSS.n1974 VSS.n1973 3.1005
R8166 VSS.n1984 VSS.n1983 3.1005
R8167 VSS.n2014 VSS.n2013 3.1005
R8168 VSS.n2037 VSS.n2036 3.1005
R8169 VSS.n2058 VSS.n2057 3.1005
R8170 VSS.n2089 VSS.n2088 3.1005
R8171 VSS.n2099 VSS.n2098 3.1005
R8172 VSS.n3065 VSS.n3064 3.1005
R8173 VSS.n3069 VSS.n3068 3.1005
R8174 VSS.n3071 VSS.n3070 3.1005
R8175 VSS.n2109 VSS.n2108 3.1005
R8176 VSS.n2068 VSS.n2067 3.1005
R8177 VSS.n2027 VSS.n2026 3.1005
R8178 VSS.n1994 VSS.n1993 3.1005
R8179 VSS.n1952 VSS.n1951 3.1005
R8180 VSS.n1912 VSS.n1911 3.1005
R8181 VSS.n1878 VSS.n1877 3.1005
R8182 VSS.n1864 VSS.n1863 3.1005
R8183 VSS.n1850 VSS.n1849 3.1005
R8184 VSS.n1238 VSS.n1237 3.1005
R8185 VSS.n1233 VSS.n1232 3.1005
R8186 VSS.n1229 VSS.n1228 3.1005
R8187 VSS.n1225 VSS.n1224 3.1005
R8188 VSS.n1221 VSS.n1220 3.1005
R8189 VSS.n1215 VSS.n1214 3.1005
R8190 VSS.n1211 VSS.n1210 3.1005
R8191 VSS.n1207 VSS.n1206 3.1005
R8192 VSS.n1203 VSS.n1202 3.1005
R8193 VSS.n1198 VSS.n1197 3.1005
R8194 VSS.n1194 VSS.n1193 3.1005
R8195 VSS.n1190 VSS.n1189 3.1005
R8196 VSS.n1186 VSS.n1185 3.1005
R8197 VSS.n1182 VSS.n1181 3.1005
R8198 VSS.n1176 VSS.n1175 3.1005
R8199 VSS.n1172 VSS.n1171 3.1005
R8200 VSS.n1168 VSS.n1167 3.1005
R8201 VSS.n1164 VSS.n1163 3.1005
R8202 VSS.n1159 VSS.n1158 3.1005
R8203 VSS.n1155 VSS.n1154 3.1005
R8204 VSS.n1150 VSS.n1149 3.1005
R8205 VSS.n1146 VSS.n137 3.1005
R8206 VSS.n1137 VSS.n1136 3.1005
R8207 VSS.n1132 VSS.n1131 3.1005
R8208 VSS.n1128 VSS.n1127 3.1005
R8209 VSS.n1124 VSS.n1123 3.1005
R8210 VSS.n1120 VSS.n1119 3.1005
R8211 VSS.n1114 VSS.n1113 3.1005
R8212 VSS.n1110 VSS.n1109 3.1005
R8213 VSS.n1106 VSS.n1105 3.1005
R8214 VSS.n1102 VSS.n1101 3.1005
R8215 VSS.n1097 VSS.n1096 3.1005
R8216 VSS.n1249 VSS.n1248 3.1005
R8217 VSS.n4124 VSS.n4123 3.1005
R8218 VSS.n3836 VSS.n3835 3.1005
R8219 VSS.n3828 VSS.n3827 3.1005
R8220 VSS.n3819 VSS.n3818 3.1005
R8221 VSS.n3815 VSS.n3814 3.1005
R8222 VSS.n3811 VSS.n3810 3.1005
R8223 VSS.n3807 VSS.n3806 3.1005
R8224 VSS.n3801 VSS.n3800 3.1005
R8225 VSS.n3797 VSS.n3796 3.1005
R8226 VSS.n3793 VSS.n3792 3.1005
R8227 VSS.n3789 VSS.n3788 3.1005
R8228 VSS.n3784 VSS.n3783 3.1005
R8229 VSS.n3780 VSS.n3779 3.1005
R8230 VSS.n3776 VSS.n3775 3.1005
R8231 VSS.n3772 VSS.n3771 3.1005
R8232 VSS.n3768 VSS.n3767 3.1005
R8233 VSS.n3762 VSS.n3761 3.1005
R8234 VSS.n3758 VSS.n3757 3.1005
R8235 VSS.n3754 VSS.n3753 3.1005
R8236 VSS.n3750 VSS.n3749 3.1005
R8237 VSS.n3740 VSS.n3739 3.1005
R8238 VSS.n3736 VSS.n3735 3.1005
R8239 VSS.n3726 VSS.n3725 3.1005
R8240 VSS.n3716 VSS.n3715 3.1005
R8241 VSS.n3714 VSS.n3713 3.1005
R8242 VSS.n3705 VSS.n3704 3.1005
R8243 VSS.n3701 VSS.n3700 3.1005
R8244 VSS.n3697 VSS.n3696 3.1005
R8245 VSS.n3693 VSS.n3692 3.1005
R8246 VSS.n3687 VSS.n3686 3.1005
R8247 VSS.n3683 VSS.n3682 3.1005
R8248 VSS.n3679 VSS.n3678 3.1005
R8249 VSS.n3675 VSS.n3674 3.1005
R8250 VSS.n3670 VSS.n3669 3.1005
R8251 VSS.n3666 VSS.n3665 3.1005
R8252 VSS.n3662 VSS.n3661 3.1005
R8253 VSS.n3658 VSS.n3657 3.1005
R8254 VSS.n3654 VSS.n3653 3.1005
R8255 VSS.n3648 VSS.n3647 3.1005
R8256 VSS.n3644 VSS.n3643 3.1005
R8257 VSS.n3640 VSS.n3639 3.1005
R8258 VSS.n3636 VSS.n3635 3.1005
R8259 VSS.n3626 VSS.n3625 3.1005
R8260 VSS.n3622 VSS.n3621 3.1005
R8261 VSS.n3612 VSS.n3611 3.1005
R8262 VSS.n3602 VSS.n3601 3.1005
R8263 VSS.n3600 VSS.n3599 3.1005
R8264 VSS.n3591 VSS.n3590 3.1005
R8265 VSS.n3587 VSS.n3586 3.1005
R8266 VSS.n3583 VSS.n3582 3.1005
R8267 VSS.n3579 VSS.n3578 3.1005
R8268 VSS.n3573 VSS.n3572 3.1005
R8269 VSS.n3569 VSS.n3568 3.1005
R8270 VSS.n3565 VSS.n3564 3.1005
R8271 VSS.n3561 VSS.n3560 3.1005
R8272 VSS.n3556 VSS.n3555 3.1005
R8273 VSS.n3552 VSS.n3551 3.1005
R8274 VSS.n3548 VSS.n3547 3.1005
R8275 VSS.n3544 VSS.n3543 3.1005
R8276 VSS.n3540 VSS.n3539 3.1005
R8277 VSS.n3534 VSS.n3533 3.1005
R8278 VSS.n3530 VSS.n3529 3.1005
R8279 VSS.n3526 VSS.n3525 3.1005
R8280 VSS.n3522 VSS.n3521 3.1005
R8281 VSS.n3512 VSS.n3511 3.1005
R8282 VSS.n3508 VSS.n3507 3.1005
R8283 VSS.n3498 VSS.n3497 3.1005
R8284 VSS.n3488 VSS.n3487 3.1005
R8285 VSS.n3486 VSS.n3485 3.1005
R8286 VSS.n3477 VSS.n3476 3.1005
R8287 VSS.n3473 VSS.n3472 3.1005
R8288 VSS.n3469 VSS.n3468 3.1005
R8289 VSS.n3465 VSS.n3464 3.1005
R8290 VSS.n3459 VSS.n3458 3.1005
R8291 VSS.n3455 VSS.n3454 3.1005
R8292 VSS.n3451 VSS.n3450 3.1005
R8293 VSS.n3447 VSS.n3446 3.1005
R8294 VSS.n3442 VSS.n3441 3.1005
R8295 VSS.n3438 VSS.n3437 3.1005
R8296 VSS.n3434 VSS.n3433 3.1005
R8297 VSS.n3430 VSS.n3429 3.1005
R8298 VSS.n3426 VSS.n3425 3.1005
R8299 VSS.n3420 VSS.n3419 3.1005
R8300 VSS.n3416 VSS.n3415 3.1005
R8301 VSS.n3412 VSS.n3411 3.1005
R8302 VSS.n3408 VSS.n3407 3.1005
R8303 VSS.n3398 VSS.n3397 3.1005
R8304 VSS.n3394 VSS.n3393 3.1005
R8305 VSS.n4238 VSS.n4237 3.1005
R8306 VSS.n4232 VSS.n0 3.1005
R8307 VSS.n4226 VSS.n4225 3.1005
R8308 VSS.n4217 VSS.n4216 3.1005
R8309 VSS.n4213 VSS.n4212 3.1005
R8310 VSS.n4209 VSS.n4208 3.1005
R8311 VSS.n4205 VSS.n4204 3.1005
R8312 VSS.n4199 VSS.n4198 3.1005
R8313 VSS.n4195 VSS.n4194 3.1005
R8314 VSS.n4191 VSS.n4190 3.1005
R8315 VSS.n4187 VSS.n4186 3.1005
R8316 VSS.n4182 VSS.n4181 3.1005
R8317 VSS.n4178 VSS.n4177 3.1005
R8318 VSS.n4174 VSS.n4173 3.1005
R8319 VSS.n4170 VSS.n4169 3.1005
R8320 VSS.n4166 VSS.n4165 3.1005
R8321 VSS.n4160 VSS.n4159 3.1005
R8322 VSS.n4156 VSS.n4155 3.1005
R8323 VSS.n4152 VSS.n4151 3.1005
R8324 VSS.n4148 VSS.n4147 3.1005
R8325 VSS.n4138 VSS.n4137 3.1005
R8326 VSS.n4134 VSS.n4133 3.1005
R8327 VSS.n4113 VSS.n4112 3.09016
R8328 VSS.n4093 VSS.n4086 3.09016
R8329 VSS.n4095 VSS.n4093 3.09016
R8330 VSS.n4079 VSS.n4073 3.09016
R8331 VSS.n4081 VSS.n4079 3.09016
R8332 VSS.n4065 VSS.n4063 3.09016
R8333 VSS.n4051 VSS.n4044 3.09016
R8334 VSS.n4053 VSS.n4051 3.09016
R8335 VSS.n4037 VSS.n4030 3.09016
R8336 VSS.n4039 VSS.n4037 3.09016
R8337 VSS.n4023 VSS.n4016 3.09016
R8338 VSS.n4025 VSS.n4023 3.09016
R8339 VSS.n36 VSS.n29 3.09016
R8340 VSS.n4008 VSS.n4006 3.09016
R8341 VSS.n3994 VSS.n3987 3.09016
R8342 VSS.n3996 VSS.n3994 3.09016
R8343 VSS.n3980 VSS.n3973 3.09016
R8344 VSS.n3982 VSS.n3980 3.09016
R8345 VSS.n3966 VSS.n3959 3.09016
R8346 VSS.n3968 VSS.n3966 3.09016
R8347 VSS.n3951 VSS.n3944 3.09016
R8348 VSS.n3954 VSS.n3951 3.09016
R8349 VSS.n3937 VSS.n3930 3.09016
R8350 VSS.n3939 VSS.n3937 3.09016
R8351 VSS.n3922 VSS.n3915 3.09016
R8352 VSS.n3925 VSS.n3922 3.09016
R8353 VSS.n3908 VSS.n3901 3.09016
R8354 VSS.n3910 VSS.n3908 3.09016
R8355 VSS.n50 VSS.n43 3.09016
R8356 VSS.n3896 VSS.n50 3.09016
R8357 VSS.n2075 VSS.n2074 2.99827
R8358 VSS.n2021 VSS.n2020 2.99827
R8359 VSS.n2001 VSS.n2000 2.8978
R8360 VSS.n26 VSS.n17 2.86947
R8361 VSS.n3048 VSS.n3047 2.7891
R8362 VSS.n2767 VSS.n2766 2.7891
R8363 VSS.n2697 VSS.n2696 2.7891
R8364 VSS.n2416 VSS.n2415 2.7891
R8365 VSS.n2346 VSS.n2345 2.7891
R8366 VSS.n151 VSS.n150 2.7891
R8367 VSS.n932 VSS.n931 2.7891
R8368 VSS.n205 VSS.n204 2.7891
R8369 VSS.n623 VSS.n622 2.7891
R8370 VSS.n259 VSS.n258 2.7891
R8371 VSS.n4115 VSS.n4105 2.7891
R8372 VSS.n27 VSS.n26 2.7891
R8373 VSS.n40 VSS.n39 2.7891
R8374 VSS.n1202 VSS.n1199 2.64878
R8375 VSS.n1101 VSS.n1098 2.64878
R8376 VSS.n1039 VSS.n1038 2.64878
R8377 VSS.n730 VSS.n729 2.64878
R8378 VSS.n421 VSS.n420 2.64878
R8379 VSS.n1784 VSS.n1781 2.64878
R8380 VSS.n1683 VSS.n1680 2.64878
R8381 VSS.n1582 VSS.n1579 2.64878
R8382 VSS.n1481 VSS.n1478 2.64878
R8383 VSS.n1380 VSS.n1377 2.64878
R8384 VSS.n4186 VSS.n4183 2.64878
R8385 VSS.n3446 VSS.n3443 2.64878
R8386 VSS.n3560 VSS.n3557 2.64878
R8387 VSS.n3674 VSS.n3671 2.64878
R8388 VSS.n3788 VSS.n3785 2.64878
R8389 VSS.n3021 VSS.n3020 2.63101
R8390 VSS.n2670 VSS.n2669 2.63101
R8391 VSS.n2319 VSS.n2318 2.63101
R8392 VSS.n195 VSS.n194 2.63101
R8393 VSS.n249 VSS.n248 2.63101
R8394 VSS.n2004 VSS.n2003 2.5203
R8395 VSS.n1133 VSS.n141 2.5203
R8396 VSS.n1234 VSS.n126 2.5203
R8397 VSS.n1412 VSS.n1314 2.5203
R8398 VSS.n1513 VSS.n1299 2.5203
R8399 VSS.n1614 VSS.n1284 2.5203
R8400 VSS.n1715 VSS.n1269 2.5203
R8401 VSS.n1816 VSS.n1254 2.5203
R8402 VSS.n3824 VSS.n3823 2.5203
R8403 VSS.n3710 VSS.n3709 2.5203
R8404 VSS.n3596 VSS.n3595 2.5203
R8405 VSS.n3482 VSS.n3481 2.5203
R8406 VSS.n4222 VSS.n4221 2.5203
R8407 VSS.n2025 VSS.n2024 2.49102
R8408 VSS.n2079 VSS.n2078 2.49102
R8409 VSS.n1856 VSS.n1855 2.49102
R8410 VSS.n3380 VSS.n3379 2.49102
R8411 VSS.n3356 VSS.n3355 2.49102
R8412 VSS.n1140 VSS.n1138 2.49102
R8413 VSS.n1160 VSS.n131 2.49102
R8414 VSS.n1242 VSS.n1239 2.49102
R8415 VSS.n3863 VSS.n3862 2.49102
R8416 VSS.n3849 VSS.n3848 2.49102
R8417 VSS.n1338 VSS.n1319 2.49102
R8418 VSS.n1419 VSS.n1417 2.49102
R8419 VSS.n1439 VSS.n1304 2.49102
R8420 VSS.n1520 VSS.n1518 2.49102
R8421 VSS.n1540 VSS.n1289 2.49102
R8422 VSS.n1621 VSS.n1619 2.49102
R8423 VSS.n1641 VSS.n1274 2.49102
R8424 VSS.n1722 VSS.n1720 2.49102
R8425 VSS.n1742 VSS.n1259 2.49102
R8426 VSS.n1823 VSS.n1821 2.49102
R8427 VSS.n3834 VSS.n3833 2.49102
R8428 VSS.n3746 VSS.n3745 2.49102
R8429 VSS.n3718 VSS.n3717 2.49102
R8430 VSS.n3632 VSS.n3631 2.49102
R8431 VSS.n3604 VSS.n3603 2.49102
R8432 VSS.n3518 VSS.n3517 2.49102
R8433 VSS.n3490 VSS.n3489 2.49102
R8434 VSS.n3404 VSS.n3403 2.49102
R8435 VSS.n4228 VSS.n4227 2.49102
R8436 VSS.n4144 VSS.n4143 2.49102
R8437 VSS.n2048 VSS.n2047 2.43201
R8438 VSS.n1842 VSS.n1841 2.43201
R8439 VSS.n1151 VSS.n136 2.43201
R8440 VSS.n1329 VSS.n1324 2.43201
R8441 VSS.n1430 VSS.n1309 2.43201
R8442 VSS.n1531 VSS.n1294 2.43201
R8443 VSS.n1632 VSS.n1279 2.43201
R8444 VSS.n1733 VSS.n1264 2.43201
R8445 VSS.n3732 VSS.n3731 2.43201
R8446 VSS.n3618 VSS.n3617 2.43201
R8447 VSS.n3504 VSS.n3503 2.43201
R8448 VSS.n6 VSS.n5 2.43201
R8449 VSS.n4130 VSS.n4129 2.43201
R8450 VSS VSS.n181 2.42809
R8451 VSS VSS.n235 2.42809
R8452 VSS.n3053 VSS.n83 2.38818
R8453 VSS.n83 VSS 2.2358
R8454 VSS.n3057 VSS.n75 2.2074
R8455 VSS.n3033 VSS.n3026 2.2074
R8456 VSS.n2921 VSS.n2914 2.2074
R8457 VSS.n2935 VSS.n2928 2.2074
R8458 VSS.n2949 VSS.n2942 2.2074
R8459 VSS.n2965 VSS.n2958 2.2074
R8460 VSS.n2979 VSS.n2972 2.2074
R8461 VSS.n2993 VSS.n2986 2.2074
R8462 VSS.n3007 VSS.n3000 2.2074
R8463 VSS.n2779 VSS.n2772 2.2074
R8464 VSS.n2793 VSS.n2786 2.2074
R8465 VSS.n2807 VSS.n2800 2.2074
R8466 VSS.n2821 VSS.n2814 2.2074
R8467 VSS.n2835 VSS.n2828 2.2074
R8468 VSS.n2851 VSS.n2844 2.2074
R8469 VSS.n2865 VSS.n2858 2.2074
R8470 VSS.n2879 VSS.n2872 2.2074
R8471 VSS.n2893 VSS.n2886 2.2074
R8472 VSS.n2738 VSS.n2731 2.2074
R8473 VSS.n2752 VSS.n2745 2.2074
R8474 VSS.n2704 VSS.n100 2.2074
R8475 VSS.n2711 VSS.n92 2.2074
R8476 VSS.n2682 VSS.n2675 2.2074
R8477 VSS.n2570 VSS.n2563 2.2074
R8478 VSS.n2584 VSS.n2577 2.2074
R8479 VSS.n2598 VSS.n2591 2.2074
R8480 VSS.n2614 VSS.n2607 2.2074
R8481 VSS.n2628 VSS.n2621 2.2074
R8482 VSS.n2642 VSS.n2635 2.2074
R8483 VSS.n2656 VSS.n2649 2.2074
R8484 VSS.n2428 VSS.n2421 2.2074
R8485 VSS.n2442 VSS.n2435 2.2074
R8486 VSS.n2456 VSS.n2449 2.2074
R8487 VSS.n2470 VSS.n2463 2.2074
R8488 VSS.n2484 VSS.n2477 2.2074
R8489 VSS.n2500 VSS.n2493 2.2074
R8490 VSS.n2514 VSS.n2507 2.2074
R8491 VSS.n2528 VSS.n2521 2.2074
R8492 VSS.n2542 VSS.n2535 2.2074
R8493 VSS.n2387 VSS.n2380 2.2074
R8494 VSS.n2401 VSS.n2394 2.2074
R8495 VSS.n2353 VSS.n112 2.2074
R8496 VSS.n2360 VSS.n104 2.2074
R8497 VSS.n2331 VSS.n2324 2.2074
R8498 VSS.n2219 VSS.n2212 2.2074
R8499 VSS.n2233 VSS.n2226 2.2074
R8500 VSS.n2247 VSS.n2240 2.2074
R8501 VSS.n2263 VSS.n2256 2.2074
R8502 VSS.n2277 VSS.n2270 2.2074
R8503 VSS.n2291 VSS.n2284 2.2074
R8504 VSS.n2305 VSS.n2298 2.2074
R8505 VSS.n2119 VSS.n2112 2.2074
R8506 VSS.n2133 VSS.n2126 2.2074
R8507 VSS.n2149 VSS.n2142 2.2074
R8508 VSS.n2163 VSS.n2156 2.2074
R8509 VSS.n2177 VSS.n2170 2.2074
R8510 VSS.n2191 VSS.n2184 2.2074
R8511 VSS.n1089 VSS.n1082 2.2074
R8512 VSS.n1091 VSS.n1089 2.2074
R8513 VSS.n1075 VSS.n1068 2.2074
R8514 VSS.n1077 VSS.n1075 2.2074
R8515 VSS.n1061 VSS.n1054 2.2074
R8516 VSS.n1063 VSS.n1061 2.2074
R8517 VSS.n1047 VSS.n1040 2.2074
R8518 VSS.n1049 VSS.n1047 2.2074
R8519 VSS.n1031 VSS.n1024 2.2074
R8520 VSS.n1033 VSS.n1031 2.2074
R8521 VSS.n1017 VSS.n1010 2.2074
R8522 VSS.n1019 VSS.n1017 2.2074
R8523 VSS.n1003 VSS.n996 2.2074
R8524 VSS.n1005 VSS.n1003 2.2074
R8525 VSS.n989 VSS.n982 2.2074
R8526 VSS.n991 VSS.n989 2.2074
R8527 VSS.n972 VSS.n965 2.2074
R8528 VSS.n974 VSS.n972 2.2074
R8529 VSS.n958 VSS.n951 2.2074
R8530 VSS.n960 VSS.n958 2.2074
R8531 VSS.n172 VSS.n165 2.2074
R8532 VSS.n943 VSS.n172 2.2074
R8533 VSS.n940 VSS.n939 2.2074
R8534 VSS.n939 VSS.n173 2.2074
R8535 VSS.n924 VSS.n917 2.2074
R8536 VSS.n926 VSS.n924 2.2074
R8537 VSS.n907 VSS.n900 2.2074
R8538 VSS.n909 VSS.n907 2.2074
R8539 VSS.n893 VSS.n886 2.2074
R8540 VSS.n895 VSS.n893 2.2074
R8541 VSS.n879 VSS.n872 2.2074
R8542 VSS.n881 VSS.n879 2.2074
R8543 VSS.n863 VSS.n857 2.2074
R8544 VSS.n867 VSS.n863 2.2074
R8545 VSS.n850 VSS.n843 2.2074
R8546 VSS.n852 VSS.n850 2.2074
R8547 VSS.n836 VSS.n829 2.2074
R8548 VSS.n838 VSS.n836 2.2074
R8549 VSS.n822 VSS.n815 2.2074
R8550 VSS.n824 VSS.n822 2.2074
R8551 VSS.n807 VSS.n800 2.2074
R8552 VSS.n810 VSS.n807 2.2074
R8553 VSS.n795 VSS.n793 2.2074
R8554 VSS.n780 VSS.n773 2.2074
R8555 VSS.n782 VSS.n780 2.2074
R8556 VSS.n766 VSS.n759 2.2074
R8557 VSS.n768 VSS.n766 2.2074
R8558 VSS.n752 VSS.n745 2.2074
R8559 VSS.n754 VSS.n752 2.2074
R8560 VSS.n738 VSS.n731 2.2074
R8561 VSS.n740 VSS.n738 2.2074
R8562 VSS.n722 VSS.n715 2.2074
R8563 VSS.n724 VSS.n722 2.2074
R8564 VSS.n708 VSS.n701 2.2074
R8565 VSS.n710 VSS.n708 2.2074
R8566 VSS.n694 VSS.n687 2.2074
R8567 VSS.n696 VSS.n694 2.2074
R8568 VSS.n680 VSS.n673 2.2074
R8569 VSS.n682 VSS.n680 2.2074
R8570 VSS.n663 VSS.n656 2.2074
R8571 VSS.n665 VSS.n663 2.2074
R8572 VSS.n649 VSS.n642 2.2074
R8573 VSS.n651 VSS.n649 2.2074
R8574 VSS.n226 VSS.n219 2.2074
R8575 VSS.n634 VSS.n226 2.2074
R8576 VSS.n631 VSS.n630 2.2074
R8577 VSS.n630 VSS.n227 2.2074
R8578 VSS.n615 VSS.n608 2.2074
R8579 VSS.n617 VSS.n615 2.2074
R8580 VSS.n598 VSS.n591 2.2074
R8581 VSS.n600 VSS.n598 2.2074
R8582 VSS.n584 VSS.n577 2.2074
R8583 VSS.n586 VSS.n584 2.2074
R8584 VSS.n570 VSS.n563 2.2074
R8585 VSS.n572 VSS.n570 2.2074
R8586 VSS.n554 VSS.n548 2.2074
R8587 VSS.n558 VSS.n554 2.2074
R8588 VSS.n541 VSS.n534 2.2074
R8589 VSS.n543 VSS.n541 2.2074
R8590 VSS.n527 VSS.n520 2.2074
R8591 VSS.n529 VSS.n527 2.2074
R8592 VSS.n513 VSS.n506 2.2074
R8593 VSS.n515 VSS.n513 2.2074
R8594 VSS.n498 VSS.n491 2.2074
R8595 VSS.n501 VSS.n498 2.2074
R8596 VSS.n486 VSS.n484 2.2074
R8597 VSS.n471 VSS.n464 2.2074
R8598 VSS.n473 VSS.n471 2.2074
R8599 VSS.n457 VSS.n450 2.2074
R8600 VSS.n459 VSS.n457 2.2074
R8601 VSS.n443 VSS.n436 2.2074
R8602 VSS.n445 VSS.n443 2.2074
R8603 VSS.n429 VSS.n422 2.2074
R8604 VSS.n431 VSS.n429 2.2074
R8605 VSS.n413 VSS.n406 2.2074
R8606 VSS.n415 VSS.n413 2.2074
R8607 VSS.n399 VSS.n392 2.2074
R8608 VSS.n401 VSS.n399 2.2074
R8609 VSS.n385 VSS.n378 2.2074
R8610 VSS.n387 VSS.n385 2.2074
R8611 VSS.n371 VSS.n364 2.2074
R8612 VSS.n373 VSS.n371 2.2074
R8613 VSS.n354 VSS.n347 2.2074
R8614 VSS.n356 VSS.n354 2.2074
R8615 VSS.n340 VSS.n333 2.2074
R8616 VSS.n342 VSS.n340 2.2074
R8617 VSS.n280 VSS.n273 2.2074
R8618 VSS.n325 VSS.n280 2.2074
R8619 VSS.n322 VSS.n321 2.2074
R8620 VSS.n321 VSS.n314 2.2074
R8621 VSS.n309 VSS.n307 2.2074
R8622 VSS.n293 VSS.n286 2.2074
R8623 VSS.n295 VSS.n293 2.2074
R8624 VSS.n3078 VSS.n67 2.2074
R8625 VSS.n3080 VSS.n3078 2.2074
R8626 VSS.n3092 VSS.n3085 2.2074
R8627 VSS.n3096 VSS.n3092 2.2074
R8628 VSS.n3108 VSS.n3101 2.2074
R8629 VSS.n3110 VSS.n3108 2.2074
R8630 VSS.n3122 VSS.n3115 2.2074
R8631 VSS.n3126 VSS.n3122 2.2074
R8632 VSS.n3137 VSS.n3131 2.2074
R8633 VSS.n3139 VSS.n3137 2.2074
R8634 VSS.n3151 VSS.n3144 2.2074
R8635 VSS.n3155 VSS.n3151 2.2074
R8636 VSS.n3167 VSS.n3160 2.2074
R8637 VSS.n3169 VSS.n3167 2.2074
R8638 VSS.n3182 VSS.n3175 2.2074
R8639 VSS.n3197 VSS.n3190 2.2074
R8640 VSS.n3199 VSS.n3197 2.2074
R8641 VSS.n3215 VSS.n3213 2.2074
R8642 VSS.n3227 VSS.n3220 2.2074
R8643 VSS.n3229 VSS.n3227 2.2074
R8644 VSS.n3243 VSS.n3236 2.2074
R8645 VSS.n3245 VSS.n3243 2.2074
R8646 VSS.n3257 VSS.n3250 2.2074
R8647 VSS.n3261 VSS.n3257 2.2074
R8648 VSS.n3273 VSS.n3266 2.2074
R8649 VSS.n3275 VSS.n3273 2.2074
R8650 VSS.n3287 VSS.n3280 2.2074
R8651 VSS.n3291 VSS.n3287 2.2074
R8652 VSS.n3303 VSS.n3296 2.2074
R8653 VSS.n3305 VSS.n3303 2.2074
R8654 VSS.n3317 VSS.n3310 2.2074
R8655 VSS.n3321 VSS.n3317 2.2074
R8656 VSS.n3333 VSS.n3326 2.2074
R8657 VSS.n3335 VSS.n3333 2.2074
R8658 VSS.n3343 VSS.n62 2.2074
R8659 VSS.n26 VSS.n25 2.2074
R8660 VSS.n3057 VSS.n3056 1.98671
R8661 VSS.n3035 VSS.n3033 1.98671
R8662 VSS.n2909 VSS.n2907 1.98671
R8663 VSS.n2923 VSS.n2921 1.98671
R8664 VSS.n2937 VSS.n2935 1.98671
R8665 VSS.n2951 VSS.n2949 1.98671
R8666 VSS.n2967 VSS.n2965 1.98671
R8667 VSS.n2981 VSS.n2979 1.98671
R8668 VSS.n2995 VSS.n2993 1.98671
R8669 VSS.n3009 VSS.n3007 1.98671
R8670 VSS.n2781 VSS.n2779 1.98671
R8671 VSS.n2795 VSS.n2793 1.98671
R8672 VSS.n2809 VSS.n2807 1.98671
R8673 VSS.n2823 VSS.n2821 1.98671
R8674 VSS.n2839 VSS.n2835 1.98671
R8675 VSS.n2853 VSS.n2851 1.98671
R8676 VSS.n2867 VSS.n2865 1.98671
R8677 VSS.n2881 VSS.n2879 1.98671
R8678 VSS.n2895 VSS.n2893 1.98671
R8679 VSS.n2740 VSS.n2738 1.98671
R8680 VSS.n2754 VSS.n2752 1.98671
R8681 VSS.n2704 VSS.n2703 1.98671
R8682 VSS.n2713 VSS.n2711 1.98671
R8683 VSS.n2684 VSS.n2682 1.98671
R8684 VSS.n2558 VSS.n2556 1.98671
R8685 VSS.n2572 VSS.n2570 1.98671
R8686 VSS.n2586 VSS.n2584 1.98671
R8687 VSS.n2600 VSS.n2598 1.98671
R8688 VSS.n2616 VSS.n2614 1.98671
R8689 VSS.n2630 VSS.n2628 1.98671
R8690 VSS.n2644 VSS.n2642 1.98671
R8691 VSS.n2658 VSS.n2656 1.98671
R8692 VSS.n2430 VSS.n2428 1.98671
R8693 VSS.n2444 VSS.n2442 1.98671
R8694 VSS.n2458 VSS.n2456 1.98671
R8695 VSS.n2472 VSS.n2470 1.98671
R8696 VSS.n2488 VSS.n2484 1.98671
R8697 VSS.n2502 VSS.n2500 1.98671
R8698 VSS.n2516 VSS.n2514 1.98671
R8699 VSS.n2530 VSS.n2528 1.98671
R8700 VSS.n2544 VSS.n2542 1.98671
R8701 VSS.n2389 VSS.n2387 1.98671
R8702 VSS.n2403 VSS.n2401 1.98671
R8703 VSS.n2353 VSS.n2352 1.98671
R8704 VSS.n2362 VSS.n2360 1.98671
R8705 VSS.n2333 VSS.n2331 1.98671
R8706 VSS.n2207 VSS.n2205 1.98671
R8707 VSS.n2221 VSS.n2219 1.98671
R8708 VSS.n2235 VSS.n2233 1.98671
R8709 VSS.n2249 VSS.n2247 1.98671
R8710 VSS.n2265 VSS.n2263 1.98671
R8711 VSS.n2279 VSS.n2277 1.98671
R8712 VSS.n2293 VSS.n2291 1.98671
R8713 VSS.n2307 VSS.n2305 1.98671
R8714 VSS.n2088 VSS.n2085 1.98671
R8715 VSS.n2098 VSS.n2095 1.98671
R8716 VSS.n2108 VSS.n2105 1.98671
R8717 VSS.n2121 VSS.n2119 1.98671
R8718 VSS.n2137 VSS.n2133 1.98671
R8719 VSS.n2151 VSS.n2149 1.98671
R8720 VSS.n2165 VSS.n2163 1.98671
R8721 VSS.n2179 VSS.n2177 1.98671
R8722 VSS.n2193 VSS.n2191 1.98671
R8723 VSS.n2057 VSS.n2054 1.98671
R8724 VSS.n2067 VSS.n2064 1.98671
R8725 VSS.n2027 VSS.n122 1.98671
R8726 VSS.n2036 VSS.n2033 1.98671
R8727 VSS.n2013 VSS.n2010 1.98671
R8728 VSS.n1921 VSS.n1918 1.98671
R8729 VSS.n1931 VSS.n1928 1.98671
R8730 VSS.n1941 VSS.n1938 1.98671
R8731 VSS.n1951 VSS.n1948 1.98671
R8732 VSS.n1963 VSS.n1960 1.98671
R8733 VSS.n1973 VSS.n1970 1.98671
R8734 VSS.n1983 VSS.n1980 1.98671
R8735 VSS.n1993 VSS.n1990 1.98671
R8736 VSS.n1891 VSS.n1888 1.98671
R8737 VSS.n1901 VSS.n1898 1.98671
R8738 VSS.n1911 VSS.n1908 1.98671
R8739 VSS.n3365 VSS.n3362 1.98671
R8740 VSS.n78 VSS.n77 1.9836
R8741 VSS.n88 VSS.n87 1.87367
R8742 VSS.n3056 VSS.n76 1.76602
R8743 VSS.n76 VSS 1.76602
R8744 VSS.n3035 VSS.n3034 1.76602
R8745 VSS.n2909 VSS.n2908 1.76602
R8746 VSS.n2923 VSS.n2922 1.76602
R8747 VSS.n2937 VSS.n2936 1.76602
R8748 VSS.n2951 VSS.n2950 1.76602
R8749 VSS.n2967 VSS.n2966 1.76602
R8750 VSS.n2981 VSS.n2980 1.76602
R8751 VSS.n2995 VSS.n2994 1.76602
R8752 VSS.n3009 VSS.n3008 1.76602
R8753 VSS.n2781 VSS.n2780 1.76602
R8754 VSS.n2795 VSS.n2794 1.76602
R8755 VSS.n2809 VSS.n2808 1.76602
R8756 VSS.n2823 VSS.n2822 1.76602
R8757 VSS.n2839 VSS.n2838 1.76602
R8758 VSS.n2853 VSS.n2852 1.76602
R8759 VSS.n2867 VSS.n2866 1.76602
R8760 VSS.n2881 VSS.n2880 1.76602
R8761 VSS.n2895 VSS.n2894 1.76602
R8762 VSS.n2740 VSS.n2739 1.76602
R8763 VSS.n2754 VSS.n2753 1.76602
R8764 VSS.n2703 VSS.n102 1.76602
R8765 VSS.n102 VSS 1.76602
R8766 VSS.n2713 VSS.n2712 1.76602
R8767 VSS.n2684 VSS.n2683 1.76602
R8768 VSS.n2558 VSS.n2557 1.76602
R8769 VSS.n2572 VSS.n2571 1.76602
R8770 VSS.n2586 VSS.n2585 1.76602
R8771 VSS.n2600 VSS.n2599 1.76602
R8772 VSS.n2616 VSS.n2615 1.76602
R8773 VSS.n2630 VSS.n2629 1.76602
R8774 VSS.n2644 VSS.n2643 1.76602
R8775 VSS.n2658 VSS.n2657 1.76602
R8776 VSS.n2430 VSS.n2429 1.76602
R8777 VSS.n2444 VSS.n2443 1.76602
R8778 VSS.n2458 VSS.n2457 1.76602
R8779 VSS.n2472 VSS.n2471 1.76602
R8780 VSS.n2488 VSS.n2487 1.76602
R8781 VSS.n2502 VSS.n2501 1.76602
R8782 VSS.n2516 VSS.n2515 1.76602
R8783 VSS.n2530 VSS.n2529 1.76602
R8784 VSS.n2544 VSS.n2543 1.76602
R8785 VSS.n2389 VSS.n2388 1.76602
R8786 VSS.n2403 VSS.n2402 1.76602
R8787 VSS.n2352 VSS.n114 1.76602
R8788 VSS.n114 VSS 1.76602
R8789 VSS.n2362 VSS.n2361 1.76602
R8790 VSS.n2333 VSS.n2332 1.76602
R8791 VSS.n2207 VSS.n2206 1.76602
R8792 VSS.n2221 VSS.n2220 1.76602
R8793 VSS.n2235 VSS.n2234 1.76602
R8794 VSS.n2249 VSS.n2248 1.76602
R8795 VSS.n2265 VSS.n2264 1.76602
R8796 VSS.n2279 VSS.n2278 1.76602
R8797 VSS.n2293 VSS.n2292 1.76602
R8798 VSS.n2307 VSS.n2306 1.76602
R8799 VSS.n2121 VSS.n2120 1.76602
R8800 VSS.n2137 VSS.n2136 1.76602
R8801 VSS.n2151 VSS.n2150 1.76602
R8802 VSS.n2165 VSS.n2164 1.76602
R8803 VSS.n2179 VSS.n2178 1.76602
R8804 VSS.n2193 VSS.n2192 1.76602
R8805 VSS.n3183 VSS.n3182 1.76602
R8806 VSS.n3213 VSS.n3206 1.76602
R8807 VSS.n39 VSS.n36 1.76602
R8808 VSS.n1841 VSS.n1839 1.72554
R8809 VSS.n1264 VSS.n1262 1.72554
R8810 VSS.n1279 VSS.n1277 1.72554
R8811 VSS.n1294 VSS.n1292 1.72554
R8812 VSS.n1309 VSS.n1307 1.72554
R8813 VSS.n1324 VSS.n1322 1.72554
R8814 VSS.n2047 VSS.n2045 1.72554
R8815 VSS.n136 VSS.n134 1.72554
R8816 VSS.n3731 VSS.n3729 1.72554
R8817 VSS.n3617 VSS.n3615 1.72554
R8818 VSS.n3503 VSS.n3501 1.72554
R8819 VSS.n5 VSS.n3 1.72554
R8820 VSS.n4129 VSS.n4127 1.72554
R8821 VSS.n3848 VSS.n3846 1.57241
R8822 VSS.n3862 VSS.n3860 1.57241
R8823 VSS.n1824 VSS.n1823 1.57241
R8824 VSS.n1259 VSS.n1257 1.57241
R8825 VSS.n1723 VSS.n1722 1.57241
R8826 VSS.n1274 VSS.n1272 1.57241
R8827 VSS.n1622 VSS.n1621 1.57241
R8828 VSS.n1289 VSS.n1287 1.57241
R8829 VSS.n1521 VSS.n1520 1.57241
R8830 VSS.n1304 VSS.n1302 1.57241
R8831 VSS.n1420 VSS.n1419 1.57241
R8832 VSS.n1319 VSS.n1317 1.57241
R8833 VSS.n3355 VSS.n3353 1.57241
R8834 VSS.n3379 VSS.n3377 1.57241
R8835 VSS.n1855 VSS.n1853 1.57241
R8836 VSS.n2024 VSS.n2022 1.57241
R8837 VSS.n2078 VSS.n2076 1.57241
R8838 VSS.n1243 VSS.n1242 1.57241
R8839 VSS.n131 VSS.n129 1.57241
R8840 VSS.n1141 VSS.n1140 1.57241
R8841 VSS.n4143 VSS.n4141 1.57241
R8842 VSS.n4229 VSS.n4228 1.57241
R8843 VSS.n3403 VSS.n3401 1.57241
R8844 VSS.n3491 VSS.n3490 1.57241
R8845 VSS.n3517 VSS.n3515 1.57241
R8846 VSS.n3605 VSS.n3604 1.57241
R8847 VSS.n3631 VSS.n3629 1.57241
R8848 VSS.n3719 VSS.n3718 1.57241
R8849 VSS.n3745 VSS.n3743 1.57241
R8850 VSS.n3833 VSS.n3831 1.57241
R8851 VSS.n75 VSS.n74 1.54533
R8852 VSS.n3026 VSS.n3025 1.54533
R8853 VSS.n2914 VSS.n2913 1.54533
R8854 VSS.n2928 VSS.n2927 1.54533
R8855 VSS.n2942 VSS.n2941 1.54533
R8856 VSS.n2958 VSS.n2957 1.54533
R8857 VSS.n2972 VSS.n2971 1.54533
R8858 VSS.n2986 VSS.n2985 1.54533
R8859 VSS.n3000 VSS.n2999 1.54533
R8860 VSS.n2772 VSS.n2771 1.54533
R8861 VSS.n2786 VSS.n2785 1.54533
R8862 VSS.n2800 VSS.n2799 1.54533
R8863 VSS.n2814 VSS.n2813 1.54533
R8864 VSS.n2828 VSS.n2827 1.54533
R8865 VSS.n2844 VSS.n2843 1.54533
R8866 VSS.n2858 VSS.n2857 1.54533
R8867 VSS.n2872 VSS.n2871 1.54533
R8868 VSS.n2886 VSS.n2885 1.54533
R8869 VSS.n2731 VSS.n2730 1.54533
R8870 VSS.n2745 VSS.n2744 1.54533
R8871 VSS.n100 VSS.n99 1.54533
R8872 VSS.n101 VSS.n92 1.54533
R8873 VSS.n2675 VSS.n2674 1.54533
R8874 VSS.n2563 VSS.n2562 1.54533
R8875 VSS.n2577 VSS.n2576 1.54533
R8876 VSS.n2591 VSS.n2590 1.54533
R8877 VSS.n2607 VSS.n2606 1.54533
R8878 VSS.n2621 VSS.n2620 1.54533
R8879 VSS.n2635 VSS.n2634 1.54533
R8880 VSS.n2649 VSS.n2648 1.54533
R8881 VSS.n2421 VSS.n2420 1.54533
R8882 VSS.n2435 VSS.n2434 1.54533
R8883 VSS.n2449 VSS.n2448 1.54533
R8884 VSS.n2463 VSS.n2462 1.54533
R8885 VSS.n2477 VSS.n2476 1.54533
R8886 VSS.n2493 VSS.n2492 1.54533
R8887 VSS.n2507 VSS.n2506 1.54533
R8888 VSS.n2521 VSS.n2520 1.54533
R8889 VSS.n2535 VSS.n2534 1.54533
R8890 VSS.n2380 VSS.n2379 1.54533
R8891 VSS.n2394 VSS.n2393 1.54533
R8892 VSS.n112 VSS.n111 1.54533
R8893 VSS.n113 VSS.n104 1.54533
R8894 VSS.n2324 VSS.n2323 1.54533
R8895 VSS.n2212 VSS.n2211 1.54533
R8896 VSS.n2226 VSS.n2225 1.54533
R8897 VSS.n2240 VSS.n2239 1.54533
R8898 VSS.n2256 VSS.n2255 1.54533
R8899 VSS.n2270 VSS.n2269 1.54533
R8900 VSS.n2284 VSS.n2283 1.54533
R8901 VSS.n2298 VSS.n2297 1.54533
R8902 VSS.n2112 VSS.n2111 1.54533
R8903 VSS.n2126 VSS.n2125 1.54533
R8904 VSS.n2142 VSS.n2141 1.54533
R8905 VSS.n2156 VSS.n2155 1.54533
R8906 VSS.n2170 VSS.n2169 1.54533
R8907 VSS.n2184 VSS.n2183 1.54533
R8908 VSS.n1082 VSS.n1081 1.54533
R8909 VSS.n1091 VSS.n1090 1.54533
R8910 VSS.n1068 VSS.n1067 1.54533
R8911 VSS.n1077 VSS.n1076 1.54533
R8912 VSS.n1054 VSS.n1053 1.54533
R8913 VSS.n1063 VSS.n1062 1.54533
R8914 VSS.n1040 VSS.n1039 1.54533
R8915 VSS.n1049 VSS.n1048 1.54533
R8916 VSS.n1024 VSS.n1023 1.54533
R8917 VSS.n1033 VSS.n1032 1.54533
R8918 VSS.n1010 VSS.n1009 1.54533
R8919 VSS.n1019 VSS.n1018 1.54533
R8920 VSS.n996 VSS.n995 1.54533
R8921 VSS.n1005 VSS.n1004 1.54533
R8922 VSS.n982 VSS.n981 1.54533
R8923 VSS.n991 VSS.n990 1.54533
R8924 VSS.n965 VSS.n964 1.54533
R8925 VSS.n974 VSS.n973 1.54533
R8926 VSS.n951 VSS.n950 1.54533
R8927 VSS.n960 VSS.n959 1.54533
R8928 VSS.n165 VSS.n164 1.54533
R8929 VSS.n943 VSS.n942 1.54533
R8930 VSS.n941 VSS.n940 1.54533
R8931 VSS.n181 VSS.n173 1.54533
R8932 VSS.n917 VSS.n916 1.54533
R8933 VSS.n926 VSS.n925 1.54533
R8934 VSS.n900 VSS.n899 1.54533
R8935 VSS.n909 VSS.n908 1.54533
R8936 VSS.n886 VSS.n885 1.54533
R8937 VSS.n895 VSS.n894 1.54533
R8938 VSS.n872 VSS.n871 1.54533
R8939 VSS.n881 VSS.n880 1.54533
R8940 VSS.n857 VSS.n856 1.54533
R8941 VSS.n867 VSS.n866 1.54533
R8942 VSS.n843 VSS.n842 1.54533
R8943 VSS.n852 VSS.n851 1.54533
R8944 VSS.n829 VSS.n828 1.54533
R8945 VSS.n838 VSS.n837 1.54533
R8946 VSS.n815 VSS.n814 1.54533
R8947 VSS.n824 VSS.n823 1.54533
R8948 VSS.n800 VSS.n799 1.54533
R8949 VSS.n810 VSS.n809 1.54533
R8950 VSS.n795 VSS.n794 1.54533
R8951 VSS.n773 VSS.n772 1.54533
R8952 VSS.n782 VSS.n781 1.54533
R8953 VSS.n759 VSS.n758 1.54533
R8954 VSS.n768 VSS.n767 1.54533
R8955 VSS.n745 VSS.n744 1.54533
R8956 VSS.n754 VSS.n753 1.54533
R8957 VSS.n731 VSS.n730 1.54533
R8958 VSS.n740 VSS.n739 1.54533
R8959 VSS.n715 VSS.n714 1.54533
R8960 VSS.n724 VSS.n723 1.54533
R8961 VSS.n701 VSS.n700 1.54533
R8962 VSS.n710 VSS.n709 1.54533
R8963 VSS.n687 VSS.n686 1.54533
R8964 VSS.n696 VSS.n695 1.54533
R8965 VSS.n673 VSS.n672 1.54533
R8966 VSS.n682 VSS.n681 1.54533
R8967 VSS.n656 VSS.n655 1.54533
R8968 VSS.n665 VSS.n664 1.54533
R8969 VSS.n642 VSS.n641 1.54533
R8970 VSS.n651 VSS.n650 1.54533
R8971 VSS.n219 VSS.n218 1.54533
R8972 VSS.n634 VSS.n633 1.54533
R8973 VSS.n632 VSS.n631 1.54533
R8974 VSS.n235 VSS.n227 1.54533
R8975 VSS.n608 VSS.n607 1.54533
R8976 VSS.n617 VSS.n616 1.54533
R8977 VSS.n591 VSS.n590 1.54533
R8978 VSS.n600 VSS.n599 1.54533
R8979 VSS.n577 VSS.n576 1.54533
R8980 VSS.n586 VSS.n585 1.54533
R8981 VSS.n563 VSS.n562 1.54533
R8982 VSS.n572 VSS.n571 1.54533
R8983 VSS.n548 VSS.n547 1.54533
R8984 VSS.n558 VSS.n557 1.54533
R8985 VSS.n534 VSS.n533 1.54533
R8986 VSS.n543 VSS.n542 1.54533
R8987 VSS.n520 VSS.n519 1.54533
R8988 VSS.n529 VSS.n528 1.54533
R8989 VSS.n506 VSS.n505 1.54533
R8990 VSS.n515 VSS.n514 1.54533
R8991 VSS.n491 VSS.n490 1.54533
R8992 VSS.n501 VSS.n500 1.54533
R8993 VSS.n486 VSS.n485 1.54533
R8994 VSS.n464 VSS.n463 1.54533
R8995 VSS.n473 VSS.n472 1.54533
R8996 VSS.n450 VSS.n449 1.54533
R8997 VSS.n459 VSS.n458 1.54533
R8998 VSS.n436 VSS.n435 1.54533
R8999 VSS.n445 VSS.n444 1.54533
R9000 VSS.n422 VSS.n421 1.54533
R9001 VSS.n431 VSS.n430 1.54533
R9002 VSS.n406 VSS.n405 1.54533
R9003 VSS.n415 VSS.n414 1.54533
R9004 VSS.n392 VSS.n391 1.54533
R9005 VSS.n401 VSS.n400 1.54533
R9006 VSS.n378 VSS.n377 1.54533
R9007 VSS.n387 VSS.n386 1.54533
R9008 VSS.n364 VSS.n363 1.54533
R9009 VSS.n373 VSS.n372 1.54533
R9010 VSS.n347 VSS.n346 1.54533
R9011 VSS.n356 VSS.n355 1.54533
R9012 VSS.n333 VSS.n332 1.54533
R9013 VSS.n342 VSS.n341 1.54533
R9014 VSS.n273 VSS.n272 1.54533
R9015 VSS.n325 VSS.n324 1.54533
R9016 VSS.n323 VSS.n322 1.54533
R9017 VSS.n314 VSS.n282 1.54533
R9018 VSS.n309 VSS.n308 1.54533
R9019 VSS.n286 VSS.n285 1.54533
R9020 VSS.n295 VSS.n294 1.54533
R9021 VSS.n67 VSS.n66 1.54533
R9022 VSS.n3080 VSS.n3079 1.54533
R9023 VSS.n3085 VSS.n3084 1.54533
R9024 VSS.n3096 VSS.n3095 1.54533
R9025 VSS.n3101 VSS.n3100 1.54533
R9026 VSS.n3110 VSS.n3109 1.54533
R9027 VSS.n3115 VSS.n3114 1.54533
R9028 VSS.n3126 VSS.n3125 1.54533
R9029 VSS.n3131 VSS.n3130 1.54533
R9030 VSS.n3139 VSS.n3138 1.54533
R9031 VSS.n3144 VSS.n3143 1.54533
R9032 VSS.n3155 VSS.n3154 1.54533
R9033 VSS.n3154 VSS.n3153 1.54533
R9034 VSS.n3160 VSS.n3159 1.54533
R9035 VSS.n3169 VSS.n3168 1.54533
R9036 VSS.n3175 VSS.n3174 1.54533
R9037 VSS.n3185 VSS.n3184 1.54533
R9038 VSS.n3190 VSS.n3189 1.54533
R9039 VSS.n3199 VSS.n3198 1.54533
R9040 VSS.n3205 VSS.n3204 1.54533
R9041 VSS.n3215 VSS.n3214 1.54533
R9042 VSS.n3220 VSS.n3219 1.54533
R9043 VSS.n3229 VSS.n3228 1.54533
R9044 VSS.n3235 VSS.n3234 1.54533
R9045 VSS.n3236 VSS.n3235 1.54533
R9046 VSS.n3245 VSS.n3244 1.54533
R9047 VSS.n3250 VSS.n3249 1.54533
R9048 VSS.n3261 VSS.n3260 1.54533
R9049 VSS.n3266 VSS.n3265 1.54533
R9050 VSS.n3275 VSS.n3274 1.54533
R9051 VSS.n3280 VSS.n3279 1.54533
R9052 VSS.n3291 VSS.n3290 1.54533
R9053 VSS.n3296 VSS.n3295 1.54533
R9054 VSS.n3305 VSS.n3304 1.54533
R9055 VSS.n3310 VSS.n3309 1.54533
R9056 VSS.n3321 VSS.n3320 1.54533
R9057 VSS.n3326 VSS.n3325 1.54533
R9058 VSS.n3335 VSS.n3334 1.54533
R9059 VSS.n62 VSS.n61 1.54533
R9060 VSS.n3341 VSS.n52 1.54533
R9061 VSS.n1254 VSS.n1253 1.49652
R9062 VSS.n1269 VSS.n1268 1.49652
R9063 VSS.n1284 VSS.n1283 1.49652
R9064 VSS.n1299 VSS.n1298 1.49652
R9065 VSS.n1314 VSS.n1313 1.49652
R9066 VSS.n2003 VSS.n2002 1.49652
R9067 VSS.n126 VSS.n125 1.49652
R9068 VSS.n141 VSS.n140 1.49652
R9069 VSS.n4221 VSS.n4220 1.49652
R9070 VSS.n3481 VSS.n3480 1.49652
R9071 VSS.n3595 VSS.n3594 1.49652
R9072 VSS.n3709 VSS.n3708 1.49652
R9073 VSS.n3823 VSS.n3822 1.49652
R9074 VSS.n2317 VSS.n2314 1.48887
R9075 VSS.n2668 VSS.n2665 1.48887
R9076 VSS.n3019 VSS.n3016 1.48887
R9077 VSS.n2344 VSS.n2341 1.48827
R9078 VSS.n2414 VSS.n2411 1.48827
R9079 VSS.n2695 VSS.n2692 1.48827
R9080 VSS.n2765 VSS.n2762 1.48827
R9081 VSS.n3046 VSS.n3043 1.48827
R9082 VSS.n160 VSS.n157 1.48702
R9083 VSS.n214 VSS.n211 1.48702
R9084 VSS.n268 VSS.n265 1.48702
R9085 VSS.n2105 VSS.n2104 1.4204
R9086 VSS.n2104 VSS.n2103 1.4204
R9087 VSS.n2095 VSS.n2094 1.4204
R9088 VSS.n2094 VSS.n2093 1.4204
R9089 VSS.n2085 VSS.n2084 1.4204
R9090 VSS.n2084 VSS.n2083 1.4204
R9091 VSS.n2074 VSS.n2073 1.4204
R9092 VSS.n2064 VSS.n2063 1.4204
R9093 VSS.n2063 VSS.n2062 1.4204
R9094 VSS.n2054 VSS.n2053 1.4204
R9095 VSS.n2053 VSS.n2052 1.4204
R9096 VSS.n2041 VSS.n2040 1.4204
R9097 VSS.n2033 VSS.n2032 1.4204
R9098 VSS.n2032 VSS.n2031 1.4204
R9099 VSS.n122 VSS.n121 1.4204
R9100 VSS.n121 VSS.n120 1.4204
R9101 VSS.n2020 VSS.n2019 1.4204
R9102 VSS.n2010 VSS.n2009 1.4204
R9103 VSS.n2009 VSS.n2008 1.4204
R9104 VSS.n2000 VSS.n1999 1.4204
R9105 VSS.n1990 VSS.n1989 1.4204
R9106 VSS.n1989 VSS.n1988 1.4204
R9107 VSS.n1980 VSS.n1979 1.4204
R9108 VSS.n1979 VSS.n1978 1.4204
R9109 VSS.n1970 VSS.n1969 1.4204
R9110 VSS.n1969 VSS.n1968 1.4204
R9111 VSS.n1960 VSS.n1959 1.4204
R9112 VSS.n1959 VSS.n1958 1.4204
R9113 VSS.n1948 VSS.n1947 1.4204
R9114 VSS.n1947 VSS.n1946 1.4204
R9115 VSS.n1938 VSS.n1937 1.4204
R9116 VSS.n1937 VSS.n1936 1.4204
R9117 VSS.n1928 VSS.n1927 1.4204
R9118 VSS.n1927 VSS.n1926 1.4204
R9119 VSS.n1918 VSS.n1917 1.4204
R9120 VSS.n1917 VSS.n1916 1.4204
R9121 VSS.n1908 VSS.n1907 1.4204
R9122 VSS.n1907 VSS.n1906 1.4204
R9123 VSS.n1898 VSS.n1897 1.4204
R9124 VSS.n1897 VSS.n1896 1.4204
R9125 VSS.n1888 VSS.n1887 1.4204
R9126 VSS.n1887 VSS.n1886 1.4204
R9127 VSS.n300 VSS.n299 1.32464
R9128 VSS.n3342 VSS.n3341 1.32464
R9129 VSS.n809 VSS.n808 1.10395
R9130 VSS.n500 VSS.n499 1.10395
R9131 VSS.n82 VSS.n78 1.08219
R9132 VSS.n307 VSS.n300 0.883259
R9133 VSS.n3343 VSS.n3342 0.883259
R9134 VSS.n3868 VSS 0.862479
R9135 VSS.n83 VSS.n82 0.821308
R9136 VSS.n89 VSS.n88 0.780988
R9137 VSS.n90 VSS.n89 0.723468
R9138 VSS.n2907 VSS.n2899 0.662569
R9139 VSS.n2556 VSS.n2548 0.662569
R9140 VSS.n2205 VSS.n2197 0.662569
R9141 VSS.n1918 VSS.n1913 0.662569
R9142 VSS.n161 VSS.n153 0.662569
R9143 VSS.n215 VSS.n207 0.662569
R9144 VSS.n269 VSS.n261 0.662569
R9145 VSS.n66 VSS.n65 0.662569
R9146 VSS.n3320 VSS.n3319 0.662569
R9147 VSS.n4114 VSS.n4113 0.662569
R9148 VSS.n4100 VSS.n4099 0.662569
R9149 VSS.n4086 VSS.n4085 0.662569
R9150 VSS.n4095 VSS.n4094 0.662569
R9151 VSS.n4073 VSS.n4072 0.662569
R9152 VSS.n4081 VSS.n4080 0.662569
R9153 VSS.n17 VSS.n16 0.662569
R9154 VSS.n25 VSS.n24 0.662569
R9155 VSS.n4065 VSS.n4064 0.662569
R9156 VSS.n4044 VSS.n4043 0.662569
R9157 VSS.n4053 VSS.n4052 0.662569
R9158 VSS.n4030 VSS.n4029 0.662569
R9159 VSS.n4039 VSS.n4038 0.662569
R9160 VSS.n4016 VSS.n4015 0.662569
R9161 VSS.n4025 VSS.n4024 0.662569
R9162 VSS.n29 VSS.n28 0.662569
R9163 VSS.n38 VSS.n37 0.662569
R9164 VSS.n4008 VSS.n4007 0.662569
R9165 VSS.n3987 VSS.n3986 0.662569
R9166 VSS.n3996 VSS.n3995 0.662569
R9167 VSS.n3973 VSS.n3972 0.662569
R9168 VSS.n3982 VSS.n3981 0.662569
R9169 VSS.n3959 VSS.n3958 0.662569
R9170 VSS.n3968 VSS.n3967 0.662569
R9171 VSS.n3944 VSS.n3943 0.662569
R9172 VSS.n3954 VSS.n3953 0.662569
R9173 VSS.n3930 VSS.n3929 0.662569
R9174 VSS.n3939 VSS.n3938 0.662569
R9175 VSS.n3915 VSS.n3914 0.662569
R9176 VSS.n3925 VSS.n3924 0.662569
R9177 VSS.n3901 VSS.n3900 0.662569
R9178 VSS.n3910 VSS.n3909 0.662569
R9179 VSS.n43 VSS.n42 0.662569
R9180 VSS.n2042 VSS.n2041 0.577409
R9181 VSS.n2022 VSS.n2021 0.535538
R9182 VSS.n2076 VSS.n2075 0.535538
R9183 VSS.n2002 VSS.n2001 0.517621
R9184 VSS.n3185 VSS.n3183 0.441879
R9185 VSS.n3206 VSS.n3205 0.441879
R9186 VSS.n3896 VSS.n3895 0.441879
R9187 VSS.n3872 VSS.n3871 0.441879
R9188 VSS.n1831 VSS.n1830 0.268864
R9189 VSS.n3348 VSS.n56 0.22119
R9190 VSS.n39 VSS.n38 0.22119
R9191 VSS.n3895 VSS.n3894 0.22119
R9192 VSS.n4124 VSS.n8 0.208232
R9193 VSS.n1836 VSS.n1831 0.188667
R9194 VSS.n1250 VSS.n1249 0.182006
R9195 VSS.n87 VSS 0.156598
R9196 VSS.n1842 VSS.n1836 0.120292
R9197 VSS.n1846 VSS.n1842 0.120292
R9198 VSS.n1850 VSS.n1846 0.120292
R9199 VSS.n1856 VSS.n1850 0.120292
R9200 VSS.n1860 VSS.n1856 0.120292
R9201 VSS.n1864 VSS.n1860 0.120292
R9202 VSS.n1868 VSS.n1864 0.120292
R9203 VSS.n1872 VSS.n1868 0.120292
R9204 VSS.n1878 VSS.n1872 0.120292
R9205 VSS.n1882 VSS.n1878 0.120292
R9206 VSS.n1892 VSS.n1882 0.120292
R9207 VSS.n1902 VSS.n1892 0.120292
R9208 VSS.n1912 VSS.n1902 0.120292
R9209 VSS.n1922 VSS.n1912 0.120292
R9210 VSS.n1932 VSS.n1922 0.120292
R9211 VSS.n1942 VSS.n1932 0.120292
R9212 VSS.n1952 VSS.n1942 0.120292
R9213 VSS.n1964 VSS.n1952 0.120292
R9214 VSS.n1974 VSS.n1964 0.120292
R9215 VSS.n1984 VSS.n1974 0.120292
R9216 VSS.n1994 VSS.n1984 0.120292
R9217 VSS.n2004 VSS.n1994 0.120292
R9218 VSS.n2014 VSS.n2004 0.120292
R9219 VSS.n2025 VSS.n2014 0.120292
R9220 VSS.n2026 VSS.n2025 0.120292
R9221 VSS.n2048 VSS.n2037 0.120292
R9222 VSS.n2058 VSS.n2048 0.120292
R9223 VSS.n2068 VSS.n2058 0.120292
R9224 VSS.n2079 VSS.n2068 0.120292
R9225 VSS.n2089 VSS.n2079 0.120292
R9226 VSS.n2099 VSS.n2089 0.120292
R9227 VSS.n2109 VSS.n2099 0.120292
R9228 VSS.n3069 VSS.n3065 0.120292
R9229 VSS.n3070 VSS.n3069 0.120292
R9230 VSS.n1249 VSS.n1239 0.120292
R9231 VSS.n1239 VSS.n1238 0.120292
R9232 VSS.n1238 VSS.n1234 0.120292
R9233 VSS.n1234 VSS.n1233 0.120292
R9234 VSS.n1233 VSS.n1229 0.120292
R9235 VSS.n1229 VSS.n1225 0.120292
R9236 VSS.n1225 VSS.n1221 0.120292
R9237 VSS.n1221 VSS.n1215 0.120292
R9238 VSS.n1215 VSS.n1211 0.120292
R9239 VSS.n1211 VSS.n1207 0.120292
R9240 VSS.n1207 VSS.n1203 0.120292
R9241 VSS.n1203 VSS.n1198 0.120292
R9242 VSS.n1198 VSS.n1194 0.120292
R9243 VSS.n1194 VSS.n1190 0.120292
R9244 VSS.n1190 VSS.n1186 0.120292
R9245 VSS.n1186 VSS.n1182 0.120292
R9246 VSS.n1182 VSS.n1176 0.120292
R9247 VSS.n1176 VSS.n1172 0.120292
R9248 VSS.n1172 VSS.n1168 0.120292
R9249 VSS.n1168 VSS.n1164 0.120292
R9250 VSS.n1164 VSS.n1160 0.120292
R9251 VSS.n1160 VSS.n1159 0.120292
R9252 VSS.n1159 VSS.n1155 0.120292
R9253 VSS.n1155 VSS.n1151 0.120292
R9254 VSS.n1151 VSS.n1150 0.120292
R9255 VSS.n1138 VSS.n137 0.120292
R9256 VSS.n1138 VSS.n1137 0.120292
R9257 VSS.n1137 VSS.n1133 0.120292
R9258 VSS.n1133 VSS.n1132 0.120292
R9259 VSS.n1132 VSS.n1128 0.120292
R9260 VSS.n1128 VSS.n1124 0.120292
R9261 VSS.n1124 VSS.n1120 0.120292
R9262 VSS.n1120 VSS.n1114 0.120292
R9263 VSS.n1114 VSS.n1110 0.120292
R9264 VSS.n1110 VSS.n1106 0.120292
R9265 VSS.n1106 VSS.n1102 0.120292
R9266 VSS.n1102 VSS.n1097 0.120292
R9267 VSS.n3350 VSS.n3349 0.120292
R9268 VSS.n3356 VSS.n3350 0.120292
R9269 VSS.n3360 VSS.n3356 0.120292
R9270 VSS.n3366 VSS.n3360 0.120292
R9271 VSS.n3367 VSS.n3366 0.120292
R9272 VSS.n3380 VSS.n3374 0.120292
R9273 VSS.n3381 VSS.n3380 0.120292
R9274 VSS.n3868 VSS.n3867 0.120292
R9275 VSS.n3867 VSS.n3863 0.120292
R9276 VSS.n3863 VSS.n3857 0.120292
R9277 VSS.n3850 VSS.n3849 0.120292
R9278 VSS.n3849 VSS.n3843 0.120292
R9279 VSS.n1821 VSS.n1820 0.120292
R9280 VSS.n1820 VSS.n1816 0.120292
R9281 VSS.n1816 VSS.n1815 0.120292
R9282 VSS.n1815 VSS.n1811 0.120292
R9283 VSS.n1811 VSS.n1807 0.120292
R9284 VSS.n1807 VSS.n1803 0.120292
R9285 VSS.n1803 VSS.n1797 0.120292
R9286 VSS.n1797 VSS.n1793 0.120292
R9287 VSS.n1793 VSS.n1789 0.120292
R9288 VSS.n1789 VSS.n1785 0.120292
R9289 VSS.n1785 VSS.n1780 0.120292
R9290 VSS.n1780 VSS.n1776 0.120292
R9291 VSS.n1776 VSS.n1772 0.120292
R9292 VSS.n1772 VSS.n1768 0.120292
R9293 VSS.n1768 VSS.n1764 0.120292
R9294 VSS.n1764 VSS.n1758 0.120292
R9295 VSS.n1758 VSS.n1754 0.120292
R9296 VSS.n1754 VSS.n1750 0.120292
R9297 VSS.n1750 VSS.n1746 0.120292
R9298 VSS.n1746 VSS.n1742 0.120292
R9299 VSS.n1742 VSS.n1741 0.120292
R9300 VSS.n1741 VSS.n1737 0.120292
R9301 VSS.n1737 VSS.n1733 0.120292
R9302 VSS.n1733 VSS.n1732 0.120292
R9303 VSS.n1720 VSS.n1719 0.120292
R9304 VSS.n1719 VSS.n1715 0.120292
R9305 VSS.n1715 VSS.n1714 0.120292
R9306 VSS.n1714 VSS.n1710 0.120292
R9307 VSS.n1710 VSS.n1706 0.120292
R9308 VSS.n1706 VSS.n1702 0.120292
R9309 VSS.n1702 VSS.n1696 0.120292
R9310 VSS.n1696 VSS.n1692 0.120292
R9311 VSS.n1692 VSS.n1688 0.120292
R9312 VSS.n1688 VSS.n1684 0.120292
R9313 VSS.n1684 VSS.n1679 0.120292
R9314 VSS.n1679 VSS.n1675 0.120292
R9315 VSS.n1675 VSS.n1671 0.120292
R9316 VSS.n1671 VSS.n1667 0.120292
R9317 VSS.n1667 VSS.n1663 0.120292
R9318 VSS.n1663 VSS.n1657 0.120292
R9319 VSS.n1657 VSS.n1653 0.120292
R9320 VSS.n1653 VSS.n1649 0.120292
R9321 VSS.n1649 VSS.n1645 0.120292
R9322 VSS.n1645 VSS.n1641 0.120292
R9323 VSS.n1641 VSS.n1640 0.120292
R9324 VSS.n1640 VSS.n1636 0.120292
R9325 VSS.n1636 VSS.n1632 0.120292
R9326 VSS.n1632 VSS.n1631 0.120292
R9327 VSS.n1619 VSS.n1618 0.120292
R9328 VSS.n1618 VSS.n1614 0.120292
R9329 VSS.n1614 VSS.n1613 0.120292
R9330 VSS.n1613 VSS.n1609 0.120292
R9331 VSS.n1609 VSS.n1605 0.120292
R9332 VSS.n1605 VSS.n1601 0.120292
R9333 VSS.n1601 VSS.n1595 0.120292
R9334 VSS.n1595 VSS.n1591 0.120292
R9335 VSS.n1591 VSS.n1587 0.120292
R9336 VSS.n1587 VSS.n1583 0.120292
R9337 VSS.n1583 VSS.n1578 0.120292
R9338 VSS.n1578 VSS.n1574 0.120292
R9339 VSS.n1574 VSS.n1570 0.120292
R9340 VSS.n1570 VSS.n1566 0.120292
R9341 VSS.n1566 VSS.n1562 0.120292
R9342 VSS.n1562 VSS.n1556 0.120292
R9343 VSS.n1556 VSS.n1552 0.120292
R9344 VSS.n1552 VSS.n1548 0.120292
R9345 VSS.n1548 VSS.n1544 0.120292
R9346 VSS.n1544 VSS.n1540 0.120292
R9347 VSS.n1540 VSS.n1539 0.120292
R9348 VSS.n1539 VSS.n1535 0.120292
R9349 VSS.n1535 VSS.n1531 0.120292
R9350 VSS.n1531 VSS.n1530 0.120292
R9351 VSS.n1518 VSS.n1517 0.120292
R9352 VSS.n1517 VSS.n1513 0.120292
R9353 VSS.n1513 VSS.n1512 0.120292
R9354 VSS.n1512 VSS.n1508 0.120292
R9355 VSS.n1508 VSS.n1504 0.120292
R9356 VSS.n1504 VSS.n1500 0.120292
R9357 VSS.n1500 VSS.n1494 0.120292
R9358 VSS.n1494 VSS.n1490 0.120292
R9359 VSS.n1490 VSS.n1486 0.120292
R9360 VSS.n1486 VSS.n1482 0.120292
R9361 VSS.n1482 VSS.n1477 0.120292
R9362 VSS.n1477 VSS.n1473 0.120292
R9363 VSS.n1473 VSS.n1469 0.120292
R9364 VSS.n1469 VSS.n1465 0.120292
R9365 VSS.n1465 VSS.n1461 0.120292
R9366 VSS.n1461 VSS.n1455 0.120292
R9367 VSS.n1455 VSS.n1451 0.120292
R9368 VSS.n1451 VSS.n1447 0.120292
R9369 VSS.n1447 VSS.n1443 0.120292
R9370 VSS.n1443 VSS.n1439 0.120292
R9371 VSS.n1439 VSS.n1438 0.120292
R9372 VSS.n1438 VSS.n1434 0.120292
R9373 VSS.n1434 VSS.n1430 0.120292
R9374 VSS.n1430 VSS.n1429 0.120292
R9375 VSS.n1417 VSS.n1416 0.120292
R9376 VSS.n1416 VSS.n1412 0.120292
R9377 VSS.n1412 VSS.n1411 0.120292
R9378 VSS.n1411 VSS.n1407 0.120292
R9379 VSS.n1407 VSS.n1403 0.120292
R9380 VSS.n1403 VSS.n1399 0.120292
R9381 VSS.n1399 VSS.n1393 0.120292
R9382 VSS.n1393 VSS.n1389 0.120292
R9383 VSS.n1389 VSS.n1385 0.120292
R9384 VSS.n1385 VSS.n1381 0.120292
R9385 VSS.n1381 VSS.n1376 0.120292
R9386 VSS.n1376 VSS.n1372 0.120292
R9387 VSS.n1372 VSS.n1368 0.120292
R9388 VSS.n1368 VSS.n1364 0.120292
R9389 VSS.n1364 VSS.n1360 0.120292
R9390 VSS.n1360 VSS.n1354 0.120292
R9391 VSS.n1354 VSS.n1350 0.120292
R9392 VSS.n1350 VSS.n1346 0.120292
R9393 VSS.n1346 VSS.n1342 0.120292
R9394 VSS.n1342 VSS.n1338 0.120292
R9395 VSS.n1338 VSS.n1337 0.120292
R9396 VSS.n1337 VSS.n1333 0.120292
R9397 VSS.n1333 VSS.n1329 0.120292
R9398 VSS.n1329 VSS.n1328 0.120292
R9399 VSS.n4130 VSS.n4124 0.120292
R9400 VSS.n4134 VSS.n4130 0.120292
R9401 VSS.n4138 VSS.n4134 0.120292
R9402 VSS.n4144 VSS.n4138 0.120292
R9403 VSS.n4148 VSS.n4144 0.120292
R9404 VSS.n4152 VSS.n4148 0.120292
R9405 VSS.n4156 VSS.n4152 0.120292
R9406 VSS.n4160 VSS.n4156 0.120292
R9407 VSS.n4166 VSS.n4160 0.120292
R9408 VSS.n4170 VSS.n4166 0.120292
R9409 VSS.n4174 VSS.n4170 0.120292
R9410 VSS.n4178 VSS.n4174 0.120292
R9411 VSS.n4182 VSS.n4178 0.120292
R9412 VSS.n4187 VSS.n4182 0.120292
R9413 VSS.n4191 VSS.n4187 0.120292
R9414 VSS.n4195 VSS.n4191 0.120292
R9415 VSS.n4199 VSS.n4195 0.120292
R9416 VSS.n4205 VSS.n4199 0.120292
R9417 VSS.n4209 VSS.n4205 0.120292
R9418 VSS.n4213 VSS.n4209 0.120292
R9419 VSS.n4217 VSS.n4213 0.120292
R9420 VSS.n4222 VSS.n4217 0.120292
R9421 VSS.n4226 VSS.n4222 0.120292
R9422 VSS.n4227 VSS.n4226 0.120292
R9423 VSS.n4227 VSS.n0 0.120292
R9424 VSS.n4238 VSS.n6 0.120292
R9425 VSS.n3394 VSS.n6 0.120292
R9426 VSS.n3398 VSS.n3394 0.120292
R9427 VSS.n3404 VSS.n3398 0.120292
R9428 VSS.n3408 VSS.n3404 0.120292
R9429 VSS.n3412 VSS.n3408 0.120292
R9430 VSS.n3416 VSS.n3412 0.120292
R9431 VSS.n3420 VSS.n3416 0.120292
R9432 VSS.n3426 VSS.n3420 0.120292
R9433 VSS.n3430 VSS.n3426 0.120292
R9434 VSS.n3434 VSS.n3430 0.120292
R9435 VSS.n3438 VSS.n3434 0.120292
R9436 VSS.n3442 VSS.n3438 0.120292
R9437 VSS.n3447 VSS.n3442 0.120292
R9438 VSS.n3451 VSS.n3447 0.120292
R9439 VSS.n3455 VSS.n3451 0.120292
R9440 VSS.n3459 VSS.n3455 0.120292
R9441 VSS.n3465 VSS.n3459 0.120292
R9442 VSS.n3469 VSS.n3465 0.120292
R9443 VSS.n3473 VSS.n3469 0.120292
R9444 VSS.n3477 VSS.n3473 0.120292
R9445 VSS.n3482 VSS.n3477 0.120292
R9446 VSS.n3486 VSS.n3482 0.120292
R9447 VSS.n3489 VSS.n3486 0.120292
R9448 VSS.n3489 VSS.n3488 0.120292
R9449 VSS.n3504 VSS.n3498 0.120292
R9450 VSS.n3508 VSS.n3504 0.120292
R9451 VSS.n3512 VSS.n3508 0.120292
R9452 VSS.n3518 VSS.n3512 0.120292
R9453 VSS.n3522 VSS.n3518 0.120292
R9454 VSS.n3526 VSS.n3522 0.120292
R9455 VSS.n3530 VSS.n3526 0.120292
R9456 VSS.n3534 VSS.n3530 0.120292
R9457 VSS.n3540 VSS.n3534 0.120292
R9458 VSS.n3544 VSS.n3540 0.120292
R9459 VSS.n3548 VSS.n3544 0.120292
R9460 VSS.n3552 VSS.n3548 0.120292
R9461 VSS.n3556 VSS.n3552 0.120292
R9462 VSS.n3561 VSS.n3556 0.120292
R9463 VSS.n3565 VSS.n3561 0.120292
R9464 VSS.n3569 VSS.n3565 0.120292
R9465 VSS.n3573 VSS.n3569 0.120292
R9466 VSS.n3579 VSS.n3573 0.120292
R9467 VSS.n3583 VSS.n3579 0.120292
R9468 VSS.n3587 VSS.n3583 0.120292
R9469 VSS.n3591 VSS.n3587 0.120292
R9470 VSS.n3596 VSS.n3591 0.120292
R9471 VSS.n3600 VSS.n3596 0.120292
R9472 VSS.n3603 VSS.n3600 0.120292
R9473 VSS.n3603 VSS.n3602 0.120292
R9474 VSS.n3618 VSS.n3612 0.120292
R9475 VSS.n3622 VSS.n3618 0.120292
R9476 VSS.n3626 VSS.n3622 0.120292
R9477 VSS.n3632 VSS.n3626 0.120292
R9478 VSS.n3636 VSS.n3632 0.120292
R9479 VSS.n3640 VSS.n3636 0.120292
R9480 VSS.n3644 VSS.n3640 0.120292
R9481 VSS.n3648 VSS.n3644 0.120292
R9482 VSS.n3654 VSS.n3648 0.120292
R9483 VSS.n3658 VSS.n3654 0.120292
R9484 VSS.n3662 VSS.n3658 0.120292
R9485 VSS.n3666 VSS.n3662 0.120292
R9486 VSS.n3670 VSS.n3666 0.120292
R9487 VSS.n3675 VSS.n3670 0.120292
R9488 VSS.n3679 VSS.n3675 0.120292
R9489 VSS.n3683 VSS.n3679 0.120292
R9490 VSS.n3687 VSS.n3683 0.120292
R9491 VSS.n3693 VSS.n3687 0.120292
R9492 VSS.n3697 VSS.n3693 0.120292
R9493 VSS.n3701 VSS.n3697 0.120292
R9494 VSS.n3705 VSS.n3701 0.120292
R9495 VSS.n3710 VSS.n3705 0.120292
R9496 VSS.n3714 VSS.n3710 0.120292
R9497 VSS.n3717 VSS.n3714 0.120292
R9498 VSS.n3717 VSS.n3716 0.120292
R9499 VSS.n3732 VSS.n3726 0.120292
R9500 VSS.n3736 VSS.n3732 0.120292
R9501 VSS.n3740 VSS.n3736 0.120292
R9502 VSS.n3746 VSS.n3740 0.120292
R9503 VSS.n3750 VSS.n3746 0.120292
R9504 VSS.n3754 VSS.n3750 0.120292
R9505 VSS.n3758 VSS.n3754 0.120292
R9506 VSS.n3762 VSS.n3758 0.120292
R9507 VSS.n3768 VSS.n3762 0.120292
R9508 VSS.n3772 VSS.n3768 0.120292
R9509 VSS.n3776 VSS.n3772 0.120292
R9510 VSS.n3780 VSS.n3776 0.120292
R9511 VSS.n3784 VSS.n3780 0.120292
R9512 VSS.n3789 VSS.n3784 0.120292
R9513 VSS.n3793 VSS.n3789 0.120292
R9514 VSS.n3797 VSS.n3793 0.120292
R9515 VSS.n3801 VSS.n3797 0.120292
R9516 VSS.n3807 VSS.n3801 0.120292
R9517 VSS.n3811 VSS.n3807 0.120292
R9518 VSS.n3815 VSS.n3811 0.120292
R9519 VSS.n3819 VSS.n3815 0.120292
R9520 VSS.n3824 VSS.n3819 0.120292
R9521 VSS.n3828 VSS.n3824 0.120292
R9522 VSS.n3834 VSS.n3828 0.120292
R9523 VSS.n3835 VSS.n3834 0.120292
R9524 VSS.n2110 VSS.n2109 0.108573
R9525 VSS.n1097 VSS.n1093 0.107271
R9526 VSS.n2124 VSS.n2123 0.0981562
R9527 VSS.n2140 VSS.n2139 0.0981562
R9528 VSS.n2154 VSS.n2153 0.0981562
R9529 VSS.n2168 VSS.n2167 0.0981562
R9530 VSS.n2182 VSS.n2181 0.0981562
R9531 VSS.n2196 VSS.n2195 0.0981562
R9532 VSS.n2210 VSS.n2209 0.0981562
R9533 VSS.n2224 VSS.n2223 0.0981562
R9534 VSS.n2238 VSS.n2237 0.0981562
R9535 VSS.n2252 VSS.n2251 0.0981562
R9536 VSS.n2268 VSS.n2267 0.0981562
R9537 VSS.n2282 VSS.n2281 0.0981562
R9538 VSS.n2296 VSS.n2295 0.0981562
R9539 VSS.n2310 VSS.n2309 0.0981562
R9540 VSS.n2322 VSS.n2321 0.0981562
R9541 VSS.n2336 VSS.n2335 0.0981562
R9542 VSS.n2349 VSS.n2348 0.0981562
R9543 VSS.n2365 VSS.n2364 0.0981562
R9544 VSS.n2378 VSS.n2377 0.0981562
R9545 VSS.n2392 VSS.n2391 0.0981562
R9546 VSS.n2406 VSS.n2405 0.0981562
R9547 VSS.n2419 VSS.n2418 0.0981562
R9548 VSS.n2433 VSS.n2432 0.0981562
R9549 VSS.n2447 VSS.n2446 0.0981562
R9550 VSS.n2461 VSS.n2460 0.0981562
R9551 VSS.n2475 VSS.n2474 0.0981562
R9552 VSS.n2491 VSS.n2490 0.0981562
R9553 VSS.n2505 VSS.n2504 0.0981562
R9554 VSS.n2519 VSS.n2518 0.0981562
R9555 VSS.n2533 VSS.n2532 0.0981562
R9556 VSS.n2547 VSS.n2546 0.0981562
R9557 VSS.n2561 VSS.n2560 0.0981562
R9558 VSS.n2575 VSS.n2574 0.0981562
R9559 VSS.n2589 VSS.n2588 0.0981562
R9560 VSS.n2603 VSS.n2602 0.0981562
R9561 VSS.n2619 VSS.n2618 0.0981562
R9562 VSS.n2633 VSS.n2632 0.0981562
R9563 VSS.n2647 VSS.n2646 0.0981562
R9564 VSS.n2661 VSS.n2660 0.0981562
R9565 VSS.n2673 VSS.n2672 0.0981562
R9566 VSS.n2687 VSS.n2686 0.0981562
R9567 VSS.n2700 VSS.n2699 0.0981562
R9568 VSS.n2716 VSS.n2715 0.0981562
R9569 VSS.n2729 VSS.n2728 0.0981562
R9570 VSS.n2743 VSS.n2742 0.0981562
R9571 VSS.n2757 VSS.n2756 0.0981562
R9572 VSS.n2770 VSS.n2769 0.0981562
R9573 VSS.n2784 VSS.n2783 0.0981562
R9574 VSS.n2798 VSS.n2797 0.0981562
R9575 VSS.n2812 VSS.n2811 0.0981562
R9576 VSS.n2826 VSS.n2825 0.0981562
R9577 VSS.n2842 VSS.n2841 0.0981562
R9578 VSS.n2856 VSS.n2855 0.0981562
R9579 VSS.n2870 VSS.n2869 0.0981562
R9580 VSS.n2884 VSS.n2883 0.0981562
R9581 VSS.n2898 VSS.n2897 0.0981562
R9582 VSS.n2912 VSS.n2911 0.0981562
R9583 VSS.n2926 VSS.n2925 0.0981562
R9584 VSS.n2940 VSS.n2939 0.0981562
R9585 VSS.n2954 VSS.n2953 0.0981562
R9586 VSS.n2970 VSS.n2969 0.0981562
R9587 VSS.n2984 VSS.n2983 0.0981562
R9588 VSS.n2998 VSS.n2997 0.0981562
R9589 VSS.n3012 VSS.n3011 0.0981562
R9590 VSS.n3024 VSS.n3023 0.0981562
R9591 VSS.n3038 VSS.n3037 0.0981562
R9592 VSS.n3052 VSS.n3051 0.0981562
R9593 VSS.n1080 VSS.n1079 0.0981562
R9594 VSS.n1066 VSS.n1065 0.0981562
R9595 VSS.n1052 VSS.n1051 0.0981562
R9596 VSS.n1036 VSS.n1035 0.0981562
R9597 VSS.n1022 VSS.n1021 0.0981562
R9598 VSS.n1008 VSS.n1007 0.0981562
R9599 VSS.n994 VSS.n993 0.0981562
R9600 VSS.n980 VSS.n979 0.0981562
R9601 VSS.n977 VSS.n976 0.0981562
R9602 VSS.n963 VSS.n962 0.0981562
R9603 VSS.n949 VSS.n948 0.0981562
R9604 VSS.n946 VSS.n945 0.0981562
R9605 VSS.n186 VSS.n185 0.0981562
R9606 VSS.n929 VSS.n928 0.0981562
R9607 VSS.n915 VSS.n914 0.0981562
R9608 VSS.n912 VSS.n911 0.0981562
R9609 VSS.n898 VSS.n897 0.0981562
R9610 VSS.n884 VSS.n883 0.0981562
R9611 VSS.n870 VSS.n869 0.0981562
R9612 VSS.n855 VSS.n854 0.0981562
R9613 VSS.n841 VSS.n840 0.0981562
R9614 VSS.n827 VSS.n826 0.0981562
R9615 VSS.n813 VSS.n812 0.0981562
R9616 VSS.n798 VSS.n797 0.0981562
R9617 VSS.n785 VSS.n784 0.0981562
R9618 VSS.n771 VSS.n770 0.0981562
R9619 VSS.n757 VSS.n756 0.0981562
R9620 VSS.n743 VSS.n742 0.0981562
R9621 VSS.n727 VSS.n726 0.0981562
R9622 VSS.n713 VSS.n712 0.0981562
R9623 VSS.n699 VSS.n698 0.0981562
R9624 VSS.n685 VSS.n684 0.0981562
R9625 VSS.n671 VSS.n670 0.0981562
R9626 VSS.n668 VSS.n667 0.0981562
R9627 VSS.n654 VSS.n653 0.0981562
R9628 VSS.n640 VSS.n639 0.0981562
R9629 VSS.n637 VSS.n636 0.0981562
R9630 VSS.n240 VSS.n239 0.0981562
R9631 VSS.n620 VSS.n619 0.0981562
R9632 VSS.n606 VSS.n605 0.0981562
R9633 VSS.n603 VSS.n602 0.0981562
R9634 VSS.n589 VSS.n588 0.0981562
R9635 VSS.n575 VSS.n574 0.0981562
R9636 VSS.n561 VSS.n560 0.0981562
R9637 VSS.n546 VSS.n545 0.0981562
R9638 VSS.n532 VSS.n531 0.0981562
R9639 VSS.n518 VSS.n517 0.0981562
R9640 VSS.n504 VSS.n503 0.0981562
R9641 VSS.n489 VSS.n488 0.0981562
R9642 VSS.n476 VSS.n475 0.0981562
R9643 VSS.n462 VSS.n461 0.0981562
R9644 VSS.n448 VSS.n447 0.0981562
R9645 VSS.n434 VSS.n433 0.0981562
R9646 VSS.n418 VSS.n417 0.0981562
R9647 VSS.n404 VSS.n403 0.0981562
R9648 VSS.n390 VSS.n389 0.0981562
R9649 VSS.n376 VSS.n375 0.0981562
R9650 VSS.n362 VSS.n361 0.0981562
R9651 VSS.n359 VSS.n358 0.0981562
R9652 VSS.n345 VSS.n344 0.0981562
R9653 VSS.n331 VSS.n330 0.0981562
R9654 VSS.n328 VSS.n327 0.0981562
R9655 VSS.n312 VSS.n311 0.0981562
R9656 VSS.n298 VSS.n297 0.0981562
R9657 VSS.n284 VSS.n63 0.0981562
R9658 VSS.n3083 VSS.n3082 0.0981562
R9659 VSS.n3099 VSS.n3098 0.0981562
R9660 VSS.n3113 VSS.n3112 0.0981562
R9661 VSS.n3129 VSS.n3128 0.0981562
R9662 VSS.n3142 VSS.n3141 0.0981562
R9663 VSS.n3158 VSS.n3157 0.0981562
R9664 VSS.n3172 VSS.n3171 0.0981562
R9665 VSS.n3188 VSS.n3187 0.0981562
R9666 VSS.n3202 VSS.n3201 0.0981562
R9667 VSS.n3218 VSS.n3217 0.0981562
R9668 VSS.n3232 VSS.n3231 0.0981562
R9669 VSS.n3248 VSS.n3247 0.0981562
R9670 VSS.n3264 VSS.n3263 0.0981562
R9671 VSS.n3278 VSS.n3277 0.0981562
R9672 VSS.n3294 VSS.n3293 0.0981562
R9673 VSS.n3308 VSS.n3307 0.0981562
R9674 VSS.n3324 VSS.n3323 0.0981562
R9675 VSS.n3338 VSS.n3337 0.0981562
R9676 VSS.n4103 VSS.n4102 0.0981562
R9677 VSS.n4098 VSS.n4097 0.0981562
R9678 VSS.n4084 VSS.n4083 0.0981562
R9679 VSS.n4071 VSS.n4070 0.0981562
R9680 VSS.n4068 VSS.n4067 0.0981562
R9681 VSS.n4056 VSS.n4055 0.0981562
R9682 VSS.n4042 VSS.n4041 0.0981562
R9683 VSS.n4028 VSS.n4027 0.0981562
R9684 VSS.n4014 VSS.n4013 0.0981562
R9685 VSS.n4011 VSS.n4010 0.0981562
R9686 VSS.n3999 VSS.n3998 0.0981562
R9687 VSS.n3985 VSS.n3984 0.0981562
R9688 VSS.n3971 VSS.n3970 0.0981562
R9689 VSS.n3957 VSS.n3956 0.0981562
R9690 VSS.n3942 VSS.n3941 0.0981562
R9691 VSS.n3928 VSS.n3927 0.0981562
R9692 VSS.n3913 VSS.n3912 0.0981562
R9693 VSS.n3899 VSS.n3898 0.0981562
R9694 VSS.n1821 VSS 0.0968542
R9695 VSS.n1720 VSS 0.0968542
R9696 VSS.n1619 VSS 0.0968542
R9697 VSS.n1518 VSS 0.0968542
R9698 VSS.n1417 VSS 0.0968542
R9699 VSS.n1831 VSS.n1250 0.0852709
R9700 VSS.n14 VSS 0.078625
R9701 VSS.n1250 VSS.n8 0.0637239
R9702 VSS.n2026 VSS 0.0603958
R9703 VSS.n2037 VSS 0.0603958
R9704 VSS.n1150 VSS 0.0603958
R9705 VSS.n137 VSS 0.0603958
R9706 VSS.n3367 VSS 0.0603958
R9707 VSS.n3374 VSS 0.0603958
R9708 VSS.n3381 VSS 0.0603958
R9709 VSS.n3857 VSS 0.0603958
R9710 VSS.n3850 VSS 0.0603958
R9711 VSS.n3843 VSS 0.0603958
R9712 VSS.n1732 VSS 0.0603958
R9713 VSS.n1265 VSS 0.0603958
R9714 VSS.n1631 VSS 0.0603958
R9715 VSS.n1280 VSS 0.0603958
R9716 VSS.n1530 VSS 0.0603958
R9717 VSS.n1295 VSS 0.0603958
R9718 VSS.n1429 VSS 0.0603958
R9719 VSS.n1310 VSS 0.0603958
R9720 VSS.n1328 VSS 0.0603958
R9721 VSS VSS.n0 0.0603958
R9722 VSS VSS.n4238 0.0603958
R9723 VSS.n3488 VSS 0.0603958
R9724 VSS.n3498 VSS 0.0603958
R9725 VSS.n3602 VSS 0.0603958
R9726 VSS.n3612 VSS 0.0603958
R9727 VSS.n3716 VSS 0.0603958
R9728 VSS.n3726 VSS 0.0603958
R9729 VSS.n3835 VSS 0.0603958
R9730 VSS VSS.n41 0.0564896
R9731 VSS.n11 VSS.n8 0.0537635
R9732 VSS VSS.n163 0.0512812
R9733 VSS VSS.n217 0.0512812
R9734 VSS VSS.n271 0.0512812
R9735 VSS.n2350 VSS 0.0499792
R9736 VSS.n2701 VSS 0.0499792
R9737 VSS.n3054 VSS 0.0499792
R9738 VSS VSS.n103 0.0486771
R9739 VSS VSS.n91 0.0486771
R9740 VSS.n183 VSS 0.047375
R9741 VSS.n237 VSS 0.047375
R9742 VSS.n283 VSS 0.047375
R9743 VSS.n3065 VSS 0.0356562
R9744 VSS.n3349 VSS 0.0343542
R9745 VSS VSS.n12 0.0239375
R9746 VSS.n1830 VSS 0.0239375
R9747 VSS VSS.n1265 0.0239375
R9748 VSS VSS.n1280 0.0239375
R9749 VSS VSS.n1295 0.0239375
R9750 VSS VSS.n1310 0.0239375
R9751 VSS.n3070 VSS 0.0226354
R9752 VSS.n4104 VSS.n14 0.0187292
R9753 VSS.n4102 VSS.n4101 0.0187292
R9754 VSS.n4097 VSS.n4096 0.0187292
R9755 VSS.n4083 VSS.n4082 0.0187292
R9756 VSS.n4070 VSS.n4069 0.0187292
R9757 VSS.n4067 VSS.n4066 0.0187292
R9758 VSS.n4055 VSS.n4054 0.0187292
R9759 VSS.n4041 VSS.n4040 0.0187292
R9760 VSS.n4027 VSS.n4026 0.0187292
R9761 VSS.n4013 VSS.n4012 0.0187292
R9762 VSS.n4010 VSS.n4009 0.0187292
R9763 VSS.n3998 VSS.n3997 0.0187292
R9764 VSS.n3984 VSS.n3983 0.0187292
R9765 VSS.n3970 VSS.n3969 0.0187292
R9766 VSS.n3956 VSS.n3955 0.0187292
R9767 VSS.n3941 VSS.n3940 0.0187292
R9768 VSS.n3927 VSS.n3926 0.0187292
R9769 VSS.n3912 VSS.n3911 0.0187292
R9770 VSS.n3898 VSS.n3897 0.0187292
R9771 VSS.n1093 VSS.n1092 0.0135208
R9772 VSS.n1079 VSS.n1078 0.0135208
R9773 VSS.n1065 VSS.n1064 0.0135208
R9774 VSS.n1051 VSS.n1050 0.0135208
R9775 VSS.n1035 VSS.n1034 0.0135208
R9776 VSS.n1021 VSS.n1020 0.0135208
R9777 VSS.n1007 VSS.n1006 0.0135208
R9778 VSS.n993 VSS.n992 0.0135208
R9779 VSS.n979 VSS.n978 0.0135208
R9780 VSS.n976 VSS.n975 0.0135208
R9781 VSS.n962 VSS.n961 0.0135208
R9782 VSS.n948 VSS.n947 0.0135208
R9783 VSS.n945 VSS.n944 0.0135208
R9784 VSS.n184 VSS.n183 0.0135208
R9785 VSS.n930 VSS.n186 0.0135208
R9786 VSS.n928 VSS.n927 0.0135208
R9787 VSS.n914 VSS.n913 0.0135208
R9788 VSS.n911 VSS.n910 0.0135208
R9789 VSS.n897 VSS.n896 0.0135208
R9790 VSS.n883 VSS.n882 0.0135208
R9791 VSS.n869 VSS.n868 0.0135208
R9792 VSS.n854 VSS.n853 0.0135208
R9793 VSS.n840 VSS.n839 0.0135208
R9794 VSS.n826 VSS.n825 0.0135208
R9795 VSS.n812 VSS.n811 0.0135208
R9796 VSS.n797 VSS.n796 0.0135208
R9797 VSS.n784 VSS.n783 0.0135208
R9798 VSS.n770 VSS.n769 0.0135208
R9799 VSS.n756 VSS.n755 0.0135208
R9800 VSS.n742 VSS.n741 0.0135208
R9801 VSS.n726 VSS.n725 0.0135208
R9802 VSS.n712 VSS.n711 0.0135208
R9803 VSS.n698 VSS.n697 0.0135208
R9804 VSS.n684 VSS.n683 0.0135208
R9805 VSS.n670 VSS.n669 0.0135208
R9806 VSS.n667 VSS.n666 0.0135208
R9807 VSS.n653 VSS.n652 0.0135208
R9808 VSS.n639 VSS.n638 0.0135208
R9809 VSS.n636 VSS.n635 0.0135208
R9810 VSS.n238 VSS.n237 0.0135208
R9811 VSS.n621 VSS.n240 0.0135208
R9812 VSS.n619 VSS.n618 0.0135208
R9813 VSS.n605 VSS.n604 0.0135208
R9814 VSS.n602 VSS.n601 0.0135208
R9815 VSS.n588 VSS.n587 0.0135208
R9816 VSS.n574 VSS.n573 0.0135208
R9817 VSS.n560 VSS.n559 0.0135208
R9818 VSS.n545 VSS.n544 0.0135208
R9819 VSS.n531 VSS.n530 0.0135208
R9820 VSS.n517 VSS.n516 0.0135208
R9821 VSS.n503 VSS.n502 0.0135208
R9822 VSS.n488 VSS.n487 0.0135208
R9823 VSS.n475 VSS.n474 0.0135208
R9824 VSS.n461 VSS.n460 0.0135208
R9825 VSS.n447 VSS.n446 0.0135208
R9826 VSS.n433 VSS.n432 0.0135208
R9827 VSS.n417 VSS.n416 0.0135208
R9828 VSS.n403 VSS.n402 0.0135208
R9829 VSS.n389 VSS.n388 0.0135208
R9830 VSS.n375 VSS.n374 0.0135208
R9831 VSS.n361 VSS.n360 0.0135208
R9832 VSS.n358 VSS.n357 0.0135208
R9833 VSS.n344 VSS.n343 0.0135208
R9834 VSS.n330 VSS.n329 0.0135208
R9835 VSS.n327 VSS.n326 0.0135208
R9836 VSS.n313 VSS.n283 0.0135208
R9837 VSS.n311 VSS.n310 0.0135208
R9838 VSS.n297 VSS.n296 0.0135208
R9839 VSS.n3081 VSS.n63 0.0135208
R9840 VSS.n3097 VSS.n3083 0.0135208
R9841 VSS.n3111 VSS.n3099 0.0135208
R9842 VSS.n3127 VSS.n3113 0.0135208
R9843 VSS.n3140 VSS.n3129 0.0135208
R9844 VSS.n3156 VSS.n3142 0.0135208
R9845 VSS.n3170 VSS.n3158 0.0135208
R9846 VSS.n3186 VSS.n3172 0.0135208
R9847 VSS.n3200 VSS.n3188 0.0135208
R9848 VSS.n3216 VSS.n3202 0.0135208
R9849 VSS.n3230 VSS.n3218 0.0135208
R9850 VSS.n3246 VSS.n3232 0.0135208
R9851 VSS.n3262 VSS.n3248 0.0135208
R9852 VSS.n3276 VSS.n3264 0.0135208
R9853 VSS.n3292 VSS.n3278 0.0135208
R9854 VSS.n3306 VSS.n3294 0.0135208
R9855 VSS.n3322 VSS.n3308 0.0135208
R9856 VSS.n3336 VSS.n3324 0.0135208
R9857 VSS.n3340 VSS.n3338 0.0135208
R9858 VSS.n2122 VSS.n2110 0.0122188
R9859 VSS.n2138 VSS.n2124 0.0122188
R9860 VSS.n2152 VSS.n2140 0.0122188
R9861 VSS.n2166 VSS.n2154 0.0122188
R9862 VSS.n2180 VSS.n2168 0.0122188
R9863 VSS.n2194 VSS.n2182 0.0122188
R9864 VSS.n2208 VSS.n2196 0.0122188
R9865 VSS.n2222 VSS.n2210 0.0122188
R9866 VSS.n2236 VSS.n2224 0.0122188
R9867 VSS.n2250 VSS.n2238 0.0122188
R9868 VSS.n2266 VSS.n2252 0.0122188
R9869 VSS.n2280 VSS.n2268 0.0122188
R9870 VSS.n2294 VSS.n2282 0.0122188
R9871 VSS.n2308 VSS.n2296 0.0122188
R9872 VSS.n2320 VSS.n2310 0.0122188
R9873 VSS.n2334 VSS.n2322 0.0122188
R9874 VSS.n2347 VSS.n2336 0.0122188
R9875 VSS.n2351 VSS.n2349 0.0122188
R9876 VSS.n2363 VSS.n103 0.0122188
R9877 VSS.n2376 VSS.n2365 0.0122188
R9878 VSS.n2390 VSS.n2378 0.0122188
R9879 VSS.n2404 VSS.n2392 0.0122188
R9880 VSS.n2417 VSS.n2406 0.0122188
R9881 VSS.n2431 VSS.n2419 0.0122188
R9882 VSS.n2445 VSS.n2433 0.0122188
R9883 VSS.n2459 VSS.n2447 0.0122188
R9884 VSS.n2473 VSS.n2461 0.0122188
R9885 VSS.n2489 VSS.n2475 0.0122188
R9886 VSS.n2503 VSS.n2491 0.0122188
R9887 VSS.n2517 VSS.n2505 0.0122188
R9888 VSS.n2531 VSS.n2519 0.0122188
R9889 VSS.n2545 VSS.n2533 0.0122188
R9890 VSS.n2559 VSS.n2547 0.0122188
R9891 VSS.n2573 VSS.n2561 0.0122188
R9892 VSS.n2587 VSS.n2575 0.0122188
R9893 VSS.n2601 VSS.n2589 0.0122188
R9894 VSS.n2617 VSS.n2603 0.0122188
R9895 VSS.n2631 VSS.n2619 0.0122188
R9896 VSS.n2645 VSS.n2633 0.0122188
R9897 VSS.n2659 VSS.n2647 0.0122188
R9898 VSS.n2671 VSS.n2661 0.0122188
R9899 VSS.n2685 VSS.n2673 0.0122188
R9900 VSS.n2698 VSS.n2687 0.0122188
R9901 VSS.n2702 VSS.n2700 0.0122188
R9902 VSS.n2714 VSS.n91 0.0122188
R9903 VSS.n2727 VSS.n2716 0.0122188
R9904 VSS.n2741 VSS.n2729 0.0122188
R9905 VSS.n2755 VSS.n2743 0.0122188
R9906 VSS.n2768 VSS.n2757 0.0122188
R9907 VSS.n2782 VSS.n2770 0.0122188
R9908 VSS.n2796 VSS.n2784 0.0122188
R9909 VSS.n2810 VSS.n2798 0.0122188
R9910 VSS.n2824 VSS.n2812 0.0122188
R9911 VSS.n2840 VSS.n2826 0.0122188
R9912 VSS.n2854 VSS.n2842 0.0122188
R9913 VSS.n2868 VSS.n2856 0.0122188
R9914 VSS.n2882 VSS.n2870 0.0122188
R9915 VSS.n2896 VSS.n2884 0.0122188
R9916 VSS.n2910 VSS.n2898 0.0122188
R9917 VSS.n2924 VSS.n2912 0.0122188
R9918 VSS.n2938 VSS.n2926 0.0122188
R9919 VSS.n2952 VSS.n2940 0.0122188
R9920 VSS.n2968 VSS.n2954 0.0122188
R9921 VSS.n2982 VSS.n2970 0.0122188
R9922 VSS.n2996 VSS.n2984 0.0122188
R9923 VSS.n3010 VSS.n2998 0.0122188
R9924 VSS.n3022 VSS.n3012 0.0122188
R9925 VSS.n3036 VSS.n3024 0.0122188
R9926 VSS.n3049 VSS.n3038 0.0122188
R9927 VSS.n3339 VSS 0.0122188
R9928 VSS.n2123 VSS.n2122 0.0109167
R9929 VSS.n2139 VSS.n2138 0.0109167
R9930 VSS.n2153 VSS.n2152 0.0109167
R9931 VSS.n2167 VSS.n2166 0.0109167
R9932 VSS.n2181 VSS.n2180 0.0109167
R9933 VSS.n2195 VSS.n2194 0.0109167
R9934 VSS.n2209 VSS.n2208 0.0109167
R9935 VSS.n2223 VSS.n2222 0.0109167
R9936 VSS.n2237 VSS.n2236 0.0109167
R9937 VSS.n2251 VSS.n2250 0.0109167
R9938 VSS.n2267 VSS.n2266 0.0109167
R9939 VSS.n2281 VSS.n2280 0.0109167
R9940 VSS.n2295 VSS.n2294 0.0109167
R9941 VSS.n2309 VSS.n2308 0.0109167
R9942 VSS.n2321 VSS.n2320 0.0109167
R9943 VSS.n2335 VSS.n2334 0.0109167
R9944 VSS.n2348 VSS.n2347 0.0109167
R9945 VSS.n2351 VSS.n2350 0.0109167
R9946 VSS.n2364 VSS.n2363 0.0109167
R9947 VSS.n2377 VSS.n2376 0.0109167
R9948 VSS.n2391 VSS.n2390 0.0109167
R9949 VSS.n2405 VSS.n2404 0.0109167
R9950 VSS.n2418 VSS.n2417 0.0109167
R9951 VSS.n2432 VSS.n2431 0.0109167
R9952 VSS.n2446 VSS.n2445 0.0109167
R9953 VSS.n2460 VSS.n2459 0.0109167
R9954 VSS.n2474 VSS.n2473 0.0109167
R9955 VSS.n2490 VSS.n2489 0.0109167
R9956 VSS.n2504 VSS.n2503 0.0109167
R9957 VSS.n2518 VSS.n2517 0.0109167
R9958 VSS.n2532 VSS.n2531 0.0109167
R9959 VSS.n2546 VSS.n2545 0.0109167
R9960 VSS.n2560 VSS.n2559 0.0109167
R9961 VSS.n2574 VSS.n2573 0.0109167
R9962 VSS.n2588 VSS.n2587 0.0109167
R9963 VSS.n2602 VSS.n2601 0.0109167
R9964 VSS.n2618 VSS.n2617 0.0109167
R9965 VSS.n2632 VSS.n2631 0.0109167
R9966 VSS.n2646 VSS.n2645 0.0109167
R9967 VSS.n2660 VSS.n2659 0.0109167
R9968 VSS.n2672 VSS.n2671 0.0109167
R9969 VSS.n2686 VSS.n2685 0.0109167
R9970 VSS.n2699 VSS.n2698 0.0109167
R9971 VSS.n2702 VSS.n2701 0.0109167
R9972 VSS.n2715 VSS.n2714 0.0109167
R9973 VSS.n2728 VSS.n2727 0.0109167
R9974 VSS.n2742 VSS.n2741 0.0109167
R9975 VSS.n2756 VSS.n2755 0.0109167
R9976 VSS.n2769 VSS.n2768 0.0109167
R9977 VSS.n2783 VSS.n2782 0.0109167
R9978 VSS.n2797 VSS.n2796 0.0109167
R9979 VSS.n2811 VSS.n2810 0.0109167
R9980 VSS.n2825 VSS.n2824 0.0109167
R9981 VSS.n2841 VSS.n2840 0.0109167
R9982 VSS.n2855 VSS.n2854 0.0109167
R9983 VSS.n2869 VSS.n2868 0.0109167
R9984 VSS.n2883 VSS.n2882 0.0109167
R9985 VSS.n2897 VSS.n2896 0.0109167
R9986 VSS.n2911 VSS.n2910 0.0109167
R9987 VSS.n2925 VSS.n2924 0.0109167
R9988 VSS.n2939 VSS.n2938 0.0109167
R9989 VSS.n2953 VSS.n2952 0.0109167
R9990 VSS.n2969 VSS.n2968 0.0109167
R9991 VSS.n2983 VSS.n2982 0.0109167
R9992 VSS.n2997 VSS.n2996 0.0109167
R9993 VSS.n3011 VSS.n3010 0.0109167
R9994 VSS.n3023 VSS.n3022 0.0109167
R9995 VSS.n3037 VSS.n3036 0.0109167
R9996 VSS.n3053 VSS.n3052 0.0109167
R9997 VSS.n3055 VSS.n3054 0.0109167
R9998 VSS.n1092 VSS.n1080 0.00961458
R9999 VSS.n1078 VSS.n1066 0.00961458
R10000 VSS.n1064 VSS.n1052 0.00961458
R10001 VSS.n1050 VSS.n1036 0.00961458
R10002 VSS.n1034 VSS.n1022 0.00961458
R10003 VSS.n1020 VSS.n1008 0.00961458
R10004 VSS.n1006 VSS.n994 0.00961458
R10005 VSS.n992 VSS.n980 0.00961458
R10006 VSS.n978 VSS.n977 0.00961458
R10007 VSS.n975 VSS.n963 0.00961458
R10008 VSS.n961 VSS.n949 0.00961458
R10009 VSS.n947 VSS.n946 0.00961458
R10010 VSS.n944 VSS.n163 0.00961458
R10011 VSS.n185 VSS.n184 0.00961458
R10012 VSS.n930 VSS.n929 0.00961458
R10013 VSS.n927 VSS.n915 0.00961458
R10014 VSS.n913 VSS.n912 0.00961458
R10015 VSS.n910 VSS.n898 0.00961458
R10016 VSS.n896 VSS.n884 0.00961458
R10017 VSS.n882 VSS.n870 0.00961458
R10018 VSS.n868 VSS.n855 0.00961458
R10019 VSS.n853 VSS.n841 0.00961458
R10020 VSS.n839 VSS.n827 0.00961458
R10021 VSS.n825 VSS.n813 0.00961458
R10022 VSS.n811 VSS.n798 0.00961458
R10023 VSS.n796 VSS.n785 0.00961458
R10024 VSS.n783 VSS.n771 0.00961458
R10025 VSS.n769 VSS.n757 0.00961458
R10026 VSS.n755 VSS.n743 0.00961458
R10027 VSS.n741 VSS.n727 0.00961458
R10028 VSS.n725 VSS.n713 0.00961458
R10029 VSS.n711 VSS.n699 0.00961458
R10030 VSS.n697 VSS.n685 0.00961458
R10031 VSS.n683 VSS.n671 0.00961458
R10032 VSS.n669 VSS.n668 0.00961458
R10033 VSS.n666 VSS.n654 0.00961458
R10034 VSS.n652 VSS.n640 0.00961458
R10035 VSS.n638 VSS.n637 0.00961458
R10036 VSS.n635 VSS.n217 0.00961458
R10037 VSS.n239 VSS.n238 0.00961458
R10038 VSS.n621 VSS.n620 0.00961458
R10039 VSS.n618 VSS.n606 0.00961458
R10040 VSS.n604 VSS.n603 0.00961458
R10041 VSS.n601 VSS.n589 0.00961458
R10042 VSS.n587 VSS.n575 0.00961458
R10043 VSS.n573 VSS.n561 0.00961458
R10044 VSS.n559 VSS.n546 0.00961458
R10045 VSS.n544 VSS.n532 0.00961458
R10046 VSS.n530 VSS.n518 0.00961458
R10047 VSS.n516 VSS.n504 0.00961458
R10048 VSS.n502 VSS.n489 0.00961458
R10049 VSS.n487 VSS.n476 0.00961458
R10050 VSS.n474 VSS.n462 0.00961458
R10051 VSS.n460 VSS.n448 0.00961458
R10052 VSS.n446 VSS.n434 0.00961458
R10053 VSS.n432 VSS.n418 0.00961458
R10054 VSS.n416 VSS.n404 0.00961458
R10055 VSS.n402 VSS.n390 0.00961458
R10056 VSS.n388 VSS.n376 0.00961458
R10057 VSS.n374 VSS.n362 0.00961458
R10058 VSS.n360 VSS.n359 0.00961458
R10059 VSS.n357 VSS.n345 0.00961458
R10060 VSS.n343 VSS.n331 0.00961458
R10061 VSS.n329 VSS.n328 0.00961458
R10062 VSS.n326 VSS.n271 0.00961458
R10063 VSS.n313 VSS.n312 0.00961458
R10064 VSS.n310 VSS.n298 0.00961458
R10065 VSS.n296 VSS.n284 0.00961458
R10066 VSS.n3082 VSS.n3081 0.00961458
R10067 VSS.n3098 VSS.n3097 0.00961458
R10068 VSS.n3112 VSS.n3111 0.00961458
R10069 VSS.n3128 VSS.n3127 0.00961458
R10070 VSS.n3141 VSS.n3140 0.00961458
R10071 VSS.n3157 VSS.n3156 0.00961458
R10072 VSS.n3171 VSS.n3170 0.00961458
R10073 VSS.n3187 VSS.n3186 0.00961458
R10074 VSS.n3201 VSS.n3200 0.00961458
R10075 VSS.n3217 VSS.n3216 0.00961458
R10076 VSS.n3231 VSS.n3230 0.00961458
R10077 VSS.n3247 VSS.n3246 0.00961458
R10078 VSS.n3263 VSS.n3262 0.00961458
R10079 VSS.n3277 VSS.n3276 0.00961458
R10080 VSS.n3293 VSS.n3292 0.00961458
R10081 VSS.n3307 VSS.n3306 0.00961458
R10082 VSS.n3323 VSS.n3322 0.00961458
R10083 VSS.n3337 VSS.n3336 0.00961458
R10084 VSS.n3340 VSS.n3339 0.00961458
R10085 VSS.n3051 VSS.n3050 0.00701042
R10086 VSS.n11 VSS 0.00673818
R10087 VSS.n3050 VSS.n3049 0.00440625
R10088 VSS.n4104 VSS.n4103 0.00440625
R10089 VSS.n4101 VSS.n4098 0.00440625
R10090 VSS.n4096 VSS.n4084 0.00440625
R10091 VSS.n4082 VSS.n4071 0.00440625
R10092 VSS.n4069 VSS.n4068 0.00440625
R10093 VSS.n4066 VSS.n4056 0.00440625
R10094 VSS.n4054 VSS.n4042 0.00440625
R10095 VSS.n4040 VSS.n4028 0.00440625
R10096 VSS.n4026 VSS.n4014 0.00440625
R10097 VSS.n4012 VSS.n4011 0.00440625
R10098 VSS.n4009 VSS.n3999 0.00440625
R10099 VSS.n3997 VSS.n3985 0.00440625
R10100 VSS.n3983 VSS.n3971 0.00440625
R10101 VSS.n3969 VSS.n3957 0.00440625
R10102 VSS.n3955 VSS.n3942 0.00440625
R10103 VSS.n3940 VSS.n3928 0.00440625
R10104 VSS.n3926 VSS.n3913 0.00440625
R10105 VSS.n3911 VSS.n3899 0.00440625
R10106 VSS.n3897 VSS.n41 0.00440625
R10107 VSS.n3055 VSS.n3053 0.00180208
R10108 x4.X.n38 x4.X.n22 585
R10109 x4.X.n24 x4.X.t66 397.144
R10110 x4.X.n31 x4.X.t50 394.462
R10111 x4.X.n39 x4.X.n37 302.474
R10112 x4.X.n124 x4.X.t41 209.331
R10113 x4.X.n89 x4.X.t36 208.625
R10114 x4.X.n178 x4.X.t59 208.013
R10115 x4.X.n96 x4.X.t33 207.919
R10116 x4.X.n62 x4.X.t58 207.919
R10117 x4.X.n69 x4.X.t55 207.919
R10118 x4.X.n117 x4.X.t42 207.915
R10119 x4.X.n144 x4.X.t56 207.911
R10120 x4.X.n171 x4.X.t47 207.853
R10121 x4.X.n152 x4.X.t53 206.475
R10122 x4.X.n134 x4.X.t61 202.565
R10123 x4.X.n106 x4.X.t49 202.565
R10124 x4.X.n111 x4.X.t67 202.565
R10125 x4.X.n83 x4.X.t60 202.565
R10126 x4.X.n164 x4.X.t62 202.163
R10127 x4.X.n139 x4.X.t43 202.163
R10128 x4.X.n78 x4.X.t39 202.163
R10129 x4.X.n152 x4.X.t40 179.695
R10130 x4.X.n178 x4.X.t44 179.094
R10131 x4.X.n144 x4.X.t35 178.258
R10132 x4.X.n117 x4.X.t64 178.256
R10133 x4.X.n96 x4.X.t63 178.252
R10134 x4.X.n62 x4.X.t45 178.252
R10135 x4.X.n69 x4.X.t51 178.252
R10136 x4.X.n165 x4.X.t48 177.588
R10137 x4.X.n170 x4.X.t68 177.588
R10138 x4.X.n140 x4.X.t65 177.588
R10139 x4.X.n79 x4.X.t34 177.588
R10140 x4.X.n89 x4.X.t57 177.536
R10141 x4.X.n135 x4.X.t46 176.834
R10142 x4.X.n107 x4.X.t69 176.834
R10143 x4.X.n112 x4.X.t52 176.834
R10144 x4.X.n84 x4.X.t54 176.834
R10145 x4.X.n124 x4.X.t38 176.816
R10146 x4.X.n19 x4.X.n17 146.811
R10147 x4.X.n40 x4.X.n39 143.149
R10148 x4.X.n24 x4.X.t32 134.986
R10149 x4.X.n31 x4.X.t37 134.484
R10150 x4.X.n19 x4.X.n18 108.412
R10151 x4.X.n21 x4.X.n20 108.412
R10152 x4.X.n45 x4.X.n13 108.412
R10153 x4.X.n44 x4.X.n14 108.412
R10154 x4.X.n43 x4.X.n15 108.412
R10155 x4.X.n42 x4.X.n16 108.412
R10156 x4.X.n48 x4.X.n46 90.8321
R10157 x4.X.n48 x4.X.n47 52.4321
R10158 x4.X.n50 x4.X.n49 52.4321
R10159 x4.X.n52 x4.X.n51 52.4321
R10160 x4.X.n54 x4.X.n53 52.4321
R10161 x4.X.n56 x4.X.n55 52.4321
R10162 x4.X.n58 x4.X.n57 52.4321
R10163 x4.X.n60 x4.X.n59 52.4321
R10164 x4.X.n50 x4.X.n48 38.4005
R10165 x4.X.n52 x4.X.n50 38.4005
R10166 x4.X.n54 x4.X.n52 38.4005
R10167 x4.X.n56 x4.X.n54 38.4005
R10168 x4.X.n58 x4.X.n56 38.4005
R10169 x4.X.n60 x4.X.n58 38.4005
R10170 x4.X.n45 x4.X.n44 38.4005
R10171 x4.X.n44 x4.X.n43 38.4005
R10172 x4.X.n43 x4.X.n42 38.4005
R10173 x4.X.n21 x4.X.n19 38.4005
R10174 x4.X.n41 x4.X.n21 38.4005
R10175 x4.X.n42 x4.X.n41 38.4005
R10176 x4.X x4.X.n45 33.7342
R10177 x4.X.n181 x4.X.n60 30.8711
R10178 x4.X.n13 x4.X.t20 26.5955
R10179 x4.X.n13 x4.X.t26 26.5955
R10180 x4.X.n14 x4.X.t19 26.5955
R10181 x4.X.n14 x4.X.t30 26.5955
R10182 x4.X.n15 x4.X.t27 26.5955
R10183 x4.X.n15 x4.X.t18 26.5955
R10184 x4.X.n16 x4.X.t23 26.5955
R10185 x4.X.n16 x4.X.t16 26.5955
R10186 x4.X.n17 x4.X.t22 26.5955
R10187 x4.X.n17 x4.X.t17 26.5955
R10188 x4.X.n18 x4.X.t24 26.5955
R10189 x4.X.n18 x4.X.t28 26.5955
R10190 x4.X.n20 x4.X.t25 26.5955
R10191 x4.X.n20 x4.X.t29 26.5955
R10192 x4.X.n46 x4.X.t2 24.9236
R10193 x4.X.n46 x4.X.t13 24.9236
R10194 x4.X.n47 x4.X.t4 24.9236
R10195 x4.X.n47 x4.X.t8 24.9236
R10196 x4.X.n49 x4.X.t5 24.9236
R10197 x4.X.n49 x4.X.t9 24.9236
R10198 x4.X.n51 x4.X.t1 24.9236
R10199 x4.X.n51 x4.X.t11 24.9236
R10200 x4.X.n53 x4.X.t3 24.9236
R10201 x4.X.n53 x4.X.t12 24.9236
R10202 x4.X.n55 x4.X.t7 24.9236
R10203 x4.X.n55 x4.X.t14 24.9236
R10204 x4.X.n57 x4.X.t15 24.9236
R10205 x4.X.n57 x4.X.t10 24.9236
R10206 x4.X.n59 x4.X.t0 24.9236
R10207 x4.X.n59 x4.X.t6 24.9236
R10208 x4.X.n23 x4.X.t21 22.6555
R10209 x4.X.n180 x4.X.n179 19.9012
R10210 x4.X.n10 x4.X.n11 3.58524
R10211 x4.X.n181 x4.X.n180 19.6126
R10212 x4.X.n38 x4.X.t31 13.7905
R10213 x4.X.n27 x4.X 13.6005
R10214 x4.X.n39 x4.X.n38 12.8055
R10215 x4.X.n142 x4.X.n141 10.4992
R10216 x4.X.n114 x4.X.n113 10.4947
R10217 x4.X.n86 x4.X.n85 10.4903
R10218 x4.X.n41 x4.X.n40 9.82233
R10219 x4.X x4.X.n181 9.6005
R10220 x4.X.n8 x4.X.n7 1.83978
R10221 x4.X.n26 x4.X.n25 9.3005
R10222 x4.X.n33 x4.X.n32 9.3005
R10223 x4.X.n166 x4.X.n165 9.3005
R10224 x4.X.n136 x4.X.n135 9.3005
R10225 x4.X.n141 x4.X.n140 9.3005
R10226 x4.X.n108 x4.X.n107 9.3005
R10227 x4.X.n113 x4.X.n112 9.3005
R10228 x4.X.n80 x4.X.n79 9.3005
R10229 x4.X.n85 x4.X.n84 9.3005
R10230 x4.X.n35 x4.X.n22 9.3005
R10231 x4.X.n23 x4.X.n22 9.3005
R10232 x4.X.n179 x4.X 9.18311
R10233 x4.X.n179 x4.X.n178 8.76429
R10234 x4.X.n87 x4.X.n75 8.41509
R10235 x4.X.n40 x4.X.n22 8.16186
R10236 x4.X.n172 x4.X.n171 7.61316
R10237 x4.X.n135 x4.X.n134 7.35553
R10238 x4.X.n107 x4.X.n106 7.35553
R10239 x4.X.n112 x4.X.n111 7.35553
R10240 x4.X.n84 x4.X.n83 7.35553
R10241 x4.X.n153 x4.X.n152 7.32997
R10242 x4.X.n97 x4.X.n96 7.28785
R10243 x4.X.n63 x4.X.n62 7.28785
R10244 x4.X.n70 x4.X.n69 7.28785
R10245 x4.X.n118 x4.X.n117 7.27968
R10246 x4.X.n145 x4.X.n144 7.27145
R10247 x4.X.n90 x4.X.n89 7.25084
R10248 x4.X.n125 x4.X.n124 7.2225
R10249 x4.X.n32 x4.X.n31 6.9915
R10250 x4.X.n26 x4.X.n24 6.95412
R10251 x4.X.n165 x4.X.n164 6.95331
R10252 x4.X.n140 x4.X.n139 6.95331
R10253 x4.X.n79 x4.X.n78 6.95331
R10254 x4.X.n115 x4.X.n103 6.17402
R10255 x4.X.n143 x4.X.n131 6.14277
R10256 x4.X.n177 x4.X.n161 6.12937
R10257 x4.X.n142 x4.X.n136 6.09927
R10258 x4.X.n86 x4.X.n80 6.09034
R10259 x4.X.n176 x4.X.n175 5.93026
R10260 x4.X.n114 x4.X.n108 5.83458
R10261 x4.X.n146 x4.X 5.56572
R10262 x4.X.n154 x4.X 5.56572
R10263 x4.X.n119 x4.X 5.28746
R10264 x4.X.n126 x4.X 5.28746
R10265 x4.X.n91 x4.X 5.28746
R10266 x4.X.n132 x4.X 5.0092
R10267 x4.X.n98 x4.X 5.0092
R10268 x4.X.n76 x4.X 5.0092
R10269 x4.X.n81 x4.X 5.0092
R10270 x4.X.n64 x4.X 5.0092
R10271 x4.X.n71 x4.X 5.0092
R10272 x4.X.n162 x4.X 4.73093
R10273 x4.X.n172 x4.X.n169 4.73093
R10274 x4.X.n137 x4.X 4.73093
R10275 x4.X.n104 x4.X 4.73093
R10276 x4.X.n109 x4.X 4.73093
R10277 x4.X.n160 x4.X.n151 4.62479
R10278 x4.X.n102 x4.X.n94 4.61713
R10279 x4.X.n130 x4.X.n122 4.6082
R10280 x4.X.n75 x4.X.n67 4.6082
R10281 x4.X.n36 x4.X.n35 4.5327
R10282 x4.X.n12 x4.X.n22 9.31609
R10283 x4.X x4.X.n11 2.9629
R10284 x4.X.n163 x4.X.n162 4.45267
R10285 x4.X.n169 x4.X 4.45267
R10286 x4.X.n138 x4.X.n137 4.45267
R10287 x4.X.n105 x4.X.n104 4.45267
R10288 x4.X.n110 x4.X.n109 4.45267
R10289 x4.X.n176 x4.X.n166 4.42753
R10290 x4.X.n161 x4.X.n143 4.25884
R10291 x4.X.n131 x4.X.n115 4.24991
R10292 x4.X.n103 x4.X.n87 4.21866
R10293 x4.X.n133 x4.X.n132 4.17441
R10294 x4.X.n77 x4.X.n76 4.17441
R10295 x4.X.n82 x4.X.n81 4.17441
R10296 x4.X.n39 x4.X.n23 3.9405
R10297 x4.X.n147 x4.X.n146 3.61789
R10298 x4.X.n155 x4.X.n154 3.33963
R10299 x4.X.n120 x4.X.n119 3.33963
R10300 x4.X.n127 x4.X.n126 3.06137
R10301 x4.X.n92 x4.X.n91 3.06137
R10302 x4.X.n99 x4.X.n98 3.06137
R10303 x4.X.n65 x4.X.n64 3.06137
R10304 x4.X.n72 x4.X.n71 3.06137
R10305 x4.X.n149 x4.X.n147 3.04032
R10306 x4.X.n174 x4.X.n173 3.035
R10307 x4.X.n157 x4.X.n155 3.035
R10308 x4.X.n5 x4.X.n120 3.03311
R10309 x4.X.n0 x4.X.n127 3.03311
R10310 x4.X.n1 x4.X.n92 3.03311
R10311 x4.X.n2 x4.X.n99 3.03311
R10312 x4.X.n3 x4.X.n65 3.03311
R10313 x4.X.n4 x4.X.n72 3.03311
R10314 x4.X.n29 x4.X.n28 3.00943
R10315 x4.X.n8 x4.X 4.1629
R10316 x4.X.n37 x4.X.n9 2.62757
R10317 x4.X.n27 x4.X.n26 2.52171
R10318 x4.X.n32 x4.X.n8 1.54783
R10319 x4.X.n12 x4.X.n36 1.50334
R10320 x4.X.n87 x4.X.n86 2.2505
R10321 x4.X.n103 x4.X.n102 2.2505
R10322 x4.X.n115 x4.X.n114 2.2505
R10323 x4.X.n131 x4.X.n130 2.2505
R10324 x4.X.n143 x4.X.n142 2.2505
R10325 x4.X.n161 x4.X.n160 2.2505
R10326 x4.X.n177 x4.X.n176 2.2505
R10327 x4.X.n175 x4.X.n174 2.23927
R10328 x4.X.n34 x4.X.n9 2.23869
R10329 x4.X.n180 x4.X.n177 2.16478
R10330 x4.X.n160 x4.X.n159 2.07162
R10331 x4.X.n75 x4.X.n74 2.045
R10332 x4.X.n102 x4.X.n101 2.04053
R10333 x4.X.n130 x4.X.n129 2.02268
R10334 x4.X.n37 x4.X.n22 1.76715
R10335 x4.X.n29 x4.X 1.72692
R10336 x4.X.n127 x4.X.n125 1.67007
R10337 x4.X.n92 x4.X.n90 1.67007
R10338 x4.X.n99 x4.X.n97 1.67007
R10339 x4.X.n65 x4.X.n63 1.67007
R10340 x4.X.n72 x4.X.n70 1.67007
R10341 x4.X.n34 x4.X.n6 1.57957
R10342 x4.X.n7 x4.X.n6 0.896263
R10343 x4.X.n121 x4.X.n5 1.50237
R10344 x4.X.n128 x4.X.n0 1.50174
R10345 x4.X.n93 x4.X.n1 1.50174
R10346 x4.X.n100 x4.X.n2 1.50174
R10347 x4.X.n66 x4.X.n3 1.50174
R10348 x4.X.n73 x4.X.n4 1.50174
R10349 x4.X.n159 x4.X.n157 1.49811
R10350 x4.X.n151 x4.X.n149 1.49801
R10351 x4.X.n155 x4.X.n153 1.3918
R10352 x4.X.n120 x4.X.n118 1.3918
R10353 x4.X.n147 x4.X.n145 1.11354
R10354 x4.X.n171 x4.X.n170 0.72374
R10355 x4.X.n136 x4.X.n133 0.557022
R10356 x4.X.n80 x4.X.n77 0.557022
R10357 x4.X.n85 x4.X.n82 0.557022
R10358 x4.X.n27 x4.X.n11 0.300347
R10359 x4.X.n166 x4.X.n163 0.278761
R10360 x4.X.n173 x4.X.n172 0.278761
R10361 x4.X.n141 x4.X.n138 0.278761
R10362 x4.X.n108 x4.X.n105 0.278761
R10363 x4.X.n113 x4.X.n110 0.278761
R10364 x4.X.n28 x4.X 0.259429
R10365 x4.X.n28 x4.X.n10 0.076587
R10366 x4.X.n25 x4.X.n10 0.0466957
R10367 x4.X.n25 x4.X 0.0358261
R10368 x4.X.n7 x4.X.n33 0.0347909
R10369 x4.X.n175 x4.X.n167 0.0291789
R10370 x4.X.n36 x4.X.n34 0.0279871
R10371 x4.X.n122 x4.X.n121 0.0269367
R10372 x4.X.n94 x4.X.n93 0.0269367
R10373 x4.X.n67 x4.X.n66 0.0269367
R10374 x4.X.n129 x4.X.n128 0.0257706
R10375 x4.X.n101 x4.X.n100 0.0257706
R10376 x4.X.n74 x4.X.n73 0.0257706
R10377 x4.X.n6 x4.X.n30 4.51062
R10378 x4.X.n5 x4.X.n116 0.0271977
R10379 x4.X.n4 x4.X.n68 0.0259313
R10380 x4.X.n3 x4.X.n61 0.0259313
R10381 x4.X.n2 x4.X.n95 0.0259313
R10382 x4.X.n1 x4.X.n88 0.0259313
R10383 x4.X.n0 x4.X.n123 0.0259313
R10384 x4.X.n149 x4.X.n148 0.0245385
R10385 x4.X.n9 x4.X.n12 0.00855895
R10386 x4.X.n33 x4.X.n30 0.0217264
R10387 x4.X.n157 x4.X.n156 0.0213333
R10388 x4.X.n30 x4.X 0.0170094
R10389 x4.X.n159 x4.X.n158 0.016693
R10390 x4.X.n174 x4.X.n168 0.0152198
R10391 x4.X.n151 x4.X.n150 0.0144347
R10392 x4.X.n35 x4.X.n9 0.0109693
R10393 x4.X x4.X.n29 0.00993396
R10394 check[5].n1 check[5].t3 331.51
R10395 check[5].n1 check[5].t2 209.403
R10396 check[5].n0 check[5].t1 207.373
R10397 check[5].n2 check[5].n1 76.0005
R10398 check[5].n4 check[5].n3 50.8596
R10399 check[5].n5 check[5].t0 31.153
R10400 check[5].n4 check[5] 18.2949
R10401 check[5].n3 check[5] 13.2142
R10402 check[5].n3 check[5] 12.3082
R10403 check[5] check[5].n0 9.01934
R10404 check[5] check[5].n2 8.58587
R10405 check[5] check[5].n5 7.78567
R10406 check[5].n0 check[5] 7.45876
R10407 check[5].n2 check[5] 2.02977
R10408 check[5].n5 check[5].n4 1.33351
R10409 check[0].n3 check[0].t5 373.283
R10410 check[0].n1 check[0].t3 331.51
R10411 check[0].n1 check[0].t2 209.403
R10412 check[0].n0 check[0].t1 207.373
R10413 check[0].n3 check[0].t4 132.282
R10414 check[0].n4 check[0].n3 84.146
R10415 check[0].n2 check[0].n1 76.0005
R10416 check[0].n8 check[0].n7 48.6767
R10417 check[0].n9 check[0].t0 33.3302
R10418 check[0].n6 check[0].n5 19.508
R10419 check[0].n8 check[0] 15.1737
R10420 check[0].n5 check[0].n4 13.3958
R10421 check[0].n7 check[0] 12.062
R10422 check[0] check[0].n9 9.55531
R10423 check[0] check[0].n0 9.01934
R10424 check[0].n6 check[0] 8.69451
R10425 check[0] check[0].n2 8.58587
R10426 check[0].n0 check[0] 7.45876
R10427 check[0].n5 check[0] 6.84701
R10428 check[0].n4 check[0] 4.07323
R10429 check[0].n7 check[0].n6 3.04048
R10430 check[0].n2 check[0] 2.02977
R10431 check[0].n9 check[0].n8 1.77306
R10432 check[2].n3 check[2].t5 331.51
R10433 check[2].n1 check[2].t3 299.377
R10434 check[2].n3 check[2].t4 209.403
R10435 check[2].n0 check[2].t1 207.373
R10436 check[2].n1 check[2].t2 206.19
R10437 check[2] check[2].n1 105.007
R10438 check[2].n4 check[2].n3 76.0005
R10439 check[2].n7 check[2].n6 49.7951
R10440 check[2].n5 check[2].n2 47.9541
R10441 check[2].n8 check[2].t0 31.8695
R10442 check[2].n7 check[2] 15.2244
R10443 check[2].n6 check[2] 11.8159
R10444 check[2].n2 check[2] 11.1489
R10445 check[2] check[2].n0 9.01934
R10446 check[2] check[2].n8 8.9196
R10447 check[2].n5 check[2] 8.84542
R10448 check[2] check[2].n4 8.58587
R10449 check[2].n0 check[2] 7.45876
R10450 check[2].n6 check[2].n5 3.04357
R10451 check[2].n2 check[2] 2.89082
R10452 check[2].n4 check[2] 2.02977
R10453 check[2].n8 check[2].n7 1.63044
R10454 D[2].n3 D[2].t2 269.921
R10455 D[2].n3 D[2].t3 234.573
R10456 D[2].n10 D[2].t1 207.373
R10457 D[2].n11 D[2] 59.1407
R10458 D[2].n13 D[2].t0 32.581
R10459 D[2] D[2].n13 9.80687
R10460 D[2] D[2].n10 9.01934
R10461 D[2].n4 D[2].n3 8.76429
R10462 D[2].n4 D[2] 7.57233
R10463 D[2].n10 D[2] 7.45876
R10464 D[2].n4 D[2] 4.68782
R10465 D[2].n12 D[2].n11 3.84831
R10466 D[2].n5 D[2].n4 3.77218
R10467 D[2].n6 D[2].n5 3.26839
R10468 D[2].n5 D[2] 3.23635
R10469 D[2].n11 D[2].n9 2.92915
R10470 D[2].n8 D[2].n1 2.26284
R10471 D[2].n7 D[2].n6 2.23869
R10472 D[2].n13 D[2].n12 0.389891
R10473 D[2].n7 D[2].n2 0.0232273
R10474 D[2].n9 D[2].n0 0.00807576
R10475 D[2].n8 D[2].n7 0.00195195
R10476 D[2].n9 D[2].n8 0.00194159
R10477 x5.X.n9 x5.X.t20 269.921
R10478 x5.X.n50 x5.X.t10 267.291
R10479 x5.X.n35 x5.X.t13 267.291
R10480 x5.X.n20 x5.X.t9 267.291
R10481 x5.X.n66 x5.X.t8 265.538
R10482 x5.X.n58 x5.X.t19 265.538
R10483 x5.X.n43 x5.X.t18 265.538
R10484 x5.X.n28 x5.X.t17 265.538
R10485 x5.X.n13 x5.X.t11 264.663
R10486 x5.X.n9 x5.X.t7 234.573
R10487 x5.X.n15 x5.X.t16 224.934
R10488 x5.X.n68 x5.X.t12 224.058
R10489 x5.X.n60 x5.X.t6 224.058
R10490 x5.X.n45 x5.X.t5 224.058
R10491 x5.X.n30 x5.X.t4 224.058
R10492 x5.X.n52 x5.X.t15 222.304
R10493 x5.X.n37 x5.X.t21 222.304
R10494 x5.X.n22 x5.X.t14 222.304
R10495 x5.X.n6 x5.X.n5 143.643
R10496 x5.X.n8 x5.X.n7 92.5005
R10497 x5.X.n10 x5.X.n9 76.0005
R10498 x5.X.n73 x5.X.n72 72.3248
R10499 x5.X.n73 x5.X.n8 36.1417
R10500 x5.X x5.X.n73 32.377
R10501 x5.X.n5 x5.X.t2 26.5955
R10502 x5.X.n5 x5.X.t3 26.5955
R10503 x5.X.n7 x5.X.t1 24.9236
R10504 x5.X.n7 x5.X.t0 24.9236
R10505 x5.X.n25 x5.X 21.2667
R10506 x5.X.n52 x5.X.n51 12.2696
R10507 x5.X.n37 x5.X.n36 12.2696
R10508 x5.X.n22 x5.X.n21 12.2696
R10509 x5.X.n40 x5.X.n25 10.5535
R10510 x5.X.n55 x5.X.n40 10.5535
R10511 x5.X.n68 x5.X.n67 10.5169
R10512 x5.X.n60 x5.X.n59 10.5169
R10513 x5.X.n45 x5.X.n44 10.5169
R10514 x5.X.n30 x5.X.n29 10.5169
R10515 x5.X.n63 x5.X.n55 10.4999
R10516 x5.X.n15 x5.X.n14 9.6405
R10517 x5.X.n46 x5.X.n45 9.3005
R10518 x5.X.n31 x5.X.n30 9.3005
R10519 x5.X x5.X.n6 9.02598
R10520 x5.X.n69 x5.X.n68 8.76429
R10521 x5.X.n61 x5.X.n60 8.76429
R10522 x5.X.n53 x5.X.n52 8.76429
R10523 x5.X.n38 x5.X.n37 8.76429
R10524 x5.X.n16 x5.X.n15 8.76429
R10525 x5.X.n23 x5.X.n22 8.76429
R10526 x5.X.n6 x5.X 7.64268
R10527 x5.X.n72 x5.X.n63 7.58473
R10528 x5.X x5.X.n10 7.57233
R10529 x5.X.n1 x5.X.n54 7.52485
R10530 x5.X.n2 x5.X.n24 7.5187
R10531 x5.X.n0 x5.X.n39 7.45404
R10532 x5.X.n72 x5.X.n4 7.19295
R10533 x5.X.n48 x5.X 7.03149
R10534 x5.X.n33 x5.X 7.03149
R10535 x5.X.n18 x5.X 7.03149
R10536 x5.X.n64 x5.X 6.67092
R10537 x5.X.n56 x5.X 6.67092
R10538 x5.X.n41 x5.X 6.67092
R10539 x5.X.n26 x5.X 6.67092
R10540 x5.X.n63 x5.X.n62 6.55969
R10541 x5.X.n11 x5.X 6.49064
R10542 x5.X.n8 x5.X 5.27109
R10543 x5.X.n4 x5.X.n70 5.26654
R10544 x5.X.n14 x5.X.n13 5.25868
R10545 x5.X.n10 x5.X 4.68782
R10546 x5.X.n40 x5.X.n0 4.38498
R10547 x5.X.n67 x5.X.n66 4.38232
R10548 x5.X.n59 x5.X.n58 4.38232
R10549 x5.X.n44 x5.X.n43 4.38232
R10550 x5.X.n29 x5.X.n28 4.38232
R10551 x5.X.n55 x5.X.n1 4.38051
R10552 x5.X.n25 x5.X.n3 4.35575
R10553 x5.X.n3 x5.X.n17 5.18552
R10554 x5.X.n0 x5.X.n32 3.49645
R10555 x5.X.n1 x5.X.n47 3.4947
R10556 x5.X.n51 x5.X.n50 2.62959
R10557 x5.X.n36 x5.X.n35 2.62959
R10558 x5.X.n21 x5.X.n20 2.62959
R10559 x5.X.n53 x5.X.n49 2.52444
R10560 x5.X.n38 x5.X.n34 2.52444
R10561 x5.X.n23 x5.X.n19 2.52444
R10562 x5.X.n70 x5.X.n69 2.27475
R10563 x5.X.n4 x5.X.n71 2.26611
R10564 x5.X.n17 x5.X.n16 2.20216
R10565 x5.X.n69 x5.X.n65 2.16388
R10566 x5.X.n61 x5.X.n57 2.16388
R10567 x5.X.n46 x5.X.n42 2.16388
R10568 x5.X.n31 x5.X.n27 2.16388
R10569 x5.X.n16 x5.X.n12 1.9836
R10570 x5.X.n32 x5.X.n31 1.45136
R10571 x5.X.n47 x5.X.n46 1.38585
R10572 x5.X.n12 x5.X.n11 1.08219
R10573 x5.X.n62 x5.X.n61 1.0658
R10574 x5.X.n62 x5.X 0.932428
R10575 x5.X.n54 x5.X 0.930853
R10576 x5.X.n24 x5.X 0.919788
R10577 x5.X.n39 x5.X 0.919522
R10578 x5.X.n65 x5.X.n64 0.901908
R10579 x5.X.n57 x5.X.n56 0.901908
R10580 x5.X.n42 x5.X.n41 0.901908
R10581 x5.X.n27 x5.X.n26 0.901908
R10582 x5.X.n39 x5.X.n38 0.850177
R10583 x5.X.n24 x5.X.n23 0.849917
R10584 x5.X.n54 x5.X.n53 0.843446
R10585 x5.X.n47 x5.X 0.801859
R10586 x5.X.n32 x5.X 0.71223
R10587 x5.X.n49 x5.X.n48 0.541345
R10588 x5.X.n34 x5.X.n33 0.541345
R10589 x5.X.n19 x5.X.n18 0.541345
R10590 x5.X.n17 x5.X 0.469125
R10591 x5.X.n70 x5.X 0.242354
R10592 x5.X.n3 x5.X.n2 0.0819394
R10593 comparator_out.n26 comparator_out.t3 331.51
R10594 comparator_out.n24 comparator_out.t12 331.51
R10595 comparator_out.n16 comparator_out.t8 331.51
R10596 comparator_out.n3 comparator_out.t9 331.51
R10597 comparator_out.n0 comparator_out.t10 331.51
R10598 comparator_out.n35 comparator_out.t1 331.51
R10599 comparator_out.n18 comparator_out.t4 328.832
R10600 comparator_out.n9 comparator_out.t2 328.832
R10601 comparator_out.n26 comparator_out.t15 209.403
R10602 comparator_out.n24 comparator_out.t11 209.403
R10603 comparator_out.n16 comparator_out.t5 209.403
R10604 comparator_out.n3 comparator_out.t6 209.403
R10605 comparator_out.n0 comparator_out.t7 209.403
R10606 comparator_out.n35 comparator_out.t13 209.403
R10607 comparator_out.n20 comparator_out.t0 196.906
R10608 comparator_out.n7 comparator_out.t14 196.906
R10609 comparator_out comparator_out.n20 152.156
R10610 comparator_out.n7 comparator_out 152.156
R10611 comparator_out.n27 comparator_out.n26 76.0005
R10612 comparator_out.n25 comparator_out.n24 76.0005
R10613 comparator_out.n17 comparator_out.n16 76.0005
R10614 comparator_out.n4 comparator_out.n3 76.0005
R10615 comparator_out.n1 comparator_out.n0 76.0005
R10616 comparator_out.n36 comparator_out.n35 76.0005
R10617 comparator_out comparator_out.n34 16.15
R10618 comparator_out.n20 comparator_out.n19 12.4968
R10619 comparator_out.n8 comparator_out.n7 12.4968
R10620 comparator_out.n28 comparator_out 11.3477
R10621 comparator_out.n29 comparator_out.n28 10.4895
R10622 comparator_out.n33 comparator_out 9.2369
R10623 comparator_out.n31 comparator_out 9.08527
R10624 comparator_out.n28 comparator_out 8.93363
R10625 comparator_out.n22 comparator_out.n18 8.76429
R10626 comparator_out.n10 comparator_out.n9 8.76429
R10627 comparator_out comparator_out.n27 8.58587
R10628 comparator_out comparator_out.n25 8.58587
R10629 comparator_out comparator_out.n17 8.58587
R10630 comparator_out comparator_out.n4 8.58587
R10631 comparator_out comparator_out.n36 8.58587
R10632 comparator_out.n29 comparator_out 8.4832
R10633 comparator_out.n2 comparator_out 7.80538
R10634 comparator_out.n34 comparator_out.n2 7.58034
R10635 comparator_out.n23 comparator_out 7.07644
R10636 comparator_out.n31 comparator_out.n30 6.98058
R10637 comparator_out.n33 comparator_out.n32 6.97165
R10638 comparator_out.n11 comparator_out 6.73582
R10639 comparator_out.n30 comparator_out.n23 6.01572
R10640 comparator_out.n32 comparator_out.n15 3.78933
R10641 comparator_out.n34 comparator_out.n33 3.51183
R10642 comparator_out.n30 comparator_out.n29 3.43148
R10643 comparator_out.n32 comparator_out.n31 3.41362
R10644 comparator_out.n19 comparator_out.n18 2.67828
R10645 comparator_out.n9 comparator_out.n8 2.67828
R10646 comparator_out.n12 comparator_out.n11 2.61902
R10647 comparator_out.n27 comparator_out 2.02977
R10648 comparator_out.n25 comparator_out 2.02977
R10649 comparator_out.n21 comparator_out 2.02977
R10650 comparator_out.n17 comparator_out 2.02977
R10651 comparator_out comparator_out.n6 2.02977
R10652 comparator_out.n4 comparator_out 2.02977
R10653 comparator_out.n1 comparator_out 2.02977
R10654 comparator_out.n36 comparator_out 2.02977
R10655 comparator_out.n14 comparator_out.n13 1.50871
R10656 comparator_out.n11 comparator_out.n10 1.08449
R10657 comparator_out.n2 comparator_out.n1 0.780988
R10658 comparator_out.n23 comparator_out.n22 0.605202
R10659 comparator_out.n22 comparator_out.n21 0.468793
R10660 comparator_out.n10 comparator_out.n6 0.468793
R10661 comparator_out.n12 comparator_out.n5 0.0341538
R10662 comparator_out.n15 comparator_out.n14 0.0226928
R10663 comparator_out.n13 comparator_out.n12 0.00372631
R10664 check[3].n7 check[3].t1 417.519
R10665 check[3].n1 check[3].t3 331.51
R10666 check[3].n1 check[3].t2 209.403
R10667 check[3].t1 check[3].n6 137.702
R10668 check[3].n2 check[3].n1 76.0005
R10669 check[3].n8 check[3] 60.7393
R10670 check[3].n9 check[3].t0 35.4919
R10671 check[3].n8 check[3] 18.329
R10672 check[3].n7 check[3].n0 12.3082
R10673 check[3].n3 check[3] 12.0607
R10674 check[3] check[3].n9 9.48284
R10675 check[3].n4 check[3].n0 9.3005
R10676 check[3].n6 check[3].n3 9.3005
R10677 check[3] check[3].n2 8.58587
R10678 check[3].n5 check[3].n4 4.59955
R10679 check[3] check[3].n0 2.70819
R10680 check[3].n2 check[3] 2.02977
R10681 check[3].n9 check[3].n8 1.84729
R10682 check[3] check[3].n7 1.72358
R10683 check[3].n5 check[3] 1.353
R10684 check[3].n6 check[3].n5 0.122715
R10685 check[3].n4 check[3].n3 0.00847872
R10686 check[6].n3 check[6].t3 331.51
R10687 check[6].n3 check[6].t2 209.403
R10688 check[6].n2 check[6].t1 207.373
R10689 check[6].n4 check[6].n3 76.0005
R10690 check[6].n6 check[6].n5 48.5667
R10691 check[6].n9 check[6].t0 31.8564
R10692 check[6].n0 check[6] 16.649
R10693 check[6].n5 check[6] 13.5264
R10694 check[6].n5 check[6] 11.8159
R10695 check[6] check[6].n2 9.01934
R10696 check[6] check[6].n9 8.94887
R10697 check[6] check[6].n4 8.58587
R10698 check[6].n2 check[6] 7.45876
R10699 check[6].n6 check[6].n1 4.3624
R10700 check[6].n8 check[6].n7 2.95435
R10701 check[6].n4 check[6] 2.02977
R10702 check[6].n7 check[6].n6 0.578192
R10703 check[6].n9 check[6].n8 0.290433
R10704 check[6].n1 check[6].n0 0.0421667
R10705 D[1].n8 D[1].t2 269.921
R10706 D[1].n8 D[1].t3 234.573
R10707 D[1].n7 D[1].t1 207.373
R10708 D[1].n9 D[1].n8 76.0005
R10709 D[1].n13 D[1].t0 33.3405
R10710 D[1].n11 D[1].n10 23.4
R10711 D[1].n10 D[1] 22.0971
R10712 D[1].n10 D[1].n9 14.9338
R10713 D[1] D[1].n13 9.32876
R10714 D[1] D[1].n7 9.01934
R10715 D[1].n9 D[1] 7.57233
R10716 D[1].n7 D[1] 7.45876
R10717 D[1].n3 D[1] 6.54947
R10718 D[1].n9 D[1] 4.68782
R10719 D[1].n12 D[1].n11 3.67573
R10720 D[1].n11 D[1].n6 2.87957
R10721 D[1].n5 D[1].n1 2.26284
R10722 D[1].n4 D[1].n3 2.23869
R10723 D[1].n13 D[1].n12 0.391757
R10724 D[1].n4 D[1].n2 0.0213333
R10725 D[1].n6 D[1].n0 0.0099697
R10726 D[1].n5 D[1].n4 0.00195195
R10727 D[1].n6 D[1].n5 0.00194159
R10728 reset.n0 reset.t0 259.634
R10729 reset.n0 reset.t1 175.183
R10730 reset.n1 reset.n0 8.19557
R10731 reset.n1 reset 2.53088
R10732 reset reset.n1 2.48048
R10733 check[4].n1 check[4].t3 331.51
R10734 check[4].n1 check[4].t2 209.403
R10735 check[4].n0 check[4].t1 207.373
R10736 check[4].n2 check[4].n1 76.0005
R10737 check[4].n4 check[4].n3 48.1851
R10738 check[4].n5 check[4].t0 34.0601
R10739 check[4].n4 check[4] 18.3315
R10740 check[4].n3 check[4] 13.0581
R10741 check[4].n3 check[4] 12.5543
R10742 check[4] check[4].n5 9.53084
R10743 check[4] check[4].n0 9.01934
R10744 check[4] check[4].n2 8.58587
R10745 check[4].n0 check[4] 7.45876
R10746 check[4].n2 check[4] 2.02977
R10747 check[4].n5 check[4].n4 1.79774
R10748 D[5].n8 D[5].t2 269.921
R10749 D[5].n8 D[5].t3 234.573
R10750 D[5].n7 D[5].t1 207.373
R10751 D[5].n9 D[5].n8 76.0005
R10752 D[5].n14 D[5].t0 34.8263
R10753 D[5].n11 D[5] 23.5855
R10754 D[5].n12 D[5].n11 23.0768
R10755 D[5].n11 D[5].n10 14.6672
R10756 D[5] D[5].n7 9.01934
R10757 D[5] D[5].n14 8.60331
R10758 D[5].n9 D[5] 7.57233
R10759 D[5].n7 D[5] 7.45876
R10760 D[5].n10 D[5] 3.78642
R10761 D[5].n13 D[5].n12 3.14374
R10762 D[5].n3 D[5] 3.01822
R10763 D[5].n12 D[5].n6 2.74043
R10764 D[5].n5 D[5].n1 2.26284
R10765 D[5].n4 D[5].n3 2.23869
R10766 D[5].n10 D[5].n9 0.901908
R10767 D[5].n14 D[5].n13 0.398471
R10768 D[5].n6 D[5].n0 0.0232273
R10769 D[5].n4 D[5].n2 0.00807576
R10770 D[5].n5 D[5].n4 0.00195195
R10771 D[5].n6 D[5].n5 0.00194159
R10772 D[4].n8 D[4].t2 269.921
R10773 D[4].n8 D[4].t3 234.573
R10774 D[4].n7 D[4].t1 207.373
R10775 D[4].n9 D[4].n8 76.0005
R10776 D[4].n14 D[4].t0 33.3509
R10777 D[4].n11 D[4] 23.2878
R10778 D[4].n12 D[4].n11 22.7446
R10779 D[4].n11 D[4].n10 14.6672
R10780 D[4] D[4].n14 9.10171
R10781 D[4] D[4].n7 9.01934
R10782 D[4].n9 D[4] 7.57233
R10783 D[4].n7 D[4] 7.45876
R10784 D[4].n10 D[4] 3.9667
R10785 D[4].n13 D[4].n12 3.32332
R10786 D[4].n12 D[4].n6 2.78529
R10787 D[4].n3 D[4] 2.75482
R10788 D[4].n5 D[4].n1 2.26284
R10789 D[4].n4 D[4].n3 2.23869
R10790 D[4].n10 D[4].n9 0.721627
R10791 D[4].n14 D[4].n13 0.379298
R10792 D[4].n6 D[4].n0 0.0251212
R10793 D[4].n4 D[4].n2 0.00618182
R10794 D[4].n5 D[4].n4 0.00195195
R10795 D[4].n6 D[4].n5 0.00194159
R10796 sel_bit[1].t1 sel_bit[1].t3 769.593
R10797 sel_bit[1].n4 sel_bit[1].t2 367.928
R10798 sel_bit[1].n2 sel_bit[1].t1 339.695
R10799 sel_bit[1].n4 sel_bit[1].t0 112.237
R10800 sel_bit[1].n5 sel_bit[1].n4 22.0348
R10801 sel_bit[1].n7 sel_bit[1] 15.3177
R10802 sel_bit[1].n5 sel_bit[1].n3 12.3948
R10803 sel_bit[1].n3 sel_bit[1].n2 11.0176
R10804 sel_bit[1].n6 sel_bit[1].n5 8.76429
R10805 sel_bit[1].n0 sel_bit[1] 5.95912
R10806 sel_bit[1] sel_bit[1].n7 3.41725
R10807 sel_bit[1].n6 sel_bit[1].n1 1.98671
R10808 sel_bit[1].n1 sel_bit[1].n0 1.76602
R10809 sel_bit[1].n7 sel_bit[1].n6 1.07617
R10810 D[7].n0 D[7].t1 207.373
R10811 D[7].n1 D[7] 66.6056
R10812 D[7].n1 D[7].t0 34.2054
R10813 D[7] D[7].n0 9.01934
R10814 D[7].n0 D[7] 7.45876
R10815 D[7].n10 D[7].n9 4.18512
R10816 D[7].n9 D[7].n8 3.02821
R10817 D[7].n4 D[7] 2.91107
R10818 D[7].n6 D[7].n2 2.26284
R10819 D[7].n5 D[7].n4 2.23869
R10820 D[7] D[7].n10 2.21588
R10821 D[7].n9 D[7].n1 0.253183
R10822 D[7].n8 D[7].n7 0.00901436
R10823 D[7].n5 D[7].n3 0.00618182
R10824 D[7].n6 D[7].n5 0.00195195
R10825 D[7].n7 D[7].n6 0.00194159
R10826 D[6].n8 D[6].t2 269.921
R10827 D[6].n8 D[6].t3 234.573
R10828 D[6].n7 D[6].t1 207.373
R10829 D[6].n9 D[6].n8 76.0005
R10830 D[6].n14 D[6].t0 34.0928
R10831 D[6].n11 D[6] 24.4785
R10832 D[6].n12 D[6].n11 21.9377
R10833 D[6].n11 D[6].n10 14.6672
R10834 D[6] D[6].n7 9.01934
R10835 D[6] D[6].n14 8.85188
R10836 D[6].n9 D[6] 7.57233
R10837 D[6].n7 D[6] 7.45876
R10838 D[6].n10 D[6] 3.24557
R10839 D[6].n13 D[6].n12 3.14374
R10840 D[6].n3 D[6] 3.01375
R10841 D[6].n12 D[6].n6 2.74043
R10842 D[6].n5 D[6].n1 2.26284
R10843 D[6].n4 D[6].n3 2.23869
R10844 D[6].n10 D[6].n9 1.44275
R10845 D[6].n14 D[6].n13 0.389863
R10846 D[6].n6 D[6].n0 0.0232273
R10847 D[6].n4 D[6].n2 0.00807576
R10848 D[6].n5 D[6].n4 0.00195195
R10849 D[6].n6 D[6].n5 0.00194159
R10850 sel_bit[0].n4 sel_bit[0].t2 445.048
R10851 sel_bit[0].n12 sel_bit[0].t0 432.193
R10852 sel_bit[0].n7 sel_bit[0].t4 287.995
R10853 sel_bit[0].n12 sel_bit[0].t3 254.389
R10854 sel_bit[0].n2 sel_bit[0].t1 252.248
R10855 sel_bit[0].n7 sel_bit[0].t5 194.809
R10856 sel_bit[0].n4 sel_bit[0].n3 152
R10857 sel_bit[0].n2 sel_bit[0].n1 152
R10858 sel_bit[0].n13 sel_bit[0].n12 76.0005
R10859 sel_bit[0].n8 sel_bit[0].n7 76.0005
R10860 sel_bit[0] sel_bit[0].n8 20.2672
R10861 sel_bit[0].n6 sel_bit[0].n5 15.6271
R10862 sel_bit[0].n5 sel_bit[0].n4 14.4605
R10863 sel_bit[0].n5 sel_bit[0].n2 12.8538
R10864 sel_bit[0].n14 sel_bit[0].n13 9.16815
R10865 sel_bit[0].n3 sel_bit[0] 9.03579
R10866 sel_bit[0].n13 sel_bit[0] 6.21226
R10867 sel_bit[0].n1 sel_bit[0] 5.64756
R10868 sel_bit[0].n10 sel_bit[0].n6 5.18664
R10869 sel_bit[0].n6 sel_bit[0].n0 4.88604
R10870 sel_bit[0].n9 sel_bit[0] 4.77729
R10871 sel_bit[0].n11 sel_bit[0] 4.25943
R10872 sel_bit[0].n8 sel_bit[0] 3.91161
R10873 sel_bit[0].n3 sel_bit[0].n0 3.01226
R10874 sel_bit[0].n1 sel_bit[0].n0 0.753441
R10875 sel_bit[0].n9 sel_bit[0] 0.563
R10876 sel_bit[0].n11 sel_bit[0] 0.259429
R10877 sel_bit[0].n10 sel_bit[0].n9 0.101633
R10878 sel_bit[0].n14 sel_bit[0].n11 0.0793043
R10879 sel_bit[0] sel_bit[0].n14 0.0793043
R10880 sel_bit[0] sel_bit[0].n10 0.0588664
R10881 clk_sar.n0 clk_sar.t0 259.031
R10882 clk_sar.n0 clk_sar.t1 175.778
R10883 clk_sar.n1 clk_sar.n0 8.08213
R10884 clk_sar.n1 clk_sar 4.54939
R10885 clk_sar clk_sar.n1 2.70993
C0 a_9322_3521# x42.Q_N 0.00203f
C1 a_6709_3521# VDD 0.00984f
C2 a_8402_3239# a_9322_3521# 1.09e-19
C3 x33.Q_N a_8803_4112# 2.89e-22
C4 a_8857_3213# a_9101_3521# 0.0104f
C5 a_7185_2366# x30.Q_N 0.0403f
C6 a_9151_3213# check[4] 1.06e-19
C7 a_9638_3213# a_10346_4801# 3.19e-20
C8 a_5561_3239# VDD 0.19f
C9 a_8998_4801# a_9370_4801# 3.34e-19
C10 a_3618_3239# x27.Q_N 3.65e-19
C11 x77.Y check[6] 3.89e-20
C12 x4.X a_6985_4112# 6.8e-19
C13 a_6375_3605# x4.X 9.07e-19
C14 a_3900_5167# a_3913_4112# 2.81e-19
C15 a_4368_4775# a_3600_4086# 0.0018f
C16 a_6845_4386# a_9238_4086# 2.9e-21
C17 a_4074_4775# a_4155_4086# 8.83e-20
C18 a_3619_4801# a_4453_4386# 7.24e-20
C19 a_3453_4801# a_4454_4086# 1.15e-19
C20 x45.Q_N a_8384_4086# 5.27e-21
C21 x20.Q_N a_4155_4086# 2.32e-19
C22 a_6410_2366# a_6780_2366# 4.11e-20
C23 check[0] a_6505_4394# 9.42e-20
C24 VDD a_4681_4801# 0.346f
C25 D[1] a_11543_3213# 1.24e-19
C26 a_9638_3213# a_9709_2550# 1.66e-21
C27 a_9464_3239# a_9441_2340# 1.03e-19
C28 a_6400_4801# check[5] 5.31e-21
C29 a_8938_2340# check[4] 1.33e-19
C30 VDD a_11857_4801# 0.343f
C31 a_11543_3213# a_11544_4775# 0.00121f
C32 a_2060_2640# eob 1.44e-19
C33 check[4] a_11184_4801# 9.44e-20
C34 a_5170_4478# a_5372_4112# 8.94e-19
C35 x77.Y a_3912_2366# 7.49e-20
C36 a_4019_4112# a_4389_4112# 4.11e-20
C37 x4.X a_3900_5167# 0.00135f
C38 a_10345_3239# x4.X 0.00275f
C39 a_7317_2550# x4.X 0.00147f
C40 check[2] a_5845_4801# 1.76e-19
C41 x4.X a_11076_5167# 0.00135f
C42 x77.Y a_4317_3521# 4.28e-20
C43 a_5089_5083# x27.Q_N 2.02e-20
C44 a_9237_2340# a_9441_2340# 0.117f
C45 a_9236_2640# a_9709_2550# 0.145f
C46 a_8938_2340# x60.Q_N 9.58e-21
C47 a_11856_3239# x66.Q_N 9.58e-21
C48 comparator_out a_5896_2340# 7.85e-19
C49 check[1] a_8803_4112# 4.26e-19
C50 a_9237_2340# x36.Q_N 1.55e-19
C51 a_11565_4112# VDD 3.47e-19
C52 a_12265_5083# x36.Q_N 2.02e-20
C53 D[7] x4.X 0.00353f
C54 check[2] a_8384_4086# 6.25e-20
C55 x5.X a_7562_4478# 1.85e-19
C56 sel_bit[0] a_2788_5674# 3.68e-19
C57 VDD a_9375_4478# 0.0163f
C58 a_3912_2366# check[6] 1.31e-20
C59 a_2060_2640# a_2777_2732# 4.45e-20
C60 a_1520_2366# D[6] 6.36e-20
C61 a_2061_2340# a_2479_2648# 0.00276f
C62 check[0] a_4926_4296# 0.00111f
C63 a_6010_3239# a_7073_4801# 6.75e-21
C64 a_7561_2366# check[0] 1.87e-20
C65 D[3] a_11629_2340# 1.1e-19
C66 check[4] a_10776_4086# 0.00416f
C67 a_12146_3239# a_12101_2550# 1.01e-20
C68 comparator_out a_4658_4086# 4.39e-21
C69 VDD a_9102_5083# 0.00984f
C70 a_12547_2366# x36.Q_N 0.0317f
C71 x4.X a_7562_4112# 6.4e-19
C72 a_6985_4112# a_7186_4112# 3.34e-19
C73 check[2] a_4855_4775# 2.07e-19
C74 a_8289_4086# a_8697_4112# 4.37e-19
C75 a_897_4112# a_1511_4112# 9.05e-20
C76 VDD a_897_4112# 0.414f
C77 a_6010_3239# a_8236_3239# 4e-20
C78 a_3599_2340# a_4154_2340# 0.197f
C79 a_4452_2640# x30.Q_N 0.00116f
C80 a_6759_3213# a_7158_3605# 0.00133f
C81 a_6291_3605# a_6605_3239# 0.0258f
C82 a_6010_3239# a_6977_3239# 0.00126f
C83 a_8237_4801# a_8858_4775# 0.117f
C84 x36.Q_N a_11331_4086# 1.3e-22
C85 comparator_out x63.Q_N 2.11e-19
C86 a_4854_3213# a_4657_2340# 2.52e-19
C87 a_4367_3213# a_4925_2550# 1.62e-19
C88 check[1] a_7481_5083# 4.45e-19
C89 a_1061_4801# a_897_4112# 0.00384f
C90 a_3504_2340# a_3505_4086# 1.07e-20
C91 x48.Q a_4318_5083# 4.61e-19
C92 a_4971_4801# a_4658_4086# 7.76e-20
C93 a_1996_2366# VDD 4.24e-19
C94 a_7317_2550# a_7186_4112# 1.72e-22
C95 a_4453_2340# a_6504_2648# 4.06e-20
C96 a_4680_3239# a_4213_3239# 0.00316f
C97 a_4367_3213# a_4585_3239# 3.73e-19
C98 VDD a_6978_4801# 0.00445f
C99 a_4073_3213# a_3913_4112# 0.00148f
C100 a_3452_3239# a_4453_4386# 6.5e-20
C101 a_3618_3239# a_4155_4086# 1.07e-20
C102 a_4854_3213# VDD 0.572f
C103 a_3453_4801# a_3807_4801# 0.0662f
C104 a_3619_4801# a_4681_4801# 0.137f
C105 a_3900_5167# a_4368_4775# 0.0633f
C106 a_5169_2366# VDD 4e-20
C107 x30.Q_N a_6846_4086# 0.0258f
C108 x5.X a_9152_4775# 0.00142f
C109 a_11089_4112# a_11630_4086# 0.125f
C110 a_11331_4086# a_11629_4386# 0.137f
C111 a_9377_4112# x39.Q_N 2.88e-20
C112 a_5991_2340# a_6780_2366# 4.2e-20
C113 a_2853_5648# a_3373_5674# 0.394f
C114 a_10345_3239# D[1] 0.0968f
C115 a_6304_2366# a_8288_2340# 8.55e-21
C116 check[1] a_3258_5648# 0.0414f
C117 a_4073_3213# x4.X 0.00798f
C118 a_9638_3213# a_10982_3239# 8.26e-21
C119 a_7073_4801# a_8403_4801# 4e-20
C120 check[1] sel_bit[1] 0.26f
C121 a_5845_4801# a_8591_4801# 3.65e-21
C122 comparator_out x5.X 6.13e-20
C123 a_9376_2366# x30.Q_N 2.98e-20
C124 x33.Q_N x39.Q_N 2.41e-20
C125 a_4367_3213# x45.Q_N 3.74e-20
C126 a_5844_3239# a_6760_4775# 9.66e-21
C127 a_11076_5167# a_11544_4775# 0.0633f
C128 a_10795_4801# a_11857_4801# 0.137f
C129 a_10629_4801# a_10983_4801# 0.0665f
C130 x77.Y D[6] 4.91e-19
C131 x75.Q_N x27.Q_N 0.02f
C132 x48.Q_N a_4113_4394# 2.02e-20
C133 a_4658_4086# a_4591_4478# 9.46e-19
C134 a_3913_4112# a_5372_4112# 1.65e-21
C135 a_4453_4386# a_4872_4394# 2.46e-19
C136 VDD a_3648_5972# 0.0123f
C137 a_8590_3239# x4.X 0.0062f
C138 VDD a_2969_6040# 0.00654f
C139 VDD a_4593_4112# 0.00494f
C140 x27.Q_N a_3913_4112# 1.32e-21
C141 a_7362_3239# x45.Q_N 0.00968f
C142 a_9465_4801# a_8697_4112# 3.76e-19
C143 a_9152_4775# a_9237_4386# 7.46e-19
C144 a_8591_4801# a_8384_4086# 3.44e-19
C145 a_8237_4801# x42.Q_N 3.67e-20
C146 a_8402_3239# a_8237_4801# 8.16e-19
C147 a_11075_3605# D[2] 3.24e-21
C148 a_11543_3213# a_12737_3239# 6.04e-19
C149 a_8236_3239# a_8403_4801# 9.04e-19
C150 a_3373_5674# a_3671_5674# 0.00489f
C151 comparator_out a_9237_4386# 2.49e-20
C152 a_11088_2366# check[4] 2.47e-20
C153 x36.Q_N a_11195_4112# 2.89e-22
C154 comparator_out a_4590_2732# 9.45e-19
C155 a_12030_3213# x36.Q_N 0.0126f
C156 x66.Q_N a_12031_4775# 4.45e-20
C157 x4.X a_5372_4112# 0.00623f
C158 a_5844_3239# a_6605_3239# 6.04e-20
C159 a_6305_4112# a_6845_4386# 0.139f
C160 a_5992_4086# a_6846_4086# 0.0492f
C161 x4.X x27.Q_N 0.425f
C162 a_9441_2340# x4.X 0.00148f
C163 a_2853_5648# eob 0.00163f
C164 x4.X x36.Q_N 0.278f
C165 a_1520_2366# a_2060_2640# 0.139f
C166 a_1207_2340# a_2061_2340# 0.0492f
C167 D[2] a_11088_2366# 5.92e-20
C168 a_5845_4801# a_6931_5083# 0.00907f
C169 a_6011_4801# a_6710_5083# 2.46e-19
C170 a_8696_2366# x63.Q_N 4.29e-21
C171 a_9237_2340# a_11629_2340# 0.00176f
C172 a_9639_4775# a_10983_4801# 8.26e-21
C173 a_11628_2640# x36.Q_N 0.572f
C174 a_5991_2340# check[6] 1.42e-21
C175 a_11630_4086# a_11767_4478# 0.00907f
C176 check[2] check[4] 0.347f
C177 D[6] a_3912_2366# 0.00221f
C178 x39.Q_N a_9954_4112# 2.57e-20
C179 a_11543_3213# a_11630_4086# 1.61e-19
C180 a_12030_3213# a_11629_4386# 3.78e-19
C181 a_10794_3239# x39.Q_N 0.348f
C182 VDD a_12102_4296# 0.317f
C183 a_11833_2340# a_12345_2732# 6.69e-20
C184 a_11629_2340# a_12547_2366# 0.0708f
C185 a_11088_2366# a_11969_2366# 0.00943f
C186 a_11330_2340# a_11768_2366# 0.00276f
C187 a_6759_3213# x30.Q_N 0.00506f
C188 a_9573_3239# x33.Q_N 1.68e-19
C189 a_4367_3213# a_6198_3239# 3.42e-20
C190 check[2] a_2883_5674# 0.0516f
C191 a_2389_5648# a_2969_6040# 0.00342f
C192 a_1338_5674# sel_bit[1] 0.0421f
C193 a_4854_3213# a_7072_3239# 1.86e-21
C194 x5.X a_4591_4478# 1.55e-19
C195 x4.X a_11629_4386# 0.0479f
C196 a_3452_3239# a_5561_3239# 1.03e-19
C197 VDD a_5170_4112# 1.14e-19
C198 a_1508_5167# a_1976_4775# 0.0627f
C199 a_9442_4086# x42.Q_N 0.00116f
C200 a_8402_3239# a_9442_4086# 2.9e-19
C201 a_8857_3213# a_9238_4086# 5.04e-19
C202 a_9638_3213# a_8697_4112# 9.49e-19
C203 a_1626_2366# VDD 0.00785f
C204 a_9151_3213# a_8939_4086# 2.12e-19
C205 a_3504_2340# x20.Q_N 6.66e-19
C206 a_6465_3213# a_6410_2366# 5.71e-21
C207 a_3912_2366# a_5991_2340# 1.15e-20
C208 a_4154_2340# a_4793_2366# 0.00316f
C209 a_5089_5083# a_5845_4801# 4.06e-20
C210 a_4452_2640# a_4592_2366# 0.00126f
C211 a_11628_2640# a_11629_4386# 1.32e-20
C212 a_11088_2366# a_11834_4086# 7.14e-22
C213 a_11330_2340# a_11630_4086# 3.47e-21
C214 a_7072_3239# a_7181_3239# 0.00707f
C215 x5.X a_11390_4801# 9.46e-19
C216 a_6546_2340# x30.Q_N 0.16f
C217 a_8403_4801# a_9370_4801# 0.00126f
C218 a_8237_4801# a_9873_5083# 1.25e-19
C219 a_9152_4775# a_9551_5167# 0.00133f
C220 a_8684_5167# a_8998_4801# 0.0258f
C221 a_4680_3239# a_3453_4801# 4.76e-21
C222 a_4367_3213# a_4074_4775# 7.57e-21
C223 reset x3.A 0.00364f
C224 a_4367_3213# x20.Q_N 1.25e-21
C225 a_1720_2648# x4.X 0.00102f
C226 x48.Q a_2993_5674# 1.96e-19
C227 a_6305_4112# a_7264_4394# 1.21e-20
C228 a_6845_4386# a_6983_4478# 1.09e-19
C229 a_6547_4086# a_6411_4112# 0.0282f
C230 a_11969_2366# check[2] 4.38e-19
C231 a_6465_3213# a_6547_4086# 1.02e-19
C232 a_6759_3213# a_5992_4086# 8.83e-19
C233 a_6291_3605# a_6305_4112# 1.61e-19
C234 a_6010_3239# a_6845_4386# 4.11e-20
C235 a_4453_2340# a_4926_4296# 6.08e-21
C236 x5.X a_7954_4801# 0.0293f
C237 a_8696_2366# a_9237_4386# 1.93e-22
C238 a_5991_2340# a_6410_2366# 0.0397f
C239 a_6304_2366# a_6982_2732# 0.00652f
C240 a_5896_2340# VDD 0.189f
C241 VDD a_1415_4801# 0.12f
C242 a_6546_2340# a_6780_2732# 0.00976f
C243 a_6466_4775# check[5] 1.71e-20
C244 a_4970_3239# x27.Q_N 0.00341f
C245 a_7362_3239# a_7049_2340# 3.49e-20
C246 check[0] a_5562_4801# 0.0162f
C247 a_10345_3239# a_10346_4801# 9.85e-20
C248 check[1] a_4926_4296# 1.97e-22
C249 check[4] a_11250_4775# 6.31e-19
C250 sel_bit[1] a_3453_4801# 0.00123f
C251 a_1061_4801# a_1415_4801# 0.0708f
C252 x4.X a_1976_4775# 0.0979f
C253 a_1227_4801# a_2289_4801# 0.137f
C254 a_3505_4086# a_4454_4086# 1.03e-19
C255 a_3600_4086# a_4453_4386# 0.0264f
C256 a_3913_4112# a_4155_4086# 0.124f
C257 a_2883_5674# x20.Q_N 5.75e-20
C258 check[2] a_11834_4086# 1.08e-19
C259 a_5991_2340# a_6547_4086# 1.3e-22
C260 a_6304_2366# a_6305_4112# 1.8e-19
C261 VDD a_1062_5674# 0.23f
C262 VDD a_4658_4086# 0.489f
C263 a_7763_2366# a_7561_2366# 3.67e-19
C264 a_3807_4801# a_4008_4801# 3.67e-19
C265 a_4681_4801# a_4586_4801# 0.00276f
C266 a_4855_4775# a_5089_5083# 0.00945f
C267 a_4368_4775# x27.Q_N 0.00773f
C268 a_8288_2340# a_8383_2340# 0.0968f
C269 a_6780_2366# a_7185_2366# 2.46e-21
C270 x57.Q_N x27.Q_N 7.46e-20
C271 a_9754_3239# VDD 4.88e-19
C272 a_11543_3213# a_10982_3239# 3.79e-20
C273 a_11075_3605# a_11159_3605# 0.00972f
C274 a_12030_3213# a_11856_3239# 0.197f
C275 D[3] check[4] 0.00432f
C276 a_10628_3239# a_11493_3521# 0.00276f
C277 D[1] x36.Q_N 1.36e-20
C278 x4.X a_4155_4086# 0.00873f
C279 a_1062_5674# a_1061_4801# 0.00165f
C280 comparator_out x30.Q_N 0.274f
C281 a_11544_4775# x36.Q_N 0.0059f
C282 a_12031_4775# a_12265_5083# 0.00945f
C283 a_10983_4801# a_11184_4801# 3.67e-19
C284 a_11857_4801# a_11762_4801# 0.00276f
C285 x4.X a_12048_4394# 8.47e-19
C286 a_4454_4086# x45.Q_N 3.85e-19
C287 a_11856_3239# x4.X 0.00481f
C288 a_8939_4086# a_10776_4086# 1.86e-21
C289 a_9238_4086# a_9377_4112# 2.56e-19
C290 a_9237_4386# a_9578_4112# 0.00118f
C291 x42.Q_N a_10156_4112# 8.23e-20
C292 check[6] a_6199_4801# 0.165f
C293 x63.Q_N VDD 0.0716f
C294 a_12030_3213# a_11629_2340# 8.72e-19
C295 a_11856_3239# a_11628_2640# 1.11e-20
C296 x33.Q_N a_9238_4086# 0.026f
C297 a_11543_3213# a_11833_2340# 0.00144f
C298 x66.Q_N D[2] 2.25e-19
C299 comparator_out a_6780_2732# 1.8e-19
C300 eob a_1616_4801# 4.1e-19
C301 check[1] x27.D 1.12e-20
C302 a_11629_2340# x4.X 0.00254f
C303 check[0] a_3876_6040# 2.26e-19
C304 a_3170_4801# a_1511_4112# 5.42e-19
C305 a_6465_3213# a_6411_4112# 3.34e-20
C306 a_5371_2366# check[6] 0.00326f
C307 a_6010_3239# a_6291_3605# 0.155f
C308 check[0] a_6305_4112# 0.00126f
C309 VDD a_3170_4801# 0.212f
C310 a_2060_2640# a_3912_2366# 1.9e-19
C311 D[3] a_11969_2366# 7.69e-20
C312 a_2265_2340# a_2401_2366# 0.07f
C313 a_2061_2340# a_3599_2340# 0.00116f
C314 comparator_out a_5992_4086# 0.00201f
C315 a_11628_2640# a_11629_2340# 0.781f
C316 a_11088_2366# a_12101_2550# 0.0633f
C317 a_5844_3239# a_6305_4112# 2.21e-19
C318 a_10775_2340# x63.Q_N 0.124f
C319 a_11330_2340# a_11833_2340# 0.00187f
C320 a_10983_4801# a_10776_4086# 3.44e-19
C321 a_8288_2340# x33.Q_N 3.7e-19
C322 a_11544_4775# a_11629_4386# 7.46e-19
C323 a_10629_4801# x39.Q_N 3.68e-20
C324 a_11857_4801# a_11089_4112# 3.76e-19
C325 x33.Q_N a_9755_4801# 3.78e-19
C326 check[1] a_6760_4775# 0.00254f
C327 a_1061_4801# a_3170_4801# 1.03e-19
C328 check[2] a_4454_4086# 2.36e-20
C329 x5.X a_1511_4112# 2.24e-19
C330 x5.A a_1338_5674# 0.263f
C331 a_1062_5674# a_2389_5648# 1.61e-20
C332 x5.X a_11289_4394# 4.41e-19
C333 D[4] x5.X 3.43e-19
C334 a_3618_3239# a_4367_3213# 0.139f
C335 a_4073_3213# a_3899_3605# 0.205f
C336 a_3452_3239# a_4854_3213# 0.0492f
C337 VDD x5.X 2.74f
C338 a_2198_2732# x20.Q_N 0.00203f
C339 a_4657_2340# a_4590_2732# 9.46e-19
C340 a_3912_2366# a_5371_2366# 9.06e-21
C341 a_6010_3239# a_6304_2366# 5.94e-19
C342 a_4452_2640# a_4871_2648# 2.46e-19
C343 a_4539_5083# check[6] 1.43e-21
C344 a_6465_3213# a_5991_2340# 2.5e-19
C345 x54.Q_N a_4112_2648# 2.02e-20
C346 a_12146_3239# x39.Q_N 0.00968f
C347 VDD a_6292_5167# 0.317f
C348 a_11761_3239# x39.Q_N 0.00399f
C349 check[1] a_9238_4086# 2.12e-19
C350 a_11565_4112# a_11089_4112# 2.87e-21
C351 x5.X a_1061_4801# 0.265f
C352 a_11715_5083# check[3] 9.55e-19
C353 x4.X a_5845_4801# 0.00422f
C354 x5.X a_7318_4296# 6.4e-19
C355 comparator_out eob 3.93e-19
C356 a_2463_4775# a_3900_5167# 7.98e-21
C357 a_7247_4775# a_6846_4086# 0.00169f
C358 a_6466_4775# x45.Q_N 2.19e-19
C359 a_12101_2550# check[2] 2.02e-19
C360 a_6760_4775# a_7050_4086# 0.00268f
C361 a_7073_4801# a_6845_4386# 1.96e-20
C362 x4.X a_12147_4801# 0.00557f
C363 a_4590_2732# VDD 0.0172f
C364 VDD a_9237_4386# 0.59f
C365 a_2289_4801# x20.Q_N 8.79e-19
C366 a_8997_3239# x42.Q_N 0.0309f
C367 a_5896_2340# a_6845_2340# 1.03e-19
C368 a_8590_3239# a_8767_3605# 8.94e-19
C369 a_7158_3605# VDD 0.00371f
C370 a_9151_3213# a_9101_3521# 1.21e-20
C371 a_8402_3239# a_8997_3239# 0.00118f
C372 x27.Q_N a_6606_4801# 1.93e-20
C373 a_8696_2366# x30.Q_N 8.85e-20
C374 comparator_out x4.A 1.12e-19
C375 a_8288_2340# check[1] 0.027f
C376 a_8998_4801# x33.Q_N 4.01e-20
C377 x75.Q_N a_4855_4775# 4.45e-20
C378 a_3899_3605# x27.Q_N 0.00192f
C379 x4.X a_8384_4086# 0.101f
C380 a_4789_3239# x4.X 1.05e-19
C381 a_2389_5648# a_3170_4801# 1.39e-19
C382 a_4368_4775# a_4155_4086# 3.72e-19
C383 a_4855_4775# a_3913_4112# 0.00161f
C384 a_6547_4086# x42.Q_N 7.23e-21
C385 a_4074_4775# a_4454_4086# 0.00336f
C386 a_3619_4801# a_4658_4086# 0.00221f
C387 x20.Q_N a_4454_4086# 1.21e-19
C388 a_6930_3521# x45.Q_N 0.00203f
C389 check[0] a_6983_4478# 6.27e-20
C390 VDD a_3984_5167# 0.0046f
C391 a_6844_2640# a_7561_2366# 0.00105f
C392 D[1] a_11856_3239# 3.54e-20
C393 x48.Q check[0] 0.0102f
C394 a_6010_3239# check[0] 0.0252f
C395 a_7481_5083# check[5] 1.93e-21
C396 a_9237_2340# check[4] 0.0399f
C397 x30.Q_N a_7954_4801# 0.182f
C398 a_12030_3213# a_12031_4775# 0.00237f
C399 comparator_out a_2777_2732# 8.11e-19
C400 VDD a_11160_5167# 0.0042f
C401 x75.Q x45.Q_N 9.42e-21
C402 a_5844_3239# a_6010_3239# 0.782f
C403 a_2265_2340# eob 9.03e-20
C404 x77.Y a_4452_2640# 4.61e-20
C405 a_1227_4801# a_3807_4801# 3.07e-21
C406 x4.X a_4855_4775# 0.102f
C407 a_2389_5648# x5.X 0.00112f
C408 sel_bit[0] a_2853_5648# 1.09f
C409 sel_bit[1] x3.A 1.43e-20
C410 check[2] a_6466_4775# 1.08e-19
C411 x4.X a_12031_4775# 0.0991f
C412 D[1] a_11629_2340# 1.09e-20
C413 a_9441_2340# a_9709_2550# 0.205f
C414 a_9237_2340# x60.Q_N 1.07e-19
C415 clk_sar reset 1.31e-20
C416 a_12737_3239# x36.Q_N 0.0107f
C417 a_11970_4112# VDD 0.0326f
C418 check[2] a_8939_4086# 5.79e-20
C419 x5.X a_8289_4086# 0.0767f
C420 a_3170_4801# a_3619_4801# 6.24e-19
C421 x27.D a_3453_4801# 0.412f
C422 a_2060_2640# D[6] 0.00655f
C423 a_2061_2340# a_2979_2366# 0.0708f
C424 a_2265_2340# a_2777_2732# 6.69e-20
C425 VDD a_9656_4394# 0.00984f
C426 a_4452_2640# check[6] 0.0327f
C427 a_9151_3213# x39.Q_N 3.3e-20
C428 D[2] a_12547_2366# 6.35e-19
C429 a_6759_3213# a_7247_4775# 1.08e-22
C430 a_7246_3213# a_6760_4775# 1.06e-20
C431 D[3] a_12101_2550# 1.91e-20
C432 VDD a_9551_5167# 0.00371f
C433 comparator_out a_8896_2648# 1.53e-19
C434 a_11768_2366# x36.Q_N 0.00473f
C435 check[1] a_5562_4801# 3.76e-20
C436 x4.X a_9173_4478# 2.12e-19
C437 x5.X a_3619_4801# 0.0076f
C438 a_8289_4086# a_9237_4386# 9.65e-21
C439 a_7764_4112# a_9238_4086# 3.65e-21
C440 x4.X a_7182_4801# 2.39e-19
C441 a_6845_2340# x5.X 2.59e-20
C442 x5.X a_2697_5083# 3.53e-19
C443 a_4368_4775# a_5845_4801# 1.72e-19
C444 a_3912_2366# a_4452_2640# 0.139f
C445 a_3599_2340# a_4453_2340# 0.0492f
C446 x5.X a_10795_4801# 0.0203f
C447 a_4970_3239# a_4789_3239# 4.11e-20
C448 a_7072_3239# a_7158_3605# 0.00976f
C449 a_6010_3239# x72.Q_N 5.46e-21
C450 a_8403_4801# a_8684_5167# 0.155f
C451 a_8237_4801# a_9152_4775# 0.125f
C452 a_10628_3239# check[3] 1.99e-20
C453 x36.Q_N a_11630_4086# 0.0255f
C454 a_11544_4775# a_12147_4801# 0.0552f
C455 a_4213_3239# a_3599_2340# 4.6e-20
C456 a_4680_3239# a_4925_2550# 1.85e-20
C457 x48.Q a_4389_4478# 3.17e-19
C458 check[6] a_6846_4086# 2.07e-22
C459 a_5371_2366# a_5991_2340# 8.26e-21
C460 a_4452_2640# a_6410_2366# 2.44e-20
C461 x48.Q a_4767_5167# 1.31e-19
C462 a_4367_3213# x75.Q_N 0.00553f
C463 a_2401_2366# VDD 0.00631f
C464 a_3806_3239# a_4007_3239# 3.67e-19
C465 a_4680_3239# a_4585_3239# 0.00276f
C466 a_4854_3213# a_5088_3521# 0.00945f
C467 D[0] a_7181_3239# 9.28e-21
C468 D[4] x30.Q_N 0.005f
C469 VDD x30.Q_N 0.444f
C470 a_3452_3239# a_4658_4086# 0.00195f
C471 a_4073_3213# a_4453_4386# 0.0015f
C472 a_3618_3239# a_4454_4086# 6.04e-20
C473 a_3899_3605# a_4155_4086# 1.7e-20
C474 a_4367_3213# a_3913_4112# 3.33e-20
C475 a_11769_4112# check[2] 3.17e-20
C476 a_3806_3239# VDD 0.117f
C477 a_3504_2340# x4.X 0.0105f
C478 check[2] a_8803_4112# 1.27e-20
C479 x4.X a_6400_4801# 8.46e-20
C480 a_4925_2550# a_4794_4112# 1.72e-22
C481 a_4074_4775# a_3807_4801# 6.99e-20
C482 a_3619_4801# a_3984_5167# 4.45e-20
C483 a_4368_4775# a_4855_4775# 0.273f
C484 a_6780_2732# VDD 0.00371f
C485 a_10776_4086# x39.Q_N 0.155f
C486 a_11629_4386# a_11630_4086# 0.782f
C487 a_6304_2366# a_6984_2366# 3.73e-19
C488 x30.Q_N a_7318_4296# 5.71e-19
C489 a_6844_2640# a_8288_2340# 6.58e-19
C490 a_11089_4112# a_12102_4296# 0.0633f
C491 x5.X a_9465_4801# 0.00117f
C492 a_6546_2340# a_6780_2366# 0.00707f
C493 x20.Q_N a_3807_4801# 1.92e-19
C494 check[2] a_9323_5083# 4.69e-19
C495 a_11331_4086# a_11834_4086# 0.00187f
C496 a_9151_3213# a_9573_3239# 2.87e-21
C497 a_9322_3521# VDD 0.0163f
C498 a_4367_3213# x4.X 0.112f
C499 a_9638_3213# a_9754_3239# 0.0397f
C500 a_8997_3239# a_9369_3239# 3.34e-19
C501 check[1] a_6305_4112# 0.00312f
C502 a_4680_3239# x45.Q_N 1.74e-21
C503 comparator_out a_1520_2366# 0.00311f
C504 a_10795_4801# a_11160_5167# 4.45e-20
C505 a_11250_4775# a_10983_4801# 6.99e-20
C506 a_11544_4775# a_12031_4775# 0.273f
C507 sel_bit[1] a_3505_4086# 1.09e-19
C508 VDD a_3373_5674# 0.353f
C509 a_3913_4112# a_4389_4112# 2.87e-21
C510 a_4454_4086# a_5170_4478# 0.0018f
C511 a_4453_4386# a_5372_4112# 0.162f
C512 a_4658_4086# a_4872_4394# 0.0104f
C513 a_7362_3239# x4.X 5.65e-19
C514 a_8384_4086# a_8897_4394# 0.00945f
C515 VDD a_5992_4086# 0.716f
C516 x4.X check[4] 0.037f
C517 x27.Q_N a_4453_4386# 0.0318f
C518 a_8383_2340# a_9172_2732# 7.71e-20
C519 a_8696_2366# a_8896_2648# 0.00185f
C520 a_10628_3239# a_10680_2340# 4.5e-19
C521 a_9152_4775# a_9442_4086# 0.00268f
C522 a_8858_4775# x42.Q_N 2.19e-19
C523 a_12030_3213# D[2] 0.00376f
C524 a_9465_4801# a_9237_4386# 1.96e-20
C525 a_9639_4775# a_9238_4086# 0.00169f
C526 a_9754_3239# a_9236_2640# 5.05e-21
C527 a_8236_3239# a_8684_5167# 8.3e-21
C528 a_8857_3213# a_8403_4801# 3.18e-21
C529 comparator_out a_4871_2648# 6.94e-19
C530 comparator_out a_9442_4086# 4.39e-21
C531 sel_bit[1] a_1227_4801# 3.62e-20
C532 a_5844_3239# a_8236_3239# 0.00176f
C533 x4.X a_4389_4112# 3.84e-19
C534 a_5844_3239# a_6977_3239# 2.56e-19
C535 D[2] x4.X 4e-19
C536 a_5992_4086# a_7318_4296# 4.7e-22
C537 a_6547_4086# a_6846_4086# 0.0334f
C538 a_6305_4112# a_7050_4086# 0.199f
C539 a_4794_4112# x45.Q_N 5.94e-20
C540 x60.Q_N x4.X 0.00784f
C541 x5.X a_6710_5083# 3.44e-19
C542 a_7561_2366# check[5] 5.2e-20
C543 a_1520_2366# a_2265_2340# 0.199f
C544 a_1762_2340# a_2061_2340# 0.0334f
C545 a_6759_3213# check[6] 8.24e-21
C546 a_1207_2340# a_2533_2550# 4.7e-22
C547 a_12737_3239# a_11629_2340# 4.83e-19
C548 D[2] a_11628_2640# 0.00729f
C549 a_12030_3213# a_11969_2366# 1.2e-20
C550 a_9236_2640# x63.Q_N 1.48e-19
C551 a_5845_4801# a_6606_4801# 6.04e-20
C552 a_6011_4801# a_7159_5167# 2.13e-19
C553 a_6466_4775# a_6931_5083# 9.46e-19
C554 check[0] a_4318_5083# 1.54e-19
C555 a_6984_2366# check[0] 3.17e-19
C556 eob a_1511_4112# 0.0585f
C557 a_3452_3239# x5.X 3.24e-20
C558 a_11833_2340# x36.Q_N 0.179f
C559 a_9152_4775# a_9574_4801# 2.87e-21
C560 a_9639_4775# a_9755_4801# 0.0397f
C561 VDD eob 2.32f
C562 x4.A a_1511_4112# 0.619f
C563 a_3453_4801# a_5562_4801# 1.03e-19
C564 VDD x4.A 0.787f
C565 D[6] a_4452_2640# 1.85e-19
C566 a_2979_2366# a_4453_2340# 3.65e-21
C567 a_11630_4086# a_12048_4394# 0.00276f
C568 a_11629_4386# a_12346_4478# 4.45e-20
C569 a_12030_3213# a_11834_4086# 2.47e-19
C570 eob a_1061_4801# 0.514f
C571 a_11075_3605# x39.Q_N 0.152f
C572 a_11543_3213# a_12102_4296# 1.71e-19
C573 a_11629_2340# a_11768_2366# 2.56e-19
C574 a_12101_2550# a_12547_2366# 0.0367f
C575 a_11628_2640# a_11969_2366# 0.00118f
C576 a_7954_4801# a_8237_4801# 8.18e-19
C577 a_7072_3239# x30.Q_N 0.00298f
C578 check[1] a_6983_4478# 9.03e-21
C579 check[2] a_3258_5648# 0.0201f
C580 check[1] x48.Q 0.0512f
C581 a_2389_5648# a_3373_5674# 0.176f
C582 a_10629_4801# a_12738_4801# 9.94e-20
C583 a_4367_3213# a_4970_3239# 0.0552f
C584 a_1061_4801# x4.A 0.00353f
C585 check[2] sel_bit[1] 0.393f
C586 x5.X a_4872_4394# 1.11e-19
C587 clk_sar sel_bit[1] 0.329f
C588 x4.X a_11834_4086# 0.00986f
C589 a_5845_4801# a_5897_4086# 6.04e-19
C590 x77.Y comparator_out 0.00119f
C591 VDD a_6781_4478# 0.00371f
C592 a_1976_4775# a_2463_4775# 0.271f
C593 a_9638_3213# a_9237_4386# 3.78e-19
C594 a_2777_2732# VDD 0.00561f
C595 a_9151_3213# a_9238_4086# 1.61e-19
C596 a_8402_3239# x42.Q_N 0.345f
C597 a_2200_2366# x20.Q_N 0.00397f
C598 a_8236_3239# a_8857_3213# 0.117f
C599 a_4452_2640# a_5991_2340# 3.67e-19
C600 a_4657_2340# a_4592_2366# 9.75e-19
C601 a_4453_2340# a_4793_2366# 6.04e-20
C602 a_11629_2340# a_11630_4086# 1.55e-19
C603 x27.Q_N a_6011_4801# 1.48e-19
C604 a_11833_2340# a_11629_4386# 1.26e-21
C605 D[7] a_897_4112# 3.76e-20
C606 a_11088_2366# x39.Q_N 6.35e-20
C607 x72.Q_N a_8236_3239# 2.94e-19
C608 a_6845_2340# x30.Q_N 0.0463f
C609 x5.X a_11762_4801# 2.61e-19
C610 comparator_out a_10156_4112# 5.5e-20
C611 a_8403_4801# x33.Q_N 2.97e-20
C612 a_9465_4801# a_9551_5167# 0.00976f
C613 a_7363_4801# a_7182_4801# 4.11e-20
C614 a_4367_3213# a_4368_4775# 0.00121f
C615 a_2198_2732# x4.X 9.81e-19
C616 x48.Q a_3877_5674# 4.02e-19
C617 x36.Q_N a_11966_4801# 7.29e-21
C618 a_7050_4086# a_6983_4478# 9.46e-19
C619 a_6845_4386# a_7264_4394# 2.46e-19
C620 x45.Q_N a_6505_4394# 2.02e-20
C621 a_6305_4112# a_7764_4112# 1.65e-21
C622 a_6759_3213# a_6547_4086# 2.12e-19
C623 a_7246_3213# a_6305_4112# 9.49e-19
C624 a_6465_3213# a_6846_4086# 5.04e-19
C625 a_6010_3239# a_7050_4086# 2.9e-19
C626 a_6304_2366# a_7263_2648# 1.21e-20
C627 a_6844_2640# a_6982_2732# 1.09e-19
C628 D[5] a_6984_2366# 8.02e-20
C629 a_8696_2366# a_9442_4086# 7.14e-22
C630 a_8938_2340# a_9238_4086# 3.47e-21
C631 a_6546_2340# a_6410_2366# 0.0282f
C632 a_9236_2640# a_9237_4386# 1.32e-20
C633 VDD a_1926_5083# 0.0117f
C634 a_4592_2366# VDD 0.00111f
C635 a_8236_3239# a_8383_2340# 8.35e-19
C636 D[7] a_1996_2366# 1.53e-19
C637 D[0] a_9754_3239# 1.61e-20
C638 a_6760_4775# check[5] 0.00406f
C639 a_7247_4775# a_7954_4801# 0.0968f
C640 D[1] check[4] 0.435f
C641 a_2389_5648# eob 0.222f
C642 a_9151_3213# a_9755_4801# 1.05e-20
C643 comparator_out check[6] 0.0236f
C644 check[4] a_11544_4775# 0.00302f
C645 a_5561_3239# x27.Q_N 0.00748f
C646 comparator_out check[3] 0.0244f
C647 a_1061_4801# a_1926_5083# 0.00276f
C648 a_1682_4775# a_1415_4801# 6.99e-20
C649 a_1227_4801# a_1592_5167# 4.45e-20
C650 x4.X a_2289_4801# 0.167f
C651 a_3913_4112# a_4454_4086# 0.125f
C652 a_4155_4086# a_4453_4386# 0.137f
C653 sel_bit[1] x20.Q_N 3.57e-20
C654 x5.X a_11089_4112# 0.00571f
C655 a_6304_2366# a_6845_4386# 1.93e-22
C656 check[2] x39.Q_N 0.0223f
C657 VDD x48.Q_N 0.0812f
C658 a_8896_2648# VDD 0.00506f
C659 check[5] a_9238_4086# 6.24e-22
C660 a_4681_4801# x27.Q_N 5.04e-19
C661 a_12030_3213# a_12548_4112# 2.07e-19
C662 a_10794_3239# a_11714_3521# 1.09e-19
C663 a_11493_3521# VDD 0.00984f
C664 a_11249_3213# a_11493_3521# 0.0104f
C665 a_12737_3239# a_12031_4775# 4.94e-20
C666 a_6606_4801# a_7182_4801# 2.46e-21
C667 comparator_out a_3912_2366# 0.00684f
C668 x5.A a_1227_4801# 6.32e-21
C669 x4.X a_4454_4086# 0.0468f
C670 check[1] a_8403_4801# 0.00119f
C671 a_11857_4801# x36.Q_N 8.57e-20
C672 x4.X a_12548_4112# 0.00434f
C673 a_11159_3605# x4.X 9.07e-19
C674 a_4926_4296# x45.Q_N 1.43e-19
C675 a_9442_4086# a_9578_4112# 0.07f
C676 x42.Q_N a_9173_4112# 0.00139f
C677 a_9238_4086# a_10776_4086# 2.98e-19
C678 a_9237_4386# a_11089_4112# 9.95e-20
C679 a_8802_2366# a_9172_2366# 4.11e-20
C680 check[6] a_4971_4801# 8.4e-20
C681 a_11856_3239# a_11833_2340# 1.03e-19
C682 a_12030_3213# a_12101_2550# 1.66e-21
C683 VDD a_8237_4801# 0.81f
C684 x33.Q_N a_9710_4296# 5.71e-19
C685 a_8236_3239# x33.Q_N 2.78e-19
C686 a_9151_3213# a_8998_4801# 1.61e-20
C687 eob a_3619_4801# 9.05e-22
C688 check[5] a_9755_4801# 1.85e-20
C689 eob a_2697_5083# 4.29e-19
C690 x77.Y a_4214_4801# 1.91e-20
C691 a_12101_2550# x4.X 0.00146f
C692 x27.D a_3505_4086# 5.09e-21
C693 D[0] x5.X 0.00133f
C694 a_2061_2340# a_4154_2340# 6.38e-20
C695 check[0] a_6845_4386# 1.56e-19
C696 a_6465_3213# a_6759_3213# 0.199f
C697 a_6010_3239# a_7246_3213# 0.0264f
C698 a_2265_2340# a_3912_2366# 9.6e-21
C699 a_2533_2550# a_3599_2340# 7.98e-21
C700 a_11629_2340# a_11833_2340# 0.117f
C701 a_11628_2640# a_12101_2550# 0.145f
C702 a_11330_2340# x63.Q_N 9.58e-21
C703 a_5844_3239# a_6845_4386# 6.5e-20
C704 a_11250_4775# x39.Q_N 2.02e-19
C705 a_11857_4801# a_11629_4386# 1.96e-20
C706 a_12031_4775# a_11630_4086# 0.00169f
C707 a_11544_4775# a_11834_4086# 0.00268f
C708 comparator_out a_10680_2340# 7.8e-19
C709 check[1] a_7073_4801# 0.00111f
C710 a_1227_4801# x27.D 4.24e-20
C711 check[2] a_4926_4296# 2.18e-22
C712 x5.X a_3600_4086# 1.13e-19
C713 x5.A check[2] 0.00137f
C714 a_1520_2366# a_1511_4112# 7.01e-19
C715 clk_sar x5.A 0.00356f
C716 x5.X a_11767_4478# 4e-19
C717 x48.Q a_3453_4801# 0.0505f
C718 a_3452_3239# a_3806_3239# 0.0662f
C719 a_3899_3605# a_4367_3213# 0.0632f
C720 a_3618_3239# a_4680_3239# 0.137f
C721 a_4452_2640# a_5371_2366# 0.159f
C722 a_4453_2340# a_5169_2732# 0.0018f
C723 a_2479_2648# x20.Q_N 0.00136f
C724 a_4657_2340# a_4871_2648# 0.0104f
C725 a_6291_3605# a_6304_2366# 1.71e-19
C726 a_6010_3239# a_6844_2640# 4.04e-20
C727 a_6465_3213# a_6546_2340# 4.18e-20
C728 a_1520_2366# VDD 0.402f
C729 a_6759_3213# a_5991_2340# 9.06e-19
C730 VDD a_7247_4775# 0.72f
C731 x66.Q_N x39.Q_N 3.91e-19
C732 check[5] a_8998_4801# 2.15e-19
C733 check[1] a_9710_4296# 3.53e-20
C734 a_8236_3239# check[1] 0.0444f
C735 a_11970_4112# a_11089_4112# 0.00943f
C736 a_11769_4112# a_11331_4086# 0.00276f
C737 x5.X a_1682_4775# 0.00283f
C738 a_11390_4801# check[3] 1.02e-20
C739 x4.X a_6466_4775# 9.39e-19
C740 a_7247_4775# a_7318_4296# 2.97e-21
C741 a_6760_4775# x45.Q_N 9.66e-21
C742 a_7073_4801# a_7050_4086# 2.59e-19
C743 a_9710_4296# a_9954_4112# 0.00812f
C744 x75.Q_N x75.Q 2.81e-20
C745 a_4871_2648# VDD 0.0102f
C746 D[7] a_1626_2366# 0.00202f
C747 VDD a_9442_4086# 0.487f
C748 a_10628_3239# x42.Q_N 1.47e-19
C749 a_5991_2340# a_6546_2340# 0.197f
C750 a_8236_3239# a_10794_3239# 2.9e-21
C751 a_8402_3239# a_10628_3239# 4e-20
C752 a_9369_3239# x42.Q_N 0.00401f
C753 a_8683_3605# a_8997_3239# 0.0258f
C754 a_9151_3213# a_9550_3605# 0.00133f
C755 a_8402_3239# a_9369_3239# 0.00126f
C756 a_8236_3239# a_9872_3521# 1.25e-19
C757 x27.Q_N a_6978_4801# 1.15e-20
C758 a_9236_2640# x30.Q_N 1.21e-20
C759 a_4854_3213# a_5372_4112# 2.07e-19
C760 a_11194_2366# check[3] 1.29e-19
C761 a_10346_4801# check[4] 0.13f
C762 a_9370_4801# x33.Q_N 4.03e-20
C763 a_4854_3213# x27.Q_N 0.0125f
C764 a_4388_2732# x4.X 4.32e-19
C765 x4.X a_8939_4086# 0.00731f
C766 a_6930_3521# x4.X 9.99e-19
C767 a_4855_4775# a_4453_4386# 6.17e-19
C768 a_4368_4775# a_4454_4086# 4.63e-19
C769 check[2] x27.D 1.63e-20
C770 a_6846_4086# x42.Q_N 2.42e-19
C771 a_6845_2340# a_8896_2648# 4.06e-20
C772 a_6605_3239# x45.Q_N 0.031f
C773 a_8237_4801# a_8289_4086# 6.04e-19
C774 a_5169_2366# x27.Q_N 0.00224f
C775 check[0] a_7264_4394# 1.47e-20
C776 VDD a_2398_4801# 6.04e-19
C777 x75.Q x4.X 8.71e-19
C778 a_6291_3605# check[0] 7.4e-20
C779 a_9709_2550# check[4] 0.00101f
C780 comparator_out D[6] 0.00566f
C781 VDD a_9574_4801# 7.87e-19
C782 comparator_out a_6465_3213# 4.84e-19
C783 a_5844_3239# a_6291_3605# 0.15f
C784 a_2784_5996# a_2883_5674# 0.00134f
C785 x77.Y a_4657_2340# 1.11e-19
C786 x4.X a_3807_4801# 2.51e-19
C787 check[2] a_6760_4775# 1.3e-19
C788 a_3452_3239# eob 3.51e-19
C789 x4.X a_10983_4801# 2.36e-19
C790 a_8696_2366# a_10680_2340# 7.33e-21
C791 a_12737_3239# D[2] 0.0747f
C792 a_5845_4801# a_6011_4801# 0.751f
C793 sel_bit[0] a_1511_4112# 3.42e-19
C794 a_8383_2340# a_9172_2366# 4.2e-20
C795 a_6304_2366# check[0] 0.00297f
C796 VDD sel_bit[0] 1.26f
C797 a_8237_4801# a_10795_4801# 2.9e-21
C798 a_8403_4801# a_10629_4801# 4e-20
C799 a_5844_3239# a_6304_2366# 1.89e-19
C800 comparator_out a_5991_2340# 0.00445f
C801 x77.Y VDD 0.423f
C802 a_12147_4801# a_11966_4801# 4.11e-20
C803 check[2] a_9238_4086# 0.439f
C804 sel_bit[0] a_1061_4801# 5.2e-20
C805 check[5] a_6305_4112# 7.68e-22
C806 x27.D a_4074_4775# 6.07e-19
C807 a_2265_2340# D[6] 1.59e-19
C808 VDD a_10156_4112# 0.109f
C809 a_2533_2550# a_2979_2366# 0.0367f
C810 x20.Q_N x27.D 0.0032f
C811 a_4657_2340# check[6] 6.83e-20
C812 x48.Q a_4790_4801# 6.64e-20
C813 a_7072_3239# a_7247_4775# 1.33e-23
C814 a_7246_3213# a_7073_4801# 4.82e-21
C815 a_11769_4112# x4.X 6.71e-19
C816 check[4] a_11630_4086# 1.46e-21
C817 comparator_out a_9374_2732# 9.52e-19
C818 a_12345_2366# x36.Q_N 0.00224f
C819 a_8791_3239# x33.Q_N 6.75e-20
C820 x4.X a_8803_4112# 0.00332f
C821 check[2] a_2579_4801# 1.13e-21
C822 a_8384_4086# a_8697_4112# 0.272f
C823 x5.X a_3900_5167# 1.6e-19
C824 a_10345_3239# x5.X 0.00125f
C825 a_4681_4801# a_5845_4801# 6.38e-20
C826 a_6759_3213# x42.Q_N 3.3e-20
C827 a_4855_4775# a_6011_4801# 1.83e-19
C828 a_4154_2340# a_4453_2340# 0.0334f
C829 a_11768_2366# a_11969_2366# 3.34e-19
C830 a_3912_2366# a_4657_2340# 0.199f
C831 a_7246_3213# a_8236_3239# 0.00116f
C832 a_3599_2340# a_4925_2550# 4.7e-22
C833 D[2] a_11630_4086# 3.53e-19
C834 a_1207_2340# x20.Q_N 0.144f
C835 a_6759_3213# a_8402_3239# 1.98e-19
C836 VDD check[6] 0.503f
C837 x5.X a_11076_5167# 0.00471f
C838 a_6759_3213# a_7480_3521# 0.00185f
C839 D[0] x30.Q_N 3.29e-19
C840 a_9172_2366# x33.Q_N 9.42e-19
C841 a_8237_4801# a_9465_4801# 0.0334f
C842 a_8403_4801# a_9639_4775# 0.0264f
C843 a_8858_4775# a_9152_4775# 0.199f
C844 check[3] a_11289_4394# 1.21e-21
C845 VDD check[3] 0.745f
C846 x36.Q_N a_12102_4296# 1.85e-19
C847 a_12031_4775# a_11966_4801# 4.2e-20
C848 a_11857_4801# a_12147_4801# 0.0282f
C849 a_5844_3239# check[0] 0.051f
C850 a_5372_4112# a_5170_4112# 3.67e-19
C851 a_3599_2340# a_3505_4086# 1.57e-20
C852 a_2389_5648# sel_bit[0] 0.137f
C853 D[5] a_6304_2366# 8.64e-19
C854 a_4018_2366# x20.Q_N 1.31e-20
C855 x48.Q a_4008_4801# 3.94e-19
C856 a_1112_2340# a_1207_2340# 0.0968f
C857 a_4680_3239# x75.Q_N 9.58e-21
C858 a_3912_2366# VDD 0.359f
C859 a_4367_3213# a_4453_4386# 5.72e-19
C860 a_3806_3239# a_3600_4086# 2.44e-19
C861 a_4680_3239# a_3913_4112# 2.16e-19
C862 a_10775_2340# check[3] 2.56e-20
C863 a_5561_3239# a_4855_4775# 4.94e-20
C864 a_4317_3521# VDD 0.0107f
C865 a_2883_5674# a_2463_4775# 6.31e-19
C866 sel_bit[1] a_1508_5167# 5.1e-20
C867 D[3] a_9238_4086# 1.26e-20
C868 a_3900_5167# a_3984_5167# 0.00972f
C869 a_4855_4775# a_4681_4801# 0.197f
C870 a_3453_4801# a_4318_5083# 0.00276f
C871 a_8857_3213# a_8802_2366# 5.71e-21
C872 a_6410_2366# VDD 4.84e-19
C873 a_11630_4086# a_11834_4086# 0.117f
C874 a_6546_2340# a_7185_2366# 0.00316f
C875 x5.X a_8768_5167# 4.18e-19
C876 x20.Q_N a_2579_4801# 0.00429f
C877 a_5896_2340# x27.Q_N 1.79e-19
C878 a_11331_4086# x39.Q_N 0.029f
C879 a_6304_2366# a_8383_2340# 7.3e-21
C880 a_6844_2640# a_6984_2366# 0.00126f
C881 a_11629_4386# a_12102_4296# 0.155f
C882 a_6010_3239# check[5] 2.24e-21
C883 a_8997_3239# VDD 5.47e-21
C884 a_9464_3239# a_9573_3239# 0.00707f
C885 a_4680_3239# x4.X 0.0059f
C886 a_7247_4775# a_9465_4801# 1.86e-21
C887 check[1] a_6845_4386# 0.163f
C888 comparator_out a_2060_2640# 0.113f
C889 comparator_out a_6199_4801# 1.97e-20
C890 a_3373_5674# a_3600_4086# 2.25e-20
C891 a_11544_4775# a_10983_4801# 3.29e-21
C892 a_11076_5167# a_11160_5167# 0.00972f
C893 a_12031_4775# a_11857_4801# 0.197f
C894 a_9172_2366# check[1] 1.35e-19
C895 a_10629_4801# a_11494_5083# 0.00276f
C896 a_6504_2648# x4.X 0.00102f
C897 VDD a_2788_5674# 6.52e-19
C898 a_4926_4296# a_5170_4478# 0.00972f
C899 a_3913_4112# a_4794_4112# 0.00943f
C900 a_4658_4086# a_5372_4112# 6.99e-20
C901 a_4454_4086# a_5897_4086# 3.23e-19
C902 a_4155_4086# a_4593_4112# 0.00276f
C903 a_9101_3521# x4.X 2.91e-19
C904 check[2] a_5562_4801# 4.53e-20
C905 a_8697_4112# a_9173_4478# 0.00133f
C906 VDD a_6547_4086# 0.34f
C907 a_8938_2340# a_9172_2732# 0.00976f
C908 a_8383_2340# a_8802_2366# 0.0397f
C909 a_8696_2366# a_9374_2732# 0.00652f
C910 a_10680_2340# VDD 0.189f
C911 a_9639_4775# a_9710_4296# 2.97e-21
C912 sel_bit[0] a_3619_4801# 8.15e-19
C913 a_9465_4801# a_9442_4086# 2.59e-19
C914 a_9152_4775# x42.Q_N 9.8e-21
C915 a_8683_3605# a_8858_4775# 1.33e-23
C916 a_9754_3239# a_9441_2340# 3.49e-20
C917 a_8857_3213# a_8684_5167# 3.52e-21
C918 D[5] check[0] 0.228f
C919 a_9151_3213# a_8403_4801# 2.05e-21
C920 a_3258_5648# x4.X 3.57e-21
C921 comparator_out x42.Q_N 0.00133f
C922 a_5844_3239# D[5] 5.19e-19
C923 sel_bit[1] x4.X 2.49e-19
C924 comparator_out a_5371_2366# 0.155f
C925 comparator_out a_8402_3239# 0.147f
C926 x77.Y a_3619_4801# 5.26e-21
C927 x4.X a_4794_4112# 0.00375f
C928 a_5844_3239# x72.Q_N 1.07e-19
C929 a_6305_4112# x45.Q_N 0.093f
C930 a_6845_4386# a_7050_4086# 0.153f
C931 a_10155_2366# a_9953_2366# 3.67e-19
C932 x5.X a_7159_5167# 1.05e-19
C933 a_1520_2366# x51.Q_N 0.00553f
C934 a_10680_2340# a_10775_2340# 0.0968f
C935 a_9172_2366# a_9577_2366# 2.46e-21
C936 a_2060_2640# a_2265_2340# 0.153f
C937 D[2] a_11833_2340# 4.68e-20
C938 a_10629_4801# a_10681_4086# 6.04e-19
C939 check[0] a_4767_5167# 1.92e-19
C940 a_6466_4775# a_6606_4801# 0.07f
C941 a_6011_4801# a_6400_4801# 0.0019f
C942 a_5845_4801# a_6978_4801# 2.56e-19
C943 a_6760_4775# a_6931_5083# 0.00652f
C944 eob a_3600_4086# 4.72e-22
C945 x63.Q_N x36.Q_N 4.08e-19
C946 a_9465_4801# a_9574_4801# 0.00707f
C947 a_3619_4801# check[6] 5.82e-21
C948 D[6] a_4657_2340# 2.71e-19
C949 a_6010_3239# a_7953_3239# 1e-20
C950 a_6845_2340# check[6] 3.11e-22
C951 x39.Q_N a_11195_4112# 0.0451f
C952 a_11834_4086# a_12346_4478# 6.69e-20
C953 eob a_1682_4775# 0.0484f
C954 a_11630_4086# a_12548_4112# 0.0708f
C955 a_11833_2340# a_11969_2366# 0.07f
C956 a_11856_3239# a_12102_4296# 2.37e-20
C957 a_12030_3213# x39.Q_N 0.144f
C958 check[5] a_8403_4801# 0.162f
C959 a_8802_2366# x33.Q_N 0.0102f
C960 comparator_out a_11564_2732# 1.8e-19
C961 check[1] a_7264_4394# 6.91e-21
C962 a_2389_5648# a_2788_5674# 2.97e-20
C963 check[4] a_11966_4801# 9.01e-21
C964 a_10795_4801# check[3] 8.42e-19
C965 a_4680_3239# a_4970_3239# 0.0282f
C966 a_4854_3213# a_4789_3239# 4.2e-20
C967 a_1682_4775# x4.A 0.00205f
C968 check[2] a_6305_4112# 1.74e-20
C969 x5.X a_5372_4112# 9.6e-19
C970 x4.X x39.Q_N 0.253f
C971 x48.Q a_3505_4086# 0.0868f
C972 VDD a_6411_4112# 0.00996f
C973 a_2463_4775# a_2289_4801# 0.197f
C974 a_4367_3213# a_5561_3239# 6.04e-19
C975 a_1508_5167# a_1592_5167# 0.00972f
C976 x5.X x27.Q_N 0.00103f
C977 a_8683_3605# x42.Q_N 0.152f
C978 a_9638_3213# a_9442_4086# 2.47e-19
C979 a_9151_3213# a_9710_4296# 1.71e-19
C980 D[6] VDD 0.28f
C981 a_3599_2340# x20.Q_N 3.36e-19
C982 a_4453_2340# a_6304_2366# 3.16e-19
C983 a_8402_3239# a_8683_3605# 0.155f
C984 a_6465_3213# VDD 0.308f
C985 a_4925_2550# a_4793_2366# 0.0258f
C986 a_4452_2640# a_6546_2340# 4.11e-20
C987 a_8236_3239# a_9151_3213# 0.126f
C988 x27.Q_N a_6292_5167# 5.48e-20
C989 a_11628_2640# x39.Q_N 4.61e-20
C990 check[4] a_8697_4112# 3.77e-22
C991 a_11629_2340# a_12102_4296# 6.08e-21
C992 a_7317_2550# x30.Q_N 0.181f
C993 x5.X x36.Q_N 0.00489f
C994 a_9152_4775# a_9873_5083# 0.00185f
C995 a_8684_5167# x33.Q_N 1.74e-20
C996 a_4854_3213# a_4855_4775# 0.00237f
C997 x4.X a_6505_4394# 1.75e-19
C998 a_6304_2366# check[1] 1.25e-21
C999 x48.Q a_1227_4801# 5.44e-21
C1000 a_2479_2648# x4.X 2.86e-19
C1001 a_6845_4386# a_7764_4112# 0.162f
C1002 a_6305_4112# a_6781_4112# 2.87e-21
C1003 a_7050_4086# a_7264_4394# 0.0104f
C1004 a_6846_4086# a_7562_4478# 0.0018f
C1005 a_7246_3213# a_6845_4386# 3.78e-19
C1006 a_6759_3213# a_6846_4086# 1.61e-19
C1007 a_6010_3239# x45.Q_N 0.346f
C1008 VDD a_2375_5167# 0.00488f
C1009 a_7049_2340# a_6982_2732# 9.46e-19
C1010 a_8696_2366# x42.Q_N 6.41e-20
C1011 x57.Q_N a_6504_2648# 2.02e-20
C1012 a_9237_2340# a_9238_4086# 1.55e-19
C1013 a_6304_2366# a_7763_2366# 5.76e-21
C1014 a_6844_2640# a_7263_2648# 2.46e-19
C1015 a_9441_2340# a_9237_4386# 1.26e-21
C1016 a_5991_2340# VDD 0.561f
C1017 a_8402_3239# a_8696_2366# 5.94e-19
C1018 a_8857_3213# a_8383_2340# 2.5e-19
C1019 D[7] a_2401_2366# 4.38e-19
C1020 a_7073_4801# check[5] 6.72e-20
C1021 x75.Q a_5897_4086# 0.00123f
C1022 check[4] a_11857_4801# 4.17e-20
C1023 a_8802_2366# check[1] 0.00244f
C1024 a_1682_4775# a_1926_5083# 0.0104f
C1025 a_1227_4801# a_2147_5083# 1.09e-19
C1026 a_4155_4086# a_4658_4086# 0.00187f
C1027 a_4453_4386# a_4454_4086# 0.75f
C1028 a_3600_4086# x48.Q_N 0.124f
C1029 a_3913_4112# a_4926_4296# 0.0633f
C1030 a_6844_2640# a_6845_4386# 1.32e-20
C1031 x5.X a_11629_4386# 0.00326f
C1032 a_6304_2366# a_7050_4086# 7.14e-22
C1033 a_6546_2340# a_6846_4086# 3.47e-21
C1034 x77.Y a_3452_3239# 0.51f
C1035 a_9374_2732# VDD 0.0163f
C1036 a_12346_4478# a_12548_4112# 8.94e-19
C1037 a_8288_2340# a_9237_2340# 1.03e-19
C1038 a_8236_3239# check[5] 0.00639f
C1039 D[0] a_8237_4801# 1.99e-20
C1040 a_10794_3239# a_11389_3239# 0.00118f
C1041 a_10982_3239# a_11159_3605# 8.94e-19
C1042 a_11543_3213# a_11493_3521# 1.21e-20
C1043 a_11942_3605# VDD 0.00371f
C1044 a_4453_2340# check[0] 0.00712f
C1045 a_12147_4801# a_12102_4296# 1.9e-20
C1046 comparator_out a_4452_2640# 0.109f
C1047 x4.X a_4926_4296# 0.0211f
C1048 check[1] check[0] 0.0116f
C1049 check[2] x48.Q 0.0879f
C1050 a_9573_3239# x4.X 1.05e-19
C1051 a_5844_3239# check[1] 2.07e-22
C1052 a_1508_5167# x27.D 4.66e-22
C1053 a_1976_4775# a_3170_4801# 6.04e-19
C1054 a_9238_4086# a_11331_4086# 1.67e-21
C1055 a_9710_4296# a_10776_4086# 7.98e-21
C1056 x42.Q_N a_9578_4112# 0.00172f
C1057 a_9638_3213# a_10156_4112# 2.07e-19
C1058 a_9236_2640# a_9953_2366# 0.00105f
C1059 check[6] a_6710_5083# 2.57e-21
C1060 VDD a_8858_4775# 0.488f
C1061 a_6984_2366# check[5] 9.43e-20
C1062 a_8857_3213# x33.Q_N 5.46e-19
C1063 comparator_out a_7561_2732# 8.23e-19
C1064 comparator_out a_10628_3239# 0.148f
C1065 a_3452_3239# check[6] 1.79e-20
C1066 check[0] a_3877_5674# 0.00787f
C1067 x5.X a_1976_4775# 0.00314f
C1068 check[0] a_7050_4086# 1.2e-19
C1069 D[1] x39.Q_N 3.4e-19
C1070 a_1520_2366# x54.Q_N 5.89e-21
C1071 a_6010_3239# a_6198_3239# 0.163f
C1072 a_6291_3605# a_7246_3213# 4.7e-22
C1073 a_6465_3213# a_7072_3239# 0.00187f
C1074 a_2061_2340# a_4453_2340# 0.00176f
C1075 a_11833_2340# a_12101_2550# 0.205f
C1076 a_11629_2340# x63.Q_N 1.07e-19
C1077 a_5844_3239# a_7050_4086# 0.00195f
C1078 comparator_out a_6846_4086# 3.21e-20
C1079 a_11544_4775# x39.Q_N 9.93e-21
C1080 a_11857_4801# a_11834_4086# 2.59e-19
C1081 a_12031_4775# a_12102_4296# 2.97e-21
C1082 a_8383_2340# x33.Q_N 0.142f
C1083 a_3618_3239# a_3599_2340# 3.73e-19
C1084 a_3452_3239# a_3912_2366# 1.89e-19
C1085 D[7] eob 2.52e-20
C1086 x4.X x27.D 0.00252f
C1087 x5.X a_4155_4086# 7.39e-20
C1088 a_2060_2640# a_1511_4112# 0.00164f
C1089 x48.Q a_4074_4775# 0.00395f
C1090 x5.X a_12048_4394# 1.32e-19
C1091 a_4073_3213# a_3806_3239# 6.99e-20
C1092 x48.Q x20.Q_N 0.0441f
C1093 a_3618_3239# a_3983_3605# 4.45e-20
C1094 a_3452_3239# a_4317_3521# 0.00276f
C1095 a_4367_3213# a_4854_3213# 0.273f
C1096 a_4657_2340# a_5371_2366# 6.99e-20
C1097 a_2979_2366# x20.Q_N 0.00156f
C1098 a_4925_2550# a_5169_2732# 0.00972f
C1099 a_4453_2340# D[5] 0.338f
C1100 a_7953_3239# a_8236_3239# 8.18e-19
C1101 VDD a_6199_4801# 0.109f
C1102 a_6759_3213# a_6546_2340# 2.17e-19
C1103 a_7246_3213# a_6304_2366# 8.4e-19
C1104 a_2060_2640# VDD 0.329f
C1105 a_6010_3239# a_7049_2340# 0.00154f
C1106 a_6465_3213# a_6845_2340# 0.00199f
C1107 check[5] a_9370_4801# 7.95e-20
C1108 a_11769_4112# a_11630_4086# 2.56e-19
C1109 a_11970_4112# a_11629_4386# 0.00118f
C1110 a_11762_4801# check[3] 7.79e-21
C1111 x72.Q_N check[1] 4.68e-20
C1112 x4.X a_6760_4775# 0.104f
C1113 a_1207_2340# x4.X 0.117f
C1114 a_2463_4775# a_3807_4801# 8.26e-21
C1115 check[2] a_8403_4801# 4.08e-19
C1116 VDD x42.Q_N 0.457f
C1117 a_11629_2340# x5.X 4.23e-20
C1118 a_9173_4112# a_9578_4112# 2.46e-21
C1119 a_10681_4086# a_10776_4086# 0.0968f
C1120 a_1822_4801# a_2194_4801# 3.34e-19
C1121 a_5371_2366# VDD 0.109f
C1122 a_6304_2366# a_6844_2640# 0.139f
C1123 a_8402_3239# VDD 0.275f
C1124 a_5991_2340# a_6845_2340# 0.0492f
C1125 x69.Q_N x42.Q_N 3.92e-19
C1126 a_8402_3239# x69.Q_N 4.5e-21
C1127 a_9464_3239# a_9550_3605# 0.00976f
C1128 a_7480_3521# VDD 0.00506f
C1129 x27.Q_N x30.Q_N 2.3e-20
C1130 a_7362_3239# a_7181_3239# 4.11e-20
C1131 a_9441_2340# x30.Q_N 9.31e-21
C1132 a_5561_3239# a_4454_4086# 4.72e-19
C1133 a_8383_2340# check[1] 0.0126f
C1134 x4.X a_9238_4086# 0.0468f
C1135 a_4018_2366# x4.X 3.78e-20
C1136 VDD a_4113_4394# 0.00555f
C1137 a_6605_3239# x4.X 0.00267f
C1138 a_4855_4775# a_4658_4086# 4.44e-19
C1139 a_4368_4775# a_4926_4296# 2.85e-19
C1140 a_7318_4296# x42.Q_N 8.46e-20
C1141 a_8236_3239# x45.Q_N 1.49e-19
C1142 a_6844_2640# a_8802_2366# 1.71e-20
C1143 a_7763_2366# a_8383_2340# 8.26e-21
C1144 VDD a_4539_5083# 0.0172f
C1145 a_6977_3239# x45.Q_N 0.00399f
C1146 D[1] a_9573_3239# 9.28e-21
C1147 check[3] a_11089_4112# 0.0033f
C1148 VDD a_11715_5083# 0.0163f
C1149 a_2883_5674# a_2969_6040# 0.0136f
C1150 a_5844_3239# a_7246_3213# 0.0492f
C1151 comparator_out a_6759_3213# 7.49e-19
C1152 x4.X a_2579_4801# 0.0171f
C1153 a_5372_4112# a_5992_4086# 8.26e-21
C1154 a_8288_2340# x4.X 0.00317f
C1155 x5.X a_5845_4801# 0.27f
C1156 check[2] a_7073_4801# 4.32e-20
C1157 x4.X a_9755_4801# 0.00557f
C1158 a_6011_4801# a_6466_4775# 0.153f
C1159 sel_bit[0] a_3600_4086# 3.59e-19
C1160 a_11564_2732# VDD 0.00371f
C1161 a_5845_4801# a_6292_5167# 0.15f
C1162 x77.Y a_5088_3521# 8.16e-21
C1163 check[0] a_3453_4801# 0.00279f
C1164 a_8938_2340# a_9172_2366# 0.00707f
C1165 a_8696_2366# a_9376_2366# 3.73e-19
C1166 a_9236_2640# a_10680_2340# 6.83e-19
C1167 x5.X a_12147_4801# 2.09e-19
C1168 a_6844_2640# check[0] 2.7e-19
C1169 a_11389_3239# a_11761_3239# 3.34e-19
C1170 x77.Y a_3600_4086# 1.36e-19
C1171 check[1] a_9377_4112# 3.4e-20
C1172 comparator_out a_6546_2340# 0.00104f
C1173 a_5844_3239# a_6844_2640# 6.01e-20
C1174 check[1] x33.Q_N 0.0011f
C1175 check[2] a_9710_4296# 0.00118f
C1176 x5.X a_8384_4086# 0.0202f
C1177 sel_bit[0] a_1682_4775# 7.55e-20
C1178 a_8236_3239# check[2] 6.24e-22
C1179 x27.D a_4368_4775# 0.00307f
C1180 check[5] a_6845_4386# 0.0306f
C1181 a_7954_4801# a_6846_4086# 6.67e-19
C1182 VDD a_9173_4112# 3.55e-19
C1183 a_10775_2340# a_11564_2732# 7.71e-20
C1184 a_11088_2366# a_11288_2648# 0.00185f
C1185 a_12346_4112# x4.X 6.38e-19
C1186 VDD a_9873_5083# 0.00506f
C1187 a_7763_2366# x33.Q_N 1.34e-20
C1188 a_10794_3239# x33.Q_N 3.79e-20
C1189 a_3618_3239# x48.Q 2.51e-19
C1190 comparator_out a_9655_2648# 7e-19
C1191 a_3452_3239# D[6] 2.82e-19
C1192 x4.X a_9954_4478# 9.15e-19
C1193 x5.X a_4855_4775# 0.00928f
C1194 a_8289_4086# x42.Q_N 0.18f
C1195 x4.X a_8998_4801# 7.25e-19
C1196 a_8697_4112# a_8939_4086# 0.124f
C1197 a_8384_4086# a_9237_4386# 0.0264f
C1198 a_4855_4775# a_6292_5167# 7.98e-21
C1199 a_3912_2366# x54.Q_N 0.00553f
C1200 x5.X a_12031_4775# 0.00483f
C1201 a_1762_2340# x20.Q_N 0.162f
C1202 a_6759_3213# a_8683_3605# 4.38e-20
C1203 a_7072_3239# a_8402_3239# 3.9e-20
C1204 a_12737_3239# x39.Q_N 3.23e-19
C1205 a_4452_2640# a_4657_2340# 0.153f
C1206 a_7246_3213# x72.Q_N 0.124f
C1207 a_8684_5167# a_9639_4775# 4.7e-22
C1208 a_8237_4801# a_8768_5167# 0.0018f
C1209 a_8403_4801# a_8591_4801# 0.162f
C1210 a_8858_4775# a_9465_4801# 0.00187f
C1211 a_9577_2366# x33.Q_N 0.0403f
C1212 a_11543_3213# check[3] 1.04e-19
C1213 a_12030_3213# a_12738_4801# 3.19e-20
C1214 x4.X a_5562_4801# 0.00612f
C1215 x48.Q a_5170_4478# 5.12e-20
C1216 a_3599_2340# a_3913_4112# 5.05e-21
C1217 a_5561_3239# x75.Q 0.0955f
C1218 x4.X a_12738_4801# 0.00262f
C1219 D[1] a_9238_4086# 3.36e-19
C1220 x48.Q a_5089_5083# 1.17e-19
C1221 a_5371_2366# a_6845_2340# 3.65e-21
C1222 D[5] a_6844_2640# 4.09e-20
C1223 D[7] a_1520_2366# 0.00164f
C1224 a_4452_2640# VDD 0.273f
C1225 D[0] a_8997_3239# 1.6e-19
C1226 a_2853_5648# a_1511_4112# 6.37e-19
C1227 a_4367_3213# a_4658_4086# 0.0014f
C1228 a_4854_3213# a_4454_4086# 7.94e-19
C1229 a_11330_2340# check[3] 1.32e-19
C1230 check[1] a_9954_4112# 5.77e-22
C1231 VDD a_2853_5648# 0.413f
C1232 a_4766_3605# VDD 0.00394f
C1233 sel_bit[1] a_2463_4775# 5.3e-20
C1234 a_3599_2340# x4.X 0.117f
C1235 x5.X a_9173_4478# 3.15e-19
C1236 check[2] a_10681_4086# 0.126f
C1237 a_4074_4775# a_4318_5083# 0.0104f
C1238 a_3619_4801# a_4539_5083# 1.09e-19
C1239 a_10628_3239# VDD 0.791f
C1240 a_7561_2732# VDD 0.0042f
C1241 x5.X a_7182_4801# 5.34e-20
C1242 a_6844_2640# a_8383_2340# 3.42e-19
C1243 a_10628_3239# a_11249_3213# 0.117f
C1244 a_11834_4086# a_12102_4296# 0.205f
C1245 a_6845_2340# a_7185_2366# 6.04e-20
C1246 a_7049_2340# a_6984_2366# 9.75e-19
C1247 a_4592_2366# x27.Q_N 0.00474f
C1248 a_11630_4086# x39.Q_N 0.00117f
C1249 a_9369_3239# VDD 6.2e-19
C1250 a_3983_3605# x4.X 0.00103f
C1251 a_6760_4775# a_7363_4801# 0.0552f
C1252 x69.Q_N a_10628_3239# 2.94e-19
C1253 check[1] a_7050_4086# 7.72e-19
C1254 comparator_out a_2265_2340# 0.00311f
C1255 a_10795_4801# a_11715_5083# 1.09e-19
C1256 a_11250_4775# a_11494_5083# 0.0104f
C1257 a_9577_2366# check[1] 4.4e-19
C1258 a_4453_4386# a_4794_4112# 0.00118f
C1259 a_6982_2732# x4.X 9.81e-19
C1260 VDD a_3671_5674# 7.34e-19
C1261 a_4155_4086# a_5992_4086# 1.86e-21
C1262 a_4454_4086# a_4593_4112# 2.56e-19
C1263 a_9550_3605# x4.X 4.4e-19
C1264 a_9238_4086# a_8897_4394# 1.25e-19
C1265 D[4] a_6846_4086# 1.26e-20
C1266 a_8697_4112# a_8803_4112# 0.051f
C1267 a_8939_4086# a_9375_4478# 0.00412f
C1268 a_9237_4386# a_9173_4478# 2.13e-19
C1269 VDD a_6846_4086# 0.805f
C1270 a_8696_2366# a_9655_2648# 1.21e-20
C1271 a_8938_2340# a_8802_2366# 0.0282f
C1272 a_9236_2640# a_9374_2732# 1.09e-19
C1273 D[4] a_9376_2366# 7.47e-20
C1274 a_9376_2366# VDD 6.2e-19
C1275 a_10628_3239# a_10775_2340# 8.35e-19
C1276 a_6304_2366# check[5] 1.15e-20
C1277 sel_bit[0] a_3900_5167# 2.68e-19
C1278 a_8402_3239# a_9465_4801# 6.75e-21
C1279 reset a_897_4112# 0.00119f
C1280 a_621_4112# x3.A 0.129f
C1281 eob a_1976_4775# 0.0525f
C1282 x77.Y a_3900_5167# 7.98e-21
C1283 comparator_out a_8683_3605# 0.0011f
C1284 x4.X a_6305_4112# 0.11f
C1285 a_6846_4086# a_7318_4296# 0.15f
C1286 a_6845_4386# x45.Q_N 0.00117f
C1287 a_11970_4112# a_12031_4775# 1.79e-20
C1288 check[0] a_4019_4112# 1.03e-20
C1289 x5.X a_6400_4801# 2.84e-19
C1290 a_2060_2640# x51.Q_N 4.18e-21
C1291 a_2061_2340# a_2533_2550# 0.15f
C1292 a_6760_4775# a_6606_4801# 0.00943f
C1293 a_5845_4801# x30.Q_N 2.24e-19
C1294 a_6466_4775# a_6978_4801# 9.75e-19
C1295 a_6292_5167# a_6400_4801# 0.00812f
C1296 a_7247_4775# a_7159_5167# 7.71e-20
C1297 a_7073_4801# a_6931_5083# 0.00412f
C1298 a_2389_5648# a_2853_5648# 0.202f
C1299 a_6844_2640# x33.Q_N 0.00104f
C1300 x33.Q_N a_10629_4801# 7.17e-19
C1301 comparator_out a_8696_2366# 0.00714f
C1302 a_4368_4775# a_5562_4801# 6.04e-19
C1303 a_3900_5167# check[6] 1.4e-21
C1304 D[6] x54.Q_N 0.00317f
C1305 x5.X check[4] 0.167f
C1306 a_6465_3213# D[0] 1.23e-20
C1307 a_12102_4296# a_12548_4112# 0.0367f
C1308 a_11389_3239# a_10776_4086# 1.16e-20
C1309 a_12101_2550# a_12345_2366# 0.00812f
C1310 a_10982_3239# x39.Q_N 7.52e-20
C1311 check[5] a_8684_5167# 0.00124f
C1312 check[1] a_7764_4112# 0.165f
C1313 check[2] a_2993_5674# 0.0021f
C1314 a_5844_3239# check[5] 1.81e-20
C1315 a_11076_5167# check[3] 5.35e-19
C1316 a_11544_4775# a_12738_4801# 6.04e-19
C1317 a_7246_3213# check[1] 0.00245f
C1318 x75.Q_N a_6010_3239# 2.12e-19
C1319 check[2] a_6845_4386# 1.41e-20
C1320 x48.Q a_3913_4112# 8.72e-19
C1321 a_5845_4801# a_5992_4086# 0.00159f
C1322 D[2] x5.X 0.0046f
C1323 VDD a_7562_4478# 0.0042f
C1324 a_1976_4775# a_1926_5083# 1.21e-20
C1325 a_4854_3213# x75.Q 0.0108f
C1326 a_6759_3213# VDD 0.353f
C1327 a_9464_3239# a_9710_4296# 2.37e-20
C1328 a_4154_2340# x20.Q_N 2.93e-20
C1329 a_9638_3213# x42.Q_N 0.144f
C1330 a_7246_3213# a_7763_2366# 2.38e-19
C1331 a_4452_2640# a_6845_2340# 2.9e-21
C1332 a_4925_2550# a_6304_2366# 9.52e-21
C1333 a_10346_4801# a_9238_4086# 6.67e-19
C1334 check[4] a_9237_4386# 0.028f
C1335 a_8857_3213# a_9151_3213# 0.199f
C1336 a_8402_3239# a_9638_3213# 0.0264f
C1337 a_8236_3239# a_9464_3239# 0.0334f
C1338 a_4453_2340# a_6844_2640# 4e-20
C1339 a_11833_2340# x39.Q_N 1.11e-19
C1340 x72.Q_N a_9151_3213# 2.97e-20
C1341 a_9639_4775# x33.Q_N 0.126f
C1342 check[1] a_3453_4801# 9.29e-20
C1343 a_2853_5648# a_3619_4801# 3.82e-19
C1344 a_6844_2640# check[1] 7.55e-20
C1345 x4.X a_6983_4478# 0.00114f
C1346 x48.Q x4.X 0.188f
C1347 a_2979_2366# x4.X 4.09e-19
C1348 a_6010_3239# x4.X 0.0446f
C1349 a_7050_4086# a_7764_4112# 6.99e-20
C1350 a_6846_4086# a_8289_4086# 3.23e-19
C1351 a_6547_4086# a_6985_4112# 0.00276f
C1352 a_7318_4296# a_7562_4478# 0.00972f
C1353 a_6305_4112# a_7186_4112# 0.00943f
C1354 a_7246_3213# a_7050_4086# 2.47e-19
C1355 a_6759_3213# a_7318_4296# 1.71e-19
C1356 a_6291_3605# x45.Q_N 0.152f
C1357 VDD a_1616_4801# 6e-19
C1358 a_9236_2640# x42.Q_N 4.61e-20
C1359 a_6844_2640# a_7763_2366# 0.159f
C1360 a_6546_2340# VDD 0.177f
C1361 a_9237_2340# a_9710_4296# 6.08e-21
C1362 a_7049_2340# a_7263_2648# 0.0104f
C1363 a_6845_2340# a_7561_2732# 0.0018f
C1364 a_9151_3213# a_8383_2340# 9.06e-19
C1365 a_8857_3213# a_8938_2340# 4.18e-20
C1366 a_8402_3239# a_9236_2640# 4.04e-20
C1367 a_8236_3239# a_9237_2340# 6.52e-20
C1368 a_8683_3605# a_8696_2366# 1.71e-19
C1369 a_10794_3239# a_10629_4801# 8.16e-19
C1370 a_10628_3239# a_10795_4801# 9.04e-19
C1371 a_1227_4801# a_1822_4801# 0.00118f
C1372 a_4454_4086# a_4658_4086# 0.117f
C1373 a_4155_4086# x48.Q_N 9.58e-21
C1374 a_4453_4386# a_4926_4296# 0.155f
C1375 x5.X a_11834_4086# 3.65e-19
C1376 a_6845_2340# a_6846_4086# 1.55e-19
C1377 a_6304_2366# x45.Q_N 6.37e-20
C1378 a_7049_2340# a_6845_4386# 1.26e-21
C1379 x77.Y a_4073_3213# 0.201f
C1380 a_9655_2648# VDD 0.00984f
C1381 a_6780_2366# x27.Q_N 9.28e-21
C1382 a_8383_2340# a_8938_2340# 0.197f
C1383 a_10628_3239# a_12264_3521# 1.25e-19
C1384 a_11543_3213# a_11942_3605# 0.00133f
C1385 x72.Q_N check[5] 0.00322f
C1386 a_11075_3605# a_11389_3239# 0.0258f
C1387 a_10794_3239# a_11761_3239# 0.00126f
C1388 x30.Q_N a_7182_4801# 7.02e-20
C1389 a_5844_3239# a_7953_3239# 1.03e-19
C1390 comparator_out a_4657_2340# 0.00586f
C1391 a_9172_2732# x4.X 4.32e-19
C1392 a_11714_3521# x4.X 9.99e-19
C1393 a_1520_2366# a_1720_2648# 0.00185f
C1394 a_2463_4775# x27.D 0.00431f
C1395 a_9238_4086# a_11630_4086# 1.37e-19
C1396 a_1207_2340# a_1996_2732# 7.71e-20
C1397 a_8697_4112# x39.Q_N 1.05e-20
C1398 a_9237_2340# a_11288_2648# 4.06e-20
C1399 a_8383_2340# check[5] 3.32e-21
C1400 comparator_out a_1511_4112# 8.67e-19
C1401 VDD a_9152_4775# 0.449f
C1402 a_9151_3213# x33.Q_N 0.00498f
C1403 comparator_out VDD 1.51f
C1404 comparator_out D[4] 0.00125f
C1405 comparator_out a_11249_3213# 4.81e-19
C1406 x77.Y x27.Q_N 0.00357f
C1407 comparator_out x69.Q_N 1.46e-19
C1408 x4.X a_8403_4801# 0.005f
C1409 x5.X a_2289_4801# 0.00166f
C1410 a_7246_3213# a_7764_4112# 2.07e-19
C1411 a_8696_2366# a_9578_4112# 1.26e-20
C1412 check[0] x45.Q_N 0.0173f
C1413 a_6291_3605# a_6198_3239# 0.0367f
C1414 a_6759_3213# a_7072_3239# 0.124f
C1415 a_6465_3213# a_6375_3605# 6.69e-20
C1416 a_2060_2640# x54.Q_N 1.48e-19
C1417 a_6010_3239# a_4970_3239# 7.73e-20
C1418 a_5844_3239# x45.Q_N 0.0434f
C1419 a_6400_4801# x30.Q_N 3.71e-20
C1420 a_8938_2340# x33.Q_N 0.16f
C1421 comparator_out a_10775_2340# 0.00442f
C1422 a_3899_3605# a_3599_2340# 3.9e-20
C1423 a_3452_3239# a_4452_2640# 6.01e-20
C1424 a_4073_3213# a_3912_2366# 0.0014f
C1425 x33.Q_N a_11184_4801# 3.99e-20
C1426 sel_bit[1] a_897_4112# 1.46e-20
C1427 x5.X a_4454_4086# 0.258f
C1428 check[6] a_5372_4112# 0.00256f
C1429 a_2265_2340# a_1511_4112# 0.00119f
C1430 x48.Q a_4368_4775# 0.0017f
C1431 x5.X a_12548_4112# 5.39e-19
C1432 D[0] x42.Q_N 3.91e-19
C1433 a_3618_3239# a_4538_3521# 1.09e-19
C1434 a_4854_3213# a_4680_3239# 0.197f
C1435 a_3899_3605# a_3983_3605# 0.00972f
C1436 a_4073_3213# a_4317_3521# 0.0104f
C1437 D[0] a_8402_3239# 0.00637f
C1438 a_2265_2340# VDD 0.326f
C1439 x27.Q_N check[6] 0.934f
C1440 VDD a_4971_4801# 0.0111f
C1441 a_7246_3213# a_6844_2640# 3.43e-19
C1442 a_6759_3213# a_6845_2340# 2.19e-19
C1443 x72.Q_N a_7953_3239# 0.178f
C1444 clk_sar a_621_4112# 9.27e-21
C1445 a_7362_3239# x30.Q_N 0.00342f
C1446 a_12737_3239# a_12738_4801# 9.85e-20
C1447 check[5] x33.Q_N 3.66e-21
C1448 x75.Q a_5896_2340# 0.00129f
C1449 a_9151_3213# check[1] 1.78e-20
C1450 a_11565_4112# x39.Q_N 0.0014f
C1451 a_11970_4112# a_11834_4086# 0.07f
C1452 x36.Q_N check[3] 1.17f
C1453 a_1762_2340# x4.X 0.00671f
C1454 x4.X a_7073_4801# 0.00316f
C1455 check[2] a_8684_5167# 1.92e-19
C1456 a_2463_4775# a_2579_4801# 0.0397f
C1457 a_1976_4775# a_2398_4801# 2.87e-21
C1458 check[2] check[0] 0.872f
C1459 a_8683_3605# VDD 0.176f
C1460 a_3912_2366# x27.Q_N 0.0928f
C1461 a_1822_4801# x20.Q_N 1.36e-19
C1462 a_5991_2340# a_7317_2550# 4.7e-22
C1463 a_5845_4801# a_8237_4801# 0.00176f
C1464 a_6304_2366# a_7049_2340# 0.199f
C1465 a_9638_3213# a_10628_3239# 0.00116f
C1466 a_9151_3213# a_10794_3239# 1.89e-19
C1467 a_6546_2340# a_6845_2340# 0.0334f
C1468 x60.Q_N x30.Q_N 8.43e-20
C1469 a_9151_3213# a_9872_3521# 0.00185f
C1470 a_4854_3213# a_4794_4112# 4.45e-20
C1471 a_11564_2366# check[3] 2.19e-20
C1472 a_8938_2340# check[1] 0.00112f
C1473 a_3600_4086# a_4113_4394# 0.00945f
C1474 x4.X a_9710_4296# 0.021f
C1475 a_5169_2732# x4.X 1.17e-19
C1476 a_8236_3239# x4.X 0.0456f
C1477 VDD a_4591_4478# 0.0172f
C1478 a_6977_3239# x4.X 4.96e-19
C1479 a_4681_4801# a_4926_4296# 3.59e-20
C1480 x72.Q_N x45.Q_N 3.9e-19
C1481 a_6410_2366# x27.Q_N 8.39e-20
C1482 a_8237_4801# a_8384_4086# 0.00159f
C1483 check[0] a_6781_4112# 9.63e-22
C1484 VDD a_4214_4801# 0.035f
C1485 a_8696_2366# VDD 0.348f
C1486 D[4] a_8696_2366# 8.79e-19
C1487 a_3648_5972# a_3258_5648# 8.72e-19
C1488 sel_bit[0] a_1976_4775# 1.72e-19
C1489 a_6198_3239# check[0] 0.00621f
C1490 comparator_out a_8289_4086# 2.05e-21
C1491 check[3] a_11629_4386# 0.138f
C1492 a_2883_5674# a_3373_5674# 4.47e-19
C1493 a_12738_4801# a_11630_4086# 6.67e-19
C1494 VDD a_11390_4801# 0.0332f
C1495 a_5844_3239# a_6198_3239# 0.0708f
C1496 comparator_out a_7072_3239# 1.93e-19
C1497 check[1] check[5] 0.343f
C1498 a_5897_4086# a_6305_4112# 4.37e-19
C1499 a_4593_4112# a_4794_4112# 3.34e-19
C1500 x5.X a_6466_4775# 0.00314f
C1501 a_11194_2366# VDD 4.84e-19
C1502 a_5845_4801# a_7247_4775# 0.0492f
C1503 a_6466_4775# a_6292_5167# 0.205f
C1504 a_6011_4801# a_6760_4775# 0.139f
C1505 a_11249_3213# a_11194_2366# 5.71e-21
C1506 a_7763_2366# check[5] 0.0034f
C1507 check[0] a_4074_4775# 5.86e-19
C1508 a_8938_2340# a_9577_2366# 0.00316f
C1509 a_9236_2640# a_9376_2366# 0.00126f
C1510 VDD a_7954_4801# 0.193f
C1511 a_8696_2366# a_10775_2340# 6.25e-21
C1512 a_7049_2340# check[0] 4.27e-19
C1513 a_9152_4775# a_10795_4801# 8.44e-20
C1514 a_9639_4775# a_10629_4801# 0.00116f
C1515 a_10680_2340# x36.Q_N 3.7e-19
C1516 x77.Y a_4155_4086# 0.00176f
C1517 comparator_out a_6845_2340# 0.182f
C1518 a_5844_3239# a_7049_2340# 4.77e-19
C1519 comparator_out a_10795_4801# 2.89e-21
C1520 a_11288_2648# x4.X 0.00102f
C1521 x5.X a_8939_4086# 0.00115f
C1522 x27.D a_4681_4801# 2.31e-21
C1523 VDD a_9578_4112# 0.0326f
C1524 a_10794_3239# a_10776_4086# 3.48e-19
C1525 a_10628_3239# a_11089_4112# 2.21e-19
C1526 a_11330_2340# a_11564_2732# 0.00976f
C1527 a_11088_2366# a_11766_2732# 0.00652f
C1528 a_10775_2340# a_11194_2366# 0.0397f
C1529 eob a_2883_5674# 6.72e-19
C1530 x75.Q x5.X 0.0011f
C1531 comparator_out a_10155_2366# 0.155f
C1532 a_11970_4112# a_12101_2550# 1.72e-22
C1533 x4.X a_10681_4086# 0.0036f
C1534 x5.X a_3807_4801# 5.48e-19
C1535 a_6985_4112# x42.Q_N 1.96e-20
C1536 a_8939_4086# a_9237_4386# 0.137f
C1537 a_8697_4112# a_9238_4086# 0.125f
C1538 x5.A a_897_4112# 5.71e-20
C1539 x4.X a_9370_4801# 5.55e-19
C1540 a_2061_2340# x20.Q_N 0.0469f
C1541 a_7246_3213# a_9151_3213# 3.71e-20
C1542 a_4452_2640# x54.Q_N 5.46e-21
C1543 a_4453_2340# a_4925_2550# 0.15f
C1544 x5.X a_10983_4801# 0.00551f
C1545 a_11088_2366# x33.Q_N 8.24e-20
C1546 check[3] a_12048_4394# 5.14e-21
C1547 a_9152_4775# a_9465_4801# 0.124f
C1548 a_8684_5167# a_8591_4801# 0.0367f
C1549 a_8858_4775# a_8768_5167# 6.69e-20
C1550 a_8403_4801# a_7363_4801# 4.14e-20
C1551 a_7953_3239# check[1] 0.00311f
C1552 a_10345_3239# x42.Q_N 3.23e-19
C1553 a_8236_3239# D[1] 7.04e-20
C1554 D[6] x27.Q_N 0.00313f
C1555 a_8402_3239# a_10345_3239# 7.94e-21
C1556 D[5] a_7049_2340# 7e-20
C1557 a_4657_2340# VDD 0.307f
C1558 a_4213_3239# a_4585_3239# 3.34e-19
C1559 D[7] a_2060_2640# 1.7e-19
C1560 D[0] a_9369_3239# 5.51e-20
C1561 a_1112_2340# a_2061_2340# 1.03e-19
C1562 a_2853_5648# a_3600_4086# 2.47e-19
C1563 a_4854_3213# a_4926_4296# 3.74e-20
C1564 a_11629_2340# check[3] 0.0405f
C1565 a_4680_3239# a_4658_4086# 4.33e-20
C1566 a_4007_3239# VDD 2.82e-19
C1567 a_4154_2340# x4.X 0.00377f
C1568 x20.Q_N a_4389_4478# 3.31e-21
C1569 check[2] a_9377_4112# 6.45e-20
C1570 VDD a_1511_4112# 1.55f
C1571 D[0] a_6846_4086# 3.2e-19
C1572 a_3807_4801# a_3984_5167# 8.94e-19
C1573 check[5] a_7764_4112# 0.00263f
C1574 a_3619_4801# a_4214_4801# 0.00118f
C1575 a_4368_4775# a_4318_5083# 1.21e-20
C1576 VDD a_11289_4394# 0.00506f
C1577 D[4] VDD 0.221f
C1578 a_10794_3239# a_11075_3605# 0.155f
C1579 a_11249_3213# VDD 0.308f
C1580 a_10628_3239# a_11543_3213# 0.126f
C1581 check[2] x33.Q_N 0.0366f
C1582 a_12102_4296# x39.Q_N 0.00244f
C1583 a_5991_2340# x27.Q_N 1.43e-19
C1584 x5.X a_9323_5083# 5.14e-19
C1585 a_7317_2550# a_7185_2366# 0.0258f
C1586 a_6844_2640# a_8938_2340# 3.87e-20
C1587 a_6845_2340# a_8696_2366# 3.1e-19
C1588 a_7246_3213# check[5] 0.00432f
C1589 a_4538_3521# x4.X 0.00211f
C1590 x69.Q_N VDD 0.0716f
C1591 a_7073_4801# a_7363_4801# 0.0282f
C1592 a_7247_4775# a_7182_4801# 4.2e-20
C1593 check[1] x45.Q_N 0.00102f
C1594 a_1061_4801# a_1511_4112# 0.00351f
C1595 a_11544_4775# a_11494_5083# 1.21e-20
C1596 a_10983_4801# a_11160_5167# 8.94e-19
C1597 a_10795_4801# a_11390_4801# 0.00118f
C1598 a_1062_5674# sel_bit[1] 0.039f
C1599 x77.Y a_4789_3239# 7.87e-19
C1600 a_7263_2648# x4.X 2.86e-19
C1601 a_4658_4086# a_4794_4112# 0.07f
C1602 a_4453_4386# a_6305_4112# 8.96e-20
C1603 VDD a_1061_4801# 0.901f
C1604 a_4454_4086# a_5992_4086# 2.98e-19
C1605 a_3618_3239# a_5844_3239# 4e-20
C1606 a_3452_3239# comparator_out 6.64e-19
C1607 a_8791_3239# x4.X 6.32e-19
C1608 x42.Q_N a_7562_4112# 2.85e-21
C1609 a_9238_4086# a_9375_4478# 0.00907f
C1610 VDD a_7318_4296# 0.317f
C1611 check[6] a_5845_4801# 0.416f
C1612 a_1207_2340# a_897_4112# 6.9e-19
C1613 a_5562_4801# a_6011_4801# 4.06e-19
C1614 a_9236_2640# a_9655_2648# 2.46e-19
C1615 a_10775_2340# VDD 0.561f
C1616 x60.Q_N a_8896_2648# 2.02e-20
C1617 a_9441_2340# a_9374_2732# 9.46e-19
C1618 a_8696_2366# a_10155_2366# 4.94e-21
C1619 a_6844_2640# check[5] 0.0314f
C1620 a_11249_3213# a_10775_2340# 2.5e-19
C1621 a_10794_3239# a_11088_2366# 5.94e-19
C1622 a_9638_3213# a_9152_4775# 1.06e-20
C1623 a_9151_3213# a_9639_4775# 1.08e-22
C1624 a_8403_4801# a_10346_4801# 9.65e-21
C1625 a_8237_4801# check[4] 8.28e-20
C1626 eob a_2289_4801# 0.0076f
C1627 comparator_out a_9638_3213# 0.00374f
C1628 x4.X a_6845_4386# 0.048f
C1629 check[3] a_12147_4801# 2.59e-19
C1630 a_7050_4086# x45.Q_N 0.00116f
C1631 D[1] a_10681_4086# 0.00123f
C1632 a_1520_2366# a_3504_2340# 9.77e-21
C1633 a_1207_2340# a_1996_2366# 4.2e-20
C1634 a_10680_2340# a_11629_2340# 1.03e-19
C1635 a_7073_4801# a_6606_4801# 0.00316f
C1636 a_10629_4801# a_10776_4086# 0.00159f
C1637 a_6466_4775# x30.Q_N 1.17e-19
C1638 a_6760_4775# a_6978_4801# 3.73e-19
C1639 check[0] a_5089_5083# 4.43e-19
C1640 check[2] check[1] 2.29f
C1641 comparator_out a_9236_2640# 0.108f
C1642 a_5561_3239# a_5562_4801# 9.85e-20
C1643 x33.Q_N a_11250_4775# 4.4e-20
C1644 a_3258_5648# a_3170_4801# 0.00133f
C1645 a_2389_5648# a_1511_4112# 0.00132f
C1646 sel_bit[1] a_3170_4801# 1.85e-19
C1647 check[2] a_9954_4112# 1.28e-19
C1648 VDD a_2389_5648# 0.696f
C1649 a_10794_3239# check[2] 0.0351f
C1650 x48.Q a_2463_4775# 9e-19
C1651 a_3599_2340# a_4112_2648# 0.00945f
C1652 a_4855_4775# check[6] 0.0103f
C1653 a_11769_4112# a_11970_4112# 3.34e-19
C1654 a_6759_3213# D[0] 4.66e-19
C1655 a_7246_3213# a_7953_3239# 0.0968f
C1656 D[3] x33.Q_N 0.00525f
C1657 check[5] a_9639_4775# 2.58e-20
C1658 check[1] a_6781_4112# 1.37e-20
C1659 comparator_out a_12345_2732# 8.26e-19
C1660 a_1338_5674# a_1227_4801# 0.00211f
C1661 x5.X a_3258_5648# 0.00256f
C1662 check[2] a_3877_5674# 8.16e-20
C1663 a_12031_4775# check[3] 0.0678f
C1664 x5.X sel_bit[1] 0.0977f
C1665 a_4926_4296# a_5170_4112# 0.00812f
C1666 check[2] a_7050_4086# 4.4e-21
C1667 x48.Q a_4453_4386# 1.14e-19
C1668 a_6466_4775# a_5992_4086# 4.54e-19
C1669 a_6011_4801# a_6305_4112# 9.06e-19
C1670 VDD a_8289_4086# 0.189f
C1671 a_1976_4775# a_2375_5167# 0.00133f
C1672 a_1415_4801# a_1592_5167# 8.94e-19
C1673 a_1508_5167# a_1822_4801# 0.0258f
C1674 a_8997_3239# a_8384_4086# 1.16e-20
C1675 a_8590_3239# x42.Q_N 8.76e-20
C1676 a_8857_3213# a_9464_3239# 0.00187f
C1677 a_8236_3239# a_8767_3605# 0.0018f
C1678 a_8402_3239# a_8590_3239# 0.163f
C1679 a_7072_3239# VDD 0.18f
C1680 a_2060_2640# x27.Q_N 0.00112f
C1681 a_8683_3605# a_9638_3213# 4.7e-22
C1682 x27.Q_N a_6199_4801# 3.25e-20
C1683 a_6605_3239# a_7181_3239# 2.46e-21
C1684 comparator_out a_11089_4112# 2.29e-20
C1685 check[1] a_4074_4775# 5.89e-20
C1686 a_8591_4801# x33.Q_N 4.33e-22
C1687 x4.X a_7264_4394# 8.47e-19
C1688 check[1] x20.Q_N 8.16e-19
C1689 a_6291_3605# x4.X 0.0177f
C1690 a_3453_4801# a_3505_4086# 6.04e-19
C1691 a_6845_4386# a_7186_4112# 0.00118f
C1692 a_6846_4086# a_6985_4112# 2.56e-19
C1693 a_6547_4086# a_8384_4086# 1.86e-21
C1694 x45.Q_N a_7764_4112# 8.17e-20
C1695 x5.A a_1415_4801# 7.6e-20
C1696 a_7072_3239# a_7318_4296# 2.37e-20
C1697 a_7246_3213# x45.Q_N 0.144f
C1698 VDD a_3619_4801# 0.617f
C1699 a_9441_2340# x42.Q_N 1.11e-19
C1700 a_10345_3239# a_10628_3239# 8.18e-19
C1701 a_5371_2366# x27.Q_N 0.0318f
C1702 a_7049_2340# a_7763_2366# 6.99e-20
C1703 VDD a_2697_5083# 0.00615f
C1704 a_6845_2340# D[4] 0.336f
C1705 a_8402_3239# a_9441_2340# 0.00154f
C1706 a_6845_2340# VDD 0.784f
C1707 a_7317_2550# a_7561_2732# 0.00972f
C1708 a_9151_3213# a_8938_2340# 2.17e-19
C1709 a_9638_3213# a_8696_2366# 8.4e-19
C1710 a_8857_3213# a_9237_2340# 0.00199f
C1711 check[6] a_7182_4801# 1.13e-20
C1712 VDD a_10795_4801# 0.593f
C1713 a_11249_3213# a_10795_4801# 3.18e-21
C1714 a_10628_3239# a_11076_5167# 8.3e-21
C1715 x77.Y a_3504_2340# 3.35e-21
C1716 a_1227_4801# a_3453_4801# 5.24e-20
C1717 a_1061_4801# a_3619_4801# 2.9e-21
C1718 a_1338_5674# check[2] 1.12e-19
C1719 a_6304_2366# x4.X 0.112f
C1720 a_1061_4801# a_2697_5083# 1.25e-19
C1721 x4.X a_1822_4801# 0.0326f
C1722 a_1227_4801# a_2194_4801# 0.00126f
C1723 eob reset 4.08e-19
C1724 a_4454_4086# x48.Q_N 1.07e-19
C1725 clk_sar a_1338_5674# 6.59e-19
C1726 a_1062_5674# x5.A 0.136f
C1727 a_4658_4086# a_4926_4296# 0.205f
C1728 a_6845_2340# a_7318_4296# 6.08e-21
C1729 a_6844_2640# x45.Q_N 4.61e-20
C1730 x5.X x39.Q_N 0.00647f
C1731 x77.Y a_4367_3213# 0.106f
C1732 a_10155_2366# VDD 0.109f
C1733 a_4214_4801# a_4586_4801# 3.34e-19
C1734 a_9151_3213# check[5] 8.29e-21
C1735 a_8696_2366# a_9236_2640# 0.139f
C1736 a_9953_2366# check[4] 5.12e-20
C1737 a_8383_2340# a_9237_2340# 0.0492f
C1738 a_9754_3239# a_9573_3239# 4.11e-20
C1739 a_12264_3521# VDD 0.00506f
C1740 reset x4.A 0.00101f
C1741 a_11856_3239# a_11942_3605# 0.00976f
C1742 a_10794_3239# x66.Q_N 3.85e-21
C1743 comparator_out D[0] 0.0253f
C1744 comparator_out x54.Q_N 0.00122f
C1745 a_11390_4801# a_11762_4801# 3.34e-19
C1746 a_8802_2366# x4.X 3.78e-20
C1747 x5.X a_6505_4394# 5.63e-19
C1748 x75.Q_N check[0] 4.68e-20
C1749 a_11389_3239# x4.X 0.00267f
C1750 x75.Q_N a_5844_3239# 2.94e-19
C1751 sel_bit[0] a_2883_5674# 0.0666f
C1752 a_1762_2340# a_1996_2732# 0.00976f
C1753 a_1520_2366# a_2198_2732# 0.00652f
C1754 x4.X a_621_4112# 9.87e-20
C1755 a_1207_2340# a_1626_2366# 0.0397f
C1756 a_9237_4386# x39.Q_N 2.03e-19
C1757 check[0] a_3913_4112# 0.00318f
C1758 a_6010_3239# a_6011_4801# 1.39e-19
C1759 a_9638_3213# a_9578_4112# 4.45e-20
C1760 a_10155_2366# a_10775_2340# 8.26e-21
C1761 a_9236_2640# a_11194_2366# 2.19e-20
C1762 check[4] a_10156_4112# 0.00259f
C1763 check[6] a_6400_4801# 1.18e-19
C1764 VDD a_9465_4801# 0.343f
C1765 comparator_out a_3600_4086# 4.69e-20
C1766 a_9464_3239# x33.Q_N 0.00295f
C1767 comparator_out a_11543_3213# 6.77e-19
C1768 a_4854_3213# a_5562_4801# 3.19e-20
C1769 a_4367_3213# check[6] 1.13e-19
C1770 check[2] a_3453_4801# 9.66e-20
C1771 x4.X a_8684_5167# 0.00132f
C1772 D[6] a_2777_2366# 1.54e-19
C1773 x5.X a_1592_5167# 4.22e-19
C1774 check[0] x4.X 0.245f
C1775 a_2200_2366# a_2401_2366# 3.34e-19
C1776 a_3504_2340# a_3912_2366# 6.04e-19
C1777 a_7363_4801# a_6845_4386# 8.84e-21
C1778 a_5844_3239# x4.X 0.0457f
C1779 check[2] a_10629_4801# 0.00307f
C1780 a_6010_3239# a_6709_3521# 2.46e-19
C1781 a_9237_2340# x33.Q_N 0.0469f
C1782 a_7481_5083# x30.Q_N 2.02e-20
C1783 comparator_out a_11330_2340# 0.00103f
C1784 a_5561_3239# a_6010_3239# 6.84e-19
C1785 a_3899_3605# a_4154_2340# 2.41e-20
C1786 check[4] check[3] 9.63e-20
C1787 a_3618_3239# a_4453_2340# 6.38e-20
C1788 a_3452_3239# a_4657_2340# 4.77e-19
C1789 a_4367_3213# a_3912_2366# 3.36e-20
C1790 a_4073_3213# a_4452_2640# 2.68e-19
C1791 check[1] a_6931_5083# 4.8e-19
C1792 x5.X a_4926_4296# 5.33e-19
C1793 x5.A x5.X 0.00793f
C1794 a_6304_2366# a_7186_4112# 1.26e-20
C1795 x48.Q a_4681_4801# 0.00128f
C1796 a_4367_3213# a_4317_3521# 1.21e-20
C1797 a_3618_3239# a_4213_3239# 0.00118f
C1798 a_7953_3239# a_9151_3213# 5.62e-20
C1799 D[0] a_8683_3605# 2.17e-19
C1800 x51.Q_N VDD 0.085f
C1801 a_6759_3213# a_7317_2550# 1.62e-19
C1802 a_7246_3213# a_7049_2340# 2.52e-19
C1803 VDD a_6710_5083# 0.00984f
C1804 D[2] check[3] 0.449f
C1805 a_3452_3239# VDD 0.821f
C1806 a_11970_4112# x39.Q_N 0.00173f
C1807 a_12346_4112# a_12102_4296# 0.00812f
C1808 a_2061_2340# x4.X 0.00458f
C1809 a_3453_4801# a_4074_4775# 0.117f
C1810 x20.Q_N a_3453_4801# 0.00252f
C1811 a_3170_4801# x27.D 0.0749f
C1812 a_10681_4086# a_11630_4086# 7e-20
C1813 a_2289_4801# a_2398_4801# 0.00707f
C1814 check[2] a_9639_4775# 0.0119f
C1815 D[0] a_8696_2366# 3.91e-20
C1816 a_6844_2640# a_7049_2340# 0.153f
C1817 a_9464_3239# a_10794_3239# 3.48e-20
C1818 a_6304_2366# x57.Q_N 0.00553f
C1819 a_4452_2640# x27.Q_N 0.569f
C1820 a_2194_4801# x20.Q_N 1.61e-19
C1821 a_8236_3239# a_10982_3239# 3.65e-21
C1822 a_9151_3213# a_11075_3605# 4.38e-20
C1823 a_9638_3213# VDD 0.569f
C1824 a_9638_3213# x69.Q_N 0.124f
C1825 a_11969_2366# check[3] 4.79e-19
C1826 a_10629_4801# a_11250_4775# 0.117f
C1827 a_9237_2340# check[1] 1.98e-19
C1828 a_3913_4112# a_4389_4478# 0.00133f
C1829 D[5] x4.X 5.17e-19
C1830 a_8857_3213# x4.X 0.00506f
C1831 x72.Q_N x4.X 0.00455f
C1832 VDD a_4872_4394# 0.0102f
C1833 x5.X x27.D 0.151f
C1834 a_4214_4801# a_3600_4086# 1.08e-19
C1835 a_8858_4775# a_8384_4086# 4.54e-19
C1836 D[4] a_9236_2640# 3.87e-20
C1837 a_8403_4801# a_8697_4112# 9.06e-19
C1838 a_7763_2366# a_9237_2340# 3.65e-21
C1839 a_7953_3239# check[5] 0.0271f
C1840 a_9236_2640# VDD 0.269f
C1841 check[0] a_7186_4112# 3.6e-20
C1842 VDD a_4586_4801# 0.00495f
C1843 D[1] a_11389_3239# 1.6e-19
C1844 a_3258_5648# a_3373_5674# 0.18f
C1845 sel_bit[1] a_3373_5674# 0.0439f
C1846 a_2883_5674# a_2788_5674# 0.00133f
C1847 check[3] a_11834_4086# 8.07e-19
C1848 a_11543_3213# a_11390_4801# 1.61e-20
C1849 a_10628_3239# x36.Q_N 2.75e-19
C1850 VDD a_11762_4801# 0.00445f
C1851 x4.X a_4389_4478# 2.12e-19
C1852 a_5372_4112# a_6846_4086# 3.65e-21
C1853 a_5897_4086# a_6845_4386# 9.02e-21
C1854 a_8383_2340# x4.X 0.111f
C1855 x5.X a_6760_4775# 0.00141f
C1856 x27.Q_N a_6846_4086# 1.92e-21
C1857 a_12345_2732# VDD 0.0042f
C1858 a_6011_4801# a_7073_4801# 0.137f
C1859 a_6292_5167# a_6760_4775# 0.0633f
C1860 a_9441_2340# a_9376_2366# 9.75e-19
C1861 a_5845_4801# a_6199_4801# 0.0663f
C1862 a_9236_2640# a_10775_2340# 3.6e-19
C1863 a_9237_2340# a_9577_2366# 6.04e-20
C1864 check[0] a_4368_4775# 0.00265f
C1865 x57.Q_N check[0] 0.0113f
C1866 comparator_out a_10345_3239# 0.00106f
C1867 x77.Y a_4454_4086# 2.63e-20
C1868 a_8237_4801# a_10983_4801# 3.65e-21
C1869 a_9465_4801# a_10795_4801# 2.57e-20
C1870 comparator_out a_7317_2550# 0.00825f
C1871 a_11766_2732# x4.X 9.81e-19
C1872 x5.X a_9238_4086# 0.261f
C1873 a_9151_3213# check[2] 2.41e-20
C1874 D[6] a_3504_2340# 0.103f
C1875 a_2060_2640# a_2777_2366# 0.0019f
C1876 check[5] x45.Q_N 5.14e-20
C1877 a_10776_4086# a_11565_4478# 7.71e-20
C1878 a_11089_4112# a_11289_4394# 0.00185f
C1879 VDD a_11089_4112# 0.448f
C1880 a_11249_3213# a_11089_4112# 0.00148f
C1881 a_10794_3239# a_11331_4086# 1.07e-20
C1882 a_10628_3239# a_11629_4386# 6.5e-20
C1883 a_11088_2366# a_12047_2648# 1.21e-20
C1884 a_11330_2340# a_11194_2366# 0.0282f
C1885 a_11628_2640# a_11766_2732# 1.09e-19
C1886 eob a_3258_5648# 3.1e-19
C1887 eob sel_bit[1] 0.317f
C1888 comparator_out D[7] 6.69e-20
C1889 a_4367_3213# a_6465_3213# 4.53e-20
C1890 a_4854_3213# a_6010_3239# 3.57e-19
C1891 sel_bit[1] x4.A 1.56e-20
C1892 x4.X a_9377_4112# 6.75e-19
C1893 a_8384_4086# x42.Q_N 0.154f
C1894 a_8697_4112# a_9710_4296# 0.0633f
C1895 a_9237_4386# a_9238_4086# 0.75f
C1896 check[6] a_4454_4086# 0.0339f
C1897 a_8939_4086# a_9442_4086# 0.00187f
C1898 a_8402_3239# a_8384_4086# 3.48e-19
C1899 x4.X x33.Q_N 0.421f
C1900 a_8236_3239# a_8697_4112# 2.21e-19
C1901 a_4855_4775# a_6199_4801# 8.26e-21
C1902 clk_sar x3.A 1.29e-20
C1903 a_10775_2340# a_11089_4112# 5.05e-21
C1904 a_7246_3213# a_9464_3239# 1.86e-21
C1905 a_2533_2550# x20.Q_N 0.153f
C1906 a_6759_3213# a_8590_3239# 3.42e-20
C1907 x5.X a_9755_4801# 2.07e-19
C1908 check[3] a_12548_4112# 0.159f
C1909 a_8403_4801# a_9102_5083# 2.46e-19
C1910 a_11628_2640# x33.Q_N 1.12e-20
C1911 a_8237_4801# a_9323_5083# 0.00907f
C1912 a_3618_3239# a_3453_4801# 8.16e-19
C1913 a_3452_3239# a_3619_4801# 9.04e-19
C1914 a_2853_5648# a_1976_4775# 1.02e-19
C1915 a_4854_3213# a_4793_2366# 1.2e-20
C1916 x48.Q a_3648_5972# 0.00114f
C1917 a_5992_4086# a_6505_4394# 0.00945f
C1918 a_4453_2340# a_3913_4112# 1.4e-21
C1919 a_4452_2640# a_4155_4086# 4.75e-21
C1920 check[2] check[5] 7.25e-20
C1921 D[0] D[4] 0.338f
C1922 D[5] x57.Q_N 0.00107f
C1923 D[0] VDD 0.301f
C1924 a_8857_3213# D[1] 1.23e-20
C1925 D[7] a_2265_2340# 2.67e-19
C1926 a_6759_3213# x27.Q_N 8.29e-21
C1927 a_7561_2366# x30.Q_N 0.00224f
C1928 x54.Q_N VDD 0.0807f
C1929 a_9755_4801# a_9237_4386# 8.84e-21
C1930 check[1] a_3913_4112# 9.87e-21
C1931 a_12101_2550# check[3] 9.97e-19
C1932 sel_bit[0] reset 8.49e-21
C1933 a_5088_3521# VDD 0.00529f
C1934 a_4074_4775# a_4019_4112# 8.14e-21
C1935 a_4453_2340# x4.X 0.00242f
C1936 x5.X a_9954_4478# 1.64e-19
C1937 check[2] a_10776_4086# 0.0128f
C1938 a_7953_3239# x45.Q_N 3.23e-19
C1939 VDD a_3600_4086# 0.741f
C1940 a_4368_4775# a_4767_5167# 0.00133f
C1941 a_3900_5167# a_4214_4801# 0.0258f
C1942 a_3453_4801# a_5089_5083# 1.25e-19
C1943 a_3619_4801# a_4586_4801# 0.00126f
C1944 a_10794_3239# a_11195_4112# 4.04e-21
C1945 VDD a_11767_4478# 0.0163f
C1946 a_9638_3213# a_10155_2366# 2.38e-19
C1947 a_6546_2340# x27.Q_N 5.08e-20
C1948 a_10628_3239# a_11856_3239# 0.0334f
C1949 a_6844_2640# a_9237_2340# 2.9e-21
C1950 x5.X a_8998_4801# 9.4e-19
C1951 a_7317_2550# a_8696_2366# 6.06e-21
C1952 a_10794_3239# a_12030_3213# 0.0264f
C1953 a_6845_2340# a_9236_2640# 4e-20
C1954 x20.Q_N a_4008_4801# 9.98e-20
C1955 a_11249_3213# a_11543_3213# 0.199f
C1956 a_11543_3213# VDD 0.352f
C1957 check[1] x4.X 0.262f
C1958 x69.Q_N a_11543_3213# 2.97e-20
C1959 a_4213_3239# x4.X 0.00268f
C1960 a_7481_5083# a_8237_4801# 4.06e-20
C1961 a_1682_4775# a_1511_4112# 0.00416f
C1962 a_10629_4801# a_12265_5083# 1.25e-19
C1963 a_10795_4801# a_11762_4801# 0.00126f
C1964 a_11076_5167# a_11390_4801# 0.0258f
C1965 a_11544_4775# a_11943_5167# 0.00133f
C1966 a_7763_2366# x4.X 8.68e-20
C1967 x4.X a_9954_4112# 6.39e-19
C1968 VDD a_1682_4775# 0.337f
C1969 a_10794_3239# x4.X 0.0425f
C1970 a_4454_4086# a_6547_4086# 1.67e-21
C1971 a_4926_4296# a_5992_4086# 7.98e-21
C1972 a_4073_3213# comparator_out 3.96e-19
C1973 a_9872_3521# x4.X 0.00103f
C1974 a_9237_4386# a_9954_4478# 4.45e-20
C1975 x5.X a_5562_4801# 0.0294f
C1976 a_8384_4086# a_9173_4112# 4.2e-20
C1977 a_9238_4086# a_9656_4394# 0.00276f
C1978 x77.Y x75.Q 3.59e-19
C1979 a_9237_2340# a_9953_2732# 0.0018f
C1980 a_9441_2340# a_9655_2648# 0.0104f
C1981 check[6] a_6466_4775# 6.88e-19
C1982 a_9236_2640# a_10155_2366# 0.159f
C1983 a_11543_3213# a_10775_2340# 9.06e-19
C1984 a_11330_2340# VDD 0.177f
C1985 a_11249_3213# a_11330_2340# 4.18e-20
C1986 a_10628_3239# a_11629_2340# 6.52e-20
C1987 a_11075_3605# a_11088_2366# 1.71e-19
C1988 a_10794_3239# a_11628_2640# 4.04e-20
C1989 a_7049_2340# check[5] 7.15e-20
C1990 x5.X a_12738_4801# 0.0161f
C1991 sel_bit[0] a_3807_4801# 7.41e-20
C1992 a_9638_3213# a_9465_4801# 4.82e-21
C1993 a_9464_3239# a_9639_4775# 1.33e-23
C1994 a_1061_4801# a_1682_4775# 0.113f
C1995 a_8858_4775# check[4] 9.03e-21
C1996 a_3877_5674# x4.X 4.83e-20
C1997 eob a_1592_5167# 5.68e-19
C1998 comparator_out a_8590_3239# 0.158f
C1999 a_11183_3239# x36.Q_N 6.74e-20
C2000 x4.X a_7050_4086# 0.00987f
C2001 a_1338_5674# a_1508_5167# 5.69e-20
C2002 a_1762_2340# a_1996_2366# 0.00707f
C2003 check[0] a_5897_4086# 0.116f
C2004 a_1520_2366# a_2200_2366# 3.73e-19
C2005 a_2060_2640# a_3504_2340# 6.83e-19
C2006 a_10775_2340# a_11330_2340# 0.197f
C2007 comparator_out a_5372_4112# 4.39e-20
C2008 a_5844_3239# a_5897_4086# 5.06e-19
C2009 a_6199_4801# a_6400_4801# 3.67e-19
C2010 a_10795_4801# a_11089_4112# 9.06e-19
C2011 a_6760_4775# x30.Q_N 0.00766f
C2012 a_7247_4775# a_7481_5083# 0.00945f
C2013 a_7073_4801# a_6978_4801# 0.00276f
C2014 a_11250_4775# a_10776_4086# 4.54e-19
C2015 D[1] x33.Q_N 3.29e-19
C2016 x5.A eob 0.0017f
C2017 comparator_out x27.Q_N 0.272f
C2018 comparator_out a_9441_2340# 0.00598f
C2019 x75.Q check[6] 0.0149f
C2020 x33.Q_N a_11544_4775# 1.35e-20
C2021 a_3373_5674# x27.D 5.58e-20
C2022 comparator_out x36.Q_N 0.267f
C2023 x5.A x4.A 5.23e-21
C2024 D[0] a_8289_4086# 0.00123f
C2025 a_11075_3605# check[2] 8.1e-20
C2026 a_3912_2366# a_4388_2732# 0.00133f
C2027 a_7072_3239# D[0] 5.18e-20
C2028 x30.Q_N a_9238_4086# 1.91e-21
C2029 a_11493_3521# x39.Q_N 0.00136f
C2030 a_6605_3239# x30.Q_N 6.1e-19
C2031 check[5] a_8591_4801# 0.165f
C2032 check[1] a_7186_4112# 2.11e-19
C2033 a_10983_4801# check[3] 1.14e-19
C2034 check[2] x45.Q_N 2.88e-21
C2035 x5.X a_6305_4112# 0.00598f
C2036 x48.Q a_4658_4086# 3.93e-19
C2037 a_5845_4801# a_6846_4086# 1.15e-19
C2038 a_6011_4801# a_6845_4386# 7.24e-20
C2039 a_6466_4775# a_6547_4086# 8.83e-20
C2040 a_6760_4775# a_5992_4086# 0.0018f
C2041 a_6292_5167# a_6305_4112# 2.81e-19
C2042 a_11088_2366# check[2] 0.00327f
C2043 VDD a_6985_4112# 0.00445f
C2044 a_2289_4801# a_2375_5167# 0.00976f
C2045 D[0] a_6845_2340# 0.0271f
C2046 a_4453_2340# x57.Q_N 2.94e-19
C2047 a_8402_3239# a_7362_3239# 1.22e-20
C2048 a_8683_3605# a_8590_3239# 0.0367f
C2049 a_6375_3605# VDD 0.0042f
C2050 a_8857_3213# a_8767_3605# 6.69e-20
C2051 a_9151_3213# a_9464_3239# 0.124f
C2052 a_8288_2340# x30.Q_N 2.02e-19
C2053 check[4] x42.Q_N 6.27e-20
C2054 x27.Q_N a_4971_4801# 0.00139f
C2055 a_3618_3239# a_4019_4112# 4.04e-21
C2056 a_8402_3239# check[4] 1.83e-21
C2057 comparator_out a_11629_4386# 2.51e-20
C2058 check[1] a_4368_4775# 1.09e-19
C2059 eob x27.D 4.69e-19
C2060 x4.X a_7764_4112# 0.00621f
C2061 a_7246_3213# x4.X 0.115f
C2062 a_6845_4386# a_8697_4112# 1.34e-19
C2063 a_3619_4801# a_3600_4086# 6.63e-19
C2064 a_7050_4086# a_7186_4112# 0.07f
C2065 x45.Q_N a_6781_4112# 0.00138f
C2066 a_6846_4086# a_8384_4086# 2.98e-19
C2067 a_3453_4801# a_3913_4112# 3.05e-19
C2068 x20.Q_N a_3505_4086# 0.00428f
C2069 a_6605_3239# a_5992_4086# 1.16e-20
C2070 a_6198_3239# x45.Q_N 7.37e-20
C2071 VDD a_3900_5167# 0.324f
C2072 a_10345_3239# VDD 0.19f
C2073 D[1] a_10794_3239# 0.00642f
C2074 a_9151_3213# a_9237_2340# 2.19e-19
C2075 a_9638_3213# a_9236_2640# 3.43e-19
C2076 a_7317_2550# VDD 0.172f
C2077 x69.Q_N a_10345_3239# 0.178f
C2078 a_11075_3605# a_11250_4775# 1.33e-23
C2079 a_11249_3213# a_11076_5167# 3.52e-21
C2080 VDD a_11076_5167# 0.317f
C2081 a_11543_3213# a_10795_4801# 2.05e-21
C2082 a_1207_2340# eob 1.75e-19
C2083 x4.X a_3453_4801# 0.00472f
C2084 x4.X a_2194_4801# 0.00509f
C2085 a_1227_4801# x20.Q_N 1.52e-19
C2086 a_6844_2640# x4.X 0.00904f
C2087 x4.X a_10629_4801# 0.00428f
C2088 a_1207_2340# x4.A 9.28e-20
C2089 a_7049_2340# x45.Q_N 1.11e-19
C2090 x48.Q a_3170_4801# 0.00244f
C2091 x77.Y a_4680_3239# 0.16f
C2092 a_12030_3213# a_12146_3239# 0.0397f
C2093 a_8938_2340# a_9237_2340# 0.0334f
C2094 a_8383_2340# a_9709_2550# 4.7e-22
C2095 a_8696_2366# a_9441_2340# 0.199f
C2096 D[7] VDD 0.225f
C2097 a_11543_3213# a_11965_3239# 2.87e-21
C2098 a_4214_4801# x27.Q_N 1.45e-19
C2099 a_11543_3213# a_12264_3521# 0.00185f
C2100 check[1] a_8897_4394# 9.73e-20
C2101 a_11390_4801# x36.Q_N 4.02e-20
C2102 a_9953_2732# x4.X 1.17e-19
C2103 a_12146_3239# x4.X 5.65e-19
C2104 x5.X a_6983_4478# 7.44e-19
C2105 x5.X x48.Q 0.203f
C2106 a_11761_3239# x4.X 4.96e-19
C2107 sel_bit[0] a_3258_5648# 0.0205f
C2108 a_6466_4775# a_6411_4112# 8.14e-21
C2109 a_1762_2340# a_1626_2366# 0.0282f
C2110 a_2060_2640# a_2198_2732# 1.09e-19
C2111 sel_bit[0] sel_bit[1] 0.428f
C2112 a_1520_2366# a_2479_2648# 1.21e-20
C2113 a_1926_5083# x27.D 3.95e-22
C2114 a_9442_4086# x39.Q_N 3.43e-20
C2115 check[0] a_4453_4386# 0.164f
C2116 a_6465_3213# a_6466_4775# 2.59e-19
C2117 a_6010_3239# a_6292_5167# 1.65e-21
C2118 D[3] a_11088_2366# 8.67e-19
C2119 a_6291_3605# a_6011_4801# 8.52e-21
C2120 a_12146_3239# a_11628_2640# 5.05e-21
C2121 a_9237_2340# check[5] 7.28e-22
C2122 VDD a_8768_5167# 0.0042f
C2123 x77.Y a_4794_4112# 7.13e-20
C2124 a_11194_2366# x36.Q_N 0.0102f
C2125 comparator_out a_11856_3239# 1.89e-19
C2126 x33.Q_N a_10346_4801# 0.184f
C2127 check[2] a_4074_4775# 1.07e-19
C2128 a_7318_4296# a_7562_4112# 0.00812f
C2129 x4.X a_9639_4775# 0.103f
C2130 x27.D x48.Q_N 8.11e-20
C2131 x5.X a_2147_5083# 4.05e-19
C2132 check[2] x20.Q_N 4.28e-20
C2133 a_7246_3213# a_7186_4112# 4.45e-20
C2134 a_11194_2366# a_11564_2366# 4.11e-20
C2135 a_3504_2340# a_4452_2640# 9.65e-21
C2136 a_7363_4801# a_7050_4086# 7.76e-20
C2137 a_6010_3239# a_7158_3605# 2.13e-19
C2138 a_6465_3213# a_6930_3521# 9.46e-19
C2139 a_9709_2550# x33.Q_N 0.181f
C2140 comparator_out a_11629_2340# 0.183f
C2141 a_4680_3239# a_3912_2366# 2.17e-19
C2142 a_4367_3213# a_4452_2640# 5.32e-19
C2143 a_3806_3239# a_3599_2340# 2.02e-19
C2144 D[3] check[2] 0.194f
C2145 x48.Q a_3984_5167# 5.76e-19
C2146 a_4367_3213# a_4766_3605# 0.00133f
C2147 a_3806_3239# a_3983_3605# 8.94e-19
C2148 a_3452_3239# a_5088_3521# 1.25e-19
C2149 a_3618_3239# a_4585_3239# 0.00126f
C2150 a_3899_3605# a_4213_3239# 0.0258f
C2151 D[0] a_9638_3213# 1.68e-20
C2152 a_7072_3239# a_7317_2550# 1.85e-20
C2153 VDD a_7159_5167# 0.00371f
C2154 a_3452_3239# a_3600_4086# 8.29e-19
C2155 a_11768_2366# x33.Q_N 2.75e-20
C2156 a_4073_3213# VDD 0.314f
C2157 a_2533_2550# x4.X 5.96e-19
C2158 x4.X a_4790_4801# 2.39e-19
C2159 a_3912_2366# a_4794_4112# 1.26e-20
C2160 a_3453_4801# a_4368_4775# 0.125f
C2161 a_3619_4801# a_3900_5167# 0.155f
C2162 a_10776_4086# a_11331_4086# 0.197f
C2163 x30.Q_N a_6305_4112# 1.32e-21
C2164 a_10156_4112# x39.Q_N 8.08e-20
C2165 x5.X a_8403_4801# 0.0201f
C2166 x20.Q_N a_4074_4775# 8.63e-20
C2167 a_9638_3213# a_11543_3213# 3.71e-20
C2168 a_6844_2640# x57.Q_N 4.82e-21
C2169 a_6845_2340# a_7317_2550# 0.15f
C2170 a_8590_3239# VDD 0.109f
C2171 a_2853_5648# a_2883_5674# 0.224f
C2172 a_4657_2340# x27.Q_N 0.179f
C2173 a_6760_4775# a_8237_4801# 1.67e-19
C2174 D[1] a_10629_4801# 1.99e-20
C2175 a_10628_3239# check[4] 0.00655f
C2176 check[0] a_6011_4801# 4.88e-19
C2177 check[1] a_5897_4086# 1.24e-21
C2178 x33.Q_N a_11630_4086# 1.91e-21
C2179 a_5844_3239# a_6011_4801# 9.04e-19
C2180 a_10629_4801# a_11544_4775# 0.125f
C2181 a_10795_4801# a_11076_5167# 0.155f
C2182 a_9709_2550# check[1] 2.04e-19
C2183 a_4454_4086# a_4113_4394# 1.25e-19
C2184 a_4007_3239# x27.Q_N 6.74e-20
C2185 a_4155_4086# a_4591_4478# 0.00412f
C2186 a_3913_4112# a_4019_4112# 0.0552f
C2187 a_4453_4386# a_4389_4478# 2.13e-19
C2188 a_9151_3213# x4.X 0.111f
C2189 VDD a_5372_4112# 0.11f
C2190 a_8858_4775# a_8939_4086# 8.83e-20
C2191 a_8684_5167# a_8697_4112# 2.81e-19
C2192 a_8237_4801# a_9238_4086# 1.15e-19
C2193 VDD x27.Q_N 0.452f
C2194 D[1] a_12146_3239# 1.57e-20
C2195 a_10628_3239# D[2] 6.24e-20
C2196 D[4] a_9441_2340# 6.5e-20
C2197 a_9152_4775# a_8384_4086# 0.0018f
C2198 a_10794_3239# a_12737_3239# 6.86e-21
C2199 a_8403_4801# a_9237_4386# 7.24e-20
C2200 a_9441_2340# VDD 0.304f
C2201 a_1112_2340# x20.Q_N 4.68e-19
C2202 a_3373_5674# a_3876_6040# 0.00336f
C2203 D[1] a_11761_3239# 5.48e-20
C2204 a_9376_2366# check[4] 9.3e-20
C2205 comparator_out a_8384_4086# 0.00194f
C2206 sel_bit[1] a_2788_5674# 2.36e-19
C2207 check[3] x39.Q_N 1.04e-19
C2208 a_11249_3213# x36.Q_N 5.36e-19
C2209 VDD x36.Q_N 0.419f
C2210 x4.X a_4019_4112# 0.00642f
C2211 a_5844_3239# a_6709_3521# 0.00276f
C2212 a_5561_3239# check[0] 0.0043f
C2213 a_5992_4086# a_6305_4112# 0.272f
C2214 x4.X a_4008_4801# 8.46e-20
C2215 a_8938_2340# x4.X 0.00706f
C2216 a_5561_3239# a_5844_3239# 8.18e-19
C2217 x4.X x3.A 2.12e-20
C2218 x5.X a_7073_4801# 0.00115f
C2219 a_1207_2340# a_1520_2366# 0.273f
C2220 x4.X a_11184_4801# 8.46e-20
C2221 x5.A sel_bit[0] 0.0448f
C2222 a_9236_2640# a_11330_2340# 4.16e-20
C2223 a_6466_4775# a_6199_4801# 6.99e-20
C2224 a_9237_2340# a_11088_2366# 3.08e-19
C2225 a_9709_2550# a_9577_2366# 0.0258f
C2226 a_6760_4775# a_7247_4775# 0.273f
C2227 a_6011_4801# a_6376_5167# 4.45e-20
C2228 check[0] a_4681_4801# 0.00122f
C2229 a_10775_2340# x36.Q_N 0.142f
C2230 x77.Y a_4926_4296# 0.00166f
C2231 a_12047_2648# x4.X 2.86e-19
C2232 x4.X check[5] 0.0317f
C2233 x5.X a_9710_4296# 6.08e-19
C2234 a_8236_3239# x5.X 9.93e-20
C2235 D[6] a_2200_2366# 1.47e-19
C2236 a_2061_2340# a_4112_2648# 4.06e-20
C2237 a_10776_4086# a_11195_4112# 0.0397f
C2238 a_11089_4112# a_11767_4478# 0.00652f
C2239 a_4388_2366# check[6] 2.11e-20
C2240 a_11331_4086# a_11565_4478# 0.00976f
C2241 a_11088_2366# a_12547_2366# 4.94e-21
C2242 a_11628_2640# a_12047_2648# 2.46e-19
C2243 x63.Q_N a_11288_2648# 2.02e-20
C2244 a_11075_3605# a_11331_4086# 1.7e-20
C2245 a_10775_2340# a_11564_2366# 4.2e-20
C2246 a_10628_3239# a_11834_4086# 0.00195f
C2247 a_10794_3239# a_11630_4086# 6.04e-20
C2248 a_11543_3213# a_11089_4112# 3.33e-20
C2249 a_11249_3213# a_11629_4386# 0.0015f
C2250 VDD a_11629_4386# 0.59f
C2251 a_11833_2340# a_11766_2732# 9.46e-19
C2252 a_6010_3239# x30.Q_N 4.02e-19
C2253 a_4367_3213# a_6759_3213# 3.6e-20
C2254 a_4854_3213# a_6291_3605# 7.98e-21
C2255 x4.X a_10776_4086# 0.1f
C2256 a_8939_4086# x42.Q_N 0.0287f
C2257 a_9238_4086# a_9442_4086# 0.117f
C2258 a_9237_4386# a_9710_4296# 0.155f
C2259 a_9237_2340# check[2] 6.22e-19
C2260 a_8857_3213# a_8697_4112# 0.00148f
C2261 a_1720_2648# VDD 0.00736f
C2262 a_8402_3239# a_8939_4086# 1.07e-20
C2263 a_8236_3239# a_9237_4386# 6.5e-20
C2264 a_3912_2366# a_4388_2366# 2.87e-21
C2265 a_8858_4775# a_8803_4112# 8.14e-21
C2266 a_4368_4775# a_4790_4801# 2.87e-21
C2267 a_4855_4775# a_4971_4801# 0.0397f
C2268 a_6759_3213# a_7362_3239# 0.0552f
C2269 x5.X a_11494_5083# 3.98e-19
C2270 sel_bit[0] x27.D 0.00108f
C2271 a_621_4112# a_897_4112# 0.00202f
C2272 a_8858_4775# a_9323_5083# 9.46e-19
C2273 a_8403_4801# a_9551_5167# 2.13e-19
C2274 a_8237_4801# a_8998_4801# 6.04e-20
C2275 a_11833_2340# x33.Q_N 8.49e-21
C2276 a_3452_3239# a_3900_5167# 8.3e-21
C2277 check[1] a_2463_4775# 0.00193f
C2278 a_5561_3239# D[5] 0.00127f
C2279 a_4073_3213# a_3619_4801# 3.18e-21
C2280 a_3618_3239# x20.Q_N 0.0017f
C2281 x48.Q a_3373_5674# 0.0679f
C2282 a_6305_4112# a_6781_4478# 0.00133f
C2283 a_1976_4775# a_1511_4112# 0.00824f
C2284 a_6010_3239# a_5992_4086# 3.48e-19
C2285 x54.Q_N a_3600_4086# 2.32e-20
C2286 a_4453_2340# a_4453_4386# 7.25e-19
C2287 a_3599_2340# x48.Q_N 9.38e-21
C2288 a_4452_2640# a_4454_4086# 7.02e-19
C2289 a_5991_2340# a_6504_2648# 0.00945f
C2290 a_8383_2340# a_8697_4112# 5.05e-21
C2291 VDD a_1976_4775# 0.489f
C2292 a_9151_3213# D[1] 4.66e-19
C2293 a_9638_3213# a_10345_3239# 0.0968f
C2294 D[7] x51.Q_N 0.00276f
C2295 a_5845_4801# a_7954_4801# 1.03e-19
C2296 a_9755_4801# a_9442_4086# 7.76e-20
C2297 check[1] a_4453_4386# 1.28e-20
C2298 a_10346_4801# a_10629_4801# 8.18e-19
C2299 a_1227_4801# a_1508_5167# 0.151f
C2300 a_1061_4801# a_1976_4775# 0.117f
C2301 a_7953_3239# x4.X 0.00272f
C2302 a_3505_4086# a_3913_4112# 6.04e-19
C2303 a_4925_2550# x4.X 0.00127f
C2304 VDD a_4155_4086# 0.348f
C2305 x5.X a_10681_4086# 0.0752f
C2306 check[2] a_11331_4086# 3.82e-19
C2307 a_2579_4801# a_2398_4801# 4.11e-20
C2308 a_4681_4801# a_4767_5167# 0.00976f
C2309 a_3619_4801# x27.Q_N 1.18e-19
C2310 a_11075_3605# a_11195_4112# 1.12e-20
C2311 VDD a_12048_4394# 0.00984f
C2312 x5.X a_9370_4801# 2.59e-19
C2313 a_10628_3239# a_11159_3605# 0.0018f
C2314 a_11249_3213# a_11856_3239# 0.00187f
C2315 a_10794_3239# a_10982_3239# 0.163f
C2316 a_11856_3239# VDD 0.18f
C2317 a_6845_2340# x27.Q_N 6.49e-21
C2318 a_11075_3605# a_12030_3213# 4.7e-22
C2319 a_8997_3239# a_9573_3239# 2.46e-21
C2320 a_4585_3239# x4.X 5e-19
C2321 x30.Q_N a_8403_4801# 2.26e-19
C2322 comparator_out a_3504_2340# 0.00285f
C2323 eob x48.Q 0.0102f
C2324 x77.Y a_4018_2366# 6.03e-20
C2325 x75.Q_N x45.Q_N 6.77e-21
C2326 x4.X a_3505_4086# 0.0122f
C2327 a_10795_4801# x36.Q_N 2.98e-20
C2328 a_11857_4801# a_11943_5167# 0.00976f
C2329 a_9755_4801# a_9574_4801# 4.11e-20
C2330 x4.X a_11565_4478# 2.12e-19
C2331 a_4854_3213# check[0] 0.00313f
C2332 a_4454_4086# a_6846_4086# 1.37e-19
C2333 a_3913_4112# x45.Q_N 1.22e-20
C2334 a_11075_3605# x4.X 0.0178f
C2335 x48.Q x4.A 1.09e-20
C2336 a_4367_3213# comparator_out 5.5e-19
C2337 a_4854_3213# a_5844_3239# 0.00116f
C2338 a_9238_4086# a_10156_4112# 0.0663f
C2339 a_9442_4086# a_9954_4478# 6.69e-20
C2340 a_8697_4112# a_9377_4112# 3.73e-19
C2341 x42.Q_N a_8803_4112# 0.0446f
C2342 a_8939_4086# a_9173_4112# 0.00707f
C2343 a_9237_4386# a_10681_4086# 3.59e-19
C2344 a_8402_3239# a_8803_4112# 4.04e-21
C2345 check[6] a_6760_4775# 0.00308f
C2346 a_9237_2340# D[3] 0.336f
C2347 a_9441_2340# a_10155_2366# 6.99e-20
C2348 a_9709_2550# a_9953_2732# 0.00972f
C2349 a_11088_2366# a_11195_4112# 8.38e-21
C2350 a_11543_3213# a_11330_2340# 2.17e-19
C2351 a_11249_3213# a_11629_2340# 0.00199f
C2352 a_11629_2340# VDD 0.784f
C2353 a_10794_3239# a_11833_2340# 0.00154f
C2354 a_12030_3213# a_11088_2366# 8.4e-19
C2355 x33.Q_N a_8697_4112# 7.32e-22
C2356 a_1227_4801# x4.X 0.311f
C2357 a_10155_2366# x36.Q_N 1.34e-20
C2358 a_9152_4775# check[4] 0.00456f
C2359 a_9639_4775# a_10346_4801# 0.0968f
C2360 eob a_2147_5083# 0.00298f
C2361 a_11965_3239# x36.Q_N 1.68e-19
C2362 x4.X x45.Q_N 0.252f
C2363 comparator_out check[4] 0.0222f
C2364 a_2389_5648# a_1976_4775# 1.09e-19
C2365 a_11088_2366# x4.X 0.112f
C2366 a_2777_2732# a_2979_2366# 8.94e-19
C2367 check[0] a_4593_4112# 5.07e-20
C2368 a_4018_2366# check[6] 1.17e-19
C2369 a_1762_2340# a_2401_2366# 0.00316f
C2370 a_1520_2366# a_3599_2340# 8.34e-21
C2371 a_2060_2640# a_2200_2366# 0.00126f
C2372 a_10775_2340# a_11629_2340# 0.0492f
C2373 a_11088_2366# a_11628_2640# 0.139f
C2374 a_7073_4801# x30.Q_N 4.49e-19
C2375 a_11076_5167# a_11089_4112# 2.81e-19
C2376 a_11250_4775# a_11331_4086# 8.83e-20
C2377 a_10795_4801# a_11629_4386# 7.24e-20
C2378 a_11544_4775# a_10776_4086# 0.0018f
C2379 a_10629_4801# a_11630_4086# 1.15e-19
C2380 comparator_out D[2] 0.0211f
C2381 check[1] a_6011_4801# 4e-19
C2382 comparator_out x60.Q_N 3.61e-19
C2383 x33.Q_N a_11857_4801# 1.75e-20
C2384 a_8998_4801# a_9574_4801# 2.46e-21
C2385 a_4367_3213# a_4971_4801# 1.05e-20
C2386 check[2] a_3913_4112# 1.35e-20
C2387 check[2] a_11195_4112# 4.22e-19
C2388 a_3452_3239# a_4073_3213# 0.115f
C2389 a_4154_2340# a_4590_2732# 0.00412f
C2390 a_4452_2640# a_4388_2732# 2.13e-19
C2391 a_3912_2366# a_4018_2366# 0.0552f
C2392 a_4453_2340# a_4112_2648# 1.25e-19
C2393 D[6] a_4388_2366# 1.34e-19
C2394 VDD a_5845_4801# 0.81f
C2395 a_4970_3239# a_4925_2550# 1.01e-20
C2396 a_11942_3605# x39.Q_N 3.64e-19
C2397 a_8236_3239# x30.Q_N 8.92e-20
C2398 check[5] a_7363_4801# 8.69e-20
C2399 VDD a_12147_4801# 0.0101f
C2400 a_6977_3239# x30.Q_N 4.04e-19
C2401 check[1] a_8697_4112# 0.00119f
C2402 check[2] x4.X 0.258f
C2403 a_5561_3239# a_4453_2340# 4.83e-19
C2404 x5.X a_6845_4386# 0.0101f
C2405 x48.Q x48.Q_N 0.00314f
C2406 a_2463_4775# a_3453_4801# 0.00116f
C2407 a_1976_4775# a_3619_4801# 2.05e-19
C2408 a_6760_4775# a_6547_4086# 3.72e-19
C2409 a_11628_2640# check[2] 3.14e-19
C2410 a_7247_4775# a_6305_4112# 0.00161f
C2411 a_9954_4478# a_10156_4112# 8.94e-19
C2412 a_6011_4801# a_7050_4086# 0.00221f
C2413 a_8803_4112# a_9173_4112# 4.11e-20
C2414 VDD a_8384_4086# 0.716f
C2415 a_6466_4775# a_6846_4086# 0.00336f
C2416 a_1976_4775# a_2697_5083# 0.00185f
C2417 a_2777_2366# VDD 8.32e-19
C2418 a_1508_5167# x20.Q_N 9.58e-20
C2419 a_5896_2340# a_6304_2366# 6.04e-19
C2420 a_4592_2366# a_4793_2366# 3.34e-19
C2421 a_9101_3521# x42.Q_N 0.00136f
C2422 a_8236_3239# a_9322_3521# 0.00907f
C2423 a_8402_3239# a_9101_3521# 2.46e-19
C2424 a_4789_3239# VDD 1.15e-19
C2425 a_6984_2366# x30.Q_N 0.00473f
C2426 a_3899_3605# a_4019_4112# 1.12e-20
C2427 comparator_out a_11834_4086# 4.39e-21
C2428 check[1] a_4681_4801# 3.58e-20
C2429 a_2853_5648# a_3807_4801# 1.57e-19
C2430 x4.X a_6781_4112# 8.67e-20
C2431 a_3452_3239# x27.Q_N 2.63e-19
C2432 a_4367_3213# a_4214_4801# 1.61e-20
C2433 a_6198_3239# x4.X 0.00604f
C2434 a_3453_4801# a_4453_4386# 9.86e-20
C2435 a_3900_5167# a_3600_4086# 4.9e-20
C2436 a_4074_4775# a_3913_4112# 0.0025f
C2437 a_7318_4296# a_8384_4086# 7.98e-21
C2438 x45.Q_N a_7186_4112# 0.00171f
C2439 a_6846_4086# a_8939_4086# 1.67e-21
C2440 x20.Q_N a_3913_4112# 7.65e-19
C2441 a_4970_3239# x45.Q_N 9.58e-21
C2442 VDD a_4855_4775# 0.723f
C2443 check[0] a_5170_4112# 8.39e-20
C2444 D[1] a_11075_3605# 2.08e-19
C2445 a_10345_3239# a_11543_3213# 5.62e-20
C2446 a_9151_3213# a_9709_2550# 1.62e-19
C2447 a_9638_3213# a_9441_2340# 2.52e-19
C2448 a_6606_4801# check[5] 1.24e-20
C2449 a_11250_4775# a_11195_4112# 8.14e-21
C2450 VDD a_12031_4775# 0.709f
C2451 a_8696_2366# check[4] 1.1e-20
C2452 a_10794_3239# a_11857_4801# 6.75e-21
C2453 check[4] a_11390_4801# 1.64e-19
C2454 a_1762_2340# eob 2.19e-19
C2455 x77.Y a_3599_2340# 2.75e-19
C2456 x4.X a_4074_4775# 0.00101f
C2457 x4.X x20.Q_N 0.274f
C2458 a_7049_2340# x4.X 0.00149f
C2459 x4.X a_11250_4775# 9.45e-19
C2460 a_1762_2340# x4.A 3.45e-19
C2461 a_5562_4801# check[6] 0.133f
C2462 D[1] a_11088_2366# 3.91e-20
C2463 a_4586_4801# x27.Q_N 1.61e-19
C2464 a_9236_2640# a_9441_2340# 0.153f
C2465 a_11856_3239# a_11965_3239# 0.00707f
C2466 a_8696_2366# x60.Q_N 0.00553f
C2467 a_5896_2340# check[0] 0.028f
C2468 a_12030_3213# x66.Q_N 0.124f
C2469 check[1] a_9375_4478# 6.38e-20
C2470 a_5844_3239# a_5896_2340# 4.5e-19
C2471 a_9236_2640# x36.Q_N 0.00112f
C2472 a_12738_4801# check[3] 0.175f
C2473 a_11762_4801# x36.Q_N 4.04e-20
C2474 x5.X a_7264_4394# 3.07e-19
C2475 D[3] x4.X 5.34e-19
C2476 a_1112_2340# x4.X 0.0104f
C2477 sel_bit[0] a_3876_6040# 0.00262f
C2478 x66.Q_N x4.X 0.00462f
C2479 VDD a_9173_4478# 0.00371f
C2480 a_2060_2640# a_2479_2648# 2.46e-19
C2481 a_1520_2366# a_2979_2366# 6.59e-21
C2482 a_2265_2340# a_2198_2732# 9.46e-19
C2483 x51.Q_N a_1720_2648# 2.02e-20
C2484 a_1207_2340# D[6] 3.57e-20
C2485 check[0] a_4658_4086# 7.37e-19
C2486 a_3599_2340# check[6] 2.38e-20
C2487 a_10155_2366# a_11629_2340# 3.65e-21
C2488 a_7072_3239# a_5845_4801# 4.76e-21
C2489 a_6759_3213# a_6466_4775# 7.57e-21
C2490 D[3] a_11628_2640# 4.01e-20
C2491 a_12146_3239# a_11833_2340# 3.49e-20
C2492 VDD a_7182_4801# 7.87e-19
C2493 comparator_out a_4454_4086# 3.22e-20
C2494 comparator_out a_12548_4112# 4.04e-20
C2495 check[2] a_4368_4775# 1.3e-19
C2496 x4.X a_8591_4801# 2.37e-19
C2497 a_6781_4112# a_7186_4112# 2.46e-21
C2498 a_8289_4086# a_8384_4086# 0.0968f
C2499 D[1] check[2] 0.171f
C2500 D[6] a_4018_2366# 0.0021f
C2501 a_3619_4801# a_5845_4801# 4e-20
C2502 a_3453_4801# a_6011_4801# 2.9e-21
C2503 a_3599_2340# a_3912_2366# 0.273f
C2504 a_6010_3239# a_6399_3239# 0.0019f
C2505 a_6465_3213# a_6605_3239# 0.07f
C2506 a_6759_3213# a_6930_3521# 0.00652f
C2507 a_8237_4801# a_8403_4801# 0.751f
C2508 x36.Q_N a_11089_4112# 1.39e-22
C2509 comparator_out a_12101_2550# 0.00818f
C2510 x75.Q a_6759_3213# 9.18e-20
C2511 a_4680_3239# a_4452_2640# 1.11e-20
C2512 a_4367_3213# a_4657_2340# 0.00144f
C2513 a_4854_3213# a_4453_2340# 8.72e-19
C2514 a_3504_2340# VDD 0.205f
C2515 D[5] a_5896_2340# 0.0999f
C2516 a_3618_3239# x75.Q_N 1.93e-21
C2517 a_4680_3239# a_4766_3605# 0.00976f
C2518 D[0] a_8590_3239# 5.04e-19
C2519 a_6605_3239# a_5991_2340# 4.6e-20
C2520 a_3618_3239# a_3913_4112# 4.9e-19
C2521 a_4073_3213# a_3600_4086# 2.45e-19
C2522 a_4367_3213# VDD 0.356f
C2523 a_4074_4775# a_4368_4775# 0.199f
C2524 a_3453_4801# a_4681_4801# 0.0334f
C2525 a_3619_4801# a_4855_4775# 0.0265f
C2526 x5.X a_8684_5167# 0.00465f
C2527 a_6606_4801# x45.Q_N 2.3e-19
C2528 x30.Q_N a_6845_4386# 0.0327f
C2529 x20.Q_N a_4368_4775# 3e-20
C2530 a_2853_5648# a_3258_5648# 0.0197f
C2531 a_10776_4086# a_11630_4086# 0.0492f
C2532 a_11089_4112# a_11629_4386# 0.139f
C2533 x5.X check[0] 0.789f
C2534 a_7362_3239# VDD 4.88e-19
C2535 a_9573_3239# x42.Q_N 7.87e-19
C2536 a_3618_3239# x4.X 0.0489f
C2537 a_9151_3213# a_10982_3239# 3.42e-20
C2538 a_9638_3213# a_11856_3239# 1.86e-21
C2539 a_7247_4775# a_8403_4801# 2.64e-19
C2540 a_7073_4801# a_8237_4801# 6.38e-20
C2541 sel_bit[0] x48.Q 0.0566f
C2542 a_2853_5648# sel_bit[1] 0.0368f
C2543 x54.Q_N x27.Q_N 4.08e-19
C2544 a_5844_3239# x5.X 8.91e-20
C2545 a_9172_2366# x30.Q_N 1.14e-20
C2546 VDD check[4] 0.5f
C2547 a_5844_3239# a_6292_5167# 8.3e-21
C2548 x69.Q_N check[4] 0.00316f
C2549 a_11250_4775# a_11544_4775# 0.199f
C2550 a_10795_4801# a_12031_4775# 0.0264f
C2551 x77.Y x48.Q 6.96e-20
C2552 a_10629_4801# a_11857_4801# 0.0334f
C2553 a_2883_5674# a_1511_4112# 1.46e-20
C2554 x77.Y a_6010_3239# 0.00188f
C2555 a_4454_4086# a_4591_4478# 0.00907f
C2556 VDD a_2883_5674# 0.172f
C2557 comparator_out reset 2.03e-20
C2558 a_9464_3239# x4.X 0.00475f
C2559 VDD a_4389_4112# 9.51e-19
C2560 D[1] D[3] 0.345f
C2561 D[2] VDD 0.29f
C2562 a_8858_4775# a_9238_4086# 0.00336f
C2563 a_8403_4801# a_9442_4086# 0.00221f
C2564 a_9639_4775# a_8697_4112# 0.00161f
C2565 a_9152_4775# a_8939_4086# 3.72e-19
C2566 D[4] x60.Q_N 0.00109f
C2567 a_11249_3213# D[2] 1.23e-20
C2568 x60.Q_N VDD 0.0716f
C2569 a_8236_3239# a_8237_4801# 6.9e-19
C2570 a_3258_5648# a_3671_5674# 3.58e-19
C2571 a_10775_2340# check[4] 7.18e-21
C2572 comparator_out a_4388_2732# 1.8e-19
C2573 a_11543_3213# x36.Q_N 0.00494f
C2574 x4.X a_5170_4478# 9.15e-19
C2575 x77.Y a_4793_2366# 5.33e-22
C2576 a_5897_4086# x45.Q_N 0.182f
C2577 a_6305_4112# a_6547_4086# 0.124f
C2578 a_5992_4086# a_6845_4386# 0.0264f
C2579 a_9237_2340# x4.X 0.00274f
C2580 x75.Q comparator_out 0.00133f
C2581 x5.X a_6376_5167# 4.16e-19
C2582 a_6010_3239# check[6] 9.27e-20
C2583 a_1207_2340# a_2060_2640# 0.0264f
C2584 a_1520_2366# a_1762_2340# 0.124f
C2585 a_12030_3213# a_12547_2366# 2.38e-19
C2586 a_6292_5167# a_6376_5167# 0.00972f
C2587 a_7247_4775# a_7073_4801# 0.197f
C2588 a_6760_4775# a_6199_4801# 8.23e-22
C2589 a_5845_4801# a_6710_5083# 0.00276f
C2590 a_9709_2550# a_11088_2366# 5.19e-21
C2591 a_9236_2640# a_11629_2340# 2.9e-21
C2592 a_9237_2340# a_11628_2640# 4e-20
C2593 a_9639_4775# a_11857_4801# 1.86e-21
C2594 a_11330_2340# x36.Q_N 0.16f
C2595 comparator_out a_10983_4801# 1.78e-20
C2596 a_12547_2366# x4.X 5.99e-20
C2597 D[5] x5.X 3.43e-19
C2598 check[2] a_10346_4801# 0.0147f
C2599 x27.D a_4539_5083# 3.01e-21
C2600 D[6] a_3599_2340# 0.0144f
C2601 a_2060_2640# a_4018_2366# 2.19e-20
C2602 a_2979_2366# a_3912_2366# 3.42e-20
C2603 a_11629_4386# a_11767_4478# 1.09e-19
C2604 a_11331_4086# a_11195_4112# 0.0282f
C2605 VDD a_11834_4086# 0.487f
C2606 a_4793_2366# check[6] 4.42e-19
C2607 a_11089_4112# a_12048_4394# 1.21e-20
C2608 eob a_2993_5674# 9.62e-20
C2609 a_11088_2366# a_11768_2366# 3.73e-19
C2610 a_11543_3213# a_11629_4386# 5.72e-19
C2611 a_10628_3239# x39.Q_N 0.0434f
C2612 a_11629_2340# a_12345_2732# 0.0018f
C2613 a_11833_2340# a_12047_2648# 0.0104f
C2614 a_10982_3239# a_10776_4086# 2.44e-19
C2615 a_11856_3239# a_11089_4112# 2.16e-19
C2616 a_11628_2640# a_12547_2366# 0.159f
C2617 a_11330_2340# a_11564_2366# 0.00707f
C2618 a_6291_3605# x30.Q_N 0.00193f
C2619 a_9754_3239# x33.Q_N 0.00342f
C2620 a_2389_5648# a_2883_5674# 0.169f
C2621 check[2] a_2784_5996# 6.63e-19
C2622 check[2] a_5897_4086# 1.35e-21
C2623 x5.X a_4389_4478# 4.04e-20
C2624 x4.X a_11331_4086# 0.00706f
C2625 a_9442_4086# a_9710_4296# 0.205f
C2626 a_9238_4086# x42.Q_N 0.00114f
C2627 a_2198_2732# VDD 0.0198f
C2628 a_8402_3239# a_9238_4086# 6.04e-20
C2629 a_9151_3213# a_8697_4112# 3.33e-20
C2630 a_8857_3213# a_9237_4386# 0.0015f
C2631 a_8683_3605# a_8939_4086# 1.7e-20
C2632 a_8236_3239# a_9442_4086# 0.00195f
C2633 a_3912_2366# a_4793_2366# 0.00943f
C2634 a_4154_2340# a_4592_2366# 0.00276f
C2635 a_4681_4801# a_4790_4801# 0.00707f
C2636 a_4453_2340# a_5896_2340# 8.18e-19
C2637 a_11629_2340# a_11089_4112# 1.4e-21
C2638 a_11628_2640# a_11331_4086# 4.75e-21
C2639 x5.X a_11943_5167# 1.78e-19
C2640 a_7072_3239# a_7362_3239# 0.0282f
C2641 a_7246_3213# a_7181_3239# 4.2e-20
C2642 a_6304_2366# x30.Q_N 0.0928f
C2643 a_8858_4775# a_8998_4801# 0.07f
C2644 a_9152_4775# a_9323_5083# 0.00652f
C2645 a_8403_4801# a_8792_4801# 0.0019f
C2646 a_8237_4801# a_9370_4801# 2.56e-19
C2647 x63.Q_N x33.Q_N 7.78e-20
C2648 a_3899_3605# a_4074_4775# 1.33e-23
C2649 a_4073_3213# a_3900_5167# 3.52e-21
C2650 a_4367_3213# a_3619_4801# 2.05e-21
C2651 a_3899_3605# x20.Q_N 2.96e-20
C2652 x48.Q a_2788_5674# 1.65e-19
C2653 a_6305_4112# a_6411_4112# 0.051f
C2654 a_6845_4386# a_6781_4478# 2.13e-19
C2655 a_6547_4086# a_6983_4478# 0.00412f
C2656 a_6846_4086# a_6505_4394# 1.25e-19
C2657 a_2289_4801# a_1511_4112# 0.00374f
C2658 a_11768_2366# check[2] 3.3e-19
C2659 a_6010_3239# a_6547_4086# 1.07e-20
C2660 a_6465_3213# a_6305_4112# 0.00148f
C2661 a_4925_2550# a_4453_4386# 6.45e-21
C2662 a_4452_2640# a_4926_4296# 6.02e-22
C2663 VDD a_2289_4801# 0.203f
C2664 a_6304_2366# a_6780_2732# 0.00133f
C2665 a_9464_3239# D[1] 5.18e-20
C2666 a_6011_4801# check[5] 1.26e-20
C2667 a_8802_2366# x30.Q_N 9.32e-20
C2668 check[1] a_4658_4086# 4.01e-21
C2669 x5.A a_2853_5648# 2.03e-20
C2670 check[4] a_10795_4801# 0.164f
C2671 a_1061_4801# a_2289_4801# 0.0334f
C2672 a_1227_4801# a_2463_4775# 0.0267f
C2673 x4.X a_1508_5167# 0.138f
C2674 a_1682_4775# a_1976_4775# 0.198f
C2675 a_1511_4112# a_4454_4086# 7.27e-20
C2676 a_3505_4086# a_4453_4386# 8.38e-21
C2677 a_3600_4086# a_4155_4086# 0.197f
C2678 check[2] a_11630_4086# 1.95e-19
C2679 VDD a_4454_4086# 0.809f
C2680 a_5991_2340# a_6305_4112# 5.05e-21
C2681 a_3900_5167# x27.Q_N 8.65e-20
C2682 a_4368_4775# a_5089_5083# 0.00185f
C2683 VDD a_12548_4112# 0.109f
C2684 D[1] a_9237_2340# 0.0263f
C2685 x5.X x33.Q_N 0.00113f
C2686 a_11159_3605# VDD 0.0042f
C2687 a_10794_3239# a_9754_3239# 9.75e-21
C2688 a_11543_3213# a_11856_3239# 0.124f
C2689 a_6845_2340# x60.Q_N 2.94e-19
C2690 a_11075_3605# a_10982_3239# 0.0367f
C2691 a_11249_3213# a_11159_3605# 6.69e-20
C2692 a_10155_2366# check[4] 0.00335f
C2693 x75.Q_N x4.X 0.00464f
C2694 check[0] x30.Q_N 0.00106f
C2695 x4.X a_3913_4112# 0.112f
C2696 a_5844_3239# x30.Q_N 2.88e-19
C2697 a_11076_5167# x36.Q_N 1.74e-20
C2698 a_11544_4775# a_12265_5083# 0.00185f
C2699 x4.X a_11195_4112# 0.00334f
C2700 a_12030_3213# x4.X 0.116f
C2701 a_4453_4386# x45.Q_N 2.05e-19
C2702 a_9237_4386# a_9377_4112# 0.00126f
C2703 a_8939_4086# a_9578_4112# 0.00316f
C2704 a_9710_4296# a_10156_4112# 0.0367f
C2705 a_4680_3239# comparator_out 1.77e-19
C2706 a_8683_3605# a_8803_4112# 1.12e-20
C2707 check[6] a_7073_4801# 4.06e-20
C2708 D[2] a_11965_3239# 9.32e-21
C2709 a_12101_2550# VDD 0.172f
C2710 a_12030_3213# a_11628_2640# 3.43e-19
C2711 a_11543_3213# a_11629_2340# 2.19e-19
C2712 a_8998_4801# x42.Q_N 2.35e-19
C2713 x33.Q_N a_9237_4386# 0.0344f
C2714 x66.Q_N a_12737_3239# 0.178f
C2715 a_9465_4801# check[4] 1.08e-19
C2716 comparator_out a_6504_2648# 1.52e-19
C2717 a_2853_5648# x27.D 3.86e-19
C2718 eob a_1822_4801# 0.00828f
C2719 a_11628_2640# x4.X 0.00712f
C2720 check[0] a_3373_5674# 0.0228f
C2721 check[2] a_2463_4775# 7.62e-20
C2722 a_2389_5648# a_2289_4801# 0.0019f
C2723 a_6010_3239# a_6411_4112# 4.04e-21
C2724 a_4453_2340# x5.X 2.59e-20
C2725 a_1822_4801# x4.A 2.88e-19
C2726 a_2979_2366# D[6] 6.09e-19
C2727 a_8696_2366# a_8803_4112# 8.38e-21
C2728 check[0] a_5992_4086# 0.0142f
C2729 a_6010_3239# a_6465_3213# 0.153f
C2730 D[3] a_11768_2366# 7.83e-20
C2731 a_2061_2340# a_2401_2366# 6.04e-20
C2732 a_2265_2340# a_2200_2366# 9.75e-19
C2733 a_2060_2640# a_3599_2340# 3.6e-19
C2734 a_11088_2366# a_11833_2340# 0.199f
C2735 a_5844_3239# a_5992_4086# 8.29e-19
C2736 a_11330_2340# a_11629_2340# 0.0334f
C2737 a_10775_2340# a_12101_2550# 4.7e-22
C2738 a_11544_4775# a_11331_4086# 3.72e-19
C2739 a_10795_4801# a_11834_4086# 0.00221f
C2740 a_11250_4775# a_11630_4086# 0.00336f
C2741 a_12031_4775# a_11089_4112# 0.00161f
C2742 check[1] x5.X 0.767f
C2743 a_3452_3239# a_3504_2340# 4.5e-19
C2744 check[1] a_6292_5167# 1.94e-19
C2745 check[2] a_4453_4386# 1.41e-20
C2746 a_1062_5674# a_1338_5674# 0.00104f
C2747 eob a_621_4112# 9.98e-19
C2748 a_10982_3239# check[2] 0.00707f
C2749 a_3452_3239# a_4367_3213# 0.125f
C2750 a_3618_3239# a_3899_3605# 0.152f
C2751 a_1996_2732# x20.Q_N 3.64e-19
C2752 a_4318_5083# check[6] 1.19e-21
C2753 D[6] a_4793_2366# 4.25e-19
C2754 a_4453_2340# a_4590_2732# 0.00907f
C2755 VDD a_6466_4775# 0.488f
C2756 a_6010_3239# a_5991_2340# 3.73e-19
C2757 D[5] x30.Q_N 0.00272f
C2758 a_621_4112# x4.A 6.66e-19
C2759 reset a_1511_4112# 1.58e-19
C2760 x3.A a_897_4112# 0.3f
C2761 x72.Q_N x30.Q_N 0.0201f
C2762 check[5] a_9102_5083# 8.63e-22
C2763 a_11543_3213# a_12147_4801# 1.05e-20
C2764 VDD reset 0.16f
C2765 check[1] a_9237_4386# 1.6e-19
C2766 a_11565_4112# a_10776_4086# 4.2e-20
C2767 a_11494_5083# check[3] 2.79e-19
C2768 x5.X a_7050_4086# 9.61e-19
C2769 a_11833_2340# check[2] 4.61e-19
C2770 a_6760_4775# a_6846_4086# 4.63e-19
C2771 a_2289_4801# a_3619_4801# 5.38e-20
C2772 a_7247_4775# a_6845_4386# 6.17e-19
C2773 a_9237_4386# a_9954_4112# 0.0019f
C2774 a_6011_4801# x45.Q_N 7.77e-20
C2775 a_4388_2732# VDD 0.00402f
C2776 VDD a_8939_4086# 0.34f
C2777 a_2463_4775# x20.Q_N 0.129f
C2778 a_9550_3605# x42.Q_N 3.64e-19
C2779 a_5896_2340# a_6844_2640# 8.38e-21
C2780 a_6930_3521# VDD 0.0163f
C2781 a_8383_2340# x30.Q_N 1.64e-19
C2782 a_8857_3213# a_9322_3521# 9.46e-19
C2783 a_8236_3239# a_8997_3239# 6.04e-20
C2784 a_8402_3239# a_9550_3605# 2.13e-19
C2785 a_9638_3213# check[4] 0.00527f
C2786 comparator_out x39.Q_N 6.03e-19
C2787 x75.Q VDD 0.216f
C2788 a_4073_3213# x27.Q_N 4.88e-19
C2789 x4.X a_7186_4112# 0.00311f
C2790 a_4970_3239# x4.X 5.69e-19
C2791 a_6846_4086# a_9238_4086# 1.37e-19
C2792 a_3900_5167# a_4155_4086# 2.46e-20
C2793 a_4368_4775# a_3913_4112# 5.67e-20
C2794 a_6305_4112# x42.Q_N 5.52e-21
C2795 a_3619_4801# a_4454_4086# 1.18e-19
C2796 a_4074_4775# a_4453_4386# 3.92e-19
C2797 a_3453_4801# a_4658_4086# 6.96e-19
C2798 x20.Q_N a_4453_4386# 1.28e-19
C2799 a_6709_3521# x45.Q_N 0.00136f
C2800 VDD a_3807_4801# 0.117f
C2801 D[1] a_12030_3213# 1.69e-20
C2802 a_9464_3239# a_9709_2550# 1.85e-20
C2803 a_9236_2640# check[4] 0.0285f
C2804 a_6978_4801# check[5] 1.84e-20
C2805 a_11543_3213# a_12031_4775# 1.08e-22
C2806 a_12030_3213# a_11544_4775# 1.06e-20
C2807 VDD a_10983_4801# 0.109f
C2808 a_5561_3239# x45.Q_N 1.19e-20
C2809 a_2061_2340# eob 0.00216f
C2810 check[4] a_11762_4801# 5.42e-20
C2811 x77.Y a_4154_2340# 0.00178f
C2812 a_1061_4801# a_3807_4801# 3.65e-21
C2813 x4.X a_4368_4775# 0.101f
C2814 a_1338_5674# x5.X 0.17f
C2815 D[1] x4.X 0.0011f
C2816 x57.Q_N x4.X 0.00786f
C2817 x27.Q_N a_5372_4112# 0.0147f
C2818 check[2] a_6011_4801# 1.18e-19
C2819 x4.X a_11544_4775# 0.105f
C2820 x77.Y a_4538_3521# 2.52e-20
C2821 a_9237_2340# a_9709_2550# 0.15f
C2822 a_9236_2640# x60.Q_N 5.14e-21
C2823 check[1] a_9656_4394# 1.56e-20
C2824 x30.Q_N x33.Q_N 2.51e-20
C2825 a_11769_4112# VDD 0.00445f
C2826 check[2] a_8697_4112# 0.00313f
C2827 x5.X a_7764_4112# 9.62e-19
C2828 a_3170_4801# a_3453_4801# 8.18e-19
C2829 VDD a_8803_4112# 0.00996f
C2830 a_2061_2340# a_2777_2732# 0.0018f
C2831 a_2265_2340# a_2479_2648# 0.0104f
C2832 a_4154_2340# check[6] 1.2e-19
C2833 a_1762_2340# D[6] 2.05e-19
C2834 a_2060_2640# a_2979_2366# 0.163f
C2835 a_6759_3213# a_6760_4775# 0.00121f
C2836 D[3] a_11833_2340# 6.82e-20
C2837 VDD a_9323_5083# 0.0163f
C2838 a_11564_2366# x36.Q_N 9.42e-19
C2839 x4.X a_8897_4394# 1.75e-19
C2840 x5.X a_3453_4801# 0.255f
C2841 check[2] a_4681_4801# 4.32e-20
C2842 x4.X a_7363_4801# 0.00557f
C2843 a_10680_2340# a_10681_4086# 1.07e-20
C2844 a_3912_2366# a_4154_2340# 0.124f
C2845 a_3599_2340# a_4452_2640# 0.0264f
C2846 x5.X a_10629_4801# 0.27f
C2847 a_3504_2340# x54.Q_N 0.178f
C2848 a_7246_3213# a_7158_3605# 7.71e-20
C2849 a_7072_3239# a_6930_3521# 0.00412f
C2850 a_6465_3213# a_6977_3239# 9.75e-19
C2851 a_6291_3605# a_6399_3239# 0.00812f
C2852 a_6759_3213# a_6605_3239# 0.00943f
C2853 a_4453_2340# x30.Q_N 1.57e-19
C2854 a_8403_4801# a_8858_4775# 0.153f
C2855 a_8237_4801# a_8684_5167# 0.15f
C2856 a_11390_4801# x39.Q_N 2.02e-19
C2857 x36.Q_N a_11629_4386# 0.0351f
C2858 a_4680_3239# a_4657_2340# 1.03e-19
C2859 a_4854_3213# a_4925_2550# 1.66e-21
C2860 check[1] x30.Q_N 0.0373f
C2861 a_1227_4801# a_897_4112# 4.21e-19
C2862 x48.Q a_4113_4394# 5.88e-19
C2863 a_3504_2340# a_3600_4086# 2.97e-20
C2864 x48.Q a_4539_5083# 6.59e-19
C2865 a_4971_4801# a_4926_4296# 1.9e-20
C2866 a_2200_2366# VDD 0.00214f
C2867 a_4925_2550# a_5169_2366# 0.00812f
C2868 a_4367_3213# a_5088_3521# 0.00185f
C2869 a_11194_2366# x39.Q_N 5e-20
C2870 D[0] a_7362_3239# 8.51e-20
C2871 a_7763_2366# x30.Q_N 0.0318f
C2872 VDD a_7481_5083# 0.00506f
C2873 a_3899_3605# a_3913_4112# 1.61e-19
C2874 a_3618_3239# a_4453_4386# 4.11e-20
C2875 a_3452_3239# a_4454_4086# 6.54e-20
C2876 a_4073_3213# a_4155_4086# 1.02e-19
C2877 a_4367_3213# a_3600_4086# 8.83e-19
C2878 a_4680_3239# VDD 0.183f
C2879 check[2] a_9375_4478# 1.05e-20
C2880 x4.X a_6606_4801# 7.25e-19
C2881 a_4074_4775# a_4681_4801# 0.00187f
C2882 a_3900_5167# a_4855_4775# 4.7e-22
C2883 a_3619_4801# a_3807_4801# 0.162f
C2884 a_3453_4801# a_3984_5167# 0.0018f
C2885 a_6504_2648# VDD 0.00506f
C2886 a_10776_4086# a_12102_4296# 4.7e-22
C2887 a_9578_4112# x39.Q_N 5.6e-20
C2888 a_1822_4801# a_2398_4801# 2.46e-21
C2889 check[2] a_9102_5083# 1.52e-19
C2890 a_11331_4086# a_11630_4086# 0.0334f
C2891 a_11089_4112# a_11834_4086# 0.199f
C2892 x5.X a_9639_4775# 0.00985f
C2893 x20.Q_N a_4681_4801# 2.69e-20
C2894 a_6304_2366# a_6780_2366# 2.87e-21
C2895 check[1] a_3373_5674# 0.027f
C2896 a_2853_5648# a_3876_6040# 0.00747f
C2897 a_9101_3521# VDD 0.00984f
C2898 a_3899_3605# x4.X 0.018f
C2899 a_9151_3213# a_9754_3239# 0.0552f
C2900 a_7247_4775# a_8684_5167# 7.98e-21
C2901 a_11543_3213# check[4] 8.39e-21
C2902 check[1] a_5992_4086# 5.87e-20
C2903 a_4854_3213# x45.Q_N 1.37e-20
C2904 comparator_out a_1207_2340# 6.22e-19
C2905 a_3258_5648# a_1511_4112# 3.06e-19
C2906 a_10795_4801# a_10983_4801# 0.162f
C2907 a_11076_5167# a_12031_4775# 4.7e-22
C2908 a_10629_4801# a_11160_5167# 0.0018f
C2909 a_11250_4775# a_11857_4801# 0.00187f
C2910 sel_bit[1] a_1511_4112# 3.24e-20
C2911 VDD a_3258_5648# 0.116f
C2912 a_4453_4386# a_5170_4478# 4.45e-20
C2913 a_3600_4086# a_4389_4112# 4.2e-20
C2914 a_4454_4086# a_4872_4394# 0.00276f
C2915 a_8767_3605# x4.X 9.07e-19
C2916 VDD sel_bit[1] 0.381f
C2917 x4.X a_10346_4801# 0.0067f
C2918 VDD a_4794_4112# 0.0336f
C2919 x27.Q_N a_4155_4086# 1.3e-22
C2920 a_7181_3239# x45.Q_N 7.87e-19
C2921 clk_sar a_897_4112# 1.96e-20
C2922 a_8383_2340# a_8896_2648# 0.00945f
C2923 a_12030_3213# a_12737_3239# 0.0968f
C2924 a_8403_4801# x42.Q_N 7.79e-20
C2925 a_9152_4775# a_9238_4086# 4.63e-19
C2926 a_9639_4775# a_9237_4386# 6.17e-19
C2927 a_11543_3213# D[2] 3.13e-19
C2928 a_8402_3239# a_8403_4801# 1.39e-19
C2929 a_3373_5674# a_3877_5674# 5.33e-19
C2930 comparator_out a_9238_4086# 3.21e-20
C2931 sel_bit[1] a_1061_4801# 7.54e-20
C2932 a_11856_3239# x36.Q_N 0.00293f
C2933 x4.X a_5897_4086# 0.00454f
C2934 a_12737_3239# x4.X 0.00277f
C2935 a_6305_4112# a_6846_4086# 0.125f
C2936 a_6547_4086# a_6845_4386# 0.137f
C2937 a_4593_4112# x45.Q_N 3.1e-20
C2938 a_9709_2550# x4.X 0.00146f
C2939 check[1] eob 0.00405f
C2940 a_1762_2340# a_2060_2640# 0.137f
C2941 a_1520_2366# a_2061_2340# 0.125f
C2942 a_6466_4775# a_6710_5083# 0.0104f
C2943 a_6011_4801# a_6931_5083# 1.09e-19
C2944 D[2] a_11330_2340# 2.3e-20
C2945 a_6780_2366# check[0] 1.28e-19
C2946 comparator_out a_8288_2340# 7.84e-19
C2947 a_11629_2340# x36.Q_N 0.0468f
C2948 a_9152_4775# a_9755_4801# 0.0552f
C2949 sel_bit[0] a_621_4112# 8.01e-21
C2950 D[6] a_4154_2340# 8.45e-19
C2951 a_11629_4386# a_12048_4394# 2.46e-19
C2952 x39.Q_N a_11289_4394# 2.02e-20
C2953 a_11834_4086# a_11767_4478# 9.46e-19
C2954 a_6304_2366# check[6] 2.39e-20
C2955 x30.Q_N a_7764_4112# 0.0147f
C2956 a_12030_3213# a_11630_4086# 7.94e-19
C2957 a_11543_3213# a_11834_4086# 0.0014f
C2958 a_11249_3213# x39.Q_N 0.194f
C2959 VDD x39.Q_N 0.458f
C2960 a_11330_2340# a_11969_2366# 0.00316f
C2961 a_11833_2340# a_12547_2366# 6.99e-20
C2962 a_12101_2550# a_12345_2732# 0.00972f
C2963 a_11628_2640# a_11768_2366# 0.00126f
C2964 x72.Q_N a_7247_4775# 4.45e-20
C2965 a_7246_3213# x30.Q_N 0.0127f
C2966 a_2853_5648# x48.Q 0.016f
C2967 a_2389_5648# a_3258_5648# 0.0296f
C2968 sel_bit[0] check[0] 0.163f
C2969 a_2389_5648# sel_bit[1] 0.0628f
C2970 a_4854_3213# a_6198_3239# 8.26e-21
C2971 x77.Y check[0] 2.24e-20
C2972 x4.X a_11630_4086# 0.0441f
C2973 VDD a_6505_4394# 0.00506f
C2974 a_3618_3239# a_5561_3239# 3.23e-21
C2975 x77.Y a_5844_3239# 2.13e-19
C2976 a_3452_3239# x75.Q 6.31e-20
C2977 a_9710_4296# x42.Q_N 0.00244f
C2978 a_8236_3239# x42.Q_N 0.0435f
C2979 a_9151_3213# a_9237_4386# 5.72e-19
C2980 a_5169_2732# a_5371_2366# 8.94e-19
C2981 a_2479_2648# VDD 0.0122f
C2982 a_9464_3239# a_8697_4112# 2.16e-19
C2983 a_8590_3239# a_8384_4086# 2.44e-19
C2984 a_8236_3239# a_8402_3239# 0.782f
C2985 a_1996_2366# x20.Q_N 7.87e-19
C2986 a_11629_2340# a_11629_4386# 7.25e-19
C2987 a_4453_2340# a_4592_2366# 2.56e-19
C2988 a_10775_2340# x39.Q_N 2.2e-19
C2989 a_4452_2640# a_4793_2366# 0.00118f
C2990 a_11628_2640# a_11630_4086# 7.02e-19
C2991 a_3912_2366# a_6304_2366# 8.41e-21
C2992 a_4154_2340# a_5991_2340# 1.86e-21
C2993 a_1112_2340# a_897_4112# 4.64e-19
C2994 x27.Q_N a_5845_4801# 4.37e-19
C2995 x63.Q_N a_10776_4086# 2.32e-20
C2996 a_7480_3521# a_8236_3239# 4.06e-20
C2997 a_6844_2640# x30.Q_N 0.57f
C2998 x5.X a_11184_4801# 2.88e-19
C2999 a_9465_4801# a_9323_5083# 0.00412f
C3000 a_8237_4801# x33.Q_N 1.26e-19
C3001 a_8684_5167# a_8792_4801# 0.00812f
C3002 a_8858_4775# a_9370_4801# 9.75e-19
C3003 a_9639_4775# a_9551_5167# 7.71e-20
C3004 a_9152_4775# a_8998_4801# 0.00943f
C3005 a_3618_3239# a_4681_4801# 6.75e-21
C3006 x48.Q a_3671_5674# 0.0017f
C3007 a_1996_2732# x4.X 4.32e-19
C3008 x36.Q_N a_12147_4801# 3.8e-19
C3009 x45.Q_N a_5170_4112# 3.4e-20
C3010 a_6846_4086# a_6983_4478# 0.00907f
C3011 a_12345_2366# check[2] 2.05e-20
C3012 a_6465_3213# a_6845_4386# 0.0015f
C3013 a_6759_3213# a_6305_4112# 3.33e-20
C3014 a_6010_3239# a_6846_4086# 6.04e-20
C3015 a_6291_3605# a_6547_4086# 1.7e-20
C3016 a_4925_2550# a_4658_4086# 2.22e-22
C3017 x5.X check[5] 0.17f
C3018 a_9236_2640# a_8939_4086# 4.75e-21
C3019 a_9237_2340# a_8697_4112# 1.4e-21
C3020 a_6845_2340# a_6504_2648# 1.25e-19
C3021 a_6304_2366# a_6410_2366# 0.0552f
C3022 VDD a_1592_5167# 0.00558f
C3023 a_4388_2366# VDD 1.64e-19
C3024 a_6546_2340# a_6982_2732# 0.00412f
C3025 a_6844_2640# a_6780_2732# 2.13e-19
C3026 D[5] a_6780_2366# 3.51e-20
C3027 a_6760_4775# a_7954_4801# 6.04e-19
C3028 a_4789_3239# x27.Q_N 1.68e-19
C3029 a_7362_3239# a_7317_2550# 1.01e-20
C3030 a_6292_5167# check[5] 7.62e-21
C3031 a_10345_3239# check[4] 0.0274f
C3032 check[0] check[6] 0.45f
C3033 a_1338_5674# eob 5.41e-19
C3034 a_5844_3239# check[6] 0.00782f
C3035 check[4] a_11076_5167# 0.0011f
C3036 a_3373_5674# a_3453_4801# 1.45e-21
C3037 a_1227_4801# a_1415_4801# 0.163f
C3038 a_1061_4801# a_1592_5167# 0.0018f
C3039 x4.X a_2463_4775# 0.148f
C3040 a_1682_4775# a_2289_4801# 0.00187f
C3041 a_3913_4112# a_4453_4386# 0.139f
C3042 a_1338_5674# x4.A 2.32e-21
C3043 a_3600_4086# a_4454_4086# 0.0492f
C3044 a_2969_6040# x20.Q_N 1.2e-20
C3045 a_4855_4775# a_5372_4112# 4.23e-19
C3046 x5.X a_10776_4086# 0.0184f
C3047 check[2] a_12102_4296# 4.54e-20
C3048 VDD a_4926_4296# 0.319f
C3049 VDD x5.A 0.23f
C3050 a_4855_4775# x27.Q_N 0.128f
C3051 a_6984_2366# a_7185_2366# 3.34e-19
C3052 a_8288_2340# a_8696_2366# 6.04e-19
C3053 a_10628_3239# a_11714_3521# 0.00907f
C3054 a_10794_3239# a_11493_3521# 2.46e-19
C3055 a_3912_2366# check[0] 2.06e-21
C3056 a_12147_4801# a_11629_4386# 8.84e-21
C3057 comparator_out a_3599_2340# 0.00328f
C3058 x4.X a_4453_4386# 0.0483f
C3059 check[1] a_8237_4801# 0.00245f
C3060 a_12031_4775# x36.Q_N 0.126f
C3061 x4.X a_12346_4478# 9.15e-19
C3062 a_10982_3239# x4.X 0.00531f
C3063 a_4658_4086# x45.Q_N 3.93e-20
C3064 a_9238_4086# a_9578_4112# 6.04e-20
C3065 a_9442_4086# a_9377_4112# 9.75e-19
C3066 x42.Q_N a_10681_4086# 1.37e-20
C3067 a_9237_4386# a_10776_4086# 1.52e-19
C3068 a_12030_3213# a_11833_2340# 2.52e-19
C3069 a_11543_3213# a_12101_2550# 1.62e-19
C3070 a_6410_2366# check[0] 0.00226f
C3071 comparator_out a_6982_2732# 9.43e-19
C3072 eob a_3453_4801# 5.9e-20
C3073 eob a_2194_4801# 0.00151f
C3074 a_11833_2340# x4.X 0.00145f
C3075 a_6291_3605# a_6411_4112# 1.12e-20
C3076 a_7953_3239# x5.X 0.00125f
C3077 D[5] check[6] 0.141f
C3078 VDD x27.D 0.294f
C3079 a_2061_2340# a_3912_2366# 3.12e-19
C3080 a_6465_3213# a_6291_3605# 0.205f
C3081 a_2060_2640# a_4154_2340# 4.16e-20
C3082 a_2533_2550# a_2401_2366# 0.0258f
C3083 check[0] a_6547_4086# 3.86e-19
C3084 a_6010_3239# a_6759_3213# 0.139f
C3085 a_11088_2366# x63.Q_N 0.00553f
C3086 a_11628_2640# a_11833_2340# 0.153f
C3087 comparator_out a_6305_4112# 2.29e-20
C3088 a_10795_4801# x39.Q_N 7.79e-20
C3089 a_12031_4775# a_11629_4386# 6.17e-19
C3090 a_11544_4775# a_11630_4086# 4.63e-19
C3091 check[1] a_7247_4775# 0.0127f
C3092 x33.Q_N a_9574_4801# 7.27e-21
C3093 a_1227_4801# a_3170_4801# 1.76e-19
C3094 a_1061_4801# x27.D 5.94e-20
C3095 x5.A a_2389_5648# 6.17e-20
C3096 x5.X a_3505_4086# 0.00259f
C3097 a_1062_5674# check[2] 1.82e-20
C3098 check[2] a_4658_4086# 4.4e-21
C3099 clk_sar a_1062_5674# 0.185f
C3100 a_1207_2340# a_1511_4112# 1.58e-19
C3101 x5.X a_11565_4478# 1.76e-19
C3102 a_6304_2366# a_6411_4112# 8.38e-21
C3103 a_4073_3213# a_4367_3213# 0.198f
C3104 a_3452_3239# a_4680_3239# 0.0334f
C3105 a_3618_3239# a_4854_3213# 0.0264f
C3106 a_1626_2366# x20.Q_N 0.00967f
C3107 a_3912_2366# D[5] 2.89e-20
C3108 a_4453_2340# a_4871_2648# 0.00276f
C3109 a_4452_2640# a_5169_2732# 4.45e-20
C3110 a_6465_3213# a_6304_2366# 0.0014f
C3111 a_6291_3605# a_5991_2340# 3.9e-20
C3112 a_1207_2340# VDD 0.608f
C3113 VDD a_6760_4775# 0.449f
C3114 a_11965_3239# x39.Q_N 7.87e-19
C3115 a_9151_3213# x30.Q_N 8.28e-21
C3116 a_9953_2366# x33.Q_N 0.00224f
C3117 a_12264_3521# x39.Q_N 2.75e-19
C3118 check[1] a_9442_4086# 1.18e-19
C3119 a_11769_4112# a_11089_4112# 3.73e-19
C3120 a_11565_4112# a_11331_4086# 0.00707f
C3121 x5.X a_1227_4801# 0.0165f
C3122 a_11943_5167# check[3] 4.39e-19
C3123 x4.X a_6011_4801# 0.00494f
C3124 x5.X x45.Q_N 0.00731f
C3125 a_6760_4775# a_7318_4296# 2.85e-19
C3126 x63.Q_N check[2] 0.0121f
C3127 a_7247_4775# a_7050_4086# 4.44e-19
C3128 a_6292_5167# x45.Q_N 9.97e-20
C3129 D[5] a_6410_2366# 5.42e-19
C3130 x75.Q_N a_5561_3239# 0.178f
C3131 a_4018_2366# VDD 0.0028f
C3132 x4.X a_11966_4801# 2.39e-19
C3133 VDD a_9238_4086# 0.805f
C3134 a_3504_2340# x27.Q_N 3.7e-19
C3135 a_8236_3239# a_10628_3239# 0.00176f
C3136 a_1415_4801# x20.Q_N 5.43e-21
C3137 a_5991_2340# a_6304_2366# 0.273f
C3138 a_8402_3239# a_8791_3239# 0.0019f
C3139 a_6605_3239# VDD 5.47e-21
C3140 a_9151_3213# a_9322_3521# 0.00652f
C3141 a_8236_3239# a_9369_3239# 2.56e-19
C3142 a_8857_3213# a_8997_3239# 0.07f
C3143 x27.Q_N a_6400_4801# 2.58e-20
C3144 x33.Q_N a_10156_4112# 0.0147f
C3145 a_8938_2340# x30.Q_N 5.93e-20
C3146 a_4367_3213# x27.Q_N 0.00484f
C3147 a_4112_2648# x4.X 0.00102f
C3148 x4.X a_8697_4112# 0.109f
C3149 a_6709_3521# x4.X 2.91e-19
C3150 a_3807_4801# a_3600_4086# 3.44e-19
C3151 a_2579_4801# a_1511_4112# 3.99e-19
C3152 check[2] a_3170_4801# 1.57e-20
C3153 a_4368_4775# a_4453_4386# 7.46e-19
C3154 a_4681_4801# a_3913_4112# 3.76e-19
C3155 a_6845_4386# x42.Q_N 1.95e-19
C3156 x20.Q_N a_4658_4086# 2.19e-20
C3157 D[4] a_8288_2340# 0.1f
C3158 a_7158_3605# x45.Q_N 3.63e-19
C3159 check[0] a_6411_4112# 4.09e-19
C3160 VDD a_2579_4801# 0.0073f
C3161 a_8288_2340# VDD 0.189f
C3162 a_5561_3239# x4.X 0.00286f
C3163 D[1] a_10982_3239# 4.96e-19
C3164 a_8997_3239# a_8383_2340# 4.6e-20
C3165 x30.Q_N check[5] 0.902f
C3166 a_9441_2340# check[4] 7.03e-20
C3167 VDD a_9755_4801# 0.0101f
C3168 a_11856_3239# a_12031_4775# 1.33e-23
C3169 a_12030_3213# a_11857_4801# 4.82e-21
C3170 comparator_out x48.Q 3.3e-20
C3171 comparator_out a_2979_2366# 0.157f
C3172 a_5844_3239# a_6465_3213# 0.117f
C3173 comparator_out a_6010_3239# 0.149f
C3174 a_9953_2366# check[1] 2.06e-20
C3175 a_2533_2550# eob 4.21e-20
C3176 x77.Y a_4453_2340# 3.65e-20
C3177 check[4] x36.Q_N 8.5e-21
C3178 x4.X a_4681_4801# 0.00584f
C3179 check[2] x5.X 0.831f
C3180 sel_bit[0] check[1] 0.583f
C3181 clk_sar x5.X 0.00891f
C3182 check[2] a_6292_5167# 5.02e-20
C3183 x4.X a_11857_4801# 0.00316f
C3184 x77.Y a_4213_3239# 0.0313f
C3185 a_5991_2340# check[0] 0.0146f
C3186 a_8237_4801# a_10629_4801# 0.00176f
C3187 D[2] x36.Q_N 0.00122f
C3188 a_5844_3239# a_5991_2340# 8.35e-19
C3189 a_11565_4112# a_11195_4112# 4.11e-20
C3190 check[2] a_9237_4386# 0.163f
C3191 sel_bit[0] a_3877_5674# 2.93e-19
C3192 a_7247_4775# a_7764_4112# 4.23e-19
C3193 x27.D a_3619_4801# 0.159f
C3194 a_10156_4112# a_9954_4112# 3.67e-19
C3195 a_2533_2550# a_2777_2732# 0.00972f
C3196 a_2265_2340# a_2979_2366# 6.99e-20
C3197 VDD a_9954_4478# 0.0042f
C3198 a_2061_2340# D[6] 0.338f
C3199 a_10628_3239# a_10681_4086# 5.06e-19
C3200 a_4453_2340# check[6] 0.0409f
C3201 x48.Q a_4971_4801# 4.12e-19
C3202 x20.Q_N a_3170_4801# 0.187f
C3203 a_2697_5083# x27.D 7.73e-21
C3204 D[3] x63.Q_N 0.00107f
C3205 a_9638_3213# x39.Q_N 3.76e-21
C3206 a_7246_3213# a_7247_4775# 0.00237f
C3207 a_11565_4112# x4.X 8.15e-20
C3208 VDD a_8998_4801# 0.0332f
C3209 comparator_out a_9172_2732# 1.81e-19
C3210 a_8997_3239# x33.Q_N 6.08e-19
C3211 a_11969_2366# x36.Q_N 0.0403f
C3212 check[1] check[6] 6.18e-20
C3213 a_11970_4112# a_11088_2366# 1.26e-20
C3214 eob x3.A 0.00123f
C3215 x4.X a_9375_4478# 0.00114f
C3216 x5.X a_4074_4775# 3.66e-19
C3217 a_2389_5648# a_2579_4801# 2.13e-20
C3218 a_8289_4086# a_9238_4086# 7e-20
C3219 x5.X x20.Q_N 0.00434f
C3220 x3.A x4.A 4.66e-19
C3221 a_4368_4775# a_6011_4801# 1.1e-19
C3222 a_4855_4775# a_5845_4801# 0.00116f
C3223 a_12547_2366# a_12345_2366# 3.67e-19
C3224 a_12737_3239# a_11630_4086# 4.72e-19
C3225 a_6759_3213# a_8236_3239# 3.41e-19
C3226 a_11564_2366# a_11969_2366# 2.46e-21
C3227 a_3912_2366# a_4453_2340# 0.125f
C3228 a_4154_2340# a_4452_2640# 0.137f
C3229 VDD a_5562_4801# 0.192f
C3230 x5.X a_11250_4775# 0.00324f
C3231 a_7953_3239# x30.Q_N 0.00834f
C3232 a_7072_3239# a_6605_3239# 0.00316f
C3233 a_6759_3213# a_6977_3239# 3.73e-19
C3234 a_10680_2340# x33.Q_N 1.87e-19
C3235 a_8237_4801# a_9639_4775# 0.0492f
C3236 a_8403_4801# a_9152_4775# 0.139f
C3237 a_8858_4775# a_8684_5167# 0.205f
C3238 a_10794_3239# check[3] 1.56e-21
C3239 VDD a_12738_4801# 0.177f
C3240 comparator_out a_8403_4801# 2.9e-21
C3241 a_12031_4775# a_12147_4801# 0.0397f
C3242 a_11544_4775# a_11966_4801# 2.87e-21
C3243 x4.X a_897_4112# 1.27e-19
C3244 x48.Q a_4591_4478# 6.11e-19
C3245 D[3] x5.X 3.43e-19
C3246 a_8288_2340# a_8289_4086# 1.07e-20
C3247 D[5] a_5991_2340# 0.0123f
C3248 a_5371_2366# a_6304_2366# 3.42e-20
C3249 x48.Q a_4214_4801# 0.00132f
C3250 a_1338_5674# sel_bit[0] 0.0446f
C3251 a_3599_2340# VDD 0.58f
C3252 a_4854_3213# x75.Q_N 0.124f
C3253 a_4073_3213# a_4454_4086# 5.04e-19
C3254 a_4367_3213# a_4155_4086# 2.12e-19
C3255 a_3618_3239# a_4658_4086# 2.9e-19
C3256 a_11970_4112# check[2] 3.49e-20
C3257 a_4854_3213# a_3913_4112# 9.49e-19
C3258 a_3983_3605# VDD 0.00494f
C3259 check[2] a_9656_4394# 7.77e-21
C3260 x4.X a_6978_4801# 5.55e-19
C3261 a_4074_4775# a_3984_5167# 6.69e-20
C3262 a_4368_4775# a_4681_4801# 0.124f
C3263 a_3619_4801# a_2579_4801# 7.73e-20
C3264 a_3900_5167# a_3807_4801# 0.0367f
C3265 a_8802_2366# x42.Q_N 4.74e-20
C3266 a_6982_2732# VDD 0.0163f
C3267 x5.X a_8591_4801# 0.00545f
C3268 a_11629_4386# a_11834_4086# 0.153f
C3269 x30.Q_N x45.Q_N 0.0041f
C3270 a_6845_2340# a_8288_2340# 8.18e-19
C3271 a_6546_2340# a_6984_2366# 0.00276f
C3272 a_11089_4112# x39.Q_N 0.0933f
C3273 check[2] a_9551_5167# 1.87e-19
C3274 a_6304_2366# a_7185_2366# 0.00943f
C3275 a_2853_5648# a_2993_5674# 1.56e-19
C3276 a_9638_3213# a_9573_3239# 4.2e-20
C3277 a_4854_3213# x4.X 0.117f
C3278 a_9550_3605# VDD 0.00371f
C3279 a_9464_3239# a_9754_3239# 0.0282f
C3280 check[1] a_6547_4086# 7.52e-20
C3281 comparator_out a_1762_2340# 1.88e-19
C3282 a_11250_4775# a_11160_5167# 6.69e-20
C3283 a_11544_4775# a_11857_4801# 0.124f
C3284 a_11076_5167# a_10983_4801# 0.0367f
C3285 a_10795_4801# a_9755_4801# 4.87e-21
C3286 a_4453_4386# a_5897_4086# 3.56e-19
C3287 a_4658_4086# a_5170_4478# 6.69e-20
C3288 a_4155_4086# a_4389_4112# 0.00707f
C3289 VDD a_3876_6040# 0.00865f
C3290 a_4454_4086# a_5372_4112# 0.0664f
C3291 a_3913_4112# a_4593_4112# 3.73e-19
C3292 a_7181_3239# x4.X 1.05e-19
C3293 a_8384_4086# a_9173_4478# 7.71e-20
C3294 a_8697_4112# a_8897_4394# 0.00185f
C3295 VDD a_6305_4112# 0.448f
C3296 x27.Q_N a_4454_4086# 0.0256f
C3297 a_8696_2366# a_9172_2732# 0.00133f
C3298 a_11856_3239# D[2] 5.2e-20
C3299 a_9152_4775# a_9710_4296# 2.85e-19
C3300 a_8684_5167# x42.Q_N 9.99e-20
C3301 a_9639_4775# a_9442_4086# 4.44e-19
C3302 sel_bit[0] a_3453_4801# 4.34e-20
C3303 a_8683_3605# a_8403_4801# 8.52e-21
C3304 a_8402_3239# a_8684_5167# 1.65e-21
C3305 a_8857_3213# a_8858_4775# 2.59e-19
C3306 a_8236_3239# a_9152_4775# 9.66e-21
C3307 a_11629_2340# check[4] 1.57e-21
C3308 comparator_out a_5169_2732# 8.25e-19
C3309 a_5844_3239# a_8402_3239# 2.9e-21
C3310 x36.Q_N a_12548_4112# 0.0133f
C3311 comparator_out a_8236_3239# 0.147f
C3312 sel_bit[1] a_1682_4775# 1.09e-19
C3313 x77.Y a_3453_4801# 9.38e-22
C3314 x4.X a_4593_4112# 0.0012f
C3315 a_5844_3239# a_7480_3521# 1.25e-19
C3316 a_5992_4086# x45.Q_N 0.154f
C3317 a_6547_4086# a_7050_4086# 0.00187f
C3318 a_6845_4386# a_6846_4086# 0.75f
C3319 a_6305_4112# a_7318_4296# 0.0633f
C3320 check[2] x30.Q_N 6.73e-21
C3321 x5.X a_6931_5083# 5.11e-19
C3322 a_2060_2640# a_2061_2340# 0.783f
C3323 a_1207_2340# x51.Q_N 0.124f
C3324 a_1520_2366# a_2533_2550# 0.0633f
C3325 a_1762_2340# a_2265_2340# 0.00187f
C3326 D[2] a_11629_2340# 0.271f
C3327 a_6760_4775# a_6710_5083# 1.21e-20
C3328 a_9237_2340# x63.Q_N 2.94e-19
C3329 a_6199_4801# a_6376_5167# 8.94e-19
C3330 a_6011_4801# a_6606_4801# 0.00118f
C3331 a_7185_2366# check[0] 4.21e-19
C3332 check[0] a_4539_5083# 4.79e-19
C3333 a_9639_4775# a_9574_4801# 4.2e-20
C3334 a_9465_4801# a_9755_4801# 0.0282f
C3335 a_12101_2550# x36.Q_N 0.181f
C3336 a_3619_4801# a_5562_4801# 1.64e-20
C3337 a_3453_4801# check[6] 8.06e-20
C3338 D[6] a_4453_2340# 2.08e-19
C3339 a_11834_4086# a_12048_4394# 0.0104f
C3340 a_11630_4086# a_12346_4478# 0.0018f
C3341 a_11629_4386# a_12548_4112# 0.163f
C3342 a_11628_2640# a_12345_2366# 0.00105f
C3343 a_11856_3239# a_11834_4086# 4.33e-20
C3344 a_11543_3213# x39.Q_N 0.0983f
C3345 eob a_1227_4801# 0.413f
C3346 a_11629_2340# a_11969_2366# 6.04e-20
C3347 a_11833_2340# a_11768_2366# 9.75e-19
C3348 a_12030_3213# a_12102_4296# 3.74e-20
C3349 check[5] a_8237_4801# 0.414f
C3350 a_7954_4801# a_8403_4801# 5.4e-19
C3351 comparator_out a_11288_2648# 1.53e-19
C3352 check[1] a_6411_4112# 1.13e-20
C3353 check[2] a_3373_5674# 0.0404f
C3354 check[4] a_12147_4801# 1.37e-20
C3355 a_10629_4801# check[3] 0.00126f
C3356 a_10795_4801# a_12738_4801# 8.38e-21
C3357 a_4854_3213# a_4970_3239# 0.0397f
C3358 a_1227_4801# x4.A 0.00377f
C3359 a_4367_3213# a_4789_3239# 2.87e-21
C3360 check[2] a_5992_4086# 3.43e-20
C3361 x5.X a_5170_4478# 1.85e-19
C3362 x4.X a_12102_4296# 0.021f
C3363 x48.Q a_1511_4112# 0.00368f
C3364 a_2979_2366# a_1511_4112# 3.09e-20
C3365 VDD a_6983_4478# 0.0163f
C3366 a_1976_4775# a_2289_4801# 0.124f
C3367 a_9237_2340# x5.X 2.59e-20
C3368 a_1508_5167# a_1415_4801# 0.0367f
C3369 a_9638_3213# a_9238_4086# 7.94e-19
C3370 VDD x48.Q 0.638f
C3371 a_9151_3213# a_9442_4086# 0.0014f
C3372 a_2979_2366# VDD 0.117f
C3373 a_8857_3213# x42.Q_N 0.194f
C3374 a_6010_3239# VDD 0.274f
C3375 a_4657_2340# a_4793_2366# 0.07f
C3376 a_4453_2340# a_5991_2340# 0.00116f
C3377 a_2401_2366# x20.Q_N 0.0313f
C3378 a_4452_2640# a_6304_2366# 1.95e-19
C3379 a_8236_3239# a_8683_3605# 0.15f
C3380 a_8402_3239# a_8857_3213# 0.153f
C3381 a_11330_2340# x39.Q_N 0.0018f
C3382 a_9639_4775# a_10156_4112# 4.23e-19
C3383 x27.Q_N a_6466_4775# 1.88e-20
C3384 a_11628_2640# a_12102_4296# 6.02e-22
C3385 a_12101_2550# a_11629_4386# 6.45e-21
C3386 x72.Q_N a_8402_3239# 9.24e-20
C3387 x5.X a_12265_5083# 1.33e-19
C3388 a_7049_2340# x30.Q_N 0.179f
C3389 a_7480_3521# x72.Q_N 2.02e-20
C3390 comparator_out a_10681_4086# 2.05e-21
C3391 a_8858_4775# x33.Q_N 2.07e-20
C3392 a_9465_4801# a_8998_4801# 0.00316f
C3393 a_9152_4775# a_9370_4801# 3.73e-19
C3394 a_4367_3213# a_4855_4775# 1.08e-22
C3395 a_4854_3213# a_4368_4775# 1.06e-20
C3396 x4.X a_5170_4112# 7.21e-19
C3397 a_3806_3239# x20.Q_N 0.00103f
C3398 x48.Q a_1061_4801# 4.14e-21
C3399 a_1626_2366# x4.X 3.78e-20
C3400 a_6845_4386# a_7562_4478# 4.45e-20
C3401 a_6846_4086# a_7264_4394# 0.00276f
C3402 a_5992_4086# a_6781_4112# 4.2e-20
C3403 a_7072_3239# a_6305_4112# 2.16e-19
C3404 a_6198_3239# a_5992_4086# 2.44e-19
C3405 a_6759_3213# a_6845_4386# 5.72e-19
C3406 a_6845_2340# a_6982_2732# 0.00907f
C3407 x60.Q_N a_8384_4086# 2.32e-20
C3408 D[5] a_7185_2366# 7.82e-20
C3409 a_9236_2640# a_9238_4086# 7.02e-19
C3410 a_9237_2340# a_9237_4386# 7.25e-19
C3411 a_8383_2340# x42.Q_N 2.17e-19
C3412 VDD a_2147_5083# 0.0199f
C3413 a_8236_3239# a_8696_2366# 1.89e-19
C3414 a_8402_3239# a_8383_2340# 3.73e-19
C3415 D[7] a_2200_2366# 3.49e-19
C3416 a_4793_2366# VDD 9.91e-19
C3417 D[0] a_9573_3239# 1.29e-20
C3418 a_7247_4775# check[5] 0.0104f
C3419 check[2] eob 0.0123f
C3420 clk_sar eob 4.74e-20
C3421 check[4] a_12031_4775# 1.91e-20
C3422 a_1061_4801# a_2147_5083# 0.00907f
C3423 a_5896_2340# x4.X 0.00507f
C3424 x4.X a_1415_4801# 9.23e-21
C3425 a_1682_4775# a_1592_5167# 6.69e-20
C3426 a_3913_4112# a_4658_4086# 0.199f
C3427 a_3600_4086# a_4926_4296# 4.7e-22
C3428 a_3505_4086# x48.Q_N 0.178f
C3429 a_4155_4086# a_4454_4086# 0.0334f
C3430 a_6845_2340# a_6305_4112# 1.4e-21
C3431 a_6844_2640# a_6547_4086# 4.75e-21
C3432 x5.X a_11331_4086# 8.88e-19
C3433 a_9172_2732# VDD 0.00371f
C3434 a_8288_2340# a_9236_2640# 9.02e-21
C3435 a_3807_4801# x27.Q_N 5.03e-21
C3436 a_10628_3239# a_11389_3239# 6.04e-20
C3437 a_11249_3213# a_11714_3521# 9.46e-19
C3438 a_10794_3239# a_11942_3605# 2.13e-19
C3439 a_11714_3521# VDD 0.0163f
C3440 a_4452_2640# check[0] 2.1e-19
C3441 a_12147_4801# a_11834_4086# 7.76e-20
C3442 comparator_out a_4154_2340# 0.00109f
C3443 x4.X a_4658_4086# 0.0102f
C3444 a_10983_4801# x36.Q_N 5.41e-22
C3445 a_2853_5648# check[0] 0.164f
C3446 a_2389_5648# x48.Q 0.00138f
C3447 a_9754_3239# x4.X 5.61e-19
C3448 a_9238_4086# a_11089_4112# 5.07e-21
C3449 x42.Q_N a_9377_4112# 0.00167f
C3450 a_9710_4296# a_9578_4112# 0.0258f
C3451 a_9237_4386# a_11331_4086# 2.53e-20
C3452 a_6780_2366# check[5] 2.23e-20
C3453 a_11856_3239# a_12101_2550# 1.85e-20
C3454 VDD a_8403_4801# 0.593f
C3455 x33.Q_N x42.Q_N 0.00395f
C3456 x77.Y a_4019_4112# 1.79e-19
C3457 a_8402_3239# x33.Q_N 3.88e-19
C3458 sel_bit[0] x3.A 6.99e-21
C3459 comparator_out a_7263_2648# 6.92e-19
C3460 check[5] a_9574_4801# 1.69e-20
C3461 eob x20.Q_N 0.365f
C3462 x63.Q_N x4.X 0.00782f
C3463 check[0] a_3671_5674# 3.04e-19
C3464 x27.D a_3600_4086# 0.00292f
C3465 x5.X a_1508_5167# 0.00288f
C3466 x20.Q_N x4.A 5.76e-19
C3467 a_7953_3239# a_7247_4775# 4.94e-20
C3468 a_6010_3239# a_7072_3239# 0.137f
C3469 a_6291_3605# a_6759_3213# 0.0633f
C3470 a_2060_2640# a_4453_2340# 2.9e-21
C3471 a_2061_2340# a_4452_2640# 4e-20
C3472 a_2533_2550# a_3912_2366# 6.92e-21
C3473 check[0] a_6846_4086# 2.15e-19
C3474 a_11629_2340# a_12101_2550# 0.15f
C3475 a_11628_2640# x63.Q_N 5.46e-21
C3476 comparator_out a_6845_4386# 2.52e-20
C3477 a_5844_3239# a_6846_4086# 6.54e-20
C3478 a_11544_4775# a_12102_4296# 2.85e-19
C3479 a_6606_4801# a_6978_4801# 3.34e-19
C3480 a_12031_4775# a_11834_4086# 4.44e-19
C3481 a_11076_5167# x39.Q_N 1e-19
C3482 a_3452_3239# a_3599_2340# 8.35e-19
C3483 a_1112_2340# eob 3.79e-20
C3484 x4.X a_3170_4801# 9.94e-19
C3485 a_1682_4775# x27.D 2.67e-21
C3486 x5.X a_3913_4112# 1.32e-19
C3487 a_1762_2340# a_1511_4112# 4.16e-20
C3488 x48.Q a_3619_4801# 0.0352f
C3489 a_3452_3239# a_3983_3605# 0.0018f
C3490 a_3618_3239# a_3806_3239# 0.159f
C3491 a_4073_3213# a_4680_3239# 0.00187f
C3492 a_3899_3605# a_4854_3213# 4.7e-22
C3493 a_1112_2340# x4.A 7.47e-22
C3494 a_2777_2732# x20.Q_N 8.48e-19
C3495 a_4452_2640# D[5] 0.00524f
C3496 a_4657_2340# a_5169_2732# 6.69e-20
C3497 a_4453_2340# a_5371_2366# 0.0708f
C3498 a_1762_2340# VDD 0.201f
C3499 VDD a_7073_4801# 0.343f
C3500 a_6291_3605# a_6546_2340# 2.41e-20
C3501 a_6465_3213# a_6844_2640# 2.68e-19
C3502 a_6010_3239# a_6845_2340# 6.38e-20
C3503 a_6759_3213# a_6304_2366# 3.36e-20
C3504 a_6605_3239# D[0] 1.08e-20
C3505 check[5] a_8792_4801# 1.67e-19
C3506 check[1] x42.Q_N 0.0239f
C3507 a_11970_4112# a_11331_4086# 0.00316f
C3508 a_11769_4112# a_11629_4386# 0.00126f
C3509 a_8402_3239# check[1] 0.0363f
C3510 x5.X x4.X 0.0429f
C3511 x4.X a_6292_5167# 0.00132f
C3512 a_3912_2366# a_4019_4112# 8.38e-21
C3513 a_7073_4801# a_7318_4296# 3.59e-20
C3514 x42.Q_N a_9954_4112# 2.4e-19
C3515 check[2] a_8237_4801# 5.48e-19
C3516 a_10156_4112# a_10776_4086# 8.26e-21
C3517 a_9237_4386# a_11195_4112# 1.71e-20
C3518 a_1976_4775# a_3807_4801# 2.23e-21
C3519 a_2463_4775# a_4681_4801# 1.86e-21
C3520 a_4970_3239# a_4658_4086# 5.48e-21
C3521 a_5169_2732# VDD 0.00436f
C3522 a_10794_3239# x42.Q_N 9.16e-19
C3523 VDD a_9710_4296# 0.317f
C3524 a_8236_3239# D[4] 5.41e-19
C3525 D[0] a_8288_2340# 0.00665f
C3526 a_5896_2340# x57.Q_N 0.178f
C3527 a_5991_2340# a_6844_2640# 0.0264f
C3528 a_6304_2366# a_6546_2340# 0.124f
C3529 a_8236_3239# VDD 0.791f
C3530 a_9872_3521# x42.Q_N 2.75e-19
C3531 a_6977_3239# VDD 6.2e-19
C3532 a_8857_3213# a_9369_3239# 9.75e-19
C3533 a_9638_3213# a_9550_3605# 7.71e-20
C3534 a_9464_3239# a_9322_3521# 0.00412f
C3535 a_9151_3213# a_8997_3239# 0.00943f
C3536 a_8683_3605# a_8791_3239# 0.00812f
C3537 a_8236_3239# x69.Q_N 1.07e-19
C3538 a_9237_2340# x30.Q_N 8.11e-21
C3539 a_9873_5083# x33.Q_N 2.02e-20
C3540 a_4680_3239# x27.Q_N 0.0029f
C3541 x4.X a_9237_4386# 0.048f
C3542 a_4590_2732# x4.X 9.81e-19
C3543 a_7158_3605# x4.X 4.4e-19
C3544 a_4855_4775# a_4454_4086# 0.00169f
C3545 a_4368_4775# a_4658_4086# 0.00268f
C3546 a_4681_4801# a_4453_4386# 1.96e-20
C3547 a_7050_4086# x42.Q_N 1.92e-20
C3548 x20.Q_N x48.Q_N 0.00138f
C3549 VDD a_4318_5083# 0.0104f
C3550 a_7317_2550# a_7561_2366# 0.00812f
C3551 a_9577_2366# x42.Q_N 5.33e-22
C3552 a_6984_2366# VDD 6.2e-19
C3553 D[1] a_9754_3239# 8.74e-20
C3554 a_6759_3213# check[0] 1.67e-20
C3555 check[3] a_10776_4086# 1.93e-20
C3556 a_12031_4775# a_12548_4112# 4.23e-19
C3557 VDD a_11494_5083# 0.00984f
C3558 a_5844_3239# a_6759_3213# 0.126f
C3559 comparator_out a_6291_3605# 0.00113f
C3560 x77.Y a_4925_2550# 0.00196f
C3561 check[2] a_7247_4775# 2.07e-19
C3562 a_11288_2648# VDD 0.00506f
C3563 a_8696_2366# a_9172_2366# 2.87e-21
C3564 x77.Y a_4585_3239# 0.00397f
C3565 a_6410_2366# check[5] 1.31e-19
C3566 a_5845_4801# a_6466_4775# 0.117f
C3567 a_6546_2340# check[0] 0.00104f
C3568 x77.Y a_3505_4086# 7.15e-21
C3569 comparator_out a_6304_2366# 0.00689f
C3570 check[1] a_9173_4112# 1.03e-21
C3571 a_11970_4112# a_12030_3213# 4.45e-20
C3572 check[2] a_9442_4086# 7.66e-19
C3573 sel_bit[0] a_1227_4801# 2.06e-20
C3574 x27.D a_3900_5167# 8.53e-19
C3575 VDD a_10681_4086# 0.189f
C3576 a_2533_2550# D[6] 0.00108f
C3577 a_10775_2340# a_11288_2648# 0.00945f
C3578 a_4925_2550# check[6] 9.23e-19
C3579 a_11970_4112# x4.X 0.00309f
C3580 VDD a_9370_4801# 0.00445f
C3581 a_10628_3239# x33.Q_N 8.92e-20
C3582 a_9369_3239# x33.Q_N 4.04e-19
C3583 a_3452_3239# x48.Q 8.21e-19
C3584 x77.Y x45.Q_N 1.27e-22
C3585 a_3452_3239# a_6010_3239# 2.9e-21
C3586 x75.Q a_5845_4801# 1.99e-20
C3587 comparator_out a_621_4112# 1.4e-20
C3588 x4.X a_9656_4394# 8.47e-19
C3589 x5.X a_4368_4775# 4.59e-19
C3590 a_7764_4112# x42.Q_N 5.48e-20
C3591 a_8384_4086# a_8939_4086# 0.197f
C3592 D[1] x5.X 0.00133f
C3593 a_8236_3239# a_8289_4086# 5.06e-19
C3594 a_3453_4801# a_6199_4801# 3.65e-21
C3595 a_4681_4801# a_6011_4801# 3.02e-20
C3596 a_10680_2340# a_10776_4086# 2.97e-20
C3597 a_7246_3213# x42.Q_N 3.76e-21
C3598 a_10775_2340# a_10681_4086# 1.57e-20
C3599 a_4452_2640# a_4453_2340# 0.781f
C3600 a_3912_2366# a_4925_2550# 0.0633f
C3601 a_7246_3213# a_8402_3239# 1.84e-19
C3602 x5.X a_11544_4775# 0.00155f
C3603 a_4154_2340# a_4657_2340# 0.00187f
C3604 a_1520_2366# x20.Q_N 0.0983f
C3605 a_7072_3239# a_8236_3239# 6.38e-20
C3606 a_6759_3213# a_8857_3213# 4.53e-20
C3607 a_3599_2340# x54.Q_N 0.124f
C3608 a_6198_3239# a_6399_3239# 3.67e-19
C3609 a_7072_3239# a_6977_3239# 0.00276f
C3610 a_7246_3213# a_7480_3521# 0.00945f
C3611 a_6759_3213# x72.Q_N 0.00553f
C3612 a_8237_4801# a_8591_4801# 0.0664f
C3613 a_9376_2366# x33.Q_N 0.00473f
C3614 a_8403_4801# a_9465_4801# 0.137f
C3615 a_8684_5167# a_9152_4775# 0.0633f
C3616 x36.Q_N x39.Q_N 0.00386f
C3617 a_11857_4801# a_11966_4801# 0.00707f
C3618 comparator_out check[0] 0.121f
C3619 a_5844_3239# comparator_out 0.147f
C3620 x48.Q a_4872_4394# 1.99e-19
C3621 a_3599_2340# a_3600_4086# 5.27e-19
C3622 check[6] x45.Q_N 6.19e-19
C3623 a_2853_5648# check[1] 0.0514f
C3624 x48.Q a_4586_4801# 3.31e-19
C3625 a_10345_3239# a_9238_4086# 4.72e-19
C3626 check[2] sel_bit[0] 0.0781f
C3627 D[5] a_6546_2340# 2.03e-19
C3628 a_7246_3213# a_7185_2366# 1.2e-20
C3629 a_4154_2340# VDD 0.182f
C3630 D[7] a_1207_2340# 0.00629f
C3631 a_1112_2340# a_1520_2366# 6.04e-19
C3632 clk_sar sel_bit[0] 0.343f
C3633 a_11088_2366# check[3] 1.09e-20
C3634 a_4367_3213# a_4454_4086# 1.61e-19
C3635 a_4854_3213# a_4453_4386# 3.78e-19
C3636 a_4538_3521# VDD 0.0174f
C3637 sel_bit[1] a_1976_4775# 8.83e-20
C3638 check[2] a_10156_4112# 0.165f
C3639 x5.X a_8897_4394# 5.64e-19
C3640 a_5896_2340# a_5897_4086# 1.07e-20
C3641 x4.X x30.Q_N 0.426f
C3642 a_3453_4801# a_4539_5083# 0.00907f
C3643 a_3619_4801# a_4318_5083# 2.46e-19
C3644 a_7561_2732# a_7763_2366# 8.94e-19
C3645 a_7263_2648# VDD 0.00984f
C3646 x20.Q_N a_2398_4801# 9.16e-20
C3647 x5.X a_7363_4801# 2.04e-19
C3648 a_4388_2366# x27.Q_N 9.43e-19
C3649 a_6304_2366# a_8696_2366# 5.35e-21
C3650 check[1] a_3671_5674# 5.38e-19
C3651 a_10628_3239# a_10794_3239# 0.782f
C3652 a_6546_2340# a_8383_2340# 1.86e-21
C3653 a_2853_5648# a_3877_5674# 8.24e-20
C3654 a_6844_2640# a_7185_2366# 0.00118f
C3655 a_6845_2340# a_6984_2366# 2.56e-19
C3656 a_11630_4086# a_12102_4296# 0.15f
C3657 a_11629_4386# x39.Q_N 0.00118f
C3658 a_3806_3239# x4.X 0.00861f
C3659 a_9872_3521# a_10628_3239# 4.06e-20
C3660 a_7247_4775# a_8591_4801# 8.26e-21
C3661 check[1] a_6846_4086# 0.441f
C3662 comparator_out a_2061_2340# 0.188f
C3663 a_10795_4801# a_11494_5083# 2.46e-19
C3664 a_9376_2366# check[1] 3.33e-19
C3665 a_10629_4801# a_11715_5083# 0.00907f
C3666 x77.Y a_6198_3239# 1.34e-20
C3667 VDD a_2993_5674# 4.34e-19
C3668 a_6780_2732# x4.X 4.32e-19
C3669 a_4155_4086# a_4794_4112# 0.00316f
C3670 a_4926_4296# a_5372_4112# 0.0367f
C3671 a_4453_4386# a_4593_4112# 0.00126f
C3672 check[2] check[6] 7.32e-20
C3673 a_9322_3521# x4.X 9.99e-19
C3674 a_8939_4086# a_9173_4478# 0.00976f
C3675 VDD a_6845_4386# 0.59f
C3676 a_8384_4086# a_8803_4112# 0.0397f
C3677 a_6410_2366# x45.Q_N 4.18e-20
C3678 a_8697_4112# a_9375_4478# 0.00652f
C3679 x27.Q_N a_4926_4296# 5.7e-19
C3680 a_8696_2366# a_8802_2366# 0.0552f
C3681 a_8938_2340# a_9374_2732# 0.00412f
C3682 D[4] a_9172_2366# 3.13e-20
C3683 a_9237_2340# a_8896_2648# 1.25e-19
C3684 a_9236_2640# a_9172_2732# 2.13e-19
C3685 sel_bit[0] a_4074_4775# 0.00112f
C3686 a_5991_2340# check[5] 2.6e-20
C3687 a_9465_4801# a_9710_4296# 3.59e-20
C3688 a_9151_3213# a_8858_4775# 7.57e-21
C3689 a_9464_3239# a_8237_4801# 4.76e-21
C3690 a_9754_3239# a_9709_2550# 1.01e-20
C3691 a_3373_5674# x4.X 5.96e-20
C3692 sel_bit[0] x20.Q_N 2.7e-20
C3693 eob a_1508_5167# 0.0514f
C3694 comparator_out D[5] 0.00123f
C3695 comparator_out a_8857_3213# 4.83e-19
C3696 x4.X a_5992_4086# 0.1f
C3697 x77.Y a_4074_4775# 5.16e-21
C3698 comparator_out x72.Q_N 1.49e-19
C3699 x77.Y x20.Q_N 0.0156f
C3700 a_6845_4386# a_7318_4296# 0.155f
C3701 a_6547_4086# x45.Q_N 0.0285f
C3702 a_6846_4086# a_7050_4086# 0.117f
C3703 a_1508_5167# x4.A 0.00373f
C3704 check[0] a_4591_4478# 1.2e-20
C3705 x5.X a_6606_4801# 9.34e-19
C3706 a_2061_2340# a_2265_2340# 0.117f
C3707 a_2060_2640# a_2533_2550# 0.155f
C3708 a_9376_2366# a_9577_2366# 3.34e-19
C3709 a_1762_2340# x51.Q_N 9.58e-21
C3710 a_10680_2340# a_11088_2366# 6.04e-19
C3711 a_5845_4801# a_7481_5083# 1.25e-19
C3712 a_6011_4801# a_6978_4801# 0.00126f
C3713 D[2] a_12101_2550# 2.21e-19
C3714 a_6760_4775# a_7159_5167# 0.00133f
C3715 a_6292_5167# a_6606_4801# 0.0258f
C3716 a_1338_5674# a_2853_5648# 5.64e-20
C3717 comparator_out a_8383_2340# 0.00434f
C3718 a_9873_5083# a_10629_4801# 4.06e-20
C3719 a_4074_4775# check[6] 4.81e-21
C3720 a_6010_3239# D[0] 5.69e-21
C3721 x5.X a_10346_4801# 0.0293f
C3722 D[6] a_4925_2550# 6.65e-20
C3723 eob x4.X 0.22f
C3724 a_12102_4296# a_12346_4478# 0.00972f
C3725 a_11834_4086# a_12548_4112# 6.99e-20
C3726 a_12101_2550# a_11969_2366# 0.0258f
C3727 a_11856_3239# x39.Q_N 0.162f
C3728 check[5] a_8858_4775# 6.94e-19
C3729 comparator_out a_11766_2732# 9.47e-19
C3730 check[2] a_2788_5674# 0.00675f
C3731 a_4073_3213# a_4018_2366# 5.71e-21
C3732 a_11250_4775# check[3] 0.00109f
C3733 a_6759_3213# check[1] 2.39e-20
C3734 x4.X x4.A 0.00766f
C3735 a_4680_3239# a_4789_3239# 0.00707f
C3736 x5.X a_5897_4086# 0.0764f
C3737 a_4453_4386# a_5170_4112# 0.0019f
C3738 x48.Q a_3600_4086# 0.00969f
C3739 VDD a_7264_4394# 0.00984f
C3740 a_10680_2340# check[2] 0.027f
C3741 a_4367_3213# x75.Q 3.3e-19
C3742 a_12737_3239# x5.X 0.00125f
C3743 a_4854_3213# a_5561_3239# 0.0968f
C3744 a_9638_3213# a_9710_4296# 3.74e-20
C3745 a_6291_3605# VDD 0.176f
C3746 a_9151_3213# x42.Q_N 0.0983f
C3747 a_9464_3239# a_9442_4086# 4.33e-20
C3748 a_4925_2550# a_5991_2340# 7.98e-21
C3749 a_8857_3213# a_8683_3605# 0.205f
C3750 a_8236_3239# a_9638_3213# 0.0492f
C3751 a_8402_3239# a_9151_3213# 0.139f
C3752 a_4453_2340# a_6546_2340# 6.38e-20
C3753 a_4657_2340# a_6304_2366# 1.32e-20
C3754 a_3912_2366# x20.Q_N 1.17e-19
C3755 x27.Q_N a_6760_4775# 6.16e-21
C3756 a_11629_2340# x39.Q_N 3.65e-20
C3757 a_12101_2550# a_11834_4086# 2.22e-22
C3758 x57.Q_N x30.Q_N 4.08e-19
C3759 a_2853_5648# a_3453_4801# 7.76e-20
C3760 a_9465_4801# a_9370_4801# 0.00276f
C3761 a_8591_4801# a_8792_4801# 3.67e-19
C3762 a_9152_4775# x33.Q_N 0.0059f
C3763 a_9639_4775# a_9873_5083# 0.00945f
C3764 a_4854_3213# a_4681_4801# 4.82e-21
C3765 x4.X a_6781_4478# 2.12e-19
C3766 a_4680_3239# a_4855_4775# 1.33e-23
C3767 x66.Q_N check[3] 0.00297f
C3768 x48.Q a_1682_4775# 4.88e-21
C3769 comparator_out x33.Q_N 0.263f
C3770 a_6845_4386# a_8289_4086# 4.36e-19
C3771 a_7050_4086# a_7562_4478# 6.69e-20
C3772 a_6547_4086# a_6781_4112# 0.00707f
C3773 a_6305_4112# a_6985_4112# 3.73e-19
C3774 x45.Q_N a_6411_4112# 0.0455f
C3775 a_6846_4086# a_7764_4112# 0.0664f
C3776 a_1822_4801# a_1511_4112# 1.33e-19
C3777 a_7246_3213# a_6846_4086# 7.94e-19
C3778 a_6465_3213# x45.Q_N 0.194f
C3779 a_6759_3213# a_7050_4086# 0.0014f
C3780 a_9709_2550# a_9237_4386# 6.45e-21
C3781 a_8938_2340# x42.Q_N 0.00179f
C3782 a_4018_2366# x27.Q_N 0.0102f
C3783 a_6845_2340# a_7263_2648# 0.00276f
C3784 a_6304_2366# D[4] 1.86e-20
C3785 a_6844_2640# a_7561_2732# 4.45e-20
C3786 VDD a_1822_4801# 0.00544f
C3787 a_9236_2640# a_9710_4296# 6.02e-22
C3788 a_6304_2366# VDD 0.348f
C3789 a_8683_3605# a_8383_2340# 3.9e-20
C3790 a_8236_3239# a_9236_2640# 6.01e-20
C3791 a_8857_3213# a_8696_2366# 0.0014f
C3792 a_10628_3239# a_10629_4801# 6.9e-19
C3793 check[4] a_10983_4801# 0.164f
C3794 a_1682_4775# a_2147_5083# 9.46e-19
C3795 a_1227_4801# a_2375_5167# 2.13e-19
C3796 a_1061_4801# a_1822_4801# 6.04e-20
C3797 a_4855_4775# a_4794_4112# 1.79e-20
C3798 a_3913_4112# x48.Q_N 0.00553f
C3799 a_4453_4386# a_4658_4086# 0.153f
C3800 x5.X a_11630_4086# 0.26f
C3801 a_6844_2640# a_6846_4086# 7.02e-19
C3802 a_5991_2340# x45.Q_N 2.01e-19
C3803 a_6845_2340# a_6845_4386# 7.25e-19
C3804 x57.Q_N a_5992_4086# 2.32e-20
C3805 x77.Y a_3618_3239# 0.528f
C3806 D[4] a_8802_2366# 5.38e-19
C3807 a_621_4112# a_1511_4112# 2.76e-19
C3808 a_8802_2366# VDD 4.84e-19
C3809 check[5] x42.Q_N 6.88e-19
C3810 a_8383_2340# a_8696_2366# 0.273f
C3811 a_11389_3239# VDD 5.47e-21
C3812 a_8402_3239# check[5] 1.82e-19
C3813 a_11249_3213# a_11389_3239# 0.07f
C3814 a_10628_3239# a_11761_3239# 2.56e-19
C3815 a_10794_3239# a_11183_3239# 0.0019f
C3816 a_11543_3213# a_11714_3521# 0.00652f
C3817 VDD a_621_4112# 0.255f
C3818 x30.Q_N a_7363_4801# 0.00129f
C3819 comparator_out a_4453_2340# 0.181f
C3820 x4.X x48.Q_N 0.00819f
C3821 a_8896_2648# x4.X 0.00102f
C3822 a_11493_3521# x4.X 2.91e-19
C3823 comparator_out check[1] 0.134f
C3824 a_1976_4775# x27.D 0.00388f
C3825 a_1207_2340# a_1720_2648# 0.00945f
C3826 a_2463_4775# a_3170_4801# 0.0968f
C3827 a_9237_4386# a_11630_4086# 2.9e-21
C3828 x42.Q_N a_10776_4086# 7.84e-21
C3829 D[3] a_10680_2340# 0.0999f
C3830 check[6] a_6931_5083# 1.5e-21
C3831 VDD a_8684_5167# 0.317f
C3832 a_7185_2366# check[5] 4.92e-19
C3833 VDD check[0] 0.685f
C3834 a_11389_3239# a_10775_2340# 4.6e-20
C3835 a_8683_3605# x33.Q_N 0.00192f
C3836 a_5844_3239# VDD 0.791f
C3837 comparator_out a_7763_2366# 0.155f
C3838 comparator_out a_10794_3239# 0.148f
C3839 a_3618_3239# check[6] 7.95e-22
C3840 a_6411_4112# a_6781_4112# 4.11e-20
C3841 a_7562_4478# a_7764_4112# 8.94e-19
C3842 x4.X a_8237_4801# 0.0043f
C3843 x5.X a_2463_4775# 0.016f
C3844 check[0] a_7318_4296# 4.24e-20
C3845 a_6465_3213# a_6198_3239# 6.99e-20
C3846 a_6010_3239# a_6375_3605# 4.45e-20
C3847 a_6759_3213# a_7246_3213# 0.273f
C3848 comparator_out a_7050_4086# 4.39e-21
C3849 a_6606_4801# x30.Q_N 1.33e-19
C3850 a_11857_4801# a_12102_4296# 3.59e-20
C3851 a_8696_2366# x33.Q_N 0.0928f
C3852 a_4073_3213# a_3599_2340# 2.5e-19
C3853 a_3618_3239# a_3912_2366# 5.94e-19
C3854 x33.Q_N a_11390_4801# 6.84e-20
C3855 x5.X a_4453_4386# 0.009f
C3856 x48.Q a_3900_5167# 0.00702f
C3857 a_2061_2340# a_1511_4112# 0.00155f
C3858 a_3899_3605# a_3806_3239# 0.0367f
C3859 a_3452_3239# a_4538_3521# 0.00907f
C3860 a_4073_3213# a_3983_3605# 6.69e-20
C3861 a_3618_3239# a_4317_3521# 2.46e-19
C3862 a_4367_3213# a_4680_3239# 0.124f
C3863 a_7953_3239# a_8402_3239# 3.93e-19
C3864 a_5089_5083# check[6] 5.84e-21
C3865 D[0] a_8236_3239# 0.348f
C3866 D[6] x20.Q_N 0.00261f
C3867 x27.Q_N a_5562_4801# 0.182f
C3868 a_2061_2340# VDD 0.853f
C3869 a_4925_2550# a_5371_2366# 0.0367f
C3870 a_7072_3239# a_6304_2366# 2.17e-19
C3871 a_6759_3213# a_6844_2640# 5.32e-19
C3872 VDD a_6376_5167# 0.0042f
C3873 a_6198_3239# a_5991_2340# 2.02e-19
C3874 a_6977_3239# D[0] 1.36e-20
C3875 a_11194_2366# x33.Q_N 8.7e-20
C3876 a_8683_3605# check[1] 8.21e-20
C3877 a_12346_4112# a_11629_4386# 0.0019f
C3878 a_11970_4112# a_11630_4086# 6.04e-20
C3879 a_11769_4112# a_11834_4086# 9.75e-19
C3880 x36.Q_N a_12738_4801# 0.184f
C3881 a_12265_5083# check[3] 0.0011f
C3882 a_1520_2366# x4.X 0.112f
C3883 x4.X a_7247_4775# 0.103f
C3884 a_6606_4801# a_5992_4086# 1.08e-19
C3885 a_1976_4775# a_2579_4801# 0.0551f
C3886 check[2] a_8858_4775# 5.69e-19
C3887 a_10681_4086# a_11089_4112# 4.37e-19
C3888 a_9377_4112# a_9578_4112# 3.34e-19
C3889 D[5] VDD 0.221f
C3890 a_8857_3213# VDD 0.308f
C3891 a_3599_2340# x27.Q_N 0.142f
C3892 a_9151_3213# a_10628_3239# 3.41e-19
C3893 a_6304_2366# a_6845_2340# 0.125f
C3894 a_6546_2340# a_6844_2640# 0.137f
C3895 x72.Q_N VDD 0.0716f
C3896 a_9151_3213# a_9369_3239# 3.73e-19
C3897 a_9464_3239# a_8997_3239# 0.00316f
C3898 a_12547_2366# check[3] 0.00323f
C3899 a_8696_2366# check[1] 0.0033f
C3900 x4.X a_9442_4086# 0.00986f
C3901 a_4871_2648# x4.X 2.86e-19
C3902 VDD a_4389_4478# 0.00402f
C3903 a_6399_3239# x4.X 6.32e-19
C3904 a_4681_4801# a_4658_4086# 2.59e-19
C3905 a_4855_4775# a_4926_4296# 2.97e-21
C3906 a_8402_3239# x45.Q_N 9.58e-19
C3907 D[4] a_8383_2340# 0.0132f
C3908 VDD a_4767_5167# 0.00394f
C3909 a_7480_3521# x45.Q_N 2.75e-19
C3910 a_8383_2340# VDD 0.561f
C3911 a_7763_2366# a_8696_2366# 3.42e-20
C3912 sel_bit[0] a_1508_5167# 3.52e-20
C3913 check[3] a_11331_4086# 4.58e-20
C3914 comparator_out a_7764_4112# 4.77e-20
C3915 a_2883_5674# a_3258_5648# 0.014f
C3916 VDD a_11943_5167# 0.00371f
C3917 a_2883_5674# sel_bit[1] 0.0353f
C3918 comparator_out a_7246_3213# 0.00381f
C3919 a_5844_3239# a_7072_3239# 0.0334f
C3920 check[1] a_7954_4801# 0.0169f
C3921 a_4389_4112# a_4794_4112# 2.46e-21
C3922 a_5897_4086# a_5992_4086# 0.0968f
C3923 x4.X a_2398_4801# 0.00124f
C3924 x5.X a_6011_4801# 0.0199f
C3925 x4.X a_9574_4801# 2.39e-19
C3926 a_7185_2366# x45.Q_N 5.33e-22
C3927 a_11766_2732# VDD 0.0163f
C3928 a_5845_4801# a_6760_4775# 0.125f
C3929 a_6011_4801# a_6292_5167# 0.155f
C3930 sel_bit[0] a_3913_4112# 5.05e-19
C3931 x77.Y x75.Q_N 3.94e-19
C3932 a_9237_2340# a_10680_2340# 8.18e-19
C3933 a_8938_2340# a_9376_2366# 0.00276f
C3934 check[0] a_3619_4801# 0.00149f
C3935 a_8696_2366# a_9577_2366# 0.00943f
C3936 x5.X a_11966_4801# 5.38e-20
C3937 a_6845_2340# check[0] 1.9e-19
C3938 a_11389_3239# a_11965_3239# 2.46e-21
C3939 x77.Y a_3913_4112# 3.94e-20
C3940 a_9152_4775# a_10629_4801# 1.67e-19
C3941 check[1] a_9578_4112# 3.76e-20
C3942 comparator_out a_6844_2640# 0.108f
C3943 a_5844_3239# a_6845_2340# 6.52e-20
C3944 check[2] x42.Q_N 8.18e-19
C3945 x5.X a_8697_4112# 0.00599f
C3946 sel_bit[0] x4.X 6.44e-20
C3947 check[5] a_6846_4086# 0.0346f
C3948 a_1626_2366# a_1996_2366# 4.11e-20
C3949 x27.D a_4855_4775# 4.69e-21
C3950 a_7247_4775# a_7186_4112# 1.79e-20
C3951 VDD a_9377_4112# 0.00445f
C3952 a_11088_2366# a_11564_2732# 0.00133f
C3953 a_10628_3239# a_10776_4086# 8.29e-19
C3954 x77.Y x4.X 0.07f
C3955 check[4] x39.Q_N 6.54e-19
C3956 VDD x33.Q_N 0.446f
C3957 D[4] x33.Q_N 0.00278f
C3958 a_5561_3239# x5.X 0.00125f
C3959 x69.Q_N x33.Q_N 0.02f
C3960 comparator_out a_9953_2732# 8.29e-19
C3961 x75.Q_N check[6] 0.00302f
C3962 x4.X a_10156_4112# 0.00621f
C3963 x5.X a_4681_4801# 1.74e-19
C3964 a_8697_4112# a_9237_4386# 0.139f
C3965 a_8384_4086# a_9238_4086# 0.0492f
C3966 check[6] a_3913_4112# 7.75e-22
C3967 x4.X a_8792_4801# 8.46e-20
C3968 a_1062_5674# a_897_4112# 9.53e-20
C3969 a_2060_2640# x20.Q_N 0.351f
C3970 D[2] x39.Q_N 0.00168f
C3971 a_4453_2340# a_4657_2340# 0.117f
C3972 x5.X a_11857_4801# 0.00141f
C3973 a_4452_2640# a_4925_2550# 0.145f
C3974 a_7246_3213# a_8683_3605# 7.98e-21
C3975 a_4154_2340# x54.Q_N 9.58e-21
C3976 a_6759_3213# a_9151_3213# 3.6e-20
C3977 a_7072_3239# x72.Q_N 9.58e-21
C3978 a_9152_4775# a_9639_4775# 0.273f
C3979 a_8858_4775# a_8591_4801# 6.99e-20
C3980 a_8403_4801# a_8768_5167# 4.45e-20
C3981 a_12030_3213# check[3] 0.00748f
C3982 a_10775_2340# x33.Q_N 1.5e-19
C3983 x4.X check[6] 0.0328f
C3984 a_3599_2340# a_4155_4086# 1.3e-22
C3985 a_3912_2366# a_3913_4112# 1.8e-19
C3986 a_8383_2340# a_8289_4086# 1.57e-20
C3987 x4.X check[3] 0.316f
C3988 a_8288_2340# a_8384_4086# 2.97e-20
C3989 a_2979_2366# x27.Q_N 1.34e-20
C3990 D[5] a_6845_2340# 1.11e-19
C3991 a_6010_3239# x27.Q_N 7.07e-20
C3992 a_8236_3239# a_10345_3239# 1.03e-19
C3993 a_4453_2340# VDD 0.788f
C3994 a_1112_2340# a_2060_2640# 7.7e-21
C3995 a_11969_2366# x39.Q_N 5.33e-22
C3996 D[7] a_1762_2340# 8.38e-19
C3997 D[0] a_8791_3239# 1.27e-19
C3998 check[1] a_1511_4112# 5.91e-22
C3999 a_4367_3213# a_4926_4296# 1.71e-19
C4000 a_4854_3213# a_4658_4086# 2.47e-19
C4001 a_11628_2640# check[3] 0.0274f
C4002 D[4] check[1] 0.194f
C4003 VDD check[1] 0.762f
C4004 a_4213_3239# VDD 0.00187f
C4005 sel_bit[1] a_2289_4801# 1.47e-20
C4006 a_3912_2366# x4.X 0.105f
C4007 x20.Q_N a_4113_4394# 6.16e-20
C4008 x5.X a_9375_4478# 7.3e-19
C4009 check[2] a_9173_4112# 1.17e-20
C4010 a_7953_3239# a_6846_4086# 4.72e-19
C4011 a_4074_4775# a_4539_5083# 9.46e-19
C4012 a_3619_4801# a_4767_5167# 2.13e-19
C4013 a_3453_4801# a_4214_4801# 6.04e-20
C4014 a_7763_2366# VDD 0.109f
C4015 a_10794_3239# VDD 0.274f
C4016 a_11834_4086# x39.Q_N 0.00118f
C4017 a_4793_2366# x27.Q_N 0.0404f
C4018 x5.X a_9102_5083# 3.46e-19
C4019 check[2] a_9873_5083# 4.31e-19
C4020 a_10794_3239# a_11249_3213# 0.153f
C4021 a_7246_3213# a_7954_4801# 3.19e-20
C4022 a_10628_3239# a_11075_3605# 0.15f
C4023 a_6845_2340# a_8383_2340# 0.00116f
C4024 a_6844_2640# a_8696_2366# 1.79e-19
C4025 a_7049_2340# a_7185_2366# 0.07f
C4026 a_6759_3213# check[5] 1.11e-19
C4027 a_4317_3521# x4.X 0.00111f
C4028 a_9872_3521# VDD 0.00506f
C4029 a_7247_4775# a_7363_4801# 0.0397f
C4030 a_6760_4775# a_7182_4801# 2.87e-21
C4031 x69.Q_N a_10794_3239# 8.64e-20
C4032 check[1] a_7318_4296# 0.0013f
C4033 a_1996_2732# eob 4.16e-20
C4034 a_9872_3521# x69.Q_N 2.02e-20
C4035 comparator_out a_2533_2550# 0.00698f
C4036 a_11250_4775# a_11715_5083# 9.46e-19
C4037 a_10629_4801# a_11390_4801# 6.04e-20
C4038 a_10795_4801# a_11943_5167# 2.13e-19
C4039 a_6410_2366# x4.X 3.78e-20
C4040 a_3452_3239# check[0] 2.98e-21
C4041 x77.Y a_4970_3239# 0.00967f
C4042 a_4454_4086# a_4794_4112# 6.04e-20
C4043 a_4658_4086# a_4593_4112# 9.75e-19
C4044 VDD a_3877_5674# 3.02e-19
C4045 a_4453_4386# a_5992_4086# 1.24e-19
C4046 a_8997_3239# x4.X 0.00265f
C4047 a_3452_3239# a_5844_3239# 0.00176f
C4048 a_8939_4086# a_8803_4112# 0.0282f
C4049 a_9237_4386# a_9375_4478# 1.09e-19
C4050 a_8697_4112# a_9656_4394# 1.21e-20
C4051 VDD a_7050_4086# 0.487f
C4052 x5.X a_897_4112# 0.00452f
C4053 a_5562_4801# a_5845_4801# 8.18e-19
C4054 D[4] a_9577_2366# 7.47e-20
C4055 a_9237_2340# a_9374_2732# 0.00907f
C4056 a_8998_4801# a_8384_4086# 1.08e-19
C4057 a_10628_3239# a_11088_2366# 1.89e-19
C4058 a_6546_2340# check[5] 1.34e-19
C4059 a_10794_3239# a_10775_2340# 3.73e-19
C4060 a_9151_3213# a_9152_4775# 0.00121f
C4061 a_8237_4801# a_10346_4801# 1.03e-19
C4062 eob a_2463_4775# 0.00567f
C4063 comparator_out a_9151_3213# 7.47e-19
C4064 x4.X a_6547_4086# 0.00727f
C4065 a_10680_2340# x4.X 0.00342f
C4066 a_7050_4086# a_7318_4296# 0.205f
C4067 a_6846_4086# x45.Q_N 0.00113f
C4068 check[0] a_4872_4394# 8.58e-21
C4069 x5.X a_6978_4801# 2.58e-19
C4070 a_2265_2340# a_2533_2550# 0.205f
C4071 a_10680_2340# a_11628_2640# 9.65e-21
C4072 a_2061_2340# x51.Q_N 1.07e-19
C4073 a_7073_4801# a_7159_5167# 0.00976f
C4074 a_4971_4801# a_4790_4801# 4.11e-20
C4075 a_6011_4801# x30.Q_N 1.04e-19
C4076 a_2389_5648# check[1] 0.0168f
C4077 a_6845_2340# x33.Q_N 1.52e-19
C4078 check[2] a_2853_5648# 0.112f
C4079 comparator_out a_8938_2340# 0.00103f
C4080 x33.Q_N a_10795_4801# 2.19e-19
C4081 comparator_out x3.A 2e-20
C4082 a_10628_3239# check[2] 0.0451f
C4083 VDD a_1338_5674# 0.255f
C4084 x48.Q a_1976_4775# 4.67e-19
C4085 a_11565_4112# a_11970_4112# 2.46e-21
C4086 a_4368_4775# check[6] 0.00421f
C4087 a_4855_4775# a_5562_4801# 0.0968f
C4088 x39.Q_N a_12548_4112# 8.27e-20
C4089 a_6759_3213# a_7953_3239# 6.04e-19
C4090 a_6291_3605# D[0] 3.23e-21
C4091 a_11159_3605# x39.Q_N 8.48e-19
C4092 check[5] a_9152_4775# 0.00306f
C4093 a_10155_2366# x33.Q_N 0.032f
C4094 check[1] a_8289_4086# 0.125f
C4095 comparator_out a_12047_2648# 6.95e-19
C4096 comparator_out check[5] 0.0221f
C4097 check[2] a_3671_5674# 0.00323f
C4098 a_1338_5674# a_1061_4801# 0.00179f
C4099 a_12031_4775# a_12738_4801# 0.0968f
C4100 a_11544_4775# check[3] 0.00913f
C4101 check[2] a_6846_4086# 2.36e-20
C4102 x48.Q a_4155_4086# 0.00101f
C4103 a_6011_4801# a_5992_4086# 6.63e-19
C4104 a_5845_4801# a_6305_4112# 3.05e-19
C4105 VDD a_7764_4112# 0.109f
C4106 a_1976_4775# a_2147_5083# 0.00652f
C4107 a_9464_3239# x42.Q_N 0.162f
C4108 sel_bit[1] reset 1.45e-20
C4109 D[0] a_6304_2366# 1.92e-21
C4110 a_7246_3213# VDD 0.569f
C4111 a_9639_4775# a_9578_4112# 1.79e-20
C4112 a_8402_3239# a_9464_3239# 0.137f
C4113 a_4453_2340# a_6845_2340# 0.00176f
C4114 a_8236_3239# a_8590_3239# 0.0708f
C4115 check[4] a_9238_4086# 0.0367f
C4116 x27.Q_N a_7073_4801# 7.65e-21
C4117 a_3912_2366# x57.Q_N 8.28e-21
C4118 a_4214_4801# a_4790_4801# 2.46e-21
C4119 a_8683_3605# a_9151_3213# 0.0633f
C4120 a_12101_2550# x39.Q_N 0.00196f
C4121 comparator_out a_10776_4086# 0.00196f
C4122 check[1] a_3619_4801# 7.46e-20
C4123 a_2853_5648# a_4074_4775# 1.12e-19
C4124 a_9465_4801# x33.Q_N 8.55e-20
C4125 a_2853_5648# x20.Q_N 2.38e-20
C4126 a_6845_2340# check[1] 6.25e-19
C4127 x4.X a_6411_4112# 0.00336f
C4128 D[6] x4.X 0.00589f
C4129 a_6465_3213# x4.X 0.00499f
C4130 a_6845_4386# a_6985_4112# 0.00126f
C4131 a_7318_4296# a_7764_4112# 0.0367f
C4132 a_6547_4086# a_7186_4112# 0.00316f
C4133 a_7072_3239# a_7050_4086# 4.33e-20
C4134 a_7246_3213# a_7318_4296# 3.74e-20
C4135 a_6759_3213# x45.Q_N 0.0983f
C4136 VDD a_3453_4801# 0.841f
C4137 a_6845_2340# a_7763_2366# 0.0708f
C4138 a_9709_2550# a_9442_4086# 2.22e-22
C4139 a_9237_2340# x42.Q_N 3.65e-20
C4140 a_6844_2640# VDD 0.269f
C4141 VDD a_2194_4801# 0.00214f
C4142 a_7049_2340# a_7561_2732# 6.69e-20
C4143 a_6844_2640# D[4] 0.00557f
C4144 a_8683_3605# a_8938_2340# 2.41e-20
C4145 a_8236_3239# a_9441_2340# 4.77e-19
C4146 a_9151_3213# a_8696_2366# 3.36e-20
C4147 a_8402_3239# a_9237_2340# 6.38e-20
C4148 a_8857_3213# a_9236_2640# 2.68e-19
C4149 a_8997_3239# D[1] 1.13e-20
C4150 check[6] a_7363_4801# 1.16e-20
C4151 a_10794_3239# a_10795_4801# 1.39e-19
C4152 VDD a_10629_4801# 0.81f
C4153 check[4] a_9755_4801# 2.75e-19
C4154 a_1061_4801# a_3453_4801# 0.00176f
C4155 a_1338_5674# a_2389_5648# 0.00356f
C4156 a_1682_4775# a_1822_4801# 0.07f
C4157 a_5991_2340# x4.X 0.111f
C4158 a_1061_4801# a_2194_4801# 2.56e-19
C4159 a_1227_4801# a_1616_4801# 0.0019f
C4160 a_4453_4386# x48.Q_N 4.82e-21
C4161 a_4454_4086# a_4926_4296# 0.15f
C4162 a_7317_2550# a_6845_4386# 6.45e-21
C4163 x5.X a_12102_4296# 1.62e-19
C4164 a_6844_2640# a_7318_4296# 6.02e-22
C4165 a_6546_2340# x45.Q_N 0.0018f
C4166 x77.Y a_3899_3605# 0.181f
C4167 a_9953_2732# VDD 0.0042f
C4168 a_6984_2366# x27.Q_N 2.64e-20
C4169 a_10628_3239# D[3] 5.2e-19
C4170 a_12146_3239# VDD 4.88e-19
C4171 D[1] a_10680_2340# 0.00635f
C4172 a_8696_2366# a_8938_2340# 0.124f
C4173 a_8288_2340# x60.Q_N 0.178f
C4174 a_8383_2340# a_9236_2640# 0.0264f
C4175 a_11761_3239# VDD 6.2e-19
C4176 a_11249_3213# a_11761_3239# 9.75e-19
C4177 a_12030_3213# a_11942_3605# 7.71e-20
C4178 a_11856_3239# a_11714_3521# 0.00412f
C4179 a_10628_3239# x66.Q_N 1.07e-19
C4180 a_11543_3213# a_11389_3239# 0.00943f
C4181 a_11075_3605# a_11183_3239# 0.00812f
C4182 a_5844_3239# D[0] 7.04e-20
C4183 comparator_out a_7953_3239# 0.00109f
C4184 comparator_out a_4925_2550# 0.0087f
C4185 a_9374_2732# x4.X 9.81e-19
C4186 a_11942_3605# x4.X 4.4e-19
C4187 a_5088_3521# a_5844_3239# 4.06e-20
C4188 sel_bit[0] a_2784_5996# 0.00164f
C4189 a_1520_2366# a_1996_2732# 0.00133f
C4190 a_8939_4086# x39.Q_N 1.36e-20
C4191 a_2289_4801# x27.D 1.17e-20
C4192 a_6010_3239# a_5845_4801# 8.16e-19
C4193 check[0] a_3600_4086# 9e-20
C4194 a_9709_2550# a_9953_2366# 0.00812f
C4195 check[6] a_6606_4801# 1.78e-19
C4196 a_8696_2366# check[5] 2.42e-20
C4197 VDD a_9639_4775# 0.72f
C4198 comparator_out a_3505_4086# 2.05e-21
C4199 a_9638_3213# x33.Q_N 0.0126f
C4200 x69.Q_N a_9639_4775# 4.45e-20
C4201 comparator_out a_11075_3605# 0.0011f
C4202 a_8998_4801# check[4] 1.23e-20
C4203 a_6845_4386# a_7562_4112# 0.0019f
C4204 x4.X a_8858_4775# 9.41e-19
C4205 x5.X a_1415_4801# 0.00367f
C4206 a_2979_2366# a_2777_2366# 3.67e-19
C4207 a_3504_2340# a_3599_2340# 0.0968f
C4208 a_1996_2366# a_2401_2366# 2.46e-21
C4209 a_6759_3213# a_6198_3239# 3.79e-20
C4210 a_7246_3213# a_7072_3239# 0.197f
C4211 a_6291_3605# a_6375_3605# 0.00972f
C4212 a_2061_2340# x54.Q_N 2.94e-19
C4213 a_7954_4801# check[5] 0.129f
C4214 comparator_out x45.Q_N 0.00129f
C4215 a_9236_2640# x33.Q_N 0.572f
C4216 a_6978_4801# x30.Q_N 1.41e-19
C4217 a_11390_4801# a_10776_4086# 1.08e-19
C4218 a_4073_3213# a_4154_2340# 4.18e-20
C4219 a_4367_3213# a_3599_2340# 9.06e-19
C4220 a_3452_3239# a_4453_2340# 6.52e-20
C4221 comparator_out a_11088_2366# 0.00716f
C4222 a_3618_3239# a_4452_2640# 4.04e-20
C4223 a_3899_3605# a_3912_2366# 1.71e-19
C4224 x33.Q_N a_11762_4801# 3.57e-20
C4225 check[1] a_6710_5083# 1.55e-19
C4226 a_1062_5674# x5.X 0.00504f
C4227 x5.X a_4658_4086# 4.53e-19
C4228 check[6] a_5897_4086# 0.00265f
C4229 a_2533_2550# a_1511_4112# 6.53e-19
C4230 x48.Q a_4855_4775# 0.00105f
C4231 a_4073_3213# a_4538_3521# 9.46e-19
C4232 a_3618_3239# a_4766_3605# 2.13e-19
C4233 a_3452_3239# a_4213_3239# 6.04e-20
C4234 D[0] a_8857_3213# 8.87e-20
C4235 a_6759_3213# a_7049_2340# 0.00144f
C4236 a_2533_2550# VDD 0.194f
C4237 a_7072_3239# a_6844_2640# 1.11e-20
C4238 a_7246_3213# a_6845_2340# 8.72e-19
C4239 VDD a_4790_4801# 9.01e-19
C4240 x72.Q_N D[0] 2.5e-19
C4241 a_7181_3239# x30.Q_N 1.68e-19
C4242 a_12737_3239# check[3] 0.0275f
C4243 a_11970_4112# a_12102_4296# 0.0258f
C4244 a_11769_4112# x39.Q_N 0.00167f
C4245 a_2060_2640# x4.X 0.00821f
C4246 x4.X a_6199_4801# 2.3e-19
C4247 a_3453_4801# a_3619_4801# 0.75f
C4248 a_10156_4112# a_11630_4086# 3.65e-21
C4249 check[2] a_9152_4775# 0.00242f
C4250 a_10681_4086# a_11629_4386# 7.74e-21
C4251 a_2697_5083# a_3453_4801# 4.06e-20
C4252 a_2463_4775# a_2398_4801# 4.2e-20
C4253 a_2289_4801# a_2579_4801# 0.0282f
C4254 a_1616_4801# x20.Q_N 4.31e-20
C4255 a_9464_3239# a_10628_3239# 6.38e-20
C4256 D[0] a_8383_2340# 0.00127f
C4257 a_9638_3213# a_10794_3239# 1.69e-19
C4258 a_9151_3213# a_11249_3213# 4.53e-20
C4259 a_4154_2340# x27.Q_N 0.16f
C4260 a_9151_3213# VDD 0.353f
C4261 a_6844_2640# a_6845_2340# 0.781f
C4262 a_6304_2366# a_7317_2550# 0.0633f
C4263 a_5991_2340# x57.Q_N 0.124f
C4264 a_6011_4801# a_8237_4801# 4e-20
C4265 a_5845_4801# a_8403_4801# 2.9e-21
C4266 a_6546_2340# a_7049_2340# 0.00187f
C4267 a_8590_3239# a_8791_3239# 3.67e-19
C4268 a_9151_3213# x69.Q_N 0.00553f
C4269 a_9464_3239# a_9369_3239# 0.00276f
C4270 a_9638_3213# a_9872_3521# 0.00945f
C4271 comparator_out check[2] 0.125f
C4272 a_11768_2366# check[3] 9.26e-20
C4273 a_10629_4801# a_10795_4801# 0.751f
C4274 eob a_897_4112# 0.00374f
C4275 a_9236_2640# check[1] 3.18e-19
C4276 a_3913_4112# a_4113_4394# 0.00185f
C4277 a_3600_4086# a_4389_4478# 7.71e-20
C4278 x4.X x42.Q_N 0.252f
C4279 a_5371_2366# x4.X 8.28e-20
C4280 a_8402_3239# x4.X 0.0429f
C4281 VDD a_4019_4112# 0.0124f
C4282 a_7480_3521# x4.X 0.00103f
C4283 x5.X a_3170_4801# 0.0367f
C4284 a_897_4112# x4.A 0.238f
C4285 a_8403_4801# a_8384_4086# 6.63e-19
C4286 a_8237_4801# a_8697_4112# 3.05e-19
C4287 check[0] a_6985_4112# 3.21e-20
C4288 a_8938_2340# VDD 0.177f
C4289 D[4] a_8938_2340# 1.94e-19
C4290 a_7953_3239# a_7954_4801# 9.85e-20
C4291 VDD a_4008_4801# 2.82e-19
C4292 a_9638_3213# a_9577_2366# 1.2e-20
C4293 VDD x3.A 0.203f
C4294 a_3648_5972# a_3373_5674# 0.0156f
C4295 sel_bit[0] a_2463_4775# 5.11e-20
C4296 sel_bit[1] a_3258_5648# 0.259f
C4297 check[3] a_11630_4086# 0.223f
C4298 comparator_out a_6198_3239# 0.158f
C4299 a_1996_2366# eob 1.64e-21
C4300 a_5844_3239# a_6375_3605# 0.0018f
C4301 x4.X a_4113_4394# 1.78e-19
C4302 x5.X a_6292_5167# 0.00462f
C4303 a_9953_2732# a_10155_2366# 8.94e-19
C4304 a_12047_2648# VDD 0.00984f
C4305 D[4] check[5] 0.00424f
C4306 a_6011_4801# a_7247_4775# 0.0264f
C4307 a_5845_4801# a_7073_4801# 0.0334f
C4308 a_6466_4775# a_6760_4775# 0.199f
C4309 a_12146_3239# a_11965_3239# 4.11e-20
C4310 a_9237_2340# a_9376_2366# 2.56e-19
C4311 VDD check[5] 0.493f
C4312 check[0] a_3900_5167# 8.76e-19
C4313 a_8696_2366# a_11088_2366# 4.59e-21
C4314 a_9236_2640# a_9577_2366# 0.00118f
C4315 a_8938_2340# a_10775_2340# 1.86e-21
C4316 D[0] x33.Q_N 1.28e-20
C4317 a_7317_2550# check[0] 1.78e-19
C4318 a_9639_4775# a_10795_4801# 1.25e-19
C4319 a_9465_4801# a_10629_4801# 6.38e-20
C4320 x77.Y a_4453_4386# 1.11e-20
C4321 comparator_out x20.Q_N 0.0881f
C4322 comparator_out a_7049_2340# 0.00589f
C4323 a_12346_4112# a_12548_4112# 3.67e-19
C4324 a_11564_2732# x4.X 4.32e-19
C4325 x5.X a_9237_4386# 0.00958f
C4326 x27.D a_3807_4801# 0.164f
C4327 a_10776_4086# a_11289_4394# 0.00945f
C4328 a_10794_3239# a_11089_4112# 4.9e-19
C4329 VDD a_10776_4086# 0.716f
C4330 a_11249_3213# a_10776_4086# 2.45e-19
C4331 a_11088_2366# a_11194_2366# 0.0552f
C4332 a_11628_2640# a_11564_2732# 2.13e-19
C4333 a_11330_2340# a_11766_2732# 0.00412f
C4334 a_11629_2340# a_11288_2648# 1.25e-19
C4335 a_11543_3213# x33.Q_N 8.28e-21
C4336 comparator_out D[3] 0.00125f
C4337 comparator_out a_1112_2340# 1.42e-19
C4338 a_4367_3213# a_6010_3239# 2.89e-19
C4339 comparator_out x66.Q_N 2.08e-20
C4340 x4.X a_9173_4112# 8.4e-20
C4341 a_7186_4112# x42.Q_N 4.05e-20
C4342 a_8384_4086# a_9710_4296# 4.7e-22
C4343 a_5562_4801# a_4454_4086# 6.67e-19
C4344 check[6] a_4453_4386# 0.0318f
C4345 a_8696_2366# check[2] 1.08e-21
C4346 a_8939_4086# a_9238_4086# 0.0334f
C4347 a_8697_4112# a_9442_4086# 0.199f
C4348 a_8236_3239# a_8384_4086# 8.29e-19
C4349 a_4855_4775# a_7073_4801# 1.86e-21
C4350 a_4368_4775# a_6199_4801# 1.49e-21
C4351 a_10775_2340# a_10776_4086# 5.27e-19
C4352 a_4453_2340# x54.Q_N 1.07e-19
C4353 a_4657_2340# a_4925_2550# 0.205f
C4354 a_2265_2340# x20.Q_N 0.194f
C4355 check[0] a_7562_4112# 5.56e-22
C4356 x5.X a_11160_5167# 4.21e-19
C4357 a_5896_2340# x30.Q_N 3.7e-19
C4358 a_9639_4775# a_9465_4801# 0.197f
C4359 a_8684_5167# a_8768_5167# 0.00972f
C4360 a_9152_4775# a_8591_4801# 2.47e-21
C4361 a_8237_4801# a_9102_5083# 0.00276f
C4362 a_11330_2340# x33.Q_N 5.36e-20
C4363 a_3452_3239# a_3453_4801# 6.9e-19
C4364 D[0] check[1] 0.169f
C4365 comparator_out a_8591_4801# 1.94e-20
C4366 a_2883_5674# x48.Q 0.00144f
C4367 a_11194_2366# check[2] 0.00242f
C4368 a_3912_2366# a_4453_4386# 1.93e-22
C4369 check[2] a_7954_4801# 4.53e-20
C4370 a_7953_3239# D[4] 0.00127f
C4371 D[1] x42.Q_N 0.00176f
C4372 a_8402_3239# D[1] 5.69e-21
C4373 a_7953_3239# VDD 0.19f
C4374 D[5] a_7317_2550# 1.96e-20
C4375 D[7] a_2061_2340# 1.85e-19
C4376 a_4925_2550# VDD 0.174f
C4377 a_2853_5648# a_3913_4112# 4.72e-21
C4378 check[1] a_3600_4086# 1.19e-20
C4379 a_4213_3239# a_3600_4086# 1.16e-20
C4380 a_4680_3239# a_4926_4296# 2.37e-20
C4381 a_11833_2340# check[3] 6.99e-20
C4382 a_4585_3239# VDD 0.00112f
C4383 a_1511_4112# a_3505_4086# 0.0121f
C4384 a_4452_2640# x4.X 0.00799f
C4385 a_5896_2340# a_5992_4086# 2.97e-20
C4386 x20.Q_N a_4591_4478# 6.94e-20
C4387 check[2] a_9578_4112# 1.87e-19
C4388 a_5991_2340# a_5897_4086# 1.57e-20
C4389 x5.X a_9656_4394# 2.97e-19
C4390 VDD a_3505_4086# 0.212f
C4391 a_3619_4801# a_4008_4801# 0.0019f
C4392 a_3453_4801# a_4586_4801# 2.56e-19
C4393 check[5] a_8289_4086# 0.00275f
C4394 a_4074_4775# a_4214_4801# 0.07f
C4395 a_4368_4775# a_4539_5083# 0.00652f
C4396 VDD a_11565_4478# 0.00371f
C4397 a_7317_2550# a_8383_2340# 7.98e-21
C4398 x20.Q_N a_4214_4801# 1.27e-19
C4399 a_6304_2366# x27.Q_N 8.23e-20
C4400 a_10628_3239# a_12030_3213# 0.0492f
C4401 a_11249_3213# a_11075_3605# 0.205f
C4402 a_11075_3605# VDD 0.176f
C4403 x5.X a_9551_5167# 1.06e-19
C4404 a_10794_3239# a_11543_3213# 0.139f
C4405 a_7049_2340# a_8696_2366# 8.4e-21
C4406 a_6845_2340# a_8938_2340# 6.38e-20
C4407 a_2853_5648# x4.X 5.73e-20
C4408 a_4766_3605# x4.X 6.48e-19
C4409 a_7073_4801# a_7182_4801# 0.00707f
C4410 a_1227_4801# a_1511_4112# 0.00301f
C4411 a_11544_4775# a_11715_5083# 0.00652f
C4412 a_10795_4801# a_11184_4801# 0.0019f
C4413 a_10629_4801# a_11762_4801# 2.56e-19
C4414 a_11250_4775# a_11390_4801# 0.07f
C4415 x5.A sel_bit[1] 0.0425f
C4416 a_7561_2732# x4.X 1.17e-19
C4417 a_10628_3239# x4.X 0.0456f
C4418 VDD a_1227_4801# 0.34f
C4419 a_4453_4386# a_6547_4086# 2.47e-20
C4420 a_4454_4086# a_6305_4112# 5.07e-21
C4421 a_4926_4296# a_4794_4112# 0.0258f
C4422 a_3618_3239# comparator_out 4.91e-19
C4423 a_9369_3239# x4.X 4.91e-19
C4424 a_8697_4112# a_10156_4112# 8.23e-22
C4425 a_9237_4386# a_9656_4394# 2.46e-19
C4426 a_9442_4086# a_9375_4478# 9.46e-19
C4427 x42.Q_N a_8897_4394# 2.02e-20
C4428 x77.Y a_5561_3239# 3.29e-19
C4429 VDD x45.Q_N 0.458f
C4430 check[6] a_6011_4801# 0.162f
C4431 a_8696_2366# D[3] 1.61e-20
C4432 a_9237_2340# a_9655_2648# 0.00276f
C4433 a_11075_3605# a_10775_2340# 3.9e-20
C4434 a_9236_2640# a_9953_2732# 4.45e-20
C4435 a_11249_3213# a_11088_2366# 0.0014f
C4436 a_11088_2366# VDD 0.348f
C4437 a_10628_3239# a_11628_2640# 6.01e-20
C4438 a_6845_2340# check[5] 0.0379f
C4439 a_9638_3213# a_9639_4775# 0.00237f
C4440 a_1061_4801# a_1227_4801# 0.619f
C4441 a_8403_4801# check[4] 1.14e-20
C4442 eob a_1415_4801# 0.151f
C4443 comparator_out a_9464_3239# 1.93e-19
C4444 a_5844_3239# a_8590_3239# 3.65e-21
C4445 a_11389_3239# x36.Q_N 6.11e-19
C4446 x4.X a_6846_4086# 0.0467f
C4447 a_7318_4296# x45.Q_N 0.00243f
C4448 check[0] a_5372_4112# 0.165f
C4449 a_1520_2366# a_1996_2366# 2.87e-21
C4450 x5.X x30.Q_N 8.83e-19
C4451 D[3] a_11194_2366# 5.39e-19
C4452 a_10775_2340# a_11088_2366# 0.273f
C4453 a_10629_4801# a_11089_4112# 3.05e-19
C4454 a_6760_4775# a_7481_5083# 0.00185f
C4455 a_6292_5167# x30.Q_N 7.29e-20
C4456 a_10795_4801# a_10776_4086# 6.63e-19
C4457 a_10345_3239# x33.Q_N 0.0101f
C4458 check[0] x27.Q_N 0.0367f
C4459 a_1062_5674# eob 2.23e-21
C4460 comparator_out a_9237_2340# 0.184f
C4461 a_5844_3239# x27.Q_N 8.96e-20
C4462 a_5561_3239# check[6] 0.027f
C4463 x33.Q_N a_11076_5167# 1.6e-19
C4464 check[2] a_1511_4112# 5.19e-20
C4465 sel_bit[1] x27.D 4.45e-19
C4466 a_1062_5674# x4.A 8.16e-22
C4467 check[2] a_11289_4394# 9.25e-20
C4468 VDD check[2] 0.713f
C4469 a_3912_2366# a_4112_2648# 0.00185f
C4470 x48.Q a_2289_4801# 8.99e-20
C4471 a_3599_2340# a_4388_2732# 7.71e-20
C4472 a_4681_4801# check[6] 4.98e-20
C4473 x69.Q_N check[2] 4.68e-20
C4474 VDD clk_sar 0.114f
C4475 a_7246_3213# D[0] 0.0116f
C4476 a_4970_3239# a_4452_2640# 5.05e-21
C4477 check[5] a_9465_4801# 6.82e-20
C4478 comparator_out a_12547_2366# 0.155f
C4479 check[1] a_6985_4112# 7.78e-20
C4480 x5.X a_3373_5674# 1.23e-19
C4481 a_2389_5648# a_1227_4801# 3.08e-19
C4482 a_11857_4801# check[3] 0.00257f
C4483 x75.Q_N a_6759_3213# 2.97e-20
C4484 clk_sar a_1061_4801# 1.18e-19
C4485 x5.X a_5992_4086# 0.0202f
C4486 a_4453_4386# a_6411_4112# 9.75e-21
C4487 check[2] a_7318_4296# 2.18e-22
C4488 x48.Q a_4454_4086# 2.06e-19
C4489 a_10775_2340# check[2] 0.0128f
C4490 a_6292_5167# a_5992_4086# 4.9e-20
C4491 a_6466_4775# a_6305_4112# 0.0025f
C4492 a_5845_4801# a_6845_4386# 9.86e-20
C4493 VDD a_6781_4112# 3.56e-19
C4494 a_2463_4775# a_2375_5167# 7.71e-20
C4495 a_2289_4801# a_2147_5083# 0.00412f
C4496 a_1508_5167# a_1616_4801# 0.00812f
C4497 a_1976_4775# a_1822_4801# 0.00943f
C4498 a_7953_3239# a_6845_2340# 4.83e-19
C4499 a_8767_3605# x42.Q_N 8.48e-19
C4500 D[0] a_6844_2640# 6.76e-19
C4501 a_6198_3239# VDD 0.109f
C4502 a_9151_3213# a_9638_3213# 0.273f
C4503 a_2061_2340# x27.Q_N 1.55e-19
C4504 a_4452_2640# x57.Q_N 1.53e-19
C4505 a_8857_3213# a_8590_3239# 6.99e-20
C4506 a_8402_3239# a_8767_3605# 4.45e-20
C4507 a_8236_3239# check[4] 1.94e-20
C4508 sel_bit[0] a_897_4112# 8.65e-21
C4509 check[1] a_3900_5167# 4.17e-20
C4510 eob a_3170_4801# 0.00132f
C4511 x4.X a_7562_4478# 9.15e-19
C4512 a_6759_3213# x4.X 0.111f
C4513 a_6845_4386# a_8384_4086# 2.16e-19
C4514 x45.Q_N a_8289_4086# 8.9e-21
C4515 a_7050_4086# a_6985_4112# 9.75e-19
C4516 a_3453_4801# a_3600_4086# 0.00159f
C4517 a_6846_4086# a_7186_4112# 6.04e-20
C4518 x20.Q_N a_1511_4112# 0.0407f
C4519 a_7072_3239# x45.Q_N 0.162f
C4520 VDD a_4074_4775# 0.494f
C4521 a_7317_2550# a_7763_2366# 0.0367f
C4522 a_10345_3239# a_10794_3239# 3.74e-19
C4523 D[5] x27.Q_N 0.00536f
C4524 a_9709_2550# x42.Q_N 0.00196f
C4525 D[1] a_10628_3239# 0.348f
C4526 a_8590_3239# a_8383_2340# 2.02e-19
C4527 a_9464_3239# a_8696_2366# 2.17e-19
C4528 VDD x20.Q_N 1.29f
C4529 a_9151_3213# a_9236_2640# 5.32e-19
C4530 a_7049_2340# VDD 0.304f
C4531 a_9369_3239# D[1] 1.36e-20
C4532 a_6710_5083# check[5] 3.95e-22
C4533 a_10794_3239# a_11076_5167# 1.65e-21
C4534 VDD a_11250_4775# 0.488f
C4535 a_11249_3213# a_11250_4775# 2.59e-19
C4536 a_11075_3605# a_10795_4801# 8.52e-21
C4537 a_10628_3239# a_11544_4775# 9.66e-21
C4538 x5.X eob 0.155f
C4539 a_1227_4801# a_3619_4801# 7.69e-21
C4540 a_2389_5648# check[2] 0.138f
C4541 a_1682_4775# a_2194_4801# 9.75e-19
C4542 a_1061_4801# x20.Q_N 2.14e-19
C4543 a_6546_2340# x4.X 0.00704f
C4544 x5.X x4.A 6.17e-19
C4545 a_6845_2340# x45.Q_N 3.65e-20
C4546 a_7317_2550# a_7050_4086# 2.22e-22
C4547 x77.Y a_4854_3213# 0.142f
C4548 D[3] VDD 0.221f
C4549 a_8938_2340# a_9236_2640# 0.137f
C4550 a_8696_2366# a_9237_2340# 0.125f
C4551 a_11543_3213# a_12146_3239# 0.0552f
C4552 a_1112_2340# VDD 0.227f
C4553 x66.Q_N VDD 0.0716f
C4554 a_11543_3213# a_11761_3239# 3.73e-19
C4555 a_11856_3239# a_11389_3239# 0.00316f
C4556 check[1] a_7562_4112# 1.69e-19
C4557 a_9655_2648# x4.X 2.86e-19
C4558 x5.X a_6781_4478# 3.2e-19
C4559 check[2] a_8289_4086# 1.35e-21
C4560 sel_bit[0] a_3648_5972# 2.6e-19
C4561 a_11183_3239# x4.X 6.32e-19
C4562 a_2061_2340# a_1720_2648# 1.25e-19
C4563 x75.Q_N comparator_out 1.48e-19
C4564 a_1520_2366# a_1626_2366# 0.0552f
C4565 a_1762_2340# a_2198_2732# 0.00412f
C4566 a_2060_2640# a_1996_2732# 2.13e-19
C4567 a_9238_4086# x39.Q_N 3.57e-19
C4568 check[0] a_4155_4086# 4.34e-20
C4569 a_10155_2366# a_11088_2366# 3.42e-20
C4570 a_6465_3213# a_6011_4801# 3.18e-21
C4571 D[3] a_10775_2340# 0.0131f
C4572 check[4] a_10681_4086# 0.00276f
C4573 check[6] a_6978_4801# 6.18e-20
C4574 comparator_out a_3913_4112# 2.29e-20
C4575 VDD a_8591_4801# 0.109f
C4576 a_9370_4801# check[4] 9.79e-21
C4577 comparator_out a_12030_3213# 0.00336f
C4578 a_4854_3213# check[6] 0.00397f
C4579 check[2] a_3619_4801# 6.48e-20
C4580 x4.X a_9152_4775# 0.104f
C4581 x5.X a_1926_5083# 3.49e-19
C4582 a_2389_5648# x20.Q_N 2.12e-20
C4583 a_5169_2366# check[6] 5.24e-20
C4584 check[2] a_10795_4801# 0.00106f
C4585 comparator_out x4.X 0.797f
C4586 a_6465_3213# a_6709_3521# 0.0104f
C4587 a_6010_3239# a_6930_3521# 1.09e-19
C4588 a_9441_2340# x33.Q_N 0.179f
C4589 comparator_out a_11628_2640# 0.108f
C4590 x75.Q a_6010_3239# 0.00207f
C4591 a_4854_3213# a_3912_2366# 8.4e-19
C4592 a_4367_3213# a_4154_2340# 2.17e-19
C4593 a_3618_3239# a_4657_2340# 0.00154f
C4594 a_4073_3213# a_4453_2340# 0.00199f
C4595 x33.Q_N x36.Q_N 2.37e-20
C4596 check[1] a_7159_5167# 1.92e-19
C4597 a_4018_2366# a_4388_2366# 4.11e-20
C4598 x48.Q a_3807_4801# 0.00791f
C4599 a_4367_3213# a_4538_3521# 0.00652f
C4600 a_3618_3239# a_4007_3239# 0.0019f
C4601 a_3452_3239# a_4585_3239# 2.56e-19
C4602 a_4073_3213# a_4213_3239# 0.07f
C4603 D[0] a_9151_3213# 1.24e-19
C4604 a_7246_3213# a_7317_2550# 1.66e-21
C4605 a_7072_3239# a_7049_2340# 1.03e-19
C4606 VDD a_6931_5083# 0.0163f
C4607 a_3452_3239# a_3505_4086# 5.06e-19
C4608 a_11564_2366# x33.Q_N 1e-20
C4609 a_3618_3239# VDD 0.291f
C4610 a_12346_4112# x39.Q_N 2.43e-19
C4611 a_8590_3239# check[1] 0.00666f
C4612 a_2265_2340# x4.X 0.00118f
C4613 x4.X a_4971_4801# 0.00557f
C4614 a_3619_4801# a_4074_4775# 0.153f
C4615 a_3453_4801# a_3900_5167# 0.15f
C4616 a_10776_4086# a_11089_4112# 0.272f
C4617 x5.X a_8237_4801# 0.27f
C4618 check[2] a_9465_4801# 0.00105f
C4619 x20.Q_N a_3619_4801# 4.85e-19
C4620 a_10982_3239# x42.Q_N 1.34e-20
C4621 a_9754_3239# a_9442_4086# 5.48e-21
C4622 a_6845_2340# a_7049_2340# 0.117f
C4623 a_9151_3213# a_11543_3213# 3.6e-20
C4624 a_2697_5083# x20.Q_N 2.02e-20
C4625 a_6546_2340# x57.Q_N 9.58e-21
C4626 a_9638_3213# a_11075_3605# 7.98e-21
C4627 a_6844_2640# a_7317_2550# 0.145f
C4628 a_4453_2340# x27.Q_N 0.0462f
C4629 a_9464_3239# VDD 0.18f
C4630 a_2853_5648# a_2784_5996# 0.00105f
C4631 a_9464_3239# x69.Q_N 9.58e-21
C4632 check[0] a_5845_4801# 0.00285f
C4633 a_12345_2366# check[3] 5.09e-20
C4634 a_5844_3239# a_5845_4801# 6.9e-19
C4635 a_10629_4801# a_11076_5167# 0.15f
C4636 a_10795_4801# a_11250_4775# 0.153f
C4637 a_9441_2340# check[1] 4.56e-19
C4638 check[1] x27.Q_N 3.1e-20
C4639 a_3600_4086# a_4019_4112# 0.0397f
C4640 a_4213_3239# x27.Q_N 6.11e-19
C4641 a_4155_4086# a_4389_4478# 0.00976f
C4642 a_3913_4112# a_4591_4478# 0.00652f
C4643 a_8683_3605# x4.X 0.0177f
C4644 a_7764_4112# a_7562_4112# 3.67e-19
C4645 VDD a_5170_4478# 0.00436f
C4646 a_8237_4801# a_9237_4386# 9.86e-20
C4647 a_8684_5167# a_8384_4086# 4.9e-20
C4648 a_8858_4775# a_8697_4112# 0.0025f
C4649 D[4] a_9237_2340# 1.09e-19
C4650 a_10628_3239# a_12737_3239# 1.03e-19
C4651 a_9237_2340# VDD 0.784f
C4652 VDD a_5089_5083# 0.00529f
C4653 D[0] check[5] 0.417f
C4654 D[1] a_11183_3239# 1.22e-19
C4655 a_6759_3213# a_7363_4801# 1.05e-20
C4656 a_9172_2366# check[4] 2.2e-20
C4657 check[3] a_12102_4296# 0.00213f
C4658 a_2883_5674# a_2993_5674# 0.00857f
C4659 VDD a_12265_5083# 0.00506f
C4660 a_10794_3239# x36.Q_N 3.85e-19
C4661 x4.X a_4591_4478# 0.00114f
C4662 a_5897_4086# a_6846_4086# 7e-20
C4663 x4.X a_4214_4801# 7.25e-19
C4664 a_8696_2366# x4.X 0.112f
C4665 x5.X a_7247_4775# 0.00983f
C4666 x4.X a_11390_4801# 7.25e-19
C4667 a_12547_2366# VDD 0.109f
C4668 a_6011_4801# a_6199_4801# 0.162f
C4669 a_9441_2340# a_9577_2366# 0.07f
C4670 a_5845_4801# a_6376_5167# 0.0018f
C4671 a_9236_2640# a_11088_2366# 1.89e-19
C4672 a_1062_5674# sel_bit[0] 0.0419f
C4673 a_9237_2340# a_10775_2340# 0.00116f
C4674 a_6466_4775# a_7073_4801# 0.00187f
C4675 a_6292_5167# a_7247_4775# 4.7e-22
C4676 check[0] a_4855_4775# 0.0127f
C4677 a_10345_3239# a_9639_4775# 4.94e-20
C4678 a_12264_3521# x66.Q_N 2.02e-20
C4679 comparator_out D[1] 0.025f
C4680 x77.Y a_4658_4086# 1.87e-21
C4681 a_9639_4775# a_11076_5167# 7.98e-21
C4682 comparator_out x57.Q_N 2.04e-19
C4683 a_11194_2366# x4.X 3.78e-20
C4684 x4.X a_7954_4801# 0.00672f
C4685 x5.X a_9442_4086# 9.38e-19
C4686 a_9638_3213# check[2] 0.0022f
C4687 D[6] a_1996_2366# 3.71e-20
C4688 a_5896_2340# check[6] 0.00282f
C4689 a_11089_4112# a_11565_4478# 0.00133f
C4690 a_11075_3605# a_11089_4112# 1.61e-19
C4691 a_11249_3213# a_11331_4086# 1.02e-19
C4692 VDD a_11331_4086# 0.34f
C4693 a_10628_3239# a_11630_4086# 6.54e-20
C4694 a_11543_3213# a_10776_4086# 8.83e-19
C4695 a_10794_3239# a_11629_4386# 4.11e-20
C4696 a_11629_2340# a_11766_2732# 0.00907f
C4697 eob a_3373_5674# 1.33e-19
C4698 a_6759_3213# a_6606_4801# 1.61e-20
C4699 a_3452_3239# a_6198_3239# 3.65e-21
C4700 a_4680_3239# a_6010_3239# 5.35e-20
C4701 a_4367_3213# a_6291_3605# 4.38e-20
C4702 x4.X a_9578_4112# 0.0031f
C4703 a_9237_4386# a_9442_4086# 0.153f
C4704 a_8697_4112# x42.Q_N 0.0927f
C4705 a_9236_2640# check[2] 8.03e-20
C4706 a_8402_3239# a_8697_4112# 4.9e-19
C4707 a_8857_3213# a_8384_4086# 2.45e-19
C4708 a_3599_2340# a_4388_2366# 4.2e-20
C4709 a_3912_2366# a_5896_2340# 1.34e-20
C4710 a_7953_3239# D[0] 0.0968f
C4711 a_4368_4775# a_4971_4801# 0.0552f
C4712 a_11088_2366# a_11089_4112# 1.8e-19
C4713 a_10775_2340# a_11331_4086# 1.3e-22
C4714 x51.Q_N x20.Q_N 4.6e-19
C4715 a_7246_3213# a_8590_3239# 8.26e-21
C4716 x5.X a_9574_4801# 5.36e-20
C4717 a_8858_4775# a_9102_5083# 0.0104f
C4718 a_11629_2340# x33.Q_N 7.03e-21
C4719 a_8403_4801# a_9323_5083# 1.09e-19
C4720 a_3618_3239# a_3619_4801# 1.39e-19
C4721 a_2853_5648# a_2463_4775# 9.54e-20
C4722 a_3452_3239# x20.Q_N 0.00411f
C4723 x77.Y a_3170_4801# 5.69e-20
C4724 x48.Q a_3258_5648# 0.00631f
C4725 sel_bit[1] x48.Q 0.173f
C4726 a_5992_4086# a_6781_4478# 7.71e-20
C4727 a_6305_4112# a_6505_4394# 0.00185f
C4728 a_1508_5167# a_1511_4112# 3.47e-19
C4729 a_4452_2640# a_4453_4386# 1.32e-20
C4730 a_3912_2366# a_4658_4086# 7.14e-22
C4731 a_4154_2340# a_4454_4086# 3.47e-21
C4732 a_8383_2340# a_8384_4086# 5.27e-19
C4733 VDD a_1508_5167# 0.197f
C4734 a_8683_3605# D[1] 3.23e-21
C4735 sel_bit[0] x5.X 0.0739f
C4736 a_9151_3213# a_10345_3239# 6.04e-19
C4737 a_1112_2340# x51.Q_N 0.178f
C4738 D[7] a_2533_2550# 6.45e-20
C4739 eob x4.A 0.0197f
C4740 x75.Q_N VDD 0.0719f
C4741 a_1061_4801# a_1508_5167# 0.138f
C4742 a_3505_4086# a_3600_4086# 0.0968f
C4743 a_1511_4112# a_3913_4112# 1e-19
C4744 a_4657_2340# x4.X 0.0013f
C4745 x5.X a_10156_4112# 9.37e-19
C4746 check[2] a_11089_4112# 0.00131f
C4747 VDD a_3913_4112# 0.46f
C4748 D[0] x45.Q_N 0.00168f
C4749 a_4368_4775# a_4214_4801# 0.00943f
C4750 a_4074_4775# a_4586_4801# 9.75e-19
C4751 a_4855_4775# a_4767_5167# 7.71e-20
C4752 a_3900_5167# a_4008_4801# 0.00812f
C4753 a_3453_4801# x27.Q_N 2.36e-19
C4754 a_4681_4801# a_4539_5083# 0.00412f
C4755 VDD a_11195_4112# 0.00996f
C4756 a_11249_3213# a_11195_4112# 3.34e-20
C4757 D[1] a_8696_2366# 1.64e-21
C4758 x5.X a_8792_4801# 2.86e-19
C4759 a_11075_3605# a_11543_3213# 0.0633f
C4760 a_10628_3239# a_10982_3239# 0.0708f
C4761 a_10794_3239# a_11856_3239# 0.137f
C4762 a_6844_2640# x27.Q_N 1.07e-20
C4763 x20.Q_N a_4586_4801# 5.69e-20
C4764 a_6304_2366# x60.Q_N 5.09e-21
C4765 a_6845_2340# a_9237_2340# 0.00176f
C4766 a_12030_3213# VDD 0.568f
C4767 a_8802_2366# check[4] 1.3e-19
C4768 a_4007_3239# x4.X 6.32e-19
C4769 x30.Q_N a_8237_4801# 3.15e-19
C4770 x4.X a_1511_4112# 1.74f
C4771 a_11250_4775# a_11762_4801# 9.75e-19
C4772 a_10629_4801# x36.Q_N 1.22e-19
C4773 a_11544_4775# a_11390_4801# 0.00943f
C4774 a_11076_5167# a_11184_4801# 0.00812f
C4775 a_11857_4801# a_11715_5083# 0.00412f
C4776 a_12031_4775# a_11943_5167# 7.71e-20
C4777 x4.X a_11289_4394# 1.75e-19
C4778 D[4] x4.X 5.2e-19
C4779 a_4367_3213# check[0] 2.58e-20
C4780 VDD x4.X 5.74f
C4781 a_4453_4386# a_6846_4086# 2.9e-21
C4782 a_11249_3213# x4.X 0.00509f
C4783 x69.Q_N x4.X 0.00454f
C4784 a_4367_3213# a_5844_3239# 3.41e-19
C4785 a_3899_3605# comparator_out 1.95e-19
C4786 a_9237_4386# a_10156_4112# 0.162f
C4787 x5.X check[6] 0.168f
C4788 a_9238_4086# a_9954_4478# 0.0018f
C4789 a_8697_4112# a_9173_4112# 2.87e-21
C4790 a_9442_4086# a_9656_4394# 0.0104f
C4791 a_9236_2640# D[3] 0.00531f
C4792 a_9441_2340# a_9953_2732# 6.69e-20
C4793 check[6] a_6292_5167# 0.00105f
C4794 a_9237_2340# a_10155_2366# 0.0708f
C4795 a_11075_3605# a_11330_2340# 2.41e-20
C4796 a_11628_2640# VDD 0.269f
C4797 a_11543_3213# a_11088_2366# 3.36e-20
C4798 a_11249_3213# a_11628_2640# 2.68e-19
C4799 a_10794_3239# a_11629_2340# 6.38e-20
C4800 a_10628_3239# a_11833_2340# 4.77e-19
C4801 a_7317_2550# check[5] 0.00103f
C4802 a_11389_3239# D[2] 1.3e-20
C4803 x5.X check[3] 0.285f
C4804 a_8684_5167# check[4] 4.29e-21
C4805 a_9152_4775# a_10346_4801# 6.04e-19
C4806 a_1227_4801# a_1682_4775# 0.145f
C4807 a_1061_4801# x4.X 0.0131f
C4808 a_12146_3239# x36.Q_N 0.00341f
C4809 eob a_1926_5083# 0.00171f
C4810 a_11761_3239# x36.Q_N 4.03e-19
C4811 x4.X a_7318_4296# 0.0211f
C4812 a_10775_2340# x4.X 0.11f
C4813 a_1626_2366# D[6] 3.23e-20
C4814 check[0] a_4389_4112# 8.48e-21
C4815 a_1762_2340# a_2200_2366# 0.00276f
C4816 a_2061_2340# a_3504_2340# 8.18e-19
C4817 a_1520_2366# a_2401_2366# 0.00943f
C4818 a_10680_2340# x63.Q_N 0.178f
C4819 a_11088_2366# a_11330_2340# 0.124f
C4820 a_10775_2340# a_11628_2640# 0.0264f
C4821 comparator_out a_5897_4086# 2.05e-21
C4822 a_7247_4775# x30.Q_N 0.126f
C4823 a_11076_5167# a_10776_4086# 4.9e-20
C4824 a_11250_4775# a_11089_4112# 0.0025f
C4825 a_10629_4801# a_11629_4386# 9.86e-20
C4826 comparator_out a_12737_3239# 1.9e-19
C4827 comparator_out a_9709_2550# 0.00825f
C4828 check[1] a_5845_4801# 5.4e-19
C4829 check[2] a_3600_4086# 1.65e-20
C4830 check[2] a_11767_4478# 5.02e-20
C4831 a_3452_3239# a_3618_3239# 0.638f
C4832 a_11543_3213# check[2] 1.77e-20
C4833 a_3599_2340# a_4018_2366# 0.0397f
C4834 a_3912_2366# a_4590_2732# 0.00652f
C4835 a_4154_2340# a_4388_2732# 0.00976f
C4836 a_4970_3239# a_4657_2340# 3.49e-20
C4837 a_11714_3521# x39.Q_N 0.00203f
C4838 a_6399_3239# x30.Q_N 6.75e-20
C4839 check[1] a_8384_4086# 0.0126f
C4840 a_2389_5648# x4.X 0.00219f
C4841 a_4854_3213# a_5371_2366# 2.38e-19
C4842 a_11160_5167# check[3] 1.13e-19
C4843 a_4213_3239# a_4789_3239# 2.46e-21
C4844 x5.X a_6547_4086# 0.00115f
C4845 a_1976_4775# a_3453_4801# 1.75e-19
C4846 x48.Q a_4926_4296# 1.36e-19
C4847 a_6760_4775# a_6305_4112# 5.67e-20
C4848 a_5371_2366# a_5169_2366# 3.67e-19
C4849 a_11330_2340# check[2] 0.00111f
C4850 a_5845_4801# a_7050_4086# 6.96e-19
C4851 a_6292_5167# a_6547_4086# 2.46e-20
C4852 a_6466_4775# a_6845_4386# 3.92e-19
C4853 a_6011_4801# a_6846_4086# 1.18e-19
C4854 VDD a_7186_4112# 0.0326f
C4855 a_2289_4801# a_1822_4801# 0.00316f
C4856 a_1976_4775# a_2194_4801# 3.73e-19
C4857 a_5896_2340# a_5991_2340# 0.0968f
C4858 a_4388_2366# a_4793_2366# 2.46e-21
C4859 a_9151_3213# a_8590_3239# 3.79e-20
C4860 a_8236_3239# a_9101_3521# 0.00276f
C4861 a_9638_3213# a_9464_3239# 0.197f
C4862 a_8683_3605# a_8767_3605# 0.00972f
C4863 a_4970_3239# VDD 0.00144f
C4864 x54.Q_N x20.Q_N 1.47e-19
C4865 x27.Q_N a_4790_4801# 8.36e-20
C4866 a_6780_2366# x30.Q_N 9.42e-19
C4867 a_4073_3213# a_4019_4112# 3.34e-20
C4868 check[1] a_4855_4775# 1.73e-19
C4869 comparator_out a_11630_4086# 3e-20
C4870 x4.X a_8289_4086# 0.00368f
C4871 a_7072_3239# x4.X 0.00457f
C4872 a_4074_4775# a_3600_4086# 4.54e-19
C4873 a_6845_4386# a_8939_4086# 3.16e-20
C4874 a_6846_4086# a_8697_4112# 5.07e-21
C4875 a_3619_4801# a_3913_4112# 9.06e-19
C4876 a_7318_4296# a_7186_4112# 0.0258f
C4877 x45.Q_N a_6985_4112# 0.00166f
C4878 x20.Q_N a_3600_4086# 0.00304f
C4879 VDD a_4368_4775# 0.453f
C4880 a_6375_3605# x45.Q_N 8.49e-19
C4881 D[1] VDD 0.3f
C4882 D[1] a_11249_3213# 8.77e-20
C4883 x57.Q_N VDD 0.0716f
C4884 a_9464_3239# a_9236_2640# 1.11e-20
C4885 a_9638_3213# a_9237_2340# 8.72e-19
C4886 a_9151_3213# a_9441_2340# 0.00144f
C4887 x69.Q_N D[1] 2.5e-19
C4888 VDD a_11544_4775# 0.449f
C4889 a_8383_2340# check[4] 2.57e-20
C4890 a_11543_3213# a_11250_4775# 7.57e-21
C4891 a_11856_3239# a_10629_4801# 4.76e-21
C4892 a_1520_2366# eob 1.2e-19
C4893 x4.X a_3619_4801# 0.00737f
C4894 a_1682_4775# x20.Q_N 1.32e-19
C4895 a_6845_2340# x4.X 0.00277f
C4896 x27.Q_N a_4019_4112# 2.89e-22
C4897 x4.X a_10795_4801# 0.00496f
C4898 a_1520_2366# x4.A 6.86e-19
C4899 x48.Q x27.D 0.0333f
C4900 a_7317_2550# x45.Q_N 0.00196f
C4901 x77.Y a_3806_3239# 0.0112f
C4902 D[1] a_10775_2340# 0.00122f
C4903 a_9236_2640# a_9237_2340# 0.781f
C4904 a_11856_3239# a_12146_3239# 0.0282f
C4905 a_8383_2340# x60.Q_N 0.124f
C4906 a_8938_2340# a_9441_2340# 0.00187f
C4907 a_4008_4801# x27.Q_N 4.32e-20
C4908 a_12030_3213# a_11965_3239# 4.2e-20
C4909 a_8696_2366# a_9709_2550# 0.0633f
C4910 a_11856_3239# a_11761_3239# 0.00276f
C4911 a_10982_3239# a_11183_3239# 3.67e-19
C4912 a_11543_3213# x66.Q_N 0.00553f
C4913 a_12030_3213# a_12264_3521# 0.00945f
C4914 a_10155_2366# x4.X 7.73e-20
C4915 a_11965_3239# x4.X 1.05e-19
C4916 sel_bit[0] a_3373_5674# 0.0563f
C4917 a_12264_3521# x4.X 0.00103f
C4918 a_2061_2340# a_2198_2732# 0.00907f
C4919 a_2147_5083# x27.D 2.85e-21
C4920 VDD a_8897_4394# 0.00506f
C4921 a_9710_4296# x39.Q_N 1.29e-19
C4922 a_6465_3213# a_6292_5167# 3.52e-21
C4923 check[0] a_4454_4086# 0.44f
C4924 a_6291_3605# a_6466_4775# 1.33e-23
C4925 a_6759_3213# a_6011_4801# 2.05e-21
C4926 D[3] a_11330_2340# 1.99e-19
C4927 check[6] x30.Q_N 1.48e-21
C4928 VDD a_7363_4801# 0.0101f
C4929 comparator_out a_4453_4386# 2.5e-20
C4930 eob a_2398_4801# 2.92e-19
C4931 x33.Q_N check[4] 0.842f
C4932 comparator_out a_10982_3239# 0.157f
C4933 check[2] a_3900_5167# 5.02e-20
C4934 x45.Q_N a_7562_4112# 2.38e-19
C4935 x4.X a_9465_4801# 0.00321f
C4936 a_7764_4112# a_8384_4086# 8.26e-21
C4937 a_6845_4386# a_8803_4112# 3.66e-20
C4938 x5.X a_2375_5167# 1.58e-19
C4939 a_10345_3239# check[2] 0.00302f
C4940 a_3453_4801# a_5845_4801# 0.00176f
C4941 a_12345_2732# a_12547_2366# 8.94e-19
C4942 a_3504_2340# a_4453_2340# 1.03e-19
C4943 a_9709_2550# a_9578_4112# 1.72e-22
C4944 a_7363_4801# a_7318_4296# 1.9e-20
C4945 a_6198_3239# a_6375_3605# 8.94e-19
C4946 a_6759_3213# a_6709_3521# 1.21e-20
C4947 a_6010_3239# a_6605_3239# 0.00118f
C4948 x60.Q_N x33.Q_N 4.08e-19
C4949 comparator_out a_11833_2340# 0.00593f
C4950 a_5561_3239# a_6759_3213# 5.62e-20
C4951 a_4854_3213# a_4452_2640# 3.43e-19
C4952 a_4367_3213# a_4453_2340# 2.19e-19
C4953 sel_bit[0] eob 0.294f
C4954 check[6] a_5992_4086# 0.00385f
C4955 x48.Q a_2579_4801# 1.65e-19
C4956 a_4452_2640# a_5169_2366# 0.00105f
C4957 a_4971_4801# a_4453_4386# 8.84e-21
C4958 x77.Y eob 0.05f
C4959 a_3452_3239# x75.Q_N 1.07e-19
C4960 a_3899_3605# a_4007_3239# 0.00812f
C4961 a_4367_3213# a_4213_3239# 0.00943f
C4962 a_4680_3239# a_4538_3521# 0.00412f
C4963 a_4854_3213# a_4766_3605# 7.71e-20
C4964 a_4073_3213# a_4585_3239# 9.75e-19
C4965 D[0] a_9464_3239# 3.72e-20
C4966 sel_bit[0] x4.A 1.17e-20
C4967 a_6410_2366# x30.Q_N 0.0102f
C4968 VDD a_6606_4801# 0.0332f
C4969 a_3452_3239# a_3913_4112# 2.21e-19
C4970 a_3618_3239# a_3600_4086# 3.48e-19
C4971 a_3899_3605# VDD 0.182f
C4972 reset a_621_4112# 0.197f
C4973 x51.Q_N x4.X 0.0098f
C4974 a_3619_4801# a_4368_4775# 0.139f
C4975 D[5] a_4454_4086# 1.26e-20
C4976 a_4074_4775# a_3900_5167# 0.205f
C4977 a_3453_4801# a_4855_4775# 0.0492f
C4978 x20.Q_N a_3900_5167# 2.13e-19
C4979 x5.X a_8858_4775# 0.00316f
C4980 a_10681_4086# x39.Q_N 0.181f
C4981 a_11089_4112# a_11331_4086# 0.124f
C4982 x30.Q_N a_6547_4086# 1.3e-22
C4983 a_10776_4086# a_11629_4386# 0.0264f
C4984 a_2853_5648# a_3648_5972# 0.00271f
C4985 a_9754_3239# x42.Q_N 0.00969f
C4986 D[0] a_9237_2340# 1.09e-20
C4987 a_7247_4775# a_8237_4801# 0.00116f
C4988 a_7049_2340# a_7317_2550# 0.205f
C4989 a_2853_5648# a_2969_6040# 0.00149f
C4990 a_6760_4775# a_8403_4801# 1.55e-19
C4991 a_8767_3605# VDD 0.0042f
C4992 a_4925_2550# x27.Q_N 0.181f
C4993 a_6845_2340# x57.Q_N 1.07e-19
C4994 check[1] a_2883_5674# 0.195f
C4995 a_3452_3239# x4.X 0.0477f
C4996 VDD a_10346_4801# 0.192f
C4997 a_10794_3239# check[4] 1.18e-19
C4998 comparator_out a_6011_4801# 2.9e-21
C4999 a_11250_4775# a_11076_5167# 0.205f
C5000 a_10629_4801# a_12031_4775# 0.0492f
C5001 a_10795_4801# a_11544_4775# 0.139f
C5002 x60.Q_N check[1] 0.0122f
C5003 a_4585_3239# x27.Q_N 4.03e-19
C5004 a_4155_4086# a_4019_4112# 0.0282f
C5005 a_4453_4386# a_4591_4478# 1.09e-19
C5006 a_3913_4112# a_4872_4394# 1.21e-20
C5007 VDD a_2784_5996# 0.00533f
C5008 a_9638_3213# x4.X 0.116f
C5009 VDD a_5897_4086# 0.189f
C5010 a_7362_3239# a_7050_4086# 5.48e-21
C5011 a_8590_3239# x45.Q_N 1.34e-20
C5012 a_10345_3239# D[3] 0.00127f
C5013 D[1] a_11965_3239# 1.23e-20
C5014 D[4] a_9709_2550# 1.83e-20
C5015 a_8684_5167# a_8939_4086# 2.46e-20
C5016 a_9152_4775# a_8697_4112# 5.67e-20
C5017 a_12737_3239# VDD 0.189f
C5018 a_10794_3239# D[2] 5.71e-21
C5019 a_8237_4801# a_9442_4086# 6.96e-19
C5020 a_8858_4775# a_9237_4386# 3.92e-19
C5021 a_8403_4801# a_9238_4086# 1.18e-19
C5022 a_9709_2550# VDD 0.172f
C5023 D[7] x20.Q_N 5.48e-19
C5024 a_9577_2366# check[4] 4.82e-19
C5025 sel_bit[1] a_2993_5674# 4.44e-19
C5026 comparator_out a_4112_2648# 1.53e-19
C5027 comparator_out a_8697_4112# 2.29e-20
C5028 x4.X a_4872_4394# 8.47e-19
C5029 a_11075_3605# x36.Q_N 0.00192f
C5030 a_5844_3239# a_6930_3521# 0.00907f
C5031 x75.Q check[0] 0.0176f
C5032 a_5992_4086# a_6547_4086# 0.197f
C5033 a_5372_4112# x45.Q_N 8.9e-20
C5034 x4.X a_4586_4801# 5.55e-19
C5035 a_9236_2640# x4.X 0.00898f
C5036 a_5561_3239# comparator_out 0.00108f
C5037 x75.Q a_5844_3239# 0.335f
C5038 x5.X a_6199_4801# 0.00541f
C5039 x4.X a_11762_4801# 5.55e-19
C5040 x27.Q_N x45.Q_N 2.8e-20
C5041 a_1207_2340# a_1762_2340# 0.197f
C5042 a_6292_5167# a_6199_4801# 0.0367f
C5043 a_11768_2366# VDD 6.2e-19
C5044 a_6011_4801# a_4971_4801# 1.71e-20
C5045 a_6466_4775# a_6376_5167# 6.69e-20
C5046 a_6760_4775# a_7073_4801# 0.124f
C5047 sel_bit[0] x48.Q_N 3.83e-20
C5048 a_1112_2340# D[7] 0.0786f
C5049 a_9237_2340# a_11330_2340# 6.38e-20
C5050 a_9709_2550# a_10775_2340# 7.98e-21
C5051 a_9441_2340# a_11088_2366# 7.2e-21
C5052 a_11088_2366# x36.Q_N 0.0928f
C5053 a_12345_2732# x4.X 1.17e-19
C5054 x5.X x42.Q_N 0.00729f
C5055 a_2979_2366# a_3599_2340# 8.26e-21
C5056 a_2533_2550# a_2777_2366# 0.00812f
C5057 D[6] a_2401_2366# 5.27e-19
C5058 x27.D a_4318_5083# 3.45e-21
C5059 a_11629_4386# a_11565_4478# 2.13e-19
C5060 a_11630_4086# a_11289_4394# 1.25e-19
C5061 a_11089_4112# a_11195_4112# 0.051f
C5062 a_4592_2366# check[6] 8.47e-20
C5063 eob a_2788_5674# 1.71e-19
C5064 x30.Q_N a_6411_4112# 2.89e-22
C5065 a_11331_4086# a_11767_4478# 0.00412f
C5066 VDD a_11630_4086# 0.809f
C5067 a_11628_2640# a_12345_2732# 4.45e-20
C5068 a_11088_2366# a_11564_2366# 2.87e-21
C5069 a_12030_3213# a_11089_4112# 9.49e-19
C5070 a_10794_3239# a_11834_4086# 2.9e-19
C5071 a_11543_3213# a_11331_4086# 2.12e-19
C5072 a_11249_3213# a_11630_4086# 5.04e-19
C5073 a_11629_2340# a_12047_2648# 0.00276f
C5074 a_6465_3213# x30.Q_N 5.84e-19
C5075 a_2389_5648# a_2784_5996# 0.0102f
C5076 a_4854_3213# a_6759_3213# 3.71e-20
C5077 x4.X a_11089_4112# 0.109f
C5078 check[2] x27.Q_N 3.57e-20
C5079 a_9238_4086# a_9710_4296# 0.15f
C5080 a_9237_4386# x42.Q_N 0.00118f
C5081 a_8857_3213# a_8939_4086# 1.02e-19
C5082 a_8402_3239# a_9237_4386# 4.11e-20
C5083 a_1996_2732# VDD 0.00483f
C5084 a_8683_3605# a_8697_4112# 1.61e-19
C5085 a_8236_3239# a_9238_4086# 6.54e-20
C5086 a_9151_3213# a_8384_4086# 8.83e-19
C5087 a_4681_4801# a_4971_4801# 0.0282f
C5088 a_4855_4775# a_4790_4801# 4.2e-20
C5089 a_4452_2640# a_5896_2340# 6.96e-19
C5090 a_4154_2340# a_4388_2366# 0.00707f
C5091 a_3912_2366# a_4592_2366# 3.73e-19
C5092 a_11088_2366# a_11629_4386# 1.93e-22
C5093 a_7246_3213# a_7362_3239# 0.0397f
C5094 a_6759_3213# a_7181_3239# 2.87e-21
C5095 x5.X a_11715_5083# 6.65e-19
C5096 check[2] x36.Q_N 0.0011f
C5097 a_5991_2340# x30.Q_N 0.142f
C5098 a_6605_3239# a_6977_3239# 3.34e-19
C5099 a_8403_4801# a_8998_4801# 0.00118f
C5100 a_8591_4801# a_8768_5167# 8.94e-19
C5101 a_9152_4775# a_9102_5083# 1.21e-20
C5102 a_3618_3239# a_3900_5167# 1.65e-21
C5103 a_4073_3213# a_4074_4775# 2.59e-19
C5104 x75.Q D[5] 9.96e-19
C5105 a_3452_3239# a_4368_4775# 9.66e-21
C5106 a_3899_3605# a_3619_4801# 8.52e-21
C5107 a_4073_3213# x20.Q_N 8.02e-21
C5108 a_11390_4801# a_11966_4801# 2.46e-21
C5109 a_6547_4086# a_6781_4478# 0.00976f
C5110 a_6305_4112# a_6983_4478# 0.00652f
C5111 a_5992_4086# a_6411_4112# 0.0397f
C5112 a_2463_4775# a_1511_4112# 0.0111f
C5113 a_6465_3213# a_5992_4086# 2.45e-19
C5114 a_11564_2366# check[2] 1.34e-19
C5115 a_6010_3239# a_6305_4112# 4.9e-19
C5116 a_4453_2340# a_4454_4086# 1.55e-19
C5117 a_4657_2340# a_4453_4386# 1.26e-21
C5118 a_5991_2340# a_6780_2732# 7.71e-20
C5119 a_8383_2340# a_8939_4086# 1.3e-22
C5120 a_6304_2366# a_6504_2648# 0.00185f
C5121 VDD a_2463_4775# 0.704f
C5122 a_8696_2366# a_8697_4112# 1.8e-19
C5123 a_8236_3239# a_8288_2340# 4.5e-19
C5124 a_5845_4801# check[5] 8.72e-20
C5125 a_6011_4801# a_7954_4801# 8.38e-21
C5126 a_9638_3213# D[1] 0.0115f
C5127 a_5088_3521# x75.Q_N 2.02e-20
C5128 a_7362_3239# a_6844_2640# 5.05e-21
C5129 a_9755_4801# a_9710_4296# 1.9e-20
C5130 check[1] a_4454_4086# 2.15e-20
C5131 a_10346_4801# a_10795_4801# 3.41e-19
C5132 check[4] a_10629_4801# 0.413f
C5133 comparator_out a_897_4112# 7.09e-20
C5134 a_1227_4801# a_1976_4775# 0.132f
C5135 a_1682_4775# a_1508_5167# 0.205f
C5136 a_1061_4801# a_2463_4775# 0.0492f
C5137 a_3600_4086# a_3913_4112# 0.273f
C5138 D[0] x4.X 0.0011f
C5139 x54.Q_N x4.X 0.00996f
C5140 check[2] a_11629_4386# 1.44e-19
C5141 VDD a_4453_4386# 0.593f
C5142 a_5991_2340# a_5992_4086# 5.27e-19
C5143 a_4681_4801# a_4214_4801# 0.00316f
C5144 a_4368_4775# a_4586_4801# 3.73e-19
C5145 a_4074_4775# x27.Q_N 1.34e-19
C5146 check[5] a_8384_4086# 0.0042f
C5147 VDD a_12346_4478# 0.0042f
C5148 x20.Q_N x27.Q_N 1.21e-20
C5149 a_10345_3239# a_9237_2340# 4.83e-19
C5150 D[1] a_9236_2640# 5.41e-19
C5151 a_10982_3239# VDD 0.109f
C5152 a_11543_3213# a_12030_3213# 0.273f
C5153 a_6844_2640# x60.Q_N 1.38e-19
C5154 a_7049_2340# x27.Q_N 8.08e-21
C5155 a_10794_3239# a_11159_3605# 4.45e-20
C5156 a_11249_3213# a_10982_3239# 6.99e-20
C5157 a_5088_3521# x4.X 0.0012f
C5158 D[6] eob 8.49e-20
C5159 x4.X a_3600_4086# 0.106f
C5160 a_11857_4801# a_11390_4801# 0.00316f
C5161 a_11544_4775# a_11762_4801# 3.73e-19
C5162 a_11250_4775# x36.Q_N 2.08e-20
C5163 x4.X a_11767_4478# 0.00114f
C5164 a_4155_4086# x45.Q_N 1.43e-20
C5165 a_11543_3213# x4.X 0.111f
C5166 a_4680_3239# a_5844_3239# 6.38e-20
C5167 a_4854_3213# comparator_out 0.00379f
C5168 a_9710_4296# a_9954_4478# 0.00972f
C5169 a_8697_4112# a_9578_4112# 0.00943f
C5170 sel_bit[1] a_621_4112# 1.03e-20
C5171 a_9442_4086# a_10156_4112# 6.99e-20
C5172 a_9238_4086# a_10681_4086# 2.08e-19
C5173 a_8939_4086# a_9377_4112# 0.00276f
C5174 a_8857_3213# a_8803_4112# 3.34e-20
C5175 check[6] a_7247_4775# 2.19e-20
C5176 a_9709_2550# a_10155_2366# 0.0367f
C5177 D[2] a_12146_3239# 9.48e-20
C5178 a_10982_3239# a_10775_2340# 2.02e-19
C5179 x33.Q_N a_8939_4086# 1.3e-22
C5180 a_11833_2340# VDD 0.304f
C5181 a_11543_3213# a_11628_2640# 5.32e-19
C5182 a_11856_3239# a_11088_2366# 2.17e-19
C5183 a_11761_3239# D[2] 1.36e-20
C5184 a_1682_4775# x4.X 0.176f
C5185 a_9639_4775# check[4] 0.0122f
C5186 D[3] x36.Q_N 0.00274f
C5187 eob a_2375_5167# 5.84e-19
C5188 x66.Q_N x36.Q_N 0.02f
C5189 a_2389_5648# a_2463_4775# 0.00225f
C5190 a_11330_2340# x4.X 0.0071f
C5191 check[2] a_1976_4775# 0.00168f
C5192 check[0] a_4794_4112# 1.51e-19
C5193 a_1762_2340# a_3599_2340# 1.86e-21
C5194 D[3] a_11564_2366# 3.38e-20
C5195 a_2060_2640# a_2401_2366# 0.00118f
C5196 a_1520_2366# a_3912_2366# 6.12e-21
C5197 a_2061_2340# a_2200_2366# 2.56e-19
C5198 a_11088_2366# a_11629_2340# 0.125f
C5199 a_11330_2340# a_11628_2640# 0.137f
C5200 a_11544_4775# a_11089_4112# 5.67e-20
C5201 a_10629_4801# a_11834_4086# 6.96e-19
C5202 a_11076_5167# a_11331_4086# 2.46e-20
C5203 a_10795_4801# a_11630_4086# 1.18e-19
C5204 a_11250_4775# a_11629_4386# 3.92e-19
C5205 a_6199_4801# x30.Q_N 4.57e-21
C5206 a_2853_5648# x5.X 6.24e-19
C5207 x33.Q_N a_10983_4801# 1e-19
C5208 check[1] a_6466_4775# 5.74e-19
C5209 check[2] a_12048_4394# 1.36e-20
C5210 a_10628_3239# x5.X 9.1e-20
C5211 a_3452_3239# a_3899_3605# 0.141f
C5212 a_3618_3239# a_4073_3213# 0.149f
C5213 D[6] a_4592_2366# 3.35e-19
C5214 a_1720_2648# x20.Q_N 2.75e-19
C5215 a_4452_2640# a_4590_2732# 1.09e-19
C5216 a_4154_2340# a_4018_2366# 0.0282f
C5217 a_3912_2366# a_4871_2648# 1.21e-20
C5218 VDD a_6011_4801# 0.593f
C5219 a_12146_3239# a_11834_4086# 5.48e-21
C5220 x30.Q_N x42.Q_N 1.63e-20
C5221 a_5371_2366# x30.Q_N 1.34e-20
C5222 a_8402_3239# x30.Q_N 3.97e-20
C5223 a_11389_3239# x39.Q_N 0.0314f
C5224 check[5] a_7182_4801# 1.11e-20
C5225 VDD a_11966_4801# 7.87e-19
C5226 check[1] a_8939_4086# 3.29e-19
C5227 x5.X a_6846_4086# 0.261f
C5228 a_5845_4801# x45.Q_N 3.67e-20
C5229 a_7073_4801# a_6305_4112# 3.76e-19
C5230 a_6760_4775# a_6845_4386# 7.46e-19
C5231 a_2463_4775# a_3619_4801# 3.31e-19
C5232 a_2289_4801# a_3453_4801# 6.38e-20
C5233 a_6199_4801# a_5992_4086# 3.44e-19
C5234 a_11629_2340# check[2] 1.99e-19
C5235 a_4112_2648# VDD 0.00555f
C5236 VDD a_8697_4112# 0.448f
C5237 a_2463_4775# a_2697_5083# 0.00945f
C5238 a_1976_4775# x20.Q_N 0.0094f
C5239 a_1415_4801# a_1616_4801# 3.67e-19
C5240 a_2289_4801# a_2194_4801# 0.00276f
C5241 a_12345_2366# VSS 8.87e-19
C5242 a_11969_2366# VSS 0.182f
C5243 a_11768_2366# VSS 0.00989f
C5244 a_11564_2366# VSS 0.00207f
C5245 a_12547_2366# VSS 0.0962f
C5246 a_12345_2732# VSS 3.33e-19
C5247 a_12047_2648# VSS 4.04e-19
C5248 a_11194_2366# VSS 0.158f
C5249 a_11766_2732# VSS 0.0011f
C5250 a_11564_2732# VSS 1.58e-19
C5251 a_11288_2648# VSS 1.45e-19
C5252 a_9953_2366# VSS 6.96e-19
C5253 x63.Q_N VSS 0.1f
C5254 a_12101_2550# VSS 0.262f
C5255 a_11833_2340# VSS 0.29f
C5256 a_11629_2340# VSS 0.606f
C5257 a_11628_2640# VSS 0.419f
C5258 a_11330_2340# VSS 0.251f
C5259 a_11088_2366# VSS 0.387f
C5260 a_10775_2340# VSS 0.458f
C5261 a_9577_2366# VSS 0.18f
C5262 a_9376_2366# VSS 0.00923f
C5263 a_9172_2366# VSS 0.00192f
C5264 a_10680_2340# VSS 0.225f
C5265 D[3] VSS 0.365f
C5266 a_10155_2366# VSS 0.0926f
C5267 a_8802_2366# VSS 0.157f
C5268 a_9374_2732# VSS 3.84e-19
C5269 a_7561_2366# VSS 6.96e-19
C5270 x60.Q_N VSS 0.1f
C5271 a_9709_2550# VSS 0.256f
C5272 a_9441_2340# VSS 0.286f
C5273 a_9237_2340# VSS 0.512f
C5274 a_9236_2640# VSS 0.4f
C5275 a_8938_2340# VSS 0.249f
C5276 a_8696_2366# VSS 0.385f
C5277 a_8383_2340# VSS 0.456f
C5278 a_7185_2366# VSS 0.18f
C5279 a_6984_2366# VSS 0.00923f
C5280 a_6780_2366# VSS 0.00192f
C5281 a_8288_2340# VSS 0.225f
C5282 D[4] VSS 0.365f
C5283 a_7763_2366# VSS 0.0926f
C5284 a_6410_2366# VSS 0.157f
C5285 a_6982_2732# VSS 3.84e-19
C5286 a_5169_2366# VSS 6.96e-19
C5287 x57.Q_N VSS 0.1f
C5288 a_7317_2550# VSS 0.256f
C5289 a_7049_2340# VSS 0.286f
C5290 a_6845_2340# VSS 0.513f
C5291 a_6844_2640# VSS 0.4f
C5292 a_6546_2340# VSS 0.249f
C5293 a_6304_2366# VSS 0.385f
C5294 a_5991_2340# VSS 0.456f
C5295 a_4793_2366# VSS 0.18f
C5296 a_4592_2366# VSS 0.00923f
C5297 a_4388_2366# VSS 0.00192f
C5298 a_5896_2340# VSS 0.225f
C5299 D[5] VSS 0.393f
C5300 a_5371_2366# VSS 0.0926f
C5301 a_4018_2366# VSS 0.157f
C5302 a_4590_2732# VSS 3.84e-19
C5303 a_2777_2366# VSS 0.00168f
C5304 x54.Q_N VSS 0.1f
C5305 a_4925_2550# VSS 0.256f
C5306 a_4657_2340# VSS 0.286f
C5307 a_4453_2340# VSS 0.513f
C5308 a_4452_2640# VSS 0.4f
C5309 a_4154_2340# VSS 0.249f
C5310 a_3912_2366# VSS 0.385f
C5311 a_3599_2340# VSS 0.458f
C5312 a_2401_2366# VSS 0.18f
C5313 a_2200_2366# VSS 0.00923f
C5314 a_1996_2366# VSS 0.00192f
C5315 a_3504_2340# VSS 0.226f
C5316 D[6] VSS 0.604f
C5317 a_2979_2366# VSS 0.0988f
C5318 a_1626_2366# VSS 0.157f
C5319 a_2198_2732# VSS 3.84e-19
C5320 x51.Q_N VSS 0.1f
C5321 a_2533_2550# VSS 0.263f
C5322 a_2265_2340# VSS 0.289f
C5323 a_2061_2340# VSS 0.517f
C5324 a_2060_2640# VSS 0.527f
C5325 a_1762_2340# VSS 0.25f
C5326 a_1520_2366# VSS 0.387f
C5327 a_1207_2340# VSS 0.469f
C5328 D[7] VSS 0.536f
C5329 a_1112_2340# VSS 0.247f
C5330 a_11965_3239# VSS 0.00208f
C5331 a_12146_3239# VSS 0.159f
C5332 D[2] VSS 1.11f
C5333 a_12737_3239# VSS 0.252f
C5334 x66.Q_N VSS 0.102f
C5335 a_12264_3521# VSS 3.9e-19
C5336 a_11761_3239# VSS 0.00967f
C5337 a_11183_3239# VSS 0.00168f
C5338 a_11389_3239# VSS 0.181f
C5339 a_11942_3605# VSS 2.25e-19
C5340 a_11714_3521# VSS 0.00103f
C5341 a_11493_3521# VSS 2.34e-19
C5342 a_9573_3239# VSS 0.00192f
C5343 a_9754_3239# VSS 0.157f
C5344 a_10982_3239# VSS 0.0988f
C5345 a_11856_3239# VSS 0.25f
C5346 a_12030_3213# VSS 0.463f
C5347 a_11543_3213# VSS 0.389f
C5348 a_11075_3605# VSS 0.259f
C5349 a_11249_3213# VSS 0.281f
C5350 a_10794_3239# VSS 0.519f
C5351 a_10628_3239# VSS 0.509f
C5352 D[1] VSS 0.467f
C5353 a_10345_3239# VSS 0.222f
C5354 x69.Q_N VSS 0.1f
C5355 a_9369_3239# VSS 0.00923f
C5356 a_8791_3239# VSS 0.00168f
C5357 a_8997_3239# VSS 0.18f
C5358 a_9322_3521# VSS 3.84e-19
C5359 a_7181_3239# VSS 0.00192f
C5360 a_7362_3239# VSS 0.157f
C5361 a_8590_3239# VSS 0.0988f
C5362 a_9464_3239# VSS 0.246f
C5363 a_9638_3213# VSS 0.446f
C5364 a_9151_3213# VSS 0.38f
C5365 a_8683_3605# VSS 0.258f
C5366 a_8857_3213# VSS 0.28f
C5367 a_8402_3239# VSS 0.519f
C5368 a_8236_3239# VSS 0.506f
C5369 D[0] VSS 0.471f
C5370 a_7953_3239# VSS 0.222f
C5371 x72.Q_N VSS 0.1f
C5372 a_6977_3239# VSS 0.00923f
C5373 a_6399_3239# VSS 0.00168f
C5374 a_6605_3239# VSS 0.18f
C5375 a_6930_3521# VSS 3.84e-19
C5376 a_4789_3239# VSS 0.00196f
C5377 a_4970_3239# VSS 0.157f
C5378 a_6198_3239# VSS 0.0988f
C5379 a_7072_3239# VSS 0.246f
C5380 a_7246_3213# VSS 0.446f
C5381 a_6759_3213# VSS 0.38f
C5382 a_6291_3605# VSS 0.258f
C5383 a_6465_3213# VSS 0.28f
C5384 a_6010_3239# VSS 0.519f
C5385 comparator_out VSS 11.6f
C5386 a_5844_3239# VSS 0.506f
C5387 x75.Q VSS 0.239f
C5388 a_5561_3239# VSS 0.222f
C5389 x75.Q_N VSS 0.1f
C5390 a_4585_3239# VSS 0.00943f
C5391 a_4007_3239# VSS 0.00202f
C5392 a_4213_3239# VSS 0.181f
C5393 a_4538_3521# VSS 3.84e-19
C5394 a_3806_3239# VSS 0.263f
C5395 a_4680_3239# VSS 0.246f
C5396 a_4854_3213# VSS 0.446f
C5397 a_4367_3213# VSS 0.379f
C5398 a_3899_3605# VSS 0.261f
C5399 a_4073_3213# VSS 0.28f
C5400 a_3618_3239# VSS 0.751f
C5401 a_3452_3239# VSS 0.888f
C5402 x77.Y VSS 1.02f
C5403 a_12346_4112# VSS 0.00226f
C5404 a_11970_4112# VSS 0.183f
C5405 a_11769_4112# VSS 0.00991f
C5406 a_11565_4112# VSS 0.00168f
C5407 a_12548_4112# VSS 0.102f
C5408 a_12346_4478# VSS 3.33e-19
C5409 a_12048_4394# VSS 3.91e-19
C5410 a_11195_4112# VSS 0.148f
C5411 a_11767_4478# VSS 0.00107f
C5412 a_11565_4478# VSS 1.58e-19
C5413 a_11289_4394# VSS 1.48e-19
C5414 a_9954_4112# VSS 0.00168f
C5415 x39.Q_N VSS 1.23f
C5416 a_12102_4296# VSS 0.261f
C5417 a_11834_4086# VSS 0.279f
C5418 a_11630_4086# VSS 0.588f
C5419 a_11629_4386# VSS 0.537f
C5420 a_11331_4086# VSS 0.238f
C5421 a_11089_4112# VSS 0.318f
C5422 a_10776_4086# VSS 0.425f
C5423 a_9578_4112# VSS 0.18f
C5424 a_9377_4112# VSS 0.00923f
C5425 a_9173_4112# VSS 0.00155f
C5426 a_10681_4086# VSS 0.207f
C5427 a_10156_4112# VSS 0.0984f
C5428 a_8803_4112# VSS 0.147f
C5429 a_9375_4478# VSS 3.84e-19
C5430 a_7562_4112# VSS 0.00168f
C5431 x42.Q_N VSS 1.22f
C5432 a_9710_4296# VSS 0.255f
C5433 a_9442_4086# VSS 0.275f
C5434 a_9238_4086# VSS 0.484f
C5435 a_9237_4386# VSS 0.515f
C5436 a_8939_4086# VSS 0.236f
C5437 a_8697_4112# VSS 0.316f
C5438 a_8384_4086# VSS 0.423f
C5439 a_7186_4112# VSS 0.18f
C5440 a_6985_4112# VSS 0.00923f
C5441 a_6781_4112# VSS 0.00157f
C5442 a_8289_4086# VSS 0.205f
C5443 a_7764_4112# VSS 0.0984f
C5444 a_6411_4112# VSS 0.147f
C5445 a_6983_4478# VSS 3.84e-19
C5446 a_5170_4112# VSS 0.00168f
C5447 x45.Q_N VSS 1.22f
C5448 a_7318_4296# VSS 0.255f
C5449 a_7050_4086# VSS 0.275f
C5450 a_6846_4086# VSS 0.484f
C5451 a_6845_4386# VSS 0.515f
C5452 a_6547_4086# VSS 0.236f
C5453 a_6305_4112# VSS 0.316f
C5454 a_5992_4086# VSS 0.423f
C5455 a_4794_4112# VSS 0.18f
C5456 a_4593_4112# VSS 0.00923f
C5457 a_4389_4112# VSS 0.00192f
C5458 a_5897_4086# VSS 0.211f
C5459 a_5372_4112# VSS 0.0984f
C5460 a_4019_4112# VSS 0.157f
C5461 a_4591_4478# VSS 3.84e-19
C5462 x48.Q_N VSS 0.1f
C5463 a_4926_4296# VSS 0.255f
C5464 a_4658_4086# VSS 0.275f
C5465 a_4454_4086# VSS 0.486f
C5466 a_4453_4386# VSS 0.515f
C5467 a_4155_4086# VSS 0.243f
C5468 a_3913_4112# VSS 0.373f
C5469 a_3600_4086# VSS 0.443f
C5470 a_3505_4086# VSS 0.225f
C5471 a_1511_4112# VSS 2.05f
C5472 x4.A VSS 0.932f
C5473 a_897_4112# VSS 0.522f
C5474 x3.A VSS 0.206f
C5475 a_621_4112# VSS 0.284f
C5476 reset VSS 0.247f
C5477 a_11966_4801# VSS 0.00215f
C5478 a_12147_4801# VSS 0.161f
C5479 check[3] VSS 1.3f
C5480 a_12738_4801# VSS 0.255f
C5481 x36.Q_N VSS 1.28f
C5482 a_12265_5083# VSS 5.88e-19
C5483 a_11762_4801# VSS 0.00989f
C5484 a_11184_4801# VSS 0.00168f
C5485 a_11390_4801# VSS 0.181f
C5486 a_11943_5167# VSS 2.29e-19
C5487 a_11715_5083# VSS 0.00114f
C5488 a_11494_5083# VSS 2.58e-19
C5489 a_9574_4801# VSS 0.00192f
C5490 a_9755_4801# VSS 0.157f
C5491 a_10983_4801# VSS 0.0987f
C5492 a_11857_4801# VSS 0.25f
C5493 a_12031_4775# VSS 0.46f
C5494 a_11544_4775# VSS 0.386f
C5495 a_11076_5167# VSS 0.257f
C5496 a_11250_4775# VSS 0.279f
C5497 a_10795_4801# VSS 0.517f
C5498 a_10629_4801# VSS 0.488f
C5499 check[4] VSS 0.823f
C5500 a_10346_4801# VSS 0.21f
C5501 x33.Q_N VSS 1.25f
C5502 a_9370_4801# VSS 0.00923f
C5503 a_8792_4801# VSS 0.00168f
C5504 a_8998_4801# VSS 0.18f
C5505 a_9323_5083# VSS 3.84e-19
C5506 a_7182_4801# VSS 0.00192f
C5507 a_7363_4801# VSS 0.157f
C5508 a_8591_4801# VSS 0.0987f
C5509 a_9465_4801# VSS 0.244f
C5510 a_9639_4775# VSS 0.435f
C5511 a_9152_4775# VSS 0.373f
C5512 a_8684_5167# VSS 0.257f
C5513 a_8858_4775# VSS 0.276f
C5514 a_8403_4801# VSS 0.515f
C5515 a_8237_4801# VSS 0.484f
C5516 check[5] VSS 0.83f
C5517 a_7954_4801# VSS 0.207f
C5518 x30.Q_N VSS 1.26f
C5519 a_6978_4801# VSS 0.00923f
C5520 a_6400_4801# VSS 0.00168f
C5521 a_6606_4801# VSS 0.18f
C5522 a_6931_5083# VSS 3.84e-19
C5523 a_4790_4801# VSS 0.00192f
C5524 a_4971_4801# VSS 0.157f
C5525 a_6199_4801# VSS 0.0987f
C5526 a_7073_4801# VSS 0.244f
C5527 a_7247_4775# VSS 0.435f
C5528 a_6760_4775# VSS 0.373f
C5529 a_6292_5167# VSS 0.257f
C5530 a_6466_4775# VSS 0.276f
C5531 a_6011_4801# VSS 0.515f
C5532 a_5845_4801# VSS 0.484f
C5533 check[6] VSS 0.845f
C5534 a_5562_4801# VSS 0.207f
C5535 x27.Q_N VSS 1.25f
C5536 a_4586_4801# VSS 0.00923f
C5537 a_4008_4801# VSS 0.00168f
C5538 a_4214_4801# VSS 0.18f
C5539 a_4539_5083# VSS 3.84e-19
C5540 a_2398_4801# VSS 0.00192f
C5541 a_2579_4801# VSS 0.157f
C5542 a_3807_4801# VSS 0.0987f
C5543 a_4681_4801# VSS 0.244f
C5544 a_4855_4775# VSS 0.435f
C5545 a_4368_4775# VSS 0.373f
C5546 a_3900_5167# VSS 0.257f
C5547 a_4074_4775# VSS 0.275f
C5548 a_3619_4801# VSS 0.513f
C5549 a_3453_4801# VSS 0.481f
C5550 x27.D VSS 0.243f
C5551 a_3170_4801# VSS 0.22f
C5552 x20.Q_N VSS 1.25f
C5553 a_2194_4801# VSS 0.00923f
C5554 a_1616_4801# VSS 0.00168f
C5555 a_1822_4801# VSS 0.18f
C5556 a_2147_5083# VSS 3.84e-19
C5557 a_1415_4801# VSS 0.0987f
C5558 a_2289_4801# VSS 0.242f
C5559 a_2463_4775# VSS 0.429f
C5560 a_1976_4775# VSS 0.37f
C5561 a_1508_5167# VSS 0.256f
C5562 x4.X VSS 16.6f
C5563 a_1682_4775# VSS 0.275f
C5564 a_1227_4801# VSS 0.516f
C5565 a_1061_4801# VSS 0.541f
C5566 a_3877_5674# VSS 0.00437f
C5567 a_3671_5674# VSS 0.00563f
C5568 a_2993_5674# VSS 0.00182f
C5569 a_2788_5674# VSS 0.00372f
C5570 a_3373_5674# VSS 0.115f
C5571 a_3258_5648# VSS 0.229f
C5572 check[0] VSS 2.45f
C5573 x48.Q VSS 0.615f
C5574 sel_bit[1] VSS 1.15f
C5575 a_2883_5674# VSS 0.185f
C5576 a_2784_5996# VSS 2.03e-19
C5577 eob VSS 2.55f
C5578 x5.X VSS 13f
C5579 check[1] VSS 2.75f
C5580 a_2853_5648# VSS 0.373f
C5581 sel_bit[0] VSS 0.54f
C5582 check[2] VSS 4.55f
C5583 a_2389_5648# VSS 0.48f
C5584 a_1338_5674# VSS 0.322f
C5585 x5.A VSS 0.226f
C5586 a_1062_5674# VSS 0.274f
C5587 clk_sar VSS 0.214f
C5588 VDD VSS 0.106p
C5589 x5.X.n0 VSS 0.112f
C5590 x5.X.n1 VSS 0.112f
C5591 x5.X.n2 VSS 0.0643f
C5592 x5.X.n3 VSS 0.0507f
C5593 x5.X.n4 VSS 0.0683f
C5594 x5.X.t2 VSS 0.00811f
C5595 x5.X.t3 VSS 0.00811f
C5596 x5.X.n5 VSS 0.0164f
C5597 x5.X.n6 VSS 8.69e-19
C5598 x5.X.t1 VSS 0.00527f
C5599 x5.X.t0 VSS 0.00527f
C5600 x5.X.n7 VSS 0.0105f
C5601 x5.X.n8 VSS 0.0106f
C5602 x5.X.t20 VSS 0.0124f
C5603 x5.X.t7 VSS 0.0096f
C5604 x5.X.n9 VSS 0.0243f
C5605 x5.X.n10 VSS 0.00725f
C5606 x5.X.n11 VSS 0.00448f
C5607 x5.X.n12 VSS 0.00181f
C5608 x5.X.t11 VSS 0.0121f
C5609 x5.X.n13 VSS 0.0125f
C5610 x5.X.n14 VSS 0.0014f
C5611 x5.X.t16 VSS 0.00914f
C5612 x5.X.n15 VSS 0.0111f
C5613 x5.X.n16 VSS 0.00251f
C5614 x5.X.n17 VSS 0.00377f
C5615 x5.X.n18 VSS 0.00447f
C5616 x5.X.n19 VSS 0.00181f
C5617 x5.X.t9 VSS 0.0122f
C5618 x5.X.n20 VSS 0.0126f
C5619 x5.X.n21 VSS 0.0014f
C5620 x5.X.t14 VSS 0.00902f
C5621 x5.X.n22 VSS 0.0109f
C5622 x5.X.n23 VSS 0.00277f
C5623 x5.X.n24 VSS 0.0479f
C5624 x5.X.n25 VSS 0.311f
C5625 x5.X.n26 VSS 0.00447f
C5626 x5.X.n27 VSS 0.00181f
C5627 x5.X.t17 VSS 0.0122f
C5628 x5.X.n28 VSS 0.0125f
C5629 x5.X.n29 VSS 0.0014f
C5630 x5.X.t4 VSS 0.0091f
C5631 x5.X.n30 VSS 0.011f
C5632 x5.X.n31 VSS 0.00263f
C5633 x5.X.n32 VSS 0.0052f
C5634 x5.X.n33 VSS 0.00447f
C5635 x5.X.n34 VSS 0.00181f
C5636 x5.X.t13 VSS 0.0122f
C5637 x5.X.n35 VSS 0.0126f
C5638 x5.X.n36 VSS 0.0014f
C5639 x5.X.t21 VSS 0.00902f
C5640 x5.X.n37 VSS 0.0109f
C5641 x5.X.n38 VSS 0.00277f
C5642 x5.X.n39 VSS 0.0472f
C5643 x5.X.n40 VSS 0.221f
C5644 x5.X.n41 VSS 0.00447f
C5645 x5.X.n42 VSS 0.00181f
C5646 x5.X.t18 VSS 0.0122f
C5647 x5.X.n43 VSS 0.0125f
C5648 x5.X.n44 VSS 0.0014f
C5649 x5.X.t5 VSS 0.0091f
C5650 x5.X.n45 VSS 0.011f
C5651 x5.X.n46 VSS 0.00256f
C5652 x5.X.n47 VSS 0.00533f
C5653 x5.X.n48 VSS 0.00447f
C5654 x5.X.n49 VSS 0.00181f
C5655 x5.X.t10 VSS 0.0122f
C5656 x5.X.n50 VSS 0.0126f
C5657 x5.X.n51 VSS 0.0014f
C5658 x5.X.t15 VSS 0.00902f
C5659 x5.X.n52 VSS 0.0109f
C5660 x5.X.n53 VSS 0.00279f
C5661 x5.X.n54 VSS 0.0466f
C5662 x5.X.n55 VSS 0.22f
C5663 x5.X.n56 VSS 0.00447f
C5664 x5.X.n57 VSS 0.00181f
C5665 x5.X.t19 VSS 0.0122f
C5666 x5.X.n58 VSS 0.0125f
C5667 x5.X.n59 VSS 0.0014f
C5668 x5.X.t6 VSS 0.0091f
C5669 x5.X.n60 VSS 0.011f
C5670 x5.X.n61 VSS 0.00265f
C5671 x5.X.n62 VSS 0.0391f
C5672 x5.X.n63 VSS 0.21f
C5673 x5.X.n64 VSS 0.00447f
C5674 x5.X.n65 VSS 0.00181f
C5675 x5.X.t8 VSS 0.0122f
C5676 x5.X.n66 VSS 0.0125f
C5677 x5.X.n67 VSS 0.0014f
C5678 x5.X.t12 VSS 0.0091f
C5679 x5.X.n68 VSS 0.011f
C5680 x5.X.n69 VSS 0.00264f
C5681 x5.X.n70 VSS 0.00429f
C5682 x5.X.n71 VSS 0.00404f
C5683 x5.X.n72 VSS 0.202f
C5684 x5.X.n73 VSS 0.0254f
C5685 check[2].t1 VSS 0.0384f
C5686 check[2].n0 VSS 0.00289f
C5687 check[2].t3 VSS 0.0197f
C5688 check[2].t2 VSS 0.0123f
C5689 check[2].n1 VSS 0.0406f
C5690 check[2].n2 VSS 0.629f
C5691 check[2].t5 VSS 0.0179f
C5692 check[2].t4 VSS 0.0125f
C5693 check[2].n3 VSS 0.0364f
C5694 check[2].n4 VSS 0.0138f
C5695 check[2].n5 VSS 0.836f
C5696 check[2].n6 VSS 0.0257f
C5697 check[2].n7 VSS 0.198f
C5698 check[2].t0 VSS 0.0144f
C5699 check[2].n8 VSS 0.0246f
C5700 x4.X.n0 VSS 0.00768f
C5701 x4.X.n1 VSS 0.00767f
C5702 x4.X.n2 VSS 0.00768f
C5703 x4.X.n3 VSS 0.00767f
C5704 x4.X.n4 VSS 0.00768f
C5705 x4.X.n5 VSS 0.00779f
C5706 x4.X.n6 VSS 0.0356f
C5707 x4.X.n7 VSS 0.00746f
C5708 x4.X.n8 VSS 0.00423f
C5709 x4.X.n9 VSS 0.00216f
C5710 x4.X.n10 VSS 0.00427f
C5711 x4.X.n11 VSS 0.0017f
C5712 x4.X.n12 VSS 0.00446f
C5713 x4.X.t20 VSS 0.00963f
C5714 x4.X.t26 VSS 0.00963f
C5715 x4.X.n13 VSS 0.0238f
C5716 x4.X.t19 VSS 0.00963f
C5717 x4.X.t30 VSS 0.00963f
C5718 x4.X.n14 VSS 0.0238f
C5719 x4.X.t27 VSS 0.00963f
C5720 x4.X.t18 VSS 0.00963f
C5721 x4.X.n15 VSS 0.0238f
C5722 x4.X.t23 VSS 0.00963f
C5723 x4.X.t16 VSS 0.00963f
C5724 x4.X.n16 VSS 0.0238f
C5725 x4.X.t22 VSS 0.00963f
C5726 x4.X.t17 VSS 0.00963f
C5727 x4.X.n17 VSS 0.0368f
C5728 x4.X.t24 VSS 0.00963f
C5729 x4.X.t28 VSS 0.00963f
C5730 x4.X.n18 VSS 0.0238f
C5731 x4.X.n19 VSS 0.0926f
C5732 x4.X.t25 VSS 0.00963f
C5733 x4.X.t29 VSS 0.00963f
C5734 x4.X.n20 VSS 0.0238f
C5735 x4.X.n21 VSS 0.0559f
C5736 x4.X.n22 VSS 0.00913f
C5737 x4.X.t21 VSS 0.00821f
C5738 x4.X.n23 VSS 0.00963f
C5739 x4.X.t66 VSS 0.0152f
C5740 x4.X.t32 VSS 0.00645f
C5741 x4.X.n24 VSS 0.0286f
C5742 x4.X.n25 VSS 0.00238f
C5743 x4.X.n26 VSS 0.0084f
C5744 x4.X.n27 VSS 0.0033f
C5745 x4.X.n28 VSS 0.0389f
C5746 x4.X.n29 VSS 0.103f
C5747 x4.X.n30 VSS 0.00153f
C5748 x4.X.t50 VSS 0.0152f
C5749 x4.X.t37 VSS 0.00644f
C5750 x4.X.n31 VSS 0.0297f
C5751 x4.X.n32 VSS 0.00977f
C5752 x4.X.n33 VSS 0.00208f
C5753 x4.X.n34 VSS 0.0273f
C5754 x4.X.n35 VSS 0.00586f
C5755 x4.X.n36 VSS 0.00803f
C5756 x4.X.n37 VSS 0.0201f
C5757 x4.X.t31 VSS 0.005f
C5758 x4.X.n38 VSS 0.00963f
C5759 x4.X.n39 VSS 0.00651f
C5760 x4.X.n40 VSS 0.00614f
C5761 x4.X.n41 VSS 0.0246f
C5762 x4.X.n42 VSS 0.0559f
C5763 x4.X.n43 VSS 0.0559f
C5764 x4.X.n44 VSS 0.0559f
C5765 x4.X.n45 VSS 0.0532f
C5766 x4.X.t2 VSS 0.00626f
C5767 x4.X.t13 VSS 0.00626f
C5768 x4.X.n46 VSS 0.0297f
C5769 x4.X.t4 VSS 0.00626f
C5770 x4.X.t8 VSS 0.00626f
C5771 x4.X.n47 VSS 0.0157f
C5772 x4.X.n48 VSS 0.0587f
C5773 x4.X.t5 VSS 0.00626f
C5774 x4.X.t9 VSS 0.00626f
C5775 x4.X.n49 VSS 0.0157f
C5776 x4.X.n50 VSS 0.0395f
C5777 x4.X.t1 VSS 0.00626f
C5778 x4.X.t11 VSS 0.00626f
C5779 x4.X.n51 VSS 0.0157f
C5780 x4.X.n52 VSS 0.0396f
C5781 x4.X.t3 VSS 0.00626f
C5782 x4.X.t12 VSS 0.00626f
C5783 x4.X.n53 VSS 0.0157f
C5784 x4.X.n54 VSS 0.0396f
C5785 x4.X.t7 VSS 0.00626f
C5786 x4.X.t14 VSS 0.00626f
C5787 x4.X.n55 VSS 0.0157f
C5788 x4.X.n56 VSS 0.0396f
C5789 x4.X.t15 VSS 0.00626f
C5790 x4.X.t10 VSS 0.00626f
C5791 x4.X.n57 VSS 0.0157f
C5792 x4.X.n58 VSS 0.0396f
C5793 x4.X.t0 VSS 0.00626f
C5794 x4.X.t6 VSS 0.00626f
C5795 x4.X.n59 VSS 0.0157f
C5796 x4.X.n60 VSS 0.0384f
C5797 x4.X.n61 VSS 0.00482f
C5798 x4.X.t58 VSS 0.009f
C5799 x4.X.t45 VSS 0.0104f
C5800 x4.X.n62 VSS 0.0242f
C5801 x4.X.n63 VSS 0.00675f
C5802 x4.X.n64 VSS 0.00238f
C5803 x4.X.n65 VSS 0.0014f
C5804 x4.X.n66 VSS 0.0083f
C5805 x4.X.n67 VSS 0.0546f
C5806 x4.X.n68 VSS 0.00482f
C5807 x4.X.t55 VSS 0.009f
C5808 x4.X.t51 VSS 0.0104f
C5809 x4.X.n69 VSS 0.0242f
C5810 x4.X.n70 VSS 0.00675f
C5811 x4.X.n71 VSS 0.00238f
C5812 x4.X.n72 VSS 0.0014f
C5813 x4.X.n73 VSS 0.00821f
C5814 x4.X.n74 VSS 0.0259f
C5815 x4.X.n75 VSS 0.113f
C5816 x4.X.n76 VSS 0.00271f
C5817 x4.X.n77 VSS 0.0014f
C5818 x4.X.t34 VSS 0.0103f
C5819 x4.X.t39 VSS 0.00868f
C5820 x4.X.n78 VSS 0.0115f
C5821 x4.X.n79 VSS 0.0128f
C5822 x4.X.n80 VSS 0.0189f
C5823 x4.X.n81 VSS 0.00271f
C5824 x4.X.n82 VSS 0.0014f
C5825 x4.X.t54 VSS 0.0103f
C5826 x4.X.t60 VSS 0.0087f
C5827 x4.X.n83 VSS 0.0117f
C5828 x4.X.n84 VSS 0.0126f
C5829 x4.X.n85 VSS 0.0588f
C5830 x4.X.n86 VSS 0.16f
C5831 x4.X.n87 VSS 0.135f
C5832 x4.X.n88 VSS 0.00482f
C5833 x4.X.t36 VSS 0.00905f
C5834 x4.X.t57 VSS 0.0103f
C5835 x4.X.n89 VSS 0.0242f
C5836 x4.X.n90 VSS 0.00661f
C5837 x4.X.n91 VSS 0.00246f
C5838 x4.X.n92 VSS 0.0014f
C5839 x4.X.n93 VSS 0.0083f
C5840 x4.X.n94 VSS 0.0547f
C5841 x4.X.n95 VSS 0.00482f
C5842 x4.X.t33 VSS 0.009f
C5843 x4.X.t63 VSS 0.0104f
C5844 x4.X.n96 VSS 0.0242f
C5845 x4.X.n97 VSS 0.00675f
C5846 x4.X.n98 VSS 0.00238f
C5847 x4.X.n99 VSS 0.0014f
C5848 x4.X.n100 VSS 0.00821f
C5849 x4.X.n101 VSS 0.0259f
C5850 x4.X.n102 VSS 0.0847f
C5851 x4.X.n103 VSS 0.125f
C5852 x4.X.n104 VSS 0.00271f
C5853 x4.X.n105 VSS 0.0014f
C5854 x4.X.t69 VSS 0.0103f
C5855 x4.X.t49 VSS 0.0087f
C5856 x4.X.n106 VSS 0.0117f
C5857 x4.X.n107 VSS 0.0126f
C5858 x4.X.n108 VSS 0.0199f
C5859 x4.X.n109 VSS 0.00271f
C5860 x4.X.n110 VSS 0.0014f
C5861 x4.X.t52 VSS 0.0103f
C5862 x4.X.t67 VSS 0.0087f
C5863 x4.X.n111 VSS 0.0117f
C5864 x4.X.n112 VSS 0.0126f
C5865 x4.X.n113 VSS 0.0589f
C5866 x4.X.n114 VSS 0.16f
C5867 x4.X.n115 VSS 0.126f
C5868 x4.X.n116 VSS 0.0047f
C5869 x4.X.t42 VSS 0.009f
C5870 x4.X.t64 VSS 0.0104f
C5871 x4.X.n117 VSS 0.0242f
C5872 x4.X.n118 VSS 0.00653f
C5873 x4.X.n119 VSS 0.00254f
C5874 x4.X.n120 VSS 0.0014f
C5875 x4.X.n121 VSS 0.0083f
C5876 x4.X.n122 VSS 0.0546f
C5877 x4.X.n123 VSS 0.00482f
C5878 x4.X.t41 VSS 0.00909f
C5879 x4.X.t38 VSS 0.0103f
C5880 x4.X.n124 VSS 0.0242f
C5881 x4.X.n125 VSS 0.00661f
C5882 x4.X.n126 VSS 0.00246f
C5883 x4.X.n127 VSS 0.0014f
C5884 x4.X.n128 VSS 0.00821f
C5885 x4.X.n129 VSS 0.0257f
C5886 x4.X.n130 VSS 0.0844f
C5887 x4.X.n131 VSS 0.125f
C5888 x4.X.n132 VSS 0.00271f
C5889 x4.X.n133 VSS 0.0014f
C5890 x4.X.t46 VSS 0.0103f
C5891 x4.X.t61 VSS 0.0087f
C5892 x4.X.n134 VSS 0.0117f
C5893 x4.X.n135 VSS 0.0126f
C5894 x4.X.n136 VSS 0.019f
C5895 x4.X.n137 VSS 0.00271f
C5896 x4.X.n138 VSS 0.0014f
C5897 x4.X.t65 VSS 0.0103f
C5898 x4.X.t43 VSS 0.00868f
C5899 x4.X.n139 VSS 0.0115f
C5900 x4.X.n140 VSS 0.0128f
C5901 x4.X.n141 VSS 0.0589f
C5902 x4.X.n142 VSS 0.161f
C5903 x4.X.n143 VSS 0.125f
C5904 x4.X.t56 VSS 0.009f
C5905 x4.X.t35 VSS 0.0104f
C5906 x4.X.n144 VSS 0.0242f
C5907 x4.X.n145 VSS 0.00631f
C5908 x4.X.n146 VSS 0.00271f
C5909 x4.X.n147 VSS 0.00141f
C5910 x4.X.n148 VSS 0.00518f
C5911 x4.X.n149 VSS 0.00686f
C5912 x4.X.n150 VSS 0.00893f
C5913 x4.X.n151 VSS 0.0541f
C5914 x4.X.t40 VSS 0.0105f
C5915 x4.X.t53 VSS 0.00892f
C5916 x4.X.n152 VSS 0.0242f
C5917 x4.X.n153 VSS 0.00639f
C5918 x4.X.n154 VSS 0.00263f
C5919 x4.X.n155 VSS 0.0014f
C5920 x4.X.n156 VSS 0.00482f
C5921 x4.X.n157 VSS 0.00769f
C5922 x4.X.n158 VSS 0.00848f
C5923 x4.X.n159 VSS 0.0259f
C5924 x4.X.n160 VSS 0.0851f
C5925 x4.X.n161 VSS 0.125f
C5926 x4.X.n162 VSS 0.00271f
C5927 x4.X.n163 VSS 0.0014f
C5928 x4.X.t48 VSS 0.0103f
C5929 x4.X.t62 VSS 0.00868f
C5930 x4.X.n164 VSS 0.0115f
C5931 x4.X.n165 VSS 0.0128f
C5932 x4.X.n166 VSS 0.0221f
C5933 x4.X.n167 VSS 0.00778f
C5934 x4.X.n168 VSS 0.0061f
C5935 x4.X.n169 VSS 0.00271f
C5936 x4.X.t47 VSS 0.009f
C5937 x4.X.t68 VSS 0.0103f
C5938 x4.X.n170 VSS 0.0128f
C5939 x4.X.n171 VSS 0.0112f
C5940 x4.X.n172 VSS 0.00148f
C5941 x4.X.n173 VSS 0.00507f
C5942 x4.X.n174 VSS 0.00813f
C5943 x4.X.n175 VSS 0.0698f
C5944 x4.X.n176 VSS 0.119f
C5945 x4.X.n177 VSS 0.103f
C5946 x4.X.t44 VSS 0.0104f
C5947 x4.X.t59 VSS 0.00899f
C5948 x4.X.n178 VSS 0.0239f
C5949 x4.X.n179 VSS 0.168f
C5950 x4.X.n180 VSS 0.304f
C5951 x4.X.n181 VSS 0.0328f
C5952 eob.t8 VSS 0.0308f
C5953 eob.t9 VSS 0.0193f
C5954 eob.n0 VSS 0.0589f
C5955 eob.t3 VSS 0.0186f
C5956 eob.t1 VSS 0.0186f
C5957 eob.n1 VSS 0.0543f
C5958 eob.t5 VSS 0.0121f
C5959 eob.t4 VSS 0.0121f
C5960 eob.n2 VSS 0.0362f
C5961 eob.n3 VSS 0.165f
C5962 eob.t0 VSS 0.0186f
C5963 eob.t2 VSS 0.0186f
C5964 eob.n4 VSS 0.0377f
C5965 eob.n5 VSS 0.0152f
C5966 eob.n6 VSS 0.0342f
C5967 eob.t7 VSS 0.0121f
C5968 eob.t6 VSS 0.0121f
C5969 eob.n7 VSS 0.0242f
C5970 eob.n8 VSS 0.0152f
C5971 eob.n9 VSS 0.0875f
C5972 eob.t11 VSS 0.025f
C5973 eob.t10 VSS 0.0174f
C5974 eob.n10 VSS 0.0508f
C5975 eob.n11 VSS 0.0192f
C5976 eob.n12 VSS 0.514f
C5977 eob.n13 VSS 0.519f
C5978 check[1].t0 VSS 0.046f
C5979 check[1].n0 VSS 0.00347f
C5980 check[1].t3 VSS 0.0153f
C5981 check[1].t2 VSS 0.0227f
C5982 check[1].n1 VSS 0.0487f
C5983 check[1].n2 VSS 0.582f
C5984 check[1].t5 VSS 0.0215f
C5985 check[1].t4 VSS 0.0149f
C5986 check[1].n3 VSS 0.0436f
C5987 check[1].n4 VSS 0.0165f
C5988 check[1].n5 VSS 0.733f
C5989 check[1].n6 VSS 0.0312f
C5990 check[1].n7 VSS 0.227f
C5991 check[1].t1 VSS 0.0177f
C5992 check[1].n8 VSS 0.0291f
C5993 VDD.n0 VSS 0.00118f
C5994 VDD.t537 VSS 3.92e-19
C5995 VDD.t406 VSS 3.92e-19
C5996 VDD.n1 VSS 8.47e-19
C5997 VDD.t536 VSS 0.00376f
C5998 VDD.n2 VSS 0.00507f
C5999 VDD.n3 VSS 7.09e-19
C6000 VDD.n4 VSS 0.00118f
C6001 VDD.t390 VSS 3.92e-19
C6002 VDD.t408 VSS 3.92e-19
C6003 VDD.n5 VSS 8.47e-19
C6004 VDD.t389 VSS 0.00376f
C6005 VDD.n6 VSS 0.00507f
C6006 VDD.n7 VSS 7.09e-19
C6007 VDD.n8 VSS 0.00118f
C6008 VDD.t521 VSS 3.92e-19
C6009 VDD.t623 VSS 3.92e-19
C6010 VDD.n9 VSS 8.47e-19
C6011 VDD.t520 VSS 0.00376f
C6012 VDD.n10 VSS 0.00507f
C6013 VDD.n11 VSS 7.09e-19
C6014 VDD.n12 VSS 0.002f
C6015 VDD.t696 VSS 5.19e-19
C6016 VDD.t49 VSS 5.19e-19
C6017 VDD.n13 VSS 0.00126f
C6018 VDD.n14 VSS 0.00238f
C6019 VDD.n15 VSS 0.00131f
C6020 VDD.n16 VSS 7.19e-19
C6021 VDD.n17 VSS 7.09e-19
C6022 VDD.n18 VSS 0.002f
C6023 VDD.t384 VSS 6.12e-19
C6024 VDD.t374 VSS 6.12e-19
C6025 VDD.n19 VSS 0.0014f
C6026 VDD.n20 VSS 0.00217f
C6027 VDD.n21 VSS 7.09e-19
C6028 VDD.t385 VSS 0.00381f
C6029 VDD.n22 VSS 7.09e-19
C6030 VDD.n23 VSS 6.7e-19
C6031 VDD.t386 VSS 6.12e-19
C6032 VDD.t382 VSS 6.12e-19
C6033 VDD.n24 VSS 0.00145f
C6034 VDD.n25 VSS 0.00249f
C6035 VDD.n26 VSS 4.73e-19
C6036 VDD.n27 VSS 3.54e-19
C6037 VDD.n28 VSS 0.00116f
C6038 VDD.n29 VSS 3.16e-19
C6039 VDD.n30 VSS 4.27e-19
C6040 VDD.t303 VSS 0.00243f
C6041 VDD.n31 VSS 0.00183f
C6042 VDD.n32 VSS 1.85e-19
C6043 VDD.n33 VSS 1.12e-19
C6044 VDD.n34 VSS 9.25e-19
C6045 VDD.n35 VSS 6.55e-20
C6046 VDD.t296 VSS 0.0031f
C6047 VDD.n36 VSS 3.28e-19
C6048 VDD.t293 VSS 6.12e-19
C6049 VDD.t297 VSS 6.12e-19
C6050 VDD.n37 VSS 0.00139f
C6051 VDD.n38 VSS 1.12e-19
C6052 VDD.n39 VSS 8.92e-19
C6053 VDD.n40 VSS 4.27e-19
C6054 VDD.n41 VSS 3.16e-19
C6055 VDD.n42 VSS 5.79e-19
C6056 VDD.n43 VSS 6.55e-20
C6057 VDD.n44 VSS 1.12e-19
C6058 VDD.n45 VSS 4.27e-19
C6059 VDD.n46 VSS 1.12e-19
C6060 VDD.n47 VSS 1.85e-19
C6061 VDD.n48 VSS 1.12e-19
C6062 VDD.t295 VSS 6.12e-19
C6063 VDD.t299 VSS 6.12e-19
C6064 VDD.n49 VSS 0.00139f
C6065 VDD.n50 VSS 3.28e-19
C6066 VDD.n51 VSS 0.00331f
C6067 VDD.n52 VSS 3.16e-19
C6068 VDD.n53 VSS 4.27e-19
C6069 VDD.n54 VSS 1.85e-19
C6070 VDD.n55 VSS 1.12e-19
C6071 VDD.n56 VSS 9.25e-19
C6072 VDD.n57 VSS 6.55e-20
C6073 VDD.t482 VSS 0.0031f
C6074 VDD.n58 VSS 3.28e-19
C6075 VDD.t483 VSS 6.12e-19
C6076 VDD.t301 VSS 6.12e-19
C6077 VDD.n59 VSS 0.00139f
C6078 VDD.n60 VSS 1.12e-19
C6079 VDD.n61 VSS 8.92e-19
C6080 VDD.n62 VSS 4.27e-19
C6081 VDD.n63 VSS 3.16e-19
C6082 VDD.n64 VSS 7.03e-19
C6083 VDD.n65 VSS 6.55e-20
C6084 VDD.n66 VSS 1.12e-19
C6085 VDD.n67 VSS 4.27e-19
C6086 VDD.n68 VSS 1.12e-19
C6087 VDD.n69 VSS 1.85e-19
C6088 VDD.n70 VSS 1.12e-19
C6089 VDD.t505 VSS 6.12e-19
C6090 VDD.t493 VSS 6.12e-19
C6091 VDD.n71 VSS 0.00139f
C6092 VDD.n72 VSS 3.28e-19
C6093 VDD.n73 VSS 0.00199f
C6094 VDD.n74 VSS 3.16e-19
C6095 VDD.n75 VSS 4.27e-19
C6096 VDD.n76 VSS 1.85e-19
C6097 VDD.t507 VSS 6.12e-19
C6098 VDD.t497 VSS 6.12e-19
C6099 VDD.n77 VSS 0.00139f
C6100 VDD.n78 VSS 0.00113f
C6101 VDD.n79 VSS 0.001f
C6102 VDD.n80 VSS 6.55e-20
C6103 VDD.t506 VSS 0.00269f
C6104 VDD.n81 VSS 2.89e-19
C6105 VDD.n82 VSS 1.77e-19
C6106 VDD.n83 VSS 0.002f
C6107 VDD.t511 VSS 6.12e-19
C6108 VDD.t499 VSS 6.12e-19
C6109 VDD.n84 VSS 0.00139f
C6110 VDD.n85 VSS 0.00167f
C6111 VDD.n86 VSS 6.05e-19
C6112 VDD.n87 VSS 1.04e-19
C6113 VDD.t490 VSS 0.00381f
C6114 VDD.n88 VSS 7.09e-19
C6115 VDD.t481 VSS 6.12e-19
C6116 VDD.t491 VSS 6.12e-19
C6117 VDD.n89 VSS 0.00139f
C6118 VDD.n90 VSS 0.00101f
C6119 VDD.n91 VSS 0.002f
C6120 VDD.n92 VSS 9.07e-19
C6121 VDD.n93 VSS 7.09e-19
C6122 VDD.n94 VSS 7.09e-19
C6123 VDD.t486 VSS 0.00381f
C6124 VDD.n95 VSS 7.09e-19
C6125 VDD.n96 VSS 8.02e-19
C6126 VDD.t509 VSS 6.12e-19
C6127 VDD.t503 VSS 6.12e-19
C6128 VDD.n97 VSS 0.00139f
C6129 VDD.n98 VSS 0.00167f
C6130 VDD.n99 VSS 0.002f
C6131 VDD.n100 VSS 6.97e-19
C6132 VDD.n101 VSS 7.09e-19
C6133 VDD.n102 VSS 0.00579f
C6134 VDD.n103 VSS 7.09e-19
C6135 VDD.n104 VSS 9.79e-19
C6136 VDD.t489 VSS 0.00227f
C6137 VDD.n105 VSS 0.00193f
C6138 VDD.n106 VSS 0.002f
C6139 VDD.t311 VSS 5.51e-19
C6140 VDD.t120 VSS -1.76e-19
C6141 VDD.n107 VSS 0.00259f
C6142 VDD.n108 VSS 7.18e-19
C6143 VDD.n109 VSS 0.00116f
C6144 VDD.n110 VSS 7.09e-19
C6145 VDD.t555 VSS 0.00381f
C6146 VDD.n111 VSS 7.09e-19
C6147 VDD.t556 VSS 5.95e-19
C6148 VDD.t307 VSS -3.29e-19
C6149 VDD.n112 VSS 0.00233f
C6150 VDD.n113 VSS 0.00159f
C6151 VDD.n114 VSS 0.002f
C6152 VDD.t141 VSS 0.0017f
C6153 VDD.n115 VSS 0.00171f
C6154 VDD.n116 VSS 0.00108f
C6155 VDD.n117 VSS 0.00414f
C6156 VDD.n118 VSS 7.09e-19
C6157 VDD.n119 VSS 0.00121f
C6158 VDD.n120 VSS 0.002f
C6159 VDD.n121 VSS 0.00121f
C6160 VDD.n122 VSS 7.09e-19
C6161 VDD.n123 VSS 0.00401f
C6162 VDD.n124 VSS 7.09e-19
C6163 VDD.t139 VSS 6.28e-19
C6164 VDD.t420 VSS 0.00141f
C6165 VDD.n125 VSS 0.00226f
C6166 VDD.n126 VSS 0.00297f
C6167 VDD.n127 VSS 0.002f
C6168 VDD.n128 VSS 7.62e-19
C6169 VDD.n129 VSS 7.09e-19
C6170 VDD.t417 VSS 0.00381f
C6171 VDD.n130 VSS 7.09e-19
C6172 VDD.n131 VSS 0.00116f
C6173 VDD.n132 VSS 0.002f
C6174 VDD.n133 VSS 9.79e-19
C6175 VDD.n134 VSS 7.09e-19
C6176 VDD.n135 VSS 0.00596f
C6177 VDD.n136 VSS 7.09e-19
C6178 VDD.n137 VSS 7.76e-19
C6179 VDD.t69 VSS 3.92e-19
C6180 VDD.t519 VSS 3.92e-19
C6181 VDD.n138 VSS 8.47e-19
C6182 VDD.n139 VSS 9.79e-19
C6183 VDD.n140 VSS 7.09e-19
C6184 VDD.t179 VSS 0.00381f
C6185 VDD.n141 VSS 7.18e-19
C6186 VDD.n142 VSS 0.0013f
C6187 VDD.n143 VSS 0.002f
C6188 VDD.n144 VSS 0.00116f
C6189 VDD.n145 VSS 7.09e-19
C6190 VDD.t645 VSS 0.00381f
C6191 VDD.n146 VSS 7.09e-19
C6192 VDD.t646 VSS 5.95e-19
C6193 VDD.t597 VSS -3.29e-19
C6194 VDD.n147 VSS 0.00233f
C6195 VDD.n148 VSS 0.00159f
C6196 VDD.n149 VSS 0.002f
C6197 VDD.t402 VSS 0.0017f
C6198 VDD.n150 VSS 0.00171f
C6199 VDD.n151 VSS 0.00108f
C6200 VDD.n152 VSS 0.00414f
C6201 VDD.n153 VSS 7.09e-19
C6202 VDD.n154 VSS 0.00121f
C6203 VDD.n155 VSS 0.002f
C6204 VDD.n156 VSS 0.00121f
C6205 VDD.n157 VSS 7.09e-19
C6206 VDD.n158 VSS 0.00401f
C6207 VDD.n159 VSS 7.09e-19
C6208 VDD.t404 VSS 6.28e-19
C6209 VDD.t574 VSS 0.00141f
C6210 VDD.n160 VSS 0.00226f
C6211 VDD.n161 VSS 0.00297f
C6212 VDD.n162 VSS 0.002f
C6213 VDD.n163 VSS 7.62e-19
C6214 VDD.n164 VSS 7.09e-19
C6215 VDD.t575 VSS 0.00381f
C6216 VDD.n165 VSS 7.09e-19
C6217 VDD.n166 VSS 0.00116f
C6218 VDD.n167 VSS 0.002f
C6219 VDD.n168 VSS 9.79e-19
C6220 VDD.n169 VSS 7.09e-19
C6221 VDD.n170 VSS 0.00596f
C6222 VDD.n171 VSS 7.09e-19
C6223 VDD.n172 VSS 7.76e-19
C6224 VDD.t71 VSS 3.92e-19
C6225 VDD.t107 VSS 3.92e-19
C6226 VDD.n173 VSS 8.47e-19
C6227 VDD.n174 VSS 9.79e-19
C6228 VDD.n175 VSS 7.09e-19
C6229 VDD.t265 VSS 0.00381f
C6230 VDD.n176 VSS 7.18e-19
C6231 VDD.n177 VSS 0.0013f
C6232 VDD.n178 VSS 0.002f
C6233 VDD.n179 VSS 0.00116f
C6234 VDD.n180 VSS 7.09e-19
C6235 VDD.t586 VSS 0.00381f
C6236 VDD.n181 VSS 7.09e-19
C6237 VDD.t587 VSS 5.95e-19
C6238 VDD.t173 VSS -3.29e-19
C6239 VDD.n182 VSS 0.00233f
C6240 VDD.n183 VSS 0.00159f
C6241 VDD.n184 VSS 0.002f
C6242 VDD.t111 VSS 0.0017f
C6243 VDD.n185 VSS 0.00171f
C6244 VDD.n186 VSS 0.00108f
C6245 VDD.n187 VSS 0.00414f
C6246 VDD.n188 VSS 7.09e-19
C6247 VDD.n189 VSS 0.00121f
C6248 VDD.n190 VSS 0.002f
C6249 VDD.n191 VSS 0.00121f
C6250 VDD.n192 VSS 7.09e-19
C6251 VDD.n193 VSS 0.00401f
C6252 VDD.n194 VSS 7.09e-19
C6253 VDD.t113 VSS 6.28e-19
C6254 VDD.t168 VSS 0.00141f
C6255 VDD.n195 VSS 0.00226f
C6256 VDD.n196 VSS 0.00297f
C6257 VDD.n197 VSS 0.002f
C6258 VDD.n198 VSS 7.62e-19
C6259 VDD.n199 VSS 7.09e-19
C6260 VDD.t165 VSS 0.00381f
C6261 VDD.n200 VSS 7.09e-19
C6262 VDD.n201 VSS 0.00116f
C6263 VDD.n202 VSS 0.002f
C6264 VDD.n203 VSS 9.79e-19
C6265 VDD.n204 VSS 7.09e-19
C6266 VDD.n205 VSS 0.00596f
C6267 VDD.n206 VSS 7.09e-19
C6268 VDD.n207 VSS 7.76e-19
C6269 VDD.t67 VSS 3.92e-19
C6270 VDD.t607 VSS 3.92e-19
C6271 VDD.n208 VSS 8.47e-19
C6272 VDD.n209 VSS 9.79e-19
C6273 VDD.n210 VSS 7.09e-19
C6274 VDD.t26 VSS 0.00381f
C6275 VDD.n211 VSS 7.18e-19
C6276 VDD.n212 VSS 0.0013f
C6277 VDD.n213 VSS 0.002f
C6278 VDD.n214 VSS 0.00116f
C6279 VDD.n215 VSS 7.09e-19
C6280 VDD.t275 VSS 0.00381f
C6281 VDD.n216 VSS 7.09e-19
C6282 VDD.t276 VSS 5.95e-19
C6283 VDD.t73 VSS -3.29e-19
C6284 VDD.n217 VSS 0.00233f
C6285 VDD.n218 VSS 0.00159f
C6286 VDD.n219 VSS 0.002f
C6287 VDD.t1 VSS 0.0017f
C6288 VDD.n220 VSS 0.00171f
C6289 VDD.n221 VSS 0.00108f
C6290 VDD.n222 VSS 0.00414f
C6291 VDD.n223 VSS 7.09e-19
C6292 VDD.n224 VSS 0.00121f
C6293 VDD.n225 VSS 0.002f
C6294 VDD.n226 VSS 0.00121f
C6295 VDD.n227 VSS 7.09e-19
C6296 VDD.n228 VSS 0.00401f
C6297 VDD.n229 VSS 7.09e-19
C6298 VDD.t3 VSS 6.28e-19
C6299 VDD.t368 VSS 0.00141f
C6300 VDD.n230 VSS 0.00226f
C6301 VDD.n231 VSS 0.00297f
C6302 VDD.n232 VSS 0.002f
C6303 VDD.n233 VSS 7.62e-19
C6304 VDD.n234 VSS 7.09e-19
C6305 VDD.t369 VSS 0.00381f
C6306 VDD.n235 VSS 7.09e-19
C6307 VDD.n236 VSS 0.00116f
C6308 VDD.n237 VSS 0.002f
C6309 VDD.n238 VSS 9.79e-19
C6310 VDD.n239 VSS 7.09e-19
C6311 VDD.n240 VSS 0.00596f
C6312 VDD.n241 VSS 7.09e-19
C6313 VDD.n242 VSS 7.76e-19
C6314 VDD.t625 VSS 3.92e-19
C6315 VDD.t471 VSS 3.92e-19
C6316 VDD.n243 VSS 8.47e-19
C6317 VDD.n244 VSS 7.19e-19
C6318 VDD.t470 VSS 0.00381f
C6319 VDD.n245 VSS 0.00347f
C6320 VDD.t624 VSS 0.00306f
C6321 VDD.n246 VSS 0.00253f
C6322 VDD.n247 VSS 9.94e-19
C6323 VDD.n248 VSS 0.00131f
C6324 VDD.n249 VSS 0.00176f
C6325 VDD.n250 VSS 0.00181f
C6326 VDD.n251 VSS 0.002f
C6327 VDD.n252 VSS 0.002f
C6328 VDD.t313 VSS 9.19e-19
C6329 VDD.n253 VSS 0.002f
C6330 VDD.n254 VSS 0.00132f
C6331 VDD.n255 VSS 7.19e-19
C6332 VDD.n256 VSS 0.00563f
C6333 VDD.t312 VSS 0.00381f
C6334 VDD.n257 VSS 0.00385f
C6335 VDD.t282 VSS 0.00381f
C6336 VDD.n258 VSS 0.00496f
C6337 VDD.t469 VSS 0.00381f
C6338 VDD.n259 VSS 0.00347f
C6339 VDD.n260 VSS 7.09e-19
C6340 VDD.n261 VSS 0.00121f
C6341 VDD.n262 VSS 0.002f
C6342 VDD.n263 VSS 0.002f
C6343 VDD.n264 VSS 0.002f
C6344 VDD.n265 VSS 0.002f
C6345 VDD.t370 VSS 3.52e-19
C6346 VDD.t244 VSS 3.71e-19
C6347 VDD.n266 VSS 7.74e-19
C6348 VDD.n267 VSS 0.0018f
C6349 VDD.n268 VSS 0.00133f
C6350 VDD.n269 VSS 7.19e-19
C6351 VDD.n270 VSS 0.00438f
C6352 VDD.t243 VSS 0.00381f
C6353 VDD.n271 VSS 0.00434f
C6354 VDD.t2 VSS 0.00368f
C6355 VDD.t29 VSS 0.0036f
C6356 VDD.n272 VSS 0.00393f
C6357 VDD.n273 VSS 7.09e-19
C6358 VDD.n274 VSS 0.00121f
C6359 VDD.n275 VSS 6.7e-19
C6360 VDD.n276 VSS 0.002f
C6361 VDD.n277 VSS 0.002f
C6362 VDD.n278 VSS 7.1e-19
C6363 VDD.n279 VSS 7.09e-19
C6364 VDD.n280 VSS 0.00546f
C6365 VDD.t367 VSS 0.00381f
C6366 VDD.n281 VSS 0.00596f
C6367 VDD.t281 VSS 0.00381f
C6368 VDD.t468 VSS 0.00728f
C6369 VDD.n282 VSS 7.09e-19
C6370 VDD.n283 VSS 0.00121f
C6371 VDD.n284 VSS 0.002f
C6372 VDD.n285 VSS 0.002f
C6373 VDD.n286 VSS 0.002f
C6374 VDD.n287 VSS 1.27e-19
C6375 VDD.t739 VSS 4.1e-19
C6376 VDD.t242 VSS 9.69e-19
C6377 VDD.n288 VSS 0.00202f
C6378 VDD.n289 VSS 3.45e-19
C6379 VDD.n290 VSS 6.83e-19
C6380 VDD.n291 VSS 0.00252f
C6381 VDD.n292 VSS 4.01e-19
C6382 VDD.n293 VSS 3.6e-19
C6383 VDD.t735 VSS 4.04e-19
C6384 VDD.n294 VSS 2.92e-19
C6385 VDD.n295 VSS 6.21e-19
C6386 VDD.n296 VSS 0.00128f
C6387 VDD.t215 VSS 0.00151f
C6388 VDD.n297 VSS 0.00114f
C6389 VDD.t75 VSS 3.71e-19
C6390 VDD.t217 VSS 3.71e-19
C6391 VDD.n298 VSS 7.82e-19
C6392 VDD.n299 VSS 0.002f
C6393 VDD.n300 VSS 0.00102f
C6394 VDD.n301 VSS 9.79e-19
C6395 VDD.n302 VSS 0.002f
C6396 VDD.n303 VSS 0.002f
C6397 VDD.n304 VSS 0.00167f
C6398 VDD.n305 VSS 9.38e-19
C6399 VDD.n306 VSS 8.61e-19
C6400 VDD.n307 VSS 9.09e-19
C6401 VDD.n308 VSS 0.00455f
C6402 VDD.t74 VSS 0.00521f
C6403 VDD.t216 VSS 0.00844f
C6404 VDD.t350 VSS 0.0062f
C6405 VDD.n309 VSS 0.00298f
C6406 VDD.t0 VSS 0.00381f
C6407 VDD.n310 VSS 0.00513f
C6408 VDD.n311 VSS 0.00687f
C6409 VDD.n312 VSS 7.09e-19
C6410 VDD.n313 VSS 0.00188f
C6411 VDD.n314 VSS 0.00272f
C6412 VDD.n315 VSS 0.002f
C6413 VDD.n316 VSS 0.002f
C6414 VDD.n317 VSS 0.00121f
C6415 VDD.n318 VSS 7.09e-19
C6416 VDD.n319 VSS 0.00401f
C6417 VDD.t72 VSS 0.00381f
C6418 VDD.n320 VSS 0.00608f
C6419 VDD.n321 VSS 0.00393f
C6420 VDD.t76 VSS 0.00381f
C6421 VDD.n322 VSS 0.0055f
C6422 VDD.n323 VSS 7.09e-19
C6423 VDD.n324 VSS 0.00105f
C6424 VDD.n325 VSS 0.002f
C6425 VDD.t77 VSS 5.51e-19
C6426 VDD.t27 VSS -1.76e-19
C6427 VDD.n326 VSS 0.00259f
C6428 VDD.n327 VSS 0.00235f
C6429 VDD.n328 VSS 0.002f
C6430 VDD.n329 VSS 6.96e-19
C6431 VDD.n330 VSS 0.0015f
C6432 VDD.n331 VSS 9.79e-19
C6433 VDD.n332 VSS 7.09e-19
C6434 VDD.n333 VSS 0.00579f
C6435 VDD.n334 VSS 0.00385f
C6436 VDD.t66 VSS 0.00306f
C6437 VDD.t606 VSS 0.00381f
C6438 VDD.n335 VSS 0.00347f
C6439 VDD.n336 VSS 7.19e-19
C6440 VDD.n337 VSS 0.00131f
C6441 VDD.n338 VSS 0.00176f
C6442 VDD.n339 VSS 0.00181f
C6443 VDD.n340 VSS 0.002f
C6444 VDD.n341 VSS 0.002f
C6445 VDD.t318 VSS 9.19e-19
C6446 VDD.n342 VSS 0.002f
C6447 VDD.n343 VSS 0.00132f
C6448 VDD.n344 VSS 7.19e-19
C6449 VDD.n345 VSS 0.00563f
C6450 VDD.t317 VSS 0.00381f
C6451 VDD.n346 VSS 0.00385f
C6452 VDD.t372 VSS 0.00381f
C6453 VDD.n347 VSS 0.00496f
C6454 VDD.t609 VSS 0.00381f
C6455 VDD.n348 VSS 0.00347f
C6456 VDD.n349 VSS 7.09e-19
C6457 VDD.n350 VSS 0.00121f
C6458 VDD.n351 VSS 0.002f
C6459 VDD.n352 VSS 0.002f
C6460 VDD.n353 VSS 0.002f
C6461 VDD.n354 VSS 0.002f
C6462 VDD.t166 VSS 3.52e-19
C6463 VDD.t247 VSS 3.71e-19
C6464 VDD.n355 VSS 7.74e-19
C6465 VDD.n356 VSS 0.0018f
C6466 VDD.n357 VSS 0.00133f
C6467 VDD.n358 VSS 7.19e-19
C6468 VDD.n359 VSS 0.00438f
C6469 VDD.t246 VSS 0.00381f
C6470 VDD.n360 VSS 0.00434f
C6471 VDD.t112 VSS 0.00368f
C6472 VDD.t456 VSS 0.0036f
C6473 VDD.n361 VSS 0.00393f
C6474 VDD.n362 VSS 7.09e-19
C6475 VDD.n363 VSS 0.00121f
C6476 VDD.n364 VSS 6.7e-19
C6477 VDD.n365 VSS 0.002f
C6478 VDD.n366 VSS 0.002f
C6479 VDD.n367 VSS 7.1e-19
C6480 VDD.n368 VSS 7.09e-19
C6481 VDD.n369 VSS 0.00546f
C6482 VDD.t167 VSS 0.00381f
C6483 VDD.n370 VSS 0.00596f
C6484 VDD.t371 VSS 0.00381f
C6485 VDD.t608 VSS 0.00728f
C6486 VDD.n371 VSS 7.09e-19
C6487 VDD.n372 VSS 0.00121f
C6488 VDD.n373 VSS 0.002f
C6489 VDD.n374 VSS 0.002f
C6490 VDD.n375 VSS 0.002f
C6491 VDD.n376 VSS 1.27e-19
C6492 VDD.t727 VSS 4.1e-19
C6493 VDD.t245 VSS 9.69e-19
C6494 VDD.n377 VSS 0.00202f
C6495 VDD.n378 VSS 3.45e-19
C6496 VDD.n379 VSS 6.83e-19
C6497 VDD.n380 VSS 0.00252f
C6498 VDD.n381 VSS 4.01e-19
C6499 VDD.n382 VSS 3.6e-19
C6500 VDD.t726 VSS 4.04e-19
C6501 VDD.n383 VSS 2.92e-19
C6502 VDD.n384 VSS 6.21e-19
C6503 VDD.n385 VSS 0.00128f
C6504 VDD.t239 VSS 0.00151f
C6505 VDD.n386 VSS 0.00114f
C6506 VDD.t175 VSS 3.71e-19
C6507 VDD.t241 VSS 3.71e-19
C6508 VDD.n387 VSS 7.82e-19
C6509 VDD.n388 VSS 0.002f
C6510 VDD.n389 VSS 0.00102f
C6511 VDD.n390 VSS 9.79e-19
C6512 VDD.n391 VSS 0.002f
C6513 VDD.n392 VSS 0.002f
C6514 VDD.n393 VSS 0.00167f
C6515 VDD.n394 VSS 9.38e-19
C6516 VDD.n395 VSS 8.61e-19
C6517 VDD.n396 VSS 9.09e-19
C6518 VDD.n397 VSS 0.00455f
C6519 VDD.t174 VSS 0.00521f
C6520 VDD.t240 VSS 0.00844f
C6521 VDD.t181 VSS 0.0062f
C6522 VDD.n398 VSS 0.00298f
C6523 VDD.t110 VSS 0.00381f
C6524 VDD.n399 VSS 0.00513f
C6525 VDD.n400 VSS 0.00687f
C6526 VDD.n401 VSS 7.09e-19
C6527 VDD.n402 VSS 0.00188f
C6528 VDD.n403 VSS 0.00272f
C6529 VDD.n404 VSS 0.002f
C6530 VDD.n405 VSS 0.002f
C6531 VDD.n406 VSS 0.00121f
C6532 VDD.n407 VSS 7.09e-19
C6533 VDD.n408 VSS 0.00401f
C6534 VDD.t172 VSS 0.00381f
C6535 VDD.n409 VSS 0.00608f
C6536 VDD.n410 VSS 0.00393f
C6537 VDD.t176 VSS 0.00381f
C6538 VDD.n411 VSS 0.0055f
C6539 VDD.n412 VSS 7.09e-19
C6540 VDD.n413 VSS 0.00105f
C6541 VDD.n414 VSS 0.002f
C6542 VDD.t177 VSS 5.51e-19
C6543 VDD.t266 VSS -1.76e-19
C6544 VDD.n415 VSS 0.00259f
C6545 VDD.n416 VSS 0.00235f
C6546 VDD.n417 VSS 0.002f
C6547 VDD.n418 VSS 6.96e-19
C6548 VDD.n419 VSS 0.0015f
C6549 VDD.n420 VSS 9.79e-19
C6550 VDD.n421 VSS 7.09e-19
C6551 VDD.n422 VSS 0.00579f
C6552 VDD.n423 VSS 0.00385f
C6553 VDD.t70 VSS 0.00306f
C6554 VDD.t106 VSS 0.00381f
C6555 VDD.n424 VSS 0.00347f
C6556 VDD.n425 VSS 7.19e-19
C6557 VDD.n426 VSS 0.00131f
C6558 VDD.n427 VSS 0.00176f
C6559 VDD.n428 VSS 0.00181f
C6560 VDD.n429 VSS 0.002f
C6561 VDD.n430 VSS 0.002f
C6562 VDD.t445 VSS 9.19e-19
C6563 VDD.n431 VSS 0.002f
C6564 VDD.n432 VSS 0.00132f
C6565 VDD.n433 VSS 7.19e-19
C6566 VDD.n434 VSS 0.00563f
C6567 VDD.t444 VSS 0.00381f
C6568 VDD.n435 VSS 0.00385f
C6569 VDD.t572 VSS 0.00381f
C6570 VDD.n436 VSS 0.00496f
C6571 VDD.t105 VSS 0.00381f
C6572 VDD.n437 VSS 0.00347f
C6573 VDD.n438 VSS 7.09e-19
C6574 VDD.n439 VSS 0.00121f
C6575 VDD.n440 VSS 0.002f
C6576 VDD.n441 VSS 0.002f
C6577 VDD.n442 VSS 0.002f
C6578 VDD.n443 VSS 0.002f
C6579 VDD.t576 VSS 3.52e-19
C6580 VDD.t226 VSS 3.71e-19
C6581 VDD.n444 VSS 7.74e-19
C6582 VDD.n445 VSS 0.0018f
C6583 VDD.n446 VSS 0.00133f
C6584 VDD.n447 VSS 7.19e-19
C6585 VDD.n448 VSS 0.00438f
C6586 VDD.t225 VSS 0.00381f
C6587 VDD.n449 VSS 0.00434f
C6588 VDD.t403 VSS 0.00368f
C6589 VDD.t388 VSS 0.0036f
C6590 VDD.n450 VSS 0.00393f
C6591 VDD.n451 VSS 7.09e-19
C6592 VDD.n452 VSS 0.00121f
C6593 VDD.n453 VSS 6.7e-19
C6594 VDD.n454 VSS 0.002f
C6595 VDD.n455 VSS 0.002f
C6596 VDD.n456 VSS 7.1e-19
C6597 VDD.n457 VSS 7.09e-19
C6598 VDD.n458 VSS 0.00546f
C6599 VDD.t573 VSS 0.00381f
C6600 VDD.n459 VSS 0.00596f
C6601 VDD.t571 VSS 0.00381f
C6602 VDD.t104 VSS 0.00728f
C6603 VDD.n460 VSS 7.09e-19
C6604 VDD.n461 VSS 0.00121f
C6605 VDD.n462 VSS 0.002f
C6606 VDD.n463 VSS 0.002f
C6607 VDD.n464 VSS 0.002f
C6608 VDD.n465 VSS 1.27e-19
C6609 VDD.t733 VSS 4.1e-19
C6610 VDD.t224 VSS 9.69e-19
C6611 VDD.n466 VSS 0.00202f
C6612 VDD.n467 VSS 3.45e-19
C6613 VDD.n468 VSS 6.83e-19
C6614 VDD.n469 VSS 0.00252f
C6615 VDD.n470 VSS 4.01e-19
C6616 VDD.n471 VSS 3.6e-19
C6617 VDD.t728 VSS 4.04e-19
C6618 VDD.n472 VSS 2.92e-19
C6619 VDD.n473 VSS 6.21e-19
C6620 VDD.n474 VSS 0.00128f
C6621 VDD.t236 VSS 0.00151f
C6622 VDD.n475 VSS 0.00114f
C6623 VDD.t599 VSS 3.71e-19
C6624 VDD.t238 VSS 3.71e-19
C6625 VDD.n476 VSS 7.82e-19
C6626 VDD.n477 VSS 0.002f
C6627 VDD.n478 VSS 0.00102f
C6628 VDD.n479 VSS 9.79e-19
C6629 VDD.n480 VSS 0.002f
C6630 VDD.n481 VSS 0.002f
C6631 VDD.n482 VSS 0.00167f
C6632 VDD.n483 VSS 9.38e-19
C6633 VDD.n484 VSS 8.61e-19
C6634 VDD.n485 VSS 9.09e-19
C6635 VDD.n486 VSS 0.00455f
C6636 VDD.t598 VSS 0.00521f
C6637 VDD.t237 VSS 0.00844f
C6638 VDD.t323 VSS 0.0062f
C6639 VDD.n487 VSS 0.00298f
C6640 VDD.t401 VSS 0.00381f
C6641 VDD.n488 VSS 0.00513f
C6642 VDD.n489 VSS 0.00687f
C6643 VDD.n490 VSS 7.09e-19
C6644 VDD.n491 VSS 0.00188f
C6645 VDD.n492 VSS 0.00272f
C6646 VDD.n493 VSS 0.002f
C6647 VDD.n494 VSS 0.002f
C6648 VDD.n495 VSS 0.00121f
C6649 VDD.n496 VSS 7.09e-19
C6650 VDD.n497 VSS 0.00401f
C6651 VDD.t596 VSS 0.00381f
C6652 VDD.n498 VSS 0.00608f
C6653 VDD.n499 VSS 0.00393f
C6654 VDD.t600 VSS 0.00381f
C6655 VDD.n500 VSS 0.0055f
C6656 VDD.n501 VSS 7.09e-19
C6657 VDD.n502 VSS 0.00105f
C6658 VDD.n503 VSS 0.002f
C6659 VDD.t601 VSS 5.51e-19
C6660 VDD.t180 VSS -1.76e-19
C6661 VDD.n504 VSS 0.00259f
C6662 VDD.n505 VSS 0.00235f
C6663 VDD.n506 VSS 0.002f
C6664 VDD.n507 VSS 6.96e-19
C6665 VDD.n508 VSS 0.0015f
C6666 VDD.n509 VSS 9.79e-19
C6667 VDD.n510 VSS 7.09e-19
C6668 VDD.n511 VSS 0.00579f
C6669 VDD.n512 VSS 0.00385f
C6670 VDD.t68 VSS 0.00306f
C6671 VDD.t518 VSS 0.00381f
C6672 VDD.n513 VSS 0.00347f
C6673 VDD.n514 VSS 7.19e-19
C6674 VDD.n515 VSS 0.00131f
C6675 VDD.n516 VSS 0.00176f
C6676 VDD.n517 VSS 0.00181f
C6677 VDD.n518 VSS 0.002f
C6678 VDD.n519 VSS 0.002f
C6679 VDD.t439 VSS 9.19e-19
C6680 VDD.n520 VSS 0.002f
C6681 VDD.n521 VSS 0.00132f
C6682 VDD.n522 VSS 7.19e-19
C6683 VDD.n523 VSS 0.00563f
C6684 VDD.t438 VSS 0.00381f
C6685 VDD.n524 VSS 0.00385f
C6686 VDD.t130 VSS 0.00381f
C6687 VDD.n525 VSS 0.00496f
C6688 VDD.t517 VSS 0.00381f
C6689 VDD.n526 VSS 0.00347f
C6690 VDD.n527 VSS 7.09e-19
C6691 VDD.n528 VSS 0.00121f
C6692 VDD.n529 VSS 0.002f
C6693 VDD.n530 VSS 0.002f
C6694 VDD.n531 VSS 0.002f
C6695 VDD.n532 VSS 0.002f
C6696 VDD.t418 VSS 3.52e-19
C6697 VDD.t211 VSS 3.71e-19
C6698 VDD.n533 VSS 7.74e-19
C6699 VDD.n534 VSS 0.0018f
C6700 VDD.n535 VSS 0.00133f
C6701 VDD.n536 VSS 7.19e-19
C6702 VDD.n537 VSS 0.00438f
C6703 VDD.t210 VSS 0.00381f
C6704 VDD.n538 VSS 0.00434f
C6705 VDD.t138 VSS 0.00368f
C6706 VDD.t642 VSS 0.0036f
C6707 VDD.n539 VSS 0.00393f
C6708 VDD.n540 VSS 7.09e-19
C6709 VDD.n541 VSS 0.00121f
C6710 VDD.n542 VSS 6.7e-19
C6711 VDD.n543 VSS 0.002f
C6712 VDD.n544 VSS 0.002f
C6713 VDD.n545 VSS 7.1e-19
C6714 VDD.n546 VSS 7.09e-19
C6715 VDD.n547 VSS 0.00546f
C6716 VDD.t419 VSS 0.00381f
C6717 VDD.n548 VSS 0.00596f
C6718 VDD.t131 VSS 0.00381f
C6719 VDD.t516 VSS 0.00728f
C6720 VDD.n549 VSS 7.09e-19
C6721 VDD.n550 VSS 0.00121f
C6722 VDD.n551 VSS 0.002f
C6723 VDD.n552 VSS 0.002f
C6724 VDD.n553 VSS 0.002f
C6725 VDD.n554 VSS 1.27e-19
C6726 VDD.t738 VSS 4.1e-19
C6727 VDD.t209 VSS 9.69e-19
C6728 VDD.n555 VSS 0.00202f
C6729 VDD.n556 VSS 3.45e-19
C6730 VDD.n557 VSS 6.83e-19
C6731 VDD.n558 VSS 0.00252f
C6732 VDD.n559 VSS 4.01e-19
C6733 VDD.n560 VSS 3.6e-19
C6734 VDD.t734 VSS 4.04e-19
C6735 VDD.n561 VSS 2.92e-19
C6736 VDD.n562 VSS 6.21e-19
C6737 VDD.n563 VSS 0.00128f
C6738 VDD.t218 VSS 0.00151f
C6739 VDD.n564 VSS 0.00114f
C6740 VDD.t309 VSS 3.71e-19
C6741 VDD.t220 VSS 3.71e-19
C6742 VDD.n565 VSS 7.82e-19
C6743 VDD.n566 VSS 0.002f
C6744 VDD.n567 VSS 0.00102f
C6745 VDD.n568 VSS 9.79e-19
C6746 VDD.n569 VSS 0.002f
C6747 VDD.n570 VSS 0.002f
C6748 VDD.n571 VSS 0.00167f
C6749 VDD.n572 VSS 9.38e-19
C6750 VDD.n573 VSS 8.61e-19
C6751 VDD.n574 VSS 9.09e-19
C6752 VDD.n575 VSS 0.00455f
C6753 VDD.t308 VSS 0.00521f
C6754 VDD.t219 VSS 0.00844f
C6755 VDD.t171 VSS 0.0062f
C6756 VDD.n576 VSS 0.00298f
C6757 VDD.t140 VSS 0.00381f
C6758 VDD.n577 VSS 0.00513f
C6759 VDD.n578 VSS 0.00687f
C6760 VDD.n579 VSS 7.09e-19
C6761 VDD.n580 VSS 0.00188f
C6762 VDD.n581 VSS 0.00272f
C6763 VDD.n582 VSS 0.002f
C6764 VDD.n583 VSS 0.002f
C6765 VDD.n584 VSS 0.002f
C6766 VDD.n585 VSS 0.00121f
C6767 VDD.n586 VSS 7.09e-19
C6768 VDD.n587 VSS 0.00401f
C6769 VDD.t306 VSS 0.00381f
C6770 VDD.n588 VSS 0.00608f
C6771 VDD.t119 VSS 0.00381f
C6772 VDD.n589 VSS 0.00393f
C6773 VDD.t310 VSS 0.00381f
C6774 VDD.n590 VSS 0.0055f
C6775 VDD.n591 VSS 7.09e-19
C6776 VDD.n592 VSS 0.00105f
C6777 VDD.n593 VSS 0.0013f
C6778 VDD.n594 VSS 0.00235f
C6779 VDD.n595 VSS 0.002f
C6780 VDD.n596 VSS 0.0015f
C6781 VDD.n597 VSS 0.0015f
C6782 VDD.n598 VSS 0.00112f
C6783 VDD.n599 VSS 7.09e-19
C6784 VDD.n600 VSS 0.00761f
C6785 VDD.n601 VSS 0.00496f
C6786 VDD.t488 VSS 0.00381f
C6787 VDD.n602 VSS 0.00347f
C6788 VDD.t500 VSS 0.00381f
C6789 VDD.n603 VSS 0.00347f
C6790 VDD.n604 VSS 7.09e-19
C6791 VDD.t501 VSS 6.12e-19
C6792 VDD.t487 VSS 6.12e-19
C6793 VDD.n605 VSS 0.00139f
C6794 VDD.n606 VSS 0.00167f
C6795 VDD.n607 VSS 0.00101f
C6796 VDD.n608 VSS 0.002f
C6797 VDD.n609 VSS 0.002f
C6798 VDD.n610 VSS 0.002f
C6799 VDD.n611 VSS 9.07e-19
C6800 VDD.n612 VSS 7.09e-19
C6801 VDD.n613 VSS 0.00347f
C6802 VDD.t508 VSS 0.00364f
C6803 VDD.t502 VSS 0.00364f
C6804 VDD.n614 VSS 0.00347f
C6805 VDD.t484 VSS 0.00381f
C6806 VDD.n615 VSS 0.00347f
C6807 VDD.t480 VSS 0.00381f
C6808 VDD.n616 VSS 0.00347f
C6809 VDD.t494 VSS 0.00381f
C6810 VDD.n617 VSS 0.00347f
C6811 VDD.n618 VSS 7.09e-19
C6812 VDD.t485 VSS 6.12e-19
C6813 VDD.t495 VSS 6.12e-19
C6814 VDD.n619 VSS 0.00139f
C6815 VDD.n620 VSS 0.00167f
C6816 VDD.n621 VSS 8.02e-19
C6817 VDD.n622 VSS 0.002f
C6818 VDD.n623 VSS 0.002f
C6819 VDD.n624 VSS 0.002f
C6820 VDD.n625 VSS 6.97e-19
C6821 VDD.n626 VSS 0.00167f
C6822 VDD.n627 VSS 0.0011f
C6823 VDD.n628 VSS 7.09e-19
C6824 VDD.n629 VSS 0.00347f
C6825 VDD.t510 VSS 0.00381f
C6826 VDD.n630 VSS 0.00347f
C6827 VDD.t498 VSS 0.00269f
C6828 VDD.n631 VSS 0.00174f
C6829 VDD.n632 VSS 0.00112f
C6830 VDD.n633 VSS 0.00174f
C6831 VDD.n634 VSS 3.16e-19
C6832 VDD.n635 VSS 5.39e-19
C6833 VDD.n636 VSS 4.4e-19
C6834 VDD.n637 VSS 0.002f
C6835 VDD.n638 VSS 0.00189f
C6836 VDD.n639 VSS 4.93e-19
C6837 VDD.n640 VSS 5.92e-20
C6838 VDD.n641 VSS 4.73e-19
C6839 VDD.n642 VSS 2.77e-19
C6840 VDD.n643 VSS 0.00165f
C6841 VDD.n644 VSS 7.03e-19
C6842 VDD.t496 VSS 0.0031f
C6843 VDD.n645 VSS 0.00182f
C6844 VDD.n646 VSS 3.28e-19
C6845 VDD.n647 VSS 1.18e-19
C6846 VDD.n648 VSS 1.12e-19
C6847 VDD.n649 VSS 4.27e-19
C6848 VDD.n650 VSS 8.92e-19
C6849 VDD.n651 VSS 9.25e-19
C6850 VDD.n652 VSS 1.31e-19
C6851 VDD.n653 VSS 1.12e-19
C6852 VDD.n654 VSS 6.55e-20
C6853 VDD.n655 VSS 7.03e-19
C6854 VDD.n656 VSS 0.00149f
C6855 VDD.t504 VSS 0.0031f
C6856 VDD.n657 VSS 0.00232f
C6857 VDD.n658 VSS 3.16e-19
C6858 VDD.n659 VSS 9.2e-20
C6859 VDD.n660 VSS 0.00145f
C6860 VDD.n661 VSS 3.81e-19
C6861 VDD.n662 VSS 8.92e-19
C6862 VDD.n663 VSS 1.85e-19
C6863 VDD.n664 VSS 9.25e-19
C6864 VDD.n665 VSS 1.31e-19
C6865 VDD.n666 VSS 3.28e-19
C6866 VDD.n667 VSS 0.00116f
C6867 VDD.t492 VSS 0.0031f
C6868 VDD.n668 VSS 0.00265f
C6869 VDD.n669 VSS 8.27e-19
C6870 VDD.n670 VSS 7.03e-19
C6871 VDD.n671 VSS 6.55e-20
C6872 VDD.n672 VSS 1.12e-19
C6873 VDD.n673 VSS 1.31e-19
C6874 VDD.n674 VSS 9.25e-19
C6875 VDD.n675 VSS 1.85e-19
C6876 VDD.n676 VSS 8.92e-19
C6877 VDD.n677 VSS 2.76e-19
C6878 VDD.n678 VSS 0.00145f
C6879 VDD.n679 VSS 1.97e-19
C6880 VDD.n680 VSS 3.16e-19
C6881 VDD.n681 VSS 0.00298f
C6882 VDD.n682 VSS 7.03e-19
C6883 VDD.t300 VSS 0.0031f
C6884 VDD.n683 VSS 4.96e-19
C6885 VDD.n684 VSS 3.28e-19
C6886 VDD.n685 VSS 1.31e-19
C6887 VDD.n686 VSS 1.12e-19
C6888 VDD.n687 VSS 4.27e-19
C6889 VDD.n688 VSS 8.92e-19
C6890 VDD.n689 VSS 9.25e-19
C6891 VDD.n690 VSS 1.31e-19
C6892 VDD.n691 VSS 1.12e-19
C6893 VDD.n692 VSS 6.55e-20
C6894 VDD.n693 VSS 4.55e-19
C6895 VDD.t294 VSS 4.14e-19
C6896 VDD.n694 VSS 0.00335f
C6897 VDD.t298 VSS 2.89e-19
C6898 VDD.n695 VSS 0.00323f
C6899 VDD.n696 VSS 3.16e-19
C6900 VDD.n697 VSS 3.02e-19
C6901 VDD.n698 VSS 0.00145f
C6902 VDD.n699 VSS 1.71e-19
C6903 VDD.n700 VSS 8.92e-19
C6904 VDD.n701 VSS 1.85e-19
C6905 VDD.n702 VSS 9.25e-19
C6906 VDD.n703 VSS 1.31e-19
C6907 VDD.n704 VSS 3.28e-19
C6908 VDD.n705 VSS 0.00331f
C6909 VDD.t292 VSS 0.0031f
C6910 VDD.n706 VSS 4.96e-19
C6911 VDD.n707 VSS 0.00298f
C6912 VDD.n708 VSS 7.03e-19
C6913 VDD.n709 VSS 6.55e-20
C6914 VDD.n710 VSS 1.12e-19
C6915 VDD.n711 VSS 1.31e-19
C6916 VDD.n712 VSS 9.25e-19
C6917 VDD.n713 VSS 1.85e-19
C6918 VDD.n714 VSS 8.92e-19
C6919 VDD.n715 VSS 6.57e-20
C6920 VDD.n716 VSS 0.00145f
C6921 VDD.n717 VSS 4.08e-19
C6922 VDD.n718 VSS 3.16e-19
C6923 VDD.n719 VSS 8.27e-19
C6924 VDD.n720 VSS 7.03e-19
C6925 VDD.t302 VSS 0.0031f
C6926 VDD.n721 VSS 0.00265f
C6927 VDD.n722 VSS 3.28e-19
C6928 VDD.n723 VSS 1.31e-19
C6929 VDD.n724 VSS 1.12e-19
C6930 VDD.n725 VSS 4.27e-19
C6931 VDD.n726 VSS 8.92e-19
C6932 VDD.n727 VSS 1.74e-19
C6933 VDD.n728 VSS 8.55e-20
C6934 VDD.n729 VSS 1.85e-19
C6935 VDD.n730 VSS 9.25e-19
C6936 VDD.n731 VSS 9.2e-20
C6937 VDD.n732 VSS 1.12e-19
C6938 VDD.n733 VSS 6.55e-20
C6939 VDD.n734 VSS 7.03e-19
C6940 VDD.n735 VSS 0.00149f
C6941 VDD.n736 VSS 0.00347f
C6942 VDD.t379 VSS 0.00381f
C6943 VDD.n737 VSS 0.00546f
C6944 VDD.n738 VSS 6.7e-19
C6945 VDD.t380 VSS 0.00256f
C6946 VDD.n739 VSS 0.00428f
C6947 VDD.n740 VSS 4.34e-19
C6948 VDD.n741 VSS 0.00128f
C6949 VDD.n742 VSS 0.002f
C6950 VDD.n743 VSS 0.002f
C6951 VDD.n744 VSS 0.002f
C6952 VDD.n745 VSS 8.41e-19
C6953 VDD.n746 VSS 0.00131f
C6954 VDD.n747 VSS 7.19e-19
C6955 VDD.n748 VSS 0.00347f
C6956 VDD.t381 VSS 0.00381f
C6957 VDD.n749 VSS 0.00347f
C6958 VDD.t383 VSS 0.00381f
C6959 VDD.n750 VSS 0.00265f
C6960 VDD.t373 VSS 0.00381f
C6961 VDD.n751 VSS 0.00347f
C6962 VDD.n752 VSS 7.09e-19
C6963 VDD.n753 VSS 6.38e-19
C6964 VDD.n754 VSS 7.1e-19
C6965 VDD.n755 VSS 0.0015f
C6966 VDD.n756 VSS 0.0015f
C6967 VDD.n757 VSS 8.87e-19
C6968 VDD.n758 VSS 7.09e-19
C6969 VDD.n759 VSS 0.00513f
C6970 VDD.t695 VSS 0.00381f
C6971 VDD.n760 VSS 0.00364f
C6972 VDD.t48 VSS 0.00381f
C6973 VDD.n761 VSS 0.00269f
C6974 VDD.n762 VSS 7.09e-19
C6975 VDD.n763 VSS 5e-19
C6976 VDD.n764 VSS 0.0015f
C6977 VDD.n765 VSS 0.002f
C6978 VDD.t196 VSS 0.00241f
C6979 VDD.n766 VSS 0.00272f
C6980 VDD.n767 VSS 7.09e-19
C6981 VDD.n768 VSS 3.54e-19
C6982 VDD.n769 VSS 4.8e-19
C6983 VDD.n770 VSS 9.27e-19
C6984 VDD.n771 VSS 9.14e-19
C6985 VDD.n772 VSS 2.5e-19
C6986 VDD.n773 VSS 3.16e-19
C6987 VDD.n774 VSS 7.09e-19
C6988 VDD.n775 VSS 7.5e-20
C6989 VDD.n776 VSS 4.01e-19
C6990 VDD.n777 VSS 9.03e-19
C6991 VDD.n778 VSS 9.14e-19
C6992 VDD.n779 VSS 3.28e-19
C6993 VDD.n780 VSS 0.00342f
C6994 VDD.n781 VSS 3.16e-19
C6995 VDD.n782 VSS 2.5e-19
C6996 VDD.n783 VSS 1.12e-19
C6997 VDD.n784 VSS 1.85e-19
C6998 VDD.n785 VSS 3.75e-19
C6999 VDD.n787 VSS 9.14e-19
C7000 VDD.n788 VSS 3.28e-19
C7001 VDD.n789 VSS 7.5e-20
C7002 VDD.n790 VSS 0.00108f
C7003 VDD.n791 VSS 3.16e-19
C7004 VDD.n792 VSS 4.27e-19
C7005 VDD.n793 VSS 1.12e-19
C7006 VDD.n794 VSS 1.85e-19
C7007 VDD.n795 VSS 1.12e-19
C7008 VDD.n796 VSS 9.14e-19
C7009 VDD.n797 VSS 6.55e-20
C7010 VDD.t199 VSS 0.00313f
C7011 VDD.n798 VSS 3.28e-19
C7012 VDD.n799 VSS 1.12e-19
C7013 VDD.n800 VSS 9.03e-19
C7014 VDD.n801 VSS 4.27e-19
C7015 VDD.n802 VSS 3.16e-19
C7016 VDD.n803 VSS 7.09e-19
C7017 VDD.n804 VSS 7.51e-20
C7018 VDD.n805 VSS 1.58e-19
C7019 VDD.n806 VSS 9.14e-19
C7020 VDD.n807 VSS 3.28e-19
C7021 VDD.n808 VSS 0.00317f
C7022 VDD.n809 VSS 3.16e-19
C7023 VDD.n810 VSS 4.27e-19
C7024 VDD.n811 VSS 1.12e-19
C7025 VDD.n812 VSS 1.85e-19
C7026 VDD.n813 VSS 1.12e-19
C7027 VDD.n814 VSS 9.14e-19
C7028 VDD.n815 VSS 6.55e-20
C7029 VDD.t557 VSS 0.00313f
C7030 VDD.n816 VSS 3.28e-19
C7031 VDD.n817 VSS 1.12e-19
C7032 VDD.n818 VSS 9.03e-19
C7033 VDD.n819 VSS 1.05e-19
C7034 VDD.n820 VSS 7.5e-20
C7035 VDD.n821 VSS 3.28e-19
C7036 VDD.n822 VSS 8.76e-19
C7037 VDD.n823 VSS 3.16e-19
C7038 VDD.n824 VSS 4.27e-19
C7039 VDD.n825 VSS 1.12e-19
C7040 VDD.n826 VSS 1.85e-19
C7041 VDD.n827 VSS 1.12e-19
C7042 VDD.n828 VSS 9.14e-19
C7043 VDD.n829 VSS 6.55e-20
C7044 VDD.t200 VSS 0.00313f
C7045 VDD.n830 VSS 3.28e-19
C7046 VDD.n831 VSS 1.12e-19
C7047 VDD.n832 VSS 9.03e-19
C7048 VDD.n833 VSS 4.27e-19
C7049 VDD.n834 VSS 3.16e-19
C7050 VDD.n835 VSS 7.09e-19
C7051 VDD.n836 VSS 6.55e-20
C7052 VDD.n837 VSS 1.12e-19
C7053 VDD.n838 VSS 4.34e-19
C7054 VDD.n839 VSS 1.12e-19
C7055 VDD.n840 VSS 1.85e-19
C7056 VDD.n841 VSS 1.12e-19
C7057 VDD.n842 VSS 3.28e-19
C7058 VDD.n843 VSS 0.00342f
C7059 VDD.n844 VSS 3.16e-19
C7060 VDD.n845 VSS 1.31e-19
C7061 VDD.n846 VSS 1.85e-19
C7062 VDD.n847 VSS 4.54e-19
C7063 VDD.n849 VSS 0.002f
C7064 VDD.n850 VSS 0.00102f
C7065 VDD.n851 VSS 7.09e-19
C7066 VDD.n852 VSS 2.81e-19
C7067 VDD.n853 VSS 0.00517f
C7068 VDD.n854 VSS 7.09e-19
C7069 VDD.n855 VSS 0.00272f
C7070 VDD.t560 VSS 0.0017f
C7071 VDD.n856 VSS 0.00171f
C7072 VDD.n857 VSS 0.002f
C7073 VDD.n858 VSS 0.00116f
C7074 VDD.n859 VSS 7.09e-19
C7075 VDD.t344 VSS 0.00384f
C7076 VDD.n860 VSS 7.18e-19
C7077 VDD.n861 VSS 0.0013f
C7078 VDD.n862 VSS 9.79e-19
C7079 VDD.n863 VSS 7.09e-19
C7080 VDD.t634 VSS 0.00384f
C7081 VDD.n864 VSS 7.09e-19
C7082 VDD.n865 VSS 7.76e-19
C7083 VDD.n866 VSS 0.002f
C7084 VDD.t451 VSS 9.19e-19
C7085 VDD.n867 VSS 9.79e-19
C7086 VDD.n868 VSS 7.09e-19
C7087 VDD.t636 VSS 0.00384f
C7088 VDD.n869 VSS 7.09e-19
C7089 VDD.n870 VSS 0.00116f
C7090 VDD.n871 VSS 0.002f
C7091 VDD.t82 VSS 3.71e-19
C7092 VDD.t532 VSS 3.52e-19
C7093 VDD.n872 VSS 7.74e-19
C7094 VDD.n873 VSS 7.62e-19
C7095 VDD.n874 VSS 7.09e-19
C7096 VDD.t314 VSS 0.00363f
C7097 VDD.n875 VSS 7.09e-19
C7098 VDD.n876 VSS 6.7e-19
C7099 VDD.n877 VSS 0.002f
C7100 VDD.n878 VSS 0.00121f
C7101 VDD.n879 VSS 7.09e-19
C7102 VDD.t17 VSS 0.00384f
C7103 VDD.n880 VSS 7.09e-19
C7104 VDD.n881 VSS 0.00121f
C7105 VDD.n882 VSS 0.002f
C7106 VDD.t80 VSS 3.71e-19
C7107 VDD.t137 VSS 3.71e-19
C7108 VDD.n883 VSS 7.84e-19
C7109 VDD.n884 VSS 0.00164f
C7110 VDD.n885 VSS 0.00133f
C7111 VDD.n886 VSS 7.19e-19
C7112 VDD.t182 VSS 0.00384f
C7113 VDD.n887 VSS 7.09e-19
C7114 VDD.n888 VSS 0.00102f
C7115 VDD.n889 VSS 0.002f
C7116 VDD.n890 VSS 0.00272f
C7117 VDD.n891 VSS 7.09e-19
C7118 VDD.t134 VSS 0.00384f
C7119 VDD.n892 VSS 7.09e-19
C7120 VDD.n893 VSS 0.00116f
C7121 VDD.t135 VSS -3.29e-19
C7122 VDD.t455 VSS 5.95e-19
C7123 VDD.n894 VSS 0.00233f
C7124 VDD.n895 VSS 0.00159f
C7125 VDD.n896 VSS 0.002f
C7126 VDD.t670 VSS -1.76e-19
C7127 VDD.t133 VSS 5.51e-19
C7128 VDD.n897 VSS 0.00259f
C7129 VDD.n898 VSS 0.00235f
C7130 VDD.n899 VSS 0.0013f
C7131 VDD.n900 VSS 7.18e-19
C7132 VDD.n901 VSS 7.09e-19
C7133 VDD.n902 VSS 9.79e-19
C7134 VDD.n903 VSS 0.002f
C7135 VDD.t270 VSS 3.92e-19
C7136 VDD.t333 VSS 3.92e-19
C7137 VDD.n904 VSS 8.47e-19
C7138 VDD.n905 VSS 7.76e-19
C7139 VDD.n906 VSS 7.09e-19
C7140 VDD.t115 VSS 0.00384f
C7141 VDD.n907 VSS 7.09e-19
C7142 VDD.n908 VSS 9.79e-19
C7143 VDD.n909 VSS 0.002f
C7144 VDD.n910 VSS 0.00116f
C7145 VDD.n911 VSS 7.09e-19
C7146 VDD.t604 VSS 0.00384f
C7147 VDD.n912 VSS 7.09e-19
C7148 VDD.n913 VSS 7.62e-19
C7149 VDD.n914 VSS 0.002f
C7150 VDD.n915 VSS 6.7e-19
C7151 VDD.n916 VSS 7.09e-19
C7152 VDD.t549 VSS 0.00384f
C7153 VDD.n917 VSS 7.09e-19
C7154 VDD.n918 VSS 0.00121f
C7155 VDD.t550 VSS 0.00141f
C7156 VDD.t564 VSS 6.28e-19
C7157 VDD.n919 VSS 0.00226f
C7158 VDD.n920 VSS 0.00297f
C7159 VDD.n921 VSS 0.002f
C7160 VDD.n922 VSS 0.00121f
C7161 VDD.n923 VSS 7.09e-19
C7162 VDD.t42 VSS 0.00384f
C7163 VDD.n924 VSS 7.19e-19
C7164 VDD.n925 VSS 0.00133f
C7165 VDD.n926 VSS 0.002f
C7166 VDD.n927 VSS 0.00102f
C7167 VDD.n928 VSS 7.09e-19
C7168 VDD.n929 VSS 0.00517f
C7169 VDD.n930 VSS 7.09e-19
C7170 VDD.n931 VSS 0.00272f
C7171 VDD.t562 VSS 0.0017f
C7172 VDD.n932 VSS 0.00171f
C7173 VDD.n933 VSS 0.002f
C7174 VDD.n934 VSS 0.00116f
C7175 VDD.n935 VSS 7.09e-19
C7176 VDD.t44 VSS 0.00384f
C7177 VDD.n936 VSS 7.18e-19
C7178 VDD.n937 VSS 0.0013f
C7179 VDD.n938 VSS 9.79e-19
C7180 VDD.n939 VSS 7.09e-19
C7181 VDD.t336 VSS 0.00384f
C7182 VDD.n940 VSS 7.09e-19
C7183 VDD.n941 VSS 7.76e-19
C7184 VDD.n942 VSS 0.002f
C7185 VDD.t184 VSS 9.19e-19
C7186 VDD.n943 VSS 9.79e-19
C7187 VDD.n944 VSS 7.09e-19
C7188 VDD.t334 VSS 0.00384f
C7189 VDD.n945 VSS 7.09e-19
C7190 VDD.n946 VSS 0.00116f
C7191 VDD.n947 VSS 0.002f
C7192 VDD.t343 VSS 3.71e-19
C7193 VDD.t186 VSS 3.52e-19
C7194 VDD.n948 VSS 7.74e-19
C7195 VDD.n949 VSS 7.62e-19
C7196 VDD.n950 VSS 7.09e-19
C7197 VDD.t83 VSS 0.00363f
C7198 VDD.n951 VSS 7.09e-19
C7199 VDD.n952 VSS 6.7e-19
C7200 VDD.n953 VSS 0.002f
C7201 VDD.n954 VSS 0.00121f
C7202 VDD.n955 VSS 7.09e-19
C7203 VDD.t38 VSS 0.00384f
C7204 VDD.n956 VSS 7.09e-19
C7205 VDD.n957 VSS 0.00121f
C7206 VDD.n958 VSS 0.002f
C7207 VDD.t341 VSS 3.71e-19
C7208 VDD.t613 VSS 3.71e-19
C7209 VDD.n959 VSS 7.84e-19
C7210 VDD.n960 VSS 0.00164f
C7211 VDD.n961 VSS 0.00133f
C7212 VDD.n962 VSS 7.19e-19
C7213 VDD.t577 VSS 0.00384f
C7214 VDD.n963 VSS 7.09e-19
C7215 VDD.n964 VSS 0.00102f
C7216 VDD.n965 VSS 0.002f
C7217 VDD.n966 VSS 0.00272f
C7218 VDD.n967 VSS 7.09e-19
C7219 VDD.t614 VSS 0.00384f
C7220 VDD.n968 VSS 7.09e-19
C7221 VDD.n969 VSS 0.00116f
C7222 VDD.t615 VSS -3.29e-19
C7223 VDD.t35 VSS 5.95e-19
C7224 VDD.n970 VSS 0.00233f
C7225 VDD.n971 VSS 0.00159f
C7226 VDD.n972 VSS 0.00628f
C7227 VDD.t611 VSS -1.76e-19
C7228 VDD.t617 VSS 5.51e-19
C7229 VDD.n973 VSS 0.00259f
C7230 VDD.n974 VSS 0.00235f
C7231 VDD.n975 VSS 0.0013f
C7232 VDD.n976 VSS 7.18e-19
C7233 VDD.n977 VSS 0.00114f
C7234 VDD.n978 VSS 0.00891f
C7235 VDD.t610 VSS 0.0044f
C7236 VDD.n979 VSS 0.00396f
C7237 VDD.t616 VSS 0.00384f
C7238 VDD.n980 VSS 0.00613f
C7239 VDD.n981 VSS 0.00555f
C7240 VDD.n982 VSS 7.09e-19
C7241 VDD.n983 VSS 0.00105f
C7242 VDD.n984 VSS 0.002f
C7243 VDD.n985 VSS 0.002f
C7244 VDD.n986 VSS 0.002f
C7245 VDD.n987 VSS 0.00121f
C7246 VDD.n988 VSS 7.09e-19
C7247 VDD.n989 VSS 0.00405f
C7248 VDD.t34 VSS 0.00384f
C7249 VDD.n990 VSS 0.00517f
C7250 VDD.n991 VSS 0.003f
C7251 VDD.t667 VSS 0.00384f
C7252 VDD.n992 VSS 0.00692f
C7253 VDD.n993 VSS 7.09e-19
C7254 VDD.t668 VSS 0.0017f
C7255 VDD.n994 VSS 0.00171f
C7256 VDD.n995 VSS 0.00188f
C7257 VDD.n996 VSS 0.002f
C7258 VDD.n997 VSS 0.002f
C7259 VDD.n998 VSS 0.002f
C7260 VDD.n999 VSS 0.00106f
C7261 VDD.n1000 VSS 7.09e-19
C7262 VDD.n1001 VSS 0.004f
C7263 VDD.t340 VSS 0.00384f
C7264 VDD.n1002 VSS 0.0045f
C7265 VDD.t612 VSS 0.00384f
C7266 VDD.n1003 VSS 0.00417f
C7267 VDD.n1004 VSS 0.00459f
C7268 VDD.n1005 VSS 7.09e-19
C7269 VDD.n1006 VSS 8.61e-19
C7270 VDD.n1007 VSS 0.002f
C7271 VDD.n1008 VSS 0.002f
C7272 VDD.n1009 VSS 0.002f
C7273 VDD.n1010 VSS 0.00121f
C7274 VDD.n1011 VSS 7.09e-19
C7275 VDD.t335 VSS 0.00734f
C7276 VDD.n1012 VSS 0.00601f
C7277 VDD.t187 VSS 0.00384f
C7278 VDD.t665 VSS 0.00371f
C7279 VDD.n1013 VSS 0.00405f
C7280 VDD.n1014 VSS 0.00551f
C7281 VDD.n1015 VSS 7.09e-19
C7282 VDD.t188 VSS 0.00141f
C7283 VDD.t666 VSS 6.28e-19
C7284 VDD.n1016 VSS 0.00226f
C7285 VDD.n1017 VSS 0.00297f
C7286 VDD.n1018 VSS 7.1e-19
C7287 VDD.n1019 VSS 0.002f
C7288 VDD.n1020 VSS 0.002f
C7289 VDD.n1021 VSS 0.002f
C7290 VDD.n1022 VSS 0.00121f
C7291 VDD.n1023 VSS 7.09e-19
C7292 VDD.n1024 VSS 0.00396f
C7293 VDD.n1025 VSS 0.00438f
C7294 VDD.t342 VSS 0.00384f
C7295 VDD.n1026 VSS 0.005f
C7296 VDD.t185 VSS 0.00384f
C7297 VDD.n1027 VSS 0.00442f
C7298 VDD.n1028 VSS 7.19e-19
C7299 VDD.n1029 VSS 0.00133f
C7300 VDD.n1030 VSS 0.0018f
C7301 VDD.n1031 VSS 0.002f
C7302 VDD.n1032 VSS 0.002f
C7303 VDD.n1033 VSS 0.002f
C7304 VDD.n1034 VSS 0.00121f
C7305 VDD.n1035 VSS 7.09e-19
C7306 VDD.n1036 VSS 0.0035f
C7307 VDD.t39 VSS 0.00384f
C7308 VDD.n1037 VSS 0.00388f
C7309 VDD.t183 VSS 0.00384f
C7310 VDD.n1038 VSS 0.00601f
C7311 VDD.n1039 VSS 0.00567f
C7312 VDD.n1040 VSS 7.19e-19
C7313 VDD.n1041 VSS 0.00132f
C7314 VDD.n1042 VSS 0.002f
C7315 VDD.n1043 VSS 0.002f
C7316 VDD.n1044 VSS 0.002f
C7317 VDD.n1045 VSS 0.00118f
C7318 VDD.n1046 VSS 0.002f
C7319 VDD.t337 VSS 3.92e-19
C7320 VDD.t339 VSS 3.92e-19
C7321 VDD.n1047 VSS 8.47e-19
C7322 VDD.n1048 VSS 0.00176f
C7323 VDD.n1049 VSS 0.00131f
C7324 VDD.n1050 VSS 7.19e-19
C7325 VDD.n1051 VSS 0.0035f
C7326 VDD.t338 VSS 0.0038f
C7327 VDD.n1052 VSS 7.09e-19
C7328 VDD.n1053 VSS 0.00396f
C7329 VDD.t458 VSS 0.00384f
C7330 VDD.n1054 VSS 0.00517f
C7331 VDD.n1055 VSS 7.09e-19
C7332 VDD.n1056 VSS 9.79e-19
C7333 VDD.n1057 VSS 0.0015f
C7334 VDD.t459 VSS -1.76e-19
C7335 VDD.t45 VSS 5.51e-19
C7336 VDD.n1058 VSS 0.00259f
C7337 VDD.n1059 VSS 0.00235f
C7338 VDD.n1060 VSS 0.002f
C7339 VDD.n1061 VSS 0.002f
C7340 VDD.n1062 VSS 0.00105f
C7341 VDD.n1063 VSS 7.09e-19
C7342 VDD.n1064 VSS 0.00555f
C7343 VDD.n1065 VSS 0.00613f
C7344 VDD.t46 VSS 0.00384f
C7345 VDD.t472 VSS 0.00384f
C7346 VDD.n1066 VSS 0.00405f
C7347 VDD.n1067 VSS 7.09e-19
C7348 VDD.t47 VSS -3.29e-19
C7349 VDD.t473 VSS 5.95e-19
C7350 VDD.n1068 VSS 0.00233f
C7351 VDD.n1069 VSS 0.00159f
C7352 VDD.n1070 VSS 0.00121f
C7353 VDD.n1071 VSS 0.002f
C7354 VDD.n1072 VSS 0.002f
C7355 VDD.n1073 VSS 0.002f
C7356 VDD.n1074 VSS 0.00188f
C7357 VDD.n1075 VSS 7.09e-19
C7358 VDD.n1076 VSS 0.00692f
C7359 VDD.t561 VSS 0.00384f
C7360 VDD.n1077 VSS 0.003f
C7361 VDD.t84 VSS 0.00384f
C7362 VDD.n1078 VSS 0.0045f
C7363 VDD.t602 VSS 0.00384f
C7364 VDD.n1079 VSS 0.004f
C7365 VDD.n1080 VSS 7.09e-19
C7366 VDD.n1081 VSS 0.00106f
C7367 VDD.n1082 VSS 0.002f
C7368 VDD.t603 VSS 3.71e-19
C7369 VDD.t43 VSS 3.71e-19
C7370 VDD.n1083 VSS 7.84e-19
C7371 VDD.n1084 VSS 0.00164f
C7372 VDD.n1085 VSS 0.002f
C7373 VDD.n1086 VSS 0.002f
C7374 VDD.n1087 VSS 8.61e-19
C7375 VDD.n1088 VSS 7.09e-19
C7376 VDD.n1089 VSS 0.00459f
C7377 VDD.n1090 VSS 0.00417f
C7378 VDD.t51 VSS 0.00384f
C7379 VDD.n1091 VSS 0.00601f
C7380 VDD.t268 VSS 0.00734f
C7381 VDD.n1092 VSS 7.09e-19
C7382 VDD.n1093 VSS 0.00121f
C7383 VDD.n1094 VSS 0.002f
C7384 VDD.n1095 VSS 0.002f
C7385 VDD.n1096 VSS 0.002f
C7386 VDD.n1097 VSS 7.1e-19
C7387 VDD.n1098 VSS 7.09e-19
C7388 VDD.n1099 VSS 0.00551f
C7389 VDD.n1100 VSS 0.00405f
C7390 VDD.t563 VSS 0.00371f
C7391 VDD.t533 VSS 0.00363f
C7392 VDD.n1101 VSS 0.00438f
C7393 VDD.n1102 VSS 0.00396f
C7394 VDD.n1103 VSS 7.09e-19
C7395 VDD.n1104 VSS 0.00121f
C7396 VDD.n1105 VSS 0.002f
C7397 VDD.n1106 VSS 0.002f
C7398 VDD.n1107 VSS 0.002f
C7399 VDD.t605 VSS 3.71e-19
C7400 VDD.t548 VSS 3.52e-19
C7401 VDD.n1108 VSS 7.74e-19
C7402 VDD.n1109 VSS 0.0018f
C7403 VDD.n1110 VSS 0.00133f
C7404 VDD.n1111 VSS 7.19e-19
C7405 VDD.n1112 VSS 0.00442f
C7406 VDD.t547 VSS 0.00384f
C7407 VDD.n1113 VSS 0.005f
C7408 VDD.t267 VSS 0.00384f
C7409 VDD.n1114 VSS 0.00388f
C7410 VDD.t50 VSS 0.00384f
C7411 VDD.n1115 VSS 0.0035f
C7412 VDD.n1116 VSS 7.09e-19
C7413 VDD.n1117 VSS 0.00121f
C7414 VDD.n1118 VSS 0.002f
C7415 VDD.n1119 VSS 0.002f
C7416 VDD.n1120 VSS 0.002f
C7417 VDD.t116 VSS 9.19e-19
C7418 VDD.n1121 VSS 0.002f
C7419 VDD.n1122 VSS 0.00132f
C7420 VDD.n1123 VSS 7.19e-19
C7421 VDD.n1124 VSS 0.00567f
C7422 VDD.n1125 VSS 0.00601f
C7423 VDD.t269 VSS 0.00384f
C7424 VDD.n1126 VSS 7.09e-19
C7425 VDD.t332 VSS 0.0038f
C7426 VDD.n1127 VSS 0.0035f
C7427 VDD.n1128 VSS 7.19e-19
C7428 VDD.n1129 VSS 0.00131f
C7429 VDD.n1130 VSS 0.00176f
C7430 VDD.n1131 VSS 0.002f
C7431 VDD.n1132 VSS 0.00118f
C7432 VDD.n1133 VSS 0.0015f
C7433 VDD.n1134 VSS 9.79e-19
C7434 VDD.n1135 VSS 7.09e-19
C7435 VDD.n1136 VSS 0.00517f
C7436 VDD.t669 VSS 0.00384f
C7437 VDD.n1137 VSS 0.00396f
C7438 VDD.t132 VSS 0.00384f
C7439 VDD.n1138 VSS 0.00613f
C7440 VDD.n1139 VSS 0.00555f
C7441 VDD.n1140 VSS 7.09e-19
C7442 VDD.n1141 VSS 0.00105f
C7443 VDD.n1142 VSS 0.002f
C7444 VDD.n1143 VSS 0.002f
C7445 VDD.n1144 VSS 0.002f
C7446 VDD.n1145 VSS 0.00121f
C7447 VDD.n1146 VSS 7.09e-19
C7448 VDD.n1147 VSS 0.00405f
C7449 VDD.t454 VSS 0.00384f
C7450 VDD.n1148 VSS 0.00517f
C7451 VDD.n1149 VSS 0.003f
C7452 VDD.t287 VSS 0.00384f
C7453 VDD.n1150 VSS 0.00692f
C7454 VDD.n1151 VSS 7.09e-19
C7455 VDD.t288 VSS 0.0017f
C7456 VDD.n1152 VSS 0.00171f
C7457 VDD.n1153 VSS 0.00188f
C7458 VDD.n1154 VSS 0.002f
C7459 VDD.n1155 VSS 0.002f
C7460 VDD.n1156 VSS 0.002f
C7461 VDD.n1157 VSS 0.00106f
C7462 VDD.n1158 VSS 7.09e-19
C7463 VDD.n1159 VSS 0.004f
C7464 VDD.t79 VSS 0.00384f
C7465 VDD.n1160 VSS 0.0045f
C7466 VDD.t136 VSS 0.00384f
C7467 VDD.n1161 VSS 0.00417f
C7468 VDD.n1162 VSS 0.00459f
C7469 VDD.n1163 VSS 7.09e-19
C7470 VDD.n1164 VSS 8.61e-19
C7471 VDD.n1165 VSS 0.002f
C7472 VDD.n1166 VSS 0.002f
C7473 VDD.n1167 VSS 0.002f
C7474 VDD.n1168 VSS 0.00121f
C7475 VDD.n1169 VSS 7.09e-19
C7476 VDD.t637 VSS 0.00734f
C7477 VDD.n1170 VSS 0.00601f
C7478 VDD.t529 VSS 0.00384f
C7479 VDD.t285 VSS 0.00371f
C7480 VDD.n1171 VSS 0.00405f
C7481 VDD.n1172 VSS 0.00551f
C7482 VDD.n1173 VSS 7.09e-19
C7483 VDD.t530 VSS 0.00141f
C7484 VDD.t286 VSS 6.28e-19
C7485 VDD.n1174 VSS 0.00226f
C7486 VDD.n1175 VSS 0.00297f
C7487 VDD.n1176 VSS 7.1e-19
C7488 VDD.n1177 VSS 0.002f
C7489 VDD.n1178 VSS 0.002f
C7490 VDD.n1179 VSS 0.002f
C7491 VDD.n1180 VSS 0.00121f
C7492 VDD.n1181 VSS 7.09e-19
C7493 VDD.n1182 VSS 0.00396f
C7494 VDD.n1183 VSS 0.00438f
C7495 VDD.t81 VSS 0.00384f
C7496 VDD.n1184 VSS 0.005f
C7497 VDD.t531 VSS 0.00384f
C7498 VDD.n1185 VSS 0.00442f
C7499 VDD.n1186 VSS 7.19e-19
C7500 VDD.n1187 VSS 0.00133f
C7501 VDD.n1188 VSS 0.0018f
C7502 VDD.n1189 VSS 0.002f
C7503 VDD.n1190 VSS 0.002f
C7504 VDD.n1191 VSS 0.002f
C7505 VDD.n1192 VSS 0.00121f
C7506 VDD.n1193 VSS 7.09e-19
C7507 VDD.n1194 VSS 0.0035f
C7508 VDD.t16 VSS 0.00384f
C7509 VDD.n1195 VSS 0.00388f
C7510 VDD.t450 VSS 0.00384f
C7511 VDD.n1196 VSS 0.00601f
C7512 VDD.n1197 VSS 0.00567f
C7513 VDD.n1198 VSS 7.19e-19
C7514 VDD.n1199 VSS 0.00132f
C7515 VDD.n1200 VSS 0.002f
C7516 VDD.n1201 VSS 0.002f
C7517 VDD.n1202 VSS 0.002f
C7518 VDD.n1203 VSS 0.00118f
C7519 VDD.n1204 VSS 0.002f
C7520 VDD.t635 VSS 3.92e-19
C7521 VDD.t170 VSS 3.92e-19
C7522 VDD.n1205 VSS 8.47e-19
C7523 VDD.n1206 VSS 0.00176f
C7524 VDD.n1207 VSS 0.00131f
C7525 VDD.n1208 VSS 7.19e-19
C7526 VDD.n1209 VSS 0.0035f
C7527 VDD.t169 VSS 0.0038f
C7528 VDD.n1210 VSS 7.09e-19
C7529 VDD.n1211 VSS 0.00396f
C7530 VDD.t122 VSS 0.00384f
C7531 VDD.n1212 VSS 0.00517f
C7532 VDD.n1213 VSS 7.09e-19
C7533 VDD.n1214 VSS 9.79e-19
C7534 VDD.n1215 VSS 0.0015f
C7535 VDD.t123 VSS -1.76e-19
C7536 VDD.t345 VSS 5.51e-19
C7537 VDD.n1216 VSS 0.00259f
C7538 VDD.n1217 VSS 0.00235f
C7539 VDD.n1218 VSS 0.002f
C7540 VDD.n1219 VSS 0.002f
C7541 VDD.n1220 VSS 0.00105f
C7542 VDD.n1221 VSS 7.09e-19
C7543 VDD.n1222 VSS 0.00555f
C7544 VDD.n1223 VSS 0.00613f
C7545 VDD.t346 VSS 0.00384f
C7546 VDD.t526 VSS 0.00384f
C7547 VDD.n1224 VSS 0.00405f
C7548 VDD.n1225 VSS 7.09e-19
C7549 VDD.t347 VSS -3.29e-19
C7550 VDD.t527 VSS 5.95e-19
C7551 VDD.n1226 VSS 0.00233f
C7552 VDD.n1227 VSS 0.00159f
C7553 VDD.n1228 VSS 0.00121f
C7554 VDD.n1229 VSS 0.002f
C7555 VDD.n1230 VSS 0.002f
C7556 VDD.n1231 VSS 0.002f
C7557 VDD.n1232 VSS 0.00188f
C7558 VDD.n1233 VSS 7.09e-19
C7559 VDD.n1234 VSS 0.00692f
C7560 VDD.t559 VSS 0.00384f
C7561 VDD.n1235 VSS 0.003f
C7562 VDD.t178 VSS 0.00384f
C7563 VDD.n1236 VSS 3.28e-19
C7564 VDD.n1237 VSS 0.00354f
C7565 VDD.n1238 VSS 7.51e-20
C7566 VDD.n1239 VSS 7.09e-19
C7567 VDD.n1240 VSS 6.26e-19
C7568 VDD.t6 VSS 0.00275f
C7569 VDD.n1241 VSS 0.004f
C7570 VDD.n1242 VSS 6.09e-19
C7571 VDD.n1243 VSS 0.00104f
C7572 VDD.n1244 VSS 0.0019f
C7573 VDD.n1245 VSS 0.001f
C7574 VDD.t7 VSS 3.71e-19
C7575 VDD.t349 VSS 3.71e-19
C7576 VDD.n1246 VSS 7.8e-19
C7577 VDD.n1247 VSS 0.00164f
C7578 VDD.n1248 VSS 7.23e-19
C7579 VDD.n1249 VSS 9.03e-19
C7580 VDD.n1250 VSS 9.14e-19
C7581 VDD.n1251 VSS 1.25e-19
C7582 VDD.n1252 VSS 1.12e-19
C7583 VDD.n1253 VSS 6.55e-20
C7584 VDD.n1254 VSS 3.34e-19
C7585 VDD.t348 VSS 4.17e-19
C7586 VDD.n1255 VSS 0.0035f
C7587 VDD.n1256 VSS 0.00342f
C7588 VDD.n1257 VSS 3.16e-19
C7589 VDD.n1258 VSS 4.27e-19
C7590 VDD.n1259 VSS 4.34e-19
C7591 VDD.n1260 VSS 9.03e-19
C7592 VDD.n1261 VSS 1.85e-19
C7593 VDD.n1262 VSS 9.14e-19
C7594 VDD.n1263 VSS 1.25e-19
C7595 VDD.n1264 VSS 3.28e-19
C7596 VDD.n1265 VSS 0.00113f
C7597 VDD.t109 VSS 0.00313f
C7598 VDD.n1266 VSS 0.00271f
C7599 VDD.n1267 VSS 7.92e-19
C7600 VDD.n1268 VSS 7.09e-19
C7601 VDD.n1269 VSS 6.55e-20
C7602 VDD.n1270 VSS 1.12e-19
C7603 VDD.n1271 VSS 1.25e-19
C7604 VDD.n1272 VSS 9.14e-19
C7605 VDD.n1273 VSS 1.85e-19
C7606 VDD.n1274 VSS 9.03e-19
C7607 VDD.n1275 VSS 4.34e-19
C7608 VDD.n1276 VSS 4.27e-19
C7609 VDD.n1277 VSS 3.16e-19
C7610 VDD.n1278 VSS 0.00304f
C7611 VDD.n1279 VSS 7.09e-19
C7612 VDD.t689 VSS 0.00313f
C7613 VDD.n1280 VSS 0.00296f
C7614 VDD.n1281 VSS 3.28e-19
C7615 VDD.n1282 VSS 1.25e-19
C7616 VDD.n1283 VSS 1.12e-19
C7617 VDD.n1284 VSS 4.34e-19
C7618 VDD.n1285 VSS 9.03e-19
C7619 VDD.n1286 VSS 1.85e-19
C7620 VDD.n1287 VSS 9.14e-19
C7621 VDD.n1288 VSS 1.25e-19
C7622 VDD.n1289 VSS 1.12e-19
C7623 VDD.n1290 VSS 6.55e-20
C7624 VDD.n1291 VSS 7.09e-19
C7625 VDD.n1292 VSS 0.00354f
C7626 VDD.n1293 VSS 0.001f
C7627 VDD.n1294 VSS 7.09e-19
C7628 VDD.n1295 VSS 0.00342f
C7629 VDD.n1296 VSS 3.16e-19
C7630 VDD.t690 VSS 0.00141f
C7631 VDD.t558 VSS 6.28e-19
C7632 VDD.n1298 VSS 0.00226f
C7633 VDD.n1299 VSS 0.00284f
C7634 VDD.n1300 VSS 6.57e-20
C7635 VDD.n1301 VSS 9.14e-19
C7636 VDD.n1302 VSS 1.85e-19
C7637 VDD.n1303 VSS 9.03e-19
C7638 VDD.n1304 VSS 4.34e-19
C7639 VDD.n1305 VSS 4.27e-19
C7640 VDD.n1306 VSS 3.16e-19
C7641 VDD.n1307 VSS 0.00284f
C7642 VDD.n1308 VSS 7.09e-19
C7643 VDD.t114 VSS 0.00313f
C7644 VDD.n1309 VSS 6.67e-19
C7645 VDD.n1310 VSS 3.28e-19
C7646 VDD.n1311 VSS 1.25e-19
C7647 VDD.n1312 VSS 1.12e-19
C7648 VDD.n1313 VSS 4.34e-19
C7649 VDD.n1314 VSS 9.03e-19
C7650 VDD.n1315 VSS 9.03e-19
C7651 VDD.n1316 VSS 1.85e-19
C7652 VDD.n1317 VSS 9.14e-19
C7653 VDD.n1318 VSS 1.25e-19
C7654 VDD.n1319 VSS 1.12e-19
C7655 VDD.n1320 VSS 6.55e-20
C7656 VDD.n1321 VSS 7.09e-19
C7657 VDD.n1322 VSS 0.00133f
C7658 VDD.t4 VSS 0.00313f
C7659 VDD.n1323 VSS 0.0025f
C7660 VDD.n1324 VSS 3.16e-19
C7661 VDD.t5 VSS 3.71e-19
C7662 VDD.t688 VSS 3.52e-19
C7663 VDD.n1325 VSS 7.7e-19
C7664 VDD.n1326 VSS 1.85e-19
C7665 VDD.n1327 VSS 0.00181f
C7666 VDD.n1328 VSS 0.0011f
C7667 VDD.n1330 VSS 3.28e-19
C7668 VDD.n1331 VSS 0.00192f
C7669 VDD.t687 VSS 0.00313f
C7670 VDD.n1332 VSS 0.00192f
C7671 VDD.n1333 VSS 0.00309f
C7672 VDD.n1334 VSS 7.09e-19
C7673 VDD.n1335 VSS 6.55e-20
C7674 VDD.n1336 VSS 1.12e-19
C7675 VDD.n1337 VSS 1.25e-19
C7676 VDD.n1338 VSS 9.14e-19
C7677 VDD.n1339 VSS 1.85e-19
C7678 VDD.n1340 VSS 9.03e-19
C7679 VDD.n1341 VSS 4.34e-19
C7680 VDD.n1342 VSS 4.27e-19
C7681 VDD.n1343 VSS 3.16e-19
C7682 VDD.n1344 VSS 7.51e-19
C7683 VDD.n1345 VSS 7.09e-19
C7684 VDD.t108 VSS 0.00313f
C7685 VDD.n1346 VSS 0.00275f
C7686 VDD.n1347 VSS 3.28e-19
C7687 VDD.n1348 VSS 1.25e-19
C7688 VDD.n1349 VSS 1.12e-19
C7689 VDD.n1350 VSS 4.34e-19
C7690 VDD.n1351 VSS 9.03e-19
C7691 VDD.n1352 VSS 9.03e-19
C7692 VDD.n1353 VSS 1.85e-19
C7693 VDD.n1354 VSS 9.14e-19
C7694 VDD.n1355 VSS 1.25e-19
C7695 VDD.n1356 VSS 1.12e-19
C7696 VDD.n1357 VSS 6.55e-20
C7697 VDD.n1358 VSS 7.09e-19
C7698 VDD.n1359 VSS 0.00279f
C7699 VDD.t283 VSS 0.00313f
C7700 VDD.n1360 VSS 3.28e-19
C7701 VDD.n1361 VSS 0.00354f
C7702 VDD.n1362 VSS 7.09e-19
C7703 VDD.n1363 VSS 0.00104f
C7704 VDD.n1364 VSS 3.16e-19
C7705 VDD.t284 VSS 9.16e-19
C7706 VDD.n1365 VSS 0.002f
C7707 VDD.n1366 VSS 0.00109f
C7708 VDD.n1367 VSS 9.03e-19
C7709 VDD.n1368 VSS 9.03e-19
C7710 VDD.n1369 VSS 1.85e-19
C7711 VDD.n1370 VSS 9.14e-19
C7712 VDD.n1371 VSS 1.25e-19
C7713 VDD.n1372 VSS 1.12e-19
C7714 VDD.n1373 VSS 6.55e-20
C7715 VDD.n1374 VSS 7.09e-19
C7716 VDD.n1375 VSS 0.00296f
C7717 VDD.t197 VSS 0.00313f
C7718 VDD.n1376 VSS 8.76e-19
C7719 VDD.n1377 VSS 3.16e-19
C7720 VDD.t198 VSS 3.92e-19
C7721 VDD.t152 VSS 3.92e-19
C7722 VDD.n1378 VSS 8.43e-19
C7723 VDD.n1379 VSS 1.85e-19
C7724 VDD.n1380 VSS 0.00176f
C7725 VDD.n1381 VSS 0.00109f
C7726 VDD.n1383 VSS 3.28e-19
C7727 VDD.n1384 VSS 0.00263f
C7728 VDD.t151 VSS 0.00313f
C7729 VDD.n1385 VSS 0.00121f
C7730 VDD.n1386 VSS 7.51e-19
C7731 VDD.n1387 VSS 7.09e-19
C7732 VDD.n1388 VSS 6.55e-20
C7733 VDD.n1389 VSS 1.12e-19
C7734 VDD.n1390 VSS 1.25e-19
C7735 VDD.n1391 VSS 1.12e-19
C7736 VDD.n1392 VSS 1.85e-19
C7737 VDD.n1393 VSS 1.74e-19
C7738 VDD.n1394 VSS 0.00129f
C7739 VDD.n1395 VSS 0.00103f
C7740 VDD.n1396 VSS 6.7e-19
C7741 VDD.n1397 VSS 0.00621f
C7742 VDD.n1398 VSS 0.00396f
C7743 VDD.t195 VSS 0.00384f
C7744 VDD.n1399 VSS 0.00442f
C7745 VDD.n1400 VSS 7.09e-19
C7746 VDD.n1401 VSS 8.87e-19
C7747 VDD.n1402 VSS 0.00119f
C7748 VDD.n1403 VSS 0.002f
C7749 VDD.t327 VSS 5.51e-19
C7750 VDD.t593 VSS -1.76e-19
C7751 VDD.n1404 VSS 0.00259f
C7752 VDD.n1405 VSS 0.00235f
C7753 VDD.n1406 VSS 0.0013f
C7754 VDD.n1407 VSS 7.18e-19
C7755 VDD.n1408 VSS 0.006f
C7756 VDD.n1409 VSS 7.09e-19
C7757 VDD.n1410 VSS 0.00116f
C7758 VDD.n1411 VSS 0.002f
C7759 VDD.t443 VSS 5.95e-19
C7760 VDD.t329 VSS -3.29e-19
C7761 VDD.n1412 VSS 0.00233f
C7762 VDD.n1413 VSS 0.00159f
C7763 VDD.n1414 VSS 7.09e-19
C7764 VDD.t691 VSS 0.00375f
C7765 VDD.n1415 VSS 7.09e-19
C7766 VDD.t692 VSS 0.0017f
C7767 VDD.n1416 VSS 0.00171f
C7768 VDD.n1417 VSS 0.00272f
C7769 VDD.n1418 VSS 0.002f
C7770 VDD.n1419 VSS 0.00133f
C7771 VDD.n1420 VSS 7.19e-19
C7772 VDD.n1421 VSS 0.00408f
C7773 VDD.n1422 VSS 7.09e-19
C7774 VDD.n1423 VSS 0.00121f
C7775 VDD.n1424 VSS 0.002f
C7776 VDD.n1425 VSS 0.00121f
C7777 VDD.n1426 VSS 7.09e-19
C7778 VDD.n1427 VSS 0.00396f
C7779 VDD.n1428 VSS 7.09e-19
C7780 VDD.t694 VSS 6.28e-19
C7781 VDD.t718 VSS 0.00141f
C7782 VDD.n1429 VSS 0.00226f
C7783 VDD.n1430 VSS 0.00297f
C7784 VDD.n1431 VSS 0.002f
C7785 VDD.n1432 VSS 7.62e-19
C7786 VDD.n1433 VSS 7.09e-19
C7787 VDD.t719 VSS 0.00375f
C7788 VDD.n1434 VSS 7.09e-19
C7789 VDD.n1435 VSS 0.00116f
C7790 VDD.n1436 VSS 0.002f
C7791 VDD.n1437 VSS 9.79e-19
C7792 VDD.n1438 VSS 7.09e-19
C7793 VDD.n1439 VSS 0.00588f
C7794 VDD.n1440 VSS 7.09e-19
C7795 VDD.n1441 VSS 7.76e-19
C7796 VDD.t41 VSS 3.92e-19
C7797 VDD.t724 VSS 3.92e-19
C7798 VDD.n1442 VSS 8.47e-19
C7799 VDD.n1443 VSS 9.79e-19
C7800 VDD.n1444 VSS 7.09e-19
C7801 VDD.t125 VSS 0.00375f
C7802 VDD.n1445 VSS 7.18e-19
C7803 VDD.n1446 VSS 0.0013f
C7804 VDD.n1447 VSS 0.002f
C7805 VDD.n1448 VSS 0.00116f
C7806 VDD.n1449 VSS 7.09e-19
C7807 VDD.t440 VSS 0.00375f
C7808 VDD.n1450 VSS 7.09e-19
C7809 VDD.t441 VSS 5.95e-19
C7810 VDD.t708 VSS -3.29e-19
C7811 VDD.n1451 VSS 0.00233f
C7812 VDD.n1452 VSS 0.00159f
C7813 VDD.n1453 VSS 0.002f
C7814 VDD.t641 VSS 0.0017f
C7815 VDD.n1454 VSS 0.00171f
C7816 VDD.n1455 VSS 7.09e-19
C7817 VDD.t545 VSS 0.00375f
C7818 VDD.n1456 VSS 7.19e-19
C7819 VDD.n1457 VSS 0.00133f
C7820 VDD.n1458 VSS 0.00102f
C7821 VDD.n1459 VSS 0.002f
C7822 VDD.n1460 VSS 0.00121f
C7823 VDD.n1461 VSS 7.09e-19
C7824 VDD.n1462 VSS 0.00588f
C7825 VDD.n1463 VSS 7.09e-19
C7826 VDD.n1464 VSS 0.00121f
C7827 VDD.n1465 VSS 0.002f
C7828 VDD.t639 VSS 6.28e-19
C7829 VDD.t11 VSS 0.00141f
C7830 VDD.n1466 VSS 0.00226f
C7831 VDD.n1467 VSS 0.00297f
C7832 VDD.n1468 VSS 7.09e-19
C7833 VDD.n1469 VSS 0.00428f
C7834 VDD.n1470 VSS 7.09e-19
C7835 VDD.n1471 VSS 7.62e-19
C7836 VDD.n1472 VSS 6.7e-19
C7837 VDD.n1473 VSS 0.002f
C7838 VDD.t9 VSS 3.52e-19
C7839 VDD.t544 VSS 3.71e-19
C7840 VDD.n1474 VSS 7.74e-19
C7841 VDD.n1475 VSS 0.00116f
C7842 VDD.n1476 VSS 7.09e-19
C7843 VDD.t103 VSS 0.00375f
C7844 VDD.n1477 VSS 7.09e-19
C7845 VDD.n1478 VSS 9.79e-19
C7846 VDD.n1479 VSS 0.002f
C7847 VDD.t436 VSS 9.19e-19
C7848 VDD.n1480 VSS 7.76e-19
C7849 VDD.n1481 VSS 7.09e-19
C7850 VDD.t675 VSS 0.00302f
C7851 VDD.n1482 VSS 7.09e-19
C7852 VDD.n1483 VSS 9.79e-19
C7853 VDD.n1484 VSS 0.002f
C7854 VDD.t58 VSS 5.51e-19
C7855 VDD.t378 VSS -1.76e-19
C7856 VDD.n1485 VSS 0.00259f
C7857 VDD.n1486 VSS 0.00235f
C7858 VDD.n1487 VSS 0.0013f
C7859 VDD.n1488 VSS 7.18e-19
C7860 VDD.n1489 VSS 0.006f
C7861 VDD.n1490 VSS 7.09e-19
C7862 VDD.n1491 VSS 0.00116f
C7863 VDD.n1492 VSS 0.002f
C7864 VDD.t627 VSS 5.95e-19
C7865 VDD.t56 VSS -3.29e-19
C7866 VDD.n1493 VSS 0.00233f
C7867 VDD.n1494 VSS 0.00159f
C7868 VDD.n1495 VSS 7.09e-19
C7869 VDD.t321 VSS 0.00375f
C7870 VDD.n1496 VSS 7.09e-19
C7871 VDD.t322 VSS 0.0017f
C7872 VDD.n1497 VSS 0.00171f
C7873 VDD.n1498 VSS 0.00272f
C7874 VDD.n1499 VSS 0.002f
C7875 VDD.n1500 VSS 0.00133f
C7876 VDD.n1501 VSS 7.19e-19
C7877 VDD.n1502 VSS 0.00408f
C7878 VDD.n1503 VSS 7.09e-19
C7879 VDD.n1504 VSS 0.00121f
C7880 VDD.n1505 VSS 0.002f
C7881 VDD.n1506 VSS 0.00121f
C7882 VDD.n1507 VSS 7.09e-19
C7883 VDD.n1508 VSS 0.00396f
C7884 VDD.n1509 VSS 7.09e-19
C7885 VDD.t320 VSS 6.28e-19
C7886 VDD.t700 VSS 0.00141f
C7887 VDD.n1510 VSS 0.00226f
C7888 VDD.n1511 VSS 0.00297f
C7889 VDD.n1512 VSS 0.002f
C7890 VDD.n1513 VSS 7.62e-19
C7891 VDD.n1514 VSS 7.09e-19
C7892 VDD.t701 VSS 0.00375f
C7893 VDD.n1515 VSS 7.09e-19
C7894 VDD.n1516 VSS 0.00116f
C7895 VDD.n1517 VSS 0.002f
C7896 VDD.n1518 VSS 9.79e-19
C7897 VDD.n1519 VSS 7.09e-19
C7898 VDD.n1520 VSS 0.00588f
C7899 VDD.n1521 VSS 7.09e-19
C7900 VDD.n1522 VSS 7.76e-19
C7901 VDD.t412 VSS 3.92e-19
C7902 VDD.t353 VSS 3.92e-19
C7903 VDD.n1523 VSS 8.47e-19
C7904 VDD.n1524 VSS 9.79e-19
C7905 VDD.n1525 VSS 7.09e-19
C7906 VDD.t565 VSS 0.00375f
C7907 VDD.n1526 VSS 7.18e-19
C7908 VDD.n1527 VSS 0.0013f
C7909 VDD.n1528 VSS 0.002f
C7910 VDD.n1529 VSS 0.00116f
C7911 VDD.n1530 VSS 7.09e-19
C7912 VDD.t36 VSS 0.00375f
C7913 VDD.n1531 VSS 7.09e-19
C7914 VDD.t37 VSS 5.95e-19
C7915 VDD.t398 VSS -3.29e-19
C7916 VDD.n1532 VSS 0.00233f
C7917 VDD.n1533 VSS 0.00159f
C7918 VDD.n1534 VSS 0.002f
C7919 VDD.t31 VSS 0.0017f
C7920 VDD.n1535 VSS 0.00171f
C7921 VDD.n1536 VSS 7.09e-19
C7922 VDD.t147 VSS 0.00375f
C7923 VDD.n1537 VSS 7.19e-19
C7924 VDD.n1538 VSS 0.00133f
C7925 VDD.n1539 VSS 0.00102f
C7926 VDD.n1540 VSS 0.002f
C7927 VDD.n1541 VSS 0.00121f
C7928 VDD.n1542 VSS 7.09e-19
C7929 VDD.n1543 VSS 0.00588f
C7930 VDD.n1544 VSS 7.09e-19
C7931 VDD.n1545 VSS 0.00121f
C7932 VDD.n1546 VSS 0.002f
C7933 VDD.t33 VSS 6.28e-19
C7934 VDD.t144 VSS 0.00141f
C7935 VDD.n1547 VSS 0.00226f
C7936 VDD.n1548 VSS 0.00297f
C7937 VDD.n1549 VSS 7.09e-19
C7938 VDD.n1550 VSS 0.00428f
C7939 VDD.n1551 VSS 7.09e-19
C7940 VDD.n1552 VSS 7.62e-19
C7941 VDD.n1553 VSS 6.7e-19
C7942 VDD.n1554 VSS 0.002f
C7943 VDD.t146 VSS 3.52e-19
C7944 VDD.t150 VSS 3.71e-19
C7945 VDD.n1555 VSS 7.74e-19
C7946 VDD.n1556 VSS 0.00116f
C7947 VDD.n1557 VSS 7.09e-19
C7948 VDD.t697 VSS 0.00375f
C7949 VDD.n1558 VSS 7.09e-19
C7950 VDD.n1559 VSS 9.79e-19
C7951 VDD.n1560 VSS 0.002f
C7952 VDD.t680 VSS 9.19e-19
C7953 VDD.n1561 VSS 7.76e-19
C7954 VDD.n1562 VSS 7.09e-19
C7955 VDD.t618 VSS 0.00302f
C7956 VDD.n1563 VSS 7.09e-19
C7957 VDD.n1564 VSS 9.79e-19
C7958 VDD.n1565 VSS 0.002f
C7959 VDD.t158 VSS 5.51e-19
C7960 VDD.t263 VSS -1.76e-19
C7961 VDD.n1566 VSS 0.00259f
C7962 VDD.n1567 VSS 0.00235f
C7963 VDD.n1568 VSS 0.0013f
C7964 VDD.n1569 VSS 7.18e-19
C7965 VDD.n1570 VSS 0.006f
C7966 VDD.n1571 VSS 7.09e-19
C7967 VDD.n1572 VSS 0.00116f
C7968 VDD.n1573 VSS 0.002f
C7969 VDD.t316 VSS 5.95e-19
C7970 VDD.t162 VSS -3.29e-19
C7971 VDD.n1574 VSS 0.00233f
C7972 VDD.n1575 VSS 0.00159f
C7973 VDD.n1576 VSS 7.09e-19
C7974 VDD.t421 VSS 0.00375f
C7975 VDD.n1577 VSS 7.09e-19
C7976 VDD.t422 VSS 0.0017f
C7977 VDD.n1578 VSS 0.00171f
C7978 VDD.n1579 VSS 0.00272f
C7979 VDD.n1580 VSS 0.002f
C7980 VDD.n1581 VSS 0.00133f
C7981 VDD.n1582 VSS 7.19e-19
C7982 VDD.n1583 VSS 0.00408f
C7983 VDD.n1584 VSS 7.09e-19
C7984 VDD.n1585 VSS 0.00121f
C7985 VDD.n1586 VSS 0.002f
C7986 VDD.n1587 VSS 0.00121f
C7987 VDD.n1588 VSS 7.09e-19
C7988 VDD.n1589 VSS 0.00396f
C7989 VDD.n1590 VSS 7.09e-19
C7990 VDD.t424 VSS 6.28e-19
C7991 VDD.t358 VSS 0.00141f
C7992 VDD.n1591 VSS 0.00226f
C7993 VDD.n1592 VSS 0.00297f
C7994 VDD.n1593 VSS 0.002f
C7995 VDD.n1594 VSS 7.62e-19
C7996 VDD.n1595 VSS 7.09e-19
C7997 VDD.t359 VSS 0.00375f
C7998 VDD.n1596 VSS 7.09e-19
C7999 VDD.n1597 VSS 0.00116f
C8000 VDD.n1598 VSS 0.002f
C8001 VDD.n1599 VSS 9.79e-19
C8002 VDD.n1600 VSS 7.09e-19
C8003 VDD.n1601 VSS 0.00588f
C8004 VDD.n1602 VSS 7.09e-19
C8005 VDD.n1603 VSS 7.76e-19
C8006 VDD.t19 VSS 3.92e-19
C8007 VDD.t463 VSS 3.92e-19
C8008 VDD.n1604 VSS 8.47e-19
C8009 VDD.n1605 VSS 7.19e-19
C8010 VDD.t462 VSS 0.00375f
C8011 VDD.n1606 VSS 0.00343f
C8012 VDD.t18 VSS 0.00302f
C8013 VDD.n1607 VSS 0.00235f
C8014 VDD.n1608 VSS 0.00102f
C8015 VDD.n1609 VSS 0.00131f
C8016 VDD.n1610 VSS 0.00176f
C8017 VDD.n1611 VSS 0.00181f
C8018 VDD.n1612 VSS 0.002f
C8019 VDD.n1613 VSS 0.002f
C8020 VDD.t376 VSS 9.19e-19
C8021 VDD.n1614 VSS 0.002f
C8022 VDD.n1615 VSS 0.00132f
C8023 VDD.n1616 VSS 7.19e-19
C8024 VDD.n1617 VSS 0.00555f
C8025 VDD.t375 VSS 0.00375f
C8026 VDD.n1618 VSS 0.00379f
C8027 VDD.t260 VSS 0.00375f
C8028 VDD.n1619 VSS 0.0049f
C8029 VDD.t461 VSS 0.00375f
C8030 VDD.n1620 VSS 0.00343f
C8031 VDD.n1621 VSS 7.09e-19
C8032 VDD.n1622 VSS 0.00121f
C8033 VDD.n1623 VSS 0.002f
C8034 VDD.n1624 VSS 0.002f
C8035 VDD.n1625 VSS 0.002f
C8036 VDD.n1626 VSS 0.002f
C8037 VDD.t360 VSS 3.52e-19
C8038 VDD.t272 VSS 3.71e-19
C8039 VDD.n1627 VSS 7.74e-19
C8040 VDD.n1628 VSS 0.0018f
C8041 VDD.n1629 VSS 0.00133f
C8042 VDD.n1630 VSS 7.19e-19
C8043 VDD.n1631 VSS 0.00432f
C8044 VDD.t271 VSS 0.00375f
C8045 VDD.n1632 VSS 0.00428f
C8046 VDD.t423 VSS 0.00363f
C8047 VDD.t202 VSS 0.00355f
C8048 VDD.n1633 VSS 0.00388f
C8049 VDD.n1634 VSS 7.09e-19
C8050 VDD.n1635 VSS 0.00121f
C8051 VDD.n1636 VSS 6.7e-19
C8052 VDD.n1637 VSS 0.002f
C8053 VDD.n1638 VSS 0.002f
C8054 VDD.n1639 VSS 7.1e-19
C8055 VDD.n1640 VSS 7.09e-19
C8056 VDD.n1641 VSS 0.00539f
C8057 VDD.t357 VSS 0.00375f
C8058 VDD.n1642 VSS 0.00588f
C8059 VDD.t261 VSS 0.00375f
C8060 VDD.t460 VSS 0.00718f
C8061 VDD.n1643 VSS 7.09e-19
C8062 VDD.n1644 VSS 0.00121f
C8063 VDD.n1645 VSS 0.002f
C8064 VDD.n1646 VSS 0.002f
C8065 VDD.t160 VSS 3.71e-19
C8066 VDD.t274 VSS 3.71e-19
C8067 VDD.n1647 VSS 7.84e-19
C8068 VDD.n1648 VSS 0.00164f
C8069 VDD.n1649 VSS 0.002f
C8070 VDD.n1650 VSS 0.002f
C8071 VDD.n1651 VSS 8.61e-19
C8072 VDD.n1652 VSS 7.09e-19
C8073 VDD.n1653 VSS 0.00449f
C8074 VDD.t159 VSS 0.00375f
C8075 VDD.n1654 VSS 0.00441f
C8076 VDD.t273 VSS 0.00375f
C8077 VDD.n1655 VSS 0.00294f
C8078 VDD.t142 VSS 0.00375f
C8079 VDD.n1656 VSS 0.00392f
C8080 VDD.n1657 VSS 7.09e-19
C8081 VDD.n1658 VSS 0.00106f
C8082 VDD.n1659 VSS 0.00102f
C8083 VDD.n1660 VSS 0.002f
C8084 VDD.n1661 VSS 0.002f
C8085 VDD.n1662 VSS 0.00188f
C8086 VDD.n1663 VSS 7.09e-19
C8087 VDD.n1664 VSS 0.00677f
C8088 VDD.n1665 VSS 0.00506f
C8089 VDD.t315 VSS 0.00375f
C8090 VDD.t161 VSS 0.00375f
C8091 VDD.n1666 VSS 0.00396f
C8092 VDD.n1667 VSS 7.09e-19
C8093 VDD.n1668 VSS 0.00121f
C8094 VDD.n1669 VSS 0.002f
C8095 VDD.n1670 VSS 0.002f
C8096 VDD.n1671 VSS 0.002f
C8097 VDD.n1672 VSS 0.00105f
C8098 VDD.n1673 VSS 7.09e-19
C8099 VDD.n1674 VSS 0.00543f
C8100 VDD.t157 VSS 0.00375f
C8101 VDD.n1675 VSS 0.00388f
C8102 VDD.t262 VSS 0.00375f
C8103 VDD.n1676 VSS 0.00379f
C8104 VDD.n1677 VSS 0.00571f
C8105 VDD.n1678 VSS 7.09e-19
C8106 VDD.n1679 VSS 9.79e-19
C8107 VDD.n1680 VSS 0.0015f
C8108 VDD.n1681 VSS 6.96e-19
C8109 VDD.n1682 VSS 0.00181f
C8110 VDD.t619 VSS 3.92e-19
C8111 VDD.t15 VSS 3.92e-19
C8112 VDD.n1683 VSS 8.47e-19
C8113 VDD.n1684 VSS 0.00176f
C8114 VDD.n1685 VSS 0.00131f
C8115 VDD.n1686 VSS 7.19e-19
C8116 VDD.n1687 VSS 0.00343f
C8117 VDD.t14 VSS 0.00375f
C8118 VDD.n1688 VSS 0.00588f
C8119 VDD.n1689 VSS 0.00379f
C8120 VDD.t679 VSS 0.00375f
C8121 VDD.n1690 VSS 0.00555f
C8122 VDD.n1691 VSS 7.19e-19
C8123 VDD.n1692 VSS 0.00132f
C8124 VDD.n1693 VSS 0.002f
C8125 VDD.n1694 VSS 0.002f
C8126 VDD.n1695 VSS 0.002f
C8127 VDD.n1696 VSS 0.002f
C8128 VDD.n1697 VSS 0.00121f
C8129 VDD.n1698 VSS 7.09e-19
C8130 VDD.n1699 VSS 0.00343f
C8131 VDD.t13 VSS 0.00375f
C8132 VDD.n1700 VSS 0.0049f
C8133 VDD.t145 VSS 0.00375f
C8134 VDD.t149 VSS 0.00375f
C8135 VDD.n1701 VSS 0.00432f
C8136 VDD.n1702 VSS 7.19e-19
C8137 VDD.n1703 VSS 0.00133f
C8138 VDD.n1704 VSS 0.0018f
C8139 VDD.n1705 VSS 0.002f
C8140 VDD.n1706 VSS 0.002f
C8141 VDD.n1707 VSS 0.002f
C8142 VDD.n1708 VSS 0.00121f
C8143 VDD.n1709 VSS 7.09e-19
C8144 VDD.n1710 VSS 0.00388f
C8145 VDD.t528 VSS 0.00355f
C8146 VDD.t32 VSS 0.00363f
C8147 VDD.n1711 VSS 0.00396f
C8148 VDD.t143 VSS 0.00375f
C8149 VDD.n1712 VSS 0.00539f
C8150 VDD.n1713 VSS 7.09e-19
C8151 VDD.n1714 VSS 7.1e-19
C8152 VDD.n1715 VSS 0.002f
C8153 VDD.n1716 VSS 0.002f
C8154 VDD.n1717 VSS 0.002f
C8155 VDD.n1718 VSS 0.00121f
C8156 VDD.n1719 VSS 7.09e-19
C8157 VDD.t12 VSS 0.00718f
C8158 VDD.t698 VSS 0.00375f
C8159 VDD.n1720 VSS 0.00408f
C8160 VDD.n1721 VSS 0.00441f
C8161 VDD.t395 VSS 0.00375f
C8162 VDD.n1722 VSS 0.00449f
C8163 VDD.n1723 VSS 7.09e-19
C8164 VDD.n1724 VSS 8.61e-19
C8165 VDD.n1725 VSS 0.002f
C8166 VDD.t396 VSS 3.71e-19
C8167 VDD.t148 VSS 3.71e-19
C8168 VDD.n1726 VSS 7.84e-19
C8169 VDD.n1727 VSS 0.00164f
C8170 VDD.n1728 VSS 0.002f
C8171 VDD.n1729 VSS 0.002f
C8172 VDD.n1730 VSS 0.002f
C8173 VDD.n1731 VSS 0.00106f
C8174 VDD.n1732 VSS 7.09e-19
C8175 VDD.n1733 VSS 0.00392f
C8176 VDD.t457 VSS 0.00375f
C8177 VDD.n1734 VSS 0.00294f
C8178 VDD.t30 VSS 0.00375f
C8179 VDD.n1735 VSS 0.00506f
C8180 VDD.n1736 VSS 0.00677f
C8181 VDD.n1737 VSS 7.09e-19
C8182 VDD.n1738 VSS 0.00188f
C8183 VDD.n1739 VSS 0.00272f
C8184 VDD.n1740 VSS 0.002f
C8185 VDD.n1741 VSS 0.002f
C8186 VDD.n1742 VSS 0.00121f
C8187 VDD.n1743 VSS 7.09e-19
C8188 VDD.n1744 VSS 0.00396f
C8189 VDD.t397 VSS 0.00375f
C8190 VDD.n1745 VSS 0.006f
C8191 VDD.n1746 VSS 0.00388f
C8192 VDD.t399 VSS 0.00375f
C8193 VDD.n1747 VSS 0.00543f
C8194 VDD.n1748 VSS 7.09e-19
C8195 VDD.n1749 VSS 0.00105f
C8196 VDD.n1750 VSS 0.002f
C8197 VDD.t400 VSS 5.51e-19
C8198 VDD.t566 VSS -1.76e-19
C8199 VDD.n1751 VSS 0.00259f
C8200 VDD.n1752 VSS 0.00235f
C8201 VDD.n1753 VSS 0.002f
C8202 VDD.n1754 VSS 6.96e-19
C8203 VDD.n1755 VSS 0.0015f
C8204 VDD.n1756 VSS 9.79e-19
C8205 VDD.n1757 VSS 7.09e-19
C8206 VDD.n1758 VSS 0.00571f
C8207 VDD.n1759 VSS 0.00379f
C8208 VDD.t411 VSS 0.00302f
C8209 VDD.t352 VSS 0.00375f
C8210 VDD.n1760 VSS 0.00343f
C8211 VDD.n1761 VSS 7.19e-19
C8212 VDD.n1762 VSS 0.00131f
C8213 VDD.n1763 VSS 0.00176f
C8214 VDD.n1764 VSS 0.00181f
C8215 VDD.n1765 VSS 0.002f
C8216 VDD.n1766 VSS 0.002f
C8217 VDD.t678 VSS 9.19e-19
C8218 VDD.n1767 VSS 0.002f
C8219 VDD.n1768 VSS 0.00132f
C8220 VDD.n1769 VSS 7.19e-19
C8221 VDD.n1770 VSS 0.00555f
C8222 VDD.t677 VSS 0.00375f
C8223 VDD.n1771 VSS 0.00379f
C8224 VDD.t633 VSS 0.00375f
C8225 VDD.n1772 VSS 0.0049f
C8226 VDD.t354 VSS 0.00375f
C8227 VDD.n1773 VSS 0.00343f
C8228 VDD.n1774 VSS 7.09e-19
C8229 VDD.n1775 VSS 0.00121f
C8230 VDD.n1776 VSS 0.002f
C8231 VDD.n1777 VSS 0.002f
C8232 VDD.n1778 VSS 0.002f
C8233 VDD.n1779 VSS 0.002f
C8234 VDD.t702 VSS 3.52e-19
C8235 VDD.t650 VSS 3.71e-19
C8236 VDD.n1780 VSS 7.74e-19
C8237 VDD.n1781 VSS 0.0018f
C8238 VDD.n1782 VSS 0.00133f
C8239 VDD.n1783 VSS 7.19e-19
C8240 VDD.n1784 VSS 0.00432f
C8241 VDD.t649 VSS 0.00375f
C8242 VDD.n1785 VSS 0.00428f
C8243 VDD.t319 VSS 0.00363f
C8244 VDD.t201 VSS 0.00355f
C8245 VDD.n1786 VSS 0.00388f
C8246 VDD.n1787 VSS 7.09e-19
C8247 VDD.n1788 VSS 0.00121f
C8248 VDD.n1789 VSS 6.7e-19
C8249 VDD.n1790 VSS 0.002f
C8250 VDD.n1791 VSS 0.002f
C8251 VDD.n1792 VSS 7.1e-19
C8252 VDD.n1793 VSS 7.09e-19
C8253 VDD.n1794 VSS 0.00539f
C8254 VDD.t699 VSS 0.00375f
C8255 VDD.n1795 VSS 0.00588f
C8256 VDD.t632 VSS 0.00375f
C8257 VDD.t351 VSS 0.00718f
C8258 VDD.n1796 VSS 7.09e-19
C8259 VDD.n1797 VSS 0.00121f
C8260 VDD.n1798 VSS 0.002f
C8261 VDD.n1799 VSS 0.002f
C8262 VDD.t54 VSS 3.71e-19
C8263 VDD.t648 VSS 3.71e-19
C8264 VDD.n1800 VSS 7.84e-19
C8265 VDD.n1801 VSS 0.00164f
C8266 VDD.n1802 VSS 0.002f
C8267 VDD.n1803 VSS 0.002f
C8268 VDD.n1804 VSS 8.61e-19
C8269 VDD.n1805 VSS 7.09e-19
C8270 VDD.n1806 VSS 0.00449f
C8271 VDD.t53 VSS 0.00375f
C8272 VDD.n1807 VSS 0.00441f
C8273 VDD.t647 VSS 0.00375f
C8274 VDD.n1808 VSS 0.00294f
C8275 VDD.t716 VSS 0.00375f
C8276 VDD.n1809 VSS 0.00392f
C8277 VDD.n1810 VSS 7.09e-19
C8278 VDD.n1811 VSS 0.00106f
C8279 VDD.n1812 VSS 0.00102f
C8280 VDD.n1813 VSS 0.002f
C8281 VDD.n1814 VSS 0.002f
C8282 VDD.n1815 VSS 0.00188f
C8283 VDD.n1816 VSS 7.09e-19
C8284 VDD.n1817 VSS 0.00677f
C8285 VDD.n1818 VSS 0.00506f
C8286 VDD.t626 VSS 0.00375f
C8287 VDD.t55 VSS 0.00375f
C8288 VDD.n1819 VSS 0.00396f
C8289 VDD.n1820 VSS 7.09e-19
C8290 VDD.n1821 VSS 0.00121f
C8291 VDD.n1822 VSS 0.002f
C8292 VDD.n1823 VSS 0.002f
C8293 VDD.n1824 VSS 0.002f
C8294 VDD.n1825 VSS 0.00105f
C8295 VDD.n1826 VSS 7.09e-19
C8296 VDD.n1827 VSS 0.00543f
C8297 VDD.t57 VSS 0.00375f
C8298 VDD.n1828 VSS 0.00388f
C8299 VDD.t377 VSS 0.00375f
C8300 VDD.n1829 VSS 0.00379f
C8301 VDD.n1830 VSS 0.00571f
C8302 VDD.n1831 VSS 7.09e-19
C8303 VDD.n1832 VSS 9.79e-19
C8304 VDD.n1833 VSS 0.0015f
C8305 VDD.n1834 VSS 6.96e-19
C8306 VDD.n1835 VSS 0.00181f
C8307 VDD.t676 VSS 3.92e-19
C8308 VDD.t431 VSS 3.92e-19
C8309 VDD.n1836 VSS 8.47e-19
C8310 VDD.n1837 VSS 0.00176f
C8311 VDD.n1838 VSS 0.00131f
C8312 VDD.n1839 VSS 7.19e-19
C8313 VDD.n1840 VSS 0.00343f
C8314 VDD.t430 VSS 0.00375f
C8315 VDD.n1841 VSS 0.00588f
C8316 VDD.n1842 VSS 0.00379f
C8317 VDD.t435 VSS 0.00375f
C8318 VDD.n1843 VSS 0.00555f
C8319 VDD.n1844 VSS 7.19e-19
C8320 VDD.n1845 VSS 0.00132f
C8321 VDD.n1846 VSS 0.002f
C8322 VDD.n1847 VSS 0.002f
C8323 VDD.n1848 VSS 0.002f
C8324 VDD.n1849 VSS 0.002f
C8325 VDD.n1850 VSS 0.00121f
C8326 VDD.n1851 VSS 7.09e-19
C8327 VDD.n1852 VSS 0.00343f
C8328 VDD.t429 VSS 0.00375f
C8329 VDD.n1853 VSS 0.0049f
C8330 VDD.t8 VSS 0.00375f
C8331 VDD.t543 VSS 0.00375f
C8332 VDD.n1854 VSS 0.00432f
C8333 VDD.n1855 VSS 7.19e-19
C8334 VDD.n1856 VSS 0.00133f
C8335 VDD.n1857 VSS 0.0018f
C8336 VDD.n1858 VSS 0.002f
C8337 VDD.n1859 VSS 0.002f
C8338 VDD.n1860 VSS 0.002f
C8339 VDD.n1861 VSS 0.00121f
C8340 VDD.n1862 VSS 7.09e-19
C8341 VDD.n1863 VSS 0.00388f
C8342 VDD.t437 VSS 0.00355f
C8343 VDD.t638 VSS 0.00363f
C8344 VDD.n1864 VSS 0.00396f
C8345 VDD.t10 VSS 0.00375f
C8346 VDD.n1865 VSS 0.00539f
C8347 VDD.n1866 VSS 7.09e-19
C8348 VDD.n1867 VSS 7.1e-19
C8349 VDD.n1868 VSS 0.002f
C8350 VDD.n1869 VSS 0.002f
C8351 VDD.n1870 VSS 0.002f
C8352 VDD.n1871 VSS 0.00121f
C8353 VDD.n1872 VSS 7.09e-19
C8354 VDD.t432 VSS 0.00718f
C8355 VDD.t102 VSS 0.00375f
C8356 VDD.n1873 VSS 0.00408f
C8357 VDD.n1874 VSS 0.00441f
C8358 VDD.t711 VSS 0.00375f
C8359 VDD.n1875 VSS 0.00449f
C8360 VDD.n1876 VSS 7.09e-19
C8361 VDD.n1877 VSS 8.61e-19
C8362 VDD.n1878 VSS 0.002f
C8363 VDD.t712 VSS 3.71e-19
C8364 VDD.t546 VSS 3.71e-19
C8365 VDD.n1879 VSS 7.84e-19
C8366 VDD.n1880 VSS 0.00164f
C8367 VDD.n1881 VSS 0.002f
C8368 VDD.n1882 VSS 0.002f
C8369 VDD.n1883 VSS 0.002f
C8370 VDD.n1884 VSS 0.00106f
C8371 VDD.n1885 VSS 7.09e-19
C8372 VDD.n1886 VSS 0.00392f
C8373 VDD.t95 VSS 0.00375f
C8374 VDD.n1887 VSS 0.00294f
C8375 VDD.t640 VSS 0.00375f
C8376 VDD.n1888 VSS 0.00506f
C8377 VDD.n1889 VSS 0.00677f
C8378 VDD.n1890 VSS 7.09e-19
C8379 VDD.n1891 VSS 0.00188f
C8380 VDD.n1892 VSS 0.00272f
C8381 VDD.n1893 VSS 0.002f
C8382 VDD.n1894 VSS 0.002f
C8383 VDD.n1895 VSS 0.00121f
C8384 VDD.n1896 VSS 7.09e-19
C8385 VDD.n1897 VSS 0.00396f
C8386 VDD.t707 VSS 0.00375f
C8387 VDD.n1898 VSS 0.006f
C8388 VDD.n1899 VSS 0.00388f
C8389 VDD.t709 VSS 0.00375f
C8390 VDD.n1900 VSS 0.00543f
C8391 VDD.n1901 VSS 7.09e-19
C8392 VDD.n1902 VSS 0.00105f
C8393 VDD.n1903 VSS 0.002f
C8394 VDD.t710 VSS 5.51e-19
C8395 VDD.t126 VSS -1.76e-19
C8396 VDD.n1904 VSS 0.00259f
C8397 VDD.n1905 VSS 0.00235f
C8398 VDD.n1906 VSS 0.002f
C8399 VDD.n1907 VSS 6.96e-19
C8400 VDD.n1908 VSS 0.0015f
C8401 VDD.n1909 VSS 9.79e-19
C8402 VDD.n1910 VSS 7.09e-19
C8403 VDD.n1911 VSS 0.00571f
C8404 VDD.n1912 VSS 0.00379f
C8405 VDD.t40 VSS 0.00302f
C8406 VDD.t723 VSS 0.00375f
C8407 VDD.n1913 VSS 0.00343f
C8408 VDD.n1914 VSS 7.19e-19
C8409 VDD.n1915 VSS 0.00131f
C8410 VDD.n1916 VSS 0.00176f
C8411 VDD.n1917 VSS 0.00181f
C8412 VDD.n1918 VSS 0.002f
C8413 VDD.n1919 VSS 0.002f
C8414 VDD.t118 VSS 9.19e-19
C8415 VDD.n1920 VSS 0.002f
C8416 VDD.n1921 VSS 0.00132f
C8417 VDD.n1922 VSS 7.19e-19
C8418 VDD.n1923 VSS 0.00555f
C8419 VDD.t117 VSS 0.00375f
C8420 VDD.n1924 VSS 0.00379f
C8421 VDD.t163 VSS 0.00375f
C8422 VDD.n1925 VSS 0.0049f
C8423 VDD.t721 VSS 0.00375f
C8424 VDD.n1926 VSS 0.00343f
C8425 VDD.n1927 VSS 7.09e-19
C8426 VDD.n1928 VSS 0.00121f
C8427 VDD.n1929 VSS 0.002f
C8428 VDD.n1930 VSS 0.002f
C8429 VDD.n1931 VSS 0.002f
C8430 VDD.n1932 VSS 0.002f
C8431 VDD.t720 VSS 3.52e-19
C8432 VDD.t568 VSS 3.71e-19
C8433 VDD.n1933 VSS 7.74e-19
C8434 VDD.n1934 VSS 0.0018f
C8435 VDD.n1935 VSS 0.00133f
C8436 VDD.n1936 VSS 7.19e-19
C8437 VDD.n1937 VSS 0.00432f
C8438 VDD.t567 VSS 0.00375f
C8439 VDD.n1938 VSS 0.00428f
C8440 VDD.t693 VSS 0.00363f
C8441 VDD.t121 VSS 0.00355f
C8442 VDD.n1939 VSS 0.00388f
C8443 VDD.n1940 VSS 7.09e-19
C8444 VDD.n1941 VSS 0.00121f
C8445 VDD.n1942 VSS 6.7e-19
C8446 VDD.n1943 VSS 0.002f
C8447 VDD.n1944 VSS 0.002f
C8448 VDD.n1945 VSS 7.1e-19
C8449 VDD.n1946 VSS 7.09e-19
C8450 VDD.n1947 VSS 0.00539f
C8451 VDD.t717 VSS 0.00375f
C8452 VDD.n1948 VSS 0.00588f
C8453 VDD.t164 VSS 0.00375f
C8454 VDD.t722 VSS 0.00718f
C8455 VDD.n1949 VSS 7.09e-19
C8456 VDD.n1950 VSS 0.00121f
C8457 VDD.n1951 VSS 0.002f
C8458 VDD.n1952 VSS 0.002f
C8459 VDD.t331 VSS 3.71e-19
C8460 VDD.t570 VSS 3.71e-19
C8461 VDD.n1953 VSS 7.84e-19
C8462 VDD.n1954 VSS 0.00164f
C8463 VDD.n1955 VSS 0.002f
C8464 VDD.n1956 VSS 0.002f
C8465 VDD.n1957 VSS 8.61e-19
C8466 VDD.n1958 VSS 7.09e-19
C8467 VDD.n1959 VSS 0.00449f
C8468 VDD.t330 VSS 0.00375f
C8469 VDD.n1960 VSS 0.00441f
C8470 VDD.t569 VSS 0.00375f
C8471 VDD.n1961 VSS 0.00294f
C8472 VDD.t387 VSS 0.00375f
C8473 VDD.n1962 VSS 0.00392f
C8474 VDD.n1963 VSS 7.09e-19
C8475 VDD.n1964 VSS 0.00106f
C8476 VDD.n1965 VSS 0.00102f
C8477 VDD.n1966 VSS 0.002f
C8478 VDD.n1967 VSS 0.002f
C8479 VDD.n1968 VSS 0.00188f
C8480 VDD.n1969 VSS 7.09e-19
C8481 VDD.n1970 VSS 0.00677f
C8482 VDD.n1971 VSS 0.00506f
C8483 VDD.t442 VSS 0.00375f
C8484 VDD.t328 VSS 0.00375f
C8485 VDD.n1972 VSS 0.00396f
C8486 VDD.n1973 VSS 7.09e-19
C8487 VDD.n1974 VSS 0.00121f
C8488 VDD.n1975 VSS 0.002f
C8489 VDD.n1976 VSS 0.002f
C8490 VDD.n1977 VSS 0.002f
C8491 VDD.n1978 VSS 0.00105f
C8492 VDD.n1979 VSS 7.09e-19
C8493 VDD.n1980 VSS 0.00543f
C8494 VDD.t326 VSS 0.00375f
C8495 VDD.n1981 VSS 0.00388f
C8496 VDD.t592 VSS 0.00429f
C8497 VDD.n1982 VSS 0.00883f
C8498 VDD.n1983 VSS 9.79e-19
C8499 VDD.n1984 VSS 0.0015f
C8500 VDD.n1985 VSS 1.62f
C8501 VDD.n1986 VSS 0.736f
C8502 VDD.n1987 VSS 0.002f
C8503 VDD.t21 VSS 5.19e-19
C8504 VDD.t656 VSS 5.19e-19
C8505 VDD.n1988 VSS 0.00126f
C8506 VDD.n1989 VSS 0.00238f
C8507 VDD.n1990 VSS 0.00131f
C8508 VDD.n1991 VSS 7.19e-19
C8509 VDD.n1992 VSS 7.09e-19
C8510 VDD.n1993 VSS 0.002f
C8511 VDD.n1994 VSS 9.47e-19
C8512 VDD.n1995 VSS 7.09e-19
C8513 VDD.n1996 VSS 0.0316f
C8514 VDD.t652 VSS 0.00247f
C8515 VDD.n1997 VSS 0.002f
C8516 VDD.n1998 VSS 0.00119f
C8517 VDD.t583 VSS 0.00285f
C8518 VDD.n1999 VSS 7.09e-19
C8519 VDD.t584 VSS 0.00377f
C8520 VDD.n2000 VSS 7.09e-19
C8521 VDD.n2001 VSS 6.38e-19
C8522 VDD.t581 VSS 9.75e-19
C8523 VDD.t579 VSS 6.12e-19
C8524 VDD.n2002 VSS 0.00204f
C8525 VDD.n2003 VSS 0.00274f
C8526 VDD.n2004 VSS 6.24e-19
C8527 VDD.n2005 VSS 0.002f
C8528 VDD.n2006 VSS 0.00121f
C8529 VDD.t129 VSS 5.8e-19
C8530 VDD.t585 VSS 2.83e-19
C8531 VDD.n2007 VSS 0.00209f
C8532 VDD.n2008 VSS 0.00167f
C8533 VDD.n2009 VSS 7.09e-19
C8534 VDD.n2010 VSS 0.00427f
C8535 VDD.n2011 VSS 7.09e-19
C8536 VDD.n2012 VSS 8.48e-19
C8537 VDD.n2013 VSS 0.002f
C8538 VDD.t447 VSS 0.00146f
C8539 VDD.n2014 VSS 0.00112f
C8540 VDD.n2015 VSS 7.09e-19
C8541 VDD.t52 VSS 0.00377f
C8542 VDD.n2016 VSS 7.09e-19
C8543 VDD.n2017 VSS 0.00121f
C8544 VDD.n2018 VSS 0.002f
C8545 VDD.t86 VSS 3.92e-19
C8546 VDD.t658 VSS 3.92e-19
C8547 VDD.n2019 VSS 8.4e-19
C8548 VDD.n2020 VSS 0.00176f
C8549 VDD.n2021 VSS 7.09e-19
C8550 VDD.t433 VSS 0.00377f
C8551 VDD.n2022 VSS 7.09e-19
C8552 VDD.n2023 VSS 0.00121f
C8553 VDD.n2024 VSS 8.48e-19
C8554 VDD.n2025 VSS 0.00181f
C8555 VDD.t704 VSS 3.92e-19
C8556 VDD.t60 VSS 3.92e-19
C8557 VDD.n2026 VSS 8.24e-19
C8558 VDD.n2027 VSS 0.00142f
C8559 VDD.n2028 VSS 0.00131f
C8560 VDD.n2029 VSS 7.19e-19
C8561 VDD.n2030 VSS 0.00102f
C8562 VDD.n2031 VSS 0.00684f
C8563 VDD.t703 VSS 0.00304f
C8564 VDD.n2032 VSS 0.00345f
C8565 VDD.t59 VSS 0.00377f
C8566 VDD.n2033 VSS 0.00345f
C8567 VDD.t671 VSS 0.00377f
C8568 VDD.n2034 VSS 0.00394f
C8569 VDD.n2035 VSS 7.09e-19
C8570 VDD.n2036 VSS 0.00101f
C8571 VDD.n2037 VSS 0.002f
C8572 VDD.n2038 VSS 0.002f
C8573 VDD.n2039 VSS 0.002f
C8574 VDD.n2040 VSS 0.00121f
C8575 VDD.n2041 VSS 7.09e-19
C8576 VDD.n2042 VSS 0.00591f
C8577 VDD.t85 VSS 0.00377f
C8578 VDD.n2043 VSS 0.00345f
C8579 VDD.t657 VSS 0.00377f
C8580 VDD.n2044 VSS 0.00722f
C8581 VDD.n2045 VSS 0.00427f
C8582 VDD.n2046 VSS 7.09e-19
C8583 VDD.n2047 VSS 9.66e-19
C8584 VDD.n2048 VSS 0.002f
C8585 VDD.n2049 VSS 0.002f
C8586 VDD.n2050 VSS 0.002f
C8587 VDD.n2051 VSS 0.00121f
C8588 VDD.n2052 VSS 7.09e-19
C8589 VDD.n2053 VSS 0.00345f
C8590 VDD.t61 VSS 0.00377f
C8591 VDD.n2054 VSS 0.00443f
C8592 VDD.t446 VSS 0.00377f
C8593 VDD.n2055 VSS 0.00706f
C8594 VDD.n2056 VSS 7.19e-19
C8595 VDD.n2057 VSS 0.00132f
C8596 VDD.n2058 VSS 0.00236f
C8597 VDD.n2059 VSS 0.002f
C8598 VDD.n2060 VSS 0.002f
C8599 VDD.n2061 VSS 0.002f
C8600 VDD.n2062 VSS 0.00121f
C8601 VDD.n2063 VSS 7.09e-19
C8602 VDD.n2064 VSS 0.00505f
C8603 VDD.t434 VSS 0.00377f
C8604 VDD.n2065 VSS 0.00345f
C8605 VDD.t672 VSS 0.00377f
C8606 VDD.n2066 VSS 0.00398f
C8607 VDD.t128 VSS 0.00377f
C8608 VDD.n2067 VSS 0.00414f
C8609 VDD.n2068 VSS 7.09e-19
C8610 VDD.n2069 VSS 0.00118f
C8611 VDD.n2070 VSS 0.002f
C8612 VDD.n2071 VSS 0.002f
C8613 VDD.n2072 VSS 0.002f
C8614 VDD.n2073 VSS 0.002f
C8615 VDD.n2074 VSS 0.00121f
C8616 VDD.n2075 VSS 7.09e-19
C8617 VDD.n2076 VSS 0.00345f
C8618 VDD.t580 VSS 0.00377f
C8619 VDD.n2077 VSS 0.0041f
C8620 VDD.t578 VSS 0.00377f
C8621 VDD.t582 VSS 0.00377f
C8622 VDD.n2078 VSS 0.00345f
C8623 VDD.n2079 VSS 7.09e-19
C8624 VDD.n2080 VSS 7.09e-19
C8625 VDD.n2081 VSS 0.00398f
C8626 VDD.n2082 VSS 0.0015f
C8627 VDD.n2083 VSS 0.002f
C8628 VDD.n2084 VSS 0.0082f
C8629 VDD.n2085 VSS 0.00386f
C8630 VDD.n2086 VSS 7.09e-19
C8631 VDD.n2087 VSS 0.0311f
C8632 VDD.t651 VSS 0.00377f
C8633 VDD.n2088 VSS 0.00345f
C8634 VDD.t653 VSS 0.00377f
C8635 VDD.n2089 VSS 0.00267f
C8636 VDD.t409 VSS 0.00377f
C8637 VDD.n2090 VSS 0.0039f
C8638 VDD.n2091 VSS 7.19e-19
C8639 VDD.t654 VSS -8.35e-21
C8640 VDD.t410 VSS 5.22e-19
C8641 VDD.n2092 VSS 0.00241f
C8642 VDD.n2093 VSS 0.00238f
C8643 VDD.n2094 VSS 0.00131f
C8644 VDD.n2095 VSS 5.46e-19
C8645 VDD.n2096 VSS 0.0015f
C8646 VDD.n2097 VSS 0.0015f
C8647 VDD.n2098 VSS 8.81e-19
C8648 VDD.n2099 VSS 7.09e-19
C8649 VDD.n2100 VSS 0.00505f
C8650 VDD.t20 VSS 0.00377f
C8651 VDD.n2101 VSS 0.00361f
C8652 VDD.t655 VSS 0.00377f
C8653 VDD.n2102 VSS 0.00267f
C8654 VDD.n2103 VSS 7.09e-19
C8655 VDD.n2104 VSS 9.93e-19
C8656 VDD.n2105 VSS 0.00119f
C8657 VDD.n2106 VSS 0.325f
C8658 VDD.n2107 VSS 0.00118f
C8659 VDD.t23 VSS 3.92e-19
C8660 VDD.t621 VSS 3.92e-19
C8661 VDD.n2108 VSS 8.47e-19
C8662 VDD.t22 VSS 0.00376f
C8663 VDD.n2109 VSS 9.79e-19
C8664 VDD.n2110 VSS 7.09e-19
C8665 VDD.n2111 VSS 6.95e-19
C8666 VDD.t620 VSS 0.00372f
C8667 VDD.n2112 VSS 0.00344f
C8668 VDD.n2113 VSS 7.19e-19
C8669 VDD.n2114 VSS 0.00131f
C8670 VDD.n2115 VSS 0.00176f
C8671 VDD.n2116 VSS 0.002f
C8672 VDD.n2117 VSS 0.00589f
C8673 VDD.n2118 VSS 7.09e-19
C8674 VDD.n2119 VSS 7.76e-19
C8675 VDD.n2120 VSS 0.002f
C8676 VDD.t595 VSS 9.19e-19
C8677 VDD.t594 VSS 0.00376f
C8678 VDD.n2121 VSS 0.00556f
C8679 VDD.n2122 VSS 7.19e-19
C8680 VDD.n2123 VSS 0.00132f
C8681 VDD.n2124 VSS 0.002f
C8682 VDD.n2125 VSS 0.002f
C8683 VDD.t714 VSS 0.00376f
C8684 VDD.n2126 VSS 0.0038f
C8685 VDD.n2127 VSS 7.09e-19
C8686 VDD.n2128 VSS 9.79e-19
C8687 VDD.n2129 VSS 0.002f
C8688 VDD.t24 VSS 0.00376f
C8689 VDD.n2130 VSS 0.00344f
C8690 VDD.n2131 VSS 7.09e-19
C8691 VDD.n2132 VSS 0.00121f
C8692 VDD.n2133 VSS 0.002f
C8693 VDD.n2134 VSS 0.00491f
C8694 VDD.n2135 VSS 7.09e-19
C8695 VDD.n2136 VSS 0.00116f
C8696 VDD.n2137 VSS 0.002f
C8697 VDD.t629 VSS 3.71e-19
C8698 VDD.t540 VSS 3.52e-19
C8699 VDD.n2138 VSS 7.74e-19
C8700 VDD.t539 VSS 0.00376f
C8701 VDD.n2139 VSS 0.00434f
C8702 VDD.n2140 VSS 7.19e-19
C8703 VDD.n2141 VSS 0.00133f
C8704 VDD.n2142 VSS 0.0018f
C8705 VDD.n2143 VSS 0.002f
C8706 VDD.t628 VSS 0.00376f
C8707 VDD.n2144 VSS 0.0043f
C8708 VDD.n2145 VSS 7.09e-19
C8709 VDD.n2146 VSS 7.62e-19
C8710 VDD.n2147 VSS 0.002f
C8711 VDD.t124 VSS 0.00356f
C8712 VDD.n2148 VSS 0.00389f
C8713 VDD.n2149 VSS 7.09e-19
C8714 VDD.n2150 VSS 0.00121f
C8715 VDD.n2151 VSS 0.002f
C8716 VDD.t542 VSS 0.00141f
C8717 VDD.t465 VSS 6.28e-19
C8718 VDD.n2152 VSS 0.00226f
C8719 VDD.n2153 VSS 0.00297f
C8720 VDD.t464 VSS 0.00364f
C8721 VDD.n2154 VSS 0.00397f
C8722 VDD.n2155 VSS 7.09e-19
C8723 VDD.n2156 VSS 6.7e-19
C8724 VDD.n2157 VSS 0.002f
C8725 VDD.t541 VSS 0.00376f
C8726 VDD.n2158 VSS 0.0054f
C8727 VDD.n2159 VSS 7.09e-19
C8728 VDD.n2160 VSS 7.1e-19
C8729 VDD.n2161 VSS 0.002f
C8730 VDD.n2162 VSS 0.00589f
C8731 VDD.n2163 VSS 7.09e-19
C8732 VDD.n2164 VSS 0.00121f
C8733 VDD.n2165 VSS 0.002f
C8734 VDD.t25 VSS 0.0072f
C8735 VDD.n2166 VSS 7.09e-19
C8736 VDD.n2167 VSS 0.00121f
C8737 VDD.n2168 VSS 0.002f
C8738 VDD.t715 VSS 0.00376f
C8739 VDD.n2169 VSS 0.00409f
C8740 VDD.n2170 VSS 7.09e-19
C8741 VDD.n2171 VSS 0.00121f
C8742 VDD.n2172 VSS 0.002f
C8743 VDD.t191 VSS 0.00376f
C8744 VDD.n2173 VSS 0.0045f
C8745 VDD.n2174 VSS 7.09e-19
C8746 VDD.n2175 VSS 8.61e-19
C8747 VDD.n2176 VSS 0.002f
C8748 VDD.t449 VSS 3.71e-19
C8749 VDD.t192 VSS 3.71e-19
C8750 VDD.n2177 VSS 7.84e-19
C8751 VDD.t448 VSS 0.00376f
C8752 VDD.n2178 VSS 0.00442f
C8753 VDD.n2179 VSS 7.19e-19
C8754 VDD.n2180 VSS 0.00133f
C8755 VDD.n2181 VSS 0.00164f
C8756 VDD.n2182 VSS 0.002f
C8757 VDD.t705 VSS 0.00376f
C8758 VDD.n2183 VSS 0.00393f
C8759 VDD.n2184 VSS 7.09e-19
C8760 VDD.n2185 VSS 0.00106f
C8761 VDD.n2186 VSS 0.002f
C8762 VDD.t466 VSS 0.00376f
C8763 VDD.n2187 VSS 0.00295f
C8764 VDD.n2188 VSS 7.09e-19
C8765 VDD.n2189 VSS 0.00102f
C8766 VDD.n2190 VSS 0.002f
C8767 VDD.t255 VSS 0.00904f
C8768 VDD.n2191 VSS 0.0081f
C8769 VDD.n2192 VSS 8.71e-19
C8770 VDD.t467 VSS 0.0017f
C8771 VDD.n2193 VSS 0.00171f
C8772 VDD.n2194 VSS 0.00185f
C8773 VDD.n2195 VSS 0.00198f
C8774 VDD.n2196 VSS 0.001f
C8775 VDD.t732 VSS 5.71e-19
C8776 VDD.n2197 VSS 0.00159f
C8777 VDD.t254 VSS 0.00104f
C8778 VDD.n2198 VSS 0.00217f
C8779 VDD.n2199 VSS 4.77e-19
C8780 VDD.n2200 VSS 0.0014f
C8781 VDD.n2201 VSS 2.58e-19
C8782 VDD.n2202 VSS 1.85e-19
C8783 VDD.n2203 VSS 0.001f
C8784 VDD.t190 VSS -3.29e-19
C8785 VDD.t256 VSS 5.95e-19
C8786 VDD.n2204 VSS 0.00233f
C8787 VDD.n2205 VSS 0.00134f
C8788 VDD.n2206 VSS 0.00121f
C8789 VDD.n2207 VSS 0.00184f
C8790 VDD.t189 VSS 0.00622f
C8791 VDD.n2208 VSS 0.00601f
C8792 VDD.n2209 VSS 0.0011f
C8793 VDD.n2210 VSS 0.00116f
C8794 VDD.n2211 VSS 0.002f
C8795 VDD.t193 VSS 0.00376f
C8796 VDD.n2212 VSS 0.00544f
C8797 VDD.n2213 VSS 7.09e-19
C8798 VDD.n2214 VSS 0.00105f
C8799 VDD.n2215 VSS 0.002f
C8800 VDD.t208 VSS -1.76e-19
C8801 VDD.t194 VSS 5.51e-19
C8802 VDD.n2216 VSS 0.00259f
C8803 VDD.t207 VSS 0.00376f
C8804 VDD.n2217 VSS 0.00389f
C8805 VDD.n2218 VSS 7.18e-19
C8806 VDD.n2219 VSS 0.0013f
C8807 VDD.n2220 VSS 0.00235f
C8808 VDD.n2221 VSS 0.002f
C8809 VDD.n2222 VSS 0.0015f
C8810 VDD.n2223 VSS 9.79e-19
C8811 VDD.n2224 VSS 9.79e-19
C8812 VDD.n2225 VSS 7.09e-19
C8813 VDD.n2226 VSS 6.95e-19
C8814 VDD.t622 VSS 0.00372f
C8815 VDD.n2227 VSS 0.00344f
C8816 VDD.n2228 VSS 7.19e-19
C8817 VDD.n2229 VSS 0.0012f
C8818 VDD.n2230 VSS 0.00176f
C8819 VDD.n2231 VSS 0.00182f
C8820 VDD.n2232 VSS 0.001f
C8821 VDD.n2233 VSS 3.68e-19
C8822 VDD.n2234 VSS 1.12e-19
C8823 VDD.n2235 VSS 3.51e-19
C8824 VDD.n2236 VSS 6.55e-20
C8825 VDD.n2237 VSS 0.00372f
C8826 VDD.n2238 VSS 6.95e-19
C8827 VDD.n2239 VSS 0.00217f
C8828 VDD.n2240 VSS 3.58e-19
C8829 VDD.n2241 VSS 4.01e-19
C8830 VDD.n2242 VSS 1.18e-19
C8831 VDD.n2243 VSS 0.00119f
C8832 VDD.t394 VSS 9.19e-19
C8833 VDD.t393 VSS 0.00376f
C8834 VDD.n2244 VSS 0.00487f
C8835 VDD.n2245 VSS 6.53e-19
C8836 VDD.n2246 VSS 0.00121f
C8837 VDD.n2247 VSS 0.002f
C8838 VDD.n2248 VSS 0.002f
C8839 VDD.t524 VSS 0.00376f
C8840 VDD.n2249 VSS 0.0038f
C8841 VDD.n2250 VSS 7.09e-19
C8842 VDD.n2251 VSS 9.79e-19
C8843 VDD.n2252 VSS 0.002f
C8844 VDD.t522 VSS 0.00376f
C8845 VDD.n2253 VSS 0.00344f
C8846 VDD.n2254 VSS 7.09e-19
C8847 VDD.n2255 VSS 0.00121f
C8848 VDD.n2256 VSS 0.002f
C8849 VDD.t62 VSS 0.007f
C8850 VDD.n2257 VSS 0.00491f
C8851 VDD.n2258 VSS 0.00124f
C8852 VDD.n2259 VSS 0.00116f
C8853 VDD.n2260 VSS 0.002f
C8854 VDD.n2261 VSS 0.00128f
C8855 VDD.t250 VSS 3.71e-19
C8856 VDD.t63 VSS 3.52e-19
C8857 VDD.n2262 VSS 7.72e-19
C8858 VDD.n2263 VSS 0.00183f
C8859 VDD.n2264 VSS 0.00193f
C8860 VDD.n2265 VSS 0.001f
C8861 VDD.n2266 VSS 6.05e-19
C8862 VDD.t251 VSS 9.65e-19
C8863 VDD.t725 VSS 4.09e-19
C8864 VDD.n2267 VSS 0.00196f
C8865 VDD.n2268 VSS 8.02e-19
C8866 VDD.n2269 VSS 0.00248f
C8867 VDD.n2270 VSS 1.83e-19
C8868 VDD.n2271 VSS 1.51e-19
C8869 VDD.n2272 VSS 8.86e-20
C8870 VDD.n2273 VSS 1.11e-19
C8871 VDD.n2274 VSS 2.1e-19
C8872 VDD.n2275 VSS 5.34e-19
C8873 VDD.t741 VSS 4.1e-19
C8874 VDD.n2276 VSS 0.00182f
C8875 VDD.t248 VSS 0.00122f
C8876 VDD.n2277 VSS 9.88e-19
C8877 VDD.n2278 VSS 1.46e-19
C8878 VDD.n2279 VSS 1.12e-19
C8879 VDD.n2280 VSS 1.85e-19
C8880 VDD.n2281 VSS 0.001f
C8881 VDD.t264 VSS 0.00356f
C8882 VDD.t249 VSS 0.00863f
C8883 VDD.n2282 VSS 0.00442f
C8884 VDD.n2283 VSS 7.48e-19
C8885 VDD.n2284 VSS 0.00114f
C8886 VDD.n2285 VSS 0.00189f
C8887 VDD.t65 VSS 0.00141f
C8888 VDD.t204 VSS 6.28e-19
C8889 VDD.n2286 VSS 0.00226f
C8890 VDD.n2287 VSS 0.00297f
C8891 VDD.t203 VSS 0.00364f
C8892 VDD.n2288 VSS 0.00397f
C8893 VDD.n2289 VSS 7.09e-19
C8894 VDD.n2290 VSS 6.7e-19
C8895 VDD.n2291 VSS 0.002f
C8896 VDD.t64 VSS 0.00376f
C8897 VDD.n2292 VSS 0.0054f
C8898 VDD.n2293 VSS 7.09e-19
C8899 VDD.n2294 VSS 7.1e-19
C8900 VDD.n2295 VSS 0.002f
C8901 VDD.n2296 VSS 0.00589f
C8902 VDD.n2297 VSS 7.09e-19
C8903 VDD.n2298 VSS 0.00121f
C8904 VDD.n2299 VSS 0.002f
C8905 VDD.t523 VSS 0.0072f
C8906 VDD.n2300 VSS 7.09e-19
C8907 VDD.n2301 VSS 0.00121f
C8908 VDD.n2302 VSS 0.002f
C8909 VDD.t525 VSS 0.00376f
C8910 VDD.n2303 VSS 0.00409f
C8911 VDD.n2304 VSS 7.09e-19
C8912 VDD.n2305 VSS 0.00121f
C8913 VDD.n2306 VSS 0.002f
C8914 VDD.t685 VSS 0.00376f
C8915 VDD.n2307 VSS 0.0045f
C8916 VDD.n2308 VSS 7.09e-19
C8917 VDD.n2309 VSS 8.61e-19
C8918 VDD.n2310 VSS 0.002f
C8919 VDD.t253 VSS 3.71e-19
C8920 VDD.t686 VSS 3.71e-19
C8921 VDD.n2311 VSS 7.84e-19
C8922 VDD.t252 VSS 0.00376f
C8923 VDD.n2312 VSS 0.00442f
C8924 VDD.n2313 VSS 7.19e-19
C8925 VDD.n2314 VSS 0.00133f
C8926 VDD.n2315 VSS 0.00164f
C8927 VDD.n2316 VSS 0.002f
C8928 VDD.t127 VSS 0.00376f
C8929 VDD.n2317 VSS 0.00393f
C8930 VDD.n2318 VSS 7.09e-19
C8931 VDD.n2319 VSS 0.00106f
C8932 VDD.n2320 VSS 0.002f
C8933 VDD.t205 VSS 0.00376f
C8934 VDD.n2321 VSS 0.00295f
C8935 VDD.n2322 VSS 7.09e-19
C8936 VDD.n2323 VSS 0.00102f
C8937 VDD.n2324 VSS 0.002f
C8938 VDD.n2325 VSS 0.00679f
C8939 VDD.n2326 VSS 7.09e-19
C8940 VDD.t206 VSS 0.0017f
C8941 VDD.n2327 VSS 0.00171f
C8942 VDD.n2328 VSS 0.00188f
C8943 VDD.n2329 VSS 0.002f
C8944 VDD.t324 VSS 0.00376f
C8945 VDD.n2330 VSS 0.00507f
C8946 VDD.n2331 VSS 7.09e-19
C8947 VDD.n2332 VSS 0.00272f
C8948 VDD.n2333 VSS 0.002f
C8949 VDD.t683 VSS 0.00376f
C8950 VDD.n2334 VSS 0.00397f
C8951 VDD.n2335 VSS 7.09e-19
C8952 VDD.t684 VSS -3.29e-19
C8953 VDD.t325 VSS 5.95e-19
C8954 VDD.n2336 VSS 0.00233f
C8955 VDD.n2337 VSS 0.00159f
C8956 VDD.n2338 VSS 0.00121f
C8957 VDD.n2339 VSS 0.002f
C8958 VDD.n2340 VSS 0.00601f
C8959 VDD.n2341 VSS 7.09e-19
C8960 VDD.n2342 VSS 0.00116f
C8961 VDD.n2343 VSS 0.002f
C8962 VDD.t681 VSS 0.00376f
C8963 VDD.n2344 VSS 0.00544f
C8964 VDD.n2345 VSS 7.09e-19
C8965 VDD.n2346 VSS 0.00105f
C8966 VDD.n2347 VSS 0.002f
C8967 VDD.t97 VSS -1.76e-19
C8968 VDD.t682 VSS 5.51e-19
C8969 VDD.n2348 VSS 0.00259f
C8970 VDD.t96 VSS 0.00376f
C8971 VDD.n2349 VSS 0.00389f
C8972 VDD.n2350 VSS 7.18e-19
C8973 VDD.n2351 VSS 0.0013f
C8974 VDD.n2352 VSS 0.00235f
C8975 VDD.n2353 VSS 0.002f
C8976 VDD.n2354 VSS 0.0015f
C8977 VDD.n2355 VSS 9.79e-19
C8978 VDD.n2356 VSS 9.79e-19
C8979 VDD.n2357 VSS 7.09e-19
C8980 VDD.n2358 VSS 6.95e-19
C8981 VDD.t407 VSS 0.00372f
C8982 VDD.n2359 VSS 0.00344f
C8983 VDD.n2360 VSS 7.19e-19
C8984 VDD.n2361 VSS 0.00131f
C8985 VDD.n2362 VSS 0.00176f
C8986 VDD.n2363 VSS 0.002f
C8987 VDD.n2364 VSS 0.00589f
C8988 VDD.n2365 VSS 7.09e-19
C8989 VDD.n2366 VSS 7.76e-19
C8990 VDD.n2367 VSS 0.002f
C8991 VDD.t674 VSS 9.19e-19
C8992 VDD.t673 VSS 0.00376f
C8993 VDD.n2368 VSS 0.00556f
C8994 VDD.n2369 VSS 7.19e-19
C8995 VDD.n2370 VSS 0.00132f
C8996 VDD.n2371 VSS 0.002f
C8997 VDD.n2372 VSS 0.002f
C8998 VDD.t588 VSS 0.00376f
C8999 VDD.n2373 VSS 0.0038f
C9000 VDD.n2374 VSS 7.09e-19
C9001 VDD.n2375 VSS 9.79e-19
C9002 VDD.n2376 VSS 0.002f
C9003 VDD.t391 VSS 0.00376f
C9004 VDD.n2377 VSS 0.00344f
C9005 VDD.n2378 VSS 7.09e-19
C9006 VDD.n2379 VSS 0.00121f
C9007 VDD.n2380 VSS 0.002f
C9008 VDD.t553 VSS 0.007f
C9009 VDD.n2381 VSS 0.00491f
C9010 VDD.n2382 VSS 0.00124f
C9011 VDD.n2383 VSS 0.00116f
C9012 VDD.n2384 VSS 0.002f
C9013 VDD.n2385 VSS 0.00128f
C9014 VDD.t214 VSS 3.71e-19
C9015 VDD.t554 VSS 3.52e-19
C9016 VDD.n2386 VSS 7.72e-19
C9017 VDD.n2387 VSS 0.00183f
C9018 VDD.n2388 VSS 0.00193f
C9019 VDD.n2389 VSS 0.001f
C9020 VDD.n2390 VSS 6.05e-19
C9021 VDD.t257 VSS 9.65e-19
C9022 VDD.t740 VSS 4.09e-19
C9023 VDD.n2391 VSS 0.00196f
C9024 VDD.n2392 VSS 8.02e-19
C9025 VDD.n2393 VSS 0.00248f
C9026 VDD.n2394 VSS 1.83e-19
C9027 VDD.n2395 VSS 1.51e-19
C9028 VDD.n2396 VSS 8.86e-20
C9029 VDD.n2397 VSS 1.11e-19
C9030 VDD.n2398 VSS 2.1e-19
C9031 VDD.n2399 VSS 5.34e-19
C9032 VDD.t737 VSS 4.1e-19
C9033 VDD.n2400 VSS 0.00182f
C9034 VDD.t212 VSS 0.00122f
C9035 VDD.n2401 VSS 9.95e-19
C9036 VDD.n2402 VSS 1.47e-19
C9037 VDD.n2403 VSS 1.12e-19
C9038 VDD.n2404 VSS 1.85e-19
C9039 VDD.n2405 VSS 0.001f
C9040 VDD.t538 VSS 0.00356f
C9041 VDD.t213 VSS 0.00863f
C9042 VDD.n2406 VSS 0.00442f
C9043 VDD.n2407 VSS 7.48e-19
C9044 VDD.n2408 VSS 0.00114f
C9045 VDD.n2409 VSS 0.00189f
C9046 VDD.t552 VSS 0.00141f
C9047 VDD.t99 VSS 6.28e-19
C9048 VDD.n2410 VSS 0.00226f
C9049 VDD.n2411 VSS 0.00297f
C9050 VDD.t98 VSS 0.00364f
C9051 VDD.n2412 VSS 0.00397f
C9052 VDD.n2413 VSS 7.09e-19
C9053 VDD.n2414 VSS 6.7e-19
C9054 VDD.n2415 VSS 0.002f
C9055 VDD.t551 VSS 0.00376f
C9056 VDD.n2416 VSS 0.0054f
C9057 VDD.n2417 VSS 7.09e-19
C9058 VDD.n2418 VSS 7.1e-19
C9059 VDD.n2419 VSS 0.002f
C9060 VDD.n2420 VSS 0.00589f
C9061 VDD.n2421 VSS 7.09e-19
C9062 VDD.n2422 VSS 0.00121f
C9063 VDD.n2423 VSS 0.002f
C9064 VDD.t392 VSS 0.0072f
C9065 VDD.n2424 VSS 7.09e-19
C9066 VDD.n2425 VSS 0.00121f
C9067 VDD.n2426 VSS 0.002f
C9068 VDD.t589 VSS 0.00376f
C9069 VDD.n2427 VSS 0.00409f
C9070 VDD.n2428 VSS 7.09e-19
C9071 VDD.n2429 VSS 0.00121f
C9072 VDD.n2430 VSS 0.002f
C9073 VDD.t365 VSS 0.00376f
C9074 VDD.n2431 VSS 0.0045f
C9075 VDD.n2432 VSS 7.09e-19
C9076 VDD.n2433 VSS 8.61e-19
C9077 VDD.n2434 VSS 0.002f
C9078 VDD.t259 VSS 3.71e-19
C9079 VDD.t366 VSS 3.71e-19
C9080 VDD.n2435 VSS 7.84e-19
C9081 VDD.t258 VSS 0.00376f
C9082 VDD.n2436 VSS 0.00442f
C9083 VDD.n2437 VSS 7.19e-19
C9084 VDD.n2438 VSS 0.00133f
C9085 VDD.n2439 VSS 0.00164f
C9086 VDD.n2440 VSS 0.002f
C9087 VDD.t289 VSS 0.00376f
C9088 VDD.n2441 VSS 0.00393f
C9089 VDD.n2442 VSS 7.09e-19
C9090 VDD.n2443 VSS 0.00106f
C9091 VDD.n2444 VSS 0.002f
C9092 VDD.t100 VSS 0.00376f
C9093 VDD.n2445 VSS 0.00295f
C9094 VDD.n2446 VSS 7.09e-19
C9095 VDD.n2447 VSS 0.00102f
C9096 VDD.n2448 VSS 0.002f
C9097 VDD.n2449 VSS 0.00679f
C9098 VDD.n2450 VSS 7.09e-19
C9099 VDD.t101 VSS 0.0017f
C9100 VDD.n2451 VSS 0.00171f
C9101 VDD.n2452 VSS 0.00188f
C9102 VDD.n2453 VSS 0.002f
C9103 VDD.t474 VSS 0.00376f
C9104 VDD.n2454 VSS 0.00507f
C9105 VDD.n2455 VSS 7.09e-19
C9106 VDD.n2456 VSS 0.00272f
C9107 VDD.n2457 VSS 0.002f
C9108 VDD.t361 VSS 0.00376f
C9109 VDD.n2458 VSS 0.00397f
C9110 VDD.n2459 VSS 7.09e-19
C9111 VDD.t362 VSS -3.29e-19
C9112 VDD.t475 VSS 5.95e-19
C9113 VDD.n2460 VSS 0.00233f
C9114 VDD.n2461 VSS 0.00159f
C9115 VDD.n2462 VSS 0.00121f
C9116 VDD.n2463 VSS 0.002f
C9117 VDD.n2464 VSS 0.00601f
C9118 VDD.n2465 VSS 7.09e-19
C9119 VDD.n2466 VSS 0.00116f
C9120 VDD.n2467 VSS 0.002f
C9121 VDD.t363 VSS 0.00376f
C9122 VDD.n2468 VSS 0.00544f
C9123 VDD.n2469 VSS 7.09e-19
C9124 VDD.n2470 VSS 0.00105f
C9125 VDD.n2471 VSS 0.002f
C9126 VDD.t591 VSS -1.76e-19
C9127 VDD.t364 VSS 5.51e-19
C9128 VDD.n2472 VSS 0.00259f
C9129 VDD.t590 VSS 0.00376f
C9130 VDD.n2473 VSS 0.00389f
C9131 VDD.n2474 VSS 7.18e-19
C9132 VDD.n2475 VSS 0.0013f
C9133 VDD.n2476 VSS 0.00235f
C9134 VDD.n2477 VSS 0.002f
C9135 VDD.n2478 VSS 0.0015f
C9136 VDD.n2479 VSS 9.79e-19
C9137 VDD.n2480 VSS 9.79e-19
C9138 VDD.n2481 VSS 7.09e-19
C9139 VDD.n2482 VSS 6.95e-19
C9140 VDD.t405 VSS 0.00372f
C9141 VDD.n2483 VSS 0.00344f
C9142 VDD.n2484 VSS 7.19e-19
C9143 VDD.n2485 VSS 0.00131f
C9144 VDD.n2486 VSS 0.00176f
C9145 VDD.n2487 VSS 0.002f
C9146 VDD.n2488 VSS 0.00589f
C9147 VDD.n2489 VSS 7.09e-19
C9148 VDD.n2490 VSS 7.76e-19
C9149 VDD.n2491 VSS 0.002f
C9150 VDD.t305 VSS 9.19e-19
C9151 VDD.t304 VSS 0.00376f
C9152 VDD.n2492 VSS 0.00556f
C9153 VDD.n2493 VSS 7.19e-19
C9154 VDD.n2494 VSS 0.00132f
C9155 VDD.n2495 VSS 0.002f
C9156 VDD.n2496 VSS 0.002f
C9157 VDD.t630 VSS 0.00376f
C9158 VDD.n2497 VSS 0.0038f
C9159 VDD.n2498 VSS 7.09e-19
C9160 VDD.n2499 VSS 9.79e-19
C9161 VDD.n2500 VSS 0.002f
C9162 VDD.t534 VSS 0.00376f
C9163 VDD.n2501 VSS 0.00344f
C9164 VDD.n2502 VSS 7.09e-19
C9165 VDD.n2503 VSS 0.00121f
C9166 VDD.n2504 VSS 0.002f
C9167 VDD.t425 VSS 0.007f
C9168 VDD.n2505 VSS 0.00491f
C9169 VDD.n2506 VSS 0.00124f
C9170 VDD.n2507 VSS 0.00116f
C9171 VDD.n2508 VSS 0.002f
C9172 VDD.n2509 VSS 0.00128f
C9173 VDD.t235 VSS 3.71e-19
C9174 VDD.t426 VSS 3.52e-19
C9175 VDD.n2510 VSS 7.72e-19
C9176 VDD.n2511 VSS 0.00183f
C9177 VDD.n2512 VSS 0.00193f
C9178 VDD.n2513 VSS 0.001f
C9179 VDD.n2514 VSS 6.05e-19
C9180 VDD.t221 VSS 9.65e-19
C9181 VDD.t736 VSS 4.09e-19
C9182 VDD.n2515 VSS 0.00196f
C9183 VDD.n2516 VSS 8.02e-19
C9184 VDD.n2517 VSS 0.00248f
C9185 VDD.n2518 VSS 1.83e-19
C9186 VDD.n2519 VSS 1.51e-19
C9187 VDD.n2520 VSS 8.86e-20
C9188 VDD.n2521 VSS 1.11e-19
C9189 VDD.n2522 VSS 2.1e-19
C9190 VDD.n2523 VSS 5.34e-19
C9191 VDD.t729 VSS 4.1e-19
C9192 VDD.n2524 VSS 0.00182f
C9193 VDD.t233 VSS 0.00122f
C9194 VDD.n2525 VSS 9.95e-19
C9195 VDD.n2526 VSS 1.47e-19
C9196 VDD.n2527 VSS 1.12e-19
C9197 VDD.n2528 VSS 1.85e-19
C9198 VDD.n2529 VSS 0.001f
C9199 VDD.t78 VSS 0.00356f
C9200 VDD.t234 VSS 0.00863f
C9201 VDD.n2530 VSS 0.00442f
C9202 VDD.n2531 VSS 7.48e-19
C9203 VDD.n2532 VSS 0.00114f
C9204 VDD.n2533 VSS 0.00189f
C9205 VDD.t428 VSS 0.00141f
C9206 VDD.t479 VSS 6.28e-19
C9207 VDD.n2534 VSS 0.00226f
C9208 VDD.n2535 VSS 0.00297f
C9209 VDD.t478 VSS 0.00364f
C9210 VDD.n2536 VSS 0.00397f
C9211 VDD.n2537 VSS 7.09e-19
C9212 VDD.n2538 VSS 6.7e-19
C9213 VDD.n2539 VSS 0.002f
C9214 VDD.t427 VSS 0.00376f
C9215 VDD.n2540 VSS 0.0054f
C9216 VDD.n2541 VSS 7.09e-19
C9217 VDD.n2542 VSS 7.1e-19
C9218 VDD.n2543 VSS 0.002f
C9219 VDD.n2544 VSS 0.00589f
C9220 VDD.n2545 VSS 7.09e-19
C9221 VDD.n2546 VSS 0.00121f
C9222 VDD.n2547 VSS 0.002f
C9223 VDD.t535 VSS 0.0072f
C9224 VDD.n2548 VSS 7.09e-19
C9225 VDD.n2549 VSS 0.00121f
C9226 VDD.n2550 VSS 0.002f
C9227 VDD.t631 VSS 0.00376f
C9228 VDD.n2551 VSS 0.00409f
C9229 VDD.n2552 VSS 7.09e-19
C9230 VDD.n2553 VSS 0.00121f
C9231 VDD.n2554 VSS 0.002f
C9232 VDD.t91 VSS 0.00376f
C9233 VDD.n2555 VSS 0.0045f
C9234 VDD.n2556 VSS 7.09e-19
C9235 VDD.n2557 VSS 8.61e-19
C9236 VDD.n2558 VSS 0.002f
C9237 VDD.t223 VSS 3.71e-19
C9238 VDD.t92 VSS 3.71e-19
C9239 VDD.n2559 VSS 7.84e-19
C9240 VDD.t222 VSS 0.00376f
C9241 VDD.n2560 VSS 0.00442f
C9242 VDD.n2561 VSS 7.19e-19
C9243 VDD.n2562 VSS 0.00133f
C9244 VDD.n2563 VSS 0.00164f
C9245 VDD.n2564 VSS 0.002f
C9246 VDD.t706 VSS 0.00376f
C9247 VDD.n2565 VSS 0.00393f
C9248 VDD.n2566 VSS 7.09e-19
C9249 VDD.n2567 VSS 0.00106f
C9250 VDD.n2568 VSS 0.002f
C9251 VDD.t476 VSS 0.00376f
C9252 VDD.n2569 VSS 0.00295f
C9253 VDD.n2570 VSS 7.09e-19
C9254 VDD.n2571 VSS 0.00102f
C9255 VDD.n2572 VSS 0.002f
C9256 VDD.n2573 VSS 0.00679f
C9257 VDD.n2574 VSS 7.09e-19
C9258 VDD.t477 VSS 0.0017f
C9259 VDD.n2575 VSS 0.00171f
C9260 VDD.n2576 VSS 0.00188f
C9261 VDD.n2577 VSS 0.002f
C9262 VDD.t413 VSS 0.00376f
C9263 VDD.n2578 VSS 0.00507f
C9264 VDD.n2579 VSS 7.09e-19
C9265 VDD.n2580 VSS 0.00272f
C9266 VDD.n2581 VSS 0.002f
C9267 VDD.t89 VSS 0.00376f
C9268 VDD.n2582 VSS 0.00397f
C9269 VDD.n2583 VSS 7.09e-19
C9270 VDD.t90 VSS -3.29e-19
C9271 VDD.t414 VSS 5.95e-19
C9272 VDD.n2584 VSS 0.00233f
C9273 VDD.n2585 VSS 0.00159f
C9274 VDD.n2586 VSS 0.00121f
C9275 VDD.n2587 VSS 0.002f
C9276 VDD.n2588 VSS 0.00601f
C9277 VDD.n2589 VSS 7.09e-19
C9278 VDD.n2590 VSS 0.00116f
C9279 VDD.n2591 VSS 0.002f
C9280 VDD.t93 VSS 0.00376f
C9281 VDD.n2592 VSS 0.00544f
C9282 VDD.n2593 VSS 7.09e-19
C9283 VDD.n2594 VSS 0.00105f
C9284 VDD.n2595 VSS 0.002f
C9285 VDD.t291 VSS -1.76e-19
C9286 VDD.t94 VSS 5.51e-19
C9287 VDD.n2596 VSS 0.00259f
C9288 VDD.t290 VSS 0.00376f
C9289 VDD.n2597 VSS 0.00389f
C9290 VDD.n2598 VSS 7.18e-19
C9291 VDD.n2599 VSS 0.0013f
C9292 VDD.n2600 VSS 0.00235f
C9293 VDD.n2601 VSS 0.002f
C9294 VDD.n2602 VSS 9.79e-19
C9295 VDD.t278 VSS 0.00376f
C9296 VDD.n2603 VSS 0.00961f
C9297 VDD.n2604 VSS 0.00108f
C9298 VDD.t356 VSS -1.76e-19
C9299 VDD.t664 VSS 5.51e-19
C9300 VDD.n2605 VSS 0.00259f
C9301 VDD.t355 VSS 0.00436f
C9302 VDD.n2606 VSS 0.00389f
C9303 VDD.n2607 VSS 7.18e-19
C9304 VDD.n2608 VSS 0.0013f
C9305 VDD.n2609 VSS 0.00235f
C9306 VDD.n2610 VSS 0.00467f
C9307 VDD.t663 VSS 0.00376f
C9308 VDD.n2611 VSS 0.00544f
C9309 VDD.n2612 VSS 7.09e-19
C9310 VDD.n2613 VSS 0.00105f
C9311 VDD.n2614 VSS 0.002f
C9312 VDD.n2615 VSS 0.00601f
C9313 VDD.n2616 VSS 7.09e-19
C9314 VDD.n2617 VSS 0.00116f
C9315 VDD.n2618 VSS 0.002f
C9316 VDD.t661 VSS 0.00376f
C9317 VDD.n2619 VSS 0.00397f
C9318 VDD.n2620 VSS 7.09e-19
C9319 VDD.t662 VSS -3.29e-19
C9320 VDD.t644 VSS 5.95e-19
C9321 VDD.n2621 VSS 0.00233f
C9322 VDD.n2622 VSS 0.00159f
C9323 VDD.n2623 VSS 0.00121f
C9324 VDD.n2624 VSS 0.002f
C9325 VDD.t643 VSS 0.00376f
C9326 VDD.n2625 VSS 0.00507f
C9327 VDD.n2626 VSS 7.09e-19
C9328 VDD.n2627 VSS 0.00272f
C9329 VDD.n2628 VSS 0.002f
C9330 VDD.n2629 VSS 0.00679f
C9331 VDD.n2630 VSS 7.09e-19
C9332 VDD.t515 VSS 0.0017f
C9333 VDD.n2631 VSS 0.00171f
C9334 VDD.n2632 VSS 0.00188f
C9335 VDD.n2633 VSS 0.002f
C9336 VDD.t514 VSS 0.00376f
C9337 VDD.n2634 VSS 0.00295f
C9338 VDD.n2635 VSS 7.09e-19
C9339 VDD.n2636 VSS 0.00102f
C9340 VDD.n2637 VSS 0.002f
C9341 VDD.t713 VSS 0.00376f
C9342 VDD.n2638 VSS 0.00393f
C9343 VDD.n2639 VSS 7.09e-19
C9344 VDD.n2640 VSS 0.00106f
C9345 VDD.n2641 VSS 0.002f
C9346 VDD.t229 VSS 3.71e-19
C9347 VDD.t660 VSS 3.71e-19
C9348 VDD.n2642 VSS 7.84e-19
C9349 VDD.t228 VSS 0.00376f
C9350 VDD.n2643 VSS 0.00442f
C9351 VDD.n2644 VSS 7.19e-19
C9352 VDD.n2645 VSS 0.00133f
C9353 VDD.n2646 VSS 0.00164f
C9354 VDD.n2647 VSS 0.002f
C9355 VDD.t659 VSS 0.00376f
C9356 VDD.n2648 VSS 0.0045f
C9357 VDD.n2649 VSS 7.09e-19
C9358 VDD.n2650 VSS 8.61e-19
C9359 VDD.n2651 VSS 0.002f
C9360 VDD.t87 VSS 0.00376f
C9361 VDD.n2652 VSS 0.00409f
C9362 VDD.n2653 VSS 7.09e-19
C9363 VDD.n2654 VSS 0.00121f
C9364 VDD.n2655 VSS 0.002f
C9365 VDD.t280 VSS 0.0072f
C9366 VDD.n2656 VSS 7.09e-19
C9367 VDD.n2657 VSS 0.00121f
C9368 VDD.n2658 VSS 0.002f
C9369 VDD.n2659 VSS 0.00589f
C9370 VDD.n2660 VSS 7.09e-19
C9371 VDD.n2661 VSS 0.00121f
C9372 VDD.n2662 VSS 0.002f
C9373 VDD.t153 VSS 0.00376f
C9374 VDD.n2663 VSS 0.0054f
C9375 VDD.n2664 VSS 7.09e-19
C9376 VDD.n2665 VSS 7.1e-19
C9377 VDD.n2666 VSS 0.002f
C9378 VDD.t154 VSS 0.00141f
C9379 VDD.t513 VSS 6.28e-19
C9380 VDD.n2667 VSS 0.00226f
C9381 VDD.n2668 VSS 0.00297f
C9382 VDD.t512 VSS 0.00364f
C9383 VDD.n2669 VSS 0.00397f
C9384 VDD.n2670 VSS 7.09e-19
C9385 VDD.n2671 VSS 6.7e-19
C9386 VDD.n2672 VSS 0.002f
C9387 VDD.t28 VSS 0.00356f
C9388 VDD.t231 VSS 0.00863f
C9389 VDD.n2673 VSS 0.00442f
C9390 VDD.n2674 VSS 7.48e-19
C9391 VDD.n2675 VSS 0.00114f
C9392 VDD.n2676 VSS 0.00189f
C9393 VDD.n2677 VSS 0.001f
C9394 VDD.n2678 VSS 6.05e-19
C9395 VDD.t227 VSS 9.65e-19
C9396 VDD.t731 VSS 4.09e-19
C9397 VDD.n2679 VSS 0.00196f
C9398 VDD.n2680 VSS 8.02e-19
C9399 VDD.n2681 VSS 0.00248f
C9400 VDD.n2682 VSS 1.83e-19
C9401 VDD.n2683 VSS 1.51e-19
C9402 VDD.n2684 VSS 8.86e-20
C9403 VDD.n2685 VSS 1.11e-19
C9404 VDD.n2686 VSS 2.1e-19
C9405 VDD.n2687 VSS 5.34e-19
C9406 VDD.t730 VSS 4.1e-19
C9407 VDD.n2688 VSS 0.00182f
C9408 VDD.t230 VSS 0.00122f
C9409 VDD.n2689 VSS 9.99e-19
C9410 VDD.n2690 VSS 1.48e-19
C9411 VDD.n2691 VSS 1.12e-19
C9412 VDD.n2692 VSS 1.85e-19
C9413 VDD.n2693 VSS 0.001f
C9414 VDD.n2694 VSS 0.00128f
C9415 VDD.t232 VSS 3.71e-19
C9416 VDD.t156 VSS 3.52e-19
C9417 VDD.n2695 VSS 7.72e-19
C9418 VDD.n2696 VSS 0.00183f
C9419 VDD.n2697 VSS 0.00193f
C9420 VDD.t155 VSS 0.007f
C9421 VDD.n2698 VSS 0.00491f
C9422 VDD.n2699 VSS 0.00124f
C9423 VDD.n2700 VSS 0.00116f
C9424 VDD.n2701 VSS 0.002f
C9425 VDD.t277 VSS 0.00376f
C9426 VDD.n2702 VSS 0.00344f
C9427 VDD.n2703 VSS 7.09e-19
C9428 VDD.n2704 VSS 0.00121f
C9429 VDD.n2705 VSS 0.002f
C9430 VDD.t88 VSS 0.00376f
C9431 VDD.n2706 VSS 0.0038f
C9432 VDD.n2707 VSS 7.09e-19
C9433 VDD.n2708 VSS 9.79e-19
C9434 VDD.n2709 VSS 0.002f
C9435 VDD.t416 VSS 9.19e-19
C9436 VDD.t415 VSS 0.00376f
C9437 VDD.n2710 VSS 0.00556f
C9438 VDD.n2711 VSS 7.19e-19
C9439 VDD.n2712 VSS 0.00132f
C9440 VDD.n2713 VSS 0.002f
C9441 VDD.n2714 VSS 0.002f
C9442 VDD.n2715 VSS 0.00589f
C9443 VDD.n2716 VSS 7.09e-19
C9444 VDD.n2717 VSS 7.76e-19
C9445 VDD.n2718 VSS 0.002f
C9446 VDD.n2719 VSS 0.00118f
C9447 VDD.n2720 VSS 0.002f
C9448 VDD.t279 VSS 3.92e-19
C9449 VDD.t453 VSS 3.92e-19
C9450 VDD.n2721 VSS 8.47e-19
C9451 VDD.n2722 VSS 0.00176f
C9452 VDD.n2723 VSS 0.00131f
C9453 VDD.n2724 VSS 7.19e-19
C9454 VDD.n2725 VSS 0.00344f
C9455 VDD.t452 VSS 0.00372f
C9456 VDD.n2726 VSS 7.09e-19
C9457 VDD.n2727 VSS 6.95e-19
C9458 VDD.n2728 VSS 0.00507f
C9459 VDD.n2729 VSS 7.09e-19
C9460 VDD.n2730 VSS 9.79e-19
C9461 VDD.n2731 VSS 0.0015f
.ends

