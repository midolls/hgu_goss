magic
tech sky130A
magscale 1 2
timestamp 1698742797
<< nwell >>
rect 415 744 437 787
rect 497 745 517 788
rect 547 745 601 786
rect 621 742 648 788
<< psubdiff >>
rect 415 204 648 208
rect 415 166 468 204
rect 506 166 556 204
rect 594 166 648 204
rect 415 162 648 166
<< nsubdiff >>
rect 415 784 648 788
rect 415 746 468 784
rect 506 746 556 784
rect 594 746 648 784
rect 415 742 648 746
<< psubdiffcont >>
rect 468 166 506 204
rect 556 166 594 204
<< nsubdiffcont >>
rect 468 746 506 784
rect 556 746 594 784
<< poly >>
rect 516 435 546 451
rect 454 419 546 435
rect 454 385 470 419
rect 504 385 546 419
rect 454 372 546 385
rect 454 369 516 372
<< polycont >>
rect 470 385 504 419
<< locali >>
rect 415 784 648 788
rect 415 746 468 784
rect 506 746 556 784
rect 594 746 648 784
rect 415 742 648 746
rect 454 385 470 419
rect 504 385 520 419
rect 558 334 592 537
rect 470 208 504 258
rect 415 204 648 208
rect 415 166 468 204
rect 506 166 556 204
rect 594 166 648 204
rect 415 162 648 166
<< viali >>
rect 468 746 506 784
rect 556 746 594 784
rect 470 385 504 419
rect 468 166 506 204
rect 556 166 594 204
<< metal1 >>
rect 415 784 648 790
rect 415 746 468 784
rect 506 746 556 784
rect 594 746 648 784
rect 415 740 648 746
rect 415 679 648 711
rect 470 646 504 679
rect 454 419 520 429
rect 454 385 470 419
rect 504 385 520 419
rect 454 375 520 385
rect 415 204 648 210
rect 415 166 468 204
rect 506 166 556 204
rect 594 166 648 204
rect 415 160 648 166
use sky130_fd_pr__nfet_01v8_L8T3GD  sky130_fd_pr__nfet_01v8_L8T3GD_0 /foss/designs/hgu_goss/hgu/mag
timestamp 1697868789
transform 1 0 531 0 1 264
box -73 -28 73 108
use sky130_fd_pr__pfet_01v8_MQX2PY  XM2
timestamp 1698734556
transform 1 0 531 0 1 592
box -152 -152 153 232
<< labels >>
flabel locali 566 388 586 424 0 FreeSans 160 0 0 0 OUT
port 15 nsew
flabel metal1 429 689 456 704 0 FreeSans 160 0 0 0 VREF
port 19 nsew
flabel metal1 422 749 457 774 0 FreeSans 160 0 0 0 VDD
port 22 nsew
flabel metal1 426 174 460 196 0 FreeSans 160 0 0 0 VSS
port 24 nsew
flabel metal1 470 385 504 419 0 FreeSans 160 0 0 0 IN
port 26 nsew
<< end >>
