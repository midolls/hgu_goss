* NGSPICE file created from hgu_cdac_8bit_array_flat.ext - technology: sky130A

.subckt hgu_cdac_8bit_array_flat SUB
C0 x1.CTOP x1.CBOT 0.647p
C1 x1.CBOT SUB 31.9f $ **FLOATING
C2 x1.CTOP SUB 56.2f $ **FLOATING
.ends

