magic
tech sky130A
magscale 1 2
timestamp 1699109888
<< nwell >>
rect 9760 2388 15943 2993
rect 9262 2021 15943 2388
rect 9760 1813 15943 2021
rect 9760 1662 15989 1813
rect 10436 1629 10654 1662
rect 11168 1629 11512 1662
rect 12380 1629 12724 1662
rect 13592 1629 13936 1662
rect 14804 1629 15148 1662
rect 15578 1644 15989 1662
rect 15578 1643 15797 1644
<< pwell >>
rect 9342 1781 9528 1963
rect 9532 1781 9718 1963
rect 9342 1777 9363 1781
rect 9329 1743 9363 1777
rect 9697 1777 9718 1781
rect 9697 1743 9731 1777
<< nmos >>
rect 10883 1477 10913 1561
rect 11615 1477 11645 1561
rect 11737 1477 11767 1561
rect 12827 1477 12857 1561
rect 12949 1477 12979 1561
rect 14165 1477 14195 1561
rect 14287 1477 14317 1561
rect 15021 1477 15051 1561
rect 15673 1478 15703 1562
rect 15765 1478 15795 1562
rect 15861 1478 15891 1562
rect 9863 1293 9893 1377
rect 9935 1293 9965 1377
rect 15673 1340 15703 1424
rect 9863 1155 9893 1239
rect 9935 1155 9965 1239
rect 9863 1017 9893 1101
rect 9935 1017 9965 1101
rect 9863 879 9893 963
rect 9935 879 9965 963
rect 9863 741 9893 825
rect 9935 741 9965 825
rect 9863 603 9893 687
rect 9935 603 9965 687
rect 9863 465 9893 549
rect 9935 465 9965 549
rect 9863 327 9893 411
rect 9935 327 9965 411
<< scnmos >>
rect 9420 1807 9450 1937
rect 9610 1807 9640 1937
<< pmos >>
rect 10530 1678 10560 1762
rect 11262 1678 11292 1762
rect 11388 1678 11418 1762
rect 12474 1678 12504 1762
rect 12600 1678 12630 1762
rect 13686 1678 13716 1762
rect 13812 1678 13842 1762
rect 14898 1678 14928 1762
rect 15024 1678 15054 1762
<< scpmoshvt >>
rect 9420 2057 9450 2257
rect 9610 2057 9640 2257
<< pmoshvt >>
rect 9888 2820 9918 2904
rect 9888 2682 9918 2766
rect 9888 2544 9918 2628
rect 9888 2406 9918 2490
rect 9888 2268 9918 2352
rect 9888 2130 9918 2214
rect 15673 1819 15703 1903
rect 15673 1681 15703 1765
rect 15765 1681 15795 1765
rect 15861 1681 15891 1765
<< ndiff >>
rect 9368 1925 9420 1937
rect 9368 1891 9376 1925
rect 9410 1891 9420 1925
rect 9368 1857 9420 1891
rect 9368 1823 9376 1857
rect 9410 1823 9420 1857
rect 9368 1807 9420 1823
rect 9450 1925 9502 1937
rect 9450 1891 9460 1925
rect 9494 1891 9502 1925
rect 9450 1857 9502 1891
rect 9450 1823 9460 1857
rect 9494 1823 9502 1857
rect 9450 1807 9502 1823
rect 9558 1925 9610 1937
rect 9558 1891 9566 1925
rect 9600 1891 9610 1925
rect 9558 1857 9610 1891
rect 9558 1823 9566 1857
rect 9600 1823 9610 1857
rect 9558 1807 9610 1823
rect 9640 1925 9692 1937
rect 9640 1891 9650 1925
rect 9684 1891 9692 1925
rect 9640 1857 9692 1891
rect 9640 1823 9650 1857
rect 9684 1823 9692 1857
rect 9640 1807 9692 1823
rect 10825 1549 10883 1561
rect 10825 1489 10837 1549
rect 10871 1489 10883 1549
rect 10825 1477 10883 1489
rect 10913 1549 10971 1561
rect 10913 1489 10927 1549
rect 10961 1489 10971 1549
rect 10913 1477 10971 1489
rect 11557 1549 11615 1561
rect 11557 1489 11569 1549
rect 11603 1489 11615 1549
rect 11557 1477 11615 1489
rect 11645 1549 11737 1561
rect 11645 1489 11676 1549
rect 11710 1489 11737 1549
rect 11645 1477 11737 1489
rect 11767 1549 11825 1561
rect 11767 1489 11779 1549
rect 11813 1489 11825 1549
rect 11767 1477 11825 1489
rect 12769 1549 12827 1561
rect 12769 1489 12781 1549
rect 12815 1489 12827 1549
rect 12769 1477 12827 1489
rect 12857 1549 12949 1561
rect 12857 1489 12887 1549
rect 12921 1489 12949 1549
rect 12857 1477 12949 1489
rect 12979 1549 13037 1561
rect 12979 1489 12991 1549
rect 13025 1489 13037 1549
rect 12979 1477 13037 1489
rect 14107 1549 14165 1561
rect 14107 1489 14119 1549
rect 14153 1489 14165 1549
rect 14107 1477 14165 1489
rect 14195 1549 14287 1561
rect 14195 1489 14227 1549
rect 14261 1489 14287 1549
rect 14195 1477 14287 1489
rect 14317 1549 14375 1561
rect 14317 1489 14329 1549
rect 14363 1489 14375 1549
rect 14317 1477 14375 1489
rect 14962 1549 15021 1561
rect 14962 1489 14974 1549
rect 15008 1489 15021 1549
rect 14962 1477 15021 1489
rect 15051 1549 15109 1561
rect 15051 1489 15063 1549
rect 15097 1489 15109 1549
rect 15051 1477 15109 1489
rect 15615 1550 15673 1562
rect 15615 1490 15627 1550
rect 15661 1490 15673 1550
rect 15615 1478 15673 1490
rect 15703 1550 15765 1562
rect 15703 1490 15715 1550
rect 15749 1490 15765 1550
rect 15703 1478 15765 1490
rect 15795 1550 15861 1562
rect 15795 1490 15811 1550
rect 15845 1490 15861 1550
rect 15795 1478 15861 1490
rect 15891 1550 15953 1562
rect 15891 1490 15907 1550
rect 15941 1490 15953 1550
rect 15891 1478 15953 1490
rect 15615 1412 15673 1424
rect 9805 1365 9863 1377
rect 9805 1305 9817 1365
rect 9851 1305 9863 1365
rect 9805 1293 9863 1305
rect 9893 1293 9935 1377
rect 9965 1365 10023 1377
rect 9965 1305 9977 1365
rect 10011 1305 10023 1365
rect 15615 1352 15627 1412
rect 15661 1352 15673 1412
rect 15615 1340 15673 1352
rect 15703 1412 15761 1424
rect 15703 1352 15715 1412
rect 15749 1352 15761 1412
rect 15703 1340 15761 1352
rect 9965 1293 10023 1305
rect 9805 1227 9863 1239
rect 9805 1167 9817 1227
rect 9851 1167 9863 1227
rect 9805 1155 9863 1167
rect 9893 1155 9935 1239
rect 9965 1227 10023 1239
rect 9965 1167 9977 1227
rect 10011 1167 10023 1227
rect 9965 1155 10023 1167
rect 9805 1089 9863 1101
rect 9805 1029 9817 1089
rect 9851 1029 9863 1089
rect 9805 1017 9863 1029
rect 9893 1017 9935 1101
rect 9965 1089 10023 1101
rect 9965 1029 9977 1089
rect 10011 1029 10023 1089
rect 9965 1017 10023 1029
rect 9805 951 9863 963
rect 9805 891 9817 951
rect 9851 891 9863 951
rect 9805 879 9863 891
rect 9893 879 9935 963
rect 9965 951 10023 963
rect 9965 891 9977 951
rect 10011 891 10023 951
rect 9965 879 10023 891
rect 9805 813 9863 825
rect 9805 753 9817 813
rect 9851 753 9863 813
rect 9805 741 9863 753
rect 9893 741 9935 825
rect 9965 813 10023 825
rect 9965 753 9977 813
rect 10011 753 10023 813
rect 9965 741 10023 753
rect 9805 675 9863 687
rect 9805 615 9817 675
rect 9851 615 9863 675
rect 9805 603 9863 615
rect 9893 603 9935 687
rect 9965 675 10023 687
rect 9965 615 9977 675
rect 10011 615 10023 675
rect 9965 603 10023 615
rect 9805 537 9863 549
rect 9805 477 9817 537
rect 9851 477 9863 537
rect 9805 465 9863 477
rect 9893 465 9935 549
rect 9965 537 10023 549
rect 9965 477 9977 537
rect 10011 477 10023 537
rect 9965 465 10023 477
rect 9805 399 9863 411
rect 9805 339 9817 399
rect 9851 339 9863 399
rect 9805 327 9863 339
rect 9893 327 9935 411
rect 9965 399 10023 411
rect 9965 339 9977 399
rect 10011 339 10023 399
rect 9965 327 10023 339
<< pdiff >>
rect 9830 2892 9888 2904
rect 9830 2832 9842 2892
rect 9876 2832 9888 2892
rect 9830 2820 9888 2832
rect 9918 2892 9976 2904
rect 9918 2832 9930 2892
rect 9964 2832 9976 2892
rect 9918 2820 9976 2832
rect 9830 2754 9888 2766
rect 9830 2694 9842 2754
rect 9876 2694 9888 2754
rect 9830 2682 9888 2694
rect 9918 2754 9976 2766
rect 9918 2694 9930 2754
rect 9964 2694 9976 2754
rect 9918 2682 9976 2694
rect 9830 2616 9888 2628
rect 9830 2556 9842 2616
rect 9876 2556 9888 2616
rect 9830 2544 9888 2556
rect 9918 2616 9976 2628
rect 9918 2556 9930 2616
rect 9964 2556 9976 2616
rect 9918 2544 9976 2556
rect 9830 2478 9888 2490
rect 9830 2418 9842 2478
rect 9876 2418 9888 2478
rect 9830 2406 9888 2418
rect 9918 2478 9976 2490
rect 9918 2418 9930 2478
rect 9964 2418 9976 2478
rect 9918 2406 9976 2418
rect 9830 2340 9888 2352
rect 9830 2280 9842 2340
rect 9876 2280 9888 2340
rect 9830 2268 9888 2280
rect 9918 2340 9976 2352
rect 9918 2280 9930 2340
rect 9964 2280 9976 2340
rect 9918 2268 9976 2280
rect 9368 2245 9420 2257
rect 9368 2211 9376 2245
rect 9410 2211 9420 2245
rect 9368 2177 9420 2211
rect 9368 2143 9376 2177
rect 9410 2143 9420 2177
rect 9368 2109 9420 2143
rect 9368 2075 9376 2109
rect 9410 2075 9420 2109
rect 9368 2057 9420 2075
rect 9450 2245 9502 2257
rect 9450 2211 9460 2245
rect 9494 2211 9502 2245
rect 9450 2177 9502 2211
rect 9450 2143 9460 2177
rect 9494 2143 9502 2177
rect 9450 2109 9502 2143
rect 9450 2075 9460 2109
rect 9494 2075 9502 2109
rect 9450 2057 9502 2075
rect 9558 2245 9610 2257
rect 9558 2211 9566 2245
rect 9600 2211 9610 2245
rect 9558 2177 9610 2211
rect 9558 2143 9566 2177
rect 9600 2143 9610 2177
rect 9558 2109 9610 2143
rect 9558 2075 9566 2109
rect 9600 2075 9610 2109
rect 9558 2057 9610 2075
rect 9640 2245 9692 2257
rect 9640 2211 9650 2245
rect 9684 2211 9692 2245
rect 9640 2177 9692 2211
rect 9640 2143 9650 2177
rect 9684 2143 9692 2177
rect 9640 2109 9692 2143
rect 9830 2202 9888 2214
rect 9830 2142 9842 2202
rect 9876 2142 9888 2202
rect 9830 2130 9888 2142
rect 9918 2202 9976 2214
rect 9918 2142 9930 2202
rect 9964 2142 9976 2202
rect 9918 2130 9976 2142
rect 9640 2075 9650 2109
rect 9684 2075 9692 2109
rect 9640 2057 9692 2075
rect 15615 1891 15673 1903
rect 15615 1831 15627 1891
rect 15661 1831 15673 1891
rect 15615 1819 15673 1831
rect 15703 1891 15761 1903
rect 15703 1831 15715 1891
rect 15749 1831 15761 1891
rect 15703 1819 15761 1831
rect 10472 1750 10530 1762
rect 10472 1690 10484 1750
rect 10518 1690 10530 1750
rect 10472 1678 10530 1690
rect 10560 1750 10618 1762
rect 10560 1690 10572 1750
rect 10606 1690 10618 1750
rect 10560 1678 10618 1690
rect 11204 1750 11262 1762
rect 11204 1690 11216 1750
rect 11250 1690 11262 1750
rect 11204 1678 11262 1690
rect 11292 1750 11388 1762
rect 11292 1690 11321 1750
rect 11355 1690 11388 1750
rect 11292 1678 11388 1690
rect 11418 1750 11476 1762
rect 11418 1690 11430 1750
rect 11464 1690 11476 1750
rect 11418 1678 11476 1690
rect 12416 1750 12474 1762
rect 12416 1690 12428 1750
rect 12462 1690 12474 1750
rect 12416 1678 12474 1690
rect 12504 1750 12600 1762
rect 12504 1690 12532 1750
rect 12566 1690 12600 1750
rect 12504 1678 12600 1690
rect 12630 1750 12688 1762
rect 12630 1690 12642 1750
rect 12676 1690 12688 1750
rect 12630 1678 12688 1690
rect 13628 1750 13686 1762
rect 13628 1690 13640 1750
rect 13674 1690 13686 1750
rect 13628 1678 13686 1690
rect 13716 1750 13812 1762
rect 13716 1690 13745 1750
rect 13779 1690 13812 1750
rect 13716 1678 13812 1690
rect 13842 1750 13900 1762
rect 13842 1690 13854 1750
rect 13888 1690 13900 1750
rect 13842 1678 13900 1690
rect 14840 1750 14898 1762
rect 14840 1690 14852 1750
rect 14886 1690 14898 1750
rect 14840 1678 14898 1690
rect 14928 1750 15024 1762
rect 14928 1690 14959 1750
rect 14993 1690 15024 1750
rect 14928 1678 15024 1690
rect 15054 1750 15112 1762
rect 15054 1690 15066 1750
rect 15100 1690 15112 1750
rect 15054 1678 15112 1690
rect 15615 1753 15673 1765
rect 15615 1693 15627 1753
rect 15661 1693 15673 1753
rect 15615 1681 15673 1693
rect 15703 1753 15765 1765
rect 15703 1693 15715 1753
rect 15749 1693 15765 1753
rect 15703 1681 15765 1693
rect 15795 1753 15861 1765
rect 15795 1693 15811 1753
rect 15845 1693 15861 1753
rect 15795 1681 15861 1693
rect 15891 1753 15953 1765
rect 15891 1693 15907 1753
rect 15941 1693 15953 1753
rect 15891 1681 15953 1693
<< ndiffc >>
rect 9376 1891 9410 1925
rect 9376 1823 9410 1857
rect 9460 1891 9494 1925
rect 9460 1823 9494 1857
rect 9566 1891 9600 1925
rect 9566 1823 9600 1857
rect 9650 1891 9684 1925
rect 9650 1823 9684 1857
rect 10837 1489 10871 1549
rect 10927 1489 10961 1549
rect 11569 1489 11603 1549
rect 11676 1489 11710 1549
rect 11779 1489 11813 1549
rect 12781 1489 12815 1549
rect 12887 1489 12921 1549
rect 12991 1489 13025 1549
rect 14119 1489 14153 1549
rect 14227 1489 14261 1549
rect 14329 1489 14363 1549
rect 14974 1489 15008 1549
rect 15063 1489 15097 1549
rect 15627 1490 15661 1550
rect 15715 1490 15749 1550
rect 15811 1490 15845 1550
rect 15907 1490 15941 1550
rect 9817 1305 9851 1365
rect 9977 1305 10011 1365
rect 15627 1352 15661 1412
rect 15715 1352 15749 1412
rect 9817 1167 9851 1227
rect 9977 1167 10011 1227
rect 9817 1029 9851 1089
rect 9977 1029 10011 1089
rect 9817 891 9851 951
rect 9977 891 10011 951
rect 9817 753 9851 813
rect 9977 753 10011 813
rect 9817 615 9851 675
rect 9977 615 10011 675
rect 9817 477 9851 537
rect 9977 477 10011 537
rect 9817 339 9851 399
rect 9977 339 10011 399
<< pdiffc >>
rect 9842 2832 9876 2892
rect 9930 2832 9964 2892
rect 9842 2694 9876 2754
rect 9930 2694 9964 2754
rect 9842 2556 9876 2616
rect 9930 2556 9964 2616
rect 9842 2418 9876 2478
rect 9930 2418 9964 2478
rect 9842 2280 9876 2340
rect 9930 2280 9964 2340
rect 9376 2211 9410 2245
rect 9376 2143 9410 2177
rect 9376 2075 9410 2109
rect 9460 2211 9494 2245
rect 9460 2143 9494 2177
rect 9460 2075 9494 2109
rect 9566 2211 9600 2245
rect 9566 2143 9600 2177
rect 9566 2075 9600 2109
rect 9650 2211 9684 2245
rect 9650 2143 9684 2177
rect 9842 2142 9876 2202
rect 9930 2142 9964 2202
rect 9650 2075 9684 2109
rect 15627 1831 15661 1891
rect 15715 1831 15749 1891
rect 10484 1690 10518 1750
rect 10572 1690 10606 1750
rect 11216 1690 11250 1750
rect 11321 1690 11355 1750
rect 11430 1690 11464 1750
rect 12428 1690 12462 1750
rect 12532 1690 12566 1750
rect 12642 1690 12676 1750
rect 13640 1690 13674 1750
rect 13745 1690 13779 1750
rect 13854 1690 13888 1750
rect 14852 1690 14886 1750
rect 14959 1690 14993 1750
rect 15066 1690 15100 1750
rect 15627 1693 15661 1753
rect 15715 1693 15749 1753
rect 15811 1693 15845 1753
rect 15907 1693 15941 1753
<< psubdiff >>
rect 9370 1714 9394 1748
rect 9428 1714 9512 1748
rect 9546 1714 9656 1748
rect 9690 1714 9732 1748
rect 9370 1712 9732 1714
rect 10492 352 10824 368
rect 10492 318 10518 352
rect 10552 318 10598 352
rect 10632 318 10678 352
rect 10712 318 10758 352
rect 10792 318 10824 352
rect 10492 300 10824 318
rect 11224 352 11556 368
rect 11224 318 11250 352
rect 11284 318 11330 352
rect 11364 318 11410 352
rect 11444 318 11490 352
rect 11524 318 11556 352
rect 11224 300 11556 318
rect 11826 352 12158 368
rect 11826 318 11858 352
rect 11892 318 11938 352
rect 11972 318 12018 352
rect 12052 318 12098 352
rect 12132 318 12158 352
rect 11826 300 12158 318
rect 12436 352 12768 368
rect 12436 318 12462 352
rect 12496 318 12542 352
rect 12576 318 12622 352
rect 12656 318 12702 352
rect 12736 318 12768 352
rect 12436 300 12768 318
rect 13038 352 13370 368
rect 13038 318 13070 352
rect 13104 318 13150 352
rect 13184 318 13230 352
rect 13264 318 13310 352
rect 13344 318 13370 352
rect 13038 300 13370 318
rect 13774 352 14106 368
rect 13774 318 13800 352
rect 13834 318 13880 352
rect 13914 318 13960 352
rect 13994 318 14040 352
rect 14074 318 14106 352
rect 13774 300 14106 318
rect 14376 352 14708 368
rect 14376 318 14408 352
rect 14442 318 14488 352
rect 14522 318 14568 352
rect 14602 318 14648 352
rect 14682 318 14708 352
rect 14376 300 14708 318
rect 15110 352 15442 368
rect 15110 318 15142 352
rect 15176 318 15222 352
rect 15256 318 15302 352
rect 15336 318 15382 352
rect 15416 318 15442 352
rect 15110 300 15442 318
<< nsubdiff >>
rect 10040 2919 10578 2939
rect 10040 2885 10088 2919
rect 10122 2885 10168 2919
rect 10202 2885 10248 2919
rect 10282 2885 10328 2919
rect 10362 2885 10408 2919
rect 10442 2885 10488 2919
rect 10522 2885 10578 2919
rect 10040 2871 10578 2885
rect 10772 2919 11310 2939
rect 10772 2885 10820 2919
rect 10854 2885 10900 2919
rect 10934 2885 10980 2919
rect 11014 2885 11060 2919
rect 11094 2885 11140 2919
rect 11174 2885 11220 2919
rect 11254 2885 11310 2919
rect 10772 2871 11310 2885
rect 11370 2919 11908 2939
rect 11370 2885 11426 2919
rect 11460 2885 11506 2919
rect 11540 2885 11586 2919
rect 11620 2885 11666 2919
rect 11700 2885 11746 2919
rect 11780 2885 11826 2919
rect 11860 2885 11908 2919
rect 11370 2871 11908 2885
rect 11984 2919 12522 2939
rect 11984 2885 12032 2919
rect 12066 2885 12112 2919
rect 12146 2885 12192 2919
rect 12226 2885 12272 2919
rect 12306 2885 12352 2919
rect 12386 2885 12432 2919
rect 12466 2885 12522 2919
rect 11984 2871 12522 2885
rect 12582 2919 13120 2939
rect 12582 2885 12638 2919
rect 12672 2885 12718 2919
rect 12752 2885 12798 2919
rect 12832 2885 12878 2919
rect 12912 2885 12958 2919
rect 12992 2885 13038 2919
rect 13072 2885 13120 2919
rect 12582 2871 13120 2885
rect 13196 2919 13734 2939
rect 13196 2885 13244 2919
rect 13278 2885 13324 2919
rect 13358 2885 13404 2919
rect 13438 2885 13484 2919
rect 13518 2885 13564 2919
rect 13598 2885 13644 2919
rect 13678 2885 13734 2919
rect 13196 2871 13734 2885
rect 13794 2919 14332 2939
rect 13794 2885 13850 2919
rect 13884 2885 13930 2919
rect 13964 2885 14010 2919
rect 14044 2885 14090 2919
rect 14124 2885 14170 2919
rect 14204 2885 14250 2919
rect 14284 2885 14332 2919
rect 13794 2871 14332 2885
rect 14408 2919 14946 2939
rect 14408 2885 14456 2919
rect 14490 2885 14536 2919
rect 14570 2885 14616 2919
rect 14650 2885 14696 2919
rect 14730 2885 14776 2919
rect 14810 2885 14856 2919
rect 14890 2885 14946 2919
rect 14408 2871 14946 2885
rect 15006 2919 15544 2939
rect 15006 2885 15062 2919
rect 15096 2885 15142 2919
rect 15176 2885 15222 2919
rect 15256 2885 15302 2919
rect 15336 2885 15382 2919
rect 15416 2885 15462 2919
rect 15496 2885 15544 2919
rect 15006 2871 15544 2885
rect 15776 2868 15862 2894
rect 15776 2834 15802 2868
rect 15836 2834 15862 2868
rect 15776 2808 15862 2834
rect 15781 2724 15867 2750
rect 15781 2690 15807 2724
rect 15841 2690 15867 2724
rect 15781 2664 15867 2690
rect 15782 2572 15868 2598
rect 15782 2538 15808 2572
rect 15842 2538 15868 2572
rect 15782 2512 15868 2538
rect 15782 2402 15868 2428
rect 15782 2368 15808 2402
rect 15842 2368 15868 2402
rect 9344 2350 9760 2352
rect 9344 2316 9374 2350
rect 9408 2316 9504 2350
rect 9538 2316 9650 2350
rect 9684 2316 9760 2350
rect 9344 2312 9760 2316
rect 15782 2342 15868 2368
rect 15781 2245 15867 2271
rect 15781 2211 15807 2245
rect 15841 2211 15867 2245
rect 15781 2185 15867 2211
<< psubdiffcont >>
rect 9394 1714 9428 1748
rect 9512 1714 9546 1748
rect 9656 1714 9690 1748
rect 10518 318 10552 352
rect 10598 318 10632 352
rect 10678 318 10712 352
rect 10758 318 10792 352
rect 11250 318 11284 352
rect 11330 318 11364 352
rect 11410 318 11444 352
rect 11490 318 11524 352
rect 11858 318 11892 352
rect 11938 318 11972 352
rect 12018 318 12052 352
rect 12098 318 12132 352
rect 12462 318 12496 352
rect 12542 318 12576 352
rect 12622 318 12656 352
rect 12702 318 12736 352
rect 13070 318 13104 352
rect 13150 318 13184 352
rect 13230 318 13264 352
rect 13310 318 13344 352
rect 13800 318 13834 352
rect 13880 318 13914 352
rect 13960 318 13994 352
rect 14040 318 14074 352
rect 14408 318 14442 352
rect 14488 318 14522 352
rect 14568 318 14602 352
rect 14648 318 14682 352
rect 15142 318 15176 352
rect 15222 318 15256 352
rect 15302 318 15336 352
rect 15382 318 15416 352
<< nsubdiffcont >>
rect 10088 2885 10122 2919
rect 10168 2885 10202 2919
rect 10248 2885 10282 2919
rect 10328 2885 10362 2919
rect 10408 2885 10442 2919
rect 10488 2885 10522 2919
rect 10820 2885 10854 2919
rect 10900 2885 10934 2919
rect 10980 2885 11014 2919
rect 11060 2885 11094 2919
rect 11140 2885 11174 2919
rect 11220 2885 11254 2919
rect 11426 2885 11460 2919
rect 11506 2885 11540 2919
rect 11586 2885 11620 2919
rect 11666 2885 11700 2919
rect 11746 2885 11780 2919
rect 11826 2885 11860 2919
rect 12032 2885 12066 2919
rect 12112 2885 12146 2919
rect 12192 2885 12226 2919
rect 12272 2885 12306 2919
rect 12352 2885 12386 2919
rect 12432 2885 12466 2919
rect 12638 2885 12672 2919
rect 12718 2885 12752 2919
rect 12798 2885 12832 2919
rect 12878 2885 12912 2919
rect 12958 2885 12992 2919
rect 13038 2885 13072 2919
rect 13244 2885 13278 2919
rect 13324 2885 13358 2919
rect 13404 2885 13438 2919
rect 13484 2885 13518 2919
rect 13564 2885 13598 2919
rect 13644 2885 13678 2919
rect 13850 2885 13884 2919
rect 13930 2885 13964 2919
rect 14010 2885 14044 2919
rect 14090 2885 14124 2919
rect 14170 2885 14204 2919
rect 14250 2885 14284 2919
rect 14456 2885 14490 2919
rect 14536 2885 14570 2919
rect 14616 2885 14650 2919
rect 14696 2885 14730 2919
rect 14776 2885 14810 2919
rect 14856 2885 14890 2919
rect 15062 2885 15096 2919
rect 15142 2885 15176 2919
rect 15222 2885 15256 2919
rect 15302 2885 15336 2919
rect 15382 2885 15416 2919
rect 15462 2885 15496 2919
rect 15802 2834 15836 2868
rect 15807 2690 15841 2724
rect 15808 2538 15842 2572
rect 15808 2368 15842 2402
rect 9374 2316 9408 2350
rect 9504 2316 9538 2350
rect 9650 2316 9684 2350
rect 15807 2211 15841 2245
<< poly >>
rect 9888 2904 9918 2934
rect 9888 2766 9918 2820
rect 9888 2628 9918 2682
rect 9888 2490 9918 2544
rect 9888 2352 9918 2406
rect 9420 2257 9450 2283
rect 9610 2257 9640 2283
rect 9888 2214 9918 2268
rect 9888 2099 9918 2130
rect 9870 2083 9936 2099
rect 9420 2025 9450 2057
rect 9364 2009 9450 2025
rect 9364 1975 9380 2009
rect 9414 1975 9450 2009
rect 9364 1959 9450 1975
rect 9420 1937 9450 1959
rect 9610 2025 9640 2057
rect 9870 2049 9886 2083
rect 9920 2049 9936 2083
rect 9870 2033 9936 2049
rect 9610 2009 9696 2025
rect 9610 1975 9646 2009
rect 9680 1975 9696 2009
rect 9610 1959 9696 1975
rect 9610 1937 9640 1959
rect 15673 1903 15703 1934
rect 10512 1843 10578 1859
rect 10512 1809 10528 1843
rect 10562 1809 10578 1843
rect 9420 1781 9450 1807
rect 9610 1781 9640 1807
rect 10512 1793 10578 1809
rect 11244 1843 11310 1859
rect 11244 1809 11260 1843
rect 11294 1809 11310 1843
rect 11244 1793 11310 1809
rect 11370 1843 11436 1859
rect 11370 1809 11386 1843
rect 11420 1809 11436 1843
rect 11370 1793 11436 1809
rect 12456 1843 12522 1859
rect 12456 1809 12472 1843
rect 12506 1809 12522 1843
rect 12456 1793 12522 1809
rect 12582 1843 12648 1859
rect 12582 1809 12598 1843
rect 12632 1809 12648 1843
rect 12582 1793 12648 1809
rect 13668 1843 13734 1859
rect 13668 1809 13684 1843
rect 13718 1809 13734 1843
rect 13668 1793 13734 1809
rect 13794 1843 13860 1859
rect 13794 1809 13810 1843
rect 13844 1809 13860 1843
rect 13794 1793 13860 1809
rect 14880 1843 14946 1859
rect 14880 1809 14896 1843
rect 14930 1809 14946 1843
rect 14880 1793 14946 1809
rect 15006 1843 15072 1859
rect 15006 1809 15022 1843
rect 15056 1809 15072 1843
rect 15006 1793 15072 1809
rect 10530 1762 10560 1793
rect 11262 1762 11292 1793
rect 11388 1762 11418 1793
rect 12474 1762 12504 1793
rect 12600 1762 12630 1793
rect 13686 1762 13716 1793
rect 13812 1762 13842 1793
rect 14898 1762 14928 1793
rect 15024 1762 15054 1793
rect 15673 1765 15703 1819
rect 15765 1765 15795 1791
rect 15861 1765 15891 1796
rect 10530 1650 10560 1678
rect 11262 1650 11292 1678
rect 11388 1650 11418 1678
rect 12474 1650 12504 1678
rect 12600 1650 12630 1678
rect 13686 1650 13716 1678
rect 13812 1650 13842 1678
rect 14898 1650 14928 1678
rect 15024 1650 15054 1678
rect 15673 1656 15703 1681
rect 15544 1636 15703 1656
rect 15765 1656 15795 1681
rect 15861 1656 15891 1681
rect 15765 1650 15891 1656
rect 15544 1602 15556 1636
rect 15590 1602 15703 1636
rect 10883 1561 10913 1587
rect 11615 1561 11645 1587
rect 11737 1561 11767 1587
rect 12827 1561 12857 1587
rect 12949 1561 12979 1587
rect 14165 1561 14195 1587
rect 14287 1561 14317 1587
rect 15021 1561 15051 1587
rect 15544 1583 15703 1602
rect 15747 1634 15891 1650
rect 15747 1600 15763 1634
rect 15797 1600 15891 1634
rect 15747 1584 15891 1600
rect 15673 1562 15703 1583
rect 15765 1577 15891 1584
rect 15765 1562 15795 1577
rect 15861 1562 15891 1577
rect 9881 1449 9947 1465
rect 10883 1455 10913 1477
rect 11615 1455 11645 1477
rect 11737 1455 11767 1477
rect 12827 1455 12857 1477
rect 12949 1455 12979 1477
rect 14165 1455 14195 1477
rect 14287 1455 14317 1477
rect 15021 1455 15051 1477
rect 9881 1422 9897 1449
rect 9863 1415 9897 1422
rect 9931 1422 9947 1449
rect 10865 1439 10931 1455
rect 9931 1415 9965 1422
rect 9863 1392 9965 1415
rect 9863 1377 9893 1392
rect 9935 1377 9965 1392
rect 10865 1405 10881 1439
rect 10915 1405 10931 1439
rect 10865 1389 10931 1405
rect 11597 1439 11663 1455
rect 11597 1405 11613 1439
rect 11647 1405 11663 1439
rect 11597 1389 11663 1405
rect 11719 1439 11785 1455
rect 11719 1405 11735 1439
rect 11769 1405 11785 1439
rect 11719 1389 11785 1405
rect 12809 1439 12875 1455
rect 12809 1405 12825 1439
rect 12859 1405 12875 1439
rect 12809 1389 12875 1405
rect 12931 1439 12997 1455
rect 12931 1405 12947 1439
rect 12981 1405 12997 1439
rect 12931 1389 12997 1405
rect 14147 1439 14213 1455
rect 14147 1405 14163 1439
rect 14197 1405 14213 1439
rect 14147 1389 14213 1405
rect 14269 1439 14335 1455
rect 14269 1405 14285 1439
rect 14319 1405 14335 1439
rect 14269 1389 14335 1405
rect 15003 1439 15069 1455
rect 15003 1405 15019 1439
rect 15053 1405 15069 1439
rect 15673 1424 15703 1478
rect 15765 1452 15795 1478
rect 15861 1452 15891 1478
rect 15003 1389 15069 1405
rect 15673 1313 15703 1340
rect 9863 1239 9893 1293
rect 9935 1239 9965 1293
rect 9863 1101 9893 1155
rect 9935 1101 9965 1155
rect 9863 963 9893 1017
rect 9935 963 9965 1017
rect 9863 825 9893 879
rect 9935 825 9965 879
rect 9863 687 9893 741
rect 9935 687 9965 741
rect 9863 549 9893 603
rect 9935 549 9965 603
rect 9863 411 9893 465
rect 9935 411 9965 465
rect 9863 301 9893 327
rect 9935 301 9965 327
<< polycont >>
rect 9380 1975 9414 2009
rect 9886 2049 9920 2083
rect 9646 1975 9680 2009
rect 10528 1809 10562 1843
rect 11260 1809 11294 1843
rect 11386 1809 11420 1843
rect 12472 1809 12506 1843
rect 12598 1809 12632 1843
rect 13684 1809 13718 1843
rect 13810 1809 13844 1843
rect 14896 1809 14930 1843
rect 15022 1809 15056 1843
rect 15556 1602 15590 1636
rect 15763 1600 15797 1634
rect 9897 1415 9931 1449
rect 10881 1405 10915 1439
rect 11613 1405 11647 1439
rect 11735 1405 11769 1439
rect 12825 1405 12859 1439
rect 12947 1405 12981 1439
rect 14163 1405 14197 1439
rect 14285 1405 14319 1439
rect 15019 1405 15053 1439
<< locali >>
rect 9972 2919 10642 2937
rect 9972 2908 10088 2919
rect 9842 2892 9876 2908
rect 9842 2816 9876 2832
rect 9930 2892 10088 2908
rect 9964 2885 10088 2892
rect 10124 2885 10168 2919
rect 10204 2885 10248 2919
rect 10284 2885 10328 2919
rect 10364 2885 10408 2919
rect 10444 2885 10488 2919
rect 10524 2885 10642 2919
rect 9964 2871 10642 2885
rect 10704 2919 15612 2937
rect 10704 2885 10820 2919
rect 10856 2885 10900 2919
rect 10936 2885 10980 2919
rect 11016 2885 11060 2919
rect 11096 2885 11140 2919
rect 11176 2885 11220 2919
rect 11256 2885 11424 2919
rect 11460 2885 11504 2919
rect 11540 2885 11584 2919
rect 11620 2885 11664 2919
rect 11700 2885 11744 2919
rect 11780 2885 11824 2919
rect 11860 2885 12032 2919
rect 12068 2885 12112 2919
rect 12148 2885 12192 2919
rect 12228 2885 12272 2919
rect 12308 2885 12352 2919
rect 12388 2885 12432 2919
rect 12468 2885 12636 2919
rect 12672 2885 12716 2919
rect 12752 2885 12796 2919
rect 12832 2885 12876 2919
rect 12912 2885 12956 2919
rect 12992 2885 13036 2919
rect 13072 2885 13244 2919
rect 13280 2885 13324 2919
rect 13360 2885 13404 2919
rect 13440 2885 13484 2919
rect 13520 2885 13564 2919
rect 13600 2885 13644 2919
rect 13680 2885 13848 2919
rect 13884 2885 13928 2919
rect 13964 2885 14008 2919
rect 14044 2885 14088 2919
rect 14124 2885 14168 2919
rect 14204 2885 14248 2919
rect 14284 2885 14456 2919
rect 14492 2885 14536 2919
rect 14572 2885 14616 2919
rect 14652 2885 14696 2919
rect 14732 2885 14776 2919
rect 14812 2885 14856 2919
rect 14892 2885 15060 2919
rect 15096 2885 15140 2919
rect 15176 2885 15220 2919
rect 15256 2885 15300 2919
rect 15336 2885 15380 2919
rect 15416 2885 15460 2919
rect 15496 2885 15612 2919
rect 10704 2871 15612 2885
rect 9930 2816 9964 2832
rect 15776 2868 15862 2894
rect 15776 2834 15802 2868
rect 15836 2834 15862 2868
rect 15776 2808 15862 2834
rect 9842 2754 9876 2770
rect 9842 2678 9876 2694
rect 9930 2754 9964 2770
rect 9930 2678 9964 2694
rect 15781 2724 15867 2750
rect 15781 2690 15807 2724
rect 15841 2690 15867 2724
rect 15781 2664 15867 2690
rect 9842 2616 9876 2632
rect 9842 2540 9876 2556
rect 9930 2616 9964 2632
rect 9930 2540 9964 2556
rect 15782 2572 15868 2598
rect 15782 2538 15808 2572
rect 15842 2538 15868 2572
rect 15782 2512 15868 2538
rect 9842 2478 9876 2494
rect 9842 2402 9876 2418
rect 9930 2478 9964 2494
rect 9930 2402 9964 2418
rect 15782 2402 15868 2428
rect 15782 2368 15808 2402
rect 15842 2368 15868 2402
rect 9358 2321 9374 2350
rect 9300 2287 9329 2321
rect 9363 2316 9374 2321
rect 9408 2321 9424 2350
rect 9488 2321 9504 2350
rect 9538 2321 9558 2350
rect 9634 2321 9650 2350
rect 9408 2316 9421 2321
rect 9363 2287 9421 2316
rect 9455 2316 9504 2321
rect 9455 2287 9513 2316
rect 9547 2287 9605 2321
rect 9639 2316 9650 2321
rect 9684 2321 9704 2350
rect 9842 2340 9876 2356
rect 9684 2316 9697 2321
rect 9639 2287 9697 2316
rect 9731 2287 9760 2321
rect 9368 2245 9410 2287
rect 9368 2211 9376 2245
rect 9368 2177 9410 2211
rect 9368 2143 9376 2177
rect 9368 2109 9410 2143
rect 9368 2075 9376 2109
rect 9368 2059 9410 2075
rect 9444 2245 9510 2253
rect 9444 2211 9460 2245
rect 9494 2211 9510 2245
rect 9444 2178 9510 2211
rect 9444 2144 9457 2178
rect 9491 2177 9510 2178
rect 9444 2143 9460 2144
rect 9494 2143 9510 2177
rect 9444 2109 9510 2143
rect 9444 2075 9460 2109
rect 9494 2075 9510 2109
rect 9444 2057 9510 2075
rect 9364 2013 9430 2023
rect 9364 1979 9376 2013
rect 9410 2009 9430 2013
rect 9364 1975 9380 1979
rect 9414 1975 9430 2009
rect 9364 1925 9410 1941
rect 9464 1937 9510 2057
rect 9364 1891 9376 1925
rect 9364 1857 9410 1891
rect 9364 1823 9376 1857
rect 9364 1777 9410 1823
rect 9444 1925 9510 1937
rect 9444 1891 9460 1925
rect 9494 1891 9510 1925
rect 9444 1857 9510 1891
rect 9444 1823 9460 1857
rect 9494 1823 9510 1857
rect 9444 1811 9510 1823
rect 9550 2245 9616 2253
rect 9550 2211 9566 2245
rect 9600 2211 9616 2245
rect 9550 2177 9616 2211
rect 9550 2143 9566 2177
rect 9600 2143 9616 2177
rect 9550 2123 9616 2143
rect 9550 2075 9566 2123
rect 9600 2075 9616 2123
rect 9550 2057 9616 2075
rect 9650 2245 9692 2287
rect 9842 2264 9876 2280
rect 9930 2340 9964 2356
rect 15782 2342 15868 2368
rect 9930 2264 9964 2280
rect 9684 2211 9692 2245
rect 15781 2245 15867 2271
rect 9650 2177 9692 2211
rect 9684 2143 9692 2177
rect 9650 2109 9692 2143
rect 9842 2202 9876 2218
rect 9842 2126 9876 2142
rect 9930 2202 9964 2218
rect 15781 2211 15807 2245
rect 15841 2211 15867 2245
rect 15781 2185 15867 2211
rect 9930 2126 9964 2142
rect 9684 2075 9692 2109
rect 9650 2059 9692 2075
rect 9550 1937 9596 2057
rect 9870 2049 9886 2083
rect 9920 2049 9936 2083
rect 9630 2012 9696 2023
rect 9630 2009 9650 2012
rect 9630 1975 9646 2009
rect 9684 1978 9696 2012
rect 9680 1975 9696 1978
rect 9780 2013 9829 2025
rect 9780 1979 9789 2013
rect 9823 2008 9829 2013
rect 9823 1979 10112 2008
rect 9780 1973 10112 1979
rect 9780 1966 9829 1973
rect 10077 1950 10112 1973
rect 9550 1925 9616 1937
rect 9550 1891 9566 1925
rect 9600 1891 9616 1925
rect 9550 1857 9616 1891
rect 9550 1823 9566 1857
rect 9600 1823 9616 1857
rect 9550 1811 9616 1823
rect 9650 1925 9696 1941
rect 10077 1938 10126 1950
rect 9684 1891 9696 1925
rect 9650 1857 9696 1891
rect 9818 1920 9867 1932
rect 9818 1886 9827 1920
rect 9861 1886 10028 1920
rect 10077 1904 10086 1938
rect 10120 1904 10126 1938
rect 10077 1891 10126 1904
rect 15627 1891 15661 1907
rect 9818 1873 9867 1886
rect 9684 1823 9696 1857
rect 9650 1777 9696 1823
rect 9987 1844 10028 1886
rect 10078 1845 10127 1857
rect 10078 1844 10087 1845
rect 9987 1811 10087 1844
rect 10121 1811 10127 1845
rect 9987 1810 10127 1811
rect 10078 1798 10127 1810
rect 10512 1809 10528 1843
rect 10562 1809 10578 1843
rect 11244 1809 11260 1843
rect 11294 1809 11310 1843
rect 11370 1809 11386 1843
rect 11420 1809 11436 1843
rect 12456 1809 12472 1843
rect 12506 1809 12522 1843
rect 12582 1809 12598 1843
rect 12632 1809 12648 1843
rect 13668 1809 13684 1843
rect 13718 1809 13734 1843
rect 13794 1809 13810 1843
rect 13844 1809 13860 1843
rect 14880 1809 14896 1843
rect 14930 1809 14946 1843
rect 15006 1809 15022 1843
rect 15056 1809 15072 1843
rect 15627 1815 15661 1831
rect 15715 1891 15749 1907
rect 15715 1815 15749 1831
rect 9300 1743 9329 1777
rect 9363 1748 9421 1777
rect 9455 1748 9513 1777
rect 9363 1743 9394 1748
rect 9455 1743 9512 1748
rect 9547 1743 9605 1777
rect 9639 1748 9697 1777
rect 9639 1743 9656 1748
rect 9378 1714 9394 1743
rect 9428 1714 9454 1743
rect 9496 1714 9512 1743
rect 9546 1714 9572 1743
rect 9638 1714 9656 1743
rect 9690 1743 9697 1748
rect 9731 1743 9760 1777
rect 10484 1750 10518 1766
rect 9690 1714 9706 1743
rect 10484 1674 10518 1690
rect 10572 1750 10606 1766
rect 10572 1674 10606 1690
rect 11216 1750 11250 1766
rect 11216 1674 11250 1690
rect 11321 1750 11355 1766
rect 11321 1674 11355 1690
rect 11430 1750 11464 1766
rect 11430 1674 11464 1690
rect 12428 1750 12462 1766
rect 12428 1674 12462 1690
rect 12532 1750 12566 1766
rect 12532 1674 12566 1690
rect 12642 1750 12676 1766
rect 12642 1674 12676 1690
rect 13640 1750 13674 1766
rect 13640 1674 13674 1690
rect 13745 1750 13779 1766
rect 13745 1674 13779 1690
rect 13854 1750 13888 1766
rect 13854 1674 13888 1690
rect 14852 1750 14886 1766
rect 14852 1674 14886 1690
rect 14959 1750 14993 1766
rect 14959 1674 14993 1690
rect 15066 1750 15100 1766
rect 15066 1674 15100 1690
rect 15627 1753 15661 1769
rect 15627 1677 15661 1693
rect 15715 1753 15749 1769
rect 15715 1677 15749 1693
rect 15811 1753 15845 1769
rect 15811 1677 15845 1693
rect 15907 1753 15941 1769
rect 15907 1677 15941 1693
rect 15540 1602 15556 1636
rect 15590 1602 15606 1636
rect 15747 1600 15763 1634
rect 15797 1600 15813 1634
rect 10837 1549 10871 1565
rect 10837 1473 10871 1489
rect 10927 1549 10961 1565
rect 10927 1473 10961 1489
rect 11569 1549 11603 1565
rect 11569 1473 11603 1489
rect 11676 1549 11710 1565
rect 11676 1473 11710 1489
rect 11779 1549 11813 1565
rect 11779 1473 11813 1489
rect 12781 1549 12815 1565
rect 12781 1473 12815 1489
rect 12887 1549 12921 1565
rect 12887 1473 12921 1489
rect 12991 1549 13025 1565
rect 12991 1473 13025 1489
rect 14119 1549 14153 1565
rect 14119 1473 14153 1489
rect 14227 1549 14261 1565
rect 14227 1473 14261 1489
rect 14329 1549 14363 1565
rect 14329 1473 14363 1489
rect 14974 1549 15008 1565
rect 14974 1473 15008 1489
rect 15063 1549 15097 1565
rect 15063 1473 15097 1489
rect 15627 1550 15661 1566
rect 15627 1474 15661 1490
rect 15715 1550 15749 1566
rect 15715 1474 15749 1490
rect 15811 1550 15845 1566
rect 15811 1474 15845 1490
rect 15907 1550 15941 1566
rect 15907 1474 15941 1490
rect 9881 1415 9897 1449
rect 9931 1415 9947 1449
rect 10865 1405 10881 1439
rect 10915 1405 10931 1439
rect 11597 1405 11613 1439
rect 11647 1405 11663 1439
rect 11719 1405 11735 1439
rect 11769 1405 11785 1439
rect 12809 1405 12825 1439
rect 12859 1405 12875 1439
rect 12931 1405 12947 1439
rect 12981 1405 12997 1439
rect 14147 1405 14163 1439
rect 14197 1405 14213 1439
rect 14269 1405 14285 1439
rect 14319 1405 14335 1439
rect 15003 1405 15019 1439
rect 15053 1405 15069 1439
rect 15627 1412 15661 1428
rect 9817 1365 9851 1381
rect 9817 1289 9851 1305
rect 9977 1365 10011 1381
rect 15627 1336 15661 1352
rect 15715 1412 15749 1428
rect 15715 1336 15749 1352
rect 9977 1289 10011 1305
rect 9817 1227 9851 1243
rect 9817 1151 9851 1167
rect 9977 1227 10011 1243
rect 9977 1151 10011 1167
rect 9817 1089 9851 1105
rect 9817 1013 9851 1029
rect 9977 1089 10011 1105
rect 9977 1013 10011 1029
rect 9817 951 9851 967
rect 9817 875 9851 891
rect 9977 951 10011 967
rect 9977 875 10011 891
rect 9817 813 9851 829
rect 9817 737 9851 753
rect 9977 813 10011 829
rect 9977 737 10011 753
rect 9817 675 9851 691
rect 9817 599 9851 615
rect 9977 675 10011 691
rect 9977 599 10011 615
rect 9817 537 9851 553
rect 9817 461 9851 477
rect 9977 537 10011 553
rect 9977 461 10011 477
rect 9817 399 9851 415
rect 9817 323 9851 339
rect 9977 399 10011 415
rect 9977 323 10011 339
rect 10492 352 10824 368
rect 10492 318 10518 352
rect 10552 318 10598 352
rect 10632 318 10678 352
rect 10712 318 10758 352
rect 10792 318 10824 352
rect 10492 300 10824 318
rect 11224 352 11556 368
rect 11224 318 11250 352
rect 11284 318 11330 352
rect 11364 318 11410 352
rect 11444 318 11490 352
rect 11524 318 11556 352
rect 11224 300 11556 318
rect 11826 352 12158 368
rect 11826 318 11858 352
rect 11892 318 11938 352
rect 11972 318 12018 352
rect 12052 318 12098 352
rect 12132 318 12158 352
rect 11826 300 12158 318
rect 12436 352 12768 368
rect 12436 318 12462 352
rect 12496 318 12542 352
rect 12576 318 12622 352
rect 12656 318 12702 352
rect 12736 318 12768 352
rect 12436 300 12768 318
rect 13038 352 13370 368
rect 13038 318 13070 352
rect 13104 318 13150 352
rect 13184 318 13230 352
rect 13264 318 13310 352
rect 13344 318 13370 352
rect 13038 300 13370 318
rect 13774 352 14106 368
rect 13774 318 13800 352
rect 13834 318 13880 352
rect 13914 318 13960 352
rect 13994 318 14040 352
rect 14074 318 14106 352
rect 13774 300 14106 318
rect 14376 352 14708 368
rect 14376 318 14408 352
rect 14442 318 14488 352
rect 14522 318 14568 352
rect 14602 318 14648 352
rect 14682 318 14708 352
rect 14376 300 14708 318
rect 15110 352 15442 368
rect 15110 318 15142 352
rect 15176 318 15222 352
rect 15256 318 15302 352
rect 15336 318 15382 352
rect 15416 318 15442 352
rect 15110 300 15442 318
<< viali >>
rect 9842 2832 9876 2892
rect 9930 2832 9964 2892
rect 10090 2885 10122 2919
rect 10122 2885 10124 2919
rect 10170 2885 10202 2919
rect 10202 2885 10204 2919
rect 10250 2885 10282 2919
rect 10282 2885 10284 2919
rect 10330 2885 10362 2919
rect 10362 2885 10364 2919
rect 10410 2885 10442 2919
rect 10442 2885 10444 2919
rect 10490 2885 10522 2919
rect 10522 2885 10524 2919
rect 10822 2885 10854 2919
rect 10854 2885 10856 2919
rect 10902 2885 10934 2919
rect 10934 2885 10936 2919
rect 10982 2885 11014 2919
rect 11014 2885 11016 2919
rect 11062 2885 11094 2919
rect 11094 2885 11096 2919
rect 11142 2885 11174 2919
rect 11174 2885 11176 2919
rect 11222 2885 11254 2919
rect 11254 2885 11256 2919
rect 11424 2885 11426 2919
rect 11426 2885 11458 2919
rect 11504 2885 11506 2919
rect 11506 2885 11538 2919
rect 11584 2885 11586 2919
rect 11586 2885 11618 2919
rect 11664 2885 11666 2919
rect 11666 2885 11698 2919
rect 11744 2885 11746 2919
rect 11746 2885 11778 2919
rect 11824 2885 11826 2919
rect 11826 2885 11858 2919
rect 12034 2885 12066 2919
rect 12066 2885 12068 2919
rect 12114 2885 12146 2919
rect 12146 2885 12148 2919
rect 12194 2885 12226 2919
rect 12226 2885 12228 2919
rect 12274 2885 12306 2919
rect 12306 2885 12308 2919
rect 12354 2885 12386 2919
rect 12386 2885 12388 2919
rect 12434 2885 12466 2919
rect 12466 2885 12468 2919
rect 12636 2885 12638 2919
rect 12638 2885 12670 2919
rect 12716 2885 12718 2919
rect 12718 2885 12750 2919
rect 12796 2885 12798 2919
rect 12798 2885 12830 2919
rect 12876 2885 12878 2919
rect 12878 2885 12910 2919
rect 12956 2885 12958 2919
rect 12958 2885 12990 2919
rect 13036 2885 13038 2919
rect 13038 2885 13070 2919
rect 13246 2885 13278 2919
rect 13278 2885 13280 2919
rect 13326 2885 13358 2919
rect 13358 2885 13360 2919
rect 13406 2885 13438 2919
rect 13438 2885 13440 2919
rect 13486 2885 13518 2919
rect 13518 2885 13520 2919
rect 13566 2885 13598 2919
rect 13598 2885 13600 2919
rect 13646 2885 13678 2919
rect 13678 2885 13680 2919
rect 13848 2885 13850 2919
rect 13850 2885 13882 2919
rect 13928 2885 13930 2919
rect 13930 2885 13962 2919
rect 14008 2885 14010 2919
rect 14010 2885 14042 2919
rect 14088 2885 14090 2919
rect 14090 2885 14122 2919
rect 14168 2885 14170 2919
rect 14170 2885 14202 2919
rect 14248 2885 14250 2919
rect 14250 2885 14282 2919
rect 14458 2885 14490 2919
rect 14490 2885 14492 2919
rect 14538 2885 14570 2919
rect 14570 2885 14572 2919
rect 14618 2885 14650 2919
rect 14650 2885 14652 2919
rect 14698 2885 14730 2919
rect 14730 2885 14732 2919
rect 14778 2885 14810 2919
rect 14810 2885 14812 2919
rect 14858 2885 14890 2919
rect 14890 2885 14892 2919
rect 15060 2885 15062 2919
rect 15062 2885 15094 2919
rect 15140 2885 15142 2919
rect 15142 2885 15174 2919
rect 15220 2885 15222 2919
rect 15222 2885 15254 2919
rect 15300 2885 15302 2919
rect 15302 2885 15334 2919
rect 15380 2885 15382 2919
rect 15382 2885 15414 2919
rect 15460 2885 15462 2919
rect 15462 2885 15494 2919
rect 15802 2834 15836 2868
rect 9842 2694 9876 2754
rect 9930 2694 9964 2754
rect 15807 2690 15841 2724
rect 9842 2556 9876 2616
rect 9930 2556 9964 2616
rect 15808 2538 15842 2572
rect 9842 2418 9876 2478
rect 9930 2418 9964 2478
rect 15808 2368 15842 2402
rect 9329 2287 9363 2321
rect 9421 2287 9455 2321
rect 9513 2316 9538 2321
rect 9538 2316 9547 2321
rect 9513 2287 9547 2316
rect 9605 2287 9639 2321
rect 9697 2287 9731 2321
rect 9457 2177 9491 2178
rect 9457 2144 9460 2177
rect 9460 2144 9491 2177
rect 9376 2009 9410 2013
rect 9376 1979 9380 2009
rect 9380 1979 9410 2009
rect 9566 2109 9600 2123
rect 9566 2089 9600 2109
rect 9842 2280 9876 2340
rect 9930 2280 9964 2340
rect 9842 2142 9876 2202
rect 9930 2142 9964 2202
rect 15807 2211 15841 2245
rect 9886 2049 9920 2083
rect 9650 2009 9684 2012
rect 9650 1978 9680 2009
rect 9680 1978 9684 2009
rect 9789 1979 9823 2013
rect 9827 1886 9861 1920
rect 10086 1904 10120 1938
rect 10087 1811 10121 1845
rect 10528 1809 10562 1843
rect 11260 1809 11294 1843
rect 11386 1809 11420 1843
rect 12472 1809 12506 1843
rect 12598 1809 12632 1843
rect 13684 1809 13718 1843
rect 13810 1809 13844 1843
rect 14896 1809 14930 1843
rect 15022 1809 15056 1843
rect 15627 1831 15661 1891
rect 15715 1831 15749 1891
rect 9329 1743 9363 1777
rect 9421 1748 9455 1777
rect 9513 1748 9547 1777
rect 9421 1743 9428 1748
rect 9428 1743 9455 1748
rect 9513 1743 9546 1748
rect 9546 1743 9547 1748
rect 9605 1743 9639 1777
rect 9697 1743 9731 1777
rect 10484 1690 10518 1750
rect 10572 1690 10606 1750
rect 11216 1690 11250 1750
rect 11321 1690 11355 1750
rect 11430 1690 11464 1750
rect 12428 1690 12462 1750
rect 12532 1690 12566 1750
rect 12642 1690 12676 1750
rect 13640 1690 13674 1750
rect 13745 1690 13779 1750
rect 13854 1690 13888 1750
rect 14852 1690 14886 1750
rect 14959 1690 14993 1750
rect 15066 1690 15100 1750
rect 15627 1693 15661 1753
rect 15715 1693 15749 1753
rect 15811 1693 15845 1753
rect 15907 1693 15941 1753
rect 15556 1602 15590 1636
rect 15763 1600 15797 1634
rect 10837 1489 10871 1549
rect 10927 1489 10961 1549
rect 11569 1489 11603 1549
rect 11676 1489 11710 1549
rect 11779 1489 11813 1549
rect 12781 1489 12815 1549
rect 12887 1489 12921 1549
rect 12991 1489 13025 1549
rect 14119 1489 14153 1549
rect 14227 1489 14261 1549
rect 14329 1489 14363 1549
rect 14974 1489 15008 1549
rect 15063 1489 15097 1549
rect 15627 1490 15661 1550
rect 15715 1490 15749 1550
rect 15811 1490 15845 1550
rect 15907 1490 15941 1550
rect 9897 1415 9931 1449
rect 10881 1405 10915 1439
rect 11613 1405 11647 1439
rect 11735 1405 11769 1439
rect 12825 1405 12859 1439
rect 12947 1405 12981 1439
rect 14163 1405 14197 1439
rect 14285 1405 14319 1439
rect 15019 1405 15053 1439
rect 9817 1305 9851 1365
rect 9977 1305 10011 1365
rect 15627 1352 15661 1412
rect 15715 1352 15749 1412
rect 9817 1167 9851 1227
rect 9977 1167 10011 1227
rect 9817 1029 9851 1089
rect 9977 1029 10011 1089
rect 9817 891 9851 951
rect 9977 891 10011 951
rect 9817 753 9851 813
rect 9977 753 10011 813
rect 9817 615 9851 675
rect 9977 615 10011 675
rect 9817 477 9851 537
rect 9977 477 10011 537
rect 9817 339 9851 399
rect 9977 339 10011 399
rect 10518 318 10552 352
rect 10598 318 10632 352
rect 10678 318 10712 352
rect 10758 318 10792 352
rect 11250 318 11284 352
rect 11330 318 11364 352
rect 11410 318 11444 352
rect 11490 318 11524 352
rect 11858 318 11892 352
rect 11938 318 11972 352
rect 12018 318 12052 352
rect 12098 318 12132 352
rect 12462 318 12496 352
rect 12542 318 12576 352
rect 12622 318 12656 352
rect 12702 318 12736 352
rect 13070 318 13104 352
rect 13150 318 13184 352
rect 13230 318 13264 352
rect 13310 318 13344 352
rect 13800 318 13834 352
rect 13880 318 13914 352
rect 13960 318 13994 352
rect 14040 318 14074 352
rect 14408 318 14442 352
rect 14488 318 14522 352
rect 14568 318 14602 352
rect 14648 318 14682 352
rect 15142 318 15176 352
rect 15222 318 15256 352
rect 15302 318 15336 352
rect 15382 318 15416 352
<< metal1 >>
rect 9963 2937 10053 2953
rect 9963 2926 9982 2937
rect 9945 2904 9982 2926
rect 9836 2892 9882 2904
rect 9836 2832 9842 2892
rect 9876 2832 9882 2892
rect 9836 2754 9882 2832
rect 9924 2892 9982 2904
rect 9924 2832 9930 2892
rect 9964 2885 9982 2892
rect 10034 2931 10642 2937
rect 10034 2885 10080 2931
rect 9964 2879 10080 2885
rect 10132 2879 10160 2931
rect 10212 2879 10240 2931
rect 10292 2879 10320 2931
rect 10372 2879 10400 2931
rect 10452 2879 10480 2931
rect 10532 2879 10642 2931
rect 9964 2871 10642 2879
rect 10704 2931 15612 2937
rect 10704 2879 10812 2931
rect 10864 2879 10892 2931
rect 10944 2879 10972 2931
rect 11024 2879 11052 2931
rect 11104 2879 11132 2931
rect 11184 2879 11212 2931
rect 11264 2879 11416 2931
rect 11468 2879 11496 2931
rect 11548 2879 11576 2931
rect 11628 2879 11656 2931
rect 11708 2879 11736 2931
rect 11788 2879 11816 2931
rect 11868 2879 12024 2931
rect 12076 2879 12104 2931
rect 12156 2879 12184 2931
rect 12236 2879 12264 2931
rect 12316 2879 12344 2931
rect 12396 2879 12424 2931
rect 12476 2879 12628 2931
rect 12680 2879 12708 2931
rect 12760 2879 12788 2931
rect 12840 2879 12868 2931
rect 12920 2879 12948 2931
rect 13000 2879 13028 2931
rect 13080 2879 13236 2931
rect 13288 2879 13316 2931
rect 13368 2879 13396 2931
rect 13448 2879 13476 2931
rect 13528 2879 13556 2931
rect 13608 2879 13636 2931
rect 13688 2879 13840 2931
rect 13892 2879 13920 2931
rect 13972 2879 14000 2931
rect 14052 2879 14080 2931
rect 14132 2879 14160 2931
rect 14212 2879 14240 2931
rect 14292 2879 14448 2931
rect 14500 2879 14528 2931
rect 14580 2879 14608 2931
rect 14660 2879 14688 2931
rect 14740 2879 14768 2931
rect 14820 2879 14848 2931
rect 14900 2879 15052 2931
rect 15104 2879 15132 2931
rect 15184 2879 15212 2931
rect 15264 2879 15292 2931
rect 15344 2879 15372 2931
rect 15424 2879 15452 2931
rect 15504 2879 15612 2931
rect 10704 2871 15612 2879
rect 15772 2875 15862 2891
rect 9964 2870 10053 2871
rect 9964 2832 9970 2870
rect 9924 2820 9970 2832
rect 15772 2823 15791 2875
rect 15843 2823 15862 2875
rect 15772 2807 15862 2823
rect 9836 2694 9842 2754
rect 9876 2694 9882 2754
rect 9836 2682 9882 2694
rect 9924 2754 9970 2766
rect 9924 2694 9930 2754
rect 9964 2694 9970 2754
rect 9836 2616 9882 2628
rect 9836 2556 9842 2616
rect 9876 2556 9882 2616
rect 9836 2478 9882 2556
rect 9924 2616 9970 2694
rect 15777 2731 15867 2747
rect 15777 2679 15796 2731
rect 15848 2679 15867 2731
rect 15777 2663 15867 2679
rect 9924 2556 9930 2616
rect 9964 2556 9970 2616
rect 9924 2544 9970 2556
rect 15778 2579 15868 2595
rect 15778 2527 15797 2579
rect 15849 2527 15868 2579
rect 15778 2511 15868 2527
rect 9836 2418 9842 2478
rect 9876 2418 9882 2478
rect 9836 2406 9882 2418
rect 9924 2478 9970 2490
rect 9924 2418 9930 2478
rect 9964 2418 9970 2478
rect 9300 2332 9760 2352
rect 9300 2321 9365 2332
rect 9300 2287 9329 2321
rect 9363 2287 9365 2321
rect 9300 2280 9365 2287
rect 9417 2331 9640 2332
rect 9417 2321 9496 2331
rect 9548 2321 9640 2331
rect 9417 2287 9421 2321
rect 9455 2287 9496 2321
rect 9548 2287 9605 2321
rect 9639 2287 9640 2321
rect 9417 2280 9496 2287
rect 9300 2279 9496 2280
rect 9548 2280 9640 2287
rect 9692 2321 9760 2332
rect 9692 2287 9697 2321
rect 9731 2287 9760 2321
rect 9692 2280 9760 2287
rect 9548 2279 9760 2280
rect 9300 2256 9760 2279
rect 9836 2340 9882 2352
rect 9836 2280 9842 2340
rect 9876 2280 9882 2340
rect 9836 2202 9882 2280
rect 9924 2340 9970 2418
rect 15778 2409 15868 2425
rect 15778 2357 15797 2409
rect 15849 2357 15868 2409
rect 15778 2341 15868 2357
rect 9924 2280 9930 2340
rect 9964 2280 9970 2340
rect 9924 2268 9970 2280
rect 15777 2252 15867 2268
rect 9445 2178 9808 2185
rect 9445 2144 9457 2178
rect 9491 2157 9808 2178
rect 9491 2144 9503 2157
rect 9445 2137 9503 2144
rect 9550 2123 9617 2129
rect 9550 2089 9566 2123
rect 9600 2110 9617 2123
rect 9600 2089 9752 2110
rect 9550 2082 9752 2089
rect 9630 2021 9696 2023
rect 9368 2016 9422 2020
rect 9367 2013 9422 2016
rect 9238 1979 9376 2013
rect 9410 1979 9422 2013
rect 9367 1976 9422 1979
rect 9367 1972 9421 1976
rect 9630 1969 9638 2021
rect 9690 1969 9696 2021
rect 9630 1968 9696 1969
rect 9724 1938 9752 2082
rect 9780 2025 9808 2157
rect 9836 2142 9842 2202
rect 9876 2142 9882 2202
rect 9836 2130 9882 2142
rect 9924 2202 10027 2214
rect 9924 2142 9930 2202
rect 9964 2142 10027 2202
rect 15777 2200 15796 2252
rect 15848 2200 15867 2252
rect 15777 2184 15867 2200
rect 9924 2130 10027 2142
rect 9874 2083 9943 2089
rect 9874 2049 9886 2083
rect 9920 2049 9943 2083
rect 9874 2043 9943 2049
rect 9780 2013 9829 2025
rect 9780 1979 9789 2013
rect 9823 1979 9829 2013
rect 9780 1966 9829 1979
rect 9724 1920 9867 1938
rect 9724 1910 9827 1920
rect 9818 1886 9827 1910
rect 9861 1886 9867 1920
rect 9818 1873 9867 1886
rect 9300 1786 9760 1808
rect 9300 1777 9383 1786
rect 9435 1777 9503 1786
rect 9555 1777 9646 1786
rect 9698 1777 9760 1786
rect 9300 1743 9329 1777
rect 9363 1743 9383 1777
rect 9455 1743 9503 1777
rect 9555 1743 9605 1777
rect 9639 1743 9646 1777
rect 9731 1743 9760 1777
rect 9300 1734 9383 1743
rect 9435 1734 9503 1743
rect 9555 1734 9646 1743
rect 9698 1734 9760 1743
rect 9300 1712 9760 1734
rect 9895 1643 9943 2043
rect 9275 1596 9943 1643
rect 9895 1455 9943 1596
rect 9885 1449 9943 1455
rect 9644 1443 9709 1444
rect 9644 1442 9650 1443
rect 9548 1440 9650 1442
rect 9546 1394 9650 1440
rect 9644 1391 9650 1394
rect 9702 1391 9709 1443
rect 9885 1415 9897 1449
rect 9931 1415 9943 1449
rect 9885 1409 9943 1415
rect 9981 1640 10027 2130
rect 15695 2010 15785 2026
rect 15695 1999 15714 2010
rect 15620 1958 15714 1999
rect 15766 1958 15785 2010
rect 10077 1943 10126 1950
rect 10077 1938 10696 1943
rect 10077 1904 10086 1938
rect 10120 1904 10696 1938
rect 10077 1896 10696 1904
rect 10077 1891 10126 1896
rect 10078 1849 10127 1857
rect 10647 1849 10696 1896
rect 15620 1940 15785 1958
rect 15620 1894 15667 1940
rect 15621 1891 15667 1894
rect 10078 1845 10579 1849
rect 10078 1811 10087 1845
rect 10121 1843 10579 1845
rect 10121 1811 10528 1843
rect 10078 1809 10528 1811
rect 10562 1809 10579 1843
rect 10078 1803 10579 1809
rect 10647 1843 15068 1849
rect 10647 1809 11260 1843
rect 11294 1809 11386 1843
rect 11420 1809 12472 1843
rect 12506 1809 12598 1843
rect 12632 1809 13684 1843
rect 13718 1809 13810 1843
rect 13844 1809 14896 1843
rect 14930 1809 15022 1843
rect 15056 1809 15068 1843
rect 15621 1831 15627 1891
rect 15661 1831 15667 1891
rect 15621 1819 15667 1831
rect 15709 1891 15755 1903
rect 15709 1831 15715 1891
rect 15749 1831 15755 1891
rect 15709 1822 15755 1831
rect 10647 1803 15068 1809
rect 10078 1802 10567 1803
rect 10647 1802 11093 1803
rect 10078 1798 10127 1802
rect 15709 1793 15947 1822
rect 10478 1754 10524 1762
rect 10455 1753 10534 1754
rect 10455 1689 10462 1753
rect 10526 1689 10534 1753
rect 10566 1750 10612 1762
rect 11210 1754 11256 1762
rect 10566 1690 10572 1750
rect 10606 1690 10612 1750
rect 10478 1678 10524 1689
rect 10566 1640 10612 1690
rect 11187 1753 11266 1754
rect 11187 1689 11194 1753
rect 11258 1689 11266 1753
rect 11315 1750 11361 1762
rect 11424 1754 11470 1762
rect 12422 1754 12468 1762
rect 11315 1690 11321 1750
rect 11355 1690 11361 1750
rect 11210 1678 11256 1689
rect 11315 1640 11361 1690
rect 11414 1753 11493 1754
rect 11414 1689 11422 1753
rect 11486 1689 11493 1753
rect 12399 1753 12478 1754
rect 12399 1689 12406 1753
rect 12470 1689 12478 1753
rect 12526 1750 12572 1762
rect 12636 1754 12682 1762
rect 13634 1754 13680 1762
rect 12526 1690 12532 1750
rect 12566 1690 12572 1750
rect 11424 1678 11470 1689
rect 12422 1678 12468 1689
rect 12526 1640 12572 1690
rect 12626 1753 12705 1754
rect 12626 1689 12634 1753
rect 12698 1689 12705 1753
rect 13611 1753 13690 1754
rect 13611 1689 13618 1753
rect 13682 1689 13690 1753
rect 13739 1750 13785 1762
rect 13848 1754 13894 1762
rect 14846 1754 14892 1762
rect 13739 1690 13745 1750
rect 13779 1690 13785 1750
rect 12636 1678 12682 1689
rect 13634 1678 13680 1689
rect 13739 1640 13785 1690
rect 13838 1753 13917 1754
rect 13838 1689 13846 1753
rect 13910 1689 13917 1753
rect 14823 1753 14902 1754
rect 14823 1689 14830 1753
rect 14894 1689 14902 1753
rect 14953 1750 14999 1762
rect 15060 1754 15106 1762
rect 14953 1690 14959 1750
rect 14993 1690 14999 1750
rect 13848 1678 13894 1689
rect 14846 1678 14892 1689
rect 14953 1640 14999 1690
rect 15050 1753 15129 1754
rect 15050 1689 15058 1753
rect 15122 1689 15129 1753
rect 15621 1753 15667 1765
rect 15621 1693 15627 1753
rect 15661 1693 15667 1753
rect 15060 1678 15106 1689
rect 15621 1681 15667 1693
rect 15709 1753 15755 1793
rect 15709 1693 15715 1753
rect 15749 1693 15755 1753
rect 15709 1681 15755 1693
rect 15783 1753 15873 1765
rect 15783 1749 15811 1753
rect 15845 1749 15873 1753
rect 15783 1697 15802 1749
rect 15854 1697 15873 1749
rect 15783 1693 15811 1697
rect 15845 1693 15873 1697
rect 15783 1681 15873 1693
rect 15901 1753 15947 1793
rect 15901 1693 15907 1753
rect 15941 1693 15947 1753
rect 15901 1681 15947 1693
rect 15540 1640 15606 1642
rect 9981 1636 15606 1640
rect 9981 1602 15556 1636
rect 15590 1602 15606 1636
rect 9981 1598 15606 1602
rect 9981 1377 10027 1598
rect 10831 1551 10877 1561
rect 10809 1487 10818 1551
rect 10882 1487 10891 1551
rect 10809 1486 10891 1487
rect 10921 1549 10967 1598
rect 11563 1551 11609 1561
rect 10921 1489 10927 1549
rect 10961 1489 10967 1549
rect 10831 1477 10877 1486
rect 10921 1477 10967 1489
rect 11541 1487 11550 1551
rect 11614 1487 11623 1551
rect 11541 1486 11623 1487
rect 11670 1549 11716 1598
rect 11773 1551 11819 1561
rect 12775 1551 12821 1561
rect 11670 1489 11676 1549
rect 11710 1489 11716 1549
rect 11563 1477 11609 1486
rect 11670 1477 11716 1489
rect 11759 1487 11768 1551
rect 11832 1487 11841 1551
rect 11759 1486 11841 1487
rect 12753 1487 12762 1551
rect 12826 1487 12835 1551
rect 12753 1486 12835 1487
rect 12881 1549 12927 1598
rect 12985 1551 13031 1561
rect 14113 1551 14159 1561
rect 12881 1489 12887 1549
rect 12921 1489 12927 1549
rect 11773 1477 11819 1486
rect 12775 1477 12821 1486
rect 12881 1477 12927 1489
rect 12971 1487 12980 1551
rect 13044 1487 13053 1551
rect 12971 1486 13053 1487
rect 14091 1487 14100 1551
rect 14164 1487 14173 1551
rect 14091 1486 14173 1487
rect 14221 1549 14267 1598
rect 14323 1551 14369 1561
rect 14221 1489 14227 1549
rect 14261 1489 14267 1549
rect 12985 1477 13031 1486
rect 14113 1477 14159 1486
rect 14221 1477 14267 1489
rect 14309 1487 14318 1551
rect 14382 1487 14391 1551
rect 14309 1486 14391 1487
rect 14968 1549 15014 1598
rect 15544 1596 15606 1598
rect 15639 1633 15667 1681
rect 15751 1634 15933 1640
rect 15751 1633 15763 1634
rect 15639 1604 15763 1633
rect 15639 1562 15667 1604
rect 15751 1600 15763 1604
rect 15797 1600 15933 1634
rect 15751 1594 15933 1600
rect 15057 1551 15103 1561
rect 14968 1489 14974 1549
rect 15008 1489 15014 1549
rect 14323 1477 14369 1486
rect 14968 1477 15014 1489
rect 15043 1487 15052 1551
rect 15116 1487 15125 1551
rect 15043 1486 15125 1487
rect 15621 1550 15667 1562
rect 15621 1490 15627 1550
rect 15661 1490 15667 1550
rect 15057 1477 15103 1486
rect 15621 1478 15667 1490
rect 15709 1550 15755 1562
rect 15709 1490 15715 1550
rect 15749 1490 15755 1550
rect 15709 1450 15755 1490
rect 15783 1550 15873 1562
rect 15783 1546 15811 1550
rect 15845 1546 15873 1550
rect 15783 1494 15802 1546
rect 15854 1494 15873 1546
rect 15783 1490 15811 1494
rect 15845 1490 15873 1494
rect 15783 1478 15873 1490
rect 15901 1550 15947 1562
rect 15901 1490 15907 1550
rect 15941 1490 15947 1550
rect 15901 1450 15947 1490
rect 15009 1445 15068 1448
rect 10131 1391 10138 1443
rect 10190 1441 10196 1443
rect 10869 1441 10927 1445
rect 10190 1439 10927 1441
rect 10190 1405 10881 1439
rect 10915 1424 10927 1439
rect 11601 1439 12997 1445
rect 10915 1405 10929 1424
rect 10190 1394 10929 1405
rect 11601 1405 11613 1439
rect 11647 1405 11735 1439
rect 11769 1405 12825 1439
rect 12859 1405 12947 1439
rect 12981 1405 12997 1439
rect 11601 1399 12997 1405
rect 14151 1439 14335 1445
rect 14151 1405 14163 1439
rect 14197 1405 14285 1439
rect 14319 1405 14335 1439
rect 14151 1399 14335 1405
rect 15007 1439 15068 1445
rect 15007 1405 15019 1439
rect 15053 1405 15068 1439
rect 15007 1399 15068 1405
rect 10190 1391 10196 1394
rect 10131 1390 10196 1391
rect 10871 1389 10929 1394
rect 9811 1365 9857 1377
rect 9811 1305 9817 1365
rect 9851 1305 9857 1365
rect 9811 1227 9857 1305
rect 9971 1365 10027 1377
rect 9971 1305 9977 1365
rect 10011 1305 10027 1365
rect 9971 1293 10027 1305
rect 9811 1167 9817 1227
rect 9851 1167 9857 1227
rect 9811 1155 9857 1167
rect 9971 1227 10017 1239
rect 9971 1167 9977 1227
rect 10011 1167 10017 1227
rect 9811 1089 9857 1101
rect 9811 1029 9817 1089
rect 9851 1029 9857 1089
rect 9811 951 9857 1029
rect 9971 1089 10017 1167
rect 9971 1029 9977 1089
rect 10011 1029 10017 1089
rect 9971 1017 10017 1029
rect 9811 891 9817 951
rect 9851 891 9857 951
rect 9811 879 9857 891
rect 9971 951 10017 963
rect 9971 891 9977 951
rect 10011 891 10017 951
rect 9811 813 9857 825
rect 9811 753 9817 813
rect 9851 753 9857 813
rect 9811 675 9857 753
rect 9971 813 10017 891
rect 9971 753 9977 813
rect 10011 753 10017 813
rect 9971 741 10017 753
rect 9811 615 9817 675
rect 9851 615 9857 675
rect 9811 603 9857 615
rect 9971 675 10017 687
rect 9971 615 9977 675
rect 10011 615 10017 675
rect 9811 537 9857 549
rect 9811 477 9817 537
rect 9851 477 9857 537
rect 9811 399 9857 477
rect 9971 537 10017 615
rect 9971 477 9977 537
rect 10011 477 10017 537
rect 9971 465 10017 477
rect 9811 339 9817 399
rect 9851 339 9857 399
rect 9971 399 10017 411
rect 9971 375 9977 399
rect 9811 327 9857 339
rect 9932 359 9977 375
rect 10011 375 10017 399
rect 10011 359 10039 375
rect 9932 307 9968 359
rect 10020 307 10039 359
rect 9932 291 10039 307
rect 10492 362 10824 368
rect 10492 310 10510 362
rect 10562 310 10590 362
rect 10642 310 10670 362
rect 10722 310 10750 362
rect 10802 310 10824 362
rect 10492 300 10824 310
rect 11224 362 11556 368
rect 11224 310 11242 362
rect 11294 310 11322 362
rect 11374 310 11402 362
rect 11454 310 11482 362
rect 11534 310 11556 362
rect 11224 300 11556 310
rect 11727 268 11785 1399
rect 11826 362 12158 368
rect 11826 310 11848 362
rect 11900 310 11928 362
rect 11980 310 12008 362
rect 12060 310 12088 362
rect 12140 310 12158 362
rect 11826 300 12158 310
rect 12436 362 12768 368
rect 12436 310 12454 362
rect 12506 310 12534 362
rect 12586 310 12614 362
rect 12666 310 12694 362
rect 12746 310 12768 362
rect 12436 300 12768 310
rect 13038 362 13370 368
rect 13038 310 13060 362
rect 13112 310 13140 362
rect 13192 310 13220 362
rect 13272 310 13300 362
rect 13352 310 13370 362
rect 13038 300 13370 310
rect 13774 362 14106 368
rect 13774 310 13792 362
rect 13844 310 13872 362
rect 13924 310 13952 362
rect 14004 310 14032 362
rect 14084 310 14106 362
rect 13774 300 14106 310
rect 14153 268 14211 1399
rect 14376 362 14708 368
rect 14376 310 14398 362
rect 14450 310 14478 362
rect 14530 310 14558 362
rect 14610 310 14638 362
rect 14690 310 14708 362
rect 14376 300 14708 310
rect 15009 267 15068 1399
rect 15621 1412 15667 1424
rect 15621 1352 15627 1412
rect 15661 1352 15667 1412
rect 15621 1300 15667 1352
rect 15709 1421 15947 1450
rect 15709 1412 15755 1421
rect 15709 1352 15715 1412
rect 15749 1352 15755 1412
rect 15709 1340 15755 1352
rect 15621 1284 15782 1300
rect 15621 1232 15711 1284
rect 15763 1232 15782 1284
rect 15621 1216 15782 1232
rect 15110 362 15442 368
rect 15110 310 15132 362
rect 15184 310 15212 362
rect 15264 310 15292 362
rect 15344 310 15372 362
rect 15424 310 15442 362
rect 15110 300 15442 310
<< via1 >>
rect 9982 2885 10034 2937
rect 10080 2919 10132 2931
rect 10080 2885 10090 2919
rect 10090 2885 10124 2919
rect 10124 2885 10132 2919
rect 10080 2879 10132 2885
rect 10160 2919 10212 2931
rect 10160 2885 10170 2919
rect 10170 2885 10204 2919
rect 10204 2885 10212 2919
rect 10160 2879 10212 2885
rect 10240 2919 10292 2931
rect 10240 2885 10250 2919
rect 10250 2885 10284 2919
rect 10284 2885 10292 2919
rect 10240 2879 10292 2885
rect 10320 2919 10372 2931
rect 10320 2885 10330 2919
rect 10330 2885 10364 2919
rect 10364 2885 10372 2919
rect 10320 2879 10372 2885
rect 10400 2919 10452 2931
rect 10400 2885 10410 2919
rect 10410 2885 10444 2919
rect 10444 2885 10452 2919
rect 10400 2879 10452 2885
rect 10480 2919 10532 2931
rect 10480 2885 10490 2919
rect 10490 2885 10524 2919
rect 10524 2885 10532 2919
rect 10480 2879 10532 2885
rect 10812 2919 10864 2931
rect 10812 2885 10822 2919
rect 10822 2885 10856 2919
rect 10856 2885 10864 2919
rect 10812 2879 10864 2885
rect 10892 2919 10944 2931
rect 10892 2885 10902 2919
rect 10902 2885 10936 2919
rect 10936 2885 10944 2919
rect 10892 2879 10944 2885
rect 10972 2919 11024 2931
rect 10972 2885 10982 2919
rect 10982 2885 11016 2919
rect 11016 2885 11024 2919
rect 10972 2879 11024 2885
rect 11052 2919 11104 2931
rect 11052 2885 11062 2919
rect 11062 2885 11096 2919
rect 11096 2885 11104 2919
rect 11052 2879 11104 2885
rect 11132 2919 11184 2931
rect 11132 2885 11142 2919
rect 11142 2885 11176 2919
rect 11176 2885 11184 2919
rect 11132 2879 11184 2885
rect 11212 2919 11264 2931
rect 11212 2885 11222 2919
rect 11222 2885 11256 2919
rect 11256 2885 11264 2919
rect 11212 2879 11264 2885
rect 11416 2919 11468 2931
rect 11416 2885 11424 2919
rect 11424 2885 11458 2919
rect 11458 2885 11468 2919
rect 11416 2879 11468 2885
rect 11496 2919 11548 2931
rect 11496 2885 11504 2919
rect 11504 2885 11538 2919
rect 11538 2885 11548 2919
rect 11496 2879 11548 2885
rect 11576 2919 11628 2931
rect 11576 2885 11584 2919
rect 11584 2885 11618 2919
rect 11618 2885 11628 2919
rect 11576 2879 11628 2885
rect 11656 2919 11708 2931
rect 11656 2885 11664 2919
rect 11664 2885 11698 2919
rect 11698 2885 11708 2919
rect 11656 2879 11708 2885
rect 11736 2919 11788 2931
rect 11736 2885 11744 2919
rect 11744 2885 11778 2919
rect 11778 2885 11788 2919
rect 11736 2879 11788 2885
rect 11816 2919 11868 2931
rect 11816 2885 11824 2919
rect 11824 2885 11858 2919
rect 11858 2885 11868 2919
rect 11816 2879 11868 2885
rect 12024 2919 12076 2931
rect 12024 2885 12034 2919
rect 12034 2885 12068 2919
rect 12068 2885 12076 2919
rect 12024 2879 12076 2885
rect 12104 2919 12156 2931
rect 12104 2885 12114 2919
rect 12114 2885 12148 2919
rect 12148 2885 12156 2919
rect 12104 2879 12156 2885
rect 12184 2919 12236 2931
rect 12184 2885 12194 2919
rect 12194 2885 12228 2919
rect 12228 2885 12236 2919
rect 12184 2879 12236 2885
rect 12264 2919 12316 2931
rect 12264 2885 12274 2919
rect 12274 2885 12308 2919
rect 12308 2885 12316 2919
rect 12264 2879 12316 2885
rect 12344 2919 12396 2931
rect 12344 2885 12354 2919
rect 12354 2885 12388 2919
rect 12388 2885 12396 2919
rect 12344 2879 12396 2885
rect 12424 2919 12476 2931
rect 12424 2885 12434 2919
rect 12434 2885 12468 2919
rect 12468 2885 12476 2919
rect 12424 2879 12476 2885
rect 12628 2919 12680 2931
rect 12628 2885 12636 2919
rect 12636 2885 12670 2919
rect 12670 2885 12680 2919
rect 12628 2879 12680 2885
rect 12708 2919 12760 2931
rect 12708 2885 12716 2919
rect 12716 2885 12750 2919
rect 12750 2885 12760 2919
rect 12708 2879 12760 2885
rect 12788 2919 12840 2931
rect 12788 2885 12796 2919
rect 12796 2885 12830 2919
rect 12830 2885 12840 2919
rect 12788 2879 12840 2885
rect 12868 2919 12920 2931
rect 12868 2885 12876 2919
rect 12876 2885 12910 2919
rect 12910 2885 12920 2919
rect 12868 2879 12920 2885
rect 12948 2919 13000 2931
rect 12948 2885 12956 2919
rect 12956 2885 12990 2919
rect 12990 2885 13000 2919
rect 12948 2879 13000 2885
rect 13028 2919 13080 2931
rect 13028 2885 13036 2919
rect 13036 2885 13070 2919
rect 13070 2885 13080 2919
rect 13028 2879 13080 2885
rect 13236 2919 13288 2931
rect 13236 2885 13246 2919
rect 13246 2885 13280 2919
rect 13280 2885 13288 2919
rect 13236 2879 13288 2885
rect 13316 2919 13368 2931
rect 13316 2885 13326 2919
rect 13326 2885 13360 2919
rect 13360 2885 13368 2919
rect 13316 2879 13368 2885
rect 13396 2919 13448 2931
rect 13396 2885 13406 2919
rect 13406 2885 13440 2919
rect 13440 2885 13448 2919
rect 13396 2879 13448 2885
rect 13476 2919 13528 2931
rect 13476 2885 13486 2919
rect 13486 2885 13520 2919
rect 13520 2885 13528 2919
rect 13476 2879 13528 2885
rect 13556 2919 13608 2931
rect 13556 2885 13566 2919
rect 13566 2885 13600 2919
rect 13600 2885 13608 2919
rect 13556 2879 13608 2885
rect 13636 2919 13688 2931
rect 13636 2885 13646 2919
rect 13646 2885 13680 2919
rect 13680 2885 13688 2919
rect 13636 2879 13688 2885
rect 13840 2919 13892 2931
rect 13840 2885 13848 2919
rect 13848 2885 13882 2919
rect 13882 2885 13892 2919
rect 13840 2879 13892 2885
rect 13920 2919 13972 2931
rect 13920 2885 13928 2919
rect 13928 2885 13962 2919
rect 13962 2885 13972 2919
rect 13920 2879 13972 2885
rect 14000 2919 14052 2931
rect 14000 2885 14008 2919
rect 14008 2885 14042 2919
rect 14042 2885 14052 2919
rect 14000 2879 14052 2885
rect 14080 2919 14132 2931
rect 14080 2885 14088 2919
rect 14088 2885 14122 2919
rect 14122 2885 14132 2919
rect 14080 2879 14132 2885
rect 14160 2919 14212 2931
rect 14160 2885 14168 2919
rect 14168 2885 14202 2919
rect 14202 2885 14212 2919
rect 14160 2879 14212 2885
rect 14240 2919 14292 2931
rect 14240 2885 14248 2919
rect 14248 2885 14282 2919
rect 14282 2885 14292 2919
rect 14240 2879 14292 2885
rect 14448 2919 14500 2931
rect 14448 2885 14458 2919
rect 14458 2885 14492 2919
rect 14492 2885 14500 2919
rect 14448 2879 14500 2885
rect 14528 2919 14580 2931
rect 14528 2885 14538 2919
rect 14538 2885 14572 2919
rect 14572 2885 14580 2919
rect 14528 2879 14580 2885
rect 14608 2919 14660 2931
rect 14608 2885 14618 2919
rect 14618 2885 14652 2919
rect 14652 2885 14660 2919
rect 14608 2879 14660 2885
rect 14688 2919 14740 2931
rect 14688 2885 14698 2919
rect 14698 2885 14732 2919
rect 14732 2885 14740 2919
rect 14688 2879 14740 2885
rect 14768 2919 14820 2931
rect 14768 2885 14778 2919
rect 14778 2885 14812 2919
rect 14812 2885 14820 2919
rect 14768 2879 14820 2885
rect 14848 2919 14900 2931
rect 14848 2885 14858 2919
rect 14858 2885 14892 2919
rect 14892 2885 14900 2919
rect 14848 2879 14900 2885
rect 15052 2919 15104 2931
rect 15052 2885 15060 2919
rect 15060 2885 15094 2919
rect 15094 2885 15104 2919
rect 15052 2879 15104 2885
rect 15132 2919 15184 2931
rect 15132 2885 15140 2919
rect 15140 2885 15174 2919
rect 15174 2885 15184 2919
rect 15132 2879 15184 2885
rect 15212 2919 15264 2931
rect 15212 2885 15220 2919
rect 15220 2885 15254 2919
rect 15254 2885 15264 2919
rect 15212 2879 15264 2885
rect 15292 2919 15344 2931
rect 15292 2885 15300 2919
rect 15300 2885 15334 2919
rect 15334 2885 15344 2919
rect 15292 2879 15344 2885
rect 15372 2919 15424 2931
rect 15372 2885 15380 2919
rect 15380 2885 15414 2919
rect 15414 2885 15424 2919
rect 15372 2879 15424 2885
rect 15452 2919 15504 2931
rect 15452 2885 15460 2919
rect 15460 2885 15494 2919
rect 15494 2885 15504 2919
rect 15452 2879 15504 2885
rect 15791 2868 15843 2875
rect 15791 2834 15802 2868
rect 15802 2834 15836 2868
rect 15836 2834 15843 2868
rect 15791 2823 15843 2834
rect 15796 2724 15848 2731
rect 15796 2690 15807 2724
rect 15807 2690 15841 2724
rect 15841 2690 15848 2724
rect 15796 2679 15848 2690
rect 15797 2572 15849 2579
rect 15797 2538 15808 2572
rect 15808 2538 15842 2572
rect 15842 2538 15849 2572
rect 15797 2527 15849 2538
rect 9365 2280 9417 2332
rect 9496 2321 9548 2331
rect 9496 2287 9513 2321
rect 9513 2287 9547 2321
rect 9547 2287 9548 2321
rect 9496 2279 9548 2287
rect 9640 2280 9692 2332
rect 15797 2402 15849 2409
rect 15797 2368 15808 2402
rect 15808 2368 15842 2402
rect 15842 2368 15849 2402
rect 15797 2357 15849 2368
rect 9638 2012 9690 2021
rect 9638 1978 9650 2012
rect 9650 1978 9684 2012
rect 9684 1978 9690 2012
rect 9638 1969 9690 1978
rect 15796 2245 15848 2252
rect 15796 2211 15807 2245
rect 15807 2211 15841 2245
rect 15841 2211 15848 2245
rect 15796 2200 15848 2211
rect 9383 1777 9435 1786
rect 9503 1777 9555 1786
rect 9646 1777 9698 1786
rect 9383 1743 9421 1777
rect 9421 1743 9435 1777
rect 9503 1743 9513 1777
rect 9513 1743 9547 1777
rect 9547 1743 9555 1777
rect 9646 1743 9697 1777
rect 9697 1743 9698 1777
rect 9383 1734 9435 1743
rect 9503 1734 9555 1743
rect 9646 1734 9698 1743
rect 9650 1391 9702 1443
rect 15714 1958 15766 2010
rect 10462 1750 10526 1753
rect 10462 1690 10484 1750
rect 10484 1690 10518 1750
rect 10518 1690 10526 1750
rect 10462 1689 10526 1690
rect 11194 1750 11258 1753
rect 11194 1690 11216 1750
rect 11216 1690 11250 1750
rect 11250 1690 11258 1750
rect 11194 1689 11258 1690
rect 11422 1750 11486 1753
rect 11422 1690 11430 1750
rect 11430 1690 11464 1750
rect 11464 1690 11486 1750
rect 11422 1689 11486 1690
rect 12406 1750 12470 1753
rect 12406 1690 12428 1750
rect 12428 1690 12462 1750
rect 12462 1690 12470 1750
rect 12406 1689 12470 1690
rect 12634 1750 12698 1753
rect 12634 1690 12642 1750
rect 12642 1690 12676 1750
rect 12676 1690 12698 1750
rect 12634 1689 12698 1690
rect 13618 1750 13682 1753
rect 13618 1690 13640 1750
rect 13640 1690 13674 1750
rect 13674 1690 13682 1750
rect 13618 1689 13682 1690
rect 13846 1750 13910 1753
rect 13846 1690 13854 1750
rect 13854 1690 13888 1750
rect 13888 1690 13910 1750
rect 13846 1689 13910 1690
rect 14830 1750 14894 1753
rect 14830 1690 14852 1750
rect 14852 1690 14886 1750
rect 14886 1690 14894 1750
rect 14830 1689 14894 1690
rect 15058 1750 15122 1753
rect 15058 1690 15066 1750
rect 15066 1690 15100 1750
rect 15100 1690 15122 1750
rect 15058 1689 15122 1690
rect 15802 1697 15811 1749
rect 15811 1697 15845 1749
rect 15845 1697 15854 1749
rect 10818 1549 10882 1551
rect 10818 1489 10837 1549
rect 10837 1489 10871 1549
rect 10871 1489 10882 1549
rect 10818 1487 10882 1489
rect 11550 1549 11614 1551
rect 11550 1489 11569 1549
rect 11569 1489 11603 1549
rect 11603 1489 11614 1549
rect 11550 1487 11614 1489
rect 11768 1549 11832 1551
rect 11768 1489 11779 1549
rect 11779 1489 11813 1549
rect 11813 1489 11832 1549
rect 11768 1487 11832 1489
rect 12762 1549 12826 1551
rect 12762 1489 12781 1549
rect 12781 1489 12815 1549
rect 12815 1489 12826 1549
rect 12762 1487 12826 1489
rect 12980 1549 13044 1551
rect 12980 1489 12991 1549
rect 12991 1489 13025 1549
rect 13025 1489 13044 1549
rect 12980 1487 13044 1489
rect 14100 1549 14164 1551
rect 14100 1489 14119 1549
rect 14119 1489 14153 1549
rect 14153 1489 14164 1549
rect 14100 1487 14164 1489
rect 14318 1549 14382 1551
rect 14318 1489 14329 1549
rect 14329 1489 14363 1549
rect 14363 1489 14382 1549
rect 14318 1487 14382 1489
rect 15052 1549 15116 1551
rect 15052 1489 15063 1549
rect 15063 1489 15097 1549
rect 15097 1489 15116 1549
rect 15052 1487 15116 1489
rect 15802 1494 15811 1546
rect 15811 1494 15845 1546
rect 15845 1494 15854 1546
rect 10138 1391 10190 1443
rect 9968 339 9977 359
rect 9977 339 10011 359
rect 10011 339 10020 359
rect 9968 307 10020 339
rect 10510 352 10562 362
rect 10510 318 10518 352
rect 10518 318 10552 352
rect 10552 318 10562 352
rect 10510 310 10562 318
rect 10590 352 10642 362
rect 10590 318 10598 352
rect 10598 318 10632 352
rect 10632 318 10642 352
rect 10590 310 10642 318
rect 10670 352 10722 362
rect 10670 318 10678 352
rect 10678 318 10712 352
rect 10712 318 10722 352
rect 10670 310 10722 318
rect 10750 352 10802 362
rect 10750 318 10758 352
rect 10758 318 10792 352
rect 10792 318 10802 352
rect 10750 310 10802 318
rect 11242 352 11294 362
rect 11242 318 11250 352
rect 11250 318 11284 352
rect 11284 318 11294 352
rect 11242 310 11294 318
rect 11322 352 11374 362
rect 11322 318 11330 352
rect 11330 318 11364 352
rect 11364 318 11374 352
rect 11322 310 11374 318
rect 11402 352 11454 362
rect 11402 318 11410 352
rect 11410 318 11444 352
rect 11444 318 11454 352
rect 11402 310 11454 318
rect 11482 352 11534 362
rect 11482 318 11490 352
rect 11490 318 11524 352
rect 11524 318 11534 352
rect 11482 310 11534 318
rect 11848 352 11900 362
rect 11848 318 11858 352
rect 11858 318 11892 352
rect 11892 318 11900 352
rect 11848 310 11900 318
rect 11928 352 11980 362
rect 11928 318 11938 352
rect 11938 318 11972 352
rect 11972 318 11980 352
rect 11928 310 11980 318
rect 12008 352 12060 362
rect 12008 318 12018 352
rect 12018 318 12052 352
rect 12052 318 12060 352
rect 12008 310 12060 318
rect 12088 352 12140 362
rect 12088 318 12098 352
rect 12098 318 12132 352
rect 12132 318 12140 352
rect 12088 310 12140 318
rect 12454 352 12506 362
rect 12454 318 12462 352
rect 12462 318 12496 352
rect 12496 318 12506 352
rect 12454 310 12506 318
rect 12534 352 12586 362
rect 12534 318 12542 352
rect 12542 318 12576 352
rect 12576 318 12586 352
rect 12534 310 12586 318
rect 12614 352 12666 362
rect 12614 318 12622 352
rect 12622 318 12656 352
rect 12656 318 12666 352
rect 12614 310 12666 318
rect 12694 352 12746 362
rect 12694 318 12702 352
rect 12702 318 12736 352
rect 12736 318 12746 352
rect 12694 310 12746 318
rect 13060 352 13112 362
rect 13060 318 13070 352
rect 13070 318 13104 352
rect 13104 318 13112 352
rect 13060 310 13112 318
rect 13140 352 13192 362
rect 13140 318 13150 352
rect 13150 318 13184 352
rect 13184 318 13192 352
rect 13140 310 13192 318
rect 13220 352 13272 362
rect 13220 318 13230 352
rect 13230 318 13264 352
rect 13264 318 13272 352
rect 13220 310 13272 318
rect 13300 352 13352 362
rect 13300 318 13310 352
rect 13310 318 13344 352
rect 13344 318 13352 352
rect 13300 310 13352 318
rect 13792 352 13844 362
rect 13792 318 13800 352
rect 13800 318 13834 352
rect 13834 318 13844 352
rect 13792 310 13844 318
rect 13872 352 13924 362
rect 13872 318 13880 352
rect 13880 318 13914 352
rect 13914 318 13924 352
rect 13872 310 13924 318
rect 13952 352 14004 362
rect 13952 318 13960 352
rect 13960 318 13994 352
rect 13994 318 14004 352
rect 13952 310 14004 318
rect 14032 352 14084 362
rect 14032 318 14040 352
rect 14040 318 14074 352
rect 14074 318 14084 352
rect 14032 310 14084 318
rect 14398 352 14450 362
rect 14398 318 14408 352
rect 14408 318 14442 352
rect 14442 318 14450 352
rect 14398 310 14450 318
rect 14478 352 14530 362
rect 14478 318 14488 352
rect 14488 318 14522 352
rect 14522 318 14530 352
rect 14478 310 14530 318
rect 14558 352 14610 362
rect 14558 318 14568 352
rect 14568 318 14602 352
rect 14602 318 14610 352
rect 14558 310 14610 318
rect 14638 352 14690 362
rect 14638 318 14648 352
rect 14648 318 14682 352
rect 14682 318 14690 352
rect 14638 310 14690 318
rect 15711 1232 15763 1284
rect 15132 352 15184 362
rect 15132 318 15142 352
rect 15142 318 15176 352
rect 15176 318 15184 352
rect 15132 310 15184 318
rect 15212 352 15264 362
rect 15212 318 15222 352
rect 15222 318 15256 352
rect 15256 318 15264 352
rect 15212 310 15264 318
rect 15292 352 15344 362
rect 15292 318 15302 352
rect 15302 318 15336 352
rect 15336 318 15344 352
rect 15292 310 15344 318
rect 15372 352 15424 362
rect 15372 318 15382 352
rect 15382 318 15416 352
rect 15416 318 15424 352
rect 15372 310 15424 318
<< metal2 >>
rect 9971 2939 10045 2943
rect 9971 2883 9980 2939
rect 10036 2937 10045 2939
rect 10036 2933 10642 2937
rect 10036 2883 10076 2933
rect 9971 2879 10076 2883
rect 9972 2877 10076 2879
rect 10132 2877 10156 2933
rect 10212 2877 10236 2933
rect 10292 2877 10316 2933
rect 10372 2877 10396 2933
rect 10452 2877 10476 2933
rect 10532 2877 10642 2933
rect 9972 2871 10642 2877
rect 10704 2933 15612 2937
rect 10704 2877 10808 2933
rect 10864 2877 10888 2933
rect 10944 2877 10968 2933
rect 11024 2877 11048 2933
rect 11104 2877 11128 2933
rect 11184 2877 11208 2933
rect 11264 2877 11416 2933
rect 11472 2877 11496 2933
rect 11552 2877 11576 2933
rect 11632 2877 11656 2933
rect 11712 2877 11736 2933
rect 11792 2877 11816 2933
rect 11872 2877 12020 2933
rect 12076 2877 12100 2933
rect 12156 2877 12180 2933
rect 12236 2877 12260 2933
rect 12316 2877 12340 2933
rect 12396 2877 12420 2933
rect 12476 2877 12628 2933
rect 12684 2877 12708 2933
rect 12764 2877 12788 2933
rect 12844 2877 12868 2933
rect 12924 2877 12948 2933
rect 13004 2877 13028 2933
rect 13084 2877 13232 2933
rect 13288 2877 13312 2933
rect 13368 2877 13392 2933
rect 13448 2877 13472 2933
rect 13528 2877 13552 2933
rect 13608 2877 13632 2933
rect 13688 2877 13840 2933
rect 13896 2877 13920 2933
rect 13976 2877 14000 2933
rect 14056 2877 14080 2933
rect 14136 2877 14160 2933
rect 14216 2877 14240 2933
rect 14296 2877 14444 2933
rect 14500 2877 14524 2933
rect 14580 2877 14604 2933
rect 14660 2877 14684 2933
rect 14740 2877 14764 2933
rect 14820 2877 14844 2933
rect 14900 2877 15052 2933
rect 15108 2877 15132 2933
rect 15188 2877 15212 2933
rect 15268 2877 15292 2933
rect 15348 2877 15372 2933
rect 15428 2877 15452 2933
rect 15508 2877 15612 2933
rect 10704 2871 15612 2877
rect 15780 2877 15854 2881
rect 15780 2821 15789 2877
rect 15845 2821 15854 2877
rect 15780 2817 15854 2821
rect 15785 2733 15859 2737
rect 15785 2677 15794 2733
rect 15850 2677 15859 2733
rect 15785 2673 15859 2677
rect 15786 2581 15860 2585
rect 15786 2525 15795 2581
rect 15851 2525 15860 2581
rect 15786 2521 15860 2525
rect 15786 2411 15860 2415
rect 15786 2355 15795 2411
rect 15851 2355 15860 2411
rect 15786 2351 15860 2355
rect 9363 2334 9419 2343
rect 9363 2269 9419 2278
rect 9494 2333 9550 2342
rect 9494 2268 9550 2277
rect 9638 2334 9694 2343
rect 9638 2269 9694 2278
rect 15785 2254 15859 2258
rect 15785 2198 15794 2254
rect 15850 2198 15859 2254
rect 15785 2194 15859 2198
rect 9630 1969 9638 2021
rect 9690 1969 9696 2021
rect 9630 1968 9696 1969
rect 15703 2012 15777 2016
rect 9648 1892 9694 1968
rect 15703 1956 15712 2012
rect 15768 1956 15777 2012
rect 15703 1952 15777 1956
rect 9648 1846 9887 1892
rect 9381 1788 9437 1797
rect 9381 1723 9437 1732
rect 9501 1788 9557 1797
rect 9501 1723 9557 1732
rect 9644 1788 9700 1797
rect 9644 1723 9700 1732
rect 9644 1443 9709 1444
rect 9644 1391 9650 1443
rect 9702 1440 9709 1443
rect 9841 1440 9887 1846
rect 10455 1753 10534 1754
rect 11187 1753 11266 1754
rect 11414 1753 11493 1754
rect 12399 1753 12478 1754
rect 12626 1753 12705 1754
rect 13611 1753 13690 1754
rect 13838 1753 13917 1754
rect 14823 1753 14902 1754
rect 15050 1753 15129 1754
rect 10452 1689 10462 1753
rect 10526 1689 10535 1753
rect 11184 1689 11194 1753
rect 11258 1689 11267 1753
rect 11413 1689 11422 1753
rect 11486 1689 11496 1753
rect 12396 1689 12406 1753
rect 12470 1689 12479 1753
rect 12625 1689 12634 1753
rect 12698 1689 12708 1753
rect 13608 1689 13618 1753
rect 13682 1689 13691 1753
rect 13837 1689 13846 1753
rect 13910 1689 13920 1753
rect 14820 1689 14830 1753
rect 14894 1689 14903 1753
rect 15049 1689 15058 1753
rect 15122 1689 15132 1753
rect 15791 1751 15865 1755
rect 15791 1695 15800 1751
rect 15856 1695 15865 1751
rect 15791 1691 15865 1695
rect 10809 1487 10818 1551
rect 10882 1487 10891 1551
rect 10809 1486 10891 1487
rect 11541 1487 11550 1551
rect 11614 1487 11623 1551
rect 11541 1486 11623 1487
rect 11759 1487 11768 1551
rect 11832 1487 11841 1551
rect 11759 1486 11841 1487
rect 12753 1487 12762 1551
rect 12826 1487 12835 1551
rect 12753 1486 12835 1487
rect 12971 1487 12980 1551
rect 13044 1487 13053 1551
rect 12971 1486 13053 1487
rect 14091 1487 14100 1551
rect 14164 1487 14173 1551
rect 14091 1486 14173 1487
rect 14309 1487 14318 1551
rect 14382 1487 14391 1551
rect 14309 1486 14391 1487
rect 15043 1487 15052 1551
rect 15116 1487 15125 1551
rect 15791 1548 15865 1552
rect 15791 1492 15800 1548
rect 15856 1492 15865 1548
rect 15791 1488 15865 1492
rect 15043 1486 15125 1487
rect 10131 1440 10138 1443
rect 9702 1394 10138 1440
rect 9702 1391 9709 1394
rect 10131 1391 10138 1394
rect 10190 1391 10196 1443
rect 10131 1390 10196 1391
rect 15700 1286 15774 1290
rect 15700 1230 15709 1286
rect 15765 1230 15774 1286
rect 15700 1226 15774 1230
rect 9957 361 10031 365
rect 9957 305 9966 361
rect 10022 305 10031 361
rect 9957 301 10031 305
rect 10492 364 10824 368
rect 10492 308 10508 364
rect 10564 308 10588 364
rect 10644 308 10668 364
rect 10724 308 10748 364
rect 10804 308 10824 364
rect 10492 300 10824 308
rect 11224 364 11556 368
rect 11224 308 11240 364
rect 11296 308 11320 364
rect 11376 308 11400 364
rect 11456 308 11480 364
rect 11536 308 11556 364
rect 11224 300 11556 308
rect 11826 364 12158 368
rect 11826 308 11846 364
rect 11902 308 11926 364
rect 11982 308 12006 364
rect 12062 308 12086 364
rect 12142 308 12158 364
rect 11826 300 12158 308
rect 12436 364 12768 368
rect 12436 308 12452 364
rect 12508 308 12532 364
rect 12588 308 12612 364
rect 12668 308 12692 364
rect 12748 308 12768 364
rect 12436 300 12768 308
rect 13038 364 13370 368
rect 13038 308 13058 364
rect 13114 308 13138 364
rect 13194 308 13218 364
rect 13274 308 13298 364
rect 13354 308 13370 364
rect 13038 300 13370 308
rect 13774 364 14106 368
rect 13774 308 13790 364
rect 13846 308 13870 364
rect 13926 308 13950 364
rect 14006 308 14030 364
rect 14086 308 14106 364
rect 13774 300 14106 308
rect 14376 364 14708 368
rect 14376 308 14396 364
rect 14452 308 14476 364
rect 14532 308 14556 364
rect 14612 308 14636 364
rect 14692 308 14708 364
rect 14376 300 14708 308
rect 15110 364 15442 368
rect 15110 308 15130 364
rect 15186 308 15210 364
rect 15266 308 15290 364
rect 15346 308 15370 364
rect 15426 308 15442 364
rect 15110 300 15442 308
<< via2 >>
rect 9980 2937 10036 2939
rect 9980 2885 9982 2937
rect 9982 2885 10034 2937
rect 10034 2885 10036 2937
rect 9980 2883 10036 2885
rect 10076 2931 10132 2933
rect 10076 2879 10080 2931
rect 10080 2879 10132 2931
rect 10076 2877 10132 2879
rect 10156 2931 10212 2933
rect 10156 2879 10160 2931
rect 10160 2879 10212 2931
rect 10156 2877 10212 2879
rect 10236 2931 10292 2933
rect 10236 2879 10240 2931
rect 10240 2879 10292 2931
rect 10236 2877 10292 2879
rect 10316 2931 10372 2933
rect 10316 2879 10320 2931
rect 10320 2879 10372 2931
rect 10316 2877 10372 2879
rect 10396 2931 10452 2933
rect 10396 2879 10400 2931
rect 10400 2879 10452 2931
rect 10396 2877 10452 2879
rect 10476 2931 10532 2933
rect 10476 2879 10480 2931
rect 10480 2879 10532 2931
rect 10476 2877 10532 2879
rect 10808 2931 10864 2933
rect 10808 2879 10812 2931
rect 10812 2879 10864 2931
rect 10808 2877 10864 2879
rect 10888 2931 10944 2933
rect 10888 2879 10892 2931
rect 10892 2879 10944 2931
rect 10888 2877 10944 2879
rect 10968 2931 11024 2933
rect 10968 2879 10972 2931
rect 10972 2879 11024 2931
rect 10968 2877 11024 2879
rect 11048 2931 11104 2933
rect 11048 2879 11052 2931
rect 11052 2879 11104 2931
rect 11048 2877 11104 2879
rect 11128 2931 11184 2933
rect 11128 2879 11132 2931
rect 11132 2879 11184 2931
rect 11128 2877 11184 2879
rect 11208 2931 11264 2933
rect 11208 2879 11212 2931
rect 11212 2879 11264 2931
rect 11208 2877 11264 2879
rect 11416 2931 11472 2933
rect 11416 2879 11468 2931
rect 11468 2879 11472 2931
rect 11416 2877 11472 2879
rect 11496 2931 11552 2933
rect 11496 2879 11548 2931
rect 11548 2879 11552 2931
rect 11496 2877 11552 2879
rect 11576 2931 11632 2933
rect 11576 2879 11628 2931
rect 11628 2879 11632 2931
rect 11576 2877 11632 2879
rect 11656 2931 11712 2933
rect 11656 2879 11708 2931
rect 11708 2879 11712 2931
rect 11656 2877 11712 2879
rect 11736 2931 11792 2933
rect 11736 2879 11788 2931
rect 11788 2879 11792 2931
rect 11736 2877 11792 2879
rect 11816 2931 11872 2933
rect 11816 2879 11868 2931
rect 11868 2879 11872 2931
rect 11816 2877 11872 2879
rect 12020 2931 12076 2933
rect 12020 2879 12024 2931
rect 12024 2879 12076 2931
rect 12020 2877 12076 2879
rect 12100 2931 12156 2933
rect 12100 2879 12104 2931
rect 12104 2879 12156 2931
rect 12100 2877 12156 2879
rect 12180 2931 12236 2933
rect 12180 2879 12184 2931
rect 12184 2879 12236 2931
rect 12180 2877 12236 2879
rect 12260 2931 12316 2933
rect 12260 2879 12264 2931
rect 12264 2879 12316 2931
rect 12260 2877 12316 2879
rect 12340 2931 12396 2933
rect 12340 2879 12344 2931
rect 12344 2879 12396 2931
rect 12340 2877 12396 2879
rect 12420 2931 12476 2933
rect 12420 2879 12424 2931
rect 12424 2879 12476 2931
rect 12420 2877 12476 2879
rect 12628 2931 12684 2933
rect 12628 2879 12680 2931
rect 12680 2879 12684 2931
rect 12628 2877 12684 2879
rect 12708 2931 12764 2933
rect 12708 2879 12760 2931
rect 12760 2879 12764 2931
rect 12708 2877 12764 2879
rect 12788 2931 12844 2933
rect 12788 2879 12840 2931
rect 12840 2879 12844 2931
rect 12788 2877 12844 2879
rect 12868 2931 12924 2933
rect 12868 2879 12920 2931
rect 12920 2879 12924 2931
rect 12868 2877 12924 2879
rect 12948 2931 13004 2933
rect 12948 2879 13000 2931
rect 13000 2879 13004 2931
rect 12948 2877 13004 2879
rect 13028 2931 13084 2933
rect 13028 2879 13080 2931
rect 13080 2879 13084 2931
rect 13028 2877 13084 2879
rect 13232 2931 13288 2933
rect 13232 2879 13236 2931
rect 13236 2879 13288 2931
rect 13232 2877 13288 2879
rect 13312 2931 13368 2933
rect 13312 2879 13316 2931
rect 13316 2879 13368 2931
rect 13312 2877 13368 2879
rect 13392 2931 13448 2933
rect 13392 2879 13396 2931
rect 13396 2879 13448 2931
rect 13392 2877 13448 2879
rect 13472 2931 13528 2933
rect 13472 2879 13476 2931
rect 13476 2879 13528 2931
rect 13472 2877 13528 2879
rect 13552 2931 13608 2933
rect 13552 2879 13556 2931
rect 13556 2879 13608 2931
rect 13552 2877 13608 2879
rect 13632 2931 13688 2933
rect 13632 2879 13636 2931
rect 13636 2879 13688 2931
rect 13632 2877 13688 2879
rect 13840 2931 13896 2933
rect 13840 2879 13892 2931
rect 13892 2879 13896 2931
rect 13840 2877 13896 2879
rect 13920 2931 13976 2933
rect 13920 2879 13972 2931
rect 13972 2879 13976 2931
rect 13920 2877 13976 2879
rect 14000 2931 14056 2933
rect 14000 2879 14052 2931
rect 14052 2879 14056 2931
rect 14000 2877 14056 2879
rect 14080 2931 14136 2933
rect 14080 2879 14132 2931
rect 14132 2879 14136 2931
rect 14080 2877 14136 2879
rect 14160 2931 14216 2933
rect 14160 2879 14212 2931
rect 14212 2879 14216 2931
rect 14160 2877 14216 2879
rect 14240 2931 14296 2933
rect 14240 2879 14292 2931
rect 14292 2879 14296 2931
rect 14240 2877 14296 2879
rect 14444 2931 14500 2933
rect 14444 2879 14448 2931
rect 14448 2879 14500 2931
rect 14444 2877 14500 2879
rect 14524 2931 14580 2933
rect 14524 2879 14528 2931
rect 14528 2879 14580 2931
rect 14524 2877 14580 2879
rect 14604 2931 14660 2933
rect 14604 2879 14608 2931
rect 14608 2879 14660 2931
rect 14604 2877 14660 2879
rect 14684 2931 14740 2933
rect 14684 2879 14688 2931
rect 14688 2879 14740 2931
rect 14684 2877 14740 2879
rect 14764 2931 14820 2933
rect 14764 2879 14768 2931
rect 14768 2879 14820 2931
rect 14764 2877 14820 2879
rect 14844 2931 14900 2933
rect 14844 2879 14848 2931
rect 14848 2879 14900 2931
rect 14844 2877 14900 2879
rect 15052 2931 15108 2933
rect 15052 2879 15104 2931
rect 15104 2879 15108 2931
rect 15052 2877 15108 2879
rect 15132 2931 15188 2933
rect 15132 2879 15184 2931
rect 15184 2879 15188 2931
rect 15132 2877 15188 2879
rect 15212 2931 15268 2933
rect 15212 2879 15264 2931
rect 15264 2879 15268 2931
rect 15212 2877 15268 2879
rect 15292 2931 15348 2933
rect 15292 2879 15344 2931
rect 15344 2879 15348 2931
rect 15292 2877 15348 2879
rect 15372 2931 15428 2933
rect 15372 2879 15424 2931
rect 15424 2879 15428 2931
rect 15372 2877 15428 2879
rect 15452 2931 15508 2933
rect 15452 2879 15504 2931
rect 15504 2879 15508 2931
rect 15452 2877 15508 2879
rect 15789 2875 15845 2877
rect 15789 2823 15791 2875
rect 15791 2823 15843 2875
rect 15843 2823 15845 2875
rect 15789 2821 15845 2823
rect 15794 2731 15850 2733
rect 15794 2679 15796 2731
rect 15796 2679 15848 2731
rect 15848 2679 15850 2731
rect 15794 2677 15850 2679
rect 15795 2579 15851 2581
rect 15795 2527 15797 2579
rect 15797 2527 15849 2579
rect 15849 2527 15851 2579
rect 15795 2525 15851 2527
rect 15795 2409 15851 2411
rect 15795 2357 15797 2409
rect 15797 2357 15849 2409
rect 15849 2357 15851 2409
rect 15795 2355 15851 2357
rect 9363 2332 9419 2334
rect 9363 2280 9365 2332
rect 9365 2280 9417 2332
rect 9417 2280 9419 2332
rect 9363 2278 9419 2280
rect 9494 2331 9550 2333
rect 9494 2279 9496 2331
rect 9496 2279 9548 2331
rect 9548 2279 9550 2331
rect 9494 2277 9550 2279
rect 9638 2332 9694 2334
rect 9638 2280 9640 2332
rect 9640 2280 9692 2332
rect 9692 2280 9694 2332
rect 9638 2278 9694 2280
rect 15794 2252 15850 2254
rect 15794 2200 15796 2252
rect 15796 2200 15848 2252
rect 15848 2200 15850 2252
rect 15794 2198 15850 2200
rect 15712 2010 15768 2012
rect 15712 1958 15714 2010
rect 15714 1958 15766 2010
rect 15766 1958 15768 2010
rect 15712 1956 15768 1958
rect 9381 1786 9437 1788
rect 9381 1734 9383 1786
rect 9383 1734 9435 1786
rect 9435 1734 9437 1786
rect 9381 1732 9437 1734
rect 9501 1786 9557 1788
rect 9501 1734 9503 1786
rect 9503 1734 9555 1786
rect 9555 1734 9557 1786
rect 9501 1732 9557 1734
rect 9644 1786 9700 1788
rect 9644 1734 9646 1786
rect 9646 1734 9698 1786
rect 9698 1734 9700 1786
rect 9644 1732 9700 1734
rect 10462 1689 10526 1753
rect 11194 1689 11258 1753
rect 11422 1689 11486 1753
rect 12406 1689 12470 1753
rect 12634 1689 12698 1753
rect 13618 1689 13682 1753
rect 13846 1689 13910 1753
rect 14830 1689 14894 1753
rect 15058 1689 15122 1753
rect 15800 1749 15856 1751
rect 15800 1697 15802 1749
rect 15802 1697 15854 1749
rect 15854 1697 15856 1749
rect 15800 1695 15856 1697
rect 10818 1487 10882 1551
rect 11550 1487 11614 1551
rect 11768 1487 11832 1551
rect 12762 1487 12826 1551
rect 12980 1487 13044 1551
rect 14100 1487 14164 1551
rect 14318 1487 14382 1551
rect 15052 1487 15116 1551
rect 15800 1546 15856 1548
rect 15800 1494 15802 1546
rect 15802 1494 15854 1546
rect 15854 1494 15856 1546
rect 15800 1492 15856 1494
rect 15709 1284 15765 1286
rect 15709 1232 15711 1284
rect 15711 1232 15763 1284
rect 15763 1232 15765 1284
rect 15709 1230 15765 1232
rect 9966 359 10022 361
rect 9966 307 9968 359
rect 9968 307 10020 359
rect 10020 307 10022 359
rect 9966 305 10022 307
rect 10508 362 10564 364
rect 10508 310 10510 362
rect 10510 310 10562 362
rect 10562 310 10564 362
rect 10508 308 10564 310
rect 10588 362 10644 364
rect 10588 310 10590 362
rect 10590 310 10642 362
rect 10642 310 10644 362
rect 10588 308 10644 310
rect 10668 362 10724 364
rect 10668 310 10670 362
rect 10670 310 10722 362
rect 10722 310 10724 362
rect 10668 308 10724 310
rect 10748 362 10804 364
rect 10748 310 10750 362
rect 10750 310 10802 362
rect 10802 310 10804 362
rect 10748 308 10804 310
rect 11240 362 11296 364
rect 11240 310 11242 362
rect 11242 310 11294 362
rect 11294 310 11296 362
rect 11240 308 11296 310
rect 11320 362 11376 364
rect 11320 310 11322 362
rect 11322 310 11374 362
rect 11374 310 11376 362
rect 11320 308 11376 310
rect 11400 362 11456 364
rect 11400 310 11402 362
rect 11402 310 11454 362
rect 11454 310 11456 362
rect 11400 308 11456 310
rect 11480 362 11536 364
rect 11480 310 11482 362
rect 11482 310 11534 362
rect 11534 310 11536 362
rect 11480 308 11536 310
rect 11846 362 11902 364
rect 11846 310 11848 362
rect 11848 310 11900 362
rect 11900 310 11902 362
rect 11846 308 11902 310
rect 11926 362 11982 364
rect 11926 310 11928 362
rect 11928 310 11980 362
rect 11980 310 11982 362
rect 11926 308 11982 310
rect 12006 362 12062 364
rect 12006 310 12008 362
rect 12008 310 12060 362
rect 12060 310 12062 362
rect 12006 308 12062 310
rect 12086 362 12142 364
rect 12086 310 12088 362
rect 12088 310 12140 362
rect 12140 310 12142 362
rect 12086 308 12142 310
rect 12452 362 12508 364
rect 12452 310 12454 362
rect 12454 310 12506 362
rect 12506 310 12508 362
rect 12452 308 12508 310
rect 12532 362 12588 364
rect 12532 310 12534 362
rect 12534 310 12586 362
rect 12586 310 12588 362
rect 12532 308 12588 310
rect 12612 362 12668 364
rect 12612 310 12614 362
rect 12614 310 12666 362
rect 12666 310 12668 362
rect 12612 308 12668 310
rect 12692 362 12748 364
rect 12692 310 12694 362
rect 12694 310 12746 362
rect 12746 310 12748 362
rect 12692 308 12748 310
rect 13058 362 13114 364
rect 13058 310 13060 362
rect 13060 310 13112 362
rect 13112 310 13114 362
rect 13058 308 13114 310
rect 13138 362 13194 364
rect 13138 310 13140 362
rect 13140 310 13192 362
rect 13192 310 13194 362
rect 13138 308 13194 310
rect 13218 362 13274 364
rect 13218 310 13220 362
rect 13220 310 13272 362
rect 13272 310 13274 362
rect 13218 308 13274 310
rect 13298 362 13354 364
rect 13298 310 13300 362
rect 13300 310 13352 362
rect 13352 310 13354 362
rect 13298 308 13354 310
rect 13790 362 13846 364
rect 13790 310 13792 362
rect 13792 310 13844 362
rect 13844 310 13846 362
rect 13790 308 13846 310
rect 13870 362 13926 364
rect 13870 310 13872 362
rect 13872 310 13924 362
rect 13924 310 13926 362
rect 13870 308 13926 310
rect 13950 362 14006 364
rect 13950 310 13952 362
rect 13952 310 14004 362
rect 14004 310 14006 362
rect 13950 308 14006 310
rect 14030 362 14086 364
rect 14030 310 14032 362
rect 14032 310 14084 362
rect 14084 310 14086 362
rect 14030 308 14086 310
rect 14396 362 14452 364
rect 14396 310 14398 362
rect 14398 310 14450 362
rect 14450 310 14452 362
rect 14396 308 14452 310
rect 14476 362 14532 364
rect 14476 310 14478 362
rect 14478 310 14530 362
rect 14530 310 14532 362
rect 14476 308 14532 310
rect 14556 362 14612 364
rect 14556 310 14558 362
rect 14558 310 14610 362
rect 14610 310 14612 362
rect 14556 308 14612 310
rect 14636 362 14692 364
rect 14636 310 14638 362
rect 14638 310 14690 362
rect 14690 310 14692 362
rect 14636 308 14692 310
rect 15130 362 15186 364
rect 15130 310 15132 362
rect 15132 310 15184 362
rect 15184 310 15186 362
rect 15130 308 15186 310
rect 15210 362 15266 364
rect 15210 310 15212 362
rect 15212 310 15264 362
rect 15264 310 15266 362
rect 15210 308 15266 310
rect 15290 362 15346 364
rect 15290 310 15292 362
rect 15292 310 15344 362
rect 15344 310 15346 362
rect 15290 308 15346 310
rect 15370 362 15426 364
rect 15370 310 15372 362
rect 15372 310 15424 362
rect 15424 310 15426 362
rect 15370 308 15426 310
<< metal3 >>
rect 9945 2943 10071 2953
rect 9945 2879 9976 2943
rect 10040 2938 10071 2943
rect 10040 2936 10641 2938
rect 10040 2879 10073 2936
rect 9945 2872 10073 2879
rect 10137 2872 10153 2936
rect 10217 2872 10233 2936
rect 10297 2872 10313 2936
rect 10377 2872 10393 2936
rect 10457 2872 10473 2936
rect 10537 2872 10641 2936
rect 9945 2870 10641 2872
rect 10701 2936 15615 2938
rect 10701 2872 10805 2936
rect 10869 2872 10885 2936
rect 10949 2872 10965 2936
rect 11029 2872 11045 2936
rect 11109 2872 11125 2936
rect 11189 2872 11205 2936
rect 11269 2872 11411 2936
rect 11475 2872 11491 2936
rect 11555 2872 11571 2936
rect 11635 2872 11651 2936
rect 11715 2872 11731 2936
rect 11795 2872 11811 2936
rect 11875 2872 12017 2936
rect 12081 2872 12097 2936
rect 12161 2872 12177 2936
rect 12241 2872 12257 2936
rect 12321 2872 12337 2936
rect 12401 2872 12417 2936
rect 12481 2872 12623 2936
rect 12687 2872 12703 2936
rect 12767 2872 12783 2936
rect 12847 2872 12863 2936
rect 12927 2872 12943 2936
rect 13007 2872 13023 2936
rect 13087 2872 13229 2936
rect 13293 2872 13309 2936
rect 13373 2872 13389 2936
rect 13453 2872 13469 2936
rect 13533 2872 13549 2936
rect 13613 2872 13629 2936
rect 13693 2872 13835 2936
rect 13899 2872 13915 2936
rect 13979 2872 13995 2936
rect 14059 2872 14075 2936
rect 14139 2872 14155 2936
rect 14219 2872 14235 2936
rect 14299 2872 14441 2936
rect 14505 2872 14521 2936
rect 14585 2872 14601 2936
rect 14665 2872 14681 2936
rect 14745 2872 14761 2936
rect 14825 2872 14841 2936
rect 14905 2872 15047 2936
rect 15111 2872 15127 2936
rect 15191 2872 15207 2936
rect 15271 2872 15287 2936
rect 15351 2872 15367 2936
rect 15431 2872 15447 2936
rect 15511 2872 15615 2936
rect 10701 2870 15615 2872
rect 15754 2881 15880 2891
rect 9969 2716 10035 2806
rect 9969 2652 9970 2716
rect 10034 2652 10035 2716
rect 9969 2636 10035 2652
rect 9969 2572 9970 2636
rect 10034 2572 10035 2636
rect 9969 2556 10035 2572
rect 9969 2492 9970 2556
rect 10034 2492 10035 2556
rect 9969 2476 10035 2492
rect 9969 2412 9970 2476
rect 10034 2412 10035 2476
rect 9969 2396 10035 2412
rect 9344 2352 9462 2353
rect 9593 2352 9737 2353
rect 9344 2338 9737 2352
rect 9344 2274 9359 2338
rect 9423 2337 9634 2338
rect 9423 2274 9490 2337
rect 9344 2273 9490 2274
rect 9554 2274 9634 2337
rect 9698 2274 9737 2338
rect 9554 2273 9737 2274
rect 9344 2257 9737 2273
rect 9969 2332 9970 2396
rect 10034 2332 10035 2396
rect 9969 2316 10035 2332
rect 9449 2256 9593 2257
rect 9969 2252 9970 2316
rect 10034 2252 10035 2316
rect 9969 2236 10035 2252
rect 9969 2172 9970 2236
rect 10034 2172 10035 2236
rect 9969 2156 10035 2172
rect 9969 2092 9970 2156
rect 10034 2092 10035 2156
rect 9969 2076 10035 2092
rect 9969 2012 9970 2076
rect 10034 2012 10035 2076
rect 9969 1996 10035 2012
rect 9969 1932 9970 1996
rect 10034 1932 10035 1996
rect 9484 1807 9576 1808
rect 9370 1792 9743 1807
rect 9370 1728 9377 1792
rect 9441 1728 9497 1792
rect 9561 1728 9640 1792
rect 9704 1728 9743 1792
rect 9370 1711 9743 1728
rect 9969 1778 10035 1932
rect 10095 1778 10155 2810
rect 10215 1840 10275 2870
rect 10335 1778 10395 2810
rect 10455 1840 10515 2870
rect 10575 2716 10641 2806
rect 10575 2652 10576 2716
rect 10640 2652 10641 2716
rect 10575 2636 10641 2652
rect 10575 2572 10576 2636
rect 10640 2572 10641 2636
rect 10575 2556 10641 2572
rect 10575 2492 10576 2556
rect 10640 2492 10641 2556
rect 10575 2476 10641 2492
rect 10575 2412 10576 2476
rect 10640 2412 10641 2476
rect 10575 2396 10641 2412
rect 10575 2332 10576 2396
rect 10640 2332 10641 2396
rect 10575 2316 10641 2332
rect 10575 2252 10576 2316
rect 10640 2252 10641 2316
rect 10575 2236 10641 2252
rect 10575 2172 10576 2236
rect 10640 2172 10641 2236
rect 10575 2156 10641 2172
rect 10575 2092 10576 2156
rect 10640 2092 10641 2156
rect 10575 2076 10641 2092
rect 10575 2012 10576 2076
rect 10640 2012 10641 2076
rect 10575 1996 10641 2012
rect 10575 1932 10576 1996
rect 10640 1932 10641 1996
rect 10575 1778 10641 1932
rect 9969 1776 10641 1778
rect 9969 1712 10073 1776
rect 10137 1712 10153 1776
rect 10217 1712 10233 1776
rect 10297 1712 10313 1776
rect 10377 1712 10393 1776
rect 10457 1753 10473 1776
rect 10457 1712 10462 1753
rect 10537 1712 10641 1776
rect 9969 1710 10462 1712
rect 10452 1689 10462 1710
rect 10526 1710 10641 1712
rect 10701 2716 10767 2806
rect 10701 2652 10702 2716
rect 10766 2652 10767 2716
rect 10701 2636 10767 2652
rect 10701 2572 10702 2636
rect 10766 2572 10767 2636
rect 10701 2556 10767 2572
rect 10701 2492 10702 2556
rect 10766 2492 10767 2556
rect 10701 2476 10767 2492
rect 10701 2412 10702 2476
rect 10766 2412 10767 2476
rect 10701 2396 10767 2412
rect 10701 2332 10702 2396
rect 10766 2332 10767 2396
rect 10701 2316 10767 2332
rect 10701 2252 10702 2316
rect 10766 2252 10767 2316
rect 10701 2236 10767 2252
rect 10701 2172 10702 2236
rect 10766 2172 10767 2236
rect 10701 2156 10767 2172
rect 10701 2092 10702 2156
rect 10766 2092 10767 2156
rect 10701 2076 10767 2092
rect 10701 2012 10702 2076
rect 10766 2012 10767 2076
rect 10701 1996 10767 2012
rect 10701 1932 10702 1996
rect 10766 1932 10767 1996
rect 10701 1778 10767 1932
rect 10827 1778 10887 2810
rect 10947 1840 11007 2870
rect 11067 1778 11127 2810
rect 11187 1840 11247 2870
rect 11307 2716 11373 2806
rect 11307 2652 11308 2716
rect 11372 2652 11373 2716
rect 11307 2636 11373 2652
rect 11307 2572 11308 2636
rect 11372 2572 11373 2636
rect 11307 2556 11373 2572
rect 11307 2492 11308 2556
rect 11372 2492 11373 2556
rect 11307 2476 11373 2492
rect 11307 2412 11308 2476
rect 11372 2412 11373 2476
rect 11307 2396 11373 2412
rect 11307 2332 11308 2396
rect 11372 2332 11373 2396
rect 11307 2316 11373 2332
rect 11307 2252 11308 2316
rect 11372 2252 11373 2316
rect 11307 2236 11373 2252
rect 11307 2172 11308 2236
rect 11372 2172 11373 2236
rect 11307 2156 11373 2172
rect 11307 2092 11308 2156
rect 11372 2092 11373 2156
rect 11307 2076 11373 2092
rect 11307 2012 11308 2076
rect 11372 2012 11373 2076
rect 11307 1996 11373 2012
rect 11307 1932 11308 1996
rect 11372 1932 11373 1996
rect 11307 1778 11373 1932
rect 11433 1840 11493 2870
rect 11553 1778 11613 2810
rect 11673 1840 11733 2870
rect 11793 1778 11853 2810
rect 11913 2716 11979 2806
rect 11913 2652 11914 2716
rect 11978 2652 11979 2716
rect 11913 2636 11979 2652
rect 11913 2572 11914 2636
rect 11978 2572 11979 2636
rect 11913 2556 11979 2572
rect 11913 2492 11914 2556
rect 11978 2492 11979 2556
rect 11913 2476 11979 2492
rect 11913 2412 11914 2476
rect 11978 2412 11979 2476
rect 11913 2396 11979 2412
rect 11913 2332 11914 2396
rect 11978 2332 11979 2396
rect 11913 2316 11979 2332
rect 11913 2252 11914 2316
rect 11978 2252 11979 2316
rect 11913 2236 11979 2252
rect 11913 2172 11914 2236
rect 11978 2172 11979 2236
rect 11913 2156 11979 2172
rect 11913 2092 11914 2156
rect 11978 2092 11979 2156
rect 11913 2076 11979 2092
rect 11913 2012 11914 2076
rect 11978 2012 11979 2076
rect 11913 1996 11979 2012
rect 11913 1932 11914 1996
rect 11978 1932 11979 1996
rect 11913 1778 11979 1932
rect 12039 1778 12099 2810
rect 12159 1840 12219 2870
rect 12279 1778 12339 2810
rect 12399 1840 12459 2870
rect 12519 2716 12585 2806
rect 12519 2652 12520 2716
rect 12584 2652 12585 2716
rect 12519 2636 12585 2652
rect 12519 2572 12520 2636
rect 12584 2572 12585 2636
rect 12519 2556 12585 2572
rect 12519 2492 12520 2556
rect 12584 2492 12585 2556
rect 12519 2476 12585 2492
rect 12519 2412 12520 2476
rect 12584 2412 12585 2476
rect 12519 2396 12585 2412
rect 12519 2332 12520 2396
rect 12584 2332 12585 2396
rect 12519 2316 12585 2332
rect 12519 2252 12520 2316
rect 12584 2252 12585 2316
rect 12519 2236 12585 2252
rect 12519 2172 12520 2236
rect 12584 2172 12585 2236
rect 12519 2156 12585 2172
rect 12519 2092 12520 2156
rect 12584 2092 12585 2156
rect 12519 2076 12585 2092
rect 12519 2012 12520 2076
rect 12584 2012 12585 2076
rect 12519 1996 12585 2012
rect 12519 1932 12520 1996
rect 12584 1932 12585 1996
rect 12519 1778 12585 1932
rect 12645 1840 12705 2870
rect 12765 1778 12825 2810
rect 12885 1840 12945 2870
rect 13005 1778 13065 2810
rect 13125 2716 13191 2806
rect 13125 2652 13126 2716
rect 13190 2652 13191 2716
rect 13125 2636 13191 2652
rect 13125 2572 13126 2636
rect 13190 2572 13191 2636
rect 13125 2556 13191 2572
rect 13125 2492 13126 2556
rect 13190 2492 13191 2556
rect 13125 2476 13191 2492
rect 13125 2412 13126 2476
rect 13190 2412 13191 2476
rect 13125 2396 13191 2412
rect 13125 2332 13126 2396
rect 13190 2332 13191 2396
rect 13125 2316 13191 2332
rect 13125 2252 13126 2316
rect 13190 2252 13191 2316
rect 13125 2236 13191 2252
rect 13125 2172 13126 2236
rect 13190 2172 13191 2236
rect 13125 2156 13191 2172
rect 13125 2092 13126 2156
rect 13190 2092 13191 2156
rect 13125 2076 13191 2092
rect 13125 2012 13126 2076
rect 13190 2012 13191 2076
rect 13125 1996 13191 2012
rect 13125 1932 13126 1996
rect 13190 1932 13191 1996
rect 13125 1778 13191 1932
rect 13251 1778 13311 2810
rect 13371 1840 13431 2870
rect 13491 1778 13551 2810
rect 13611 1840 13671 2870
rect 13731 2716 13797 2806
rect 13731 2652 13732 2716
rect 13796 2652 13797 2716
rect 13731 2636 13797 2652
rect 13731 2572 13732 2636
rect 13796 2572 13797 2636
rect 13731 2556 13797 2572
rect 13731 2492 13732 2556
rect 13796 2492 13797 2556
rect 13731 2476 13797 2492
rect 13731 2412 13732 2476
rect 13796 2412 13797 2476
rect 13731 2396 13797 2412
rect 13731 2332 13732 2396
rect 13796 2332 13797 2396
rect 13731 2316 13797 2332
rect 13731 2252 13732 2316
rect 13796 2252 13797 2316
rect 13731 2236 13797 2252
rect 13731 2172 13732 2236
rect 13796 2172 13797 2236
rect 13731 2156 13797 2172
rect 13731 2092 13732 2156
rect 13796 2092 13797 2156
rect 13731 2076 13797 2092
rect 13731 2012 13732 2076
rect 13796 2012 13797 2076
rect 13731 1996 13797 2012
rect 13731 1932 13732 1996
rect 13796 1932 13797 1996
rect 13731 1778 13797 1932
rect 13857 1840 13917 2870
rect 13977 1778 14037 2810
rect 14097 1840 14157 2870
rect 14217 1778 14277 2810
rect 14337 2716 14403 2806
rect 14337 2652 14338 2716
rect 14402 2652 14403 2716
rect 14337 2636 14403 2652
rect 14337 2572 14338 2636
rect 14402 2572 14403 2636
rect 14337 2556 14403 2572
rect 14337 2492 14338 2556
rect 14402 2492 14403 2556
rect 14337 2476 14403 2492
rect 14337 2412 14338 2476
rect 14402 2412 14403 2476
rect 14337 2396 14403 2412
rect 14337 2332 14338 2396
rect 14402 2332 14403 2396
rect 14337 2316 14403 2332
rect 14337 2252 14338 2316
rect 14402 2252 14403 2316
rect 14337 2236 14403 2252
rect 14337 2172 14338 2236
rect 14402 2172 14403 2236
rect 14337 2156 14403 2172
rect 14337 2092 14338 2156
rect 14402 2092 14403 2156
rect 14337 2076 14403 2092
rect 14337 2012 14338 2076
rect 14402 2012 14403 2076
rect 14337 1996 14403 2012
rect 14337 1932 14338 1996
rect 14402 1932 14403 1996
rect 14337 1778 14403 1932
rect 14463 1778 14523 2810
rect 14583 1840 14643 2870
rect 14703 1778 14763 2810
rect 14823 1840 14883 2870
rect 14943 2716 15009 2806
rect 14943 2652 14944 2716
rect 15008 2652 15009 2716
rect 14943 2636 15009 2652
rect 14943 2572 14944 2636
rect 15008 2572 15009 2636
rect 14943 2556 15009 2572
rect 14943 2492 14944 2556
rect 15008 2492 15009 2556
rect 14943 2476 15009 2492
rect 14943 2412 14944 2476
rect 15008 2412 15009 2476
rect 14943 2396 15009 2412
rect 14943 2332 14944 2396
rect 15008 2332 15009 2396
rect 14943 2316 15009 2332
rect 14943 2252 14944 2316
rect 15008 2252 15009 2316
rect 14943 2236 15009 2252
rect 14943 2172 14944 2236
rect 15008 2172 15009 2236
rect 14943 2156 15009 2172
rect 14943 2092 14944 2156
rect 15008 2092 15009 2156
rect 14943 2076 15009 2092
rect 14943 2012 14944 2076
rect 15008 2012 15009 2076
rect 14943 1996 15009 2012
rect 14943 1932 14944 1996
rect 15008 1932 15009 1996
rect 14943 1778 15009 1932
rect 15069 1840 15129 2870
rect 15189 1778 15249 2810
rect 15309 1840 15369 2870
rect 15754 2817 15785 2881
rect 15849 2817 15880 2881
rect 15429 1778 15489 2810
rect 15754 2807 15880 2817
rect 15549 2716 15615 2806
rect 15549 2652 15550 2716
rect 15614 2652 15615 2716
rect 15759 2737 15885 2747
rect 15759 2673 15790 2737
rect 15854 2673 15885 2737
rect 15759 2663 15885 2673
rect 15549 2636 15615 2652
rect 15549 2572 15550 2636
rect 15614 2572 15615 2636
rect 15549 2556 15615 2572
rect 15549 2492 15550 2556
rect 15614 2492 15615 2556
rect 15760 2585 15886 2595
rect 15760 2521 15791 2585
rect 15855 2521 15886 2585
rect 15760 2511 15886 2521
rect 15549 2476 15615 2492
rect 15549 2412 15550 2476
rect 15614 2412 15615 2476
rect 15549 2396 15615 2412
rect 15549 2332 15550 2396
rect 15614 2332 15615 2396
rect 15760 2415 15886 2425
rect 15760 2351 15791 2415
rect 15855 2351 15886 2415
rect 15760 2341 15886 2351
rect 15549 2316 15615 2332
rect 15549 2252 15550 2316
rect 15614 2252 15615 2316
rect 15549 2236 15615 2252
rect 15549 2172 15550 2236
rect 15614 2172 15615 2236
rect 15759 2258 15885 2268
rect 15759 2194 15790 2258
rect 15854 2194 15885 2258
rect 15759 2184 15885 2194
rect 15549 2156 15615 2172
rect 15549 2092 15550 2156
rect 15614 2092 15615 2156
rect 15549 2076 15615 2092
rect 15549 2012 15550 2076
rect 15614 2012 15615 2076
rect 15549 1996 15615 2012
rect 15549 1932 15550 1996
rect 15614 1932 15615 1996
rect 15677 2016 15803 2026
rect 15677 1952 15708 2016
rect 15772 1952 15803 2016
rect 15677 1942 15803 1952
rect 15549 1778 15615 1932
rect 10701 1776 15615 1778
rect 10701 1712 10805 1776
rect 10869 1712 10885 1776
rect 10949 1712 10965 1776
rect 11029 1712 11045 1776
rect 11109 1712 11125 1776
rect 11189 1753 11205 1776
rect 11189 1712 11194 1753
rect 11269 1712 11411 1776
rect 11475 1753 11491 1776
rect 11486 1712 11491 1753
rect 11555 1712 11571 1776
rect 11635 1712 11651 1776
rect 11715 1712 11731 1776
rect 11795 1712 11811 1776
rect 11875 1712 12017 1776
rect 12081 1712 12097 1776
rect 12161 1712 12177 1776
rect 12241 1712 12257 1776
rect 12321 1712 12337 1776
rect 12401 1753 12417 1776
rect 12401 1712 12406 1753
rect 12481 1712 12623 1776
rect 12687 1753 12703 1776
rect 12698 1712 12703 1753
rect 12767 1712 12783 1776
rect 12847 1712 12863 1776
rect 12927 1712 12943 1776
rect 13007 1712 13023 1776
rect 13087 1712 13229 1776
rect 13293 1712 13309 1776
rect 13373 1712 13389 1776
rect 13453 1712 13469 1776
rect 13533 1712 13549 1776
rect 13613 1753 13629 1776
rect 13613 1712 13618 1753
rect 13693 1712 13835 1776
rect 13899 1753 13915 1776
rect 13910 1712 13915 1753
rect 13979 1712 13995 1776
rect 14059 1712 14075 1776
rect 14139 1712 14155 1776
rect 14219 1712 14235 1776
rect 14299 1712 14441 1776
rect 14505 1712 14521 1776
rect 14585 1712 14601 1776
rect 14665 1712 14681 1776
rect 14745 1712 14761 1776
rect 14825 1753 14841 1776
rect 14825 1712 14830 1753
rect 14905 1712 15047 1776
rect 15111 1753 15127 1776
rect 15122 1712 15127 1753
rect 15191 1712 15207 1776
rect 15271 1712 15287 1776
rect 15351 1712 15367 1776
rect 15431 1712 15447 1776
rect 15511 1712 15615 1776
rect 10701 1710 11194 1712
rect 10526 1689 10535 1710
rect 10452 1684 10535 1689
rect 11184 1689 11194 1710
rect 11258 1710 11422 1712
rect 11258 1689 11267 1710
rect 11184 1684 11267 1689
rect 11413 1689 11422 1710
rect 11486 1710 12406 1712
rect 11486 1689 11496 1710
rect 11413 1684 11496 1689
rect 12396 1689 12406 1710
rect 12470 1710 12634 1712
rect 12470 1689 12479 1710
rect 12396 1684 12479 1689
rect 12625 1689 12634 1710
rect 12698 1710 13618 1712
rect 12698 1689 12708 1710
rect 12625 1684 12708 1689
rect 13608 1689 13618 1710
rect 13682 1710 13846 1712
rect 13682 1689 13691 1710
rect 13608 1684 13691 1689
rect 13837 1689 13846 1710
rect 13910 1710 14830 1712
rect 13910 1689 13920 1710
rect 13837 1684 13920 1689
rect 14820 1689 14830 1710
rect 14894 1710 15058 1712
rect 14894 1689 14903 1710
rect 14820 1684 14903 1689
rect 15049 1689 15058 1710
rect 15122 1710 15615 1712
rect 15765 1755 15891 1765
rect 15122 1689 15132 1710
rect 15049 1684 15132 1689
rect 15765 1691 15796 1755
rect 15860 1691 15891 1755
rect 15765 1681 15891 1691
rect 10809 1551 10891 1557
rect 10809 1530 10818 1551
rect 10320 1528 10818 1530
rect 10882 1530 10891 1551
rect 11541 1551 11623 1557
rect 11541 1530 11550 1551
rect 10882 1528 10992 1530
rect 10320 1464 10424 1528
rect 10488 1464 10504 1528
rect 10568 1464 10584 1528
rect 10648 1464 10664 1528
rect 10728 1464 10744 1528
rect 10808 1487 10818 1528
rect 10808 1464 10824 1487
rect 10888 1464 10992 1528
rect 10320 1462 10992 1464
rect 10320 1308 10386 1462
rect 10320 1244 10321 1308
rect 10385 1244 10386 1308
rect 10320 1228 10386 1244
rect 10320 1164 10321 1228
rect 10385 1164 10386 1228
rect 10320 1148 10386 1164
rect 10320 1084 10321 1148
rect 10385 1084 10386 1148
rect 10320 1068 10386 1084
rect 10320 1004 10321 1068
rect 10385 1004 10386 1068
rect 10320 988 10386 1004
rect 10320 924 10321 988
rect 10385 924 10386 988
rect 10320 908 10386 924
rect 10320 844 10321 908
rect 10385 844 10386 908
rect 10320 828 10386 844
rect 10320 764 10321 828
rect 10385 764 10386 828
rect 10320 748 10386 764
rect 10320 684 10321 748
rect 10385 684 10386 748
rect 10320 668 10386 684
rect 10320 604 10321 668
rect 10385 604 10386 668
rect 10320 588 10386 604
rect 10320 524 10321 588
rect 10385 524 10386 588
rect 10320 434 10386 524
rect 10446 430 10506 1462
rect 9932 365 10057 375
rect 10566 370 10626 1400
rect 10686 430 10746 1462
rect 10806 370 10866 1400
rect 10926 1308 10992 1462
rect 10926 1244 10927 1308
rect 10991 1244 10992 1308
rect 10926 1228 10992 1244
rect 10926 1164 10927 1228
rect 10991 1164 10992 1228
rect 10926 1148 10992 1164
rect 10926 1084 10927 1148
rect 10991 1084 10992 1148
rect 10926 1068 10992 1084
rect 10926 1004 10927 1068
rect 10991 1004 10992 1068
rect 10926 988 10992 1004
rect 10926 924 10927 988
rect 10991 924 10992 988
rect 10926 908 10992 924
rect 10926 844 10927 908
rect 10991 844 10992 908
rect 10926 828 10992 844
rect 10926 764 10927 828
rect 10991 764 10992 828
rect 10926 748 10992 764
rect 10926 684 10927 748
rect 10991 684 10992 748
rect 10926 668 10992 684
rect 10926 604 10927 668
rect 10991 604 10992 668
rect 10926 588 10992 604
rect 10926 524 10927 588
rect 10991 524 10992 588
rect 10926 434 10992 524
rect 11052 1528 11550 1530
rect 11614 1530 11623 1551
rect 11759 1551 11841 1557
rect 11759 1530 11768 1551
rect 11614 1528 11768 1530
rect 11832 1530 11841 1551
rect 12753 1551 12835 1557
rect 12753 1530 12762 1551
rect 11832 1528 12762 1530
rect 12826 1530 12835 1551
rect 12971 1551 13053 1557
rect 12971 1530 12980 1551
rect 12826 1528 12980 1530
rect 13044 1530 13053 1551
rect 14091 1551 14173 1557
rect 14091 1530 14100 1551
rect 13044 1528 13542 1530
rect 11052 1464 11156 1528
rect 11220 1464 11236 1528
rect 11300 1464 11316 1528
rect 11380 1464 11396 1528
rect 11460 1464 11476 1528
rect 11540 1487 11550 1528
rect 11540 1464 11556 1487
rect 11620 1464 11762 1528
rect 11832 1487 11842 1528
rect 11826 1464 11842 1487
rect 11906 1464 11922 1528
rect 11986 1464 12002 1528
rect 12066 1464 12082 1528
rect 12146 1464 12162 1528
rect 12226 1464 12368 1528
rect 12432 1464 12448 1528
rect 12512 1464 12528 1528
rect 12592 1464 12608 1528
rect 12672 1464 12688 1528
rect 12752 1487 12762 1528
rect 12752 1464 12768 1487
rect 12832 1464 12974 1528
rect 13044 1487 13054 1528
rect 13038 1464 13054 1487
rect 13118 1464 13134 1528
rect 13198 1464 13214 1528
rect 13278 1464 13294 1528
rect 13358 1464 13374 1528
rect 13438 1464 13542 1528
rect 11052 1462 13542 1464
rect 11052 1308 11118 1462
rect 11052 1244 11053 1308
rect 11117 1244 11118 1308
rect 11052 1228 11118 1244
rect 11052 1164 11053 1228
rect 11117 1164 11118 1228
rect 11052 1148 11118 1164
rect 11052 1084 11053 1148
rect 11117 1084 11118 1148
rect 11052 1068 11118 1084
rect 11052 1004 11053 1068
rect 11117 1004 11118 1068
rect 11052 988 11118 1004
rect 11052 924 11053 988
rect 11117 924 11118 988
rect 11052 908 11118 924
rect 11052 844 11053 908
rect 11117 844 11118 908
rect 11052 828 11118 844
rect 11052 764 11053 828
rect 11117 764 11118 828
rect 11052 748 11118 764
rect 11052 684 11053 748
rect 11117 684 11118 748
rect 11052 668 11118 684
rect 11052 604 11053 668
rect 11117 604 11118 668
rect 11052 588 11118 604
rect 11052 524 11053 588
rect 11117 524 11118 588
rect 11052 434 11118 524
rect 11178 430 11238 1462
rect 11298 370 11358 1400
rect 11418 430 11478 1462
rect 11538 370 11598 1400
rect 11658 1308 11724 1462
rect 11658 1244 11659 1308
rect 11723 1244 11724 1308
rect 11658 1228 11724 1244
rect 11658 1164 11659 1228
rect 11723 1164 11724 1228
rect 11658 1148 11724 1164
rect 11658 1084 11659 1148
rect 11723 1084 11724 1148
rect 11658 1068 11724 1084
rect 11658 1004 11659 1068
rect 11723 1004 11724 1068
rect 11658 988 11724 1004
rect 11658 924 11659 988
rect 11723 924 11724 988
rect 11658 908 11724 924
rect 11658 844 11659 908
rect 11723 844 11724 908
rect 11658 828 11724 844
rect 11658 764 11659 828
rect 11723 764 11724 828
rect 11658 748 11724 764
rect 11658 684 11659 748
rect 11723 684 11724 748
rect 11658 668 11724 684
rect 11658 604 11659 668
rect 11723 604 11724 668
rect 11658 588 11724 604
rect 11658 524 11659 588
rect 11723 524 11724 588
rect 11658 434 11724 524
rect 11784 370 11844 1400
rect 11904 430 11964 1462
rect 12024 370 12084 1400
rect 12144 430 12204 1462
rect 12264 1308 12330 1462
rect 12264 1244 12265 1308
rect 12329 1244 12330 1308
rect 12264 1228 12330 1244
rect 12264 1164 12265 1228
rect 12329 1164 12330 1228
rect 12264 1148 12330 1164
rect 12264 1084 12265 1148
rect 12329 1084 12330 1148
rect 12264 1068 12330 1084
rect 12264 1004 12265 1068
rect 12329 1004 12330 1068
rect 12264 988 12330 1004
rect 12264 924 12265 988
rect 12329 924 12330 988
rect 12264 908 12330 924
rect 12264 844 12265 908
rect 12329 844 12330 908
rect 12264 828 12330 844
rect 12264 764 12265 828
rect 12329 764 12330 828
rect 12264 748 12330 764
rect 12264 684 12265 748
rect 12329 684 12330 748
rect 12264 668 12330 684
rect 12264 604 12265 668
rect 12329 604 12330 668
rect 12264 588 12330 604
rect 12264 524 12265 588
rect 12329 524 12330 588
rect 12264 434 12330 524
rect 12390 430 12450 1462
rect 12510 370 12570 1400
rect 12630 430 12690 1462
rect 12750 370 12810 1400
rect 12870 1308 12936 1462
rect 12870 1244 12871 1308
rect 12935 1244 12936 1308
rect 12870 1228 12936 1244
rect 12870 1164 12871 1228
rect 12935 1164 12936 1228
rect 12870 1148 12936 1164
rect 12870 1084 12871 1148
rect 12935 1084 12936 1148
rect 12870 1068 12936 1084
rect 12870 1004 12871 1068
rect 12935 1004 12936 1068
rect 12870 988 12936 1004
rect 12870 924 12871 988
rect 12935 924 12936 988
rect 12870 908 12936 924
rect 12870 844 12871 908
rect 12935 844 12936 908
rect 12870 828 12936 844
rect 12870 764 12871 828
rect 12935 764 12936 828
rect 12870 748 12936 764
rect 12870 684 12871 748
rect 12935 684 12936 748
rect 12870 668 12936 684
rect 12870 604 12871 668
rect 12935 604 12936 668
rect 12870 588 12936 604
rect 12870 524 12871 588
rect 12935 524 12936 588
rect 12870 434 12936 524
rect 12996 370 13056 1400
rect 13116 430 13176 1462
rect 13236 370 13296 1400
rect 13356 430 13416 1462
rect 13476 1308 13542 1462
rect 13476 1244 13477 1308
rect 13541 1244 13542 1308
rect 13476 1228 13542 1244
rect 13476 1164 13477 1228
rect 13541 1164 13542 1228
rect 13476 1148 13542 1164
rect 13476 1084 13477 1148
rect 13541 1084 13542 1148
rect 13476 1068 13542 1084
rect 13476 1004 13477 1068
rect 13541 1004 13542 1068
rect 13476 988 13542 1004
rect 13476 924 13477 988
rect 13541 924 13542 988
rect 13476 908 13542 924
rect 13476 844 13477 908
rect 13541 844 13542 908
rect 13476 828 13542 844
rect 13476 764 13477 828
rect 13541 764 13542 828
rect 13476 748 13542 764
rect 13476 684 13477 748
rect 13541 684 13542 748
rect 13476 668 13542 684
rect 13476 604 13477 668
rect 13541 604 13542 668
rect 13476 588 13542 604
rect 13476 524 13477 588
rect 13541 524 13542 588
rect 13476 434 13542 524
rect 13602 1528 14100 1530
rect 14164 1530 14173 1551
rect 14309 1551 14391 1557
rect 14309 1530 14318 1551
rect 14164 1528 14318 1530
rect 14382 1530 14391 1551
rect 15043 1551 15125 1557
rect 15043 1530 15052 1551
rect 14382 1528 14880 1530
rect 13602 1464 13706 1528
rect 13770 1464 13786 1528
rect 13850 1464 13866 1528
rect 13930 1464 13946 1528
rect 14010 1464 14026 1528
rect 14090 1487 14100 1528
rect 14090 1464 14106 1487
rect 14170 1464 14312 1528
rect 14382 1487 14392 1528
rect 14376 1464 14392 1487
rect 14456 1464 14472 1528
rect 14536 1464 14552 1528
rect 14616 1464 14632 1528
rect 14696 1464 14712 1528
rect 14776 1464 14880 1528
rect 13602 1462 14880 1464
rect 13602 1308 13668 1462
rect 13602 1244 13603 1308
rect 13667 1244 13668 1308
rect 13602 1228 13668 1244
rect 13602 1164 13603 1228
rect 13667 1164 13668 1228
rect 13602 1148 13668 1164
rect 13602 1084 13603 1148
rect 13667 1084 13668 1148
rect 13602 1068 13668 1084
rect 13602 1004 13603 1068
rect 13667 1004 13668 1068
rect 13602 988 13668 1004
rect 13602 924 13603 988
rect 13667 924 13668 988
rect 13602 908 13668 924
rect 13602 844 13603 908
rect 13667 844 13668 908
rect 13602 828 13668 844
rect 13602 764 13603 828
rect 13667 764 13668 828
rect 13602 748 13668 764
rect 13602 684 13603 748
rect 13667 684 13668 748
rect 13602 668 13668 684
rect 13602 604 13603 668
rect 13667 604 13668 668
rect 13602 588 13668 604
rect 13602 524 13603 588
rect 13667 524 13668 588
rect 13602 434 13668 524
rect 13728 430 13788 1462
rect 13848 370 13908 1400
rect 13968 430 14028 1462
rect 14088 370 14148 1400
rect 14208 1308 14274 1462
rect 14208 1244 14209 1308
rect 14273 1244 14274 1308
rect 14208 1228 14274 1244
rect 14208 1164 14209 1228
rect 14273 1164 14274 1228
rect 14208 1148 14274 1164
rect 14208 1084 14209 1148
rect 14273 1084 14274 1148
rect 14208 1068 14274 1084
rect 14208 1004 14209 1068
rect 14273 1004 14274 1068
rect 14208 988 14274 1004
rect 14208 924 14209 988
rect 14273 924 14274 988
rect 14208 908 14274 924
rect 14208 844 14209 908
rect 14273 844 14274 908
rect 14208 828 14274 844
rect 14208 764 14209 828
rect 14273 764 14274 828
rect 14208 748 14274 764
rect 14208 684 14209 748
rect 14273 684 14274 748
rect 14208 668 14274 684
rect 14208 604 14209 668
rect 14273 604 14274 668
rect 14208 588 14274 604
rect 14208 524 14209 588
rect 14273 524 14274 588
rect 14208 434 14274 524
rect 14334 370 14394 1400
rect 14454 430 14514 1462
rect 14574 370 14634 1400
rect 14694 430 14754 1462
rect 14814 1308 14880 1462
rect 14814 1244 14815 1308
rect 14879 1244 14880 1308
rect 14814 1228 14880 1244
rect 14814 1164 14815 1228
rect 14879 1164 14880 1228
rect 14814 1148 14880 1164
rect 14814 1084 14815 1148
rect 14879 1084 14880 1148
rect 14814 1068 14880 1084
rect 14814 1004 14815 1068
rect 14879 1004 14880 1068
rect 14814 988 14880 1004
rect 14814 924 14815 988
rect 14879 924 14880 988
rect 14814 908 14880 924
rect 14814 844 14815 908
rect 14879 844 14880 908
rect 14814 828 14880 844
rect 14814 764 14815 828
rect 14879 764 14880 828
rect 14814 748 14880 764
rect 14814 684 14815 748
rect 14879 684 14880 748
rect 14814 668 14880 684
rect 14814 604 14815 668
rect 14879 604 14880 668
rect 14814 588 14880 604
rect 14814 524 14815 588
rect 14879 524 14880 588
rect 14814 434 14880 524
rect 14942 1528 15052 1530
rect 15116 1530 15125 1551
rect 15765 1552 15891 1562
rect 15116 1528 15614 1530
rect 14942 1464 15046 1528
rect 15116 1487 15126 1528
rect 15110 1464 15126 1487
rect 15190 1464 15206 1528
rect 15270 1464 15286 1528
rect 15350 1464 15366 1528
rect 15430 1464 15446 1528
rect 15510 1464 15614 1528
rect 15765 1488 15796 1552
rect 15860 1488 15891 1552
rect 15765 1478 15891 1488
rect 15791 1477 15865 1478
rect 14942 1462 15614 1464
rect 14942 1308 15008 1462
rect 14942 1244 14943 1308
rect 15007 1244 15008 1308
rect 14942 1228 15008 1244
rect 14942 1164 14943 1228
rect 15007 1164 15008 1228
rect 14942 1148 15008 1164
rect 14942 1084 14943 1148
rect 15007 1084 15008 1148
rect 14942 1068 15008 1084
rect 14942 1004 14943 1068
rect 15007 1004 15008 1068
rect 14942 988 15008 1004
rect 14942 924 14943 988
rect 15007 924 15008 988
rect 14942 908 15008 924
rect 14942 844 14943 908
rect 15007 844 15008 908
rect 14942 828 15008 844
rect 14942 764 14943 828
rect 15007 764 15008 828
rect 14942 748 15008 764
rect 14942 684 14943 748
rect 15007 684 15008 748
rect 14942 668 15008 684
rect 14942 604 14943 668
rect 15007 604 15008 668
rect 14942 588 15008 604
rect 14942 524 14943 588
rect 15007 524 15008 588
rect 14942 434 15008 524
rect 15068 370 15128 1400
rect 15188 430 15248 1462
rect 15308 370 15368 1400
rect 15428 430 15488 1462
rect 15548 1308 15614 1462
rect 15548 1244 15549 1308
rect 15613 1244 15614 1308
rect 15548 1228 15614 1244
rect 15548 1164 15549 1228
rect 15613 1164 15614 1228
rect 15675 1290 15800 1300
rect 15675 1226 15705 1290
rect 15769 1226 15800 1290
rect 15675 1216 15800 1226
rect 15548 1148 15614 1164
rect 15548 1084 15549 1148
rect 15613 1084 15614 1148
rect 15548 1068 15614 1084
rect 15548 1004 15549 1068
rect 15613 1004 15614 1068
rect 15548 988 15614 1004
rect 15548 924 15549 988
rect 15613 924 15614 988
rect 15548 908 15614 924
rect 15548 844 15549 908
rect 15613 844 15614 908
rect 15548 828 15614 844
rect 15548 764 15549 828
rect 15613 764 15614 828
rect 15548 748 15614 764
rect 15548 684 15549 748
rect 15613 684 15614 748
rect 15548 668 15614 684
rect 15548 604 15549 668
rect 15613 604 15614 668
rect 15548 588 15614 604
rect 15548 524 15549 588
rect 15613 524 15614 588
rect 15548 434 15614 524
rect 9932 301 9962 365
rect 10026 301 10057 365
rect 10320 368 10992 370
rect 10320 304 10504 368
rect 10568 304 10584 368
rect 10648 304 10664 368
rect 10728 304 10744 368
rect 10808 304 10992 368
rect 10320 302 10992 304
rect 11052 368 13542 370
rect 11052 304 11236 368
rect 11300 304 11316 368
rect 11380 304 11396 368
rect 11460 304 11476 368
rect 11540 304 11842 368
rect 11906 304 11922 368
rect 11986 304 12002 368
rect 12066 304 12082 368
rect 12146 304 12448 368
rect 12512 304 12528 368
rect 12592 304 12608 368
rect 12672 304 12688 368
rect 12752 304 13054 368
rect 13118 304 13134 368
rect 13198 304 13214 368
rect 13278 304 13294 368
rect 13358 304 13542 368
rect 11052 302 13542 304
rect 13602 368 14880 370
rect 13602 304 13786 368
rect 13850 304 13866 368
rect 13930 304 13946 368
rect 14010 304 14026 368
rect 14090 304 14392 368
rect 14456 304 14472 368
rect 14536 304 14552 368
rect 14616 304 14632 368
rect 14696 304 14880 368
rect 13602 302 14880 304
rect 14942 368 15614 370
rect 14942 304 15126 368
rect 15190 304 15206 368
rect 15270 304 15286 368
rect 15350 304 15366 368
rect 15430 304 15614 368
rect 14942 302 15614 304
rect 9932 291 10057 301
<< via3 >>
rect 9976 2939 10040 2943
rect 9976 2883 9980 2939
rect 9980 2883 10036 2939
rect 10036 2883 10040 2939
rect 9976 2879 10040 2883
rect 10073 2933 10137 2936
rect 10073 2877 10076 2933
rect 10076 2877 10132 2933
rect 10132 2877 10137 2933
rect 10073 2872 10137 2877
rect 10153 2933 10217 2936
rect 10153 2877 10156 2933
rect 10156 2877 10212 2933
rect 10212 2877 10217 2933
rect 10153 2872 10217 2877
rect 10233 2933 10297 2936
rect 10233 2877 10236 2933
rect 10236 2877 10292 2933
rect 10292 2877 10297 2933
rect 10233 2872 10297 2877
rect 10313 2933 10377 2936
rect 10313 2877 10316 2933
rect 10316 2877 10372 2933
rect 10372 2877 10377 2933
rect 10313 2872 10377 2877
rect 10393 2933 10457 2936
rect 10393 2877 10396 2933
rect 10396 2877 10452 2933
rect 10452 2877 10457 2933
rect 10393 2872 10457 2877
rect 10473 2933 10537 2936
rect 10473 2877 10476 2933
rect 10476 2877 10532 2933
rect 10532 2877 10537 2933
rect 10473 2872 10537 2877
rect 10805 2933 10869 2936
rect 10805 2877 10808 2933
rect 10808 2877 10864 2933
rect 10864 2877 10869 2933
rect 10805 2872 10869 2877
rect 10885 2933 10949 2936
rect 10885 2877 10888 2933
rect 10888 2877 10944 2933
rect 10944 2877 10949 2933
rect 10885 2872 10949 2877
rect 10965 2933 11029 2936
rect 10965 2877 10968 2933
rect 10968 2877 11024 2933
rect 11024 2877 11029 2933
rect 10965 2872 11029 2877
rect 11045 2933 11109 2936
rect 11045 2877 11048 2933
rect 11048 2877 11104 2933
rect 11104 2877 11109 2933
rect 11045 2872 11109 2877
rect 11125 2933 11189 2936
rect 11125 2877 11128 2933
rect 11128 2877 11184 2933
rect 11184 2877 11189 2933
rect 11125 2872 11189 2877
rect 11205 2933 11269 2936
rect 11205 2877 11208 2933
rect 11208 2877 11264 2933
rect 11264 2877 11269 2933
rect 11205 2872 11269 2877
rect 11411 2933 11475 2936
rect 11411 2877 11416 2933
rect 11416 2877 11472 2933
rect 11472 2877 11475 2933
rect 11411 2872 11475 2877
rect 11491 2933 11555 2936
rect 11491 2877 11496 2933
rect 11496 2877 11552 2933
rect 11552 2877 11555 2933
rect 11491 2872 11555 2877
rect 11571 2933 11635 2936
rect 11571 2877 11576 2933
rect 11576 2877 11632 2933
rect 11632 2877 11635 2933
rect 11571 2872 11635 2877
rect 11651 2933 11715 2936
rect 11651 2877 11656 2933
rect 11656 2877 11712 2933
rect 11712 2877 11715 2933
rect 11651 2872 11715 2877
rect 11731 2933 11795 2936
rect 11731 2877 11736 2933
rect 11736 2877 11792 2933
rect 11792 2877 11795 2933
rect 11731 2872 11795 2877
rect 11811 2933 11875 2936
rect 11811 2877 11816 2933
rect 11816 2877 11872 2933
rect 11872 2877 11875 2933
rect 11811 2872 11875 2877
rect 12017 2933 12081 2936
rect 12017 2877 12020 2933
rect 12020 2877 12076 2933
rect 12076 2877 12081 2933
rect 12017 2872 12081 2877
rect 12097 2933 12161 2936
rect 12097 2877 12100 2933
rect 12100 2877 12156 2933
rect 12156 2877 12161 2933
rect 12097 2872 12161 2877
rect 12177 2933 12241 2936
rect 12177 2877 12180 2933
rect 12180 2877 12236 2933
rect 12236 2877 12241 2933
rect 12177 2872 12241 2877
rect 12257 2933 12321 2936
rect 12257 2877 12260 2933
rect 12260 2877 12316 2933
rect 12316 2877 12321 2933
rect 12257 2872 12321 2877
rect 12337 2933 12401 2936
rect 12337 2877 12340 2933
rect 12340 2877 12396 2933
rect 12396 2877 12401 2933
rect 12337 2872 12401 2877
rect 12417 2933 12481 2936
rect 12417 2877 12420 2933
rect 12420 2877 12476 2933
rect 12476 2877 12481 2933
rect 12417 2872 12481 2877
rect 12623 2933 12687 2936
rect 12623 2877 12628 2933
rect 12628 2877 12684 2933
rect 12684 2877 12687 2933
rect 12623 2872 12687 2877
rect 12703 2933 12767 2936
rect 12703 2877 12708 2933
rect 12708 2877 12764 2933
rect 12764 2877 12767 2933
rect 12703 2872 12767 2877
rect 12783 2933 12847 2936
rect 12783 2877 12788 2933
rect 12788 2877 12844 2933
rect 12844 2877 12847 2933
rect 12783 2872 12847 2877
rect 12863 2933 12927 2936
rect 12863 2877 12868 2933
rect 12868 2877 12924 2933
rect 12924 2877 12927 2933
rect 12863 2872 12927 2877
rect 12943 2933 13007 2936
rect 12943 2877 12948 2933
rect 12948 2877 13004 2933
rect 13004 2877 13007 2933
rect 12943 2872 13007 2877
rect 13023 2933 13087 2936
rect 13023 2877 13028 2933
rect 13028 2877 13084 2933
rect 13084 2877 13087 2933
rect 13023 2872 13087 2877
rect 13229 2933 13293 2936
rect 13229 2877 13232 2933
rect 13232 2877 13288 2933
rect 13288 2877 13293 2933
rect 13229 2872 13293 2877
rect 13309 2933 13373 2936
rect 13309 2877 13312 2933
rect 13312 2877 13368 2933
rect 13368 2877 13373 2933
rect 13309 2872 13373 2877
rect 13389 2933 13453 2936
rect 13389 2877 13392 2933
rect 13392 2877 13448 2933
rect 13448 2877 13453 2933
rect 13389 2872 13453 2877
rect 13469 2933 13533 2936
rect 13469 2877 13472 2933
rect 13472 2877 13528 2933
rect 13528 2877 13533 2933
rect 13469 2872 13533 2877
rect 13549 2933 13613 2936
rect 13549 2877 13552 2933
rect 13552 2877 13608 2933
rect 13608 2877 13613 2933
rect 13549 2872 13613 2877
rect 13629 2933 13693 2936
rect 13629 2877 13632 2933
rect 13632 2877 13688 2933
rect 13688 2877 13693 2933
rect 13629 2872 13693 2877
rect 13835 2933 13899 2936
rect 13835 2877 13840 2933
rect 13840 2877 13896 2933
rect 13896 2877 13899 2933
rect 13835 2872 13899 2877
rect 13915 2933 13979 2936
rect 13915 2877 13920 2933
rect 13920 2877 13976 2933
rect 13976 2877 13979 2933
rect 13915 2872 13979 2877
rect 13995 2933 14059 2936
rect 13995 2877 14000 2933
rect 14000 2877 14056 2933
rect 14056 2877 14059 2933
rect 13995 2872 14059 2877
rect 14075 2933 14139 2936
rect 14075 2877 14080 2933
rect 14080 2877 14136 2933
rect 14136 2877 14139 2933
rect 14075 2872 14139 2877
rect 14155 2933 14219 2936
rect 14155 2877 14160 2933
rect 14160 2877 14216 2933
rect 14216 2877 14219 2933
rect 14155 2872 14219 2877
rect 14235 2933 14299 2936
rect 14235 2877 14240 2933
rect 14240 2877 14296 2933
rect 14296 2877 14299 2933
rect 14235 2872 14299 2877
rect 14441 2933 14505 2936
rect 14441 2877 14444 2933
rect 14444 2877 14500 2933
rect 14500 2877 14505 2933
rect 14441 2872 14505 2877
rect 14521 2933 14585 2936
rect 14521 2877 14524 2933
rect 14524 2877 14580 2933
rect 14580 2877 14585 2933
rect 14521 2872 14585 2877
rect 14601 2933 14665 2936
rect 14601 2877 14604 2933
rect 14604 2877 14660 2933
rect 14660 2877 14665 2933
rect 14601 2872 14665 2877
rect 14681 2933 14745 2936
rect 14681 2877 14684 2933
rect 14684 2877 14740 2933
rect 14740 2877 14745 2933
rect 14681 2872 14745 2877
rect 14761 2933 14825 2936
rect 14761 2877 14764 2933
rect 14764 2877 14820 2933
rect 14820 2877 14825 2933
rect 14761 2872 14825 2877
rect 14841 2933 14905 2936
rect 14841 2877 14844 2933
rect 14844 2877 14900 2933
rect 14900 2877 14905 2933
rect 14841 2872 14905 2877
rect 15047 2933 15111 2936
rect 15047 2877 15052 2933
rect 15052 2877 15108 2933
rect 15108 2877 15111 2933
rect 15047 2872 15111 2877
rect 15127 2933 15191 2936
rect 15127 2877 15132 2933
rect 15132 2877 15188 2933
rect 15188 2877 15191 2933
rect 15127 2872 15191 2877
rect 15207 2933 15271 2936
rect 15207 2877 15212 2933
rect 15212 2877 15268 2933
rect 15268 2877 15271 2933
rect 15207 2872 15271 2877
rect 15287 2933 15351 2936
rect 15287 2877 15292 2933
rect 15292 2877 15348 2933
rect 15348 2877 15351 2933
rect 15287 2872 15351 2877
rect 15367 2933 15431 2936
rect 15367 2877 15372 2933
rect 15372 2877 15428 2933
rect 15428 2877 15431 2933
rect 15367 2872 15431 2877
rect 15447 2933 15511 2936
rect 15447 2877 15452 2933
rect 15452 2877 15508 2933
rect 15508 2877 15511 2933
rect 15447 2872 15511 2877
rect 9970 2652 10034 2716
rect 9970 2572 10034 2636
rect 9970 2492 10034 2556
rect 9970 2412 10034 2476
rect 9359 2334 9423 2338
rect 9359 2278 9363 2334
rect 9363 2278 9419 2334
rect 9419 2278 9423 2334
rect 9359 2274 9423 2278
rect 9490 2333 9554 2337
rect 9490 2277 9494 2333
rect 9494 2277 9550 2333
rect 9550 2277 9554 2333
rect 9490 2273 9554 2277
rect 9634 2334 9698 2338
rect 9634 2278 9638 2334
rect 9638 2278 9694 2334
rect 9694 2278 9698 2334
rect 9634 2274 9698 2278
rect 9970 2332 10034 2396
rect 9970 2252 10034 2316
rect 9970 2172 10034 2236
rect 9970 2092 10034 2156
rect 9970 2012 10034 2076
rect 9970 1932 10034 1996
rect 9377 1788 9441 1792
rect 9377 1732 9381 1788
rect 9381 1732 9437 1788
rect 9437 1732 9441 1788
rect 9377 1728 9441 1732
rect 9497 1788 9561 1792
rect 9497 1732 9501 1788
rect 9501 1732 9557 1788
rect 9557 1732 9561 1788
rect 9497 1728 9561 1732
rect 9640 1788 9704 1792
rect 9640 1732 9644 1788
rect 9644 1732 9700 1788
rect 9700 1732 9704 1788
rect 9640 1728 9704 1732
rect 10576 2652 10640 2716
rect 10576 2572 10640 2636
rect 10576 2492 10640 2556
rect 10576 2412 10640 2476
rect 10576 2332 10640 2396
rect 10576 2252 10640 2316
rect 10576 2172 10640 2236
rect 10576 2092 10640 2156
rect 10576 2012 10640 2076
rect 10576 1932 10640 1996
rect 10073 1712 10137 1776
rect 10153 1712 10217 1776
rect 10233 1712 10297 1776
rect 10313 1712 10377 1776
rect 10393 1712 10457 1776
rect 10473 1753 10537 1776
rect 10473 1712 10526 1753
rect 10526 1712 10537 1753
rect 10702 2652 10766 2716
rect 10702 2572 10766 2636
rect 10702 2492 10766 2556
rect 10702 2412 10766 2476
rect 10702 2332 10766 2396
rect 10702 2252 10766 2316
rect 10702 2172 10766 2236
rect 10702 2092 10766 2156
rect 10702 2012 10766 2076
rect 10702 1932 10766 1996
rect 11308 2652 11372 2716
rect 11308 2572 11372 2636
rect 11308 2492 11372 2556
rect 11308 2412 11372 2476
rect 11308 2332 11372 2396
rect 11308 2252 11372 2316
rect 11308 2172 11372 2236
rect 11308 2092 11372 2156
rect 11308 2012 11372 2076
rect 11308 1932 11372 1996
rect 11914 2652 11978 2716
rect 11914 2572 11978 2636
rect 11914 2492 11978 2556
rect 11914 2412 11978 2476
rect 11914 2332 11978 2396
rect 11914 2252 11978 2316
rect 11914 2172 11978 2236
rect 11914 2092 11978 2156
rect 11914 2012 11978 2076
rect 11914 1932 11978 1996
rect 12520 2652 12584 2716
rect 12520 2572 12584 2636
rect 12520 2492 12584 2556
rect 12520 2412 12584 2476
rect 12520 2332 12584 2396
rect 12520 2252 12584 2316
rect 12520 2172 12584 2236
rect 12520 2092 12584 2156
rect 12520 2012 12584 2076
rect 12520 1932 12584 1996
rect 13126 2652 13190 2716
rect 13126 2572 13190 2636
rect 13126 2492 13190 2556
rect 13126 2412 13190 2476
rect 13126 2332 13190 2396
rect 13126 2252 13190 2316
rect 13126 2172 13190 2236
rect 13126 2092 13190 2156
rect 13126 2012 13190 2076
rect 13126 1932 13190 1996
rect 13732 2652 13796 2716
rect 13732 2572 13796 2636
rect 13732 2492 13796 2556
rect 13732 2412 13796 2476
rect 13732 2332 13796 2396
rect 13732 2252 13796 2316
rect 13732 2172 13796 2236
rect 13732 2092 13796 2156
rect 13732 2012 13796 2076
rect 13732 1932 13796 1996
rect 14338 2652 14402 2716
rect 14338 2572 14402 2636
rect 14338 2492 14402 2556
rect 14338 2412 14402 2476
rect 14338 2332 14402 2396
rect 14338 2252 14402 2316
rect 14338 2172 14402 2236
rect 14338 2092 14402 2156
rect 14338 2012 14402 2076
rect 14338 1932 14402 1996
rect 14944 2652 15008 2716
rect 14944 2572 15008 2636
rect 14944 2492 15008 2556
rect 14944 2412 15008 2476
rect 14944 2332 15008 2396
rect 14944 2252 15008 2316
rect 14944 2172 15008 2236
rect 14944 2092 15008 2156
rect 14944 2012 15008 2076
rect 14944 1932 15008 1996
rect 15785 2877 15849 2881
rect 15785 2821 15789 2877
rect 15789 2821 15845 2877
rect 15845 2821 15849 2877
rect 15785 2817 15849 2821
rect 15550 2652 15614 2716
rect 15790 2733 15854 2737
rect 15790 2677 15794 2733
rect 15794 2677 15850 2733
rect 15850 2677 15854 2733
rect 15790 2673 15854 2677
rect 15550 2572 15614 2636
rect 15550 2492 15614 2556
rect 15791 2581 15855 2585
rect 15791 2525 15795 2581
rect 15795 2525 15851 2581
rect 15851 2525 15855 2581
rect 15791 2521 15855 2525
rect 15550 2412 15614 2476
rect 15550 2332 15614 2396
rect 15791 2411 15855 2415
rect 15791 2355 15795 2411
rect 15795 2355 15851 2411
rect 15851 2355 15855 2411
rect 15791 2351 15855 2355
rect 15550 2252 15614 2316
rect 15550 2172 15614 2236
rect 15790 2254 15854 2258
rect 15790 2198 15794 2254
rect 15794 2198 15850 2254
rect 15850 2198 15854 2254
rect 15790 2194 15854 2198
rect 15550 2092 15614 2156
rect 15550 2012 15614 2076
rect 15550 1932 15614 1996
rect 15708 2012 15772 2016
rect 15708 1956 15712 2012
rect 15712 1956 15768 2012
rect 15768 1956 15772 2012
rect 15708 1952 15772 1956
rect 10805 1712 10869 1776
rect 10885 1712 10949 1776
rect 10965 1712 11029 1776
rect 11045 1712 11109 1776
rect 11125 1712 11189 1776
rect 11205 1753 11269 1776
rect 11205 1712 11258 1753
rect 11258 1712 11269 1753
rect 11411 1753 11475 1776
rect 11411 1712 11422 1753
rect 11422 1712 11475 1753
rect 11491 1712 11555 1776
rect 11571 1712 11635 1776
rect 11651 1712 11715 1776
rect 11731 1712 11795 1776
rect 11811 1712 11875 1776
rect 12017 1712 12081 1776
rect 12097 1712 12161 1776
rect 12177 1712 12241 1776
rect 12257 1712 12321 1776
rect 12337 1712 12401 1776
rect 12417 1753 12481 1776
rect 12417 1712 12470 1753
rect 12470 1712 12481 1753
rect 12623 1753 12687 1776
rect 12623 1712 12634 1753
rect 12634 1712 12687 1753
rect 12703 1712 12767 1776
rect 12783 1712 12847 1776
rect 12863 1712 12927 1776
rect 12943 1712 13007 1776
rect 13023 1712 13087 1776
rect 13229 1712 13293 1776
rect 13309 1712 13373 1776
rect 13389 1712 13453 1776
rect 13469 1712 13533 1776
rect 13549 1712 13613 1776
rect 13629 1753 13693 1776
rect 13629 1712 13682 1753
rect 13682 1712 13693 1753
rect 13835 1753 13899 1776
rect 13835 1712 13846 1753
rect 13846 1712 13899 1753
rect 13915 1712 13979 1776
rect 13995 1712 14059 1776
rect 14075 1712 14139 1776
rect 14155 1712 14219 1776
rect 14235 1712 14299 1776
rect 14441 1712 14505 1776
rect 14521 1712 14585 1776
rect 14601 1712 14665 1776
rect 14681 1712 14745 1776
rect 14761 1712 14825 1776
rect 14841 1753 14905 1776
rect 14841 1712 14894 1753
rect 14894 1712 14905 1753
rect 15047 1753 15111 1776
rect 15047 1712 15058 1753
rect 15058 1712 15111 1753
rect 15127 1712 15191 1776
rect 15207 1712 15271 1776
rect 15287 1712 15351 1776
rect 15367 1712 15431 1776
rect 15447 1712 15511 1776
rect 15796 1751 15860 1755
rect 15796 1695 15800 1751
rect 15800 1695 15856 1751
rect 15856 1695 15860 1751
rect 15796 1691 15860 1695
rect 10424 1464 10488 1528
rect 10504 1464 10568 1528
rect 10584 1464 10648 1528
rect 10664 1464 10728 1528
rect 10744 1464 10808 1528
rect 10824 1487 10882 1528
rect 10882 1487 10888 1528
rect 10824 1464 10888 1487
rect 10321 1244 10385 1308
rect 10321 1164 10385 1228
rect 10321 1084 10385 1148
rect 10321 1004 10385 1068
rect 10321 924 10385 988
rect 10321 844 10385 908
rect 10321 764 10385 828
rect 10321 684 10385 748
rect 10321 604 10385 668
rect 10321 524 10385 588
rect 10927 1244 10991 1308
rect 10927 1164 10991 1228
rect 10927 1084 10991 1148
rect 10927 1004 10991 1068
rect 10927 924 10991 988
rect 10927 844 10991 908
rect 10927 764 10991 828
rect 10927 684 10991 748
rect 10927 604 10991 668
rect 10927 524 10991 588
rect 11156 1464 11220 1528
rect 11236 1464 11300 1528
rect 11316 1464 11380 1528
rect 11396 1464 11460 1528
rect 11476 1464 11540 1528
rect 11556 1487 11614 1528
rect 11614 1487 11620 1528
rect 11556 1464 11620 1487
rect 11762 1487 11768 1528
rect 11768 1487 11826 1528
rect 11762 1464 11826 1487
rect 11842 1464 11906 1528
rect 11922 1464 11986 1528
rect 12002 1464 12066 1528
rect 12082 1464 12146 1528
rect 12162 1464 12226 1528
rect 12368 1464 12432 1528
rect 12448 1464 12512 1528
rect 12528 1464 12592 1528
rect 12608 1464 12672 1528
rect 12688 1464 12752 1528
rect 12768 1487 12826 1528
rect 12826 1487 12832 1528
rect 12768 1464 12832 1487
rect 12974 1487 12980 1528
rect 12980 1487 13038 1528
rect 12974 1464 13038 1487
rect 13054 1464 13118 1528
rect 13134 1464 13198 1528
rect 13214 1464 13278 1528
rect 13294 1464 13358 1528
rect 13374 1464 13438 1528
rect 11053 1244 11117 1308
rect 11053 1164 11117 1228
rect 11053 1084 11117 1148
rect 11053 1004 11117 1068
rect 11053 924 11117 988
rect 11053 844 11117 908
rect 11053 764 11117 828
rect 11053 684 11117 748
rect 11053 604 11117 668
rect 11053 524 11117 588
rect 11659 1244 11723 1308
rect 11659 1164 11723 1228
rect 11659 1084 11723 1148
rect 11659 1004 11723 1068
rect 11659 924 11723 988
rect 11659 844 11723 908
rect 11659 764 11723 828
rect 11659 684 11723 748
rect 11659 604 11723 668
rect 11659 524 11723 588
rect 12265 1244 12329 1308
rect 12265 1164 12329 1228
rect 12265 1084 12329 1148
rect 12265 1004 12329 1068
rect 12265 924 12329 988
rect 12265 844 12329 908
rect 12265 764 12329 828
rect 12265 684 12329 748
rect 12265 604 12329 668
rect 12265 524 12329 588
rect 12871 1244 12935 1308
rect 12871 1164 12935 1228
rect 12871 1084 12935 1148
rect 12871 1004 12935 1068
rect 12871 924 12935 988
rect 12871 844 12935 908
rect 12871 764 12935 828
rect 12871 684 12935 748
rect 12871 604 12935 668
rect 12871 524 12935 588
rect 13477 1244 13541 1308
rect 13477 1164 13541 1228
rect 13477 1084 13541 1148
rect 13477 1004 13541 1068
rect 13477 924 13541 988
rect 13477 844 13541 908
rect 13477 764 13541 828
rect 13477 684 13541 748
rect 13477 604 13541 668
rect 13477 524 13541 588
rect 13706 1464 13770 1528
rect 13786 1464 13850 1528
rect 13866 1464 13930 1528
rect 13946 1464 14010 1528
rect 14026 1464 14090 1528
rect 14106 1487 14164 1528
rect 14164 1487 14170 1528
rect 14106 1464 14170 1487
rect 14312 1487 14318 1528
rect 14318 1487 14376 1528
rect 14312 1464 14376 1487
rect 14392 1464 14456 1528
rect 14472 1464 14536 1528
rect 14552 1464 14616 1528
rect 14632 1464 14696 1528
rect 14712 1464 14776 1528
rect 13603 1244 13667 1308
rect 13603 1164 13667 1228
rect 13603 1084 13667 1148
rect 13603 1004 13667 1068
rect 13603 924 13667 988
rect 13603 844 13667 908
rect 13603 764 13667 828
rect 13603 684 13667 748
rect 13603 604 13667 668
rect 13603 524 13667 588
rect 14209 1244 14273 1308
rect 14209 1164 14273 1228
rect 14209 1084 14273 1148
rect 14209 1004 14273 1068
rect 14209 924 14273 988
rect 14209 844 14273 908
rect 14209 764 14273 828
rect 14209 684 14273 748
rect 14209 604 14273 668
rect 14209 524 14273 588
rect 14815 1244 14879 1308
rect 14815 1164 14879 1228
rect 14815 1084 14879 1148
rect 14815 1004 14879 1068
rect 14815 924 14879 988
rect 14815 844 14879 908
rect 14815 764 14879 828
rect 14815 684 14879 748
rect 14815 604 14879 668
rect 14815 524 14879 588
rect 15046 1487 15052 1528
rect 15052 1487 15110 1528
rect 15046 1464 15110 1487
rect 15126 1464 15190 1528
rect 15206 1464 15270 1528
rect 15286 1464 15350 1528
rect 15366 1464 15430 1528
rect 15446 1464 15510 1528
rect 15796 1548 15860 1552
rect 15796 1492 15800 1548
rect 15800 1492 15856 1548
rect 15856 1492 15860 1548
rect 15796 1488 15860 1492
rect 14943 1244 15007 1308
rect 14943 1164 15007 1228
rect 14943 1084 15007 1148
rect 14943 1004 15007 1068
rect 14943 924 15007 988
rect 14943 844 15007 908
rect 14943 764 15007 828
rect 14943 684 15007 748
rect 14943 604 15007 668
rect 14943 524 15007 588
rect 15549 1244 15613 1308
rect 15549 1164 15613 1228
rect 15705 1286 15769 1290
rect 15705 1230 15709 1286
rect 15709 1230 15765 1286
rect 15765 1230 15769 1286
rect 15705 1226 15769 1230
rect 15549 1084 15613 1148
rect 15549 1004 15613 1068
rect 15549 924 15613 988
rect 15549 844 15613 908
rect 15549 764 15613 828
rect 15549 684 15613 748
rect 15549 604 15613 668
rect 15549 524 15613 588
rect 9962 361 10026 365
rect 9962 305 9966 361
rect 9966 305 10022 361
rect 10022 305 10026 361
rect 9962 301 10026 305
rect 10504 364 10568 368
rect 10504 308 10508 364
rect 10508 308 10564 364
rect 10564 308 10568 364
rect 10504 304 10568 308
rect 10584 364 10648 368
rect 10584 308 10588 364
rect 10588 308 10644 364
rect 10644 308 10648 364
rect 10584 304 10648 308
rect 10664 364 10728 368
rect 10664 308 10668 364
rect 10668 308 10724 364
rect 10724 308 10728 364
rect 10664 304 10728 308
rect 10744 364 10808 368
rect 10744 308 10748 364
rect 10748 308 10804 364
rect 10804 308 10808 364
rect 10744 304 10808 308
rect 11236 364 11300 368
rect 11236 308 11240 364
rect 11240 308 11296 364
rect 11296 308 11300 364
rect 11236 304 11300 308
rect 11316 364 11380 368
rect 11316 308 11320 364
rect 11320 308 11376 364
rect 11376 308 11380 364
rect 11316 304 11380 308
rect 11396 364 11460 368
rect 11396 308 11400 364
rect 11400 308 11456 364
rect 11456 308 11460 364
rect 11396 304 11460 308
rect 11476 364 11540 368
rect 11476 308 11480 364
rect 11480 308 11536 364
rect 11536 308 11540 364
rect 11476 304 11540 308
rect 11842 364 11906 368
rect 11842 308 11846 364
rect 11846 308 11902 364
rect 11902 308 11906 364
rect 11842 304 11906 308
rect 11922 364 11986 368
rect 11922 308 11926 364
rect 11926 308 11982 364
rect 11982 308 11986 364
rect 11922 304 11986 308
rect 12002 364 12066 368
rect 12002 308 12006 364
rect 12006 308 12062 364
rect 12062 308 12066 364
rect 12002 304 12066 308
rect 12082 364 12146 368
rect 12082 308 12086 364
rect 12086 308 12142 364
rect 12142 308 12146 364
rect 12082 304 12146 308
rect 12448 364 12512 368
rect 12448 308 12452 364
rect 12452 308 12508 364
rect 12508 308 12512 364
rect 12448 304 12512 308
rect 12528 364 12592 368
rect 12528 308 12532 364
rect 12532 308 12588 364
rect 12588 308 12592 364
rect 12528 304 12592 308
rect 12608 364 12672 368
rect 12608 308 12612 364
rect 12612 308 12668 364
rect 12668 308 12672 364
rect 12608 304 12672 308
rect 12688 364 12752 368
rect 12688 308 12692 364
rect 12692 308 12748 364
rect 12748 308 12752 364
rect 12688 304 12752 308
rect 13054 364 13118 368
rect 13054 308 13058 364
rect 13058 308 13114 364
rect 13114 308 13118 364
rect 13054 304 13118 308
rect 13134 364 13198 368
rect 13134 308 13138 364
rect 13138 308 13194 364
rect 13194 308 13198 364
rect 13134 304 13198 308
rect 13214 364 13278 368
rect 13214 308 13218 364
rect 13218 308 13274 364
rect 13274 308 13278 364
rect 13214 304 13278 308
rect 13294 364 13358 368
rect 13294 308 13298 364
rect 13298 308 13354 364
rect 13354 308 13358 364
rect 13294 304 13358 308
rect 13786 364 13850 368
rect 13786 308 13790 364
rect 13790 308 13846 364
rect 13846 308 13850 364
rect 13786 304 13850 308
rect 13866 364 13930 368
rect 13866 308 13870 364
rect 13870 308 13926 364
rect 13926 308 13930 364
rect 13866 304 13930 308
rect 13946 364 14010 368
rect 13946 308 13950 364
rect 13950 308 14006 364
rect 14006 308 14010 364
rect 13946 304 14010 308
rect 14026 364 14090 368
rect 14026 308 14030 364
rect 14030 308 14086 364
rect 14086 308 14090 364
rect 14026 304 14090 308
rect 14392 364 14456 368
rect 14392 308 14396 364
rect 14396 308 14452 364
rect 14452 308 14456 364
rect 14392 304 14456 308
rect 14472 364 14536 368
rect 14472 308 14476 364
rect 14476 308 14532 364
rect 14532 308 14536 364
rect 14472 304 14536 308
rect 14552 364 14616 368
rect 14552 308 14556 364
rect 14556 308 14612 364
rect 14612 308 14616 364
rect 14552 304 14616 308
rect 14632 364 14696 368
rect 14632 308 14636 364
rect 14636 308 14692 364
rect 14692 308 14696 364
rect 14632 304 14696 308
rect 15126 364 15190 368
rect 15126 308 15130 364
rect 15130 308 15186 364
rect 15186 308 15190 364
rect 15126 304 15190 308
rect 15206 364 15270 368
rect 15206 308 15210 364
rect 15210 308 15266 364
rect 15266 308 15270 364
rect 15206 304 15270 308
rect 15286 364 15350 368
rect 15286 308 15290 364
rect 15290 308 15346 364
rect 15346 308 15350 364
rect 15286 304 15350 308
rect 15366 364 15430 368
rect 15366 308 15370 364
rect 15370 308 15426 364
rect 15426 308 15430 364
rect 15366 304 15430 308
<< metal4 >>
rect 9945 2948 10071 2953
rect 9344 2943 15993 2948
rect 9344 2879 9976 2943
rect 10040 2936 15993 2943
rect 10040 2879 10073 2936
rect 9344 2872 10073 2879
rect 10137 2872 10153 2936
rect 10217 2872 10233 2936
rect 10297 2872 10313 2936
rect 10377 2872 10393 2936
rect 10457 2872 10473 2936
rect 10537 2872 10805 2936
rect 10869 2872 10885 2936
rect 10949 2872 10965 2936
rect 11029 2872 11045 2936
rect 11109 2872 11125 2936
rect 11189 2872 11205 2936
rect 11269 2872 11411 2936
rect 11475 2872 11491 2936
rect 11555 2872 11571 2936
rect 11635 2872 11651 2936
rect 11715 2872 11731 2936
rect 11795 2872 11811 2936
rect 11875 2872 12017 2936
rect 12081 2872 12097 2936
rect 12161 2872 12177 2936
rect 12241 2872 12257 2936
rect 12321 2872 12337 2936
rect 12401 2872 12417 2936
rect 12481 2872 12623 2936
rect 12687 2872 12703 2936
rect 12767 2872 12783 2936
rect 12847 2872 12863 2936
rect 12927 2872 12943 2936
rect 13007 2872 13023 2936
rect 13087 2872 13229 2936
rect 13293 2872 13309 2936
rect 13373 2872 13389 2936
rect 13453 2872 13469 2936
rect 13533 2872 13549 2936
rect 13613 2872 13629 2936
rect 13693 2872 13835 2936
rect 13899 2872 13915 2936
rect 13979 2872 13995 2936
rect 14059 2872 14075 2936
rect 14139 2872 14155 2936
rect 14219 2872 14235 2936
rect 14299 2872 14441 2936
rect 14505 2872 14521 2936
rect 14585 2872 14601 2936
rect 14665 2872 14681 2936
rect 14745 2872 14761 2936
rect 14825 2872 14841 2936
rect 14905 2872 15047 2936
rect 15111 2872 15127 2936
rect 15191 2872 15207 2936
rect 15271 2872 15287 2936
rect 15351 2872 15367 2936
rect 15431 2872 15447 2936
rect 15511 2881 15993 2936
rect 15511 2872 15785 2881
rect 9344 2870 15785 2872
rect 9344 2338 9762 2870
rect 9344 2274 9359 2338
rect 9423 2337 9634 2338
rect 9423 2274 9490 2337
rect 9344 2273 9490 2274
rect 9554 2274 9634 2337
rect 9698 2332 9762 2338
rect 9969 2716 10035 2806
rect 9969 2652 9970 2716
rect 10034 2652 10035 2716
rect 9969 2636 10035 2652
rect 9969 2572 9970 2636
rect 10034 2572 10035 2636
rect 9969 2556 10035 2572
rect 9969 2492 9970 2556
rect 10034 2492 10035 2556
rect 9969 2476 10035 2492
rect 9969 2412 9970 2476
rect 10034 2412 10035 2476
rect 9969 2396 10035 2412
rect 9969 2332 9970 2396
rect 10034 2332 10035 2396
rect 9698 2274 9761 2332
rect 9554 2273 9761 2274
rect 9344 2255 9761 2273
rect 9969 2316 10035 2332
rect 9969 2252 9970 2316
rect 10034 2252 10035 2316
rect 9969 2236 10035 2252
rect 9969 2172 9970 2236
rect 10034 2172 10035 2236
rect 9969 2156 10035 2172
rect 9969 2092 9970 2156
rect 10034 2092 10035 2156
rect 9969 2076 10035 2092
rect 9969 2012 9970 2076
rect 10034 2012 10035 2076
rect 9969 1996 10035 2012
rect 9969 1932 9970 1996
rect 10034 1932 10035 1996
rect 9370 1792 9747 1807
rect 9370 1728 9377 1792
rect 9441 1728 9497 1792
rect 9561 1728 9640 1792
rect 9704 1728 9747 1792
rect 9969 1778 10035 1932
rect 10095 1840 10155 2870
rect 10215 1778 10275 2810
rect 10335 1840 10395 2870
rect 10455 1778 10515 2810
rect 10575 2716 10641 2806
rect 10575 2652 10576 2716
rect 10640 2652 10641 2716
rect 10575 2636 10641 2652
rect 10575 2572 10576 2636
rect 10640 2572 10641 2636
rect 10575 2556 10641 2572
rect 10575 2492 10576 2556
rect 10640 2492 10641 2556
rect 10575 2476 10641 2492
rect 10575 2412 10576 2476
rect 10640 2412 10641 2476
rect 10575 2396 10641 2412
rect 10575 2332 10576 2396
rect 10640 2332 10641 2396
rect 10575 2316 10641 2332
rect 10575 2252 10576 2316
rect 10640 2252 10641 2316
rect 10575 2236 10641 2252
rect 10575 2172 10576 2236
rect 10640 2172 10641 2236
rect 10575 2156 10641 2172
rect 10575 2092 10576 2156
rect 10640 2092 10641 2156
rect 10575 2076 10641 2092
rect 10575 2012 10576 2076
rect 10640 2012 10641 2076
rect 10575 1996 10641 2012
rect 10575 1932 10576 1996
rect 10640 1932 10641 1996
rect 10575 1778 10641 1932
rect 9969 1776 10641 1778
rect 9372 369 9748 1728
rect 9969 1712 10073 1776
rect 10137 1712 10153 1776
rect 10217 1712 10233 1776
rect 10297 1712 10313 1776
rect 10377 1712 10393 1776
rect 10457 1712 10473 1776
rect 10537 1712 10641 1776
rect 9969 1710 10641 1712
rect 10701 2716 10767 2806
rect 10701 2652 10702 2716
rect 10766 2652 10767 2716
rect 10701 2636 10767 2652
rect 10701 2572 10702 2636
rect 10766 2572 10767 2636
rect 10701 2556 10767 2572
rect 10701 2492 10702 2556
rect 10766 2492 10767 2556
rect 10701 2476 10767 2492
rect 10701 2412 10702 2476
rect 10766 2412 10767 2476
rect 10701 2396 10767 2412
rect 10701 2332 10702 2396
rect 10766 2332 10767 2396
rect 10701 2316 10767 2332
rect 10701 2252 10702 2316
rect 10766 2252 10767 2316
rect 10701 2236 10767 2252
rect 10701 2172 10702 2236
rect 10766 2172 10767 2236
rect 10701 2156 10767 2172
rect 10701 2092 10702 2156
rect 10766 2092 10767 2156
rect 10701 2076 10767 2092
rect 10701 2012 10702 2076
rect 10766 2012 10767 2076
rect 10701 1996 10767 2012
rect 10701 1932 10702 1996
rect 10766 1932 10767 1996
rect 10701 1778 10767 1932
rect 10827 1840 10887 2870
rect 10947 1778 11007 2810
rect 11067 1840 11127 2870
rect 11187 1778 11247 2810
rect 11307 2716 11373 2806
rect 11307 2652 11308 2716
rect 11372 2652 11373 2716
rect 11307 2636 11373 2652
rect 11307 2572 11308 2636
rect 11372 2572 11373 2636
rect 11307 2556 11373 2572
rect 11307 2492 11308 2556
rect 11372 2492 11373 2556
rect 11307 2476 11373 2492
rect 11307 2412 11308 2476
rect 11372 2412 11373 2476
rect 11307 2396 11373 2412
rect 11307 2332 11308 2396
rect 11372 2332 11373 2396
rect 11307 2316 11373 2332
rect 11307 2252 11308 2316
rect 11372 2252 11373 2316
rect 11307 2236 11373 2252
rect 11307 2172 11308 2236
rect 11372 2172 11373 2236
rect 11307 2156 11373 2172
rect 11307 2092 11308 2156
rect 11372 2092 11373 2156
rect 11307 2076 11373 2092
rect 11307 2012 11308 2076
rect 11372 2012 11373 2076
rect 11307 1996 11373 2012
rect 11307 1932 11308 1996
rect 11372 1932 11373 1996
rect 11307 1778 11373 1932
rect 11433 1778 11493 2810
rect 11553 1840 11613 2870
rect 11673 1778 11733 2810
rect 11793 1840 11853 2870
rect 11913 2716 11979 2806
rect 11913 2652 11914 2716
rect 11978 2652 11979 2716
rect 11913 2636 11979 2652
rect 11913 2572 11914 2636
rect 11978 2572 11979 2636
rect 11913 2556 11979 2572
rect 11913 2492 11914 2556
rect 11978 2492 11979 2556
rect 11913 2476 11979 2492
rect 11913 2412 11914 2476
rect 11978 2412 11979 2476
rect 11913 2396 11979 2412
rect 11913 2332 11914 2396
rect 11978 2332 11979 2396
rect 11913 2316 11979 2332
rect 11913 2252 11914 2316
rect 11978 2252 11979 2316
rect 11913 2236 11979 2252
rect 11913 2172 11914 2236
rect 11978 2172 11979 2236
rect 11913 2156 11979 2172
rect 11913 2092 11914 2156
rect 11978 2092 11979 2156
rect 11913 2076 11979 2092
rect 11913 2012 11914 2076
rect 11978 2012 11979 2076
rect 11913 1996 11979 2012
rect 11913 1932 11914 1996
rect 11978 1932 11979 1996
rect 11913 1778 11979 1932
rect 12039 1840 12099 2870
rect 12159 1778 12219 2810
rect 12279 1840 12339 2870
rect 12399 1778 12459 2810
rect 12519 2716 12585 2806
rect 12519 2652 12520 2716
rect 12584 2652 12585 2716
rect 12519 2636 12585 2652
rect 12519 2572 12520 2636
rect 12584 2572 12585 2636
rect 12519 2556 12585 2572
rect 12519 2492 12520 2556
rect 12584 2492 12585 2556
rect 12519 2476 12585 2492
rect 12519 2412 12520 2476
rect 12584 2412 12585 2476
rect 12519 2396 12585 2412
rect 12519 2332 12520 2396
rect 12584 2332 12585 2396
rect 12519 2316 12585 2332
rect 12519 2252 12520 2316
rect 12584 2252 12585 2316
rect 12519 2236 12585 2252
rect 12519 2172 12520 2236
rect 12584 2172 12585 2236
rect 12519 2156 12585 2172
rect 12519 2092 12520 2156
rect 12584 2092 12585 2156
rect 12519 2076 12585 2092
rect 12519 2012 12520 2076
rect 12584 2012 12585 2076
rect 12519 1996 12585 2012
rect 12519 1932 12520 1996
rect 12584 1932 12585 1996
rect 12519 1778 12585 1932
rect 12645 1778 12705 2810
rect 12765 1840 12825 2870
rect 12885 1778 12945 2810
rect 13005 1840 13065 2870
rect 13125 2716 13191 2806
rect 13125 2652 13126 2716
rect 13190 2652 13191 2716
rect 13125 2636 13191 2652
rect 13125 2572 13126 2636
rect 13190 2572 13191 2636
rect 13125 2556 13191 2572
rect 13125 2492 13126 2556
rect 13190 2492 13191 2556
rect 13125 2476 13191 2492
rect 13125 2412 13126 2476
rect 13190 2412 13191 2476
rect 13125 2396 13191 2412
rect 13125 2332 13126 2396
rect 13190 2332 13191 2396
rect 13125 2316 13191 2332
rect 13125 2252 13126 2316
rect 13190 2252 13191 2316
rect 13125 2236 13191 2252
rect 13125 2172 13126 2236
rect 13190 2172 13191 2236
rect 13125 2156 13191 2172
rect 13125 2092 13126 2156
rect 13190 2092 13191 2156
rect 13125 2076 13191 2092
rect 13125 2012 13126 2076
rect 13190 2012 13191 2076
rect 13125 1996 13191 2012
rect 13125 1932 13126 1996
rect 13190 1932 13191 1996
rect 13125 1778 13191 1932
rect 13251 1840 13311 2870
rect 13371 1778 13431 2810
rect 13491 1840 13551 2870
rect 13611 1778 13671 2810
rect 13731 2716 13797 2806
rect 13731 2652 13732 2716
rect 13796 2652 13797 2716
rect 13731 2636 13797 2652
rect 13731 2572 13732 2636
rect 13796 2572 13797 2636
rect 13731 2556 13797 2572
rect 13731 2492 13732 2556
rect 13796 2492 13797 2556
rect 13731 2476 13797 2492
rect 13731 2412 13732 2476
rect 13796 2412 13797 2476
rect 13731 2396 13797 2412
rect 13731 2332 13732 2396
rect 13796 2332 13797 2396
rect 13731 2316 13797 2332
rect 13731 2252 13732 2316
rect 13796 2252 13797 2316
rect 13731 2236 13797 2252
rect 13731 2172 13732 2236
rect 13796 2172 13797 2236
rect 13731 2156 13797 2172
rect 13731 2092 13732 2156
rect 13796 2092 13797 2156
rect 13731 2076 13797 2092
rect 13731 2012 13732 2076
rect 13796 2012 13797 2076
rect 13731 1996 13797 2012
rect 13731 1932 13732 1996
rect 13796 1932 13797 1996
rect 13731 1778 13797 1932
rect 13857 1778 13917 2810
rect 13977 1840 14037 2870
rect 14097 1778 14157 2810
rect 14217 1840 14277 2870
rect 14337 2716 14403 2806
rect 14337 2652 14338 2716
rect 14402 2652 14403 2716
rect 14337 2636 14403 2652
rect 14337 2572 14338 2636
rect 14402 2572 14403 2636
rect 14337 2556 14403 2572
rect 14337 2492 14338 2556
rect 14402 2492 14403 2556
rect 14337 2476 14403 2492
rect 14337 2412 14338 2476
rect 14402 2412 14403 2476
rect 14337 2396 14403 2412
rect 14337 2332 14338 2396
rect 14402 2332 14403 2396
rect 14337 2316 14403 2332
rect 14337 2252 14338 2316
rect 14402 2252 14403 2316
rect 14337 2236 14403 2252
rect 14337 2172 14338 2236
rect 14402 2172 14403 2236
rect 14337 2156 14403 2172
rect 14337 2092 14338 2156
rect 14402 2092 14403 2156
rect 14337 2076 14403 2092
rect 14337 2012 14338 2076
rect 14402 2012 14403 2076
rect 14337 1996 14403 2012
rect 14337 1932 14338 1996
rect 14402 1932 14403 1996
rect 14337 1778 14403 1932
rect 14463 1840 14523 2870
rect 14583 1778 14643 2810
rect 14703 1840 14763 2870
rect 14823 1778 14883 2810
rect 14943 2716 15009 2806
rect 14943 2652 14944 2716
rect 15008 2652 15009 2716
rect 14943 2636 15009 2652
rect 14943 2572 14944 2636
rect 15008 2572 15009 2636
rect 14943 2556 15009 2572
rect 14943 2492 14944 2556
rect 15008 2492 15009 2556
rect 14943 2476 15009 2492
rect 14943 2412 14944 2476
rect 15008 2412 15009 2476
rect 14943 2396 15009 2412
rect 14943 2332 14944 2396
rect 15008 2332 15009 2396
rect 14943 2316 15009 2332
rect 14943 2252 14944 2316
rect 15008 2252 15009 2316
rect 14943 2236 15009 2252
rect 14943 2172 14944 2236
rect 15008 2172 15009 2236
rect 14943 2156 15009 2172
rect 14943 2092 14944 2156
rect 15008 2092 15009 2156
rect 14943 2076 15009 2092
rect 14943 2012 14944 2076
rect 15008 2012 15009 2076
rect 14943 1996 15009 2012
rect 14943 1932 14944 1996
rect 15008 1932 15009 1996
rect 14943 1778 15009 1932
rect 15069 1778 15129 2810
rect 15189 1840 15249 2870
rect 15309 1778 15369 2810
rect 15429 1840 15489 2870
rect 15675 2817 15785 2870
rect 15849 2817 15993 2881
rect 15549 2716 15615 2806
rect 15549 2652 15550 2716
rect 15614 2652 15615 2716
rect 15549 2636 15615 2652
rect 15549 2572 15550 2636
rect 15614 2572 15615 2636
rect 15549 2556 15615 2572
rect 15549 2492 15550 2556
rect 15614 2492 15615 2556
rect 15549 2476 15615 2492
rect 15549 2412 15550 2476
rect 15614 2412 15615 2476
rect 15549 2396 15615 2412
rect 15549 2332 15550 2396
rect 15614 2332 15615 2396
rect 15549 2316 15615 2332
rect 15549 2252 15550 2316
rect 15614 2252 15615 2316
rect 15549 2236 15615 2252
rect 15549 2172 15550 2236
rect 15614 2172 15615 2236
rect 15549 2156 15615 2172
rect 15549 2092 15550 2156
rect 15614 2092 15615 2156
rect 15549 2076 15615 2092
rect 15549 2012 15550 2076
rect 15614 2012 15615 2076
rect 15549 1996 15615 2012
rect 15549 1932 15550 1996
rect 15614 1932 15615 1996
rect 15675 2737 15993 2817
rect 15675 2673 15790 2737
rect 15854 2673 15993 2737
rect 15675 2585 15993 2673
rect 15675 2521 15791 2585
rect 15855 2521 15993 2585
rect 15675 2415 15993 2521
rect 15675 2351 15791 2415
rect 15855 2351 15993 2415
rect 15675 2258 15993 2351
rect 15675 2194 15790 2258
rect 15854 2194 15993 2258
rect 15675 2016 15993 2194
rect 15675 1952 15708 2016
rect 15772 1952 15993 2016
rect 15675 1940 15993 1952
rect 15549 1778 15615 1932
rect 10701 1776 15615 1778
rect 10701 1712 10805 1776
rect 10869 1712 10885 1776
rect 10949 1712 10965 1776
rect 11029 1712 11045 1776
rect 11109 1712 11125 1776
rect 11189 1712 11205 1776
rect 11269 1712 11411 1776
rect 11475 1712 11491 1776
rect 11555 1712 11571 1776
rect 11635 1712 11651 1776
rect 11715 1712 11731 1776
rect 11795 1712 11811 1776
rect 11875 1712 12017 1776
rect 12081 1712 12097 1776
rect 12161 1712 12177 1776
rect 12241 1712 12257 1776
rect 12321 1712 12337 1776
rect 12401 1712 12417 1776
rect 12481 1712 12623 1776
rect 12687 1712 12703 1776
rect 12767 1712 12783 1776
rect 12847 1712 12863 1776
rect 12927 1712 12943 1776
rect 13007 1712 13023 1776
rect 13087 1712 13229 1776
rect 13293 1712 13309 1776
rect 13373 1712 13389 1776
rect 13453 1712 13469 1776
rect 13533 1712 13549 1776
rect 13613 1712 13629 1776
rect 13693 1712 13835 1776
rect 13899 1712 13915 1776
rect 13979 1712 13995 1776
rect 14059 1712 14075 1776
rect 14139 1712 14155 1776
rect 14219 1712 14235 1776
rect 14299 1712 14441 1776
rect 14505 1712 14521 1776
rect 14585 1712 14601 1776
rect 14665 1712 14681 1776
rect 14745 1712 14761 1776
rect 14825 1712 14841 1776
rect 14905 1712 15047 1776
rect 15111 1712 15127 1776
rect 15191 1712 15207 1776
rect 15271 1712 15287 1776
rect 15351 1712 15367 1776
rect 15431 1712 15447 1776
rect 15511 1712 15615 1776
rect 10701 1710 15615 1712
rect 15675 1755 15873 1765
rect 15675 1691 15796 1755
rect 15860 1691 15873 1755
rect 15675 1681 15873 1691
rect 10320 1528 10992 1530
rect 10320 1464 10424 1528
rect 10488 1464 10504 1528
rect 10568 1464 10584 1528
rect 10648 1464 10664 1528
rect 10728 1464 10744 1528
rect 10808 1464 10824 1528
rect 10888 1464 10992 1528
rect 10320 1462 10992 1464
rect 10320 1308 10386 1462
rect 10320 1244 10321 1308
rect 10385 1244 10386 1308
rect 10320 1228 10386 1244
rect 10320 1164 10321 1228
rect 10385 1164 10386 1228
rect 10320 1148 10386 1164
rect 10320 1084 10321 1148
rect 10385 1084 10386 1148
rect 10320 1068 10386 1084
rect 10320 1004 10321 1068
rect 10385 1004 10386 1068
rect 10320 988 10386 1004
rect 10320 924 10321 988
rect 10385 924 10386 988
rect 10320 908 10386 924
rect 10320 844 10321 908
rect 10385 844 10386 908
rect 10320 828 10386 844
rect 10320 764 10321 828
rect 10385 764 10386 828
rect 10320 748 10386 764
rect 10320 684 10321 748
rect 10385 684 10386 748
rect 10320 668 10386 684
rect 10320 604 10321 668
rect 10385 604 10386 668
rect 10320 588 10386 604
rect 10320 524 10321 588
rect 10385 524 10386 588
rect 10320 434 10386 524
rect 9932 369 10057 375
rect 10446 370 10506 1400
rect 10566 430 10626 1462
rect 10686 370 10746 1400
rect 10806 430 10866 1462
rect 10926 1308 10992 1462
rect 10926 1244 10927 1308
rect 10991 1244 10992 1308
rect 10926 1228 10992 1244
rect 10926 1164 10927 1228
rect 10991 1164 10992 1228
rect 10926 1148 10992 1164
rect 10926 1084 10927 1148
rect 10991 1084 10992 1148
rect 10926 1068 10992 1084
rect 10926 1004 10927 1068
rect 10991 1004 10992 1068
rect 10926 988 10992 1004
rect 10926 924 10927 988
rect 10991 924 10992 988
rect 10926 908 10992 924
rect 10926 844 10927 908
rect 10991 844 10992 908
rect 10926 828 10992 844
rect 10926 764 10927 828
rect 10991 764 10992 828
rect 10926 748 10992 764
rect 10926 684 10927 748
rect 10991 684 10992 748
rect 10926 668 10992 684
rect 10926 604 10927 668
rect 10991 604 10992 668
rect 10926 588 10992 604
rect 10926 524 10927 588
rect 10991 524 10992 588
rect 10926 434 10992 524
rect 11052 1528 13542 1530
rect 11052 1464 11156 1528
rect 11220 1464 11236 1528
rect 11300 1464 11316 1528
rect 11380 1464 11396 1528
rect 11460 1464 11476 1528
rect 11540 1464 11556 1528
rect 11620 1464 11762 1528
rect 11826 1464 11842 1528
rect 11906 1464 11922 1528
rect 11986 1464 12002 1528
rect 12066 1464 12082 1528
rect 12146 1464 12162 1528
rect 12226 1464 12368 1528
rect 12432 1464 12448 1528
rect 12512 1464 12528 1528
rect 12592 1464 12608 1528
rect 12672 1464 12688 1528
rect 12752 1464 12768 1528
rect 12832 1464 12974 1528
rect 13038 1464 13054 1528
rect 13118 1464 13134 1528
rect 13198 1464 13214 1528
rect 13278 1464 13294 1528
rect 13358 1464 13374 1528
rect 13438 1464 13542 1528
rect 11052 1462 13542 1464
rect 11052 1308 11118 1462
rect 11052 1244 11053 1308
rect 11117 1244 11118 1308
rect 11052 1228 11118 1244
rect 11052 1164 11053 1228
rect 11117 1164 11118 1228
rect 11052 1148 11118 1164
rect 11052 1084 11053 1148
rect 11117 1084 11118 1148
rect 11052 1068 11118 1084
rect 11052 1004 11053 1068
rect 11117 1004 11118 1068
rect 11052 988 11118 1004
rect 11052 924 11053 988
rect 11117 924 11118 988
rect 11052 908 11118 924
rect 11052 844 11053 908
rect 11117 844 11118 908
rect 11052 828 11118 844
rect 11052 764 11053 828
rect 11117 764 11118 828
rect 11052 748 11118 764
rect 11052 684 11053 748
rect 11117 684 11118 748
rect 11052 668 11118 684
rect 11052 604 11053 668
rect 11117 604 11118 668
rect 11052 588 11118 604
rect 11052 524 11053 588
rect 11117 524 11118 588
rect 11052 434 11118 524
rect 11178 370 11238 1400
rect 11298 430 11358 1462
rect 11418 370 11478 1400
rect 11538 430 11598 1462
rect 11658 1308 11724 1462
rect 11658 1244 11659 1308
rect 11723 1244 11724 1308
rect 11658 1228 11724 1244
rect 11658 1164 11659 1228
rect 11723 1164 11724 1228
rect 11658 1148 11724 1164
rect 11658 1084 11659 1148
rect 11723 1084 11724 1148
rect 11658 1068 11724 1084
rect 11658 1004 11659 1068
rect 11723 1004 11724 1068
rect 11658 988 11724 1004
rect 11658 924 11659 988
rect 11723 924 11724 988
rect 11658 908 11724 924
rect 11658 844 11659 908
rect 11723 844 11724 908
rect 11658 828 11724 844
rect 11658 764 11659 828
rect 11723 764 11724 828
rect 11658 748 11724 764
rect 11658 684 11659 748
rect 11723 684 11724 748
rect 11658 668 11724 684
rect 11658 604 11659 668
rect 11723 604 11724 668
rect 11658 588 11724 604
rect 11658 524 11659 588
rect 11723 524 11724 588
rect 11658 434 11724 524
rect 11784 430 11844 1462
rect 11904 370 11964 1400
rect 12024 430 12084 1462
rect 12144 370 12204 1400
rect 12264 1308 12330 1462
rect 12264 1244 12265 1308
rect 12329 1244 12330 1308
rect 12264 1228 12330 1244
rect 12264 1164 12265 1228
rect 12329 1164 12330 1228
rect 12264 1148 12330 1164
rect 12264 1084 12265 1148
rect 12329 1084 12330 1148
rect 12264 1068 12330 1084
rect 12264 1004 12265 1068
rect 12329 1004 12330 1068
rect 12264 988 12330 1004
rect 12264 924 12265 988
rect 12329 924 12330 988
rect 12264 908 12330 924
rect 12264 844 12265 908
rect 12329 844 12330 908
rect 12264 828 12330 844
rect 12264 764 12265 828
rect 12329 764 12330 828
rect 12264 748 12330 764
rect 12264 684 12265 748
rect 12329 684 12330 748
rect 12264 668 12330 684
rect 12264 604 12265 668
rect 12329 604 12330 668
rect 12264 588 12330 604
rect 12264 524 12265 588
rect 12329 524 12330 588
rect 12264 434 12330 524
rect 12390 370 12450 1400
rect 12510 430 12570 1462
rect 12630 370 12690 1400
rect 12750 430 12810 1462
rect 12870 1308 12936 1462
rect 12870 1244 12871 1308
rect 12935 1244 12936 1308
rect 12870 1228 12936 1244
rect 12870 1164 12871 1228
rect 12935 1164 12936 1228
rect 12870 1148 12936 1164
rect 12870 1084 12871 1148
rect 12935 1084 12936 1148
rect 12870 1068 12936 1084
rect 12870 1004 12871 1068
rect 12935 1004 12936 1068
rect 12870 988 12936 1004
rect 12870 924 12871 988
rect 12935 924 12936 988
rect 12870 908 12936 924
rect 12870 844 12871 908
rect 12935 844 12936 908
rect 12870 828 12936 844
rect 12870 764 12871 828
rect 12935 764 12936 828
rect 12870 748 12936 764
rect 12870 684 12871 748
rect 12935 684 12936 748
rect 12870 668 12936 684
rect 12870 604 12871 668
rect 12935 604 12936 668
rect 12870 588 12936 604
rect 12870 524 12871 588
rect 12935 524 12936 588
rect 12870 434 12936 524
rect 12996 430 13056 1462
rect 13116 370 13176 1400
rect 13236 430 13296 1462
rect 13356 370 13416 1400
rect 13476 1308 13542 1462
rect 13476 1244 13477 1308
rect 13541 1244 13542 1308
rect 13476 1228 13542 1244
rect 13476 1164 13477 1228
rect 13541 1164 13542 1228
rect 13476 1148 13542 1164
rect 13476 1084 13477 1148
rect 13541 1084 13542 1148
rect 13476 1068 13542 1084
rect 13476 1004 13477 1068
rect 13541 1004 13542 1068
rect 13476 988 13542 1004
rect 13476 924 13477 988
rect 13541 924 13542 988
rect 13476 908 13542 924
rect 13476 844 13477 908
rect 13541 844 13542 908
rect 13476 828 13542 844
rect 13476 764 13477 828
rect 13541 764 13542 828
rect 13476 748 13542 764
rect 13476 684 13477 748
rect 13541 684 13542 748
rect 13476 668 13542 684
rect 13476 604 13477 668
rect 13541 604 13542 668
rect 13476 588 13542 604
rect 13476 524 13477 588
rect 13541 524 13542 588
rect 13476 434 13542 524
rect 13602 1528 14880 1530
rect 13602 1464 13706 1528
rect 13770 1464 13786 1528
rect 13850 1464 13866 1528
rect 13930 1464 13946 1528
rect 14010 1464 14026 1528
rect 14090 1464 14106 1528
rect 14170 1464 14312 1528
rect 14376 1464 14392 1528
rect 14456 1464 14472 1528
rect 14536 1464 14552 1528
rect 14616 1464 14632 1528
rect 14696 1464 14712 1528
rect 14776 1464 14880 1528
rect 13602 1462 14880 1464
rect 13602 1308 13668 1462
rect 13602 1244 13603 1308
rect 13667 1244 13668 1308
rect 13602 1228 13668 1244
rect 13602 1164 13603 1228
rect 13667 1164 13668 1228
rect 13602 1148 13668 1164
rect 13602 1084 13603 1148
rect 13667 1084 13668 1148
rect 13602 1068 13668 1084
rect 13602 1004 13603 1068
rect 13667 1004 13668 1068
rect 13602 988 13668 1004
rect 13602 924 13603 988
rect 13667 924 13668 988
rect 13602 908 13668 924
rect 13602 844 13603 908
rect 13667 844 13668 908
rect 13602 828 13668 844
rect 13602 764 13603 828
rect 13667 764 13668 828
rect 13602 748 13668 764
rect 13602 684 13603 748
rect 13667 684 13668 748
rect 13602 668 13668 684
rect 13602 604 13603 668
rect 13667 604 13668 668
rect 13602 588 13668 604
rect 13602 524 13603 588
rect 13667 524 13668 588
rect 13602 434 13668 524
rect 13728 370 13788 1400
rect 13848 430 13908 1462
rect 13968 370 14028 1400
rect 14088 430 14148 1462
rect 14208 1308 14274 1462
rect 14208 1244 14209 1308
rect 14273 1244 14274 1308
rect 14208 1228 14274 1244
rect 14208 1164 14209 1228
rect 14273 1164 14274 1228
rect 14208 1148 14274 1164
rect 14208 1084 14209 1148
rect 14273 1084 14274 1148
rect 14208 1068 14274 1084
rect 14208 1004 14209 1068
rect 14273 1004 14274 1068
rect 14208 988 14274 1004
rect 14208 924 14209 988
rect 14273 924 14274 988
rect 14208 908 14274 924
rect 14208 844 14209 908
rect 14273 844 14274 908
rect 14208 828 14274 844
rect 14208 764 14209 828
rect 14273 764 14274 828
rect 14208 748 14274 764
rect 14208 684 14209 748
rect 14273 684 14274 748
rect 14208 668 14274 684
rect 14208 604 14209 668
rect 14273 604 14274 668
rect 14208 588 14274 604
rect 14208 524 14209 588
rect 14273 524 14274 588
rect 14208 434 14274 524
rect 14334 430 14394 1462
rect 14454 370 14514 1400
rect 14574 430 14634 1462
rect 14694 370 14754 1400
rect 14814 1308 14880 1462
rect 14814 1244 14815 1308
rect 14879 1244 14880 1308
rect 14814 1228 14880 1244
rect 14814 1164 14815 1228
rect 14879 1164 14880 1228
rect 14814 1148 14880 1164
rect 14814 1084 14815 1148
rect 14879 1084 14880 1148
rect 14814 1068 14880 1084
rect 14814 1004 14815 1068
rect 14879 1004 14880 1068
rect 14814 988 14880 1004
rect 14814 924 14815 988
rect 14879 924 14880 988
rect 14814 908 14880 924
rect 14814 844 14815 908
rect 14879 844 14880 908
rect 14814 828 14880 844
rect 14814 764 14815 828
rect 14879 764 14880 828
rect 14814 748 14880 764
rect 14814 684 14815 748
rect 14879 684 14880 748
rect 14814 668 14880 684
rect 14814 604 14815 668
rect 14879 604 14880 668
rect 14814 588 14880 604
rect 14814 524 14815 588
rect 14879 524 14880 588
rect 14814 434 14880 524
rect 14942 1528 15614 1530
rect 14942 1464 15046 1528
rect 15110 1464 15126 1528
rect 15190 1464 15206 1528
rect 15270 1464 15286 1528
rect 15350 1464 15366 1528
rect 15430 1464 15446 1528
rect 15510 1464 15614 1528
rect 14942 1462 15614 1464
rect 14942 1308 15008 1462
rect 14942 1244 14943 1308
rect 15007 1244 15008 1308
rect 14942 1228 15008 1244
rect 14942 1164 14943 1228
rect 15007 1164 15008 1228
rect 14942 1148 15008 1164
rect 14942 1084 14943 1148
rect 15007 1084 15008 1148
rect 14942 1068 15008 1084
rect 14942 1004 14943 1068
rect 15007 1004 15008 1068
rect 14942 988 15008 1004
rect 14942 924 14943 988
rect 15007 924 15008 988
rect 14942 908 15008 924
rect 14942 844 14943 908
rect 15007 844 15008 908
rect 14942 828 15008 844
rect 14942 764 14943 828
rect 15007 764 15008 828
rect 14942 748 15008 764
rect 14942 684 14943 748
rect 15007 684 15008 748
rect 14942 668 15008 684
rect 14942 604 14943 668
rect 15007 604 15008 668
rect 14942 588 15008 604
rect 14942 524 14943 588
rect 15007 524 15008 588
rect 14942 434 15008 524
rect 15068 430 15128 1462
rect 15188 370 15248 1400
rect 15308 430 15368 1462
rect 15428 370 15488 1400
rect 15548 1308 15614 1462
rect 15548 1244 15549 1308
rect 15613 1244 15614 1308
rect 15548 1228 15614 1244
rect 15548 1164 15549 1228
rect 15613 1164 15614 1228
rect 15548 1148 15614 1164
rect 15548 1084 15549 1148
rect 15613 1084 15614 1148
rect 15548 1068 15614 1084
rect 15548 1004 15549 1068
rect 15613 1004 15614 1068
rect 15548 988 15614 1004
rect 15548 924 15549 988
rect 15613 924 15614 988
rect 15548 908 15614 924
rect 15548 844 15549 908
rect 15613 844 15614 908
rect 15548 828 15614 844
rect 15548 764 15549 828
rect 15613 764 15614 828
rect 15548 748 15614 764
rect 15548 684 15549 748
rect 15613 684 15614 748
rect 15548 668 15614 684
rect 15548 604 15549 668
rect 15613 604 15614 668
rect 15548 588 15614 604
rect 15548 524 15549 588
rect 15613 524 15614 588
rect 15548 434 15614 524
rect 15675 1300 15735 1681
rect 15933 1562 15993 1940
rect 15795 1552 15993 1562
rect 15795 1488 15796 1552
rect 15860 1488 15993 1552
rect 15795 1478 15993 1488
rect 15675 1290 15993 1300
rect 15675 1226 15705 1290
rect 15769 1226 15993 1290
rect 10320 369 10992 370
rect 11052 369 13542 370
rect 13602 369 14880 370
rect 14942 369 15614 370
rect 15675 369 15993 1226
rect 9372 368 15993 369
rect 9372 365 10504 368
rect 9372 301 9962 365
rect 10026 304 10504 365
rect 10568 304 10584 368
rect 10648 304 10664 368
rect 10728 304 10744 368
rect 10808 304 11236 368
rect 11300 304 11316 368
rect 11380 304 11396 368
rect 11460 304 11476 368
rect 11540 304 11842 368
rect 11906 304 11922 368
rect 11986 304 12002 368
rect 12066 304 12082 368
rect 12146 304 12448 368
rect 12512 304 12528 368
rect 12592 304 12608 368
rect 12672 304 12688 368
rect 12752 304 13054 368
rect 13118 304 13134 368
rect 13198 304 13214 368
rect 13278 304 13294 368
rect 13358 304 13786 368
rect 13850 304 13866 368
rect 13930 304 13946 368
rect 14010 304 14026 368
rect 14090 304 14392 368
rect 14456 304 14472 368
rect 14536 304 14552 368
rect 14616 304 14632 368
rect 14696 304 15126 368
rect 15190 304 15206 368
rect 15270 304 15286 368
rect 15350 304 15366 368
rect 15430 304 15993 368
rect 10026 301 15993 304
rect 9372 291 15993 301
<< labels >>
flabel metal1 9275 1596 9943 1643 0 FreeSans 320 0 0 0 IN
port 1 nsew
flabel metal1 15751 1594 15933 1640 0 FreeSans 320 0 0 0 OUT
port 2 nsew
flabel metal1 9238 1979 9376 2013 0 FreeSans 320 0 0 0 code[3]
port 5 nsew
flabel metal1 14153 268 14211 1445 0 FreeSans 320 0 0 0 code[1]
port 8 nsew
flabel metal1 11727 268 11785 1445 0 FreeSans 320 0 0 0 code[2]
port 10 nsew
flabel metal4 9344 2338 9762 2948 0 FreeSans 320 0 0 0 VDD
port 17 nsew
flabel metal4 9372 291 9748 1728 0 FreeSans 320 0 0 0 VSS
port 19 nsew
flabel metal2 9702 1394 10138 1440 0 FreeSans 320 0 0 0 code_offset
port 21 nsew
flabel metal1 15009 267 15068 1448 0 FreeSans 320 0 0 0 code[0]
port 22 nsew
flabel metal1 10120 1896 10696 1943 0 FreeSans 320 0 0 0 code[0]
port 23 nsew
flabel locali 9464 2049 9498 2083 0 FreeSans 340 0 0 0 x1.Y
flabel locali 9464 1981 9498 2015 0 FreeSans 340 0 0 0 x1.Y
flabel locali 9372 1981 9406 2015 0 FreeSans 340 0 0 0 x1.A
flabel metal1 9329 1743 9363 1777 0 FreeSans 200 0 0 0 x1.VGND
flabel metal1 9329 2287 9363 2321 0 FreeSans 200 0 0 0 x1.VPWR
rlabel comment 9300 1760 9300 1760 4 x1.inv_1
rlabel metal1 9300 1712 9576 1808 1 x1.VGND
rlabel metal1 9300 2256 9576 2352 1 x1.VPWR
flabel pwell 9329 1743 9363 1777 0 FreeSans 200 0 0 0 x1.VNB
flabel nwell 9329 2287 9363 2321 0 FreeSans 200 0 0 0 x1.VPB
flabel locali 9562 2049 9596 2083 0 FreeSans 340 0 0 0 x5.Y
flabel locali 9562 1981 9596 2015 0 FreeSans 340 0 0 0 x5.Y
flabel locali 9654 1981 9688 2015 0 FreeSans 340 0 0 0 x5.A
flabel metal1 9697 1743 9731 1777 0 FreeSans 200 0 0 0 x5.VGND
flabel metal1 9697 2287 9731 2321 0 FreeSans 200 0 0 0 x5.VPWR
rlabel comment 9760 1760 9760 1760 6 x5.inv_1
rlabel metal1 9484 1712 9760 1808 1 x5.VGND
rlabel metal1 9484 2256 9760 2352 1 x5.VPWR
flabel pwell 9697 1743 9731 1777 0 FreeSans 200 0 0 0 x5.VNB
flabel nwell 9697 2287 9731 2321 0 FreeSans 200 0 0 0 x5.VPB
flabel metal1 9886 2049 9920 2083 0 FreeSans 320 0 0 0 x8.input_stack
flabel space 9930 2832 9964 2892 0 FreeSans 320 0 0 0 x8.vdd
flabel space 9930 2142 9964 2202 0 FreeSans 320 0 0 0 x8.output_stack
flabel poly 9863 1392 9965 1422 0 FreeSans 320 0 0 0 x9.input_stack
flabel space 9977 1305 10011 1365 0 FreeSans 320 0 0 0 x9.output_stack
flabel space 9977 339 10011 399 0 FreeSans 320 0 0 0 x9.vss
flabel metal1 10528 1809 10562 1843 0 FreeSans 320 0 0 0 x6.SW
flabel pdiff 10560 1678 10618 1762 0 FreeSans 320 0 0 0 x6.delay_signal
flabel metal4 9972 2871 10642 2939 0 FreeSans 320 0 0 0 x6.CTOP
flabel metal1 10881 1405 10915 1439 0 FreeSans 320 0 0 0 x7.SW
flabel ndiff 10913 1477 10971 1561 0 FreeSans 320 0 0 0 x7.delay_signal
flabel metal4 10320 300 10992 368 0 FreeSans 320 0 0 0 x7.CTOP
flabel metal1 11386 1809 11420 1843 0 FreeSans 320 0 0 0 x5[6].SW
flabel pdiff 11330 1678 11388 1762 0 FreeSans 320 0 0 0 x5[6].delay_signal
flabel metal4 11306 2871 11976 2939 0 FreeSans 320 0 0 0 x5[6].CTOP
flabel metal1 11260 1809 11294 1843 0 FreeSans 320 0 0 0 x5[7].SW
flabel pdiff 11292 1678 11350 1762 0 FreeSans 320 0 0 0 x5[7].delay_signal
flabel metal4 10704 2871 11374 2939 0 FreeSans 320 0 0 0 x5[7].CTOP
flabel metal1 11613 1405 11647 1439 0 FreeSans 320 0 0 0 x4[3].SW
flabel ndiff 11645 1477 11703 1561 0 FreeSans 320 0 0 0 x4[3].delay_signal
flabel metal4 11052 300 11724 368 0 FreeSans 320 0 0 0 x4[3].CTOP
flabel metal1 12472 1809 12506 1843 0 FreeSans 320 0 0 0 x5[5].SW
flabel pdiff 12504 1678 12562 1762 0 FreeSans 320 0 0 0 x5[5].delay_signal
flabel metal4 11916 2871 12586 2939 0 FreeSans 320 0 0 0 x5[5].CTOP
flabel metal1 11735 1405 11769 1439 0 FreeSans 320 0 0 0 x4[2].SW
flabel ndiff 11679 1477 11737 1561 0 FreeSans 320 0 0 0 x4[2].delay_signal
flabel metal4 11658 300 12330 368 0 FreeSans 320 0 0 0 x4[2].CTOP
flabel metal1 12598 1809 12632 1843 0 FreeSans 320 0 0 0 x5[4].SW
flabel pdiff 12542 1678 12600 1762 0 FreeSans 320 0 0 0 x5[4].delay_signal
flabel metal4 12518 2871 13188 2939 0 FreeSans 320 0 0 0 x5[4].CTOP
flabel metal1 12825 1405 12859 1439 0 FreeSans 320 0 0 0 x4[1].SW
flabel ndiff 12857 1477 12915 1561 0 FreeSans 320 0 0 0 x4[1].delay_signal
flabel metal4 12264 300 12936 368 0 FreeSans 320 0 0 0 x4[1].CTOP
flabel metal1 13684 1809 13718 1843 0 FreeSans 320 0 0 0 x5[3].SW
flabel pdiff 13716 1678 13774 1762 0 FreeSans 320 0 0 0 x5[3].delay_signal
flabel metal4 13128 2871 13798 2939 0 FreeSans 320 0 0 0 x5[3].CTOP
flabel metal1 12947 1405 12981 1439 0 FreeSans 320 0 0 0 x4[0].SW
flabel ndiff 12891 1477 12949 1561 0 FreeSans 320 0 0 0 x4[0].delay_signal
flabel metal4 12870 300 13542 368 0 FreeSans 320 0 0 0 x4[0].CTOP
flabel metal1 13810 1809 13844 1843 0 FreeSans 320 0 0 0 x5[2].SW
flabel pdiff 13754 1678 13812 1762 0 FreeSans 320 0 0 0 x5[2].delay_signal
flabel metal4 13730 2871 14400 2939 0 FreeSans 320 0 0 0 x5[2].CTOP
flabel metal1 14163 1405 14197 1439 0 FreeSans 320 0 0 0 x3[1].SW
flabel ndiff 14195 1477 14253 1561 0 FreeSans 320 0 0 0 x3[1].delay_signal
flabel metal4 13602 300 14274 368 0 FreeSans 320 0 0 0 x3[1].CTOP
flabel metal1 14896 1809 14930 1843 0 FreeSans 320 0 0 0 x5[1].SW
flabel pdiff 14928 1678 14986 1762 0 FreeSans 320 0 0 0 x5[1].delay_signal
flabel metal4 14340 2871 15010 2939 0 FreeSans 320 0 0 0 x5[1].CTOP
flabel metal1 14285 1405 14319 1439 0 FreeSans 320 0 0 0 x3[0].SW
flabel ndiff 14229 1477 14287 1561 0 FreeSans 320 0 0 0 x3[0].delay_signal
flabel metal4 14208 300 14880 368 0 FreeSans 320 0 0 0 x3[0].CTOP
flabel metal1 15022 1809 15056 1843 0 FreeSans 320 0 0 0 x5[0].SW
flabel pdiff 14966 1678 15024 1762 0 FreeSans 320 0 0 0 x5[0].delay_signal
flabel metal4 14942 2871 15612 2939 0 FreeSans 320 0 0 0 x5[0].CTOP
flabel metal1 15019 1405 15053 1439 0 FreeSans 320 0 0 0 x2.SW
flabel ndiff 14963 1477 15021 1561 0 FreeSans 320 0 0 0 x2.delay_signal
flabel metal4 14942 300 15614 368 0 FreeSans 320 0 0 0 x2.CTOP
<< end >>
