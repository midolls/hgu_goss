magic
tech sky130A
magscale 1 2
timestamp 1699320260
<< checkpaint >>
rect -944 2490 1998 2596
rect -944 -766 2736 2490
rect -206 -872 2736 -766
<< error_s >>
rect 316 1317 369 1336
rect 298 1300 369 1317
rect 316 1266 387 1300
rect 129 1215 187 1221
rect 129 1181 141 1215
rect 129 1175 187 1181
rect 129 1021 187 1027
rect 129 987 141 1021
rect 129 981 187 987
rect 129 913 187 919
rect 129 879 141 913
rect 129 873 187 879
rect 129 719 187 725
rect 129 685 141 719
rect 129 679 187 685
rect 316 583 386 1266
rect 668 1247 702 1265
rect 668 1211 738 1247
rect 498 1198 556 1204
rect 498 1164 510 1198
rect 685 1177 756 1211
rect 498 1158 556 1164
rect 498 986 556 992
rect 498 952 510 986
rect 498 946 556 952
rect 498 878 556 884
rect 498 844 510 878
rect 498 838 556 844
rect 498 666 556 672
rect 498 632 510 666
rect 498 626 556 632
rect 316 547 369 583
rect 685 530 755 1177
rect 867 1109 925 1115
rect 867 1075 879 1109
rect 867 1069 925 1075
rect 867 915 925 921
rect 867 881 879 915
rect 867 875 925 881
rect 867 807 925 813
rect 867 773 879 807
rect 867 767 925 773
rect 867 613 925 619
rect 867 579 879 613
rect 867 573 925 579
rect 685 494 738 530
use sky130_fd_pr__nfet_01v8_PTX3GD  XM1
timestamp 0
transform 1 0 158 0 1 950
box -211 -403 211 403
use sky130_fd_pr__nfet_01v8_PTX3GD  XM13
timestamp 0
transform 1 0 896 0 1 844
box -211 -403 211 403
use sky130_fd_pr__pfet_01v8_hvt_M47XPL  XM46
timestamp 0
transform 1 0 1265 0 1 809
box -211 -421 211 421
use sky130_fd_pr__pfet_01v8_hvt_M47XPL  XM48
timestamp 0
transform 1 0 527 0 1 915
box -211 -421 211 421
<< end >>
