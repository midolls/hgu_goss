* NGSPICE file created from hgu_sarlogic_8bit_logic.ext - technology: sky130A

.subckt sky130_fd_sc_hd__buf_1 A VGND VPWR X VNB VPB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_4 A VGND VPWR X VNB VPB
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_16 A VGND VPWR X VNB VPB
X0 VGND A a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 a_109_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 VPWR A a_109_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 a_109_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X17 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X18 VPWR A a_109_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 VGND A a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X21 VGND A a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X22 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X23 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X24 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X25 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X26 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X27 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X28 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X29 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X30 a_109_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X31 a_109_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X32 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X33 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X34 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X35 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X36 VPWR A a_109_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X37 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X38 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X39 a_109_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X40 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X41 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X42 a_109_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X43 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_2 A VGND VPWR X VNB VPB
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X2 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X3 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X4 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfbbp_1 CLK D RESET_B SET_B VGND VPWR Q Q_N VNB VPB
X0 a_788_47# a_942_21# a_648_21# VNB sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1 VPWR RESET_B a_942_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X2 VGND a_1429_21# a_1364_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X3 VPWR a_942_21# a_1663_329# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X4 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X6 VPWR a_1429_21# a_1341_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X7 a_474_413# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X8 a_1545_47# a_942_21# a_1429_21# VNB sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X9 VPWR a_1429_21# a_2136_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X10 a_582_47# a_193_47# a_474_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X11 a_1429_21# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X12 a_648_21# a_474_413# a_788_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X13 a_1341_413# a_193_47# a_1255_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X14 a_1663_329# a_1255_47# a_1429_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X15 a_1160_47# a_648_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X16 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X17 a_1255_47# a_27_47# a_1113_329# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X18 Q a_2136_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X19 a_648_21# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X20 a_788_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X21 Q_N a_1429_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X22 VGND RESET_B a_942_21# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X23 Q a_2136_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X24 VPWR a_942_21# a_892_329# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X25 a_558_413# a_27_47# a_474_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X26 VGND a_648_21# a_582_47# VNB sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X27 a_892_329# a_474_413# a_648_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X28 VGND a_1429_21# a_2136_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X29 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X30 a_474_413# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X31 a_1364_47# a_27_47# a_1255_47# VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X32 a_1255_47# a_193_47# a_1160_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X33 Q_N a_1429_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X34 a_1545_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X35 VPWR a_648_21# a_558_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X36 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X37 a_1113_329# a_648_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X38 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X39 a_1429_21# a_1255_47# a_1545_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
.ends

.subckt sky130_fd_sc_hd__mux4_4 A0 A1 A2 A3 S0 S1 VGND VPWR X VNB VPB
X0 X a_789_316# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X1 X a_789_316# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.154 ps=1.34 w=1 l=0.15
X2 VPWR A0 a_1280_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.105 ps=0.995 w=0.64 l=0.15
X3 a_873_316# a_601_345# a_789_316# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X4 a_601_345# S1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5 VPWR S0 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6 VGND a_789_316# X VNB sky130_fd_pr__nfet_01v8 ad=0.218 pd=1.97 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 VGND a_789_316# X VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 VPWR A3 a_373_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.164 ps=1.33 w=0.64 l=0.15
X9 a_1282_47# a_27_47# a_873_316# VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.072 ps=0.76 w=0.36 l=0.15
X10 a_1280_413# S0 a_873_316# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=0.995 as=0.0567 ps=0.69 w=0.42 l=0.15
X11 a_1065_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0786 pd=0.805 as=0.109 ps=1.36 w=0.42 l=0.15
X12 a_193_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X13 a_873_316# S0 a_1065_47# VNB sky130_fd_pr__nfet_01v8 ad=0.072 pd=0.76 as=0.0786 ps=0.805 w=0.36 l=0.15
X14 X a_789_316# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=1 w=0.65 l=0.15
X15 a_1061_369# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.16 as=0.166 ps=1.8 w=0.64 l=0.15
X16 a_873_316# a_27_47# a_1061_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.138 ps=1.16 w=0.42 l=0.15
X17 VPWR a_789_316# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.335 pd=2.67 as=0.135 ps=1.27 w=1 l=0.15
X18 X a_789_316# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.175 ps=1.35 w=1 l=0.15
X19 VGND A3 a_398_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0819 pd=0.81 as=0.0671 ps=0.75 w=0.42 l=0.15
X20 a_601_345# S1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.38 as=0.0819 ps=0.81 w=0.42 l=0.15
X21 a_873_316# S1 a_789_316# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.6 as=0.0729 ps=0.81 w=0.54 l=0.15
X22 a_193_369# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0974 pd=0.97 as=0.0864 ps=0.91 w=0.64 l=0.15
X23 a_789_316# a_601_345# a_288_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0729 pd=0.81 as=0.14 ps=1.6 w=0.54 l=0.15
X24 a_398_47# S0 a_288_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.072 ps=0.76 w=0.36 l=0.15
X25 VGND A0 a_1282_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=1 as=0.066 ps=0.745 w=0.42 l=0.15
X26 a_373_413# a_27_47# a_288_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.164 pd=1.33 as=0.0567 ps=0.69 w=0.42 l=0.15
X27 a_288_47# a_27_47# a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0.072 pd=0.76 as=0.066 ps=0.745 w=0.36 l=0.15
X28 VPWR a_789_316# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X29 a_288_47# S0 a_193_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0974 ps=0.97 w=0.42 l=0.15
X30 VGND S0 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X31 a_789_316# S1 a_288_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__inv_1 A VGND VPWR Y VNB VPB
X0 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
.ends

.subckt hgu_sarlogic_8bit_logic sel_bit[0] sel_bit[1] reset eob comparator_out D[7]
+ D[6] check[6] D[5] check[0] check[5] check[1] check[4] check[2] check[3] D[2] D[3]
+ D[1] D[4] D[0] clk_sar VSS VDD
Xx1 reset VSS VDD x3/A VSS VDD sky130_fd_sc_hd__buf_1
Xx2 clk_sar VSS VDD x5/A VSS VDD sky130_fd_sc_hd__buf_1
Xx3 x3/A VSS VDD x4/A VSS VDD sky130_fd_sc_hd__buf_4
Xx4 x4/A VSS VDD x4/X VSS VDD sky130_fd_sc_hd__buf_16
Xx5 x5/A VSS VDD x5/X VSS VDD sky130_fd_sc_hd__buf_2
Xx60 D[3] comparator_out x4/X x33/Q_N VSS VDD D[4] x60/Q_N VSS VDD sky130_fd_sc_hd__dfbbp_1
Xx72 x75/Q comparator_out x4/X x45/Q_N VSS VDD D[0] x72/Q_N VSS VDD sky130_fd_sc_hd__dfbbp_1
Xx51 D[6] comparator_out x4/X x20/Q_N VSS VDD D[7] x51/Q_N VSS VDD sky130_fd_sc_hd__dfbbp_1
Xx30 x5/X check[6] x4/X VDD VSS VDD check[5] x30/Q_N VSS VDD sky130_fd_sc_hd__dfbbp_1
Xx63 D[2] comparator_out x4/X x36/Q_N VSS VDD D[3] x63/Q_N VSS VDD sky130_fd_sc_hd__dfbbp_1
Xx20 x5/X eob VDD x4/X VSS VDD x27/D x20/Q_N VSS VDD sky130_fd_sc_hd__dfbbp_1
Xx42 x5/X check[2] x4/X VDD VSS VDD check[1] x42/Q_N VSS VDD sky130_fd_sc_hd__dfbbp_1
Xx75 VSS VSS x4/X x77/Y VSS VDD x75/Q x75/Q_N VSS VDD sky130_fd_sc_hd__dfbbp_1
Xsky130_fd_sc_hd__mux4_4_0 check[2] check[1] check[0] x48/Q sel_bit[0] sel_bit[1]
+ VSS VDD eob VSS VDD sky130_fd_sc_hd__mux4_4
Xx54 D[5] comparator_out x4/X x27/Q_N VSS VDD D[6] x54/Q_N VSS VDD sky130_fd_sc_hd__dfbbp_1
Xx33 x5/X check[5] x4/X VDD VSS VDD check[4] x33/Q_N VSS VDD sky130_fd_sc_hd__dfbbp_1
Xx66 D[1] comparator_out x4/X x39/Q_N VSS VDD D[2] x66/Q_N VSS VDD sky130_fd_sc_hd__dfbbp_1
Xx77 eob VSS VDD x77/Y VSS VDD sky130_fd_sc_hd__inv_1
Xx45 x5/X check[1] x4/X VDD VSS VDD check[0] x45/Q_N VSS VDD sky130_fd_sc_hd__dfbbp_1
Xx57 D[4] comparator_out x4/X x30/Q_N VSS VDD D[5] x57/Q_N VSS VDD sky130_fd_sc_hd__dfbbp_1
Xx36 x5/X check[4] x4/X VDD VSS VDD check[3] x36/Q_N VSS VDD sky130_fd_sc_hd__dfbbp_1
Xx48 x5/X check[0] x4/X VDD VSS VDD x48/Q x48/Q_N VSS VDD sky130_fd_sc_hd__dfbbp_1
Xx69 D[0] comparator_out x4/X x42/Q_N VSS VDD D[1] x69/Q_N VSS VDD sky130_fd_sc_hd__dfbbp_1
Xx27 x5/X x27/D x4/X VDD VSS VDD check[6] x27/Q_N VSS VDD sky130_fd_sc_hd__dfbbp_1
Xx39 x5/X check[3] x4/X VDD VSS VDD check[2] x39/Q_N VSS VDD sky130_fd_sc_hd__dfbbp_1
.ends

