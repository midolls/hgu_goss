magic
tech sky130A
magscale 1 2
timestamp 1698045514
<< checkpaint >>
rect -944 -766 1998 2360
<< error_s >>
rect 129 913 187 919
rect 129 879 141 913
rect 129 873 187 879
rect 129 719 187 725
rect 129 685 141 719
rect 129 679 187 685
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
use sky130_fd_pr__nfet_01v8_L7T3GD  XM1
timestamp 0
transform 1 0 158 0 1 799
box -211 -252 211 252
use sky130_fd_pr__pfet_01v8_MQX2PY  XM2
timestamp 0
transform 1 0 527 0 1 797
box -211 -303 211 303
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 IN
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 OUT
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 VSS
port 3 nsew
<< end >>
