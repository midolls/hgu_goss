magic
tech sky130A
magscale 1 2
timestamp 1699633464
<< nmos >>
rect -63 -275 -33 275
rect 33 -275 63 275
<< ndiff >>
rect -125 263 -63 275
rect -125 -263 -113 263
rect -79 -263 -63 263
rect -125 -275 -63 -263
rect -33 263 33 275
rect -33 -263 -17 263
rect 17 -263 33 263
rect -33 -275 33 -263
rect 63 263 125 275
rect 63 -263 79 263
rect 113 -263 125 263
rect 63 -275 125 -263
<< ndiffc >>
rect -113 -263 -79 263
rect -17 -263 17 263
rect 79 -263 113 263
<< psubdiff >>
rect -145 448 -121 482
rect -71 448 -25 482
rect 25 448 71 482
rect 121 448 227 482
rect 193 375 227 448
rect 193 -393 227 -331
rect -145 -427 -121 -393
rect -71 -427 -25 -393
rect 25 -427 71 -393
rect 121 -427 227 -393
<< psubdiffcont >>
rect -121 448 -71 482
rect -25 448 25 482
rect 71 448 121 482
rect 193 -331 227 375
rect -121 -427 -71 -393
rect -25 -427 25 -393
rect 71 -427 121 -393
<< poly >>
rect -63 275 -33 301
rect 33 275 63 301
rect -63 -301 -33 -275
rect 33 -301 63 -275
<< locali >>
rect -145 448 -121 482
rect -71 448 -25 482
rect 25 448 71 482
rect 121 448 227 482
rect 193 375 227 448
rect -113 263 -79 279
rect -113 -279 -79 -263
rect -17 263 17 279
rect -17 -279 17 -263
rect 79 263 113 279
rect 79 -279 113 -263
rect 193 -393 227 -331
rect -145 -427 -121 -393
rect -71 -427 -25 -393
rect 25 -427 71 -393
rect 121 -427 227 -393
<< viali >>
rect -113 -263 -79 263
rect -17 -263 17 263
rect 79 -263 113 263
<< metal1 >>
rect -119 263 -73 275
rect -119 -263 -113 263
rect -79 -263 -73 263
rect -119 -275 -73 -263
rect -23 263 23 275
rect -23 -263 -17 263
rect 17 -263 23 263
rect -23 -275 23 -263
rect 73 263 119 275
rect 73 -263 79 263
rect 113 -263 119 263
rect 73 -275 119 -263
<< properties >>
string FIXED_BBOX -210 -432 210 432
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2.75 l 0.15 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
