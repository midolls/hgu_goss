magic
tech sky130A
magscale 1 2
timestamp 1698619433
<< pwell >>
rect 1224 9352 1250 9384
rect 1830 9352 1856 9384
rect 2436 9352 2462 9384
rect 3042 9352 3068 9384
rect 3648 9352 3674 9384
rect 4254 9352 4280 9384
rect 4860 9352 4886 9384
rect 5466 9352 5492 9384
rect 3646 8848 3682 8882
rect 1224 8192 1250 8224
rect 1830 8192 1856 8224
rect 2436 8192 2462 8224
rect 3042 8192 3068 8224
rect 3648 8192 3674 8224
rect 4254 8192 4280 8224
rect 4860 8192 4886 8224
rect 5466 8192 5492 8224
<< metal3 >>
rect 904 10162 5818 10164
rect 904 10098 1008 10162
rect 1072 10098 1088 10162
rect 1152 10098 1168 10162
rect 1232 10098 1248 10162
rect 1312 10098 1328 10162
rect 1392 10098 1408 10162
rect 1472 10098 1614 10162
rect 1678 10098 1694 10162
rect 1758 10098 1774 10162
rect 1838 10098 1854 10162
rect 1918 10098 1934 10162
rect 1998 10098 2014 10162
rect 2078 10098 2220 10162
rect 2284 10098 2300 10162
rect 2364 10098 2380 10162
rect 2444 10098 2460 10162
rect 2524 10098 2540 10162
rect 2604 10098 2620 10162
rect 2684 10098 2826 10162
rect 2890 10098 2906 10162
rect 2970 10098 2986 10162
rect 3050 10098 3066 10162
rect 3130 10098 3146 10162
rect 3210 10098 3226 10162
rect 3290 10098 3432 10162
rect 3496 10098 3512 10162
rect 3576 10098 3592 10162
rect 3656 10098 3672 10162
rect 3736 10098 3752 10162
rect 3816 10098 3832 10162
rect 3896 10098 4038 10162
rect 4102 10098 4118 10162
rect 4182 10098 4198 10162
rect 4262 10098 4278 10162
rect 4342 10098 4358 10162
rect 4422 10098 4438 10162
rect 4502 10098 4644 10162
rect 4708 10098 4724 10162
rect 4788 10098 4804 10162
rect 4868 10098 4884 10162
rect 4948 10098 4964 10162
rect 5028 10098 5044 10162
rect 5108 10098 5250 10162
rect 5314 10098 5330 10162
rect 5394 10098 5410 10162
rect 5474 10098 5490 10162
rect 5554 10098 5570 10162
rect 5634 10098 5650 10162
rect 5714 10098 5818 10162
rect 904 10096 5818 10098
rect 904 9942 970 10096
rect 904 9878 905 9942
rect 969 9878 970 9942
rect 904 9862 970 9878
rect 904 9798 905 9862
rect 969 9798 970 9862
rect 904 9782 970 9798
rect 904 9718 905 9782
rect 969 9718 970 9782
rect 904 9702 970 9718
rect 904 9638 905 9702
rect 969 9638 970 9702
rect 904 9622 970 9638
rect 904 9558 905 9622
rect 969 9558 970 9622
rect 904 9542 970 9558
rect 904 9478 905 9542
rect 969 9478 970 9542
rect 904 9462 970 9478
rect 904 9398 905 9462
rect 969 9398 970 9462
rect 904 9382 970 9398
rect 904 9318 905 9382
rect 969 9318 970 9382
rect 904 9302 970 9318
rect 904 9238 905 9302
rect 969 9238 970 9302
rect 904 9222 970 9238
rect 904 9158 905 9222
rect 969 9158 970 9222
rect 904 9068 970 9158
rect 1030 9064 1090 10096
rect 1150 9004 1210 10034
rect 1270 9064 1330 10096
rect 1390 9004 1450 10034
rect 1510 9942 1576 10096
rect 1510 9878 1511 9942
rect 1575 9878 1576 9942
rect 1510 9862 1576 9878
rect 1510 9798 1511 9862
rect 1575 9798 1576 9862
rect 1510 9782 1576 9798
rect 1510 9718 1511 9782
rect 1575 9718 1576 9782
rect 1510 9702 1576 9718
rect 1510 9638 1511 9702
rect 1575 9638 1576 9702
rect 1510 9622 1576 9638
rect 1510 9558 1511 9622
rect 1575 9558 1576 9622
rect 1510 9542 1576 9558
rect 1510 9478 1511 9542
rect 1575 9478 1576 9542
rect 1510 9462 1576 9478
rect 1510 9398 1511 9462
rect 1575 9398 1576 9462
rect 1510 9382 1576 9398
rect 1510 9318 1511 9382
rect 1575 9318 1576 9382
rect 1510 9302 1576 9318
rect 1510 9238 1511 9302
rect 1575 9238 1576 9302
rect 1510 9222 1576 9238
rect 1510 9158 1511 9222
rect 1575 9158 1576 9222
rect 1510 9068 1576 9158
rect 1636 9064 1696 10096
rect 1756 9004 1816 10034
rect 1876 9064 1936 10096
rect 1996 9004 2056 10034
rect 2116 9942 2182 10096
rect 2116 9878 2117 9942
rect 2181 9878 2182 9942
rect 2116 9862 2182 9878
rect 2116 9798 2117 9862
rect 2181 9798 2182 9862
rect 2116 9782 2182 9798
rect 2116 9718 2117 9782
rect 2181 9718 2182 9782
rect 2116 9702 2182 9718
rect 2116 9638 2117 9702
rect 2181 9638 2182 9702
rect 2116 9622 2182 9638
rect 2116 9558 2117 9622
rect 2181 9558 2182 9622
rect 2116 9542 2182 9558
rect 2116 9478 2117 9542
rect 2181 9478 2182 9542
rect 2116 9462 2182 9478
rect 2116 9398 2117 9462
rect 2181 9398 2182 9462
rect 2116 9382 2182 9398
rect 2116 9318 2117 9382
rect 2181 9318 2182 9382
rect 2116 9302 2182 9318
rect 2116 9238 2117 9302
rect 2181 9238 2182 9302
rect 2116 9222 2182 9238
rect 2116 9158 2117 9222
rect 2181 9158 2182 9222
rect 2116 9068 2182 9158
rect 2242 9064 2302 10096
rect 2362 9004 2422 10034
rect 2482 9064 2542 10096
rect 2602 9004 2662 10034
rect 2722 9942 2788 10096
rect 2722 9878 2723 9942
rect 2787 9878 2788 9942
rect 2722 9862 2788 9878
rect 2722 9798 2723 9862
rect 2787 9798 2788 9862
rect 2722 9782 2788 9798
rect 2722 9718 2723 9782
rect 2787 9718 2788 9782
rect 2722 9702 2788 9718
rect 2722 9638 2723 9702
rect 2787 9638 2788 9702
rect 2722 9622 2788 9638
rect 2722 9558 2723 9622
rect 2787 9558 2788 9622
rect 2722 9542 2788 9558
rect 2722 9478 2723 9542
rect 2787 9478 2788 9542
rect 2722 9462 2788 9478
rect 2722 9398 2723 9462
rect 2787 9398 2788 9462
rect 2722 9382 2788 9398
rect 2722 9318 2723 9382
rect 2787 9318 2788 9382
rect 2722 9302 2788 9318
rect 2722 9238 2723 9302
rect 2787 9238 2788 9302
rect 2722 9222 2788 9238
rect 2722 9158 2723 9222
rect 2787 9158 2788 9222
rect 2722 9068 2788 9158
rect 2848 9064 2908 10096
rect 2968 9004 3028 10034
rect 3088 9064 3148 10096
rect 3208 9004 3268 10034
rect 3328 9942 3394 10096
rect 3328 9878 3329 9942
rect 3393 9878 3394 9942
rect 3328 9862 3394 9878
rect 3328 9798 3329 9862
rect 3393 9798 3394 9862
rect 3328 9782 3394 9798
rect 3328 9718 3329 9782
rect 3393 9718 3394 9782
rect 3328 9702 3394 9718
rect 3328 9638 3329 9702
rect 3393 9638 3394 9702
rect 3328 9622 3394 9638
rect 3328 9558 3329 9622
rect 3393 9558 3394 9622
rect 3328 9542 3394 9558
rect 3328 9478 3329 9542
rect 3393 9478 3394 9542
rect 3328 9462 3394 9478
rect 3328 9398 3329 9462
rect 3393 9398 3394 9462
rect 3328 9382 3394 9398
rect 3328 9318 3329 9382
rect 3393 9318 3394 9382
rect 3328 9302 3394 9318
rect 3328 9238 3329 9302
rect 3393 9238 3394 9302
rect 3328 9222 3394 9238
rect 3328 9158 3329 9222
rect 3393 9158 3394 9222
rect 3328 9068 3394 9158
rect 3454 9064 3514 10096
rect 3574 9004 3634 10034
rect 3694 9064 3754 10096
rect 3814 9004 3874 10034
rect 3934 9942 4000 10096
rect 3934 9878 3935 9942
rect 3999 9878 4000 9942
rect 3934 9862 4000 9878
rect 3934 9798 3935 9862
rect 3999 9798 4000 9862
rect 3934 9782 4000 9798
rect 3934 9718 3935 9782
rect 3999 9718 4000 9782
rect 3934 9702 4000 9718
rect 3934 9638 3935 9702
rect 3999 9638 4000 9702
rect 3934 9622 4000 9638
rect 3934 9558 3935 9622
rect 3999 9558 4000 9622
rect 3934 9542 4000 9558
rect 3934 9478 3935 9542
rect 3999 9478 4000 9542
rect 3934 9462 4000 9478
rect 3934 9398 3935 9462
rect 3999 9398 4000 9462
rect 3934 9382 4000 9398
rect 3934 9318 3935 9382
rect 3999 9318 4000 9382
rect 3934 9302 4000 9318
rect 3934 9238 3935 9302
rect 3999 9238 4000 9302
rect 3934 9222 4000 9238
rect 3934 9158 3935 9222
rect 3999 9158 4000 9222
rect 3934 9068 4000 9158
rect 4060 9064 4120 10096
rect 4180 9004 4240 10034
rect 4300 9064 4360 10096
rect 4420 9004 4480 10034
rect 4540 9942 4606 10096
rect 4540 9878 4541 9942
rect 4605 9878 4606 9942
rect 4540 9862 4606 9878
rect 4540 9798 4541 9862
rect 4605 9798 4606 9862
rect 4540 9782 4606 9798
rect 4540 9718 4541 9782
rect 4605 9718 4606 9782
rect 4540 9702 4606 9718
rect 4540 9638 4541 9702
rect 4605 9638 4606 9702
rect 4540 9622 4606 9638
rect 4540 9558 4541 9622
rect 4605 9558 4606 9622
rect 4540 9542 4606 9558
rect 4540 9478 4541 9542
rect 4605 9478 4606 9542
rect 4540 9462 4606 9478
rect 4540 9398 4541 9462
rect 4605 9398 4606 9462
rect 4540 9382 4606 9398
rect 4540 9318 4541 9382
rect 4605 9318 4606 9382
rect 4540 9302 4606 9318
rect 4540 9238 4541 9302
rect 4605 9238 4606 9302
rect 4540 9222 4606 9238
rect 4540 9158 4541 9222
rect 4605 9158 4606 9222
rect 4540 9068 4606 9158
rect 4666 9064 4726 10096
rect 4786 9004 4846 10034
rect 4906 9064 4966 10096
rect 5026 9004 5086 10034
rect 5146 9942 5212 10096
rect 5146 9878 5147 9942
rect 5211 9878 5212 9942
rect 5146 9862 5212 9878
rect 5146 9798 5147 9862
rect 5211 9798 5212 9862
rect 5146 9782 5212 9798
rect 5146 9718 5147 9782
rect 5211 9718 5212 9782
rect 5146 9702 5212 9718
rect 5146 9638 5147 9702
rect 5211 9638 5212 9702
rect 5146 9622 5212 9638
rect 5146 9558 5147 9622
rect 5211 9558 5212 9622
rect 5146 9542 5212 9558
rect 5146 9478 5147 9542
rect 5211 9478 5212 9542
rect 5146 9462 5212 9478
rect 5146 9398 5147 9462
rect 5211 9398 5212 9462
rect 5146 9382 5212 9398
rect 5146 9318 5147 9382
rect 5211 9318 5212 9382
rect 5146 9302 5212 9318
rect 5146 9238 5147 9302
rect 5211 9238 5212 9302
rect 5146 9222 5212 9238
rect 5146 9158 5147 9222
rect 5211 9158 5212 9222
rect 5146 9068 5212 9158
rect 5272 9064 5332 10096
rect 5392 9004 5452 10034
rect 5512 9064 5572 10096
rect 5632 9004 5692 10034
rect 5752 9942 5818 10096
rect 5752 9878 5753 9942
rect 5817 9878 5818 9942
rect 5752 9862 5818 9878
rect 5752 9798 5753 9862
rect 5817 9798 5818 9862
rect 5752 9782 5818 9798
rect 5752 9718 5753 9782
rect 5817 9718 5818 9782
rect 5752 9702 5818 9718
rect 5752 9638 5753 9702
rect 5817 9638 5818 9702
rect 5752 9622 5818 9638
rect 5752 9558 5753 9622
rect 5817 9558 5818 9622
rect 5752 9542 5818 9558
rect 5752 9478 5753 9542
rect 5817 9478 5818 9542
rect 5752 9462 5818 9478
rect 5752 9398 5753 9462
rect 5817 9398 5818 9462
rect 5752 9382 5818 9398
rect 5752 9318 5753 9382
rect 5817 9318 5818 9382
rect 5752 9302 5818 9318
rect 5752 9238 5753 9302
rect 5817 9238 5818 9302
rect 5752 9222 5818 9238
rect 5752 9158 5753 9222
rect 5817 9158 5818 9222
rect 5752 9068 5818 9158
rect 904 9002 5818 9004
rect 904 8938 1008 9002
rect 1072 8938 1088 9002
rect 1152 8938 1168 9002
rect 1232 8938 1248 9002
rect 1312 8938 1328 9002
rect 1392 8938 1408 9002
rect 1472 8938 1614 9002
rect 1678 8938 1694 9002
rect 1758 8938 1774 9002
rect 1838 8938 1854 9002
rect 1918 8938 1934 9002
rect 1998 8938 2014 9002
rect 2078 8938 2220 9002
rect 2284 8938 2300 9002
rect 2364 8938 2380 9002
rect 2444 8938 2460 9002
rect 2524 8938 2540 9002
rect 2604 8938 2620 9002
rect 2684 8938 2826 9002
rect 2890 8938 2906 9002
rect 2970 8938 2986 9002
rect 3050 8938 3066 9002
rect 3130 8938 3146 9002
rect 3210 8938 3226 9002
rect 3290 8938 3432 9002
rect 3496 8938 3512 9002
rect 3576 8938 3592 9002
rect 3656 8938 3672 9002
rect 3736 8938 3752 9002
rect 3816 8938 3832 9002
rect 3896 8938 4038 9002
rect 4102 8938 4118 9002
rect 4182 8938 4198 9002
rect 4262 8938 4278 9002
rect 4342 8938 4358 9002
rect 4422 8938 4438 9002
rect 4502 8938 4644 9002
rect 4708 8938 4724 9002
rect 4788 8938 4804 9002
rect 4868 8938 4884 9002
rect 4948 8938 4964 9002
rect 5028 8938 5044 9002
rect 5108 8938 5250 9002
rect 5314 8938 5330 9002
rect 5394 8938 5410 9002
rect 5474 8938 5490 9002
rect 5554 8938 5570 9002
rect 5634 8938 5650 9002
rect 5714 8938 5818 9002
rect 904 8936 5818 8938
rect 904 8782 970 8936
rect 904 8718 905 8782
rect 969 8718 970 8782
rect 904 8702 970 8718
rect 904 8638 905 8702
rect 969 8638 970 8702
rect 904 8622 970 8638
rect 904 8558 905 8622
rect 969 8558 970 8622
rect 904 8542 970 8558
rect 904 8478 905 8542
rect 969 8478 970 8542
rect 904 8462 970 8478
rect 904 8398 905 8462
rect 969 8398 970 8462
rect 904 8382 970 8398
rect 904 8318 905 8382
rect 969 8318 970 8382
rect 904 8302 970 8318
rect 904 8238 905 8302
rect 969 8238 970 8302
rect 904 8222 970 8238
rect 904 8158 905 8222
rect 969 8158 970 8222
rect 904 8142 970 8158
rect 904 8078 905 8142
rect 969 8078 970 8142
rect 904 8062 970 8078
rect 904 7998 905 8062
rect 969 7998 970 8062
rect 904 7908 970 7998
rect 1030 7904 1090 8936
rect 1150 7844 1210 8874
rect 1270 7904 1330 8936
rect 1390 7844 1450 8874
rect 1510 8782 1576 8936
rect 1510 8718 1511 8782
rect 1575 8718 1576 8782
rect 1510 8702 1576 8718
rect 1510 8638 1511 8702
rect 1575 8638 1576 8702
rect 1510 8622 1576 8638
rect 1510 8558 1511 8622
rect 1575 8558 1576 8622
rect 1510 8542 1576 8558
rect 1510 8478 1511 8542
rect 1575 8478 1576 8542
rect 1510 8462 1576 8478
rect 1510 8398 1511 8462
rect 1575 8398 1576 8462
rect 1510 8382 1576 8398
rect 1510 8318 1511 8382
rect 1575 8318 1576 8382
rect 1510 8302 1576 8318
rect 1510 8238 1511 8302
rect 1575 8238 1576 8302
rect 1510 8222 1576 8238
rect 1510 8158 1511 8222
rect 1575 8158 1576 8222
rect 1510 8142 1576 8158
rect 1510 8078 1511 8142
rect 1575 8078 1576 8142
rect 1510 8062 1576 8078
rect 1510 7998 1511 8062
rect 1575 7998 1576 8062
rect 1510 7908 1576 7998
rect 1636 7904 1696 8936
rect 1756 7844 1816 8874
rect 1876 7904 1936 8936
rect 1996 7844 2056 8874
rect 2116 8782 2182 8936
rect 2116 8718 2117 8782
rect 2181 8718 2182 8782
rect 2116 8702 2182 8718
rect 2116 8638 2117 8702
rect 2181 8638 2182 8702
rect 2116 8622 2182 8638
rect 2116 8558 2117 8622
rect 2181 8558 2182 8622
rect 2116 8542 2182 8558
rect 2116 8478 2117 8542
rect 2181 8478 2182 8542
rect 2116 8462 2182 8478
rect 2116 8398 2117 8462
rect 2181 8398 2182 8462
rect 2116 8382 2182 8398
rect 2116 8318 2117 8382
rect 2181 8318 2182 8382
rect 2116 8302 2182 8318
rect 2116 8238 2117 8302
rect 2181 8238 2182 8302
rect 2116 8222 2182 8238
rect 2116 8158 2117 8222
rect 2181 8158 2182 8222
rect 2116 8142 2182 8158
rect 2116 8078 2117 8142
rect 2181 8078 2182 8142
rect 2116 8062 2182 8078
rect 2116 7998 2117 8062
rect 2181 7998 2182 8062
rect 2116 7908 2182 7998
rect 2242 7904 2302 8936
rect 2362 7844 2422 8874
rect 2482 7904 2542 8936
rect 2602 7844 2662 8874
rect 2722 8782 2788 8936
rect 2722 8718 2723 8782
rect 2787 8718 2788 8782
rect 2722 8702 2788 8718
rect 2722 8638 2723 8702
rect 2787 8638 2788 8702
rect 2722 8622 2788 8638
rect 2722 8558 2723 8622
rect 2787 8558 2788 8622
rect 2722 8542 2788 8558
rect 2722 8478 2723 8542
rect 2787 8478 2788 8542
rect 2722 8462 2788 8478
rect 2722 8398 2723 8462
rect 2787 8398 2788 8462
rect 2722 8382 2788 8398
rect 2722 8318 2723 8382
rect 2787 8318 2788 8382
rect 2722 8302 2788 8318
rect 2722 8238 2723 8302
rect 2787 8238 2788 8302
rect 2722 8222 2788 8238
rect 2722 8158 2723 8222
rect 2787 8158 2788 8222
rect 2722 8142 2788 8158
rect 2722 8078 2723 8142
rect 2787 8078 2788 8142
rect 2722 8062 2788 8078
rect 2722 7998 2723 8062
rect 2787 7998 2788 8062
rect 2722 7908 2788 7998
rect 2848 7904 2908 8936
rect 2968 7844 3028 8874
rect 3088 7904 3148 8936
rect 3208 7844 3268 8874
rect 3328 8782 3394 8936
rect 3328 8718 3329 8782
rect 3393 8718 3394 8782
rect 3328 8702 3394 8718
rect 3328 8638 3329 8702
rect 3393 8638 3394 8702
rect 3328 8622 3394 8638
rect 3328 8558 3329 8622
rect 3393 8558 3394 8622
rect 3328 8542 3394 8558
rect 3328 8478 3329 8542
rect 3393 8478 3394 8542
rect 3328 8462 3394 8478
rect 3328 8398 3329 8462
rect 3393 8398 3394 8462
rect 3328 8382 3394 8398
rect 3328 8318 3329 8382
rect 3393 8318 3394 8382
rect 3328 8302 3394 8318
rect 3328 8238 3329 8302
rect 3393 8238 3394 8302
rect 3328 8222 3394 8238
rect 3328 8158 3329 8222
rect 3393 8158 3394 8222
rect 3328 8142 3394 8158
rect 3328 8078 3329 8142
rect 3393 8078 3394 8142
rect 3328 8062 3394 8078
rect 3328 7998 3329 8062
rect 3393 7998 3394 8062
rect 3328 7908 3394 7998
rect 3454 7904 3514 8936
rect 3574 7844 3634 8874
rect 3694 7904 3754 8936
rect 3814 7844 3874 8874
rect 3934 8782 4000 8936
rect 3934 8718 3935 8782
rect 3999 8718 4000 8782
rect 3934 8702 4000 8718
rect 3934 8638 3935 8702
rect 3999 8638 4000 8702
rect 3934 8622 4000 8638
rect 3934 8558 3935 8622
rect 3999 8558 4000 8622
rect 3934 8542 4000 8558
rect 3934 8478 3935 8542
rect 3999 8478 4000 8542
rect 3934 8462 4000 8478
rect 3934 8398 3935 8462
rect 3999 8398 4000 8462
rect 3934 8382 4000 8398
rect 3934 8318 3935 8382
rect 3999 8318 4000 8382
rect 3934 8302 4000 8318
rect 3934 8238 3935 8302
rect 3999 8238 4000 8302
rect 3934 8222 4000 8238
rect 3934 8158 3935 8222
rect 3999 8158 4000 8222
rect 3934 8142 4000 8158
rect 3934 8078 3935 8142
rect 3999 8078 4000 8142
rect 3934 8062 4000 8078
rect 3934 7998 3935 8062
rect 3999 7998 4000 8062
rect 3934 7908 4000 7998
rect 4060 7904 4120 8936
rect 4180 7844 4240 8874
rect 4300 7904 4360 8936
rect 4420 7844 4480 8874
rect 4540 8782 4606 8936
rect 4540 8718 4541 8782
rect 4605 8718 4606 8782
rect 4540 8702 4606 8718
rect 4540 8638 4541 8702
rect 4605 8638 4606 8702
rect 4540 8622 4606 8638
rect 4540 8558 4541 8622
rect 4605 8558 4606 8622
rect 4540 8542 4606 8558
rect 4540 8478 4541 8542
rect 4605 8478 4606 8542
rect 4540 8462 4606 8478
rect 4540 8398 4541 8462
rect 4605 8398 4606 8462
rect 4540 8382 4606 8398
rect 4540 8318 4541 8382
rect 4605 8318 4606 8382
rect 4540 8302 4606 8318
rect 4540 8238 4541 8302
rect 4605 8238 4606 8302
rect 4540 8222 4606 8238
rect 4540 8158 4541 8222
rect 4605 8158 4606 8222
rect 4540 8142 4606 8158
rect 4540 8078 4541 8142
rect 4605 8078 4606 8142
rect 4540 8062 4606 8078
rect 4540 7998 4541 8062
rect 4605 7998 4606 8062
rect 4540 7908 4606 7998
rect 4666 7904 4726 8936
rect 4786 7844 4846 8874
rect 4906 7904 4966 8936
rect 5026 7844 5086 8874
rect 5146 8782 5212 8936
rect 5146 8718 5147 8782
rect 5211 8718 5212 8782
rect 5146 8702 5212 8718
rect 5146 8638 5147 8702
rect 5211 8638 5212 8702
rect 5146 8622 5212 8638
rect 5146 8558 5147 8622
rect 5211 8558 5212 8622
rect 5146 8542 5212 8558
rect 5146 8478 5147 8542
rect 5211 8478 5212 8542
rect 5146 8462 5212 8478
rect 5146 8398 5147 8462
rect 5211 8398 5212 8462
rect 5146 8382 5212 8398
rect 5146 8318 5147 8382
rect 5211 8318 5212 8382
rect 5146 8302 5212 8318
rect 5146 8238 5147 8302
rect 5211 8238 5212 8302
rect 5146 8222 5212 8238
rect 5146 8158 5147 8222
rect 5211 8158 5212 8222
rect 5146 8142 5212 8158
rect 5146 8078 5147 8142
rect 5211 8078 5212 8142
rect 5146 8062 5212 8078
rect 5146 7998 5147 8062
rect 5211 7998 5212 8062
rect 5146 7908 5212 7998
rect 5272 7904 5332 8936
rect 5392 7844 5452 8874
rect 5512 7904 5572 8936
rect 5632 7844 5692 8874
rect 5752 8782 5818 8936
rect 5752 8718 5753 8782
rect 5817 8718 5818 8782
rect 5752 8702 5818 8718
rect 5752 8638 5753 8702
rect 5817 8638 5818 8702
rect 5752 8622 5818 8638
rect 5752 8558 5753 8622
rect 5817 8558 5818 8622
rect 5752 8542 5818 8558
rect 5752 8478 5753 8542
rect 5817 8478 5818 8542
rect 5752 8462 5818 8478
rect 5752 8398 5753 8462
rect 5817 8398 5818 8462
rect 5752 8382 5818 8398
rect 5752 8318 5753 8382
rect 5817 8318 5818 8382
rect 5752 8302 5818 8318
rect 5752 8238 5753 8302
rect 5817 8238 5818 8302
rect 5752 8222 5818 8238
rect 5752 8158 5753 8222
rect 5817 8158 5818 8222
rect 5752 8142 5818 8158
rect 5752 8078 5753 8142
rect 5817 8078 5818 8142
rect 5752 8062 5818 8078
rect 5752 7998 5753 8062
rect 5817 7998 5818 8062
rect 5752 7908 5818 7998
rect 904 7842 5818 7844
rect 904 7778 1008 7842
rect 1072 7778 1088 7842
rect 1152 7778 1168 7842
rect 1232 7778 1248 7842
rect 1312 7778 1328 7842
rect 1392 7778 1408 7842
rect 1472 7778 1614 7842
rect 1678 7778 1694 7842
rect 1758 7778 1774 7842
rect 1838 7778 1854 7842
rect 1918 7778 1934 7842
rect 1998 7778 2014 7842
rect 2078 7778 2220 7842
rect 2284 7778 2300 7842
rect 2364 7778 2380 7842
rect 2444 7778 2460 7842
rect 2524 7778 2540 7842
rect 2604 7778 2620 7842
rect 2684 7778 2826 7842
rect 2890 7778 2906 7842
rect 2970 7778 2986 7842
rect 3050 7778 3066 7842
rect 3130 7778 3146 7842
rect 3210 7778 3226 7842
rect 3290 7778 3432 7842
rect 3496 7778 3512 7842
rect 3576 7778 3592 7842
rect 3656 7778 3672 7842
rect 3736 7778 3752 7842
rect 3816 7778 3832 7842
rect 3896 7778 4038 7842
rect 4102 7778 4118 7842
rect 4182 7778 4198 7842
rect 4262 7778 4278 7842
rect 4342 7778 4358 7842
rect 4422 7778 4438 7842
rect 4502 7778 4644 7842
rect 4708 7778 4724 7842
rect 4788 7778 4804 7842
rect 4868 7778 4884 7842
rect 4948 7778 4964 7842
rect 5028 7778 5044 7842
rect 5108 7778 5250 7842
rect 5314 7778 5330 7842
rect 5394 7778 5410 7842
rect 5474 7778 5490 7842
rect 5554 7778 5570 7842
rect 5634 7778 5650 7842
rect 5714 7778 5818 7842
rect 904 7776 5818 7778
<< via3 >>
rect 1008 10098 1072 10162
rect 1088 10098 1152 10162
rect 1168 10098 1232 10162
rect 1248 10098 1312 10162
rect 1328 10098 1392 10162
rect 1408 10098 1472 10162
rect 1614 10098 1678 10162
rect 1694 10098 1758 10162
rect 1774 10098 1838 10162
rect 1854 10098 1918 10162
rect 1934 10098 1998 10162
rect 2014 10098 2078 10162
rect 2220 10098 2284 10162
rect 2300 10098 2364 10162
rect 2380 10098 2444 10162
rect 2460 10098 2524 10162
rect 2540 10098 2604 10162
rect 2620 10098 2684 10162
rect 2826 10098 2890 10162
rect 2906 10098 2970 10162
rect 2986 10098 3050 10162
rect 3066 10098 3130 10162
rect 3146 10098 3210 10162
rect 3226 10098 3290 10162
rect 3432 10098 3496 10162
rect 3512 10098 3576 10162
rect 3592 10098 3656 10162
rect 3672 10098 3736 10162
rect 3752 10098 3816 10162
rect 3832 10098 3896 10162
rect 4038 10098 4102 10162
rect 4118 10098 4182 10162
rect 4198 10098 4262 10162
rect 4278 10098 4342 10162
rect 4358 10098 4422 10162
rect 4438 10098 4502 10162
rect 4644 10098 4708 10162
rect 4724 10098 4788 10162
rect 4804 10098 4868 10162
rect 4884 10098 4948 10162
rect 4964 10098 5028 10162
rect 5044 10098 5108 10162
rect 5250 10098 5314 10162
rect 5330 10098 5394 10162
rect 5410 10098 5474 10162
rect 5490 10098 5554 10162
rect 5570 10098 5634 10162
rect 5650 10098 5714 10162
rect 905 9878 969 9942
rect 905 9798 969 9862
rect 905 9718 969 9782
rect 905 9638 969 9702
rect 905 9558 969 9622
rect 905 9478 969 9542
rect 905 9398 969 9462
rect 905 9318 969 9382
rect 905 9238 969 9302
rect 905 9158 969 9222
rect 1511 9878 1575 9942
rect 1511 9798 1575 9862
rect 1511 9718 1575 9782
rect 1511 9638 1575 9702
rect 1511 9558 1575 9622
rect 1511 9478 1575 9542
rect 1511 9398 1575 9462
rect 1511 9318 1575 9382
rect 1511 9238 1575 9302
rect 1511 9158 1575 9222
rect 2117 9878 2181 9942
rect 2117 9798 2181 9862
rect 2117 9718 2181 9782
rect 2117 9638 2181 9702
rect 2117 9558 2181 9622
rect 2117 9478 2181 9542
rect 2117 9398 2181 9462
rect 2117 9318 2181 9382
rect 2117 9238 2181 9302
rect 2117 9158 2181 9222
rect 2723 9878 2787 9942
rect 2723 9798 2787 9862
rect 2723 9718 2787 9782
rect 2723 9638 2787 9702
rect 2723 9558 2787 9622
rect 2723 9478 2787 9542
rect 2723 9398 2787 9462
rect 2723 9318 2787 9382
rect 2723 9238 2787 9302
rect 2723 9158 2787 9222
rect 3329 9878 3393 9942
rect 3329 9798 3393 9862
rect 3329 9718 3393 9782
rect 3329 9638 3393 9702
rect 3329 9558 3393 9622
rect 3329 9478 3393 9542
rect 3329 9398 3393 9462
rect 3329 9318 3393 9382
rect 3329 9238 3393 9302
rect 3329 9158 3393 9222
rect 3935 9878 3999 9942
rect 3935 9798 3999 9862
rect 3935 9718 3999 9782
rect 3935 9638 3999 9702
rect 3935 9558 3999 9622
rect 3935 9478 3999 9542
rect 3935 9398 3999 9462
rect 3935 9318 3999 9382
rect 3935 9238 3999 9302
rect 3935 9158 3999 9222
rect 4541 9878 4605 9942
rect 4541 9798 4605 9862
rect 4541 9718 4605 9782
rect 4541 9638 4605 9702
rect 4541 9558 4605 9622
rect 4541 9478 4605 9542
rect 4541 9398 4605 9462
rect 4541 9318 4605 9382
rect 4541 9238 4605 9302
rect 4541 9158 4605 9222
rect 5147 9878 5211 9942
rect 5147 9798 5211 9862
rect 5147 9718 5211 9782
rect 5147 9638 5211 9702
rect 5147 9558 5211 9622
rect 5147 9478 5211 9542
rect 5147 9398 5211 9462
rect 5147 9318 5211 9382
rect 5147 9238 5211 9302
rect 5147 9158 5211 9222
rect 5753 9878 5817 9942
rect 5753 9798 5817 9862
rect 5753 9718 5817 9782
rect 5753 9638 5817 9702
rect 5753 9558 5817 9622
rect 5753 9478 5817 9542
rect 5753 9398 5817 9462
rect 5753 9318 5817 9382
rect 5753 9238 5817 9302
rect 5753 9158 5817 9222
rect 1008 8938 1072 9002
rect 1088 8938 1152 9002
rect 1168 8938 1232 9002
rect 1248 8938 1312 9002
rect 1328 8938 1392 9002
rect 1408 8938 1472 9002
rect 1614 8938 1678 9002
rect 1694 8938 1758 9002
rect 1774 8938 1838 9002
rect 1854 8938 1918 9002
rect 1934 8938 1998 9002
rect 2014 8938 2078 9002
rect 2220 8938 2284 9002
rect 2300 8938 2364 9002
rect 2380 8938 2444 9002
rect 2460 8938 2524 9002
rect 2540 8938 2604 9002
rect 2620 8938 2684 9002
rect 2826 8938 2890 9002
rect 2906 8938 2970 9002
rect 2986 8938 3050 9002
rect 3066 8938 3130 9002
rect 3146 8938 3210 9002
rect 3226 8938 3290 9002
rect 3432 8938 3496 9002
rect 3512 8938 3576 9002
rect 3592 8938 3656 9002
rect 3672 8938 3736 9002
rect 3752 8938 3816 9002
rect 3832 8938 3896 9002
rect 4038 8938 4102 9002
rect 4118 8938 4182 9002
rect 4198 8938 4262 9002
rect 4278 8938 4342 9002
rect 4358 8938 4422 9002
rect 4438 8938 4502 9002
rect 4644 8938 4708 9002
rect 4724 8938 4788 9002
rect 4804 8938 4868 9002
rect 4884 8938 4948 9002
rect 4964 8938 5028 9002
rect 5044 8938 5108 9002
rect 5250 8938 5314 9002
rect 5330 8938 5394 9002
rect 5410 8938 5474 9002
rect 5490 8938 5554 9002
rect 5570 8938 5634 9002
rect 5650 8938 5714 9002
rect 905 8718 969 8782
rect 905 8638 969 8702
rect 905 8558 969 8622
rect 905 8478 969 8542
rect 905 8398 969 8462
rect 905 8318 969 8382
rect 905 8238 969 8302
rect 905 8158 969 8222
rect 905 8078 969 8142
rect 905 7998 969 8062
rect 1511 8718 1575 8782
rect 1511 8638 1575 8702
rect 1511 8558 1575 8622
rect 1511 8478 1575 8542
rect 1511 8398 1575 8462
rect 1511 8318 1575 8382
rect 1511 8238 1575 8302
rect 1511 8158 1575 8222
rect 1511 8078 1575 8142
rect 1511 7998 1575 8062
rect 2117 8718 2181 8782
rect 2117 8638 2181 8702
rect 2117 8558 2181 8622
rect 2117 8478 2181 8542
rect 2117 8398 2181 8462
rect 2117 8318 2181 8382
rect 2117 8238 2181 8302
rect 2117 8158 2181 8222
rect 2117 8078 2181 8142
rect 2117 7998 2181 8062
rect 2723 8718 2787 8782
rect 2723 8638 2787 8702
rect 2723 8558 2787 8622
rect 2723 8478 2787 8542
rect 2723 8398 2787 8462
rect 2723 8318 2787 8382
rect 2723 8238 2787 8302
rect 2723 8158 2787 8222
rect 2723 8078 2787 8142
rect 2723 7998 2787 8062
rect 3329 8718 3393 8782
rect 3329 8638 3393 8702
rect 3329 8558 3393 8622
rect 3329 8478 3393 8542
rect 3329 8398 3393 8462
rect 3329 8318 3393 8382
rect 3329 8238 3393 8302
rect 3329 8158 3393 8222
rect 3329 8078 3393 8142
rect 3329 7998 3393 8062
rect 3935 8718 3999 8782
rect 3935 8638 3999 8702
rect 3935 8558 3999 8622
rect 3935 8478 3999 8542
rect 3935 8398 3999 8462
rect 3935 8318 3999 8382
rect 3935 8238 3999 8302
rect 3935 8158 3999 8222
rect 3935 8078 3999 8142
rect 3935 7998 3999 8062
rect 4541 8718 4605 8782
rect 4541 8638 4605 8702
rect 4541 8558 4605 8622
rect 4541 8478 4605 8542
rect 4541 8398 4605 8462
rect 4541 8318 4605 8382
rect 4541 8238 4605 8302
rect 4541 8158 4605 8222
rect 4541 8078 4605 8142
rect 4541 7998 4605 8062
rect 5147 8718 5211 8782
rect 5147 8638 5211 8702
rect 5147 8558 5211 8622
rect 5147 8478 5211 8542
rect 5147 8398 5211 8462
rect 5147 8318 5211 8382
rect 5147 8238 5211 8302
rect 5147 8158 5211 8222
rect 5147 8078 5211 8142
rect 5147 7998 5211 8062
rect 5753 8718 5817 8782
rect 5753 8638 5817 8702
rect 5753 8558 5817 8622
rect 5753 8478 5817 8542
rect 5753 8398 5817 8462
rect 5753 8318 5817 8382
rect 5753 8238 5817 8302
rect 5753 8158 5817 8222
rect 5753 8078 5817 8142
rect 5753 7998 5817 8062
rect 1008 7778 1072 7842
rect 1088 7778 1152 7842
rect 1168 7778 1232 7842
rect 1248 7778 1312 7842
rect 1328 7778 1392 7842
rect 1408 7778 1472 7842
rect 1614 7778 1678 7842
rect 1694 7778 1758 7842
rect 1774 7778 1838 7842
rect 1854 7778 1918 7842
rect 1934 7778 1998 7842
rect 2014 7778 2078 7842
rect 2220 7778 2284 7842
rect 2300 7778 2364 7842
rect 2380 7778 2444 7842
rect 2460 7778 2524 7842
rect 2540 7778 2604 7842
rect 2620 7778 2684 7842
rect 2826 7778 2890 7842
rect 2906 7778 2970 7842
rect 2986 7778 3050 7842
rect 3066 7778 3130 7842
rect 3146 7778 3210 7842
rect 3226 7778 3290 7842
rect 3432 7778 3496 7842
rect 3512 7778 3576 7842
rect 3592 7778 3656 7842
rect 3672 7778 3736 7842
rect 3752 7778 3816 7842
rect 3832 7778 3896 7842
rect 4038 7778 4102 7842
rect 4118 7778 4182 7842
rect 4198 7778 4262 7842
rect 4278 7778 4342 7842
rect 4358 7778 4422 7842
rect 4438 7778 4502 7842
rect 4644 7778 4708 7842
rect 4724 7778 4788 7842
rect 4804 7778 4868 7842
rect 4884 7778 4948 7842
rect 4964 7778 5028 7842
rect 5044 7778 5108 7842
rect 5250 7778 5314 7842
rect 5330 7778 5394 7842
rect 5410 7778 5474 7842
rect 5490 7778 5554 7842
rect 5570 7778 5634 7842
rect 5650 7778 5714 7842
<< metal4 >>
rect 904 10162 5818 10164
rect 904 10098 1008 10162
rect 1072 10098 1088 10162
rect 1152 10098 1168 10162
rect 1232 10098 1248 10162
rect 1312 10098 1328 10162
rect 1392 10098 1408 10162
rect 1472 10098 1614 10162
rect 1678 10098 1694 10162
rect 1758 10098 1774 10162
rect 1838 10098 1854 10162
rect 1918 10098 1934 10162
rect 1998 10098 2014 10162
rect 2078 10098 2220 10162
rect 2284 10098 2300 10162
rect 2364 10098 2380 10162
rect 2444 10098 2460 10162
rect 2524 10098 2540 10162
rect 2604 10098 2620 10162
rect 2684 10098 2826 10162
rect 2890 10098 2906 10162
rect 2970 10098 2986 10162
rect 3050 10098 3066 10162
rect 3130 10098 3146 10162
rect 3210 10098 3226 10162
rect 3290 10098 3432 10162
rect 3496 10098 3512 10162
rect 3576 10098 3592 10162
rect 3656 10098 3672 10162
rect 3736 10098 3752 10162
rect 3816 10098 3832 10162
rect 3896 10098 4038 10162
rect 4102 10098 4118 10162
rect 4182 10098 4198 10162
rect 4262 10098 4278 10162
rect 4342 10098 4358 10162
rect 4422 10098 4438 10162
rect 4502 10098 4644 10162
rect 4708 10098 4724 10162
rect 4788 10098 4804 10162
rect 4868 10098 4884 10162
rect 4948 10098 4964 10162
rect 5028 10098 5044 10162
rect 5108 10098 5250 10162
rect 5314 10098 5330 10162
rect 5394 10098 5410 10162
rect 5474 10098 5490 10162
rect 5554 10098 5570 10162
rect 5634 10098 5650 10162
rect 5714 10098 5818 10162
rect 904 10096 5818 10098
rect 904 9942 970 10096
rect 904 9878 905 9942
rect 969 9878 970 9942
rect 904 9862 970 9878
rect 904 9798 905 9862
rect 969 9798 970 9862
rect 904 9782 970 9798
rect 904 9718 905 9782
rect 969 9718 970 9782
rect 904 9702 970 9718
rect 904 9638 905 9702
rect 969 9638 970 9702
rect 904 9622 970 9638
rect 904 9558 905 9622
rect 969 9558 970 9622
rect 904 9542 970 9558
rect 904 9478 905 9542
rect 969 9478 970 9542
rect 904 9462 970 9478
rect 904 9398 905 9462
rect 969 9398 970 9462
rect 904 9382 970 9398
rect 904 9318 905 9382
rect 969 9318 970 9382
rect 904 9302 970 9318
rect 904 9238 905 9302
rect 969 9238 970 9302
rect 904 9222 970 9238
rect 904 9158 905 9222
rect 969 9158 970 9222
rect 904 9068 970 9158
rect 1030 9004 1090 10034
rect 1150 9064 1210 10096
rect 1270 9004 1330 10034
rect 1390 9064 1450 10096
rect 1510 9942 1576 10096
rect 1510 9878 1511 9942
rect 1575 9878 1576 9942
rect 1510 9862 1576 9878
rect 1510 9798 1511 9862
rect 1575 9798 1576 9862
rect 1510 9782 1576 9798
rect 1510 9718 1511 9782
rect 1575 9718 1576 9782
rect 1510 9702 1576 9718
rect 1510 9638 1511 9702
rect 1575 9638 1576 9702
rect 1510 9622 1576 9638
rect 1510 9558 1511 9622
rect 1575 9558 1576 9622
rect 1510 9542 1576 9558
rect 1510 9478 1511 9542
rect 1575 9478 1576 9542
rect 1510 9462 1576 9478
rect 1510 9398 1511 9462
rect 1575 9398 1576 9462
rect 1510 9382 1576 9398
rect 1510 9318 1511 9382
rect 1575 9318 1576 9382
rect 1510 9302 1576 9318
rect 1510 9238 1511 9302
rect 1575 9238 1576 9302
rect 1510 9222 1576 9238
rect 1510 9158 1511 9222
rect 1575 9158 1576 9222
rect 1510 9068 1576 9158
rect 1636 9004 1696 10034
rect 1756 9064 1816 10096
rect 1876 9004 1936 10034
rect 1996 9064 2056 10096
rect 2116 9942 2182 10096
rect 2116 9878 2117 9942
rect 2181 9878 2182 9942
rect 2116 9862 2182 9878
rect 2116 9798 2117 9862
rect 2181 9798 2182 9862
rect 2116 9782 2182 9798
rect 2116 9718 2117 9782
rect 2181 9718 2182 9782
rect 2116 9702 2182 9718
rect 2116 9638 2117 9702
rect 2181 9638 2182 9702
rect 2116 9622 2182 9638
rect 2116 9558 2117 9622
rect 2181 9558 2182 9622
rect 2116 9542 2182 9558
rect 2116 9478 2117 9542
rect 2181 9478 2182 9542
rect 2116 9462 2182 9478
rect 2116 9398 2117 9462
rect 2181 9398 2182 9462
rect 2116 9382 2182 9398
rect 2116 9318 2117 9382
rect 2181 9318 2182 9382
rect 2116 9302 2182 9318
rect 2116 9238 2117 9302
rect 2181 9238 2182 9302
rect 2116 9222 2182 9238
rect 2116 9158 2117 9222
rect 2181 9158 2182 9222
rect 2116 9068 2182 9158
rect 2242 9004 2302 10034
rect 2362 9064 2422 10096
rect 2482 9004 2542 10034
rect 2602 9064 2662 10096
rect 2722 9942 2788 10096
rect 2722 9878 2723 9942
rect 2787 9878 2788 9942
rect 2722 9862 2788 9878
rect 2722 9798 2723 9862
rect 2787 9798 2788 9862
rect 2722 9782 2788 9798
rect 2722 9718 2723 9782
rect 2787 9718 2788 9782
rect 2722 9702 2788 9718
rect 2722 9638 2723 9702
rect 2787 9638 2788 9702
rect 2722 9622 2788 9638
rect 2722 9558 2723 9622
rect 2787 9558 2788 9622
rect 2722 9542 2788 9558
rect 2722 9478 2723 9542
rect 2787 9478 2788 9542
rect 2722 9462 2788 9478
rect 2722 9398 2723 9462
rect 2787 9398 2788 9462
rect 2722 9382 2788 9398
rect 2722 9318 2723 9382
rect 2787 9318 2788 9382
rect 2722 9302 2788 9318
rect 2722 9238 2723 9302
rect 2787 9238 2788 9302
rect 2722 9222 2788 9238
rect 2722 9158 2723 9222
rect 2787 9158 2788 9222
rect 2722 9068 2788 9158
rect 2848 9004 2908 10034
rect 2968 9064 3028 10096
rect 3088 9004 3148 10034
rect 3208 9064 3268 10096
rect 3328 9942 3394 10096
rect 3328 9878 3329 9942
rect 3393 9878 3394 9942
rect 3328 9862 3394 9878
rect 3328 9798 3329 9862
rect 3393 9798 3394 9862
rect 3328 9782 3394 9798
rect 3328 9718 3329 9782
rect 3393 9718 3394 9782
rect 3328 9702 3394 9718
rect 3328 9638 3329 9702
rect 3393 9638 3394 9702
rect 3328 9622 3394 9638
rect 3328 9558 3329 9622
rect 3393 9558 3394 9622
rect 3328 9542 3394 9558
rect 3328 9478 3329 9542
rect 3393 9478 3394 9542
rect 3328 9462 3394 9478
rect 3328 9398 3329 9462
rect 3393 9398 3394 9462
rect 3328 9382 3394 9398
rect 3328 9318 3329 9382
rect 3393 9318 3394 9382
rect 3328 9302 3394 9318
rect 3328 9238 3329 9302
rect 3393 9238 3394 9302
rect 3328 9222 3394 9238
rect 3328 9158 3329 9222
rect 3393 9158 3394 9222
rect 3328 9068 3394 9158
rect 3454 9004 3514 10034
rect 3574 9064 3634 10096
rect 3694 9004 3754 10034
rect 3814 9064 3874 10096
rect 3934 9942 4000 10096
rect 3934 9878 3935 9942
rect 3999 9878 4000 9942
rect 3934 9862 4000 9878
rect 3934 9798 3935 9862
rect 3999 9798 4000 9862
rect 3934 9782 4000 9798
rect 3934 9718 3935 9782
rect 3999 9718 4000 9782
rect 3934 9702 4000 9718
rect 3934 9638 3935 9702
rect 3999 9638 4000 9702
rect 3934 9622 4000 9638
rect 3934 9558 3935 9622
rect 3999 9558 4000 9622
rect 3934 9542 4000 9558
rect 3934 9478 3935 9542
rect 3999 9478 4000 9542
rect 3934 9462 4000 9478
rect 3934 9398 3935 9462
rect 3999 9398 4000 9462
rect 3934 9382 4000 9398
rect 3934 9318 3935 9382
rect 3999 9318 4000 9382
rect 3934 9302 4000 9318
rect 3934 9238 3935 9302
rect 3999 9238 4000 9302
rect 3934 9222 4000 9238
rect 3934 9158 3935 9222
rect 3999 9158 4000 9222
rect 3934 9068 4000 9158
rect 4060 9004 4120 10034
rect 4180 9064 4240 10096
rect 4300 9004 4360 10034
rect 4420 9064 4480 10096
rect 4540 9942 4606 10096
rect 4540 9878 4541 9942
rect 4605 9878 4606 9942
rect 4540 9862 4606 9878
rect 4540 9798 4541 9862
rect 4605 9798 4606 9862
rect 4540 9782 4606 9798
rect 4540 9718 4541 9782
rect 4605 9718 4606 9782
rect 4540 9702 4606 9718
rect 4540 9638 4541 9702
rect 4605 9638 4606 9702
rect 4540 9622 4606 9638
rect 4540 9558 4541 9622
rect 4605 9558 4606 9622
rect 4540 9542 4606 9558
rect 4540 9478 4541 9542
rect 4605 9478 4606 9542
rect 4540 9462 4606 9478
rect 4540 9398 4541 9462
rect 4605 9398 4606 9462
rect 4540 9382 4606 9398
rect 4540 9318 4541 9382
rect 4605 9318 4606 9382
rect 4540 9302 4606 9318
rect 4540 9238 4541 9302
rect 4605 9238 4606 9302
rect 4540 9222 4606 9238
rect 4540 9158 4541 9222
rect 4605 9158 4606 9222
rect 4540 9068 4606 9158
rect 4666 9004 4726 10034
rect 4786 9064 4846 10096
rect 4906 9004 4966 10034
rect 5026 9064 5086 10096
rect 5146 9942 5212 10096
rect 5146 9878 5147 9942
rect 5211 9878 5212 9942
rect 5146 9862 5212 9878
rect 5146 9798 5147 9862
rect 5211 9798 5212 9862
rect 5146 9782 5212 9798
rect 5146 9718 5147 9782
rect 5211 9718 5212 9782
rect 5146 9702 5212 9718
rect 5146 9638 5147 9702
rect 5211 9638 5212 9702
rect 5146 9622 5212 9638
rect 5146 9558 5147 9622
rect 5211 9558 5212 9622
rect 5146 9542 5212 9558
rect 5146 9478 5147 9542
rect 5211 9478 5212 9542
rect 5146 9462 5212 9478
rect 5146 9398 5147 9462
rect 5211 9398 5212 9462
rect 5146 9382 5212 9398
rect 5146 9318 5147 9382
rect 5211 9318 5212 9382
rect 5146 9302 5212 9318
rect 5146 9238 5147 9302
rect 5211 9238 5212 9302
rect 5146 9222 5212 9238
rect 5146 9158 5147 9222
rect 5211 9158 5212 9222
rect 5146 9068 5212 9158
rect 5272 9004 5332 10034
rect 5392 9064 5452 10096
rect 5512 9004 5572 10034
rect 5632 9064 5692 10096
rect 5752 9942 5818 10096
rect 5752 9878 5753 9942
rect 5817 9878 5818 9942
rect 5752 9862 5818 9878
rect 5752 9798 5753 9862
rect 5817 9798 5818 9862
rect 5752 9782 5818 9798
rect 5752 9718 5753 9782
rect 5817 9718 5818 9782
rect 5752 9702 5818 9718
rect 5752 9638 5753 9702
rect 5817 9638 5818 9702
rect 5752 9622 5818 9638
rect 5752 9558 5753 9622
rect 5817 9558 5818 9622
rect 5752 9542 5818 9558
rect 5752 9478 5753 9542
rect 5817 9478 5818 9542
rect 5752 9462 5818 9478
rect 5752 9398 5753 9462
rect 5817 9398 5818 9462
rect 5752 9382 5818 9398
rect 5752 9318 5753 9382
rect 5817 9318 5818 9382
rect 5752 9302 5818 9318
rect 5752 9238 5753 9302
rect 5817 9238 5818 9302
rect 5752 9222 5818 9238
rect 5752 9158 5753 9222
rect 5817 9158 5818 9222
rect 5752 9068 5818 9158
rect 904 9002 5818 9004
rect 904 8938 1008 9002
rect 1072 8938 1088 9002
rect 1152 8938 1168 9002
rect 1232 8938 1248 9002
rect 1312 8938 1328 9002
rect 1392 8938 1408 9002
rect 1472 8938 1614 9002
rect 1678 8938 1694 9002
rect 1758 8938 1774 9002
rect 1838 8938 1854 9002
rect 1918 8938 1934 9002
rect 1998 8938 2014 9002
rect 2078 8938 2220 9002
rect 2284 8938 2300 9002
rect 2364 8938 2380 9002
rect 2444 8938 2460 9002
rect 2524 8938 2540 9002
rect 2604 8938 2620 9002
rect 2684 8938 2826 9002
rect 2890 8938 2906 9002
rect 2970 8938 2986 9002
rect 3050 8938 3066 9002
rect 3130 8938 3146 9002
rect 3210 8938 3226 9002
rect 3290 8938 3432 9002
rect 3496 8938 3512 9002
rect 3576 8938 3592 9002
rect 3656 8938 3672 9002
rect 3736 8938 3752 9002
rect 3816 8938 3832 9002
rect 3896 8938 4038 9002
rect 4102 8938 4118 9002
rect 4182 8938 4198 9002
rect 4262 8938 4278 9002
rect 4342 8938 4358 9002
rect 4422 8938 4438 9002
rect 4502 8938 4644 9002
rect 4708 8938 4724 9002
rect 4788 8938 4804 9002
rect 4868 8938 4884 9002
rect 4948 8938 4964 9002
rect 5028 8938 5044 9002
rect 5108 8938 5250 9002
rect 5314 8938 5330 9002
rect 5394 8938 5410 9002
rect 5474 8938 5490 9002
rect 5554 8938 5570 9002
rect 5634 8938 5650 9002
rect 5714 8938 5818 9002
rect 904 8936 5818 8938
rect 904 8782 970 8936
rect 904 8718 905 8782
rect 969 8718 970 8782
rect 904 8702 970 8718
rect 904 8638 905 8702
rect 969 8638 970 8702
rect 904 8622 970 8638
rect 904 8558 905 8622
rect 969 8558 970 8622
rect 904 8542 970 8558
rect 904 8478 905 8542
rect 969 8478 970 8542
rect 904 8462 970 8478
rect 904 8398 905 8462
rect 969 8398 970 8462
rect 904 8382 970 8398
rect 904 8318 905 8382
rect 969 8318 970 8382
rect 904 8302 970 8318
rect 904 8238 905 8302
rect 969 8238 970 8302
rect 904 8222 970 8238
rect 904 8158 905 8222
rect 969 8158 970 8222
rect 904 8142 970 8158
rect 904 8078 905 8142
rect 969 8078 970 8142
rect 904 8062 970 8078
rect 904 7998 905 8062
rect 969 7998 970 8062
rect 904 7908 970 7998
rect 1030 7844 1090 8874
rect 1150 7904 1210 8936
rect 1270 7844 1330 8874
rect 1390 7904 1450 8936
rect 1510 8782 1576 8936
rect 1510 8718 1511 8782
rect 1575 8718 1576 8782
rect 1510 8702 1576 8718
rect 1510 8638 1511 8702
rect 1575 8638 1576 8702
rect 1510 8622 1576 8638
rect 1510 8558 1511 8622
rect 1575 8558 1576 8622
rect 1510 8542 1576 8558
rect 1510 8478 1511 8542
rect 1575 8478 1576 8542
rect 1510 8462 1576 8478
rect 1510 8398 1511 8462
rect 1575 8398 1576 8462
rect 1510 8382 1576 8398
rect 1510 8318 1511 8382
rect 1575 8318 1576 8382
rect 1510 8302 1576 8318
rect 1510 8238 1511 8302
rect 1575 8238 1576 8302
rect 1510 8222 1576 8238
rect 1510 8158 1511 8222
rect 1575 8158 1576 8222
rect 1510 8142 1576 8158
rect 1510 8078 1511 8142
rect 1575 8078 1576 8142
rect 1510 8062 1576 8078
rect 1510 7998 1511 8062
rect 1575 7998 1576 8062
rect 1510 7908 1576 7998
rect 1636 7844 1696 8874
rect 1756 7904 1816 8936
rect 1876 7844 1936 8874
rect 1996 7904 2056 8936
rect 2116 8782 2182 8936
rect 2116 8718 2117 8782
rect 2181 8718 2182 8782
rect 2116 8702 2182 8718
rect 2116 8638 2117 8702
rect 2181 8638 2182 8702
rect 2116 8622 2182 8638
rect 2116 8558 2117 8622
rect 2181 8558 2182 8622
rect 2116 8542 2182 8558
rect 2116 8478 2117 8542
rect 2181 8478 2182 8542
rect 2116 8462 2182 8478
rect 2116 8398 2117 8462
rect 2181 8398 2182 8462
rect 2116 8382 2182 8398
rect 2116 8318 2117 8382
rect 2181 8318 2182 8382
rect 2116 8302 2182 8318
rect 2116 8238 2117 8302
rect 2181 8238 2182 8302
rect 2116 8222 2182 8238
rect 2116 8158 2117 8222
rect 2181 8158 2182 8222
rect 2116 8142 2182 8158
rect 2116 8078 2117 8142
rect 2181 8078 2182 8142
rect 2116 8062 2182 8078
rect 2116 7998 2117 8062
rect 2181 7998 2182 8062
rect 2116 7908 2182 7998
rect 2242 7844 2302 8874
rect 2362 7904 2422 8936
rect 2482 7844 2542 8874
rect 2602 7904 2662 8936
rect 2722 8782 2788 8936
rect 2722 8718 2723 8782
rect 2787 8718 2788 8782
rect 2722 8702 2788 8718
rect 2722 8638 2723 8702
rect 2787 8638 2788 8702
rect 2722 8622 2788 8638
rect 2722 8558 2723 8622
rect 2787 8558 2788 8622
rect 2722 8542 2788 8558
rect 2722 8478 2723 8542
rect 2787 8478 2788 8542
rect 2722 8462 2788 8478
rect 2722 8398 2723 8462
rect 2787 8398 2788 8462
rect 2722 8382 2788 8398
rect 2722 8318 2723 8382
rect 2787 8318 2788 8382
rect 2722 8302 2788 8318
rect 2722 8238 2723 8302
rect 2787 8238 2788 8302
rect 2722 8222 2788 8238
rect 2722 8158 2723 8222
rect 2787 8158 2788 8222
rect 2722 8142 2788 8158
rect 2722 8078 2723 8142
rect 2787 8078 2788 8142
rect 2722 8062 2788 8078
rect 2722 7998 2723 8062
rect 2787 7998 2788 8062
rect 2722 7908 2788 7998
rect 2848 7844 2908 8874
rect 2968 7904 3028 8936
rect 3088 7844 3148 8874
rect 3208 7904 3268 8936
rect 3328 8782 3394 8936
rect 3328 8718 3329 8782
rect 3393 8718 3394 8782
rect 3328 8702 3394 8718
rect 3328 8638 3329 8702
rect 3393 8638 3394 8702
rect 3328 8622 3394 8638
rect 3328 8558 3329 8622
rect 3393 8558 3394 8622
rect 3328 8542 3394 8558
rect 3328 8478 3329 8542
rect 3393 8478 3394 8542
rect 3328 8462 3394 8478
rect 3328 8398 3329 8462
rect 3393 8398 3394 8462
rect 3328 8382 3394 8398
rect 3328 8318 3329 8382
rect 3393 8318 3394 8382
rect 3328 8302 3394 8318
rect 3328 8238 3329 8302
rect 3393 8238 3394 8302
rect 3328 8222 3394 8238
rect 3328 8158 3329 8222
rect 3393 8158 3394 8222
rect 3328 8142 3394 8158
rect 3328 8078 3329 8142
rect 3393 8078 3394 8142
rect 3328 8062 3394 8078
rect 3328 7998 3329 8062
rect 3393 7998 3394 8062
rect 3328 7908 3394 7998
rect 3454 7844 3514 8874
rect 3574 7904 3634 8936
rect 3694 7844 3754 8874
rect 3814 7904 3874 8936
rect 3934 8782 4000 8936
rect 3934 8718 3935 8782
rect 3999 8718 4000 8782
rect 3934 8702 4000 8718
rect 3934 8638 3935 8702
rect 3999 8638 4000 8702
rect 3934 8622 4000 8638
rect 3934 8558 3935 8622
rect 3999 8558 4000 8622
rect 3934 8542 4000 8558
rect 3934 8478 3935 8542
rect 3999 8478 4000 8542
rect 3934 8462 4000 8478
rect 3934 8398 3935 8462
rect 3999 8398 4000 8462
rect 3934 8382 4000 8398
rect 3934 8318 3935 8382
rect 3999 8318 4000 8382
rect 3934 8302 4000 8318
rect 3934 8238 3935 8302
rect 3999 8238 4000 8302
rect 3934 8222 4000 8238
rect 3934 8158 3935 8222
rect 3999 8158 4000 8222
rect 3934 8142 4000 8158
rect 3934 8078 3935 8142
rect 3999 8078 4000 8142
rect 3934 8062 4000 8078
rect 3934 7998 3935 8062
rect 3999 7998 4000 8062
rect 3934 7908 4000 7998
rect 4060 7844 4120 8874
rect 4180 7904 4240 8936
rect 4300 7844 4360 8874
rect 4420 7904 4480 8936
rect 4540 8782 4606 8936
rect 4540 8718 4541 8782
rect 4605 8718 4606 8782
rect 4540 8702 4606 8718
rect 4540 8638 4541 8702
rect 4605 8638 4606 8702
rect 4540 8622 4606 8638
rect 4540 8558 4541 8622
rect 4605 8558 4606 8622
rect 4540 8542 4606 8558
rect 4540 8478 4541 8542
rect 4605 8478 4606 8542
rect 4540 8462 4606 8478
rect 4540 8398 4541 8462
rect 4605 8398 4606 8462
rect 4540 8382 4606 8398
rect 4540 8318 4541 8382
rect 4605 8318 4606 8382
rect 4540 8302 4606 8318
rect 4540 8238 4541 8302
rect 4605 8238 4606 8302
rect 4540 8222 4606 8238
rect 4540 8158 4541 8222
rect 4605 8158 4606 8222
rect 4540 8142 4606 8158
rect 4540 8078 4541 8142
rect 4605 8078 4606 8142
rect 4540 8062 4606 8078
rect 4540 7998 4541 8062
rect 4605 7998 4606 8062
rect 4540 7908 4606 7998
rect 4666 7844 4726 8874
rect 4786 7904 4846 8936
rect 4906 7844 4966 8874
rect 5026 7904 5086 8936
rect 5146 8782 5212 8936
rect 5146 8718 5147 8782
rect 5211 8718 5212 8782
rect 5146 8702 5212 8718
rect 5146 8638 5147 8702
rect 5211 8638 5212 8702
rect 5146 8622 5212 8638
rect 5146 8558 5147 8622
rect 5211 8558 5212 8622
rect 5146 8542 5212 8558
rect 5146 8478 5147 8542
rect 5211 8478 5212 8542
rect 5146 8462 5212 8478
rect 5146 8398 5147 8462
rect 5211 8398 5212 8462
rect 5146 8382 5212 8398
rect 5146 8318 5147 8382
rect 5211 8318 5212 8382
rect 5146 8302 5212 8318
rect 5146 8238 5147 8302
rect 5211 8238 5212 8302
rect 5146 8222 5212 8238
rect 5146 8158 5147 8222
rect 5211 8158 5212 8222
rect 5146 8142 5212 8158
rect 5146 8078 5147 8142
rect 5211 8078 5212 8142
rect 5146 8062 5212 8078
rect 5146 7998 5147 8062
rect 5211 7998 5212 8062
rect 5146 7908 5212 7998
rect 5272 7844 5332 8874
rect 5392 7904 5452 8936
rect 5512 7844 5572 8874
rect 5632 7904 5692 8936
rect 5752 8782 5818 8936
rect 5752 8718 5753 8782
rect 5817 8718 5818 8782
rect 5752 8702 5818 8718
rect 5752 8638 5753 8702
rect 5817 8638 5818 8702
rect 5752 8622 5818 8638
rect 5752 8558 5753 8622
rect 5817 8558 5818 8622
rect 5752 8542 5818 8558
rect 5752 8478 5753 8542
rect 5817 8478 5818 8542
rect 5752 8462 5818 8478
rect 5752 8398 5753 8462
rect 5817 8398 5818 8462
rect 5752 8382 5818 8398
rect 5752 8318 5753 8382
rect 5817 8318 5818 8382
rect 5752 8302 5818 8318
rect 5752 8238 5753 8302
rect 5817 8238 5818 8302
rect 5752 8222 5818 8238
rect 5752 8158 5753 8222
rect 5817 8158 5818 8222
rect 5752 8142 5818 8158
rect 5752 8078 5753 8142
rect 5817 8078 5818 8142
rect 5752 8062 5818 8078
rect 5752 7998 5753 8062
rect 5817 7998 5818 8062
rect 5752 7908 5818 7998
rect 904 7842 5818 7844
rect 904 7778 1008 7842
rect 1072 7778 1088 7842
rect 1152 7778 1168 7842
rect 1232 7778 1248 7842
rect 1312 7778 1328 7842
rect 1392 7778 1408 7842
rect 1472 7778 1614 7842
rect 1678 7778 1694 7842
rect 1758 7778 1774 7842
rect 1838 7778 1854 7842
rect 1918 7778 1934 7842
rect 1998 7778 2014 7842
rect 2078 7778 2220 7842
rect 2284 7778 2300 7842
rect 2364 7778 2380 7842
rect 2444 7778 2460 7842
rect 2524 7778 2540 7842
rect 2604 7778 2620 7842
rect 2684 7778 2826 7842
rect 2890 7778 2906 7842
rect 2970 7778 2986 7842
rect 3050 7778 3066 7842
rect 3130 7778 3146 7842
rect 3210 7778 3226 7842
rect 3290 7778 3432 7842
rect 3496 7778 3512 7842
rect 3576 7778 3592 7842
rect 3656 7778 3672 7842
rect 3736 7778 3752 7842
rect 3816 7778 3832 7842
rect 3896 7778 4038 7842
rect 4102 7778 4118 7842
rect 4182 7778 4198 7842
rect 4262 7778 4278 7842
rect 4342 7778 4358 7842
rect 4422 7778 4438 7842
rect 4502 7778 4644 7842
rect 4708 7778 4724 7842
rect 4788 7778 4804 7842
rect 4868 7778 4884 7842
rect 4948 7778 4964 7842
rect 5028 7778 5044 7842
rect 5108 7778 5250 7842
rect 5314 7778 5330 7842
rect 5394 7778 5410 7842
rect 5474 7778 5490 7842
rect 5554 7778 5570 7842
rect 5634 7778 5650 7842
rect 5714 7778 5818 7842
rect 904 7776 5818 7778
<< labels >>
flabel pwell 3646 8848 3682 8882 0 FreeSans 160 0 0 0 SUB
port 1 nsew
flabel pwell 2436 8192 2462 8224 0 FreeSans 160 0 0 0 x1[4].SUB
flabel metal4 2378 8526 2404 8558 0 FreeSans 320 0 0 0 x1[4].CBOT
flabel metal4 2496 7936 2522 7968 0 FreeSans 320 0 0 0 x1[4].CTOP
flabel pwell 2436 9352 2462 9384 0 FreeSans 160 0 0 0 x1[5].SUB
flabel metal4 2378 9686 2404 9718 0 FreeSans 320 0 0 0 x1[5].CBOT
flabel metal4 2496 9096 2522 9128 0 FreeSans 320 0 0 0 x1[5].CTOP
flabel pwell 1830 9352 1856 9384 0 FreeSans 160 0 0 0 x1[3].SUB
flabel metal4 1772 9686 1798 9718 0 FreeSans 320 0 0 0 x1[3].CBOT
flabel metal4 1890 9096 1916 9128 0 FreeSans 320 0 0 0 x1[3].CTOP
flabel pwell 1830 8192 1856 8224 0 FreeSans 160 0 0 0 x1[2].SUB
flabel metal4 1772 8526 1798 8558 0 FreeSans 320 0 0 0 x1[2].CBOT
flabel metal4 1890 7936 1916 7968 0 FreeSans 320 0 0 0 x1[2].CTOP
flabel pwell 1224 9352 1250 9384 0 FreeSans 160 0 0 0 x1[1].SUB
flabel metal4 1166 9686 1192 9718 0 FreeSans 320 0 0 0 x1[1].CBOT
flabel metal4 1284 9096 1310 9128 0 FreeSans 320 0 0 0 x1[1].CTOP
flabel pwell 1224 8192 1250 8224 0 FreeSans 160 0 0 0 x1[0].SUB
flabel metal4 1166 8526 1192 8558 0 FreeSans 320 0 0 0 x1[0].CBOT
flabel metal4 1284 7936 1310 7968 0 FreeSans 320 0 0 0 x1[0].CTOP
flabel pwell 3648 8192 3674 8224 0 FreeSans 160 0 0 0 x1[8].SUB
flabel metal4 3590 8526 3616 8558 0 FreeSans 320 0 0 0 x1[8].CBOT
flabel metal4 3708 7936 3734 7968 0 FreeSans 320 0 0 0 x1[8].CTOP
flabel pwell 3648 9352 3674 9384 0 FreeSans 160 0 0 0 x1[9].SUB
flabel metal4 3590 9686 3616 9718 0 FreeSans 320 0 0 0 x1[9].CBOT
flabel metal4 3708 9096 3734 9128 0 FreeSans 320 0 0 0 x1[9].CTOP
flabel pwell 3042 8192 3068 8224 0 FreeSans 160 0 0 0 x1[6].SUB
flabel metal4 2984 8526 3010 8558 0 FreeSans 320 0 0 0 x1[6].CBOT
flabel metal4 3102 7936 3128 7968 0 FreeSans 320 0 0 0 x1[6].CTOP
flabel pwell 3042 9352 3068 9384 0 FreeSans 160 0 0 0 x1[7].SUB
flabel metal4 2984 9686 3010 9718 0 FreeSans 320 0 0 0 x1[7].CBOT
flabel metal4 3102 9096 3128 9128 0 FreeSans 320 0 0 0 x1[7].CTOP
flabel pwell 5466 8192 5492 8224 0 FreeSans 160 0 0 0 x1[14].SUB
flabel metal4 5408 8526 5434 8558 0 FreeSans 320 0 0 0 x1[14].CBOT
flabel metal4 5526 7936 5552 7968 0 FreeSans 320 0 0 0 x1[14].CTOP
flabel pwell 5466 9352 5492 9384 0 FreeSans 160 0 0 0 x1[15].SUB
flabel metal4 5408 9686 5434 9718 0 FreeSans 320 0 0 0 x1[15].CBOT
flabel metal4 5526 9096 5552 9128 0 FreeSans 320 0 0 0 x1[15].CTOP
flabel pwell 4860 8192 4886 8224 0 FreeSans 160 0 0 0 x1[12].SUB
flabel metal4 4802 8526 4828 8558 0 FreeSans 320 0 0 0 x1[12].CBOT
flabel metal4 4920 7936 4946 7968 0 FreeSans 320 0 0 0 x1[12].CTOP
flabel pwell 4860 9352 4886 9384 0 FreeSans 160 0 0 0 x1[13].SUB
flabel metal4 4802 9686 4828 9718 0 FreeSans 320 0 0 0 x1[13].CBOT
flabel metal4 4920 9096 4946 9128 0 FreeSans 320 0 0 0 x1[13].CTOP
flabel pwell 4254 8192 4280 8224 0 FreeSans 160 0 0 0 x1[10].SUB
flabel metal4 4196 8526 4222 8558 0 FreeSans 320 0 0 0 x1[10].CBOT
flabel metal4 4314 7936 4340 7968 0 FreeSans 320 0 0 0 x1[10].CTOP
flabel pwell 4254 9352 4280 9384 0 FreeSans 160 0 0 0 x1[11].SUB
flabel metal4 4196 9686 4222 9718 0 FreeSans 320 0 0 0 x1[11].CBOT
flabel metal4 4314 9096 4340 9128 0 FreeSans 320 0 0 0 x1[11].CTOP
<< end >>
