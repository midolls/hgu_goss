magic
tech sky130A
magscale 1 2
timestamp 1701054579
<< nwell >>
rect -3314 8582 -3207 8954
rect -3419 7301 -3156 7964
<< metal1 >>
rect -8588 14613 -8582 14665
rect -8530 14663 -8524 14665
rect -8530 14616 -8469 14663
rect -8530 14613 -8524 14616
rect -50095 10792 -49983 10799
rect -50095 10690 -50089 10792
rect -49990 10690 -49983 10792
rect -50095 10685 -49983 10690
rect -50079 9932 -49998 10685
rect -6380 10156 -6374 10208
rect -6322 10156 -6316 10208
rect -972 9906 -966 9916
rect -6221 9876 -966 9906
rect -972 9864 -966 9876
rect -914 9906 -908 9916
rect -914 9876 -899 9906
rect -914 9864 -908 9876
rect -1065 9836 -1059 9846
rect -6221 9806 -1059 9836
rect -1065 9794 -1059 9806
rect -1007 9836 -1001 9846
rect -1007 9806 -899 9836
rect -1007 9794 -1001 9806
rect -1527 9766 -1521 9778
rect -6221 9736 -1521 9766
rect -1527 9726 -1521 9736
rect -1469 9766 -1463 9778
rect -1469 9736 -899 9766
rect -1469 9726 -1463 9736
rect -1805 9697 -1799 9708
rect -2399 9696 -1799 9697
rect -6221 9666 -1799 9696
rect -1805 9656 -1799 9666
rect -1747 9697 -1741 9708
rect -1747 9696 -1109 9697
rect -1747 9666 -899 9696
rect -1747 9656 -1741 9666
rect -1655 9627 -1649 9638
rect -6221 9597 -1649 9627
rect -1655 9586 -1649 9597
rect -1597 9627 -1591 9638
rect -1597 9597 -899 9627
rect -1597 9586 -1591 9597
rect -2319 9557 -2313 9568
rect -6221 9527 -2313 9557
rect -2319 9516 -2313 9527
rect -2261 9557 -2255 9568
rect -2261 9527 -899 9557
rect -2261 9516 -2255 9527
rect -1247 9488 -1241 9498
rect -6221 9458 -1241 9488
rect -1247 9446 -1241 9458
rect -1189 9488 -1183 9498
rect -1189 9458 -899 9488
rect -1189 9446 -1183 9458
rect -3256 9418 -3250 9429
rect -6221 9388 -3250 9418
rect -3256 9377 -3250 9388
rect -3198 9418 -3192 9429
rect -3198 9388 -899 9418
rect -3198 9377 -3192 9388
rect -3343 9348 -3337 9358
rect -6221 9318 -3337 9348
rect -3343 9306 -3337 9318
rect -3285 9348 -3279 9358
rect -3285 9318 -899 9348
rect -3285 9306 -3279 9318
rect -3705 9278 -3699 9290
rect -6221 9248 -3699 9278
rect -3705 9238 -3699 9248
rect -3647 9278 -3641 9290
rect -3647 9248 -899 9278
rect -3647 9238 -3641 9248
rect -3983 9209 -3977 9220
rect -6221 9179 -3977 9209
rect -3983 9168 -3977 9179
rect -3925 9209 -3919 9220
rect -3925 9179 -899 9209
rect -3925 9168 -3919 9179
rect -3833 9139 -3827 9150
rect -6221 9109 -3827 9139
rect -3833 9098 -3827 9109
rect -3775 9139 -3769 9150
rect -3775 9109 -899 9139
rect -3775 9098 -3769 9109
rect -4497 9069 -4491 9080
rect -6221 9039 -4491 9069
rect -4497 9028 -4491 9039
rect -4439 9069 -4433 9080
rect -4439 9039 -899 9069
rect -4439 9028 -4433 9039
rect -3430 9000 -3424 9010
rect -6221 8970 -3424 9000
rect -3430 8958 -3424 8970
rect -3372 9000 -3366 9010
rect -3372 8970 -899 9000
rect -3372 8958 -3366 8970
rect -8587 8776 -8581 8828
rect -8529 8814 -8523 8828
rect -3356 8816 -3180 8912
rect -8529 8786 -5992 8814
rect -8529 8776 -8523 8786
rect -6020 6724 -5992 8786
rect -3469 8176 -3172 8368
rect -3465 7536 -3168 7728
rect -3443 6992 -3182 7088
rect -5419 6783 -5413 6799
rect -5444 6748 -5413 6783
rect -5419 6747 -5413 6748
rect -5361 6783 -5355 6799
rect -5361 6748 142 6783
rect -5361 6747 -5355 6748
rect -6033 6672 -6027 6724
rect -5975 6672 -5969 6724
rect -1336 6590 -1330 6642
rect -1278 6631 -1272 6642
rect -1150 6631 -1144 6641
rect -1278 6601 -1144 6631
rect -1278 6590 -1272 6601
rect -1150 6589 -1144 6601
rect -1092 6589 -1086 6641
rect -1611 6521 -1605 6573
rect -1553 6561 -1547 6573
rect -1236 6561 -1230 6571
rect -1553 6531 -1230 6561
rect -1553 6521 -1547 6531
rect -1236 6519 -1230 6531
rect -1178 6519 -1172 6571
rect -1886 6451 -1880 6503
rect -1828 6491 -1822 6503
rect -1323 6491 -1317 6502
rect -1828 6461 -1317 6491
rect -1828 6451 -1822 6461
rect -1323 6450 -1317 6461
rect -1265 6450 -1259 6502
rect -2428 6381 -2422 6433
rect -2370 6422 -2364 6433
rect -1409 6422 -1403 6432
rect -2370 6392 -1403 6422
rect -2370 6381 -2364 6392
rect -1409 6380 -1403 6392
rect -1351 6380 -1345 6432
rect -2993 6312 -2987 6364
rect -2935 6352 -2929 6364
rect -1496 6352 -1490 6363
rect -2935 6322 -1490 6352
rect -2935 6312 -2929 6322
rect -1496 6311 -1490 6322
rect -1438 6311 -1432 6363
rect -3257 6242 -3251 6294
rect -3199 6283 -3193 6294
rect -1582 6283 -1576 6293
rect -3199 6253 -1576 6283
rect -3199 6242 -3193 6253
rect -1582 6241 -1576 6253
rect -1524 6241 -1518 6293
rect -3345 6172 -3339 6224
rect -3287 6213 -3281 6224
rect -1668 6213 -1662 6223
rect -3287 6183 -1662 6213
rect -3287 6172 -3281 6183
rect -1668 6171 -1662 6183
rect -1610 6171 -1604 6223
rect -3519 6102 -3513 6154
rect -3461 6143 -3455 6154
rect -1754 6143 -1748 6153
rect -3461 6113 -1748 6143
rect -3461 6102 -3455 6113
rect -1754 6101 -1748 6113
rect -1696 6101 -1690 6153
rect -3792 6033 -3786 6085
rect -3734 6073 -3728 6085
rect -1841 6073 -1835 6084
rect -3734 6043 -1835 6073
rect -3734 6033 -3728 6043
rect -1841 6032 -1835 6043
rect -1783 6032 -1777 6084
rect -4071 5963 -4065 6015
rect -4013 6004 -4007 6015
rect -1927 6004 -1921 6014
rect -4013 5974 -1921 6004
rect -4013 5963 -4007 5974
rect -1927 5962 -1921 5974
rect -1869 5962 -1863 6014
rect -4618 5894 -4612 5946
rect -4560 5934 -4554 5946
rect -2013 5934 -2007 5944
rect -4560 5904 -2007 5934
rect -4560 5894 -4554 5904
rect -2013 5892 -2007 5904
rect -1955 5892 -1949 5944
rect -5169 5824 -5163 5876
rect -5111 5864 -5105 5876
rect -2100 5864 -2094 5875
rect -5111 5834 -2094 5864
rect -5111 5824 -5105 5834
rect -2100 5823 -2094 5834
rect -2042 5823 -2036 5875
rect -50079 4516 -49998 5205
rect -50094 4511 -49982 4516
rect -50094 4409 -50087 4511
rect -49988 4409 -49982 4511
rect -50094 4402 -49982 4409
rect -1374 972 -1368 1024
rect -1316 1014 -1310 1024
rect -1316 984 14462 1014
rect -1316 972 -1310 984
rect -826 902 -820 954
rect -768 944 -762 954
rect -768 914 14462 944
rect -768 902 -762 914
rect -559 833 -553 885
rect -501 874 -495 885
rect -501 844 14462 874
rect -501 833 -495 844
rect -273 763 -267 815
rect -215 805 -209 815
rect -215 775 14462 805
rect -215 763 -209 775
rect -46 694 -40 746
rect 12 735 18 746
rect 12 705 14462 735
rect 12 694 18 705
rect 90 624 96 676
rect 148 666 154 676
rect 148 636 14462 666
rect 148 624 154 636
rect 426 554 432 606
rect 484 596 490 606
rect 484 566 14462 596
rect 484 554 490 566
rect 972 484 978 536
rect 1030 526 1036 536
rect 1030 496 14462 526
rect 1030 484 1036 496
rect 1519 415 1525 467
rect 1577 456 1583 467
rect 1577 426 14462 456
rect 1577 415 1583 426
rect 1805 345 1811 397
rect 1863 387 1869 397
rect 1863 357 14462 387
rect 1863 345 1869 357
rect 2071 275 2077 327
rect 2129 317 2135 327
rect 2129 287 14462 317
rect 2129 275 2135 287
rect 2316 206 2322 258
rect 2374 247 2380 258
rect 2374 217 14462 247
rect 2374 206 2380 217
rect 2454 137 2460 189
rect 2512 178 2518 189
rect 2512 148 14462 178
rect 2512 137 2518 148
rect -186 -1922 -180 -1910
rect -2431 -1952 -180 -1922
rect -186 -1962 -180 -1952
rect -128 -1922 -122 -1910
rect -128 -1952 2620 -1922
rect -128 -1962 -122 -1952
rect -1258 -1991 -1252 -1980
rect -2431 -2021 -1252 -1991
rect -1258 -2032 -1252 -2021
rect -1200 -1991 -1194 -1980
rect -1200 -2021 2620 -1991
rect -1200 -2032 -1194 -2021
rect -594 -2061 -588 -2050
rect -2431 -2091 -588 -2061
rect -594 -2102 -588 -2091
rect -536 -2061 -530 -2050
rect -536 -2091 2620 -2061
rect -536 -2102 -530 -2091
rect -744 -2131 -738 -2120
rect -2431 -2161 -738 -2131
rect -744 -2172 -738 -2161
rect -686 -2131 -680 -2120
rect -686 -2161 2620 -2131
rect -686 -2172 -680 -2161
rect -466 -2200 -460 -2190
rect -2431 -2230 -460 -2200
rect -466 -2242 -460 -2230
rect -408 -2200 -402 -2190
rect -408 -2230 2620 -2200
rect -408 -2242 -402 -2230
rect -44 -2270 -38 -2258
rect -2431 -2300 -38 -2270
rect -44 -2310 -38 -2300
rect 14 -2270 20 -2258
rect 14 -2300 2620 -2270
rect 14 -2310 20 -2300
rect 90 -2340 96 -2328
rect -2431 -2370 96 -2340
rect 90 -2380 96 -2370
rect 148 -2340 154 -2328
rect 148 -2370 2620 -2340
rect 148 -2380 154 -2370
rect 2168 -2410 2174 -2398
rect -2431 -2440 2174 -2410
rect 2168 -2450 2174 -2440
rect 2226 -2410 2232 -2398
rect 2226 -2440 2620 -2410
rect 2226 -2450 2232 -2440
rect 1096 -2479 1102 -2468
rect -2431 -2509 1102 -2479
rect 1096 -2520 1102 -2509
rect 1154 -2479 1160 -2468
rect 1154 -2509 2620 -2479
rect 1154 -2520 1160 -2509
rect 1760 -2549 1766 -2538
rect -2431 -2579 1766 -2549
rect 1760 -2590 1766 -2579
rect 1818 -2549 1824 -2538
rect 1818 -2579 2620 -2549
rect 1818 -2590 1824 -2579
rect 1610 -2618 1616 -2608
rect -2431 -2648 1616 -2618
rect 1016 -2649 1616 -2648
rect 1610 -2660 1616 -2649
rect 1668 -2618 1674 -2608
rect 1668 -2648 2620 -2618
rect 1668 -2649 2306 -2648
rect 1668 -2660 1674 -2649
rect 1888 -2688 1894 -2678
rect -2431 -2718 1894 -2688
rect 1888 -2730 1894 -2718
rect 1946 -2688 1952 -2678
rect 1946 -2718 2620 -2688
rect 1946 -2730 1952 -2718
rect 2315 -2758 2321 -2746
rect -2431 -2788 2321 -2758
rect 2315 -2798 2321 -2788
rect 2373 -2758 2379 -2746
rect 2373 -2788 2620 -2758
rect 2373 -2798 2379 -2788
rect 2459 -2828 2465 -2816
rect -2432 -2858 2465 -2828
rect 2459 -2868 2465 -2858
rect 2517 -2828 2523 -2816
rect 2517 -2858 2619 -2828
rect 2517 -2868 2523 -2858
<< via1 >>
rect -8582 14613 -8530 14665
rect -50089 10690 -49990 10792
rect -6374 10156 -6322 10208
rect -966 9864 -914 9916
rect -1059 9794 -1007 9846
rect -1521 9726 -1469 9778
rect -1799 9656 -1747 9708
rect -1649 9586 -1597 9638
rect -2313 9516 -2261 9568
rect -1241 9446 -1189 9498
rect -3250 9377 -3198 9429
rect -3337 9306 -3285 9358
rect -3699 9238 -3647 9290
rect -3977 9168 -3925 9220
rect -3827 9098 -3775 9150
rect -4491 9028 -4439 9080
rect -3424 8958 -3372 9010
rect -8581 8776 -8529 8828
rect -5413 6747 -5361 6799
rect -6027 6672 -5975 6724
rect -1330 6590 -1278 6642
rect -1144 6589 -1092 6641
rect -1605 6521 -1553 6573
rect -1230 6519 -1178 6571
rect -1880 6451 -1828 6503
rect -1317 6450 -1265 6502
rect -2422 6381 -2370 6433
rect -1403 6380 -1351 6432
rect -2987 6312 -2935 6364
rect -1490 6311 -1438 6363
rect -3251 6242 -3199 6294
rect -1576 6241 -1524 6293
rect -3339 6172 -3287 6224
rect -1662 6171 -1610 6223
rect -3513 6102 -3461 6154
rect -1748 6101 -1696 6153
rect -3786 6033 -3734 6085
rect -1835 6032 -1783 6084
rect -4065 5963 -4013 6015
rect -1921 5962 -1869 6014
rect -4612 5894 -4560 5946
rect -2007 5892 -1955 5944
rect -5163 5824 -5111 5876
rect -2094 5823 -2042 5875
rect -50087 4409 -49988 4511
rect -1368 972 -1316 1024
rect -820 902 -768 954
rect -553 833 -501 885
rect -267 763 -215 815
rect -40 694 12 746
rect 96 624 148 676
rect 432 554 484 606
rect 978 484 1030 536
rect 1525 415 1577 467
rect 1811 345 1863 397
rect 2077 275 2129 327
rect 2322 206 2374 258
rect 2460 137 2512 189
rect -180 -1962 -128 -1910
rect -1252 -2032 -1200 -1980
rect -588 -2102 -536 -2050
rect -738 -2172 -686 -2120
rect -460 -2242 -408 -2190
rect -38 -2310 14 -2258
rect 96 -2380 148 -2328
rect 2174 -2450 2226 -2398
rect 1102 -2520 1154 -2468
rect 1766 -2590 1818 -2538
rect 1616 -2660 1668 -2608
rect 1894 -2730 1946 -2678
rect 2321 -2798 2373 -2746
rect 2465 -2868 2517 -2816
<< metal2 >>
rect -8588 14613 -8582 14665
rect -8530 14613 -8524 14665
rect -50109 10801 -49970 10811
rect -50109 10680 -50099 10801
rect -49979 10680 -49970 10801
rect -50109 10670 -49970 10680
rect -8574 8828 -8546 14613
rect -6380 10156 -6374 10208
rect -6322 10156 -6316 10208
rect -8587 8776 -8581 8828
rect -8529 8776 -8523 8828
rect -6360 8739 -6332 10156
rect -972 9864 -966 9916
rect -914 9864 -908 9916
rect -1065 9794 -1059 9846
rect -1007 9794 -1001 9846
rect -1527 9726 -1521 9778
rect -1469 9726 -1463 9778
rect -1805 9656 -1799 9708
rect -1747 9656 -1741 9708
rect -2319 9516 -2313 9568
rect -2261 9516 -2255 9568
rect -3256 9377 -3250 9429
rect -3198 9377 -3192 9429
rect -3343 9306 -3337 9358
rect -3285 9306 -3279 9358
rect -3705 9238 -3699 9290
rect -3647 9238 -3641 9290
rect -3983 9168 -3977 9220
rect -3925 9168 -3919 9220
rect -4497 9028 -4491 9080
rect -4439 9028 -4433 9080
rect -4486 8944 -4445 9028
rect -3967 8944 -3926 9168
rect -3833 9098 -3827 9150
rect -3775 9098 -3769 9150
rect -3823 8944 -3782 9098
rect -3691 8944 -3650 9238
rect -3430 8958 -3424 9010
rect -3372 8958 -3366 9010
rect -3413 8944 -3372 8958
rect -5419 6747 -5413 6799
rect -5361 6747 -5355 6799
rect -6033 6672 -6027 6724
rect -5975 6672 -5969 6724
rect -5157 5876 -5115 6958
rect -4608 5946 -4566 6953
rect -4060 6015 -4018 6955
rect -3780 6085 -3738 6956
rect -3508 6154 -3466 6952
rect -3334 6224 -3292 9306
rect -3245 6294 -3203 9377
rect -2308 8944 -2267 9516
rect -1789 8944 -1748 9656
rect -1655 9586 -1649 9638
rect -1597 9586 -1591 9638
rect -1645 8944 -1604 9586
rect -1513 8944 -1472 9726
rect -1247 9446 -1241 9498
rect -1189 9446 -1183 9498
rect -1235 8944 -1194 9446
rect -2981 6364 -2939 6949
rect -2417 6433 -2375 6954
rect -1874 6503 -1832 6957
rect -1600 6573 -1558 6957
rect -1325 6642 -1283 6965
rect -1336 6590 -1330 6642
rect -1278 6590 -1272 6642
rect -1150 6589 -1144 6641
rect -1092 6589 -1086 6641
rect -1611 6521 -1605 6573
rect -1553 6521 -1547 6573
rect -1236 6519 -1230 6571
rect -1178 6519 -1172 6571
rect -1886 6451 -1880 6503
rect -1828 6451 -1822 6503
rect -1323 6450 -1317 6502
rect -1265 6450 -1259 6502
rect -2428 6381 -2422 6433
rect -2370 6381 -2364 6433
rect -1409 6380 -1403 6432
rect -1351 6380 -1345 6432
rect -2993 6312 -2987 6364
rect -2935 6312 -2929 6364
rect -1496 6311 -1490 6363
rect -1438 6311 -1432 6363
rect -3257 6242 -3251 6294
rect -3199 6242 -3193 6294
rect -1582 6241 -1576 6293
rect -1524 6241 -1518 6293
rect -3345 6172 -3339 6224
rect -3287 6172 -3281 6224
rect -1668 6171 -1662 6223
rect -1610 6171 -1604 6223
rect -3519 6102 -3513 6154
rect -3461 6102 -3455 6154
rect -1754 6101 -1748 6153
rect -1696 6101 -1690 6153
rect -3792 6033 -3786 6085
rect -3734 6033 -3728 6085
rect -1841 6032 -1835 6084
rect -1783 6032 -1777 6084
rect -4071 5963 -4065 6015
rect -4013 5963 -4007 6015
rect -1927 5962 -1921 6014
rect -1869 5962 -1863 6014
rect -4618 5894 -4612 5946
rect -4560 5894 -4554 5946
rect -2013 5892 -2007 5944
rect -1955 5892 -1949 5944
rect -5169 5824 -5163 5876
rect -5111 5824 -5105 5876
rect -2100 5823 -2094 5875
rect -2042 5823 -2036 5875
rect -2084 5715 -2042 5823
rect -2002 5715 -1960 5892
rect -1918 5715 -1876 5962
rect -1830 5715 -1788 6032
rect -1743 5715 -1701 6101
rect -1657 5715 -1615 6171
rect -1571 5715 -1529 6241
rect -1484 5715 -1442 6311
rect -1398 5715 -1356 6380
rect -1312 5715 -1270 6450
rect -1225 5715 -1183 6519
rect -1140 5715 -1098 6589
rect -1053 5716 -1011 9794
rect -966 5716 -924 9864
rect -50107 4521 -49968 4531
rect -50107 4400 -50098 4521
rect -49978 4400 -49968 4521
rect -50107 4390 -49968 4400
rect -1374 972 -1368 1024
rect -1316 972 -1310 1024
rect -1924 138 -1882 906
rect -1362 93 -1320 972
rect -826 902 -820 954
rect -768 902 -762 954
rect -816 93 -774 902
rect -559 833 -553 885
rect -501 833 -495 885
rect -548 93 -506 833
rect -273 763 -267 815
rect -215 763 -209 815
rect -261 93 -219 763
rect -46 694 -40 746
rect 12 694 18 746
rect -1247 -1980 -1206 -1718
rect -1258 -2032 -1252 -1980
rect -1200 -2032 -1194 -1980
rect -728 -2120 -687 -1838
rect -584 -2050 -543 -1791
rect -594 -2102 -588 -2050
rect -536 -2102 -530 -2050
rect -744 -2172 -738 -2120
rect -686 -2172 -680 -2120
rect -452 -2190 -411 -1903
rect -186 -1962 -180 -1910
rect -128 -1962 -122 -1910
rect -466 -2242 -460 -2190
rect -408 -2242 -402 -2190
rect -35 -2258 7 694
rect 90 624 96 676
rect 148 624 154 676
rect -44 -2310 -38 -2258
rect 14 -2310 20 -2258
rect 101 -2328 143 624
rect 426 554 432 606
rect 484 554 490 606
rect 438 93 480 554
rect 972 484 978 536
rect 1030 484 1036 536
rect 984 93 1026 484
rect 1519 415 1525 467
rect 1577 415 1583 467
rect 1530 93 1572 415
rect 1805 345 1811 397
rect 1863 345 1869 397
rect 1817 93 1859 345
rect 2071 275 2077 327
rect 2129 275 2135 327
rect 2082 93 2124 275
rect 2316 206 2322 258
rect 2374 206 2380 258
rect 90 -2380 96 -2328
rect 148 -2380 154 -2328
rect 1107 -2468 1148 -1625
rect 1096 -2520 1102 -2468
rect 1154 -2520 1160 -2468
rect 1626 -2608 1667 -1766
rect 1770 -2538 1811 -1680
rect 1760 -2590 1766 -2538
rect 1818 -2590 1824 -2538
rect 1610 -2660 1616 -2608
rect 1668 -2660 1674 -2608
rect 1902 -2678 1943 -1820
rect 2180 -2398 2221 -1892
rect 2168 -2450 2174 -2398
rect 2226 -2450 2232 -2398
rect 1888 -2730 1894 -2678
rect 1946 -2730 1952 -2678
rect 2327 -2746 2369 206
rect 2454 137 2460 189
rect 2512 137 2518 189
rect 2315 -2798 2321 -2746
rect 2373 -2798 2379 -2746
rect 2465 -2816 2507 137
rect 2459 -2868 2465 -2816
rect 2517 -2868 2523 -2816
<< via2 >>
rect -50099 10792 -49979 10801
rect -50099 10690 -50089 10792
rect -50089 10690 -49990 10792
rect -49990 10690 -49979 10792
rect -50099 10680 -49979 10690
rect -50098 4511 -49978 4521
rect -50098 4409 -50087 4511
rect -50087 4409 -49988 4511
rect -49988 4409 -49978 4511
rect -50098 4400 -49978 4409
<< metal3 >>
rect -50133 10828 -49945 10835
rect -50133 10652 -50127 10828
rect -49950 10652 -49945 10828
rect -50133 10646 -49945 10652
rect -9304 7723 -9294 7791
rect -9230 7787 -9220 7791
rect -9230 7727 -8766 7787
rect -9230 7723 -9220 7727
rect -9304 7405 -9294 7473
rect -9230 7469 -9220 7473
rect -9230 7409 -8766 7469
rect -9230 7405 -9220 7409
rect -50132 4549 -49944 4555
rect -50132 4373 -50127 4549
rect -49950 4373 -49944 4549
rect -50132 4366 -49944 4373
<< via3 >>
rect -50127 10801 -49950 10828
rect -50127 10680 -50099 10801
rect -50099 10680 -49979 10801
rect -49979 10680 -49950 10801
rect -50127 10652 -49950 10680
rect -9294 7723 -9230 7791
rect -9294 7405 -9230 7473
rect -50127 4521 -49950 4549
rect -50127 4400 -50098 4521
rect -50098 4400 -49978 4521
rect -49978 4400 -49950 4521
rect -50127 4373 -49950 4400
<< metal4 >>
rect -50084 12269 -49569 12337
rect -50084 10859 -50006 12269
rect -9312 10856 -9208 10902
rect -9312 7791 -9209 10620
rect -5368 10334 -4404 10340
rect -9312 7723 -9294 7791
rect -9230 7723 -9209 7791
rect -9312 7712 -9209 7723
rect -5778 10155 -4404 10334
rect -5778 10063 -5590 10155
rect -5400 10153 -4404 10155
rect -5400 10063 -5196 10153
rect -5778 10061 -5196 10063
rect -5006 10151 -4404 10153
rect -5006 10061 -4789 10151
rect -5778 10059 -4789 10061
rect -4599 10059 -4404 10151
rect -5778 8895 -4404 10059
rect -3193 10143 -2229 10302
rect -3193 10051 -3064 10143
rect -2874 10139 -2229 10143
rect -2874 10051 -2638 10139
rect -3193 10047 -2638 10051
rect -2448 10047 -2229 10139
rect -5778 8889 -4814 8895
rect -9312 7473 -9209 7483
rect -9312 7405 -9294 7473
rect -9230 7405 -9209 7473
rect -9312 4676 -9209 7405
rect -5778 6995 -5366 8889
rect -3193 8858 -2229 10047
rect -6166 5674 -5884 6314
rect -4322 5674 -3345 7099
rect -1193 6988 -721 8917
rect -6166 5380 -2607 5674
rect -6166 5376 -5884 5380
rect -9312 4580 -9208 4676
rect -50084 2927 -50006 4342
rect -50084 2859 -49569 2927
<< via4 >>
rect -50157 10828 -49920 10859
rect -50157 10652 -50127 10828
rect -50127 10652 -49950 10828
rect -49950 10652 -49920 10828
rect -50157 10623 -49920 10652
rect -9380 10620 -9144 10856
rect -50157 4549 -49920 4578
rect -50157 4373 -50127 4549
rect -50127 4373 -49950 4549
rect -49950 4373 -49920 4549
rect -50157 4342 -49920 4373
rect -9380 4344 -9144 4580
<< metal5 >>
rect -50203 10903 -49852 10904
rect -50203 10902 -49437 10903
rect -50203 10859 -9105 10902
rect -50203 10623 -50157 10859
rect -49920 10856 -9105 10859
rect -49920 10623 -9380 10856
rect -50203 10620 -9380 10623
rect -9144 10620 -9105 10856
rect -50203 10570 -9105 10620
rect -50137 10569 -49437 10570
rect -50202 4580 -9105 4626
rect -50202 4578 -9380 4580
rect -50202 4342 -50157 4578
rect -49920 4344 -9380 4578
rect -9144 4344 -9105 4580
rect -49920 4342 -9105 4344
rect -50202 4294 -9105 4342
rect -50202 4292 -49508 4294
use hgu_cdac_half  hgu_cdac_half_0
timestamp 1700938627
transform 1 0 -49110 0 -1 6793
box -459 -645 39606 6322
use hgu_cdac_half  hgu_cdac_half_1
timestamp 1700938627
transform 1 0 -49110 0 1 8403
box -459 -645 39606 6322
use hgu_cdac_sw_buffer  hgu_cdac_sw_buffer_0
timestamp 1699539897
transform -1 0 -337 0 -1 -2647
box -270 -2798 1830 -714
use hgu_cdac_sw_buffer  hgu_cdac_sw_buffer_1
timestamp 1699539897
transform -1 0 2017 0 -1 -2643
box -270 -2798 1830 -714
use hgu_cdac_sw_buffer  hgu_cdac_sw_buffer_2
timestamp 1699539897
transform -1 0 -1398 0 1 9721
box -270 -2798 1830 -714
use hgu_cdac_sw_buffer  hgu_cdac_sw_buffer_3
timestamp 1699539897
transform -1 0 -3576 0 1 9720
box -270 -2798 1830 -714
use hgu_comp_flat  hgu_comp_flat_0
timestamp 1698719859
transform 1 0 -9104 0 1 8167
box 338 -1940 3788 618
use hgu_sarlogic_flat  hgu_sarlogic_flat_0
timestamp 1700302578
transform 1 0 -10800 0 1 2806
box 2064 -1908 31250 13749
use hgu_tah  hgu_tah_0
timestamp 1699832401
transform 1 0 -51706 0 1 4757
box 711 297 1858 5355
use hgu_vgen_vref  hgu_vgen_vref_0
timestamp 1701018915
transform -1 0 -50750 0 1 -30367
box 0 0 22370 76000
<< end >>
