* NGSPICE file created from hgu_cdac_unit_flat.ext - technology: sky130A

.subckt hgu_cdac_unit_flat C1 C0
C0 C1 C0 4.38f
C1 C1 VSUBS 1.24f
.ends

