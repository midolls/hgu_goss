magic
tech sky130A
timestamp 1698674462
<< end >>
