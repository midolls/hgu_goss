magic
tech sky130A
magscale 1 2
timestamp 1698843163
<< error_s >>
rect 298 981 333 1015
rect 299 962 333 981
rect 129 913 187 919
rect 129 879 141 913
rect 129 873 187 879
rect 129 719 187 725
rect 129 685 141 719
rect 129 679 187 685
rect 318 583 333 962
rect 352 928 387 962
rect 667 928 702 962
rect 352 583 386 928
rect 668 909 702 928
rect 498 860 556 866
rect 498 826 510 860
rect 498 820 556 826
rect 498 666 556 672
rect 498 632 510 666
rect 498 626 556 632
rect 352 549 367 583
rect 687 530 702 909
rect 721 875 756 909
rect 1036 875 1071 909
rect 721 530 755 875
rect 1037 856 1071 875
rect 867 807 925 813
rect 867 773 879 807
rect 867 767 925 773
rect 867 613 925 619
rect 867 579 879 613
rect 867 573 925 579
rect 721 496 736 530
rect 1056 477 1071 856
rect 1090 822 1125 856
rect 1405 822 1440 856
rect 1090 477 1124 822
rect 1406 803 1440 822
rect 1236 754 1294 760
rect 1236 720 1248 754
rect 1236 714 1294 720
rect 1236 560 1294 566
rect 1236 526 1248 560
rect 1236 520 1294 526
rect 1090 443 1105 477
rect 1425 424 1440 803
rect 1459 769 1494 803
rect 1774 769 1809 803
rect 1459 424 1493 769
rect 1775 750 1809 769
rect 1605 701 1663 707
rect 1605 667 1617 701
rect 1605 661 1663 667
rect 1605 507 1663 513
rect 1605 473 1617 507
rect 1605 467 1663 473
rect 1459 390 1474 424
rect 1794 371 1809 750
rect 1828 716 1863 750
rect 2143 716 2178 750
rect 1828 371 1862 716
rect 2144 697 2178 716
rect 1974 648 2032 654
rect 1974 614 1986 648
rect 1974 608 2032 614
rect 1974 454 2032 460
rect 1974 420 1986 454
rect 1974 414 2032 420
rect 1828 337 1843 371
rect 2163 318 2178 697
rect 2197 663 2232 697
rect 2512 663 2547 697
rect 2197 318 2231 663
rect 2513 644 2547 663
rect 2343 595 2401 601
rect 2343 561 2355 595
rect 2343 555 2401 561
rect 2343 401 2401 407
rect 2343 367 2355 401
rect 2343 361 2401 367
rect 2197 284 2212 318
rect 2532 265 2547 644
rect 2566 610 2601 644
rect 2881 610 2916 644
rect 2566 265 2600 610
rect 2882 591 2916 610
rect 2712 542 2770 548
rect 2712 508 2724 542
rect 2712 502 2770 508
rect 2712 348 2770 354
rect 2712 314 2724 348
rect 2712 308 2770 314
rect 2566 231 2581 265
rect 2901 212 2916 591
rect 2935 557 2970 591
rect 3250 557 3285 591
rect 2935 212 2969 557
rect 3251 538 3285 557
rect 3081 489 3139 495
rect 3081 455 3093 489
rect 3081 449 3139 455
rect 3081 295 3139 301
rect 3081 261 3093 295
rect 3081 255 3139 261
rect 2935 178 2950 212
rect 3270 159 3285 538
rect 3304 504 3339 538
rect 3619 504 3654 538
rect 3304 159 3338 504
rect 3620 485 3654 504
rect 3450 436 3508 442
rect 3450 402 3462 436
rect 3450 396 3508 402
rect 3450 242 3508 248
rect 3450 208 3462 242
rect 3450 202 3508 208
rect 3304 125 3319 159
rect 3639 106 3654 485
rect 3673 451 3708 485
rect 3988 451 4023 485
rect 3673 106 3707 451
rect 3989 432 4023 451
rect 3819 383 3877 389
rect 3819 349 3831 383
rect 3819 343 3877 349
rect 3819 189 3877 195
rect 3819 155 3831 189
rect 3819 149 3877 155
rect 3673 72 3688 106
rect 4008 53 4023 432
rect 4042 398 4077 432
rect 4357 398 4392 432
rect 4042 53 4076 398
rect 4358 379 4392 398
rect 4188 330 4246 336
rect 4188 296 4200 330
rect 4188 290 4246 296
rect 4188 136 4246 142
rect 4188 102 4200 136
rect 4188 96 4246 102
rect 4042 19 4057 53
rect 4377 0 4392 379
rect 4411 345 4446 379
rect 4726 345 4761 379
rect 4411 0 4445 345
rect 4727 326 4761 345
rect 4557 277 4615 283
rect 4557 243 4569 277
rect 4557 237 4615 243
rect 4557 83 4615 89
rect 4557 49 4569 83
rect 4557 43 4615 49
rect 4411 -34 4426 0
rect 4746 -53 4761 326
rect 4780 292 4815 326
rect 5095 292 5130 326
rect 4780 -53 4814 292
rect 5096 273 5130 292
rect 4926 224 4984 230
rect 4926 190 4938 224
rect 4926 184 4984 190
rect 4926 30 4984 36
rect 4926 -4 4938 30
rect 4926 -10 4984 -4
rect 4780 -87 4795 -53
rect 5115 -106 5130 273
rect 5149 239 5184 273
rect 5464 239 5499 273
rect 5149 -106 5183 239
rect 5465 220 5499 239
rect 5295 171 5353 177
rect 5295 137 5307 171
rect 5295 131 5353 137
rect 5295 -23 5353 -17
rect 5295 -57 5307 -23
rect 5295 -63 5353 -57
rect 5149 -140 5164 -106
rect 5484 -159 5499 220
rect 5518 186 5553 220
rect 5518 -159 5552 186
rect 5664 118 5722 124
rect 5664 84 5676 118
rect 5664 78 5722 84
rect 5664 -76 5722 -70
rect 5664 -110 5676 -76
rect 5664 -116 5722 -110
rect 5518 -193 5533 -159
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
use sky130_fd_pr__nfet_01v8_L7T3GD  XM1
timestamp 0
transform 1 0 158 0 1 799
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_L7T3GD  XM2
timestamp 0
transform 1 0 527 0 1 746
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_L7T3GD  XM3
timestamp 0
transform 1 0 896 0 1 693
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_L7T3GD  XM4
timestamp 0
transform 1 0 1265 0 1 640
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_L7T3GD  XM5
timestamp 0
transform 1 0 1634 0 1 587
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_L7T3GD  XM6
timestamp 0
transform 1 0 2003 0 1 534
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_L7T3GD  XM7
timestamp 0
transform 1 0 2372 0 1 481
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_L7T3GD  XM8
timestamp 0
transform 1 0 2741 0 1 428
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_L7T3GD  XM9
timestamp 0
transform 1 0 3110 0 1 375
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_L7T3GD  XM10
timestamp 0
transform 1 0 3479 0 1 322
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_L7T3GD  XM11
timestamp 0
transform 1 0 3848 0 1 269
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_L7T3GD  XM12
timestamp 0
transform 1 0 4217 0 1 216
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_L7T3GD  XM13
timestamp 0
transform 1 0 4586 0 1 163
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_L7T3GD  XM14
timestamp 0
transform 1 0 4955 0 1 110
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_L7T3GD  XM15
timestamp 0
transform 1 0 5324 0 1 57
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_L7T3GD  XM16
timestamp 0
transform 1 0 5693 0 1 4
box -211 -252 211 252
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 input_stack
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 output_stack
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 VSS
port 2 nsew
<< end >>
