magic
tech sky130A
magscale 1 2
timestamp 1699538049
<< nwell >>
rect 18434 9634 18880 10661
rect 18545 9622 18673 9634
rect 18745 9622 18873 9634
rect 13332 6954 18192 6996
rect 13332 5670 18192 5724
<< psubdiff >>
rect 18473 9040 18593 9041
rect 18473 9006 18501 9040
rect 18535 9007 18593 9040
rect 18627 9007 18685 9041
rect 18719 9007 18778 9041
rect 18812 9007 18842 9041
rect 18535 9006 18842 9007
rect 18473 9005 18842 9006
rect 13370 7581 13399 7615
rect 13433 7581 13491 7615
rect 13525 7581 13583 7615
rect 13617 7581 13675 7615
rect 13709 7581 13767 7615
rect 13801 7581 13859 7615
rect 13893 7581 13951 7615
rect 13985 7581 14043 7615
rect 14077 7581 14135 7615
rect 14169 7581 14226 7615
rect 14260 7581 14319 7615
rect 14353 7581 14411 7615
rect 14445 7581 14503 7615
rect 14537 7581 14595 7615
rect 14629 7581 14687 7615
rect 14721 7581 14779 7615
rect 14813 7581 14871 7615
rect 14905 7581 14963 7615
rect 14997 7581 15055 7615
rect 15089 7581 15147 7615
rect 15181 7581 15239 7615
rect 15273 7581 15331 7615
rect 15365 7581 15423 7615
rect 15457 7581 15515 7615
rect 15549 7581 15607 7615
rect 15641 7581 15699 7615
rect 15733 7581 15791 7615
rect 15825 7581 15883 7615
rect 15917 7581 15975 7615
rect 16009 7581 16067 7615
rect 16101 7581 16159 7615
rect 16193 7581 16251 7615
rect 16285 7581 16343 7615
rect 16377 7581 16435 7615
rect 16469 7581 16527 7615
rect 16561 7581 16619 7615
rect 16653 7581 16711 7615
rect 16745 7581 16803 7615
rect 16837 7581 16895 7615
rect 16929 7581 16987 7615
rect 17021 7581 17079 7615
rect 17113 7581 17171 7615
rect 17205 7581 17263 7615
rect 17297 7581 17355 7615
rect 17389 7581 17447 7615
rect 17481 7581 17539 7615
rect 17573 7581 17631 7615
rect 17665 7581 17723 7615
rect 17757 7581 17815 7615
rect 17849 7581 17907 7615
rect 17941 7581 17999 7615
rect 18033 7581 18091 7615
rect 18125 7581 18154 7615
rect 13370 6316 13399 6350
rect 13433 6316 13491 6350
rect 13525 6316 13583 6350
rect 13617 6316 13675 6350
rect 13709 6316 13767 6350
rect 13801 6316 13859 6350
rect 13893 6316 13951 6350
rect 13985 6316 14043 6350
rect 14077 6316 14135 6350
rect 14169 6316 14227 6350
rect 14261 6316 14319 6350
rect 14353 6316 14411 6350
rect 14445 6316 14503 6350
rect 14537 6316 14595 6350
rect 14629 6316 14687 6350
rect 14721 6316 14779 6350
rect 14813 6316 14871 6350
rect 14905 6316 14964 6350
rect 14998 6316 15055 6350
rect 15089 6316 15147 6350
rect 15181 6316 15239 6350
rect 15273 6316 15332 6350
rect 15366 6316 15423 6350
rect 15457 6316 15515 6350
rect 15549 6316 15607 6350
rect 15641 6316 15699 6350
rect 15733 6316 15791 6350
rect 15825 6316 15883 6350
rect 15917 6316 15975 6350
rect 16009 6316 16067 6350
rect 16101 6316 16159 6350
rect 16193 6316 16251 6350
rect 16285 6316 16343 6350
rect 16377 6316 16435 6350
rect 16469 6316 16526 6350
rect 16560 6316 16618 6350
rect 16652 6316 16711 6350
rect 16745 6316 16803 6350
rect 16837 6316 16895 6350
rect 16929 6316 16986 6350
rect 17020 6316 17079 6350
rect 17113 6316 17170 6350
rect 17204 6316 17263 6350
rect 17297 6316 17355 6350
rect 17389 6316 17447 6350
rect 17481 6316 17539 6350
rect 17573 6316 17631 6350
rect 17665 6316 17723 6350
rect 17757 6316 17815 6350
rect 17849 6316 17907 6350
rect 17941 6316 17999 6350
rect 18033 6316 18091 6350
rect 18125 6316 18154 6350
rect 13370 5049 13399 5083
rect 13433 5049 13491 5083
rect 13525 5049 13583 5083
rect 13617 5049 13675 5083
rect 13709 5049 13767 5083
rect 13801 5049 13859 5083
rect 13893 5049 13951 5083
rect 13985 5049 14043 5083
rect 14077 5049 14135 5083
rect 14169 5049 14227 5083
rect 14261 5049 14319 5083
rect 14353 5049 14411 5083
rect 14445 5049 14503 5083
rect 14537 5049 14595 5083
rect 14629 5049 14687 5083
rect 14721 5049 14779 5083
rect 14813 5049 14871 5083
rect 14905 5049 14963 5083
rect 14997 5049 15055 5083
rect 15089 5049 15147 5083
rect 15181 5049 15239 5083
rect 15273 5049 15331 5083
rect 15365 5049 15423 5083
rect 15457 5049 15515 5083
rect 15549 5049 15607 5083
rect 15641 5049 15699 5083
rect 15733 5049 15791 5083
rect 15825 5049 15883 5083
rect 15917 5049 15975 5083
rect 16009 5049 16067 5083
rect 16101 5049 16159 5083
rect 16193 5049 16251 5083
rect 16285 5049 16343 5083
rect 16377 5049 16435 5083
rect 16469 5049 16527 5083
rect 16561 5049 16619 5083
rect 16653 5049 16711 5083
rect 16745 5049 16803 5083
rect 16837 5049 16895 5083
rect 16929 5049 16987 5083
rect 17021 5049 17079 5083
rect 17113 5049 17171 5083
rect 17205 5049 17263 5083
rect 17297 5049 17355 5083
rect 17389 5049 17447 5083
rect 17481 5049 17539 5083
rect 17573 5049 17631 5083
rect 17665 5049 17723 5083
rect 17757 5049 17815 5083
rect 17849 5049 17907 5083
rect 17941 5049 17999 5083
rect 18033 5049 18091 5083
rect 18125 5049 18154 5083
<< nsubdiff >>
rect 18472 9652 18841 9654
rect 18472 9618 18501 9652
rect 18535 9618 18684 9652
rect 18718 9618 18841 9652
rect 13370 6955 13400 6989
rect 13434 6955 13491 6989
rect 13525 6955 13584 6989
rect 13618 6955 13675 6989
rect 13709 6955 13766 6989
rect 13800 6955 13860 6989
rect 13894 6955 13951 6989
rect 13985 6955 14044 6989
rect 14078 6955 14135 6989
rect 14169 6955 14227 6989
rect 14261 6955 14318 6989
rect 14352 6955 14411 6989
rect 14445 6955 14504 6989
rect 14538 6955 14595 6989
rect 14629 6955 14687 6989
rect 14721 6955 14779 6989
rect 14813 6955 14871 6989
rect 14905 6955 14963 6989
rect 14997 6955 15055 6989
rect 15089 6955 15147 6989
rect 15181 6955 15240 6989
rect 15274 6955 15330 6989
rect 15364 6955 15423 6989
rect 15457 6955 15516 6989
rect 15550 6955 15608 6989
rect 15642 6955 15699 6989
rect 15733 6955 15792 6989
rect 15826 6955 15884 6989
rect 15918 6955 15976 6989
rect 16010 6955 16068 6989
rect 16102 6955 16160 6989
rect 16194 6955 16252 6989
rect 16286 6955 16343 6989
rect 16377 6955 16434 6989
rect 16468 6955 16527 6989
rect 16561 6955 16620 6989
rect 16654 6955 16712 6989
rect 16746 6955 16803 6989
rect 16837 6955 16897 6989
rect 16931 6955 16987 6989
rect 17021 6955 17078 6989
rect 17112 6955 17171 6989
rect 17205 6955 17264 6989
rect 17298 6955 17356 6989
rect 17390 6955 17447 6989
rect 17481 6955 17539 6989
rect 17573 6955 17631 6989
rect 17665 6955 17722 6989
rect 17756 6955 17814 6989
rect 17848 6955 17907 6989
rect 17941 6955 17999 6989
rect 18033 6955 18091 6989
rect 18125 6955 18154 6989
rect 13370 5674 13402 5708
rect 13436 5674 13492 5708
rect 13526 5674 13585 5708
rect 13619 5674 13675 5708
rect 13709 5674 13766 5708
rect 13800 5674 13860 5708
rect 13894 5674 13951 5708
rect 13985 5674 14043 5708
rect 14077 5674 14135 5708
rect 14169 5674 14228 5708
rect 14262 5674 14319 5708
rect 14353 5674 14411 5708
rect 14445 5674 14503 5708
rect 14537 5674 14595 5708
rect 14629 5674 14688 5708
rect 14722 5674 14779 5708
rect 14813 5674 14870 5708
rect 14904 5674 14963 5708
rect 14997 5674 15056 5708
rect 15090 5674 15147 5708
rect 15181 5674 15239 5708
rect 15273 5674 15331 5708
rect 15365 5674 15423 5708
rect 15457 5674 15516 5708
rect 15550 5674 15606 5708
rect 15640 5674 15699 5708
rect 15733 5674 15791 5708
rect 15825 5674 15884 5708
rect 15918 5674 15978 5708
rect 16012 5674 16067 5708
rect 16101 5674 16159 5708
rect 16193 5674 16251 5708
rect 16285 5674 16343 5708
rect 16377 5674 16435 5708
rect 16469 5674 16527 5708
rect 16561 5674 16619 5708
rect 16653 5674 16711 5708
rect 16745 5674 16803 5708
rect 16837 5674 16895 5708
rect 16929 5674 16987 5708
rect 17021 5674 17079 5708
rect 17113 5674 17171 5708
rect 17205 5674 17263 5708
rect 17297 5674 17355 5708
rect 17389 5674 17447 5708
rect 17481 5674 17539 5708
rect 17573 5674 17631 5708
rect 17665 5674 17723 5708
rect 17757 5674 17815 5708
rect 17849 5674 17907 5708
rect 17941 5674 18000 5708
rect 18034 5674 18091 5708
rect 18125 5674 18154 5708
<< psubdiffcont >>
rect 18501 9006 18535 9040
rect 18593 9007 18627 9041
rect 18685 9007 18719 9041
rect 18778 9007 18812 9041
rect 13399 7581 13433 7615
rect 13491 7581 13525 7615
rect 13583 7581 13617 7615
rect 13675 7581 13709 7615
rect 13767 7581 13801 7615
rect 13859 7581 13893 7615
rect 13951 7581 13985 7615
rect 14043 7581 14077 7615
rect 14135 7581 14169 7615
rect 14226 7581 14260 7615
rect 14319 7581 14353 7615
rect 14411 7581 14445 7615
rect 14503 7581 14537 7615
rect 14595 7581 14629 7615
rect 14687 7581 14721 7615
rect 14779 7581 14813 7615
rect 14871 7581 14905 7615
rect 14963 7581 14997 7615
rect 15055 7581 15089 7615
rect 15147 7581 15181 7615
rect 15239 7581 15273 7615
rect 15331 7581 15365 7615
rect 15423 7581 15457 7615
rect 15515 7581 15549 7615
rect 15607 7581 15641 7615
rect 15699 7581 15733 7615
rect 15791 7581 15825 7615
rect 15883 7581 15917 7615
rect 15975 7581 16009 7615
rect 16067 7581 16101 7615
rect 16159 7581 16193 7615
rect 16251 7581 16285 7615
rect 16343 7581 16377 7615
rect 16435 7581 16469 7615
rect 16527 7581 16561 7615
rect 16619 7581 16653 7615
rect 16711 7581 16745 7615
rect 16803 7581 16837 7615
rect 16895 7581 16929 7615
rect 16987 7581 17021 7615
rect 17079 7581 17113 7615
rect 17171 7581 17205 7615
rect 17263 7581 17297 7615
rect 17355 7581 17389 7615
rect 17447 7581 17481 7615
rect 17539 7581 17573 7615
rect 17631 7581 17665 7615
rect 17723 7581 17757 7615
rect 17815 7581 17849 7615
rect 17907 7581 17941 7615
rect 17999 7581 18033 7615
rect 18091 7581 18125 7615
rect 13399 6316 13433 6350
rect 13491 6316 13525 6350
rect 13583 6316 13617 6350
rect 13675 6316 13709 6350
rect 13767 6316 13801 6350
rect 13859 6316 13893 6350
rect 13951 6316 13985 6350
rect 14043 6316 14077 6350
rect 14135 6316 14169 6350
rect 14227 6316 14261 6350
rect 14319 6316 14353 6350
rect 14411 6316 14445 6350
rect 14503 6316 14537 6350
rect 14595 6316 14629 6350
rect 14687 6316 14721 6350
rect 14779 6316 14813 6350
rect 14871 6316 14905 6350
rect 14964 6316 14998 6350
rect 15055 6316 15089 6350
rect 15147 6316 15181 6350
rect 15239 6316 15273 6350
rect 15332 6316 15366 6350
rect 15423 6316 15457 6350
rect 15515 6316 15549 6350
rect 15607 6316 15641 6350
rect 15699 6316 15733 6350
rect 15791 6316 15825 6350
rect 15883 6316 15917 6350
rect 15975 6316 16009 6350
rect 16067 6316 16101 6350
rect 16159 6316 16193 6350
rect 16251 6316 16285 6350
rect 16343 6316 16377 6350
rect 16435 6316 16469 6350
rect 16526 6316 16560 6350
rect 16618 6316 16652 6350
rect 16711 6316 16745 6350
rect 16803 6316 16837 6350
rect 16895 6316 16929 6350
rect 16986 6316 17020 6350
rect 17079 6316 17113 6350
rect 17170 6316 17204 6350
rect 17263 6316 17297 6350
rect 17355 6316 17389 6350
rect 17447 6316 17481 6350
rect 17539 6316 17573 6350
rect 17631 6316 17665 6350
rect 17723 6316 17757 6350
rect 17815 6316 17849 6350
rect 17907 6316 17941 6350
rect 17999 6316 18033 6350
rect 18091 6316 18125 6350
rect 13399 5049 13433 5083
rect 13491 5049 13525 5083
rect 13583 5049 13617 5083
rect 13675 5049 13709 5083
rect 13767 5049 13801 5083
rect 13859 5049 13893 5083
rect 13951 5049 13985 5083
rect 14043 5049 14077 5083
rect 14135 5049 14169 5083
rect 14227 5049 14261 5083
rect 14319 5049 14353 5083
rect 14411 5049 14445 5083
rect 14503 5049 14537 5083
rect 14595 5049 14629 5083
rect 14687 5049 14721 5083
rect 14779 5049 14813 5083
rect 14871 5049 14905 5083
rect 14963 5049 14997 5083
rect 15055 5049 15089 5083
rect 15147 5049 15181 5083
rect 15239 5049 15273 5083
rect 15331 5049 15365 5083
rect 15423 5049 15457 5083
rect 15515 5049 15549 5083
rect 15607 5049 15641 5083
rect 15699 5049 15733 5083
rect 15791 5049 15825 5083
rect 15883 5049 15917 5083
rect 15975 5049 16009 5083
rect 16067 5049 16101 5083
rect 16159 5049 16193 5083
rect 16251 5049 16285 5083
rect 16343 5049 16377 5083
rect 16435 5049 16469 5083
rect 16527 5049 16561 5083
rect 16619 5049 16653 5083
rect 16711 5049 16745 5083
rect 16803 5049 16837 5083
rect 16895 5049 16929 5083
rect 16987 5049 17021 5083
rect 17079 5049 17113 5083
rect 17171 5049 17205 5083
rect 17263 5049 17297 5083
rect 17355 5049 17389 5083
rect 17447 5049 17481 5083
rect 17539 5049 17573 5083
rect 17631 5049 17665 5083
rect 17723 5049 17757 5083
rect 17815 5049 17849 5083
rect 17907 5049 17941 5083
rect 17999 5049 18033 5083
rect 18091 5049 18125 5083
<< nsubdiffcont >>
rect 18501 9618 18535 9652
rect 18684 9618 18718 9652
rect 13400 6955 13434 6989
rect 13491 6955 13525 6989
rect 13584 6955 13618 6989
rect 13675 6955 13709 6989
rect 13766 6955 13800 6989
rect 13860 6955 13894 6989
rect 13951 6955 13985 6989
rect 14044 6955 14078 6989
rect 14135 6955 14169 6989
rect 14227 6955 14261 6989
rect 14318 6955 14352 6989
rect 14411 6955 14445 6989
rect 14504 6955 14538 6989
rect 14595 6955 14629 6989
rect 14687 6955 14721 6989
rect 14779 6955 14813 6989
rect 14871 6955 14905 6989
rect 14963 6955 14997 6989
rect 15055 6955 15089 6989
rect 15147 6955 15181 6989
rect 15240 6955 15274 6989
rect 15330 6955 15364 6989
rect 15423 6955 15457 6989
rect 15516 6955 15550 6989
rect 15608 6955 15642 6989
rect 15699 6955 15733 6989
rect 15792 6955 15826 6989
rect 15884 6955 15918 6989
rect 15976 6955 16010 6989
rect 16068 6955 16102 6989
rect 16160 6955 16194 6989
rect 16252 6955 16286 6989
rect 16343 6955 16377 6989
rect 16434 6955 16468 6989
rect 16527 6955 16561 6989
rect 16620 6955 16654 6989
rect 16712 6955 16746 6989
rect 16803 6955 16837 6989
rect 16897 6955 16931 6989
rect 16987 6955 17021 6989
rect 17078 6955 17112 6989
rect 17171 6955 17205 6989
rect 17264 6955 17298 6989
rect 17356 6955 17390 6989
rect 17447 6955 17481 6989
rect 17539 6955 17573 6989
rect 17631 6955 17665 6989
rect 17722 6955 17756 6989
rect 17814 6955 17848 6989
rect 17907 6955 17941 6989
rect 17999 6955 18033 6989
rect 18091 6955 18125 6989
rect 13402 5674 13436 5708
rect 13492 5674 13526 5708
rect 13585 5674 13619 5708
rect 13675 5674 13709 5708
rect 13766 5674 13800 5708
rect 13860 5674 13894 5708
rect 13951 5674 13985 5708
rect 14043 5674 14077 5708
rect 14135 5674 14169 5708
rect 14228 5674 14262 5708
rect 14319 5674 14353 5708
rect 14411 5674 14445 5708
rect 14503 5674 14537 5708
rect 14595 5674 14629 5708
rect 14688 5674 14722 5708
rect 14779 5674 14813 5708
rect 14870 5674 14904 5708
rect 14963 5674 14997 5708
rect 15056 5674 15090 5708
rect 15147 5674 15181 5708
rect 15239 5674 15273 5708
rect 15331 5674 15365 5708
rect 15423 5674 15457 5708
rect 15516 5674 15550 5708
rect 15606 5674 15640 5708
rect 15699 5674 15733 5708
rect 15791 5674 15825 5708
rect 15884 5674 15918 5708
rect 15978 5674 16012 5708
rect 16067 5674 16101 5708
rect 16159 5674 16193 5708
rect 16251 5674 16285 5708
rect 16343 5674 16377 5708
rect 16435 5674 16469 5708
rect 16527 5674 16561 5708
rect 16619 5674 16653 5708
rect 16711 5674 16745 5708
rect 16803 5674 16837 5708
rect 16895 5674 16929 5708
rect 16987 5674 17021 5708
rect 17079 5674 17113 5708
rect 17171 5674 17205 5708
rect 17263 5674 17297 5708
rect 17355 5674 17389 5708
rect 17447 5674 17481 5708
rect 17539 5674 17573 5708
rect 17631 5674 17665 5708
rect 17723 5674 17757 5708
rect 17815 5674 17849 5708
rect 17907 5674 17941 5708
rect 18000 5674 18034 5708
rect 18091 5674 18125 5708
<< locali >>
rect 18472 9652 18841 9654
rect 18472 9618 18501 9652
rect 18535 9618 18684 9652
rect 18718 9618 18841 9652
rect 18473 9040 18593 9041
rect 18473 9006 18501 9040
rect 18535 9007 18593 9040
rect 18627 9007 18685 9041
rect 18719 9007 18778 9041
rect 18812 9007 18842 9041
rect 18535 9006 18842 9007
rect 18473 9005 18842 9006
rect 13370 7581 13399 7615
rect 13433 7581 13491 7615
rect 13525 7581 13583 7615
rect 13617 7581 13675 7615
rect 13709 7581 13767 7615
rect 13801 7581 13859 7615
rect 13893 7581 13951 7615
rect 13985 7581 14043 7615
rect 14077 7581 14135 7615
rect 14169 7581 14226 7615
rect 14260 7581 14319 7615
rect 14353 7581 14411 7615
rect 14445 7581 14503 7615
rect 14537 7581 14595 7615
rect 14629 7581 14687 7615
rect 14721 7581 14779 7615
rect 14813 7581 14871 7615
rect 14905 7581 14963 7615
rect 14997 7581 15055 7615
rect 15089 7581 15147 7615
rect 15181 7581 15239 7615
rect 15273 7581 15331 7615
rect 15365 7581 15423 7615
rect 15457 7581 15515 7615
rect 15549 7581 15607 7615
rect 15641 7581 15699 7615
rect 15733 7581 15791 7615
rect 15825 7581 15883 7615
rect 15917 7581 15975 7615
rect 16009 7581 16067 7615
rect 16101 7581 16159 7615
rect 16193 7581 16251 7615
rect 16285 7581 16343 7615
rect 16377 7581 16435 7615
rect 16469 7581 16527 7615
rect 16561 7581 16619 7615
rect 16653 7581 16711 7615
rect 16745 7581 16803 7615
rect 16837 7581 16895 7615
rect 16929 7581 16987 7615
rect 17021 7581 17079 7615
rect 17113 7581 17171 7615
rect 17205 7581 17263 7615
rect 17297 7581 17355 7615
rect 17389 7581 17447 7615
rect 17481 7581 17539 7615
rect 17573 7581 17631 7615
rect 17665 7581 17723 7615
rect 17757 7581 17815 7615
rect 17849 7581 17907 7615
rect 17941 7581 17999 7615
rect 18033 7581 18091 7615
rect 18125 7581 18154 7615
rect 13370 6989 18154 7008
rect 13370 6955 13400 6989
rect 13434 6955 13491 6989
rect 13525 6955 13584 6989
rect 13618 6955 13675 6989
rect 13709 6955 13766 6989
rect 13800 6955 13860 6989
rect 13894 6955 13951 6989
rect 13985 6955 14044 6989
rect 14078 6955 14135 6989
rect 14169 6955 14227 6989
rect 14261 6955 14318 6989
rect 14352 6955 14411 6989
rect 14445 6955 14504 6989
rect 14538 6955 14595 6989
rect 14629 6955 14687 6989
rect 14721 6955 14779 6989
rect 14813 6955 14871 6989
rect 14905 6955 14963 6989
rect 14997 6955 15055 6989
rect 15089 6955 15147 6989
rect 15181 6955 15240 6989
rect 15274 6955 15330 6989
rect 15364 6955 15423 6989
rect 15457 6955 15516 6989
rect 15550 6955 15608 6989
rect 15642 6955 15699 6989
rect 15733 6955 15792 6989
rect 15826 6955 15884 6989
rect 15918 6955 15976 6989
rect 16010 6955 16068 6989
rect 16102 6955 16160 6989
rect 16194 6955 16252 6989
rect 16286 6955 16343 6989
rect 16377 6955 16434 6989
rect 16468 6955 16527 6989
rect 16561 6955 16620 6989
rect 16654 6955 16712 6989
rect 16746 6955 16803 6989
rect 16837 6955 16897 6989
rect 16931 6955 16987 6989
rect 17021 6955 17078 6989
rect 17112 6955 17171 6989
rect 17205 6955 17264 6989
rect 17298 6955 17356 6989
rect 17390 6955 17447 6989
rect 17481 6955 17539 6989
rect 17573 6955 17631 6989
rect 17665 6955 17722 6989
rect 17756 6955 17814 6989
rect 17848 6955 17907 6989
rect 17941 6955 17999 6989
rect 18033 6955 18091 6989
rect 18125 6955 18154 6989
rect 13370 6933 18154 6955
rect 13370 6350 18154 6367
rect 13370 6316 13399 6350
rect 13433 6316 13491 6350
rect 13525 6316 13583 6350
rect 13617 6316 13675 6350
rect 13709 6316 13767 6350
rect 13801 6316 13859 6350
rect 13893 6316 13951 6350
rect 13985 6316 14043 6350
rect 14077 6316 14135 6350
rect 14169 6316 14227 6350
rect 14261 6316 14319 6350
rect 14353 6316 14411 6350
rect 14445 6316 14503 6350
rect 14537 6316 14595 6350
rect 14629 6316 14687 6350
rect 14721 6316 14779 6350
rect 14813 6316 14871 6350
rect 14905 6316 14964 6350
rect 14998 6316 15055 6350
rect 15089 6316 15147 6350
rect 15181 6316 15239 6350
rect 15273 6316 15332 6350
rect 15366 6316 15423 6350
rect 15457 6316 15515 6350
rect 15549 6316 15607 6350
rect 15641 6316 15699 6350
rect 15733 6316 15791 6350
rect 15825 6316 15883 6350
rect 15917 6316 15975 6350
rect 16009 6316 16067 6350
rect 16101 6316 16159 6350
rect 16193 6316 16251 6350
rect 16285 6316 16343 6350
rect 16377 6316 16435 6350
rect 16469 6316 16526 6350
rect 16560 6316 16618 6350
rect 16652 6316 16711 6350
rect 16745 6316 16803 6350
rect 16837 6316 16895 6350
rect 16929 6316 16986 6350
rect 17020 6316 17079 6350
rect 17113 6316 17170 6350
rect 17204 6316 17263 6350
rect 17297 6316 17355 6350
rect 17389 6316 17447 6350
rect 17481 6316 17539 6350
rect 17573 6316 17631 6350
rect 17665 6316 17723 6350
rect 17757 6316 17815 6350
rect 17849 6316 17907 6350
rect 17941 6316 17999 6350
rect 18033 6316 18091 6350
rect 18125 6316 18154 6350
rect 13370 6292 18154 6316
rect 13370 5708 18154 5726
rect 13370 5674 13402 5708
rect 13436 5674 13492 5708
rect 13526 5674 13585 5708
rect 13619 5674 13675 5708
rect 13709 5674 13766 5708
rect 13800 5674 13860 5708
rect 13894 5674 13951 5708
rect 13985 5674 14043 5708
rect 14077 5674 14135 5708
rect 14169 5674 14228 5708
rect 14262 5674 14319 5708
rect 14353 5674 14411 5708
rect 14445 5674 14503 5708
rect 14537 5674 14595 5708
rect 14629 5674 14688 5708
rect 14722 5674 14779 5708
rect 14813 5674 14870 5708
rect 14904 5674 14963 5708
rect 14997 5674 15056 5708
rect 15090 5674 15147 5708
rect 15181 5674 15239 5708
rect 15273 5674 15331 5708
rect 15365 5674 15423 5708
rect 15457 5674 15516 5708
rect 15550 5674 15606 5708
rect 15640 5674 15699 5708
rect 15733 5674 15791 5708
rect 15825 5674 15884 5708
rect 15918 5674 15978 5708
rect 16012 5674 16067 5708
rect 16101 5674 16159 5708
rect 16193 5674 16251 5708
rect 16285 5674 16343 5708
rect 16377 5674 16435 5708
rect 16469 5674 16527 5708
rect 16561 5674 16619 5708
rect 16653 5674 16711 5708
rect 16745 5674 16803 5708
rect 16837 5674 16895 5708
rect 16929 5674 16987 5708
rect 17021 5674 17079 5708
rect 17113 5674 17171 5708
rect 17205 5674 17263 5708
rect 17297 5674 17355 5708
rect 17389 5674 17447 5708
rect 17481 5674 17539 5708
rect 17573 5674 17631 5708
rect 17665 5674 17723 5708
rect 17757 5674 17815 5708
rect 17849 5674 17907 5708
rect 17941 5674 18000 5708
rect 18034 5674 18091 5708
rect 18125 5674 18154 5708
rect 13370 5651 18154 5674
rect 13370 5049 13399 5083
rect 13433 5049 13491 5083
rect 13525 5049 13583 5083
rect 13617 5049 13675 5083
rect 13709 5049 13767 5083
rect 13801 5049 13859 5083
rect 13893 5049 13951 5083
rect 13985 5049 14043 5083
rect 14077 5049 14135 5083
rect 14169 5049 14227 5083
rect 14261 5049 14319 5083
rect 14353 5049 14411 5083
rect 14445 5049 14503 5083
rect 14537 5049 14595 5083
rect 14629 5049 14687 5083
rect 14721 5049 14779 5083
rect 14813 5049 14871 5083
rect 14905 5049 14963 5083
rect 14997 5049 15055 5083
rect 15089 5049 15147 5083
rect 15181 5049 15239 5083
rect 15273 5049 15331 5083
rect 15365 5049 15423 5083
rect 15457 5049 15515 5083
rect 15549 5049 15607 5083
rect 15641 5049 15699 5083
rect 15733 5049 15791 5083
rect 15825 5049 15883 5083
rect 15917 5049 15975 5083
rect 16009 5049 16067 5083
rect 16101 5049 16159 5083
rect 16193 5049 16251 5083
rect 16285 5049 16343 5083
rect 16377 5049 16435 5083
rect 16469 5049 16527 5083
rect 16561 5049 16619 5083
rect 16653 5049 16711 5083
rect 16745 5049 16803 5083
rect 16837 5049 16895 5083
rect 16929 5049 16987 5083
rect 17021 5049 17079 5083
rect 17113 5049 17171 5083
rect 17205 5049 17263 5083
rect 17297 5049 17355 5083
rect 17389 5049 17447 5083
rect 17481 5049 17539 5083
rect 17573 5049 17631 5083
rect 17665 5049 17723 5083
rect 17757 5049 17815 5083
rect 17849 5049 17907 5083
rect 17941 5049 17999 5083
rect 18033 5049 18091 5083
rect 18125 5049 18154 5083
<< viali >>
rect 18495 9275 18529 9309
rect 18702 9275 18736 9309
rect 18091 7426 18125 7460
rect 13416 7321 13450 7355
rect 15255 7306 15289 7340
rect 13736 7247 13770 7281
rect 15805 7276 15839 7310
rect 16138 7309 16172 7343
rect 17654 7310 17688 7344
rect 15703 7109 15737 7143
rect 15702 6797 15736 6831
rect 13411 6671 13445 6705
rect 13741 6601 13775 6635
rect 15256 6599 15290 6633
rect 15806 6628 15840 6662
rect 16139 6600 16173 6634
rect 17649 6600 17683 6634
rect 18092 6468 18126 6502
rect 18086 6145 18120 6179
rect 13419 6055 13453 6089
rect 15265 6029 15299 6063
rect 15803 6011 15837 6045
rect 16140 6028 16174 6062
rect 17649 6031 17683 6065
rect 13746 5971 13780 6005
rect 15699 5834 15733 5868
rect 15699 5519 15733 5553
rect 13743 5379 13777 5413
rect 13415 5295 13449 5329
rect 15257 5319 15291 5353
rect 15804 5325 15838 5359
rect 16141 5320 16175 5354
rect 17649 5320 17683 5354
rect 18087 5186 18121 5220
<< metal1 >>
rect 18564 9693 18654 9709
rect 11730 9654 11784 9688
rect 18564 9682 18583 9693
rect 18545 9641 18583 9682
rect 18635 9641 18654 9693
rect 18764 9693 18854 9709
rect 18764 9682 18783 9693
rect 18545 9623 18654 9641
rect 18745 9641 18783 9682
rect 18835 9641 18854 9693
rect 18745 9623 18854 9641
rect 11767 9271 11864 9318
rect 18424 9309 18542 9315
rect 18424 9275 18495 9309
rect 18529 9275 18542 9309
rect 18424 9269 18542 9275
rect 18690 9309 18748 9315
rect 18690 9275 18702 9309
rect 18736 9306 18748 9309
rect 18736 9278 18897 9306
rect 18736 9275 18748 9278
rect 18690 9269 18748 9275
rect 12030 9069 12142 9117
rect 18358 9051 18841 9067
rect 18358 8999 18394 9051
rect 18446 8999 18841 9051
rect 18358 8983 18841 8999
rect 17602 7984 17899 7991
rect 13338 7918 14277 7946
rect 16645 7890 16703 7963
rect 13338 7862 16703 7890
rect 17501 7834 17560 7954
rect 13338 7806 17560 7834
rect 17602 7778 17934 7984
rect 13285 7750 17934 7778
rect 13285 7612 13339 7750
rect 13409 7655 13415 7707
rect 13467 7695 13473 7707
rect 15803 7695 15809 7707
rect 13467 7667 15809 7695
rect 13467 7655 13473 7667
rect 15803 7655 15809 7667
rect 15861 7695 15867 7707
rect 18869 7695 18897 9278
rect 15861 7667 18897 7695
rect 15861 7655 15867 7667
rect 13285 7516 13400 7612
rect 13491 7589 13525 7615
rect 13491 7581 13507 7589
rect 13500 7537 13507 7581
rect 13559 7537 13566 7589
rect 13583 7581 13617 7615
rect 13675 7588 13709 7615
rect 13674 7536 13681 7588
rect 13733 7536 13740 7588
rect 13767 7581 13801 7615
rect 13859 7581 13893 7615
rect 13951 7590 13985 7615
rect 13899 7538 13906 7590
rect 13958 7581 13985 7590
rect 14043 7581 14077 7615
rect 14135 7592 14169 7615
rect 13958 7538 13965 7581
rect 14100 7540 14107 7592
rect 14159 7581 14169 7592
rect 14226 7581 14260 7615
rect 14319 7590 14353 7615
rect 14319 7581 14330 7590
rect 14159 7540 14166 7581
rect 14323 7538 14330 7581
rect 14382 7538 14389 7590
rect 14411 7581 14445 7615
rect 14503 7595 14537 7615
rect 14595 7595 14629 7615
rect 14503 7581 14539 7595
rect 14532 7543 14539 7581
rect 14591 7581 14629 7595
rect 14687 7581 14721 7615
rect 14779 7588 14813 7615
rect 14591 7543 14598 7581
rect 14760 7536 14767 7588
rect 14819 7536 14826 7588
rect 14871 7581 14905 7615
rect 14963 7592 14997 7615
rect 14950 7540 14957 7592
rect 15009 7540 15016 7592
rect 15055 7581 15089 7615
rect 15147 7595 15181 7615
rect 15147 7581 15162 7595
rect 15155 7543 15162 7581
rect 15214 7543 15221 7595
rect 15239 7581 15273 7615
rect 15331 7595 15365 7615
rect 15331 7581 15361 7595
rect 15354 7543 15361 7581
rect 15413 7543 15420 7595
rect 15423 7581 15457 7615
rect 15515 7581 15549 7615
rect 15607 7590 15641 7615
rect 15570 7538 15577 7590
rect 15629 7581 15641 7590
rect 15699 7581 15733 7615
rect 15791 7581 15825 7615
rect 15883 7581 15917 7615
rect 15975 7595 16009 7615
rect 15629 7538 15636 7581
rect 15958 7543 15965 7595
rect 16017 7543 16024 7595
rect 16067 7581 16101 7615
rect 16159 7590 16193 7615
rect 16251 7590 16285 7615
rect 16159 7581 16200 7590
rect 16193 7538 16200 7581
rect 16252 7581 16285 7590
rect 16343 7581 16377 7615
rect 16435 7592 16469 7615
rect 16252 7538 16259 7581
rect 16435 7540 16442 7592
rect 16494 7540 16501 7592
rect 16527 7581 16561 7615
rect 16619 7581 16653 7615
rect 16711 7593 16745 7615
rect 16667 7541 16674 7593
rect 16726 7581 16745 7593
rect 16803 7581 16837 7615
rect 16895 7596 16929 7615
rect 16895 7581 16903 7596
rect 16726 7541 16733 7581
rect 16896 7544 16903 7581
rect 16955 7544 16962 7596
rect 16987 7581 17021 7615
rect 17079 7581 17113 7615
rect 17171 7588 17205 7615
rect 17145 7536 17152 7588
rect 17204 7536 17211 7588
rect 17263 7581 17297 7615
rect 17355 7592 17389 7615
rect 17355 7581 17370 7592
rect 17363 7540 17370 7581
rect 17422 7540 17429 7592
rect 17447 7581 17481 7615
rect 17539 7581 17573 7615
rect 17631 7588 17665 7615
rect 17592 7536 17599 7588
rect 17651 7581 17665 7588
rect 17723 7581 17757 7615
rect 17815 7590 17849 7615
rect 17651 7536 17658 7581
rect 17813 7538 17820 7590
rect 17872 7538 17879 7590
rect 17907 7581 17941 7615
rect 17999 7595 18033 7615
rect 18091 7595 18125 7615
rect 17999 7581 18036 7595
rect 18029 7543 18036 7581
rect 18088 7581 18125 7595
rect 18088 7543 18095 7581
rect 13289 7476 13334 7486
rect 13289 7448 15907 7476
rect 18207 7466 18252 7476
rect 18078 7460 18252 7466
rect 13289 7438 13334 7448
rect 13406 7364 13458 7370
rect 14858 7350 14865 7402
rect 14917 7350 14924 7402
rect 13406 7306 13458 7312
rect 15243 7299 15250 7351
rect 15302 7299 15309 7351
rect 15878 7342 15906 7448
rect 18078 7426 18091 7460
rect 18125 7437 18252 7460
rect 18125 7426 18137 7437
rect 18207 7428 18252 7437
rect 18078 7420 18137 7426
rect 16120 7343 16187 7352
rect 17253 7349 17260 7401
rect 17312 7349 17319 7401
rect 16120 7342 16138 7343
rect 15798 7322 15850 7328
rect 15878 7314 16138 7342
rect 13721 7281 13782 7287
rect 13297 7269 13342 7280
rect 13721 7269 13736 7281
rect 13297 7247 13736 7269
rect 13770 7247 13782 7281
rect 16120 7309 16138 7314
rect 16172 7309 16187 7343
rect 16120 7301 16187 7309
rect 17638 7300 17645 7352
rect 17697 7300 17704 7352
rect 15798 7264 15850 7270
rect 13297 7241 13782 7247
rect 13297 7232 13342 7241
rect 15691 7143 15749 7150
rect 15691 7109 15703 7143
rect 15737 7136 15749 7143
rect 18207 7136 18252 7146
rect 15737 7109 18252 7136
rect 15691 7108 18252 7109
rect 15691 7102 15749 7108
rect 18207 7098 18252 7108
rect 13502 6988 13509 7006
rect 13491 6954 13509 6988
rect 13561 6954 13568 7006
rect 13584 6955 13618 6989
rect 13677 6952 13684 7004
rect 13736 6952 13743 7004
rect 13874 6954 13881 7006
rect 13933 6954 13940 7006
rect 14093 6957 14100 7009
rect 14152 6957 14159 7009
rect 14325 6953 14332 7005
rect 14384 6953 14391 7005
rect 14549 6960 14556 7012
rect 14608 6960 14615 7012
rect 14761 6948 14768 7000
rect 14820 6948 14827 7000
rect 14983 6944 14990 6996
rect 15042 6944 15049 6996
rect 15206 6941 15213 6993
rect 15265 6941 15272 6993
rect 15416 6941 15423 6993
rect 15475 6941 15482 6993
rect 15629 6941 15636 6993
rect 15688 6941 15695 6993
rect 15792 6954 15826 6988
rect 15946 6934 15953 6986
rect 16005 6934 16012 6986
rect 16148 6937 16155 6989
rect 16207 6937 16214 6989
rect 16349 6938 16356 6990
rect 16408 6938 16415 6990
rect 16528 6939 16535 6991
rect 16587 6939 16594 6991
rect 16720 6943 16727 6995
rect 16779 6943 16786 6995
rect 16905 6940 16912 6992
rect 16964 6940 16971 6992
rect 17137 6939 17144 6991
rect 17196 6939 17203 6991
rect 17342 6941 17349 6993
rect 17401 6941 17408 6993
rect 17548 6943 17555 6995
rect 17607 6943 17614 6995
rect 17649 6940 17655 6992
rect 17707 6940 17713 6992
rect 17756 6950 17763 7002
rect 17815 6950 17822 7002
rect 17978 6951 17985 7003
rect 18037 6951 18044 7003
rect 18207 6837 18252 6847
rect 15689 6831 18252 6837
rect 15689 6797 15702 6831
rect 15736 6809 18252 6831
rect 15736 6797 15750 6809
rect 18207 6799 18252 6809
rect 15689 6790 15750 6797
rect 13401 6715 13453 6721
rect 13401 6657 13453 6663
rect 15797 6673 15849 6679
rect 13307 6629 13352 6639
rect 13723 6635 13790 6644
rect 13723 6629 13741 6635
rect 13307 6601 13741 6629
rect 13775 6601 13790 6635
rect 13307 6591 13352 6601
rect 13723 6593 13790 6601
rect 15242 6588 15248 6640
rect 15300 6588 15306 6640
rect 16121 6634 16188 6643
rect 16121 6629 16139 6634
rect 15797 6615 15849 6621
rect 15885 6601 16139 6629
rect 14484 6524 14490 6576
rect 14542 6524 14548 6576
rect 14484 6523 14548 6524
rect 13310 6495 13355 6505
rect 15885 6495 15913 6601
rect 16121 6600 16139 6601
rect 16173 6600 16188 6634
rect 16121 6592 16188 6600
rect 17635 6589 17641 6641
rect 17693 6589 17699 6641
rect 16879 6524 16885 6576
rect 16937 6524 16943 6576
rect 18080 6502 18137 6514
rect 13310 6467 15914 6495
rect 18080 6468 18092 6502
rect 18126 6499 18137 6502
rect 18212 6499 18257 6505
rect 18126 6468 18257 6499
rect 13310 6457 13355 6467
rect 18080 6465 18257 6468
rect 18080 6462 18137 6465
rect 18212 6457 18257 6465
rect 13399 6315 13433 6349
rect 13491 6316 13525 6350
rect 13529 6305 13536 6357
rect 13588 6350 13595 6357
rect 13588 6316 13617 6350
rect 13675 6316 13709 6350
rect 13588 6305 13595 6316
rect 13745 6310 13752 6362
rect 13804 6310 13811 6362
rect 13859 6316 13893 6350
rect 13951 6311 13958 6363
rect 14010 6311 14017 6363
rect 14153 6350 14160 6355
rect 14043 6316 14077 6350
rect 14135 6316 14160 6350
rect 14153 6303 14160 6316
rect 14212 6303 14219 6355
rect 14349 6350 14356 6357
rect 14227 6316 14261 6350
rect 14319 6316 14356 6350
rect 14349 6305 14356 6316
rect 14408 6350 14415 6357
rect 14408 6316 14445 6350
rect 14503 6316 14537 6350
rect 14408 6305 14415 6316
rect 14574 6307 14581 6359
rect 14633 6307 14640 6359
rect 14789 6350 14796 6355
rect 14687 6316 14721 6350
rect 14779 6316 14796 6350
rect 14789 6303 14796 6316
rect 14848 6303 14855 6355
rect 14871 6316 14905 6350
rect 14964 6316 14998 6350
rect 15024 6303 15031 6355
rect 15083 6303 15090 6355
rect 15147 6316 15181 6350
rect 15232 6306 15239 6358
rect 15291 6306 15298 6358
rect 15332 6316 15366 6350
rect 15423 6316 15457 6350
rect 15474 6306 15481 6358
rect 15533 6350 15540 6358
rect 15533 6316 15549 6350
rect 15607 6316 15641 6350
rect 15533 6306 15540 6316
rect 15672 6307 15679 6359
rect 15731 6307 15738 6359
rect 15979 6350 15986 6359
rect 15791 6316 15825 6350
rect 15883 6316 15917 6350
rect 15975 6316 15986 6350
rect 15979 6307 15986 6316
rect 16038 6307 16045 6359
rect 16067 6316 16101 6350
rect 16159 6316 16193 6350
rect 16204 6308 16211 6360
rect 16263 6350 16270 6360
rect 16263 6316 16285 6350
rect 16343 6316 16377 6350
rect 16263 6308 16270 6316
rect 16433 6307 16440 6359
rect 16492 6307 16499 6359
rect 16649 6350 16656 6363
rect 16526 6316 16560 6350
rect 16618 6316 16656 6350
rect 16649 6311 16656 6316
rect 16708 6350 16715 6363
rect 16708 6316 16745 6350
rect 16803 6316 16837 6350
rect 16708 6311 16715 6316
rect 16872 6314 16879 6366
rect 16931 6314 16938 6366
rect 17096 6350 17103 6362
rect 16986 6316 17020 6350
rect 17079 6316 17103 6350
rect 17096 6310 17103 6316
rect 17155 6310 17162 6362
rect 17170 6316 17204 6350
rect 17263 6316 17297 6350
rect 17323 6299 17330 6351
rect 17382 6299 17389 6351
rect 17747 6350 17754 6354
rect 17447 6316 17481 6350
rect 17536 6298 17543 6350
rect 17595 6298 17602 6350
rect 17631 6316 17665 6350
rect 17723 6316 17754 6350
rect 17747 6302 17754 6316
rect 17806 6302 17813 6354
rect 17815 6316 17849 6350
rect 17907 6316 17941 6350
rect 17974 6303 17981 6355
rect 18033 6303 18040 6355
rect 18091 6316 18125 6350
rect 13297 6196 13342 6205
rect 13297 6168 15928 6196
rect 18203 6189 18248 6195
rect 18070 6179 18248 6189
rect 13297 6157 13342 6168
rect 13409 6100 13461 6106
rect 14863 6076 14870 6128
rect 14922 6076 14929 6128
rect 13409 6042 13461 6048
rect 15246 6017 15253 6069
rect 15305 6017 15312 6069
rect 15796 6057 15848 6063
rect 13728 6005 13795 6014
rect 13298 5990 13343 6002
rect 13728 5990 13746 6005
rect 13298 5971 13746 5990
rect 13780 5971 13795 6005
rect 15899 6062 15927 6168
rect 18070 6145 18086 6179
rect 18120 6155 18248 6179
rect 18120 6145 18137 6155
rect 18203 6147 18248 6155
rect 18070 6135 18137 6145
rect 17255 6078 17262 6130
rect 17314 6078 17321 6130
rect 16122 6062 16189 6071
rect 15899 6034 16140 6062
rect 16122 6028 16140 6034
rect 16174 6028 16189 6062
rect 16122 6020 16189 6028
rect 17632 6024 17639 6076
rect 17691 6024 17698 6076
rect 15796 5999 15848 6005
rect 13298 5963 13795 5971
rect 13298 5962 13744 5963
rect 13298 5954 13343 5962
rect 15684 5868 15747 5874
rect 15684 5834 15699 5868
rect 15733 5855 15747 5868
rect 18206 5855 18251 5864
rect 15733 5834 18251 5855
rect 15684 5827 18251 5834
rect 18206 5816 18251 5827
rect 13555 5660 13562 5712
rect 13614 5660 13621 5712
rect 13780 5669 13787 5721
rect 13839 5669 13846 5721
rect 14057 5666 14064 5718
rect 14116 5666 14123 5718
rect 14278 5669 14285 5721
rect 14337 5669 14344 5721
rect 14523 5666 14530 5718
rect 14582 5666 14589 5718
rect 14749 5670 14756 5722
rect 14808 5670 14815 5722
rect 14961 5668 14968 5720
rect 15020 5668 15027 5720
rect 15181 5674 15188 5726
rect 15240 5674 15247 5726
rect 15419 5676 15426 5728
rect 15478 5676 15485 5728
rect 15632 5678 15639 5730
rect 15691 5678 15698 5730
rect 16019 5668 16026 5720
rect 16078 5668 16085 5720
rect 16366 5669 16373 5721
rect 16425 5669 16432 5721
rect 16602 5664 16609 5716
rect 16661 5664 16668 5716
rect 16786 5664 16793 5716
rect 16845 5664 16852 5716
rect 17025 5666 17032 5718
rect 17084 5666 17091 5718
rect 17228 5662 17235 5714
rect 17287 5662 17294 5714
rect 17413 5659 17420 5711
rect 17472 5659 17479 5711
rect 17604 5661 17611 5713
rect 17663 5661 17670 5713
rect 17795 5665 17802 5717
rect 17854 5665 17861 5717
rect 17981 5661 17988 5713
rect 18040 5661 18047 5713
rect 18209 5560 18254 5568
rect 15687 5553 18254 5560
rect 15687 5519 15699 5553
rect 15733 5532 18254 5553
rect 15733 5519 15745 5532
rect 18209 5520 18254 5532
rect 15687 5512 15745 5519
rect 13285 5412 13330 5424
rect 13725 5413 13792 5422
rect 13725 5412 13743 5413
rect 13285 5384 13743 5412
rect 13285 5376 13330 5384
rect 13725 5379 13743 5384
rect 13777 5379 13792 5413
rect 13725 5371 13792 5379
rect 15797 5370 15849 5376
rect 15242 5361 15307 5362
rect 13404 5340 13456 5346
rect 15242 5309 15248 5361
rect 15300 5309 15307 5361
rect 16123 5354 16190 5363
rect 16123 5349 16141 5354
rect 15797 5312 15849 5318
rect 15886 5321 16141 5349
rect 13404 5282 13456 5288
rect 14491 5244 14499 5296
rect 14551 5244 14557 5296
rect 13282 5215 13327 5225
rect 15886 5215 15914 5321
rect 16123 5320 16141 5321
rect 16175 5320 16190 5354
rect 16123 5312 16190 5320
rect 17634 5362 17698 5363
rect 17634 5310 17640 5362
rect 17692 5310 17698 5362
rect 16882 5244 16889 5296
rect 16942 5244 16949 5296
rect 18075 5220 18133 5227
rect 13282 5187 15915 5215
rect 13282 5177 13327 5187
rect 18075 5186 18087 5220
rect 18121 5218 18133 5220
rect 18205 5218 18250 5224
rect 18121 5186 18250 5218
rect 18075 5184 18250 5186
rect 18075 5180 18133 5184
rect 18205 5176 18250 5184
rect 13428 5083 13435 5130
rect 13399 5078 13435 5083
rect 13487 5083 13494 5130
rect 13487 5078 13525 5083
rect 13399 5049 13433 5078
rect 13491 5049 13525 5078
rect 13583 5049 13617 5083
rect 13633 5074 13640 5126
rect 13692 5083 13699 5126
rect 13692 5074 13709 5083
rect 13675 5049 13709 5074
rect 13767 5049 13801 5083
rect 13819 5079 13826 5131
rect 13878 5083 13885 5131
rect 13878 5079 13893 5083
rect 13859 5049 13893 5079
rect 13951 5049 13985 5083
rect 14013 5072 14020 5124
rect 14072 5072 14079 5124
rect 14232 5083 14239 5129
rect 14043 5049 14077 5072
rect 14135 5049 14169 5083
rect 14227 5077 14239 5083
rect 14291 5077 14298 5129
rect 14442 5083 14449 5129
rect 14227 5049 14261 5077
rect 14319 5049 14353 5083
rect 14411 5077 14449 5083
rect 14501 5083 14508 5129
rect 14501 5077 14537 5083
rect 14411 5049 14445 5077
rect 14503 5049 14537 5077
rect 14595 5049 14629 5083
rect 14671 5074 14678 5126
rect 14730 5074 14737 5126
rect 14687 5049 14721 5074
rect 14779 5049 14813 5083
rect 14871 5049 14905 5083
rect 14917 5074 14924 5126
rect 14976 5083 14983 5126
rect 14976 5074 14997 5083
rect 14963 5049 14997 5074
rect 15055 5049 15089 5083
rect 15147 5049 15181 5083
rect 15191 5074 15198 5126
rect 15250 5083 15257 5126
rect 15250 5074 15273 5083
rect 15239 5049 15273 5074
rect 15331 5049 15365 5083
rect 15423 5049 15457 5083
rect 15466 5074 15473 5126
rect 15525 5083 15532 5126
rect 15702 5083 15709 5126
rect 15525 5074 15549 5083
rect 15515 5049 15549 5074
rect 15607 5049 15641 5083
rect 15699 5074 15709 5083
rect 15761 5074 15768 5126
rect 15699 5049 15733 5074
rect 15791 5049 15825 5083
rect 15883 5049 15917 5083
rect 15925 5077 15932 5129
rect 15984 5083 15991 5129
rect 15984 5077 16009 5083
rect 15975 5049 16009 5077
rect 16067 5049 16101 5083
rect 16143 5080 16150 5132
rect 16202 5080 16209 5132
rect 16159 5049 16193 5080
rect 16251 5049 16285 5083
rect 16321 5071 16328 5123
rect 16380 5071 16387 5123
rect 16560 5083 16567 5125
rect 16343 5049 16377 5071
rect 16435 5049 16469 5083
rect 16527 5073 16567 5083
rect 16619 5083 16626 5125
rect 16527 5049 16561 5073
rect 16619 5049 16653 5083
rect 16711 5049 16745 5083
rect 16757 5073 16764 5125
rect 16816 5083 16823 5125
rect 16816 5073 16837 5083
rect 16803 5049 16837 5073
rect 16895 5049 16929 5083
rect 16955 5073 16962 5125
rect 17014 5073 17021 5125
rect 16987 5049 17021 5073
rect 17079 5049 17113 5083
rect 17168 5074 17175 5126
rect 17227 5074 17234 5126
rect 17171 5049 17205 5074
rect 17263 5049 17297 5083
rect 17355 5049 17389 5083
rect 17391 5073 17398 5125
rect 17450 5083 17457 5125
rect 17450 5073 17481 5083
rect 17447 5049 17481 5073
rect 17539 5049 17573 5083
rect 17588 5078 17595 5130
rect 17647 5083 17654 5130
rect 17647 5078 17665 5083
rect 17631 5049 17665 5078
rect 17723 5049 17757 5083
rect 17804 5076 17811 5128
rect 17863 5076 17870 5128
rect 18013 5083 18020 5128
rect 17815 5049 17849 5076
rect 17907 5049 17941 5083
rect 17999 5076 18020 5083
rect 18072 5076 18079 5128
rect 17999 5049 18033 5076
rect 18091 5049 18125 5083
<< via1 >>
rect 18583 9641 18635 9693
rect 18783 9641 18835 9693
rect 18394 8999 18446 9051
rect 13415 7655 13467 7707
rect 15809 7655 15861 7707
rect 13507 7537 13559 7589
rect 13681 7536 13733 7588
rect 13906 7538 13958 7590
rect 14107 7540 14159 7592
rect 14330 7538 14382 7590
rect 14539 7543 14591 7595
rect 14767 7536 14819 7588
rect 14957 7540 15009 7592
rect 15162 7543 15214 7595
rect 15361 7543 15413 7595
rect 15577 7538 15629 7590
rect 15965 7543 16017 7595
rect 16200 7538 16252 7590
rect 16442 7540 16494 7592
rect 16674 7541 16726 7593
rect 16903 7544 16955 7596
rect 17152 7536 17204 7588
rect 17370 7540 17422 7592
rect 17599 7536 17651 7588
rect 17820 7538 17872 7590
rect 18036 7543 18088 7595
rect 13406 7355 13458 7364
rect 13406 7321 13416 7355
rect 13416 7321 13450 7355
rect 13450 7321 13458 7355
rect 14865 7350 14917 7402
rect 13406 7312 13458 7321
rect 15250 7340 15302 7351
rect 15250 7306 15255 7340
rect 15255 7306 15289 7340
rect 15289 7306 15302 7340
rect 15250 7299 15302 7306
rect 17260 7349 17312 7401
rect 15798 7310 15850 7322
rect 15798 7276 15805 7310
rect 15805 7276 15839 7310
rect 15839 7276 15850 7310
rect 17645 7344 17697 7352
rect 17645 7310 17654 7344
rect 17654 7310 17688 7344
rect 17688 7310 17697 7344
rect 17645 7300 17697 7310
rect 15798 7270 15850 7276
rect 13509 6954 13561 7006
rect 13684 6952 13736 7004
rect 13881 6954 13933 7006
rect 14100 6957 14152 7009
rect 14332 6953 14384 7005
rect 14556 6960 14608 7012
rect 14768 6948 14820 7000
rect 14990 6944 15042 6996
rect 15213 6941 15265 6993
rect 15423 6941 15475 6993
rect 15636 6941 15688 6993
rect 15953 6934 16005 6986
rect 16155 6937 16207 6989
rect 16356 6938 16408 6990
rect 16535 6939 16587 6991
rect 16727 6943 16779 6995
rect 16912 6940 16964 6992
rect 17144 6939 17196 6991
rect 17349 6941 17401 6993
rect 17555 6943 17607 6995
rect 17655 6940 17707 6992
rect 17763 6950 17815 7002
rect 17985 6951 18037 7003
rect 13401 6705 13453 6715
rect 13401 6671 13411 6705
rect 13411 6671 13445 6705
rect 13445 6671 13453 6705
rect 13401 6663 13453 6671
rect 15797 6662 15849 6673
rect 15248 6633 15300 6640
rect 15248 6599 15256 6633
rect 15256 6599 15290 6633
rect 15290 6599 15300 6633
rect 15248 6588 15300 6599
rect 15797 6628 15806 6662
rect 15806 6628 15840 6662
rect 15840 6628 15849 6662
rect 15797 6621 15849 6628
rect 14490 6524 14542 6576
rect 17641 6634 17693 6641
rect 17641 6600 17649 6634
rect 17649 6600 17683 6634
rect 17683 6600 17693 6634
rect 17641 6589 17693 6600
rect 16885 6524 16937 6576
rect 13536 6305 13588 6357
rect 13752 6310 13804 6362
rect 13958 6311 14010 6363
rect 14160 6303 14212 6355
rect 14356 6305 14408 6357
rect 14581 6307 14633 6359
rect 14796 6303 14848 6355
rect 15031 6303 15083 6355
rect 15239 6306 15291 6358
rect 15481 6306 15533 6358
rect 15679 6307 15731 6359
rect 15986 6307 16038 6359
rect 16211 6308 16263 6360
rect 16440 6307 16492 6359
rect 16656 6311 16708 6363
rect 16879 6314 16931 6366
rect 17103 6310 17155 6362
rect 17330 6299 17382 6351
rect 17543 6298 17595 6350
rect 17754 6302 17806 6354
rect 17981 6303 18033 6355
rect 13409 6089 13461 6100
rect 13409 6055 13419 6089
rect 13419 6055 13453 6089
rect 13453 6055 13461 6089
rect 14870 6076 14922 6128
rect 13409 6048 13461 6055
rect 15253 6063 15305 6069
rect 15253 6029 15265 6063
rect 15265 6029 15299 6063
rect 15299 6029 15305 6063
rect 15253 6017 15305 6029
rect 15796 6045 15848 6057
rect 15796 6011 15803 6045
rect 15803 6011 15837 6045
rect 15837 6011 15848 6045
rect 17262 6078 17314 6130
rect 17639 6065 17691 6076
rect 17639 6031 17649 6065
rect 17649 6031 17683 6065
rect 17683 6031 17691 6065
rect 17639 6024 17691 6031
rect 15796 6005 15848 6011
rect 13562 5660 13614 5712
rect 13787 5669 13839 5721
rect 14064 5666 14116 5718
rect 14285 5669 14337 5721
rect 14530 5666 14582 5718
rect 14756 5670 14808 5722
rect 14968 5668 15020 5720
rect 15188 5674 15240 5726
rect 15426 5676 15478 5728
rect 15639 5678 15691 5730
rect 16026 5668 16078 5720
rect 16373 5669 16425 5721
rect 16609 5664 16661 5716
rect 16793 5664 16845 5716
rect 17032 5666 17084 5718
rect 17235 5662 17287 5714
rect 17420 5659 17472 5711
rect 17611 5661 17663 5713
rect 17802 5665 17854 5717
rect 17988 5661 18040 5713
rect 13404 5329 13456 5340
rect 13404 5295 13415 5329
rect 13415 5295 13449 5329
rect 13449 5295 13456 5329
rect 15248 5353 15300 5361
rect 15248 5319 15257 5353
rect 15257 5319 15291 5353
rect 15291 5319 15300 5353
rect 15248 5309 15300 5319
rect 15797 5359 15849 5370
rect 15797 5325 15804 5359
rect 15804 5325 15838 5359
rect 15838 5325 15849 5359
rect 15797 5318 15849 5325
rect 13404 5288 13456 5295
rect 14499 5244 14551 5296
rect 17640 5354 17692 5362
rect 17640 5320 17649 5354
rect 17649 5320 17683 5354
rect 17683 5320 17692 5354
rect 17640 5310 17692 5320
rect 16889 5244 16942 5296
rect 13435 5078 13487 5130
rect 13640 5074 13692 5126
rect 13826 5079 13878 5131
rect 14020 5072 14072 5124
rect 14239 5077 14291 5129
rect 14449 5077 14501 5129
rect 14678 5074 14730 5126
rect 14924 5074 14976 5126
rect 15198 5074 15250 5126
rect 15473 5074 15525 5126
rect 15709 5074 15761 5126
rect 15932 5077 15984 5129
rect 16150 5080 16202 5132
rect 16328 5071 16380 5123
rect 16567 5073 16619 5125
rect 16764 5073 16816 5125
rect 16962 5073 17014 5125
rect 17175 5074 17227 5126
rect 17398 5073 17450 5125
rect 17595 5078 17647 5130
rect 17811 5076 17863 5128
rect 18020 5076 18072 5128
<< metal2 >>
rect 18572 9695 18646 9699
rect 18572 9639 18581 9695
rect 18637 9639 18646 9695
rect 18572 9635 18646 9639
rect 18772 9695 18846 9699
rect 18772 9639 18781 9695
rect 18837 9639 18846 9695
rect 18772 9635 18846 9639
rect 18383 9053 18457 9057
rect 18383 8997 18392 9053
rect 18448 8997 18457 9053
rect 18383 8993 18457 8997
rect 13409 7655 13415 7707
rect 13467 7655 13473 7707
rect 15803 7655 15809 7707
rect 15861 7655 15867 7707
rect 13428 7370 13456 7655
rect 13496 7535 13505 7591
rect 13561 7535 13571 7591
rect 13496 7534 13571 7535
rect 13670 7534 13679 7590
rect 13735 7534 13745 7590
rect 13895 7536 13904 7592
rect 13960 7536 13970 7592
rect 14096 7538 14105 7594
rect 14161 7538 14171 7594
rect 14096 7537 14171 7538
rect 13895 7535 13970 7536
rect 14319 7536 14328 7592
rect 14384 7536 14394 7592
rect 14528 7541 14537 7597
rect 14593 7541 14603 7597
rect 14528 7540 14603 7541
rect 14319 7535 14394 7536
rect 13670 7533 13745 7534
rect 14756 7534 14765 7590
rect 14821 7534 14831 7590
rect 14946 7538 14955 7594
rect 15011 7538 15021 7594
rect 15151 7541 15160 7597
rect 15216 7541 15226 7597
rect 15151 7540 15226 7541
rect 15350 7541 15359 7597
rect 15415 7541 15425 7597
rect 15350 7540 15425 7541
rect 14946 7537 15021 7538
rect 15566 7536 15575 7592
rect 15631 7536 15641 7592
rect 15566 7535 15641 7536
rect 14756 7533 14831 7534
rect 13406 7364 13458 7370
rect 14854 7348 14863 7404
rect 14919 7348 14929 7404
rect 14854 7347 14929 7348
rect 13406 7306 13458 7312
rect 13428 6721 13456 7306
rect 15239 7297 15248 7353
rect 15304 7297 15314 7353
rect 15822 7328 15850 7655
rect 15954 7541 15963 7597
rect 16019 7541 16029 7597
rect 15954 7540 16029 7541
rect 16189 7536 16198 7592
rect 16254 7536 16264 7592
rect 16431 7538 16440 7594
rect 16496 7538 16506 7594
rect 16663 7539 16672 7595
rect 16728 7539 16738 7595
rect 16892 7542 16901 7598
rect 16957 7542 16967 7598
rect 16892 7541 16967 7542
rect 16663 7538 16738 7539
rect 16431 7537 16506 7538
rect 16189 7535 16264 7536
rect 17141 7534 17150 7590
rect 17206 7534 17216 7590
rect 17359 7538 17368 7594
rect 17424 7538 17434 7594
rect 17359 7537 17434 7538
rect 17141 7533 17216 7534
rect 17588 7534 17597 7590
rect 17653 7534 17663 7590
rect 17809 7536 17818 7592
rect 17874 7536 17884 7592
rect 18025 7541 18034 7597
rect 18090 7541 18100 7597
rect 18025 7540 18100 7541
rect 17809 7535 17884 7536
rect 17588 7533 17663 7534
rect 17249 7347 17258 7403
rect 17314 7347 17324 7403
rect 17249 7346 17324 7347
rect 15239 7296 15314 7297
rect 15798 7322 15850 7328
rect 17634 7298 17643 7354
rect 17699 7298 17709 7354
rect 17634 7297 17709 7298
rect 15798 7264 15850 7270
rect 13498 6952 13507 7008
rect 13563 6952 13573 7008
rect 13498 6951 13573 6952
rect 13673 6950 13682 7006
rect 13738 6950 13748 7006
rect 13870 6952 13879 7008
rect 13935 6952 13945 7008
rect 14089 6955 14098 7011
rect 14154 6955 14164 7011
rect 14089 6954 14164 6955
rect 13870 6951 13945 6952
rect 14321 6951 14330 7007
rect 14386 6951 14396 7007
rect 14321 6950 14396 6951
rect 14505 6958 14554 7014
rect 14610 6958 14620 7014
rect 13673 6949 13748 6950
rect 13401 6715 13456 6721
rect 13453 6663 13456 6715
rect 13401 6657 13456 6663
rect 13428 6106 13456 6657
rect 14505 6905 14620 6958
rect 14757 6946 14766 7002
rect 14822 6946 14832 7002
rect 14757 6945 14832 6946
rect 14979 6942 14988 6998
rect 15044 6942 15054 6998
rect 14979 6941 15054 6942
rect 15201 6995 15289 7000
rect 15201 6939 15211 6995
rect 15267 6939 15289 6995
rect 15201 6919 15289 6939
rect 15412 6939 15421 6995
rect 15477 6939 15487 6995
rect 15412 6938 15487 6939
rect 15625 6939 15634 6995
rect 15690 6939 15700 6995
rect 15625 6938 15700 6939
rect 14505 6576 14549 6905
rect 15253 6640 15289 6919
rect 15822 6679 15850 7264
rect 15942 6932 15951 6988
rect 16007 6932 16017 6988
rect 16144 6935 16153 6991
rect 16209 6935 16219 6991
rect 16345 6936 16354 6992
rect 16410 6936 16420 6992
rect 16524 6937 16533 6993
rect 16589 6937 16599 6993
rect 16716 6941 16725 6997
rect 16781 6941 16791 6997
rect 16716 6940 16791 6941
rect 16889 6994 16977 6998
rect 16524 6936 16599 6937
rect 16889 6938 16910 6994
rect 16966 6938 16977 6994
rect 16345 6935 16420 6936
rect 16144 6934 16219 6935
rect 15942 6931 16017 6932
rect 15797 6673 15850 6679
rect 15242 6588 15248 6640
rect 15300 6588 15306 6640
rect 15849 6621 15850 6673
rect 15797 6615 15850 6621
rect 14484 6524 14490 6576
rect 14542 6559 14549 6576
rect 14542 6524 14548 6559
rect 14484 6523 14548 6524
rect 13525 6303 13534 6359
rect 13590 6303 13600 6359
rect 13741 6308 13750 6364
rect 13806 6308 13816 6364
rect 13947 6309 13956 6365
rect 14012 6309 14022 6365
rect 13947 6308 14022 6309
rect 13741 6307 13816 6308
rect 13525 6302 13600 6303
rect 14149 6301 14158 6357
rect 14214 6301 14224 6357
rect 14345 6303 14354 6359
rect 14410 6303 14420 6359
rect 14570 6305 14579 6361
rect 14635 6305 14645 6361
rect 14570 6304 14645 6305
rect 14345 6302 14420 6303
rect 14149 6300 14224 6301
rect 14785 6301 14794 6357
rect 14850 6301 14860 6357
rect 14785 6300 14860 6301
rect 15020 6301 15029 6357
rect 15085 6301 15095 6357
rect 15228 6304 15237 6360
rect 15293 6304 15303 6360
rect 15228 6303 15303 6304
rect 15470 6304 15479 6360
rect 15535 6304 15545 6360
rect 15668 6305 15677 6361
rect 15733 6305 15743 6361
rect 15668 6304 15743 6305
rect 15470 6303 15545 6304
rect 15020 6300 15095 6301
rect 13409 6100 13461 6106
rect 14859 6074 14868 6130
rect 14924 6074 14934 6130
rect 14859 6073 14934 6074
rect 13409 6042 13461 6048
rect 13428 5346 13456 6042
rect 15242 6015 15251 6071
rect 15307 6015 15317 6071
rect 15822 6063 15850 6615
rect 16889 6923 16977 6938
rect 17133 6937 17142 6993
rect 17198 6937 17208 6993
rect 17338 6939 17347 6995
rect 17403 6939 17413 6995
rect 17544 6941 17553 6997
rect 17609 6941 17619 6997
rect 17544 6940 17619 6941
rect 17649 6940 17655 6992
rect 17707 6940 17713 6992
rect 17752 6948 17761 7004
rect 17817 6948 17827 7004
rect 17974 6949 17983 7005
rect 18039 6949 18049 7005
rect 17974 6948 18049 6949
rect 17752 6947 17827 6948
rect 17338 6938 17413 6939
rect 17133 6936 17208 6937
rect 16889 6576 16933 6923
rect 17649 6641 17699 6940
rect 17635 6589 17641 6641
rect 17693 6589 17699 6641
rect 16879 6524 16885 6576
rect 16937 6524 16943 6576
rect 15975 6305 15984 6361
rect 16040 6305 16050 6361
rect 16200 6306 16209 6362
rect 16265 6306 16275 6362
rect 16200 6305 16275 6306
rect 16429 6305 16438 6361
rect 16494 6305 16504 6361
rect 16645 6309 16654 6365
rect 16710 6309 16720 6365
rect 16868 6312 16877 6368
rect 16933 6312 16943 6368
rect 16868 6311 16943 6312
rect 16645 6308 16720 6309
rect 17092 6308 17101 6364
rect 17157 6308 17167 6364
rect 17092 6307 17167 6308
rect 15975 6304 16050 6305
rect 16429 6304 16504 6305
rect 17319 6297 17328 6353
rect 17384 6297 17394 6353
rect 17319 6296 17394 6297
rect 17532 6296 17541 6352
rect 17597 6296 17607 6352
rect 17743 6300 17752 6356
rect 17808 6300 17818 6356
rect 17970 6301 17979 6357
rect 18035 6301 18045 6357
rect 17970 6300 18045 6301
rect 17743 6299 17818 6300
rect 17532 6295 17607 6296
rect 17251 6076 17260 6132
rect 17316 6076 17326 6132
rect 17251 6075 17326 6076
rect 15242 6014 15317 6015
rect 15796 6057 15850 6063
rect 15848 6005 15850 6057
rect 17628 6022 17637 6078
rect 17693 6022 17703 6078
rect 17628 6021 17703 6022
rect 15796 5999 15850 6005
rect 13551 5658 13560 5714
rect 13616 5658 13626 5714
rect 13776 5667 13785 5723
rect 13841 5667 13851 5723
rect 13776 5666 13851 5667
rect 14053 5664 14062 5720
rect 14118 5664 14128 5720
rect 14274 5667 14283 5723
rect 14339 5667 14349 5723
rect 14274 5666 14349 5667
rect 14490 5720 14558 5722
rect 14053 5663 14128 5664
rect 14490 5664 14528 5720
rect 14584 5664 14594 5720
rect 14745 5668 14754 5724
rect 14810 5668 14820 5724
rect 14745 5667 14820 5668
rect 14957 5666 14966 5722
rect 15022 5666 15032 5722
rect 15177 5672 15186 5728
rect 15242 5725 15252 5728
rect 15242 5672 15291 5725
rect 15415 5674 15424 5730
rect 15480 5674 15490 5730
rect 15628 5676 15637 5732
rect 15693 5676 15703 5732
rect 15628 5675 15703 5676
rect 15415 5673 15490 5674
rect 15177 5671 15291 5672
rect 14957 5665 15032 5666
rect 14490 5663 14594 5664
rect 13551 5657 13626 5658
rect 13404 5340 13456 5346
rect 14507 5296 14543 5663
rect 15246 5362 15291 5671
rect 15822 5376 15850 5999
rect 16015 5666 16024 5722
rect 16080 5666 16090 5722
rect 16362 5667 16371 5723
rect 16427 5667 16437 5723
rect 16779 5720 17096 5726
rect 16779 5718 17030 5720
rect 16362 5666 16437 5667
rect 16015 5665 16090 5666
rect 16598 5662 16607 5718
rect 16663 5662 16673 5718
rect 16598 5661 16673 5662
rect 16779 5662 16791 5718
rect 16847 5664 17030 5718
rect 17086 5664 17096 5720
rect 16847 5662 17096 5664
rect 16779 5651 17096 5662
rect 17224 5660 17233 5716
rect 17289 5660 17299 5716
rect 17224 5659 17299 5660
rect 17409 5657 17418 5713
rect 17474 5657 17484 5713
rect 17600 5659 17609 5715
rect 17665 5712 17675 5715
rect 17665 5659 17688 5712
rect 17791 5663 17800 5719
rect 17856 5663 17866 5719
rect 17791 5662 17866 5663
rect 17600 5658 17688 5659
rect 17977 5659 17986 5715
rect 18042 5659 18052 5715
rect 17977 5658 18052 5659
rect 17409 5656 17484 5657
rect 15797 5370 15850 5376
rect 15242 5361 15307 5362
rect 15242 5309 15248 5361
rect 15300 5309 15307 5361
rect 15849 5318 15850 5370
rect 15797 5312 15850 5318
rect 13404 5282 13456 5288
rect 13428 5281 13456 5282
rect 14490 5257 14499 5296
rect 14491 5244 14499 5257
rect 14551 5257 14558 5296
rect 15822 5294 15850 5312
rect 16900 5296 16936 5651
rect 17651 5363 17688 5658
rect 17634 5362 17698 5363
rect 17634 5310 17640 5362
rect 17692 5310 17698 5362
rect 14551 5244 14557 5257
rect 16882 5244 16889 5296
rect 16942 5244 16949 5296
rect 13424 5076 13433 5132
rect 13489 5076 13499 5132
rect 13424 5075 13499 5076
rect 13629 5072 13638 5128
rect 13694 5072 13704 5128
rect 13815 5077 13824 5133
rect 13880 5077 13890 5133
rect 13815 5076 13890 5077
rect 13629 5071 13704 5072
rect 14009 5070 14018 5126
rect 14074 5070 14084 5126
rect 14228 5075 14237 5131
rect 14293 5075 14303 5131
rect 14228 5074 14303 5075
rect 14438 5075 14447 5131
rect 14503 5075 14513 5131
rect 14438 5074 14513 5075
rect 14667 5072 14676 5128
rect 14732 5072 14742 5128
rect 14667 5071 14742 5072
rect 14913 5072 14922 5128
rect 14978 5072 14988 5128
rect 14913 5071 14988 5072
rect 15187 5072 15196 5128
rect 15252 5072 15262 5128
rect 15187 5071 15262 5072
rect 15462 5072 15471 5128
rect 15527 5072 15537 5128
rect 15462 5071 15537 5072
rect 15698 5072 15707 5128
rect 15763 5072 15773 5128
rect 15921 5075 15930 5131
rect 15986 5075 15996 5131
rect 16139 5078 16148 5134
rect 16204 5078 16214 5134
rect 16139 5077 16214 5078
rect 15921 5074 15996 5075
rect 15698 5071 15773 5072
rect 14009 5069 14084 5070
rect 16317 5069 16326 5125
rect 16382 5069 16392 5125
rect 16556 5071 16565 5127
rect 16621 5071 16631 5127
rect 16556 5070 16631 5071
rect 16753 5071 16762 5127
rect 16818 5071 16828 5127
rect 16753 5070 16828 5071
rect 16951 5071 16960 5127
rect 17016 5071 17026 5127
rect 17164 5072 17173 5128
rect 17229 5072 17239 5128
rect 17164 5071 17239 5072
rect 17387 5071 17396 5127
rect 17452 5071 17462 5127
rect 17584 5076 17593 5132
rect 17649 5076 17659 5132
rect 17584 5075 17659 5076
rect 17800 5074 17809 5130
rect 17865 5074 17875 5130
rect 17800 5073 17875 5074
rect 18009 5074 18018 5130
rect 18074 5074 18084 5130
rect 18009 5073 18084 5074
rect 16951 5070 17026 5071
rect 17387 5070 17462 5071
rect 16317 5068 16392 5069
<< via2 >>
rect 18581 9693 18637 9695
rect 18581 9641 18583 9693
rect 18583 9641 18635 9693
rect 18635 9641 18637 9693
rect 18581 9639 18637 9641
rect 18781 9693 18837 9695
rect 18781 9641 18783 9693
rect 18783 9641 18835 9693
rect 18835 9641 18837 9693
rect 18781 9639 18837 9641
rect 18392 9051 18448 9053
rect 18392 8999 18394 9051
rect 18394 8999 18446 9051
rect 18446 8999 18448 9051
rect 18392 8997 18448 8999
rect 13505 7589 13561 7591
rect 13505 7537 13507 7589
rect 13507 7537 13559 7589
rect 13559 7537 13561 7589
rect 13505 7535 13561 7537
rect 13679 7588 13735 7590
rect 13679 7536 13681 7588
rect 13681 7536 13733 7588
rect 13733 7536 13735 7588
rect 13679 7534 13735 7536
rect 13904 7590 13960 7592
rect 13904 7538 13906 7590
rect 13906 7538 13958 7590
rect 13958 7538 13960 7590
rect 13904 7536 13960 7538
rect 14105 7592 14161 7594
rect 14105 7540 14107 7592
rect 14107 7540 14159 7592
rect 14159 7540 14161 7592
rect 14105 7538 14161 7540
rect 14328 7590 14384 7592
rect 14328 7538 14330 7590
rect 14330 7538 14382 7590
rect 14382 7538 14384 7590
rect 14328 7536 14384 7538
rect 14537 7595 14593 7597
rect 14537 7543 14539 7595
rect 14539 7543 14591 7595
rect 14591 7543 14593 7595
rect 14537 7541 14593 7543
rect 14765 7588 14821 7590
rect 14765 7536 14767 7588
rect 14767 7536 14819 7588
rect 14819 7536 14821 7588
rect 14765 7534 14821 7536
rect 14955 7592 15011 7594
rect 14955 7540 14957 7592
rect 14957 7540 15009 7592
rect 15009 7540 15011 7592
rect 14955 7538 15011 7540
rect 15160 7595 15216 7597
rect 15160 7543 15162 7595
rect 15162 7543 15214 7595
rect 15214 7543 15216 7595
rect 15160 7541 15216 7543
rect 15359 7595 15415 7597
rect 15359 7543 15361 7595
rect 15361 7543 15413 7595
rect 15413 7543 15415 7595
rect 15359 7541 15415 7543
rect 15575 7590 15631 7592
rect 15575 7538 15577 7590
rect 15577 7538 15629 7590
rect 15629 7538 15631 7590
rect 15575 7536 15631 7538
rect 14863 7402 14919 7404
rect 14863 7350 14865 7402
rect 14865 7350 14917 7402
rect 14917 7350 14919 7402
rect 14863 7348 14919 7350
rect 15248 7351 15304 7353
rect 15248 7299 15250 7351
rect 15250 7299 15302 7351
rect 15302 7299 15304 7351
rect 15248 7297 15304 7299
rect 15963 7595 16019 7597
rect 15963 7543 15965 7595
rect 15965 7543 16017 7595
rect 16017 7543 16019 7595
rect 15963 7541 16019 7543
rect 16198 7590 16254 7592
rect 16198 7538 16200 7590
rect 16200 7538 16252 7590
rect 16252 7538 16254 7590
rect 16198 7536 16254 7538
rect 16440 7592 16496 7594
rect 16440 7540 16442 7592
rect 16442 7540 16494 7592
rect 16494 7540 16496 7592
rect 16440 7538 16496 7540
rect 16672 7593 16728 7595
rect 16672 7541 16674 7593
rect 16674 7541 16726 7593
rect 16726 7541 16728 7593
rect 16672 7539 16728 7541
rect 16901 7596 16957 7598
rect 16901 7544 16903 7596
rect 16903 7544 16955 7596
rect 16955 7544 16957 7596
rect 16901 7542 16957 7544
rect 17150 7588 17206 7590
rect 17150 7536 17152 7588
rect 17152 7536 17204 7588
rect 17204 7536 17206 7588
rect 17150 7534 17206 7536
rect 17368 7592 17424 7594
rect 17368 7540 17370 7592
rect 17370 7540 17422 7592
rect 17422 7540 17424 7592
rect 17368 7538 17424 7540
rect 17597 7588 17653 7590
rect 17597 7536 17599 7588
rect 17599 7536 17651 7588
rect 17651 7536 17653 7588
rect 17597 7534 17653 7536
rect 17818 7590 17874 7592
rect 17818 7538 17820 7590
rect 17820 7538 17872 7590
rect 17872 7538 17874 7590
rect 17818 7536 17874 7538
rect 18034 7595 18090 7597
rect 18034 7543 18036 7595
rect 18036 7543 18088 7595
rect 18088 7543 18090 7595
rect 18034 7541 18090 7543
rect 17258 7401 17314 7403
rect 17258 7349 17260 7401
rect 17260 7349 17312 7401
rect 17312 7349 17314 7401
rect 17258 7347 17314 7349
rect 17643 7352 17699 7354
rect 17643 7300 17645 7352
rect 17645 7300 17697 7352
rect 17697 7300 17699 7352
rect 17643 7298 17699 7300
rect 13507 7006 13563 7008
rect 13507 6954 13509 7006
rect 13509 6954 13561 7006
rect 13561 6954 13563 7006
rect 13507 6952 13563 6954
rect 13682 7004 13738 7006
rect 13682 6952 13684 7004
rect 13684 6952 13736 7004
rect 13736 6952 13738 7004
rect 13682 6950 13738 6952
rect 13879 7006 13935 7008
rect 13879 6954 13881 7006
rect 13881 6954 13933 7006
rect 13933 6954 13935 7006
rect 13879 6952 13935 6954
rect 14098 7009 14154 7011
rect 14098 6957 14100 7009
rect 14100 6957 14152 7009
rect 14152 6957 14154 7009
rect 14098 6955 14154 6957
rect 14330 7005 14386 7007
rect 14330 6953 14332 7005
rect 14332 6953 14384 7005
rect 14384 6953 14386 7005
rect 14330 6951 14386 6953
rect 14554 7012 14610 7014
rect 14554 6960 14556 7012
rect 14556 6960 14608 7012
rect 14608 6960 14610 7012
rect 14554 6958 14610 6960
rect 14766 7000 14822 7002
rect 14766 6948 14768 7000
rect 14768 6948 14820 7000
rect 14820 6948 14822 7000
rect 14766 6946 14822 6948
rect 14988 6996 15044 6998
rect 14988 6944 14990 6996
rect 14990 6944 15042 6996
rect 15042 6944 15044 6996
rect 14988 6942 15044 6944
rect 15211 6993 15267 6995
rect 15211 6941 15213 6993
rect 15213 6941 15265 6993
rect 15265 6941 15267 6993
rect 15211 6939 15267 6941
rect 15421 6993 15477 6995
rect 15421 6941 15423 6993
rect 15423 6941 15475 6993
rect 15475 6941 15477 6993
rect 15421 6939 15477 6941
rect 15634 6993 15690 6995
rect 15634 6941 15636 6993
rect 15636 6941 15688 6993
rect 15688 6941 15690 6993
rect 15634 6939 15690 6941
rect 15951 6986 16007 6988
rect 15951 6934 15953 6986
rect 15953 6934 16005 6986
rect 16005 6934 16007 6986
rect 15951 6932 16007 6934
rect 16153 6989 16209 6991
rect 16153 6937 16155 6989
rect 16155 6937 16207 6989
rect 16207 6937 16209 6989
rect 16153 6935 16209 6937
rect 16354 6990 16410 6992
rect 16354 6938 16356 6990
rect 16356 6938 16408 6990
rect 16408 6938 16410 6990
rect 16354 6936 16410 6938
rect 16533 6991 16589 6993
rect 16533 6939 16535 6991
rect 16535 6939 16587 6991
rect 16587 6939 16589 6991
rect 16533 6937 16589 6939
rect 16725 6995 16781 6997
rect 16725 6943 16727 6995
rect 16727 6943 16779 6995
rect 16779 6943 16781 6995
rect 16725 6941 16781 6943
rect 16910 6992 16966 6994
rect 16910 6940 16912 6992
rect 16912 6940 16964 6992
rect 16964 6940 16966 6992
rect 16910 6938 16966 6940
rect 13534 6357 13590 6359
rect 13534 6305 13536 6357
rect 13536 6305 13588 6357
rect 13588 6305 13590 6357
rect 13534 6303 13590 6305
rect 13750 6362 13806 6364
rect 13750 6310 13752 6362
rect 13752 6310 13804 6362
rect 13804 6310 13806 6362
rect 13750 6308 13806 6310
rect 13956 6363 14012 6365
rect 13956 6311 13958 6363
rect 13958 6311 14010 6363
rect 14010 6311 14012 6363
rect 13956 6309 14012 6311
rect 14158 6355 14214 6357
rect 14158 6303 14160 6355
rect 14160 6303 14212 6355
rect 14212 6303 14214 6355
rect 14158 6301 14214 6303
rect 14354 6357 14410 6359
rect 14354 6305 14356 6357
rect 14356 6305 14408 6357
rect 14408 6305 14410 6357
rect 14354 6303 14410 6305
rect 14579 6359 14635 6361
rect 14579 6307 14581 6359
rect 14581 6307 14633 6359
rect 14633 6307 14635 6359
rect 14579 6305 14635 6307
rect 14794 6355 14850 6357
rect 14794 6303 14796 6355
rect 14796 6303 14848 6355
rect 14848 6303 14850 6355
rect 14794 6301 14850 6303
rect 15029 6355 15085 6357
rect 15029 6303 15031 6355
rect 15031 6303 15083 6355
rect 15083 6303 15085 6355
rect 15029 6301 15085 6303
rect 15237 6358 15293 6360
rect 15237 6306 15239 6358
rect 15239 6306 15291 6358
rect 15291 6306 15293 6358
rect 15237 6304 15293 6306
rect 15479 6358 15535 6360
rect 15479 6306 15481 6358
rect 15481 6306 15533 6358
rect 15533 6306 15535 6358
rect 15479 6304 15535 6306
rect 15677 6359 15733 6361
rect 15677 6307 15679 6359
rect 15679 6307 15731 6359
rect 15731 6307 15733 6359
rect 15677 6305 15733 6307
rect 14868 6128 14924 6130
rect 14868 6076 14870 6128
rect 14870 6076 14922 6128
rect 14922 6076 14924 6128
rect 14868 6074 14924 6076
rect 15251 6069 15307 6071
rect 15251 6017 15253 6069
rect 15253 6017 15305 6069
rect 15305 6017 15307 6069
rect 15251 6015 15307 6017
rect 17142 6991 17198 6993
rect 17142 6939 17144 6991
rect 17144 6939 17196 6991
rect 17196 6939 17198 6991
rect 17142 6937 17198 6939
rect 17347 6993 17403 6995
rect 17347 6941 17349 6993
rect 17349 6941 17401 6993
rect 17401 6941 17403 6993
rect 17347 6939 17403 6941
rect 17553 6995 17609 6997
rect 17553 6943 17555 6995
rect 17555 6943 17607 6995
rect 17607 6943 17609 6995
rect 17553 6941 17609 6943
rect 17761 7002 17817 7004
rect 17761 6950 17763 7002
rect 17763 6950 17815 7002
rect 17815 6950 17817 7002
rect 17761 6948 17817 6950
rect 17983 7003 18039 7005
rect 17983 6951 17985 7003
rect 17985 6951 18037 7003
rect 18037 6951 18039 7003
rect 17983 6949 18039 6951
rect 15984 6359 16040 6361
rect 15984 6307 15986 6359
rect 15986 6307 16038 6359
rect 16038 6307 16040 6359
rect 15984 6305 16040 6307
rect 16209 6360 16265 6362
rect 16209 6308 16211 6360
rect 16211 6308 16263 6360
rect 16263 6308 16265 6360
rect 16209 6306 16265 6308
rect 16438 6359 16494 6361
rect 16438 6307 16440 6359
rect 16440 6307 16492 6359
rect 16492 6307 16494 6359
rect 16438 6305 16494 6307
rect 16654 6363 16710 6365
rect 16654 6311 16656 6363
rect 16656 6311 16708 6363
rect 16708 6311 16710 6363
rect 16654 6309 16710 6311
rect 16877 6366 16933 6368
rect 16877 6314 16879 6366
rect 16879 6314 16931 6366
rect 16931 6314 16933 6366
rect 16877 6312 16933 6314
rect 17101 6362 17157 6364
rect 17101 6310 17103 6362
rect 17103 6310 17155 6362
rect 17155 6310 17157 6362
rect 17101 6308 17157 6310
rect 17328 6351 17384 6353
rect 17328 6299 17330 6351
rect 17330 6299 17382 6351
rect 17382 6299 17384 6351
rect 17328 6297 17384 6299
rect 17541 6350 17597 6352
rect 17541 6298 17543 6350
rect 17543 6298 17595 6350
rect 17595 6298 17597 6350
rect 17541 6296 17597 6298
rect 17752 6354 17808 6356
rect 17752 6302 17754 6354
rect 17754 6302 17806 6354
rect 17806 6302 17808 6354
rect 17752 6300 17808 6302
rect 17979 6355 18035 6357
rect 17979 6303 17981 6355
rect 17981 6303 18033 6355
rect 18033 6303 18035 6355
rect 17979 6301 18035 6303
rect 17260 6130 17316 6132
rect 17260 6078 17262 6130
rect 17262 6078 17314 6130
rect 17314 6078 17316 6130
rect 17260 6076 17316 6078
rect 17637 6076 17693 6078
rect 17637 6024 17639 6076
rect 17639 6024 17691 6076
rect 17691 6024 17693 6076
rect 17637 6022 17693 6024
rect 13560 5712 13616 5714
rect 13560 5660 13562 5712
rect 13562 5660 13614 5712
rect 13614 5660 13616 5712
rect 13560 5658 13616 5660
rect 13785 5721 13841 5723
rect 13785 5669 13787 5721
rect 13787 5669 13839 5721
rect 13839 5669 13841 5721
rect 13785 5667 13841 5669
rect 14062 5718 14118 5720
rect 14062 5666 14064 5718
rect 14064 5666 14116 5718
rect 14116 5666 14118 5718
rect 14062 5664 14118 5666
rect 14283 5721 14339 5723
rect 14283 5669 14285 5721
rect 14285 5669 14337 5721
rect 14337 5669 14339 5721
rect 14283 5667 14339 5669
rect 14528 5718 14584 5720
rect 14528 5666 14530 5718
rect 14530 5666 14582 5718
rect 14582 5666 14584 5718
rect 14528 5664 14584 5666
rect 14754 5722 14810 5724
rect 14754 5670 14756 5722
rect 14756 5670 14808 5722
rect 14808 5670 14810 5722
rect 14754 5668 14810 5670
rect 14966 5720 15022 5722
rect 14966 5668 14968 5720
rect 14968 5668 15020 5720
rect 15020 5668 15022 5720
rect 14966 5666 15022 5668
rect 15186 5726 15242 5728
rect 15186 5674 15188 5726
rect 15188 5674 15240 5726
rect 15240 5674 15242 5726
rect 15186 5672 15242 5674
rect 15424 5728 15480 5730
rect 15424 5676 15426 5728
rect 15426 5676 15478 5728
rect 15478 5676 15480 5728
rect 15424 5674 15480 5676
rect 15637 5730 15693 5732
rect 15637 5678 15639 5730
rect 15639 5678 15691 5730
rect 15691 5678 15693 5730
rect 15637 5676 15693 5678
rect 16024 5720 16080 5722
rect 16024 5668 16026 5720
rect 16026 5668 16078 5720
rect 16078 5668 16080 5720
rect 16024 5666 16080 5668
rect 16371 5721 16427 5723
rect 16371 5669 16373 5721
rect 16373 5669 16425 5721
rect 16425 5669 16427 5721
rect 16371 5667 16427 5669
rect 17030 5718 17086 5720
rect 16607 5716 16663 5718
rect 16607 5664 16609 5716
rect 16609 5664 16661 5716
rect 16661 5664 16663 5716
rect 16607 5662 16663 5664
rect 16791 5716 16847 5718
rect 16791 5664 16793 5716
rect 16793 5664 16845 5716
rect 16845 5664 16847 5716
rect 17030 5666 17032 5718
rect 17032 5666 17084 5718
rect 17084 5666 17086 5718
rect 17030 5664 17086 5666
rect 16791 5662 16847 5664
rect 17233 5714 17289 5716
rect 17233 5662 17235 5714
rect 17235 5662 17287 5714
rect 17287 5662 17289 5714
rect 17233 5660 17289 5662
rect 17418 5711 17474 5713
rect 17418 5659 17420 5711
rect 17420 5659 17472 5711
rect 17472 5659 17474 5711
rect 17418 5657 17474 5659
rect 17609 5713 17665 5715
rect 17609 5661 17611 5713
rect 17611 5661 17663 5713
rect 17663 5661 17665 5713
rect 17609 5659 17665 5661
rect 17800 5717 17856 5719
rect 17800 5665 17802 5717
rect 17802 5665 17854 5717
rect 17854 5665 17856 5717
rect 17800 5663 17856 5665
rect 17986 5713 18042 5715
rect 17986 5661 17988 5713
rect 17988 5661 18040 5713
rect 18040 5661 18042 5713
rect 17986 5659 18042 5661
rect 13433 5130 13489 5132
rect 13433 5078 13435 5130
rect 13435 5078 13487 5130
rect 13487 5078 13489 5130
rect 13433 5076 13489 5078
rect 13638 5126 13694 5128
rect 13638 5074 13640 5126
rect 13640 5074 13692 5126
rect 13692 5074 13694 5126
rect 13638 5072 13694 5074
rect 13824 5131 13880 5133
rect 13824 5079 13826 5131
rect 13826 5079 13878 5131
rect 13878 5079 13880 5131
rect 13824 5077 13880 5079
rect 14018 5124 14074 5126
rect 14018 5072 14020 5124
rect 14020 5072 14072 5124
rect 14072 5072 14074 5124
rect 14018 5070 14074 5072
rect 14237 5129 14293 5131
rect 14237 5077 14239 5129
rect 14239 5077 14291 5129
rect 14291 5077 14293 5129
rect 14237 5075 14293 5077
rect 14447 5129 14503 5131
rect 14447 5077 14449 5129
rect 14449 5077 14501 5129
rect 14501 5077 14503 5129
rect 14447 5075 14503 5077
rect 14676 5126 14732 5128
rect 14676 5074 14678 5126
rect 14678 5074 14730 5126
rect 14730 5074 14732 5126
rect 14676 5072 14732 5074
rect 14922 5126 14978 5128
rect 14922 5074 14924 5126
rect 14924 5074 14976 5126
rect 14976 5074 14978 5126
rect 14922 5072 14978 5074
rect 15196 5126 15252 5128
rect 15196 5074 15198 5126
rect 15198 5074 15250 5126
rect 15250 5074 15252 5126
rect 15196 5072 15252 5074
rect 15471 5126 15527 5128
rect 15471 5074 15473 5126
rect 15473 5074 15525 5126
rect 15525 5074 15527 5126
rect 15471 5072 15527 5074
rect 15707 5126 15763 5128
rect 15707 5074 15709 5126
rect 15709 5074 15761 5126
rect 15761 5074 15763 5126
rect 15707 5072 15763 5074
rect 15930 5129 15986 5131
rect 15930 5077 15932 5129
rect 15932 5077 15984 5129
rect 15984 5077 15986 5129
rect 15930 5075 15986 5077
rect 16148 5132 16204 5134
rect 16148 5080 16150 5132
rect 16150 5080 16202 5132
rect 16202 5080 16204 5132
rect 16148 5078 16204 5080
rect 16326 5123 16382 5125
rect 16326 5071 16328 5123
rect 16328 5071 16380 5123
rect 16380 5071 16382 5123
rect 16326 5069 16382 5071
rect 16565 5125 16621 5127
rect 16565 5073 16567 5125
rect 16567 5073 16619 5125
rect 16619 5073 16621 5125
rect 16565 5071 16621 5073
rect 16762 5125 16818 5127
rect 16762 5073 16764 5125
rect 16764 5073 16816 5125
rect 16816 5073 16818 5125
rect 16762 5071 16818 5073
rect 16960 5125 17016 5127
rect 16960 5073 16962 5125
rect 16962 5073 17014 5125
rect 17014 5073 17016 5125
rect 16960 5071 17016 5073
rect 17173 5126 17229 5128
rect 17173 5074 17175 5126
rect 17175 5074 17227 5126
rect 17227 5074 17229 5126
rect 17173 5072 17229 5074
rect 17396 5125 17452 5127
rect 17396 5073 17398 5125
rect 17398 5073 17450 5125
rect 17450 5073 17452 5125
rect 17396 5071 17452 5073
rect 17593 5130 17649 5132
rect 17593 5078 17595 5130
rect 17595 5078 17647 5130
rect 17647 5078 17649 5130
rect 17593 5076 17649 5078
rect 17809 5128 17865 5130
rect 17809 5076 17811 5128
rect 17811 5076 17863 5128
rect 17863 5076 17865 5128
rect 17809 5074 17865 5076
rect 18018 5128 18074 5130
rect 18018 5076 18020 5128
rect 18020 5076 18072 5128
rect 18072 5076 18074 5128
rect 18018 5074 18074 5076
<< metal3 >>
rect 18546 9699 18672 9709
rect 18546 9635 18577 9699
rect 18641 9635 18672 9699
rect 18546 9625 18672 9635
rect 18746 9699 18872 9709
rect 18746 9635 18777 9699
rect 18841 9635 18872 9699
rect 18746 9625 18872 9635
rect 18358 9057 18483 9067
rect 18358 8993 18388 9057
rect 18452 8993 18483 9057
rect 18358 8983 18483 8993
rect 13478 7595 13592 7608
rect 13478 7531 13501 7595
rect 13565 7531 13592 7595
rect 13478 7521 13592 7531
rect 13652 7594 13766 7607
rect 13652 7530 13675 7594
rect 13739 7530 13766 7594
rect 13652 7520 13766 7530
rect 13877 7596 13991 7609
rect 13877 7532 13900 7596
rect 13964 7532 13991 7596
rect 13877 7522 13991 7532
rect 14078 7598 14192 7611
rect 14078 7534 14101 7598
rect 14165 7534 14192 7598
rect 14078 7524 14192 7534
rect 14301 7596 14415 7609
rect 14301 7532 14324 7596
rect 14388 7532 14415 7596
rect 14301 7522 14415 7532
rect 14510 7601 14624 7614
rect 14510 7537 14533 7601
rect 14597 7537 14624 7601
rect 14510 7527 14624 7537
rect 14738 7594 14852 7607
rect 14738 7530 14761 7594
rect 14825 7530 14852 7594
rect 14738 7520 14852 7530
rect 14928 7598 15042 7611
rect 14928 7534 14951 7598
rect 15015 7534 15042 7598
rect 14928 7524 15042 7534
rect 15133 7601 15247 7614
rect 15133 7537 15156 7601
rect 15220 7537 15247 7601
rect 15133 7527 15247 7537
rect 15332 7601 15446 7614
rect 15332 7537 15355 7601
rect 15419 7537 15446 7601
rect 15332 7527 15446 7537
rect 15548 7596 15662 7609
rect 15548 7532 15571 7596
rect 15635 7532 15662 7596
rect 15548 7522 15662 7532
rect 15936 7601 16050 7614
rect 15936 7537 15959 7601
rect 16023 7537 16050 7601
rect 15936 7527 16050 7537
rect 16171 7596 16285 7609
rect 16171 7532 16194 7596
rect 16258 7532 16285 7596
rect 16171 7522 16285 7532
rect 16413 7598 16527 7611
rect 16413 7534 16436 7598
rect 16500 7534 16527 7598
rect 16413 7524 16527 7534
rect 16645 7599 16759 7612
rect 16645 7535 16668 7599
rect 16732 7535 16759 7599
rect 16645 7525 16759 7535
rect 16874 7602 16988 7615
rect 16874 7538 16897 7602
rect 16961 7538 16988 7602
rect 16874 7528 16988 7538
rect 17123 7594 17237 7607
rect 17123 7530 17146 7594
rect 17210 7530 17237 7594
rect 17123 7520 17237 7530
rect 17341 7598 17455 7611
rect 17341 7534 17364 7598
rect 17428 7534 17455 7598
rect 17341 7524 17455 7534
rect 17570 7594 17684 7607
rect 17570 7530 17593 7594
rect 17657 7530 17684 7594
rect 17570 7520 17684 7530
rect 17791 7596 17905 7609
rect 17791 7532 17814 7596
rect 17878 7532 17905 7596
rect 17791 7522 17905 7532
rect 18007 7601 18121 7614
rect 18007 7537 18030 7601
rect 18094 7537 18121 7601
rect 18007 7527 18121 7537
rect 14836 7408 14950 7421
rect 14836 7344 14859 7408
rect 14923 7344 14950 7408
rect 17231 7407 17345 7420
rect 14836 7334 14950 7344
rect 15221 7357 15335 7370
rect 15221 7293 15244 7357
rect 15308 7293 15335 7357
rect 17231 7343 17254 7407
rect 17318 7343 17345 7407
rect 17231 7333 17345 7343
rect 17616 7358 17730 7371
rect 15221 7283 15335 7293
rect 17616 7294 17639 7358
rect 17703 7294 17730 7358
rect 17616 7284 17730 7294
rect 13480 7012 13594 7025
rect 13480 6948 13503 7012
rect 13567 6948 13594 7012
rect 13480 6938 13594 6948
rect 13655 7010 13769 7023
rect 13655 6946 13678 7010
rect 13742 6946 13769 7010
rect 13655 6936 13769 6946
rect 13852 7012 13966 7025
rect 13852 6948 13875 7012
rect 13939 6948 13966 7012
rect 13852 6938 13966 6948
rect 14071 7015 14185 7028
rect 14071 6951 14094 7015
rect 14158 6951 14185 7015
rect 14071 6941 14185 6951
rect 14303 7011 14417 7024
rect 14303 6947 14326 7011
rect 14390 6947 14417 7011
rect 14303 6937 14417 6947
rect 14527 7018 14641 7031
rect 14527 6954 14550 7018
rect 14614 6954 14641 7018
rect 14527 6944 14641 6954
rect 14739 7006 14853 7019
rect 14739 6942 14762 7006
rect 14826 6942 14853 7006
rect 14739 6932 14853 6942
rect 14961 7002 15075 7015
rect 14961 6938 14984 7002
rect 15048 6938 15075 7002
rect 14961 6928 15075 6938
rect 15184 6999 15298 7012
rect 15184 6935 15207 6999
rect 15271 6935 15298 6999
rect 15184 6925 15298 6935
rect 15394 6999 15508 7012
rect 15394 6935 15417 6999
rect 15481 6935 15508 6999
rect 15394 6925 15508 6935
rect 15607 6999 15721 7012
rect 15607 6935 15630 6999
rect 15694 6935 15721 6999
rect 15607 6925 15721 6935
rect 15924 6992 16038 7005
rect 15924 6928 15947 6992
rect 16011 6928 16038 6992
rect 15924 6918 16038 6928
rect 16126 6995 16240 7008
rect 16126 6931 16149 6995
rect 16213 6931 16240 6995
rect 16126 6921 16240 6931
rect 16327 6996 16441 7009
rect 16327 6932 16350 6996
rect 16414 6932 16441 6996
rect 16327 6922 16441 6932
rect 16506 6997 16620 7010
rect 16506 6933 16529 6997
rect 16593 6933 16620 6997
rect 16506 6923 16620 6933
rect 16698 7001 16812 7014
rect 16698 6937 16721 7001
rect 16785 6937 16812 7001
rect 16698 6927 16812 6937
rect 16883 6998 16997 7011
rect 16883 6934 16906 6998
rect 16970 6934 16997 6998
rect 16883 6924 16997 6934
rect 17115 6997 17229 7010
rect 17115 6933 17138 6997
rect 17202 6933 17229 6997
rect 17115 6923 17229 6933
rect 17320 6999 17434 7012
rect 17320 6935 17343 6999
rect 17407 6935 17434 6999
rect 17320 6925 17434 6935
rect 17526 7001 17640 7014
rect 17526 6937 17549 7001
rect 17613 6937 17640 7001
rect 17526 6927 17640 6937
rect 17734 7008 17848 7021
rect 17734 6944 17757 7008
rect 17821 6944 17848 7008
rect 17734 6934 17848 6944
rect 17956 7009 18070 7022
rect 17956 6945 17979 7009
rect 18043 6945 18070 7009
rect 17956 6935 18070 6945
rect 13507 6363 13621 6376
rect 13507 6299 13530 6363
rect 13594 6299 13621 6363
rect 13507 6289 13621 6299
rect 13723 6368 13837 6381
rect 13723 6304 13746 6368
rect 13810 6304 13837 6368
rect 13723 6294 13837 6304
rect 13929 6369 14043 6382
rect 13929 6305 13952 6369
rect 14016 6305 14043 6369
rect 13929 6295 14043 6305
rect 14131 6361 14245 6374
rect 14131 6297 14154 6361
rect 14218 6297 14245 6361
rect 14131 6287 14245 6297
rect 14327 6363 14441 6376
rect 14327 6299 14350 6363
rect 14414 6299 14441 6363
rect 14327 6289 14441 6299
rect 14552 6365 14666 6378
rect 14552 6301 14575 6365
rect 14639 6301 14666 6365
rect 14552 6291 14666 6301
rect 14767 6361 14881 6374
rect 14767 6297 14790 6361
rect 14854 6297 14881 6361
rect 14767 6287 14881 6297
rect 15002 6361 15116 6374
rect 15002 6297 15025 6361
rect 15089 6297 15116 6361
rect 15002 6287 15116 6297
rect 15210 6364 15324 6377
rect 15210 6300 15233 6364
rect 15297 6300 15324 6364
rect 15210 6290 15324 6300
rect 15452 6364 15566 6377
rect 15452 6300 15475 6364
rect 15539 6300 15566 6364
rect 15452 6290 15566 6300
rect 15650 6365 15764 6378
rect 15650 6301 15673 6365
rect 15737 6301 15764 6365
rect 15650 6291 15764 6301
rect 15957 6365 16071 6378
rect 15957 6301 15980 6365
rect 16044 6301 16071 6365
rect 15957 6291 16071 6301
rect 16182 6366 16296 6379
rect 16182 6302 16205 6366
rect 16269 6302 16296 6366
rect 16182 6292 16296 6302
rect 16411 6365 16525 6378
rect 16411 6301 16434 6365
rect 16498 6301 16525 6365
rect 16411 6291 16525 6301
rect 16627 6369 16741 6382
rect 16627 6305 16650 6369
rect 16714 6305 16741 6369
rect 16627 6295 16741 6305
rect 16850 6372 16964 6385
rect 16850 6308 16873 6372
rect 16937 6308 16964 6372
rect 16850 6298 16964 6308
rect 17074 6368 17188 6381
rect 17074 6304 17097 6368
rect 17161 6304 17188 6368
rect 17074 6294 17188 6304
rect 17301 6357 17415 6370
rect 17301 6293 17324 6357
rect 17388 6293 17415 6357
rect 17301 6283 17415 6293
rect 17514 6356 17628 6369
rect 17514 6292 17537 6356
rect 17601 6292 17628 6356
rect 17514 6282 17628 6292
rect 17725 6360 17839 6373
rect 17725 6296 17748 6360
rect 17812 6296 17839 6360
rect 17725 6286 17839 6296
rect 17952 6361 18066 6374
rect 17952 6297 17975 6361
rect 18039 6297 18066 6361
rect 17952 6287 18066 6297
rect 14841 6134 14955 6147
rect 14841 6070 14864 6134
rect 14928 6070 14955 6134
rect 17233 6136 17347 6149
rect 14841 6060 14955 6070
rect 15224 6075 15338 6088
rect 15224 6011 15247 6075
rect 15311 6011 15338 6075
rect 17233 6072 17256 6136
rect 17320 6072 17347 6136
rect 17233 6062 17347 6072
rect 17610 6082 17724 6095
rect 15224 6001 15338 6011
rect 17610 6018 17633 6082
rect 17697 6018 17724 6082
rect 17610 6008 17724 6018
rect 13533 5718 13647 5731
rect 13533 5654 13556 5718
rect 13620 5654 13647 5718
rect 13533 5644 13647 5654
rect 13758 5727 13872 5740
rect 13758 5663 13781 5727
rect 13845 5663 13872 5727
rect 13758 5653 13872 5663
rect 14035 5724 14149 5737
rect 14035 5660 14058 5724
rect 14122 5660 14149 5724
rect 14035 5650 14149 5660
rect 14256 5727 14370 5740
rect 14256 5663 14279 5727
rect 14343 5663 14370 5727
rect 14256 5653 14370 5663
rect 14501 5724 14615 5737
rect 14501 5660 14524 5724
rect 14588 5660 14615 5724
rect 14501 5650 14615 5660
rect 14727 5728 14841 5741
rect 14727 5664 14750 5728
rect 14814 5664 14841 5728
rect 14727 5654 14841 5664
rect 14939 5726 15053 5739
rect 14939 5662 14962 5726
rect 15026 5662 15053 5726
rect 14939 5652 15053 5662
rect 15159 5732 15273 5745
rect 15159 5668 15182 5732
rect 15246 5668 15273 5732
rect 15159 5658 15273 5668
rect 15397 5734 15511 5747
rect 15397 5670 15420 5734
rect 15484 5670 15511 5734
rect 15397 5660 15511 5670
rect 15610 5736 15724 5749
rect 15610 5672 15633 5736
rect 15697 5672 15724 5736
rect 15610 5662 15724 5672
rect 15997 5726 16111 5739
rect 15997 5662 16020 5726
rect 16084 5662 16111 5726
rect 15997 5652 16111 5662
rect 16344 5727 16458 5740
rect 16344 5663 16367 5727
rect 16431 5663 16458 5727
rect 16344 5653 16458 5663
rect 16580 5722 16694 5735
rect 16580 5658 16603 5722
rect 16667 5658 16694 5722
rect 16580 5648 16694 5658
rect 16764 5722 16878 5735
rect 16764 5658 16787 5722
rect 16851 5658 16878 5722
rect 16764 5648 16878 5658
rect 17003 5724 17117 5737
rect 17003 5660 17026 5724
rect 17090 5660 17117 5724
rect 17003 5650 17117 5660
rect 17206 5720 17320 5733
rect 17206 5656 17229 5720
rect 17293 5656 17320 5720
rect 17206 5646 17320 5656
rect 17391 5717 17505 5730
rect 17391 5653 17414 5717
rect 17478 5653 17505 5717
rect 17391 5643 17505 5653
rect 17582 5719 17696 5732
rect 17582 5655 17605 5719
rect 17669 5655 17696 5719
rect 17582 5645 17696 5655
rect 17773 5723 17887 5736
rect 17773 5659 17796 5723
rect 17860 5659 17887 5723
rect 17773 5649 17887 5659
rect 17959 5719 18073 5732
rect 17959 5655 17982 5719
rect 18046 5655 18073 5719
rect 17959 5645 18073 5655
rect 13406 5136 13520 5149
rect 13406 5072 13429 5136
rect 13493 5072 13520 5136
rect 13406 5062 13520 5072
rect 13611 5132 13725 5145
rect 13611 5068 13634 5132
rect 13698 5068 13725 5132
rect 13611 5058 13725 5068
rect 13797 5137 13911 5150
rect 13797 5073 13820 5137
rect 13884 5073 13911 5137
rect 13797 5063 13911 5073
rect 13991 5130 14105 5143
rect 13991 5066 14014 5130
rect 14078 5066 14105 5130
rect 13991 5056 14105 5066
rect 14210 5135 14324 5148
rect 14210 5071 14233 5135
rect 14297 5071 14324 5135
rect 14210 5061 14324 5071
rect 14420 5135 14534 5148
rect 14420 5071 14443 5135
rect 14507 5071 14534 5135
rect 14420 5061 14534 5071
rect 14649 5132 14763 5145
rect 14649 5068 14672 5132
rect 14736 5068 14763 5132
rect 14649 5058 14763 5068
rect 14895 5132 15009 5145
rect 14895 5068 14918 5132
rect 14982 5068 15009 5132
rect 14895 5058 15009 5068
rect 15169 5132 15283 5145
rect 15169 5068 15192 5132
rect 15256 5068 15283 5132
rect 15169 5058 15283 5068
rect 15444 5132 15558 5145
rect 15444 5068 15467 5132
rect 15531 5068 15558 5132
rect 15444 5058 15558 5068
rect 15680 5132 15794 5145
rect 15680 5068 15703 5132
rect 15767 5068 15794 5132
rect 15680 5058 15794 5068
rect 15903 5135 16017 5148
rect 15903 5071 15926 5135
rect 15990 5071 16017 5135
rect 15903 5061 16017 5071
rect 16121 5138 16235 5151
rect 16121 5074 16144 5138
rect 16208 5074 16235 5138
rect 16121 5064 16235 5074
rect 16299 5129 16413 5142
rect 16299 5065 16322 5129
rect 16386 5065 16413 5129
rect 16299 5055 16413 5065
rect 16538 5131 16652 5144
rect 16538 5067 16561 5131
rect 16625 5067 16652 5131
rect 16538 5057 16652 5067
rect 16735 5131 16849 5144
rect 16735 5067 16758 5131
rect 16822 5067 16849 5131
rect 16735 5057 16849 5067
rect 16933 5131 17047 5144
rect 16933 5067 16956 5131
rect 17020 5067 17047 5131
rect 16933 5057 17047 5067
rect 17146 5132 17260 5145
rect 17146 5068 17169 5132
rect 17233 5068 17260 5132
rect 17146 5058 17260 5068
rect 17369 5131 17483 5144
rect 17369 5067 17392 5131
rect 17456 5067 17483 5131
rect 17369 5057 17483 5067
rect 17566 5136 17680 5149
rect 17566 5072 17589 5136
rect 17653 5072 17680 5136
rect 17566 5062 17680 5072
rect 17782 5134 17896 5147
rect 17782 5070 17805 5134
rect 17869 5070 17896 5134
rect 17782 5060 17896 5070
rect 17991 5134 18105 5147
rect 17991 5070 18014 5134
rect 18078 5070 18105 5134
rect 17991 5060 18105 5070
<< via3 >>
rect 18577 9695 18641 9699
rect 18577 9639 18581 9695
rect 18581 9639 18637 9695
rect 18637 9639 18641 9695
rect 18577 9635 18641 9639
rect 18777 9695 18841 9699
rect 18777 9639 18781 9695
rect 18781 9639 18837 9695
rect 18837 9639 18841 9695
rect 18777 9635 18841 9639
rect 18388 9053 18452 9057
rect 18388 8997 18392 9053
rect 18392 8997 18448 9053
rect 18448 8997 18452 9053
rect 18388 8993 18452 8997
rect 13501 7591 13565 7595
rect 13501 7535 13505 7591
rect 13505 7535 13561 7591
rect 13561 7535 13565 7591
rect 13501 7531 13565 7535
rect 13675 7590 13739 7594
rect 13675 7534 13679 7590
rect 13679 7534 13735 7590
rect 13735 7534 13739 7590
rect 13675 7530 13739 7534
rect 13900 7592 13964 7596
rect 13900 7536 13904 7592
rect 13904 7536 13960 7592
rect 13960 7536 13964 7592
rect 13900 7532 13964 7536
rect 14101 7594 14165 7598
rect 14101 7538 14105 7594
rect 14105 7538 14161 7594
rect 14161 7538 14165 7594
rect 14101 7534 14165 7538
rect 14324 7592 14388 7596
rect 14324 7536 14328 7592
rect 14328 7536 14384 7592
rect 14384 7536 14388 7592
rect 14324 7532 14388 7536
rect 14533 7597 14597 7601
rect 14533 7541 14537 7597
rect 14537 7541 14593 7597
rect 14593 7541 14597 7597
rect 14533 7537 14597 7541
rect 14761 7590 14825 7594
rect 14761 7534 14765 7590
rect 14765 7534 14821 7590
rect 14821 7534 14825 7590
rect 14761 7530 14825 7534
rect 14951 7594 15015 7598
rect 14951 7538 14955 7594
rect 14955 7538 15011 7594
rect 15011 7538 15015 7594
rect 14951 7534 15015 7538
rect 15156 7597 15220 7601
rect 15156 7541 15160 7597
rect 15160 7541 15216 7597
rect 15216 7541 15220 7597
rect 15156 7537 15220 7541
rect 15355 7597 15419 7601
rect 15355 7541 15359 7597
rect 15359 7541 15415 7597
rect 15415 7541 15419 7597
rect 15355 7537 15419 7541
rect 15571 7592 15635 7596
rect 15571 7536 15575 7592
rect 15575 7536 15631 7592
rect 15631 7536 15635 7592
rect 15571 7532 15635 7536
rect 15959 7597 16023 7601
rect 15959 7541 15963 7597
rect 15963 7541 16019 7597
rect 16019 7541 16023 7597
rect 15959 7537 16023 7541
rect 16194 7592 16258 7596
rect 16194 7536 16198 7592
rect 16198 7536 16254 7592
rect 16254 7536 16258 7592
rect 16194 7532 16258 7536
rect 16436 7594 16500 7598
rect 16436 7538 16440 7594
rect 16440 7538 16496 7594
rect 16496 7538 16500 7594
rect 16436 7534 16500 7538
rect 16668 7595 16732 7599
rect 16668 7539 16672 7595
rect 16672 7539 16728 7595
rect 16728 7539 16732 7595
rect 16668 7535 16732 7539
rect 16897 7598 16961 7602
rect 16897 7542 16901 7598
rect 16901 7542 16957 7598
rect 16957 7542 16961 7598
rect 16897 7538 16961 7542
rect 17146 7590 17210 7594
rect 17146 7534 17150 7590
rect 17150 7534 17206 7590
rect 17206 7534 17210 7590
rect 17146 7530 17210 7534
rect 17364 7594 17428 7598
rect 17364 7538 17368 7594
rect 17368 7538 17424 7594
rect 17424 7538 17428 7594
rect 17364 7534 17428 7538
rect 17593 7590 17657 7594
rect 17593 7534 17597 7590
rect 17597 7534 17653 7590
rect 17653 7534 17657 7590
rect 17593 7530 17657 7534
rect 17814 7592 17878 7596
rect 17814 7536 17818 7592
rect 17818 7536 17874 7592
rect 17874 7536 17878 7592
rect 17814 7532 17878 7536
rect 18030 7597 18094 7601
rect 18030 7541 18034 7597
rect 18034 7541 18090 7597
rect 18090 7541 18094 7597
rect 18030 7537 18094 7541
rect 14859 7404 14923 7408
rect 14859 7348 14863 7404
rect 14863 7348 14919 7404
rect 14919 7348 14923 7404
rect 14859 7344 14923 7348
rect 15244 7353 15308 7357
rect 15244 7297 15248 7353
rect 15248 7297 15304 7353
rect 15304 7297 15308 7353
rect 15244 7293 15308 7297
rect 17254 7403 17318 7407
rect 17254 7347 17258 7403
rect 17258 7347 17314 7403
rect 17314 7347 17318 7403
rect 17254 7343 17318 7347
rect 17639 7354 17703 7358
rect 17639 7298 17643 7354
rect 17643 7298 17699 7354
rect 17699 7298 17703 7354
rect 17639 7294 17703 7298
rect 13503 7008 13567 7012
rect 13503 6952 13507 7008
rect 13507 6952 13563 7008
rect 13563 6952 13567 7008
rect 13503 6948 13567 6952
rect 13678 7006 13742 7010
rect 13678 6950 13682 7006
rect 13682 6950 13738 7006
rect 13738 6950 13742 7006
rect 13678 6946 13742 6950
rect 13875 7008 13939 7012
rect 13875 6952 13879 7008
rect 13879 6952 13935 7008
rect 13935 6952 13939 7008
rect 13875 6948 13939 6952
rect 14094 7011 14158 7015
rect 14094 6955 14098 7011
rect 14098 6955 14154 7011
rect 14154 6955 14158 7011
rect 14094 6951 14158 6955
rect 14326 7007 14390 7011
rect 14326 6951 14330 7007
rect 14330 6951 14386 7007
rect 14386 6951 14390 7007
rect 14326 6947 14390 6951
rect 14550 7014 14614 7018
rect 14550 6958 14554 7014
rect 14554 6958 14610 7014
rect 14610 6958 14614 7014
rect 14550 6954 14614 6958
rect 14762 7002 14826 7006
rect 14762 6946 14766 7002
rect 14766 6946 14822 7002
rect 14822 6946 14826 7002
rect 14762 6942 14826 6946
rect 14984 6998 15048 7002
rect 14984 6942 14988 6998
rect 14988 6942 15044 6998
rect 15044 6942 15048 6998
rect 14984 6938 15048 6942
rect 15207 6995 15271 6999
rect 15207 6939 15211 6995
rect 15211 6939 15267 6995
rect 15267 6939 15271 6995
rect 15207 6935 15271 6939
rect 15417 6995 15481 6999
rect 15417 6939 15421 6995
rect 15421 6939 15477 6995
rect 15477 6939 15481 6995
rect 15417 6935 15481 6939
rect 15630 6995 15694 6999
rect 15630 6939 15634 6995
rect 15634 6939 15690 6995
rect 15690 6939 15694 6995
rect 15630 6935 15694 6939
rect 15947 6988 16011 6992
rect 15947 6932 15951 6988
rect 15951 6932 16007 6988
rect 16007 6932 16011 6988
rect 15947 6928 16011 6932
rect 16149 6991 16213 6995
rect 16149 6935 16153 6991
rect 16153 6935 16209 6991
rect 16209 6935 16213 6991
rect 16149 6931 16213 6935
rect 16350 6992 16414 6996
rect 16350 6936 16354 6992
rect 16354 6936 16410 6992
rect 16410 6936 16414 6992
rect 16350 6932 16414 6936
rect 16529 6993 16593 6997
rect 16529 6937 16533 6993
rect 16533 6937 16589 6993
rect 16589 6937 16593 6993
rect 16529 6933 16593 6937
rect 16721 6997 16785 7001
rect 16721 6941 16725 6997
rect 16725 6941 16781 6997
rect 16781 6941 16785 6997
rect 16721 6937 16785 6941
rect 16906 6994 16970 6998
rect 16906 6938 16910 6994
rect 16910 6938 16966 6994
rect 16966 6938 16970 6994
rect 16906 6934 16970 6938
rect 17138 6993 17202 6997
rect 17138 6937 17142 6993
rect 17142 6937 17198 6993
rect 17198 6937 17202 6993
rect 17138 6933 17202 6937
rect 17343 6995 17407 6999
rect 17343 6939 17347 6995
rect 17347 6939 17403 6995
rect 17403 6939 17407 6995
rect 17343 6935 17407 6939
rect 17549 6997 17613 7001
rect 17549 6941 17553 6997
rect 17553 6941 17609 6997
rect 17609 6941 17613 6997
rect 17549 6937 17613 6941
rect 17757 7004 17821 7008
rect 17757 6948 17761 7004
rect 17761 6948 17817 7004
rect 17817 6948 17821 7004
rect 17757 6944 17821 6948
rect 17979 7005 18043 7009
rect 17979 6949 17983 7005
rect 17983 6949 18039 7005
rect 18039 6949 18043 7005
rect 17979 6945 18043 6949
rect 13530 6359 13594 6363
rect 13530 6303 13534 6359
rect 13534 6303 13590 6359
rect 13590 6303 13594 6359
rect 13530 6299 13594 6303
rect 13746 6364 13810 6368
rect 13746 6308 13750 6364
rect 13750 6308 13806 6364
rect 13806 6308 13810 6364
rect 13746 6304 13810 6308
rect 13952 6365 14016 6369
rect 13952 6309 13956 6365
rect 13956 6309 14012 6365
rect 14012 6309 14016 6365
rect 13952 6305 14016 6309
rect 14154 6357 14218 6361
rect 14154 6301 14158 6357
rect 14158 6301 14214 6357
rect 14214 6301 14218 6357
rect 14154 6297 14218 6301
rect 14350 6359 14414 6363
rect 14350 6303 14354 6359
rect 14354 6303 14410 6359
rect 14410 6303 14414 6359
rect 14350 6299 14414 6303
rect 14575 6361 14639 6365
rect 14575 6305 14579 6361
rect 14579 6305 14635 6361
rect 14635 6305 14639 6361
rect 14575 6301 14639 6305
rect 14790 6357 14854 6361
rect 14790 6301 14794 6357
rect 14794 6301 14850 6357
rect 14850 6301 14854 6357
rect 14790 6297 14854 6301
rect 15025 6357 15089 6361
rect 15025 6301 15029 6357
rect 15029 6301 15085 6357
rect 15085 6301 15089 6357
rect 15025 6297 15089 6301
rect 15233 6360 15297 6364
rect 15233 6304 15237 6360
rect 15237 6304 15293 6360
rect 15293 6304 15297 6360
rect 15233 6300 15297 6304
rect 15475 6360 15539 6364
rect 15475 6304 15479 6360
rect 15479 6304 15535 6360
rect 15535 6304 15539 6360
rect 15475 6300 15539 6304
rect 15673 6361 15737 6365
rect 15673 6305 15677 6361
rect 15677 6305 15733 6361
rect 15733 6305 15737 6361
rect 15673 6301 15737 6305
rect 15980 6361 16044 6365
rect 15980 6305 15984 6361
rect 15984 6305 16040 6361
rect 16040 6305 16044 6361
rect 15980 6301 16044 6305
rect 16205 6362 16269 6366
rect 16205 6306 16209 6362
rect 16209 6306 16265 6362
rect 16265 6306 16269 6362
rect 16205 6302 16269 6306
rect 16434 6361 16498 6365
rect 16434 6305 16438 6361
rect 16438 6305 16494 6361
rect 16494 6305 16498 6361
rect 16434 6301 16498 6305
rect 16650 6365 16714 6369
rect 16650 6309 16654 6365
rect 16654 6309 16710 6365
rect 16710 6309 16714 6365
rect 16650 6305 16714 6309
rect 16873 6368 16937 6372
rect 16873 6312 16877 6368
rect 16877 6312 16933 6368
rect 16933 6312 16937 6368
rect 16873 6308 16937 6312
rect 17097 6364 17161 6368
rect 17097 6308 17101 6364
rect 17101 6308 17157 6364
rect 17157 6308 17161 6364
rect 17097 6304 17161 6308
rect 17324 6353 17388 6357
rect 17324 6297 17328 6353
rect 17328 6297 17384 6353
rect 17384 6297 17388 6353
rect 17324 6293 17388 6297
rect 17537 6352 17601 6356
rect 17537 6296 17541 6352
rect 17541 6296 17597 6352
rect 17597 6296 17601 6352
rect 17537 6292 17601 6296
rect 17748 6356 17812 6360
rect 17748 6300 17752 6356
rect 17752 6300 17808 6356
rect 17808 6300 17812 6356
rect 17748 6296 17812 6300
rect 17975 6357 18039 6361
rect 17975 6301 17979 6357
rect 17979 6301 18035 6357
rect 18035 6301 18039 6357
rect 17975 6297 18039 6301
rect 14864 6130 14928 6134
rect 14864 6074 14868 6130
rect 14868 6074 14924 6130
rect 14924 6074 14928 6130
rect 14864 6070 14928 6074
rect 15247 6071 15311 6075
rect 15247 6015 15251 6071
rect 15251 6015 15307 6071
rect 15307 6015 15311 6071
rect 15247 6011 15311 6015
rect 17256 6132 17320 6136
rect 17256 6076 17260 6132
rect 17260 6076 17316 6132
rect 17316 6076 17320 6132
rect 17256 6072 17320 6076
rect 17633 6078 17697 6082
rect 17633 6022 17637 6078
rect 17637 6022 17693 6078
rect 17693 6022 17697 6078
rect 17633 6018 17697 6022
rect 13556 5714 13620 5718
rect 13556 5658 13560 5714
rect 13560 5658 13616 5714
rect 13616 5658 13620 5714
rect 13556 5654 13620 5658
rect 13781 5723 13845 5727
rect 13781 5667 13785 5723
rect 13785 5667 13841 5723
rect 13841 5667 13845 5723
rect 13781 5663 13845 5667
rect 14058 5720 14122 5724
rect 14058 5664 14062 5720
rect 14062 5664 14118 5720
rect 14118 5664 14122 5720
rect 14058 5660 14122 5664
rect 14279 5723 14343 5727
rect 14279 5667 14283 5723
rect 14283 5667 14339 5723
rect 14339 5667 14343 5723
rect 14279 5663 14343 5667
rect 14524 5720 14588 5724
rect 14524 5664 14528 5720
rect 14528 5664 14584 5720
rect 14584 5664 14588 5720
rect 14524 5660 14588 5664
rect 14750 5724 14814 5728
rect 14750 5668 14754 5724
rect 14754 5668 14810 5724
rect 14810 5668 14814 5724
rect 14750 5664 14814 5668
rect 14962 5722 15026 5726
rect 14962 5666 14966 5722
rect 14966 5666 15022 5722
rect 15022 5666 15026 5722
rect 14962 5662 15026 5666
rect 15182 5728 15246 5732
rect 15182 5672 15186 5728
rect 15186 5672 15242 5728
rect 15242 5672 15246 5728
rect 15182 5668 15246 5672
rect 15420 5730 15484 5734
rect 15420 5674 15424 5730
rect 15424 5674 15480 5730
rect 15480 5674 15484 5730
rect 15420 5670 15484 5674
rect 15633 5732 15697 5736
rect 15633 5676 15637 5732
rect 15637 5676 15693 5732
rect 15693 5676 15697 5732
rect 15633 5672 15697 5676
rect 16020 5722 16084 5726
rect 16020 5666 16024 5722
rect 16024 5666 16080 5722
rect 16080 5666 16084 5722
rect 16020 5662 16084 5666
rect 16367 5723 16431 5727
rect 16367 5667 16371 5723
rect 16371 5667 16427 5723
rect 16427 5667 16431 5723
rect 16367 5663 16431 5667
rect 16603 5718 16667 5722
rect 16603 5662 16607 5718
rect 16607 5662 16663 5718
rect 16663 5662 16667 5718
rect 16603 5658 16667 5662
rect 16787 5718 16851 5722
rect 16787 5662 16791 5718
rect 16791 5662 16847 5718
rect 16847 5662 16851 5718
rect 16787 5658 16851 5662
rect 17026 5720 17090 5724
rect 17026 5664 17030 5720
rect 17030 5664 17086 5720
rect 17086 5664 17090 5720
rect 17026 5660 17090 5664
rect 17229 5716 17293 5720
rect 17229 5660 17233 5716
rect 17233 5660 17289 5716
rect 17289 5660 17293 5716
rect 17229 5656 17293 5660
rect 17414 5713 17478 5717
rect 17414 5657 17418 5713
rect 17418 5657 17474 5713
rect 17474 5657 17478 5713
rect 17414 5653 17478 5657
rect 17605 5715 17669 5719
rect 17605 5659 17609 5715
rect 17609 5659 17665 5715
rect 17665 5659 17669 5715
rect 17605 5655 17669 5659
rect 17796 5719 17860 5723
rect 17796 5663 17800 5719
rect 17800 5663 17856 5719
rect 17856 5663 17860 5719
rect 17796 5659 17860 5663
rect 17982 5715 18046 5719
rect 17982 5659 17986 5715
rect 17986 5659 18042 5715
rect 18042 5659 18046 5715
rect 17982 5655 18046 5659
rect 13429 5132 13493 5136
rect 13429 5076 13433 5132
rect 13433 5076 13489 5132
rect 13489 5076 13493 5132
rect 13429 5072 13493 5076
rect 13634 5128 13698 5132
rect 13634 5072 13638 5128
rect 13638 5072 13694 5128
rect 13694 5072 13698 5128
rect 13634 5068 13698 5072
rect 13820 5133 13884 5137
rect 13820 5077 13824 5133
rect 13824 5077 13880 5133
rect 13880 5077 13884 5133
rect 13820 5073 13884 5077
rect 14014 5126 14078 5130
rect 14014 5070 14018 5126
rect 14018 5070 14074 5126
rect 14074 5070 14078 5126
rect 14014 5066 14078 5070
rect 14233 5131 14297 5135
rect 14233 5075 14237 5131
rect 14237 5075 14293 5131
rect 14293 5075 14297 5131
rect 14233 5071 14297 5075
rect 14443 5131 14507 5135
rect 14443 5075 14447 5131
rect 14447 5075 14503 5131
rect 14503 5075 14507 5131
rect 14443 5071 14507 5075
rect 14672 5128 14736 5132
rect 14672 5072 14676 5128
rect 14676 5072 14732 5128
rect 14732 5072 14736 5128
rect 14672 5068 14736 5072
rect 14918 5128 14982 5132
rect 14918 5072 14922 5128
rect 14922 5072 14978 5128
rect 14978 5072 14982 5128
rect 14918 5068 14982 5072
rect 15192 5128 15256 5132
rect 15192 5072 15196 5128
rect 15196 5072 15252 5128
rect 15252 5072 15256 5128
rect 15192 5068 15256 5072
rect 15467 5128 15531 5132
rect 15467 5072 15471 5128
rect 15471 5072 15527 5128
rect 15527 5072 15531 5128
rect 15467 5068 15531 5072
rect 15703 5128 15767 5132
rect 15703 5072 15707 5128
rect 15707 5072 15763 5128
rect 15763 5072 15767 5128
rect 15703 5068 15767 5072
rect 15926 5131 15990 5135
rect 15926 5075 15930 5131
rect 15930 5075 15986 5131
rect 15986 5075 15990 5131
rect 15926 5071 15990 5075
rect 16144 5134 16208 5138
rect 16144 5078 16148 5134
rect 16148 5078 16204 5134
rect 16204 5078 16208 5134
rect 16144 5074 16208 5078
rect 16322 5125 16386 5129
rect 16322 5069 16326 5125
rect 16326 5069 16382 5125
rect 16382 5069 16386 5125
rect 16322 5065 16386 5069
rect 16561 5127 16625 5131
rect 16561 5071 16565 5127
rect 16565 5071 16621 5127
rect 16621 5071 16625 5127
rect 16561 5067 16625 5071
rect 16758 5127 16822 5131
rect 16758 5071 16762 5127
rect 16762 5071 16818 5127
rect 16818 5071 16822 5127
rect 16758 5067 16822 5071
rect 16956 5127 17020 5131
rect 16956 5071 16960 5127
rect 16960 5071 17016 5127
rect 17016 5071 17020 5127
rect 16956 5067 17020 5071
rect 17169 5128 17233 5132
rect 17169 5072 17173 5128
rect 17173 5072 17229 5128
rect 17229 5072 17233 5128
rect 17169 5068 17233 5072
rect 17392 5127 17456 5131
rect 17392 5071 17396 5127
rect 17396 5071 17452 5127
rect 17452 5071 17456 5127
rect 17392 5067 17456 5071
rect 17589 5132 17653 5136
rect 17589 5076 17593 5132
rect 17593 5076 17649 5132
rect 17649 5076 17653 5132
rect 17589 5072 17653 5076
rect 17805 5130 17869 5134
rect 17805 5074 17809 5130
rect 17809 5074 17865 5130
rect 17865 5074 17869 5130
rect 17805 5070 17869 5074
rect 18014 5130 18078 5134
rect 18014 5074 18018 5130
rect 18018 5074 18074 5130
rect 18074 5074 18078 5130
rect 18014 5070 18078 5074
<< metal4 >>
rect 11836 10013 12254 10623
rect 18267 10492 19041 10623
rect 18267 10217 18493 10492
rect 18590 10217 19041 10492
rect 18267 9699 19041 10217
rect 18267 9636 18577 9699
rect 18545 9635 18577 9636
rect 18641 9635 18777 9699
rect 18841 9635 19041 9699
rect 11864 7966 12240 9403
rect 18197 9057 18483 9093
rect 18197 8993 18388 9057
rect 18452 8993 18483 9057
rect 18197 8890 18483 8993
rect 11864 7602 18154 7966
rect 11864 7601 16897 7602
rect 11864 7598 14533 7601
rect 11864 7596 14101 7598
rect 11864 7595 13900 7596
rect 11864 7531 13501 7595
rect 13565 7594 13900 7595
rect 13565 7531 13675 7594
rect 11864 7530 13675 7531
rect 13739 7532 13900 7594
rect 13964 7534 14101 7596
rect 14165 7596 14533 7598
rect 14165 7534 14324 7596
rect 13964 7532 14324 7534
rect 14388 7537 14533 7596
rect 14597 7598 15156 7601
rect 14597 7594 14951 7598
rect 14597 7537 14761 7594
rect 14388 7532 14761 7537
rect 13739 7530 14761 7532
rect 14825 7534 14951 7594
rect 15015 7537 15156 7598
rect 15220 7537 15355 7601
rect 15419 7596 15959 7601
rect 15419 7537 15571 7596
rect 15015 7534 15571 7537
rect 14825 7532 15571 7534
rect 15635 7537 15959 7596
rect 16023 7599 16897 7601
rect 16023 7598 16668 7599
rect 16023 7596 16436 7598
rect 16023 7537 16194 7596
rect 15635 7532 16194 7537
rect 16258 7534 16436 7596
rect 16500 7535 16668 7598
rect 16732 7538 16897 7599
rect 16961 7601 18154 7602
rect 16961 7598 18030 7601
rect 16961 7594 17364 7598
rect 16961 7538 17146 7594
rect 16732 7535 17146 7538
rect 16500 7534 17146 7535
rect 16258 7532 17146 7534
rect 14825 7530 17146 7532
rect 17210 7534 17364 7594
rect 17428 7596 18030 7598
rect 17428 7594 17814 7596
rect 17428 7534 17593 7594
rect 17210 7530 17593 7534
rect 17657 7532 17814 7594
rect 17878 7537 18030 7596
rect 18094 7537 18154 7601
rect 17878 7532 18154 7537
rect 17657 7530 18154 7532
rect 11864 7481 18154 7530
rect 12771 6704 13267 7481
rect 14836 7408 14950 7421
rect 14836 7351 14859 7408
rect 13330 7344 14859 7351
rect 14923 7351 14950 7408
rect 17231 7407 17345 7420
rect 15221 7357 15335 7370
rect 15221 7351 15244 7357
rect 14923 7344 15244 7351
rect 13330 7293 15244 7344
rect 15308 7351 15335 7357
rect 17231 7351 17254 7407
rect 15308 7343 17254 7351
rect 17318 7351 17345 7407
rect 17616 7358 17730 7371
rect 17616 7351 17639 7358
rect 17318 7343 17639 7351
rect 15308 7294 17639 7343
rect 17703 7351 17730 7358
rect 18545 7351 19041 9635
rect 17703 7294 19043 7351
rect 15308 7293 19043 7294
rect 13330 7146 19043 7293
rect 13330 7018 19042 7146
rect 13330 7015 14550 7018
rect 13330 7012 14094 7015
rect 13330 6948 13503 7012
rect 13567 7010 13875 7012
rect 13567 6948 13678 7010
rect 13330 6946 13678 6948
rect 13742 6948 13875 7010
rect 13939 6951 14094 7012
rect 14158 7011 14550 7015
rect 14158 6951 14326 7011
rect 13939 6948 14326 6951
rect 13742 6947 14326 6948
rect 14390 6954 14550 7011
rect 14614 7009 19042 7018
rect 14614 7008 17979 7009
rect 14614 7006 17757 7008
rect 14614 6954 14762 7006
rect 14390 6947 14762 6954
rect 13742 6946 14762 6947
rect 13330 6942 14762 6946
rect 14826 7002 17757 7006
rect 14826 6942 14984 7002
rect 13330 6938 14984 6942
rect 15048 7001 17757 7002
rect 15048 6999 16721 7001
rect 15048 6938 15207 6999
rect 13330 6935 15207 6938
rect 15271 6935 15417 6999
rect 15481 6935 15630 6999
rect 15694 6997 16721 6999
rect 15694 6996 16529 6997
rect 15694 6995 16350 6996
rect 15694 6992 16149 6995
rect 15694 6935 15947 6992
rect 13330 6928 15947 6935
rect 16011 6931 16149 6992
rect 16213 6932 16350 6995
rect 16414 6933 16529 6996
rect 16593 6937 16721 6997
rect 16785 6999 17549 7001
rect 16785 6998 17343 6999
rect 16785 6937 16906 6998
rect 16593 6934 16906 6937
rect 16970 6997 17343 6998
rect 16970 6934 17138 6997
rect 16593 6933 17138 6934
rect 17202 6935 17343 6997
rect 17407 6937 17549 6999
rect 17613 6944 17757 7001
rect 17821 6945 17979 7008
rect 18043 6945 19042 7009
rect 17821 6944 19042 6945
rect 17613 6937 19042 6944
rect 17407 6935 19042 6937
rect 17202 6933 19042 6935
rect 16414 6932 19042 6933
rect 16213 6931 19042 6932
rect 16011 6928 19042 6931
rect 13330 6866 19042 6928
rect 12771 6372 18193 6704
rect 12771 6369 16873 6372
rect 12771 6368 13952 6369
rect 12771 6363 13746 6368
rect 12771 6299 13530 6363
rect 13594 6304 13746 6363
rect 13810 6305 13952 6368
rect 14016 6366 16650 6369
rect 14016 6365 16205 6366
rect 14016 6363 14575 6365
rect 14016 6361 14350 6363
rect 14016 6305 14154 6361
rect 13810 6304 14154 6305
rect 13594 6299 14154 6304
rect 12771 6297 14154 6299
rect 14218 6299 14350 6361
rect 14414 6301 14575 6363
rect 14639 6364 15673 6365
rect 14639 6361 15233 6364
rect 14639 6301 14790 6361
rect 14414 6299 14790 6301
rect 14218 6297 14790 6299
rect 14854 6297 15025 6361
rect 15089 6300 15233 6361
rect 15297 6300 15475 6364
rect 15539 6301 15673 6364
rect 15737 6301 15980 6365
rect 16044 6302 16205 6365
rect 16269 6365 16650 6366
rect 16269 6302 16434 6365
rect 16044 6301 16434 6302
rect 16498 6305 16650 6365
rect 16714 6308 16873 6369
rect 16937 6368 18193 6372
rect 16937 6308 17097 6368
rect 16714 6305 17097 6308
rect 16498 6304 17097 6305
rect 17161 6361 18193 6368
rect 17161 6360 17975 6361
rect 17161 6357 17748 6360
rect 17161 6304 17324 6357
rect 16498 6301 17324 6304
rect 15539 6300 17324 6301
rect 15089 6297 17324 6300
rect 12771 6293 17324 6297
rect 17388 6356 17748 6357
rect 17388 6293 17537 6356
rect 12771 6292 17537 6293
rect 17601 6296 17748 6356
rect 17812 6297 17975 6360
rect 18039 6297 18193 6361
rect 17812 6296 18193 6297
rect 17601 6292 18193 6296
rect 12771 6219 18193 6292
rect 12771 5525 13267 6219
rect 14841 6134 14955 6147
rect 14841 6076 14864 6134
rect 13327 6070 14864 6076
rect 14928 6076 14955 6134
rect 17233 6136 17347 6149
rect 15224 6076 15338 6088
rect 17233 6076 17256 6136
rect 14928 6075 17256 6076
rect 14928 6070 15247 6075
rect 13327 6011 15247 6070
rect 15311 6072 17256 6075
rect 17320 6076 17347 6136
rect 17610 6082 17724 6095
rect 17610 6076 17633 6082
rect 17320 6072 17633 6076
rect 15311 6018 17633 6072
rect 17697 6076 17724 6082
rect 18545 6076 19041 6866
rect 17697 6018 19043 6076
rect 15311 6011 19043 6018
rect 13327 5894 19043 6011
rect 13327 5785 19042 5894
rect 13327 5736 19043 5785
rect 13327 5734 15633 5736
rect 13327 5732 15420 5734
rect 13327 5728 15182 5732
rect 13327 5727 14750 5728
rect 13327 5718 13781 5727
rect 13327 5654 13556 5718
rect 13620 5663 13781 5718
rect 13845 5724 14279 5727
rect 13845 5663 14058 5724
rect 13620 5660 14058 5663
rect 14122 5663 14279 5724
rect 14343 5724 14750 5727
rect 14343 5663 14524 5724
rect 14122 5660 14524 5663
rect 14588 5664 14750 5724
rect 14814 5726 15182 5728
rect 14814 5664 14962 5726
rect 14588 5662 14962 5664
rect 15026 5668 15182 5726
rect 15246 5670 15420 5732
rect 15484 5672 15633 5734
rect 15697 5727 19043 5736
rect 15697 5726 16367 5727
rect 15697 5672 16020 5726
rect 15484 5670 16020 5672
rect 15246 5668 16020 5670
rect 15026 5662 16020 5668
rect 16084 5663 16367 5726
rect 16431 5724 19043 5727
rect 16431 5722 17026 5724
rect 16431 5663 16603 5722
rect 16084 5662 16603 5663
rect 14588 5660 16603 5662
rect 13620 5658 16603 5660
rect 16667 5658 16787 5722
rect 16851 5660 17026 5722
rect 17090 5723 19043 5724
rect 17090 5720 17796 5723
rect 17090 5660 17229 5720
rect 16851 5658 17229 5660
rect 13620 5656 17229 5658
rect 17293 5719 17796 5720
rect 17293 5717 17605 5719
rect 17293 5656 17414 5717
rect 13620 5654 17414 5656
rect 13327 5653 17414 5654
rect 17478 5655 17605 5717
rect 17669 5659 17796 5719
rect 17860 5719 19043 5723
rect 17860 5659 17982 5719
rect 17669 5655 17982 5659
rect 18046 5655 19043 5719
rect 17478 5653 19043 5655
rect 13327 5591 19043 5653
rect 12771 5138 18195 5525
rect 12771 5137 16144 5138
rect 12771 5136 13820 5137
rect 12771 5072 13429 5136
rect 13493 5132 13820 5136
rect 13493 5072 13634 5132
rect 12771 5068 13634 5072
rect 13698 5073 13820 5132
rect 13884 5135 16144 5137
rect 13884 5130 14233 5135
rect 13884 5073 14014 5130
rect 13698 5068 14014 5073
rect 12771 5066 14014 5068
rect 14078 5071 14233 5130
rect 14297 5071 14443 5135
rect 14507 5132 15926 5135
rect 14507 5071 14672 5132
rect 14078 5068 14672 5071
rect 14736 5068 14918 5132
rect 14982 5068 15192 5132
rect 15256 5068 15467 5132
rect 15531 5068 15703 5132
rect 15767 5071 15926 5132
rect 15990 5074 16144 5135
rect 16208 5136 18195 5138
rect 16208 5132 17589 5136
rect 16208 5131 17169 5132
rect 16208 5129 16561 5131
rect 16208 5074 16322 5129
rect 15990 5071 16322 5074
rect 15767 5068 16322 5071
rect 14078 5066 16322 5068
rect 12771 5065 16322 5066
rect 16386 5067 16561 5129
rect 16625 5067 16758 5131
rect 16822 5067 16956 5131
rect 17020 5068 17169 5131
rect 17233 5131 17589 5132
rect 17233 5068 17392 5131
rect 17020 5067 17392 5068
rect 17456 5072 17589 5131
rect 17653 5134 18195 5136
rect 17653 5072 17805 5134
rect 17456 5070 17805 5072
rect 17869 5070 18014 5134
rect 18078 5070 18195 5134
rect 17456 5067 18195 5070
rect 16386 5065 18195 5067
rect 12771 5040 18195 5065
use sky130_fd_sc_hd__dfbbp_1  x1[0] $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1699530450
transform 1 0 13370 0 -1 7564
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbp_1  x1[1]
timestamp 1699530450
transform 1 0 15762 0 -1 7564
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbp_1  x1[2]
timestamp 1699530450
transform 1 0 13370 0 1 6380
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbp_1  x1[3]
timestamp 1699530450
transform 1 0 15762 0 1 6380
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbp_1  x1[4]
timestamp 1699530450
transform 1 0 13370 0 -1 6284
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbp_1  x1[5]
timestamp 1699530450
transform 1 0 15762 0 -1 6284
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbp_1  x1[6]
timestamp 1699530450
transform 1 0 13370 0 1 5100
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbp_1  x1[7]
timestamp 1699530450
transform 1 0 15762 0 1 5100
box -38 -48 2430 592
use hgu_delay_no_code  x2
timestamp 1699326296
transform 1 0 2492 0 1 7675
box 9238 267 15997 2986
use sky130_fd_sc_hd__buf_2  x3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1699535479
transform 1 0 18472 0 1 9058
box -38 -48 406 592
<< labels >>
flabel metal4 11864 7966 12240 9403 0 FreeSans 320 0 0 0 VSS
port 31 nsew
flabel metal4 11836 10013 12254 10623 0 FreeSans 320 0 0 0 VDD
port 2 nsew
flabel metal1 11767 9271 11864 9318 0 FreeSans 320 0 0 0 eob
port 4 nsew
flabel metal1 13338 7918 14277 7946 0 FreeSans 320 0 0 0 delay_code[2]
port 6 nsew
flabel metal1 13338 7862 16703 7890 0 FreeSans 320 0 0 0 delay_code[1]
port 7 nsew
flabel metal1 13338 7806 17560 7834 0 FreeSans 320 0 0 0 delay_code[0]
port 8 nsew
flabel metal1 11730 9654 11784 9688 0 FreeSans 320 0 0 0 delay_code[3]
port 9 nsew
flabel metal1 13297 7232 13342 7280 0 FreeSans 320 0 0 0 sar_logic[0]
port 29 nsew
flabel metal1 13289 7438 13334 7486 0 FreeSans 320 0 0 0 sar_logic[1]
port 10 nsew
flabel metal1 13307 6591 13352 6639 0 FreeSans 320 0 0 0 sar_logic[2]
port 11 nsew
flabel metal1 13298 5954 13343 6002 0 FreeSans 320 0 0 0 sar_logic[4]
port 14 nsew
flabel metal1 13297 6157 13342 6205 0 FreeSans 320 0 0 0 sar_logic[5]
port 13 nsew
flabel metal1 18207 7428 18252 7476 0 FreeSans 320 0 0 0 sar_retimer[1]
port 17 nsew
flabel metal1 18207 7098 18252 7146 0 FreeSans 320 0 0 0 sar_retimer[0]
port 18 nsew
flabel metal1 18212 6457 18257 6505 0 FreeSans 320 0 0 0 sar_retimer[3]
port 19 nsew
flabel metal1 18207 6799 18252 6847 0 FreeSans 320 0 0 0 sar_retimer[2]
port 20 nsew
flabel metal1 18203 6147 18248 6195 0 FreeSans 320 0 0 0 sar_retimer[5]
port 21 nsew
flabel metal1 18206 5816 18251 5864 0 FreeSans 320 0 0 0 sar_retimer[4]
port 22 nsew
flabel metal1 18205 5176 18250 5224 0 FreeSans 320 0 0 0 sar_retimer[7]
port 23 nsew
flabel metal1 18209 5520 18254 5568 0 FreeSans 320 0 0 0 sar_retimer[6]
port 25 nsew
flabel metal1 13310 6457 13355 6505 0 FreeSans 320 0 0 0 sar_logic[3]
port 28 nsew
flabel metal1 13285 5376 13330 5424 0 FreeSans 320 0 0 0 sar_logic[6]
port 26 nsew
flabel metal1 13282 5177 13327 5225 0 FreeSans 320 0 0 0 sar_logic[7]
port 27 nsew
flabel metal1 12030 9069 12142 9117 0 FreeSans 320 0 0 0 delay_offset
port 32 nsew
<< end >>
