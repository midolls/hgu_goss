magic
tech sky130A
magscale 1 2
timestamp 1698581447
<< nmos >>
rect 143 757 173 841
rect 215 757 245 841
rect 287 757 317 841
rect 390 757 420 843
rect 462 757 492 843
rect 534 757 564 843
rect 606 757 636 843
rect 678 757 708 843
rect 750 757 780 843
<< ndiff >>
rect 332 841 390 843
rect 85 827 143 841
rect 85 771 94 827
rect 128 771 143 827
rect 85 757 143 771
rect 173 757 215 841
rect 245 757 287 841
rect 317 757 390 841
rect 420 757 462 843
rect 492 757 534 843
rect 564 757 606 843
rect 636 757 678 843
rect 708 757 750 843
rect 780 827 838 843
rect 780 771 791 827
rect 825 771 838 827
rect 780 757 838 771
<< ndiffc >>
rect 94 771 128 827
rect 791 771 825 827
<< poly >>
rect 742 888 786 903
rect 143 858 786 888
rect 143 841 173 858
rect 215 841 245 858
rect 287 841 317 858
rect 390 843 420 858
rect 462 843 492 858
rect 534 843 564 858
rect 606 843 636 858
rect 678 843 708 858
rect 750 843 780 858
rect 143 731 173 757
rect 215 731 245 757
rect 287 731 317 757
rect 390 731 420 757
rect 462 731 492 757
rect 534 731 564 757
rect 606 731 636 757
rect 678 731 708 757
rect 750 731 780 757
<< locali >>
rect 94 827 128 843
rect 94 755 128 771
rect 791 827 825 843
rect 791 755 825 771
<< end >>
