magic
tech sky130A
magscale 1 2
timestamp 1699706918
<< nwell >>
rect 984 3863 1018 3872
rect 984 3845 1039 3863
rect 984 3838 1018 3845
<< nsubdiff >>
rect 984 3863 1018 3872
rect 984 3845 1039 3863
rect 984 3838 1018 3845
<< poly >>
rect 1148 5162 1466 5192
rect 1532 5162 1658 5192
rect 1148 3979 1475 4010
rect 1440 3966 1475 3979
rect 1628 3989 1694 4010
rect 1440 3950 1507 3966
rect 1440 3916 1457 3950
rect 1491 3916 1507 3950
rect 1628 3955 1644 3989
rect 1678 3955 1694 3989
rect 1628 3943 1694 3955
rect 1440 3900 1507 3916
rect 1476 3631 1543 3647
rect 1476 3611 1493 3631
rect 1436 3597 1493 3611
rect 1527 3597 1543 3631
rect 1436 3581 1543 3597
rect 1617 3626 1684 3642
rect 1617 3592 1633 3626
rect 1667 3592 1684 3626
rect 1436 3568 1466 3581
rect 1617 3576 1684 3592
rect 1148 3537 1466 3568
rect 1628 3536 1658 3576
rect 1532 2905 1658 2935
rect 1532 2717 1658 2747
rect 1148 2084 1466 2115
rect 1436 2071 1466 2084
rect 1628 2076 1658 2116
rect 1436 2055 1543 2071
rect 1436 2041 1493 2055
rect 1476 2021 1493 2041
rect 1527 2021 1543 2055
rect 1476 2005 1543 2021
rect 1617 2060 1684 2076
rect 1617 2026 1633 2060
rect 1667 2026 1684 2060
rect 1617 2010 1684 2026
rect 1440 1736 1507 1752
rect 1440 1702 1457 1736
rect 1491 1702 1507 1736
rect 1440 1686 1507 1702
rect 1628 1697 1694 1709
rect 1440 1673 1475 1686
rect 1148 1642 1475 1673
rect 1628 1663 1644 1697
rect 1678 1663 1694 1697
rect 1628 1642 1694 1663
rect 1148 460 1466 491
rect 1532 460 1658 490
<< polycont >>
rect 1457 3916 1491 3950
rect 1644 3955 1678 3989
rect 1493 3597 1527 3631
rect 1633 3592 1667 3626
rect 1493 2021 1527 2055
rect 1633 2026 1667 2060
rect 1457 1702 1491 1736
rect 1644 1663 1678 1697
<< locali >>
rect 1628 3955 1644 3989
rect 1678 3955 1694 3989
rect 1441 3916 1457 3950
rect 1491 3916 1507 3950
rect 1018 3845 1039 3863
rect 1477 3597 1493 3631
rect 1527 3597 1543 3631
rect 1633 3626 1667 3642
rect 1633 3576 1667 3592
rect 995 2819 1026 2838
rect 1633 2060 1667 2076
rect 1477 2021 1493 2055
rect 1527 2021 1543 2055
rect 1633 2010 1667 2026
rect 1441 1702 1457 1736
rect 1491 1702 1507 1736
rect 1628 1663 1644 1697
rect 1678 1663 1694 1697
<< viali >>
rect 1644 3955 1678 3989
rect 1457 3916 1491 3950
rect 984 3838 1018 3872
rect 1493 3597 1527 3631
rect 1633 3592 1667 3626
rect 1493 2021 1527 2055
rect 1633 2026 1667 2060
rect 984 1783 1018 1817
rect 1457 1702 1491 1736
rect 1644 1663 1678 1697
<< metal1 >>
rect 1098 5175 1708 5209
rect 1098 5124 1132 5175
rect 1290 5124 1324 5175
rect 1482 5124 1516 5175
rect 1578 5124 1612 5175
rect 1674 5124 1708 5175
rect 1709 4036 1799 4070
rect 1635 4002 1687 4008
rect 1289 3975 1323 3980
rect 751 3903 877 3913
rect 751 3797 761 3903
rect 867 3879 877 3903
rect 867 3872 1030 3879
rect 867 3838 984 3872
rect 1018 3838 1030 3872
rect 867 3831 1030 3838
rect 867 3797 877 3831
rect 751 3787 877 3797
rect 1289 3573 1323 3974
rect 1448 3959 1500 3965
rect 1631 3955 1635 3989
rect 1687 3955 1691 3989
rect 1444 3916 1448 3950
rect 1500 3916 1504 3950
rect 1635 3944 1687 3950
rect 1448 3901 1500 3907
rect 1484 3640 1536 3646
rect 1633 3635 1667 3639
rect 1480 3597 1484 3631
rect 1536 3597 1540 3631
rect 1484 3582 1536 3588
rect 1618 3583 1624 3635
rect 1676 3583 1682 3635
rect 1633 3579 1667 3583
rect 1194 3539 1420 3573
rect 1765 3511 1799 4036
rect 1708 3477 1799 3511
rect 1714 3476 1799 3477
rect 1578 2888 1612 2973
rect 1674 2888 1708 2973
rect 1578 2679 1612 2764
rect 1674 2679 1708 2764
rect 1708 2141 1785 2175
rect 1194 2079 1420 2113
rect 748 1847 874 1857
rect 748 1741 758 1847
rect 864 1829 874 1847
rect 864 1817 1030 1829
rect 864 1783 984 1817
rect 1018 1783 1030 1817
rect 864 1771 1030 1783
rect 864 1741 874 1771
rect 748 1731 874 1741
rect 1289 1678 1323 2079
rect 1484 2064 1536 2070
rect 1633 2069 1667 2073
rect 1480 2021 1484 2055
rect 1536 2021 1540 2055
rect 1618 2017 1624 2069
rect 1676 2017 1682 2069
rect 1633 2013 1667 2017
rect 1484 2006 1536 2012
rect 1448 1745 1500 1751
rect 1444 1702 1448 1736
rect 1500 1702 1504 1736
rect 1635 1702 1687 1708
rect 1448 1687 1500 1693
rect 1289 1672 1323 1677
rect 1631 1663 1635 1697
rect 1687 1663 1691 1697
rect 1635 1644 1687 1650
rect 1751 1616 1785 2141
rect 1714 1582 1785 1616
rect 1098 477 1132 528
rect 1290 477 1324 528
rect 1482 477 1516 528
rect 1578 477 1612 528
rect 1674 477 1708 529
rect 1098 444 1708 477
rect 1098 443 1674 444
<< via1 >>
rect 1635 3989 1687 4002
rect 761 3797 867 3903
rect 1448 3950 1500 3959
rect 1635 3955 1644 3989
rect 1644 3955 1678 3989
rect 1678 3955 1687 3989
rect 1635 3950 1687 3955
rect 1448 3916 1457 3950
rect 1457 3916 1491 3950
rect 1491 3916 1500 3950
rect 1448 3907 1500 3916
rect 1484 3631 1536 3640
rect 1484 3597 1493 3631
rect 1493 3597 1527 3631
rect 1527 3597 1536 3631
rect 1484 3588 1536 3597
rect 1624 3626 1676 3635
rect 1624 3592 1633 3626
rect 1633 3592 1667 3626
rect 1667 3592 1676 3626
rect 1624 3583 1676 3592
rect 758 1741 864 1847
rect 1484 2055 1536 2064
rect 1484 2021 1493 2055
rect 1493 2021 1527 2055
rect 1527 2021 1536 2055
rect 1484 2012 1536 2021
rect 1624 2060 1676 2069
rect 1624 2026 1633 2060
rect 1633 2026 1667 2060
rect 1667 2026 1676 2060
rect 1624 2017 1676 2026
rect 1448 1736 1500 1745
rect 1448 1702 1457 1736
rect 1457 1702 1491 1736
rect 1491 1702 1500 1736
rect 1448 1693 1500 1702
rect 1635 1697 1687 1702
rect 1635 1663 1644 1697
rect 1644 1663 1678 1697
rect 1678 1663 1687 1697
rect 1635 1650 1687 1663
<< metal2 >>
rect 1629 4002 1694 4009
rect 1442 3959 1506 3965
rect 741 3787 751 3913
rect 877 3787 887 3913
rect 1442 3907 1448 3959
rect 1500 3907 1506 3959
rect 1629 3950 1635 4002
rect 1687 3972 1694 4002
rect 1687 3950 1701 3972
rect 1629 3944 1701 3950
rect 1442 3901 1506 3907
rect 1442 3738 1476 3901
rect 1667 3873 1701 3944
rect 1508 3864 1564 3873
rect 1508 3799 1564 3808
rect 1673 3864 1729 3873
rect 1673 3799 1729 3808
rect 1406 3682 1415 3738
rect 1471 3682 1480 3738
rect 1508 3646 1542 3799
rect 1570 3682 1580 3738
rect 1636 3721 1645 3738
rect 1636 3682 1660 3721
rect 1478 3640 1542 3646
rect 1626 3641 1660 3682
rect 1478 3588 1484 3640
rect 1536 3588 1542 3640
rect 1478 3582 1542 3588
rect 1618 3635 1682 3641
rect 1618 3583 1624 3635
rect 1676 3583 1682 3635
rect 1618 3577 1682 3583
rect 1478 2064 1542 2070
rect 1478 2012 1484 2064
rect 1536 2012 1542 2064
rect 1478 2006 1542 2012
rect 1618 2069 1682 2075
rect 1618 2017 1624 2069
rect 1676 2017 1682 2069
rect 1618 2011 1682 2017
rect 1406 1915 1415 1971
rect 1471 1915 1480 1971
rect 738 1731 748 1857
rect 874 1731 884 1857
rect 1442 1751 1476 1915
rect 1508 1853 1542 2006
rect 1626 1971 1660 2011
rect 1570 1915 1580 1971
rect 1636 1934 1660 1971
rect 1636 1915 1645 1934
rect 1508 1844 1564 1853
rect 1508 1779 1564 1788
rect 1673 1844 1729 1853
rect 1673 1779 1729 1788
rect 1442 1745 1506 1751
rect 1442 1693 1448 1745
rect 1500 1693 1506 1745
rect 1667 1708 1701 1779
rect 1442 1687 1506 1693
rect 1629 1702 1701 1708
rect 1629 1650 1635 1702
rect 1687 1680 1701 1702
rect 1687 1650 1694 1680
rect 1629 1643 1694 1650
<< via2 >>
rect 751 3903 877 3913
rect 751 3797 761 3903
rect 761 3797 867 3903
rect 867 3797 877 3903
rect 751 3787 877 3797
rect 1508 3808 1564 3864
rect 1673 3808 1729 3864
rect 1415 3682 1471 3738
rect 1580 3682 1636 3738
rect 1415 1915 1471 1971
rect 748 1847 874 1857
rect 748 1741 758 1847
rect 758 1741 864 1847
rect 864 1741 874 1847
rect 748 1731 874 1741
rect 1580 1915 1636 1971
rect 1508 1788 1564 1844
rect 1673 1788 1729 1844
<< metal3 >>
rect 735 3780 741 3920
rect 887 3780 893 3920
rect 1503 3864 1734 3869
rect 1503 3808 1508 3864
rect 1564 3808 1673 3864
rect 1729 3808 1734 3864
rect 1503 3803 1734 3808
rect 1406 3738 1641 3743
rect 1406 3682 1415 3738
rect 1471 3682 1580 3738
rect 1636 3682 1641 3738
rect 1406 3677 1641 3682
rect 1410 1971 1641 1977
rect 1410 1915 1415 1971
rect 1471 1915 1580 1971
rect 1636 1915 1641 1971
rect 1410 1909 1641 1915
rect 732 1724 738 1864
rect 884 1724 890 1864
rect 1503 1844 1734 1849
rect 1503 1788 1508 1844
rect 1564 1788 1673 1844
rect 1729 1788 1734 1844
rect 1503 1783 1734 1788
<< via3 >>
rect 741 3913 887 3920
rect 741 3787 751 3913
rect 751 3787 877 3913
rect 877 3787 887 3913
rect 741 3780 887 3787
rect 738 1857 884 1864
rect 738 1731 748 1857
rect 748 1731 874 1857
rect 874 1731 884 1857
rect 738 1724 884 1731
<< metal4 >>
rect 711 3920 917 3935
rect 711 3780 741 3920
rect 887 3780 917 3920
rect 711 1864 917 3780
rect 711 1724 738 1864
rect 884 1724 917 1864
rect 711 1688 917 1724
use sky130_fd_pr__nfet_01v8_5AY3TR  sky130_fd_pr__nfet_01v8_5AY3TR_0
timestamp 1699633464
transform 1 0 1595 0 1 3236
box -145 -427 227 482
use sky130_fd_pr__nfet_01v8_5AY3TR  sky130_fd_pr__nfet_01v8_5AY3TR_1
timestamp 1699633464
transform 1 0 1595 0 -1 2416
box -145 -427 227 482
use sky130_fd_pr__nfet_01v8_YCY3T5  sky130_fd_pr__nfet_01v8_YCY3T5_0
timestamp 1699631965
transform 1 0 1307 0 -1 2416
box -323 -427 401 482
use sky130_fd_pr__nfet_01v8_YCY3T5  sky130_fd_pr__nfet_01v8_YCY3T5_1
timestamp 1699631965
transform 1 0 1307 0 1 3236
box -323 -427 401 482
use sky130_fd_pr__pfet_01v8_UJB66J  sky130_fd_pr__pfet_01v8_UJB66J_0
timestamp 1699598487
transform 1 0 1595 0 -1 1066
box -399 -787 263 769
use sky130_fd_pr__pfet_01v8_UJB66J  sky130_fd_pr__pfet_01v8_UJB66J_1
timestamp 1699598487
transform 1 0 1595 0 1 4586
box -399 -787 263 769
use sky130_fd_pr__pfet_01v8_UJKTUG  sky130_fd_pr__pfet_01v8_UJKTUG_0
timestamp 1699600097
transform 1 0 1307 0 1 4586
box -359 -787 359 769
use sky130_fd_pr__pfet_01v8_UJKTUG  sky130_fd_pr__pfet_01v8_UJKTUG_1
timestamp 1699600097
transform 1 0 1307 0 -1 1066
box -359 -787 359 769
<< labels >>
flabel metal1 1293 3796 1316 3825 0 FreeSans 320 0 0 0 vip
port 3 nsew
flabel metal2 1632 3650 1656 3672 0 FreeSans 320 0 0 0 sw_n
port 8 nsew
flabel metal2 1674 3886 1698 3916 0 FreeSans 320 0 0 0 sw
port 10 nsew
flabel metal1 1770 3739 1795 3781 0 FreeSans 320 0 0 0 tah_vp
port 12 nsew
flabel metal1 1756 1869 1780 1907 0 FreeSans 320 0 0 0 tah_vn
port 14 nsew
flabel metal1 1292 1862 1320 1901 0 FreeSans 320 0 0 0 vin
port 16 nsew
flabel metal4 744 2724 881 2933 0 FreeSans 640 0 0 0 VDD
port 24 nsew
flabel metal2 1674 1728 1695 1760 0 FreeSans 320 0 0 0 sw
port 27 nsew
flabel metal2 1631 1982 1656 2002 0 FreeSans 320 0 0 0 sw_n
port 29 nsew
flabel locali 995 2819 1026 2838 0 FreeSans 320 0 0 0 VSS
port 35 nsew
<< end >>
