magic
tech sky130A
magscale 1 2
timestamp 1700485439
<< psubdiff >>
rect -87 5794 436 5840
rect 818 5794 1345 5840
rect 1983 5794 2878 5840
rect 4028 5794 5429 5840
rect 14738 5794 20301 5840
rect -109 5106 565 5152
rect 4598 5106 8013 5152
rect 10187 5106 15171 5152
rect 19393 5106 20225 5152
rect 20308 5106 20314 5152
<< poly >>
rect -249 5978 -179 6110
rect 656 5978 726 6110
rect 1437 6023 1891 6093
rect 2970 6023 3936 6093
rect 5521 6023 7511 6093
rect 10608 6023 14646 6093
rect 20393 6023 28527 6093
rect -271 5290 -201 5422
rect 657 5290 727 5422
rect 1921 5335 2375 5405
rect 3540 5335 4506 5405
rect 8105 5335 10095 5405
rect 15263 5335 19301 5405
rect 20317 5335 28451 5405
<< locali >>
rect -87 6374 436 6420
rect 818 6374 1345 6420
rect 1983 6374 2878 6420
rect 4028 6374 5429 6420
rect 7603 6374 10516 6420
rect 14738 6374 20301 6420
rect -87 5794 436 5840
rect 818 5794 1345 5840
rect 1983 5794 2878 5840
rect 4028 5794 5429 5840
rect 7603 5794 10516 5840
rect 14738 5794 20301 5840
rect -109 5686 565 5732
rect 947 5686 1829 5732
rect 2467 5686 3448 5732
rect 4598 5686 8013 5732
rect 10187 5686 15171 5732
rect 19393 5686 20264 5732
rect -109 5106 565 5152
rect 947 5106 1829 5152
rect 2467 5106 3448 5152
rect 4598 5106 8013 5152
rect 10187 5106 15171 5152
rect 19393 5106 20225 5152
rect 20308 5106 20314 5152
<< metal1 >>
rect 29502 6422 29566 6426
rect -95 6372 440 6422
rect 818 6372 1345 6422
rect 1983 6372 2878 6422
rect 4028 6372 5429 6422
rect 7603 6372 10516 6422
rect 14738 6372 20301 6422
rect 28616 6420 29566 6422
rect 28616 6372 29508 6420
rect 29502 6368 29508 6372
rect 29560 6368 29566 6420
rect 29502 6362 29566 6368
rect -87 6311 436 6343
rect 818 6311 1345 6343
rect 1983 6311 2878 6343
rect 4028 6311 5429 6343
rect 7603 6311 10516 6343
rect 14738 6311 20301 6343
rect 28619 6337 28783 6343
rect 28619 6311 28725 6337
rect 28719 6285 28725 6311
rect 28777 6285 28783 6337
rect 28719 6279 28783 6285
rect -95 6083 -31 6089
rect -95 6073 -89 6083
rect -133 6040 -89 6073
rect -95 6031 -89 6040
rect -37 6031 -31 6083
rect -95 6025 -31 6031
rect 357 6061 421 6067
rect 357 6009 363 6061
rect 415 6053 421 6061
rect 1268 6061 1332 6067
rect 415 6017 643 6053
rect 415 6009 421 6017
rect 357 6003 421 6009
rect 1268 6009 1274 6061
rect 1326 6050 1332 6061
rect 1326 6019 1553 6050
rect 2803 6049 2867 6055
rect 1326 6009 1332 6019
rect 1268 6003 1332 6009
rect 2803 5997 2809 6049
rect 2861 6038 2867 6049
rect 5353 6047 5417 6053
rect 2861 6009 3052 6038
rect 2861 5997 2867 6009
rect 2803 5991 2867 5997
rect 5353 5995 5359 6047
rect 5411 6036 5417 6047
rect 10326 6047 10390 6053
rect 5411 6007 5603 6036
rect 5411 5995 5417 6007
rect 5353 5989 5417 5995
rect 10326 5995 10332 6047
rect 10384 6036 10390 6047
rect 28631 6047 28695 6053
rect 28631 6036 28637 6047
rect 10384 6006 10690 6036
rect 28445 6007 28637 6036
rect 10384 5995 10390 6006
rect 10326 5989 10390 5995
rect 28631 5995 28637 6007
rect 28689 5995 28695 6047
rect 28631 5989 28695 5995
rect 28824 5843 28888 5849
rect 28824 5842 28830 5843
rect -87 5792 436 5842
rect 818 5792 1345 5842
rect 1983 5792 2878 5842
rect 4028 5792 5429 5842
rect 7603 5792 10516 5842
rect 14738 5792 20301 5842
rect 28619 5792 28830 5842
rect 28824 5791 28830 5792
rect 28882 5791 28888 5843
rect 28824 5785 28888 5791
rect 29504 5736 29568 5742
rect 29504 5734 29510 5736
rect -109 5684 565 5734
rect 947 5684 1829 5734
rect 2467 5684 3448 5734
rect 4598 5684 8013 5734
rect 10187 5684 15171 5734
rect 19393 5684 20264 5734
rect 28543 5684 29510 5734
rect 29562 5684 29568 5736
rect 29504 5678 29568 5684
rect -109 5623 565 5655
rect 947 5623 1829 5655
rect 2467 5623 3448 5655
rect 4598 5623 8013 5655
rect 10187 5623 15171 5655
rect 19393 5623 20264 5655
rect 28543 5649 28783 5655
rect 28543 5623 28725 5649
rect 28719 5597 28725 5623
rect 28777 5597 28783 5649
rect 28719 5591 28783 5597
rect 962 5401 1026 5407
rect 962 5394 968 5401
rect -95 5363 -31 5369
rect -95 5356 -89 5363
rect -173 5322 -89 5356
rect -95 5311 -89 5322
rect -37 5311 -31 5363
rect 773 5358 968 5394
rect 962 5349 968 5358
rect 1020 5349 1026 5401
rect 2480 5364 2544 5370
rect 2480 5354 2486 5364
rect 962 5343 1026 5349
rect 2293 5323 2486 5354
rect -95 5305 -31 5311
rect 2480 5312 2486 5323
rect 2538 5312 2544 5364
rect 4620 5359 4684 5365
rect 4620 5348 4626 5359
rect 4424 5319 4626 5348
rect 2480 5306 2544 5312
rect 4620 5307 4626 5319
rect 4678 5307 4684 5359
rect 10200 5362 10264 5368
rect 10200 5353 10206 5362
rect 10013 5324 10206 5353
rect 4620 5301 4684 5307
rect 10200 5310 10206 5324
rect 10258 5310 10264 5362
rect 19416 5358 19480 5364
rect 19416 5347 19422 5358
rect 19219 5318 19422 5347
rect 10200 5304 10264 5310
rect 19416 5306 19422 5318
rect 19474 5306 19480 5358
rect 19416 5300 19480 5306
rect 20149 5358 20213 5364
rect 20149 5306 20155 5358
rect 20207 5348 20213 5358
rect 20207 5319 20399 5348
rect 20207 5306 20213 5319
rect 20149 5300 20213 5306
rect 28825 5158 28889 5164
rect 28825 5154 28831 5158
rect -109 5104 565 5154
rect 947 5104 1829 5154
rect 2467 5104 3448 5154
rect 4598 5104 8013 5154
rect 10187 5104 15171 5154
rect 19393 5104 20225 5154
rect 28543 5106 28831 5154
rect 28883 5106 28889 5158
rect 28543 5104 28889 5106
rect 28825 5100 28889 5104
rect 150 4070 210 4078
rect 150 4018 154 4070
rect 206 4018 210 4070
rect 150 4007 210 4018
rect 162 3998 196 4007
rect 10327 3271 10391 3282
rect 10327 3219 10332 3271
rect 10384 3219 10391 3271
rect 10327 3208 10391 3219
rect 10341 3204 10375 3208
rect 28633 3177 28697 3183
rect 5352 3163 5418 3174
rect 2804 3131 2864 3137
rect 2804 3079 2808 3131
rect 2860 3079 2864 3131
rect 5352 3111 5358 3163
rect 5410 3111 5418 3163
rect 28633 3125 28639 3177
rect 28691 3125 28697 3177
rect 28633 3119 28697 3125
rect 28647 3114 28681 3119
rect 5352 3100 5418 3111
rect 5367 3096 5401 3100
rect 2804 3070 2864 3079
rect 2816 3059 2850 3070
rect 358 2914 418 2920
rect 358 2862 362 2914
rect 414 2862 418 2914
rect 358 2853 418 2862
rect 1270 2914 1330 2920
rect 1270 2862 1274 2914
rect 1326 2862 1330 2914
rect 1270 2853 1330 2862
rect 370 2842 404 2853
rect 1282 2842 1316 2853
rect -93 1954 -33 1960
rect -93 1902 -89 1954
rect -37 1902 -33 1954
rect -93 1896 -33 1902
rect -81 1882 -47 1896
rect 964 1815 1024 1821
rect 964 1763 968 1815
rect 1020 1763 1024 1815
rect 964 1754 1024 1763
rect 2482 1815 2542 1821
rect 2482 1763 2486 1815
rect 2538 1763 2542 1815
rect 2482 1754 2542 1763
rect 4620 1805 4684 1811
rect 976 1743 1010 1754
rect 2494 1743 2528 1754
rect 4620 1753 4626 1805
rect 4678 1753 4684 1805
rect 4620 1747 4684 1753
rect 10200 1807 10266 1818
rect 10200 1755 10206 1807
rect 10258 1755 10266 1807
rect 19417 1815 19481 1821
rect 19417 1763 19423 1815
rect 19475 1763 19481 1815
rect 19417 1757 19481 1763
rect 20149 1816 20213 1822
rect 20149 1764 20155 1816
rect 20207 1764 20213 1816
rect 20149 1758 20213 1764
rect 4634 1733 4668 1747
rect 10200 1744 10266 1755
rect 19431 1752 19465 1757
rect 20163 1753 20197 1758
rect 10215 1735 10249 1744
<< via1 >>
rect 29508 6368 29560 6420
rect 28725 6285 28777 6337
rect -89 6031 -37 6083
rect 363 6009 415 6061
rect 1274 6009 1326 6061
rect 2809 5997 2861 6049
rect 5359 5995 5411 6047
rect 10332 5995 10384 6047
rect 28637 5995 28689 6047
rect 28830 5791 28882 5843
rect 29510 5684 29562 5736
rect 28725 5597 28777 5649
rect -89 5311 -37 5363
rect 968 5349 1020 5401
rect 2486 5312 2538 5364
rect 4626 5307 4678 5359
rect 10206 5310 10258 5362
rect 19422 5306 19474 5358
rect 20155 5306 20207 5358
rect 28831 5106 28883 5158
rect 154 4018 206 4070
rect 10332 3219 10384 3271
rect 2808 3079 2860 3131
rect 5358 3111 5410 3163
rect 28639 3125 28691 3177
rect 362 2862 414 2914
rect 1274 2862 1326 2914
rect -89 1902 -37 1954
rect 968 1763 1020 1815
rect 2486 1763 2538 1815
rect 4626 1753 4678 1805
rect 10206 1755 10258 1807
rect 19423 1763 19475 1815
rect 20155 1764 20207 1816
<< metal2 >>
rect 29502 6420 29566 6426
rect 29502 6368 29508 6420
rect 29560 6368 29566 6420
rect 29502 6362 29566 6368
rect 28719 6337 28783 6343
rect 28719 6285 28725 6337
rect 28777 6285 28783 6337
rect -79 6248 196 6281
rect 28719 6279 28783 6285
rect -79 6089 -46 6248
rect -95 6083 -31 6089
rect -95 6031 -89 6083
rect -37 6031 -31 6083
rect -95 6025 -31 6031
rect -95 5363 -31 5369
rect -95 5311 -89 5363
rect -37 5311 -31 5363
rect -95 5305 -31 5311
rect -80 1965 -47 5305
rect 163 4081 196 6248
rect 357 6061 421 6067
rect 357 6009 363 6061
rect 415 6009 421 6061
rect 357 6003 421 6009
rect 1268 6061 1332 6067
rect 1268 6009 1274 6061
rect 1326 6009 1332 6061
rect 28734 6058 28768 6279
rect 29518 6060 29552 6362
rect 29753 6061 29828 6063
rect 29749 6060 29828 6061
rect 28946 6058 29021 6060
rect 1268 6003 1332 6009
rect 2803 6049 2867 6055
rect 371 5734 405 6003
rect 372 5684 405 5734
rect 150 4072 210 4081
rect 150 4016 152 4072
rect 208 4016 210 4072
rect 150 4007 210 4016
rect 371 2925 405 5684
rect 962 5401 1026 5407
rect 962 5349 968 5401
rect 1020 5349 1026 5401
rect 962 5343 1026 5349
rect 358 2916 418 2925
rect 358 2860 360 2916
rect 416 2860 418 2916
rect 358 2851 418 2860
rect -93 1956 -33 1965
rect -93 1900 -91 1956
rect -35 1900 -33 1956
rect -93 1891 -33 1900
rect 977 1826 1011 5343
rect 1283 2925 1317 6003
rect 2803 5997 2809 6049
rect 2861 5997 2867 6049
rect 2803 5991 2867 5997
rect 5353 6047 5417 6053
rect 5353 5995 5359 6047
rect 5411 5995 5417 6047
rect 1449 5173 1483 5603
rect 2480 5364 2544 5370
rect 2480 5312 2486 5364
rect 2538 5312 2544 5364
rect 2480 5306 2544 5312
rect 1270 2916 1330 2925
rect 1270 2860 1272 2916
rect 1328 2860 1330 2916
rect 1270 2851 1330 2860
rect 2495 1826 2529 5306
rect 2817 3142 2850 5991
rect 5353 5989 5417 5995
rect 10326 6047 10390 6053
rect 10326 5995 10332 6047
rect 10384 5995 10390 6047
rect 10326 5989 10390 5995
rect 28631 6047 28695 6053
rect 28631 5995 28637 6047
rect 28689 5995 28695 6047
rect 28631 5989 28695 5995
rect 28734 6051 29021 6058
rect 28734 5995 28955 6051
rect 29011 5995 29021 6051
rect 4620 5359 4684 5365
rect 4620 5307 4626 5359
rect 4678 5307 4684 5359
rect 4620 5301 4684 5307
rect 2804 3133 2864 3142
rect 2804 3077 2806 3133
rect 2862 3077 2864 3133
rect 2804 3068 2864 3077
rect 964 1817 1024 1826
rect 964 1761 966 1817
rect 1022 1761 1024 1817
rect 964 1752 1024 1761
rect 2482 1817 2542 1826
rect 2482 1761 2484 1817
rect 2540 1761 2542 1817
rect 4635 1816 4669 5301
rect 5367 3174 5401 5989
rect 10200 5362 10264 5368
rect 10200 5310 10206 5362
rect 10258 5310 10264 5362
rect 10200 5304 10264 5310
rect 5352 3165 5418 3174
rect 5352 3109 5357 3165
rect 5413 3109 5418 3165
rect 5352 3100 5418 3109
rect 10215 1818 10249 5304
rect 10341 3282 10375 5989
rect 19416 5358 19480 5364
rect 19416 5306 19422 5358
rect 19474 5306 19480 5358
rect 19416 5300 19480 5306
rect 20149 5358 20213 5364
rect 20149 5306 20155 5358
rect 20207 5306 20213 5358
rect 20149 5300 20213 5306
rect 10327 3273 10391 3282
rect 10327 3217 10331 3273
rect 10387 3217 10391 3273
rect 10327 3208 10391 3217
rect 19431 1826 19465 5300
rect 20163 1827 20197 5300
rect 28647 3188 28681 5989
rect 28734 5988 29021 5995
rect 28734 5655 28768 5988
rect 28946 5986 29021 5988
rect 29518 6054 29828 6060
rect 29518 5998 29762 6054
rect 29818 5998 29828 6054
rect 29518 5992 29828 5998
rect 28824 5843 28888 5849
rect 28824 5791 28830 5843
rect 28882 5791 28888 5843
rect 28824 5785 28888 5791
rect 28719 5649 28783 5655
rect 28719 5597 28725 5649
rect 28777 5597 28783 5649
rect 28719 5591 28783 5597
rect 28839 5429 28873 5785
rect 29518 5742 29552 5992
rect 29749 5991 29828 5992
rect 29753 5989 29828 5991
rect 29504 5736 29568 5742
rect 29504 5684 29510 5736
rect 29562 5684 29568 5736
rect 29504 5678 29568 5684
rect 28839 5425 28874 5429
rect 29142 5426 29217 5428
rect 29138 5425 29217 5426
rect 28839 5419 29217 5425
rect 28839 5363 29151 5419
rect 29207 5363 29217 5419
rect 28839 5357 29217 5363
rect 28839 5352 28874 5357
rect 29138 5356 29217 5357
rect 29142 5354 29217 5356
rect 28839 5164 28873 5352
rect 28825 5158 28889 5164
rect 28825 5106 28831 5158
rect 28883 5106 28889 5158
rect 28825 5100 28889 5106
rect 28633 3179 28697 3188
rect 28633 3123 28637 3179
rect 28693 3123 28697 3179
rect 28633 3114 28697 3123
rect 2482 1752 2542 1761
rect 4620 1807 4684 1816
rect 4620 1751 4624 1807
rect 4680 1751 4684 1807
rect 4620 1742 4684 1751
rect 10200 1809 10266 1818
rect 10200 1753 10205 1809
rect 10261 1753 10266 1809
rect 10200 1744 10266 1753
rect 19417 1817 19481 1826
rect 19417 1761 19421 1817
rect 19477 1761 19481 1817
rect 19417 1752 19481 1761
rect 20149 1818 20213 1827
rect 20149 1762 20153 1818
rect 20209 1762 20213 1818
rect 20149 1753 20213 1762
<< via2 >>
rect 152 4070 208 4072
rect 152 4018 154 4070
rect 154 4018 206 4070
rect 206 4018 208 4070
rect 152 4016 208 4018
rect 360 2914 416 2916
rect 360 2862 362 2914
rect 362 2862 414 2914
rect 414 2862 416 2914
rect 360 2860 416 2862
rect -91 1954 -35 1956
rect -91 1902 -89 1954
rect -89 1902 -37 1954
rect -37 1902 -35 1954
rect -91 1900 -35 1902
rect 1272 2914 1328 2916
rect 1272 2862 1274 2914
rect 1274 2862 1326 2914
rect 1326 2862 1328 2914
rect 1272 2860 1328 2862
rect 28955 5995 29011 6051
rect 2806 3131 2862 3133
rect 2806 3079 2808 3131
rect 2808 3079 2860 3131
rect 2860 3079 2862 3131
rect 2806 3077 2862 3079
rect 966 1815 1022 1817
rect 966 1763 968 1815
rect 968 1763 1020 1815
rect 1020 1763 1022 1815
rect 966 1761 1022 1763
rect 2484 1815 2540 1817
rect 2484 1763 2486 1815
rect 2486 1763 2538 1815
rect 2538 1763 2540 1815
rect 2484 1761 2540 1763
rect 5357 3163 5413 3165
rect 5357 3111 5358 3163
rect 5358 3111 5410 3163
rect 5410 3111 5413 3163
rect 5357 3109 5413 3111
rect 10331 3271 10387 3273
rect 10331 3219 10332 3271
rect 10332 3219 10384 3271
rect 10384 3219 10387 3271
rect 10331 3217 10387 3219
rect 29762 5998 29818 6054
rect 29151 5363 29207 5419
rect 28637 3177 28693 3179
rect 28637 3125 28639 3177
rect 28639 3125 28691 3177
rect 28691 3125 28693 3177
rect 28637 3123 28693 3125
rect 4624 1805 4680 1807
rect 4624 1753 4626 1805
rect 4626 1753 4678 1805
rect 4678 1753 4680 1805
rect 4624 1751 4680 1753
rect 10205 1807 10261 1809
rect 10205 1755 10206 1807
rect 10206 1755 10258 1807
rect 10258 1755 10261 1807
rect 10205 1753 10261 1755
rect 19421 1815 19477 1817
rect 19421 1763 19423 1815
rect 19423 1763 19475 1815
rect 19475 1763 19477 1815
rect 19421 1761 19477 1763
rect 20153 1816 20209 1818
rect 20153 1764 20155 1816
rect 20155 1764 20207 1816
rect 20207 1764 20209 1816
rect 20153 1762 20209 1764
<< metal3 >>
rect 28942 6055 29039 6075
rect 28942 5991 28951 6055
rect 29015 5991 29039 6055
rect 28942 5971 29039 5991
rect 29749 6058 29846 6078
rect 29749 5994 29758 6058
rect 29822 5994 29846 6058
rect 29749 5974 29846 5994
rect 29138 5423 29235 5443
rect 29138 5359 29147 5423
rect 29211 5359 29235 5423
rect 29138 5339 29235 5359
rect 150 4072 210 4087
rect 150 4016 152 4072
rect 208 4016 210 4072
rect 150 4007 210 4016
rect 10327 3203 10391 3213
rect 5352 3165 5367 3186
rect 5401 3165 5418 3186
rect 2804 3133 2864 3137
rect 2804 3077 2806 3133
rect 2862 3077 2864 3133
rect 5352 3109 5357 3165
rect 5413 3109 5418 3165
rect 5352 3096 5418 3109
rect 28632 3183 28633 3192
rect 28697 3183 28698 3192
rect 28632 3179 28698 3183
rect 28632 3157 28637 3179
rect 28632 3156 28636 3157
rect 28632 3123 28637 3156
rect 28693 3158 28698 3179
rect 28694 3157 28698 3158
rect 28693 3123 28698 3157
rect 28632 3122 28642 3123
rect 28643 3122 28698 3123
rect 28632 3102 28698 3122
rect 2804 3071 2864 3077
rect 2866 3059 2867 3060
rect 10205 2984 10261 2987
rect 358 2929 418 2931
rect 355 2916 421 2929
rect 355 2860 360 2916
rect 416 2860 421 2916
rect 355 2840 421 2860
rect 1267 2916 1333 2925
rect 1267 2860 1272 2916
rect 1328 2860 1333 2916
rect 1267 2850 1333 2860
rect 1268 2845 1332 2850
rect -93 1961 -33 1971
rect 2442 1894 2545 1904
rect 964 1821 1024 1832
rect 2482 1830 2542 1832
rect 2479 1821 2545 1830
rect 2479 1757 2480 1821
rect 2544 1757 2545 1821
rect 964 1752 1024 1757
rect 2479 1740 2545 1757
rect 4620 1812 4685 1828
rect 19416 1821 19482 1826
rect 4620 1748 4621 1812
rect 10200 1809 10266 1818
rect 10200 1753 10205 1809
rect 10261 1753 10266 1809
rect 4620 1733 4685 1748
rect 10200 1744 10266 1753
rect 19416 1757 19417 1821
rect 19481 1757 19482 1821
rect 19416 1740 19482 1757
<< via3 >>
rect 28951 6051 29015 6055
rect 28951 5995 28955 6051
rect 28955 5995 29011 6051
rect 29011 5995 29015 6051
rect 28951 5991 29015 5995
rect 29758 6054 29822 6058
rect 29758 5998 29762 6054
rect 29762 5998 29818 6054
rect 29818 5998 29822 6054
rect 29758 5994 29822 5998
rect 29147 5419 29211 5423
rect 29147 5363 29151 5419
rect 29151 5363 29207 5419
rect 29207 5363 29211 5419
rect 29147 5359 29211 5363
rect 962 1817 1026 1821
rect 962 1761 966 1817
rect 966 1761 1022 1817
rect 1022 1761 1026 1817
rect 962 1757 1026 1761
rect 2480 1817 2544 1821
rect 2480 1761 2484 1817
rect 2484 1761 2540 1817
rect 2540 1761 2544 1817
rect 2480 1757 2544 1761
<< metal4 >>
rect 29171 6320 29404 6321
rect 28942 6055 29404 6320
rect 28942 5991 28951 6055
rect 29015 5991 29404 6055
rect 28942 5756 29404 5991
rect 29171 5755 29404 5756
rect 29745 6058 30233 6365
rect 29745 5994 29758 6058
rect 29822 5994 30233 6058
rect 29745 5731 30233 5994
rect 29133 5423 29572 5639
rect 29133 5359 29147 5423
rect 29211 5359 29572 5423
rect 29133 5154 29572 5359
rect -209 4434 -158 4641
rect 150 3994 210 4087
rect 10327 3203 10391 3282
rect 5352 3163 5367 3186
rect 5401 3163 5418 3186
rect 5352 3096 5418 3163
rect 355 2840 421 2929
rect 8383 2928 8447 2992
rect 1267 2842 1333 2925
rect -93 1961 -33 1971
rect -93 1882 -33 1897
rect 964 1821 1024 1830
rect 2479 1821 2545 1830
rect 2479 1757 2480 1821
rect 2544 1757 2545 1821
rect 964 1740 1024 1757
rect 2479 1740 2545 1757
rect 4620 1812 4685 1828
rect 19417 1821 19481 1825
rect 4620 1748 4621 1812
rect 4620 1733 4685 1748
rect 10200 1744 10266 1818
rect 20148 1741 20214 1831
rect -205 1413 -161 1543
<< metal5 >>
rect 245 4094 565 5026
rect 1675 4100 1995 5026
rect 3259 4132 3579 5026
rect 5352 4142 5672 5026
rect 10326 4154 10646 5026
rect 39256 4154 39576 5026
rect 287 -595 524 -359
rect 1717 -595 1954 -359
rect 3301 -595 3538 -359
rect 5394 -595 5631 -359
rect 10368 -595 10605 -359
rect 39298 -595 39534 -359
use hgu_cdac_8bit_array  hgu_cdac_8bit_array_2
timestamp 1700482620
transform 1 0 4202 0 -1 -5445
box -4661 -7612 35404 -4800
use hgu_cdac_8bit_array  hgu_cdac_8bit_array_3
timestamp 1700482620
transform 1 0 4202 0 -1 -2312
box -4661 -7612 35404 -4800
use hgu_cdac_unit  hgu_cdac_unit_0
timestamp 1699890160
transform 1 0 -1145 0 -1 1399
box 686 598 1358 1826
use hgu_cdac_unit  hgu_cdac_unit_1
timestamp 1699890160
transform 1 0 -1145 0 -1 4532
box 686 598 1358 1826
use hgu_inverter  hgu_inverter_0
timestamp 1699345134
transform 1 0 -747 0 1 4944
box 347 160 675 824
use hgu_inverter  hgu_inverter_1
timestamp 1699345134
transform 1 0 -725 0 1 5632
box 347 160 675 824
use inv_2_test  inv_2_test_0
timestamp 1699782319
transform 1 0 128 0 1 2744
box 400 2360 856 3024
use inv_2_test  inv_2_test_1
timestamp 1699782319
transform 1 0 -1 0 1 3432
box 400 2360 856 3024
use inv_4_test  inv_4_test_1
timestamp 1699782319
transform 1 0 2239 0 1 3780
box -447 1324 265 1988
use inv_4_test  inv_4_test_2
timestamp 1699782319
transform 1 0 1755 0 1 4468
box -447 1324 265 1988
use inv_8_test  inv_8_test_0
timestamp 1699782319
transform 1 0 3315 0 1 2784
box 96 2320 1320 2984
use inv_8_test  inv_8_test_1
timestamp 1699782319
transform 1 0 2745 0 1 3472
box 96 2320 1320 2984
use inv_16_test  inv_16_test_0
timestamp 1699782319
transform 1 0 8625 0 1 5144
box -649 -40 1599 624
use inv_16_test  inv_16_test_1
timestamp 1699782319
transform 1 0 6041 0 1 5832
box -649 -40 1599 624
use inv_32_test  inv_32_test_0
timestamp 1699782319
transform 1 0 12782 0 1 8194
box -2303 -2402 1993 -1738
use inv_32_test  inv_32_test_1
timestamp 1699782319
transform 1 0 17437 0 1 7506
box -2303 -2402 1993 -1738
use inv_64_test  inv_64_test_0
timestamp 1699782319
transform 1 0 23771 0 1 7506
box -3583 -2402 4809 -1738
use inv_64_test  inv_64_test_1
timestamp 1699782319
transform 1 0 23847 0 1 8194
box -3583 -2402 4809 -1738
<< labels >>
flabel metal4 -209 4434 -158 4641 0 FreeSans 480 0 0 0 t<0>
port 27 nsew
flabel poly 2970 6023 3936 6093 0 FreeSans 320 0 0 0 d<3>
port 102 nsew
flabel poly 1437 6023 1891 6093 0 FreeSans 320 0 0 0 d<2>
port 104 nsew
flabel poly 656 5978 726 6110 0 FreeSans 320 0 0 0 d<1>
port 106 nsew
flabel poly -249 5978 -179 6110 0 FreeSans 320 0 0 0 d<0>
port 109 nsew
flabel poly 5521 6023 7511 6093 0 FreeSans 320 0 0 0 d<4>
port 111 nsew
flabel poly 10608 6023 14646 6093 0 FreeSans 320 0 0 0 d<5>
port 113 nsew
flabel poly 20393 6023 28527 6093 0 FreeSans 320 0 0 0 d<6>
port 115 nsew
flabel poly -271 5290 -201 5422 0 FreeSans 320 0 0 0 db<0>
port 117 nsew
flabel poly 657 5290 727 5422 0 FreeSans 320 0 0 0 db<1>
port 119 nsew
flabel poly 1921 5335 2375 5405 0 FreeSans 320 0 0 0 db<2>
port 121 nsew
flabel poly 3540 5335 4506 5405 0 FreeSans 320 0 0 0 db<3>
port 123 nsew
flabel poly 8105 5335 10095 5405 0 FreeSans 320 0 0 0 db<4>
port 125 nsew
flabel poly 15263 5335 19301 5405 0 FreeSans 320 0 0 0 db<5>
port 127 nsew
flabel poly 20317 5335 28451 5405 0 FreeSans 320 0 0 0 db<6>
port 133 nsew
flabel metal4 29211 5154 29572 5639 0 FreeSans 1600 0 0 0 VSS
port 159 nsew
flabel metal4 29822 5731 30233 6365 0 FreeSans 1600 0 0 0 VDD
port 161 nsew
flabel metal4 29015 5756 29404 6320 0 FreeSans 1600 0 0 0 VREF
port 163 nsew
flabel metal5 245 4094 565 5026 0 FreeSans 800 0 0 0 t<1>
port 166 nsew
flabel metal5 1675 4100 1995 5026 0 FreeSans 800 0 0 0 t<2>
port 168 nsew
flabel metal5 3259 4132 3579 5026 0 FreeSans 800 0 0 0 t<3>
port 170 nsew
flabel metal5 5352 4142 5672 5026 0 FreeSans 800 0 0 0 t<4>
port 172 nsew
flabel metal5 10326 4154 10646 5026 0 FreeSans 800 0 0 0 t<5>
port 176 nsew
flabel metal5 39256 4154 39576 5026 0 FreeSans 800 0 0 0 t<6>
port 178 nsew
flabel metal4 -205 1413 -161 1543 0 FreeSans 320 0 0 0 tb<0>
port 76 nsew
flabel metal5 287 -595 524 -359 0 FreeSans 480 0 0 0 tb<1>
port 147 nsew
flabel metal5 1717 -595 1954 -359 0 FreeSans 480 0 0 0 tb<2>
port 149 nsew
flabel metal5 3301 -595 3538 -359 0 FreeSans 480 0 0 0 tb<3>
port 151 nsew
flabel metal5 5394 -595 5631 -359 0 FreeSans 480 0 0 0 tb<4>
port 153 nsew
flabel metal5 10368 -595 10605 -359 0 FreeSans 480 0 0 0 tb<5>
port 155 nsew
flabel metal5 39298 -595 39534 -359 0 FreeSans 480 0 0 0 tb<6>
port 157 nsew
<< end >>
