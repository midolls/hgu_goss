magic
tech sky130A
timestamp 1699890160
<< psubdiff >>
rect 11352 1633 11373 1678
<< metal4 >>
rect 11260 1605 11283 1640
rect 11380 1403 11403 1438
rect 11319 1268 11342 1303
use hgu_cdac_unit  x1[0]
timestamp 1699890160
transform -1 0 7570 0 -1 2395
box 343 299 679 913
use hgu_cdac_unit  x1[1]
timestamp 1699890160
transform 1 0 6548 0 1 603
box 343 299 679 913
use hgu_cdac_unit  x1[2]
timestamp 1699890160
transform -1 0 7873 0 -1 2395
box 343 299 679 913
use hgu_cdac_unit  x1[3]
timestamp 1699890160
transform 1 0 6851 0 1 603
box 343 299 679 913
use hgu_cdac_unit  x1[4]
timestamp 1699890160
transform -1 0 8176 0 -1 2395
box 343 299 679 913
use hgu_cdac_unit  x1[5]
timestamp 1699890160
transform 1 0 7154 0 1 603
box 343 299 679 913
use hgu_cdac_unit  x1[6]
timestamp 1699890160
transform -1 0 8479 0 -1 2395
box 343 299 679 913
use hgu_cdac_unit  x1[7]
timestamp 1699890160
transform 1 0 7457 0 1 603
box 343 299 679 913
use hgu_cdac_unit  x1[8]
timestamp 1699890160
transform -1 0 8782 0 -1 2395
box 343 299 679 913
use hgu_cdac_unit  x1[9]
timestamp 1699890160
transform 1 0 7760 0 1 603
box 343 299 679 913
use hgu_cdac_unit  x1[10]
timestamp 1699890160
transform -1 0 9085 0 -1 2395
box 343 299 679 913
use hgu_cdac_unit  x1[11]
timestamp 1699890160
transform 1 0 8063 0 1 603
box 343 299 679 913
use hgu_cdac_unit  x1[12]
timestamp 1699890160
transform -1 0 9388 0 -1 2395
box 343 299 679 913
use hgu_cdac_unit  x1[13]
timestamp 1699890160
transform 1 0 8366 0 1 603
box 343 299 679 913
use hgu_cdac_unit  x1[14]
timestamp 1699890160
transform -1 0 9691 0 -1 2395
box 343 299 679 913
use hgu_cdac_unit  x1[15]
timestamp 1699890160
transform 1 0 8669 0 1 603
box 343 299 679 913
use hgu_cdac_unit  x1[16]
timestamp 1699890160
transform -1 0 9994 0 -1 2395
box 343 299 679 913
use hgu_cdac_unit  x1[17]
timestamp 1699890160
transform 1 0 8972 0 1 603
box 343 299 679 913
use hgu_cdac_unit  x1[18]
timestamp 1699890160
transform -1 0 10297 0 -1 2395
box 343 299 679 913
use hgu_cdac_unit  x1[19]
timestamp 1699890160
transform 1 0 9275 0 1 603
box 343 299 679 913
use hgu_cdac_unit  x1[20]
timestamp 1699890160
transform -1 0 10600 0 -1 2395
box 343 299 679 913
use hgu_cdac_unit  x1[21]
timestamp 1699890160
transform 1 0 9578 0 1 603
box 343 299 679 913
use hgu_cdac_unit  x1[22]
timestamp 1699890160
transform -1 0 10903 0 -1 2395
box 343 299 679 913
use hgu_cdac_unit  x1[23]
timestamp 1699890160
transform 1 0 9881 0 1 603
box 343 299 679 913
use hgu_cdac_unit  x1[24]
timestamp 1699890160
transform -1 0 11206 0 -1 2395
box 343 299 679 913
use hgu_cdac_unit  x1[25]
timestamp 1699890160
transform 1 0 10184 0 1 603
box 343 299 679 913
use hgu_cdac_unit  x1[26]
timestamp 1699890160
transform -1 0 11509 0 -1 2395
box 343 299 679 913
use hgu_cdac_unit  x1[27]
timestamp 1699890160
transform 1 0 10487 0 1 603
box 343 299 679 913
use hgu_cdac_unit  x1[28]
timestamp 1699890160
transform -1 0 11812 0 -1 2395
box 343 299 679 913
use hgu_cdac_unit  x1[29]
timestamp 1699890160
transform 1 0 10790 0 1 603
box 343 299 679 913
use hgu_cdac_unit  x1[30]
timestamp 1699890160
transform -1 0 12115 0 -1 2395
box 343 299 679 913
use hgu_cdac_unit  x1[31]
timestamp 1699890160
transform 1 0 11093 0 1 603
box 343 299 679 913
use hgu_cdac_unit  x1[32]
timestamp 1699890160
transform -1 0 12418 0 -1 2395
box 343 299 679 913
use hgu_cdac_unit  x1[33]
timestamp 1699890160
transform 1 0 11396 0 1 603
box 343 299 679 913
use hgu_cdac_unit  x1[34]
timestamp 1699890160
transform -1 0 12721 0 -1 2395
box 343 299 679 913
use hgu_cdac_unit  x1[35]
timestamp 1699890160
transform 1 0 11699 0 1 603
box 343 299 679 913
use hgu_cdac_unit  x1[36]
timestamp 1699890160
transform -1 0 13024 0 -1 2395
box 343 299 679 913
use hgu_cdac_unit  x1[37]
timestamp 1699890160
transform 1 0 12002 0 1 603
box 343 299 679 913
use hgu_cdac_unit  x1[38]
timestamp 1699890160
transform -1 0 13327 0 -1 2395
box 343 299 679 913
use hgu_cdac_unit  x1[39]
timestamp 1699890160
transform 1 0 12305 0 1 603
box 343 299 679 913
use hgu_cdac_unit  x1[40]
timestamp 1699890160
transform -1 0 13630 0 -1 2395
box 343 299 679 913
use hgu_cdac_unit  x1[41]
timestamp 1699890160
transform 1 0 12608 0 1 603
box 343 299 679 913
use hgu_cdac_unit  x1[42]
timestamp 1699890160
transform -1 0 13933 0 -1 2395
box 343 299 679 913
use hgu_cdac_unit  x1[43]
timestamp 1699890160
transform 1 0 12911 0 1 603
box 343 299 679 913
use hgu_cdac_unit  x1[44]
timestamp 1699890160
transform -1 0 14236 0 -1 2395
box 343 299 679 913
use hgu_cdac_unit  x1[45]
timestamp 1699890160
transform 1 0 13214 0 1 603
box 343 299 679 913
use hgu_cdac_unit  x1[46]
timestamp 1699890160
transform -1 0 14539 0 -1 2395
box 343 299 679 913
use hgu_cdac_unit  x1[47]
timestamp 1699890160
transform 1 0 13517 0 1 603
box 343 299 679 913
use hgu_cdac_unit  x1[48]
timestamp 1699890160
transform -1 0 14842 0 -1 2395
box 343 299 679 913
use hgu_cdac_unit  x1[49]
timestamp 1699890160
transform 1 0 13820 0 1 603
box 343 299 679 913
use hgu_cdac_unit  x1[50]
timestamp 1699890160
transform -1 0 15145 0 -1 2395
box 343 299 679 913
use hgu_cdac_unit  x1[51]
timestamp 1699890160
transform 1 0 14123 0 1 603
box 343 299 679 913
use hgu_cdac_unit  x1[52]
timestamp 1699890160
transform -1 0 15448 0 -1 2395
box 343 299 679 913
use hgu_cdac_unit  x1[53]
timestamp 1699890160
transform 1 0 14426 0 1 603
box 343 299 679 913
use hgu_cdac_unit  x1[54]
timestamp 1699890160
transform -1 0 15751 0 -1 2395
box 343 299 679 913
use hgu_cdac_unit  x1[55]
timestamp 1699890160
transform 1 0 14729 0 1 603
box 343 299 679 913
use hgu_cdac_unit  x1[56]
timestamp 1699890160
transform -1 0 16054 0 -1 2395
box 343 299 679 913
use hgu_cdac_unit  x1[57]
timestamp 1699890160
transform 1 0 15032 0 1 603
box 343 299 679 913
use hgu_cdac_unit  x1[58]
timestamp 1699890160
transform -1 0 16357 0 -1 2395
box 343 299 679 913
use hgu_cdac_unit  x1[59]
timestamp 1699890160
transform 1 0 15335 0 1 603
box 343 299 679 913
use hgu_cdac_unit  x1[60]
timestamp 1699890160
transform -1 0 16660 0 -1 2395
box 343 299 679 913
use hgu_cdac_unit  x1[61]
timestamp 1699890160
transform 1 0 15638 0 1 603
box 343 299 679 913
use hgu_cdac_unit  x1[62]
timestamp 1699890160
transform -1 0 16963 0 -1 2395
box 343 299 679 913
use hgu_cdac_unit  x1[63]
timestamp 1699890160
transform 1 0 15941 0 1 603
box 343 299 679 913
<< labels >>
flabel psubdiff 11352 1633 11373 1678 0 FreeSans 160 0 0 0 SUB
port 1 nsew
flabel metal4 11260 1605 11283 1640 0 FreeSans 160 0 0 0 CTOP
port 3 nsew
flabel metal4 11319 1268 11342 1303 0 FreeSans 160 0 0 0 CTOP
port 5 nsew
flabel metal4 11380 1403 11403 1438 0 FreeSans 160 0 0 0 CBOT
port 7 nsew
<< end >>
