* NGSPICE file created from hgu_cdac_half_flat.ext - technology: sky130A

.subckt hgu_cdac_half_flat d<3> d<2> d<1> d<0> d<4> d<5> d<6> db<0> db<1> db<2> db<3>
+ db<4> db<5> db<6> tb<1> tb<2> tb<3> tb<4> tb<5> VREF t<1> t<2> t<3> t<4> t<5> tb<0>
+ t<0> t<6> VDD tb<6> VSS
X0 hgu_cdac_8bit_array_3.drv<7:0> d<3> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1 VREF db<3> hgu_cdac_8bit_array_2.drv<7:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.35
X2 VREF d<5> hgu_cdac_8bit_array_3.drv<31:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3 VREF db<6> hgu_cdac_8bit_array_2.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X4 hgu_cdac_8bit_array_3.drv<31:0> d<5> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X5 hgu_cdac_8bit_array_2.drv<63:0> db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X6 VSS d<5> hgu_cdac_8bit_array_3.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X7 hgu_cdac_8bit_array_2.drv<31:0> db<5> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X8 hgu_cdac_8bit_array_3.drv<63:0> d<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X9 hgu_cdac_8bit_array_2.drv<63:0> db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X10 hgu_cdac_8bit_array_2.drv<63:0> db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X11 VREF d<6> hgu_cdac_8bit_array_3.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X12 VSS d<6> hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X13 VSS d<1> hgu_cdac_8bit_array_3.drv<1:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.35
X14 hgu_cdac_8bit_array_3.drv<63:0> d<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X15 hgu_cdac_8bit_array_3.drv<31:0> d<5> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X16 VREF db<6> hgu_cdac_8bit_array_2.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X17 VSS d<5> hgu_cdac_8bit_array_3.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X18 hgu_cdac_8bit_array_2.drv<31:0> db<5> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X19 hgu_cdac_8bit_array_2.drv<63:0> db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X20 hgu_cdac_8bit_array_2.drv<15:0> db<4> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X21 hgu_cdac_8bit_array_3.drv<63:0> d<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X22 VSS d<6> hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.35
X23 VSS db<4> hgu_cdac_8bit_array_2.drv<15:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X24 hgu_cdac_8bit_array_2.drv<63:0> db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X25 hgu_cdac_8bit_array_3.drv<15:0> d<4> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X26 VSS d<6> hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X27 VREF d<5> hgu_cdac_8bit_array_3.drv<31:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X28 VSS db<5> hgu_cdac_8bit_array_2.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X29 hgu_cdac_8bit_array_2.drv<63:0> db<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X30 VSS db<6> hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X31 hgu_cdac_8bit_array_2.drv<1:0> db<1> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.122 ps=1.42 w=0.42 l=0.35
X32 hgu_cdac_8bit_array_3.drv<31:0> d<5> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X33 VSS d<5> hgu_cdac_8bit_array_3.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X34 hgu_cdac_8bit_array_3.drv<63:0> d<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X35 VSS db<6> hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X36 hgu_cdac_8bit_array_2.drv<7:0> db<3> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X37 VREF db<6> hgu_cdac_8bit_array_2.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X38 hgu_cdac_8bit_array_2.drv<31:0> db<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X39 hgu_cdac_8bit_array_3.drv<63:0> d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X40 hgu_cdac_8bit_array_3.drv<15:0> d<4> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X41 VSS db<5> hgu_cdac_8bit_array_2.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X42 hgu_cdac_8bit_array_2.drv<63:0> db<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X43 VSS d<6> hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X44 VREF db<5> hgu_cdac_8bit_array_2.drv<31:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X45 hgu_cdac_8bit_array_2.drv<7:0> db<3> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.35
X46 VREF d<6> hgu_cdac_8bit_array_3.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X47 VREF db<2> hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X48 VSS d<4> hgu_cdac_8bit_array_3.drv<15:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.35
X49 hgu_cdac_8bit_array_3.drv<31:0> d<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X50 VREF db<6> hgu_cdac_8bit_array_2.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X51 VREF db<5> hgu_cdac_8bit_array_2.drv<31:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X52 VREF d<6> hgu_cdac_8bit_array_3.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X53 VREF db<6> hgu_cdac_8bit_array_2.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X54 hgu_cdac_8bit_array_2.drv<31:0> db<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X55 hgu_cdac_8bit_array_3.drv<63:0> d<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X56 VSS d<6> hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X57 hgu_cdac_8bit_array_3.drv<15:0> d<4> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X58 VREF d<6> hgu_cdac_8bit_array_3.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X59 hgu_cdac_8bit_array_2.drv<63:0> db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X60 VSS d<6> hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X61 hgu_cdac_8bit_array_3.drv<31:0> d<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X62 VSS d<3> hgu_cdac_8bit_array_3.drv<7:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X63 VREF db<6> hgu_cdac_8bit_array_2.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X64 hgu_cdac_8bit_array_2.drv<31:0> db<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X65 hgu_cdac_8bit_array_3.drv<63:0> d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X66 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT db<2> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X67 hgu_cdac_8bit_array_3.drv<63:0> d<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X68 hgu_cdac_8bit_array_2.drv<0> db<0> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.35
X69 hgu_cdac_8bit_array_3.drv<7:0> d<3> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X70 VSS d<3> hgu_cdac_8bit_array_3.drv<7:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X71 hgu_cdac_8bit_array_2.drv<63:0> db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X72 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT d<2> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X73 hgu_cdac_8bit_array_2.drv<31:0> db<5> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X74 VSS d<6> hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X75 VREF d<5> hgu_cdac_8bit_array_3.drv<31:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X76 VSS d<6> hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X77 VREF db<4> hgu_cdac_8bit_array_2.drv<15:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X78 hgu_cdac_8bit_array_2.drv<63:0> db<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X79 hgu_cdac_8bit_array_3.drv<31:0> d<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X80 VSS db<6> hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X81 VSS db<6> hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X82 VREF d<6> hgu_cdac_8bit_array_3.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X83 VREF db<6> hgu_cdac_8bit_array_2.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X84 VREF d<1> hgu_cdac_8bit_array_3.drv<1:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.35
X85 hgu_cdac_8bit_array_2.drv<15:0> db<4> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X86 hgu_cdac_8bit_array_2.drv<31:0> db<5> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.35
X87 VREF d<5> hgu_cdac_8bit_array_3.drv<31:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X88 hgu_cdac_8bit_array_2.drv<63:0> db<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X89 VSS d<6> hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X90 VREF db<6> hgu_cdac_8bit_array_2.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X91 VREF db<4> hgu_cdac_8bit_array_2.drv<15:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X92 hgu_cdac_8bit_array_2.drv<63:0> db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X93 VREF d<6> hgu_cdac_8bit_array_3.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.35
X94 hgu_cdac_8bit_array_3.drv<31:0> d<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X95 VSS db<6> hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X96 VREF d<6> hgu_cdac_8bit_array_3.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X97 hgu_cdac_8bit_array_2.drv<15:0> db<4> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.122 ps=1.42 w=0.42 l=0.35
X98 VREF db<6> hgu_cdac_8bit_array_2.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X99 hgu_cdac_8bit_array_2.drv<15:0> db<4> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X100 VREF db<3> hgu_cdac_8bit_array_2.drv<7:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X101 VREF d<5> hgu_cdac_8bit_array_3.drv<31:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X102 VREF db<6> hgu_cdac_8bit_array_2.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X103 hgu_cdac_8bit_array_3.drv<63:0> d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X104 hgu_cdac_8bit_array_2.drv<63:0> db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X105 hgu_cdac_8bit_array_3.drv<63:0> d<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X106 VSS d<6> hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X107 VSS db<5> hgu_cdac_8bit_array_2.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X108 VREF db<5> hgu_cdac_8bit_array_2.drv<31:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.35
X109 VSS db<6> hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.35
X110 VREF db<6> hgu_cdac_8bit_array_2.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X111 VREF d<6> hgu_cdac_8bit_array_3.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X112 hgu_cdac_8bit_array_2.drv<31:0> db<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X113 VSS db<5> hgu_cdac_8bit_array_2.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X114 hgu_cdac_8bit_array_2.drv<15:0> db<4> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X115 hgu_cdac_8bit_array_2.drv<63:0> db<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X116 VREF d<4> hgu_cdac_8bit_array_3.drv<15:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.35
X117 hgu_cdac_8bit_array_3.drv<15:0> d<4> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X118 VSS d<4> hgu_cdac_8bit_array_3.drv<15:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X119 hgu_cdac_8bit_array_3.drv<31:0> d<5> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X120 VSS d<5> hgu_cdac_8bit_array_3.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X121 hgu_cdac_8bit_array_2.drv<31:0> db<5> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X122 hgu_cdac_8bit_array_3.drv<7:0> d<3> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X123 hgu_cdac_8bit_array_2.drv<15:0> db<4> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X124 VSS d<6> hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X125 hgu_cdac_8bit_array_2.drv<7:0> db<3> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X126 hgu_cdac_8bit_array_3.drv<31:0> d<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X127 VREF d<6> hgu_cdac_8bit_array_3.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X128 hgu_cdac_8bit_array_2.drv<63:0> db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X129 hgu_cdac_8bit_array_3.drv<15:0> d<4> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X130 VSS db<5> hgu_cdac_8bit_array_2.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X131 hgu_cdac_8bit_array_2.drv<63:0> db<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X132 VSS d<6> hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X133 VSS db<2> hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT VSS sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.35
X134 VREF d<6> hgu_cdac_8bit_array_3.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X135 hgu_cdac_8bit_array_3.drv<31:0> d<5> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X136 VREF d<3> hgu_cdac_8bit_array_3.drv<7:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X137 hgu_cdac_8bit_array_3.drv<7:0> d<3> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X138 hgu_cdac_8bit_array_2.drv<31:0> db<5> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X139 VSS d<2> hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT VSS sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.35
X140 VREF db<5> hgu_cdac_8bit_array_2.drv<31:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X141 hgu_cdac_8bit_array_2.drv<15:0> db<4> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X142 hgu_cdac_8bit_array_3.drv<63:0> d<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X143 VSS d<6> hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X144 VREF db<6> hgu_cdac_8bit_array_2.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X145 VSS d<6> hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X146 VREF d<3> hgu_cdac_8bit_array_3.drv<7:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X147 hgu_cdac_8bit_array_2.drv<63:0> db<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X148 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT d<2> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X149 VSS db<5> hgu_cdac_8bit_array_2.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X150 VREF d<6> hgu_cdac_8bit_array_3.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X151 VREF d<6> hgu_cdac_8bit_array_3.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X152 VSS d<4> hgu_cdac_8bit_array_3.drv<15:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X153 VSS db<6> hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X154 hgu_cdac_8bit_array_3.drv<31:0> d<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X155 VREF db<6> hgu_cdac_8bit_array_2.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X156 hgu_cdac_8bit_array_3.drv<63:0> d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X157 hgu_cdac_8bit_array_3.drv<31:0> d<5> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X158 hgu_cdac_8bit_array_2.drv<63:0> db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X159 hgu_cdac_8bit_array_2.drv<63:0> db<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X160 VSS db<5> hgu_cdac_8bit_array_2.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X161 hgu_cdac_8bit_array_2.drv<7:0> db<3> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X162 hgu_cdac_8bit_array_2.drv<63:0> db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X163 VREF d<6> hgu_cdac_8bit_array_3.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X164 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT db<2> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.122 ps=1.42 w=0.42 l=0.35
X165 VSS d<4> hgu_cdac_8bit_array_3.drv<15:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X166 VSS db<5> hgu_cdac_8bit_array_2.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X167 hgu_cdac_8bit_array_2.drv<63:0> db<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X168 VSS d<6> hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X169 VREF db<5> hgu_cdac_8bit_array_2.drv<31:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X170 hgu_cdac_8bit_array_3.drv<63:0> d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X171 hgu_cdac_8bit_array_3.drv<31:0> d<5> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X172 hgu_cdac_8bit_array_3.drv<63:0> d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X173 hgu_cdac_8bit_array_2.drv<63:0> db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X174 hgu_cdac_8bit_array_3.drv<63:0> d<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X175 VSS db<5> hgu_cdac_8bit_array_2.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X176 hgu_cdac_8bit_array_2.drv<63:0> db<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X177 VSS d<6> hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X178 VSS db<4> hgu_cdac_8bit_array_2.drv<15:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X179 hgu_cdac_8bit_array_2.drv<63:0> db<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X180 VREF d<6> hgu_cdac_8bit_array_3.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X181 hgu_cdac_8bit_array_3.drv<63:0> d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X182 hgu_cdac_8bit_array_2.drv<63:0> db<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X183 VSS db<6> hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X184 hgu_cdac_8bit_array_3.drv<63:0> d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X185 VSS db<3> hgu_cdac_8bit_array_2.drv<7:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X186 VSS d<5> hgu_cdac_8bit_array_3.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X187 hgu_cdac_8bit_array_3.drv<15:0> d<4> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X188 VSS db<6> hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X189 VREF d<4> hgu_cdac_8bit_array_3.drv<15:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X190 VSS db<4> hgu_cdac_8bit_array_2.drv<15:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X191 hgu_cdac_8bit_array_2.drv<63:0> db<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X192 hgu_cdac_8bit_array_3.drv<7:0> d<3> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X193 VREF d<5> hgu_cdac_8bit_array_3.drv<31:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X194 VREF db<4> hgu_cdac_8bit_array_2.drv<15:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X195 VREF d<6> hgu_cdac_8bit_array_3.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X196 hgu_cdac_8bit_array_3.drv<31:0> d<5> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X197 hgu_cdac_8bit_array_2.drv<63:0> db<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X198 VSS db<6> hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X199 hgu_cdac_8bit_array_3.drv<31:0> d<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X200 VREF db<6> hgu_cdac_8bit_array_2.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X201 VREF db<5> hgu_cdac_8bit_array_2.drv<31:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X202 VREF d<6> hgu_cdac_8bit_array_3.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X203 hgu_cdac_8bit_array_3.drv<63:0> d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X204 hgu_cdac_8bit_array_2.drv<1:0> db<1> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.35
X205 VSS db<6> hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X206 hgu_cdac_8bit_array_3.drv<7:0> d<3> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X207 hgu_cdac_8bit_array_2.drv<31:0> db<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X208 VREF db<6> hgu_cdac_8bit_array_2.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X209 hgu_cdac_8bit_array_3.drv<63:0> d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X210 VREF d<2> hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT VDD sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.35
X211 hgu_cdac_8bit_array_2.drv<7:0> db<3> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X212 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT d<2> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.122 ps=1.42 w=0.42 l=0.35
X213 hgu_cdac_8bit_array_2.drv<63:0> db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X214 hgu_cdac_8bit_array_2.drv<31:0> db<5> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X215 VREF d<6> hgu_cdac_8bit_array_3.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X216 hgu_cdac_8bit_array_3.drv<15:0> d<4> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X217 hgu_cdac_8bit_array_3.drv<31:0> d<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X218 VREF db<5> hgu_cdac_8bit_array_2.drv<31:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X219 VREF d<6> hgu_cdac_8bit_array_3.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X220 VREF d<4> hgu_cdac_8bit_array_3.drv<15:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X221 hgu_cdac_8bit_array_2.drv<31:0> db<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X222 hgu_cdac_8bit_array_3.drv<63:0> d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X223 hgu_cdac_8bit_array_3.drv<15:0> d<4> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X224 hgu_cdac_8bit_array_3.drv<31:0> d<5> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X225 hgu_cdac_8bit_array_2.drv<63:0> db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X226 hgu_cdac_8bit_array_3.drv<63:0> d<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X227 hgu_cdac_8bit_array_2.drv<31:0> db<5> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X228 VSS d<6> hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X229 VSS db<1> hgu_cdac_8bit_array_2.drv<1:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.35
X230 hgu_cdac_8bit_array_3.drv<63:0> d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X231 VSS db<3> hgu_cdac_8bit_array_2.drv<7:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X232 hgu_cdac_8bit_array_2.drv<63:0> db<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X233 VSS d<6> hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X234 VSS db<5> hgu_cdac_8bit_array_2.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X235 VSS d<6> hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X236 VREF d<4> hgu_cdac_8bit_array_3.drv<15:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X237 VREF d<6> hgu_cdac_8bit_array_3.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X238 hgu_cdac_8bit_array_2.drv<31:0> db<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X239 hgu_cdac_8bit_array_3.drv<63:0> d<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X240 hgu_cdac_8bit_array_2.drv<31:0> db<5> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X241 hgu_cdac_8bit_array_3.drv<63:0> d<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X242 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT db<2> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X243 hgu_cdac_8bit_array_2.drv<0> db<0> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.244 ps=2.26 w=0.84 l=0.35
X244 VSS db<4> hgu_cdac_8bit_array_2.drv<15:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.35
X245 VSS d<5> hgu_cdac_8bit_array_3.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X246 hgu_cdac_8bit_array_2.drv<63:0> db<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X247 VSS db<6> hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X248 hgu_cdac_8bit_array_3.drv<31:0> d<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X249 VREF d<6> hgu_cdac_8bit_array_3.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X250 hgu_cdac_8bit_array_2.drv<63:0> db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X251 hgu_cdac_8bit_array_2.drv<15:0> db<4> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X252 hgu_cdac_8bit_array_3.drv<63:0> d<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X253 VSS db<6> hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X254 VREF db<6> hgu_cdac_8bit_array_2.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X255 VREF db<6> hgu_cdac_8bit_array_2.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X256 hgu_cdac_8bit_array_3.drv<63:0> d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X257 hgu_cdac_8bit_array_2.drv<15:0> db<4> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X258 hgu_cdac_8bit_array_3.drv<63:0> d<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X259 VREF d<5> hgu_cdac_8bit_array_3.drv<31:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X260 hgu_cdac_8bit_array_2.drv<63:0> db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.122 ps=1.42 w=0.42 l=0.35
X261 hgu_cdac_8bit_array_2.drv<63:0> db<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X262 VSS db<6> hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X263 hgu_cdac_8bit_array_2.drv<31:0> db<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X264 VREF db<6> hgu_cdac_8bit_array_2.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X265 hgu_cdac_8bit_array_3.drv<63:0> d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X266 VSS d<4> hgu_cdac_8bit_array_3.drv<15:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X267 hgu_cdac_8bit_array_3.drv<31:0> d<5> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X268 hgu_cdac_8bit_array_2.drv<15:0> db<4> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.35
X269 hgu_cdac_8bit_array_3.drv<63:0> d<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X270 hgu_cdac_8bit_array_2.drv<15:0> db<4> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X271 hgu_cdac_8bit_array_2.drv<63:0> db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X272 hgu_cdac_8bit_array_2.drv<63:0> db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X273 hgu_cdac_8bit_array_3.drv<63:0> d<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X274 hgu_cdac_8bit_array_2.drv<63:0> db<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X275 VSS d<6> hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X276 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT d<2> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.35
X277 VSS db<5> hgu_cdac_8bit_array_2.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X278 VSS db<4> hgu_cdac_8bit_array_2.drv<15:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X279 VREF db<5> hgu_cdac_8bit_array_2.drv<31:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X280 hgu_cdac_8bit_array_3.drv<15:0> d<4> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X281 VSS d<4> hgu_cdac_8bit_array_3.drv<15:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X282 hgu_cdac_8bit_array_3.drv<31:0> d<5> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X283 VREF db<6> hgu_cdac_8bit_array_2.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.35
X284 hgu_cdac_8bit_array_2.drv<31:0> db<5> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X285 hgu_cdac_8bit_array_3.drv<31:0> d<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.122 ps=1.42 w=0.42 l=0.35
X286 VREF db<5> hgu_cdac_8bit_array_2.drv<31:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X287 hgu_cdac_8bit_array_2.drv<15:0> db<4> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X288 VSS d<5> hgu_cdac_8bit_array_3.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X289 hgu_cdac_8bit_array_2.drv<63:0> db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X290 hgu_cdac_8bit_array_3.drv<15:0> d<4> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X291 VSS d<6> hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X292 hgu_cdac_8bit_array_3.drv<63:0> d<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X293 VSS d<6> hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X294 VSS db<4> hgu_cdac_8bit_array_2.drv<15:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X295 hgu_cdac_8bit_array_3.drv<63:0> d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X296 VREF d<6> hgu_cdac_8bit_array_3.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X297 hgu_cdac_8bit_array_2.drv<7:0> db<3> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X298 hgu_cdac_8bit_array_2.drv<63:0> db<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X299 VREF db<5> hgu_cdac_8bit_array_2.drv<31:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X300 hgu_cdac_8bit_array_3.drv<63:0> d<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X301 VSS db<6> hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X302 hgu_cdac_8bit_array_3.drv<31:0> d<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X303 VREF d<6> hgu_cdac_8bit_array_3.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X304 VREF d<6> hgu_cdac_8bit_array_3.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X305 VREF db<2> hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT VDD sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.35
X306 hgu_cdac_8bit_array_3.drv<63:0> d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X307 VSS d<5> hgu_cdac_8bit_array_3.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X308 hgu_cdac_8bit_array_2.drv<63:0> db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X309 VSS d<4> hgu_cdac_8bit_array_3.drv<15:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X310 VREF d<5> hgu_cdac_8bit_array_3.drv<31:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X311 VSS db<6> hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X312 hgu_cdac_8bit_array_3.drv<31:0> d<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X313 VREF db<5> hgu_cdac_8bit_array_2.drv<31:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X314 VSS d<3> hgu_cdac_8bit_array_3.drv<7:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.35
X315 hgu_cdac_8bit_array_2.drv<63:0> db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X316 hgu_cdac_8bit_array_3.drv<63:0> d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X317 hgu_cdac_8bit_array_3.drv<31:0> d<5> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X318 hgu_cdac_8bit_array_2.drv<31:0> db<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X319 VREF db<6> hgu_cdac_8bit_array_2.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X320 hgu_cdac_8bit_array_3.drv<63:0> d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X321 hgu_cdac_8bit_array_2.drv<63:0> db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X322 hgu_cdac_8bit_array_3.drv<63:0> d<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X323 hgu_cdac_8bit_array_2.drv<63:0> db<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X324 hgu_cdac_8bit_array_3.drv<15:0> d<4> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.122 ps=1.42 w=0.42 l=0.35
X325 VSS d<3> hgu_cdac_8bit_array_3.drv<7:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X326 VREF db<5> hgu_cdac_8bit_array_2.drv<31:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X327 hgu_cdac_8bit_array_2.drv<7:0> db<3> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X328 hgu_cdac_8bit_array_2.drv<63:0> db<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X329 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT db<2> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.35
X330 VREF db<5> hgu_cdac_8bit_array_2.drv<31:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X331 VSS db<6> hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X332 hgu_cdac_8bit_array_2.drv<31:0> db<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X333 hgu_cdac_8bit_array_3.drv<63:0> d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X334 VSS db<6> hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X335 hgu_cdac_8bit_array_3.drv<63:0> d<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X336 VREF d<4> hgu_cdac_8bit_array_3.drv<15:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X337 hgu_cdac_8bit_array_3.drv<1:0> d<1> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.122 ps=1.42 w=0.42 l=0.35
X338 VSS d<5> hgu_cdac_8bit_array_3.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X339 hgu_cdac_8bit_array_2.drv<63:0> db<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X340 VSS d<6> hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X341 VREF db<5> hgu_cdac_8bit_array_2.drv<31:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X342 VSS db<6> hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X343 VREF db<4> hgu_cdac_8bit_array_2.drv<15:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X344 VREF d<6> hgu_cdac_8bit_array_3.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X345 hgu_cdac_8bit_array_3.drv<63:0> d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X346 VSS db<3> hgu_cdac_8bit_array_2.drv<7:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.35
X347 VSS db<6> hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X348 VREF d<4> hgu_cdac_8bit_array_3.drv<15:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X349 hgu_cdac_8bit_array_3.drv<31:0> d<5> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.35
X350 hgu_cdac_8bit_array_2.drv<31:0> db<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X351 VREF db<6> hgu_cdac_8bit_array_2.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X352 hgu_cdac_8bit_array_3.drv<63:0> d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X353 VREF db<3> hgu_cdac_8bit_array_2.drv<7:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X354 hgu_cdac_8bit_array_3.drv<7:0> d<3> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.122 ps=1.42 w=0.42 l=0.35
X355 VREF db<6> hgu_cdac_8bit_array_2.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X356 VREF d<5> hgu_cdac_8bit_array_3.drv<31:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X357 hgu_cdac_8bit_array_3.drv<31:0> d<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X358 hgu_cdac_8bit_array_3.drv<0> d<0> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.35
X359 VREF db<4> hgu_cdac_8bit_array_2.drv<15:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X360 VREF d<6> hgu_cdac_8bit_array_3.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X361 VREF d<6> hgu_cdac_8bit_array_3.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X362 hgu_cdac_8bit_array_3.drv<63:0> d<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X363 VSS db<6> hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X364 hgu_cdac_8bit_array_2.drv<31:0> db<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X365 VREF db<6> hgu_cdac_8bit_array_2.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X366 hgu_cdac_8bit_array_3.drv<63:0> d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X367 hgu_cdac_8bit_array_3.drv<31:0> d<5> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X368 hgu_cdac_8bit_array_2.drv<15:0> db<4> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X369 hgu_cdac_8bit_array_3.drv<63:0> d<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X370 hgu_cdac_8bit_array_3.drv<15:0> d<4> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X371 VREF d<5> hgu_cdac_8bit_array_3.drv<31:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X372 VREF db<6> hgu_cdac_8bit_array_2.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X373 VSS d<5> hgu_cdac_8bit_array_3.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X374 hgu_cdac_8bit_array_2.drv<31:0> db<5> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X375 hgu_cdac_8bit_array_2.drv<63:0> db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X376 hgu_cdac_8bit_array_2.drv<63:0> db<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X377 VSS d<6> hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X378 VREF d<4> hgu_cdac_8bit_array_3.drv<15:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X379 VSS d<6> hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X380 VSS d<4> hgu_cdac_8bit_array_3.drv<15:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X381 VREF d<3> hgu_cdac_8bit_array_3.drv<7:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.35
X382 hgu_cdac_8bit_array_3.drv<31:0> d<5> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X383 hgu_cdac_8bit_array_3.drv<63:0> d<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X384 VSS db<6> hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X385 hgu_cdac_8bit_array_2.drv<31:0> db<5> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X386 hgu_cdac_8bit_array_2.drv<63:0> db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X387 VSS d<5> hgu_cdac_8bit_array_3.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X388 hgu_cdac_8bit_array_2.drv<63:0> db<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X389 hgu_cdac_8bit_array_3.drv<63:0> d<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X390 VSS db<5> hgu_cdac_8bit_array_2.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X391 VSS d<6> hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X392 VSS d<6> hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X393 hgu_cdac_8bit_array_2.drv<7:0> db<3> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.122 ps=1.42 w=0.42 l=0.35
X394 VSS db<2> hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X395 VREF db<1> hgu_cdac_8bit_array_2.drv<1:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.35
X396 hgu_cdac_8bit_array_3.drv<15:0> d<4> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.35
X397 VREF d<3> hgu_cdac_8bit_array_3.drv<7:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X398 VSS db<5> hgu_cdac_8bit_array_2.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X399 VSS db<6> hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X400 VREF db<3> hgu_cdac_8bit_array_2.drv<7:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X401 VSS d<2> hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X402 VSS db<6> hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X403 VREF db<5> hgu_cdac_8bit_array_2.drv<31:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X404 hgu_cdac_8bit_array_3.drv<63:0> d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X405 VSS d<5> hgu_cdac_8bit_array_3.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X406 hgu_cdac_8bit_array_2.drv<31:0> db<5> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X407 hgu_cdac_8bit_array_3.drv<63:0> d<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X408 VSS d<5> hgu_cdac_8bit_array_3.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X409 hgu_cdac_8bit_array_3.drv<1:0> d<1> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.35
X410 VREF db<4> hgu_cdac_8bit_array_2.drv<15:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.35
X411 VREF d<5> hgu_cdac_8bit_array_3.drv<31:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X412 VSS db<6> hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X413 VREF d<6> hgu_cdac_8bit_array_3.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X414 VREF db<6> hgu_cdac_8bit_array_2.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X415 hgu_cdac_8bit_array_3.drv<63:0> d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X416 hgu_cdac_8bit_array_2.drv<63:0> db<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X417 hgu_cdac_8bit_array_2.drv<15:0> db<4> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X418 hgu_cdac_8bit_array_3.drv<63:0> d<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X419 VREF db<6> hgu_cdac_8bit_array_2.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X420 hgu_cdac_8bit_array_2.drv<31:0> db<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X421 hgu_cdac_8bit_array_3.drv<63:0> d<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X422 hgu_cdac_8bit_array_3.drv<7:0> d<3> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.35
X423 VSS db<4> hgu_cdac_8bit_array_2.drv<15:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X424 hgu_cdac_8bit_array_2.drv<63:0> db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X425 hgu_cdac_8bit_array_3.drv<0> d<0> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.244 ps=2.26 w=0.84 l=0.35
X426 hgu_cdac_8bit_array_3.drv<31:0> d<5> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X427 hgu_cdac_8bit_array_2.drv<63:0> db<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.35
X428 VSS db<6> hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X429 VREF db<6> hgu_cdac_8bit_array_2.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X430 hgu_cdac_8bit_array_2.drv<31:0> db<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.122 ps=1.42 w=0.42 l=0.35
X431 hgu_cdac_8bit_array_3.drv<63:0> d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.122 ps=1.42 w=0.42 l=0.35
X432 hgu_cdac_8bit_array_2.drv<31:0> db<5> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X433 hgu_cdac_8bit_array_2.drv<63:0> db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X434 VSS d<5> hgu_cdac_8bit_array_3.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.35
X435 hgu_cdac_8bit_array_3.drv<63:0> d<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X436 VSS db<6> hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X437 VSS db<4> hgu_cdac_8bit_array_2.drv<15:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X438 hgu_cdac_8bit_array_3.drv<63:0> d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X439 hgu_cdac_8bit_array_3.drv<15:0> d<4> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X440 hgu_cdac_8bit_array_2.drv<63:0> db<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X441 VREF d<5> hgu_cdac_8bit_array_3.drv<31:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X442 hgu_cdac_8bit_array_2.drv<63:0> db<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X443 VSS d<6> hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X444 VREF db<5> hgu_cdac_8bit_array_2.drv<31:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X445 VSS db<6> hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X446 VREF db<4> hgu_cdac_8bit_array_2.drv<15:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X447 VREF d<6> hgu_cdac_8bit_array_3.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X448 VSS db<3> hgu_cdac_8bit_array_2.drv<7:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X449 VSS d<5> hgu_cdac_8bit_array_3.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X450 hgu_cdac_8bit_array_3.drv<31:0> d<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X451 VSS db<6> hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X452 VREF d<4> hgu_cdac_8bit_array_3.drv<15:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X453 VREF d<6> hgu_cdac_8bit_array_3.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X454 hgu_cdac_8bit_array_3.drv<63:0> d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X455 VSS db<5> hgu_cdac_8bit_array_2.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.35
X456 hgu_cdac_8bit_array_2.drv<63:0> db<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X457 VSS d<6> hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X458 VREF d<5> hgu_cdac_8bit_array_3.drv<31:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X459 VSS db<6> hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X460 VREF db<4> hgu_cdac_8bit_array_2.drv<15:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X461 VREF d<6> hgu_cdac_8bit_array_3.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X462 VREF d<6> hgu_cdac_8bit_array_3.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X463 hgu_cdac_8bit_array_2.drv<63:0> db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X464 hgu_cdac_8bit_array_3.drv<63:0> d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X465 hgu_cdac_8bit_array_3.drv<31:0> d<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X466 VREF db<6> hgu_cdac_8bit_array_2.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X467 hgu_cdac_8bit_array_3.drv<63:0> d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X468 VREF d<2> hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X469 hgu_cdac_8bit_array_2.drv<31:0> db<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X470 hgu_cdac_8bit_array_2.drv<15:0> db<4> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X471 hgu_cdac_8bit_array_3.drv<63:0> d<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X472 hgu_cdac_8bit_array_3.drv<15:0> d<4> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X473 VREF d<5> hgu_cdac_8bit_array_3.drv<31:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X474 hgu_cdac_8bit_array_2.drv<63:0> db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X475 VSS d<5> hgu_cdac_8bit_array_3.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X476 hgu_cdac_8bit_array_2.drv<63:0> db<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X477 VREF d<5> hgu_cdac_8bit_array_3.drv<31:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X478 hgu_cdac_8bit_array_3.drv<31:0> d<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X479 VREF db<6> hgu_cdac_8bit_array_2.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X480 hgu_cdac_8bit_array_2.drv<31:0> db<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X481 hgu_cdac_8bit_array_3.drv<63:0> d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X482 VSS db<5> hgu_cdac_8bit_array_2.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X483 hgu_cdac_8bit_array_2.drv<15:0> db<4> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X484 hgu_cdac_8bit_array_2.drv<63:0> db<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X485 VSS db<6> hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X486 hgu_cdac_8bit_array_3.drv<63:0> d<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X487 hgu_cdac_8bit_array_3.drv<15:0> d<4> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X488 hgu_cdac_8bit_array_2.drv<31:0> db<5> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X489 hgu_cdac_8bit_array_2.drv<63:0> db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X490 hgu_cdac_8bit_array_2.drv<63:0> db<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X491 VSS d<6> hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X492 VSS d<6> hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X493 VSS db<6> hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X494 hgu_cdac_8bit_array_3.drv<63:0> d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X495 VREF db<6> hgu_cdac_8bit_array_2.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X496 hgu_cdac_8bit_array_2.drv<63:0> db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X497 hgu_cdac_8bit_array_2.drv<31:0> db<5> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X498 hgu_cdac_8bit_array_3.drv<63:0> d<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.35
X499 VSS d<6> hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X500 VREF db<6> hgu_cdac_8bit_array_2.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X501 VREF d<5> hgu_cdac_8bit_array_3.drv<31:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.35
X502 hgu_cdac_8bit_array_2.drv<63:0> db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X503 hgu_cdac_8bit_array_3.drv<63:0> d<6> VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X504 VSS db<5> hgu_cdac_8bit_array_2.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X505 VREF d<6> hgu_cdac_8bit_array_3.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X506 VREF db<6> hgu_cdac_8bit_array_2.drv<63:0> VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X507 hgu_cdac_8bit_array_3.drv<63:0> d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
.ends

