magic
tech sky130A
timestamp 1698381494
use hgu_cdac_unit  x1[0]
timestamp 1698381206
transform 1 0 0 0 1 1100
box 343 299 679 912
use hgu_cdac_unit  x1[1]
timestamp 1698381206
transform 1 0 0 0 1 1679
box 343 299 679 912
use hgu_cdac_unit  x1[2]
timestamp 1698381206
transform 1 0 303 0 1 1100
box 343 299 679 912
use hgu_cdac_unit  x1[3]
timestamp 1698381206
transform 1 0 303 0 1 1679
box 343 299 679 912
<< end >>
