magic
tech sky130A
magscale 1 2
timestamp 1698742797
<< nwell >>
rect 379 440 684 824
<< nmos >>
rect 516 262 546 346
<< pmos >>
rect 516 478 546 646
<< ndiff >>
rect 458 334 516 346
rect 458 274 470 334
rect 504 274 516 334
rect 458 262 516 274
rect 546 334 604 346
rect 546 274 558 334
rect 592 274 604 334
rect 546 262 604 274
<< pdiff >>
rect 458 634 516 646
rect 458 581 470 634
rect 504 581 516 634
rect 458 543 516 581
rect 458 490 470 543
rect 504 490 516 543
rect 458 478 516 490
rect 546 634 604 646
rect 546 581 558 634
rect 592 581 604 634
rect 546 543 604 581
rect 546 490 558 543
rect 592 490 604 543
rect 546 478 604 490
<< ndiffc >>
rect 470 274 504 334
rect 558 274 592 334
<< pdiffc >>
rect 470 581 504 634
rect 470 490 504 543
rect 558 581 592 634
rect 558 490 592 543
<< psubdiff >>
rect 415 204 648 208
rect 415 166 468 204
rect 506 166 556 204
rect 594 166 648 204
rect 415 162 648 166
<< nsubdiff >>
rect 415 784 648 788
rect 415 746 468 784
rect 506 746 556 784
rect 594 746 648 784
rect 415 742 648 746
<< psubdiffcont >>
rect 468 166 506 204
rect 556 166 594 204
<< nsubdiffcont >>
rect 468 746 506 784
rect 556 746 594 784
<< poly >>
rect 516 646 546 677
rect 516 435 546 478
rect 454 419 546 435
rect 454 385 470 419
rect 504 385 546 419
rect 454 369 546 385
rect 516 346 546 369
rect 516 236 546 262
<< polycont >>
rect 470 385 504 419
<< locali >>
rect 415 784 648 788
rect 415 746 468 784
rect 506 746 556 784
rect 594 746 648 784
rect 415 742 648 746
rect 470 634 504 650
rect 470 543 504 581
rect 470 474 504 490
rect 558 634 592 650
rect 558 543 592 581
rect 454 385 470 419
rect 504 385 520 419
rect 470 334 504 350
rect 470 208 504 274
rect 558 334 592 490
rect 558 258 592 274
rect 415 204 648 208
rect 415 166 468 204
rect 506 166 556 204
rect 594 166 648 204
rect 415 162 648 166
<< viali >>
rect 468 746 506 784
rect 556 746 594 784
rect 470 581 504 634
rect 470 490 504 543
rect 558 581 592 634
rect 558 490 592 543
rect 470 385 504 419
rect 470 274 504 334
rect 558 274 592 334
rect 468 166 506 204
rect 556 166 594 204
<< metal1 >>
rect 415 784 648 790
rect 415 746 468 784
rect 506 746 556 784
rect 594 746 648 784
rect 415 740 648 746
rect 415 679 648 711
rect 470 646 504 679
rect 464 634 510 646
rect 464 581 470 634
rect 504 581 510 634
rect 464 543 510 581
rect 464 490 470 543
rect 504 490 510 543
rect 464 478 510 490
rect 552 634 598 646
rect 552 581 558 634
rect 592 581 598 634
rect 552 543 598 581
rect 552 490 558 543
rect 592 490 598 543
rect 552 478 598 490
rect 454 419 520 429
rect 454 385 470 419
rect 504 385 520 419
rect 454 375 520 385
rect 464 334 510 346
rect 464 274 470 334
rect 504 274 510 334
rect 464 262 510 274
rect 552 334 598 346
rect 552 274 558 334
rect 592 274 598 334
rect 552 262 598 274
rect 415 204 648 210
rect 415 166 468 204
rect 506 166 556 204
rect 594 166 648 204
rect 415 160 648 166
<< labels >>
flabel locali 566 388 586 424 0 FreeSans 160 0 0 0 OUT
port 15 nsew
flabel metal1 429 689 456 704 0 FreeSans 160 0 0 0 VREF
port 19 nsew
flabel metal1 422 749 457 774 0 FreeSans 160 0 0 0 VDD
port 22 nsew
flabel metal1 426 174 460 196 0 FreeSans 160 0 0 0 VSS
port 24 nsew
flabel metal1 470 385 504 419 0 FreeSans 160 0 0 0 IN
port 26 nsew
<< end >>
