magic
tech sky130A
magscale 1 2
timestamp 1697025759
<< error_p >>
rect -29 161 29 167
rect -29 127 -17 161
rect -29 121 29 127
rect -29 -127 29 -121
rect -29 -161 -17 -127
rect -29 -167 29 -161
<< nwell >>
rect -211 -299 211 299
<< pmos >>
rect -15 -80 15 80
<< pdiff >>
rect -73 68 -15 80
rect -73 -68 -61 68
rect -27 -68 -15 68
rect -73 -80 -15 -68
rect 15 68 73 80
rect 15 -68 27 68
rect 61 -68 73 68
rect 15 -80 73 -68
<< pdiffc >>
rect -61 -68 -27 68
rect 27 -68 61 68
<< nsubdiff >>
rect -175 229 -79 263
rect 79 229 175 263
rect -175 167 -141 229
rect 141 167 175 229
rect -175 -229 -141 -167
rect 141 -229 175 -167
rect -175 -263 -79 -229
rect 79 -263 175 -229
<< nsubdiffcont >>
rect -79 229 79 263
rect -175 -167 -141 167
rect 141 -167 175 167
rect -79 -263 79 -229
<< poly >>
rect -33 161 33 177
rect -33 127 -17 161
rect 17 127 33 161
rect -33 111 33 127
rect -15 80 15 111
rect -15 -111 15 -80
rect -33 -127 33 -111
rect -33 -161 -17 -127
rect 17 -161 33 -127
rect -33 -177 33 -161
<< polycont >>
rect -17 127 17 161
rect -17 -161 17 -127
<< locali >>
rect -175 229 -79 263
rect 79 229 175 263
rect -175 167 -141 229
rect 141 167 175 229
rect -33 127 -17 161
rect 17 127 33 161
rect -61 68 -27 84
rect -61 -84 -27 -68
rect 27 68 61 84
rect 27 -84 61 -68
rect -33 -161 -17 -127
rect 17 -161 33 -127
rect -175 -229 -141 -167
rect 141 -229 175 -167
rect -175 -263 -79 -229
rect 79 -263 175 -229
<< viali >>
rect -17 127 17 161
rect -61 -68 -27 68
rect 27 -68 61 68
rect -17 -161 17 -127
<< metal1 >>
rect -29 161 29 167
rect -29 127 -17 161
rect 17 127 29 161
rect -29 121 29 127
rect -67 68 -21 80
rect -67 -68 -61 68
rect -27 -68 -21 68
rect -67 -80 -21 -68
rect 21 68 67 80
rect 21 -68 27 68
rect 61 -68 67 68
rect 21 -80 67 -68
rect -29 -127 29 -121
rect -29 -161 -17 -127
rect 17 -161 29 -127
rect -29 -167 29 -161
<< properties >>
string FIXED_BBOX -158 -246 158 246
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.8 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
