magic
tech sky130A
magscale 1 2
timestamp 1700647327
<< nwell >>
rect -98 1296 408 2272
<< pwell >>
rect -176 -206 498 1048
<< psubdiff >>
rect -135 944 -31 979
rect -135 910 -104 944
rect -70 910 -31 944
rect -135 882 -31 910
rect 329 876 433 911
rect 329 842 360 876
rect 394 842 433 876
rect 329 814 433 842
rect -151 738 -47 773
rect -151 704 -120 738
rect -86 704 -47 738
rect -151 676 -47 704
rect 321 724 425 759
rect 321 690 352 724
rect 386 690 425 724
rect 321 662 425 690
rect -147 546 -43 581
rect -147 512 -116 546
rect -82 512 -43 546
rect -147 484 -43 512
rect 329 534 433 569
rect 329 500 360 534
rect 394 500 433 534
rect 329 472 433 500
rect -129 390 -25 425
rect -129 356 -98 390
rect -64 356 -25 390
rect -129 328 -25 356
rect 345 382 449 417
rect 345 348 376 382
rect 410 348 449 382
rect 345 320 449 348
rect -131 236 -27 271
rect -131 202 -100 236
rect -66 202 -27 236
rect -131 174 -27 202
rect -133 60 -29 95
rect -133 26 -102 60
rect -68 26 -29 60
rect -133 -2 -29 26
rect 333 46 437 81
rect 333 12 364 46
rect 398 12 437 46
rect 333 -16 437 12
rect -115 -104 -11 -69
rect -115 -138 -84 -104
rect -50 -138 -11 -104
rect -115 -166 -11 -138
rect 111 -104 215 -69
rect 111 -138 142 -104
rect 176 -138 215 -104
rect 111 -166 215 -138
rect 323 -110 427 -75
rect 323 -144 354 -110
rect 388 -144 427 -110
rect 323 -172 427 -144
<< nsubdiff >>
rect 276 2203 359 2228
rect 276 2168 301 2203
rect 335 2168 359 2203
rect -60 2139 23 2164
rect 276 2144 359 2168
rect -60 2104 -35 2139
rect -1 2104 23 2139
rect -60 2080 23 2104
rect 288 2065 371 2090
rect 288 2030 313 2065
rect 347 2030 371 2065
rect -54 1983 29 2008
rect 288 2006 371 2030
rect -54 1948 -29 1983
rect 5 1948 29 1983
rect -54 1924 29 1948
rect -54 1799 29 1824
rect -54 1764 -29 1799
rect 5 1764 29 1799
rect -54 1740 29 1764
rect 284 1769 367 1794
rect 284 1734 309 1769
rect 343 1734 367 1769
rect 284 1710 367 1734
rect -58 1653 25 1678
rect -58 1618 -33 1653
rect 1 1618 25 1653
rect -58 1594 25 1618
rect 286 1623 369 1648
rect 286 1588 311 1623
rect 345 1588 369 1623
rect 286 1564 369 1588
rect -54 1471 29 1496
rect -54 1436 -29 1471
rect 5 1436 29 1471
rect -54 1412 29 1436
rect 286 1471 369 1496
rect 286 1436 311 1471
rect 345 1436 369 1471
rect 286 1412 369 1436
<< psubdiffcont >>
rect -104 910 -70 944
rect 360 842 394 876
rect -120 704 -86 738
rect 352 690 386 724
rect -116 512 -82 546
rect 360 500 394 534
rect -98 356 -64 390
rect 376 348 410 382
rect -100 202 -66 236
rect -102 26 -68 60
rect 364 12 398 46
rect -84 -138 -50 -104
rect 142 -138 176 -104
rect 354 -144 388 -110
<< nsubdiffcont >>
rect 301 2168 335 2203
rect -35 2104 -1 2139
rect 313 2030 347 2065
rect -29 1948 5 1983
rect -29 1764 5 1799
rect 309 1734 343 1769
rect -33 1618 1 1653
rect 311 1588 345 1623
rect -29 1436 5 1471
rect 311 1436 345 1471
<< poly >>
rect 124 1098 190 1222
<< locali >>
rect -18 2256 32 2258
rect 298 2256 348 2258
rect -18 2248 356 2256
rect -18 2228 358 2248
rect -18 2210 359 2228
rect -18 2164 32 2210
rect -60 2139 32 2164
rect 276 2203 359 2210
rect 276 2168 301 2203
rect 335 2168 359 2203
rect 276 2144 359 2168
rect -60 2104 -35 2139
rect -1 2104 32 2139
rect -60 2080 32 2104
rect 292 2090 358 2144
rect -18 2008 32 2080
rect 288 2065 371 2090
rect 288 2030 313 2065
rect 347 2030 371 2065
rect -54 1983 29 2008
rect 288 2006 371 2030
rect -54 1948 -29 1983
rect 5 1948 29 1983
rect -54 1924 29 1948
rect -18 1824 32 1924
rect 96 1912 130 1996
rect -54 1799 29 1824
rect -54 1764 -29 1799
rect 5 1764 29 1799
rect 184 1796 218 1880
rect 298 1794 348 2006
rect -54 1740 29 1764
rect 284 1769 367 1794
rect -18 1678 32 1740
rect -58 1653 32 1678
rect 96 1656 130 1740
rect 284 1734 309 1769
rect 343 1734 367 1769
rect 284 1710 367 1734
rect -58 1618 -33 1653
rect 1 1618 32 1653
rect 298 1648 348 1710
rect -58 1594 32 1618
rect 286 1623 369 1648
rect -18 1496 32 1594
rect 184 1510 218 1594
rect 286 1588 311 1623
rect 345 1588 369 1623
rect 286 1564 369 1588
rect 298 1496 348 1564
rect -54 1471 32 1496
rect -54 1436 -29 1471
rect 5 1436 32 1471
rect 286 1471 369 1496
rect -54 1412 32 1436
rect -18 1302 32 1412
rect 96 1362 130 1446
rect 286 1436 311 1471
rect 345 1436 369 1471
rect 286 1412 369 1436
rect 298 1302 348 1412
rect 116 1126 162 1144
rect 116 1092 122 1126
rect 156 1092 162 1126
rect 116 1080 162 1092
rect -94 980 -44 1062
rect -114 979 -44 980
rect -136 944 -31 979
rect -136 910 -104 944
rect -70 910 -31 944
rect 42 928 76 1012
rect 340 912 390 1044
rect 340 911 400 912
rect -136 882 -31 910
rect -94 774 -44 882
rect 202 794 236 878
rect 328 876 433 911
rect 328 842 360 876
rect 394 842 433 876
rect 328 814 433 842
rect -130 773 -44 774
rect -152 738 -44 773
rect 340 760 390 814
rect 340 759 392 760
rect -152 704 -120 738
rect -86 704 -44 738
rect -152 676 -44 704
rect -94 582 -44 676
rect 42 658 76 742
rect 320 724 425 759
rect 320 690 352 724
rect 386 690 425 724
rect 320 662 425 690
rect -126 581 -44 582
rect -148 546 -43 581
rect -148 512 -116 546
rect -82 512 -43 546
rect 202 520 236 604
rect 340 570 390 662
rect 340 569 400 570
rect 328 534 433 569
rect -148 484 -43 512
rect 328 500 360 534
rect 394 500 433 534
rect -94 426 -44 484
rect 328 472 433 500
rect -108 425 -44 426
rect -130 390 -25 425
rect -130 356 -98 390
rect -64 356 -25 390
rect 42 382 76 466
rect 340 418 390 472
rect 340 417 416 418
rect 340 382 449 417
rect -130 328 -25 356
rect 340 348 376 382
rect 410 348 449 382
rect -94 272 -44 328
rect -110 271 -44 272
rect -132 236 -27 271
rect 202 242 236 326
rect 340 320 449 348
rect -132 202 -100 236
rect -66 202 -27 236
rect -132 174 -27 202
rect -94 96 -44 174
rect 42 106 76 190
rect -112 95 -44 96
rect -134 60 -29 95
rect 340 88 390 320
rect 348 82 384 88
rect 348 81 404 82
rect -134 26 -102 60
rect -68 26 -29 60
rect 332 46 437 81
rect 332 44 364 46
rect -134 -2 -29 26
rect 324 12 364 44
rect 398 12 437 46
rect -94 -69 -44 -2
rect 324 -16 437 12
rect 132 -69 182 -68
rect -116 -88 -11 -69
rect 110 -88 215 -69
rect 324 -75 410 -16
rect 322 -88 427 -75
rect -116 -104 427 -88
rect -116 -138 -84 -104
rect -50 -132 142 -104
rect -50 -138 -11 -132
rect -116 -166 -11 -138
rect 110 -138 142 -132
rect 176 -110 427 -104
rect 176 -132 354 -110
rect 176 -138 215 -132
rect 110 -166 215 -138
rect 322 -144 354 -132
rect 388 -144 427 -110
rect 322 -172 427 -144
<< viali >>
rect 122 1092 156 1126
<< metal1 >>
rect 158 2140 252 2190
rect 178 2078 224 2140
rect 184 1796 218 1880
rect 96 1656 130 1740
rect 184 1510 218 1594
rect 96 1362 130 1446
rect 180 1334 528 1336
rect 180 1312 548 1334
rect 178 1294 548 1312
rect 280 1292 548 1294
rect -62 1172 -6 1192
rect 116 1172 160 1260
rect 502 1208 548 1292
rect 594 1208 688 1226
rect 502 1174 688 1208
rect -62 1126 186 1172
rect -62 1104 -6 1126
rect 116 1092 122 1126
rect 156 1092 162 1126
rect 502 1096 548 1174
rect 594 1136 688 1174
rect 116 1080 162 1092
rect 196 1054 548 1096
rect 196 1052 544 1054
rect 196 -10 242 34
rect 182 -60 264 -10
use hgu_nfet_hvt_stack_in_delay  hgu_nfet_hvt_stack_in_delay_0
timestamp 1699184006
transform -1 0 333 0 1 235
box -90 -235 303 886
use hgu_pfet_hvt_stack_in_delay  hgu_pfet_hvt_stack_in_delay_0
timestamp 1699184006
transform -1 0 315 0 -1 2157
box -98 40 268 947
<< labels >>
flabel metal1 182 -60 264 -10 0 FreeSans 320 0 0 0 vss
port 1 nsew
flabel metal1 -62 1104 -6 1192 0 FreeSans 320 0 0 0 input
port 2 nsew
flabel metal1 158 2140 252 2190 0 FreeSans 320 0 0 0 vdd
port 0 nsew
flabel metal1 594 1136 688 1226 0 FreeSans 320 0 0 0 output
port 4 nsew
<< end >>
