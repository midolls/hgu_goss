magic
tech sky130A
timestamp 1698619350
<< end >>
