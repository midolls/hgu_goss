magic
tech sky130A
timestamp 1697519636
<< checkpaint >>
rect -630 -1030 730 730
<< metal1 >>
rect 0 0 100 100
rect 0 -200 100 -100
rect 0 -400 100 -300
<< labels >>
flabel metal1 0 0 100 100 0 FreeSans 128 0 0 0 C0
port 0 nsew
flabel metal1 0 -200 100 -100 0 FreeSans 128 0 0 0 C1
port 1 nsew
flabel metal1 0 -400 100 -300 0 FreeSans 128 0 0 0 SUB
port 2 nsew
<< end >>
