magic
tech sky130A
magscale 1 2
timestamp 1698286991
use inv_2_test  inv_2_test_0
timestamp 1698286991
transform 1 0 -591 0 1 -1036
box 425 2360 831 3025
use inv_2_test  inv_2_test_1
timestamp 1698286991
transform 1 0 -767 0 1 -1036
box 425 2360 831 3025
<< end >>
