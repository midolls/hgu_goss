magic
tech sky130A
magscale 1 2
timestamp 1698671623
<< error_s >>
rect 10671 4108 10729 4114
rect 10671 4074 10683 4108
rect 10671 4068 10729 4074
rect 10671 3896 10729 3902
rect 10671 3862 10683 3896
rect 10671 3856 10729 3862
rect 11161 3724 11165 4246
rect 11343 4108 11401 4114
rect 11343 4074 11355 4108
rect 11343 4068 11401 4074
rect 11343 3896 11401 3902
rect 11343 3862 11355 3896
rect 11343 3856 11401 3862
rect 11833 3724 11837 4246
rect 12015 4108 12073 4114
rect 12015 4074 12027 4108
rect 12015 4068 12073 4074
rect 12015 3896 12073 3902
rect 12015 3862 12027 3896
rect 12015 3856 12073 3862
rect 12505 3724 12509 4246
rect 12687 4108 12745 4114
rect 12687 4074 12699 4108
rect 12687 4068 12745 4074
rect 12687 3896 12745 3902
rect 12687 3862 12699 3896
rect 12687 3856 12745 3862
rect 13177 3724 13181 4246
rect 13359 4108 13417 4114
rect 13359 4074 13371 4108
rect 13359 4068 13417 4074
rect 13359 3896 13417 3902
rect 13359 3862 13371 3896
rect 13359 3856 13417 3862
rect 13849 3724 13853 4246
rect 14031 4108 14089 4114
rect 14031 4074 14043 4108
rect 14031 4068 14089 4074
rect 14031 3896 14089 3902
rect 14031 3862 14043 3896
rect 14031 3856 14089 3862
rect 14521 3724 14525 4246
rect 14703 4108 14761 4114
rect 14703 4074 14715 4108
rect 14703 4068 14761 4074
rect 14703 3896 14761 3902
rect 14703 3862 14715 3896
rect 14703 3856 14761 3862
rect 15193 3724 15197 4246
rect 15375 4108 15433 4114
rect 15375 4074 15387 4108
rect 15375 4068 15433 4074
rect 15375 3896 15433 3902
rect 15375 3862 15387 3896
rect 15375 3856 15433 3862
rect 11051 3443 11065 3507
rect 11723 3443 11737 3507
rect 12395 3443 12409 3507
rect 13067 3443 13081 3507
rect 13739 3443 13753 3507
rect 14411 3443 14425 3507
rect 15083 3443 15097 3507
rect 11051 3363 11065 3427
rect 11723 3363 11737 3427
rect 12395 3363 12409 3427
rect 13067 3363 13081 3427
rect 13739 3363 13753 3427
rect 14411 3363 14425 3427
rect 15083 3363 15097 3427
rect 11051 3283 11065 3347
rect 11723 3283 11737 3347
rect 12395 3283 12409 3347
rect 13067 3283 13081 3347
rect 13739 3283 13753 3347
rect 14411 3283 14425 3347
rect 15083 3283 15097 3347
rect 11051 3203 11065 3267
rect 11723 3203 11737 3267
rect 12395 3203 12409 3267
rect 13067 3203 13081 3267
rect 13739 3203 13753 3267
rect 14411 3203 14425 3267
rect 15083 3203 15097 3267
rect 11051 3123 11065 3187
rect 11723 3123 11737 3187
rect 12395 3123 12409 3187
rect 13067 3123 13081 3187
rect 13739 3123 13753 3187
rect 14411 3123 14425 3187
rect 15083 3123 15097 3187
rect 11051 3043 11065 3107
rect 11723 3043 11737 3107
rect 12395 3043 12409 3107
rect 13067 3043 13081 3107
rect 13739 3043 13753 3107
rect 14411 3043 14425 3107
rect 15083 3043 15097 3107
rect 11051 2963 11065 3027
rect 11723 2963 11737 3027
rect 12395 2963 12409 3027
rect 13067 2963 13081 3027
rect 13739 2963 13753 3027
rect 14411 2963 14425 3027
rect 15083 2963 15097 3027
rect 11051 2883 11065 2947
rect 11723 2883 11737 2947
rect 12395 2883 12409 2947
rect 13067 2883 13081 2947
rect 13739 2883 13753 2947
rect 14411 2883 14425 2947
rect 15083 2883 15097 2947
rect 11051 2803 11065 2867
rect 11723 2803 11737 2867
rect 12395 2803 12409 2867
rect 13067 2803 13081 2867
rect 13739 2803 13753 2867
rect 14411 2803 14425 2867
rect 15083 2803 15097 2867
rect 11051 2723 11065 2787
rect 11723 2723 11737 2787
rect 12395 2723 12409 2787
rect 13067 2723 13081 2787
rect 13739 2723 13753 2787
rect 14411 2723 14425 2787
rect 15083 2723 15097 2787
rect 10637 2068 11059 2394
rect 11243 2068 11665 2394
rect 11849 2068 12271 2394
rect 12455 2068 12877 2394
rect 13187 2068 13609 2394
rect 13793 2068 14215 2394
rect 14525 2068 14947 2394
rect 10637 2024 10746 2068
rect 10819 2062 10877 2068
rect 10819 2028 10831 2062
rect 10608 2014 10666 2020
rect 10673 2014 10704 2024
rect 10819 2022 10877 2028
rect 10608 1980 10620 2014
rect 10639 1990 10704 2014
rect 11035 2007 11059 2068
rect 11425 2062 11483 2068
rect 11425 2028 11437 2062
rect 11425 2022 11483 2028
rect 11641 2007 11665 2068
rect 12031 2062 12089 2068
rect 12031 2028 12043 2062
rect 12031 2022 12089 2028
rect 12247 2007 12271 2068
rect 12637 2062 12695 2068
rect 12637 2028 12649 2062
rect 12637 2022 12695 2028
rect 12853 2007 12877 2068
rect 13369 2062 13427 2068
rect 13369 2028 13381 2062
rect 13369 2022 13427 2028
rect 13459 2007 13609 2068
rect 13975 2062 14033 2068
rect 13975 2028 13987 2062
rect 13975 2022 14033 2028
rect 14065 2007 14215 2068
rect 14671 2007 14855 2068
rect 10673 1980 10701 1990
rect 10608 1974 10666 1980
rect 10673 1956 10697 1980
rect 10671 1928 10697 1956
rect 10673 1926 10701 1928
<< nwell >>
rect 10637 2195 11059 2394
rect 10644 2192 11059 2195
rect 10746 2068 11059 2192
rect 11243 2068 11665 2394
rect 11849 2068 12271 2394
rect 12455 2068 12877 2394
rect 13187 2068 13609 2394
rect 13793 2068 14215 2394
rect 14525 2068 14947 2394
rect 11035 2007 11059 2068
rect 11641 2007 11665 2068
rect 12247 2007 12271 2068
rect 12853 2007 12877 2068
rect 13459 2007 13609 2068
rect 14065 2007 14215 2068
rect 14671 2007 14855 2068
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
rect 0 -2400 200 -2200
rect 0 -2800 200 -2600
use hgu_sw_cap  x2
timestamp 1698575955
transform -1 0 11543 0 1 154
box 369 547 1041 2240
use hgu_pfet_hvt_stack_in_delay  x3
timestamp 1698575910
transform 1 0 10303 0 1 1295
box 49 669 443 910
use hgu_sw_cap  x3[0]
timestamp 1698575955
transform -1 0 12755 0 1 154
box 369 547 1041 2240
use hgu_sw_cap  x3[1]
timestamp 1698575955
transform -1 0 12149 0 1 154
box 369 547 1041 2240
use hgu_nfet_hvt_stack_in_delay  x4
timestamp 1698575851
transform 1 0 9863 0 1 1085
box 85 693 838 905
use hgu_sw_cap  x4[0]
timestamp 1698575955
transform -1 0 15431 0 1 154
box 369 547 1041 2240
use hgu_sw_cap  x4[1]
timestamp 1698575955
transform -1 0 14699 0 1 154
box 369 547 1041 2240
use hgu_sw_cap  x4[2]
timestamp 1698575955
transform -1 0 14093 0 1 154
box 369 547 1041 2240
use hgu_sw_cap  x4[3]
timestamp 1698575955
transform -1 0 13361 0 1 154
box 369 547 1041 2240
use hgu_sw_cap_pmos  x5[0]
timestamp 1698575999
transform 1 0 14713 0 1 1954
box 369 547 1041 2292
use hgu_sw_cap_pmos  x5[1]
timestamp 1698575999
transform 1 0 14041 0 1 1954
box 369 547 1041 2292
use hgu_sw_cap_pmos  x5[2]
timestamp 1698575999
transform 1 0 13369 0 1 1954
box 369 547 1041 2292
use hgu_sw_cap_pmos  x5[3]
timestamp 1698575999
transform 1 0 12697 0 1 1954
box 369 547 1041 2292
use hgu_sw_cap_pmos  x5[4]
timestamp 1698575999
transform 1 0 12025 0 1 1954
box 369 547 1041 2292
use hgu_sw_cap_pmos  x5[5]
timestamp 1698575999
transform 1 0 11353 0 1 1954
box 369 547 1041 2292
use hgu_sw_cap_pmos  x5[6]
timestamp 1698575999
transform 1 0 10681 0 1 1954
box 369 547 1041 2292
use hgu_sw_cap_pmos  x5[7]
timestamp 1698575999
transform 1 0 10009 0 1 1954
box 369 547 1041 2292
use sky130_fd_pr__nfet_01v8_ZPNSVB  XM13
timestamp 1698581447
transform -1 0 15671 0 -1 1651
box -73 -106 73 107
use sky130_fd_pr__nfet_01v8_ZPNSVB  XM15
timestamp 1698581447
transform -1 0 15583 0 -1 1651
box -73 -106 73 107
use sky130_fd_pr__pfet_01v8_hvt_M479BZ  XM46
timestamp 1698581447
transform -1 0 15671 0 -1 2300
box -109 -78 110 90
use sky130_fd_pr__pfet_01v8_hvt_M479BZ  XM47
timestamp 1698581447
transform -1 0 15583 0 -1 2300
box -109 -78 110 90
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 128 0 0 0 IN
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 128 0 0 0 VDD
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 128 0 0 0 VSS
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 128 0 0 0 OUT
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 128 0 0 0 {code\[0\]}
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 128 0 0 0 {code\[1\]}
port 5 nsew
flabel metal1 0 -2400 200 -2200 0 FreeSans 128 0 0 0 {code\[2\]}
port 6 nsew
flabel metal1 0 -2800 200 -2600 0 FreeSans 128 0 0 0 {code\[3\]}
port 7 nsew
<< end >>
