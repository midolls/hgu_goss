magic
tech sky130A
magscale 1 2
timestamp 1698625662
<< pwell >>
rect 32592 4404 32618 4436
rect 33198 4404 33224 4436
rect 33804 4404 33830 4436
rect 34410 4404 34436 4436
rect 35016 4404 35042 4436
rect 35622 4404 35648 4436
rect 36228 4404 36254 4436
rect 36834 4404 36860 4436
rect 37440 4404 37466 4436
rect 38046 4404 38072 4436
rect 38652 4404 38678 4436
rect 39258 4404 39284 4436
rect 39864 4404 39890 4436
rect 40470 4404 40496 4436
rect 41076 4404 41102 4436
rect 41682 4404 41708 4436
rect 42288 4404 42314 4436
rect 42894 4404 42920 4436
rect 43500 4404 43526 4436
rect 44106 4404 44132 4436
rect 44712 4404 44738 4436
rect 45318 4404 45344 4436
rect 45924 4404 45950 4436
rect 46530 4404 46556 4436
rect 47136 4404 47162 4436
rect 47742 4404 47768 4436
rect 48348 4404 48374 4436
rect 48954 4404 48980 4436
rect 49560 4404 49586 4436
rect 50166 4404 50192 4436
rect 50772 4404 50798 4436
rect 51378 4404 51404 4436
rect 42298 4090 42322 4112
rect 32592 3244 32618 3276
rect 33198 3244 33224 3276
rect 33804 3244 33830 3276
rect 34410 3244 34436 3276
rect 35016 3244 35042 3276
rect 35622 3244 35648 3276
rect 36228 3244 36254 3276
rect 36834 3244 36860 3276
rect 37440 3244 37466 3276
rect 38046 3244 38072 3276
rect 38652 3244 38678 3276
rect 39258 3244 39284 3276
rect 39864 3244 39890 3276
rect 40470 3244 40496 3276
rect 41076 3244 41102 3276
rect 41682 3244 41708 3276
rect 42288 3244 42314 3276
rect 42894 3244 42920 3276
rect 43500 3244 43526 3276
rect 44106 3244 44132 3276
rect 44712 3244 44738 3276
rect 45318 3244 45344 3276
rect 45924 3244 45950 3276
rect 46530 3244 46556 3276
rect 47136 3244 47162 3276
rect 47742 3244 47768 3276
rect 48348 3244 48374 3276
rect 48954 3244 48980 3276
rect 49560 3244 49586 3276
rect 50166 3244 50192 3276
rect 50772 3244 50798 3276
rect 51378 3244 51404 3276
<< metal3 >>
rect 32272 5214 51730 5216
rect 32272 5150 32376 5214
rect 32440 5150 32456 5214
rect 32520 5150 32536 5214
rect 32600 5150 32616 5214
rect 32680 5150 32696 5214
rect 32760 5150 32776 5214
rect 32840 5150 32982 5214
rect 33046 5150 33062 5214
rect 33126 5150 33142 5214
rect 33206 5150 33222 5214
rect 33286 5150 33302 5214
rect 33366 5150 33382 5214
rect 33446 5150 33588 5214
rect 33652 5150 33668 5214
rect 33732 5150 33748 5214
rect 33812 5150 33828 5214
rect 33892 5150 33908 5214
rect 33972 5150 33988 5214
rect 34052 5150 34194 5214
rect 34258 5150 34274 5214
rect 34338 5150 34354 5214
rect 34418 5150 34434 5214
rect 34498 5150 34514 5214
rect 34578 5150 34594 5214
rect 34658 5150 34800 5214
rect 34864 5150 34880 5214
rect 34944 5150 34960 5214
rect 35024 5150 35040 5214
rect 35104 5150 35120 5214
rect 35184 5150 35200 5214
rect 35264 5150 35406 5214
rect 35470 5150 35486 5214
rect 35550 5150 35566 5214
rect 35630 5150 35646 5214
rect 35710 5150 35726 5214
rect 35790 5150 35806 5214
rect 35870 5150 36012 5214
rect 36076 5150 36092 5214
rect 36156 5150 36172 5214
rect 36236 5150 36252 5214
rect 36316 5150 36332 5214
rect 36396 5150 36412 5214
rect 36476 5150 36618 5214
rect 36682 5150 36698 5214
rect 36762 5150 36778 5214
rect 36842 5150 36858 5214
rect 36922 5150 36938 5214
rect 37002 5150 37018 5214
rect 37082 5150 37224 5214
rect 37288 5150 37304 5214
rect 37368 5150 37384 5214
rect 37448 5150 37464 5214
rect 37528 5150 37544 5214
rect 37608 5150 37624 5214
rect 37688 5150 37830 5214
rect 37894 5150 37910 5214
rect 37974 5150 37990 5214
rect 38054 5150 38070 5214
rect 38134 5150 38150 5214
rect 38214 5150 38230 5214
rect 38294 5150 38436 5214
rect 38500 5150 38516 5214
rect 38580 5150 38596 5214
rect 38660 5150 38676 5214
rect 38740 5150 38756 5214
rect 38820 5150 38836 5214
rect 38900 5150 39042 5214
rect 39106 5150 39122 5214
rect 39186 5150 39202 5214
rect 39266 5150 39282 5214
rect 39346 5150 39362 5214
rect 39426 5150 39442 5214
rect 39506 5150 39648 5214
rect 39712 5150 39728 5214
rect 39792 5150 39808 5214
rect 39872 5150 39888 5214
rect 39952 5150 39968 5214
rect 40032 5150 40048 5214
rect 40112 5150 40254 5214
rect 40318 5150 40334 5214
rect 40398 5150 40414 5214
rect 40478 5150 40494 5214
rect 40558 5150 40574 5214
rect 40638 5150 40654 5214
rect 40718 5150 40860 5214
rect 40924 5150 40940 5214
rect 41004 5150 41020 5214
rect 41084 5150 41100 5214
rect 41164 5150 41180 5214
rect 41244 5150 41260 5214
rect 41324 5150 41466 5214
rect 41530 5150 41546 5214
rect 41610 5150 41626 5214
rect 41690 5150 41706 5214
rect 41770 5150 41786 5214
rect 41850 5150 41866 5214
rect 41930 5150 42072 5214
rect 42136 5150 42152 5214
rect 42216 5150 42232 5214
rect 42296 5150 42312 5214
rect 42376 5150 42392 5214
rect 42456 5150 42472 5214
rect 42536 5150 42678 5214
rect 42742 5150 42758 5214
rect 42822 5150 42838 5214
rect 42902 5150 42918 5214
rect 42982 5150 42998 5214
rect 43062 5150 43078 5214
rect 43142 5150 43284 5214
rect 43348 5150 43364 5214
rect 43428 5150 43444 5214
rect 43508 5150 43524 5214
rect 43588 5150 43604 5214
rect 43668 5150 43684 5214
rect 43748 5150 43890 5214
rect 43954 5150 43970 5214
rect 44034 5150 44050 5214
rect 44114 5150 44130 5214
rect 44194 5150 44210 5214
rect 44274 5150 44290 5214
rect 44354 5150 44496 5214
rect 44560 5150 44576 5214
rect 44640 5150 44656 5214
rect 44720 5150 44736 5214
rect 44800 5150 44816 5214
rect 44880 5150 44896 5214
rect 44960 5150 45102 5214
rect 45166 5150 45182 5214
rect 45246 5150 45262 5214
rect 45326 5150 45342 5214
rect 45406 5150 45422 5214
rect 45486 5150 45502 5214
rect 45566 5150 45708 5214
rect 45772 5150 45788 5214
rect 45852 5150 45868 5214
rect 45932 5150 45948 5214
rect 46012 5150 46028 5214
rect 46092 5150 46108 5214
rect 46172 5150 46314 5214
rect 46378 5150 46394 5214
rect 46458 5150 46474 5214
rect 46538 5150 46554 5214
rect 46618 5150 46634 5214
rect 46698 5150 46714 5214
rect 46778 5150 46920 5214
rect 46984 5150 47000 5214
rect 47064 5150 47080 5214
rect 47144 5150 47160 5214
rect 47224 5150 47240 5214
rect 47304 5150 47320 5214
rect 47384 5150 47526 5214
rect 47590 5150 47606 5214
rect 47670 5150 47686 5214
rect 47750 5150 47766 5214
rect 47830 5150 47846 5214
rect 47910 5150 47926 5214
rect 47990 5150 48132 5214
rect 48196 5150 48212 5214
rect 48276 5150 48292 5214
rect 48356 5150 48372 5214
rect 48436 5150 48452 5214
rect 48516 5150 48532 5214
rect 48596 5150 48738 5214
rect 48802 5150 48818 5214
rect 48882 5150 48898 5214
rect 48962 5150 48978 5214
rect 49042 5150 49058 5214
rect 49122 5150 49138 5214
rect 49202 5150 49344 5214
rect 49408 5150 49424 5214
rect 49488 5150 49504 5214
rect 49568 5150 49584 5214
rect 49648 5150 49664 5214
rect 49728 5150 49744 5214
rect 49808 5150 49950 5214
rect 50014 5150 50030 5214
rect 50094 5150 50110 5214
rect 50174 5150 50190 5214
rect 50254 5150 50270 5214
rect 50334 5150 50350 5214
rect 50414 5150 50556 5214
rect 50620 5150 50636 5214
rect 50700 5150 50716 5214
rect 50780 5150 50796 5214
rect 50860 5150 50876 5214
rect 50940 5150 50956 5214
rect 51020 5150 51162 5214
rect 51226 5150 51242 5214
rect 51306 5150 51322 5214
rect 51386 5150 51402 5214
rect 51466 5150 51482 5214
rect 51546 5150 51562 5214
rect 51626 5150 51730 5214
rect 32272 5148 51730 5150
rect 32272 4994 32338 5148
rect 32272 4930 32273 4994
rect 32337 4930 32338 4994
rect 32272 4914 32338 4930
rect 32272 4850 32273 4914
rect 32337 4850 32338 4914
rect 32272 4834 32338 4850
rect 32272 4770 32273 4834
rect 32337 4770 32338 4834
rect 32272 4754 32338 4770
rect 32272 4690 32273 4754
rect 32337 4690 32338 4754
rect 32272 4674 32338 4690
rect 32272 4610 32273 4674
rect 32337 4610 32338 4674
rect 32272 4594 32338 4610
rect 32272 4530 32273 4594
rect 32337 4530 32338 4594
rect 32272 4514 32338 4530
rect 32272 4450 32273 4514
rect 32337 4450 32338 4514
rect 32272 4434 32338 4450
rect 32272 4370 32273 4434
rect 32337 4370 32338 4434
rect 32272 4354 32338 4370
rect 32272 4290 32273 4354
rect 32337 4290 32338 4354
rect 32272 4274 32338 4290
rect 32272 4210 32273 4274
rect 32337 4210 32338 4274
rect 32272 4120 32338 4210
rect 32398 4116 32458 5148
rect 32518 4056 32578 5086
rect 32638 4116 32698 5148
rect 32758 4056 32818 5086
rect 32878 4994 32944 5148
rect 32878 4930 32879 4994
rect 32943 4930 32944 4994
rect 32878 4914 32944 4930
rect 32878 4850 32879 4914
rect 32943 4850 32944 4914
rect 32878 4834 32944 4850
rect 32878 4770 32879 4834
rect 32943 4770 32944 4834
rect 32878 4754 32944 4770
rect 32878 4690 32879 4754
rect 32943 4690 32944 4754
rect 32878 4674 32944 4690
rect 32878 4610 32879 4674
rect 32943 4610 32944 4674
rect 32878 4594 32944 4610
rect 32878 4530 32879 4594
rect 32943 4530 32944 4594
rect 32878 4514 32944 4530
rect 32878 4450 32879 4514
rect 32943 4450 32944 4514
rect 32878 4434 32944 4450
rect 32878 4370 32879 4434
rect 32943 4370 32944 4434
rect 32878 4354 32944 4370
rect 32878 4290 32879 4354
rect 32943 4290 32944 4354
rect 32878 4274 32944 4290
rect 32878 4210 32879 4274
rect 32943 4210 32944 4274
rect 32878 4120 32944 4210
rect 33004 4116 33064 5148
rect 33124 4056 33184 5086
rect 33244 4116 33304 5148
rect 33364 4056 33424 5086
rect 33484 4994 33550 5148
rect 33484 4930 33485 4994
rect 33549 4930 33550 4994
rect 33484 4914 33550 4930
rect 33484 4850 33485 4914
rect 33549 4850 33550 4914
rect 33484 4834 33550 4850
rect 33484 4770 33485 4834
rect 33549 4770 33550 4834
rect 33484 4754 33550 4770
rect 33484 4690 33485 4754
rect 33549 4690 33550 4754
rect 33484 4674 33550 4690
rect 33484 4610 33485 4674
rect 33549 4610 33550 4674
rect 33484 4594 33550 4610
rect 33484 4530 33485 4594
rect 33549 4530 33550 4594
rect 33484 4514 33550 4530
rect 33484 4450 33485 4514
rect 33549 4450 33550 4514
rect 33484 4434 33550 4450
rect 33484 4370 33485 4434
rect 33549 4370 33550 4434
rect 33484 4354 33550 4370
rect 33484 4290 33485 4354
rect 33549 4290 33550 4354
rect 33484 4274 33550 4290
rect 33484 4210 33485 4274
rect 33549 4210 33550 4274
rect 33484 4120 33550 4210
rect 33610 4116 33670 5148
rect 33730 4056 33790 5086
rect 33850 4116 33910 5148
rect 33970 4056 34030 5086
rect 34090 4994 34156 5148
rect 34090 4930 34091 4994
rect 34155 4930 34156 4994
rect 34090 4914 34156 4930
rect 34090 4850 34091 4914
rect 34155 4850 34156 4914
rect 34090 4834 34156 4850
rect 34090 4770 34091 4834
rect 34155 4770 34156 4834
rect 34090 4754 34156 4770
rect 34090 4690 34091 4754
rect 34155 4690 34156 4754
rect 34090 4674 34156 4690
rect 34090 4610 34091 4674
rect 34155 4610 34156 4674
rect 34090 4594 34156 4610
rect 34090 4530 34091 4594
rect 34155 4530 34156 4594
rect 34090 4514 34156 4530
rect 34090 4450 34091 4514
rect 34155 4450 34156 4514
rect 34090 4434 34156 4450
rect 34090 4370 34091 4434
rect 34155 4370 34156 4434
rect 34090 4354 34156 4370
rect 34090 4290 34091 4354
rect 34155 4290 34156 4354
rect 34090 4274 34156 4290
rect 34090 4210 34091 4274
rect 34155 4210 34156 4274
rect 34090 4120 34156 4210
rect 34216 4116 34276 5148
rect 34336 4056 34396 5086
rect 34456 4116 34516 5148
rect 34576 4056 34636 5086
rect 34696 4994 34762 5148
rect 34696 4930 34697 4994
rect 34761 4930 34762 4994
rect 34696 4914 34762 4930
rect 34696 4850 34697 4914
rect 34761 4850 34762 4914
rect 34696 4834 34762 4850
rect 34696 4770 34697 4834
rect 34761 4770 34762 4834
rect 34696 4754 34762 4770
rect 34696 4690 34697 4754
rect 34761 4690 34762 4754
rect 34696 4674 34762 4690
rect 34696 4610 34697 4674
rect 34761 4610 34762 4674
rect 34696 4594 34762 4610
rect 34696 4530 34697 4594
rect 34761 4530 34762 4594
rect 34696 4514 34762 4530
rect 34696 4450 34697 4514
rect 34761 4450 34762 4514
rect 34696 4434 34762 4450
rect 34696 4370 34697 4434
rect 34761 4370 34762 4434
rect 34696 4354 34762 4370
rect 34696 4290 34697 4354
rect 34761 4290 34762 4354
rect 34696 4274 34762 4290
rect 34696 4210 34697 4274
rect 34761 4210 34762 4274
rect 34696 4120 34762 4210
rect 34822 4116 34882 5148
rect 34942 4056 35002 5086
rect 35062 4116 35122 5148
rect 35182 4056 35242 5086
rect 35302 4994 35368 5148
rect 35302 4930 35303 4994
rect 35367 4930 35368 4994
rect 35302 4914 35368 4930
rect 35302 4850 35303 4914
rect 35367 4850 35368 4914
rect 35302 4834 35368 4850
rect 35302 4770 35303 4834
rect 35367 4770 35368 4834
rect 35302 4754 35368 4770
rect 35302 4690 35303 4754
rect 35367 4690 35368 4754
rect 35302 4674 35368 4690
rect 35302 4610 35303 4674
rect 35367 4610 35368 4674
rect 35302 4594 35368 4610
rect 35302 4530 35303 4594
rect 35367 4530 35368 4594
rect 35302 4514 35368 4530
rect 35302 4450 35303 4514
rect 35367 4450 35368 4514
rect 35302 4434 35368 4450
rect 35302 4370 35303 4434
rect 35367 4370 35368 4434
rect 35302 4354 35368 4370
rect 35302 4290 35303 4354
rect 35367 4290 35368 4354
rect 35302 4274 35368 4290
rect 35302 4210 35303 4274
rect 35367 4210 35368 4274
rect 35302 4120 35368 4210
rect 35428 4116 35488 5148
rect 35548 4056 35608 5086
rect 35668 4116 35728 5148
rect 35788 4056 35848 5086
rect 35908 4994 35974 5148
rect 35908 4930 35909 4994
rect 35973 4930 35974 4994
rect 35908 4914 35974 4930
rect 35908 4850 35909 4914
rect 35973 4850 35974 4914
rect 35908 4834 35974 4850
rect 35908 4770 35909 4834
rect 35973 4770 35974 4834
rect 35908 4754 35974 4770
rect 35908 4690 35909 4754
rect 35973 4690 35974 4754
rect 35908 4674 35974 4690
rect 35908 4610 35909 4674
rect 35973 4610 35974 4674
rect 35908 4594 35974 4610
rect 35908 4530 35909 4594
rect 35973 4530 35974 4594
rect 35908 4514 35974 4530
rect 35908 4450 35909 4514
rect 35973 4450 35974 4514
rect 35908 4434 35974 4450
rect 35908 4370 35909 4434
rect 35973 4370 35974 4434
rect 35908 4354 35974 4370
rect 35908 4290 35909 4354
rect 35973 4290 35974 4354
rect 35908 4274 35974 4290
rect 35908 4210 35909 4274
rect 35973 4210 35974 4274
rect 35908 4120 35974 4210
rect 36034 4116 36094 5148
rect 36154 4056 36214 5086
rect 36274 4116 36334 5148
rect 36394 4056 36454 5086
rect 36514 4994 36580 5148
rect 36514 4930 36515 4994
rect 36579 4930 36580 4994
rect 36514 4914 36580 4930
rect 36514 4850 36515 4914
rect 36579 4850 36580 4914
rect 36514 4834 36580 4850
rect 36514 4770 36515 4834
rect 36579 4770 36580 4834
rect 36514 4754 36580 4770
rect 36514 4690 36515 4754
rect 36579 4690 36580 4754
rect 36514 4674 36580 4690
rect 36514 4610 36515 4674
rect 36579 4610 36580 4674
rect 36514 4594 36580 4610
rect 36514 4530 36515 4594
rect 36579 4530 36580 4594
rect 36514 4514 36580 4530
rect 36514 4450 36515 4514
rect 36579 4450 36580 4514
rect 36514 4434 36580 4450
rect 36514 4370 36515 4434
rect 36579 4370 36580 4434
rect 36514 4354 36580 4370
rect 36514 4290 36515 4354
rect 36579 4290 36580 4354
rect 36514 4274 36580 4290
rect 36514 4210 36515 4274
rect 36579 4210 36580 4274
rect 36514 4120 36580 4210
rect 36640 4116 36700 5148
rect 36760 4056 36820 5086
rect 36880 4116 36940 5148
rect 37000 4056 37060 5086
rect 37120 4994 37186 5148
rect 37120 4930 37121 4994
rect 37185 4930 37186 4994
rect 37120 4914 37186 4930
rect 37120 4850 37121 4914
rect 37185 4850 37186 4914
rect 37120 4834 37186 4850
rect 37120 4770 37121 4834
rect 37185 4770 37186 4834
rect 37120 4754 37186 4770
rect 37120 4690 37121 4754
rect 37185 4690 37186 4754
rect 37120 4674 37186 4690
rect 37120 4610 37121 4674
rect 37185 4610 37186 4674
rect 37120 4594 37186 4610
rect 37120 4530 37121 4594
rect 37185 4530 37186 4594
rect 37120 4514 37186 4530
rect 37120 4450 37121 4514
rect 37185 4450 37186 4514
rect 37120 4434 37186 4450
rect 37120 4370 37121 4434
rect 37185 4370 37186 4434
rect 37120 4354 37186 4370
rect 37120 4290 37121 4354
rect 37185 4290 37186 4354
rect 37120 4274 37186 4290
rect 37120 4210 37121 4274
rect 37185 4210 37186 4274
rect 37120 4120 37186 4210
rect 37246 4116 37306 5148
rect 37366 4056 37426 5086
rect 37486 4116 37546 5148
rect 37606 4056 37666 5086
rect 37726 4994 37792 5148
rect 37726 4930 37727 4994
rect 37791 4930 37792 4994
rect 37726 4914 37792 4930
rect 37726 4850 37727 4914
rect 37791 4850 37792 4914
rect 37726 4834 37792 4850
rect 37726 4770 37727 4834
rect 37791 4770 37792 4834
rect 37726 4754 37792 4770
rect 37726 4690 37727 4754
rect 37791 4690 37792 4754
rect 37726 4674 37792 4690
rect 37726 4610 37727 4674
rect 37791 4610 37792 4674
rect 37726 4594 37792 4610
rect 37726 4530 37727 4594
rect 37791 4530 37792 4594
rect 37726 4514 37792 4530
rect 37726 4450 37727 4514
rect 37791 4450 37792 4514
rect 37726 4434 37792 4450
rect 37726 4370 37727 4434
rect 37791 4370 37792 4434
rect 37726 4354 37792 4370
rect 37726 4290 37727 4354
rect 37791 4290 37792 4354
rect 37726 4274 37792 4290
rect 37726 4210 37727 4274
rect 37791 4210 37792 4274
rect 37726 4120 37792 4210
rect 37852 4116 37912 5148
rect 37972 4056 38032 5086
rect 38092 4116 38152 5148
rect 38212 4056 38272 5086
rect 38332 4994 38398 5148
rect 38332 4930 38333 4994
rect 38397 4930 38398 4994
rect 38332 4914 38398 4930
rect 38332 4850 38333 4914
rect 38397 4850 38398 4914
rect 38332 4834 38398 4850
rect 38332 4770 38333 4834
rect 38397 4770 38398 4834
rect 38332 4754 38398 4770
rect 38332 4690 38333 4754
rect 38397 4690 38398 4754
rect 38332 4674 38398 4690
rect 38332 4610 38333 4674
rect 38397 4610 38398 4674
rect 38332 4594 38398 4610
rect 38332 4530 38333 4594
rect 38397 4530 38398 4594
rect 38332 4514 38398 4530
rect 38332 4450 38333 4514
rect 38397 4450 38398 4514
rect 38332 4434 38398 4450
rect 38332 4370 38333 4434
rect 38397 4370 38398 4434
rect 38332 4354 38398 4370
rect 38332 4290 38333 4354
rect 38397 4290 38398 4354
rect 38332 4274 38398 4290
rect 38332 4210 38333 4274
rect 38397 4210 38398 4274
rect 38332 4120 38398 4210
rect 38458 4116 38518 5148
rect 38578 4056 38638 5086
rect 38698 4116 38758 5148
rect 38818 4056 38878 5086
rect 38938 4994 39004 5148
rect 38938 4930 38939 4994
rect 39003 4930 39004 4994
rect 38938 4914 39004 4930
rect 38938 4850 38939 4914
rect 39003 4850 39004 4914
rect 38938 4834 39004 4850
rect 38938 4770 38939 4834
rect 39003 4770 39004 4834
rect 38938 4754 39004 4770
rect 38938 4690 38939 4754
rect 39003 4690 39004 4754
rect 38938 4674 39004 4690
rect 38938 4610 38939 4674
rect 39003 4610 39004 4674
rect 38938 4594 39004 4610
rect 38938 4530 38939 4594
rect 39003 4530 39004 4594
rect 38938 4514 39004 4530
rect 38938 4450 38939 4514
rect 39003 4450 39004 4514
rect 38938 4434 39004 4450
rect 38938 4370 38939 4434
rect 39003 4370 39004 4434
rect 38938 4354 39004 4370
rect 38938 4290 38939 4354
rect 39003 4290 39004 4354
rect 38938 4274 39004 4290
rect 38938 4210 38939 4274
rect 39003 4210 39004 4274
rect 38938 4120 39004 4210
rect 39064 4116 39124 5148
rect 39184 4056 39244 5086
rect 39304 4116 39364 5148
rect 39424 4056 39484 5086
rect 39544 4994 39610 5148
rect 39544 4930 39545 4994
rect 39609 4930 39610 4994
rect 39544 4914 39610 4930
rect 39544 4850 39545 4914
rect 39609 4850 39610 4914
rect 39544 4834 39610 4850
rect 39544 4770 39545 4834
rect 39609 4770 39610 4834
rect 39544 4754 39610 4770
rect 39544 4690 39545 4754
rect 39609 4690 39610 4754
rect 39544 4674 39610 4690
rect 39544 4610 39545 4674
rect 39609 4610 39610 4674
rect 39544 4594 39610 4610
rect 39544 4530 39545 4594
rect 39609 4530 39610 4594
rect 39544 4514 39610 4530
rect 39544 4450 39545 4514
rect 39609 4450 39610 4514
rect 39544 4434 39610 4450
rect 39544 4370 39545 4434
rect 39609 4370 39610 4434
rect 39544 4354 39610 4370
rect 39544 4290 39545 4354
rect 39609 4290 39610 4354
rect 39544 4274 39610 4290
rect 39544 4210 39545 4274
rect 39609 4210 39610 4274
rect 39544 4120 39610 4210
rect 39670 4116 39730 5148
rect 39790 4056 39850 5086
rect 39910 4116 39970 5148
rect 40030 4056 40090 5086
rect 40150 4994 40216 5148
rect 40150 4930 40151 4994
rect 40215 4930 40216 4994
rect 40150 4914 40216 4930
rect 40150 4850 40151 4914
rect 40215 4850 40216 4914
rect 40150 4834 40216 4850
rect 40150 4770 40151 4834
rect 40215 4770 40216 4834
rect 40150 4754 40216 4770
rect 40150 4690 40151 4754
rect 40215 4690 40216 4754
rect 40150 4674 40216 4690
rect 40150 4610 40151 4674
rect 40215 4610 40216 4674
rect 40150 4594 40216 4610
rect 40150 4530 40151 4594
rect 40215 4530 40216 4594
rect 40150 4514 40216 4530
rect 40150 4450 40151 4514
rect 40215 4450 40216 4514
rect 40150 4434 40216 4450
rect 40150 4370 40151 4434
rect 40215 4370 40216 4434
rect 40150 4354 40216 4370
rect 40150 4290 40151 4354
rect 40215 4290 40216 4354
rect 40150 4274 40216 4290
rect 40150 4210 40151 4274
rect 40215 4210 40216 4274
rect 40150 4120 40216 4210
rect 40276 4116 40336 5148
rect 40396 4056 40456 5086
rect 40516 4116 40576 5148
rect 40636 4056 40696 5086
rect 40756 4994 40822 5148
rect 40756 4930 40757 4994
rect 40821 4930 40822 4994
rect 40756 4914 40822 4930
rect 40756 4850 40757 4914
rect 40821 4850 40822 4914
rect 40756 4834 40822 4850
rect 40756 4770 40757 4834
rect 40821 4770 40822 4834
rect 40756 4754 40822 4770
rect 40756 4690 40757 4754
rect 40821 4690 40822 4754
rect 40756 4674 40822 4690
rect 40756 4610 40757 4674
rect 40821 4610 40822 4674
rect 40756 4594 40822 4610
rect 40756 4530 40757 4594
rect 40821 4530 40822 4594
rect 40756 4514 40822 4530
rect 40756 4450 40757 4514
rect 40821 4450 40822 4514
rect 40756 4434 40822 4450
rect 40756 4370 40757 4434
rect 40821 4370 40822 4434
rect 40756 4354 40822 4370
rect 40756 4290 40757 4354
rect 40821 4290 40822 4354
rect 40756 4274 40822 4290
rect 40756 4210 40757 4274
rect 40821 4210 40822 4274
rect 40756 4120 40822 4210
rect 40882 4116 40942 5148
rect 41002 4056 41062 5086
rect 41122 4116 41182 5148
rect 41242 4056 41302 5086
rect 41362 4994 41428 5148
rect 41362 4930 41363 4994
rect 41427 4930 41428 4994
rect 41362 4914 41428 4930
rect 41362 4850 41363 4914
rect 41427 4850 41428 4914
rect 41362 4834 41428 4850
rect 41362 4770 41363 4834
rect 41427 4770 41428 4834
rect 41362 4754 41428 4770
rect 41362 4690 41363 4754
rect 41427 4690 41428 4754
rect 41362 4674 41428 4690
rect 41362 4610 41363 4674
rect 41427 4610 41428 4674
rect 41362 4594 41428 4610
rect 41362 4530 41363 4594
rect 41427 4530 41428 4594
rect 41362 4514 41428 4530
rect 41362 4450 41363 4514
rect 41427 4450 41428 4514
rect 41362 4434 41428 4450
rect 41362 4370 41363 4434
rect 41427 4370 41428 4434
rect 41362 4354 41428 4370
rect 41362 4290 41363 4354
rect 41427 4290 41428 4354
rect 41362 4274 41428 4290
rect 41362 4210 41363 4274
rect 41427 4210 41428 4274
rect 41362 4120 41428 4210
rect 41488 4116 41548 5148
rect 41608 4056 41668 5086
rect 41728 4116 41788 5148
rect 41848 4056 41908 5086
rect 41968 4994 42034 5148
rect 41968 4930 41969 4994
rect 42033 4930 42034 4994
rect 41968 4914 42034 4930
rect 41968 4850 41969 4914
rect 42033 4850 42034 4914
rect 41968 4834 42034 4850
rect 41968 4770 41969 4834
rect 42033 4770 42034 4834
rect 41968 4754 42034 4770
rect 41968 4690 41969 4754
rect 42033 4690 42034 4754
rect 41968 4674 42034 4690
rect 41968 4610 41969 4674
rect 42033 4610 42034 4674
rect 41968 4594 42034 4610
rect 41968 4530 41969 4594
rect 42033 4530 42034 4594
rect 41968 4514 42034 4530
rect 41968 4450 41969 4514
rect 42033 4450 42034 4514
rect 41968 4434 42034 4450
rect 41968 4370 41969 4434
rect 42033 4370 42034 4434
rect 41968 4354 42034 4370
rect 41968 4290 41969 4354
rect 42033 4290 42034 4354
rect 41968 4274 42034 4290
rect 41968 4210 41969 4274
rect 42033 4210 42034 4274
rect 41968 4120 42034 4210
rect 42094 4116 42154 5148
rect 42214 4056 42274 5086
rect 42334 4116 42394 5148
rect 42454 4056 42514 5086
rect 42574 4994 42640 5148
rect 42574 4930 42575 4994
rect 42639 4930 42640 4994
rect 42574 4914 42640 4930
rect 42574 4850 42575 4914
rect 42639 4850 42640 4914
rect 42574 4834 42640 4850
rect 42574 4770 42575 4834
rect 42639 4770 42640 4834
rect 42574 4754 42640 4770
rect 42574 4690 42575 4754
rect 42639 4690 42640 4754
rect 42574 4674 42640 4690
rect 42574 4610 42575 4674
rect 42639 4610 42640 4674
rect 42574 4594 42640 4610
rect 42574 4530 42575 4594
rect 42639 4530 42640 4594
rect 42574 4514 42640 4530
rect 42574 4450 42575 4514
rect 42639 4450 42640 4514
rect 42574 4434 42640 4450
rect 42574 4370 42575 4434
rect 42639 4370 42640 4434
rect 42574 4354 42640 4370
rect 42574 4290 42575 4354
rect 42639 4290 42640 4354
rect 42574 4274 42640 4290
rect 42574 4210 42575 4274
rect 42639 4210 42640 4274
rect 42574 4120 42640 4210
rect 42700 4116 42760 5148
rect 42820 4056 42880 5086
rect 42940 4116 43000 5148
rect 43060 4056 43120 5086
rect 43180 4994 43246 5148
rect 43180 4930 43181 4994
rect 43245 4930 43246 4994
rect 43180 4914 43246 4930
rect 43180 4850 43181 4914
rect 43245 4850 43246 4914
rect 43180 4834 43246 4850
rect 43180 4770 43181 4834
rect 43245 4770 43246 4834
rect 43180 4754 43246 4770
rect 43180 4690 43181 4754
rect 43245 4690 43246 4754
rect 43180 4674 43246 4690
rect 43180 4610 43181 4674
rect 43245 4610 43246 4674
rect 43180 4594 43246 4610
rect 43180 4530 43181 4594
rect 43245 4530 43246 4594
rect 43180 4514 43246 4530
rect 43180 4450 43181 4514
rect 43245 4450 43246 4514
rect 43180 4434 43246 4450
rect 43180 4370 43181 4434
rect 43245 4370 43246 4434
rect 43180 4354 43246 4370
rect 43180 4290 43181 4354
rect 43245 4290 43246 4354
rect 43180 4274 43246 4290
rect 43180 4210 43181 4274
rect 43245 4210 43246 4274
rect 43180 4120 43246 4210
rect 43306 4116 43366 5148
rect 43426 4056 43486 5086
rect 43546 4116 43606 5148
rect 43666 4056 43726 5086
rect 43786 4994 43852 5148
rect 43786 4930 43787 4994
rect 43851 4930 43852 4994
rect 43786 4914 43852 4930
rect 43786 4850 43787 4914
rect 43851 4850 43852 4914
rect 43786 4834 43852 4850
rect 43786 4770 43787 4834
rect 43851 4770 43852 4834
rect 43786 4754 43852 4770
rect 43786 4690 43787 4754
rect 43851 4690 43852 4754
rect 43786 4674 43852 4690
rect 43786 4610 43787 4674
rect 43851 4610 43852 4674
rect 43786 4594 43852 4610
rect 43786 4530 43787 4594
rect 43851 4530 43852 4594
rect 43786 4514 43852 4530
rect 43786 4450 43787 4514
rect 43851 4450 43852 4514
rect 43786 4434 43852 4450
rect 43786 4370 43787 4434
rect 43851 4370 43852 4434
rect 43786 4354 43852 4370
rect 43786 4290 43787 4354
rect 43851 4290 43852 4354
rect 43786 4274 43852 4290
rect 43786 4210 43787 4274
rect 43851 4210 43852 4274
rect 43786 4120 43852 4210
rect 43912 4116 43972 5148
rect 44032 4056 44092 5086
rect 44152 4116 44212 5148
rect 44272 4056 44332 5086
rect 44392 4994 44458 5148
rect 44392 4930 44393 4994
rect 44457 4930 44458 4994
rect 44392 4914 44458 4930
rect 44392 4850 44393 4914
rect 44457 4850 44458 4914
rect 44392 4834 44458 4850
rect 44392 4770 44393 4834
rect 44457 4770 44458 4834
rect 44392 4754 44458 4770
rect 44392 4690 44393 4754
rect 44457 4690 44458 4754
rect 44392 4674 44458 4690
rect 44392 4610 44393 4674
rect 44457 4610 44458 4674
rect 44392 4594 44458 4610
rect 44392 4530 44393 4594
rect 44457 4530 44458 4594
rect 44392 4514 44458 4530
rect 44392 4450 44393 4514
rect 44457 4450 44458 4514
rect 44392 4434 44458 4450
rect 44392 4370 44393 4434
rect 44457 4370 44458 4434
rect 44392 4354 44458 4370
rect 44392 4290 44393 4354
rect 44457 4290 44458 4354
rect 44392 4274 44458 4290
rect 44392 4210 44393 4274
rect 44457 4210 44458 4274
rect 44392 4120 44458 4210
rect 44518 4116 44578 5148
rect 44638 4056 44698 5086
rect 44758 4116 44818 5148
rect 44878 4056 44938 5086
rect 44998 4994 45064 5148
rect 44998 4930 44999 4994
rect 45063 4930 45064 4994
rect 44998 4914 45064 4930
rect 44998 4850 44999 4914
rect 45063 4850 45064 4914
rect 44998 4834 45064 4850
rect 44998 4770 44999 4834
rect 45063 4770 45064 4834
rect 44998 4754 45064 4770
rect 44998 4690 44999 4754
rect 45063 4690 45064 4754
rect 44998 4674 45064 4690
rect 44998 4610 44999 4674
rect 45063 4610 45064 4674
rect 44998 4594 45064 4610
rect 44998 4530 44999 4594
rect 45063 4530 45064 4594
rect 44998 4514 45064 4530
rect 44998 4450 44999 4514
rect 45063 4450 45064 4514
rect 44998 4434 45064 4450
rect 44998 4370 44999 4434
rect 45063 4370 45064 4434
rect 44998 4354 45064 4370
rect 44998 4290 44999 4354
rect 45063 4290 45064 4354
rect 44998 4274 45064 4290
rect 44998 4210 44999 4274
rect 45063 4210 45064 4274
rect 44998 4120 45064 4210
rect 45124 4116 45184 5148
rect 45244 4056 45304 5086
rect 45364 4116 45424 5148
rect 45484 4056 45544 5086
rect 45604 4994 45670 5148
rect 45604 4930 45605 4994
rect 45669 4930 45670 4994
rect 45604 4914 45670 4930
rect 45604 4850 45605 4914
rect 45669 4850 45670 4914
rect 45604 4834 45670 4850
rect 45604 4770 45605 4834
rect 45669 4770 45670 4834
rect 45604 4754 45670 4770
rect 45604 4690 45605 4754
rect 45669 4690 45670 4754
rect 45604 4674 45670 4690
rect 45604 4610 45605 4674
rect 45669 4610 45670 4674
rect 45604 4594 45670 4610
rect 45604 4530 45605 4594
rect 45669 4530 45670 4594
rect 45604 4514 45670 4530
rect 45604 4450 45605 4514
rect 45669 4450 45670 4514
rect 45604 4434 45670 4450
rect 45604 4370 45605 4434
rect 45669 4370 45670 4434
rect 45604 4354 45670 4370
rect 45604 4290 45605 4354
rect 45669 4290 45670 4354
rect 45604 4274 45670 4290
rect 45604 4210 45605 4274
rect 45669 4210 45670 4274
rect 45604 4120 45670 4210
rect 45730 4116 45790 5148
rect 45850 4056 45910 5086
rect 45970 4116 46030 5148
rect 46090 4056 46150 5086
rect 46210 4994 46276 5148
rect 46210 4930 46211 4994
rect 46275 4930 46276 4994
rect 46210 4914 46276 4930
rect 46210 4850 46211 4914
rect 46275 4850 46276 4914
rect 46210 4834 46276 4850
rect 46210 4770 46211 4834
rect 46275 4770 46276 4834
rect 46210 4754 46276 4770
rect 46210 4690 46211 4754
rect 46275 4690 46276 4754
rect 46210 4674 46276 4690
rect 46210 4610 46211 4674
rect 46275 4610 46276 4674
rect 46210 4594 46276 4610
rect 46210 4530 46211 4594
rect 46275 4530 46276 4594
rect 46210 4514 46276 4530
rect 46210 4450 46211 4514
rect 46275 4450 46276 4514
rect 46210 4434 46276 4450
rect 46210 4370 46211 4434
rect 46275 4370 46276 4434
rect 46210 4354 46276 4370
rect 46210 4290 46211 4354
rect 46275 4290 46276 4354
rect 46210 4274 46276 4290
rect 46210 4210 46211 4274
rect 46275 4210 46276 4274
rect 46210 4120 46276 4210
rect 46336 4116 46396 5148
rect 46456 4056 46516 5086
rect 46576 4116 46636 5148
rect 46696 4056 46756 5086
rect 46816 4994 46882 5148
rect 46816 4930 46817 4994
rect 46881 4930 46882 4994
rect 46816 4914 46882 4930
rect 46816 4850 46817 4914
rect 46881 4850 46882 4914
rect 46816 4834 46882 4850
rect 46816 4770 46817 4834
rect 46881 4770 46882 4834
rect 46816 4754 46882 4770
rect 46816 4690 46817 4754
rect 46881 4690 46882 4754
rect 46816 4674 46882 4690
rect 46816 4610 46817 4674
rect 46881 4610 46882 4674
rect 46816 4594 46882 4610
rect 46816 4530 46817 4594
rect 46881 4530 46882 4594
rect 46816 4514 46882 4530
rect 46816 4450 46817 4514
rect 46881 4450 46882 4514
rect 46816 4434 46882 4450
rect 46816 4370 46817 4434
rect 46881 4370 46882 4434
rect 46816 4354 46882 4370
rect 46816 4290 46817 4354
rect 46881 4290 46882 4354
rect 46816 4274 46882 4290
rect 46816 4210 46817 4274
rect 46881 4210 46882 4274
rect 46816 4120 46882 4210
rect 46942 4116 47002 5148
rect 47062 4056 47122 5086
rect 47182 4116 47242 5148
rect 47302 4056 47362 5086
rect 47422 4994 47488 5148
rect 47422 4930 47423 4994
rect 47487 4930 47488 4994
rect 47422 4914 47488 4930
rect 47422 4850 47423 4914
rect 47487 4850 47488 4914
rect 47422 4834 47488 4850
rect 47422 4770 47423 4834
rect 47487 4770 47488 4834
rect 47422 4754 47488 4770
rect 47422 4690 47423 4754
rect 47487 4690 47488 4754
rect 47422 4674 47488 4690
rect 47422 4610 47423 4674
rect 47487 4610 47488 4674
rect 47422 4594 47488 4610
rect 47422 4530 47423 4594
rect 47487 4530 47488 4594
rect 47422 4514 47488 4530
rect 47422 4450 47423 4514
rect 47487 4450 47488 4514
rect 47422 4434 47488 4450
rect 47422 4370 47423 4434
rect 47487 4370 47488 4434
rect 47422 4354 47488 4370
rect 47422 4290 47423 4354
rect 47487 4290 47488 4354
rect 47422 4274 47488 4290
rect 47422 4210 47423 4274
rect 47487 4210 47488 4274
rect 47422 4120 47488 4210
rect 47548 4116 47608 5148
rect 47668 4056 47728 5086
rect 47788 4116 47848 5148
rect 47908 4056 47968 5086
rect 48028 4994 48094 5148
rect 48028 4930 48029 4994
rect 48093 4930 48094 4994
rect 48028 4914 48094 4930
rect 48028 4850 48029 4914
rect 48093 4850 48094 4914
rect 48028 4834 48094 4850
rect 48028 4770 48029 4834
rect 48093 4770 48094 4834
rect 48028 4754 48094 4770
rect 48028 4690 48029 4754
rect 48093 4690 48094 4754
rect 48028 4674 48094 4690
rect 48028 4610 48029 4674
rect 48093 4610 48094 4674
rect 48028 4594 48094 4610
rect 48028 4530 48029 4594
rect 48093 4530 48094 4594
rect 48028 4514 48094 4530
rect 48028 4450 48029 4514
rect 48093 4450 48094 4514
rect 48028 4434 48094 4450
rect 48028 4370 48029 4434
rect 48093 4370 48094 4434
rect 48028 4354 48094 4370
rect 48028 4290 48029 4354
rect 48093 4290 48094 4354
rect 48028 4274 48094 4290
rect 48028 4210 48029 4274
rect 48093 4210 48094 4274
rect 48028 4120 48094 4210
rect 48154 4116 48214 5148
rect 48274 4056 48334 5086
rect 48394 4116 48454 5148
rect 48514 4056 48574 5086
rect 48634 4994 48700 5148
rect 48634 4930 48635 4994
rect 48699 4930 48700 4994
rect 48634 4914 48700 4930
rect 48634 4850 48635 4914
rect 48699 4850 48700 4914
rect 48634 4834 48700 4850
rect 48634 4770 48635 4834
rect 48699 4770 48700 4834
rect 48634 4754 48700 4770
rect 48634 4690 48635 4754
rect 48699 4690 48700 4754
rect 48634 4674 48700 4690
rect 48634 4610 48635 4674
rect 48699 4610 48700 4674
rect 48634 4594 48700 4610
rect 48634 4530 48635 4594
rect 48699 4530 48700 4594
rect 48634 4514 48700 4530
rect 48634 4450 48635 4514
rect 48699 4450 48700 4514
rect 48634 4434 48700 4450
rect 48634 4370 48635 4434
rect 48699 4370 48700 4434
rect 48634 4354 48700 4370
rect 48634 4290 48635 4354
rect 48699 4290 48700 4354
rect 48634 4274 48700 4290
rect 48634 4210 48635 4274
rect 48699 4210 48700 4274
rect 48634 4120 48700 4210
rect 48760 4116 48820 5148
rect 48880 4056 48940 5086
rect 49000 4116 49060 5148
rect 49120 4056 49180 5086
rect 49240 4994 49306 5148
rect 49240 4930 49241 4994
rect 49305 4930 49306 4994
rect 49240 4914 49306 4930
rect 49240 4850 49241 4914
rect 49305 4850 49306 4914
rect 49240 4834 49306 4850
rect 49240 4770 49241 4834
rect 49305 4770 49306 4834
rect 49240 4754 49306 4770
rect 49240 4690 49241 4754
rect 49305 4690 49306 4754
rect 49240 4674 49306 4690
rect 49240 4610 49241 4674
rect 49305 4610 49306 4674
rect 49240 4594 49306 4610
rect 49240 4530 49241 4594
rect 49305 4530 49306 4594
rect 49240 4514 49306 4530
rect 49240 4450 49241 4514
rect 49305 4450 49306 4514
rect 49240 4434 49306 4450
rect 49240 4370 49241 4434
rect 49305 4370 49306 4434
rect 49240 4354 49306 4370
rect 49240 4290 49241 4354
rect 49305 4290 49306 4354
rect 49240 4274 49306 4290
rect 49240 4210 49241 4274
rect 49305 4210 49306 4274
rect 49240 4120 49306 4210
rect 49366 4116 49426 5148
rect 49486 4056 49546 5086
rect 49606 4116 49666 5148
rect 49726 4056 49786 5086
rect 49846 4994 49912 5148
rect 49846 4930 49847 4994
rect 49911 4930 49912 4994
rect 49846 4914 49912 4930
rect 49846 4850 49847 4914
rect 49911 4850 49912 4914
rect 49846 4834 49912 4850
rect 49846 4770 49847 4834
rect 49911 4770 49912 4834
rect 49846 4754 49912 4770
rect 49846 4690 49847 4754
rect 49911 4690 49912 4754
rect 49846 4674 49912 4690
rect 49846 4610 49847 4674
rect 49911 4610 49912 4674
rect 49846 4594 49912 4610
rect 49846 4530 49847 4594
rect 49911 4530 49912 4594
rect 49846 4514 49912 4530
rect 49846 4450 49847 4514
rect 49911 4450 49912 4514
rect 49846 4434 49912 4450
rect 49846 4370 49847 4434
rect 49911 4370 49912 4434
rect 49846 4354 49912 4370
rect 49846 4290 49847 4354
rect 49911 4290 49912 4354
rect 49846 4274 49912 4290
rect 49846 4210 49847 4274
rect 49911 4210 49912 4274
rect 49846 4120 49912 4210
rect 49972 4116 50032 5148
rect 50092 4056 50152 5086
rect 50212 4116 50272 5148
rect 50332 4056 50392 5086
rect 50452 4994 50518 5148
rect 50452 4930 50453 4994
rect 50517 4930 50518 4994
rect 50452 4914 50518 4930
rect 50452 4850 50453 4914
rect 50517 4850 50518 4914
rect 50452 4834 50518 4850
rect 50452 4770 50453 4834
rect 50517 4770 50518 4834
rect 50452 4754 50518 4770
rect 50452 4690 50453 4754
rect 50517 4690 50518 4754
rect 50452 4674 50518 4690
rect 50452 4610 50453 4674
rect 50517 4610 50518 4674
rect 50452 4594 50518 4610
rect 50452 4530 50453 4594
rect 50517 4530 50518 4594
rect 50452 4514 50518 4530
rect 50452 4450 50453 4514
rect 50517 4450 50518 4514
rect 50452 4434 50518 4450
rect 50452 4370 50453 4434
rect 50517 4370 50518 4434
rect 50452 4354 50518 4370
rect 50452 4290 50453 4354
rect 50517 4290 50518 4354
rect 50452 4274 50518 4290
rect 50452 4210 50453 4274
rect 50517 4210 50518 4274
rect 50452 4120 50518 4210
rect 50578 4116 50638 5148
rect 50698 4056 50758 5086
rect 50818 4116 50878 5148
rect 50938 4056 50998 5086
rect 51058 4994 51124 5148
rect 51058 4930 51059 4994
rect 51123 4930 51124 4994
rect 51058 4914 51124 4930
rect 51058 4850 51059 4914
rect 51123 4850 51124 4914
rect 51058 4834 51124 4850
rect 51058 4770 51059 4834
rect 51123 4770 51124 4834
rect 51058 4754 51124 4770
rect 51058 4690 51059 4754
rect 51123 4690 51124 4754
rect 51058 4674 51124 4690
rect 51058 4610 51059 4674
rect 51123 4610 51124 4674
rect 51058 4594 51124 4610
rect 51058 4530 51059 4594
rect 51123 4530 51124 4594
rect 51058 4514 51124 4530
rect 51058 4450 51059 4514
rect 51123 4450 51124 4514
rect 51058 4434 51124 4450
rect 51058 4370 51059 4434
rect 51123 4370 51124 4434
rect 51058 4354 51124 4370
rect 51058 4290 51059 4354
rect 51123 4290 51124 4354
rect 51058 4274 51124 4290
rect 51058 4210 51059 4274
rect 51123 4210 51124 4274
rect 51058 4120 51124 4210
rect 51184 4116 51244 5148
rect 51304 4056 51364 5086
rect 51424 4116 51484 5148
rect 51544 4056 51604 5086
rect 51664 4994 51730 5148
rect 51664 4930 51665 4994
rect 51729 4930 51730 4994
rect 51664 4914 51730 4930
rect 51664 4850 51665 4914
rect 51729 4850 51730 4914
rect 51664 4834 51730 4850
rect 51664 4770 51665 4834
rect 51729 4770 51730 4834
rect 51664 4754 51730 4770
rect 51664 4690 51665 4754
rect 51729 4690 51730 4754
rect 51664 4674 51730 4690
rect 51664 4610 51665 4674
rect 51729 4610 51730 4674
rect 51664 4594 51730 4610
rect 51664 4530 51665 4594
rect 51729 4530 51730 4594
rect 51664 4514 51730 4530
rect 51664 4450 51665 4514
rect 51729 4450 51730 4514
rect 51664 4434 51730 4450
rect 51664 4370 51665 4434
rect 51729 4370 51730 4434
rect 51664 4354 51730 4370
rect 51664 4290 51665 4354
rect 51729 4290 51730 4354
rect 51664 4274 51730 4290
rect 51664 4210 51665 4274
rect 51729 4210 51730 4274
rect 51664 4120 51730 4210
rect 32272 4054 51730 4056
rect 32272 3990 32376 4054
rect 32440 3990 32456 4054
rect 32520 3990 32536 4054
rect 32600 3990 32616 4054
rect 32680 3990 32696 4054
rect 32760 3990 32776 4054
rect 32840 3990 32982 4054
rect 33046 3990 33062 4054
rect 33126 3990 33142 4054
rect 33206 3990 33222 4054
rect 33286 3990 33302 4054
rect 33366 3990 33382 4054
rect 33446 3990 33588 4054
rect 33652 3990 33668 4054
rect 33732 3990 33748 4054
rect 33812 3990 33828 4054
rect 33892 3990 33908 4054
rect 33972 3990 33988 4054
rect 34052 3990 34194 4054
rect 34258 3990 34274 4054
rect 34338 3990 34354 4054
rect 34418 3990 34434 4054
rect 34498 3990 34514 4054
rect 34578 3990 34594 4054
rect 34658 3990 34800 4054
rect 34864 3990 34880 4054
rect 34944 3990 34960 4054
rect 35024 3990 35040 4054
rect 35104 3990 35120 4054
rect 35184 3990 35200 4054
rect 35264 3990 35406 4054
rect 35470 3990 35486 4054
rect 35550 3990 35566 4054
rect 35630 3990 35646 4054
rect 35710 3990 35726 4054
rect 35790 3990 35806 4054
rect 35870 3990 36012 4054
rect 36076 3990 36092 4054
rect 36156 3990 36172 4054
rect 36236 3990 36252 4054
rect 36316 3990 36332 4054
rect 36396 3990 36412 4054
rect 36476 3990 36618 4054
rect 36682 3990 36698 4054
rect 36762 3990 36778 4054
rect 36842 3990 36858 4054
rect 36922 3990 36938 4054
rect 37002 3990 37018 4054
rect 37082 3990 37224 4054
rect 37288 3990 37304 4054
rect 37368 3990 37384 4054
rect 37448 3990 37464 4054
rect 37528 3990 37544 4054
rect 37608 3990 37624 4054
rect 37688 3990 37830 4054
rect 37894 3990 37910 4054
rect 37974 3990 37990 4054
rect 38054 3990 38070 4054
rect 38134 3990 38150 4054
rect 38214 3990 38230 4054
rect 38294 3990 38436 4054
rect 38500 3990 38516 4054
rect 38580 3990 38596 4054
rect 38660 3990 38676 4054
rect 38740 3990 38756 4054
rect 38820 3990 38836 4054
rect 38900 3990 39042 4054
rect 39106 3990 39122 4054
rect 39186 3990 39202 4054
rect 39266 3990 39282 4054
rect 39346 3990 39362 4054
rect 39426 3990 39442 4054
rect 39506 3990 39648 4054
rect 39712 3990 39728 4054
rect 39792 3990 39808 4054
rect 39872 3990 39888 4054
rect 39952 3990 39968 4054
rect 40032 3990 40048 4054
rect 40112 3990 40254 4054
rect 40318 3990 40334 4054
rect 40398 3990 40414 4054
rect 40478 3990 40494 4054
rect 40558 3990 40574 4054
rect 40638 3990 40654 4054
rect 40718 3990 40860 4054
rect 40924 3990 40940 4054
rect 41004 3990 41020 4054
rect 41084 3990 41100 4054
rect 41164 3990 41180 4054
rect 41244 3990 41260 4054
rect 41324 3990 41466 4054
rect 41530 3990 41546 4054
rect 41610 3990 41626 4054
rect 41690 3990 41706 4054
rect 41770 3990 41786 4054
rect 41850 3990 41866 4054
rect 41930 3990 42072 4054
rect 42136 3990 42152 4054
rect 42216 3990 42232 4054
rect 42296 3990 42312 4054
rect 42376 3990 42392 4054
rect 42456 3990 42472 4054
rect 42536 3990 42678 4054
rect 42742 3990 42758 4054
rect 42822 3990 42838 4054
rect 42902 3990 42918 4054
rect 42982 3990 42998 4054
rect 43062 3990 43078 4054
rect 43142 3990 43284 4054
rect 43348 3990 43364 4054
rect 43428 3990 43444 4054
rect 43508 3990 43524 4054
rect 43588 3990 43604 4054
rect 43668 3990 43684 4054
rect 43748 3990 43890 4054
rect 43954 3990 43970 4054
rect 44034 3990 44050 4054
rect 44114 3990 44130 4054
rect 44194 3990 44210 4054
rect 44274 3990 44290 4054
rect 44354 3990 44496 4054
rect 44560 3990 44576 4054
rect 44640 3990 44656 4054
rect 44720 3990 44736 4054
rect 44800 3990 44816 4054
rect 44880 3990 44896 4054
rect 44960 3990 45102 4054
rect 45166 3990 45182 4054
rect 45246 3990 45262 4054
rect 45326 3990 45342 4054
rect 45406 3990 45422 4054
rect 45486 3990 45502 4054
rect 45566 3990 45708 4054
rect 45772 3990 45788 4054
rect 45852 3990 45868 4054
rect 45932 3990 45948 4054
rect 46012 3990 46028 4054
rect 46092 3990 46108 4054
rect 46172 3990 46314 4054
rect 46378 3990 46394 4054
rect 46458 3990 46474 4054
rect 46538 3990 46554 4054
rect 46618 3990 46634 4054
rect 46698 3990 46714 4054
rect 46778 3990 46920 4054
rect 46984 3990 47000 4054
rect 47064 3990 47080 4054
rect 47144 3990 47160 4054
rect 47224 3990 47240 4054
rect 47304 3990 47320 4054
rect 47384 3990 47526 4054
rect 47590 3990 47606 4054
rect 47670 3990 47686 4054
rect 47750 3990 47766 4054
rect 47830 3990 47846 4054
rect 47910 3990 47926 4054
rect 47990 3990 48132 4054
rect 48196 3990 48212 4054
rect 48276 3990 48292 4054
rect 48356 3990 48372 4054
rect 48436 3990 48452 4054
rect 48516 3990 48532 4054
rect 48596 3990 48738 4054
rect 48802 3990 48818 4054
rect 48882 3990 48898 4054
rect 48962 3990 48978 4054
rect 49042 3990 49058 4054
rect 49122 3990 49138 4054
rect 49202 3990 49344 4054
rect 49408 3990 49424 4054
rect 49488 3990 49504 4054
rect 49568 3990 49584 4054
rect 49648 3990 49664 4054
rect 49728 3990 49744 4054
rect 49808 3990 49950 4054
rect 50014 3990 50030 4054
rect 50094 3990 50110 4054
rect 50174 3990 50190 4054
rect 50254 3990 50270 4054
rect 50334 3990 50350 4054
rect 50414 3990 50556 4054
rect 50620 3990 50636 4054
rect 50700 3990 50716 4054
rect 50780 3990 50796 4054
rect 50860 3990 50876 4054
rect 50940 3990 50956 4054
rect 51020 3990 51162 4054
rect 51226 3990 51242 4054
rect 51306 3990 51322 4054
rect 51386 3990 51402 4054
rect 51466 3990 51482 4054
rect 51546 3990 51562 4054
rect 51626 3990 51730 4054
rect 32272 3988 51730 3990
rect 32272 3834 32338 3988
rect 32272 3770 32273 3834
rect 32337 3770 32338 3834
rect 32272 3754 32338 3770
rect 32272 3690 32273 3754
rect 32337 3690 32338 3754
rect 32272 3674 32338 3690
rect 32272 3610 32273 3674
rect 32337 3610 32338 3674
rect 32272 3594 32338 3610
rect 32272 3530 32273 3594
rect 32337 3530 32338 3594
rect 32272 3514 32338 3530
rect 32272 3450 32273 3514
rect 32337 3450 32338 3514
rect 32272 3434 32338 3450
rect 32272 3370 32273 3434
rect 32337 3370 32338 3434
rect 32272 3354 32338 3370
rect 32272 3290 32273 3354
rect 32337 3290 32338 3354
rect 32272 3274 32338 3290
rect 32272 3210 32273 3274
rect 32337 3210 32338 3274
rect 32272 3194 32338 3210
rect 32272 3130 32273 3194
rect 32337 3130 32338 3194
rect 32272 3114 32338 3130
rect 32272 3050 32273 3114
rect 32337 3050 32338 3114
rect 32272 2960 32338 3050
rect 32398 2956 32458 3988
rect 32518 2896 32578 3926
rect 32638 2956 32698 3988
rect 32758 2896 32818 3926
rect 32878 3834 32944 3988
rect 32878 3770 32879 3834
rect 32943 3770 32944 3834
rect 32878 3754 32944 3770
rect 32878 3690 32879 3754
rect 32943 3690 32944 3754
rect 32878 3674 32944 3690
rect 32878 3610 32879 3674
rect 32943 3610 32944 3674
rect 32878 3594 32944 3610
rect 32878 3530 32879 3594
rect 32943 3530 32944 3594
rect 32878 3514 32944 3530
rect 32878 3450 32879 3514
rect 32943 3450 32944 3514
rect 32878 3434 32944 3450
rect 32878 3370 32879 3434
rect 32943 3370 32944 3434
rect 32878 3354 32944 3370
rect 32878 3290 32879 3354
rect 32943 3290 32944 3354
rect 32878 3274 32944 3290
rect 32878 3210 32879 3274
rect 32943 3210 32944 3274
rect 32878 3194 32944 3210
rect 32878 3130 32879 3194
rect 32943 3130 32944 3194
rect 32878 3114 32944 3130
rect 32878 3050 32879 3114
rect 32943 3050 32944 3114
rect 32878 2960 32944 3050
rect 33004 2956 33064 3988
rect 33124 2896 33184 3926
rect 33244 2956 33304 3988
rect 33364 2896 33424 3926
rect 33484 3834 33550 3988
rect 33484 3770 33485 3834
rect 33549 3770 33550 3834
rect 33484 3754 33550 3770
rect 33484 3690 33485 3754
rect 33549 3690 33550 3754
rect 33484 3674 33550 3690
rect 33484 3610 33485 3674
rect 33549 3610 33550 3674
rect 33484 3594 33550 3610
rect 33484 3530 33485 3594
rect 33549 3530 33550 3594
rect 33484 3514 33550 3530
rect 33484 3450 33485 3514
rect 33549 3450 33550 3514
rect 33484 3434 33550 3450
rect 33484 3370 33485 3434
rect 33549 3370 33550 3434
rect 33484 3354 33550 3370
rect 33484 3290 33485 3354
rect 33549 3290 33550 3354
rect 33484 3274 33550 3290
rect 33484 3210 33485 3274
rect 33549 3210 33550 3274
rect 33484 3194 33550 3210
rect 33484 3130 33485 3194
rect 33549 3130 33550 3194
rect 33484 3114 33550 3130
rect 33484 3050 33485 3114
rect 33549 3050 33550 3114
rect 33484 2960 33550 3050
rect 33610 2956 33670 3988
rect 33730 2896 33790 3926
rect 33850 2956 33910 3988
rect 33970 2896 34030 3926
rect 34090 3834 34156 3988
rect 34090 3770 34091 3834
rect 34155 3770 34156 3834
rect 34090 3754 34156 3770
rect 34090 3690 34091 3754
rect 34155 3690 34156 3754
rect 34090 3674 34156 3690
rect 34090 3610 34091 3674
rect 34155 3610 34156 3674
rect 34090 3594 34156 3610
rect 34090 3530 34091 3594
rect 34155 3530 34156 3594
rect 34090 3514 34156 3530
rect 34090 3450 34091 3514
rect 34155 3450 34156 3514
rect 34090 3434 34156 3450
rect 34090 3370 34091 3434
rect 34155 3370 34156 3434
rect 34090 3354 34156 3370
rect 34090 3290 34091 3354
rect 34155 3290 34156 3354
rect 34090 3274 34156 3290
rect 34090 3210 34091 3274
rect 34155 3210 34156 3274
rect 34090 3194 34156 3210
rect 34090 3130 34091 3194
rect 34155 3130 34156 3194
rect 34090 3114 34156 3130
rect 34090 3050 34091 3114
rect 34155 3050 34156 3114
rect 34090 2960 34156 3050
rect 34216 2956 34276 3988
rect 34336 2896 34396 3926
rect 34456 2956 34516 3988
rect 34576 2896 34636 3926
rect 34696 3834 34762 3988
rect 34696 3770 34697 3834
rect 34761 3770 34762 3834
rect 34696 3754 34762 3770
rect 34696 3690 34697 3754
rect 34761 3690 34762 3754
rect 34696 3674 34762 3690
rect 34696 3610 34697 3674
rect 34761 3610 34762 3674
rect 34696 3594 34762 3610
rect 34696 3530 34697 3594
rect 34761 3530 34762 3594
rect 34696 3514 34762 3530
rect 34696 3450 34697 3514
rect 34761 3450 34762 3514
rect 34696 3434 34762 3450
rect 34696 3370 34697 3434
rect 34761 3370 34762 3434
rect 34696 3354 34762 3370
rect 34696 3290 34697 3354
rect 34761 3290 34762 3354
rect 34696 3274 34762 3290
rect 34696 3210 34697 3274
rect 34761 3210 34762 3274
rect 34696 3194 34762 3210
rect 34696 3130 34697 3194
rect 34761 3130 34762 3194
rect 34696 3114 34762 3130
rect 34696 3050 34697 3114
rect 34761 3050 34762 3114
rect 34696 2960 34762 3050
rect 34822 2956 34882 3988
rect 34942 2896 35002 3926
rect 35062 2956 35122 3988
rect 35182 2896 35242 3926
rect 35302 3834 35368 3988
rect 35302 3770 35303 3834
rect 35367 3770 35368 3834
rect 35302 3754 35368 3770
rect 35302 3690 35303 3754
rect 35367 3690 35368 3754
rect 35302 3674 35368 3690
rect 35302 3610 35303 3674
rect 35367 3610 35368 3674
rect 35302 3594 35368 3610
rect 35302 3530 35303 3594
rect 35367 3530 35368 3594
rect 35302 3514 35368 3530
rect 35302 3450 35303 3514
rect 35367 3450 35368 3514
rect 35302 3434 35368 3450
rect 35302 3370 35303 3434
rect 35367 3370 35368 3434
rect 35302 3354 35368 3370
rect 35302 3290 35303 3354
rect 35367 3290 35368 3354
rect 35302 3274 35368 3290
rect 35302 3210 35303 3274
rect 35367 3210 35368 3274
rect 35302 3194 35368 3210
rect 35302 3130 35303 3194
rect 35367 3130 35368 3194
rect 35302 3114 35368 3130
rect 35302 3050 35303 3114
rect 35367 3050 35368 3114
rect 35302 2960 35368 3050
rect 35428 2956 35488 3988
rect 35548 2896 35608 3926
rect 35668 2956 35728 3988
rect 35788 2896 35848 3926
rect 35908 3834 35974 3988
rect 35908 3770 35909 3834
rect 35973 3770 35974 3834
rect 35908 3754 35974 3770
rect 35908 3690 35909 3754
rect 35973 3690 35974 3754
rect 35908 3674 35974 3690
rect 35908 3610 35909 3674
rect 35973 3610 35974 3674
rect 35908 3594 35974 3610
rect 35908 3530 35909 3594
rect 35973 3530 35974 3594
rect 35908 3514 35974 3530
rect 35908 3450 35909 3514
rect 35973 3450 35974 3514
rect 35908 3434 35974 3450
rect 35908 3370 35909 3434
rect 35973 3370 35974 3434
rect 35908 3354 35974 3370
rect 35908 3290 35909 3354
rect 35973 3290 35974 3354
rect 35908 3274 35974 3290
rect 35908 3210 35909 3274
rect 35973 3210 35974 3274
rect 35908 3194 35974 3210
rect 35908 3130 35909 3194
rect 35973 3130 35974 3194
rect 35908 3114 35974 3130
rect 35908 3050 35909 3114
rect 35973 3050 35974 3114
rect 35908 2960 35974 3050
rect 36034 2956 36094 3988
rect 36154 2896 36214 3926
rect 36274 2956 36334 3988
rect 36394 2896 36454 3926
rect 36514 3834 36580 3988
rect 36514 3770 36515 3834
rect 36579 3770 36580 3834
rect 36514 3754 36580 3770
rect 36514 3690 36515 3754
rect 36579 3690 36580 3754
rect 36514 3674 36580 3690
rect 36514 3610 36515 3674
rect 36579 3610 36580 3674
rect 36514 3594 36580 3610
rect 36514 3530 36515 3594
rect 36579 3530 36580 3594
rect 36514 3514 36580 3530
rect 36514 3450 36515 3514
rect 36579 3450 36580 3514
rect 36514 3434 36580 3450
rect 36514 3370 36515 3434
rect 36579 3370 36580 3434
rect 36514 3354 36580 3370
rect 36514 3290 36515 3354
rect 36579 3290 36580 3354
rect 36514 3274 36580 3290
rect 36514 3210 36515 3274
rect 36579 3210 36580 3274
rect 36514 3194 36580 3210
rect 36514 3130 36515 3194
rect 36579 3130 36580 3194
rect 36514 3114 36580 3130
rect 36514 3050 36515 3114
rect 36579 3050 36580 3114
rect 36514 2960 36580 3050
rect 36640 2956 36700 3988
rect 36760 2896 36820 3926
rect 36880 2956 36940 3988
rect 37000 2896 37060 3926
rect 37120 3834 37186 3988
rect 37120 3770 37121 3834
rect 37185 3770 37186 3834
rect 37120 3754 37186 3770
rect 37120 3690 37121 3754
rect 37185 3690 37186 3754
rect 37120 3674 37186 3690
rect 37120 3610 37121 3674
rect 37185 3610 37186 3674
rect 37120 3594 37186 3610
rect 37120 3530 37121 3594
rect 37185 3530 37186 3594
rect 37120 3514 37186 3530
rect 37120 3450 37121 3514
rect 37185 3450 37186 3514
rect 37120 3434 37186 3450
rect 37120 3370 37121 3434
rect 37185 3370 37186 3434
rect 37120 3354 37186 3370
rect 37120 3290 37121 3354
rect 37185 3290 37186 3354
rect 37120 3274 37186 3290
rect 37120 3210 37121 3274
rect 37185 3210 37186 3274
rect 37120 3194 37186 3210
rect 37120 3130 37121 3194
rect 37185 3130 37186 3194
rect 37120 3114 37186 3130
rect 37120 3050 37121 3114
rect 37185 3050 37186 3114
rect 37120 2960 37186 3050
rect 37246 2956 37306 3988
rect 37366 2896 37426 3926
rect 37486 2956 37546 3988
rect 37606 2896 37666 3926
rect 37726 3834 37792 3988
rect 37726 3770 37727 3834
rect 37791 3770 37792 3834
rect 37726 3754 37792 3770
rect 37726 3690 37727 3754
rect 37791 3690 37792 3754
rect 37726 3674 37792 3690
rect 37726 3610 37727 3674
rect 37791 3610 37792 3674
rect 37726 3594 37792 3610
rect 37726 3530 37727 3594
rect 37791 3530 37792 3594
rect 37726 3514 37792 3530
rect 37726 3450 37727 3514
rect 37791 3450 37792 3514
rect 37726 3434 37792 3450
rect 37726 3370 37727 3434
rect 37791 3370 37792 3434
rect 37726 3354 37792 3370
rect 37726 3290 37727 3354
rect 37791 3290 37792 3354
rect 37726 3274 37792 3290
rect 37726 3210 37727 3274
rect 37791 3210 37792 3274
rect 37726 3194 37792 3210
rect 37726 3130 37727 3194
rect 37791 3130 37792 3194
rect 37726 3114 37792 3130
rect 37726 3050 37727 3114
rect 37791 3050 37792 3114
rect 37726 2960 37792 3050
rect 37852 2956 37912 3988
rect 37972 2896 38032 3926
rect 38092 2956 38152 3988
rect 38212 2896 38272 3926
rect 38332 3834 38398 3988
rect 38332 3770 38333 3834
rect 38397 3770 38398 3834
rect 38332 3754 38398 3770
rect 38332 3690 38333 3754
rect 38397 3690 38398 3754
rect 38332 3674 38398 3690
rect 38332 3610 38333 3674
rect 38397 3610 38398 3674
rect 38332 3594 38398 3610
rect 38332 3530 38333 3594
rect 38397 3530 38398 3594
rect 38332 3514 38398 3530
rect 38332 3450 38333 3514
rect 38397 3450 38398 3514
rect 38332 3434 38398 3450
rect 38332 3370 38333 3434
rect 38397 3370 38398 3434
rect 38332 3354 38398 3370
rect 38332 3290 38333 3354
rect 38397 3290 38398 3354
rect 38332 3274 38398 3290
rect 38332 3210 38333 3274
rect 38397 3210 38398 3274
rect 38332 3194 38398 3210
rect 38332 3130 38333 3194
rect 38397 3130 38398 3194
rect 38332 3114 38398 3130
rect 38332 3050 38333 3114
rect 38397 3050 38398 3114
rect 38332 2960 38398 3050
rect 38458 2956 38518 3988
rect 38578 2896 38638 3926
rect 38698 2956 38758 3988
rect 38818 2896 38878 3926
rect 38938 3834 39004 3988
rect 38938 3770 38939 3834
rect 39003 3770 39004 3834
rect 38938 3754 39004 3770
rect 38938 3690 38939 3754
rect 39003 3690 39004 3754
rect 38938 3674 39004 3690
rect 38938 3610 38939 3674
rect 39003 3610 39004 3674
rect 38938 3594 39004 3610
rect 38938 3530 38939 3594
rect 39003 3530 39004 3594
rect 38938 3514 39004 3530
rect 38938 3450 38939 3514
rect 39003 3450 39004 3514
rect 38938 3434 39004 3450
rect 38938 3370 38939 3434
rect 39003 3370 39004 3434
rect 38938 3354 39004 3370
rect 38938 3290 38939 3354
rect 39003 3290 39004 3354
rect 38938 3274 39004 3290
rect 38938 3210 38939 3274
rect 39003 3210 39004 3274
rect 38938 3194 39004 3210
rect 38938 3130 38939 3194
rect 39003 3130 39004 3194
rect 38938 3114 39004 3130
rect 38938 3050 38939 3114
rect 39003 3050 39004 3114
rect 38938 2960 39004 3050
rect 39064 2956 39124 3988
rect 39184 2896 39244 3926
rect 39304 2956 39364 3988
rect 39424 2896 39484 3926
rect 39544 3834 39610 3988
rect 39544 3770 39545 3834
rect 39609 3770 39610 3834
rect 39544 3754 39610 3770
rect 39544 3690 39545 3754
rect 39609 3690 39610 3754
rect 39544 3674 39610 3690
rect 39544 3610 39545 3674
rect 39609 3610 39610 3674
rect 39544 3594 39610 3610
rect 39544 3530 39545 3594
rect 39609 3530 39610 3594
rect 39544 3514 39610 3530
rect 39544 3450 39545 3514
rect 39609 3450 39610 3514
rect 39544 3434 39610 3450
rect 39544 3370 39545 3434
rect 39609 3370 39610 3434
rect 39544 3354 39610 3370
rect 39544 3290 39545 3354
rect 39609 3290 39610 3354
rect 39544 3274 39610 3290
rect 39544 3210 39545 3274
rect 39609 3210 39610 3274
rect 39544 3194 39610 3210
rect 39544 3130 39545 3194
rect 39609 3130 39610 3194
rect 39544 3114 39610 3130
rect 39544 3050 39545 3114
rect 39609 3050 39610 3114
rect 39544 2960 39610 3050
rect 39670 2956 39730 3988
rect 39790 2896 39850 3926
rect 39910 2956 39970 3988
rect 40030 2896 40090 3926
rect 40150 3834 40216 3988
rect 40150 3770 40151 3834
rect 40215 3770 40216 3834
rect 40150 3754 40216 3770
rect 40150 3690 40151 3754
rect 40215 3690 40216 3754
rect 40150 3674 40216 3690
rect 40150 3610 40151 3674
rect 40215 3610 40216 3674
rect 40150 3594 40216 3610
rect 40150 3530 40151 3594
rect 40215 3530 40216 3594
rect 40150 3514 40216 3530
rect 40150 3450 40151 3514
rect 40215 3450 40216 3514
rect 40150 3434 40216 3450
rect 40150 3370 40151 3434
rect 40215 3370 40216 3434
rect 40150 3354 40216 3370
rect 40150 3290 40151 3354
rect 40215 3290 40216 3354
rect 40150 3274 40216 3290
rect 40150 3210 40151 3274
rect 40215 3210 40216 3274
rect 40150 3194 40216 3210
rect 40150 3130 40151 3194
rect 40215 3130 40216 3194
rect 40150 3114 40216 3130
rect 40150 3050 40151 3114
rect 40215 3050 40216 3114
rect 40150 2960 40216 3050
rect 40276 2956 40336 3988
rect 40396 2896 40456 3926
rect 40516 2956 40576 3988
rect 40636 2896 40696 3926
rect 40756 3834 40822 3988
rect 40756 3770 40757 3834
rect 40821 3770 40822 3834
rect 40756 3754 40822 3770
rect 40756 3690 40757 3754
rect 40821 3690 40822 3754
rect 40756 3674 40822 3690
rect 40756 3610 40757 3674
rect 40821 3610 40822 3674
rect 40756 3594 40822 3610
rect 40756 3530 40757 3594
rect 40821 3530 40822 3594
rect 40756 3514 40822 3530
rect 40756 3450 40757 3514
rect 40821 3450 40822 3514
rect 40756 3434 40822 3450
rect 40756 3370 40757 3434
rect 40821 3370 40822 3434
rect 40756 3354 40822 3370
rect 40756 3290 40757 3354
rect 40821 3290 40822 3354
rect 40756 3274 40822 3290
rect 40756 3210 40757 3274
rect 40821 3210 40822 3274
rect 40756 3194 40822 3210
rect 40756 3130 40757 3194
rect 40821 3130 40822 3194
rect 40756 3114 40822 3130
rect 40756 3050 40757 3114
rect 40821 3050 40822 3114
rect 40756 2960 40822 3050
rect 40882 2956 40942 3988
rect 41002 2896 41062 3926
rect 41122 2956 41182 3988
rect 41242 2896 41302 3926
rect 41362 3834 41428 3988
rect 41362 3770 41363 3834
rect 41427 3770 41428 3834
rect 41362 3754 41428 3770
rect 41362 3690 41363 3754
rect 41427 3690 41428 3754
rect 41362 3674 41428 3690
rect 41362 3610 41363 3674
rect 41427 3610 41428 3674
rect 41362 3594 41428 3610
rect 41362 3530 41363 3594
rect 41427 3530 41428 3594
rect 41362 3514 41428 3530
rect 41362 3450 41363 3514
rect 41427 3450 41428 3514
rect 41362 3434 41428 3450
rect 41362 3370 41363 3434
rect 41427 3370 41428 3434
rect 41362 3354 41428 3370
rect 41362 3290 41363 3354
rect 41427 3290 41428 3354
rect 41362 3274 41428 3290
rect 41362 3210 41363 3274
rect 41427 3210 41428 3274
rect 41362 3194 41428 3210
rect 41362 3130 41363 3194
rect 41427 3130 41428 3194
rect 41362 3114 41428 3130
rect 41362 3050 41363 3114
rect 41427 3050 41428 3114
rect 41362 2960 41428 3050
rect 41488 2956 41548 3988
rect 41608 2896 41668 3926
rect 41728 2956 41788 3988
rect 41848 2896 41908 3926
rect 41968 3834 42034 3988
rect 41968 3770 41969 3834
rect 42033 3770 42034 3834
rect 41968 3754 42034 3770
rect 41968 3690 41969 3754
rect 42033 3690 42034 3754
rect 41968 3674 42034 3690
rect 41968 3610 41969 3674
rect 42033 3610 42034 3674
rect 41968 3594 42034 3610
rect 41968 3530 41969 3594
rect 42033 3530 42034 3594
rect 41968 3514 42034 3530
rect 41968 3450 41969 3514
rect 42033 3450 42034 3514
rect 41968 3434 42034 3450
rect 41968 3370 41969 3434
rect 42033 3370 42034 3434
rect 41968 3354 42034 3370
rect 41968 3290 41969 3354
rect 42033 3290 42034 3354
rect 41968 3274 42034 3290
rect 41968 3210 41969 3274
rect 42033 3210 42034 3274
rect 41968 3194 42034 3210
rect 41968 3130 41969 3194
rect 42033 3130 42034 3194
rect 41968 3114 42034 3130
rect 41968 3050 41969 3114
rect 42033 3050 42034 3114
rect 41968 2960 42034 3050
rect 42094 2956 42154 3988
rect 42214 2896 42274 3926
rect 42334 2956 42394 3988
rect 42454 2896 42514 3926
rect 42574 3834 42640 3988
rect 42574 3770 42575 3834
rect 42639 3770 42640 3834
rect 42574 3754 42640 3770
rect 42574 3690 42575 3754
rect 42639 3690 42640 3754
rect 42574 3674 42640 3690
rect 42574 3610 42575 3674
rect 42639 3610 42640 3674
rect 42574 3594 42640 3610
rect 42574 3530 42575 3594
rect 42639 3530 42640 3594
rect 42574 3514 42640 3530
rect 42574 3450 42575 3514
rect 42639 3450 42640 3514
rect 42574 3434 42640 3450
rect 42574 3370 42575 3434
rect 42639 3370 42640 3434
rect 42574 3354 42640 3370
rect 42574 3290 42575 3354
rect 42639 3290 42640 3354
rect 42574 3274 42640 3290
rect 42574 3210 42575 3274
rect 42639 3210 42640 3274
rect 42574 3194 42640 3210
rect 42574 3130 42575 3194
rect 42639 3130 42640 3194
rect 42574 3114 42640 3130
rect 42574 3050 42575 3114
rect 42639 3050 42640 3114
rect 42574 2960 42640 3050
rect 42700 2956 42760 3988
rect 42820 2896 42880 3926
rect 42940 2956 43000 3988
rect 43060 2896 43120 3926
rect 43180 3834 43246 3988
rect 43180 3770 43181 3834
rect 43245 3770 43246 3834
rect 43180 3754 43246 3770
rect 43180 3690 43181 3754
rect 43245 3690 43246 3754
rect 43180 3674 43246 3690
rect 43180 3610 43181 3674
rect 43245 3610 43246 3674
rect 43180 3594 43246 3610
rect 43180 3530 43181 3594
rect 43245 3530 43246 3594
rect 43180 3514 43246 3530
rect 43180 3450 43181 3514
rect 43245 3450 43246 3514
rect 43180 3434 43246 3450
rect 43180 3370 43181 3434
rect 43245 3370 43246 3434
rect 43180 3354 43246 3370
rect 43180 3290 43181 3354
rect 43245 3290 43246 3354
rect 43180 3274 43246 3290
rect 43180 3210 43181 3274
rect 43245 3210 43246 3274
rect 43180 3194 43246 3210
rect 43180 3130 43181 3194
rect 43245 3130 43246 3194
rect 43180 3114 43246 3130
rect 43180 3050 43181 3114
rect 43245 3050 43246 3114
rect 43180 2960 43246 3050
rect 43306 2956 43366 3988
rect 43426 2896 43486 3926
rect 43546 2956 43606 3988
rect 43666 2896 43726 3926
rect 43786 3834 43852 3988
rect 43786 3770 43787 3834
rect 43851 3770 43852 3834
rect 43786 3754 43852 3770
rect 43786 3690 43787 3754
rect 43851 3690 43852 3754
rect 43786 3674 43852 3690
rect 43786 3610 43787 3674
rect 43851 3610 43852 3674
rect 43786 3594 43852 3610
rect 43786 3530 43787 3594
rect 43851 3530 43852 3594
rect 43786 3514 43852 3530
rect 43786 3450 43787 3514
rect 43851 3450 43852 3514
rect 43786 3434 43852 3450
rect 43786 3370 43787 3434
rect 43851 3370 43852 3434
rect 43786 3354 43852 3370
rect 43786 3290 43787 3354
rect 43851 3290 43852 3354
rect 43786 3274 43852 3290
rect 43786 3210 43787 3274
rect 43851 3210 43852 3274
rect 43786 3194 43852 3210
rect 43786 3130 43787 3194
rect 43851 3130 43852 3194
rect 43786 3114 43852 3130
rect 43786 3050 43787 3114
rect 43851 3050 43852 3114
rect 43786 2960 43852 3050
rect 43912 2956 43972 3988
rect 44032 2896 44092 3926
rect 44152 2956 44212 3988
rect 44272 2896 44332 3926
rect 44392 3834 44458 3988
rect 44392 3770 44393 3834
rect 44457 3770 44458 3834
rect 44392 3754 44458 3770
rect 44392 3690 44393 3754
rect 44457 3690 44458 3754
rect 44392 3674 44458 3690
rect 44392 3610 44393 3674
rect 44457 3610 44458 3674
rect 44392 3594 44458 3610
rect 44392 3530 44393 3594
rect 44457 3530 44458 3594
rect 44392 3514 44458 3530
rect 44392 3450 44393 3514
rect 44457 3450 44458 3514
rect 44392 3434 44458 3450
rect 44392 3370 44393 3434
rect 44457 3370 44458 3434
rect 44392 3354 44458 3370
rect 44392 3290 44393 3354
rect 44457 3290 44458 3354
rect 44392 3274 44458 3290
rect 44392 3210 44393 3274
rect 44457 3210 44458 3274
rect 44392 3194 44458 3210
rect 44392 3130 44393 3194
rect 44457 3130 44458 3194
rect 44392 3114 44458 3130
rect 44392 3050 44393 3114
rect 44457 3050 44458 3114
rect 44392 2960 44458 3050
rect 44518 2956 44578 3988
rect 44638 2896 44698 3926
rect 44758 2956 44818 3988
rect 44878 2896 44938 3926
rect 44998 3834 45064 3988
rect 44998 3770 44999 3834
rect 45063 3770 45064 3834
rect 44998 3754 45064 3770
rect 44998 3690 44999 3754
rect 45063 3690 45064 3754
rect 44998 3674 45064 3690
rect 44998 3610 44999 3674
rect 45063 3610 45064 3674
rect 44998 3594 45064 3610
rect 44998 3530 44999 3594
rect 45063 3530 45064 3594
rect 44998 3514 45064 3530
rect 44998 3450 44999 3514
rect 45063 3450 45064 3514
rect 44998 3434 45064 3450
rect 44998 3370 44999 3434
rect 45063 3370 45064 3434
rect 44998 3354 45064 3370
rect 44998 3290 44999 3354
rect 45063 3290 45064 3354
rect 44998 3274 45064 3290
rect 44998 3210 44999 3274
rect 45063 3210 45064 3274
rect 44998 3194 45064 3210
rect 44998 3130 44999 3194
rect 45063 3130 45064 3194
rect 44998 3114 45064 3130
rect 44998 3050 44999 3114
rect 45063 3050 45064 3114
rect 44998 2960 45064 3050
rect 45124 2956 45184 3988
rect 45244 2896 45304 3926
rect 45364 2956 45424 3988
rect 45484 2896 45544 3926
rect 45604 3834 45670 3988
rect 45604 3770 45605 3834
rect 45669 3770 45670 3834
rect 45604 3754 45670 3770
rect 45604 3690 45605 3754
rect 45669 3690 45670 3754
rect 45604 3674 45670 3690
rect 45604 3610 45605 3674
rect 45669 3610 45670 3674
rect 45604 3594 45670 3610
rect 45604 3530 45605 3594
rect 45669 3530 45670 3594
rect 45604 3514 45670 3530
rect 45604 3450 45605 3514
rect 45669 3450 45670 3514
rect 45604 3434 45670 3450
rect 45604 3370 45605 3434
rect 45669 3370 45670 3434
rect 45604 3354 45670 3370
rect 45604 3290 45605 3354
rect 45669 3290 45670 3354
rect 45604 3274 45670 3290
rect 45604 3210 45605 3274
rect 45669 3210 45670 3274
rect 45604 3194 45670 3210
rect 45604 3130 45605 3194
rect 45669 3130 45670 3194
rect 45604 3114 45670 3130
rect 45604 3050 45605 3114
rect 45669 3050 45670 3114
rect 45604 2960 45670 3050
rect 45730 2956 45790 3988
rect 45850 2896 45910 3926
rect 45970 2956 46030 3988
rect 46090 2896 46150 3926
rect 46210 3834 46276 3988
rect 46210 3770 46211 3834
rect 46275 3770 46276 3834
rect 46210 3754 46276 3770
rect 46210 3690 46211 3754
rect 46275 3690 46276 3754
rect 46210 3674 46276 3690
rect 46210 3610 46211 3674
rect 46275 3610 46276 3674
rect 46210 3594 46276 3610
rect 46210 3530 46211 3594
rect 46275 3530 46276 3594
rect 46210 3514 46276 3530
rect 46210 3450 46211 3514
rect 46275 3450 46276 3514
rect 46210 3434 46276 3450
rect 46210 3370 46211 3434
rect 46275 3370 46276 3434
rect 46210 3354 46276 3370
rect 46210 3290 46211 3354
rect 46275 3290 46276 3354
rect 46210 3274 46276 3290
rect 46210 3210 46211 3274
rect 46275 3210 46276 3274
rect 46210 3194 46276 3210
rect 46210 3130 46211 3194
rect 46275 3130 46276 3194
rect 46210 3114 46276 3130
rect 46210 3050 46211 3114
rect 46275 3050 46276 3114
rect 46210 2960 46276 3050
rect 46336 2956 46396 3988
rect 46456 2896 46516 3926
rect 46576 2956 46636 3988
rect 46696 2896 46756 3926
rect 46816 3834 46882 3988
rect 46816 3770 46817 3834
rect 46881 3770 46882 3834
rect 46816 3754 46882 3770
rect 46816 3690 46817 3754
rect 46881 3690 46882 3754
rect 46816 3674 46882 3690
rect 46816 3610 46817 3674
rect 46881 3610 46882 3674
rect 46816 3594 46882 3610
rect 46816 3530 46817 3594
rect 46881 3530 46882 3594
rect 46816 3514 46882 3530
rect 46816 3450 46817 3514
rect 46881 3450 46882 3514
rect 46816 3434 46882 3450
rect 46816 3370 46817 3434
rect 46881 3370 46882 3434
rect 46816 3354 46882 3370
rect 46816 3290 46817 3354
rect 46881 3290 46882 3354
rect 46816 3274 46882 3290
rect 46816 3210 46817 3274
rect 46881 3210 46882 3274
rect 46816 3194 46882 3210
rect 46816 3130 46817 3194
rect 46881 3130 46882 3194
rect 46816 3114 46882 3130
rect 46816 3050 46817 3114
rect 46881 3050 46882 3114
rect 46816 2960 46882 3050
rect 46942 2956 47002 3988
rect 47062 2896 47122 3926
rect 47182 2956 47242 3988
rect 47302 2896 47362 3926
rect 47422 3834 47488 3988
rect 47422 3770 47423 3834
rect 47487 3770 47488 3834
rect 47422 3754 47488 3770
rect 47422 3690 47423 3754
rect 47487 3690 47488 3754
rect 47422 3674 47488 3690
rect 47422 3610 47423 3674
rect 47487 3610 47488 3674
rect 47422 3594 47488 3610
rect 47422 3530 47423 3594
rect 47487 3530 47488 3594
rect 47422 3514 47488 3530
rect 47422 3450 47423 3514
rect 47487 3450 47488 3514
rect 47422 3434 47488 3450
rect 47422 3370 47423 3434
rect 47487 3370 47488 3434
rect 47422 3354 47488 3370
rect 47422 3290 47423 3354
rect 47487 3290 47488 3354
rect 47422 3274 47488 3290
rect 47422 3210 47423 3274
rect 47487 3210 47488 3274
rect 47422 3194 47488 3210
rect 47422 3130 47423 3194
rect 47487 3130 47488 3194
rect 47422 3114 47488 3130
rect 47422 3050 47423 3114
rect 47487 3050 47488 3114
rect 47422 2960 47488 3050
rect 47548 2956 47608 3988
rect 47668 2896 47728 3926
rect 47788 2956 47848 3988
rect 47908 2896 47968 3926
rect 48028 3834 48094 3988
rect 48028 3770 48029 3834
rect 48093 3770 48094 3834
rect 48028 3754 48094 3770
rect 48028 3690 48029 3754
rect 48093 3690 48094 3754
rect 48028 3674 48094 3690
rect 48028 3610 48029 3674
rect 48093 3610 48094 3674
rect 48028 3594 48094 3610
rect 48028 3530 48029 3594
rect 48093 3530 48094 3594
rect 48028 3514 48094 3530
rect 48028 3450 48029 3514
rect 48093 3450 48094 3514
rect 48028 3434 48094 3450
rect 48028 3370 48029 3434
rect 48093 3370 48094 3434
rect 48028 3354 48094 3370
rect 48028 3290 48029 3354
rect 48093 3290 48094 3354
rect 48028 3274 48094 3290
rect 48028 3210 48029 3274
rect 48093 3210 48094 3274
rect 48028 3194 48094 3210
rect 48028 3130 48029 3194
rect 48093 3130 48094 3194
rect 48028 3114 48094 3130
rect 48028 3050 48029 3114
rect 48093 3050 48094 3114
rect 48028 2960 48094 3050
rect 48154 2956 48214 3988
rect 48274 2896 48334 3926
rect 48394 2956 48454 3988
rect 48514 2896 48574 3926
rect 48634 3834 48700 3988
rect 48634 3770 48635 3834
rect 48699 3770 48700 3834
rect 48634 3754 48700 3770
rect 48634 3690 48635 3754
rect 48699 3690 48700 3754
rect 48634 3674 48700 3690
rect 48634 3610 48635 3674
rect 48699 3610 48700 3674
rect 48634 3594 48700 3610
rect 48634 3530 48635 3594
rect 48699 3530 48700 3594
rect 48634 3514 48700 3530
rect 48634 3450 48635 3514
rect 48699 3450 48700 3514
rect 48634 3434 48700 3450
rect 48634 3370 48635 3434
rect 48699 3370 48700 3434
rect 48634 3354 48700 3370
rect 48634 3290 48635 3354
rect 48699 3290 48700 3354
rect 48634 3274 48700 3290
rect 48634 3210 48635 3274
rect 48699 3210 48700 3274
rect 48634 3194 48700 3210
rect 48634 3130 48635 3194
rect 48699 3130 48700 3194
rect 48634 3114 48700 3130
rect 48634 3050 48635 3114
rect 48699 3050 48700 3114
rect 48634 2960 48700 3050
rect 48760 2956 48820 3988
rect 48880 2896 48940 3926
rect 49000 2956 49060 3988
rect 49120 2896 49180 3926
rect 49240 3834 49306 3988
rect 49240 3770 49241 3834
rect 49305 3770 49306 3834
rect 49240 3754 49306 3770
rect 49240 3690 49241 3754
rect 49305 3690 49306 3754
rect 49240 3674 49306 3690
rect 49240 3610 49241 3674
rect 49305 3610 49306 3674
rect 49240 3594 49306 3610
rect 49240 3530 49241 3594
rect 49305 3530 49306 3594
rect 49240 3514 49306 3530
rect 49240 3450 49241 3514
rect 49305 3450 49306 3514
rect 49240 3434 49306 3450
rect 49240 3370 49241 3434
rect 49305 3370 49306 3434
rect 49240 3354 49306 3370
rect 49240 3290 49241 3354
rect 49305 3290 49306 3354
rect 49240 3274 49306 3290
rect 49240 3210 49241 3274
rect 49305 3210 49306 3274
rect 49240 3194 49306 3210
rect 49240 3130 49241 3194
rect 49305 3130 49306 3194
rect 49240 3114 49306 3130
rect 49240 3050 49241 3114
rect 49305 3050 49306 3114
rect 49240 2960 49306 3050
rect 49366 2956 49426 3988
rect 49486 2896 49546 3926
rect 49606 2956 49666 3988
rect 49726 2896 49786 3926
rect 49846 3834 49912 3988
rect 49846 3770 49847 3834
rect 49911 3770 49912 3834
rect 49846 3754 49912 3770
rect 49846 3690 49847 3754
rect 49911 3690 49912 3754
rect 49846 3674 49912 3690
rect 49846 3610 49847 3674
rect 49911 3610 49912 3674
rect 49846 3594 49912 3610
rect 49846 3530 49847 3594
rect 49911 3530 49912 3594
rect 49846 3514 49912 3530
rect 49846 3450 49847 3514
rect 49911 3450 49912 3514
rect 49846 3434 49912 3450
rect 49846 3370 49847 3434
rect 49911 3370 49912 3434
rect 49846 3354 49912 3370
rect 49846 3290 49847 3354
rect 49911 3290 49912 3354
rect 49846 3274 49912 3290
rect 49846 3210 49847 3274
rect 49911 3210 49912 3274
rect 49846 3194 49912 3210
rect 49846 3130 49847 3194
rect 49911 3130 49912 3194
rect 49846 3114 49912 3130
rect 49846 3050 49847 3114
rect 49911 3050 49912 3114
rect 49846 2960 49912 3050
rect 49972 2956 50032 3988
rect 50092 2896 50152 3926
rect 50212 2956 50272 3988
rect 50332 2896 50392 3926
rect 50452 3834 50518 3988
rect 50452 3770 50453 3834
rect 50517 3770 50518 3834
rect 50452 3754 50518 3770
rect 50452 3690 50453 3754
rect 50517 3690 50518 3754
rect 50452 3674 50518 3690
rect 50452 3610 50453 3674
rect 50517 3610 50518 3674
rect 50452 3594 50518 3610
rect 50452 3530 50453 3594
rect 50517 3530 50518 3594
rect 50452 3514 50518 3530
rect 50452 3450 50453 3514
rect 50517 3450 50518 3514
rect 50452 3434 50518 3450
rect 50452 3370 50453 3434
rect 50517 3370 50518 3434
rect 50452 3354 50518 3370
rect 50452 3290 50453 3354
rect 50517 3290 50518 3354
rect 50452 3274 50518 3290
rect 50452 3210 50453 3274
rect 50517 3210 50518 3274
rect 50452 3194 50518 3210
rect 50452 3130 50453 3194
rect 50517 3130 50518 3194
rect 50452 3114 50518 3130
rect 50452 3050 50453 3114
rect 50517 3050 50518 3114
rect 50452 2960 50518 3050
rect 50578 2956 50638 3988
rect 50698 2896 50758 3926
rect 50818 2956 50878 3988
rect 50938 2896 50998 3926
rect 51058 3834 51124 3988
rect 51058 3770 51059 3834
rect 51123 3770 51124 3834
rect 51058 3754 51124 3770
rect 51058 3690 51059 3754
rect 51123 3690 51124 3754
rect 51058 3674 51124 3690
rect 51058 3610 51059 3674
rect 51123 3610 51124 3674
rect 51058 3594 51124 3610
rect 51058 3530 51059 3594
rect 51123 3530 51124 3594
rect 51058 3514 51124 3530
rect 51058 3450 51059 3514
rect 51123 3450 51124 3514
rect 51058 3434 51124 3450
rect 51058 3370 51059 3434
rect 51123 3370 51124 3434
rect 51058 3354 51124 3370
rect 51058 3290 51059 3354
rect 51123 3290 51124 3354
rect 51058 3274 51124 3290
rect 51058 3210 51059 3274
rect 51123 3210 51124 3274
rect 51058 3194 51124 3210
rect 51058 3130 51059 3194
rect 51123 3130 51124 3194
rect 51058 3114 51124 3130
rect 51058 3050 51059 3114
rect 51123 3050 51124 3114
rect 51058 2960 51124 3050
rect 51184 2956 51244 3988
rect 51304 2896 51364 3926
rect 51424 2956 51484 3988
rect 51544 2896 51604 3926
rect 51664 3834 51730 3988
rect 51664 3770 51665 3834
rect 51729 3770 51730 3834
rect 51664 3754 51730 3770
rect 51664 3690 51665 3754
rect 51729 3690 51730 3754
rect 51664 3674 51730 3690
rect 51664 3610 51665 3674
rect 51729 3610 51730 3674
rect 51664 3594 51730 3610
rect 51664 3530 51665 3594
rect 51729 3530 51730 3594
rect 51664 3514 51730 3530
rect 51664 3450 51665 3514
rect 51729 3450 51730 3514
rect 51664 3434 51730 3450
rect 51664 3370 51665 3434
rect 51729 3370 51730 3434
rect 51664 3354 51730 3370
rect 51664 3290 51665 3354
rect 51729 3290 51730 3354
rect 51664 3274 51730 3290
rect 51664 3210 51665 3274
rect 51729 3210 51730 3274
rect 51664 3194 51730 3210
rect 51664 3130 51665 3194
rect 51729 3130 51730 3194
rect 51664 3114 51730 3130
rect 51664 3050 51665 3114
rect 51729 3050 51730 3114
rect 51664 2960 51730 3050
rect 32272 2894 51730 2896
rect 32272 2830 32376 2894
rect 32440 2830 32456 2894
rect 32520 2830 32536 2894
rect 32600 2830 32616 2894
rect 32680 2830 32696 2894
rect 32760 2830 32776 2894
rect 32840 2830 32982 2894
rect 33046 2830 33062 2894
rect 33126 2830 33142 2894
rect 33206 2830 33222 2894
rect 33286 2830 33302 2894
rect 33366 2830 33382 2894
rect 33446 2830 33588 2894
rect 33652 2830 33668 2894
rect 33732 2830 33748 2894
rect 33812 2830 33828 2894
rect 33892 2830 33908 2894
rect 33972 2830 33988 2894
rect 34052 2830 34194 2894
rect 34258 2830 34274 2894
rect 34338 2830 34354 2894
rect 34418 2830 34434 2894
rect 34498 2830 34514 2894
rect 34578 2830 34594 2894
rect 34658 2830 34800 2894
rect 34864 2830 34880 2894
rect 34944 2830 34960 2894
rect 35024 2830 35040 2894
rect 35104 2830 35120 2894
rect 35184 2830 35200 2894
rect 35264 2830 35406 2894
rect 35470 2830 35486 2894
rect 35550 2830 35566 2894
rect 35630 2830 35646 2894
rect 35710 2830 35726 2894
rect 35790 2830 35806 2894
rect 35870 2830 36012 2894
rect 36076 2830 36092 2894
rect 36156 2830 36172 2894
rect 36236 2830 36252 2894
rect 36316 2830 36332 2894
rect 36396 2830 36412 2894
rect 36476 2830 36618 2894
rect 36682 2830 36698 2894
rect 36762 2830 36778 2894
rect 36842 2830 36858 2894
rect 36922 2830 36938 2894
rect 37002 2830 37018 2894
rect 37082 2830 37224 2894
rect 37288 2830 37304 2894
rect 37368 2830 37384 2894
rect 37448 2830 37464 2894
rect 37528 2830 37544 2894
rect 37608 2830 37624 2894
rect 37688 2830 37830 2894
rect 37894 2830 37910 2894
rect 37974 2830 37990 2894
rect 38054 2830 38070 2894
rect 38134 2830 38150 2894
rect 38214 2830 38230 2894
rect 38294 2830 38436 2894
rect 38500 2830 38516 2894
rect 38580 2830 38596 2894
rect 38660 2830 38676 2894
rect 38740 2830 38756 2894
rect 38820 2830 38836 2894
rect 38900 2830 39042 2894
rect 39106 2830 39122 2894
rect 39186 2830 39202 2894
rect 39266 2830 39282 2894
rect 39346 2830 39362 2894
rect 39426 2830 39442 2894
rect 39506 2830 39648 2894
rect 39712 2830 39728 2894
rect 39792 2830 39808 2894
rect 39872 2830 39888 2894
rect 39952 2830 39968 2894
rect 40032 2830 40048 2894
rect 40112 2830 40254 2894
rect 40318 2830 40334 2894
rect 40398 2830 40414 2894
rect 40478 2830 40494 2894
rect 40558 2830 40574 2894
rect 40638 2830 40654 2894
rect 40718 2830 40860 2894
rect 40924 2830 40940 2894
rect 41004 2830 41020 2894
rect 41084 2830 41100 2894
rect 41164 2830 41180 2894
rect 41244 2830 41260 2894
rect 41324 2830 41466 2894
rect 41530 2830 41546 2894
rect 41610 2830 41626 2894
rect 41690 2830 41706 2894
rect 41770 2830 41786 2894
rect 41850 2830 41866 2894
rect 41930 2830 42072 2894
rect 42136 2830 42152 2894
rect 42216 2830 42232 2894
rect 42296 2830 42312 2894
rect 42376 2830 42392 2894
rect 42456 2830 42472 2894
rect 42536 2830 42678 2894
rect 42742 2830 42758 2894
rect 42822 2830 42838 2894
rect 42902 2830 42918 2894
rect 42982 2830 42998 2894
rect 43062 2830 43078 2894
rect 43142 2830 43284 2894
rect 43348 2830 43364 2894
rect 43428 2830 43444 2894
rect 43508 2830 43524 2894
rect 43588 2830 43604 2894
rect 43668 2830 43684 2894
rect 43748 2830 43890 2894
rect 43954 2830 43970 2894
rect 44034 2830 44050 2894
rect 44114 2830 44130 2894
rect 44194 2830 44210 2894
rect 44274 2830 44290 2894
rect 44354 2830 44496 2894
rect 44560 2830 44576 2894
rect 44640 2830 44656 2894
rect 44720 2830 44736 2894
rect 44800 2830 44816 2894
rect 44880 2830 44896 2894
rect 44960 2830 45102 2894
rect 45166 2830 45182 2894
rect 45246 2830 45262 2894
rect 45326 2830 45342 2894
rect 45406 2830 45422 2894
rect 45486 2830 45502 2894
rect 45566 2830 45708 2894
rect 45772 2830 45788 2894
rect 45852 2830 45868 2894
rect 45932 2830 45948 2894
rect 46012 2830 46028 2894
rect 46092 2830 46108 2894
rect 46172 2830 46314 2894
rect 46378 2830 46394 2894
rect 46458 2830 46474 2894
rect 46538 2830 46554 2894
rect 46618 2830 46634 2894
rect 46698 2830 46714 2894
rect 46778 2830 46920 2894
rect 46984 2830 47000 2894
rect 47064 2830 47080 2894
rect 47144 2830 47160 2894
rect 47224 2830 47240 2894
rect 47304 2830 47320 2894
rect 47384 2830 47526 2894
rect 47590 2830 47606 2894
rect 47670 2830 47686 2894
rect 47750 2830 47766 2894
rect 47830 2830 47846 2894
rect 47910 2830 47926 2894
rect 47990 2830 48132 2894
rect 48196 2830 48212 2894
rect 48276 2830 48292 2894
rect 48356 2830 48372 2894
rect 48436 2830 48452 2894
rect 48516 2830 48532 2894
rect 48596 2830 48738 2894
rect 48802 2830 48818 2894
rect 48882 2830 48898 2894
rect 48962 2830 48978 2894
rect 49042 2830 49058 2894
rect 49122 2830 49138 2894
rect 49202 2830 49344 2894
rect 49408 2830 49424 2894
rect 49488 2830 49504 2894
rect 49568 2830 49584 2894
rect 49648 2830 49664 2894
rect 49728 2830 49744 2894
rect 49808 2830 49950 2894
rect 50014 2830 50030 2894
rect 50094 2830 50110 2894
rect 50174 2830 50190 2894
rect 50254 2830 50270 2894
rect 50334 2830 50350 2894
rect 50414 2830 50556 2894
rect 50620 2830 50636 2894
rect 50700 2830 50716 2894
rect 50780 2830 50796 2894
rect 50860 2830 50876 2894
rect 50940 2830 50956 2894
rect 51020 2830 51162 2894
rect 51226 2830 51242 2894
rect 51306 2830 51322 2894
rect 51386 2830 51402 2894
rect 51466 2830 51482 2894
rect 51546 2830 51562 2894
rect 51626 2830 51730 2894
rect 32272 2828 51730 2830
<< via3 >>
rect 32376 5150 32440 5214
rect 32456 5150 32520 5214
rect 32536 5150 32600 5214
rect 32616 5150 32680 5214
rect 32696 5150 32760 5214
rect 32776 5150 32840 5214
rect 32982 5150 33046 5214
rect 33062 5150 33126 5214
rect 33142 5150 33206 5214
rect 33222 5150 33286 5214
rect 33302 5150 33366 5214
rect 33382 5150 33446 5214
rect 33588 5150 33652 5214
rect 33668 5150 33732 5214
rect 33748 5150 33812 5214
rect 33828 5150 33892 5214
rect 33908 5150 33972 5214
rect 33988 5150 34052 5214
rect 34194 5150 34258 5214
rect 34274 5150 34338 5214
rect 34354 5150 34418 5214
rect 34434 5150 34498 5214
rect 34514 5150 34578 5214
rect 34594 5150 34658 5214
rect 34800 5150 34864 5214
rect 34880 5150 34944 5214
rect 34960 5150 35024 5214
rect 35040 5150 35104 5214
rect 35120 5150 35184 5214
rect 35200 5150 35264 5214
rect 35406 5150 35470 5214
rect 35486 5150 35550 5214
rect 35566 5150 35630 5214
rect 35646 5150 35710 5214
rect 35726 5150 35790 5214
rect 35806 5150 35870 5214
rect 36012 5150 36076 5214
rect 36092 5150 36156 5214
rect 36172 5150 36236 5214
rect 36252 5150 36316 5214
rect 36332 5150 36396 5214
rect 36412 5150 36476 5214
rect 36618 5150 36682 5214
rect 36698 5150 36762 5214
rect 36778 5150 36842 5214
rect 36858 5150 36922 5214
rect 36938 5150 37002 5214
rect 37018 5150 37082 5214
rect 37224 5150 37288 5214
rect 37304 5150 37368 5214
rect 37384 5150 37448 5214
rect 37464 5150 37528 5214
rect 37544 5150 37608 5214
rect 37624 5150 37688 5214
rect 37830 5150 37894 5214
rect 37910 5150 37974 5214
rect 37990 5150 38054 5214
rect 38070 5150 38134 5214
rect 38150 5150 38214 5214
rect 38230 5150 38294 5214
rect 38436 5150 38500 5214
rect 38516 5150 38580 5214
rect 38596 5150 38660 5214
rect 38676 5150 38740 5214
rect 38756 5150 38820 5214
rect 38836 5150 38900 5214
rect 39042 5150 39106 5214
rect 39122 5150 39186 5214
rect 39202 5150 39266 5214
rect 39282 5150 39346 5214
rect 39362 5150 39426 5214
rect 39442 5150 39506 5214
rect 39648 5150 39712 5214
rect 39728 5150 39792 5214
rect 39808 5150 39872 5214
rect 39888 5150 39952 5214
rect 39968 5150 40032 5214
rect 40048 5150 40112 5214
rect 40254 5150 40318 5214
rect 40334 5150 40398 5214
rect 40414 5150 40478 5214
rect 40494 5150 40558 5214
rect 40574 5150 40638 5214
rect 40654 5150 40718 5214
rect 40860 5150 40924 5214
rect 40940 5150 41004 5214
rect 41020 5150 41084 5214
rect 41100 5150 41164 5214
rect 41180 5150 41244 5214
rect 41260 5150 41324 5214
rect 41466 5150 41530 5214
rect 41546 5150 41610 5214
rect 41626 5150 41690 5214
rect 41706 5150 41770 5214
rect 41786 5150 41850 5214
rect 41866 5150 41930 5214
rect 42072 5150 42136 5214
rect 42152 5150 42216 5214
rect 42232 5150 42296 5214
rect 42312 5150 42376 5214
rect 42392 5150 42456 5214
rect 42472 5150 42536 5214
rect 42678 5150 42742 5214
rect 42758 5150 42822 5214
rect 42838 5150 42902 5214
rect 42918 5150 42982 5214
rect 42998 5150 43062 5214
rect 43078 5150 43142 5214
rect 43284 5150 43348 5214
rect 43364 5150 43428 5214
rect 43444 5150 43508 5214
rect 43524 5150 43588 5214
rect 43604 5150 43668 5214
rect 43684 5150 43748 5214
rect 43890 5150 43954 5214
rect 43970 5150 44034 5214
rect 44050 5150 44114 5214
rect 44130 5150 44194 5214
rect 44210 5150 44274 5214
rect 44290 5150 44354 5214
rect 44496 5150 44560 5214
rect 44576 5150 44640 5214
rect 44656 5150 44720 5214
rect 44736 5150 44800 5214
rect 44816 5150 44880 5214
rect 44896 5150 44960 5214
rect 45102 5150 45166 5214
rect 45182 5150 45246 5214
rect 45262 5150 45326 5214
rect 45342 5150 45406 5214
rect 45422 5150 45486 5214
rect 45502 5150 45566 5214
rect 45708 5150 45772 5214
rect 45788 5150 45852 5214
rect 45868 5150 45932 5214
rect 45948 5150 46012 5214
rect 46028 5150 46092 5214
rect 46108 5150 46172 5214
rect 46314 5150 46378 5214
rect 46394 5150 46458 5214
rect 46474 5150 46538 5214
rect 46554 5150 46618 5214
rect 46634 5150 46698 5214
rect 46714 5150 46778 5214
rect 46920 5150 46984 5214
rect 47000 5150 47064 5214
rect 47080 5150 47144 5214
rect 47160 5150 47224 5214
rect 47240 5150 47304 5214
rect 47320 5150 47384 5214
rect 47526 5150 47590 5214
rect 47606 5150 47670 5214
rect 47686 5150 47750 5214
rect 47766 5150 47830 5214
rect 47846 5150 47910 5214
rect 47926 5150 47990 5214
rect 48132 5150 48196 5214
rect 48212 5150 48276 5214
rect 48292 5150 48356 5214
rect 48372 5150 48436 5214
rect 48452 5150 48516 5214
rect 48532 5150 48596 5214
rect 48738 5150 48802 5214
rect 48818 5150 48882 5214
rect 48898 5150 48962 5214
rect 48978 5150 49042 5214
rect 49058 5150 49122 5214
rect 49138 5150 49202 5214
rect 49344 5150 49408 5214
rect 49424 5150 49488 5214
rect 49504 5150 49568 5214
rect 49584 5150 49648 5214
rect 49664 5150 49728 5214
rect 49744 5150 49808 5214
rect 49950 5150 50014 5214
rect 50030 5150 50094 5214
rect 50110 5150 50174 5214
rect 50190 5150 50254 5214
rect 50270 5150 50334 5214
rect 50350 5150 50414 5214
rect 50556 5150 50620 5214
rect 50636 5150 50700 5214
rect 50716 5150 50780 5214
rect 50796 5150 50860 5214
rect 50876 5150 50940 5214
rect 50956 5150 51020 5214
rect 51162 5150 51226 5214
rect 51242 5150 51306 5214
rect 51322 5150 51386 5214
rect 51402 5150 51466 5214
rect 51482 5150 51546 5214
rect 51562 5150 51626 5214
rect 32273 4930 32337 4994
rect 32273 4850 32337 4914
rect 32273 4770 32337 4834
rect 32273 4690 32337 4754
rect 32273 4610 32337 4674
rect 32273 4530 32337 4594
rect 32273 4450 32337 4514
rect 32273 4370 32337 4434
rect 32273 4290 32337 4354
rect 32273 4210 32337 4274
rect 32879 4930 32943 4994
rect 32879 4850 32943 4914
rect 32879 4770 32943 4834
rect 32879 4690 32943 4754
rect 32879 4610 32943 4674
rect 32879 4530 32943 4594
rect 32879 4450 32943 4514
rect 32879 4370 32943 4434
rect 32879 4290 32943 4354
rect 32879 4210 32943 4274
rect 33485 4930 33549 4994
rect 33485 4850 33549 4914
rect 33485 4770 33549 4834
rect 33485 4690 33549 4754
rect 33485 4610 33549 4674
rect 33485 4530 33549 4594
rect 33485 4450 33549 4514
rect 33485 4370 33549 4434
rect 33485 4290 33549 4354
rect 33485 4210 33549 4274
rect 34091 4930 34155 4994
rect 34091 4850 34155 4914
rect 34091 4770 34155 4834
rect 34091 4690 34155 4754
rect 34091 4610 34155 4674
rect 34091 4530 34155 4594
rect 34091 4450 34155 4514
rect 34091 4370 34155 4434
rect 34091 4290 34155 4354
rect 34091 4210 34155 4274
rect 34697 4930 34761 4994
rect 34697 4850 34761 4914
rect 34697 4770 34761 4834
rect 34697 4690 34761 4754
rect 34697 4610 34761 4674
rect 34697 4530 34761 4594
rect 34697 4450 34761 4514
rect 34697 4370 34761 4434
rect 34697 4290 34761 4354
rect 34697 4210 34761 4274
rect 35303 4930 35367 4994
rect 35303 4850 35367 4914
rect 35303 4770 35367 4834
rect 35303 4690 35367 4754
rect 35303 4610 35367 4674
rect 35303 4530 35367 4594
rect 35303 4450 35367 4514
rect 35303 4370 35367 4434
rect 35303 4290 35367 4354
rect 35303 4210 35367 4274
rect 35909 4930 35973 4994
rect 35909 4850 35973 4914
rect 35909 4770 35973 4834
rect 35909 4690 35973 4754
rect 35909 4610 35973 4674
rect 35909 4530 35973 4594
rect 35909 4450 35973 4514
rect 35909 4370 35973 4434
rect 35909 4290 35973 4354
rect 35909 4210 35973 4274
rect 36515 4930 36579 4994
rect 36515 4850 36579 4914
rect 36515 4770 36579 4834
rect 36515 4690 36579 4754
rect 36515 4610 36579 4674
rect 36515 4530 36579 4594
rect 36515 4450 36579 4514
rect 36515 4370 36579 4434
rect 36515 4290 36579 4354
rect 36515 4210 36579 4274
rect 37121 4930 37185 4994
rect 37121 4850 37185 4914
rect 37121 4770 37185 4834
rect 37121 4690 37185 4754
rect 37121 4610 37185 4674
rect 37121 4530 37185 4594
rect 37121 4450 37185 4514
rect 37121 4370 37185 4434
rect 37121 4290 37185 4354
rect 37121 4210 37185 4274
rect 37727 4930 37791 4994
rect 37727 4850 37791 4914
rect 37727 4770 37791 4834
rect 37727 4690 37791 4754
rect 37727 4610 37791 4674
rect 37727 4530 37791 4594
rect 37727 4450 37791 4514
rect 37727 4370 37791 4434
rect 37727 4290 37791 4354
rect 37727 4210 37791 4274
rect 38333 4930 38397 4994
rect 38333 4850 38397 4914
rect 38333 4770 38397 4834
rect 38333 4690 38397 4754
rect 38333 4610 38397 4674
rect 38333 4530 38397 4594
rect 38333 4450 38397 4514
rect 38333 4370 38397 4434
rect 38333 4290 38397 4354
rect 38333 4210 38397 4274
rect 38939 4930 39003 4994
rect 38939 4850 39003 4914
rect 38939 4770 39003 4834
rect 38939 4690 39003 4754
rect 38939 4610 39003 4674
rect 38939 4530 39003 4594
rect 38939 4450 39003 4514
rect 38939 4370 39003 4434
rect 38939 4290 39003 4354
rect 38939 4210 39003 4274
rect 39545 4930 39609 4994
rect 39545 4850 39609 4914
rect 39545 4770 39609 4834
rect 39545 4690 39609 4754
rect 39545 4610 39609 4674
rect 39545 4530 39609 4594
rect 39545 4450 39609 4514
rect 39545 4370 39609 4434
rect 39545 4290 39609 4354
rect 39545 4210 39609 4274
rect 40151 4930 40215 4994
rect 40151 4850 40215 4914
rect 40151 4770 40215 4834
rect 40151 4690 40215 4754
rect 40151 4610 40215 4674
rect 40151 4530 40215 4594
rect 40151 4450 40215 4514
rect 40151 4370 40215 4434
rect 40151 4290 40215 4354
rect 40151 4210 40215 4274
rect 40757 4930 40821 4994
rect 40757 4850 40821 4914
rect 40757 4770 40821 4834
rect 40757 4690 40821 4754
rect 40757 4610 40821 4674
rect 40757 4530 40821 4594
rect 40757 4450 40821 4514
rect 40757 4370 40821 4434
rect 40757 4290 40821 4354
rect 40757 4210 40821 4274
rect 41363 4930 41427 4994
rect 41363 4850 41427 4914
rect 41363 4770 41427 4834
rect 41363 4690 41427 4754
rect 41363 4610 41427 4674
rect 41363 4530 41427 4594
rect 41363 4450 41427 4514
rect 41363 4370 41427 4434
rect 41363 4290 41427 4354
rect 41363 4210 41427 4274
rect 41969 4930 42033 4994
rect 41969 4850 42033 4914
rect 41969 4770 42033 4834
rect 41969 4690 42033 4754
rect 41969 4610 42033 4674
rect 41969 4530 42033 4594
rect 41969 4450 42033 4514
rect 41969 4370 42033 4434
rect 41969 4290 42033 4354
rect 41969 4210 42033 4274
rect 42575 4930 42639 4994
rect 42575 4850 42639 4914
rect 42575 4770 42639 4834
rect 42575 4690 42639 4754
rect 42575 4610 42639 4674
rect 42575 4530 42639 4594
rect 42575 4450 42639 4514
rect 42575 4370 42639 4434
rect 42575 4290 42639 4354
rect 42575 4210 42639 4274
rect 43181 4930 43245 4994
rect 43181 4850 43245 4914
rect 43181 4770 43245 4834
rect 43181 4690 43245 4754
rect 43181 4610 43245 4674
rect 43181 4530 43245 4594
rect 43181 4450 43245 4514
rect 43181 4370 43245 4434
rect 43181 4290 43245 4354
rect 43181 4210 43245 4274
rect 43787 4930 43851 4994
rect 43787 4850 43851 4914
rect 43787 4770 43851 4834
rect 43787 4690 43851 4754
rect 43787 4610 43851 4674
rect 43787 4530 43851 4594
rect 43787 4450 43851 4514
rect 43787 4370 43851 4434
rect 43787 4290 43851 4354
rect 43787 4210 43851 4274
rect 44393 4930 44457 4994
rect 44393 4850 44457 4914
rect 44393 4770 44457 4834
rect 44393 4690 44457 4754
rect 44393 4610 44457 4674
rect 44393 4530 44457 4594
rect 44393 4450 44457 4514
rect 44393 4370 44457 4434
rect 44393 4290 44457 4354
rect 44393 4210 44457 4274
rect 44999 4930 45063 4994
rect 44999 4850 45063 4914
rect 44999 4770 45063 4834
rect 44999 4690 45063 4754
rect 44999 4610 45063 4674
rect 44999 4530 45063 4594
rect 44999 4450 45063 4514
rect 44999 4370 45063 4434
rect 44999 4290 45063 4354
rect 44999 4210 45063 4274
rect 45605 4930 45669 4994
rect 45605 4850 45669 4914
rect 45605 4770 45669 4834
rect 45605 4690 45669 4754
rect 45605 4610 45669 4674
rect 45605 4530 45669 4594
rect 45605 4450 45669 4514
rect 45605 4370 45669 4434
rect 45605 4290 45669 4354
rect 45605 4210 45669 4274
rect 46211 4930 46275 4994
rect 46211 4850 46275 4914
rect 46211 4770 46275 4834
rect 46211 4690 46275 4754
rect 46211 4610 46275 4674
rect 46211 4530 46275 4594
rect 46211 4450 46275 4514
rect 46211 4370 46275 4434
rect 46211 4290 46275 4354
rect 46211 4210 46275 4274
rect 46817 4930 46881 4994
rect 46817 4850 46881 4914
rect 46817 4770 46881 4834
rect 46817 4690 46881 4754
rect 46817 4610 46881 4674
rect 46817 4530 46881 4594
rect 46817 4450 46881 4514
rect 46817 4370 46881 4434
rect 46817 4290 46881 4354
rect 46817 4210 46881 4274
rect 47423 4930 47487 4994
rect 47423 4850 47487 4914
rect 47423 4770 47487 4834
rect 47423 4690 47487 4754
rect 47423 4610 47487 4674
rect 47423 4530 47487 4594
rect 47423 4450 47487 4514
rect 47423 4370 47487 4434
rect 47423 4290 47487 4354
rect 47423 4210 47487 4274
rect 48029 4930 48093 4994
rect 48029 4850 48093 4914
rect 48029 4770 48093 4834
rect 48029 4690 48093 4754
rect 48029 4610 48093 4674
rect 48029 4530 48093 4594
rect 48029 4450 48093 4514
rect 48029 4370 48093 4434
rect 48029 4290 48093 4354
rect 48029 4210 48093 4274
rect 48635 4930 48699 4994
rect 48635 4850 48699 4914
rect 48635 4770 48699 4834
rect 48635 4690 48699 4754
rect 48635 4610 48699 4674
rect 48635 4530 48699 4594
rect 48635 4450 48699 4514
rect 48635 4370 48699 4434
rect 48635 4290 48699 4354
rect 48635 4210 48699 4274
rect 49241 4930 49305 4994
rect 49241 4850 49305 4914
rect 49241 4770 49305 4834
rect 49241 4690 49305 4754
rect 49241 4610 49305 4674
rect 49241 4530 49305 4594
rect 49241 4450 49305 4514
rect 49241 4370 49305 4434
rect 49241 4290 49305 4354
rect 49241 4210 49305 4274
rect 49847 4930 49911 4994
rect 49847 4850 49911 4914
rect 49847 4770 49911 4834
rect 49847 4690 49911 4754
rect 49847 4610 49911 4674
rect 49847 4530 49911 4594
rect 49847 4450 49911 4514
rect 49847 4370 49911 4434
rect 49847 4290 49911 4354
rect 49847 4210 49911 4274
rect 50453 4930 50517 4994
rect 50453 4850 50517 4914
rect 50453 4770 50517 4834
rect 50453 4690 50517 4754
rect 50453 4610 50517 4674
rect 50453 4530 50517 4594
rect 50453 4450 50517 4514
rect 50453 4370 50517 4434
rect 50453 4290 50517 4354
rect 50453 4210 50517 4274
rect 51059 4930 51123 4994
rect 51059 4850 51123 4914
rect 51059 4770 51123 4834
rect 51059 4690 51123 4754
rect 51059 4610 51123 4674
rect 51059 4530 51123 4594
rect 51059 4450 51123 4514
rect 51059 4370 51123 4434
rect 51059 4290 51123 4354
rect 51059 4210 51123 4274
rect 51665 4930 51729 4994
rect 51665 4850 51729 4914
rect 51665 4770 51729 4834
rect 51665 4690 51729 4754
rect 51665 4610 51729 4674
rect 51665 4530 51729 4594
rect 51665 4450 51729 4514
rect 51665 4370 51729 4434
rect 51665 4290 51729 4354
rect 51665 4210 51729 4274
rect 32376 3990 32440 4054
rect 32456 3990 32520 4054
rect 32536 3990 32600 4054
rect 32616 3990 32680 4054
rect 32696 3990 32760 4054
rect 32776 3990 32840 4054
rect 32982 3990 33046 4054
rect 33062 3990 33126 4054
rect 33142 3990 33206 4054
rect 33222 3990 33286 4054
rect 33302 3990 33366 4054
rect 33382 3990 33446 4054
rect 33588 3990 33652 4054
rect 33668 3990 33732 4054
rect 33748 3990 33812 4054
rect 33828 3990 33892 4054
rect 33908 3990 33972 4054
rect 33988 3990 34052 4054
rect 34194 3990 34258 4054
rect 34274 3990 34338 4054
rect 34354 3990 34418 4054
rect 34434 3990 34498 4054
rect 34514 3990 34578 4054
rect 34594 3990 34658 4054
rect 34800 3990 34864 4054
rect 34880 3990 34944 4054
rect 34960 3990 35024 4054
rect 35040 3990 35104 4054
rect 35120 3990 35184 4054
rect 35200 3990 35264 4054
rect 35406 3990 35470 4054
rect 35486 3990 35550 4054
rect 35566 3990 35630 4054
rect 35646 3990 35710 4054
rect 35726 3990 35790 4054
rect 35806 3990 35870 4054
rect 36012 3990 36076 4054
rect 36092 3990 36156 4054
rect 36172 3990 36236 4054
rect 36252 3990 36316 4054
rect 36332 3990 36396 4054
rect 36412 3990 36476 4054
rect 36618 3990 36682 4054
rect 36698 3990 36762 4054
rect 36778 3990 36842 4054
rect 36858 3990 36922 4054
rect 36938 3990 37002 4054
rect 37018 3990 37082 4054
rect 37224 3990 37288 4054
rect 37304 3990 37368 4054
rect 37384 3990 37448 4054
rect 37464 3990 37528 4054
rect 37544 3990 37608 4054
rect 37624 3990 37688 4054
rect 37830 3990 37894 4054
rect 37910 3990 37974 4054
rect 37990 3990 38054 4054
rect 38070 3990 38134 4054
rect 38150 3990 38214 4054
rect 38230 3990 38294 4054
rect 38436 3990 38500 4054
rect 38516 3990 38580 4054
rect 38596 3990 38660 4054
rect 38676 3990 38740 4054
rect 38756 3990 38820 4054
rect 38836 3990 38900 4054
rect 39042 3990 39106 4054
rect 39122 3990 39186 4054
rect 39202 3990 39266 4054
rect 39282 3990 39346 4054
rect 39362 3990 39426 4054
rect 39442 3990 39506 4054
rect 39648 3990 39712 4054
rect 39728 3990 39792 4054
rect 39808 3990 39872 4054
rect 39888 3990 39952 4054
rect 39968 3990 40032 4054
rect 40048 3990 40112 4054
rect 40254 3990 40318 4054
rect 40334 3990 40398 4054
rect 40414 3990 40478 4054
rect 40494 3990 40558 4054
rect 40574 3990 40638 4054
rect 40654 3990 40718 4054
rect 40860 3990 40924 4054
rect 40940 3990 41004 4054
rect 41020 3990 41084 4054
rect 41100 3990 41164 4054
rect 41180 3990 41244 4054
rect 41260 3990 41324 4054
rect 41466 3990 41530 4054
rect 41546 3990 41610 4054
rect 41626 3990 41690 4054
rect 41706 3990 41770 4054
rect 41786 3990 41850 4054
rect 41866 3990 41930 4054
rect 42072 3990 42136 4054
rect 42152 3990 42216 4054
rect 42232 3990 42296 4054
rect 42312 3990 42376 4054
rect 42392 3990 42456 4054
rect 42472 3990 42536 4054
rect 42678 3990 42742 4054
rect 42758 3990 42822 4054
rect 42838 3990 42902 4054
rect 42918 3990 42982 4054
rect 42998 3990 43062 4054
rect 43078 3990 43142 4054
rect 43284 3990 43348 4054
rect 43364 3990 43428 4054
rect 43444 3990 43508 4054
rect 43524 3990 43588 4054
rect 43604 3990 43668 4054
rect 43684 3990 43748 4054
rect 43890 3990 43954 4054
rect 43970 3990 44034 4054
rect 44050 3990 44114 4054
rect 44130 3990 44194 4054
rect 44210 3990 44274 4054
rect 44290 3990 44354 4054
rect 44496 3990 44560 4054
rect 44576 3990 44640 4054
rect 44656 3990 44720 4054
rect 44736 3990 44800 4054
rect 44816 3990 44880 4054
rect 44896 3990 44960 4054
rect 45102 3990 45166 4054
rect 45182 3990 45246 4054
rect 45262 3990 45326 4054
rect 45342 3990 45406 4054
rect 45422 3990 45486 4054
rect 45502 3990 45566 4054
rect 45708 3990 45772 4054
rect 45788 3990 45852 4054
rect 45868 3990 45932 4054
rect 45948 3990 46012 4054
rect 46028 3990 46092 4054
rect 46108 3990 46172 4054
rect 46314 3990 46378 4054
rect 46394 3990 46458 4054
rect 46474 3990 46538 4054
rect 46554 3990 46618 4054
rect 46634 3990 46698 4054
rect 46714 3990 46778 4054
rect 46920 3990 46984 4054
rect 47000 3990 47064 4054
rect 47080 3990 47144 4054
rect 47160 3990 47224 4054
rect 47240 3990 47304 4054
rect 47320 3990 47384 4054
rect 47526 3990 47590 4054
rect 47606 3990 47670 4054
rect 47686 3990 47750 4054
rect 47766 3990 47830 4054
rect 47846 3990 47910 4054
rect 47926 3990 47990 4054
rect 48132 3990 48196 4054
rect 48212 3990 48276 4054
rect 48292 3990 48356 4054
rect 48372 3990 48436 4054
rect 48452 3990 48516 4054
rect 48532 3990 48596 4054
rect 48738 3990 48802 4054
rect 48818 3990 48882 4054
rect 48898 3990 48962 4054
rect 48978 3990 49042 4054
rect 49058 3990 49122 4054
rect 49138 3990 49202 4054
rect 49344 3990 49408 4054
rect 49424 3990 49488 4054
rect 49504 3990 49568 4054
rect 49584 3990 49648 4054
rect 49664 3990 49728 4054
rect 49744 3990 49808 4054
rect 49950 3990 50014 4054
rect 50030 3990 50094 4054
rect 50110 3990 50174 4054
rect 50190 3990 50254 4054
rect 50270 3990 50334 4054
rect 50350 3990 50414 4054
rect 50556 3990 50620 4054
rect 50636 3990 50700 4054
rect 50716 3990 50780 4054
rect 50796 3990 50860 4054
rect 50876 3990 50940 4054
rect 50956 3990 51020 4054
rect 51162 3990 51226 4054
rect 51242 3990 51306 4054
rect 51322 3990 51386 4054
rect 51402 3990 51466 4054
rect 51482 3990 51546 4054
rect 51562 3990 51626 4054
rect 32273 3770 32337 3834
rect 32273 3690 32337 3754
rect 32273 3610 32337 3674
rect 32273 3530 32337 3594
rect 32273 3450 32337 3514
rect 32273 3370 32337 3434
rect 32273 3290 32337 3354
rect 32273 3210 32337 3274
rect 32273 3130 32337 3194
rect 32273 3050 32337 3114
rect 32879 3770 32943 3834
rect 32879 3690 32943 3754
rect 32879 3610 32943 3674
rect 32879 3530 32943 3594
rect 32879 3450 32943 3514
rect 32879 3370 32943 3434
rect 32879 3290 32943 3354
rect 32879 3210 32943 3274
rect 32879 3130 32943 3194
rect 32879 3050 32943 3114
rect 33485 3770 33549 3834
rect 33485 3690 33549 3754
rect 33485 3610 33549 3674
rect 33485 3530 33549 3594
rect 33485 3450 33549 3514
rect 33485 3370 33549 3434
rect 33485 3290 33549 3354
rect 33485 3210 33549 3274
rect 33485 3130 33549 3194
rect 33485 3050 33549 3114
rect 34091 3770 34155 3834
rect 34091 3690 34155 3754
rect 34091 3610 34155 3674
rect 34091 3530 34155 3594
rect 34091 3450 34155 3514
rect 34091 3370 34155 3434
rect 34091 3290 34155 3354
rect 34091 3210 34155 3274
rect 34091 3130 34155 3194
rect 34091 3050 34155 3114
rect 34697 3770 34761 3834
rect 34697 3690 34761 3754
rect 34697 3610 34761 3674
rect 34697 3530 34761 3594
rect 34697 3450 34761 3514
rect 34697 3370 34761 3434
rect 34697 3290 34761 3354
rect 34697 3210 34761 3274
rect 34697 3130 34761 3194
rect 34697 3050 34761 3114
rect 35303 3770 35367 3834
rect 35303 3690 35367 3754
rect 35303 3610 35367 3674
rect 35303 3530 35367 3594
rect 35303 3450 35367 3514
rect 35303 3370 35367 3434
rect 35303 3290 35367 3354
rect 35303 3210 35367 3274
rect 35303 3130 35367 3194
rect 35303 3050 35367 3114
rect 35909 3770 35973 3834
rect 35909 3690 35973 3754
rect 35909 3610 35973 3674
rect 35909 3530 35973 3594
rect 35909 3450 35973 3514
rect 35909 3370 35973 3434
rect 35909 3290 35973 3354
rect 35909 3210 35973 3274
rect 35909 3130 35973 3194
rect 35909 3050 35973 3114
rect 36515 3770 36579 3834
rect 36515 3690 36579 3754
rect 36515 3610 36579 3674
rect 36515 3530 36579 3594
rect 36515 3450 36579 3514
rect 36515 3370 36579 3434
rect 36515 3290 36579 3354
rect 36515 3210 36579 3274
rect 36515 3130 36579 3194
rect 36515 3050 36579 3114
rect 37121 3770 37185 3834
rect 37121 3690 37185 3754
rect 37121 3610 37185 3674
rect 37121 3530 37185 3594
rect 37121 3450 37185 3514
rect 37121 3370 37185 3434
rect 37121 3290 37185 3354
rect 37121 3210 37185 3274
rect 37121 3130 37185 3194
rect 37121 3050 37185 3114
rect 37727 3770 37791 3834
rect 37727 3690 37791 3754
rect 37727 3610 37791 3674
rect 37727 3530 37791 3594
rect 37727 3450 37791 3514
rect 37727 3370 37791 3434
rect 37727 3290 37791 3354
rect 37727 3210 37791 3274
rect 37727 3130 37791 3194
rect 37727 3050 37791 3114
rect 38333 3770 38397 3834
rect 38333 3690 38397 3754
rect 38333 3610 38397 3674
rect 38333 3530 38397 3594
rect 38333 3450 38397 3514
rect 38333 3370 38397 3434
rect 38333 3290 38397 3354
rect 38333 3210 38397 3274
rect 38333 3130 38397 3194
rect 38333 3050 38397 3114
rect 38939 3770 39003 3834
rect 38939 3690 39003 3754
rect 38939 3610 39003 3674
rect 38939 3530 39003 3594
rect 38939 3450 39003 3514
rect 38939 3370 39003 3434
rect 38939 3290 39003 3354
rect 38939 3210 39003 3274
rect 38939 3130 39003 3194
rect 38939 3050 39003 3114
rect 39545 3770 39609 3834
rect 39545 3690 39609 3754
rect 39545 3610 39609 3674
rect 39545 3530 39609 3594
rect 39545 3450 39609 3514
rect 39545 3370 39609 3434
rect 39545 3290 39609 3354
rect 39545 3210 39609 3274
rect 39545 3130 39609 3194
rect 39545 3050 39609 3114
rect 40151 3770 40215 3834
rect 40151 3690 40215 3754
rect 40151 3610 40215 3674
rect 40151 3530 40215 3594
rect 40151 3450 40215 3514
rect 40151 3370 40215 3434
rect 40151 3290 40215 3354
rect 40151 3210 40215 3274
rect 40151 3130 40215 3194
rect 40151 3050 40215 3114
rect 40757 3770 40821 3834
rect 40757 3690 40821 3754
rect 40757 3610 40821 3674
rect 40757 3530 40821 3594
rect 40757 3450 40821 3514
rect 40757 3370 40821 3434
rect 40757 3290 40821 3354
rect 40757 3210 40821 3274
rect 40757 3130 40821 3194
rect 40757 3050 40821 3114
rect 41363 3770 41427 3834
rect 41363 3690 41427 3754
rect 41363 3610 41427 3674
rect 41363 3530 41427 3594
rect 41363 3450 41427 3514
rect 41363 3370 41427 3434
rect 41363 3290 41427 3354
rect 41363 3210 41427 3274
rect 41363 3130 41427 3194
rect 41363 3050 41427 3114
rect 41969 3770 42033 3834
rect 41969 3690 42033 3754
rect 41969 3610 42033 3674
rect 41969 3530 42033 3594
rect 41969 3450 42033 3514
rect 41969 3370 42033 3434
rect 41969 3290 42033 3354
rect 41969 3210 42033 3274
rect 41969 3130 42033 3194
rect 41969 3050 42033 3114
rect 42575 3770 42639 3834
rect 42575 3690 42639 3754
rect 42575 3610 42639 3674
rect 42575 3530 42639 3594
rect 42575 3450 42639 3514
rect 42575 3370 42639 3434
rect 42575 3290 42639 3354
rect 42575 3210 42639 3274
rect 42575 3130 42639 3194
rect 42575 3050 42639 3114
rect 43181 3770 43245 3834
rect 43181 3690 43245 3754
rect 43181 3610 43245 3674
rect 43181 3530 43245 3594
rect 43181 3450 43245 3514
rect 43181 3370 43245 3434
rect 43181 3290 43245 3354
rect 43181 3210 43245 3274
rect 43181 3130 43245 3194
rect 43181 3050 43245 3114
rect 43787 3770 43851 3834
rect 43787 3690 43851 3754
rect 43787 3610 43851 3674
rect 43787 3530 43851 3594
rect 43787 3450 43851 3514
rect 43787 3370 43851 3434
rect 43787 3290 43851 3354
rect 43787 3210 43851 3274
rect 43787 3130 43851 3194
rect 43787 3050 43851 3114
rect 44393 3770 44457 3834
rect 44393 3690 44457 3754
rect 44393 3610 44457 3674
rect 44393 3530 44457 3594
rect 44393 3450 44457 3514
rect 44393 3370 44457 3434
rect 44393 3290 44457 3354
rect 44393 3210 44457 3274
rect 44393 3130 44457 3194
rect 44393 3050 44457 3114
rect 44999 3770 45063 3834
rect 44999 3690 45063 3754
rect 44999 3610 45063 3674
rect 44999 3530 45063 3594
rect 44999 3450 45063 3514
rect 44999 3370 45063 3434
rect 44999 3290 45063 3354
rect 44999 3210 45063 3274
rect 44999 3130 45063 3194
rect 44999 3050 45063 3114
rect 45605 3770 45669 3834
rect 45605 3690 45669 3754
rect 45605 3610 45669 3674
rect 45605 3530 45669 3594
rect 45605 3450 45669 3514
rect 45605 3370 45669 3434
rect 45605 3290 45669 3354
rect 45605 3210 45669 3274
rect 45605 3130 45669 3194
rect 45605 3050 45669 3114
rect 46211 3770 46275 3834
rect 46211 3690 46275 3754
rect 46211 3610 46275 3674
rect 46211 3530 46275 3594
rect 46211 3450 46275 3514
rect 46211 3370 46275 3434
rect 46211 3290 46275 3354
rect 46211 3210 46275 3274
rect 46211 3130 46275 3194
rect 46211 3050 46275 3114
rect 46817 3770 46881 3834
rect 46817 3690 46881 3754
rect 46817 3610 46881 3674
rect 46817 3530 46881 3594
rect 46817 3450 46881 3514
rect 46817 3370 46881 3434
rect 46817 3290 46881 3354
rect 46817 3210 46881 3274
rect 46817 3130 46881 3194
rect 46817 3050 46881 3114
rect 47423 3770 47487 3834
rect 47423 3690 47487 3754
rect 47423 3610 47487 3674
rect 47423 3530 47487 3594
rect 47423 3450 47487 3514
rect 47423 3370 47487 3434
rect 47423 3290 47487 3354
rect 47423 3210 47487 3274
rect 47423 3130 47487 3194
rect 47423 3050 47487 3114
rect 48029 3770 48093 3834
rect 48029 3690 48093 3754
rect 48029 3610 48093 3674
rect 48029 3530 48093 3594
rect 48029 3450 48093 3514
rect 48029 3370 48093 3434
rect 48029 3290 48093 3354
rect 48029 3210 48093 3274
rect 48029 3130 48093 3194
rect 48029 3050 48093 3114
rect 48635 3770 48699 3834
rect 48635 3690 48699 3754
rect 48635 3610 48699 3674
rect 48635 3530 48699 3594
rect 48635 3450 48699 3514
rect 48635 3370 48699 3434
rect 48635 3290 48699 3354
rect 48635 3210 48699 3274
rect 48635 3130 48699 3194
rect 48635 3050 48699 3114
rect 49241 3770 49305 3834
rect 49241 3690 49305 3754
rect 49241 3610 49305 3674
rect 49241 3530 49305 3594
rect 49241 3450 49305 3514
rect 49241 3370 49305 3434
rect 49241 3290 49305 3354
rect 49241 3210 49305 3274
rect 49241 3130 49305 3194
rect 49241 3050 49305 3114
rect 49847 3770 49911 3834
rect 49847 3690 49911 3754
rect 49847 3610 49911 3674
rect 49847 3530 49911 3594
rect 49847 3450 49911 3514
rect 49847 3370 49911 3434
rect 49847 3290 49911 3354
rect 49847 3210 49911 3274
rect 49847 3130 49911 3194
rect 49847 3050 49911 3114
rect 50453 3770 50517 3834
rect 50453 3690 50517 3754
rect 50453 3610 50517 3674
rect 50453 3530 50517 3594
rect 50453 3450 50517 3514
rect 50453 3370 50517 3434
rect 50453 3290 50517 3354
rect 50453 3210 50517 3274
rect 50453 3130 50517 3194
rect 50453 3050 50517 3114
rect 51059 3770 51123 3834
rect 51059 3690 51123 3754
rect 51059 3610 51123 3674
rect 51059 3530 51123 3594
rect 51059 3450 51123 3514
rect 51059 3370 51123 3434
rect 51059 3290 51123 3354
rect 51059 3210 51123 3274
rect 51059 3130 51123 3194
rect 51059 3050 51123 3114
rect 51665 3770 51729 3834
rect 51665 3690 51729 3754
rect 51665 3610 51729 3674
rect 51665 3530 51729 3594
rect 51665 3450 51729 3514
rect 51665 3370 51729 3434
rect 51665 3290 51729 3354
rect 51665 3210 51729 3274
rect 51665 3130 51729 3194
rect 51665 3050 51729 3114
rect 32376 2830 32440 2894
rect 32456 2830 32520 2894
rect 32536 2830 32600 2894
rect 32616 2830 32680 2894
rect 32696 2830 32760 2894
rect 32776 2830 32840 2894
rect 32982 2830 33046 2894
rect 33062 2830 33126 2894
rect 33142 2830 33206 2894
rect 33222 2830 33286 2894
rect 33302 2830 33366 2894
rect 33382 2830 33446 2894
rect 33588 2830 33652 2894
rect 33668 2830 33732 2894
rect 33748 2830 33812 2894
rect 33828 2830 33892 2894
rect 33908 2830 33972 2894
rect 33988 2830 34052 2894
rect 34194 2830 34258 2894
rect 34274 2830 34338 2894
rect 34354 2830 34418 2894
rect 34434 2830 34498 2894
rect 34514 2830 34578 2894
rect 34594 2830 34658 2894
rect 34800 2830 34864 2894
rect 34880 2830 34944 2894
rect 34960 2830 35024 2894
rect 35040 2830 35104 2894
rect 35120 2830 35184 2894
rect 35200 2830 35264 2894
rect 35406 2830 35470 2894
rect 35486 2830 35550 2894
rect 35566 2830 35630 2894
rect 35646 2830 35710 2894
rect 35726 2830 35790 2894
rect 35806 2830 35870 2894
rect 36012 2830 36076 2894
rect 36092 2830 36156 2894
rect 36172 2830 36236 2894
rect 36252 2830 36316 2894
rect 36332 2830 36396 2894
rect 36412 2830 36476 2894
rect 36618 2830 36682 2894
rect 36698 2830 36762 2894
rect 36778 2830 36842 2894
rect 36858 2830 36922 2894
rect 36938 2830 37002 2894
rect 37018 2830 37082 2894
rect 37224 2830 37288 2894
rect 37304 2830 37368 2894
rect 37384 2830 37448 2894
rect 37464 2830 37528 2894
rect 37544 2830 37608 2894
rect 37624 2830 37688 2894
rect 37830 2830 37894 2894
rect 37910 2830 37974 2894
rect 37990 2830 38054 2894
rect 38070 2830 38134 2894
rect 38150 2830 38214 2894
rect 38230 2830 38294 2894
rect 38436 2830 38500 2894
rect 38516 2830 38580 2894
rect 38596 2830 38660 2894
rect 38676 2830 38740 2894
rect 38756 2830 38820 2894
rect 38836 2830 38900 2894
rect 39042 2830 39106 2894
rect 39122 2830 39186 2894
rect 39202 2830 39266 2894
rect 39282 2830 39346 2894
rect 39362 2830 39426 2894
rect 39442 2830 39506 2894
rect 39648 2830 39712 2894
rect 39728 2830 39792 2894
rect 39808 2830 39872 2894
rect 39888 2830 39952 2894
rect 39968 2830 40032 2894
rect 40048 2830 40112 2894
rect 40254 2830 40318 2894
rect 40334 2830 40398 2894
rect 40414 2830 40478 2894
rect 40494 2830 40558 2894
rect 40574 2830 40638 2894
rect 40654 2830 40718 2894
rect 40860 2830 40924 2894
rect 40940 2830 41004 2894
rect 41020 2830 41084 2894
rect 41100 2830 41164 2894
rect 41180 2830 41244 2894
rect 41260 2830 41324 2894
rect 41466 2830 41530 2894
rect 41546 2830 41610 2894
rect 41626 2830 41690 2894
rect 41706 2830 41770 2894
rect 41786 2830 41850 2894
rect 41866 2830 41930 2894
rect 42072 2830 42136 2894
rect 42152 2830 42216 2894
rect 42232 2830 42296 2894
rect 42312 2830 42376 2894
rect 42392 2830 42456 2894
rect 42472 2830 42536 2894
rect 42678 2830 42742 2894
rect 42758 2830 42822 2894
rect 42838 2830 42902 2894
rect 42918 2830 42982 2894
rect 42998 2830 43062 2894
rect 43078 2830 43142 2894
rect 43284 2830 43348 2894
rect 43364 2830 43428 2894
rect 43444 2830 43508 2894
rect 43524 2830 43588 2894
rect 43604 2830 43668 2894
rect 43684 2830 43748 2894
rect 43890 2830 43954 2894
rect 43970 2830 44034 2894
rect 44050 2830 44114 2894
rect 44130 2830 44194 2894
rect 44210 2830 44274 2894
rect 44290 2830 44354 2894
rect 44496 2830 44560 2894
rect 44576 2830 44640 2894
rect 44656 2830 44720 2894
rect 44736 2830 44800 2894
rect 44816 2830 44880 2894
rect 44896 2830 44960 2894
rect 45102 2830 45166 2894
rect 45182 2830 45246 2894
rect 45262 2830 45326 2894
rect 45342 2830 45406 2894
rect 45422 2830 45486 2894
rect 45502 2830 45566 2894
rect 45708 2830 45772 2894
rect 45788 2830 45852 2894
rect 45868 2830 45932 2894
rect 45948 2830 46012 2894
rect 46028 2830 46092 2894
rect 46108 2830 46172 2894
rect 46314 2830 46378 2894
rect 46394 2830 46458 2894
rect 46474 2830 46538 2894
rect 46554 2830 46618 2894
rect 46634 2830 46698 2894
rect 46714 2830 46778 2894
rect 46920 2830 46984 2894
rect 47000 2830 47064 2894
rect 47080 2830 47144 2894
rect 47160 2830 47224 2894
rect 47240 2830 47304 2894
rect 47320 2830 47384 2894
rect 47526 2830 47590 2894
rect 47606 2830 47670 2894
rect 47686 2830 47750 2894
rect 47766 2830 47830 2894
rect 47846 2830 47910 2894
rect 47926 2830 47990 2894
rect 48132 2830 48196 2894
rect 48212 2830 48276 2894
rect 48292 2830 48356 2894
rect 48372 2830 48436 2894
rect 48452 2830 48516 2894
rect 48532 2830 48596 2894
rect 48738 2830 48802 2894
rect 48818 2830 48882 2894
rect 48898 2830 48962 2894
rect 48978 2830 49042 2894
rect 49058 2830 49122 2894
rect 49138 2830 49202 2894
rect 49344 2830 49408 2894
rect 49424 2830 49488 2894
rect 49504 2830 49568 2894
rect 49584 2830 49648 2894
rect 49664 2830 49728 2894
rect 49744 2830 49808 2894
rect 49950 2830 50014 2894
rect 50030 2830 50094 2894
rect 50110 2830 50174 2894
rect 50190 2830 50254 2894
rect 50270 2830 50334 2894
rect 50350 2830 50414 2894
rect 50556 2830 50620 2894
rect 50636 2830 50700 2894
rect 50716 2830 50780 2894
rect 50796 2830 50860 2894
rect 50876 2830 50940 2894
rect 50956 2830 51020 2894
rect 51162 2830 51226 2894
rect 51242 2830 51306 2894
rect 51322 2830 51386 2894
rect 51402 2830 51466 2894
rect 51482 2830 51546 2894
rect 51562 2830 51626 2894
<< metal4 >>
rect 32272 5214 51730 5216
rect 32272 5150 32376 5214
rect 32440 5150 32456 5214
rect 32520 5150 32536 5214
rect 32600 5150 32616 5214
rect 32680 5150 32696 5214
rect 32760 5150 32776 5214
rect 32840 5150 32982 5214
rect 33046 5150 33062 5214
rect 33126 5150 33142 5214
rect 33206 5150 33222 5214
rect 33286 5150 33302 5214
rect 33366 5150 33382 5214
rect 33446 5150 33588 5214
rect 33652 5150 33668 5214
rect 33732 5150 33748 5214
rect 33812 5150 33828 5214
rect 33892 5150 33908 5214
rect 33972 5150 33988 5214
rect 34052 5150 34194 5214
rect 34258 5150 34274 5214
rect 34338 5150 34354 5214
rect 34418 5150 34434 5214
rect 34498 5150 34514 5214
rect 34578 5150 34594 5214
rect 34658 5150 34800 5214
rect 34864 5150 34880 5214
rect 34944 5150 34960 5214
rect 35024 5150 35040 5214
rect 35104 5150 35120 5214
rect 35184 5150 35200 5214
rect 35264 5150 35406 5214
rect 35470 5150 35486 5214
rect 35550 5150 35566 5214
rect 35630 5150 35646 5214
rect 35710 5150 35726 5214
rect 35790 5150 35806 5214
rect 35870 5150 36012 5214
rect 36076 5150 36092 5214
rect 36156 5150 36172 5214
rect 36236 5150 36252 5214
rect 36316 5150 36332 5214
rect 36396 5150 36412 5214
rect 36476 5150 36618 5214
rect 36682 5150 36698 5214
rect 36762 5150 36778 5214
rect 36842 5150 36858 5214
rect 36922 5150 36938 5214
rect 37002 5150 37018 5214
rect 37082 5150 37224 5214
rect 37288 5150 37304 5214
rect 37368 5150 37384 5214
rect 37448 5150 37464 5214
rect 37528 5150 37544 5214
rect 37608 5150 37624 5214
rect 37688 5150 37830 5214
rect 37894 5150 37910 5214
rect 37974 5150 37990 5214
rect 38054 5150 38070 5214
rect 38134 5150 38150 5214
rect 38214 5150 38230 5214
rect 38294 5150 38436 5214
rect 38500 5150 38516 5214
rect 38580 5150 38596 5214
rect 38660 5150 38676 5214
rect 38740 5150 38756 5214
rect 38820 5150 38836 5214
rect 38900 5150 39042 5214
rect 39106 5150 39122 5214
rect 39186 5150 39202 5214
rect 39266 5150 39282 5214
rect 39346 5150 39362 5214
rect 39426 5150 39442 5214
rect 39506 5150 39648 5214
rect 39712 5150 39728 5214
rect 39792 5150 39808 5214
rect 39872 5150 39888 5214
rect 39952 5150 39968 5214
rect 40032 5150 40048 5214
rect 40112 5150 40254 5214
rect 40318 5150 40334 5214
rect 40398 5150 40414 5214
rect 40478 5150 40494 5214
rect 40558 5150 40574 5214
rect 40638 5150 40654 5214
rect 40718 5150 40860 5214
rect 40924 5150 40940 5214
rect 41004 5150 41020 5214
rect 41084 5150 41100 5214
rect 41164 5150 41180 5214
rect 41244 5150 41260 5214
rect 41324 5150 41466 5214
rect 41530 5150 41546 5214
rect 41610 5150 41626 5214
rect 41690 5150 41706 5214
rect 41770 5150 41786 5214
rect 41850 5150 41866 5214
rect 41930 5150 42072 5214
rect 42136 5150 42152 5214
rect 42216 5150 42232 5214
rect 42296 5150 42312 5214
rect 42376 5150 42392 5214
rect 42456 5150 42472 5214
rect 42536 5150 42678 5214
rect 42742 5150 42758 5214
rect 42822 5150 42838 5214
rect 42902 5150 42918 5214
rect 42982 5150 42998 5214
rect 43062 5150 43078 5214
rect 43142 5150 43284 5214
rect 43348 5150 43364 5214
rect 43428 5150 43444 5214
rect 43508 5150 43524 5214
rect 43588 5150 43604 5214
rect 43668 5150 43684 5214
rect 43748 5150 43890 5214
rect 43954 5150 43970 5214
rect 44034 5150 44050 5214
rect 44114 5150 44130 5214
rect 44194 5150 44210 5214
rect 44274 5150 44290 5214
rect 44354 5150 44496 5214
rect 44560 5150 44576 5214
rect 44640 5150 44656 5214
rect 44720 5150 44736 5214
rect 44800 5150 44816 5214
rect 44880 5150 44896 5214
rect 44960 5150 45102 5214
rect 45166 5150 45182 5214
rect 45246 5150 45262 5214
rect 45326 5150 45342 5214
rect 45406 5150 45422 5214
rect 45486 5150 45502 5214
rect 45566 5150 45708 5214
rect 45772 5150 45788 5214
rect 45852 5150 45868 5214
rect 45932 5150 45948 5214
rect 46012 5150 46028 5214
rect 46092 5150 46108 5214
rect 46172 5150 46314 5214
rect 46378 5150 46394 5214
rect 46458 5150 46474 5214
rect 46538 5150 46554 5214
rect 46618 5150 46634 5214
rect 46698 5150 46714 5214
rect 46778 5150 46920 5214
rect 46984 5150 47000 5214
rect 47064 5150 47080 5214
rect 47144 5150 47160 5214
rect 47224 5150 47240 5214
rect 47304 5150 47320 5214
rect 47384 5150 47526 5214
rect 47590 5150 47606 5214
rect 47670 5150 47686 5214
rect 47750 5150 47766 5214
rect 47830 5150 47846 5214
rect 47910 5150 47926 5214
rect 47990 5150 48132 5214
rect 48196 5150 48212 5214
rect 48276 5150 48292 5214
rect 48356 5150 48372 5214
rect 48436 5150 48452 5214
rect 48516 5150 48532 5214
rect 48596 5150 48738 5214
rect 48802 5150 48818 5214
rect 48882 5150 48898 5214
rect 48962 5150 48978 5214
rect 49042 5150 49058 5214
rect 49122 5150 49138 5214
rect 49202 5150 49344 5214
rect 49408 5150 49424 5214
rect 49488 5150 49504 5214
rect 49568 5150 49584 5214
rect 49648 5150 49664 5214
rect 49728 5150 49744 5214
rect 49808 5150 49950 5214
rect 50014 5150 50030 5214
rect 50094 5150 50110 5214
rect 50174 5150 50190 5214
rect 50254 5150 50270 5214
rect 50334 5150 50350 5214
rect 50414 5150 50556 5214
rect 50620 5150 50636 5214
rect 50700 5150 50716 5214
rect 50780 5150 50796 5214
rect 50860 5150 50876 5214
rect 50940 5150 50956 5214
rect 51020 5150 51162 5214
rect 51226 5150 51242 5214
rect 51306 5150 51322 5214
rect 51386 5150 51402 5214
rect 51466 5150 51482 5214
rect 51546 5150 51562 5214
rect 51626 5150 51730 5214
rect 32272 5148 51730 5150
rect 32272 4994 32338 5148
rect 32272 4930 32273 4994
rect 32337 4930 32338 4994
rect 32272 4914 32338 4930
rect 32272 4850 32273 4914
rect 32337 4850 32338 4914
rect 32272 4834 32338 4850
rect 32272 4770 32273 4834
rect 32337 4770 32338 4834
rect 32272 4754 32338 4770
rect 32272 4690 32273 4754
rect 32337 4690 32338 4754
rect 32272 4674 32338 4690
rect 32272 4610 32273 4674
rect 32337 4610 32338 4674
rect 32272 4594 32338 4610
rect 32272 4530 32273 4594
rect 32337 4530 32338 4594
rect 32272 4514 32338 4530
rect 32272 4450 32273 4514
rect 32337 4450 32338 4514
rect 32272 4434 32338 4450
rect 32272 4370 32273 4434
rect 32337 4370 32338 4434
rect 32272 4354 32338 4370
rect 32272 4290 32273 4354
rect 32337 4290 32338 4354
rect 32272 4274 32338 4290
rect 32272 4210 32273 4274
rect 32337 4210 32338 4274
rect 32272 4120 32338 4210
rect 32398 4056 32458 5086
rect 32518 4116 32578 5148
rect 32638 4056 32698 5086
rect 32758 4116 32818 5148
rect 32878 4994 32944 5148
rect 32878 4930 32879 4994
rect 32943 4930 32944 4994
rect 32878 4914 32944 4930
rect 32878 4850 32879 4914
rect 32943 4850 32944 4914
rect 32878 4834 32944 4850
rect 32878 4770 32879 4834
rect 32943 4770 32944 4834
rect 32878 4754 32944 4770
rect 32878 4690 32879 4754
rect 32943 4690 32944 4754
rect 32878 4674 32944 4690
rect 32878 4610 32879 4674
rect 32943 4610 32944 4674
rect 32878 4594 32944 4610
rect 32878 4530 32879 4594
rect 32943 4530 32944 4594
rect 32878 4514 32944 4530
rect 32878 4450 32879 4514
rect 32943 4450 32944 4514
rect 32878 4434 32944 4450
rect 32878 4370 32879 4434
rect 32943 4370 32944 4434
rect 32878 4354 32944 4370
rect 32878 4290 32879 4354
rect 32943 4290 32944 4354
rect 32878 4274 32944 4290
rect 32878 4210 32879 4274
rect 32943 4210 32944 4274
rect 32878 4120 32944 4210
rect 33004 4056 33064 5086
rect 33124 4116 33184 5148
rect 33244 4056 33304 5086
rect 33364 4116 33424 5148
rect 33484 4994 33550 5148
rect 33484 4930 33485 4994
rect 33549 4930 33550 4994
rect 33484 4914 33550 4930
rect 33484 4850 33485 4914
rect 33549 4850 33550 4914
rect 33484 4834 33550 4850
rect 33484 4770 33485 4834
rect 33549 4770 33550 4834
rect 33484 4754 33550 4770
rect 33484 4690 33485 4754
rect 33549 4690 33550 4754
rect 33484 4674 33550 4690
rect 33484 4610 33485 4674
rect 33549 4610 33550 4674
rect 33484 4594 33550 4610
rect 33484 4530 33485 4594
rect 33549 4530 33550 4594
rect 33484 4514 33550 4530
rect 33484 4450 33485 4514
rect 33549 4450 33550 4514
rect 33484 4434 33550 4450
rect 33484 4370 33485 4434
rect 33549 4370 33550 4434
rect 33484 4354 33550 4370
rect 33484 4290 33485 4354
rect 33549 4290 33550 4354
rect 33484 4274 33550 4290
rect 33484 4210 33485 4274
rect 33549 4210 33550 4274
rect 33484 4120 33550 4210
rect 33610 4056 33670 5086
rect 33730 4116 33790 5148
rect 33850 4056 33910 5086
rect 33970 4116 34030 5148
rect 34090 4994 34156 5148
rect 34090 4930 34091 4994
rect 34155 4930 34156 4994
rect 34090 4914 34156 4930
rect 34090 4850 34091 4914
rect 34155 4850 34156 4914
rect 34090 4834 34156 4850
rect 34090 4770 34091 4834
rect 34155 4770 34156 4834
rect 34090 4754 34156 4770
rect 34090 4690 34091 4754
rect 34155 4690 34156 4754
rect 34090 4674 34156 4690
rect 34090 4610 34091 4674
rect 34155 4610 34156 4674
rect 34090 4594 34156 4610
rect 34090 4530 34091 4594
rect 34155 4530 34156 4594
rect 34090 4514 34156 4530
rect 34090 4450 34091 4514
rect 34155 4450 34156 4514
rect 34090 4434 34156 4450
rect 34090 4370 34091 4434
rect 34155 4370 34156 4434
rect 34090 4354 34156 4370
rect 34090 4290 34091 4354
rect 34155 4290 34156 4354
rect 34090 4274 34156 4290
rect 34090 4210 34091 4274
rect 34155 4210 34156 4274
rect 34090 4120 34156 4210
rect 34216 4056 34276 5086
rect 34336 4116 34396 5148
rect 34456 4056 34516 5086
rect 34576 4116 34636 5148
rect 34696 4994 34762 5148
rect 34696 4930 34697 4994
rect 34761 4930 34762 4994
rect 34696 4914 34762 4930
rect 34696 4850 34697 4914
rect 34761 4850 34762 4914
rect 34696 4834 34762 4850
rect 34696 4770 34697 4834
rect 34761 4770 34762 4834
rect 34696 4754 34762 4770
rect 34696 4690 34697 4754
rect 34761 4690 34762 4754
rect 34696 4674 34762 4690
rect 34696 4610 34697 4674
rect 34761 4610 34762 4674
rect 34696 4594 34762 4610
rect 34696 4530 34697 4594
rect 34761 4530 34762 4594
rect 34696 4514 34762 4530
rect 34696 4450 34697 4514
rect 34761 4450 34762 4514
rect 34696 4434 34762 4450
rect 34696 4370 34697 4434
rect 34761 4370 34762 4434
rect 34696 4354 34762 4370
rect 34696 4290 34697 4354
rect 34761 4290 34762 4354
rect 34696 4274 34762 4290
rect 34696 4210 34697 4274
rect 34761 4210 34762 4274
rect 34696 4120 34762 4210
rect 34822 4056 34882 5086
rect 34942 4116 35002 5148
rect 35062 4056 35122 5086
rect 35182 4116 35242 5148
rect 35302 4994 35368 5148
rect 35302 4930 35303 4994
rect 35367 4930 35368 4994
rect 35302 4914 35368 4930
rect 35302 4850 35303 4914
rect 35367 4850 35368 4914
rect 35302 4834 35368 4850
rect 35302 4770 35303 4834
rect 35367 4770 35368 4834
rect 35302 4754 35368 4770
rect 35302 4690 35303 4754
rect 35367 4690 35368 4754
rect 35302 4674 35368 4690
rect 35302 4610 35303 4674
rect 35367 4610 35368 4674
rect 35302 4594 35368 4610
rect 35302 4530 35303 4594
rect 35367 4530 35368 4594
rect 35302 4514 35368 4530
rect 35302 4450 35303 4514
rect 35367 4450 35368 4514
rect 35302 4434 35368 4450
rect 35302 4370 35303 4434
rect 35367 4370 35368 4434
rect 35302 4354 35368 4370
rect 35302 4290 35303 4354
rect 35367 4290 35368 4354
rect 35302 4274 35368 4290
rect 35302 4210 35303 4274
rect 35367 4210 35368 4274
rect 35302 4120 35368 4210
rect 35428 4056 35488 5086
rect 35548 4116 35608 5148
rect 35668 4056 35728 5086
rect 35788 4116 35848 5148
rect 35908 4994 35974 5148
rect 35908 4930 35909 4994
rect 35973 4930 35974 4994
rect 35908 4914 35974 4930
rect 35908 4850 35909 4914
rect 35973 4850 35974 4914
rect 35908 4834 35974 4850
rect 35908 4770 35909 4834
rect 35973 4770 35974 4834
rect 35908 4754 35974 4770
rect 35908 4690 35909 4754
rect 35973 4690 35974 4754
rect 35908 4674 35974 4690
rect 35908 4610 35909 4674
rect 35973 4610 35974 4674
rect 35908 4594 35974 4610
rect 35908 4530 35909 4594
rect 35973 4530 35974 4594
rect 35908 4514 35974 4530
rect 35908 4450 35909 4514
rect 35973 4450 35974 4514
rect 35908 4434 35974 4450
rect 35908 4370 35909 4434
rect 35973 4370 35974 4434
rect 35908 4354 35974 4370
rect 35908 4290 35909 4354
rect 35973 4290 35974 4354
rect 35908 4274 35974 4290
rect 35908 4210 35909 4274
rect 35973 4210 35974 4274
rect 35908 4120 35974 4210
rect 36034 4056 36094 5086
rect 36154 4116 36214 5148
rect 36274 4056 36334 5086
rect 36394 4116 36454 5148
rect 36514 4994 36580 5148
rect 36514 4930 36515 4994
rect 36579 4930 36580 4994
rect 36514 4914 36580 4930
rect 36514 4850 36515 4914
rect 36579 4850 36580 4914
rect 36514 4834 36580 4850
rect 36514 4770 36515 4834
rect 36579 4770 36580 4834
rect 36514 4754 36580 4770
rect 36514 4690 36515 4754
rect 36579 4690 36580 4754
rect 36514 4674 36580 4690
rect 36514 4610 36515 4674
rect 36579 4610 36580 4674
rect 36514 4594 36580 4610
rect 36514 4530 36515 4594
rect 36579 4530 36580 4594
rect 36514 4514 36580 4530
rect 36514 4450 36515 4514
rect 36579 4450 36580 4514
rect 36514 4434 36580 4450
rect 36514 4370 36515 4434
rect 36579 4370 36580 4434
rect 36514 4354 36580 4370
rect 36514 4290 36515 4354
rect 36579 4290 36580 4354
rect 36514 4274 36580 4290
rect 36514 4210 36515 4274
rect 36579 4210 36580 4274
rect 36514 4120 36580 4210
rect 36640 4056 36700 5086
rect 36760 4116 36820 5148
rect 36880 4056 36940 5086
rect 37000 4116 37060 5148
rect 37120 4994 37186 5148
rect 37120 4930 37121 4994
rect 37185 4930 37186 4994
rect 37120 4914 37186 4930
rect 37120 4850 37121 4914
rect 37185 4850 37186 4914
rect 37120 4834 37186 4850
rect 37120 4770 37121 4834
rect 37185 4770 37186 4834
rect 37120 4754 37186 4770
rect 37120 4690 37121 4754
rect 37185 4690 37186 4754
rect 37120 4674 37186 4690
rect 37120 4610 37121 4674
rect 37185 4610 37186 4674
rect 37120 4594 37186 4610
rect 37120 4530 37121 4594
rect 37185 4530 37186 4594
rect 37120 4514 37186 4530
rect 37120 4450 37121 4514
rect 37185 4450 37186 4514
rect 37120 4434 37186 4450
rect 37120 4370 37121 4434
rect 37185 4370 37186 4434
rect 37120 4354 37186 4370
rect 37120 4290 37121 4354
rect 37185 4290 37186 4354
rect 37120 4274 37186 4290
rect 37120 4210 37121 4274
rect 37185 4210 37186 4274
rect 37120 4120 37186 4210
rect 37246 4056 37306 5086
rect 37366 4116 37426 5148
rect 37486 4056 37546 5086
rect 37606 4116 37666 5148
rect 37726 4994 37792 5148
rect 37726 4930 37727 4994
rect 37791 4930 37792 4994
rect 37726 4914 37792 4930
rect 37726 4850 37727 4914
rect 37791 4850 37792 4914
rect 37726 4834 37792 4850
rect 37726 4770 37727 4834
rect 37791 4770 37792 4834
rect 37726 4754 37792 4770
rect 37726 4690 37727 4754
rect 37791 4690 37792 4754
rect 37726 4674 37792 4690
rect 37726 4610 37727 4674
rect 37791 4610 37792 4674
rect 37726 4594 37792 4610
rect 37726 4530 37727 4594
rect 37791 4530 37792 4594
rect 37726 4514 37792 4530
rect 37726 4450 37727 4514
rect 37791 4450 37792 4514
rect 37726 4434 37792 4450
rect 37726 4370 37727 4434
rect 37791 4370 37792 4434
rect 37726 4354 37792 4370
rect 37726 4290 37727 4354
rect 37791 4290 37792 4354
rect 37726 4274 37792 4290
rect 37726 4210 37727 4274
rect 37791 4210 37792 4274
rect 37726 4120 37792 4210
rect 37852 4056 37912 5086
rect 37972 4116 38032 5148
rect 38092 4056 38152 5086
rect 38212 4116 38272 5148
rect 38332 4994 38398 5148
rect 38332 4930 38333 4994
rect 38397 4930 38398 4994
rect 38332 4914 38398 4930
rect 38332 4850 38333 4914
rect 38397 4850 38398 4914
rect 38332 4834 38398 4850
rect 38332 4770 38333 4834
rect 38397 4770 38398 4834
rect 38332 4754 38398 4770
rect 38332 4690 38333 4754
rect 38397 4690 38398 4754
rect 38332 4674 38398 4690
rect 38332 4610 38333 4674
rect 38397 4610 38398 4674
rect 38332 4594 38398 4610
rect 38332 4530 38333 4594
rect 38397 4530 38398 4594
rect 38332 4514 38398 4530
rect 38332 4450 38333 4514
rect 38397 4450 38398 4514
rect 38332 4434 38398 4450
rect 38332 4370 38333 4434
rect 38397 4370 38398 4434
rect 38332 4354 38398 4370
rect 38332 4290 38333 4354
rect 38397 4290 38398 4354
rect 38332 4274 38398 4290
rect 38332 4210 38333 4274
rect 38397 4210 38398 4274
rect 38332 4120 38398 4210
rect 38458 4056 38518 5086
rect 38578 4116 38638 5148
rect 38698 4056 38758 5086
rect 38818 4116 38878 5148
rect 38938 4994 39004 5148
rect 38938 4930 38939 4994
rect 39003 4930 39004 4994
rect 38938 4914 39004 4930
rect 38938 4850 38939 4914
rect 39003 4850 39004 4914
rect 38938 4834 39004 4850
rect 38938 4770 38939 4834
rect 39003 4770 39004 4834
rect 38938 4754 39004 4770
rect 38938 4690 38939 4754
rect 39003 4690 39004 4754
rect 38938 4674 39004 4690
rect 38938 4610 38939 4674
rect 39003 4610 39004 4674
rect 38938 4594 39004 4610
rect 38938 4530 38939 4594
rect 39003 4530 39004 4594
rect 38938 4514 39004 4530
rect 38938 4450 38939 4514
rect 39003 4450 39004 4514
rect 38938 4434 39004 4450
rect 38938 4370 38939 4434
rect 39003 4370 39004 4434
rect 38938 4354 39004 4370
rect 38938 4290 38939 4354
rect 39003 4290 39004 4354
rect 38938 4274 39004 4290
rect 38938 4210 38939 4274
rect 39003 4210 39004 4274
rect 38938 4120 39004 4210
rect 39064 4056 39124 5086
rect 39184 4116 39244 5148
rect 39304 4056 39364 5086
rect 39424 4116 39484 5148
rect 39544 4994 39610 5148
rect 39544 4930 39545 4994
rect 39609 4930 39610 4994
rect 39544 4914 39610 4930
rect 39544 4850 39545 4914
rect 39609 4850 39610 4914
rect 39544 4834 39610 4850
rect 39544 4770 39545 4834
rect 39609 4770 39610 4834
rect 39544 4754 39610 4770
rect 39544 4690 39545 4754
rect 39609 4690 39610 4754
rect 39544 4674 39610 4690
rect 39544 4610 39545 4674
rect 39609 4610 39610 4674
rect 39544 4594 39610 4610
rect 39544 4530 39545 4594
rect 39609 4530 39610 4594
rect 39544 4514 39610 4530
rect 39544 4450 39545 4514
rect 39609 4450 39610 4514
rect 39544 4434 39610 4450
rect 39544 4370 39545 4434
rect 39609 4370 39610 4434
rect 39544 4354 39610 4370
rect 39544 4290 39545 4354
rect 39609 4290 39610 4354
rect 39544 4274 39610 4290
rect 39544 4210 39545 4274
rect 39609 4210 39610 4274
rect 39544 4120 39610 4210
rect 39670 4056 39730 5086
rect 39790 4116 39850 5148
rect 39910 4056 39970 5086
rect 40030 4116 40090 5148
rect 40150 4994 40216 5148
rect 40150 4930 40151 4994
rect 40215 4930 40216 4994
rect 40150 4914 40216 4930
rect 40150 4850 40151 4914
rect 40215 4850 40216 4914
rect 40150 4834 40216 4850
rect 40150 4770 40151 4834
rect 40215 4770 40216 4834
rect 40150 4754 40216 4770
rect 40150 4690 40151 4754
rect 40215 4690 40216 4754
rect 40150 4674 40216 4690
rect 40150 4610 40151 4674
rect 40215 4610 40216 4674
rect 40150 4594 40216 4610
rect 40150 4530 40151 4594
rect 40215 4530 40216 4594
rect 40150 4514 40216 4530
rect 40150 4450 40151 4514
rect 40215 4450 40216 4514
rect 40150 4434 40216 4450
rect 40150 4370 40151 4434
rect 40215 4370 40216 4434
rect 40150 4354 40216 4370
rect 40150 4290 40151 4354
rect 40215 4290 40216 4354
rect 40150 4274 40216 4290
rect 40150 4210 40151 4274
rect 40215 4210 40216 4274
rect 40150 4120 40216 4210
rect 40276 4056 40336 5086
rect 40396 4116 40456 5148
rect 40516 4056 40576 5086
rect 40636 4116 40696 5148
rect 40756 4994 40822 5148
rect 40756 4930 40757 4994
rect 40821 4930 40822 4994
rect 40756 4914 40822 4930
rect 40756 4850 40757 4914
rect 40821 4850 40822 4914
rect 40756 4834 40822 4850
rect 40756 4770 40757 4834
rect 40821 4770 40822 4834
rect 40756 4754 40822 4770
rect 40756 4690 40757 4754
rect 40821 4690 40822 4754
rect 40756 4674 40822 4690
rect 40756 4610 40757 4674
rect 40821 4610 40822 4674
rect 40756 4594 40822 4610
rect 40756 4530 40757 4594
rect 40821 4530 40822 4594
rect 40756 4514 40822 4530
rect 40756 4450 40757 4514
rect 40821 4450 40822 4514
rect 40756 4434 40822 4450
rect 40756 4370 40757 4434
rect 40821 4370 40822 4434
rect 40756 4354 40822 4370
rect 40756 4290 40757 4354
rect 40821 4290 40822 4354
rect 40756 4274 40822 4290
rect 40756 4210 40757 4274
rect 40821 4210 40822 4274
rect 40756 4120 40822 4210
rect 40882 4056 40942 5086
rect 41002 4116 41062 5148
rect 41122 4056 41182 5086
rect 41242 4116 41302 5148
rect 41362 4994 41428 5148
rect 41362 4930 41363 4994
rect 41427 4930 41428 4994
rect 41362 4914 41428 4930
rect 41362 4850 41363 4914
rect 41427 4850 41428 4914
rect 41362 4834 41428 4850
rect 41362 4770 41363 4834
rect 41427 4770 41428 4834
rect 41362 4754 41428 4770
rect 41362 4690 41363 4754
rect 41427 4690 41428 4754
rect 41362 4674 41428 4690
rect 41362 4610 41363 4674
rect 41427 4610 41428 4674
rect 41362 4594 41428 4610
rect 41362 4530 41363 4594
rect 41427 4530 41428 4594
rect 41362 4514 41428 4530
rect 41362 4450 41363 4514
rect 41427 4450 41428 4514
rect 41362 4434 41428 4450
rect 41362 4370 41363 4434
rect 41427 4370 41428 4434
rect 41362 4354 41428 4370
rect 41362 4290 41363 4354
rect 41427 4290 41428 4354
rect 41362 4274 41428 4290
rect 41362 4210 41363 4274
rect 41427 4210 41428 4274
rect 41362 4120 41428 4210
rect 41488 4056 41548 5086
rect 41608 4116 41668 5148
rect 41728 4056 41788 5086
rect 41848 4116 41908 5148
rect 41968 4994 42034 5148
rect 41968 4930 41969 4994
rect 42033 4930 42034 4994
rect 41968 4914 42034 4930
rect 41968 4850 41969 4914
rect 42033 4850 42034 4914
rect 41968 4834 42034 4850
rect 41968 4770 41969 4834
rect 42033 4770 42034 4834
rect 41968 4754 42034 4770
rect 41968 4690 41969 4754
rect 42033 4690 42034 4754
rect 41968 4674 42034 4690
rect 41968 4610 41969 4674
rect 42033 4610 42034 4674
rect 41968 4594 42034 4610
rect 41968 4530 41969 4594
rect 42033 4530 42034 4594
rect 41968 4514 42034 4530
rect 41968 4450 41969 4514
rect 42033 4450 42034 4514
rect 41968 4434 42034 4450
rect 41968 4370 41969 4434
rect 42033 4370 42034 4434
rect 41968 4354 42034 4370
rect 41968 4290 41969 4354
rect 42033 4290 42034 4354
rect 41968 4274 42034 4290
rect 41968 4210 41969 4274
rect 42033 4210 42034 4274
rect 41968 4120 42034 4210
rect 42094 4056 42154 5086
rect 42214 4116 42274 5148
rect 42334 4056 42394 5086
rect 42454 4116 42514 5148
rect 42574 4994 42640 5148
rect 42574 4930 42575 4994
rect 42639 4930 42640 4994
rect 42574 4914 42640 4930
rect 42574 4850 42575 4914
rect 42639 4850 42640 4914
rect 42574 4834 42640 4850
rect 42574 4770 42575 4834
rect 42639 4770 42640 4834
rect 42574 4754 42640 4770
rect 42574 4690 42575 4754
rect 42639 4690 42640 4754
rect 42574 4674 42640 4690
rect 42574 4610 42575 4674
rect 42639 4610 42640 4674
rect 42574 4594 42640 4610
rect 42574 4530 42575 4594
rect 42639 4530 42640 4594
rect 42574 4514 42640 4530
rect 42574 4450 42575 4514
rect 42639 4450 42640 4514
rect 42574 4434 42640 4450
rect 42574 4370 42575 4434
rect 42639 4370 42640 4434
rect 42574 4354 42640 4370
rect 42574 4290 42575 4354
rect 42639 4290 42640 4354
rect 42574 4274 42640 4290
rect 42574 4210 42575 4274
rect 42639 4210 42640 4274
rect 42574 4120 42640 4210
rect 42700 4056 42760 5086
rect 42820 4116 42880 5148
rect 42940 4056 43000 5086
rect 43060 4116 43120 5148
rect 43180 4994 43246 5148
rect 43180 4930 43181 4994
rect 43245 4930 43246 4994
rect 43180 4914 43246 4930
rect 43180 4850 43181 4914
rect 43245 4850 43246 4914
rect 43180 4834 43246 4850
rect 43180 4770 43181 4834
rect 43245 4770 43246 4834
rect 43180 4754 43246 4770
rect 43180 4690 43181 4754
rect 43245 4690 43246 4754
rect 43180 4674 43246 4690
rect 43180 4610 43181 4674
rect 43245 4610 43246 4674
rect 43180 4594 43246 4610
rect 43180 4530 43181 4594
rect 43245 4530 43246 4594
rect 43180 4514 43246 4530
rect 43180 4450 43181 4514
rect 43245 4450 43246 4514
rect 43180 4434 43246 4450
rect 43180 4370 43181 4434
rect 43245 4370 43246 4434
rect 43180 4354 43246 4370
rect 43180 4290 43181 4354
rect 43245 4290 43246 4354
rect 43180 4274 43246 4290
rect 43180 4210 43181 4274
rect 43245 4210 43246 4274
rect 43180 4120 43246 4210
rect 43306 4056 43366 5086
rect 43426 4116 43486 5148
rect 43546 4056 43606 5086
rect 43666 4116 43726 5148
rect 43786 4994 43852 5148
rect 43786 4930 43787 4994
rect 43851 4930 43852 4994
rect 43786 4914 43852 4930
rect 43786 4850 43787 4914
rect 43851 4850 43852 4914
rect 43786 4834 43852 4850
rect 43786 4770 43787 4834
rect 43851 4770 43852 4834
rect 43786 4754 43852 4770
rect 43786 4690 43787 4754
rect 43851 4690 43852 4754
rect 43786 4674 43852 4690
rect 43786 4610 43787 4674
rect 43851 4610 43852 4674
rect 43786 4594 43852 4610
rect 43786 4530 43787 4594
rect 43851 4530 43852 4594
rect 43786 4514 43852 4530
rect 43786 4450 43787 4514
rect 43851 4450 43852 4514
rect 43786 4434 43852 4450
rect 43786 4370 43787 4434
rect 43851 4370 43852 4434
rect 43786 4354 43852 4370
rect 43786 4290 43787 4354
rect 43851 4290 43852 4354
rect 43786 4274 43852 4290
rect 43786 4210 43787 4274
rect 43851 4210 43852 4274
rect 43786 4120 43852 4210
rect 43912 4056 43972 5086
rect 44032 4116 44092 5148
rect 44152 4056 44212 5086
rect 44272 4116 44332 5148
rect 44392 4994 44458 5148
rect 44392 4930 44393 4994
rect 44457 4930 44458 4994
rect 44392 4914 44458 4930
rect 44392 4850 44393 4914
rect 44457 4850 44458 4914
rect 44392 4834 44458 4850
rect 44392 4770 44393 4834
rect 44457 4770 44458 4834
rect 44392 4754 44458 4770
rect 44392 4690 44393 4754
rect 44457 4690 44458 4754
rect 44392 4674 44458 4690
rect 44392 4610 44393 4674
rect 44457 4610 44458 4674
rect 44392 4594 44458 4610
rect 44392 4530 44393 4594
rect 44457 4530 44458 4594
rect 44392 4514 44458 4530
rect 44392 4450 44393 4514
rect 44457 4450 44458 4514
rect 44392 4434 44458 4450
rect 44392 4370 44393 4434
rect 44457 4370 44458 4434
rect 44392 4354 44458 4370
rect 44392 4290 44393 4354
rect 44457 4290 44458 4354
rect 44392 4274 44458 4290
rect 44392 4210 44393 4274
rect 44457 4210 44458 4274
rect 44392 4120 44458 4210
rect 44518 4056 44578 5086
rect 44638 4116 44698 5148
rect 44758 4056 44818 5086
rect 44878 4116 44938 5148
rect 44998 4994 45064 5148
rect 44998 4930 44999 4994
rect 45063 4930 45064 4994
rect 44998 4914 45064 4930
rect 44998 4850 44999 4914
rect 45063 4850 45064 4914
rect 44998 4834 45064 4850
rect 44998 4770 44999 4834
rect 45063 4770 45064 4834
rect 44998 4754 45064 4770
rect 44998 4690 44999 4754
rect 45063 4690 45064 4754
rect 44998 4674 45064 4690
rect 44998 4610 44999 4674
rect 45063 4610 45064 4674
rect 44998 4594 45064 4610
rect 44998 4530 44999 4594
rect 45063 4530 45064 4594
rect 44998 4514 45064 4530
rect 44998 4450 44999 4514
rect 45063 4450 45064 4514
rect 44998 4434 45064 4450
rect 44998 4370 44999 4434
rect 45063 4370 45064 4434
rect 44998 4354 45064 4370
rect 44998 4290 44999 4354
rect 45063 4290 45064 4354
rect 44998 4274 45064 4290
rect 44998 4210 44999 4274
rect 45063 4210 45064 4274
rect 44998 4120 45064 4210
rect 45124 4056 45184 5086
rect 45244 4116 45304 5148
rect 45364 4056 45424 5086
rect 45484 4116 45544 5148
rect 45604 4994 45670 5148
rect 45604 4930 45605 4994
rect 45669 4930 45670 4994
rect 45604 4914 45670 4930
rect 45604 4850 45605 4914
rect 45669 4850 45670 4914
rect 45604 4834 45670 4850
rect 45604 4770 45605 4834
rect 45669 4770 45670 4834
rect 45604 4754 45670 4770
rect 45604 4690 45605 4754
rect 45669 4690 45670 4754
rect 45604 4674 45670 4690
rect 45604 4610 45605 4674
rect 45669 4610 45670 4674
rect 45604 4594 45670 4610
rect 45604 4530 45605 4594
rect 45669 4530 45670 4594
rect 45604 4514 45670 4530
rect 45604 4450 45605 4514
rect 45669 4450 45670 4514
rect 45604 4434 45670 4450
rect 45604 4370 45605 4434
rect 45669 4370 45670 4434
rect 45604 4354 45670 4370
rect 45604 4290 45605 4354
rect 45669 4290 45670 4354
rect 45604 4274 45670 4290
rect 45604 4210 45605 4274
rect 45669 4210 45670 4274
rect 45604 4120 45670 4210
rect 45730 4056 45790 5086
rect 45850 4116 45910 5148
rect 45970 4056 46030 5086
rect 46090 4116 46150 5148
rect 46210 4994 46276 5148
rect 46210 4930 46211 4994
rect 46275 4930 46276 4994
rect 46210 4914 46276 4930
rect 46210 4850 46211 4914
rect 46275 4850 46276 4914
rect 46210 4834 46276 4850
rect 46210 4770 46211 4834
rect 46275 4770 46276 4834
rect 46210 4754 46276 4770
rect 46210 4690 46211 4754
rect 46275 4690 46276 4754
rect 46210 4674 46276 4690
rect 46210 4610 46211 4674
rect 46275 4610 46276 4674
rect 46210 4594 46276 4610
rect 46210 4530 46211 4594
rect 46275 4530 46276 4594
rect 46210 4514 46276 4530
rect 46210 4450 46211 4514
rect 46275 4450 46276 4514
rect 46210 4434 46276 4450
rect 46210 4370 46211 4434
rect 46275 4370 46276 4434
rect 46210 4354 46276 4370
rect 46210 4290 46211 4354
rect 46275 4290 46276 4354
rect 46210 4274 46276 4290
rect 46210 4210 46211 4274
rect 46275 4210 46276 4274
rect 46210 4120 46276 4210
rect 46336 4056 46396 5086
rect 46456 4116 46516 5148
rect 46576 4056 46636 5086
rect 46696 4116 46756 5148
rect 46816 4994 46882 5148
rect 46816 4930 46817 4994
rect 46881 4930 46882 4994
rect 46816 4914 46882 4930
rect 46816 4850 46817 4914
rect 46881 4850 46882 4914
rect 46816 4834 46882 4850
rect 46816 4770 46817 4834
rect 46881 4770 46882 4834
rect 46816 4754 46882 4770
rect 46816 4690 46817 4754
rect 46881 4690 46882 4754
rect 46816 4674 46882 4690
rect 46816 4610 46817 4674
rect 46881 4610 46882 4674
rect 46816 4594 46882 4610
rect 46816 4530 46817 4594
rect 46881 4530 46882 4594
rect 46816 4514 46882 4530
rect 46816 4450 46817 4514
rect 46881 4450 46882 4514
rect 46816 4434 46882 4450
rect 46816 4370 46817 4434
rect 46881 4370 46882 4434
rect 46816 4354 46882 4370
rect 46816 4290 46817 4354
rect 46881 4290 46882 4354
rect 46816 4274 46882 4290
rect 46816 4210 46817 4274
rect 46881 4210 46882 4274
rect 46816 4120 46882 4210
rect 46942 4056 47002 5086
rect 47062 4116 47122 5148
rect 47182 4056 47242 5086
rect 47302 4116 47362 5148
rect 47422 4994 47488 5148
rect 47422 4930 47423 4994
rect 47487 4930 47488 4994
rect 47422 4914 47488 4930
rect 47422 4850 47423 4914
rect 47487 4850 47488 4914
rect 47422 4834 47488 4850
rect 47422 4770 47423 4834
rect 47487 4770 47488 4834
rect 47422 4754 47488 4770
rect 47422 4690 47423 4754
rect 47487 4690 47488 4754
rect 47422 4674 47488 4690
rect 47422 4610 47423 4674
rect 47487 4610 47488 4674
rect 47422 4594 47488 4610
rect 47422 4530 47423 4594
rect 47487 4530 47488 4594
rect 47422 4514 47488 4530
rect 47422 4450 47423 4514
rect 47487 4450 47488 4514
rect 47422 4434 47488 4450
rect 47422 4370 47423 4434
rect 47487 4370 47488 4434
rect 47422 4354 47488 4370
rect 47422 4290 47423 4354
rect 47487 4290 47488 4354
rect 47422 4274 47488 4290
rect 47422 4210 47423 4274
rect 47487 4210 47488 4274
rect 47422 4120 47488 4210
rect 47548 4056 47608 5086
rect 47668 4116 47728 5148
rect 47788 4056 47848 5086
rect 47908 4116 47968 5148
rect 48028 4994 48094 5148
rect 48028 4930 48029 4994
rect 48093 4930 48094 4994
rect 48028 4914 48094 4930
rect 48028 4850 48029 4914
rect 48093 4850 48094 4914
rect 48028 4834 48094 4850
rect 48028 4770 48029 4834
rect 48093 4770 48094 4834
rect 48028 4754 48094 4770
rect 48028 4690 48029 4754
rect 48093 4690 48094 4754
rect 48028 4674 48094 4690
rect 48028 4610 48029 4674
rect 48093 4610 48094 4674
rect 48028 4594 48094 4610
rect 48028 4530 48029 4594
rect 48093 4530 48094 4594
rect 48028 4514 48094 4530
rect 48028 4450 48029 4514
rect 48093 4450 48094 4514
rect 48028 4434 48094 4450
rect 48028 4370 48029 4434
rect 48093 4370 48094 4434
rect 48028 4354 48094 4370
rect 48028 4290 48029 4354
rect 48093 4290 48094 4354
rect 48028 4274 48094 4290
rect 48028 4210 48029 4274
rect 48093 4210 48094 4274
rect 48028 4120 48094 4210
rect 48154 4056 48214 5086
rect 48274 4116 48334 5148
rect 48394 4056 48454 5086
rect 48514 4116 48574 5148
rect 48634 4994 48700 5148
rect 48634 4930 48635 4994
rect 48699 4930 48700 4994
rect 48634 4914 48700 4930
rect 48634 4850 48635 4914
rect 48699 4850 48700 4914
rect 48634 4834 48700 4850
rect 48634 4770 48635 4834
rect 48699 4770 48700 4834
rect 48634 4754 48700 4770
rect 48634 4690 48635 4754
rect 48699 4690 48700 4754
rect 48634 4674 48700 4690
rect 48634 4610 48635 4674
rect 48699 4610 48700 4674
rect 48634 4594 48700 4610
rect 48634 4530 48635 4594
rect 48699 4530 48700 4594
rect 48634 4514 48700 4530
rect 48634 4450 48635 4514
rect 48699 4450 48700 4514
rect 48634 4434 48700 4450
rect 48634 4370 48635 4434
rect 48699 4370 48700 4434
rect 48634 4354 48700 4370
rect 48634 4290 48635 4354
rect 48699 4290 48700 4354
rect 48634 4274 48700 4290
rect 48634 4210 48635 4274
rect 48699 4210 48700 4274
rect 48634 4120 48700 4210
rect 48760 4056 48820 5086
rect 48880 4116 48940 5148
rect 49000 4056 49060 5086
rect 49120 4116 49180 5148
rect 49240 4994 49306 5148
rect 49240 4930 49241 4994
rect 49305 4930 49306 4994
rect 49240 4914 49306 4930
rect 49240 4850 49241 4914
rect 49305 4850 49306 4914
rect 49240 4834 49306 4850
rect 49240 4770 49241 4834
rect 49305 4770 49306 4834
rect 49240 4754 49306 4770
rect 49240 4690 49241 4754
rect 49305 4690 49306 4754
rect 49240 4674 49306 4690
rect 49240 4610 49241 4674
rect 49305 4610 49306 4674
rect 49240 4594 49306 4610
rect 49240 4530 49241 4594
rect 49305 4530 49306 4594
rect 49240 4514 49306 4530
rect 49240 4450 49241 4514
rect 49305 4450 49306 4514
rect 49240 4434 49306 4450
rect 49240 4370 49241 4434
rect 49305 4370 49306 4434
rect 49240 4354 49306 4370
rect 49240 4290 49241 4354
rect 49305 4290 49306 4354
rect 49240 4274 49306 4290
rect 49240 4210 49241 4274
rect 49305 4210 49306 4274
rect 49240 4120 49306 4210
rect 49366 4056 49426 5086
rect 49486 4116 49546 5148
rect 49606 4056 49666 5086
rect 49726 4116 49786 5148
rect 49846 4994 49912 5148
rect 49846 4930 49847 4994
rect 49911 4930 49912 4994
rect 49846 4914 49912 4930
rect 49846 4850 49847 4914
rect 49911 4850 49912 4914
rect 49846 4834 49912 4850
rect 49846 4770 49847 4834
rect 49911 4770 49912 4834
rect 49846 4754 49912 4770
rect 49846 4690 49847 4754
rect 49911 4690 49912 4754
rect 49846 4674 49912 4690
rect 49846 4610 49847 4674
rect 49911 4610 49912 4674
rect 49846 4594 49912 4610
rect 49846 4530 49847 4594
rect 49911 4530 49912 4594
rect 49846 4514 49912 4530
rect 49846 4450 49847 4514
rect 49911 4450 49912 4514
rect 49846 4434 49912 4450
rect 49846 4370 49847 4434
rect 49911 4370 49912 4434
rect 49846 4354 49912 4370
rect 49846 4290 49847 4354
rect 49911 4290 49912 4354
rect 49846 4274 49912 4290
rect 49846 4210 49847 4274
rect 49911 4210 49912 4274
rect 49846 4120 49912 4210
rect 49972 4056 50032 5086
rect 50092 4116 50152 5148
rect 50212 4056 50272 5086
rect 50332 4116 50392 5148
rect 50452 4994 50518 5148
rect 50452 4930 50453 4994
rect 50517 4930 50518 4994
rect 50452 4914 50518 4930
rect 50452 4850 50453 4914
rect 50517 4850 50518 4914
rect 50452 4834 50518 4850
rect 50452 4770 50453 4834
rect 50517 4770 50518 4834
rect 50452 4754 50518 4770
rect 50452 4690 50453 4754
rect 50517 4690 50518 4754
rect 50452 4674 50518 4690
rect 50452 4610 50453 4674
rect 50517 4610 50518 4674
rect 50452 4594 50518 4610
rect 50452 4530 50453 4594
rect 50517 4530 50518 4594
rect 50452 4514 50518 4530
rect 50452 4450 50453 4514
rect 50517 4450 50518 4514
rect 50452 4434 50518 4450
rect 50452 4370 50453 4434
rect 50517 4370 50518 4434
rect 50452 4354 50518 4370
rect 50452 4290 50453 4354
rect 50517 4290 50518 4354
rect 50452 4274 50518 4290
rect 50452 4210 50453 4274
rect 50517 4210 50518 4274
rect 50452 4120 50518 4210
rect 50578 4056 50638 5086
rect 50698 4116 50758 5148
rect 50818 4056 50878 5086
rect 50938 4116 50998 5148
rect 51058 4994 51124 5148
rect 51058 4930 51059 4994
rect 51123 4930 51124 4994
rect 51058 4914 51124 4930
rect 51058 4850 51059 4914
rect 51123 4850 51124 4914
rect 51058 4834 51124 4850
rect 51058 4770 51059 4834
rect 51123 4770 51124 4834
rect 51058 4754 51124 4770
rect 51058 4690 51059 4754
rect 51123 4690 51124 4754
rect 51058 4674 51124 4690
rect 51058 4610 51059 4674
rect 51123 4610 51124 4674
rect 51058 4594 51124 4610
rect 51058 4530 51059 4594
rect 51123 4530 51124 4594
rect 51058 4514 51124 4530
rect 51058 4450 51059 4514
rect 51123 4450 51124 4514
rect 51058 4434 51124 4450
rect 51058 4370 51059 4434
rect 51123 4370 51124 4434
rect 51058 4354 51124 4370
rect 51058 4290 51059 4354
rect 51123 4290 51124 4354
rect 51058 4274 51124 4290
rect 51058 4210 51059 4274
rect 51123 4210 51124 4274
rect 51058 4120 51124 4210
rect 51184 4056 51244 5086
rect 51304 4116 51364 5148
rect 51424 4056 51484 5086
rect 51544 4116 51604 5148
rect 51664 4994 51730 5148
rect 51664 4930 51665 4994
rect 51729 4930 51730 4994
rect 51664 4914 51730 4930
rect 51664 4850 51665 4914
rect 51729 4850 51730 4914
rect 51664 4834 51730 4850
rect 51664 4770 51665 4834
rect 51729 4770 51730 4834
rect 51664 4754 51730 4770
rect 51664 4690 51665 4754
rect 51729 4690 51730 4754
rect 51664 4674 51730 4690
rect 51664 4610 51665 4674
rect 51729 4610 51730 4674
rect 51664 4594 51730 4610
rect 51664 4530 51665 4594
rect 51729 4530 51730 4594
rect 51664 4514 51730 4530
rect 51664 4450 51665 4514
rect 51729 4450 51730 4514
rect 51664 4434 51730 4450
rect 51664 4370 51665 4434
rect 51729 4370 51730 4434
rect 51664 4354 51730 4370
rect 51664 4290 51665 4354
rect 51729 4290 51730 4354
rect 51664 4274 51730 4290
rect 51664 4210 51665 4274
rect 51729 4210 51730 4274
rect 51664 4120 51730 4210
rect 32272 4054 51730 4056
rect 32272 3990 32376 4054
rect 32440 3990 32456 4054
rect 32520 3990 32536 4054
rect 32600 3990 32616 4054
rect 32680 3990 32696 4054
rect 32760 3990 32776 4054
rect 32840 3990 32982 4054
rect 33046 3990 33062 4054
rect 33126 3990 33142 4054
rect 33206 3990 33222 4054
rect 33286 3990 33302 4054
rect 33366 3990 33382 4054
rect 33446 3990 33588 4054
rect 33652 3990 33668 4054
rect 33732 3990 33748 4054
rect 33812 3990 33828 4054
rect 33892 3990 33908 4054
rect 33972 3990 33988 4054
rect 34052 3990 34194 4054
rect 34258 3990 34274 4054
rect 34338 3990 34354 4054
rect 34418 3990 34434 4054
rect 34498 3990 34514 4054
rect 34578 3990 34594 4054
rect 34658 3990 34800 4054
rect 34864 3990 34880 4054
rect 34944 3990 34960 4054
rect 35024 3990 35040 4054
rect 35104 3990 35120 4054
rect 35184 3990 35200 4054
rect 35264 3990 35406 4054
rect 35470 3990 35486 4054
rect 35550 3990 35566 4054
rect 35630 3990 35646 4054
rect 35710 3990 35726 4054
rect 35790 3990 35806 4054
rect 35870 3990 36012 4054
rect 36076 3990 36092 4054
rect 36156 3990 36172 4054
rect 36236 3990 36252 4054
rect 36316 3990 36332 4054
rect 36396 3990 36412 4054
rect 36476 3990 36618 4054
rect 36682 3990 36698 4054
rect 36762 3990 36778 4054
rect 36842 3990 36858 4054
rect 36922 3990 36938 4054
rect 37002 3990 37018 4054
rect 37082 3990 37224 4054
rect 37288 3990 37304 4054
rect 37368 3990 37384 4054
rect 37448 3990 37464 4054
rect 37528 3990 37544 4054
rect 37608 3990 37624 4054
rect 37688 3990 37830 4054
rect 37894 3990 37910 4054
rect 37974 3990 37990 4054
rect 38054 3990 38070 4054
rect 38134 3990 38150 4054
rect 38214 3990 38230 4054
rect 38294 3990 38436 4054
rect 38500 3990 38516 4054
rect 38580 3990 38596 4054
rect 38660 3990 38676 4054
rect 38740 3990 38756 4054
rect 38820 3990 38836 4054
rect 38900 3990 39042 4054
rect 39106 3990 39122 4054
rect 39186 3990 39202 4054
rect 39266 3990 39282 4054
rect 39346 3990 39362 4054
rect 39426 3990 39442 4054
rect 39506 3990 39648 4054
rect 39712 3990 39728 4054
rect 39792 3990 39808 4054
rect 39872 3990 39888 4054
rect 39952 3990 39968 4054
rect 40032 3990 40048 4054
rect 40112 3990 40254 4054
rect 40318 3990 40334 4054
rect 40398 3990 40414 4054
rect 40478 3990 40494 4054
rect 40558 3990 40574 4054
rect 40638 3990 40654 4054
rect 40718 3990 40860 4054
rect 40924 3990 40940 4054
rect 41004 3990 41020 4054
rect 41084 3990 41100 4054
rect 41164 3990 41180 4054
rect 41244 3990 41260 4054
rect 41324 3990 41466 4054
rect 41530 3990 41546 4054
rect 41610 3990 41626 4054
rect 41690 3990 41706 4054
rect 41770 3990 41786 4054
rect 41850 3990 41866 4054
rect 41930 3990 42072 4054
rect 42136 3990 42152 4054
rect 42216 3990 42232 4054
rect 42296 3990 42312 4054
rect 42376 3990 42392 4054
rect 42456 3990 42472 4054
rect 42536 3990 42678 4054
rect 42742 3990 42758 4054
rect 42822 3990 42838 4054
rect 42902 3990 42918 4054
rect 42982 3990 42998 4054
rect 43062 3990 43078 4054
rect 43142 3990 43284 4054
rect 43348 3990 43364 4054
rect 43428 3990 43444 4054
rect 43508 3990 43524 4054
rect 43588 3990 43604 4054
rect 43668 3990 43684 4054
rect 43748 3990 43890 4054
rect 43954 3990 43970 4054
rect 44034 3990 44050 4054
rect 44114 3990 44130 4054
rect 44194 3990 44210 4054
rect 44274 3990 44290 4054
rect 44354 3990 44496 4054
rect 44560 3990 44576 4054
rect 44640 3990 44656 4054
rect 44720 3990 44736 4054
rect 44800 3990 44816 4054
rect 44880 3990 44896 4054
rect 44960 3990 45102 4054
rect 45166 3990 45182 4054
rect 45246 3990 45262 4054
rect 45326 3990 45342 4054
rect 45406 3990 45422 4054
rect 45486 3990 45502 4054
rect 45566 3990 45708 4054
rect 45772 3990 45788 4054
rect 45852 3990 45868 4054
rect 45932 3990 45948 4054
rect 46012 3990 46028 4054
rect 46092 3990 46108 4054
rect 46172 3990 46314 4054
rect 46378 3990 46394 4054
rect 46458 3990 46474 4054
rect 46538 3990 46554 4054
rect 46618 3990 46634 4054
rect 46698 3990 46714 4054
rect 46778 3990 46920 4054
rect 46984 3990 47000 4054
rect 47064 3990 47080 4054
rect 47144 3990 47160 4054
rect 47224 3990 47240 4054
rect 47304 3990 47320 4054
rect 47384 3990 47526 4054
rect 47590 3990 47606 4054
rect 47670 3990 47686 4054
rect 47750 3990 47766 4054
rect 47830 3990 47846 4054
rect 47910 3990 47926 4054
rect 47990 3990 48132 4054
rect 48196 3990 48212 4054
rect 48276 3990 48292 4054
rect 48356 3990 48372 4054
rect 48436 3990 48452 4054
rect 48516 3990 48532 4054
rect 48596 3990 48738 4054
rect 48802 3990 48818 4054
rect 48882 3990 48898 4054
rect 48962 3990 48978 4054
rect 49042 3990 49058 4054
rect 49122 3990 49138 4054
rect 49202 3990 49344 4054
rect 49408 3990 49424 4054
rect 49488 3990 49504 4054
rect 49568 3990 49584 4054
rect 49648 3990 49664 4054
rect 49728 3990 49744 4054
rect 49808 3990 49950 4054
rect 50014 3990 50030 4054
rect 50094 3990 50110 4054
rect 50174 3990 50190 4054
rect 50254 3990 50270 4054
rect 50334 3990 50350 4054
rect 50414 3990 50556 4054
rect 50620 3990 50636 4054
rect 50700 3990 50716 4054
rect 50780 3990 50796 4054
rect 50860 3990 50876 4054
rect 50940 3990 50956 4054
rect 51020 3990 51162 4054
rect 51226 3990 51242 4054
rect 51306 3990 51322 4054
rect 51386 3990 51402 4054
rect 51466 3990 51482 4054
rect 51546 3990 51562 4054
rect 51626 3990 51730 4054
rect 32272 3988 51730 3990
rect 32272 3834 32338 3988
rect 32272 3770 32273 3834
rect 32337 3770 32338 3834
rect 32272 3754 32338 3770
rect 32272 3690 32273 3754
rect 32337 3690 32338 3754
rect 32272 3674 32338 3690
rect 32272 3610 32273 3674
rect 32337 3610 32338 3674
rect 32272 3594 32338 3610
rect 32272 3530 32273 3594
rect 32337 3530 32338 3594
rect 32272 3514 32338 3530
rect 32272 3450 32273 3514
rect 32337 3450 32338 3514
rect 32272 3434 32338 3450
rect 32272 3370 32273 3434
rect 32337 3370 32338 3434
rect 32272 3354 32338 3370
rect 32272 3290 32273 3354
rect 32337 3290 32338 3354
rect 32272 3274 32338 3290
rect 32272 3210 32273 3274
rect 32337 3210 32338 3274
rect 32272 3194 32338 3210
rect 32272 3130 32273 3194
rect 32337 3130 32338 3194
rect 32272 3114 32338 3130
rect 32272 3050 32273 3114
rect 32337 3050 32338 3114
rect 32272 2960 32338 3050
rect 32398 2896 32458 3926
rect 32518 2956 32578 3988
rect 32638 2896 32698 3926
rect 32758 2956 32818 3988
rect 32878 3834 32944 3988
rect 32878 3770 32879 3834
rect 32943 3770 32944 3834
rect 32878 3754 32944 3770
rect 32878 3690 32879 3754
rect 32943 3690 32944 3754
rect 32878 3674 32944 3690
rect 32878 3610 32879 3674
rect 32943 3610 32944 3674
rect 32878 3594 32944 3610
rect 32878 3530 32879 3594
rect 32943 3530 32944 3594
rect 32878 3514 32944 3530
rect 32878 3450 32879 3514
rect 32943 3450 32944 3514
rect 32878 3434 32944 3450
rect 32878 3370 32879 3434
rect 32943 3370 32944 3434
rect 32878 3354 32944 3370
rect 32878 3290 32879 3354
rect 32943 3290 32944 3354
rect 32878 3274 32944 3290
rect 32878 3210 32879 3274
rect 32943 3210 32944 3274
rect 32878 3194 32944 3210
rect 32878 3130 32879 3194
rect 32943 3130 32944 3194
rect 32878 3114 32944 3130
rect 32878 3050 32879 3114
rect 32943 3050 32944 3114
rect 32878 2960 32944 3050
rect 33004 2896 33064 3926
rect 33124 2956 33184 3988
rect 33244 2896 33304 3926
rect 33364 2956 33424 3988
rect 33484 3834 33550 3988
rect 33484 3770 33485 3834
rect 33549 3770 33550 3834
rect 33484 3754 33550 3770
rect 33484 3690 33485 3754
rect 33549 3690 33550 3754
rect 33484 3674 33550 3690
rect 33484 3610 33485 3674
rect 33549 3610 33550 3674
rect 33484 3594 33550 3610
rect 33484 3530 33485 3594
rect 33549 3530 33550 3594
rect 33484 3514 33550 3530
rect 33484 3450 33485 3514
rect 33549 3450 33550 3514
rect 33484 3434 33550 3450
rect 33484 3370 33485 3434
rect 33549 3370 33550 3434
rect 33484 3354 33550 3370
rect 33484 3290 33485 3354
rect 33549 3290 33550 3354
rect 33484 3274 33550 3290
rect 33484 3210 33485 3274
rect 33549 3210 33550 3274
rect 33484 3194 33550 3210
rect 33484 3130 33485 3194
rect 33549 3130 33550 3194
rect 33484 3114 33550 3130
rect 33484 3050 33485 3114
rect 33549 3050 33550 3114
rect 33484 2960 33550 3050
rect 33610 2896 33670 3926
rect 33730 2956 33790 3988
rect 33850 2896 33910 3926
rect 33970 2956 34030 3988
rect 34090 3834 34156 3988
rect 34090 3770 34091 3834
rect 34155 3770 34156 3834
rect 34090 3754 34156 3770
rect 34090 3690 34091 3754
rect 34155 3690 34156 3754
rect 34090 3674 34156 3690
rect 34090 3610 34091 3674
rect 34155 3610 34156 3674
rect 34090 3594 34156 3610
rect 34090 3530 34091 3594
rect 34155 3530 34156 3594
rect 34090 3514 34156 3530
rect 34090 3450 34091 3514
rect 34155 3450 34156 3514
rect 34090 3434 34156 3450
rect 34090 3370 34091 3434
rect 34155 3370 34156 3434
rect 34090 3354 34156 3370
rect 34090 3290 34091 3354
rect 34155 3290 34156 3354
rect 34090 3274 34156 3290
rect 34090 3210 34091 3274
rect 34155 3210 34156 3274
rect 34090 3194 34156 3210
rect 34090 3130 34091 3194
rect 34155 3130 34156 3194
rect 34090 3114 34156 3130
rect 34090 3050 34091 3114
rect 34155 3050 34156 3114
rect 34090 2960 34156 3050
rect 34216 2896 34276 3926
rect 34336 2956 34396 3988
rect 34456 2896 34516 3926
rect 34576 2956 34636 3988
rect 34696 3834 34762 3988
rect 34696 3770 34697 3834
rect 34761 3770 34762 3834
rect 34696 3754 34762 3770
rect 34696 3690 34697 3754
rect 34761 3690 34762 3754
rect 34696 3674 34762 3690
rect 34696 3610 34697 3674
rect 34761 3610 34762 3674
rect 34696 3594 34762 3610
rect 34696 3530 34697 3594
rect 34761 3530 34762 3594
rect 34696 3514 34762 3530
rect 34696 3450 34697 3514
rect 34761 3450 34762 3514
rect 34696 3434 34762 3450
rect 34696 3370 34697 3434
rect 34761 3370 34762 3434
rect 34696 3354 34762 3370
rect 34696 3290 34697 3354
rect 34761 3290 34762 3354
rect 34696 3274 34762 3290
rect 34696 3210 34697 3274
rect 34761 3210 34762 3274
rect 34696 3194 34762 3210
rect 34696 3130 34697 3194
rect 34761 3130 34762 3194
rect 34696 3114 34762 3130
rect 34696 3050 34697 3114
rect 34761 3050 34762 3114
rect 34696 2960 34762 3050
rect 34822 2896 34882 3926
rect 34942 2956 35002 3988
rect 35062 2896 35122 3926
rect 35182 2956 35242 3988
rect 35302 3834 35368 3988
rect 35302 3770 35303 3834
rect 35367 3770 35368 3834
rect 35302 3754 35368 3770
rect 35302 3690 35303 3754
rect 35367 3690 35368 3754
rect 35302 3674 35368 3690
rect 35302 3610 35303 3674
rect 35367 3610 35368 3674
rect 35302 3594 35368 3610
rect 35302 3530 35303 3594
rect 35367 3530 35368 3594
rect 35302 3514 35368 3530
rect 35302 3450 35303 3514
rect 35367 3450 35368 3514
rect 35302 3434 35368 3450
rect 35302 3370 35303 3434
rect 35367 3370 35368 3434
rect 35302 3354 35368 3370
rect 35302 3290 35303 3354
rect 35367 3290 35368 3354
rect 35302 3274 35368 3290
rect 35302 3210 35303 3274
rect 35367 3210 35368 3274
rect 35302 3194 35368 3210
rect 35302 3130 35303 3194
rect 35367 3130 35368 3194
rect 35302 3114 35368 3130
rect 35302 3050 35303 3114
rect 35367 3050 35368 3114
rect 35302 2960 35368 3050
rect 35428 2896 35488 3926
rect 35548 2956 35608 3988
rect 35668 2896 35728 3926
rect 35788 2956 35848 3988
rect 35908 3834 35974 3988
rect 35908 3770 35909 3834
rect 35973 3770 35974 3834
rect 35908 3754 35974 3770
rect 35908 3690 35909 3754
rect 35973 3690 35974 3754
rect 35908 3674 35974 3690
rect 35908 3610 35909 3674
rect 35973 3610 35974 3674
rect 35908 3594 35974 3610
rect 35908 3530 35909 3594
rect 35973 3530 35974 3594
rect 35908 3514 35974 3530
rect 35908 3450 35909 3514
rect 35973 3450 35974 3514
rect 35908 3434 35974 3450
rect 35908 3370 35909 3434
rect 35973 3370 35974 3434
rect 35908 3354 35974 3370
rect 35908 3290 35909 3354
rect 35973 3290 35974 3354
rect 35908 3274 35974 3290
rect 35908 3210 35909 3274
rect 35973 3210 35974 3274
rect 35908 3194 35974 3210
rect 35908 3130 35909 3194
rect 35973 3130 35974 3194
rect 35908 3114 35974 3130
rect 35908 3050 35909 3114
rect 35973 3050 35974 3114
rect 35908 2960 35974 3050
rect 36034 2896 36094 3926
rect 36154 2956 36214 3988
rect 36274 2896 36334 3926
rect 36394 2956 36454 3988
rect 36514 3834 36580 3988
rect 36514 3770 36515 3834
rect 36579 3770 36580 3834
rect 36514 3754 36580 3770
rect 36514 3690 36515 3754
rect 36579 3690 36580 3754
rect 36514 3674 36580 3690
rect 36514 3610 36515 3674
rect 36579 3610 36580 3674
rect 36514 3594 36580 3610
rect 36514 3530 36515 3594
rect 36579 3530 36580 3594
rect 36514 3514 36580 3530
rect 36514 3450 36515 3514
rect 36579 3450 36580 3514
rect 36514 3434 36580 3450
rect 36514 3370 36515 3434
rect 36579 3370 36580 3434
rect 36514 3354 36580 3370
rect 36514 3290 36515 3354
rect 36579 3290 36580 3354
rect 36514 3274 36580 3290
rect 36514 3210 36515 3274
rect 36579 3210 36580 3274
rect 36514 3194 36580 3210
rect 36514 3130 36515 3194
rect 36579 3130 36580 3194
rect 36514 3114 36580 3130
rect 36514 3050 36515 3114
rect 36579 3050 36580 3114
rect 36514 2960 36580 3050
rect 36640 2896 36700 3926
rect 36760 2956 36820 3988
rect 36880 2896 36940 3926
rect 37000 2956 37060 3988
rect 37120 3834 37186 3988
rect 37120 3770 37121 3834
rect 37185 3770 37186 3834
rect 37120 3754 37186 3770
rect 37120 3690 37121 3754
rect 37185 3690 37186 3754
rect 37120 3674 37186 3690
rect 37120 3610 37121 3674
rect 37185 3610 37186 3674
rect 37120 3594 37186 3610
rect 37120 3530 37121 3594
rect 37185 3530 37186 3594
rect 37120 3514 37186 3530
rect 37120 3450 37121 3514
rect 37185 3450 37186 3514
rect 37120 3434 37186 3450
rect 37120 3370 37121 3434
rect 37185 3370 37186 3434
rect 37120 3354 37186 3370
rect 37120 3290 37121 3354
rect 37185 3290 37186 3354
rect 37120 3274 37186 3290
rect 37120 3210 37121 3274
rect 37185 3210 37186 3274
rect 37120 3194 37186 3210
rect 37120 3130 37121 3194
rect 37185 3130 37186 3194
rect 37120 3114 37186 3130
rect 37120 3050 37121 3114
rect 37185 3050 37186 3114
rect 37120 2960 37186 3050
rect 37246 2896 37306 3926
rect 37366 2956 37426 3988
rect 37486 2896 37546 3926
rect 37606 2956 37666 3988
rect 37726 3834 37792 3988
rect 37726 3770 37727 3834
rect 37791 3770 37792 3834
rect 37726 3754 37792 3770
rect 37726 3690 37727 3754
rect 37791 3690 37792 3754
rect 37726 3674 37792 3690
rect 37726 3610 37727 3674
rect 37791 3610 37792 3674
rect 37726 3594 37792 3610
rect 37726 3530 37727 3594
rect 37791 3530 37792 3594
rect 37726 3514 37792 3530
rect 37726 3450 37727 3514
rect 37791 3450 37792 3514
rect 37726 3434 37792 3450
rect 37726 3370 37727 3434
rect 37791 3370 37792 3434
rect 37726 3354 37792 3370
rect 37726 3290 37727 3354
rect 37791 3290 37792 3354
rect 37726 3274 37792 3290
rect 37726 3210 37727 3274
rect 37791 3210 37792 3274
rect 37726 3194 37792 3210
rect 37726 3130 37727 3194
rect 37791 3130 37792 3194
rect 37726 3114 37792 3130
rect 37726 3050 37727 3114
rect 37791 3050 37792 3114
rect 37726 2960 37792 3050
rect 37852 2896 37912 3926
rect 37972 2956 38032 3988
rect 38092 2896 38152 3926
rect 38212 2956 38272 3988
rect 38332 3834 38398 3988
rect 38332 3770 38333 3834
rect 38397 3770 38398 3834
rect 38332 3754 38398 3770
rect 38332 3690 38333 3754
rect 38397 3690 38398 3754
rect 38332 3674 38398 3690
rect 38332 3610 38333 3674
rect 38397 3610 38398 3674
rect 38332 3594 38398 3610
rect 38332 3530 38333 3594
rect 38397 3530 38398 3594
rect 38332 3514 38398 3530
rect 38332 3450 38333 3514
rect 38397 3450 38398 3514
rect 38332 3434 38398 3450
rect 38332 3370 38333 3434
rect 38397 3370 38398 3434
rect 38332 3354 38398 3370
rect 38332 3290 38333 3354
rect 38397 3290 38398 3354
rect 38332 3274 38398 3290
rect 38332 3210 38333 3274
rect 38397 3210 38398 3274
rect 38332 3194 38398 3210
rect 38332 3130 38333 3194
rect 38397 3130 38398 3194
rect 38332 3114 38398 3130
rect 38332 3050 38333 3114
rect 38397 3050 38398 3114
rect 38332 2960 38398 3050
rect 38458 2896 38518 3926
rect 38578 2956 38638 3988
rect 38698 2896 38758 3926
rect 38818 2956 38878 3988
rect 38938 3834 39004 3988
rect 38938 3770 38939 3834
rect 39003 3770 39004 3834
rect 38938 3754 39004 3770
rect 38938 3690 38939 3754
rect 39003 3690 39004 3754
rect 38938 3674 39004 3690
rect 38938 3610 38939 3674
rect 39003 3610 39004 3674
rect 38938 3594 39004 3610
rect 38938 3530 38939 3594
rect 39003 3530 39004 3594
rect 38938 3514 39004 3530
rect 38938 3450 38939 3514
rect 39003 3450 39004 3514
rect 38938 3434 39004 3450
rect 38938 3370 38939 3434
rect 39003 3370 39004 3434
rect 38938 3354 39004 3370
rect 38938 3290 38939 3354
rect 39003 3290 39004 3354
rect 38938 3274 39004 3290
rect 38938 3210 38939 3274
rect 39003 3210 39004 3274
rect 38938 3194 39004 3210
rect 38938 3130 38939 3194
rect 39003 3130 39004 3194
rect 38938 3114 39004 3130
rect 38938 3050 38939 3114
rect 39003 3050 39004 3114
rect 38938 2960 39004 3050
rect 39064 2896 39124 3926
rect 39184 2956 39244 3988
rect 39304 2896 39364 3926
rect 39424 2956 39484 3988
rect 39544 3834 39610 3988
rect 39544 3770 39545 3834
rect 39609 3770 39610 3834
rect 39544 3754 39610 3770
rect 39544 3690 39545 3754
rect 39609 3690 39610 3754
rect 39544 3674 39610 3690
rect 39544 3610 39545 3674
rect 39609 3610 39610 3674
rect 39544 3594 39610 3610
rect 39544 3530 39545 3594
rect 39609 3530 39610 3594
rect 39544 3514 39610 3530
rect 39544 3450 39545 3514
rect 39609 3450 39610 3514
rect 39544 3434 39610 3450
rect 39544 3370 39545 3434
rect 39609 3370 39610 3434
rect 39544 3354 39610 3370
rect 39544 3290 39545 3354
rect 39609 3290 39610 3354
rect 39544 3274 39610 3290
rect 39544 3210 39545 3274
rect 39609 3210 39610 3274
rect 39544 3194 39610 3210
rect 39544 3130 39545 3194
rect 39609 3130 39610 3194
rect 39544 3114 39610 3130
rect 39544 3050 39545 3114
rect 39609 3050 39610 3114
rect 39544 2960 39610 3050
rect 39670 2896 39730 3926
rect 39790 2956 39850 3988
rect 39910 2896 39970 3926
rect 40030 2956 40090 3988
rect 40150 3834 40216 3988
rect 40150 3770 40151 3834
rect 40215 3770 40216 3834
rect 40150 3754 40216 3770
rect 40150 3690 40151 3754
rect 40215 3690 40216 3754
rect 40150 3674 40216 3690
rect 40150 3610 40151 3674
rect 40215 3610 40216 3674
rect 40150 3594 40216 3610
rect 40150 3530 40151 3594
rect 40215 3530 40216 3594
rect 40150 3514 40216 3530
rect 40150 3450 40151 3514
rect 40215 3450 40216 3514
rect 40150 3434 40216 3450
rect 40150 3370 40151 3434
rect 40215 3370 40216 3434
rect 40150 3354 40216 3370
rect 40150 3290 40151 3354
rect 40215 3290 40216 3354
rect 40150 3274 40216 3290
rect 40150 3210 40151 3274
rect 40215 3210 40216 3274
rect 40150 3194 40216 3210
rect 40150 3130 40151 3194
rect 40215 3130 40216 3194
rect 40150 3114 40216 3130
rect 40150 3050 40151 3114
rect 40215 3050 40216 3114
rect 40150 2960 40216 3050
rect 40276 2896 40336 3926
rect 40396 2956 40456 3988
rect 40516 2896 40576 3926
rect 40636 2956 40696 3988
rect 40756 3834 40822 3988
rect 40756 3770 40757 3834
rect 40821 3770 40822 3834
rect 40756 3754 40822 3770
rect 40756 3690 40757 3754
rect 40821 3690 40822 3754
rect 40756 3674 40822 3690
rect 40756 3610 40757 3674
rect 40821 3610 40822 3674
rect 40756 3594 40822 3610
rect 40756 3530 40757 3594
rect 40821 3530 40822 3594
rect 40756 3514 40822 3530
rect 40756 3450 40757 3514
rect 40821 3450 40822 3514
rect 40756 3434 40822 3450
rect 40756 3370 40757 3434
rect 40821 3370 40822 3434
rect 40756 3354 40822 3370
rect 40756 3290 40757 3354
rect 40821 3290 40822 3354
rect 40756 3274 40822 3290
rect 40756 3210 40757 3274
rect 40821 3210 40822 3274
rect 40756 3194 40822 3210
rect 40756 3130 40757 3194
rect 40821 3130 40822 3194
rect 40756 3114 40822 3130
rect 40756 3050 40757 3114
rect 40821 3050 40822 3114
rect 40756 2960 40822 3050
rect 40882 2896 40942 3926
rect 41002 2956 41062 3988
rect 41122 2896 41182 3926
rect 41242 2956 41302 3988
rect 41362 3834 41428 3988
rect 41362 3770 41363 3834
rect 41427 3770 41428 3834
rect 41362 3754 41428 3770
rect 41362 3690 41363 3754
rect 41427 3690 41428 3754
rect 41362 3674 41428 3690
rect 41362 3610 41363 3674
rect 41427 3610 41428 3674
rect 41362 3594 41428 3610
rect 41362 3530 41363 3594
rect 41427 3530 41428 3594
rect 41362 3514 41428 3530
rect 41362 3450 41363 3514
rect 41427 3450 41428 3514
rect 41362 3434 41428 3450
rect 41362 3370 41363 3434
rect 41427 3370 41428 3434
rect 41362 3354 41428 3370
rect 41362 3290 41363 3354
rect 41427 3290 41428 3354
rect 41362 3274 41428 3290
rect 41362 3210 41363 3274
rect 41427 3210 41428 3274
rect 41362 3194 41428 3210
rect 41362 3130 41363 3194
rect 41427 3130 41428 3194
rect 41362 3114 41428 3130
rect 41362 3050 41363 3114
rect 41427 3050 41428 3114
rect 41362 2960 41428 3050
rect 41488 2896 41548 3926
rect 41608 2956 41668 3988
rect 41728 2896 41788 3926
rect 41848 2956 41908 3988
rect 41968 3834 42034 3988
rect 41968 3770 41969 3834
rect 42033 3770 42034 3834
rect 41968 3754 42034 3770
rect 41968 3690 41969 3754
rect 42033 3690 42034 3754
rect 41968 3674 42034 3690
rect 41968 3610 41969 3674
rect 42033 3610 42034 3674
rect 41968 3594 42034 3610
rect 41968 3530 41969 3594
rect 42033 3530 42034 3594
rect 41968 3514 42034 3530
rect 41968 3450 41969 3514
rect 42033 3450 42034 3514
rect 41968 3434 42034 3450
rect 41968 3370 41969 3434
rect 42033 3370 42034 3434
rect 41968 3354 42034 3370
rect 41968 3290 41969 3354
rect 42033 3290 42034 3354
rect 41968 3274 42034 3290
rect 41968 3210 41969 3274
rect 42033 3210 42034 3274
rect 41968 3194 42034 3210
rect 41968 3130 41969 3194
rect 42033 3130 42034 3194
rect 41968 3114 42034 3130
rect 41968 3050 41969 3114
rect 42033 3050 42034 3114
rect 41968 2960 42034 3050
rect 42094 2896 42154 3926
rect 42214 2956 42274 3988
rect 42334 2896 42394 3926
rect 42454 2956 42514 3988
rect 42574 3834 42640 3988
rect 42574 3770 42575 3834
rect 42639 3770 42640 3834
rect 42574 3754 42640 3770
rect 42574 3690 42575 3754
rect 42639 3690 42640 3754
rect 42574 3674 42640 3690
rect 42574 3610 42575 3674
rect 42639 3610 42640 3674
rect 42574 3594 42640 3610
rect 42574 3530 42575 3594
rect 42639 3530 42640 3594
rect 42574 3514 42640 3530
rect 42574 3450 42575 3514
rect 42639 3450 42640 3514
rect 42574 3434 42640 3450
rect 42574 3370 42575 3434
rect 42639 3370 42640 3434
rect 42574 3354 42640 3370
rect 42574 3290 42575 3354
rect 42639 3290 42640 3354
rect 42574 3274 42640 3290
rect 42574 3210 42575 3274
rect 42639 3210 42640 3274
rect 42574 3194 42640 3210
rect 42574 3130 42575 3194
rect 42639 3130 42640 3194
rect 42574 3114 42640 3130
rect 42574 3050 42575 3114
rect 42639 3050 42640 3114
rect 42574 2960 42640 3050
rect 42700 2896 42760 3926
rect 42820 2956 42880 3988
rect 42940 2896 43000 3926
rect 43060 2956 43120 3988
rect 43180 3834 43246 3988
rect 43180 3770 43181 3834
rect 43245 3770 43246 3834
rect 43180 3754 43246 3770
rect 43180 3690 43181 3754
rect 43245 3690 43246 3754
rect 43180 3674 43246 3690
rect 43180 3610 43181 3674
rect 43245 3610 43246 3674
rect 43180 3594 43246 3610
rect 43180 3530 43181 3594
rect 43245 3530 43246 3594
rect 43180 3514 43246 3530
rect 43180 3450 43181 3514
rect 43245 3450 43246 3514
rect 43180 3434 43246 3450
rect 43180 3370 43181 3434
rect 43245 3370 43246 3434
rect 43180 3354 43246 3370
rect 43180 3290 43181 3354
rect 43245 3290 43246 3354
rect 43180 3274 43246 3290
rect 43180 3210 43181 3274
rect 43245 3210 43246 3274
rect 43180 3194 43246 3210
rect 43180 3130 43181 3194
rect 43245 3130 43246 3194
rect 43180 3114 43246 3130
rect 43180 3050 43181 3114
rect 43245 3050 43246 3114
rect 43180 2960 43246 3050
rect 43306 2896 43366 3926
rect 43426 2956 43486 3988
rect 43546 2896 43606 3926
rect 43666 2956 43726 3988
rect 43786 3834 43852 3988
rect 43786 3770 43787 3834
rect 43851 3770 43852 3834
rect 43786 3754 43852 3770
rect 43786 3690 43787 3754
rect 43851 3690 43852 3754
rect 43786 3674 43852 3690
rect 43786 3610 43787 3674
rect 43851 3610 43852 3674
rect 43786 3594 43852 3610
rect 43786 3530 43787 3594
rect 43851 3530 43852 3594
rect 43786 3514 43852 3530
rect 43786 3450 43787 3514
rect 43851 3450 43852 3514
rect 43786 3434 43852 3450
rect 43786 3370 43787 3434
rect 43851 3370 43852 3434
rect 43786 3354 43852 3370
rect 43786 3290 43787 3354
rect 43851 3290 43852 3354
rect 43786 3274 43852 3290
rect 43786 3210 43787 3274
rect 43851 3210 43852 3274
rect 43786 3194 43852 3210
rect 43786 3130 43787 3194
rect 43851 3130 43852 3194
rect 43786 3114 43852 3130
rect 43786 3050 43787 3114
rect 43851 3050 43852 3114
rect 43786 2960 43852 3050
rect 43912 2896 43972 3926
rect 44032 2956 44092 3988
rect 44152 2896 44212 3926
rect 44272 2956 44332 3988
rect 44392 3834 44458 3988
rect 44392 3770 44393 3834
rect 44457 3770 44458 3834
rect 44392 3754 44458 3770
rect 44392 3690 44393 3754
rect 44457 3690 44458 3754
rect 44392 3674 44458 3690
rect 44392 3610 44393 3674
rect 44457 3610 44458 3674
rect 44392 3594 44458 3610
rect 44392 3530 44393 3594
rect 44457 3530 44458 3594
rect 44392 3514 44458 3530
rect 44392 3450 44393 3514
rect 44457 3450 44458 3514
rect 44392 3434 44458 3450
rect 44392 3370 44393 3434
rect 44457 3370 44458 3434
rect 44392 3354 44458 3370
rect 44392 3290 44393 3354
rect 44457 3290 44458 3354
rect 44392 3274 44458 3290
rect 44392 3210 44393 3274
rect 44457 3210 44458 3274
rect 44392 3194 44458 3210
rect 44392 3130 44393 3194
rect 44457 3130 44458 3194
rect 44392 3114 44458 3130
rect 44392 3050 44393 3114
rect 44457 3050 44458 3114
rect 44392 2960 44458 3050
rect 44518 2896 44578 3926
rect 44638 2956 44698 3988
rect 44758 2896 44818 3926
rect 44878 2956 44938 3988
rect 44998 3834 45064 3988
rect 44998 3770 44999 3834
rect 45063 3770 45064 3834
rect 44998 3754 45064 3770
rect 44998 3690 44999 3754
rect 45063 3690 45064 3754
rect 44998 3674 45064 3690
rect 44998 3610 44999 3674
rect 45063 3610 45064 3674
rect 44998 3594 45064 3610
rect 44998 3530 44999 3594
rect 45063 3530 45064 3594
rect 44998 3514 45064 3530
rect 44998 3450 44999 3514
rect 45063 3450 45064 3514
rect 44998 3434 45064 3450
rect 44998 3370 44999 3434
rect 45063 3370 45064 3434
rect 44998 3354 45064 3370
rect 44998 3290 44999 3354
rect 45063 3290 45064 3354
rect 44998 3274 45064 3290
rect 44998 3210 44999 3274
rect 45063 3210 45064 3274
rect 44998 3194 45064 3210
rect 44998 3130 44999 3194
rect 45063 3130 45064 3194
rect 44998 3114 45064 3130
rect 44998 3050 44999 3114
rect 45063 3050 45064 3114
rect 44998 2960 45064 3050
rect 45124 2896 45184 3926
rect 45244 2956 45304 3988
rect 45364 2896 45424 3926
rect 45484 2956 45544 3988
rect 45604 3834 45670 3988
rect 45604 3770 45605 3834
rect 45669 3770 45670 3834
rect 45604 3754 45670 3770
rect 45604 3690 45605 3754
rect 45669 3690 45670 3754
rect 45604 3674 45670 3690
rect 45604 3610 45605 3674
rect 45669 3610 45670 3674
rect 45604 3594 45670 3610
rect 45604 3530 45605 3594
rect 45669 3530 45670 3594
rect 45604 3514 45670 3530
rect 45604 3450 45605 3514
rect 45669 3450 45670 3514
rect 45604 3434 45670 3450
rect 45604 3370 45605 3434
rect 45669 3370 45670 3434
rect 45604 3354 45670 3370
rect 45604 3290 45605 3354
rect 45669 3290 45670 3354
rect 45604 3274 45670 3290
rect 45604 3210 45605 3274
rect 45669 3210 45670 3274
rect 45604 3194 45670 3210
rect 45604 3130 45605 3194
rect 45669 3130 45670 3194
rect 45604 3114 45670 3130
rect 45604 3050 45605 3114
rect 45669 3050 45670 3114
rect 45604 2960 45670 3050
rect 45730 2896 45790 3926
rect 45850 2956 45910 3988
rect 45970 2896 46030 3926
rect 46090 2956 46150 3988
rect 46210 3834 46276 3988
rect 46210 3770 46211 3834
rect 46275 3770 46276 3834
rect 46210 3754 46276 3770
rect 46210 3690 46211 3754
rect 46275 3690 46276 3754
rect 46210 3674 46276 3690
rect 46210 3610 46211 3674
rect 46275 3610 46276 3674
rect 46210 3594 46276 3610
rect 46210 3530 46211 3594
rect 46275 3530 46276 3594
rect 46210 3514 46276 3530
rect 46210 3450 46211 3514
rect 46275 3450 46276 3514
rect 46210 3434 46276 3450
rect 46210 3370 46211 3434
rect 46275 3370 46276 3434
rect 46210 3354 46276 3370
rect 46210 3290 46211 3354
rect 46275 3290 46276 3354
rect 46210 3274 46276 3290
rect 46210 3210 46211 3274
rect 46275 3210 46276 3274
rect 46210 3194 46276 3210
rect 46210 3130 46211 3194
rect 46275 3130 46276 3194
rect 46210 3114 46276 3130
rect 46210 3050 46211 3114
rect 46275 3050 46276 3114
rect 46210 2960 46276 3050
rect 46336 2896 46396 3926
rect 46456 2956 46516 3988
rect 46576 2896 46636 3926
rect 46696 2956 46756 3988
rect 46816 3834 46882 3988
rect 46816 3770 46817 3834
rect 46881 3770 46882 3834
rect 46816 3754 46882 3770
rect 46816 3690 46817 3754
rect 46881 3690 46882 3754
rect 46816 3674 46882 3690
rect 46816 3610 46817 3674
rect 46881 3610 46882 3674
rect 46816 3594 46882 3610
rect 46816 3530 46817 3594
rect 46881 3530 46882 3594
rect 46816 3514 46882 3530
rect 46816 3450 46817 3514
rect 46881 3450 46882 3514
rect 46816 3434 46882 3450
rect 46816 3370 46817 3434
rect 46881 3370 46882 3434
rect 46816 3354 46882 3370
rect 46816 3290 46817 3354
rect 46881 3290 46882 3354
rect 46816 3274 46882 3290
rect 46816 3210 46817 3274
rect 46881 3210 46882 3274
rect 46816 3194 46882 3210
rect 46816 3130 46817 3194
rect 46881 3130 46882 3194
rect 46816 3114 46882 3130
rect 46816 3050 46817 3114
rect 46881 3050 46882 3114
rect 46816 2960 46882 3050
rect 46942 2896 47002 3926
rect 47062 2956 47122 3988
rect 47182 2896 47242 3926
rect 47302 2956 47362 3988
rect 47422 3834 47488 3988
rect 47422 3770 47423 3834
rect 47487 3770 47488 3834
rect 47422 3754 47488 3770
rect 47422 3690 47423 3754
rect 47487 3690 47488 3754
rect 47422 3674 47488 3690
rect 47422 3610 47423 3674
rect 47487 3610 47488 3674
rect 47422 3594 47488 3610
rect 47422 3530 47423 3594
rect 47487 3530 47488 3594
rect 47422 3514 47488 3530
rect 47422 3450 47423 3514
rect 47487 3450 47488 3514
rect 47422 3434 47488 3450
rect 47422 3370 47423 3434
rect 47487 3370 47488 3434
rect 47422 3354 47488 3370
rect 47422 3290 47423 3354
rect 47487 3290 47488 3354
rect 47422 3274 47488 3290
rect 47422 3210 47423 3274
rect 47487 3210 47488 3274
rect 47422 3194 47488 3210
rect 47422 3130 47423 3194
rect 47487 3130 47488 3194
rect 47422 3114 47488 3130
rect 47422 3050 47423 3114
rect 47487 3050 47488 3114
rect 47422 2960 47488 3050
rect 47548 2896 47608 3926
rect 47668 2956 47728 3988
rect 47788 2896 47848 3926
rect 47908 2956 47968 3988
rect 48028 3834 48094 3988
rect 48028 3770 48029 3834
rect 48093 3770 48094 3834
rect 48028 3754 48094 3770
rect 48028 3690 48029 3754
rect 48093 3690 48094 3754
rect 48028 3674 48094 3690
rect 48028 3610 48029 3674
rect 48093 3610 48094 3674
rect 48028 3594 48094 3610
rect 48028 3530 48029 3594
rect 48093 3530 48094 3594
rect 48028 3514 48094 3530
rect 48028 3450 48029 3514
rect 48093 3450 48094 3514
rect 48028 3434 48094 3450
rect 48028 3370 48029 3434
rect 48093 3370 48094 3434
rect 48028 3354 48094 3370
rect 48028 3290 48029 3354
rect 48093 3290 48094 3354
rect 48028 3274 48094 3290
rect 48028 3210 48029 3274
rect 48093 3210 48094 3274
rect 48028 3194 48094 3210
rect 48028 3130 48029 3194
rect 48093 3130 48094 3194
rect 48028 3114 48094 3130
rect 48028 3050 48029 3114
rect 48093 3050 48094 3114
rect 48028 2960 48094 3050
rect 48154 2896 48214 3926
rect 48274 2956 48334 3988
rect 48394 2896 48454 3926
rect 48514 2956 48574 3988
rect 48634 3834 48700 3988
rect 48634 3770 48635 3834
rect 48699 3770 48700 3834
rect 48634 3754 48700 3770
rect 48634 3690 48635 3754
rect 48699 3690 48700 3754
rect 48634 3674 48700 3690
rect 48634 3610 48635 3674
rect 48699 3610 48700 3674
rect 48634 3594 48700 3610
rect 48634 3530 48635 3594
rect 48699 3530 48700 3594
rect 48634 3514 48700 3530
rect 48634 3450 48635 3514
rect 48699 3450 48700 3514
rect 48634 3434 48700 3450
rect 48634 3370 48635 3434
rect 48699 3370 48700 3434
rect 48634 3354 48700 3370
rect 48634 3290 48635 3354
rect 48699 3290 48700 3354
rect 48634 3274 48700 3290
rect 48634 3210 48635 3274
rect 48699 3210 48700 3274
rect 48634 3194 48700 3210
rect 48634 3130 48635 3194
rect 48699 3130 48700 3194
rect 48634 3114 48700 3130
rect 48634 3050 48635 3114
rect 48699 3050 48700 3114
rect 48634 2960 48700 3050
rect 48760 2896 48820 3926
rect 48880 2956 48940 3988
rect 49000 2896 49060 3926
rect 49120 2956 49180 3988
rect 49240 3834 49306 3988
rect 49240 3770 49241 3834
rect 49305 3770 49306 3834
rect 49240 3754 49306 3770
rect 49240 3690 49241 3754
rect 49305 3690 49306 3754
rect 49240 3674 49306 3690
rect 49240 3610 49241 3674
rect 49305 3610 49306 3674
rect 49240 3594 49306 3610
rect 49240 3530 49241 3594
rect 49305 3530 49306 3594
rect 49240 3514 49306 3530
rect 49240 3450 49241 3514
rect 49305 3450 49306 3514
rect 49240 3434 49306 3450
rect 49240 3370 49241 3434
rect 49305 3370 49306 3434
rect 49240 3354 49306 3370
rect 49240 3290 49241 3354
rect 49305 3290 49306 3354
rect 49240 3274 49306 3290
rect 49240 3210 49241 3274
rect 49305 3210 49306 3274
rect 49240 3194 49306 3210
rect 49240 3130 49241 3194
rect 49305 3130 49306 3194
rect 49240 3114 49306 3130
rect 49240 3050 49241 3114
rect 49305 3050 49306 3114
rect 49240 2960 49306 3050
rect 49366 2896 49426 3926
rect 49486 2956 49546 3988
rect 49606 2896 49666 3926
rect 49726 2956 49786 3988
rect 49846 3834 49912 3988
rect 49846 3770 49847 3834
rect 49911 3770 49912 3834
rect 49846 3754 49912 3770
rect 49846 3690 49847 3754
rect 49911 3690 49912 3754
rect 49846 3674 49912 3690
rect 49846 3610 49847 3674
rect 49911 3610 49912 3674
rect 49846 3594 49912 3610
rect 49846 3530 49847 3594
rect 49911 3530 49912 3594
rect 49846 3514 49912 3530
rect 49846 3450 49847 3514
rect 49911 3450 49912 3514
rect 49846 3434 49912 3450
rect 49846 3370 49847 3434
rect 49911 3370 49912 3434
rect 49846 3354 49912 3370
rect 49846 3290 49847 3354
rect 49911 3290 49912 3354
rect 49846 3274 49912 3290
rect 49846 3210 49847 3274
rect 49911 3210 49912 3274
rect 49846 3194 49912 3210
rect 49846 3130 49847 3194
rect 49911 3130 49912 3194
rect 49846 3114 49912 3130
rect 49846 3050 49847 3114
rect 49911 3050 49912 3114
rect 49846 2960 49912 3050
rect 49972 2896 50032 3926
rect 50092 2956 50152 3988
rect 50212 2896 50272 3926
rect 50332 2956 50392 3988
rect 50452 3834 50518 3988
rect 50452 3770 50453 3834
rect 50517 3770 50518 3834
rect 50452 3754 50518 3770
rect 50452 3690 50453 3754
rect 50517 3690 50518 3754
rect 50452 3674 50518 3690
rect 50452 3610 50453 3674
rect 50517 3610 50518 3674
rect 50452 3594 50518 3610
rect 50452 3530 50453 3594
rect 50517 3530 50518 3594
rect 50452 3514 50518 3530
rect 50452 3450 50453 3514
rect 50517 3450 50518 3514
rect 50452 3434 50518 3450
rect 50452 3370 50453 3434
rect 50517 3370 50518 3434
rect 50452 3354 50518 3370
rect 50452 3290 50453 3354
rect 50517 3290 50518 3354
rect 50452 3274 50518 3290
rect 50452 3210 50453 3274
rect 50517 3210 50518 3274
rect 50452 3194 50518 3210
rect 50452 3130 50453 3194
rect 50517 3130 50518 3194
rect 50452 3114 50518 3130
rect 50452 3050 50453 3114
rect 50517 3050 50518 3114
rect 50452 2960 50518 3050
rect 50578 2896 50638 3926
rect 50698 2956 50758 3988
rect 50818 2896 50878 3926
rect 50938 2956 50998 3988
rect 51058 3834 51124 3988
rect 51058 3770 51059 3834
rect 51123 3770 51124 3834
rect 51058 3754 51124 3770
rect 51058 3690 51059 3754
rect 51123 3690 51124 3754
rect 51058 3674 51124 3690
rect 51058 3610 51059 3674
rect 51123 3610 51124 3674
rect 51058 3594 51124 3610
rect 51058 3530 51059 3594
rect 51123 3530 51124 3594
rect 51058 3514 51124 3530
rect 51058 3450 51059 3514
rect 51123 3450 51124 3514
rect 51058 3434 51124 3450
rect 51058 3370 51059 3434
rect 51123 3370 51124 3434
rect 51058 3354 51124 3370
rect 51058 3290 51059 3354
rect 51123 3290 51124 3354
rect 51058 3274 51124 3290
rect 51058 3210 51059 3274
rect 51123 3210 51124 3274
rect 51058 3194 51124 3210
rect 51058 3130 51059 3194
rect 51123 3130 51124 3194
rect 51058 3114 51124 3130
rect 51058 3050 51059 3114
rect 51123 3050 51124 3114
rect 51058 2960 51124 3050
rect 51184 2896 51244 3926
rect 51304 2956 51364 3988
rect 51424 2896 51484 3926
rect 51544 2956 51604 3988
rect 51664 3834 51730 3988
rect 51664 3770 51665 3834
rect 51729 3770 51730 3834
rect 51664 3754 51730 3770
rect 51664 3690 51665 3754
rect 51729 3690 51730 3754
rect 51664 3674 51730 3690
rect 51664 3610 51665 3674
rect 51729 3610 51730 3674
rect 51664 3594 51730 3610
rect 51664 3530 51665 3594
rect 51729 3530 51730 3594
rect 51664 3514 51730 3530
rect 51664 3450 51665 3514
rect 51729 3450 51730 3514
rect 51664 3434 51730 3450
rect 51664 3370 51665 3434
rect 51729 3370 51730 3434
rect 51664 3354 51730 3370
rect 51664 3290 51665 3354
rect 51729 3290 51730 3354
rect 51664 3274 51730 3290
rect 51664 3210 51665 3274
rect 51729 3210 51730 3274
rect 51664 3194 51730 3210
rect 51664 3130 51665 3194
rect 51729 3130 51730 3194
rect 51664 3114 51730 3130
rect 51664 3050 51665 3114
rect 51729 3050 51730 3114
rect 51664 2960 51730 3050
rect 32272 2894 51730 2896
rect 32272 2830 32376 2894
rect 32440 2830 32456 2894
rect 32520 2830 32536 2894
rect 32600 2830 32616 2894
rect 32680 2830 32696 2894
rect 32760 2830 32776 2894
rect 32840 2830 32982 2894
rect 33046 2830 33062 2894
rect 33126 2830 33142 2894
rect 33206 2830 33222 2894
rect 33286 2830 33302 2894
rect 33366 2830 33382 2894
rect 33446 2830 33588 2894
rect 33652 2830 33668 2894
rect 33732 2830 33748 2894
rect 33812 2830 33828 2894
rect 33892 2830 33908 2894
rect 33972 2830 33988 2894
rect 34052 2830 34194 2894
rect 34258 2830 34274 2894
rect 34338 2830 34354 2894
rect 34418 2830 34434 2894
rect 34498 2830 34514 2894
rect 34578 2830 34594 2894
rect 34658 2830 34800 2894
rect 34864 2830 34880 2894
rect 34944 2830 34960 2894
rect 35024 2830 35040 2894
rect 35104 2830 35120 2894
rect 35184 2830 35200 2894
rect 35264 2830 35406 2894
rect 35470 2830 35486 2894
rect 35550 2830 35566 2894
rect 35630 2830 35646 2894
rect 35710 2830 35726 2894
rect 35790 2830 35806 2894
rect 35870 2830 36012 2894
rect 36076 2830 36092 2894
rect 36156 2830 36172 2894
rect 36236 2830 36252 2894
rect 36316 2830 36332 2894
rect 36396 2830 36412 2894
rect 36476 2830 36618 2894
rect 36682 2830 36698 2894
rect 36762 2830 36778 2894
rect 36842 2830 36858 2894
rect 36922 2830 36938 2894
rect 37002 2830 37018 2894
rect 37082 2830 37224 2894
rect 37288 2830 37304 2894
rect 37368 2830 37384 2894
rect 37448 2830 37464 2894
rect 37528 2830 37544 2894
rect 37608 2830 37624 2894
rect 37688 2830 37830 2894
rect 37894 2830 37910 2894
rect 37974 2830 37990 2894
rect 38054 2830 38070 2894
rect 38134 2830 38150 2894
rect 38214 2830 38230 2894
rect 38294 2830 38436 2894
rect 38500 2830 38516 2894
rect 38580 2830 38596 2894
rect 38660 2830 38676 2894
rect 38740 2830 38756 2894
rect 38820 2830 38836 2894
rect 38900 2830 39042 2894
rect 39106 2830 39122 2894
rect 39186 2830 39202 2894
rect 39266 2830 39282 2894
rect 39346 2830 39362 2894
rect 39426 2830 39442 2894
rect 39506 2830 39648 2894
rect 39712 2830 39728 2894
rect 39792 2830 39808 2894
rect 39872 2830 39888 2894
rect 39952 2830 39968 2894
rect 40032 2830 40048 2894
rect 40112 2830 40254 2894
rect 40318 2830 40334 2894
rect 40398 2830 40414 2894
rect 40478 2830 40494 2894
rect 40558 2830 40574 2894
rect 40638 2830 40654 2894
rect 40718 2830 40860 2894
rect 40924 2830 40940 2894
rect 41004 2830 41020 2894
rect 41084 2830 41100 2894
rect 41164 2830 41180 2894
rect 41244 2830 41260 2894
rect 41324 2830 41466 2894
rect 41530 2830 41546 2894
rect 41610 2830 41626 2894
rect 41690 2830 41706 2894
rect 41770 2830 41786 2894
rect 41850 2830 41866 2894
rect 41930 2830 42072 2894
rect 42136 2830 42152 2894
rect 42216 2830 42232 2894
rect 42296 2830 42312 2894
rect 42376 2830 42392 2894
rect 42456 2830 42472 2894
rect 42536 2830 42678 2894
rect 42742 2830 42758 2894
rect 42822 2830 42838 2894
rect 42902 2830 42918 2894
rect 42982 2830 42998 2894
rect 43062 2830 43078 2894
rect 43142 2830 43284 2894
rect 43348 2830 43364 2894
rect 43428 2830 43444 2894
rect 43508 2830 43524 2894
rect 43588 2830 43604 2894
rect 43668 2830 43684 2894
rect 43748 2830 43890 2894
rect 43954 2830 43970 2894
rect 44034 2830 44050 2894
rect 44114 2830 44130 2894
rect 44194 2830 44210 2894
rect 44274 2830 44290 2894
rect 44354 2830 44496 2894
rect 44560 2830 44576 2894
rect 44640 2830 44656 2894
rect 44720 2830 44736 2894
rect 44800 2830 44816 2894
rect 44880 2830 44896 2894
rect 44960 2830 45102 2894
rect 45166 2830 45182 2894
rect 45246 2830 45262 2894
rect 45326 2830 45342 2894
rect 45406 2830 45422 2894
rect 45486 2830 45502 2894
rect 45566 2830 45708 2894
rect 45772 2830 45788 2894
rect 45852 2830 45868 2894
rect 45932 2830 45948 2894
rect 46012 2830 46028 2894
rect 46092 2830 46108 2894
rect 46172 2830 46314 2894
rect 46378 2830 46394 2894
rect 46458 2830 46474 2894
rect 46538 2830 46554 2894
rect 46618 2830 46634 2894
rect 46698 2830 46714 2894
rect 46778 2830 46920 2894
rect 46984 2830 47000 2894
rect 47064 2830 47080 2894
rect 47144 2830 47160 2894
rect 47224 2830 47240 2894
rect 47304 2830 47320 2894
rect 47384 2830 47526 2894
rect 47590 2830 47606 2894
rect 47670 2830 47686 2894
rect 47750 2830 47766 2894
rect 47830 2830 47846 2894
rect 47910 2830 47926 2894
rect 47990 2830 48132 2894
rect 48196 2830 48212 2894
rect 48276 2830 48292 2894
rect 48356 2830 48372 2894
rect 48436 2830 48452 2894
rect 48516 2830 48532 2894
rect 48596 2830 48738 2894
rect 48802 2830 48818 2894
rect 48882 2830 48898 2894
rect 48962 2830 48978 2894
rect 49042 2830 49058 2894
rect 49122 2830 49138 2894
rect 49202 2830 49344 2894
rect 49408 2830 49424 2894
rect 49488 2830 49504 2894
rect 49568 2830 49584 2894
rect 49648 2830 49664 2894
rect 49728 2830 49744 2894
rect 49808 2830 49950 2894
rect 50014 2830 50030 2894
rect 50094 2830 50110 2894
rect 50174 2830 50190 2894
rect 50254 2830 50270 2894
rect 50334 2830 50350 2894
rect 50414 2830 50556 2894
rect 50620 2830 50636 2894
rect 50700 2830 50716 2894
rect 50780 2830 50796 2894
rect 50860 2830 50876 2894
rect 50940 2830 50956 2894
rect 51020 2830 51162 2894
rect 51226 2830 51242 2894
rect 51306 2830 51322 2894
rect 51386 2830 51402 2894
rect 51466 2830 51482 2894
rect 51546 2830 51562 2894
rect 51626 2830 51730 2894
rect 32272 2828 51730 2830
<< labels >>
flabel pwell 32592 4404 32618 4436 0 FreeSans 160 0 0 0 x1[1].SUB
flabel metal4 32534 4738 32560 4770 0 FreeSans 320 0 0 0 x1[1].CBOT
flabel metal4 32652 4148 32678 4180 0 FreeSans 320 0 0 0 x1[1].CTOP
flabel pwell 32592 3244 32618 3276 0 FreeSans 160 0 0 0 x1[0].SUB
flabel metal4 32534 3578 32560 3610 0 FreeSans 320 0 0 0 x1[0].CBOT
flabel metal4 32652 2988 32678 3020 0 FreeSans 320 0 0 0 x1[0].CTOP
flabel pwell 33804 3244 33830 3276 0 FreeSans 160 0 0 0 x1[4].SUB
flabel metal4 33746 3578 33772 3610 0 FreeSans 320 0 0 0 x1[4].CBOT
flabel metal4 33864 2988 33890 3020 0 FreeSans 320 0 0 0 x1[4].CTOP
flabel pwell 33198 3244 33224 3276 0 FreeSans 160 0 0 0 x1[2].SUB
flabel metal4 33140 3578 33166 3610 0 FreeSans 320 0 0 0 x1[2].CBOT
flabel metal4 33258 2988 33284 3020 0 FreeSans 320 0 0 0 x1[2].CTOP
flabel pwell 34410 3244 34436 3276 0 FreeSans 160 0 0 0 x1[6].SUB
flabel metal4 34352 3578 34378 3610 0 FreeSans 320 0 0 0 x1[6].CBOT
flabel metal4 34470 2988 34496 3020 0 FreeSans 320 0 0 0 x1[6].CTOP
flabel pwell 35016 3244 35042 3276 0 FreeSans 160 0 0 0 x1[8].SUB
flabel metal4 34958 3578 34984 3610 0 FreeSans 320 0 0 0 x1[8].CBOT
flabel metal4 35076 2988 35102 3020 0 FreeSans 320 0 0 0 x1[8].CTOP
flabel pwell 35622 3244 35648 3276 0 FreeSans 160 0 0 0 x1[10].SUB
flabel metal4 35564 3578 35590 3610 0 FreeSans 320 0 0 0 x1[10].CBOT
flabel metal4 35682 2988 35708 3020 0 FreeSans 320 0 0 0 x1[10].CTOP
flabel pwell 36228 3244 36254 3276 0 FreeSans 160 0 0 0 x1[12].SUB
flabel metal4 36170 3578 36196 3610 0 FreeSans 320 0 0 0 x1[12].CBOT
flabel metal4 36288 2988 36314 3020 0 FreeSans 320 0 0 0 x1[12].CTOP
flabel pwell 33804 4404 33830 4436 0 FreeSans 160 0 0 0 x1[5].SUB
flabel metal4 33746 4738 33772 4770 0 FreeSans 320 0 0 0 x1[5].CBOT
flabel metal4 33864 4148 33890 4180 0 FreeSans 320 0 0 0 x1[5].CTOP
flabel pwell 33198 4404 33224 4436 0 FreeSans 160 0 0 0 x1[3].SUB
flabel metal4 33140 4738 33166 4770 0 FreeSans 320 0 0 0 x1[3].CBOT
flabel metal4 33258 4148 33284 4180 0 FreeSans 320 0 0 0 x1[3].CTOP
flabel pwell 34410 4404 34436 4436 0 FreeSans 160 0 0 0 x1[7].SUB
flabel metal4 34352 4738 34378 4770 0 FreeSans 320 0 0 0 x1[7].CBOT
flabel metal4 34470 4148 34496 4180 0 FreeSans 320 0 0 0 x1[7].CTOP
flabel pwell 35016 4404 35042 4436 0 FreeSans 160 0 0 0 x1[9].SUB
flabel metal4 34958 4738 34984 4770 0 FreeSans 320 0 0 0 x1[9].CBOT
flabel metal4 35076 4148 35102 4180 0 FreeSans 320 0 0 0 x1[9].CTOP
flabel pwell 35622 4404 35648 4436 0 FreeSans 160 0 0 0 x1[11].SUB
flabel metal4 35564 4738 35590 4770 0 FreeSans 320 0 0 0 x1[11].CBOT
flabel metal4 35682 4148 35708 4180 0 FreeSans 320 0 0 0 x1[11].CTOP
flabel pwell 36228 4404 36254 4436 0 FreeSans 160 0 0 0 x1[13].SUB
flabel metal4 36170 4738 36196 4770 0 FreeSans 320 0 0 0 x1[13].CBOT
flabel metal4 36288 4148 36314 4180 0 FreeSans 320 0 0 0 x1[13].CTOP
flabel pwell 37440 3244 37466 3276 0 FreeSans 160 0 0 0 x1[16].SUB
flabel metal4 37382 3578 37408 3610 0 FreeSans 320 0 0 0 x1[16].CBOT
flabel metal4 37500 2988 37526 3020 0 FreeSans 320 0 0 0 x1[16].CTOP
flabel pwell 36834 3244 36860 3276 0 FreeSans 160 0 0 0 x1[14].SUB
flabel metal4 36776 3578 36802 3610 0 FreeSans 320 0 0 0 x1[14].CBOT
flabel metal4 36894 2988 36920 3020 0 FreeSans 320 0 0 0 x1[14].CTOP
flabel pwell 38046 3244 38072 3276 0 FreeSans 160 0 0 0 x1[18].SUB
flabel metal4 37988 3578 38014 3610 0 FreeSans 320 0 0 0 x1[18].CBOT
flabel metal4 38106 2988 38132 3020 0 FreeSans 320 0 0 0 x1[18].CTOP
flabel pwell 38652 3244 38678 3276 0 FreeSans 160 0 0 0 x1[20].SUB
flabel metal4 38594 3578 38620 3610 0 FreeSans 320 0 0 0 x1[20].CBOT
flabel metal4 38712 2988 38738 3020 0 FreeSans 320 0 0 0 x1[20].CTOP
flabel pwell 39258 3244 39284 3276 0 FreeSans 160 0 0 0 x1[22].SUB
flabel metal4 39200 3578 39226 3610 0 FreeSans 320 0 0 0 x1[22].CBOT
flabel metal4 39318 2988 39344 3020 0 FreeSans 320 0 0 0 x1[22].CTOP
flabel pwell 39864 3244 39890 3276 0 FreeSans 160 0 0 0 x1[24].SUB
flabel metal4 39806 3578 39832 3610 0 FreeSans 320 0 0 0 x1[24].CBOT
flabel metal4 39924 2988 39950 3020 0 FreeSans 320 0 0 0 x1[24].CTOP
flabel pwell 37440 4404 37466 4436 0 FreeSans 160 0 0 0 x1[17].SUB
flabel metal4 37382 4738 37408 4770 0 FreeSans 320 0 0 0 x1[17].CBOT
flabel metal4 37500 4148 37526 4180 0 FreeSans 320 0 0 0 x1[17].CTOP
flabel pwell 36834 4404 36860 4436 0 FreeSans 160 0 0 0 x1[15].SUB
flabel metal4 36776 4738 36802 4770 0 FreeSans 320 0 0 0 x1[15].CBOT
flabel metal4 36894 4148 36920 4180 0 FreeSans 320 0 0 0 x1[15].CTOP
flabel pwell 38046 4404 38072 4436 0 FreeSans 160 0 0 0 x1[19].SUB
flabel metal4 37988 4738 38014 4770 0 FreeSans 320 0 0 0 x1[19].CBOT
flabel metal4 38106 4148 38132 4180 0 FreeSans 320 0 0 0 x1[19].CTOP
flabel pwell 38652 4404 38678 4436 0 FreeSans 160 0 0 0 x1[21].SUB
flabel metal4 38594 4738 38620 4770 0 FreeSans 320 0 0 0 x1[21].CBOT
flabel metal4 38712 4148 38738 4180 0 FreeSans 320 0 0 0 x1[21].CTOP
flabel pwell 39258 4404 39284 4436 0 FreeSans 160 0 0 0 x1[23].SUB
flabel metal4 39200 4738 39226 4770 0 FreeSans 320 0 0 0 x1[23].CBOT
flabel metal4 39318 4148 39344 4180 0 FreeSans 320 0 0 0 x1[23].CTOP
flabel pwell 39864 4404 39890 4436 0 FreeSans 160 0 0 0 x1[25].SUB
flabel metal4 39806 4738 39832 4770 0 FreeSans 320 0 0 0 x1[25].CBOT
flabel metal4 39924 4148 39950 4180 0 FreeSans 320 0 0 0 x1[25].CTOP
flabel pwell 41682 3244 41708 3276 0 FreeSans 160 0 0 0 x1[30].SUB
flabel metal4 41624 3578 41650 3610 0 FreeSans 320 0 0 0 x1[30].CBOT
flabel metal4 41742 2988 41768 3020 0 FreeSans 320 0 0 0 x1[30].CTOP
flabel pwell 40470 3244 40496 3276 0 FreeSans 160 0 0 0 x1[26].SUB
flabel metal4 40412 3578 40438 3610 0 FreeSans 320 0 0 0 x1[26].CBOT
flabel metal4 40530 2988 40556 3020 0 FreeSans 320 0 0 0 x1[26].CTOP
flabel pwell 41076 3244 41102 3276 0 FreeSans 160 0 0 0 x1[28].SUB
flabel metal4 41018 3578 41044 3610 0 FreeSans 320 0 0 0 x1[28].CBOT
flabel metal4 41136 2988 41162 3020 0 FreeSans 320 0 0 0 x1[28].CTOP
flabel pwell 44106 3244 44132 3276 0 FreeSans 160 0 0 0 x1[38].SUB
flabel metal4 44048 3578 44074 3610 0 FreeSans 320 0 0 0 x1[38].CBOT
flabel metal4 44166 2988 44192 3020 0 FreeSans 320 0 0 0 x1[38].CTOP
flabel pwell 43500 3244 43526 3276 0 FreeSans 160 0 0 0 x1[36].SUB
flabel metal4 43442 3578 43468 3610 0 FreeSans 320 0 0 0 x1[36].CBOT
flabel metal4 43560 2988 43586 3020 0 FreeSans 320 0 0 0 x1[36].CTOP
flabel pwell 42894 3244 42920 3276 0 FreeSans 160 0 0 0 x1[34].SUB
flabel metal4 42836 3578 42862 3610 0 FreeSans 320 0 0 0 x1[34].CBOT
flabel metal4 42954 2988 42980 3020 0 FreeSans 320 0 0 0 x1[34].CTOP
flabel pwell 42288 3244 42314 3276 0 FreeSans 160 0 0 0 x1[32].SUB
flabel metal4 42230 3578 42256 3610 0 FreeSans 320 0 0 0 x1[32].CBOT
flabel metal4 42348 2988 42374 3020 0 FreeSans 320 0 0 0 x1[32].CTOP
flabel pwell 41682 4404 41708 4436 0 FreeSans 160 0 0 0 x1[31].SUB
flabel metal4 41624 4738 41650 4770 0 FreeSans 320 0 0 0 x1[31].CBOT
flabel metal4 41742 4148 41768 4180 0 FreeSans 320 0 0 0 x1[31].CTOP
flabel pwell 40470 4404 40496 4436 0 FreeSans 160 0 0 0 x1[27].SUB
flabel metal4 40412 4738 40438 4770 0 FreeSans 320 0 0 0 x1[27].CBOT
flabel metal4 40530 4148 40556 4180 0 FreeSans 320 0 0 0 x1[27].CTOP
flabel pwell 41076 4404 41102 4436 0 FreeSans 160 0 0 0 x1[29].SUB
flabel metal4 41018 4738 41044 4770 0 FreeSans 320 0 0 0 x1[29].CBOT
flabel metal4 41136 4148 41162 4180 0 FreeSans 320 0 0 0 x1[29].CTOP
flabel pwell 44106 4404 44132 4436 0 FreeSans 160 0 0 0 x1[39].SUB
flabel metal4 44048 4738 44074 4770 0 FreeSans 320 0 0 0 x1[39].CBOT
flabel metal4 44166 4148 44192 4180 0 FreeSans 320 0 0 0 x1[39].CTOP
flabel pwell 43500 4404 43526 4436 0 FreeSans 160 0 0 0 x1[37].SUB
flabel metal4 43442 4738 43468 4770 0 FreeSans 320 0 0 0 x1[37].CBOT
flabel metal4 43560 4148 43586 4180 0 FreeSans 320 0 0 0 x1[37].CTOP
flabel pwell 42894 4404 42920 4436 0 FreeSans 160 0 0 0 x1[35].SUB
flabel metal4 42836 4738 42862 4770 0 FreeSans 320 0 0 0 x1[35].CBOT
flabel metal4 42954 4148 42980 4180 0 FreeSans 320 0 0 0 x1[35].CTOP
flabel pwell 42288 4404 42314 4436 0 FreeSans 160 0 0 0 x1[33].SUB
flabel metal4 42230 4738 42256 4770 0 FreeSans 320 0 0 0 x1[33].CBOT
flabel metal4 42348 4148 42374 4180 0 FreeSans 320 0 0 0 x1[33].CTOP
flabel pwell 45318 3244 45344 3276 0 FreeSans 160 0 0 0 x1[42].SUB
flabel metal4 45260 3578 45286 3610 0 FreeSans 320 0 0 0 x1[42].CBOT
flabel metal4 45378 2988 45404 3020 0 FreeSans 320 0 0 0 x1[42].CTOP
flabel pwell 44712 3244 44738 3276 0 FreeSans 160 0 0 0 x1[40].SUB
flabel metal4 44654 3578 44680 3610 0 FreeSans 320 0 0 0 x1[40].CBOT
flabel metal4 44772 2988 44798 3020 0 FreeSans 320 0 0 0 x1[40].CTOP
flabel pwell 46530 3244 46556 3276 0 FreeSans 160 0 0 0 x1[46].SUB
flabel metal4 46472 3578 46498 3610 0 FreeSans 320 0 0 0 x1[46].CBOT
flabel metal4 46590 2988 46616 3020 0 FreeSans 320 0 0 0 x1[46].CTOP
flabel pwell 45924 3244 45950 3276 0 FreeSans 160 0 0 0 x1[44].SUB
flabel metal4 45866 3578 45892 3610 0 FreeSans 320 0 0 0 x1[44].CBOT
flabel metal4 45984 2988 46010 3020 0 FreeSans 320 0 0 0 x1[44].CTOP
flabel pwell 47742 3244 47768 3276 0 FreeSans 160 0 0 0 x1[50].SUB
flabel metal4 47684 3578 47710 3610 0 FreeSans 320 0 0 0 x1[50].CBOT
flabel metal4 47802 2988 47828 3020 0 FreeSans 320 0 0 0 x1[50].CTOP
flabel pwell 47136 3244 47162 3276 0 FreeSans 160 0 0 0 x1[48].SUB
flabel metal4 47078 3578 47104 3610 0 FreeSans 320 0 0 0 x1[48].CBOT
flabel metal4 47196 2988 47222 3020 0 FreeSans 320 0 0 0 x1[48].CTOP
flabel pwell 45318 4404 45344 4436 0 FreeSans 160 0 0 0 x1[43].SUB
flabel metal4 45260 4738 45286 4770 0 FreeSans 320 0 0 0 x1[43].CBOT
flabel metal4 45378 4148 45404 4180 0 FreeSans 320 0 0 0 x1[43].CTOP
flabel pwell 44712 4404 44738 4436 0 FreeSans 160 0 0 0 x1[41].SUB
flabel metal4 44654 4738 44680 4770 0 FreeSans 320 0 0 0 x1[41].CBOT
flabel metal4 44772 4148 44798 4180 0 FreeSans 320 0 0 0 x1[41].CTOP
flabel pwell 46530 4404 46556 4436 0 FreeSans 160 0 0 0 x1[47].SUB
flabel metal4 46472 4738 46498 4770 0 FreeSans 320 0 0 0 x1[47].CBOT
flabel metal4 46590 4148 46616 4180 0 FreeSans 320 0 0 0 x1[47].CTOP
flabel pwell 45924 4404 45950 4436 0 FreeSans 160 0 0 0 x1[45].SUB
flabel metal4 45866 4738 45892 4770 0 FreeSans 320 0 0 0 x1[45].CBOT
flabel metal4 45984 4148 46010 4180 0 FreeSans 320 0 0 0 x1[45].CTOP
flabel pwell 47742 4404 47768 4436 0 FreeSans 160 0 0 0 x1[51].SUB
flabel metal4 47684 4738 47710 4770 0 FreeSans 320 0 0 0 x1[51].CBOT
flabel metal4 47802 4148 47828 4180 0 FreeSans 320 0 0 0 x1[51].CTOP
flabel pwell 47136 4404 47162 4436 0 FreeSans 160 0 0 0 x1[49].SUB
flabel metal4 47078 4738 47104 4770 0 FreeSans 320 0 0 0 x1[49].CBOT
flabel metal4 47196 4148 47222 4180 0 FreeSans 320 0 0 0 x1[49].CTOP
flabel pwell 48954 3244 48980 3276 0 FreeSans 160 0 0 0 x1[54].SUB
flabel metal4 48896 3578 48922 3610 0 FreeSans 320 0 0 0 x1[54].CBOT
flabel metal4 49014 2988 49040 3020 0 FreeSans 320 0 0 0 x1[54].CTOP
flabel pwell 48348 3244 48374 3276 0 FreeSans 160 0 0 0 x1[52].SUB
flabel metal4 48290 3578 48316 3610 0 FreeSans 320 0 0 0 x1[52].CBOT
flabel metal4 48408 2988 48434 3020 0 FreeSans 320 0 0 0 x1[52].CTOP
flabel pwell 50166 3244 50192 3276 0 FreeSans 160 0 0 0 x1[58].SUB
flabel metal4 50108 3578 50134 3610 0 FreeSans 320 0 0 0 x1[58].CBOT
flabel metal4 50226 2988 50252 3020 0 FreeSans 320 0 0 0 x1[58].CTOP
flabel pwell 49560 3244 49586 3276 0 FreeSans 160 0 0 0 x1[56].SUB
flabel metal4 49502 3578 49528 3610 0 FreeSans 320 0 0 0 x1[56].CBOT
flabel metal4 49620 2988 49646 3020 0 FreeSans 320 0 0 0 x1[56].CTOP
flabel pwell 51378 3244 51404 3276 0 FreeSans 160 0 0 0 x1[62].SUB
flabel metal4 51320 3578 51346 3610 0 FreeSans 320 0 0 0 x1[62].CBOT
flabel metal4 51438 2988 51464 3020 0 FreeSans 320 0 0 0 x1[62].CTOP
flabel pwell 50772 3244 50798 3276 0 FreeSans 160 0 0 0 x1[60].SUB
flabel metal4 50714 3578 50740 3610 0 FreeSans 320 0 0 0 x1[60].CBOT
flabel metal4 50832 2988 50858 3020 0 FreeSans 320 0 0 0 x1[60].CTOP
flabel pwell 48954 4404 48980 4436 0 FreeSans 160 0 0 0 x1[55].SUB
flabel metal4 48896 4738 48922 4770 0 FreeSans 320 0 0 0 x1[55].CBOT
flabel metal4 49014 4148 49040 4180 0 FreeSans 320 0 0 0 x1[55].CTOP
flabel pwell 48348 4404 48374 4436 0 FreeSans 160 0 0 0 x1[53].SUB
flabel metal4 48290 4738 48316 4770 0 FreeSans 320 0 0 0 x1[53].CBOT
flabel metal4 48408 4148 48434 4180 0 FreeSans 320 0 0 0 x1[53].CTOP
flabel pwell 50166 4404 50192 4436 0 FreeSans 160 0 0 0 x1[59].SUB
flabel metal4 50108 4738 50134 4770 0 FreeSans 320 0 0 0 x1[59].CBOT
flabel metal4 50226 4148 50252 4180 0 FreeSans 320 0 0 0 x1[59].CTOP
flabel pwell 49560 4404 49586 4436 0 FreeSans 160 0 0 0 x1[57].SUB
flabel metal4 49502 4738 49528 4770 0 FreeSans 320 0 0 0 x1[57].CBOT
flabel metal4 49620 4148 49646 4180 0 FreeSans 320 0 0 0 x1[57].CTOP
flabel pwell 51378 4404 51404 4436 0 FreeSans 160 0 0 0 x1[63].SUB
flabel metal4 51320 4738 51346 4770 0 FreeSans 320 0 0 0 x1[63].CBOT
flabel metal4 51438 4148 51464 4180 0 FreeSans 320 0 0 0 x1[63].CTOP
flabel pwell 50772 4404 50798 4436 0 FreeSans 160 0 0 0 x1[61].SUB
flabel metal4 50714 4738 50740 4770 0 FreeSans 320 0 0 0 x1[61].CBOT
flabel metal4 50832 4148 50858 4180 0 FreeSans 320 0 0 0 x1[61].CTOP
flabel pwell 42298 4090 42322 4112 0 FreeSans 160 0 0 0 SUB
port 2 nsew
<< end >>
