* NGSPICE file created from hgu_cdac_cap_32.ext - technology: sky130A

.subckt hgu_cdac_cap_32 SUB
C0 x1[9].CTOP x1[9].CBOT 80.7f
C1 x1[9].CTOP x1[8].CTOP 80.7f
.ends

