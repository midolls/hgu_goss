magic
tech sky130A
magscale 1 2
timestamp 1699773655
<< nwell >>
rect 5466 7675 5573 8047
rect 5361 6394 5624 7057
<< metal1 >>
rect 192 13707 198 13759
rect 250 13757 256 13759
rect 250 13710 311 13757
rect 250 13707 256 13710
rect 2400 9250 2406 9302
rect 2458 9250 2464 9302
rect 2700 9026 7880 9056
rect 2700 8957 7880 8987
rect 2700 8887 7880 8917
rect 2700 8817 7880 8847
rect 2700 8748 7880 8778
rect 2700 8678 7880 8708
rect 2700 8608 7880 8638
rect 2700 8538 7880 8568
rect 2700 8469 7880 8499
rect 2700 8399 7880 8429
rect 2700 8330 7880 8360
rect 2700 8260 7880 8290
rect 2700 8190 7880 8220
rect 193 7870 199 7922
rect 251 7908 257 7922
rect 5424 7910 5600 8006
rect 251 7880 2788 7908
rect 251 7870 257 7880
rect 2760 5818 2788 7880
rect 5311 7270 5608 7462
rect 5315 6630 5612 6822
rect 5337 6086 5598 6182
rect 3361 5877 3367 5893
rect 3336 5842 3367 5877
rect 3361 5841 3367 5842
rect 3419 5877 3425 5893
rect 3419 5842 8922 5877
rect 3419 5841 3425 5842
rect 2747 5766 2753 5818
rect 2805 5766 2811 5818
rect 7444 5684 7450 5736
rect 7502 5725 7508 5736
rect 7630 5725 7636 5735
rect 7502 5695 7636 5725
rect 7502 5684 7508 5695
rect 7630 5683 7636 5695
rect 7688 5683 7694 5735
rect 7169 5615 7175 5667
rect 7227 5655 7233 5667
rect 7544 5655 7550 5665
rect 7227 5625 7550 5655
rect 7227 5615 7233 5625
rect 7544 5613 7550 5625
rect 7602 5613 7608 5665
rect 6894 5545 6900 5597
rect 6952 5585 6958 5597
rect 7457 5585 7463 5596
rect 6952 5555 7463 5585
rect 6952 5545 6958 5555
rect 7457 5544 7463 5555
rect 7515 5544 7521 5596
rect 6352 5475 6358 5527
rect 6410 5516 6416 5527
rect 7371 5516 7377 5526
rect 6410 5486 7377 5516
rect 6410 5475 6416 5486
rect 7371 5474 7377 5486
rect 7429 5474 7435 5526
rect 5787 5406 5793 5458
rect 5845 5446 5851 5458
rect 7284 5446 7290 5457
rect 5845 5416 7290 5446
rect 5845 5406 5851 5416
rect 7284 5405 7290 5416
rect 7342 5405 7348 5457
rect 5494 5336 5500 5388
rect 5552 5377 5558 5388
rect 7198 5377 7204 5387
rect 5552 5347 7204 5377
rect 5552 5336 5558 5347
rect 7198 5335 7204 5347
rect 7256 5335 7262 5387
rect 5408 5266 5414 5318
rect 5466 5307 5472 5318
rect 7112 5307 7118 5317
rect 5466 5277 7118 5307
rect 5466 5266 5472 5277
rect 7112 5265 7118 5277
rect 7170 5265 7176 5317
rect 5261 5196 5267 5248
rect 5319 5237 5325 5248
rect 7026 5237 7032 5247
rect 5319 5207 7032 5237
rect 5319 5196 5325 5207
rect 7026 5195 7032 5207
rect 7084 5195 7090 5247
rect 4988 5127 4994 5179
rect 5046 5167 5052 5179
rect 6939 5167 6945 5178
rect 5046 5137 6945 5167
rect 5046 5127 5052 5137
rect 6939 5126 6945 5137
rect 6997 5126 7003 5178
rect 4709 5057 4715 5109
rect 4767 5098 4773 5109
rect 6853 5098 6859 5108
rect 4767 5068 6859 5098
rect 4767 5057 4773 5068
rect 6853 5056 6859 5068
rect 6911 5056 6917 5108
rect 4162 4988 4168 5040
rect 4220 5028 4226 5040
rect 6767 5028 6773 5038
rect 4220 4998 6773 5028
rect 4220 4988 4226 4998
rect 6767 4986 6773 4998
rect 6825 4986 6831 5038
rect 3611 4918 3617 4970
rect 3669 4958 3675 4970
rect 6680 4958 6686 4969
rect 3669 4928 6686 4958
rect 3669 4918 3675 4928
rect 6680 4917 6686 4928
rect 6738 4917 6744 4969
rect 7406 66 7412 118
rect 7464 108 7470 118
rect 7464 78 23242 108
rect 7464 66 7470 78
rect 7954 -4 7960 48
rect 8012 38 8018 48
rect 8012 8 23242 38
rect 8012 -4 8018 8
rect 8221 -73 8227 -21
rect 8279 -32 8285 -21
rect 8279 -62 23242 -32
rect 8279 -73 8285 -62
rect 8507 -143 8513 -91
rect 8565 -101 8571 -91
rect 8565 -131 23242 -101
rect 8565 -143 8571 -131
rect 8734 -212 8740 -160
rect 8792 -171 8798 -160
rect 8792 -201 23242 -171
rect 8792 -212 8798 -201
rect 8820 -282 8826 -230
rect 8878 -240 8884 -230
rect 8878 -270 23242 -240
rect 8878 -282 8884 -270
rect 9206 -352 9212 -300
rect 9264 -310 9270 -300
rect 9264 -340 23242 -310
rect 9264 -352 9270 -340
rect 9752 -422 9758 -370
rect 9810 -380 9816 -370
rect 9810 -410 23242 -380
rect 9810 -422 9816 -410
rect 10299 -491 10305 -439
rect 10357 -450 10363 -439
rect 10357 -480 23242 -450
rect 10357 -491 10363 -480
rect 10585 -561 10591 -509
rect 10643 -519 10649 -509
rect 10643 -549 23242 -519
rect 10643 -561 10649 -549
rect 10851 -631 10857 -579
rect 10909 -589 10915 -579
rect 10909 -619 23242 -589
rect 10909 -631 10915 -619
rect 10998 -700 11004 -648
rect 11056 -659 11062 -648
rect 11056 -689 23242 -659
rect 11056 -700 11062 -689
rect 11085 -769 11091 -717
rect 11143 -728 11149 -717
rect 11143 -758 23242 -728
rect 11143 -769 11149 -758
rect 6349 -2874 11400 -2844
rect 6349 -2943 11400 -2913
rect 6349 -3013 11400 -2983
rect 6349 -3083 11400 -3053
rect 6349 -3152 11400 -3122
rect 6349 -3222 11400 -3192
rect 6349 -3292 11400 -3262
rect 6349 -3362 11400 -3332
rect 6349 -3431 11400 -3401
rect 6349 -3501 11400 -3471
rect 6349 -3570 11400 -3540
rect 6349 -3640 11400 -3610
rect 6349 -3710 11400 -3680
<< via1 >>
rect 198 13707 250 13759
rect 2406 9250 2458 9302
rect 199 7870 251 7922
rect 3367 5841 3419 5893
rect 2753 5766 2805 5818
rect 7450 5684 7502 5736
rect 7636 5683 7688 5735
rect 7175 5615 7227 5667
rect 7550 5613 7602 5665
rect 6900 5545 6952 5597
rect 7463 5544 7515 5596
rect 6358 5475 6410 5527
rect 7377 5474 7429 5526
rect 5793 5406 5845 5458
rect 7290 5405 7342 5457
rect 5500 5336 5552 5388
rect 7204 5335 7256 5387
rect 5414 5266 5466 5318
rect 7118 5265 7170 5317
rect 5267 5196 5319 5248
rect 7032 5195 7084 5247
rect 4994 5127 5046 5179
rect 6945 5126 6997 5178
rect 4715 5057 4767 5109
rect 6859 5056 6911 5108
rect 4168 4988 4220 5040
rect 6773 4986 6825 5038
rect 3617 4918 3669 4970
rect 6686 4917 6738 4969
rect 7412 66 7464 118
rect 7960 -4 8012 48
rect 8227 -73 8279 -21
rect 8513 -143 8565 -91
rect 8740 -212 8792 -160
rect 8826 -282 8878 -230
rect 9212 -352 9264 -300
rect 9758 -422 9810 -370
rect 10305 -491 10357 -439
rect 10591 -561 10643 -509
rect 10857 -631 10909 -579
rect 11004 -700 11056 -648
rect 11091 -769 11143 -717
<< metal2 >>
rect 192 13707 198 13759
rect 250 13707 256 13759
rect 206 7922 234 13707
rect 2400 9250 2406 9302
rect 2458 9250 2464 9302
rect 193 7870 199 7922
rect 251 7870 257 7922
rect 2420 7833 2448 9250
rect 3361 5841 3367 5893
rect 3419 5841 3425 5893
rect 2747 5766 2753 5818
rect 2805 5766 2811 5818
rect 3623 4970 3665 5750
rect 4172 5040 4214 5750
rect 4720 5109 4762 5750
rect 5000 5179 5042 5750
rect 5272 5248 5314 5750
rect 5419 5318 5461 5750
rect 5506 5388 5548 5750
rect 5799 5458 5841 5750
rect 6363 5527 6405 5750
rect 6906 5597 6948 5750
rect 7180 5667 7222 5750
rect 7455 5736 7497 5750
rect 7444 5684 7450 5736
rect 7502 5684 7508 5736
rect 7630 5683 7636 5735
rect 7688 5683 7694 5735
rect 7169 5615 7175 5667
rect 7227 5615 7233 5667
rect 7544 5613 7550 5665
rect 7602 5613 7608 5665
rect 6894 5545 6900 5597
rect 6952 5545 6958 5597
rect 7457 5544 7463 5596
rect 7515 5544 7521 5596
rect 6352 5475 6358 5527
rect 6410 5475 6416 5527
rect 7371 5474 7377 5526
rect 7429 5474 7435 5526
rect 5787 5406 5793 5458
rect 5845 5406 5851 5458
rect 7284 5405 7290 5457
rect 7342 5405 7348 5457
rect 5494 5336 5500 5388
rect 5552 5336 5558 5388
rect 7198 5335 7204 5387
rect 7256 5335 7262 5387
rect 5408 5266 5414 5318
rect 5466 5266 5472 5318
rect 7112 5265 7118 5317
rect 7170 5265 7176 5317
rect 5261 5196 5267 5248
rect 5319 5196 5325 5248
rect 7026 5195 7032 5247
rect 7084 5195 7090 5247
rect 4988 5127 4994 5179
rect 5046 5127 5052 5179
rect 6939 5126 6945 5178
rect 6997 5126 7003 5178
rect 4709 5057 4715 5109
rect 4767 5057 4773 5109
rect 6853 5056 6859 5108
rect 6911 5056 6917 5108
rect 4162 4988 4168 5040
rect 4220 4988 4226 5040
rect 6767 4986 6773 5038
rect 6825 4986 6831 5038
rect 3611 4918 3617 4970
rect 3669 4918 3675 4970
rect 6680 4917 6686 4969
rect 6738 4917 6744 4969
rect 6696 4809 6738 4917
rect 6778 4809 6820 4986
rect 6862 4809 6904 5056
rect 6950 4809 6992 5126
rect 7037 4809 7079 5195
rect 7123 4809 7165 5265
rect 7209 4809 7251 5335
rect 7296 4809 7338 5405
rect 7382 4809 7424 5474
rect 7468 4809 7510 5544
rect 7555 4809 7597 5613
rect 7640 4809 7682 5683
rect 7727 4810 7769 9120
rect 7814 4810 7856 9120
rect 7406 66 7412 118
rect 7464 66 7470 118
rect 7418 -813 7460 66
rect 7954 -4 7960 48
rect 8012 -4 8018 48
rect 7964 -813 8006 -4
rect 8221 -73 8227 -21
rect 8279 -73 8285 -21
rect 8232 -813 8274 -73
rect 8507 -143 8513 -91
rect 8565 -143 8571 -91
rect 8519 -813 8561 -143
rect 8734 -212 8740 -160
rect 8792 -212 8798 -160
rect 8745 -813 8787 -212
rect 8820 -282 8826 -230
rect 8878 -282 8884 -230
rect 8831 -813 8873 -282
rect 9206 -352 9212 -300
rect 9264 -352 9270 -300
rect 9218 -813 9260 -352
rect 9752 -422 9758 -370
rect 9810 -422 9816 -370
rect 9764 -813 9806 -422
rect 10299 -491 10305 -439
rect 10357 -491 10363 -439
rect 10310 -813 10352 -491
rect 10585 -561 10591 -509
rect 10643 -561 10649 -509
rect 10597 -813 10639 -561
rect 10851 -631 10857 -579
rect 10909 -631 10915 -579
rect 10862 -813 10904 -631
rect 10998 -700 11004 -648
rect 11056 -700 11062 -648
rect 11009 -813 11051 -700
rect 11085 -769 11091 -717
rect 11143 -769 11149 -717
rect 11096 -813 11138 -769
<< metal4 >>
rect 3412 9427 4376 9433
rect 3002 9248 4376 9427
rect 3002 9156 3190 9248
rect 3380 9246 4376 9248
rect 3380 9156 3584 9246
rect 3002 9154 3584 9156
rect 3774 9244 4376 9246
rect 3774 9154 3991 9244
rect 3002 9152 3991 9154
rect 4181 9152 4376 9244
rect 3002 7988 4376 9152
rect 5587 9236 6551 9395
rect 5587 9144 5716 9236
rect 5906 9232 6551 9236
rect 5906 9144 6142 9232
rect 5587 9140 6142 9144
rect 6332 9140 6551 9232
rect 3002 7982 3966 7988
rect 3002 6088 3414 7982
rect 5587 7951 6551 9140
rect 2614 4767 2896 5407
rect 4458 4767 5435 6192
rect 7587 6081 8059 8010
rect 2614 4473 6173 4767
rect 2614 4469 2896 4473
use hgu_cdac_sw_buffer  hgu_cdac_sw_buffer_0
timestamp 1699539897
transform -1 0 8443 0 -1 -3553
box -270 -2798 1830 -714
use hgu_cdac_sw_buffer  hgu_cdac_sw_buffer_1
timestamp 1699539897
transform -1 0 10797 0 -1 -3549
box -270 -2798 1830 -714
use hgu_cdac_sw_buffer  hgu_cdac_sw_buffer_2
timestamp 1699539897
transform -1 0 7382 0 1 8814
box -270 -2798 1830 -714
use hgu_cdac_sw_buffer  hgu_cdac_sw_buffer_3
timestamp 1699539897
transform -1 0 5204 0 1 8814
box -270 -2798 1830 -714
use hgu_comp_flat  hgu_comp_flat_0
timestamp 1698719859
transform 1 0 -324 0 1 7260
box 338 -1940 3788 618
use hgu_sarlogic_flat  hgu_sarlogic_flat_0
timestamp 1699766314
transform 1 0 -2020 0 1 1900
box 2064 -1908 31250 13749
use hgu_vgen_vref  hgu_vgen_vref_0
timestamp 1699773655
transform -1 0 -50750 0 1 -30367
box 0 -13 22370 76000
<< end >>
