* NGSPICE file created from hgu_sarlogic_retimer_flat.ext - technology: sky130A

.subckt hgu_sarlogic_retimer_RC VDD VSS sar_logic[0] sar_logic[1] sar_logic[2] sar_logic[3] sar_logic[4] sar_logic[5] sar_logic[6] sar_logic[7]
+ eob delay_code[0] delay_code[1] delay_code[2] delay_code[3] delay_offset
+ sar_retimer[0] sar_retimer[1] sar_retimer[2] sar_retimer[3] sar_retimer[4] sar_retimer[5] sar_retimer[6] sar_retimer[7]
X0 a_14018_6401# a_13844_6793# a_14158_6427# VSS.t214 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X1 sar_retimer[3].t1 a_17898_6427# VDD.t149 VDD.t148 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X2 a_16654_5787# a_16236_5787# a_16410_5761# VDD.t136 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X3 a_16410_7041# a_16236_7067# a_16550_7433# VSS.t184 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X4 VSS.t179 a_17191_5121# a_17126_5147# VSS.t178 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X5 a_13751_5147# sar_logic[6].t0 VSS.t48 VSS.t47 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X6 a_16922_6109# a_16410_5761# VSS.t63 VSS.t29 sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X7 VSS.t167 a_16410_5121# a_16344_5147# VSS.t166 sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X8 VSS.t107 eob.t0 a_12385_8002# VSS.t87 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X9 a_14530_7389# a_14018_7041# VSS.t163 VSS.t162 sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X10 sar_retimer[2].t1 a_15506_6427# VDD.t192 VDD.t49 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X11 a_14483_5787# a_14018_5761# VDD.t191 VDD.t23 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X12 a_16410_5761# VDD.t119 VDD.t120 VDD.t99 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X13 a_18195_9356# x2.x9.output_stack VDD.t174 VDD.t173 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X14 x3.X a_18499_9105# VDD.t189 VDD.t187 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X15 VDD.t171 a_16704_7267# a_16654_7067# VDD.t47 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X16 VDD.t169 a_17191_7041# a_17898_7083# VDD.t168 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X17 x2.x3[1].floating delay_code[1].t0 x2.x9.output_stack VSS.t215 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X18 VSS.t152 x3.X a_13397_7073# VSS.t151 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X19 x1[0].Q_N a_14799_7041# VDD.t161 VDD.t153 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X20 VDD.t118 VDD.t117 a_14312_6401# VDD.t96 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X21 a_16236_5787# a_15955_5793# a_16143_5787# VDD.t57 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X22 VDD.t186 x3.X a_13397_5147# VDD.t183 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X23 a_14262_7067# a_13844_7067# a_14018_7041# VDD.t34 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X24 a_16143_6427# sar_logic[3].t0 VDD.t197 VDD.t127 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X25 a_14734_7445# a_13397_7073# a_14625_7445# VSS.t126 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X26 a_14915_6153# a_14312_5987# a_14799_5761# VSS.t34 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X27 a_13928_5513# a_13397_5147# a_13844_5513# VDD.t140 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X28 VSS.t161 a_14018_7041# a_13952_7445# VSS.t160 sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X29 a_16236_7067# a_15789_7073# a_16143_7067# VSS.t221 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X30 VSS.t105 a_14799_5761# a_14734_6165# VSS.t104 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X31 a_13844_5787# a_13563_5793# a_13751_5787# VDD.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X32 VDD.t116 VDD.t115 a_16704_7267# VDD.t86 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X33 VDD.t229 a_17191_5761# a_17898_5803# VDD.t207 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X34 a_14018_7041# VDD.t113 VDD.t114 VDD.t89 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X35 a_13751_6427# sar_logic[2].t0 VDD.t131 VDD.t130 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X36 a_16654_6709# a_16236_6793# a_16410_6401# VDD.t213 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X37 VDD.t226 a_17191_6401# a_17103_6793# VDD.t166 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X38 VSS.t150 x3.X a_13397_5147# VSS.t149 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X39 a_14018_7041# a_13844_7067# a_14158_7433# VSS.t44 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X40 a_15033_7067# a_14625_7445# a_14799_7041# VDD.t147 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X41 VDD.t30 a_16410_6401# a_16320_6793# VDD.t29 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X42 VDD.t185 x3.X a_15789_5793# VDD.t175 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X43 a_16410_5761# a_16236_5787# a_16550_6153# VSS.t97 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X44 a_16875_5429# a_16410_5121# VDD.t196 VDD.t53 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X45 a_13844_7067# a_13397_7073# a_13751_7067# VSS.t125 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X46 VSS.t212 VDD.t239 a_16704_7267# VSS.t211 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X47 sar_retimer[1].t1 a_17898_7083# VDD.t163 VDD.t148 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X48 a_14483_6709# a_14018_6401# VDD.t125 VDD.t124 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X49 a_17103_5787# a_15955_5793# a_17017_6165# VDD.t56 sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X50 VDD.t170 a_16704_7267# a_17425_7067# VDD.t45 sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X51 a_14530_6109# a_14018_5761# VSS.t158 VSS.t77 sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X52 a_17307_6153# VDD.t240 VSS.t206 VSS.t197 sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X53 VSS.t28 a_14018_5121# a_13952_5147# VSS.t27 sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X54 a_16550_6427# VDD.t241 VSS.t207 VSS.t191 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X55 VDD.t160 a_14799_7041# a_15506_7083# VDD.t157 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X56 a_15955_7073# a_15789_7073# VDD.t219 VDD.t218 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X57 a_16922_5147# a_16410_5121# VSS.t165 VSS.t164 sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X58 VDD.t60 a_14312_5121# a_14262_5429# VDD.t40 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X59 sar_retimer[0].t1 a_15506_7083# VDD.t50 VDD.t49 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X60 a_17191_6401# a_17017_6427# a_17307_6427# VSS.t9 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X61 a_14711_5787# a_13563_5793# a_14625_6165# VDD.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X62 x2.x9.output_stack x2.x10.Y.t2 x2.x5[7].floating.t7 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X63 a_12385_8278# eob.t1 a_12297_8278# VSS.t72 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X64 a_14915_6153# VDD.t242 VSS.t208 VSS.t199 sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X65 VSS.t210 VDD.t243 a_16704_5121# VSS.t209 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X66 VDD.t112 VDD.t111 a_14312_5121# VDD.t77 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X67 VSS.t201 VDD.t244 a_14312_6401# VSS.t42 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X68 VSS.t231 a_17191_6401# a_17898_6427# VSS.t230 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X69 a_16143_5147# sar_logic[7].t0 VDD.t221 VDD.t21 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X70 a_17017_6165# a_15789_5793# a_16875_5787# VDD.t132 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X71 a_18195_9015# x2.x9.output_stack VSS.t138 VSS.t137 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X72 a_16320_6793# a_15789_6427# a_16236_6793# VDD.t217 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X73 VDD.t146 a_14799_5761# a_15506_5803# VDD.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X74 x1[7].Q_N a_17191_5121# VSS.t177 VSS.t176 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X75 VDD.t210 a_17191_5121# a_17103_5513# VDD.t209 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X76 a_14915_5147# a_14312_5121# a_14799_5121# VSS.t70 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X77 a_13751_5147# sar_logic[6].t1 VDD.t214 VDD.t150 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X78 a_17191_7041# VDD.t101 VDD.t102 VDD.t74 sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X79 VDD.t123 a_14018_6401# a_13928_6793# VDD.t122 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X80 x1[2].Q_N a_14799_6401# VSS.t116 VSS.t102 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X81 VDD.t184 x3.X a_13397_5793# VDD.t183 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X82 a_14018_5761# a_13844_5787# a_14158_6153# VSS.t214 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X83 VDD.t195 a_16410_5121# a_16320_5513# VDD.t51 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X84 a_16550_6427# a_16704_6401# a_16410_6401# VSS.t59 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X85 x2.x10.Y.t1 delay_code[3].t0 VDD.t231 VDD.t230 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X86 a_14158_6427# VDD.t245 VSS.t202 VSS.t85 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X87 a_16410_5121# a_16236_5513# a_16550_5147# VSS.t113 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X88 VDD.t59 a_14312_5121# a_15033_5429# VDD.t38 sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X89 a_17017_7445# a_15955_7073# a_16922_7389# VSS.t22 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X90 a_16344_5147# a_15955_5147# a_16236_5513# VSS.t66 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X91 a_18195_9356# x2.x9.output_stack x3.A VDD.t172 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.122 ps=1.42 w=0.42 l=0.15
X92 a_14625_7445# a_13397_7073# a_14483_7067# VDD.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X93 VDD.t159 a_14799_7041# a_14711_7067# VDD.t155 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X94 a_14530_5147# a_14018_5121# VSS.t26 VSS.t25 sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X95 a_12385_8692# eob.t2 a_12297_8554# VSS.t72 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X96 a_15955_7073# a_15789_7073# VSS.t220 VSS.t219 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X97 a_17191_7041# a_17017_7445# a_17307_7433# VSS.t76 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X98 a_14799_6401# a_14625_6427# a_14915_6427# VSS.t8 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X99 x1[6].Q_N a_14799_5121# VDD.t18 VDD.t17 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X100 a_13952_5147# a_13563_5147# a_13844_5513# VSS.t7 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X101 x1[1].Q_N a_17191_7041# VSS.t134 VSS.t133 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X102 VSS.t115 a_14799_6401# a_15506_6427# VSS.t100 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X103 a_14799_5761# VDD.t109 VDD.t110 VDD.t83 sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X104 sar_retimer[3].t0 a_17898_6427# VSS.t108 VSS.t45 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X105 VSS.t148 x3.X a_15789_5793# VSS.t145 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X106 a_16143_5787# sar_logic[5].t0 VSS.t52 VSS.t51 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X107 a_15955_5147# a_15789_5147# VDD.t135 VDD.t134 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X108 a_17425_5787# a_17017_6165# a_17191_5761# VDD.t55 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X109 x2.x9.output_stack x2.x10.Y.t3 x2.x5[7].floating.t6 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X110 x2.x9.output_stack delay_code[2].t0 x2.x4[3].floating VSS.t109 sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X111 a_14625_5147# a_13563_5147# a_14530_5147# VSS.t6 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X112 a_12385_8968# eob.t3 a_12297_8830# VSS.t72 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X113 a_12457_8140# eob.t4 a_12385_8278# VSS.t87 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X114 a_17126_7445# a_15789_7073# a_17017_7445# VSS.t218 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X115 a_13563_6427# a_13397_6427# VDD.t8 VDD.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X116 a_13751_5787# sar_logic[4].t0 VSS.t55 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X117 VSS.t234 a_17191_5761# a_17126_6165# VSS.t228 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X118 a_16320_5513# a_15789_5147# a_16236_5513# VDD.t133 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X119 x2.x9.output_stack delay_offset.t0 x2.x7.floating VSS.t12 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X120 a_18195_9015# x3.A VDD.t237 VSS.t240 sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X121 sar_retimer[2].t0 a_15506_6427# VSS.t159 VSS.t67 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X122 VDD.t26 a_14018_5121# a_13928_5513# VDD.t25 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X123 a_16410_6401# VDD.t107 VDD.t108 VDD.t80 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X124 VSS.t62 a_16410_5761# a_16344_6165# VSS.t31 sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X125 a_15955_5147# a_15789_5147# VSS.t96 VSS.t95 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X126 x3.X a_18499_9105# VSS.t156 VSS.t155 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X127 a_16550_7433# a_16704_7267# a_16410_7041# VSS.t136 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X128 VDD.t223 a_16704_5987# a_16654_5787# VDD.t203 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X129 x2.x9.output_stack x2.x10.Y.t4 x2.x5[7].floating.t5 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X130 a_13563_6427# a_13397_6427# VSS.t5 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X131 x1[4].Q_N a_14799_5761# VDD.t145 VDD.t17 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X132 sar_retimer[7].t1 a_17898_5147# VDD.t152 VDD.t35 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X133 a_14018_5121# a_13844_5513# a_14158_5147# VSS.t33 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X134 a_16236_6793# a_15955_6427# a_16143_6427# VDD.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X135 a_16875_7067# a_16410_7041# VDD.t212 VDD.t27 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X136 a_14262_5787# a_13844_5787# a_14018_5761# VDD.t31 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X137 a_13928_7067# a_13397_7073# a_13844_7067# VDD.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X138 sar_retimer[6].t1 a_15506_5147# VDD.t44 VDD.t43 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X139 a_17191_5761# a_17017_6165# a_17307_6153# VSS.t9 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X140 VDD.t233 delay_offset.t1 x2.x6.SW VDD.t232 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X141 a_14799_7041# a_14625_7445# a_14915_7433# VSS.t106 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X142 VDD.t143 eob.t5 a_12322_10357# VDD.t142 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X143 a_13844_6793# a_13563_6427# a_13751_6427# VDD.t199 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X144 a_17425_6709# a_17017_6427# a_17191_6401# VDD.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X145 VDD.t106 VDD.t105 a_16704_5987# VDD.t71 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X146 x1[5].Q_N a_17191_5761# VSS.t233 VSS.t226 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X147 VDD.t4 a_14312_7267# a_14262_7067# VDD.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X148 VSS.t147 x3.X a_13397_5793# VSS.t143 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X149 a_14018_5761# VDD.t103 VDD.t104 VDD.t68 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X150 x2.x9.output_stack delay_code[1].t1 x2.x3[1].floating VSS.t213 sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X151 a_14734_6427# a_13397_6427# a_14625_6427# VSS.t3 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X152 a_15033_5787# a_14625_6165# a_14799_5761# VDD.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X153 a_12457_8692# eob.t6 a_12385_8692# VSS.t87 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X154 a_16236_6793# a_15789_6427# a_16143_6427# VSS.t171 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X155 sar_retimer[5].t1 a_17898_5803# VDD.t36 VDD.t35 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X156 a_12410_9943# eob.t7 a_12322_9805# VDD.t42 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X157 VDD.t48 a_16704_6401# a_16654_6709# VDD.t47 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X158 a_17103_6793# a_15955_6427# a_17017_6427# VDD.t19 sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X159 a_14734_6165# a_13397_5793# a_14625_6165# VSS.t3 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X160 VDD.t222 a_16704_5987# a_17425_5787# VDD.t201 sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X161 a_16550_7433# VDD.t246 VSS.t204 VSS.t203 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X162 VSS.t114 a_14799_6401# a_14734_6427# VSS.t104 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X163 VSS.t157 a_14018_5761# a_13952_6165# VSS.t79 sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X164 a_16236_5787# a_15789_5793# a_16143_5787# VSS.t171 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X165 a_16410_5121# VDD.t98 VDD.t100 VDD.t99 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X166 a_13844_6793# a_13397_6427# a_13751_6427# VSS.t2 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X167 VDD.t225 a_17191_6401# a_17898_6427# VDD.t168 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X168 a_15955_5793# a_15789_5793# VDD.t200 VDD.t134 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X169 a_16550_6153# a_16704_5987# a_16410_5761# VSS.t59 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X170 a_16654_5429# a_16236_5513# a_16410_5121# VDD.t136 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X171 x2.x9.output_stack eob.t8 a_12385_8968# VSS.t87 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X172 a_14711_6793# a_13563_6427# a_14625_6427# VDD.t198 sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X173 sar_retimer[4].t1 a_15506_5803# VDD.t58 VDD.t43 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X174 VDD.t97 VDD.t95 a_14312_7267# VDD.t96 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X175 a_13844_5787# a_13397_5793# a_13751_5787# VSS.t2 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X176 VSS.t205 VDD.t247 a_16704_5987# VSS.t40 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X177 a_14262_6709# a_13844_6793# a_14018_6401# VDD.t34 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X178 a_16236_5513# a_15955_5147# a_16143_5147# VDD.t57 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X179 a_16143_7067# sar_logic[1].t0 VDD.t128 VDD.t127 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X180 VSS.t132 a_17191_7041# a_17898_7083# VSS.t131 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X181 a_14483_5429# a_14018_5121# VDD.t24 VDD.t23 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X182 VSS.t194 VDD.t248 a_14312_7267# VSS.t193 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X183 a_16550_5147# VDD.t249 VSS.t196 VSS.t195 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X184 a_12385_8554# eob.t9 a_12297_8554# VSS.t72 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X185 a_17307_6427# VDD.t250 VSS.t198 VSS.t197 sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X186 a_17307_6427# a_16704_6401# a_17191_6401# VSS.t58 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X187 a_14799_5761# a_14625_6165# a_14915_6153# VSS.t8 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X188 a_13844_5513# a_13563_5147# a_13751_5147# VDD.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X189 a_13751_7067# sar_logic[0].t0 VDD.t137 VDD.t130 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X190 VDD.t2 a_14312_7267# a_15033_7067# VDD.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X191 VDD.t167 a_17191_7041# a_17103_7067# VDD.t166 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X192 a_15033_6709# a_14625_6427# a_14799_6401# VDD.t147 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X193 a_17017_6427# a_15789_6427# a_16875_6709# VDD.t216 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X194 a_13563_7073# a_13397_7073# VDD.t162 VDD.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X195 a_17191_5121# a_17017_5147# a_17307_5147# VSS.t64 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X196 a_17191_5761# VDD.t93 VDD.t94 VDD.t65 sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X197 VDD.t211 a_16410_7041# a_16320_7067# VDD.t29 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X198 a_14915_6427# VDD.t251 VSS.t200 VSS.t199 sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X199 VSS.t175 a_17191_5121# a_17898_5147# VSS.t174 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X200 VDD.t46 a_16704_6401# a_17425_6709# VDD.t45 sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X201 a_17103_5513# a_15955_5147# a_17017_5147# VDD.t56 sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X202 VSS.t186 VDD.t252 a_14312_5121# VSS.t185 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X203 x2.x5[7].floating.t4 x2.x10.Y.t5 x2.x9.output_stack VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X204 VDD.t236 x3.A a_18499_9105# VDD.t235 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X205 VDD.t234 x3.A a_18195_9015# VSS.t239 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0651 ps=0.73 w=0.42 l=0.15
X206 a_14158_7433# VDD.t253 VSS.t188 VSS.t187 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X207 VSS.t238 x3.A a_18499_9105# VSS.t237 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X208 VDD.t158 a_14799_6401# a_15506_6427# VDD.t157 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X209 x2.x5[7].floating.t3 x2.x10.Y.t6 x2.x9.output_stack VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X210 x1[3].Q_N a_17191_6401# VDD.t224 VDD.t164 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X211 a_14625_6165# a_13397_5793# a_14483_5787# VDD.t141 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X212 x1[6].Q_N a_14799_5121# VSS.t20 VSS.t19 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X213 a_14711_5513# a_13563_5147# a_14625_5147# VDD.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X214 a_12410_9943# eob.t10 a_12322_10081# VDD.t121 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X215 a_16344_7445# a_15955_7073# a_16236_7067# VSS.t21 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X216 VDD.t144 a_14799_5761# a_14711_5787# VDD.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X217 a_16550_5147# a_16704_5121# a_16410_5121# VSS.t173 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X218 a_18195_9356# x3.A VSS.t236 VDD.t172 sky130_fd_pr__pfet_01v8_hvt ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X219 a_17017_6427# a_15955_6427# a_16922_6427# VSS.t75 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X220 VSS.t122 a_14799_7041# a_15506_7083# VSS.t121 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X221 a_14799_6401# VDD.t91 VDD.t92 VDD.t62 sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X222 a_14158_6427# a_14312_6401# a_14018_6401# VSS.t35 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X223 a_14158_5147# VDD.t254 VSS.t190 VSS.t189 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X224 a_12410_10219# eob.t11 a_12322_10357# VDD.t215 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X225 a_13952_7445# a_13563_7073# a_13844_7067# VSS.t217 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X226 a_16320_7067# a_15789_7073# a_16236_7067# VDD.t217 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X227 a_17307_7433# a_16704_7267# a_17191_7041# VSS.t135 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X228 a_17017_6165# a_15955_5793# a_16922_6109# VSS.t75 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X229 a_17017_5147# a_15789_5147# a_16875_5429# VDD.t132 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X230 VDD.t182 x3.X a_15789_6427# VDD.t179 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X231 x2.x5[7].floating.t2 x2.x10.Y.t7 x2.x9.output_stack VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X232 a_14625_7445# a_13563_7073# a_14530_7389# VSS.t216 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X233 VDD.t194 a_14018_7041# a_13928_7067# VDD.t122 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X234 a_15955_5793# a_15789_5793# VSS.t170 VSS.t169 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X235 a_14799_5121# a_14625_5147# a_14915_5147# VSS.t242 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X236 VDD.t188 a_18499_9105# x3.X VDD.t187 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X237 a_12457_8416# eob.t12 a_12385_8554# VSS.t87 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X238 a_17126_6427# a_15789_6427# a_17017_6427# VSS.t168 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X239 VSS.t18 a_14799_5121# a_15506_5147# VSS.t17 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X240 a_13563_7073# a_13397_7073# VSS.t124 VSS.t123 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X241 a_16143_6427# sar_logic[3].t1 VSS.t71 VSS.t51 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X242 sar_retimer[7].t0 a_17898_5147# VSS.t112 VSS.t111 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X243 x2.x9.output_stack eob.t13 a_12322_9805# VDD.t37 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X244 x1[0].Q_N a_14799_7041# VSS.t120 VSS.t119 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X245 VSS.t146 x3.X a_15789_6427# VSS.t145 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X246 a_17126_6165# a_15789_5793# a_17017_6165# VSS.t168 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X247 a_13563_5147# a_13397_5147# VDD.t220 VDD.t138 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X248 a_16875_5787# a_16410_5761# VDD.t54 VDD.t53 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X249 sar_retimer[6].t0 a_15506_5147# VSS.t57 VSS.t56 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X250 a_12385_8140# eob.t14 a_12297_8002# VSS.t72 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X251 a_13751_6427# sar_logic[2].t1 VSS.t11 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X252 VSS.t229 a_17191_6401# a_17126_6427# VSS.t228 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X253 a_13928_5787# a_13397_5793# a_13844_5787# VDD.t140 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X254 VSS.t32 a_16410_6401# a_16344_6427# VSS.t31 sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X255 x1[1].Q_N a_17191_7041# VDD.t165 VDD.t164 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X256 a_13563_5147# a_13397_5147# VSS.t225 VSS.t224 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X257 a_14018_6401# VDD.t88 VDD.t90 VDD.t89 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X258 VDD.t87 VDD.t85 a_16704_6401# VDD.t86 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X259 a_14799_5121# VDD.t82 VDD.t84 VDD.t83 sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X260 a_12385_8416# eob.t15 a_12297_8278# VSS.t72 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X261 a_14158_7433# a_14312_7267# a_14018_7041# VSS.t1 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X262 a_16654_7067# a_16236_7067# a_16410_7041# VDD.t213 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X263 VDD.t41 a_14312_5987# a_14262_5787# VDD.t40 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X264 a_17307_6153# a_16704_5987# a_17191_5761# VSS.t58 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X265 VDD.t181 x3.X a_13397_6427# VDD.t177 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X266 a_14483_7067# a_14018_7041# VDD.t193 VDD.t124 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X267 sar_retimer[1].t0 a_17898_7083# VSS.t128 VSS.t127 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X268 x2.x9.output_stack x2.x10.Y.t8 x2.x5[7].floating.t1 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X269 VSS.t118 a_14799_7041# a_14734_7445# VSS.t117 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X270 a_16410_7041# VDD.t79 VDD.t81 VDD.t80 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X271 a_17425_5429# a_17017_5147# a_17191_5121# VDD.t55 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X272 sar_retimer[0].t0 a_15506_7083# VSS.t61 VSS.t60 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X273 VSS.t144 x3.X a_13397_6427# VSS.t143 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X274 a_16875_6709# a_16410_6401# VDD.t28 VDD.t27 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X275 x1[4].Q_N a_14799_5761# VSS.t103 VSS.t102 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X276 VDD.t78 VDD.t76 a_14312_5987# VDD.t77 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X277 a_14734_5147# a_13397_5147# a_14625_5147# VSS.t223 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X278 x2.x10.Y.t0 delay_code[3].t1 VSS.t50 VSS.t49 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X279 a_16236_7067# a_15955_7073# a_16143_7067# VDD.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X280 a_16236_5513# a_15789_5147# a_16143_5147# VSS.t94 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X281 a_16143_5787# sar_logic[5].t1 VDD.t22 VDD.t21 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X282 x2.x2.floating delay_code[0].t0 x2.x9.output_stack VSS.t90 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.124 ps=1.43 w=0.42 l=0.15
X283 a_16550_6153# VDD.t255 VSS.t192 VSS.t191 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X284 VDD.t204 a_16704_5121# a_16654_5429# VDD.t203 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X285 VSS.t16 a_14799_5121# a_14734_5147# VSS.t15 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X286 a_13844_7067# a_13563_7073# a_13751_7067# VDD.t199 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X287 a_17307_7433# VDD.t256 VSS.t37 VSS.t36 sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X288 VSS.t80 a_14018_6401# a_13952_6427# VSS.t79 sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X289 VSS.t235 x3.A a_18195_9356# VDD.t172 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0651 ps=0.73 w=0.42 l=0.15
X290 VDD.t33 a_14312_6401# a_14262_6709# VDD.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X291 a_13751_5787# sar_logic[4].t1 VDD.t151 VDD.t150 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X292 VDD.t39 a_14312_5987# a_15033_5787# VDD.t38 sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X293 VDD.t208 a_17191_5121# a_17898_5147# VDD.t207 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X294 a_13844_5513# a_13397_5147# a_13751_5147# VSS.t222 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X295 VDD.t228 a_17191_5761# a_17103_5787# VDD.t209 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X296 a_17191_6401# VDD.t73 VDD.t75 VDD.t74 sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X297 a_16922_6427# a_16410_6401# VSS.t30 VSS.t29 sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X298 VDD.t72 VDD.t70 a_16704_5121# VDD.t71 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X299 a_14018_5121# VDD.t67 VDD.t69 VDD.t68 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X300 a_14915_7433# VDD.t257 VSS.t39 VSS.t38 sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X301 VDD.t180 x3.X a_15789_7073# VDD.t179 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X302 VSS.t41 VDD.t258 a_16704_6401# VSS.t40 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X303 a_13563_5793# a_13397_5793# VDD.t139 VDD.t138 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X304 a_14158_6153# a_14312_5987# a_14018_5761# VSS.t35 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X305 VDD.t52 a_16410_5761# a_16320_5787# VDD.t51 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X306 a_14262_5429# a_13844_5513# a_14018_5121# VDD.t31 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X307 a_12410_10219# eob.t16 a_12322_10081# VDD.t126 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X308 x2.x9.output_stack x2.x6.SW x2.x6.floating VDD.t129 sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X309 x2.x4[3].floating delay_code[2].t1 x2.x9.output_stack VSS.t110 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X310 a_12385_8830# eob.t17 a_12297_8830# VSS.t72 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X311 a_12457_8140# eob.t18 a_12385_8140# VSS.t87 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X312 VSS.t232 a_17191_5761# a_17898_5803# VSS.t230 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X313 a_17103_7067# a_15955_7073# a_17017_7445# VDD.t19 sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X314 VSS.t43 VDD.t259 a_14312_5987# VSS.t42 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X315 a_17307_5147# a_16704_5121# a_17191_5121# VSS.t172 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X316 a_17307_5147# VDD.t260 VSS.t82 VSS.t81 sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X317 sar_retimer[5].t0 a_17898_5803# VSS.t46 VSS.t45 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X318 a_12457_8416# eob.t19 a_12385_8416# VSS.t87 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X319 x1[3].Q_N a_17191_6401# VSS.t227 VSS.t226 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X320 a_15033_5429# a_14625_5147# a_14799_5121# VDD.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X321 a_14711_7067# a_13563_7073# a_14625_7445# VDD.t198 sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X322 a_14915_6427# a_14312_6401# a_14799_6401# VSS.t34 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X323 sar_retimer[4].t0 a_15506_5803# VSS.t68 VSS.t67 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X324 a_14625_6427# a_13397_6427# a_14483_6709# VDD.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X325 VDD.t156 a_14799_6401# a_14711_6793# VDD.t155 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X326 a_14915_5147# VDD.t261 VSS.t84 VSS.t83 sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X327 VDD.t202 a_16704_5121# a_17425_5429# VDD.t201 sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X328 a_12385_8002# eob.t20 a_12297_8002# VSS.t72 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X329 a_16410_6401# a_16236_6793# a_16550_6427# VSS.t97 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X330 a_14158_6153# VDD.t262 VSS.t86 VSS.t85 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X331 a_17017_7445# a_15789_7073# a_16875_7067# VDD.t216 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X332 VDD.t32 a_14312_6401# a_15033_6709# VDD.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X333 a_16344_6427# a_15955_6427# a_16236_6793# VSS.t74 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X334 a_16320_5787# a_15789_5793# a_16236_5787# VDD.t133 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X335 VDD.t16 a_14799_5121# a_15506_5147# VDD.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X336 x1[7].Q_N a_17191_5121# VDD.t206 VDD.t205 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X337 VSS.t89 delay_offset.t2 x2.x6.SW VSS.t88 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X338 x2.x9.output_stack delay_code[2].t2 x2.x4[3].floating VSS.t98 sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X339 a_16922_7389# a_16410_7041# VSS.t183 VSS.t182 sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X340 a_14530_6427# a_14018_6401# VSS.t78 VSS.t77 sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X341 VDD.t190 a_14018_5761# a_13928_5787# VDD.t25 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X342 a_17191_5121# VDD.t64 VDD.t66 VDD.t65 sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X343 VSS.t154 a_18499_9105# x3.X VSS.t153 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X344 VDD.t178 x3.X a_13397_7073# VDD.t177 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X345 a_16344_6165# a_15955_5793# a_16236_5787# VSS.t74 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X346 x2.x5[7].floating.t0 x2.x10.Y.t9 x2.x9.output_stack VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X347 a_13952_6427# a_13563_6427# a_13844_6793# VSS.t54 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X348 x1[2].Q_N a_14799_6401# VDD.t154 VDD.t153 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X349 VSS.t101 a_14799_5761# a_15506_5803# VSS.t100 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X350 a_17017_5147# a_15955_5147# a_16922_5147# VSS.t65 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X351 a_16143_7067# sar_logic[1].t1 VSS.t92 VSS.t91 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X352 a_15955_6427# a_15789_6427# VDD.t238 VDD.t218 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X353 a_14158_5147# a_14312_5121# a_14018_5121# VSS.t69 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X354 x2.x4[3].floating delay_code[2].t3 x2.x9.output_stack VSS.t73 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X355 VSS.t142 x3.X a_15789_7073# VSS.t141 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X356 a_14625_6427# a_13563_6427# a_14530_6427# VSS.t53 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X357 a_13952_6165# a_13563_5793# a_13844_5787# VSS.t54 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X358 VDD.t176 x3.X a_15789_5147# VDD.t175 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X359 a_12457_8692# eob.t21 a_12385_8830# VSS.t87 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X360 a_13751_7067# sar_logic[0].t1 VSS.t14 VSS.t13 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X361 a_14915_7433# a_14312_7267# a_14799_7041# VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X362 VSS.t130 a_17191_7041# a_17126_7445# VSS.t129 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X363 a_13928_6793# a_13397_6427# a_13844_6793# VDD.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X364 a_14625_6165# a_13563_5793# a_14530_6109# VSS.t53 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X365 a_14625_5147# a_13397_5147# a_14483_5429# VDD.t141 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X366 VSS.t181 a_16410_7041# a_16344_7445# VSS.t180 sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X367 a_15955_6427# a_15789_6427# VSS.t241 VSS.t169 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X368 a_17126_5147# a_15789_5147# a_17017_5147# VSS.t93 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X369 VDD.t14 a_14799_5121# a_14711_5513# VDD.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X370 a_14799_7041# VDD.t61 VDD.t63 VDD.t62 sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X371 x1[5].Q_N a_17191_5761# VDD.t227 VDD.t205 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X372 a_18195_9015# x2.x9.output_stack x3.A VSS.t137 sky130_fd_pr__nfet_01v8 ad=0.0651 pd=0.73 as=0.122 ps=1.42 w=0.42 l=0.15
X373 a_17425_7067# a_17017_7445# a_17191_7041# VDD.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X374 a_13563_5793# a_13397_5793# VSS.t99 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X375 a_16143_5147# sar_logic[7].t1 VSS.t24 VSS.t23 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X376 VSS.t140 x3.X a_15789_5147# VSS.t139 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
R0 VSS.n751 VSS 23902
R1 VSS.n1054 VSS.n1053 5020.45
R2 VSS.n752 VSS.n751 3808.6
R3 VSS.n2175 VSS 1043.16
R4 VSS.n507 VSS 1041.74
R5 VSS.t139 VSS 644.237
R6 VSS.t149 VSS 644.237
R7 VSS.n2147 VSS.t88 641.946
R8 VSS.n262 VSS.t94 616.822
R9 VSS.n703 VSS.t222 616.822
R10 VSS.n287 VSS.t111 603.115
R11 VSS.n482 VSS.t23 603.115
R12 VSS.n499 VSS.t139 603.115
R13 VSS.n525 VSS.t56 603.115
R14 VSS.n228 VSS.t47 603.115
R15 VSS.n742 VSS.t149 603.115
R16 VSS.n1053 VSS.n1052 598.058
R17 VSS.n280 VSS.t174 561.995
R18 VSS.n532 VSS.t17 561.995
R19 VSS.n499 VSS.t95 548.288
R20 VSS.n742 VSS.t224 548.288
R21 VSS.n912 VSS 541.101
R22 VSS.n1685 VSS.n1594 538.854
R23 VSS.n1084 VSS.n51 533.059
R24 VSS.n1089 VSS.n51 533.059
R25 VSS.n1089 VSS.n33 533.059
R26 VSS.n1125 VSS.n33 533.059
R27 VSS.n1125 VSS.n20 533.059
R28 VSS.n2048 VSS.n20 533.059
R29 VSS.n2048 VSS.n21 533.059
R30 VSS.n2044 VSS.n21 533.059
R31 VSS.n2044 VSS.n1146 533.059
R32 VSS.n2035 VSS.n1146 533.059
R33 VSS.n2035 VSS.n1154 533.059
R34 VSS.n2018 VSS.n1154 533.059
R35 VSS.n2018 VSS.n1184 533.059
R36 VSS.n1269 VSS.n1184 533.059
R37 VSS.n1269 VSS.n1203 533.059
R38 VSS.n2001 VSS.n1203 533.059
R39 VSS.n2001 VSS.n1204 533.059
R40 VSS.n1980 VSS.n1204 533.059
R41 VSS.n1980 VSS.n1298 533.059
R42 VSS.n1346 VSS.n1298 533.059
R43 VSS.n1953 VSS.n1346 533.059
R44 VSS.n1953 VSS.n1347 533.059
R45 VSS.n1949 VSS.n1347 533.059
R46 VSS.n1949 VSS.n1350 533.059
R47 VSS.n1435 VSS.n1350 533.059
R48 VSS.n1445 VSS.n1435 533.059
R49 VSS.n1445 VSS.n1392 533.059
R50 VSS.n1916 VSS.n1392 533.059
R51 VSS.n1916 VSS.n1393 533.059
R52 VSS.n1510 VSS.n1393 533.059
R53 VSS.n1510 VSS.n1468 533.059
R54 VSS.n1897 VSS.n1468 533.059
R55 VSS.n1897 VSS.n1469 533.059
R56 VSS.n1890 VSS.n1469 533.059
R57 VSS.n1890 VSS.n1476 533.059
R58 VSS.n1618 VSS.n1476 533.059
R59 VSS.n1618 VSS.n1613 533.059
R60 VSS.n1627 VSS.n1613 533.059
R61 VSS.n1627 VSS.n1593 533.059
R62 VSS.n1843 VSS.n1593 533.059
R63 VSS.n1843 VSS.n1594 533.059
R64 VSS.n1681 VSS.n1667 533.059
R65 VSS.n1822 VSS.n1667 533.059
R66 VSS.n1822 VSS.n1668 533.059
R67 VSS.n1800 VSS.n1668 533.059
R68 VSS.n1800 VSS.n1738 533.059
R69 VSS.n1780 VSS.n1738 533.059
R70 VSS.n1780 VSS.n7 533.059
R71 VSS.n2061 VSS.n7 533.059
R72 VSS.n1685 VSS.n1681 527.265
R73 VSS.n359 VSS.t64 520.872
R74 VSS.n597 VSS.t242 520.872
R75 VSS.n307 VSS.t176 507.166
R76 VSS.n554 VSS.t19 507.166
R77 VSS VSS.n752 484.142
R78 VSS.n330 VSS.t209 466.045
R79 VSS.n561 VSS.t185 466.045
R80 VSS.n256 VSS.t66 424.923
R81 VSS.n686 VSS.t7 424.923
R82 VSS.n354 VSS.t172 411.216
R83 VSS.n590 VSS.t70 411.216
R84 VSS.n2111 VSS.n2110 405.82
R85 VSS.t153 VSS.n87 402.445
R86 VSS.n251 VSS.t166 370.094
R87 VSS.n681 VSS.t27 370.094
R88 VSS.t145 VSS 334.628
R89 VSS.t143 VSS 334.628
R90 VSS.n2147 VSS 320.974
R91 VSS.n938 VSS.t171 320.389
R92 VSS.n769 VSS.t2 320.389
R93 VSS.n1046 VSS.t45 313.269
R94 VSS.n890 VSS.t51 313.269
R95 VSS.n904 VSS.t145 313.269
R96 VSS.n919 VSS.t67 313.269
R97 VSS.n777 VSS.t10 313.269
R98 VSS.n756 VSS.t143 313.269
R99 VSS.n230 VSS.n229 295.61
R100 VSS.n1740 VSS.n1738 295.61
R101 VSS.n1347 VSS.n1344 295.61
R102 VSS.n484 VSS.n483 295.61
R103 VSS.n2149 VSS.n2148 292.5
R104 VSS.n2148 VSS.n2147 292.5
R105 VSS.n1051 VSS.n1050 292.5
R106 VSS.n1052 VSS.n1051 292.5
R107 VSS.n1048 VSS.n1047 292.5
R108 VSS.n1047 VSS.n1046 292.5
R109 VSS.n1040 VSS.n1039 292.5
R110 VSS.n1039 VSS.n1038 292.5
R111 VSS.n1036 VSS.n1035 292.5
R112 VSS.n1035 VSS.n1034 292.5
R113 VSS.n1031 VSS.n1030 292.5
R114 VSS.n1030 VSS.n1029 292.5
R115 VSS.n1024 VSS.n1023 292.5
R116 VSS.n1023 VSS.n1022 292.5
R117 VSS.n1017 VSS.n1016 292.5
R118 VSS.n1016 VSS.n1015 292.5
R119 VSS.n1010 VSS.n1009 292.5
R120 VSS.n1009 VSS.n1008 292.5
R121 VSS.n1005 VSS.n1004 292.5
R122 VSS.n1004 VSS.n1003 292.5
R123 VSS.n112 VSS.n111 292.5
R124 VSS.n111 VSS.n110 292.5
R125 VSS.n116 VSS.n115 292.5
R126 VSS.n115 VSS.n114 292.5
R127 VSS.n126 VSS.n125 292.5
R128 VSS.n125 VSS.n124 292.5
R129 VSS.n121 VSS.n120 292.5
R130 VSS.n120 VSS.n119 292.5
R131 VSS.n961 VSS.n960 292.5
R132 VSS.n960 VSS.n959 292.5
R133 VSS.n967 VSS.n966 292.5
R134 VSS.n966 VSS.n965 292.5
R135 VSS.n971 VSS.n970 292.5
R136 VSS.n970 VSS.n969 292.5
R137 VSS.n974 VSS.n973 292.5
R138 VSS.n973 VSS.t97 292.5
R139 VSS.n142 VSS.n141 292.5
R140 VSS.n141 VSS.n140 292.5
R141 VSS.n150 VSS.n149 292.5
R142 VSS.n149 VSS.n148 292.5
R143 VSS.n936 VSS.n935 292.5
R144 VSS.n935 VSS.n934 292.5
R145 VSS.n940 VSS.n939 292.5
R146 VSS.n939 VSS.n938 292.5
R147 VSS.n944 VSS.n943 292.5
R148 VSS.n943 VSS.n942 292.5
R149 VSS.n892 VSS.n891 292.5
R150 VSS.n891 VSS.n890 292.5
R151 VSS.n899 VSS.n898 292.5
R152 VSS.n898 VSS.n897 292.5
R153 VSS.n906 VSS.n905 292.5
R154 VSS.n905 VSS.n904 292.5
R155 VSS.n910 VSS.n909 292.5
R156 VSS.n911 VSS.n910 292.5
R157 VSS.n914 VSS.n913 292.5
R158 VSS.n913 VSS.n912 292.5
R159 VSS.n921 VSS.n920 292.5
R160 VSS.n920 VSS.n919 292.5
R161 VSS.n876 VSS.n875 292.5
R162 VSS.n875 VSS.n874 292.5
R163 VSS.n880 VSS.n879 292.5
R164 VSS.n879 VSS.n878 292.5
R165 VSS.n856 VSS.n855 292.5
R166 VSS.n855 VSS.n854 292.5
R167 VSS.n864 VSS.n863 292.5
R168 VSS.n863 VSS.n862 292.5
R169 VSS.n161 VSS.n160 292.5
R170 VSS.n160 VSS.n159 292.5
R171 VSS.n165 VSS.n164 292.5
R172 VSS.n164 VSS.n163 292.5
R173 VSS.n169 VSS.n168 292.5
R174 VSS.n168 VSS.n167 292.5
R175 VSS.n182 VSS.n181 292.5
R176 VSS.n181 VSS.n180 292.5
R177 VSS.n186 VSS.n185 292.5
R178 VSS.n185 VSS.n184 292.5
R179 VSS.n830 VSS.n829 292.5
R180 VSS.n829 VSS.n828 292.5
R181 VSS.n834 VSS.n833 292.5
R182 VSS.n833 VSS.n832 292.5
R183 VSS.n838 VSS.n837 292.5
R184 VSS.n837 VSS.n836 292.5
R185 VSS.n814 VSS.n813 292.5
R186 VSS.n813 VSS.n812 292.5
R187 VSS.n818 VSS.n817 292.5
R188 VSS.n817 VSS.n816 292.5
R189 VSS.n195 VSS.n194 292.5
R190 VSS.n194 VSS.n193 292.5
R191 VSS.n199 VSS.n198 292.5
R192 VSS.n198 VSS.n197 292.5
R193 VSS.n794 VSS.n793 292.5
R194 VSS.n793 VSS.n792 292.5
R195 VSS.n798 VSS.n797 292.5
R196 VSS.n797 VSS.n796 292.5
R197 VSS.n771 VSS.n770 292.5
R198 VSS.n770 VSS.n769 292.5
R199 VSS.n775 VSS.n774 292.5
R200 VSS.n774 VSS.n773 292.5
R201 VSS.n779 VSS.n778 292.5
R202 VSS.n778 VSS.n777 292.5
R203 VSS.n208 VSS.n207 292.5
R204 VSS.n207 VSS.n206 292.5
R205 VSS.n758 VSS.n757 292.5
R206 VSS.n757 VSS.n756 292.5
R207 VSS.n754 VSS.n753 292.5
R208 VSS.n755 VSS.n754 292.5
R209 VSS.n1059 VSS.n1058 292.5
R210 VSS.n1058 VSS.n1057 292.5
R211 VSS.n1056 VSS.n1055 292.5
R212 VSS.n89 VSS.n88 292.5
R213 VSS.n1084 VSS.n1083 292.5
R214 VSS.n1085 VSS.n1084 292.5
R215 VSS.n2061 VSS.n2060 292.5
R216 VSS.n2062 VSS.n2061 292.5
R217 VSS.n1784 VSS.n7 292.5
R218 VSS.n1778 VSS.n7 292.5
R219 VSS.n1781 VSS.n1780 292.5
R220 VSS.n1780 VSS.n1779 292.5
R221 VSS.n1777 VSS.n1738 292.5
R222 VSS.n1800 VSS.n1799 292.5
R223 VSS.n1801 VSS.n1800 292.5
R224 VSS.n1739 VSS.n1668 292.5
R225 VSS.n1736 VSS.n1668 292.5
R226 VSS.n1822 VSS.n1821 292.5
R227 VSS.n1823 VSS.n1822 292.5
R228 VSS.n1681 VSS.n1673 292.5
R229 VSS.n1684 VSS.n1681 292.5
R230 VSS.n1702 VSS.n1667 292.5
R231 VSS.n1683 VSS.n1667 292.5
R232 VSS.n1686 VSS.n1685 292.5
R233 VSS.n1685 VSS.t44 292.5
R234 VSS.n1675 VSS.n1594 292.5
R235 VSS.n1682 VSS.n1594 292.5
R236 VSS.n1843 VSS.n1842 292.5
R237 VSS.n1844 VSS.n1843 292.5
R238 VSS.n1629 VSS.n1593 292.5
R239 VSS.n1621 VSS.n1593 292.5
R240 VSS.n1628 VSS.n1627 292.5
R241 VSS.n1627 VSS.n1626 292.5
R242 VSS.n1613 VSS.n1609 292.5
R243 VSS.n1620 VSS.n1613 292.5
R244 VSS.n1618 VSS.n1617 292.5
R245 VSS.n1619 VSS.n1618 292.5
R246 VSS.n1476 VSS.n1474 292.5
R247 VSS.n1614 VSS.n1476 292.5
R248 VSS.n1891 VSS.n1890 292.5
R249 VSS.n1890 VSS.n1889 292.5
R250 VSS.n1892 VSS.n1469 292.5
R251 VSS.n1477 VSS.n1469 292.5
R252 VSS.n1897 VSS.n1896 292.5
R253 VSS.n1898 VSS.n1897 292.5
R254 VSS.n1514 VSS.n1468 292.5
R255 VSS.n1468 VSS.n1466 292.5
R256 VSS.n1511 VSS.n1510 292.5
R257 VSS.n1510 VSS.n1509 292.5
R258 VSS.n1395 VSS.n1393 292.5
R259 VSS.n1508 VSS.n1393 292.5
R260 VSS.n1916 VSS.n1915 292.5
R261 VSS.n1917 VSS.n1916 292.5
R262 VSS.n1449 VSS.n1392 292.5
R263 VSS.n1392 VSS.n1391 292.5
R264 VSS.n1435 VSS.n1434 292.5
R265 VSS.n1438 VSS.n1435 292.5
R266 VSS.n1446 VSS.n1445 292.5
R267 VSS.n1445 VSS.n1444 292.5
R268 VSS.n1351 VSS.n1350 292.5
R269 VSS.n1437 VSS.n1350 292.5
R270 VSS.n1949 VSS.n1948 292.5
R271 VSS.n1950 VSS.n1949 292.5
R272 VSS.n1951 VSS.n1347 292.5
R273 VSS.n1954 VSS.n1953 292.5
R274 VSS.n1953 VSS.n1952 292.5
R275 VSS.n1346 VSS.n1343 292.5
R276 VSS.n1349 VSS.n1346 292.5
R277 VSS.n1342 VSS.n1298 292.5
R278 VSS.n1300 VSS.n1298 292.5
R279 VSS.n1981 VSS.n1980 292.5
R280 VSS.n1980 VSS.n1979 292.5
R281 VSS.n1204 VSS.n1201 292.5
R282 VSS.n1272 VSS.n1204 292.5
R283 VSS.n2002 VSS.n2001 292.5
R284 VSS.n2001 VSS.n2000 292.5
R285 VSS.n1203 VSS.n1200 292.5
R286 VSS.n1271 VSS.n1203 292.5
R287 VSS.n1269 VSS.n1268 292.5
R288 VSS.n1270 VSS.n1269 292.5
R289 VSS.n1263 VSS.n1184 292.5
R290 VSS.n1188 VSS.n1184 292.5
R291 VSS.n2019 VSS.n2018 292.5
R292 VSS.n2018 VSS.n2017 292.5
R293 VSS.n2020 VSS.n1154 292.5
R294 VSS.n1185 VSS.n1154 292.5
R295 VSS.n2036 VSS.n2035 292.5
R296 VSS.n2035 VSS.n2034 292.5
R297 VSS.n2039 VSS.n1146 292.5
R298 VSS.n1155 VSS.n1146 292.5
R299 VSS.n21 VSS.n19 292.5
R300 VSS.n2046 VSS.n21 292.5
R301 VSS.n2044 VSS.n2043 292.5
R302 VSS.n2045 VSS.n2044 292.5
R303 VSS.n2049 VSS.n2048 292.5
R304 VSS.n2048 VSS.n2047 292.5
R305 VSS.n1126 VSS.n1125 292.5
R306 VSS.n1125 VSS.n1124 292.5
R307 VSS.n1129 VSS.n20 292.5
R308 VSS.n1145 VSS.n20 292.5
R309 VSS.n1091 VSS.n33 292.5
R310 VSS.n34 VSS.n33 292.5
R311 VSS.n51 VSS.n49 292.5
R312 VSS.n1086 VSS.n51 292.5
R313 VSS.n1090 VSS.n1089 292.5
R314 VSS.n1089 VSS.n1088 292.5
R315 VSS.n437 VSS.n436 292.5
R316 VSS.n436 VSS.n435 292.5
R317 VSS.n744 VSS.n743 292.5
R318 VSS.n743 VSS.n742 292.5
R319 VSS.n749 VSS.n748 292.5
R320 VSS.n750 VSS.n749 292.5
R321 VSS.n738 VSS.n737 292.5
R322 VSS.n737 VSS.n736 292.5
R323 VSS.n229 VSS.n228 292.5
R324 VSS.n247 VSS.n246 292.5
R325 VSS.n246 VSS.n245 292.5
R326 VSS.n253 VSS.n252 292.5
R327 VSS.n252 VSS.n251 292.5
R328 VSS.n258 VSS.n257 292.5
R329 VSS.n257 VSS.n256 292.5
R330 VSS.n264 VSS.n263 292.5
R331 VSS.n263 VSS.n262 292.5
R332 VSS.n269 VSS.n268 292.5
R333 VSS.n268 VSS.n267 292.5
R334 VSS.n278 VSS.n277 292.5
R335 VSS.n277 VSS.n276 292.5
R336 VSS.n290 VSS.n288 292.5
R337 VSS.n288 VSS.n287 292.5
R338 VSS.n282 VSS.n281 292.5
R339 VSS.n281 VSS.n280 292.5
R340 VSS.n314 VSS.n313 292.5
R341 VSS.n313 VSS.n312 292.5
R342 VSS.n309 VSS.n308 292.5
R343 VSS.n308 VSS.n307 292.5
R344 VSS.n332 VSS.n331 292.5
R345 VSS.n331 VSS.n330 292.5
R346 VSS.n337 VSS.n336 292.5
R347 VSS.n336 VSS.n335 292.5
R348 VSS.n356 VSS.n355 292.5
R349 VSS.n355 VSS.n354 292.5
R350 VSS.n361 VSS.n360 292.5
R351 VSS.n360 VSS.n359 292.5
R352 VSS.n377 VSS.n376 292.5
R353 VSS.n376 VSS.n375 292.5
R354 VSS.n385 VSS.n383 292.5
R355 VSS.n383 VSS.n382 292.5
R356 VSS.n401 VSS.n400 292.5
R357 VSS.n400 VSS.n399 292.5
R358 VSS.n408 VSS.n407 292.5
R359 VSS.n407 VSS.n406 292.5
R360 VSS.n414 VSS.n413 292.5
R361 VSS.n413 VSS.n412 292.5
R362 VSS.n432 VSS.n431 292.5
R363 VSS.n431 VSS.n430 292.5
R364 VSS.n441 VSS.n440 292.5
R365 VSS.n440 VSS.n439 292.5
R366 VSS.n483 VSS.n482 292.5
R367 VSS.n674 VSS.n673 292.5
R368 VSS.n673 VSS.n672 292.5
R369 VSS.n683 VSS.n682 292.5
R370 VSS.n682 VSS.n681 292.5
R371 VSS.n688 VSS.n687 292.5
R372 VSS.n687 VSS.n686 292.5
R373 VSS.n705 VSS.n704 292.5
R374 VSS.n704 VSS.n703 292.5
R375 VSS.n710 VSS.n709 292.5
R376 VSS.n709 VSS.n708 292.5
R377 VSS.n659 VSS.n657 292.5
R378 VSS.n657 VSS.n656 292.5
R379 VSS.n651 VSS.n650 292.5
R380 VSS.n650 VSS.n649 292.5
R381 VSS.n626 VSS.n625 292.5
R382 VSS.n625 VSS.n624 292.5
R383 VSS.n621 VSS.n620 292.5
R384 VSS.n620 VSS.n619 292.5
R385 VSS.n492 VSS.n491 292.5
R386 VSS.n491 VSS.n490 292.5
R387 VSS.n501 VSS.n500 292.5
R388 VSS.n500 VSS.n499 292.5
R389 VSS.n505 VSS.n504 292.5
R390 VSS.n506 VSS.n505 292.5
R391 VSS.n510 VSS.n508 292.5
R392 VSS.n508 VSS.n507 292.5
R393 VSS.n527 VSS.n526 292.5
R394 VSS.n526 VSS.n525 292.5
R395 VSS.n534 VSS.n533 292.5
R396 VSS.n533 VSS.n532 292.5
R397 VSS.n539 VSS.n538 292.5
R398 VSS.n538 VSS.n537 292.5
R399 VSS.n556 VSS.n555 292.5
R400 VSS.n555 VSS.n554 292.5
R401 VSS.n563 VSS.n562 292.5
R402 VSS.n562 VSS.n561 292.5
R403 VSS.n568 VSS.n567 292.5
R404 VSS.n567 VSS.n566 292.5
R405 VSS.n592 VSS.n591 292.5
R406 VSS.n591 VSS.n590 292.5
R407 VSS.n599 VSS.n598 292.5
R408 VSS.n598 VSS.n597 292.5
R409 VSS.n608 VSS.n607 292.5
R410 VSS.n607 VSS.n606 292.5
R411 VSS.n612 VSS.n611 292.5
R412 VSS.n611 VSS.n610 292.5
R413 VSS.n617 VSS.n616 292.5
R414 VSS.n616 VSS.n615 292.5
R415 VSS.n630 VSS.n629 292.5
R416 VSS.n629 VSS.n628 292.5
R417 VSS VSS.t240 292.454
R418 VSS.n1038 VSS.t230 291.909
R419 VSS.n874 VSS.t100 291.909
R420 VSS.n904 VSS.t169 284.791
R421 VSS.n756 VSS.t4 284.791
R422 VSS.n1003 VSS.t9 270.55
R423 VSS.n2064 VSS.t12 270.466
R424 VSS.n1029 VSS.t226 263.43
R425 VSS.n167 VSS.t8 263.43
R426 VSS.n854 VSS.t102 256.312
R427 VSS.n382 VSS.t178 246.73
R428 VSS.n610 VSS.t15 246.73
R429 VSS.n1022 VSS.t40 242.071
R430 VSS.n862 VSS.t42 242.071
R431 VSS.n1121 VSS.n35 231.766
R432 VSS.n1121 VSS.n22 231.766
R433 VSS.n1143 VSS.n22 231.766
R434 VSS.n2032 VSS.n1156 231.766
R435 VSS.n1187 VSS.n1156 231.766
R436 VSS.n2014 VSS.n1187 231.766
R437 VSS.n1998 VSS.n1273 231.766
R438 VSS.n1977 VSS.n1273 231.766
R439 VSS.n1977 VSS.n1301 231.766
R440 VSS.n1441 VSS.n1440 231.766
R441 VSS.n1441 VSS.n1389 231.766
R442 VSS.n1919 VSS.n1389 231.766
R443 VSS.n1900 VSS.n1465 231.766
R444 VSS.n1479 VSS.n1465 231.766
R445 VSS.n1887 VSS.n1479 231.766
R446 VSS.n1624 VSS.n1590 231.766
R447 VSS.n1846 VSS.n1590 231.766
R448 VSS.n1846 VSS.n1591 231.766
R449 VSS.n1825 VSS.n1666 231.766
R450 VSS.n1803 VSS.n1666 231.766
R451 VSS.n1803 VSS.n1734 231.766
R452 VSS.n934 VSS.t74 220.713
R453 VSS.n796 VSS.t54 220.713
R454 VSS VSS.n506 219.315
R455 VSS VSS.n750 219.315
R456 VSS.n1008 VSS.t58 213.593
R457 VSS.n163 VSS.t34 213.593
R458 VSS.t240 VSS.t239 211.095
R459 VSS.n399 VSS.t93 205.607
R460 VSS.n615 VSS.t223 205.607
R461 VSS.t239 VSS.t137 202.299
R462 VSS.n2047 VSS.n1145 202.299
R463 VSS.n1951 VSS.n1950 202.299
R464 VSS.n1626 VSS.n1620 202.299
R465 VSS.n1779 VSS.n1777 202.299
R466 VSS.n2136 VSS.n2135 200.608
R467 VSS.t44 VSS.n1684 200.101
R468 VSS.n2110 VSS.t87 198.263
R469 VSS.n148 VSS.t31 192.233
R470 VSS.n792 VSS.t79 192.233
R471 VSS.n1270 VSS.t182 191.304
R472 VSS.t184 VSS.n1999 189.106
R473 VSS.n1205 VSS.t183 184.713
R474 VSS.n1595 VSS.t163 184.713
R475 VSS.n958 VSS.t30 184.713
R476 VSS.n958 VSS.t63 184.713
R477 VSS.n811 VSS.t78 184.713
R478 VSS.n811 VSS.t158 184.713
R479 VSS.n411 VSS.t165 184.713
R480 VSS.n618 VSS.t26 184.713
R481 VSS.t73 VSS.t1 182.51
R482 VSS.n2045 VSS.t36 175.912
R483 VSS.n2016 VSS.n2015 175.912
R484 VSS.n1625 VSS.n1622 175.912
R485 VSS.n2177 VSS.n2176 173.861
R486 VSS.t126 VSS.n1619 169.315
R487 VSS.n1917 VSS.t110 167.117
R488 VSS.n375 VSS.t81 164.487
R489 VSS.n606 VSS.t83 164.487
R490 VSS.t129 VSS.n1155 162.72
R491 VSS.t117 VSS.n1614 162.72
R492 VSS.n2017 VSS.n1186 160.52
R493 VSS.n1085 VSS.t137 158.321
R494 VSS.n1888 VSS.t38 156.123
R495 VSS.n1845 VSS.t162 149.525
R496 VSS.n2177 VSS.t49 147.113
R497 VSS.n1271 VSS.t215 145.127
R498 VSS.n1299 VSS.t203 145.127
R499 VSS.n231 VSS.t48 144.97
R500 VSS.n1771 VSS.t14 144.97
R501 VSS.n1352 VSS.t92 144.97
R502 VSS.n485 VSS.t24 144.97
R503 VSS.n779 VSS.t11 141.861
R504 VSS.n779 VSS.t55 141.861
R505 VSS.n892 VSS.t71 141.861
R506 VSS.n892 VSS.t52 141.861
R507 VSS.t109 VSS.n1683 136.333
R508 VSS.n114 VSS.t228 135.275
R509 VSS.n1844 VSS.n1592 134.133
R510 VSS.n1087 VSS.n34 129.736
R511 VSS.n184 VSS.t104 128.155
R512 VSS.n439 VSS.t173 123.365
R513 VSS.n245 VSS.t195 123.365
R514 VSS.n649 VSS.t69 123.365
R515 VSS.n672 VSS.t189 123.365
R516 VSS.t119 VSS.n1508 120.941
R517 VSS.n2046 VSS.t76 118.742
R518 VSS.n1442 VSS 116.543
R519 VSS.n1950 VSS.t219 114.344
R520 VSS.n1779 VSS.t123 114.344
R521 VSS VSS.n911 113.916
R522 VSS.n755 VSS 113.916
R523 VSS.n1296 VSS.n1295 113.207
R524 VSS.n1701 VSS.n1672 113.207
R525 VSS.n147 VSS.n145 113.207
R526 VSS.n147 VSS.n146 113.207
R527 VSS.n791 VSS.n789 113.207
R528 VSS.n791 VSS.n790 113.207
R529 VSS.n250 VSS.n249 113.207
R530 VSS.n679 VSS.n678 113.207
R531 VSS.t131 VSS.n1086 112.144
R532 VSS.n1123 VSS.t211 107.746
R533 VSS.n2149 VSS.t89 107.195
R534 VSS.n2170 VSS.t50 107.195
R535 VSS.n124 VSS.t168 106.796
R536 VSS.n828 VSS.t3 106.796
R537 VSS.n2038 VSS.n1151 106.038
R538 VSS.n1616 VSS.n1615 106.038
R539 VSS.n109 VSS.n107 106.038
R540 VSS.n109 VSS.n108 106.038
R541 VSS.n179 VSS.n177 106.038
R542 VSS.n179 VSS.n178 106.038
R543 VSS.n374 VSS.n373 106.038
R544 VSS.n605 VSS.n604 106.038
R545 VSS.t237 VSS.n1056 105.547
R546 VSS.t127 VSS.n1085 105.547
R547 VSS.n1952 VSS.t91 105.547
R548 VSS.n1444 VSS.t60 105.547
R549 VSS.n53 VSS.n52 105.3
R550 VSS.n1448 VSS.n1428 105.3
R551 VSS.n1045 VSS.n1043 105.3
R552 VSS.n1045 VSS.n1044 105.3
R553 VSS.n918 VSS.n916 105.3
R554 VSS.n918 VSS.n917 105.3
R555 VSS.n291 VSS.n286 105.3
R556 VSS.n524 VSS.n523 105.3
R557 VSS.n82 VSS.t154 104.15
R558 VSS.n741 VSS.n740 103.942
R559 VSS.n1783 VSS.n1782 103.942
R560 VSS.n1127 VSS.n30 103.942
R561 VSS.n1513 VSS.n1504 103.942
R562 VSS.n1431 VSS.n1430 103.942
R563 VSS.n86 VSS.n85 103.942
R564 VSS.n1028 VSS.n1026 103.942
R565 VSS.n1028 VSS.n1027 103.942
R566 VSS.n903 VSS.n901 103.942
R567 VSS.n903 VSS.n902 103.942
R568 VSS.n859 VSS.n857 103.942
R569 VSS.n859 VSS.n858 103.942
R570 VSS.n213 VSS.n211 103.942
R571 VSS.n213 VSS.n212 103.942
R572 VSS.n306 VSS.n305 103.942
R573 VSS.n498 VSS.n497 103.942
R574 VSS.n553 VSS.n552 103.942
R575 VSS.t213 VSS.t136 103.349
R576 VSS.n1952 VSS.t221 103.349
R577 VSS.n1899 VSS.n1898 103.349
R578 VSS.t125 VSS.n1801 103.349
R579 VSS.t151 VSS 103.349
R580 VSS.n2033 VSS.t218 101.15
R581 VSS.t221 VSS.n1349 98.951
R582 VSS.n1918 VSS.n1391 98.951
R583 VSS.n1899 VSS.n1466 98.951
R584 VSS.n1054 VSS.t155 96.7521
R585 VSS.n1057 VSS.t237 96.7521
R586 VSS.n1086 VSS.t127 96.7521
R587 VSS.t91 VSS.n1951 96.7521
R588 VSS.t141 VSS.n1437 96.7521
R589 VSS.t98 VSS.t193 96.7521
R590 VSS.n1777 VSS.t13 96.7521
R591 VSS.n1778 VSS.t151 96.7521
R592 VSS.n89 VSS.t153 94.5532
R593 VSS.n1736 VSS.n1735 94.5532
R594 VSS.n2137 VSS.n2133 93.0283
R595 VSS.t155 VSS.n89 90.1554
R596 VSS.n1088 VSS.t131 90.1554
R597 VSS.n1349 VSS.n1348 90.1554
R598 VSS.t121 VSS.n1917 90.1554
R599 VSS.n1437 VSS.t219 87.9565
R600 VSS.t123 VSS.n1778 87.9565
R601 VSS.n110 VSS.t197 85.4374
R602 VSS.n180 VSS.t199 85.4374
R603 VSS.t76 VSS.n2045 83.5587
R604 VSS.n1889 VSS.t106 83.5587
R605 VSS.n1124 VSS.t133 81.3598
R606 VSS.n1439 VSS.t141 81.3598
R607 VSS.n1509 VSS.t119 81.3598
R608 VSS.n1802 VSS.n1736 81.3598
R609 VSS.n2000 VSS.t213 79.1609
R610 VSS.t180 VSS.n1978 79.1609
R611 VSS.n1066 VSS.t236 77.3934
R612 VSS.n1066 VSS.t235 77.3934
R613 VSS.n1443 VSS.n1391 76.962
R614 VSS.n1295 VSS.t181 75.7148
R615 VSS.n1672 VSS.t161 75.7148
R616 VSS.n146 VSS.t62 75.7148
R617 VSS.n145 VSS.t32 75.7148
R618 VSS.n790 VSS.t157 75.7148
R619 VSS.n789 VSS.t80 75.7148
R620 VSS.n249 VSS.t167 75.7148
R621 VSS.n678 VSS.t28 75.7148
R622 VSS.t133 VSS.n1122 74.7631
R623 VSS.t90 VSS.t135 74.7631
R624 VSS.t193 VSS.n1466 74.7631
R625 VSS.n1824 VSS.t160 74.7631
R626 VSS.t87 VSS.t72 74.3492
R627 VSS.n1088 VSS.n1087 72.5642
R628 VSS.n1898 VSS.n1467 72.5642
R629 VSS.n1478 VSS.t106 72.5642
R630 VSS.n2178 VSS.n2174 71.1394
R631 VSS.n412 VSS.t164 68.5363
R632 VSS.n624 VSS.t25 68.5363
R633 VSS.n1144 VSS.t211 68.1664
R634 VSS.n2034 VSS.n2033 68.1664
R635 VSS.t21 VSS.n1300 68.1664
R636 VSS.n1682 VSS.n1592 68.1664
R637 VSS.n1824 VSS.n1823 68.1664
R638 VSS.n1823 VSS.t217 68.1664
R639 VSS.t135 VSS.n2046 65.9675
R640 VSS.n1477 VSS.t0 65.9675
R641 VSS.n969 VSS.t59 64.0782
R642 VSS.n816 VSS.t35 64.0782
R643 VSS.n197 VSS.t85 64.0782
R644 VSS.n1978 VSS.n1300 63.7686
R645 VSS.t0 VSS.n1467 63.7686
R646 VSS.n2047 VSS.t90 61.5697
R647 VSS.n2064 VSS.n2063 61.5697
R648 VSS.n1979 VSS.t180 59.3708
R649 VSS.n1683 VSS.t160 59.3708
R650 VSS.t215 VSS.n1270 57.1719
R651 VSS.n140 VSS.t191 56.9584
R652 VSS.n1801 VSS.n1737 54.973
R653 VSS.n30 VSS.t212 54.2862
R654 VSS.n52 VSS.t132 54.2862
R655 VSS.n1504 VSS.t194 54.2862
R656 VSS.n1428 VSS.t122 54.2862
R657 VSS.n1044 VSS.t232 54.2862
R658 VSS.n1043 VSS.t231 54.2862
R659 VSS.n1027 VSS.t205 54.2862
R660 VSS.n1026 VSS.t41 54.2862
R661 VSS.n917 VSS.t101 54.2862
R662 VSS.n916 VSS.t115 54.2862
R663 VSS.n858 VSS.t43 54.2862
R664 VSS.n857 VSS.t201 54.2862
R665 VSS.n286 VSS.t175 54.2862
R666 VSS.n305 VSS.t210 54.2862
R667 VSS.n523 VSS.t18 54.2862
R668 VSS.n552 VSS.t186 54.2862
R669 VSS.n2176 VSS.n2175 53.4959
R670 VSS.n85 VSS.t238 51.4291
R671 VSS.n1444 VSS.n1442 50.5752
R672 VSS.t13 VSS.n1737 50.5752
R673 VSS.n1122 VSS.n34 46.1774
R674 VSS.n1478 VSS.n1477 46.1774
R675 VSS.t187 VSS.t109 46.1774
R676 VSS.n1348 VSS.t21 43.9785
R677 VSS.n80 VSS.t138 43.7547
R678 VSS.n1186 VSS.n1185 41.7796
R679 VSS.n1845 VSS.n1844 41.7796
R680 VSS.n2197 VSS.t107 41.4448
R681 VSS.n1151 VSS.t130 41.4291
R682 VSS.n1615 VSS.t118 41.4291
R683 VSS.n108 VSS.t234 41.4291
R684 VSS.n107 VSS.t229 41.4291
R685 VSS.n178 VSS.t105 41.4291
R686 VSS.n177 VSS.t114 41.4291
R687 VSS.n373 VSS.t179 41.4291
R688 VSS.n604 VSS.t16 41.4291
R689 VSS.n751 VSS.n227 40.2727
R690 VSS.n2034 VSS.t129 39.5807
R691 VSS.n1619 VSS.t117 39.5807
R692 VSS.n1735 VSS.t217 39.5807
R693 VSS.n740 VSS.t225 38.5719
R694 VSS.n740 VSS.t150 38.5719
R695 VSS.n1782 VSS.t124 38.5719
R696 VSS.n1782 VSS.t152 38.5719
R697 VSS.n1295 VSS.t204 38.5719
R698 VSS.n1151 VSS.t37 38.5719
R699 VSS.n1672 VSS.t188 38.5719
R700 VSS.n1615 VSS.t39 38.5719
R701 VSS.n1430 VSS.t220 38.5719
R702 VSS.n1430 VSS.t142 38.5719
R703 VSS.n108 VSS.t206 38.5719
R704 VSS.n107 VSS.t198 38.5719
R705 VSS.n146 VSS.t192 38.5719
R706 VSS.n145 VSS.t207 38.5719
R707 VSS.n902 VSS.t170 38.5719
R708 VSS.n902 VSS.t148 38.5719
R709 VSS.n901 VSS.t241 38.5719
R710 VSS.n901 VSS.t146 38.5719
R711 VSS.n178 VSS.t208 38.5719
R712 VSS.n177 VSS.t200 38.5719
R713 VSS.n790 VSS.t86 38.5719
R714 VSS.n789 VSS.t202 38.5719
R715 VSS.n212 VSS.t99 38.5719
R716 VSS.n212 VSS.t147 38.5719
R717 VSS.n211 VSS.t5 38.5719
R718 VSS.n211 VSS.t144 38.5719
R719 VSS.n373 VSS.t82 38.5719
R720 VSS.n249 VSS.t196 38.5719
R721 VSS.n497 VSS.t96 38.5719
R722 VSS.n497 VSS.t140 38.5719
R723 VSS.n604 VSS.t84 38.5719
R724 VSS.n678 VSS.t190 38.5719
R725 VSS.n1056 VSS 37.3818
R726 VSS.n1979 VSS.n1299 37.3818
R727 VSS.n959 VSS.t29 35.5992
R728 VSS.n836 VSS.t77 35.5992
R729 VSS.n1438 VSS 35.1829
R730 VSS.n1508 VSS.t110 35.1829
R731 VSS VSS.n2062 35.1829
R732 VSS.n1185 VSS.t218 32.984
R733 VSS.n1620 VSS.t126 32.984
R734 VSS.n1509 VSS.t98 30.7851
R735 VSS.n85 VSS.t156 28.7917
R736 VSS.n406 VSS.t65 27.4148
R737 VSS.n628 VSS.t6 27.4148
R738 VSS.n2135 VSS.n2134 26.7482
R739 VSS.n1155 VSS.t36 26.3873
R740 VSS.n1614 VSS.t38 26.3873
R741 VSS.n30 VSS.t134 25.9346
R742 VSS.n52 VSS.t128 25.9346
R743 VSS.n1504 VSS.t120 25.9346
R744 VSS.n1428 VSS.t61 25.9346
R745 VSS.n1044 VSS.t46 25.9346
R746 VSS.n1043 VSS.t108 25.9346
R747 VSS.n1027 VSS.t233 25.9346
R748 VSS.n1026 VSS.t227 25.9346
R749 VSS.n917 VSS.t68 25.9346
R750 VSS.n916 VSS.t159 25.9346
R751 VSS.n858 VSS.t103 25.9346
R752 VSS.n857 VSS.t116 25.9346
R753 VSS.n286 VSS.t112 25.9346
R754 VSS.n305 VSS.t177 25.9346
R755 VSS.n523 VSS.t57 25.9346
R756 VSS.n552 VSS.t20 25.9346
R757 VSS.n1439 VSS 21.9895
R758 VSS.t12 VSS 21.9895
R759 VSS.n2174 VSS.n2173 21.8894
R760 VSS.n1124 VSS.n1123 19.7906
R761 VSS.t136 VSS.n1271 19.7906
R762 VSS.t203 VSS.n1272 19.7906
R763 VSS.t60 VSS.n1443 19.7906
R764 VSS.n1889 VSS.n1888 19.7906
R765 VSS.t1 VSS.n1682 19.7906
R766 VSS.n1684 VSS.t187 19.7906
R767 VSS VSS.n2058 19.4706
R768 VSS.n1802 VSS.t125 17.5917
R769 VSS.n1090 VSS.n49 17.3181
R770 VSS.n2049 VSS.n19 17.3181
R771 VSS.n2020 VSS.n2019 17.3181
R772 VSS.n2002 VSS.n1201 17.3181
R773 VSS.n1343 VSS.n1342 17.3181
R774 VSS.n1948 VSS.n1351 17.3181
R775 VSS.n1915 VSS.n1395 17.3181
R776 VSS.n1892 VSS.n1891 17.3181
R777 VSS.n1891 VSS.n1474 17.3181
R778 VSS.n1617 VSS.n1609 17.3181
R779 VSS.n1628 VSS.n1609 17.3181
R780 VSS.n1629 VSS.n1628 17.3181
R781 VSS.n1799 VSS.n1739 17.3181
R782 VSS.n2020 VSS.n1152 17.1299
R783 VSS.n1092 VSS.n1090 16.9417
R784 VSS.n1434 VSS.n1431 16.9417
R785 VSS.n1702 VSS.n1669 16.7534
R786 VSS.n2019 VSS.n1183 16.5652
R787 VSS.n1083 VSS.n53 16.377
R788 VSS.n1514 VSS.n1513 16.377
R789 VSS.n1842 VSS.n1596 16.377
R790 VSS.n1915 VSS.n1394 16.1887
R791 VSS.n2049 VSS.n18 16.0005
R792 VSS.n1147 VSS.n19 16.0005
R793 VSS.n1268 VSS.n1206 16.0005
R794 VSS.n1514 VSS.n1470 16.0005
R795 VSS.n1785 VSS.n1781 15.8123
R796 VSS.n2060 VSS.n8 15.624
R797 VSS.n2039 VSS.n1148 15.4358
R798 VSS.n2003 VSS.n2002 15.4358
R799 VSS.n1892 VSS.n1471 15.4358
R800 VSS.n1057 VSS.n1054 15.3928
R801 VSS.n1622 VSS.n1621 15.3928
R802 VSS.n1447 VSS.n1446 15.2476
R803 VSS.n1680 VSS.n1679 15.0593
R804 VSS.n1436 VSS.n1388 15.0593
R805 VSS.n1921 VSS.n1388 15.0593
R806 VSS.n1921 VSS.n1920 15.0593
R807 VSS.n1901 VSS.n1464 15.0593
R808 VSS.n1480 VSS.n1464 15.0593
R809 VSS.n1886 VSS.n1480 15.0593
R810 VSS.n1623 VSS.n1588 15.0593
R811 VSS.n1847 VSS.n1588 15.0593
R812 VSS.n1847 VSS.n1589 15.0593
R813 VSS.n1826 VSS.n1665 15.0593
R814 VSS.n1804 VSS.n1665 15.0593
R815 VSS.n1804 VSS.n1733 15.0593
R816 VSS.n2031 VSS.n1157 15.0593
R817 VSS.n1189 VSS.n1157 15.0593
R818 VSS.n2013 VSS.n1189 15.0593
R819 VSS.n1997 VSS.n1274 15.0593
R820 VSS.n1976 VSS.n1274 15.0593
R821 VSS.n1976 VSS.n1302 15.0593
R822 VSS.n1120 VSS.n36 15.0593
R823 VSS.n1120 VSS.n23 15.0593
R824 VSS.n1142 VSS.n23 15.0593
R825 VSS.n1687 VSS.n1686 14.8711
R826 VSS.n1342 VSS.n1297 14.6829
R827 VSS.n1739 VSS.n1670 14.6829
R828 VSS.n1126 VSS.n31 14.4946
R829 VSS.n1128 VSS.n1127 14.4946
R830 VSS.n1505 VSS.n1395 14.4946
R831 VSS.n1446 VSS 14.3064
R832 VSS.n832 VSS.t53 14.24
R833 VSS.n1955 VSS.n1954 14.1181
R834 VSS.n435 VSS.t113 13.7077
R835 VSS.n506 VSS 13.7077
R836 VSS.n656 VSS.t33 13.7077
R837 VSS.n750 VSS 13.7077
R838 VSS.n1918 VSS.t121 13.1939
R839 VSS.n2150 VSS.n2149 13.1351
R840 VSS.t22 VSS.n2016 10.995
R841 VSS.n2015 VSS.n1188 10.995
R842 VSS.t182 VSS.n1188 10.995
R843 VSS.n1999 VSS.n1272 10.995
R844 VSS.n1621 VSS.t162 10.995
R845 VSS.n1781 VSS.n1740 10.7299
R846 VSS.n1954 VSS.n1344 10.7299
R847 VSS.n1948 VSS.n1344 10.7299
R848 VSS.n1799 VSS.n1740 10.7299
R849 VSS.n1617 VSS.n1616 9.97697
R850 VSS.n1296 VSS.n1201 9.6005
R851 VSS.n1128 VSS.n29 9.3005
R852 VSS.n1130 VSS.n1129 9.3005
R853 VSS.n2043 VSS.n2042 9.3005
R854 VSS.n2037 VSS.n1150 9.3005
R855 VSS.n1340 VSS.n1297 9.3005
R856 VSS.n1265 VSS.n1264 9.3005
R857 VSS.n1266 VSS.n1206 9.3005
R858 VSS.n1200 VSS.n1198 9.3005
R859 VSS.n1447 VSS.n1427 9.3005
R860 VSS.n1896 VSS.n1895 9.3005
R861 VSS.n1677 VSS.n1675 9.3005
R862 VSS.n9 VSS.n8 9.3005
R863 VSS.n1784 VSS.n1774 9.3005
R864 VSS.n1704 VSS.n1669 9.3005
R865 VSS.n1821 VSS.n1820 9.3005
R866 VSS.n1689 VSS.n1673 9.3005
R867 VSS.n1688 VSS.n1687 9.3005
R868 VSS.n1679 VSS.n1678 9.3005
R869 VSS.n1894 VSS.n1471 9.3005
R870 VSS.n1511 VSS.n1507 9.3005
R871 VSS.n1512 VSS.n1503 9.3005
R872 VSS.n1450 VSS.n1449 9.3005
R873 VSS.n1981 VSS.n1293 9.3005
R874 VSS.n2036 VSS.n1153 9.3005
R875 VSS.n1263 VSS.n1262 9.3005
R876 VSS.n2041 VSS.n1148 9.3005
R877 VSS.n47 VSS.n31 9.3005
R878 VSS.n1091 VSS.n48 9.3005
R879 VSS.n2167 VSS.n2166 9.3005
R880 VSS.n2165 VSS.n2164 9.3005
R881 VSS.n2179 VSS.n2178 9.3005
R882 VSS.n2178 VSS.n2177 9.3005
R883 VSS.n226 VSS.n225 9.15497
R884 VSS.n227 VSS.n226 9.15497
R885 VSS.n2113 VSS.n2112 9.15497
R886 VSS.n2112 VSS.n2111 9.15497
R887 VSS.n2066 VSS.n2065 9.15497
R888 VSS.n2065 VSS.n2064 9.15497
R889 VSS.n218 VSS.n217 9.15497
R890 VSS.n217 VSS.n216 9.15497
R891 VSS.n1666 VSS.n1665 9.15497
R892 VSS.n1735 VSS.n1666 9.15497
R893 VSS.n1804 VSS.n1803 9.15497
R894 VSS.n1803 VSS.n1802 9.15497
R895 VSS.n1734 VSS.n1733 9.15497
R896 VSS.n1737 VSS.n1734 9.15497
R897 VSS.n1826 VSS.n1825 9.15497
R898 VSS.n1825 VSS.n1824 9.15497
R899 VSS.n1590 VSS.n1588 9.15497
R900 VSS.n1622 VSS.n1590 9.15497
R901 VSS.n1847 VSS.n1846 9.15497
R902 VSS.n1846 VSS.n1845 9.15497
R903 VSS.n1591 VSS.n1589 9.15497
R904 VSS.n1592 VSS.n1591 9.15497
R905 VSS.n1624 VSS.n1623 9.15497
R906 VSS.n1625 VSS.n1624 9.15497
R907 VSS.n1465 VSS.n1464 9.15497
R908 VSS.n1467 VSS.n1465 9.15497
R909 VSS.n1480 VSS.n1479 9.15497
R910 VSS.n1479 VSS.n1478 9.15497
R911 VSS.n1887 VSS.n1886 9.15497
R912 VSS.n1888 VSS.n1887 9.15497
R913 VSS.n1901 VSS.n1900 9.15497
R914 VSS.n1900 VSS.n1899 9.15497
R915 VSS.n1921 VSS.n1389 9.15497
R916 VSS.n1443 VSS.n1389 9.15497
R917 VSS.n1920 VSS.n1919 9.15497
R918 VSS.n1919 VSS.n1918 9.15497
R919 VSS.n1440 VSS.n1436 9.15497
R920 VSS.n1440 VSS.n1439 9.15497
R921 VSS.n1441 VSS.n1388 9.15497
R922 VSS.n1442 VSS.n1441 9.15497
R923 VSS.n1274 VSS.n1273 9.15497
R924 VSS.n1299 VSS.n1273 9.15497
R925 VSS.n1977 VSS.n1976 9.15497
R926 VSS.n1978 VSS.n1977 9.15497
R927 VSS.n1302 VSS.n1301 9.15497
R928 VSS.n1348 VSS.n1301 9.15497
R929 VSS.n1998 VSS.n1997 9.15497
R930 VSS.n1999 VSS.n1998 9.15497
R931 VSS.n1189 VSS.n1187 9.15497
R932 VSS.n2016 VSS.n1187 9.15497
R933 VSS.n2014 VSS.n2013 9.15497
R934 VSS.n2015 VSS.n2014 9.15497
R935 VSS.n2032 VSS.n2031 9.15497
R936 VSS.n2033 VSS.n2032 9.15497
R937 VSS.n1157 VSS.n1156 9.15497
R938 VSS.n1186 VSS.n1156 9.15497
R939 VSS.n36 VSS.n35 9.15497
R940 VSS.n1087 VSS.n35 9.15497
R941 VSS.n1121 VSS.n1120 9.15497
R942 VSS.n1122 VSS.n1121 9.15497
R943 VSS.n23 VSS.n22 9.15497
R944 VSS.n1123 VSS.n22 9.15497
R945 VSS.n1143 VSS.n1142 9.15497
R946 VSS.n1144 VSS.n1143 9.15497
R947 VSS.n2138 VSS.n2137 9.01392
R948 VSS.n2137 VSS.n2136 9.01392
R949 VSS.n1629 VSS.n1595 8.84756
R950 VSS.n414 VSS.n411 8.84756
R951 VSS.n1701 VSS.n1700 8.65932
R952 VSS.n1268 VSS.n1205 8.47109
R953 VSS.n1842 VSS.n1595 8.47109
R954 VSS.n621 VSS.n618 8.47109
R955 VSS.n2149 VSS 7.93155
R956 VSS.n1702 VSS.n1701 7.71815
R957 VSS.n253 VSS.n250 7.71815
R958 VSS.n2171 VSS.n2170 7.52991
R959 VSS.n914 VSS 7.48358
R960 VSS.n2039 VSS.n2038 7.34168
R961 VSS.n1616 VSS.n1474 7.34168
R962 VSS.n377 VSS.n374 7.34168
R963 VSS.n608 VSS.n605 7.34168
R964 VSS.n1982 VSS.n1296 7.15344
R965 VSS.n119 VSS.t75 7.12024
R966 VSS.n911 VSS 7.12024
R967 VSS.n193 VSS.t214 7.12024
R968 VSS VSS.n755 7.12024
R969 VSS.n2038 VSS.n2037 6.96521
R970 VSS.n1145 VSS.n1144 6.5972
R971 VSS.t216 VSS.n1625 6.5972
R972 VSS.n1264 VSS.n1205 6.4005
R973 VSS.n680 VSS.n679 5.08285
R974 VSS.n279 VSS.n278 4.72342
R975 VSS.n1083 VSS.n1082 4.7104
R976 VSS.n1081 VSS.n49 4.6505
R977 VSS.n1090 VSS.n50 4.6505
R978 VSS.n1292 VSS.n1201 4.6505
R979 VSS.n1342 VSS.n1341 4.6505
R980 VSS.n1954 VSS.n1345 4.6505
R981 VSS.n1446 VSS.n1429 4.6505
R982 VSS.n1611 VSS.n1609 4.6505
R983 VSS.n1781 VSS.n1773 4.6505
R984 VSS.n2060 VSS.n2059 4.6505
R985 VSS.n1703 VSS.n1702 4.6505
R986 VSS.n1742 VSS.n1739 4.6505
R987 VSS.n1799 VSS.n1798 4.6505
R988 VSS.n1680 VSS.n1674 4.6505
R989 VSS.n1630 VSS.n1629 4.6505
R990 VSS.n1842 VSS.n1841 4.6505
R991 VSS.n1628 VSS.n1612 4.6505
R992 VSS.n1876 VSS.n1474 4.6505
R993 VSS.n1893 VSS.n1892 4.6505
R994 VSS.n1515 VSS.n1514 4.6505
R995 VSS.n1915 VSS.n1914 4.6505
R996 VSS.n1913 VSS.n1395 4.6505
R997 VSS.n1434 VSS.n1433 4.6505
R998 VSS.n1432 VSS.n1351 4.6505
R999 VSS.n1353 VSS.n1352 4.6505
R1000 VSS.n1343 VSS.n1338 4.6505
R1001 VSS.n2002 VSS.n1202 4.6505
R1002 VSS.n1268 VSS.n1267 4.6505
R1003 VSS.n2021 VSS.n2020 4.6505
R1004 VSS.n2019 VSS.n1182 4.6505
R1005 VSS.n2040 VSS.n2039 4.6505
R1006 VSS.n19 VSS.n17 4.6505
R1007 VSS.n2050 VSS.n2049 4.6505
R1008 VSS.n1126 VSS.n32 4.6505
R1009 VSS.n1060 VSS.n1059 4.6505
R1010 VSS.n1062 VSS.n1061 4.6505
R1011 VSS.n2151 VSS.n2150 4.6505
R1012 VSS.n283 VSS.n282 4.6505
R1013 VSS.n310 VSS.n309 4.6505
R1014 VSS.n338 VSS.n337 4.6505
R1015 VSS.n362 VSS.n361 4.6505
R1016 VSS.n378 VSS.n377 4.6505
R1017 VSS.n631 VSS.n630 4.6505
R1018 VSS.n622 VSS.n621 4.6505
R1019 VSS.n748 VSS.n747 4.6505
R1020 VSS.n739 VSS.n738 4.6505
R1021 VSS.n745 VSS.n744 4.6505
R1022 VSS.n711 VSS.n710 4.6505
R1023 VSS.n689 VSS.n688 4.6505
R1024 VSS.n675 VSS.n674 4.6505
R1025 VSS.n652 VSS.n651 4.6505
R1026 VSS.n442 VSS.n441 4.6505
R1027 VSS.n415 VSS.n414 4.6505
R1028 VSS.n402 VSS.n401 4.6505
R1029 VSS.n486 VSS.n485 4.6505
R1030 VSS.n502 VSS.n501 4.6505
R1031 VSS.n504 VSS.n503 4.6505
R1032 VSS.n613 VSS.n612 4.6505
R1033 VSS.n609 VSS.n608 4.6505
R1034 VSS.n593 VSS.n592 4.6505
R1035 VSS.n569 VSS.n568 4.6505
R1036 VSS.n557 VSS.n556 4.6505
R1037 VSS.n540 VSS.n539 4.6505
R1038 VSS.n528 VSS.n527 4.6505
R1039 VSS.n265 VSS.n264 4.6505
R1040 VSS.n254 VSS.n253 4.6505
R1041 VSS.n248 VSS.n247 4.6505
R1042 VSS.n627 VSS.n626 4.6505
R1043 VSS.n438 VSS.n437 4.6505
R1044 VSS.n961 VSS.n958 4.62819
R1045 VSS.n1068 VSS.n1067 4.5005
R1046 VSS.n1936 VSS.n1369 4.5005
R1047 VSS.n1386 VSS.n1373 4.5005
R1048 VSS.n1418 VSS.n1417 4.5005
R1049 VSS.n1924 VSS.n1923 4.5005
R1050 VSS.n1922 VSS.n1385 4.5005
R1051 VSS.n1416 VSS.n1415 4.5005
R1052 VSS.n1413 VSS.n1390 4.5005
R1053 VSS.n1933 VSS.n1370 4.5005
R1054 VSS.n1935 VSS.n1934 4.5005
R1055 VSS.n1529 VSS.n1528 4.5005
R1056 VSS.n1534 VSS.n1533 4.5005
R1057 VSS.n1532 VSS.n1531 4.5005
R1058 VSS.n1497 VSS.n1463 4.5005
R1059 VSS.n1550 VSS.n1549 4.5005
R1060 VSS.n1544 VSS.n1491 4.5005
R1061 VSS.n1547 VSS.n1490 4.5005
R1062 VSS.n1548 VSS.n1483 4.5005
R1063 VSS.n1902 VSS.n1462 4.5005
R1064 VSS.n1861 VSS.n1860 4.5005
R1065 VSS.n1859 VSS.n1575 4.5005
R1066 VSS.n1586 VSS.n1578 4.5005
R1067 VSS.n1863 VSS.n1862 4.5005
R1068 VSS.n1642 VSS.n1641 4.5005
R1069 VSS.n1850 VSS.n1849 4.5005
R1070 VSS.n1848 VSS.n1585 4.5005
R1071 VSS.n1653 VSS.n1639 4.5005
R1072 VSS.n1655 VSS.n1654 4.5005
R1073 VSS.n1717 VSS.n1716 4.5005
R1074 VSS.n1728 VSS.n1715 4.5005
R1075 VSS.n1730 VSS.n1729 4.5005
R1076 VSS.n1664 VSS.n1663 4.5005
R1077 VSS.n1750 VSS.n1732 4.5005
R1078 VSS.n1808 VSS.n1807 4.5005
R1079 VSS.n1805 VSS.n1731 4.5005
R1080 VSS.n1762 VSS.n1761 4.5005
R1081 VSS.n1828 VSS.n1827 4.5005
R1082 VSS.n1160 VSS.n1159 4.5005
R1083 VSS.n1220 VSS.n1219 4.5005
R1084 VSS.n1251 VSS.n1190 4.5005
R1085 VSS.n1243 VSS.n1242 4.5005
R1086 VSS.n1244 VSS.n1218 4.5005
R1087 VSS.n1245 VSS.n1214 4.5005
R1088 VSS.n2012 VSS.n1191 4.5005
R1089 VSS.n1228 VSS.n1225 4.5005
R1090 VSS.n1230 VSS.n1229 4.5005
R1091 VSS.n1317 VSS.n1277 4.5005
R1092 VSS.n1323 VSS.n1316 4.5005
R1093 VSS.n1325 VSS.n1324 4.5005
R1094 VSS.n1995 VSS.n1994 4.5005
R1095 VSS.n1974 VSS.n1973 4.5005
R1096 VSS.n1327 VSS.n1326 4.5005
R1097 VSS.n1975 VSS.n1304 4.5005
R1098 VSS.n1961 VSS.n1305 4.5005
R1099 VSS.n1996 VSS.n1276 4.5005
R1100 VSS.n1139 VSS.n24 4.5005
R1101 VSS.n71 VSS.n70 4.5005
R1102 VSS.n40 VSS.n39 4.5005
R1103 VSS.n58 VSS.n37 4.5005
R1104 VSS.n1119 VSS.n38 4.5005
R1105 VSS.n1104 VSS.n1103 4.5005
R1106 VSS.n1109 VSS.n1108 4.5005
R1107 VSS.n1107 VSS.n1102 4.5005
R1108 VSS.n1141 VSS.n1140 4.5005
R1109 VSS.n2058 VSS.n2057 4.5005
R1110 VSS.n1819 VSS.n1818 4.5005
R1111 VSS.n1819 VSS.n1670 4.5005
R1112 VSS.n1741 VSS.n1707 4.5005
R1113 VSS.n1840 VSS.n1839 4.5005
R1114 VSS.n1676 VSS.n1633 4.5005
R1115 VSS.n1676 VSS.n1596 4.5005
R1116 VSS.n1875 VSS.n1874 4.5005
R1117 VSS.n1873 VSS.n1563 4.5005
R1118 VSS.n1610 VSS.n1566 4.5005
R1119 VSS.n1180 VSS.n1179 4.5005
R1120 VSS.n1180 VSS.n1152 4.5005
R1121 VSS.n2023 VSS.n2022 4.5005
R1122 VSS.n1132 VSS.n1131 4.5005
R1123 VSS.n1131 VSS.n18 4.5005
R1124 VSS.n2052 VSS.n2051 4.5005
R1125 VSS.n62 VSS.n61 4.5005
R1126 VSS.n1094 VSS.n1093 4.5005
R1127 VSS.n1093 VSS.n1092 4.5005
R1128 VSS.n1358 VSS.n1354 4.5005
R1129 VSS.n1947 VSS.n1355 4.5005
R1130 VSS.n1357 VSS.n1356 4.5005
R1131 VSS.n1361 VSS.n1360 4.5005
R1132 VSS.n1957 VSS.n1956 4.5005
R1133 VSS.n1956 VSS.n1955 4.5005
R1134 VSS.n1983 VSS.n1294 4.5005
R1135 VSS.n1983 VSS.n1982 4.5005
R1136 VSS.n1986 VSS.n1985 4.5005
R1137 VSS.n2005 VSS.n2004 4.5005
R1138 VSS.n2004 VSS.n2003 4.5005
R1139 VSS.n1284 VSS.n1283 4.5005
R1140 VSS.n1210 VSS.n1209 4.5005
R1141 VSS.n1454 VSS.n1396 4.5005
R1142 VSS.n1912 VSS.n1911 4.5005
R1143 VSS.n1506 VSS.n1399 4.5005
R1144 VSS.n1506 VSS.n1505 4.5005
R1145 VSS.n1516 VSS.n1502 4.5005
R1146 VSS.n1559 VSS.n1473 4.5005
R1147 VSS.n1562 VSS.n1475 4.5005
R1148 VSS.n1699 VSS.n1698 4.5005
R1149 VSS.n1700 VSS.n1699 4.5005
R1150 VSS.n1770 VSS.n1745 4.5005
R1151 VSS.n1789 VSS.n1788 4.5005
R1152 VSS.n1786 VSS.n1776 4.5005
R1153 VSS.n1786 VSS.n1785 4.5005
R1154 VSS.n1692 VSS.n1671 4.5005
R1155 VSS.n1797 VSS.n1796 4.5005
R1156 VSS.n1878 VSS.n1877 4.5005
R1157 VSS.n1518 VSS.n1472 4.5005
R1158 VSS.n1472 VSS.n1470 4.5005
R1159 VSS.n1451 VSS.n1426 4.5005
R1160 VSS.n1451 VSS.n1394 4.5005
R1161 VSS.n1261 VSS.n1260 4.5005
R1162 VSS.n1261 VSS.n1183 4.5005
R1163 VSS.n1170 VSS.n1169 4.5005
R1164 VSS.n1173 VSS.n1149 4.5005
R1165 VSS.n1149 VSS.n1147 4.5005
R1166 VSS VSS.n2145 4.5005
R1167 VSS.n2181 VSS.n2180 4.5005
R1168 VSS.n707 VSS.n706 4.5005
R1169 VSS.n685 VSS.n684 4.5005
R1170 VSS.n293 VSS.n292 4.5005
R1171 VSS.n334 VSS.n333 4.5005
R1172 VSS.n387 VSS.n386 4.5005
R1173 VSS.n661 VSS.n660 4.5005
R1174 VSS.n434 VSS.n433 4.5005
R1175 VSS.n410 VSS.n409 4.5005
R1176 VSS.n494 VSS.n493 4.5005
R1177 VSS.n601 VSS.n600 4.5005
R1178 VSS.n565 VSS.n564 4.5005
R1179 VSS.n536 VSS.n535 4.5005
R1180 VSS.n512 VSS.n511 4.5005
R1181 VSS.n358 VSS.n357 4.5005
R1182 VSS.n814 VSS.n811 4.43127
R1183 VSS.n2017 VSS.t22 4.3983
R1184 VSS.n1626 VSS.t216 4.3983
R1185 VSS.n150 VSS.n147 4.03742
R1186 VSS.n794 VSS.n791 4.03742
R1187 VSS.n112 VSS.n109 3.8405
R1188 VSS.n182 VSS.n179 3.8405
R1189 VSS.n2180 VSS.n2169 3.76521
R1190 VSS.n1080 VSS.n54 3.46971
R1191 VSS.n1607 VSS.n1597 3.46971
R1192 VSS.n1362 VSS.n1361 3.46752
R1193 VSS.n1911 VSS.n1398 3.46532
R1194 VSS.n81 VSS.n80 3.46323
R1195 VSS.n1070 VSS.n1069 3.46321
R1196 VSS.n1169 VSS.n1168 3.46272
R1197 VSS.n1815 VSS.n1707 3.46094
R1198 VSS.n2138 VSS.n2132 3.45447
R1199 VSS.n1411 VSS.n1402 3.45291
R1200 VSS.n1657 VSS.n1656 3.45291
R1201 VSS.n2011 VSS.n2010 3.45291
R1202 VSS.n1285 VSS.n1284 3.45217
R1203 VSS.n1904 VSS.n1903 3.45156
R1204 VSS.n1662 VSS.n1658 3.45156
R1205 VSS.n1279 VSS.n1275 3.45156
R1206 VSS.n1502 VSS.n1500 3.44997
R1207 VSS.n1179 VSS.n1178 3.44997
R1208 VSS.n1790 VSS.n1789 3.44997
R1209 VSS.n2053 VSS.n2052 3.44778
R1210 VSS.n1455 VSS.n1454 3.44559
R1211 VSS.n1839 VSS.n1632 3.44559
R1212 VSS.n1776 VSS.n1775 3.44457
R1213 VSS.n1095 VSS.n1094 3.44339
R1214 VSS.n1693 VSS.n1692 3.44339
R1215 VSS.n1746 VSS.n1745 3.44339
R1216 VSS.n1987 VSS.n1986 3.4412
R1217 VSS.n1309 VSS.n1294 3.4412
R1218 VSS.n1211 VSS.n1210 3.4412
R1219 VSS.n1260 VSS.n1259 3.4412
R1220 VSS.n1940 VSS.n1939 3.43949
R1221 VSS.n1884 VSS.n1482 3.43949
R1222 VSS.n1866 VSS.n1865 3.43949
R1223 VSS.n1766 VSS.n1765 3.43949
R1224 VSS.n1161 VSS.n1158 3.43949
R1225 VSS.n1965 VSS.n1964 3.43949
R1226 VSS.n75 VSS.n74 3.43943
R1227 VSS.n63 VSS.n62 3.43901
R1228 VSS.n1698 VSS.n1691 3.43901
R1229 VSS.n1796 VSS.n1744 3.43901
R1230 VSS.n1067 VSS.n1063 3.43687
R1231 VSS.n1426 VSS.n1425 3.43682
R1232 VSS.n1634 VSS.n1633 3.43682
R1233 VSS.n1133 VSS.n1132 3.43462
R1234 VSS.n1518 VSS.n1501 3.43243
R1235 VSS.n2024 VSS.n2023 3.43243
R1236 VSS.n1174 VSS.n1173 3.43243
R1237 VSS.n2006 VSS.n2005 3.43024
R1238 VSS.n1606 VSS.n1581 3.42639
R1239 VSS.n1559 VSS.n1558 3.42585
R1240 VSS.n1567 VSS.n1566 3.42585
R1241 VSS.n1079 VSS.n77 3.42429
R1242 VSS.n1943 VSS.n1357 3.42366
R1243 VSS.n2057 VSS.n2056 3.42153
R1244 VSS.n1359 VSS.n1358 3.42146
R1245 VSS.n1818 VSS.n1706 3.42146
R1246 VSS.n1879 VSS.n1878 3.41927
R1247 VSS.n1874 VSS.n1564 3.41927
R1248 VSS.n1908 VSS.n1399 3.41708
R1249 VSS.n1958 VSS.n1957 3.41489
R1250 VSS.n1941 VSS.n1940 3.41257
R1251 VSS.n1767 VSS.n1766 3.41257
R1252 VSS.n1176 VSS.n1161 3.41257
R1253 VSS.n1966 VSS.n1965 3.41257
R1254 VSS.n76 VSS.n75 3.41257
R1255 VSS.n2056 VSS.n2055 3.41257
R1256 VSS.n1071 VSS.n1070 3.41218
R1257 VSS.n81 VSS.n78 3.41218
R1258 VSS.n1076 VSS.n54 3.41212
R1259 VSS.n64 VSS.n63 3.41212
R1260 VSS.n1096 VSS.n1095 3.41212
R1261 VSS.n1134 VSS.n1133 3.41212
R1262 VSS.n2054 VSS.n2053 3.41212
R1263 VSS.n1694 VSS.n1691 3.41212
R1264 VSS.n1693 VSS.n1659 3.41212
R1265 VSS.n1558 VSS.n1557 3.41212
R1266 VSS.n1880 VSS.n1879 3.41212
R1267 VSS.n1500 VSS.n1401 3.41212
R1268 VSS.n1501 VSS.n1494 3.41212
R1269 VSS.n1457 VSS.n1398 3.41212
R1270 VSS.n1908 VSS.n1907 3.41212
R1271 VSS.n1425 VSS.n1424 3.41212
R1272 VSS.n1456 VSS.n1455 3.41212
R1273 VSS.n1364 VSS.n1359 3.41212
R1274 VSS.n1943 VSS.n1942 3.41212
R1275 VSS.n1598 VSS.n1597 3.41212
R1276 VSS.n1648 VSS.n1632 3.41212
R1277 VSS.n1636 VSS.n1634 3.41212
R1278 VSS.n1747 VSS.n1744 3.41212
R1279 VSS.n1792 VSS.n1746 3.41212
R1280 VSS.n1568 VSS.n1564 3.41212
R1281 VSS.n1869 VSS.n1567 3.41212
R1282 VSS.n1959 VSS.n1958 3.41212
R1283 VSS.n1363 VSS.n1362 3.41212
R1284 VSS.n1988 VSS.n1987 3.41212
R1285 VSS.n1310 VSS.n1309 3.41212
R1286 VSS.n2007 VSS.n2006 3.41212
R1287 VSS.n1286 VSS.n1285 3.41212
R1288 VSS.n1178 VSS.n1177 3.41212
R1289 VSS.n2025 VSS.n2024 3.41212
R1290 VSS.n1212 VSS.n1211 3.41212
R1291 VSS.n1259 VSS.n1195 3.41212
R1292 VSS.n1791 VSS.n1790 3.41212
R1293 VSS.n1720 VSS.n1706 3.41212
R1294 VSS.n1815 VSS.n1814 3.41212
R1295 VSS.n1175 VSS.n1174 3.41212
R1296 VSS.n1723 VSS.n1661 3.4105
R1297 VSS.n1713 VSS.n1711 3.4105
R1298 VSS.n1752 VSS.n1751 3.4105
R1299 VSS.n1810 VSS.n1809 3.4105
R1300 VSS.n1760 VSS.n1759 3.4105
R1301 VSS.n1725 VSS.n1724 3.4105
R1302 VSS.n1600 VSS.n1574 3.4105
R1303 VSS.n1584 VSS.n1580 3.4105
R1304 VSS.n1644 VSS.n1643 3.4105
R1305 VSS.n1852 VSS.n1851 3.4105
R1306 VSS.n1652 VSS.n1651 3.4105
R1307 VSS.n1579 VSS.n1576 3.4105
R1308 VSS.n1526 VSS.n1525 3.4105
R1309 VSS.n1496 VSS.n1492 3.4105
R1310 VSS.n1553 VSS.n1552 3.4105
R1311 VSS.n1543 VSS.n1542 3.4105
R1312 VSS.n1551 VSS.n1484 3.4105
R1313 VSS.n1527 VSS.n1495 3.4105
R1314 VSS.n1374 VSS.n1371 3.4105
R1315 VSS.n1384 VSS.n1375 3.4105
R1316 VSS.n1378 VSS.n1377 3.4105
R1317 VSS.n1410 VSS.n1408 3.4105
R1318 VSS.n1926 VSS.n1925 3.4105
R1319 VSS.n1420 VSS.n1419 3.4105
R1320 VSS.n1993 VSS.n1992 3.4105
R1321 VSS.n1320 VSS.n1314 3.4105
R1322 VSS.n1972 VSS.n1971 3.4105
R1323 VSS.n1329 VSS.n1328 3.4105
R1324 VSS.n1333 VSS.n1306 3.4105
R1325 VSS.n1319 VSS.n1278 3.4105
R1326 VSS.n1232 VSS.n1231 3.4105
R1327 VSS.n1240 VSS.n1239 3.4105
R1328 VSS.n1224 VSS.n1162 3.4105
R1329 VSS.n1250 VSS.n1249 3.4105
R1330 VSS.n1241 VSS.n1215 3.4105
R1331 VSS.n1253 VSS.n1252 3.4105
R1332 VSS.n1223 VSS.n1164 3.4105
R1333 VSS.n1991 VSS.n1990 3.4105
R1334 VSS.n1970 VSS.n1969 3.4105
R1335 VSS.n1331 VSS.n1330 3.4105
R1336 VSS.n1968 VSS.n1308 3.4105
R1337 VSS.n1313 VSS.n1312 3.4105
R1338 VSS.n1989 VSS.n1282 3.4105
R1339 VSS.n1287 VSS.n1194 3.4105
R1340 VSS.n1238 VSS.n1237 3.4105
R1341 VSS.n1216 VSS.n1213 3.4105
R1342 VSS.n1236 VSS.n1222 3.4105
R1343 VSS.n2009 VSS.n2008 3.4105
R1344 VSS.n1255 VSS.n1254 3.4105
R1345 VSS.n1234 VSS.n1233 3.4105
R1346 VSS.n1379 VSS.n1376 3.4105
R1347 VSS.n1719 VSS.n1660 3.4105
R1348 VSS.n1755 VSS.n1753 3.4105
R1349 VSS.n1811 VSS.n1710 3.4105
R1350 VSS.n1758 VSS.n1757 3.4105
R1351 VSS.n1813 VSS.n1812 3.4105
R1352 VSS.n1722 VSS.n1721 3.4105
R1353 VSS.n1833 VSS.n1832 3.4105
R1354 VSS.n1601 VSS.n1599 3.4105
R1355 VSS.n1647 VSS.n1645 3.4105
R1356 VSS.n1853 VSS.n1582 3.4105
R1357 VSS.n1835 VSS.n1834 3.4105
R1358 VSS.n1650 VSS.n1649 3.4105
R1359 VSS.n1855 VSS.n1854 3.4105
R1360 VSS.n1603 VSS.n1602 3.4105
R1361 VSS.n1868 VSS.n1867 3.4105
R1362 VSS.n1524 VSS.n1523 3.4105
R1363 VSS.n1554 VSS.n1488 3.4105
R1364 VSS.n1541 VSS.n1540 3.4105
R1365 VSS.n1570 VSS.n1486 3.4105
R1366 VSS.n1556 VSS.n1555 3.4105
R1367 VSS.n1538 VSS.n1493 3.4105
R1368 VSS.n1522 VSS.n1498 3.4105
R1369 VSS.n1906 VSS.n1905 3.4105
R1370 VSS.n1929 VSS.n1928 3.4105
R1371 VSS.n1423 VSS.n1422 3.4105
R1372 VSS.n1927 VSS.n1382 3.4105
R1373 VSS.n1459 VSS.n1458 3.4105
R1374 VSS.n1421 VSS.n1407 3.4105
R1375 VSS.n1381 VSS.n1380 3.4105
R1376 VSS.n1138 VSS.n1137 3.4105
R1377 VSS.n69 VSS.n68 3.4105
R1378 VSS.n1098 VSS.n25 3.4105
R1379 VSS.n1111 VSS.n1110 3.4105
R1380 VSS.n1101 VSS.n42 3.4105
R1381 VSS.n59 VSS.n41 3.4105
R1382 VSS.n27 VSS.n26 3.4105
R1383 VSS.n1112 VSS.n1097 3.4105
R1384 VSS.n1114 VSS.n1113 3.4105
R1385 VSS.n60 VSS.n43 3.4105
R1386 VSS.n67 VSS.n66 3.4105
R1387 VSS.n1136 VSS.n1135 3.4105
R1388 VSS.n1074 VSS.n1073 3.4105
R1389 VSS.n1075 VSS.n1074 3.4105
R1390 VSS.n2172 VSS.n2171 3.38874
R1391 VSS.n2139 VSS.n2131 3.25129
R1392 VSS.n84 VSS.n82 3.22773
R1393 VSS.n1955 VSS.n1343 3.2005
R1394 VSS.n1072 VSS 3.19575
R1395 VSS.n231 VSS.n230 3.10907
R1396 VSS.n1771 VSS.n1740 3.10907
R1397 VSS.n1352 VSS.n1344 3.10907
R1398 VSS.n1061 VSS 3.10907
R1399 VSS.n485 VSS.n484 3.10907
R1400 VSS.n1042 VSS.n997 3.10177
R1401 VSS.n1436 VSS.n1368 3.03311
R1402 VSS.n1533 VSS.n1464 3.03311
R1403 VSS.n1588 VSS.n1575 3.03311
R1404 VSS.n1715 VSS.n1665 3.03311
R1405 VSS.n2031 VSS.n2030 3.03311
R1406 VSS.n1316 VSS.n1274 3.03311
R1407 VSS.n57 VSS.n36 3.03311
R1408 VSS.n1948 VSS.n1947 3.03311
R1409 VSS.n1617 VSS.n1563 3.03311
R1410 VSS.n1891 VSS.n1475 3.03311
R1411 VSS.n225 VSS.n224 3.03311
R1412 VSS.n2140 VSS.n2139 3.03311
R1413 VSS.n2114 VSS.n2113 3.03311
R1414 VSS.n2067 VSS.n2066 3.03311
R1415 VSS.n219 VSS.n218 3.03311
R1416 VSS.n1805 VSS.n1804 3.03311
R1417 VSS.n1749 VSS.n1733 3.03311
R1418 VSS.n1827 VSS.n1826 3.03311
R1419 VSS.n1848 VSS.n1847 3.03311
R1420 VSS.n1655 VSS.n1589 3.03311
R1421 VSS.n1623 VSS.n1572 3.03311
R1422 VSS.n1547 VSS.n1480 3.03311
R1423 VSS.n1886 VSS.n1885 3.03311
R1424 VSS.n1902 VSS.n1901 3.03311
R1425 VSS.n1922 VSS.n1921 3.03311
R1426 VSS.n1920 VSS.n1390 3.03311
R1427 VSS.n1388 VSS.n1370 3.03311
R1428 VSS.n1976 VSS.n1975 3.03311
R1429 VSS.n1960 VSS.n1302 3.03311
R1430 VSS.n1997 VSS.n1996 3.03311
R1431 VSS.n1244 VSS.n1189 3.03311
R1432 VSS.n2013 VSS.n2012 3.03311
R1433 VSS.n1228 VSS.n1157 3.03311
R1434 VSS.n1120 VSS.n1119 3.03311
R1435 VSS.n1107 VSS.n23 3.03311
R1436 VSS.n1142 VSS.n1141 3.03311
R1437 VSS.n315 VSS.n314 3.03311
R1438 VSS.n480 VSS.n269 3.03311
R1439 VSS.n633 VSS.n617 3.03311
R1440 VSS.n259 VSS.n258 3.03311
R1441 VSS.n2060 VSS 3.01226
R1442 VSS.n2037 VSS.n2036 3.01226
R1443 VSS.n1434 VSS 3.01226
R1444 VSS.n2179 VSS.n2172 3.01226
R1445 VSS.n357 VSS.n356 3.01226
R1446 VSS.n84 VSS.n83 2.98487
R1447 VSS.n1091 VSS.n31 2.82403
R1448 VSS.n1511 VSS.n1505 2.82403
R1449 VSS.n385 VSS.n384 2.82403
R1450 VSS.n1981 VSS.n1297 2.63579
R1451 VSS.n1821 VSS.n1670 2.63579
R1452 VSS.n683 VSS.n680 2.63579
R1453 VSS.n1264 VSS.n1263 2.44756
R1454 VSS.n408 VSS.n405 2.44756
R1455 VSS.n493 VSS.n492 2.44756
R1456 VSS.n1050 VSS.n1049 2.3854
R1457 VSS.n1049 VSS.n1048 2.3255
R1458 VSS.n1041 VSS.n1040 2.3255
R1459 VSS.n1037 VSS.n1036 2.3255
R1460 VSS.n1032 VSS.n1031 2.3255
R1461 VSS.n1025 VSS.n1024 2.3255
R1462 VSS.n1018 VSS.n1017 2.3255
R1463 VSS.n1011 VSS.n1010 2.3255
R1464 VSS.n1006 VSS.n1005 2.3255
R1465 VSS.n113 VSS.n112 2.3255
R1466 VSS.n118 VSS.n117 2.3255
R1467 VSS.n127 VSS.n126 2.3255
R1468 VSS.n123 VSS.n122 2.3255
R1469 VSS.n968 VSS.n967 2.3255
R1470 VSS.n972 VSS.n971 2.3255
R1471 VSS.n976 VSS.n975 2.3255
R1472 VSS.n144 VSS.n143 2.3255
R1473 VSS.n151 VSS.n150 2.3255
R1474 VSS.n937 VSS.n936 2.3255
R1475 VSS.n941 VSS.n940 2.3255
R1476 VSS.n945 VSS.n944 2.3255
R1477 VSS.n893 VSS.n892 2.3255
R1478 VSS.n900 VSS.n899 2.3255
R1479 VSS.n907 VSS.n906 2.3255
R1480 VSS.n909 VSS.n908 2.3255
R1481 VSS.n915 VSS.n914 2.3255
R1482 VSS.n922 VSS.n921 2.3255
R1483 VSS.n877 VSS.n876 2.3255
R1484 VSS.n881 VSS.n880 2.3255
R1485 VSS.n861 VSS.n860 2.3255
R1486 VSS.n865 VSS.n864 2.3255
R1487 VSS.n162 VSS.n161 2.3255
R1488 VSS.n166 VSS.n165 2.3255
R1489 VSS.n171 VSS.n170 2.3255
R1490 VSS.n183 VSS.n182 2.3255
R1491 VSS.n187 VSS.n186 2.3255
R1492 VSS.n831 VSS.n830 2.3255
R1493 VSS.n835 VSS.n834 2.3255
R1494 VSS.n839 VSS.n838 2.3255
R1495 VSS.n815 VSS.n814 2.3255
R1496 VSS.n819 VSS.n818 2.3255
R1497 VSS.n196 VSS.n195 2.3255
R1498 VSS.n200 VSS.n199 2.3255
R1499 VSS.n795 VSS.n794 2.3255
R1500 VSS.n799 VSS.n798 2.3255
R1501 VSS.n772 VSS.n771 2.3255
R1502 VSS.n776 VSS.n775 2.3255
R1503 VSS.n780 VSS.n779 2.3255
R1504 VSS.n209 VSS.n208 2.3255
R1505 VSS.n759 VSS.n758 2.3255
R1506 VSS.n753 VSS.n210 2.3255
R1507 VSS.n1772 VSS.n1771 2.28373
R1508 VSS.n232 VSS.n231 2.28323
R1509 VSS.n1679 VSS.n1675 2.25932
R1510 VSS.n1687 VSS.n1673 2.25932
R1511 VSS.n510 VSS.n509 2.25932
R1512 VSS.n535 VSS.n534 2.25932
R1513 VSS.n564 VSS.n563 2.25932
R1514 VSS.n1939 VSS.n1368 2.251
R1515 VSS.n1885 VSS.n1884 2.251
R1516 VSS.n1865 VSS.n1572 2.251
R1517 VSS.n1765 VSS.n1749 2.251
R1518 VSS.n2030 VSS.n1158 2.251
R1519 VSS.n1964 VSS.n1960 2.251
R1520 VSS.n74 VSS.n57 2.24363
R1521 VSS.n2200 VSS.n2199 2.24031
R1522 VSS.n2000 VSS.t184 2.1994
R1523 VSS VSS.n1438 2.1994
R1524 VSS.t44 VSS.t73 2.1994
R1525 VSS.n2062 VSS 2.1994
R1526 VSS.n433 VSS.n432 2.07109
R1527 VSS.n600 VSS.n599 2.07109
R1528 VSS.n659 VSS.n658 2.07109
R1529 VSS.n2201 VSS 1.94963
R1530 VSS.n1082 VSS.n1080 1.94045
R1531 VSS.n1608 VSS.n1607 1.94045
R1532 VSS.n801 VSS.n800 1.94045
R1533 VSS.n761 VSS.n760 1.94045
R1534 VSS.n841 VSS.n840 1.94045
R1535 VSS.n821 VSS.n820 1.94045
R1536 VSS.n867 VSS.n866 1.94045
R1537 VSS.n883 VSS.n882 1.94045
R1538 VSS.n924 VSS.n923 1.94045
R1539 VSS.n896 VSS.n895 1.94045
R1540 VSS.n947 VSS.n946 1.94045
R1541 VSS.n978 VSS.n977 1.94045
R1542 VSS.n153 VSS.n152 1.94045
R1543 VSS.n129 VSS.n128 1.94045
R1544 VSS.n173 VSS.n172 1.94045
R1545 VSS.n189 VSS.n188 1.94045
R1546 VSS.n202 VSS.n201 1.94045
R1547 VSS.n782 VSS.n781 1.94045
R1548 VSS.n1129 VSS.n1128 1.88285
R1549 VSS.n2043 VSS.n1148 1.88285
R1550 VSS.n2003 VSS.n1200 1.88285
R1551 VSS.n1896 VSS.n1471 1.88285
R1552 VSS.n333 VSS.n332 1.69462
R1553 VSS.n705 VSS.n702 1.69462
R1554 VSS.n909 VSS 1.57588
R1555 VSS.n753 VSS 1.57588
R1556 VSS.n962 VSS.n961 1.53347
R1557 VSS.n1785 VSS.n1784 1.50638
R1558 VSS.n2180 VSS.n2179 1.50638
R1559 VSS.n332 VSS.n329 1.50638
R1560 VSS.n706 VSS.n705 1.50638
R1561 VSS.n1017 VSS.n1014 1.47742
R1562 VSS.n73 VSS.n72 1.35607
R1563 VSS.n1697 VSS.n1690 1.35607
R1564 VSS.n1453 VSS.n1452 1.35607
R1565 VSS.n1199 VSS.n1197 1.35607
R1566 VSS.n1208 VSS.n1207 1.35607
R1567 VSS.n1181 VSS.n1166 1.35607
R1568 VSS.n1519 VSS.n1517 1.35607
R1569 VSS.n1872 VSS.n1565 1.35607
R1570 VSS.n1838 VSS.n1631 1.35607
R1571 VSS.n1795 VSS.n1743 1.35607
R1572 VSS.n1787 VSS.n1769 1.35607
R1573 VSS.n1984 VSS.n1291 1.35607
R1574 VSS.n46 VSS.n45 1.35607
R1575 VSS.n16 VSS.n15 1.35607
R1576 VSS.n1172 VSS.n1171 1.35607
R1577 VSS.n2186 VSS.n2185 1.35607
R1578 VSS.n2162 VSS.n2161 1.35607
R1579 VSS.n514 VSS.n513 1.35607
R1580 VSS.n543 VSS.n542 1.35607
R1581 VSS.n572 VSS.n571 1.35607
R1582 VSS.n365 VSS.n364 1.35607
R1583 VSS.n418 VSS.n417 1.35607
R1584 VSS.n445 VSS.n444 1.35607
R1585 VSS.n664 VSS.n662 1.35607
R1586 VSS.n390 VSS.n388 1.35607
R1587 VSS.n342 VSS.n340 1.35607
R1588 VSS.n319 VSS.n316 1.35607
R1589 VSS.n296 VSS.n294 1.35607
R1590 VSS.n693 VSS.n691 1.35607
R1591 VSS.n1806 VSS.n1714 1.35607
R1592 VSS.n1764 VSS.n1763 1.35607
R1593 VSS.n1727 VSS.n1718 1.35607
R1594 VSS.n1864 VSS.n1573 1.35607
R1595 VSS.n1640 VSS.n1587 1.35607
R1596 VSS.n1858 VSS.n1577 1.35607
R1597 VSS.n1546 VSS.n1545 1.35607
R1598 VSS.n1883 VSS.n1481 1.35607
R1599 VSS.n1535 VSS.n1530 1.35607
R1600 VSS.n1932 VSS.n1372 1.35607
R1601 VSS.n1414 VSS.n1387 1.35607
R1602 VSS.n1938 VSS.n1937 1.35607
R1603 VSS.n1315 VSS.n1303 1.35607
R1604 VSS.n1963 VSS.n1962 1.35607
R1605 VSS.n1322 VSS.n1318 1.35607
R1606 VSS.n1227 VSS.n1226 1.35607
R1607 VSS.n1247 VSS.n1246 1.35607
R1608 VSS.n2029 VSS.n2028 1.35607
R1609 VSS.n1106 VSS.n1105 1.35607
R1610 VSS.n1118 VSS.n1117 1.35607
R1611 VSS.n11 VSS.n10 1.35607
R1612 VSS.n1561 VSS.n1560 1.35607
R1613 VSS.n1910 VSS.n1397 1.35607
R1614 VSS.n1946 VSS.n1945 1.35607
R1615 VSS.n1339 VSS.n1337 1.35607
R1616 VSS.n1817 VSS.n1705 1.35607
R1617 VSS.n2117 VSS.n2115 1.35607
R1618 VSS.n2154 VSS.n2153 1.35607
R1619 VSS.n734 VSS.n733 1.35607
R1620 VSS.n715 VSS.n713 1.35607
R1621 VSS.n1783 VSS.n8 1.31815
R1622 VSS.n1129 VSS.n18 1.31815
R1623 VSS.n2043 VSS.n1147 1.31815
R1624 VSS.n1206 VSS.n1200 1.31815
R1625 VSS.n1896 VSS.n1470 1.31815
R1626 VSS.n290 VSS.n289 1.31815
R1627 VSS.n1059 VSS.n86 1.2805
R1628 VSS.n1005 VSS.n1001 1.2805
R1629 VSS.n79 VSS.n78 1.13981
R1630 VSS.n1448 VSS.n1447 1.12991
R1631 VSS.n1449 VSS.n1394 1.12991
R1632 VSS.n432 VSS.n429 1.12991
R1633 VSS.n599 VSS.n596 1.12991
R1634 VSS.n660 VSS.n659 1.12991
R1635 VSS.n634 VSS.n633 1.04225
R1636 VSS.n480 VSS.n479 1.04225
R1637 VSS.n1411 VSS.n1390 1.04008
R1638 VSS.n1656 VSS.n1655 1.04008
R1639 VSS.n2012 VSS.n2011 1.04008
R1640 VSS.n1903 VSS.n1902 1.03985
R1641 VSS.n1827 VSS.n1662 1.03985
R1642 VSS.n1996 VSS.n1275 1.03985
R1643 VSS.n2068 VSS.n2067 1.03985
R1644 VSS.n53 VSS.n49 0.941676
R1645 VSS.n1127 VSS.n1126 0.941676
R1646 VSS.n1449 VSS.n1448 0.941676
R1647 VSS.n1675 VSS.n1596 0.941676
R1648 VSS.n1700 VSS.n1673 0.941676
R1649 VSS.n292 VSS.n291 0.941676
R1650 VSS.n291 VSS.n290 0.941676
R1651 VSS.n309 VSS.n306 0.941676
R1652 VSS.n511 VSS.n510 0.941676
R1653 VSS.n527 VSS.n524 0.941676
R1654 VSS.n534 VSS.n531 0.941676
R1655 VSS.n556 VSS.n553 0.941676
R1656 VSS.n563 VSS.n560 0.941676
R1657 VSS.n1060 VSS.n84 0.935851
R1658 VSS.n472 VSS.n471 0.853
R1659 VSS.n733 VSS.n731 0.853
R1660 VSS.n665 VSS.n664 0.853
R1661 VSS.n391 VSS.n390 0.853
R1662 VSS.n343 VSS.n342 0.853
R1663 VSS.n320 VSS.n319 0.853
R1664 VSS.n297 VSS.n296 0.853
R1665 VSS.n446 VSS.n445 0.853
R1666 VSS.n419 VSS.n418 0.853
R1667 VSS.n366 VSS.n365 0.853
R1668 VSS.n463 VSS.n462 0.853
R1669 VSS.n635 VSS.n634 0.853
R1670 VSS.n582 VSS.n581 0.853
R1671 VSS.n573 VSS.n572 0.853
R1672 VSS.n544 VSS.n543 0.853
R1673 VSS.n515 VSS.n514 0.853
R1674 VSS.n694 VSS.n693 0.853
R1675 VSS.n1065 VSS.n1064 0.853
R1676 VSS.n45 VSS.n44 0.853
R1677 VSS.n15 VSS.n14 0.853
R1678 VSS.n1697 VSS.n1696 0.853
R1679 VSS.n1520 VSS.n1519 0.853
R1680 VSS.n1453 VSS.n1404 0.853
R1681 VSS.n1838 VSS.n1837 0.853
R1682 VSS.n1795 VSS.n1794 0.853
R1683 VSS.n1872 VSS.n1871 0.853
R1684 VSS.n1764 VSS.n1748 0.853
R1685 VSS.n1291 VSS.n1290 0.853
R1686 VSS.n1197 VSS.n1196 0.853
R1687 VSS.n1166 VSS.n1165 0.853
R1688 VSS.n1258 VSS.n1208 0.853
R1689 VSS.n1963 VSS.n1334 0.853
R1690 VSS.n1967 VSS.n1334 0.853
R1691 VSS.n2028 VSS.n2027 0.853
R1692 VSS.n1332 VSS.n1307 0.853
R1693 VSS.n1315 VSS.n1307 0.853
R1694 VSS.n1321 VSS.n1289 0.853
R1695 VSS.n1322 VSS.n1321 0.853
R1696 VSS.n1288 VSS.n1281 0.853
R1697 VSS.n1281 VSS.n1280 0.853
R1698 VSS.n1248 VSS.n1217 0.853
R1699 VSS.n1248 VSS.n1247 0.853
R1700 VSS.n1256 VSS.n1193 0.853
R1701 VSS.n1193 VSS.n1192 0.853
R1702 VSS.n1226 VSS.n1221 0.853
R1703 VSS.n1235 VSS.n1221 0.853
R1704 VSS.n2027 VSS.n2026 0.853
R1705 VSS.n1258 VSS.n1257 0.853
R1706 VSS.n1165 VSS.n1163 0.853
R1707 VSS.n1196 VSS 0.853
R1708 VSS.n1311 VSS.n1290 0.853
R1709 VSS.n1336 VSS.n1335 0.853
R1710 VSS.n1769 VSS.n1768 0.853
R1711 VSS.n1756 VSS.n1748 0.853
R1712 VSS.n1938 VSS.n1367 0.853
R1713 VSS.n1754 VSS.n1712 0.853
R1714 VSS.n1714 VSS.n1712 0.853
R1715 VSS.n1726 VSS.n1709 0.853
R1716 VSS.n1727 VSS.n1726 0.853
R1717 VSS.n1831 VSS.n1830 0.853
R1718 VSS.n1830 VSS.n1829 0.853
R1719 VSS.n1646 VSS.n1583 0.853
R1720 VSS.n1640 VSS.n1583 0.853
R1721 VSS.n1637 VSS.n1635 0.853
R1722 VSS.n1638 VSS.n1637 0.853
R1723 VSS.n1857 VSS.n1856 0.853
R1724 VSS.n1858 VSS.n1857 0.853
R1725 VSS.n1571 VSS.n1569 0.853
R1726 VSS.n1864 VSS.n1571 0.853
R1727 VSS.n1539 VSS.n1489 0.853
R1728 VSS.n1545 VSS.n1489 0.853
R1729 VSS.n1882 VSS.n1881 0.853
R1730 VSS.n1883 VSS.n1882 0.853
R1731 VSS.n1537 VSS.n1536 0.853
R1732 VSS.n1536 VSS.n1535 0.853
R1733 VSS.n1499 VSS.n1460 0.853
R1734 VSS.n1461 VSS.n1460 0.853
R1735 VSS.n1405 VSS.n1383 0.853
R1736 VSS.n1414 VSS.n1383 0.853
R1737 VSS.n1409 VSS.n1403 0.853
R1738 VSS.n1412 VSS.n1409 0.853
R1739 VSS.n1932 VSS.n1931 0.853
R1740 VSS.n1931 VSS.n1930 0.853
R1741 VSS.n1367 VSS.n1366 0.853
R1742 VSS.n1871 VSS.n1870 0.853
R1743 VSS.n1794 VSS.n1793 0.853
R1744 VSS.n1837 VSS.n1836 0.853
R1745 VSS.n1406 VSS.n1404 0.853
R1746 VSS.n1521 VSS.n1520 0.853
R1747 VSS.n1696 VSS.n1695 0.853
R1748 VSS.n1487 VSS.n1485 0.853
R1749 VSS.n1909 VSS.n1400 0.853
R1750 VSS.n1944 VSS.n1365 0.853
R1751 VSS.n1605 VSS.n1604 0.853
R1752 VSS.n1816 VSS.n1708 0.853
R1753 VSS.n12 VSS.n11 0.853
R1754 VSS.n73 VSS.n56 0.853
R1755 VSS.n1561 VSS.n1487 0.853
R1756 VSS.n1910 VSS.n1909 0.853
R1757 VSS.n1945 VSS.n1944 0.853
R1758 VSS.n1337 VSS.n1336 0.853
R1759 VSS.n1817 VSS.n1816 0.853
R1760 VSS.n1172 VSS.n1167 0.853
R1761 VSS.n28 VSS.n12 0.853
R1762 VSS.n1078 VSS.n1077 0.853
R1763 VSS.n65 VSS.n44 0.853
R1764 VSS.n14 VSS.n13 0.853
R1765 VSS.n1105 VSS.n1100 0.853
R1766 VSS.n1117 VSS.n1116 0.853
R1767 VSS.n56 VSS.n55 0.853
R1768 VSS.n1116 VSS.n1115 0.853
R1769 VSS.n1100 VSS.n1099 0.853
R1770 VSS.n2203 VSS.n2201 0.853
R1771 VSS.n2161 VSS.n2160 0.853
R1772 VSS.n2187 VSS.n2186 0.853
R1773 VSS.n2155 VSS.n2154 0.853
R1774 VSS.n99 VSS.n98 0.853
R1775 VSS.n138 VSS.n137 0.853
R1776 VSS.n984 VSS.n138 0.853
R1777 VSS.n987 VSS.n131 0.853
R1778 VSS.n996 VSS.n93 0.853
R1779 VSS.n993 VSS.n99 0.853
R1780 VSS.n990 VSS.n105 0.853
R1781 VSS.n850 VSS.n175 0.853
R1782 VSS.n847 VSS.n191 0.853
R1783 VSS.n807 VSS.n204 0.853
R1784 VSS.n765 VSS.n763 0.853
R1785 VSS.n953 VSS.n155 0.853
R1786 VSS.n930 VSS.n157 0.853
R1787 VSS.n844 VSS.n843 0.853
R1788 VSS.n824 VSS.n823 0.853
R1789 VSS.n870 VSS.n869 0.853
R1790 VSS.n886 VSS.n885 0.853
R1791 VSS.n927 VSS.n926 0.853
R1792 VSS.n950 VSS.n949 0.853
R1793 VSS.n981 VSS.n980 0.853
R1794 VSS.n785 VSS.n784 0.853
R1795 VSS.n804 VSS.n803 0.853
R1796 VSS.n105 VSS.n103 0.853
R1797 VSS.n479 VSS.n478 0.853
R1798 VSS.n478 VSS.n477 0.853
R1799 VSS.n344 VSS.n343 0.853
R1800 VSS.n321 VSS.n320 0.853
R1801 VSS.n367 VSS.n366 0.853
R1802 VSS.n420 VSS.n419 0.853
R1803 VSS.n447 VSS.n446 0.853
R1804 VSS.n454 VSS.n453 0.853
R1805 VSS.n464 VSS.n463 0.853
R1806 VSS.n695 VSS.n694 0.853
R1807 VSS.n731 VSS.n729 0.853
R1808 VSS.n726 VSS.n724 0.853
R1809 VSS.n392 VSS.n391 0.853
R1810 VSS.n474 VSS.n472 0.853
R1811 VSS.n666 VSS.n665 0.853
R1812 VSS.n643 VSS.n642 0.853
R1813 VSS.n636 VSS.n635 0.853
R1814 VSS.n583 VSS.n582 0.853
R1815 VSS.n574 VSS.n573 0.853
R1816 VSS.n545 VSS.n544 0.853
R1817 VSS.n516 VSS.n515 0.853
R1818 VSS.n717 VSS.n715 0.853
R1819 VSS.n718 VSS.n717 0.853
R1820 VSS.n2072 VSS.n2069 0.853
R1821 VSS.n2101 VSS.n2100 0.853
R1822 VSS.n2100 VSS.n2099 0.853
R1823 VSS.n2119 VSS.n2118 0.853
R1824 VSS.n2118 VSS.n2117 0.853
R1825 VSS.n2086 VSS.n2085 0.853
R1826 VSS.n2087 VSS.n2086 0.853
R1827 VSS.n2073 VSS.n2072 0.853
R1828 VSS.n2204 VSS.n2203 0.853
R1829 VSS.n1775 VSS 0.830206
R1830 VSS.n1168 VSS 0.822548
R1831 VSS.n1263 VSS.n1183 0.753441
R1832 VSS.n409 VSS.n408 0.753441
R1833 VSS.n492 VSS.n489 0.753441
R1834 VSS.n2144 VSS.n2122 0.699777
R1835 VSS.n2189 VSS.n2188 0.699516
R1836 VSS.n1071 VSS.n1063 0.698382
R1837 VSS.n80 VSS.n79 0.684595
R1838 VSS.n299 VSS.n298 0.683764
R1839 VSS.n1607 VSS.n1606 0.683294
R1840 VSS.n979 VSS.n978 0.683294
R1841 VSS.n925 VSS.n924 0.683294
R1842 VSS.n884 VSS.n883 0.683294
R1843 VSS.n868 VSS.n867 0.683294
R1844 VSS.n822 VSS.n821 0.683294
R1845 VSS.n842 VSS.n841 0.683294
R1846 VSS.n948 VSS.n947 0.683294
R1847 VSS.n783 VSS.n782 0.683294
R1848 VSS.n452 VSS.n451 0.683034
R1849 VSS.n641 VSS.n640 0.683034
R1850 VSS.n723 VSS.n722 0.683034
R1851 VSS.n1080 VSS.n1079 0.683034
R1852 VSS.n895 VSS.n894 0.683034
R1853 VSS.n154 VSS.n153 0.683034
R1854 VSS.n762 VSS.n761 0.683034
R1855 VSS.n203 VSS.n202 0.683034
R1856 VSS.n190 VSS.n189 0.683034
R1857 VSS.n174 VSS.n173 0.683034
R1858 VSS.n92 VSS.n91 0.683034
R1859 VSS.n130 VSS.n129 0.683034
R1860 VSS.n802 VSS.n801 0.683034
R1861 VSS.n1982 VSS.n1981 0.565206
R1862 VSS.n1513 VSS.n1512 0.565206
R1863 VSS.n1821 VSS.n1669 0.565206
R1864 VSS.n684 VSS.n683 0.565206
R1865 VSS.n1048 VSS.n1045 0.492808
R1866 VSS.n1031 VSS.n1028 0.492808
R1867 VSS.n921 VSS.n918 0.492808
R1868 VSS.n860 VSS.n859 0.492808
R1869 VSS.n1005 VSS.n1002 0.394346
R1870 VSS.n1076 VSS.n1075 0.380161
R1871 VSS.n744 VSS.n741 0.376971
R1872 VSS.n1784 VSS.n1783 0.376971
R1873 VSS.n1092 VSS.n1091 0.376971
R1874 VSS.n1431 VSS.n1351 0.376971
R1875 VSS.n1512 VSS.n1511 0.376971
R1876 VSS.n386 VSS.n385 0.376971
R1877 VSS.n501 VSS.n498 0.376971
R1878 VSS.n1072 VSS.n1071 0.309535
R1879 VSS.n1905 VSS.n1459 0.212
R1880 VSS.n1867 VSS.n1570 0.212
R1881 VSS.n1834 VSS.n1833 0.212
R1882 VSS.n2009 VSS.n1194 0.212
R1883 VSS.n2139 VSS.n2138 0.203675
R1884 VSS.n1017 VSS.n1013 0.197423
R1885 VSS.n906 VSS.n903 0.197423
R1886 VSS.n758 VSS.n213 0.197423
R1887 VSS.n2036 VSS.n1152 0.188735
R1888 VSS.n1686 VSS.n1680 0.188735
R1889 VSS.n356 VSS.n353 0.188735
R1890 VSS.n2193 VSS.n2192 0.170375
R1891 VSS.n725 VSS.n0 0.128113
R1892 VSS.n1081 VSS.n50 0.120292
R1893 VSS.n2050 VSS.n17 0.120292
R1894 VSS.n2021 VSS.n1182 0.120292
R1895 VSS.n1292 VSS.n1202 0.120292
R1896 VSS.n1341 VSS.n1338 0.120292
R1897 VSS.n1353 VSS.n1345 0.120292
R1898 VSS.n1433 VSS.n1432 0.120292
R1899 VSS.n1914 VSS.n1913 0.120292
R1900 VSS.n1612 VSS.n1611 0.120292
R1901 VSS.n1841 VSS.n1630 0.120292
R1902 VSS.n1798 VSS.n1742 0.120292
R1903 VSS.n442 VSS.n438 0.120292
R1904 VSS.n254 VSS.n248 0.120292
R1905 VSS.n503 VSS.n502 0.120292
R1906 VSS.n613 VSS.n609 0.120292
R1907 VSS.n631 VSS.n627 0.120292
R1908 VSS.n745 VSS.n739 0.120292
R1909 VSS.n1773 VSS.n1772 0.118643
R1910 VSS.n1515 VSS.n1503 0.117688
R1911 VSS.n1704 VSS.n1703 0.116385
R1912 VSS.n487 VSS.n486 0.115083
R1913 VSS.n529 VSS.n528 0.113781
R1914 VSS.n558 VSS.n557 0.113781
R1915 VSS.n594 VSS.n593 0.112479
R1916 VSS.n1267 VSS.n1266 0.111177
R1917 VSS.n284 VSS.n283 0.111177
R1918 VSS.n2059 VSS.n9 0.108573
R1919 VSS.n32 VSS.n29 0.107271
R1920 VSS.n2041 VSS.n2040 0.107271
R1921 VSS.n1894 VSS.n1893 0.107271
R1922 VSS.n1429 VSS.n1427 0.105969
R1923 VSS.n2198 VSS 0.104812
R1924 VSS.n1688 VSS.n1674 0.104667
R1925 VSS.n1678 VSS.n1674 0.104667
R1926 VSS.n1267 VSS.n1265 0.103365
R1927 VSS.n403 VSS.n402 0.103365
R1928 VSS.n1341 VSS.n1340 0.102062
R1929 VSS.n676 VSS.n675 0.102062
R1930 VSS.n47 VSS.n32 0.10076
R1931 VSS.n2040 VSS.n1150 0.0994583
R1932 VSS.n117 VSS.n116 0.0989615
R1933 VSS.n122 VSS.n121 0.0989615
R1934 VSS.n975 VSS.n974 0.0989615
R1935 VSS.n143 VSS.n142 0.0989615
R1936 VSS.n860 VSS.n856 0.0989615
R1937 VSS.n170 VSS.n169 0.0989615
R1938 VSS.n2120 VSS.n0 0.0971532
R1939 VSS.n255 VSS.n254 0.0968542
R1940 VSS.n311 VSS.n310 0.0955521
R1941 VSS.n1877 VSS.n1876 0.09425
R1942 VSS.n1876 VSS.n1875 0.09425
R1943 VSS.n1062 VSS.n1060 0.0939959
R1944 VSS.n1354 VSS.n1353 0.0929479
R1945 VSS.n266 VSS.n265 0.0929479
R1946 VSS.n614 VSS.n613 0.0929479
R1947 VSS.n1432 VSS.n1356 0.0916458
R1948 VSS.n486 VSS.n481 0.0916458
R1949 VSS.n632 VSS.n631 0.0916458
R1950 VSS.n1893 VSS.n1473 0.0903438
R1951 VSS.n1611 VSS.n1610 0.0903438
R1952 VSS.n265 VSS.n261 0.0877396
R1953 VSS.n2022 VSS.n2021 0.0851354
R1954 VSS.n61 VSS.n50 0.0838333
R1955 VSS.n379 VSS.n378 0.0838333
R1956 VSS.n1985 VSS.n1292 0.0825312
R1957 VSS.n1798 VSS.n1797 0.0825312
R1958 VSS.n690 VSS.n689 0.0825312
R1959 VSS.n1209 VSS.n1182 0.0812292
R1960 VSS.n416 VSS.n415 0.0812292
R1961 VSS.n1841 VSS.n1840 0.0799271
R1962 VSS.n1703 VSS.n1671 0.0799271
R1963 VSS.n1914 VSS.n1396 0.078625
R1964 VSS.n653 VSS.n652 0.078625
R1965 VSS.n2051 VSS.n2050 0.0773229
R1966 VSS.n1170 VSS.n17 0.0773229
R1967 VSS.n1516 VSS.n1515 0.0773229
R1968 VSS.n1788 VSS.n1773 0.0760208
R1969 VSS.n712 VSS.n711 0.0760208
R1970 VSS.n339 VSS.n338 0.0747188
R1971 VSS.n739 VSS.n735 0.0747188
R1972 VSS.n1283 VSS.n1202 0.0734167
R1973 VSS.n2184 VSS.n2183 0.0734167
R1974 VSS.n443 VSS.n442 0.0721146
R1975 VSS.n609 VSS.n603 0.0721146
R1976 VSS.n541 VSS.n540 0.0708125
R1977 VSS.n570 VSS.n569 0.0708125
R1978 VSS.n502 VSS.n496 0.0695104
R1979 VSS.n1936 VSS.n1935 0.0685147
R1980 VSS.n1923 VSS.n1386 0.0685147
R1981 VSS.n1417 VSS.n1416 0.0685147
R1982 VSS.n1529 VSS.n1463 0.0685147
R1983 VSS.n1532 VSS.n1491 0.0685147
R1984 VSS.n1549 VSS.n1548 0.0685147
R1985 VSS.n1862 VSS.n1861 0.0685147
R1986 VSS.n1849 VSS.n1586 0.0685147
R1987 VSS.n1641 VSS.n1639 0.0685147
R1988 VSS.n1717 VSS.n1664 0.0685147
R1989 VSS.n1807 VSS.n1730 0.0685147
R1990 VSS.n1762 VSS.n1732 0.0685147
R1991 VSS.n1229 VSS.n1159 0.0685147
R1992 VSS.n1243 VSS.n1219 0.0685147
R1993 VSS.n1245 VSS.n1190 0.0685147
R1994 VSS.n1995 VSS.n1277 0.0685147
R1995 VSS.n1326 VSS.n1325 0.0685147
R1996 VSS.n1974 VSS.n1305 0.0685147
R1997 VSS.n214 VSS.n6 0.0685147
R1998 VSS.n221 VSS.n220 0.0685147
R1999 VSS.n1742 VSS.n1741 0.0682083
R2000 VSS.n1913 VSS.n1912 0.0669062
R2001 VSS.n363 VSS.n362 0.0656042
R2002 VSS.n1360 VSS.n1345 0.0643021
R2003 VSS.n2152 VSS.n2151 0.0643021
R2004 VSS.n248 VSS.n244 0.0643021
R2005 VSS.n1612 VSS.n1608 0.0616979
R2006 VSS.n623 VSS.n622 0.0616979
R2007 VSS.n746 VSS.n745 0.0616979
R2008 VSS.n1082 VSS.n1081 0.0603958
R2009 VSS.n1433 VSS 0.0603958
R2010 VSS VSS.n1429 0.0603958
R2011 VSS.n2059 VSS 0.0603958
R2012 VSS.n1041 VSS.n1037 0.0603958
R2013 VSS.n1032 VSS.n1025 0.0603958
R2014 VSS.n118 VSS.n113 0.0603958
R2015 VSS.n127 VSS.n123 0.0603958
R2016 VSS.n972 VSS.n968 0.0603958
R2017 VSS.n941 VSS.n937 0.0603958
R2018 VSS.n907 VSS.n900 0.0603958
R2019 VSS.n908 VSS.n907 0.0603958
R2020 VSS.n166 VSS.n162 0.0603958
R2021 VSS.n835 VSS.n831 0.0603958
R2022 VSS.n776 VSS.n772 0.0603958
R2023 VSS.n759 VSS.n210 0.0603958
R2024 VSS.n1630 VSS.n1608 0.0590938
R2025 VSS.n627 VSS.n623 0.0590938
R2026 VSS.n747 VSS.n746 0.0590938
R2027 VSS.n840 VSS.n839 0.0571406
R2028 VSS.n781 VSS.n780 0.0564896
R2029 VSS.n1957 VSS.n1337 0.0553246
R2030 VSS.n1042 VSS.n1041 0.0545365
R2031 VSS.n866 VSS.n861 0.0545365
R2032 VSS.n923 VSS.n922 0.0532344
R2033 VSS.n365 VSS.n349 0.0531316
R2034 VSS.n1910 VSS.n1399 0.0531316
R2035 VSS.n1011 VSS.n1007 0.0519323
R2036 VSS.n2165 VSS 0.0512812
R2037 VSS.n152 VSS.n144 0.0512812
R2038 VSS.n1012 VSS.n1011 0.0506302
R2039 VSS.n172 VSS.n171 0.0506302
R2040 VSS.n800 VSS.n795 0.0499792
R2041 VSS.n2192 VSS.n2122 0.0498797
R2042 VSS.n634 VSS.n589 0.0487456
R2043 VSS.n1818 VSS.n1817 0.0487456
R2044 VSS.n479 VSS.n271 0.0487456
R2045 VSS.n1377 VSS.n1371 0.0482941
R2046 VSS.n1925 VSS.n1384 0.0482941
R2047 VSS.n1419 VSS.n1410 0.0482941
R2048 VSS.n1527 VSS.n1526 0.0482941
R2049 VSS.n1543 VSS.n1492 0.0482941
R2050 VSS.n1552 VSS.n1551 0.0482941
R2051 VSS.n1576 VSS.n1574 0.0482941
R2052 VSS.n1851 VSS.n1584 0.0482941
R2053 VSS.n1652 VSS.n1643 0.0482941
R2054 VSS.n1724 VSS.n1723 0.0482941
R2055 VSS.n1809 VSS.n1713 0.0482941
R2056 VSS.n1760 VSS.n1751 0.0482941
R2057 VSS.n1231 VSS.n1224 0.0482941
R2058 VSS.n1241 VSS.n1240 0.0482941
R2059 VSS.n1252 VSS.n1250 0.0482941
R2060 VSS.n1993 VSS.n1278 0.0482941
R2061 VSS.n1328 VSS.n1314 0.0482941
R2062 VSS.n1972 VSS.n1306 0.0482941
R2063 VSS.n69 VSS.n59 0.0482941
R2064 VSS.n1110 VSS.n1101 0.0482941
R2065 VSS.n1138 VSS.n25 0.0482941
R2066 VSS.n896 VSS.n893 0.047375
R2067 VSS VSS.n1062 0.047248
R2068 VSS.n471 VSS.n469 0.0465526
R2069 VSS.n634 VSS.n588 0.0465526
R2070 VSS.n543 VSS.n521 0.0465526
R2071 VSS.n1358 VSS.n1355 0.0465526
R2072 VSS.n1945 VSS.n1357 0.0465526
R2073 VSS.n479 VSS.n270 0.0465526
R2074 VSS.n296 VSS.n295 0.0443596
R2075 VSS.n572 VSS.n550 0.0443596
R2076 VSS.n1561 VSS.n1559 0.0443596
R2077 VSS.n1878 VSS.n1562 0.0443596
R2078 VSS.n1874 VSS.n1873 0.0443596
R2079 VSS.n1872 VSS.n1566 0.0443596
R2080 VSS.n968 VSS.n964 0.0441198
R2081 VSS.n882 VSS.n881 0.0441198
R2082 VSS.n188 VSS.n183 0.0434688
R2083 VSS.n2154 VSS.n2145 0.0427297
R2084 VSS.n319 VSS.n303 0.0421667
R2085 VSS.n318 VSS.n317 0.0421667
R2086 VSS.n445 VSS.n425 0.0421667
R2087 VSS.n462 VSS.n461 0.0421667
R2088 VSS.n581 VSS.n579 0.0421667
R2089 VSS.n1025 VSS.n1021 0.0421667
R2090 VSS.n1067 VSS.n1065 0.0415156
R2091 VSS.n2201 VSS.n2196 0.0415156
R2092 VSS.n2158 VSS.n2157 0.0411354
R2093 VSS.n946 VSS.n945 0.0402135
R2094 VSS.n342 VSS.n326 0.0399737
R2095 VSS.n460 VSS.n459 0.0399737
R2096 VSS.n2005 VSS.n1197 0.0399737
R2097 VSS.n135 VSS.n134 0.0399737
R2098 VSS.n137 VSS.n136 0.0399737
R2099 VSS.n1937 VSS.n1936 0.0391029
R2100 VSS.n1935 VSS.n1370 0.0391029
R2101 VSS.n1386 VSS.n1372 0.0391029
R2102 VSS.n1923 VSS.n1922 0.0391029
R2103 VSS.n1416 VSS.n1387 0.0391029
R2104 VSS.n1417 VSS.n1390 0.0391029
R2105 VSS.n1938 VSS.n1369 0.0391029
R2106 VSS.n1934 VSS.n1933 0.0391029
R2107 VSS.n1932 VSS.n1373 0.0391029
R2108 VSS.n1924 VSS.n1385 0.0391029
R2109 VSS.n1415 VSS.n1414 0.0391029
R2110 VSS.n1418 VSS.n1413 0.0391029
R2111 VSS.n1902 VSS.n1463 0.0391029
R2112 VSS.n1530 VSS.n1529 0.0391029
R2113 VSS.n1533 VSS.n1532 0.0391029
R2114 VSS.n1546 VSS.n1491 0.0391029
R2115 VSS.n1549 VSS.n1547 0.0391029
R2116 VSS.n1548 VSS.n1481 0.0391029
R2117 VSS.n1497 VSS.n1462 0.0391029
R2118 VSS.n1535 VSS.n1528 0.0391029
R2119 VSS.n1534 VSS.n1531 0.0391029
R2120 VSS.n1545 VSS.n1544 0.0391029
R2121 VSS.n1550 VSS.n1490 0.0391029
R2122 VSS.n1883 VSS.n1483 0.0391029
R2123 VSS.n1862 VSS.n1573 0.0391029
R2124 VSS.n1861 VSS.n1575 0.0391029
R2125 VSS.n1586 VSS.n1577 0.0391029
R2126 VSS.n1849 VSS.n1848 0.0391029
R2127 VSS.n1641 VSS.n1587 0.0391029
R2128 VSS.n1655 VSS.n1639 0.0391029
R2129 VSS.n1864 VSS.n1863 0.0391029
R2130 VSS.n1860 VSS.n1859 0.0391029
R2131 VSS.n1858 VSS.n1578 0.0391029
R2132 VSS.n1850 VSS.n1585 0.0391029
R2133 VSS.n1642 VSS.n1640 0.0391029
R2134 VSS.n1654 VSS.n1653 0.0391029
R2135 VSS.n1827 VSS.n1664 0.0391029
R2136 VSS.n1718 VSS.n1717 0.0391029
R2137 VSS.n1730 VSS.n1715 0.0391029
R2138 VSS.n1807 VSS.n1806 0.0391029
R2139 VSS.n1805 VSS.n1732 0.0391029
R2140 VSS.n1763 VSS.n1762 0.0391029
R2141 VSS.n1828 VSS.n1663 0.0391029
R2142 VSS.n1727 VSS.n1716 0.0391029
R2143 VSS.n1729 VSS.n1728 0.0391029
R2144 VSS.n1808 VSS.n1714 0.0391029
R2145 VSS.n1750 VSS.n1731 0.0391029
R2146 VSS.n1764 VSS.n1761 0.0391029
R2147 VSS.n2029 VSS.n1159 0.0391029
R2148 VSS.n1229 VSS.n1228 0.0391029
R2149 VSS.n1227 VSS.n1219 0.0391029
R2150 VSS.n1244 VSS.n1243 0.0391029
R2151 VSS.n1246 VSS.n1245 0.0391029
R2152 VSS.n2012 VSS.n1190 0.0391029
R2153 VSS.n2028 VSS.n1160 0.0391029
R2154 VSS.n1230 VSS.n1225 0.0391029
R2155 VSS.n1226 VSS.n1220 0.0391029
R2156 VSS.n1242 VSS.n1218 0.0391029
R2157 VSS.n1247 VSS.n1214 0.0391029
R2158 VSS.n1251 VSS.n1191 0.0391029
R2159 VSS.n1996 VSS.n1995 0.0391029
R2160 VSS.n1318 VSS.n1277 0.0391029
R2161 VSS.n1325 VSS.n1316 0.0391029
R2162 VSS.n1326 VSS.n1303 0.0391029
R2163 VSS.n1975 VSS.n1974 0.0391029
R2164 VSS.n1962 VSS.n1305 0.0391029
R2165 VSS.n1994 VSS.n1276 0.0391029
R2166 VSS.n1322 VSS.n1317 0.0391029
R2167 VSS.n1324 VSS.n1323 0.0391029
R2168 VSS.n1327 VSS.n1315 0.0391029
R2169 VSS.n1973 VSS.n1304 0.0391029
R2170 VSS.n1963 VSS.n1961 0.0391029
R2171 VSS.n73 VSS.n70 0.0391029
R2172 VSS.n58 VSS.n38 0.0391029
R2173 VSS.n1117 VSS.n40 0.0391029
R2174 VSS.n1109 VSS.n1102 0.0391029
R2175 VSS.n1105 VSS.n1104 0.0391029
R2176 VSS.n1140 VSS.n1139 0.0391029
R2177 VSS.n2057 VSS.n11 0.0391029
R2178 VSS.n2067 VSS.n6 0.0391029
R2179 VSS.n215 VSS.n214 0.0391029
R2180 VSS.n220 VSS.n219 0.0391029
R2181 VSS.n222 VSS.n221 0.0391029
R2182 VSS.n224 VSS.n223 0.0391029
R2183 VSS.n2115 VSS.n2109 0.0391029
R2184 VSS.n5 VSS.n4 0.0391029
R2185 VSS.n2085 VSS.n2081 0.0391029
R2186 VSS.n2084 VSS.n2083 0.0391029
R2187 VSS.n2099 VSS.n2095 0.0391029
R2188 VSS.n2098 VSS.n2097 0.0391029
R2189 VSS.n2117 VSS.n2108 0.0391029
R2190 VSS.n128 VSS.n118 0.0389115
R2191 VSS.n201 VSS.n196 0.0382604
R2192 VSS.n733 VSS.n234 0.0377807
R2193 VSS.n1519 VSS.n1518 0.0377807
R2194 VSS.n2023 VSS.n1166 0.0377807
R2195 VSS.n1776 VSS.n1769 0.0377807
R2196 VSS.n1173 VSS.n1172 0.0377807
R2197 VSS.n2190 VSS.n2189 0.0361962
R2198 VSS.n2142 VSS.n2141 0.035973
R2199 VSS.n2161 VSS.n2143 0.035973
R2200 VSS.n760 VSS.n759 0.0356562
R2201 VSS.n1132 VSS.n15 0.0355877
R2202 VSS.n715 VSS.n699 0.0355877
R2203 VSS.n1037 VSS.n1033 0.0343542
R2204 VSS.n2194 VSS.n2193 0.0342265
R2205 VSS.n664 VSS.n663 0.0333947
R2206 VSS.n390 VSS.n372 0.0333947
R2207 VSS.n693 VSS.n692 0.0333947
R2208 VSS.n1453 VSS.n1426 0.0333947
R2209 VSS.n1838 VSS.n1633 0.0333947
R2210 VSS.n98 VSS.n96 0.0333947
R2211 VSS.n1956 VSS.n1339 0.0330521
R2212 VSS.n2153 VSS 0.0330521
R2213 VSS.n2186 VSS.n2127 0.0325946
R2214 VSS.n1506 VSS.n1397 0.03175
R2215 VSS VSS.n2163 0.03175
R2216 VSS.n364 VSS.n358 0.03175
R2217 VSS.n418 VSS.n398 0.0312018
R2218 VSS.n514 VSS.n240 0.0312018
R2219 VSS.n62 VSS.n45 0.0312018
R2220 VSS.n1698 VSS.n1697 0.0312018
R2221 VSS.n1796 VSS.n1795 0.0312018
R2222 VSS.n103 VSS.n102 0.0312018
R2223 VSS.n977 VSS.n972 0.0304479
R2224 VSS.n977 VSS.n976 0.0304479
R2225 VSS.n908 VSS 0.0304479
R2226 VSS.n915 VSS 0.0304479
R2227 VSS.n820 VSS.n815 0.0304479
R2228 VSS.n820 VSS.n819 0.0304479
R2229 VSS.n210 VSS 0.0304479
R2230 VSS.n2125 VSS.n2124 0.029875
R2231 VSS.n1819 VSS.n1705 0.0291458
R2232 VSS.n481 VSS.n480 0.0291458
R2233 VSS.n633 VSS.n632 0.0291458
R2234 VSS.n1986 VSS.n1291 0.0290088
R2235 VSS.n1294 VSS.n1291 0.0290088
R2236 VSS.n1210 VSS.n1208 0.0290088
R2237 VSS.n1260 VSS.n1208 0.0290088
R2238 VSS.n1947 VSS.n1354 0.0278438
R2239 VSS.n1946 VSS.n1356 0.0278438
R2240 VSS.n2163 VSS.n2162 0.0278438
R2241 VSS.n480 VSS.n266 0.0278438
R2242 VSS.n495 VSS.n494 0.0278438
R2243 VSS.n542 VSS.n536 0.0278438
R2244 VSS.n633 VSS.n614 0.0278438
R2245 VSS.n418 VSS.n397 0.0268158
R2246 VSS.n514 VSS.n239 0.0268158
R2247 VSS.n1094 VSS.n45 0.0268158
R2248 VSS.n1697 VSS.n1692 0.0268158
R2249 VSS.n1795 VSS.n1745 0.0268158
R2250 VSS.n103 VSS.n101 0.0268158
R2251 VSS.n1560 VSS.n1473 0.0265417
R2252 VSS.n1877 VSS.n1475 0.0265417
R2253 VSS.n1875 VSS.n1563 0.0265417
R2254 VSS.n1610 VSS.n1565 0.0265417
R2255 VSS.n1033 VSS.n1032 0.0265417
R2256 VSS.n294 VSS.n293 0.0265417
R2257 VSS.n571 VSS.n565 0.0265417
R2258 VSS.n764 VSS.n0 0.0261804
R2259 VSS.n2199 VSS.n2198 0.0257686
R2260 VSS.n760 VSS.n209 0.0252396
R2261 VSS.n316 VSS.n304 0.0252396
R2262 VSS.n315 VSS.n311 0.0252396
R2263 VSS.n444 VSS.n434 0.0252396
R2264 VSS.n261 VSS.n260 0.0252396
R2265 VSS.n602 VSS.n601 0.0252396
R2266 VSS VSS.n2205 0.0252105
R2267 VSS.n664 VSS.n648 0.0246228
R2268 VSS.n390 VSS.n389 0.0246228
R2269 VSS.n693 VSS.n671 0.0246228
R2270 VSS.n1454 VSS.n1453 0.0246228
R2271 VSS.n1839 VSS.n1838 0.0246228
R2272 VSS.n98 VSS.n97 0.0246228
R2273 VSS.n929 VSS.n928 0.0244361
R2274 VSS.n1068 VSS.n1066 0.024008
R2275 VSS.n2004 VSS.n1199 0.0239375
R2276 VSS.n340 VSS.n334 0.0239375
R2277 VSS.n259 VSS.n255 0.0239375
R2278 VSS.n1171 VSS.n1149 0.0226354
R2279 VSS.n2022 VSS.n1181 0.0226354
R2280 VSS.n1956 VSS.n1338 0.0226354
R2281 VSS.n1517 VSS.n1472 0.0226354
R2282 VSS.n1787 VSS.n1786 0.0226354
R2283 VSS.n2183 VSS 0.0226354
R2284 VSS.n201 VSS.n200 0.0226354
R2285 VSS.n734 VSS.n233 0.0226354
R2286 VSS.n2052 VSS.n15 0.0224298
R2287 VSS.n715 VSS.n714 0.0224298
R2288 VSS.n2201 VSS.n2200 0.0223823
R2289 VSS.n74 VSS.n73 0.0220382
R2290 VSS.n128 VSS.n127 0.0219844
R2291 VSS.n1939 VSS.n1938 0.0219755
R2292 VSS.n1884 VSS.n1883 0.0219755
R2293 VSS.n1865 VSS.n1864 0.0219755
R2294 VSS.n1765 VSS.n1764 0.0219755
R2295 VSS.n2028 VSS.n1158 0.0219755
R2296 VSS.n1964 VSS.n1963 0.0219755
R2297 VSS.n2117 VSS.n2116 0.0219755
R2298 VSS.n547 VSS.n546 0.0213351
R2299 VSS.n1131 VSS.n16 0.0213333
R2300 VSS.n1153 VSS.n1150 0.0213333
R2301 VSS.n2140 VSS.n2130 0.0213333
R2302 VSS.n358 VSS.n352 0.0213333
R2303 VSS.n503 VSS 0.0213333
R2304 VSS.n713 VSS.n707 0.0213333
R2305 VSS.n747 VSS 0.0213333
R2306 VSS.n576 VSS.n575 0.0212381
R2307 VSS.n946 VSS.n941 0.0206823
R2308 VSS.n733 VSS.n732 0.0202368
R2309 VSS.n1519 VSS.n1502 0.0202368
R2310 VSS.n1179 VSS.n1166 0.0202368
R2311 VSS.n1789 VSS.n1769 0.0202368
R2312 VSS.n1172 VSS.n1169 0.0202368
R2313 VSS.n48 VSS.n47 0.0200312
R2314 VSS.n1452 VSS.n1451 0.0200312
R2315 VSS.n1507 VSS.n1506 0.0200312
R2316 VSS.n1676 VSS.n1631 0.0200312
R2317 VSS.n2185 VSS.n2182 0.0200312
R2318 VSS.n388 VSS.n379 0.0200312
R2319 VSS.n381 VSS.n380 0.0200312
R2320 VSS VSS.n241 0.0200312
R2321 VSS.n662 VSS.n661 0.0200312
R2322 VSS.n691 VSS.n690 0.0200312
R2323 VSS.n1940 VSS.n1367 0.0191618
R2324 VSS.n1378 VSS.n1367 0.0191618
R2325 VSS.n1931 VSS.n1374 0.0191618
R2326 VSS.n1931 VSS.n1375 0.0191618
R2327 VSS.n1926 VSS.n1383 0.0191618
R2328 VSS.n1408 VSS.n1383 0.0191618
R2329 VSS.n1420 VSS.n1409 0.0191618
R2330 VSS.n1409 VSS.n1402 0.0191618
R2331 VSS.n1904 VSS.n1460 0.0191618
R2332 VSS.n1525 VSS.n1460 0.0191618
R2333 VSS.n1536 VSS.n1495 0.0191618
R2334 VSS.n1536 VSS.n1496 0.0191618
R2335 VSS.n1542 VSS.n1489 0.0191618
R2336 VSS.n1553 VSS.n1489 0.0191618
R2337 VSS.n1882 VSS.n1484 0.0191618
R2338 VSS.n1882 VSS.n1482 0.0191618
R2339 VSS.n1866 VSS.n1571 0.0191618
R2340 VSS.n1600 VSS.n1571 0.0191618
R2341 VSS.n1857 VSS.n1579 0.0191618
R2342 VSS.n1857 VSS.n1580 0.0191618
R2343 VSS.n1852 VSS.n1583 0.0191618
R2344 VSS.n1644 VSS.n1583 0.0191618
R2345 VSS.n1651 VSS.n1637 0.0191618
R2346 VSS.n1657 VSS.n1637 0.0191618
R2347 VSS.n1830 VSS.n1658 0.0191618
R2348 VSS.n1830 VSS.n1661 0.0191618
R2349 VSS.n1726 VSS.n1725 0.0191618
R2350 VSS.n1726 VSS.n1711 0.0191618
R2351 VSS.n1810 VSS.n1712 0.0191618
R2352 VSS.n1752 VSS.n1712 0.0191618
R2353 VSS.n1759 VSS.n1748 0.0191618
R2354 VSS.n1766 VSS.n1748 0.0191618
R2355 VSS.n2027 VSS.n1161 0.0191618
R2356 VSS.n2027 VSS.n1162 0.0191618
R2357 VSS.n1232 VSS.n1221 0.0191618
R2358 VSS.n1239 VSS.n1221 0.0191618
R2359 VSS.n1248 VSS.n1215 0.0191618
R2360 VSS.n1249 VSS.n1248 0.0191618
R2361 VSS.n1253 VSS.n1193 0.0191618
R2362 VSS.n2010 VSS.n1193 0.0191618
R2363 VSS.n1281 VSS.n1279 0.0191618
R2364 VSS.n1992 VSS.n1281 0.0191618
R2365 VSS.n1321 VSS.n1319 0.0191618
R2366 VSS.n1321 VSS.n1320 0.0191618
R2367 VSS.n1329 VSS.n1307 0.0191618
R2368 VSS.n1971 VSS.n1307 0.0191618
R2369 VSS.n1334 VSS.n1333 0.0191618
R2370 VSS.n1965 VSS.n1334 0.0191618
R2371 VSS.n75 VSS.n56 0.0191618
R2372 VSS.n68 VSS.n56 0.0191618
R2373 VSS.n1116 VSS.n41 0.0191618
R2374 VSS.n1116 VSS.n42 0.0191618
R2375 VSS.n1111 VSS.n1100 0.0191618
R2376 VSS.n1100 VSS.n1098 0.0191618
R2377 VSS.n1137 VSS.n12 0.0191618
R2378 VSS.n2056 VSS.n12 0.0191618
R2379 VSS.n2072 VSS.n2 0.0191618
R2380 VSS.n2072 VSS.n2071 0.0191618
R2381 VSS.n2086 VSS.n2077 0.0191618
R2382 VSS.n2086 VSS.n2079 0.0191618
R2383 VSS.n2100 VSS.n2091 0.0191618
R2384 VSS.n2100 VSS.n2093 0.0191618
R2385 VSS.n2118 VSS.n2105 0.0191618
R2386 VSS.n2118 VSS.n2106 0.0191618
R2387 VSS.n61 VSS.n46 0.0187292
R2388 VSS.n1340 VSS.n1293 0.0187292
R2389 VSS.n1699 VSS.n1690 0.0187292
R2390 VSS.n1820 VSS.n1819 0.0187292
R2391 VSS.n1797 VSS.n1743 0.0187292
R2392 VSS.n417 VSS.n416 0.0187292
R2393 VSS.n513 VSS.n512 0.0187292
R2394 VSS.n677 VSS.n676 0.0187292
R2395 VSS.n585 VSS.n584 0.0185247
R2396 VSS.n2192 VSS.n2191 0.0183481
R2397 VSS.n2191 VSS.n2190 0.0183481
R2398 VSS.n872 VSS.n871 0.0181371
R2399 VSS.n342 VSS.n341 0.0180439
R2400 VSS.n1284 VSS.n1197 0.0180439
R2401 VSS.n456 VSS.n455 0.0178464
R2402 VSS.n518 VSS.n517 0.0175557
R2403 VSS.n849 VSS.n848 0.0174588
R2404 VSS.n1209 VSS.n1207 0.0174271
R2405 VSS.n1261 VSS.n1207 0.0174271
R2406 VSS.n1265 VSS.n1262 0.0174271
R2407 VSS.n1985 VSS.n1984 0.0174271
R2408 VSS.n1984 VSS.n1983 0.0174271
R2409 VSS.n188 VSS.n187 0.0174271
R2410 VSS.n404 VSS.n403 0.0174271
R2411 VSS.n494 VSS.n488 0.0174271
R2412 VSS.n952 VSS.n951 0.0168773
R2413 VSS.n638 VSS.n637 0.0168773
R2414 VSS.n882 VSS.n877 0.016776
R2415 VSS.n989 VSS.n988 0.0166835
R2416 VSS.n932 VSS.n931 0.0164897
R2417 VSS.n826 VSS.n825 0.0164897
R2418 VSS.n986 VSS.n985 0.0163928
R2419 VSS.n983 VSS.n982 0.0162959
R2420 VSS.n369 VSS.n368 0.0162959
R2421 VSS.n473 VSS.n236 0.0162959
R2422 VSS.n71 VSS.n37 0.016285
R2423 VSS.n1108 VSS.n39 0.016285
R2424 VSS.n1103 VSS.n24 0.016285
R2425 VSS.n2193 VSS 0.0161945
R2426 VSS.n1093 VSS.n46 0.016125
R2427 VSS.n1678 VSS.n1677 0.016125
R2428 VSS.n1689 VSS.n1688 0.016125
R2429 VSS.n1690 VSS.n1671 0.016125
R2430 VSS.n1770 VSS.n1743 0.016125
R2431 VSS.n417 VSS.n410 0.016125
R2432 VSS.n513 VSS.n241 0.016125
R2433 VSS.n243 VSS.n242 0.016125
R2434 VSS.n536 VSS.n530 0.016125
R2435 VSS.n565 VSS.n559 0.016125
R2436 VSS VSS.n1 0.0160275
R2437 VSS VSS.n2121 0.0160275
R2438 VSS.n668 VSS.n667 0.0159082
R2439 VSS.n445 VSS.n426 0.0158509
R2440 VSS.n581 VSS.n580 0.0158509
R2441 VSS.n137 VSS.n135 0.0158509
R2442 VSS.n476 VSS.n475 0.0158113
R2443 VSS.n955 VSS.n954 0.0156175
R2444 VSS.n767 VSS.n766 0.0156175
R2445 VSS.n323 VSS.n322 0.0156175
R2446 VSS.n1070 VSS.n1064 0.0156071
R2447 VSS.n1074 VSS.n81 0.0156071
R2448 VSS.n2203 VSS.n2195 0.0156071
R2449 VSS.n2203 VSS.n2202 0.0156071
R2450 VSS.n846 VSS.n845 0.0155206
R2451 VSS.n992 VSS.n991 0.0153268
R2452 VSS.n394 VSS.n393 0.0153268
R2453 VSS.n995 VSS.n994 0.015133
R2454 VSS.n453 VSS.n450 0.0150862
R2455 VSS.n642 VSS.n639 0.0150862
R2456 VSS.n472 VSS.n467 0.0150862
R2457 VSS.n472 VSS.n468 0.0150862
R2458 VSS.n724 VSS.n721 0.0150862
R2459 VSS.n731 VSS.n235 0.0150862
R2460 VSS.n731 VSS.n730 0.0150862
R2461 VSS.n665 VSS.n646 0.0150862
R2462 VSS.n665 VSS.n647 0.0150862
R2463 VSS.n391 VSS.n370 0.0150862
R2464 VSS.n391 VSS.n371 0.0150862
R2465 VSS.n343 VSS.n324 0.0150862
R2466 VSS.n343 VSS.n325 0.0150862
R2467 VSS.n320 VSS.n301 0.0150862
R2468 VSS.n320 VSS.n302 0.0150862
R2469 VSS.n297 VSS.n274 0.0150862
R2470 VSS.n446 VSS.n423 0.0150862
R2471 VSS.n446 VSS.n424 0.0150862
R2472 VSS.n419 VSS.n395 0.0150862
R2473 VSS.n419 VSS.n396 0.0150862
R2474 VSS.n366 VSS.n347 0.0150862
R2475 VSS.n366 VSS.n348 0.0150862
R2476 VSS.n463 VSS.n457 0.0150862
R2477 VSS.n463 VSS.n458 0.0150862
R2478 VSS.n635 VSS.n586 0.0150862
R2479 VSS.n635 VSS.n587 0.0150862
R2480 VSS.n582 VSS.n577 0.0150862
R2481 VSS.n582 VSS.n578 0.0150862
R2482 VSS.n573 VSS.n548 0.0150862
R2483 VSS.n573 VSS.n549 0.0150862
R2484 VSS.n544 VSS.n519 0.0150862
R2485 VSS.n544 VSS.n520 0.0150862
R2486 VSS.n515 VSS.n237 0.0150862
R2487 VSS.n515 VSS.n238 0.0150862
R2488 VSS.n694 VSS.n669 0.0150862
R2489 VSS.n694 VSS.n670 0.0150862
R2490 VSS.n1078 VSS.n54 0.0150862
R2491 VSS.n63 VSS.n44 0.0150862
R2492 VSS.n1095 VSS.n44 0.0150862
R2493 VSS.n1133 VSS.n14 0.0150862
R2494 VSS.n2053 VSS.n14 0.0150862
R2495 VSS.n1696 VSS.n1691 0.0150862
R2496 VSS.n1696 VSS.n1693 0.0150862
R2497 VSS.n1558 VSS.n1487 0.0150862
R2498 VSS.n1879 VSS.n1487 0.0150862
R2499 VSS.n1520 VSS.n1500 0.0150862
R2500 VSS.n1520 VSS.n1501 0.0150862
R2501 VSS.n1909 VSS.n1398 0.0150862
R2502 VSS.n1909 VSS.n1908 0.0150862
R2503 VSS.n1425 VSS.n1404 0.0150862
R2504 VSS.n1455 VSS.n1404 0.0150862
R2505 VSS.n1944 VSS.n1359 0.0150862
R2506 VSS.n1944 VSS.n1943 0.0150862
R2507 VSS.n1605 VSS.n1597 0.0150862
R2508 VSS.n1837 VSS.n1632 0.0150862
R2509 VSS.n1837 VSS.n1634 0.0150862
R2510 VSS.n1794 VSS.n1744 0.0150862
R2511 VSS.n1794 VSS.n1746 0.0150862
R2512 VSS.n1871 VSS.n1564 0.0150862
R2513 VSS.n1871 VSS.n1567 0.0150862
R2514 VSS.n1958 VSS.n1336 0.0150862
R2515 VSS.n1362 VSS.n1336 0.0150862
R2516 VSS.n1987 VSS.n1290 0.0150862
R2517 VSS.n1309 VSS.n1290 0.0150862
R2518 VSS.n2006 VSS.n1196 0.0150862
R2519 VSS.n1285 VSS.n1196 0.0150862
R2520 VSS.n1178 VSS.n1165 0.0150862
R2521 VSS.n2024 VSS.n1165 0.0150862
R2522 VSS.n1258 VSS.n1211 0.0150862
R2523 VSS.n1259 VSS.n1258 0.0150862
R2524 VSS.n1790 VSS.n1768 0.0150862
R2525 VSS.n1816 VSS.n1706 0.0150862
R2526 VSS.n1816 VSS.n1815 0.0150862
R2527 VSS.n1174 VSS.n1167 0.0150862
R2528 VSS.n980 VSS.n956 0.0150862
R2529 VSS.n926 VSS.n889 0.0150862
R2530 VSS.n885 VSS.n873 0.0150862
R2531 VSS.n869 VSS.n853 0.0150862
R2532 VSS.n823 VSS.n810 0.0150862
R2533 VSS.n843 VSS.n827 0.0150862
R2534 VSS.n157 VSS.n156 0.0150862
R2535 VSS.n949 VSS.n933 0.0150862
R2536 VSS.n155 VSS.n139 0.0150862
R2537 VSS.n784 VSS.n768 0.0150862
R2538 VSS.n763 VSS.n205 0.0150862
R2539 VSS.n204 VSS.n192 0.0150862
R2540 VSS.n191 VSS.n176 0.0150862
R2541 VSS.n175 VSS.n158 0.0150862
R2542 VSS.n105 VSS.n100 0.0150862
R2543 VSS.n105 VSS.n104 0.0150862
R2544 VSS.n99 VSS.n94 0.0150862
R2545 VSS.n99 VSS.n95 0.0150862
R2546 VSS.n93 VSS.n90 0.0150862
R2547 VSS.n131 VSS.n106 0.0150862
R2548 VSS.n138 VSS.n132 0.0150862
R2549 VSS.n138 VSS.n133 0.0150862
R2550 VSS.n803 VSS.n788 0.0150862
R2551 VSS.n717 VSS.n698 0.0150862
R2552 VSS.n717 VSS.n716 0.0150862
R2553 VSS.n478 VSS.n272 0.0150862
R2554 VSS.n478 VSS.n273 0.0150862
R2555 VSS.n645 VSS.n644 0.0150361
R2556 VSS.n300 VSS.n299 0.0149392
R2557 VSS.n852 VSS.n851 0.0148423
R2558 VSS.n1450 VSS.n1427 0.0148229
R2559 VSS.n1452 VSS.n1396 0.0148229
R2560 VSS.n1840 VSS.n1631 0.0148229
R2561 VSS.n388 VSS.n387 0.0148229
R2562 VSS.n434 VSS.n428 0.0148229
R2563 VSS.n601 VSS.n595 0.0148229
R2564 VSS.n662 VSS.n653 0.0148229
R2565 VSS.n655 VSS.n654 0.0148229
R2566 VSS.n691 VSS.n685 0.0148229
R2567 VSS.n787 VSS.n786 0.0146485
R2568 VSS.n728 VSS.n727 0.0145515
R2569 VSS.n1380 VSS.n1379 0.0143235
R2570 VSS.n1928 VSS.n1927 0.0143235
R2571 VSS.n1422 VSS.n1421 0.0143235
R2572 VSS.n1524 VSS.n1498 0.0143235
R2573 VSS.n1541 VSS.n1493 0.0143235
R2574 VSS.n1555 VSS.n1554 0.0143235
R2575 VSS.n1602 VSS.n1601 0.0143235
R2576 VSS.n1854 VSS.n1853 0.0143235
R2577 VSS.n1650 VSS.n1645 0.0143235
R2578 VSS.n1722 VSS.n1719 0.0143235
R2579 VSS.n1812 VSS.n1811 0.0143235
R2580 VSS.n1758 VSS.n1753 0.0143235
R2581 VSS.n1233 VSS.n1223 0.0143235
R2582 VSS.n1238 VSS.n1222 0.0143235
R2583 VSS.n1254 VSS.n1213 0.0143235
R2584 VSS.n1991 VSS.n1282 0.0143235
R2585 VSS.n1330 VSS.n1313 0.0143235
R2586 VSS.n1970 VSS.n1308 0.0143235
R2587 VSS.n67 VSS.n60 0.0143235
R2588 VSS.n1113 VSS.n1112 0.0143235
R2589 VSS.n1136 VSS.n26 0.0143235
R2590 VSS.n2198 VSS.n2197 0.0142993
R2591 VSS.n806 VSS.n805 0.0142608
R2592 VSS.n1694 VSS.n1636 0.0140833
R2593 VSS.n2054 VSS 0.0139167
R2594 VSS.n888 VSS.n887 0.0138732
R2595 VSS.n422 VSS.n421 0.0138732
R2596 VSS.n346 VSS.n345 0.0137763
R2597 VSS.n449 VSS.n448 0.0137763
R2598 VSS.n1069 VSS.n1068 0.0137243
R2599 VSS.n2156 VSS.n2155 0.0137188
R2600 VSS.n2160 VSS.n2159 0.0137188
R2601 VSS.n2187 VSS.n2126 0.0137188
R2602 VSS.n809 VSS.n808 0.0136794
R2603 VSS.n1177 VSS.n1175 0.0136667
R2604 VSS.n296 VSS.n275 0.0136579
R2605 VSS.n462 VSS.n460 0.0136579
R2606 VSS.n572 VSS.n551 0.0136579
R2607 VSS.n1130 VSS.n29 0.0135208
R2608 VSS.n2051 VSS.n16 0.0135208
R2609 VSS.n2042 VSS.n2041 0.0135208
R2610 VSS.n2004 VSS.n1198 0.0135208
R2611 VSS.n1895 VSS.n1894 0.0135208
R2612 VSS.n2181 VSS.n2168 0.0135208
R2613 VSS.n900 VSS.n896 0.0135208
R2614 VSS.n293 VSS.n285 0.0135208
R2615 VSS.n713 VSS.n712 0.0135208
R2616 VSS.n2008 VSS.n2007 0.0135
R2617 VSS.n697 VSS.n696 0.0134856
R2618 VSS.n720 VSS.n719 0.0127103
R2619 VSS.n2186 VSS.n2128 0.0123243
R2620 VSS.n1171 VSS.n1170 0.0122188
R2621 VSS.n1181 VSS.n1180 0.0122188
R2622 VSS.n1517 VSS.n1516 0.0122188
R2623 VSS.n1788 VSS.n1787 0.0122188
R2624 VSS.n1774 VSS.n9 0.0122188
R2625 VSS.n962 VSS.n957 0.0122188
R2626 VSS.n964 VSS.n963 0.0122188
R2627 VSS.n334 VSS.n328 0.0122188
R2628 VSS.n701 VSS.n700 0.0122188
R2629 VSS.n735 VSS.n734 0.0122188
R2630 VSS.n2199 VSS 0.0121822
R2631 VSS.n466 VSS.n465 0.0119351
R2632 VSS.n1377 VSS.n1369 0.0115294
R2633 VSS.n1384 VSS.n1373 0.0115294
R2634 VSS.n1415 VSS.n1410 0.0115294
R2635 VSS.n1528 VSS.n1527 0.0115294
R2636 VSS.n1544 VSS.n1543 0.0115294
R2637 VSS.n1551 VSS.n1483 0.0115294
R2638 VSS.n1863 VSS.n1574 0.0115294
R2639 VSS.n1584 VSS.n1578 0.0115294
R2640 VSS.n1643 VSS.n1642 0.0115294
R2641 VSS.n1724 VSS.n1716 0.0115294
R2642 VSS.n1809 VSS.n1808 0.0115294
R2643 VSS.n1761 VSS.n1760 0.0115294
R2644 VSS.n1224 VSS.n1160 0.0115294
R2645 VSS.n1240 VSS.n1220 0.0115294
R2646 VSS.n1250 VSS.n1214 0.0115294
R2647 VSS.n1317 VSS.n1278 0.0115294
R2648 VSS.n1328 VSS.n1327 0.0115294
R2649 VSS.n1961 VSS.n1306 0.0115294
R2650 VSS.n70 VSS.n69 0.0115294
R2651 VSS.n1101 VSS.n40 0.0115294
R2652 VSS.n1104 VSS.n25 0.0115294
R2653 VSS.n2081 VSS.n2080 0.0115294
R2654 VSS.n2095 VSS.n2094 0.0115294
R2655 VSS.n2108 VSS.n2107 0.0115294
R2656 VSS.n471 VSS.n470 0.0114649
R2657 VSS.n319 VSS.n318 0.0114649
R2658 VSS.n543 VSS.n522 0.0114649
R2659 VSS.n1458 VSS.n1457 0.0114167
R2660 VSS.n1283 VSS.n1199 0.0109167
R2661 VSS.n1786 VSS.n1774 0.0109167
R2662 VSS.n800 VSS.n799 0.0109167
R2663 VSS.n328 VSS.n327 0.0109167
R2664 VSS.n340 VSS.n339 0.0109167
R2665 VSS.n707 VSS.n701 0.0109167
R2666 VSS VSS.n1868 0.0105
R2667 VSS.n1412 VSS.n1411 0.0104679
R2668 VSS.n1656 VSS.n1638 0.0104679
R2669 VSS.n2011 VSS.n1192 0.0104679
R2670 VSS.n1568 VSS.n1486 0.0104167
R2671 VSS.n1021 VSS.n1020 0.0102656
R2672 VSS.n1018 VSS.n1012 0.0102656
R2673 VSS.n172 VSS.n166 0.0102656
R2674 VSS.n2193 VSS 0.01025
R2675 VSS.n1907 VSS.n1906 0.0100833
R2676 VSS.n1792 VSS.n1791 0.01
R2677 VSS.n233 VSS.n232 0.00993343
R2678 VSS.n1942 VSS.n1941 0.00991667
R2679 VSS.n77 VSS.n76 0.00983333
R2680 VSS.n1829 VSS.n1662 0.0098203
R2681 VSS.n1903 VSS.n1461 0.0098203
R2682 VSS.n1280 VSS.n1275 0.0098203
R2683 VSS.n2069 VSS.n2068 0.0098203
R2684 VSS.n1934 VSS.n1371 0.00969118
R2685 VSS.n1925 VSS.n1924 0.00969118
R2686 VSS.n1419 VSS.n1418 0.00969118
R2687 VSS.n1526 VSS.n1497 0.00969118
R2688 VSS.n1531 VSS.n1492 0.00969118
R2689 VSS.n1552 VSS.n1550 0.00969118
R2690 VSS.n1860 VSS.n1576 0.00969118
R2691 VSS.n1851 VSS.n1850 0.00969118
R2692 VSS.n1653 VSS.n1652 0.00969118
R2693 VSS.n1723 VSS.n1663 0.00969118
R2694 VSS.n1729 VSS.n1713 0.00969118
R2695 VSS.n1751 VSS.n1750 0.00969118
R2696 VSS.n1231 VSS.n1230 0.00969118
R2697 VSS.n1242 VSS.n1241 0.00969118
R2698 VSS.n1252 VSS.n1251 0.00969118
R2699 VSS.n1994 VSS.n1993 0.00969118
R2700 VSS.n1324 VSS.n1314 0.00969118
R2701 VSS.n1973 VSS.n1972 0.00969118
R2702 VSS.n59 VSS.n58 0.00969118
R2703 VSS.n1110 VSS.n1109 0.00969118
R2704 VSS.n1139 VSS.n1138 0.00969118
R2705 VSS.n4 VSS.n3 0.00969118
R2706 VSS.n2083 VSS.n2082 0.00969118
R2707 VSS.n2097 VSS.n2096 0.00969118
R2708 VSS.n1131 VSS.n1130 0.00961458
R2709 VSS.n2042 VSS.n1149 0.00961458
R2710 VSS.n1266 VSS.n1198 0.00961458
R2711 VSS.n1895 VSS.n1472 0.00961458
R2712 VSS.n2185 VSS.n2184 0.00961458
R2713 VSS.n999 VSS.n998 0.00961458
R2714 VSS.n152 VSS.n151 0.00961458
R2715 VSS.n285 VSS.n284 0.00961458
R2716 VSS.n444 VSS.n443 0.00961458
R2717 VSS.n603 VSS.n602 0.00961458
R2718 VSS.n72 VSS.n71 0.00945904
R2719 VSS.n1119 VSS.n37 0.00945904
R2720 VSS.n1118 VSS.n39 0.00945904
R2721 VSS.n1108 VSS.n1107 0.00945904
R2722 VSS.n1106 VSS.n1103 0.00945904
R2723 VSS.n1141 VSS.n24 0.00945904
R2724 VSS.n2058 VSS.n10 0.00945904
R2725 VSS.n1817 VSS.n1707 0.00927193
R2726 VSS VSS.n1363 0.009
R2727 VSS.n1007 VSS.n1006 0.00896354
R2728 VSS.n1451 VSS.n1450 0.0083125
R2729 VSS.n1000 VSS.n999 0.0083125
R2730 VSS.n294 VSS.n279 0.0083125
R2731 VSS.n428 VSS.n427 0.0083125
R2732 VSS.n260 VSS.n259 0.0083125
R2733 VSS.n571 VSS.n570 0.0083125
R2734 VSS.n595 VSS.n594 0.0083125
R2735 VSS.n661 VSS.n655 0.0083125
R2736 VSS.n1772 VSS.n1770 0.00801655
R2737 VSS.n1287 VSS.n1286 0.008
R2738 VSS.n1020 VSS.n1019 0.00766146
R2739 VSS.n923 VSS.n915 0.00766146
R2740 VSS.n1562 VSS.n1561 0.00707895
R2741 VSS.n1873 VSS.n1872 0.00707895
R2742 VSS.n1677 VSS.n1676 0.00701042
R2743 VSS.n1699 VSS.n1689 0.00701042
R2744 VSS.n2130 VSS.n2129 0.00701042
R2745 VSS.n316 VSS.n315 0.00701042
R2746 VSS.n496 VSS.n495 0.00701042
R2747 VSS.n512 VSS.n243 0.00701042
R2748 VSS.n530 VSS.n529 0.00701042
R2749 VSS.n542 VSS.n541 0.00701042
R2750 VSS.n559 VSS.n558 0.00701042
R2751 VSS.n1364 VSS 0.00659221
R2752 VSS.n1832 VSS.n1659 0.00658333
R2753 VSS.n1049 VSS.n1042 0.00635938
R2754 VSS.n866 VSS.n865 0.00635938
R2755 VSS.n1262 VSS.n1261 0.00570833
R2756 VSS.n1741 VSS.n1705 0.00570833
R2757 VSS.n2167 VSS.n2165 0.00570833
R2758 VSS.n2182 VSS.n2181 0.00570833
R2759 VSS.n410 VSS.n404 0.00570833
R2760 VSS.n488 VSS.n487 0.00570833
R2761 VSS.n963 VSS.n962 0.00505729
R2762 VSS.n1073 VSS.n78 0.00493396
R2763 VSS.n1075 VSS.n78 0.00493396
R2764 VSS.n1064 VSS.n1063 0.00489326
R2765 VSS.n365 VSS.n350 0.00488596
R2766 VSS.n1911 VSS.n1910 0.00488596
R2767 VSS.n1606 VSS.n1605 0.00476179
R2768 VSS.n843 VSS.n842 0.00476179
R2769 VSS.n823 VSS.n822 0.00476179
R2770 VSS.n869 VSS.n868 0.00476179
R2771 VSS.n885 VSS.n884 0.00476179
R2772 VSS.n926 VSS.n925 0.00476179
R2773 VSS.n949 VSS.n948 0.00476179
R2774 VSS.n980 VSS.n979 0.00476179
R2775 VSS.n784 VSS.n783 0.00476179
R2776 VSS.n2155 VSS.n2144 0.00451955
R2777 VSS.n1983 VSS.n1293 0.00440625
R2778 VSS.n1560 VSS.n1475 0.00440625
R2779 VSS.n1565 VSS.n1563 0.00440625
R2780 VSS.n1820 VSS.n1704 0.00440625
R2781 VSS.n2168 VSS.n2167 0.00440625
R2782 VSS.n781 VSS.n776 0.00440625
R2783 VSS.n685 VSS.n677 0.00440625
R2784 VSS.n1168 VSS.n1167 0.00429297
R2785 VSS.n298 VSS.n297 0.00390422
R2786 VSS.n1775 VSS.n1768 0.00389678
R2787 VSS.n453 VSS.n452 0.00386759
R2788 VSS.n642 VSS.n641 0.00386759
R2789 VSS.n724 VSS.n723 0.00386759
R2790 VSS.n1079 VSS.n1078 0.00386759
R2791 VSS.n894 VSS.n157 0.00386759
R2792 VSS.n155 VSS.n154 0.00386759
R2793 VSS.n763 VSS.n762 0.00386759
R2794 VSS.n204 VSS.n203 0.00386759
R2795 VSS.n191 VSS.n190 0.00386759
R2796 VSS.n175 VSS.n174 0.00386759
R2797 VSS.n93 VSS.n92 0.00386759
R2798 VSS.n131 VSS.n130 0.00386759
R2799 VSS.n803 VSS.n802 0.00386759
R2800 VSS.n840 VSS.n835 0.00375521
R2801 VSS.n2188 VSS.n2187 0.00362372
R2802 VSS.n997 VSS.n996 0.00340722
R2803 VSS.n996 VSS.n995 0.00340722
R2804 VSS.n994 VSS.n993 0.00340722
R2805 VSS.n993 VSS.n992 0.00340722
R2806 VSS.n991 VSS.n990 0.00340722
R2807 VSS.n990 VSS.n989 0.00340722
R2808 VSS.n988 VSS.n987 0.00340722
R2809 VSS.n987 VSS.n986 0.00340722
R2810 VSS.n985 VSS.n984 0.00340722
R2811 VSS.n984 VSS.n983 0.00340722
R2812 VSS.n982 VSS.n981 0.00340722
R2813 VSS.n981 VSS.n955 0.00340722
R2814 VSS.n954 VSS.n953 0.00340722
R2815 VSS.n953 VSS.n952 0.00340722
R2816 VSS.n951 VSS.n950 0.00340722
R2817 VSS.n950 VSS.n932 0.00340722
R2818 VSS.n931 VSS.n930 0.00340722
R2819 VSS.n930 VSS.n929 0.00340722
R2820 VSS.n928 VSS.n927 0.00340722
R2821 VSS.n927 VSS.n888 0.00340722
R2822 VSS.n887 VSS.n886 0.00340722
R2823 VSS.n886 VSS.n872 0.00340722
R2824 VSS.n871 VSS.n870 0.00340722
R2825 VSS.n870 VSS.n852 0.00340722
R2826 VSS.n851 VSS.n850 0.00340722
R2827 VSS.n850 VSS.n849 0.00340722
R2828 VSS.n848 VSS.n847 0.00340722
R2829 VSS.n847 VSS.n846 0.00340722
R2830 VSS.n845 VSS.n844 0.00340722
R2831 VSS.n844 VSS.n826 0.00340722
R2832 VSS.n825 VSS.n824 0.00340722
R2833 VSS.n824 VSS.n809 0.00340722
R2834 VSS.n808 VSS.n807 0.00340722
R2835 VSS.n807 VSS.n806 0.00340722
R2836 VSS.n805 VSS.n804 0.00340722
R2837 VSS.n804 VSS.n787 0.00340722
R2838 VSS.n786 VSS.n785 0.00340722
R2839 VSS.n785 VSS.n767 0.00340722
R2840 VSS.n766 VSS.n765 0.00340722
R2841 VSS.n765 VSS.n764 0.00340722
R2842 VSS.n321 VSS.n300 0.00340722
R2843 VSS.n322 VSS.n321 0.00340722
R2844 VSS.n344 VSS.n323 0.00340722
R2845 VSS.n345 VSS.n344 0.00340722
R2846 VSS.n367 VSS.n346 0.00340722
R2847 VSS.n368 VSS.n367 0.00340722
R2848 VSS.n392 VSS.n369 0.00340722
R2849 VSS.n393 VSS.n392 0.00340722
R2850 VSS.n420 VSS.n394 0.00340722
R2851 VSS.n421 VSS.n420 0.00340722
R2852 VSS.n447 VSS.n422 0.00340722
R2853 VSS.n448 VSS.n447 0.00340722
R2854 VSS.n454 VSS.n449 0.00340722
R2855 VSS.n455 VSS.n454 0.00340722
R2856 VSS.n464 VSS.n456 0.00340722
R2857 VSS.n465 VSS.n464 0.00340722
R2858 VSS.n477 VSS.n466 0.00340722
R2859 VSS.n477 VSS.n476 0.00340722
R2860 VSS.n475 VSS.n474 0.00340722
R2861 VSS.n474 VSS.n473 0.00340722
R2862 VSS.n516 VSS.n236 0.00340722
R2863 VSS.n517 VSS.n516 0.00340722
R2864 VSS.n545 VSS.n518 0.00340722
R2865 VSS.n546 VSS.n545 0.00340722
R2866 VSS.n574 VSS.n547 0.00340722
R2867 VSS.n575 VSS.n574 0.00340722
R2868 VSS.n583 VSS.n576 0.00340722
R2869 VSS.n584 VSS.n583 0.00340722
R2870 VSS.n636 VSS.n585 0.00340722
R2871 VSS.n637 VSS.n636 0.00340722
R2872 VSS.n643 VSS.n638 0.00340722
R2873 VSS.n644 VSS.n643 0.00340722
R2874 VSS.n666 VSS.n645 0.00340722
R2875 VSS.n667 VSS.n666 0.00340722
R2876 VSS.n695 VSS.n668 0.00340722
R2877 VSS.n696 VSS.n695 0.00340722
R2878 VSS.n718 VSS.n697 0.00340722
R2879 VSS.n719 VSS.n718 0.00340722
R2880 VSS.n729 VSS.n720 0.00340722
R2881 VSS.n729 VSS.n728 0.00340722
R2882 VSS.n727 VSS.n726 0.00340722
R2883 VSS.n726 VSS.n725 0.00340722
R2884 VSS.n1093 VSS.n48 0.00310417
R2885 VSS.n1912 VSS.n1397 0.00310417
R2886 VSS.n1507 VSS.n1503 0.00310417
R2887 VSS.n1006 VSS.n1000 0.00310417
R2888 VSS.n364 VSS.n363 0.00310417
R2889 VSS.n387 VSS.n381 0.00310417
R2890 VSS.n2073 VSS.n1 0.00300444
R2891 VSS.n2074 VSS.n2073 0.00300444
R2892 VSS.n2087 VSS.n2075 0.00300444
R2893 VSS.n2088 VSS.n2087 0.00300444
R2894 VSS.n2101 VSS.n2089 0.00300444
R2895 VSS.n2102 VSS.n2101 0.00300444
R2896 VSS.n2119 VSS.n2103 0.00300444
R2897 VSS.n2205 VSS.n2204 0.00300444
R2898 VSS.n2204 VSS.n2194 0.00300444
R2899 VSS.n1235 VSS.n1234 0.003
R2900 VSS.n1237 VSS.n1235 0.003
R2901 VSS.n1236 VSS.n1217 0.003
R2902 VSS.n1217 VSS.n1216 0.003
R2903 VSS.n2007 VSS 0.003
R2904 VSS.n1286 VSS 0.003
R2905 VSS.n1288 VSS.n1287 0.003
R2906 VSS.n1990 VSS.n1288 0.003
R2907 VSS.n1332 VSS.n1331 0.003
R2908 VSS.n1969 VSS.n1332 0.003
R2909 VSS.n1968 VSS.n1967 0.003
R2910 VSS.n1967 VSS.n1966 0.003
R2911 VSS.n1959 VSS.n1335 0.003
R2912 VSS.n1363 VSS.n1335 0.003
R2913 VSS.n1365 VSS.n1364 0.003
R2914 VSS.n1942 VSS.n1365 0.003
R2915 VSS.n1941 VSS.n1366 0.003
R2916 VSS.n1376 VSS.n1366 0.003
R2917 VSS.n1930 VSS.n1381 0.003
R2918 VSS.n1930 VSS.n1929 0.003
R2919 VSS.n1405 VSS.n1382 0.003
R2920 VSS.n1457 VSS.n1400 0.003
R2921 VSS.n1538 VSS.n1537 0.003
R2922 VSS.n1540 VSS.n1539 0.003
R2923 VSS.n1539 VSS.n1488 0.003
R2924 VSS.n1870 VSS.n1568 0.003
R2925 VSS.n1870 VSS.n1869 0.003
R2926 VSS.n1868 VSS.n1569 0.003
R2927 VSS.n1856 VSS.n1855 0.003
R2928 VSS.n1646 VSS.n1582 0.003
R2929 VSS.n1647 VSS.n1646 0.003
R2930 VSS.n1695 VSS.n1659 0.003
R2931 VSS.n1832 VSS.n1831 0.003
R2932 VSS.n1831 VSS.n1660 0.003
R2933 VSS.n1754 VSS.n1710 0.003
R2934 VSS.n1755 VSS.n1754 0.003
R2935 VSS.n1757 VSS.n1756 0.003
R2936 VSS.n1793 VSS.n1792 0.003
R2937 VSS.n1077 VSS.n1076 0.003
R2938 VSS.n1077 VSS.n77 0.003
R2939 VSS.n76 VSS.n55 0.003
R2940 VSS.n1115 VSS.n1114 0.003
R2941 VSS.n1099 VSS.n1097 0.003
R2942 VSS.n1099 VSS.n27 0.003
R2943 VSS.n1988 VSS.n1289 0.00283333
R2944 VSS.n1312 VSS.n1311 0.00283333
R2945 VSS.n1945 VSS.n1355 0.00269298
R2946 VSS.n1361 VSS.n1337 0.00269298
R2947 VSS.n1537 VSS.n1494 0.00266667
R2948 VSS.n1424 VSS.n1405 0.00258333
R2949 VSS.n1406 VSS.n1403 0.00258333
R2950 VSS.n1458 VSS.n1456 0.00258333
R2951 VSS VSS.n1400 0.00258333
R2952 VSS.n1135 VSS.n1134 0.00258333
R2953 VSS.n28 VSS.n13 0.00258333
R2954 VSS.n2055 VSS.n2054 0.00258333
R2955 VSS.n1379 VSS.n1378 0.00257353
R2956 VSS.n1380 VSS.n1374 0.00257353
R2957 VSS.n1928 VSS.n1375 0.00257353
R2958 VSS.n1927 VSS.n1926 0.00257353
R2959 VSS.n1422 VSS.n1408 0.00257353
R2960 VSS.n1421 VSS.n1420 0.00257353
R2961 VSS.n1459 VSS.n1402 0.00257353
R2962 VSS.n1905 VSS.n1904 0.00257353
R2963 VSS.n1525 VSS.n1524 0.00257353
R2964 VSS.n1498 VSS.n1495 0.00257353
R2965 VSS.n1496 VSS.n1493 0.00257353
R2966 VSS.n1542 VSS.n1541 0.00257353
R2967 VSS.n1554 VSS.n1553 0.00257353
R2968 VSS.n1555 VSS.n1484 0.00257353
R2969 VSS.n1570 VSS.n1482 0.00257353
R2970 VSS.n1867 VSS.n1866 0.00257353
R2971 VSS.n1601 VSS.n1600 0.00257353
R2972 VSS.n1602 VSS.n1579 0.00257353
R2973 VSS.n1854 VSS.n1580 0.00257353
R2974 VSS.n1853 VSS.n1852 0.00257353
R2975 VSS.n1645 VSS.n1644 0.00257353
R2976 VSS.n1651 VSS.n1650 0.00257353
R2977 VSS.n1834 VSS.n1657 0.00257353
R2978 VSS.n1833 VSS.n1658 0.00257353
R2979 VSS.n1719 VSS.n1661 0.00257353
R2980 VSS.n1725 VSS.n1722 0.00257353
R2981 VSS.n1812 VSS.n1711 0.00257353
R2982 VSS.n1811 VSS.n1810 0.00257353
R2983 VSS.n1753 VSS.n1752 0.00257353
R2984 VSS.n1759 VSS.n1758 0.00257353
R2985 VSS.n1223 VSS.n1162 0.00257353
R2986 VSS.n1233 VSS.n1232 0.00257353
R2987 VSS.n1239 VSS.n1238 0.00257353
R2988 VSS.n1222 VSS.n1215 0.00257353
R2989 VSS.n1249 VSS.n1213 0.00257353
R2990 VSS.n1254 VSS.n1253 0.00257353
R2991 VSS.n2010 VSS.n2009 0.00257353
R2992 VSS.n1279 VSS.n1194 0.00257353
R2993 VSS.n1992 VSS.n1991 0.00257353
R2994 VSS.n1319 VSS.n1282 0.00257353
R2995 VSS.n1320 VSS.n1313 0.00257353
R2996 VSS.n1330 VSS.n1329 0.00257353
R2997 VSS.n1971 VSS.n1970 0.00257353
R2998 VSS.n1333 VSS.n1308 0.00257353
R2999 VSS.n68 VSS.n67 0.00257353
R3000 VSS.n60 VSS.n41 0.00257353
R3001 VSS.n1113 VSS.n42 0.00257353
R3002 VSS.n1112 VSS.n1111 0.00257353
R3003 VSS.n1098 VSS.n26 0.00257353
R3004 VSS.n1137 VSS.n1136 0.00257353
R3005 VSS.n2071 VSS.n2070 0.00257353
R3006 VSS.n2077 VSS.n2076 0.00257353
R3007 VSS.n2079 VSS.n2078 0.00257353
R3008 VSS.n2091 VSS.n2090 0.00257353
R3009 VSS.n2093 VSS.n2092 0.00257353
R3010 VSS.n2105 VSS.n2104 0.00257353
R3011 VSS.n1966 VSS.n1959 0.0025
R3012 VSS.n1906 VSS.n1401 0.0025
R3013 VSS.n1521 VSS.n1499 0.0025
R3014 VSS.n1096 VSS.n43 0.0025
R3015 VSS.n1756 VSS.n1747 0.00241667
R3016 VSS.n1793 VSS.n1767 0.00241667
R3017 VSS.n1937 VSS.n1368 0.00233824
R3018 VSS.n1372 VSS.n1370 0.00233824
R3019 VSS.n1922 VSS.n1387 0.00233824
R3020 VSS.n1933 VSS.n1932 0.00233824
R3021 VSS.n1414 VSS.n1385 0.00233824
R3022 VSS.n1413 VSS.n1412 0.00233824
R3023 VSS.n1533 VSS.n1530 0.00233824
R3024 VSS.n1547 VSS.n1546 0.00233824
R3025 VSS.n1885 VSS.n1481 0.00233824
R3026 VSS.n1462 VSS.n1461 0.00233824
R3027 VSS.n1535 VSS.n1534 0.00233824
R3028 VSS.n1545 VSS.n1490 0.00233824
R3029 VSS.n1573 VSS.n1572 0.00233824
R3030 VSS.n1577 VSS.n1575 0.00233824
R3031 VSS.n1848 VSS.n1587 0.00233824
R3032 VSS.n1859 VSS.n1858 0.00233824
R3033 VSS.n1640 VSS.n1585 0.00233824
R3034 VSS.n1654 VSS.n1638 0.00233824
R3035 VSS.n1718 VSS.n1715 0.00233824
R3036 VSS.n1806 VSS.n1805 0.00233824
R3037 VSS.n1763 VSS.n1749 0.00233824
R3038 VSS.n1829 VSS.n1828 0.00233824
R3039 VSS.n1728 VSS.n1727 0.00233824
R3040 VSS.n1731 VSS.n1714 0.00233824
R3041 VSS.n2030 VSS.n2029 0.00233824
R3042 VSS.n1228 VSS.n1227 0.00233824
R3043 VSS.n1246 VSS.n1244 0.00233824
R3044 VSS.n1226 VSS.n1225 0.00233824
R3045 VSS.n1247 VSS.n1218 0.00233824
R3046 VSS.n1192 VSS.n1191 0.00233824
R3047 VSS.n1318 VSS.n1316 0.00233824
R3048 VSS.n1975 VSS.n1303 0.00233824
R3049 VSS.n1962 VSS.n1960 0.00233824
R3050 VSS.n1280 VSS.n1276 0.00233824
R3051 VSS.n1323 VSS.n1322 0.00233824
R3052 VSS.n1315 VSS.n1304 0.00233824
R3053 VSS.n1117 VSS.n38 0.00233824
R3054 VSS.n1105 VSS.n1102 0.00233824
R3055 VSS.n1140 VSS.n11 0.00233824
R3056 VSS.n219 VSS.n215 0.00233824
R3057 VSS.n224 VSS.n222 0.00233824
R3058 VSS.n2115 VSS.n2114 0.00233824
R3059 VSS.n2069 VSS.n5 0.00233824
R3060 VSS.n2085 VSS.n2084 0.00233824
R3061 VSS.n2099 VSS.n2098 0.00233824
R3062 VSS.n1177 VSS.n1176 0.00233333
R3063 VSS.n2026 VSS.n1163 0.00233333
R3064 VSS.n2025 VSS.n1164 0.00233333
R3065 VSS.n1073 VSS.n1072 0.00227358
R3066 VSS.n2121 VSS.n2120 0.00225311
R3067 VSS.n1603 VSS.n1581 0.00225
R3068 VSS.n2154 VSS.n2146 0.00218919
R3069 VSS.n2161 VSS.n2142 0.00218919
R3070 VSS.n2075 VSS.n2074 0.00216963
R3071 VSS.n2089 VSS.n2088 0.00216963
R3072 VSS.n2103 VSS.n2102 0.00216963
R3073 VSS.n1234 VSS.n1164 0.00216667
R3074 VSS.n1237 VSS.n1236 0.00216667
R3075 VSS.n1990 VSS.n1989 0.00216667
R3076 VSS.n1969 VSS.n1968 0.00216667
R3077 VSS.n1381 VSS.n1376 0.00216667
R3078 VSS.n1929 VSS.n1382 0.00216667
R3079 VSS.n1423 VSS.n1407 0.00216667
R3080 VSS.n1523 VSS.n1522 0.00216667
R3081 VSS.n1540 VSS.n1538 0.00216667
R3082 VSS.n1855 VSS.n1582 0.00216667
R3083 VSS.n1649 VSS.n1647 0.00216667
R3084 VSS.n1648 VSS.n1635 0.00216667
R3085 VSS.n1836 VSS.n1835 0.00216667
R3086 VSS.n1813 VSS.n1710 0.00216667
R3087 VSS.n1757 VSS.n1755 0.00216667
R3088 VSS.n1114 VSS.n1097 0.00216667
R3089 VSS.n1135 VSS.n27 0.00216667
R3090 VSS.n1074 VSS.n79 0.0021514
R3091 VSS.n1556 VSS.n1485 0.00208333
R3092 VSS.n1881 VSS.n1880 0.00208333
R3093 VSS.n1599 VSS.n1598 0.00208333
R3094 VSS.n1791 VSS 0.00208333
R3095 VSS.n1331 VSS.n1310 0.002
R3096 VSS.n1721 VSS.n1708 0.002
R3097 VSS.n1814 VSS.n1709 0.002
R3098 VSS.n2157 VSS.n2156 0.00196875
R3099 VSS.n2159 VSS.n2158 0.00196875
R3100 VSS.n2124 VSS.n2123 0.00196875
R3101 VSS.n2126 VSS.n2125 0.00196875
R3102 VSS.n1257 VSS.n1255 0.00191667
R3103 VSS.n1256 VSS.n1195 0.00191667
R3104 VSS.n1695 VSS 0.00191667
R3105 VSS.n66 VSS.n64 0.00183333
R3106 VSS.n1180 VSS.n1153 0.00180208
R3107 VSS.n1360 VSS.n1339 0.00180208
R3108 VSS.n1947 VSS.n1946 0.00180208
R3109 VSS.n2153 VSS.n2152 0.00180208
R3110 VSS.n2162 VSS.n2140 0.00180208
R3111 VSS.n1019 VSS.n1018 0.00180208
R3112 VSS.n352 VSS.n351 0.00180208
R3113 VSS.n64 VSS.n55 0.00166667
R3114 VSS.n66 VSS.n65 0.00166667
R3115 VSS.n1255 VSS.n1212 0.00158333
R3116 VSS.n1257 VSS.n1256 0.00158333
R3117 VSS.n2008 VSS.n1195 0.00158333
R3118 VSS VSS.n1694 0.00158333
R3119 VSS.n1721 VSS.n1720 0.0015
R3120 VSS.n1709 VSS.n1708 0.0015
R3121 VSS.n1814 VSS.n1813 0.0015
R3122 VSS.n1557 VSS.n1556 0.00141667
R3123 VSS.n1881 VSS.n1485 0.00141667
R3124 VSS.n1880 VSS.n1486 0.00141667
R3125 VSS.n1598 VSS.n1569 0.00141667
R3126 VSS.n1604 VSS.n1599 0.00141667
R3127 VSS.n1649 VSS.n1648 0.00133333
R3128 VSS.n1836 VSS.n1635 0.00133333
R3129 VSS.n1835 VSS.n1636 0.00133333
R3130 VSS.n2120 VSS.n2119 0.00125133
R3131 VSS.n1557 VSS.n1488 0.00125
R3132 VSS.n1604 VSS.n1603 0.00125
R3133 VSS.n1856 VSS.n1581 0.00125
R3134 VSS.n1176 VSS.n1163 0.00116667
R3135 VSS.n2026 VSS.n2025 0.00116667
R3136 VSS.n1720 VSS.n1660 0.00116667
R3137 VSS.n1069 VSS.n1065 0.0011215
R3138 VSS.n1216 VSS.n1212 0.00108333
R3139 VSS.n1869 VSS 0.00108333
R3140 VSS.n1767 VSS.n1747 0.00108333
R3141 VSS.n1175 VSS 0.001
R3142 VSS.n1499 VSS.n1401 0.001
R3143 VSS.n1523 VSS.n1521 0.001
R3144 VSS.n65 VSS.n43 0.001
R3145 VSS.n1115 VSS.n1096 0.001
R3146 VSS.n72 VSS.n57 0.000926621
R3147 VSS.n1119 VSS.n1118 0.000926621
R3148 VSS.n1107 VSS.n1106 0.000926621
R3149 VSS.n1141 VSS.n10 0.000926621
R3150 VSS.n1424 VSS.n1423 0.000916667
R3151 VSS.n1407 VSS.n1406 0.000916667
R3152 VSS.n1456 VSS.n1403 0.000916667
R3153 VSS.n1907 VSS 0.000916667
R3154 VSS.n1134 VSS.n28 0.000916667
R3155 VSS.n2055 VSS.n13 0.000916667
R3156 VSS.n1522 VSS.n1494 0.000833333
R3157 VSS.n1989 VSS.n1988 0.000666667
R3158 VSS.n1311 VSS.n1289 0.000666667
R3159 VSS.n1312 VSS.n1310 0.000666667
R3160 VDD.n32 VDD.n31 1340.43
R3161 VDD.n2990 VDD.n35 553.333
R3162 VDD.n721 VDD.t202 500.865
R3163 VDD.n721 VDD.t222 500.865
R3164 VDD.n1165 VDD.t39 500.865
R3165 VDD.n1165 VDD.t59 500.865
R3166 VDD.n354 VDD.t32 500.865
R3167 VDD.n354 VDD.t2 500.865
R3168 VDD.n73 VDD.t170 500.865
R3169 VDD.n73 VDD.t46 500.865
R3170 VDD.n744 VDD.n742 440.25
R3171 VDD.n744 VDD.n743 440.25
R3172 VDD.n929 VDD.n927 440.25
R3173 VDD.n929 VDD.n928 440.25
R3174 VDD.n574 VDD.n262 440.25
R3175 VDD.n574 VDD.n263 440.25
R3176 VDD.n116 VDD.n114 440.25
R3177 VDD.n116 VDD.n115 440.25
R3178 VDD.n2995 VDD.n4 426
R3179 VDD.n1074 VDD.t67 397.144
R3180 VDD.n814 VDD.t98 397.144
R3181 VDD.n156 VDD.t107 397.144
R3182 VDD.n515 VDD.t88 397.144
R3183 VDD.n1070 VDD.t82 394.462
R3184 VDD.n810 VDD.t64 394.462
R3185 VDD.n152 VDD.t73 394.462
R3186 VDD.n511 VDD.t91 394.462
R3187 VDD.n846 VDD.t119 391.623
R3188 VDD.n1050 VDD.t103 391.623
R3189 VDD.n647 VDD.t79 391.623
R3190 VDD.n539 VDD.t113 391.623
R3191 VDD.n857 VDD.t93 384.286
R3192 VDD.n1043 VDD.t109 384.286
R3193 VDD.n658 VDD.t101 384.286
R3194 VDD.n551 VDD.t61 384.286
R3195 VDD.n1126 VDD.t151 371
R3196 VDD.n1126 VDD.t214 371
R3197 VDD.n1206 VDD.t22 371
R3198 VDD.n1206 VDD.t221 371
R3199 VDD.n237 VDD.t128 371
R3200 VDD.n237 VDD.t197 371
R3201 VDD.n390 VDD.t137 371
R3202 VDD.n390 VDD.t131 371
R3203 VDD.n3019 VDD.n2 351
R3204 VDD.n1201 VDD.n788 331.765
R3205 VDD.n978 VDD.n970 331.765
R3206 VDD.n631 VDD.n134 331.765
R3207 VDD.n487 VDD.n385 331.765
R3208 VDD.n737 VDD.n726 328.236
R3209 VDD.n1201 VDD.n790 328.236
R3210 VDD.n922 VDD.n797 328.236
R3211 VDD.n1179 VDD.n909 328.236
R3212 VDD.n1163 VDD.n942 328.236
R3213 VDD.n1159 VDD.n942 328.236
R3214 VDD.n1150 VDD.n952 328.236
R3215 VDD.n1138 VDD.n956 328.236
R3216 VDD.n1121 VDD.n979 328.236
R3217 VDD.n106 VDD.n90 328.236
R3218 VDD.n131 VDD.n130 328.236
R3219 VDD.n131 VDD.n69 328.236
R3220 VDD.n209 VDD.n136 328.236
R3221 VDD.n209 VDD.n206 328.236
R3222 VDD.n587 VDD.n242 328.236
R3223 VDD.n580 VDD.n258 328.236
R3224 VDD.n576 VDD.n258 328.236
R3225 VDD.n353 VDD.n260 328.236
R3226 VDD.n504 VDD.n339 328.236
R3227 VDD.n504 VDD.n340 328.236
R3228 VDD.n491 VDD.n384 328.236
R3229 VDD.n466 VDD.n454 328.236
R3230 VDD.n737 VDD.n724 324.707
R3231 VDD.n747 VDD.n724 324.707
R3232 VDD.n747 VDD.n722 324.707
R3233 VDD.n1246 VDD.n722 324.707
R3234 VDD.n1246 VDD.n723 324.707
R3235 VDD.n1242 VDD.n723 324.707
R3236 VDD.n1242 VDD.n750 324.707
R3237 VDD.n1235 VDD.n750 324.707
R3238 VDD.n1235 VDD.n760 324.707
R3239 VDD.n1232 VDD.n760 324.707
R3240 VDD.n1232 VDD.n763 324.707
R3241 VDD.n1226 VDD.n763 324.707
R3242 VDD.n1226 VDD.n770 324.707
R3243 VDD.n1222 VDD.n770 324.707
R3244 VDD.n1222 VDD.n772 324.707
R3245 VDD.n1215 VDD.n772 324.707
R3246 VDD.n1215 VDD.n782 324.707
R3247 VDD.n1211 VDD.n782 324.707
R3248 VDD.n1211 VDD.n783 324.707
R3249 VDD.n1205 VDD.n783 324.707
R3250 VDD.n797 VDD.n790 324.707
R3251 VDD.n1179 VDD.n910 324.707
R3252 VDD.n1175 VDD.n910 324.707
R3253 VDD.n1175 VDD.n926 324.707
R3254 VDD.n1150 VDD.n1149 324.707
R3255 VDD.n1149 VDD.n955 324.707
R3256 VDD.n1145 VDD.n955 324.707
R3257 VDD.n1138 VDD.n968 324.707
R3258 VDD.n1134 VDD.n968 324.707
R3259 VDD.n97 VDD.n92 324.707
R3260 VDD.n106 VDD.n92 324.707
R3261 VDD.n112 VDD.n90 324.707
R3262 VDD.n91 VDD.n72 324.707
R3263 VDD.n126 VDD.n72 324.707
R3264 VDD.n130 VDD.n70 324.707
R3265 VDD.n627 VDD.n136 324.707
R3266 VDD.n604 VDD.n207 324.707
R3267 VDD.n604 VDD.n212 324.707
R3268 VDD.n241 VDD.n212 324.707
R3269 VDD.n590 VDD.n241 324.707
R3270 VDD.n590 VDD.n242 324.707
R3271 VDD.n580 VDD.n245 324.707
R3272 VDD.n357 VDD.n353 324.707
R3273 VDD.n357 VDD.n350 324.707
R3274 VDD.n363 VDD.n350 324.707
R3275 VDD.n363 VDD.n347 324.707
R3276 VDD.n347 VDD.n341 324.707
R3277 VDD.n373 VDD.n341 324.707
R3278 VDD.n500 VDD.n376 324.707
R3279 VDD.n733 VDD.n726 321.176
R3280 VDD.n1163 VDD.n926 321.176
R3281 VDD.n1159 VDD.n943 321.176
R3282 VDD.n952 VDD.n943 321.176
R3283 VDD.n1145 VDD.n956 321.176
R3284 VDD.n1134 VDD.n970 321.176
R3285 VDD.n1125 VDD.n978 321.176
R3286 VDD.n112 VDD.n91 321.176
R3287 VDD.n126 VDD.n70 321.176
R3288 VDD.n632 VDD.n69 321.176
R3289 VDD.n627 VDD.n134 321.176
R3290 VDD.n608 VDD.n206 321.176
R3291 VDD.n608 VDD.n207 321.176
R3292 VDD.n587 VDD.n245 321.176
R3293 VDD.n373 VDD.n339 321.176
R3294 VDD.n500 VDD.n340 321.176
R3295 VDD.n491 VDD.n376 321.176
R3296 VDD.n487 VDD.n384 321.176
R3297 VDD.n462 VDD.n385 321.176
R3298 VDD.n462 VDD.n454 321.176
R3299 VDD.n466 VDD.n460 321.176
R3300 VDD.n922 VDD.n909 317.647
R3301 VDD.n1125 VDD.n979 317.647
R3302 VDD.n1121 VDD.n983 317.647
R3303 VDD.n632 VDD.n631 317.647
R3304 VDD.n576 VDD.n260 317.647
R3305 VDD.n1205 VDD.n788 314.118
R3306 VDD.n987 VDD.n985 308.598
R3307 VDD.n987 VDD.n986 308.598
R3308 VDD.n794 VDD.n792 308.598
R3309 VDD.n794 VDD.n793 308.598
R3310 VDD.n248 VDD.n246 308.598
R3311 VDD.n248 VDD.n247 308.598
R3312 VDD.n450 VDD.n448 308.598
R3313 VDD.n450 VDD.n449 308.598
R3314 VDD.n967 VDD.n965 304.122
R3315 VDD.n967 VDD.n966 304.122
R3316 VDD.n780 VDD.n778 304.122
R3317 VDD.n780 VDD.n779 304.122
R3318 VDD.n202 VDD.n198 304.122
R3319 VDD.n202 VDD.n199 304.122
R3320 VDD.n493 VDD.n381 304.122
R3321 VDD.n493 VDD.n382 304.122
R3322 VDD.n1157 VDD.n945 302.438
R3323 VDD.n1157 VDD.n946 302.438
R3324 VDD.n758 VDD.n756 302.438
R3325 VDD.n758 VDD.n757 302.438
R3326 VDD.n78 VDD.n75 302.438
R3327 VDD.n78 VDD.n76 302.438
R3328 VDD.n346 VDD.n344 302.438
R3329 VDD.n346 VDD.n345 302.438
R3330 VDD.t232 VDD.n3 258.856
R3331 VDD VDD.n2993 242.981
R3332 VDD.n284 VDD.t248 208.607
R3333 VDD.n935 VDD.t252 208.013
R3334 VDD.n1256 VDD.t247 208.013
R3335 VDD.n271 VDD.t244 208.013
R3336 VDD.n714 VDD.t243 206.459
R3337 VDD.n85 VDD.t258 206.459
R3338 VDD.n1014 VDD.t259 201.76
R3339 VDD.n683 VDD.t239 201.76
R3340 VDD.n2540 VDD.n2539 198.118
R3341 VDD.n2314 VDD.n2313 198.118
R3342 VDD.n2088 VDD.n2087 198.118
R3343 VDD.n1297 VDD.n1282 198.118
R3344 VDD.n2090 VDD.n2089 198.118
R3345 VDD.n2316 VDD.n2315 198.118
R3346 VDD.n2542 VDD.n2541 198.118
R3347 VDD.t230 VDD.n3017 188.965
R3348 VDD.n2795 VDD.n2794 185
R3349 VDD.n1334 VDD.n1333 185
R3350 VDD.n1323 VDD.n1322 185
R3351 VDD.n1312 VDD.n1311 185
R3352 VDD.n1300 VDD.n1299 185
R3353 VDD.n2814 VDD.n2813 185
R3354 VDD.n2814 VDD.n1298 185
R3355 VDD.n2833 VDD.n2832 185
R3356 VDD.n2833 VDD.n1298 185
R3357 VDD.n2852 VDD.n2851 185
R3358 VDD.n2852 VDD.n1298 185
R3359 VDD.n2872 VDD.n2871 185
R3360 VDD.n1296 VDD.n1295 185
R3361 VDD.n2776 VDD.n1345 185
R3362 VDD.n1893 VDD.n1892 185
R3363 VDD.n1851 VDD.n1850 185
R3364 VDD.n1942 VDD.n1941 185
R3365 VDD.n1961 VDD.n1838 185
R3366 VDD.n1979 VDD.n1978 185
R3367 VDD.n1998 VDD.n1803 185
R3368 VDD.n1997 VDD.n1806 185
R3369 VDD.n2001 VDD.n1805 185
R3370 VDD.n1804 VDD.n1789 185
R3371 VDD.n2037 VDD.n2036 185
R3372 VDD.n2034 VDD.n1788 185
R3373 VDD.n2064 VDD.n2063 185
R3374 VDD.n2066 VDD.n1770 185
R3375 VDD.n2085 VDD.n2084 185
R3376 VDD.n1760 VDD.n1759 185
R3377 VDD.n2091 VDD.n1758 185
R3378 VDD.n1732 VDD.n1731 185
R3379 VDD.n1717 VDD.n1716 185
R3380 VDD.n2168 VDD.n2167 185
R3381 VDD.n2187 VDD.n1704 185
R3382 VDD.n2205 VDD.n2204 185
R3383 VDD.n2224 VDD.n1669 185
R3384 VDD.n2223 VDD.n1672 185
R3385 VDD.n2227 VDD.n1671 185
R3386 VDD.n1670 VDD.n1655 185
R3387 VDD.n2263 VDD.n2262 185
R3388 VDD.n2260 VDD.n1654 185
R3389 VDD.n2290 VDD.n2289 185
R3390 VDD.n2292 VDD.n1636 185
R3391 VDD.n2311 VDD.n2310 185
R3392 VDD.n1626 VDD.n1625 185
R3393 VDD.n2317 VDD.n1624 185
R3394 VDD.n1598 VDD.n1597 185
R3395 VDD.n1583 VDD.n1582 185
R3396 VDD.n2394 VDD.n2393 185
R3397 VDD.n2413 VDD.n1570 185
R3398 VDD.n2431 VDD.n2430 185
R3399 VDD.n2450 VDD.n1535 185
R3400 VDD.n2449 VDD.n1538 185
R3401 VDD.n2453 VDD.n1537 185
R3402 VDD.n1536 VDD.n1521 185
R3403 VDD.n2489 VDD.n2488 185
R3404 VDD.n2486 VDD.n1520 185
R3405 VDD.n2516 VDD.n2515 185
R3406 VDD.n2518 VDD.n1502 185
R3407 VDD.n2537 VDD.n2536 185
R3408 VDD.n1492 VDD.n1491 185
R3409 VDD.n2543 VDD.n1490 185
R3410 VDD.n1464 VDD.n1463 185
R3411 VDD.n1449 VDD.n1448 185
R3412 VDD.n2620 VDD.n2619 185
R3413 VDD.n2639 VDD.n1436 185
R3414 VDD.n2657 VDD.n2656 185
R3415 VDD.n2676 VDD.n1401 185
R3416 VDD.n2675 VDD.n1404 185
R3417 VDD.n2679 VDD.n1403 185
R3418 VDD.n1402 VDD.n1387 185
R3419 VDD.n2715 VDD.n2714 185
R3420 VDD.n2712 VDD.n1386 185
R3421 VDD.n2742 VDD.n2741 185
R3422 VDD.n2744 VDD.n1368 185
R3423 VDD.n2768 VDD.n2767 185
R3424 VDD.n1357 VDD.n1356 185
R3425 VDD.n2637 VDD.n2636 185
R3426 VDD.n2617 VDD.n1447 185
R3427 VDD.n2592 VDD.n2591 185
R3428 VDD.n2571 VDD.n2570 185
R3429 VDD.n2658 VDD.n1416 185
R3430 VDD.n1475 VDD.n1474 185
R3431 VDD.n2411 VDD.n2410 185
R3432 VDD.n2391 VDD.n1581 185
R3433 VDD.n2366 VDD.n2365 185
R3434 VDD.n2345 VDD.n2344 185
R3435 VDD.n2432 VDD.n1550 185
R3436 VDD.n1609 VDD.n1608 185
R3437 VDD.n2185 VDD.n2184 185
R3438 VDD.n2165 VDD.n1715 185
R3439 VDD.n2140 VDD.n2139 185
R3440 VDD.n2119 VDD.n2118 185
R3441 VDD.n2206 VDD.n1684 185
R3442 VDD.n1743 VDD.n1742 185
R3443 VDD.n1959 VDD.n1958 185
R3444 VDD.n1939 VDD.n1849 185
R3445 VDD.n1914 VDD.n1913 185
R3446 VDD.n1980 VDD.n1818 185
R3447 VDD.n1891 VDD.n1866 185
R3448 VDD.n2969 VDD.n35 185
R3449 VDD.n3013 VDD.n2 185
R3450 VDD.n3017 VDD.n2 185
R3451 VDD.n714 VDD.t70 179.706
R3452 VDD.n85 VDD.t85 179.706
R3453 VDD.n935 VDD.t111 179.094
R3454 VDD.n1256 VDD.t105 179.094
R3455 VDD.n271 VDD.t117 179.094
R3456 VDD.n1016 VDD.t76 178.34
R3457 VDD.n685 VDD.t115 178.34
R3458 VDD.n284 VDD.t95 177.549
R3459 VDD.n730 VDD.n727 165.252
R3460 VDD.n730 VDD.n728 165.252
R3461 VDD.n915 VDD.n913 165.252
R3462 VDD.n915 VDD.n914 165.252
R3463 VDD.n95 VDD.n93 165.252
R3464 VDD.n95 VDD.n94 165.252
R3465 VDD.n253 VDD.n251 165.252
R3466 VDD.n253 VDD.n252 165.252
R3467 VDD.n2968 VDD.n2967 162.47
R3468 VDD.t35 VDD.n733 161.382
R3469 VDD.n97 VDD.t148 161.382
R3470 VDD.n959 VDD.n957 160.918
R3471 VDD.n959 VDD.n958 160.918
R3472 VDD.n769 VDD.n767 160.918
R3473 VDD.n769 VDD.n768 160.918
R3474 VDD.n139 VDD.n137 160.918
R3475 VDD.n139 VDD.n138 160.918
R3476 VDD.n338 VDD.n336 160.918
R3477 VDD.n338 VDD.n337 160.918
R3478 VDD.n3018 VDD 160.49
R3479 VDD.n3021 VDD.t231 152.88
R3480 VDD.n28 VDD.t233 152.879
R3481 VDD.n1016 VDD.n1015 152
R3482 VDD.n857 VDD.n856 152
R3483 VDD.n859 VDD.n858 152
R3484 VDD.n1045 VDD.n1044 152
R3485 VDD.n1043 VDD.n1042 152
R3486 VDD.n685 VDD.n684 152
R3487 VDD.n660 VDD.n659 152
R3488 VDD.n658 VDD.n657 152
R3489 VDD.n551 VDD.n550 152
R3490 VDD.n553 VDD.n552 152
R3491 VDD.n2965 VDD.t188 147.82
R3492 VDD.n1074 VDD.t254 134.986
R3493 VDD.n814 VDD.t249 134.986
R3494 VDD.n156 VDD.t241 134.986
R3495 VDD.n515 VDD.t245 134.986
R3496 VDD.n1070 VDD.t261 134.484
R3497 VDD.n810 VDD.t260 134.484
R3498 VDD.n152 VDD.t250 134.484
R3499 VDD.n511 VDD.t251 134.484
R3500 VDD.n847 VDD.t255 133.957
R3501 VDD.n1051 VDD.t262 133.957
R3502 VDD.n648 VDD.t246 133.957
R3503 VDD.n540 VDD.t253 133.957
R3504 VDD.n855 VDD.t240 133.5
R3505 VDD.n1041 VDD.t242 133.5
R3506 VDD.n656 VDD.t256 133.5
R3507 VDD.n548 VDD.t257 133.5
R3508 VDD.n1178 VDD.n924 133.459
R3509 VDD.n1137 VDD.n969 133.459
R3510 VDD.n108 VDD.n107 133.459
R3511 VDD.n133 VDD.n132 133.459
R3512 VDD.n210 VDD.n208 133.459
R3513 VDD.n579 VDD.n578 133.459
R3514 VDD.n352 VDD.n351 133.459
R3515 VDD.n503 VDD.n502 133.459
R3516 VDD.n736 VDD.n735 132.024
R3517 VDD.n1245 VDD.n749 132.024
R3518 VDD.n1234 VDD.n1233 132.024
R3519 VDD.t132 VDD.n762 132.024
R3520 VDD.n1225 VDD.n1224 132.024
R3521 VDD.n1223 VDD.n771 132.024
R3522 VDD.n1176 VDD.n925 132.024
R3523 VDD.n1148 VDD.t141 132.024
R3524 VDD.n1147 VDD.n1146 132.024
R3525 VDD.n110 VDD.n109 132.024
R3526 VDD.n244 VDD.n243 132.024
R3527 VDD.n361 VDD.n360 132.024
R3528 VDD.n501 VDD.n375 132.024
R3529 VDD.n954 VDD.n953 130.589
R3530 VDD.n629 VDD.n628 130.589
R3531 VDD.n374 VDD.t6 130.589
R3532 VDD.n464 VDD.n463 130.589
R3533 VDD.n1124 VDD.n1123 129.155
R3534 VDD.n630 VDD.t216 129.155
R3535 VDD.n1204 VDD.n1203 127.719
R3536 VDD.t56 VDD.t132 120.544
R3537 VDD.t203 VDD.t136 120.544
R3538 VDD.t141 VDD.t9 120.544
R3539 VDD.t31 VDD.t40 120.544
R3540 VDD.t216 VDD.t19 120.544
R3541 VDD.t213 VDD.t47 120.544
R3542 VDD.t6 VDD.t198 120.544
R3543 VDD.t3 VDD.t34 120.544
R3544 VDD.n211 VDD.t80 114.805
R3545 VDD.n3018 VDD.t230 113.897
R3546 VDD.n1214 VDD.t99 113.37
R3547 VDD.t68 VDD.n1136 113.37
R3548 VDD.n490 VDD.t89 111.934
R3549 VDD.n2710 VDD.n1387 111.177
R3550 VDD.n2746 VDD.n2744 111.177
R3551 VDD.n2570 VDD.n2568 111.177
R3552 VDD.n2591 VDD.n2589 111.177
R3553 VDD.n2617 VDD.n2616 111.177
R3554 VDD.n2637 VDD.n1437 111.177
R3555 VDD.n2484 VDD.n1521 111.177
R3556 VDD.n2520 VDD.n2518 111.177
R3557 VDD.n2344 VDD.n2342 111.177
R3558 VDD.n2365 VDD.n2363 111.177
R3559 VDD.n2391 VDD.n2390 111.177
R3560 VDD.n2411 VDD.n1571 111.177
R3561 VDD.n2258 VDD.n1655 111.177
R3562 VDD.n2294 VDD.n2292 111.177
R3563 VDD.n2118 VDD.n2116 111.177
R3564 VDD.n2139 VDD.n2137 111.177
R3565 VDD.n2165 VDD.n2164 111.177
R3566 VDD.n2185 VDD.n1705 111.177
R3567 VDD.n2032 VDD.n1789 111.177
R3568 VDD.n2068 VDD.n2066 111.177
R3569 VDD.n1913 VDD.n1911 111.177
R3570 VDD.n1939 VDD.n1938 111.177
R3571 VDD.n1959 VDD.n1839 111.177
R3572 VDD.n2797 VDD.n2795 111.177
R3573 VDD.n2816 VDD.n2814 111.177
R3574 VDD.n2835 VDD.n2833 111.177
R3575 VDD.n2854 VDD.n2852 111.177
R3576 VDD.n912 VDD 109.064
R3577 VDD VDD.n588 109.064
R3578 VDD.n2994 VDD.t232 108.719
R3579 VDD.n129 VDD.t166 107.629
R3580 VDD.n1245 VDD.t201 106.194
R3581 VDD.t209 VDD.n761 106.194
R3582 VDD.t38 VDD.n925 106.194
R3583 VDD.n109 VDD.t45 106.194
R3584 VDD.n352 VDD.t1 106.194
R3585 VDD.n362 VDD.t155 106.194
R3586 VDD.n1160 VDD.t13 104.758
R3587 VDD.t51 VDD.n1213 93.2784
R3588 VDD.t25 VDD.n1135 93.2784
R3589 VDD.n607 VDD.t29 93.2784
R3590 VDD.t122 VDD.n489 93.2784
R3591 VDD.n1116 VDD.n983 92.5005
R3592 VDD.n983 VDD.n982 92.5005
R3593 VDD.n1150 VDD.t141 92.5005
R3594 VDD.n1121 VDD.n1120 92.5005
R3595 VDD.n1122 VDD.n1121 92.5005
R3596 VDD.n1106 VDD.n979 92.5005
R3597 VDD.n1123 VDD.n979 92.5005
R3598 VDD.n1126 VDD.n1125 92.5005
R3599 VDD.n1125 VDD.n1124 92.5005
R3600 VDD.n978 VDD.n975 92.5005
R3601 VDD.n981 VDD.n978 92.5005
R3602 VDD.n972 VDD.n970 92.5005
R3603 VDD.n980 VDD.n970 92.5005
R3604 VDD.n1134 VDD.n1133 92.5005
R3605 VDD.n1135 VDD.n1134 92.5005
R3606 VDD.n971 VDD.n968 92.5005
R3607 VDD.n1136 VDD.n968 92.5005
R3608 VDD.n1139 VDD.n1138 92.5005
R3609 VDD.n1138 VDD.n1137 92.5005
R3610 VDD.n960 VDD.n956 92.5005
R3611 VDD.n969 VDD.n956 92.5005
R3612 VDD.n1145 VDD.n1144 92.5005
R3613 VDD.n1146 VDD.n1145 92.5005
R3614 VDD.n961 VDD.n955 92.5005
R3615 VDD.n1147 VDD.n955 92.5005
R3616 VDD.n1149 VDD.n951 92.5005
R3617 VDD.n1149 VDD.n1148 92.5005
R3618 VDD.n1151 VDD.n1150 92.5005
R3619 VDD.n952 VDD.n947 92.5005
R3620 VDD.n954 VDD.n952 92.5005
R3621 VDD.n1156 VDD.n943 92.5005
R3622 VDD.n953 VDD.n943 92.5005
R3623 VDD.n1159 VDD.n1158 92.5005
R3624 VDD.n1160 VDD.n1159 92.5005
R3625 VDD.n1028 VDD.n942 92.5005
R3626 VDD.n1161 VDD.n942 92.5005
R3627 VDD.n1164 VDD.n1163 92.5005
R3628 VDD.n1163 VDD.n1162 92.5005
R3629 VDD.n1166 VDD.n926 92.5005
R3630 VDD.n926 VDD.n925 92.5005
R3631 VDD.n1175 VDD.n1174 92.5005
R3632 VDD.n1176 VDD.n1175 92.5005
R3633 VDD.n932 VDD.n910 92.5005
R3634 VDD.n1177 VDD.n910 92.5005
R3635 VDD.n741 VDD.n724 92.5005
R3636 VDD.n735 VDD.n724 92.5005
R3637 VDD.n738 VDD.n737 92.5005
R3638 VDD.n737 VDD.n736 92.5005
R3639 VDD.n729 VDD.n726 92.5005
R3640 VDD.n734 VDD.n726 92.5005
R3641 VDD.n733 VDD.n732 92.5005
R3642 VDD.n1247 VDD.n1246 92.5005
R3643 VDD.n1246 VDD.n1245 92.5005
R3644 VDD.n722 VDD.n720 92.5005
R3645 VDD.n749 VDD.n722 92.5005
R3646 VDD.n747 VDD.n746 92.5005
R3647 VDD.n748 VDD.n747 92.5005
R3648 VDD.t132 VDD.n1232 92.5005
R3649 VDD.n1180 VDD.n1179 92.5005
R3650 VDD.n1179 VDD.n1178 92.5005
R3651 VDD.n917 VDD.n909 92.5005
R3652 VDD.n924 VDD.n909 92.5005
R3653 VDD.n922 VDD.n921 92.5005
R3654 VDD.n923 VDD.n922 92.5005
R3655 VDD.n1195 VDD.n797 92.5005
R3656 VDD.n912 VDD.n797 92.5005
R3657 VDD.n1196 VDD.n790 92.5005
R3658 VDD.n911 VDD.n790 92.5005
R3659 VDD.n1201 VDD.n1200 92.5005
R3660 VDD.n1202 VDD.n1201 92.5005
R3661 VDD.n788 VDD.n787 92.5005
R3662 VDD.n1203 VDD.n788 92.5005
R3663 VDD.n1206 VDD.n1205 92.5005
R3664 VDD.n1205 VDD.n1204 92.5005
R3665 VDD.n784 VDD.n783 92.5005
R3666 VDD.n789 VDD.n783 92.5005
R3667 VDD.n1211 VDD.n1210 92.5005
R3668 VDD.n1212 VDD.n1211 92.5005
R3669 VDD.n782 VDD.n781 92.5005
R3670 VDD.n1213 VDD.n782 92.5005
R3671 VDD.n1216 VDD.n1215 92.5005
R3672 VDD.n1215 VDD.n1214 92.5005
R3673 VDD.n774 VDD.n772 92.5005
R3674 VDD.n772 VDD.n771 92.5005
R3675 VDD.n1222 VDD.n1221 92.5005
R3676 VDD.n1223 VDD.n1222 92.5005
R3677 VDD.n773 VDD.n770 92.5005
R3678 VDD.n1224 VDD.n770 92.5005
R3679 VDD.n1227 VDD.n1226 92.5005
R3680 VDD.n1226 VDD.n1225 92.5005
R3681 VDD.n764 VDD.n763 92.5005
R3682 VDD.n763 VDD.n762 92.5005
R3683 VDD.n1232 VDD.n1231 92.5005
R3684 VDD.n760 VDD.n759 92.5005
R3685 VDD.n1233 VDD.n760 92.5005
R3686 VDD.n1236 VDD.n1235 92.5005
R3687 VDD.n1235 VDD.n1234 92.5005
R3688 VDD.n752 VDD.n750 92.5005
R3689 VDD.n761 VDD.n750 92.5005
R3690 VDD.n1242 VDD.n1241 92.5005
R3691 VDD.n1243 VDD.n1242 92.5005
R3692 VDD.n831 VDD.n723 92.5005
R3693 VDD.n1244 VDD.n723 92.5005
R3694 VDD.n101 VDD.n90 92.5005
R3695 VDD.n108 VDD.n90 92.5005
R3696 VDD.n106 VDD.n105 92.5005
R3697 VDD.n107 VDD.n106 92.5005
R3698 VDD.n100 VDD.n92 92.5005
R3699 VDD.n96 VDD.n92 92.5005
R3700 VDD.n98 VDD.n97 92.5005
R3701 VDD.n122 VDD.n72 92.5005
R3702 VDD.n109 VDD.n72 92.5005
R3703 VDD.n91 VDD.n84 92.5005
R3704 VDD.n110 VDD.n91 92.5005
R3705 VDD.n113 VDD.n112 92.5005
R3706 VDD.n112 VDD.n111 92.5005
R3707 VDD.n632 VDD.t216 92.5005
R3708 VDD.n301 VDD.n258 92.5005
R3709 VDD.n578 VDD.n258 92.5005
R3710 VDD.n581 VDD.n580 92.5005
R3711 VDD.n580 VDD.n579 92.5005
R3712 VDD.n256 VDD.n245 92.5005
R3713 VDD.n259 VDD.n245 92.5005
R3714 VDD.n587 VDD.n586 92.5005
R3715 VDD.n588 VDD.n587 92.5005
R3716 VDD.n249 VDD.n242 92.5005
R3717 VDD VDD.n242 92.5005
R3718 VDD.n591 VDD.n590 92.5005
R3719 VDD.n590 VDD.n589 92.5005
R3720 VDD.n241 VDD.n240 92.5005
R3721 VDD.n244 VDD.n241 92.5005
R3722 VDD.n215 VDD.n212 92.5005
R3723 VDD.n243 VDD.n212 92.5005
R3724 VDD.n604 VDD.n603 92.5005
R3725 VDD.n605 VDD.n604 92.5005
R3726 VDD.n213 VDD.n207 92.5005
R3727 VDD.n606 VDD.n207 92.5005
R3728 VDD.n609 VDD.n608 92.5005
R3729 VDD.n608 VDD.n607 92.5005
R3730 VDD.n206 VDD.n204 92.5005
R3731 VDD.n211 VDD.n206 92.5005
R3732 VDD.n209 VDD.n143 92.5005
R3733 VDD.n210 VDD.n209 92.5005
R3734 VDD.n140 VDD.n136 92.5005
R3735 VDD.n208 VDD.n136 92.5005
R3736 VDD.n627 VDD.n626 92.5005
R3737 VDD.n628 VDD.n627 92.5005
R3738 VDD.n174 VDD.n134 92.5005
R3739 VDD.n629 VDD.n134 92.5005
R3740 VDD.n631 VDD.n135 92.5005
R3741 VDD.n631 VDD.n630 92.5005
R3742 VDD.n633 VDD.n632 92.5005
R3743 VDD.n69 VDD.n65 92.5005
R3744 VDD.n133 VDD.n69 92.5005
R3745 VDD.n131 VDD.n64 92.5005
R3746 VDD.n132 VDD.n131 92.5005
R3747 VDD.n130 VDD.n71 92.5005
R3748 VDD.n130 VDD.n129 92.5005
R3749 VDD.n83 VDD.n70 92.5005
R3750 VDD.n128 VDD.n70 92.5005
R3751 VDD.n126 VDD.n125 92.5005
R3752 VDD.n127 VDD.n126 92.5005
R3753 VDD.n353 VDD.n264 92.5005
R3754 VDD.n353 VDD.n352 92.5005
R3755 VDD.n573 VDD.n260 92.5005
R3756 VDD.n351 VDD.n260 92.5005
R3757 VDD.n576 VDD.n575 92.5005
R3758 VDD.n577 VDD.n576 92.5005
R3759 VDD.t6 VDD.n373 92.5005
R3760 VDD.n460 VDD.n459 92.5005
R3761 VDD VDD.n460 92.5005
R3762 VDD.n467 VDD.n466 92.5005
R3763 VDD.n466 VDD.n465 92.5005
R3764 VDD.n454 VDD.n453 92.5005
R3765 VDD.n464 VDD.n454 92.5005
R3766 VDD.n462 VDD.n390 92.5005
R3767 VDD.n463 VDD.n462 92.5005
R3768 VDD.n480 VDD.n385 92.5005
R3769 VDD.n461 VDD.n385 92.5005
R3770 VDD.n487 VDD.n486 92.5005
R3771 VDD.n488 VDD.n487 92.5005
R3772 VDD.n429 VDD.n384 92.5005
R3773 VDD.n489 VDD.n384 92.5005
R3774 VDD.n492 VDD.n491 92.5005
R3775 VDD.n491 VDD.n490 92.5005
R3776 VDD.n495 VDD.n376 92.5005
R3777 VDD.n376 VDD.n375 92.5005
R3778 VDD.n500 VDD.n499 92.5005
R3779 VDD.n501 VDD.n500 92.5005
R3780 VDD.n411 VDD.n340 92.5005
R3781 VDD.n502 VDD.n340 92.5005
R3782 VDD.n505 VDD.n504 92.5005
R3783 VDD.n504 VDD.n503 92.5005
R3784 VDD.n339 VDD.n335 92.5005
R3785 VDD.n374 VDD.n339 92.5005
R3786 VDD.n373 VDD.n372 92.5005
R3787 VDD.n368 VDD.n341 92.5005
R3788 VDD.n360 VDD.n341 92.5005
R3789 VDD.n367 VDD.n347 92.5005
R3790 VDD.n361 VDD.n347 92.5005
R3791 VDD.n364 VDD.n363 92.5005
R3792 VDD.n363 VDD.n362 92.5005
R3793 VDD.n350 VDD.n349 92.5005
R3794 VDD.n359 VDD.n350 92.5005
R3795 VDD.n357 VDD.n356 92.5005
R3796 VDD.n358 VDD.n357 92.5005
R3797 VDD.n2992 VDD.n30 92.5005
R3798 VDD.n3020 VDD.n3019 92.5005
R3799 VDD.n3019 VDD.n3018 92.5005
R3800 VDD.n2996 VDD.n2995 92.5005
R3801 VDD.n2995 VDD.n2994 92.5005
R3802 VDD.n3015 VDD.n3014 92.5005
R3803 VDD.n3016 VDD.n3015 92.5005
R3804 VDD.n946 VDD.t84 91.4648
R3805 VDD.n946 VDD.t14 91.4648
R3806 VDD.n945 VDD.t110 91.4648
R3807 VDD.n945 VDD.t144 91.4648
R3808 VDD.n966 VDD.t69 91.4648
R3809 VDD.n965 VDD.t104 91.4648
R3810 VDD.n757 VDD.t66 91.4648
R3811 VDD.n757 VDD.t210 91.4648
R3812 VDD.n756 VDD.t94 91.4648
R3813 VDD.n756 VDD.t228 91.4648
R3814 VDD.n779 VDD.t100 91.4648
R3815 VDD.n778 VDD.t120 91.4648
R3816 VDD.n76 VDD.t75 91.4648
R3817 VDD.n76 VDD.t226 91.4648
R3818 VDD.n75 VDD.t102 91.4648
R3819 VDD.n75 VDD.t167 91.4648
R3820 VDD.n199 VDD.t108 91.4648
R3821 VDD.n198 VDD.t81 91.4648
R3822 VDD.n345 VDD.t92 91.4648
R3823 VDD.n345 VDD.t156 91.4648
R3824 VDD.n344 VDD.t63 91.4648
R3825 VDD.n344 VDD.t159 91.4648
R3826 VDD.n382 VDD.t90 91.4648
R3827 VDD.n381 VDD.t114 91.4648
R3828 VDD.n958 VDD.t24 86.7743
R3829 VDD.n957 VDD.t191 86.7743
R3830 VDD.n966 VDD.t26 86.7743
R3831 VDD.n965 VDD.t190 86.7743
R3832 VDD.n768 VDD.t196 86.7743
R3833 VDD.n767 VDD.t54 86.7743
R3834 VDD.n779 VDD.t195 86.7743
R3835 VDD.n778 VDD.t52 86.7743
R3836 VDD.n138 VDD.t28 86.7743
R3837 VDD.n137 VDD.t212 86.7743
R3838 VDD.n199 VDD.t30 86.7743
R3839 VDD.n198 VDD.t211 86.7743
R3840 VDD.n337 VDD.t125 86.7743
R3841 VDD.n336 VDD.t193 86.7743
R3842 VDD.n382 VDD.t123 86.7743
R3843 VDD.n381 VDD.t194 86.7743
R3844 VDD.t71 VDD.n748 86.1032
R3845 VDD.n1177 VDD.t77 86.1032
R3846 VDD.n1344 VDD.n1298 85.9427
R3847 VDD.n1298 VDD.n1297 85.9427
R3848 VDD.n1912 VDD.n1355 85.9427
R3849 VDD.n1940 VDD.n1355 85.9427
R3850 VDD.n1960 VDD.n1355 85.9427
R3851 VDD.n2000 VDD.n1355 85.9427
R3852 VDD.n2065 VDD.n1355 85.9427
R3853 VDD.n2090 VDD.n1355 85.9427
R3854 VDD.n2087 VDD.n1355 85.9427
R3855 VDD.n2117 VDD.n1355 85.9427
R3856 VDD.n2138 VDD.n1355 85.9427
R3857 VDD.n2166 VDD.n1355 85.9427
R3858 VDD.n2186 VDD.n1355 85.9427
R3859 VDD.n2226 VDD.n1355 85.9427
R3860 VDD.n2291 VDD.n1355 85.9427
R3861 VDD.n2316 VDD.n1355 85.9427
R3862 VDD.n2313 VDD.n1355 85.9427
R3863 VDD.n2343 VDD.n1355 85.9427
R3864 VDD.n2364 VDD.n1355 85.9427
R3865 VDD.n2392 VDD.n1355 85.9427
R3866 VDD.n2412 VDD.n1355 85.9427
R3867 VDD.n2452 VDD.n1355 85.9427
R3868 VDD.n2517 VDD.n1355 85.9427
R3869 VDD.n2542 VDD.n1355 85.9427
R3870 VDD.n2539 VDD.n1355 85.9427
R3871 VDD.n2569 VDD.n1355 85.9427
R3872 VDD.n2590 VDD.n1355 85.9427
R3873 VDD.n2618 VDD.n1355 85.9427
R3874 VDD.n2638 VDD.n1355 85.9427
R3875 VDD.n2678 VDD.n1355 85.9427
R3876 VDD.n2743 VDD.n1355 85.9427
R3877 VDD.n111 VDD.t86 84.6682
R3878 VDD.t74 VDD.n128 84.6682
R3879 VDD.n577 VDD.t96 84.6682
R3880 VDD.n1243 VDD.t65 83.2331
R3881 VDD.n1161 VDD.t83 83.2331
R3882 VDD.t62 VDD.n359 83.2331
R3883 VDD.n735 VDD.t205 78.928
R3884 VDD.n1213 VDD.t133 78.928
R3885 VDD.n1203 VDD.t134 78.928
R3886 VDD.n1178 VDD.t17 78.928
R3887 VDD.n1162 VDD.t11 78.928
R3888 VDD.n1135 VDD.t140 78.928
R3889 VDD.n607 VDD.t217 78.928
R3890 VDD.n578 VDD.t153 78.928
R3891 VDD.n489 VDD.t5 78.928
R3892 VDD.n2994 VDD 77.6572
R3893 VDD.n1244 VDD.t55 77.4929
R3894 VDD.n1123 VDD.t138 77.4929
R3895 VDD.t164 VDD.n108 77.4929
R3896 VDD.t12 VDD.n127 77.4929
R3897 VDD.n630 VDD.t27 77.4929
R3898 VDD.t147 VDD.n358 77.4929
R3899 VDD.t218 VDD.n244 76.0579
R3900 VDD.t124 VDD.n374 76.0579
R3901 VDD.t7 VDD.n464 76.0579
R3902 VDD.t207 VDD.n734 74.6229
R3903 VDD.t53 VDD.n762 74.6229
R3904 VDD.n1148 VDD.t23 74.6229
R3905 VDD.t157 VDD.n259 74.6229
R3906 VDD.n96 VDD.t168 73.1878
R3907 VDD.n1014 VDD.n1013 73.1034
R3908 VDD.n683 VDD.n50 73.1034
R3909 VDD.t15 VDD.n923 71.7528
R3910 VDD.n2927 VDD.t174 70.3649
R3911 VDD.n605 VDD.t127 70.3177
R3912 VDD.t21 VDD.n789 68.8827
R3913 VDD.t43 VDD.n912 68.8827
R3914 VDD.t10 VDD.n980 68.8827
R3915 VDD.n606 VDD.t20 68.8827
R3916 VDD.n588 VDD.t49 68.8827
R3917 VDD.n488 VDD.t199 68.8827
R3918 VDD.n2892 VDD.t143 68.0287
R3919 VDD.n1892 VDD.n1890 67.5405
R3920 VDD.n2769 VDD.n2768 67.5405
R3921 VDD.n1212 VDD.t57 67.4476
R3922 VDD VDD.t175 67.4476
R3923 VDD.t150 VDD.n981 67.4476
R3924 VDD.t179 VDD 67.4476
R3925 VDD.t130 VDD.n461 67.4476
R3926 VDD.t177 VDD 67.4476
R3927 VDD.n2657 VDD.n1426 67.3307
R3928 VDD.n2431 VDD.n1560 67.3307
R3929 VDD.n2205 VDD.n1694 67.3307
R3930 VDD.n1979 VDD.n1828 67.3307
R3931 VDD.n2873 VDD.n2872 67.3307
R3932 VDD.n1999 VDD.n1998 67.3307
R3933 VDD.n2036 VDD.n2035 67.3307
R3934 VDD.n2086 VDD.n2085 67.3307
R3935 VDD.n2225 VDD.n2224 67.3307
R3936 VDD.n2262 VDD.n2261 67.3307
R3937 VDD.n2312 VDD.n2311 67.3307
R3938 VDD.n2451 VDD.n2450 67.3307
R3939 VDD.n2488 VDD.n2487 67.3307
R3940 VDD.n2538 VDD.n2537 67.3307
R3941 VDD.n2677 VDD.n2676 67.3307
R3942 VDD.n2714 VDD.n2713 67.3307
R3943 VDD.n981 VDD.t10 66.0126
R3944 VDD.n461 VDD.t199 66.0126
R3945 VDD.n789 VDD.t57 64.5775
R3946 VDD.n1202 VDD.t175 64.5775
R3947 VDD.n923 VDD.t43 64.5775
R3948 VDD.n1122 VDD.t183 64.5775
R3949 VDD.n982 VDD.t183 64.5775
R3950 VDD.n589 VDD.t179 64.5775
R3951 VDD.n1204 VDD.t21 63.1425
R3952 VDD.n1124 VDD.t150 63.1425
R3953 VDD.t148 VDD.n96 63.1425
R3954 VDD.t20 VDD.n605 63.1425
R3955 VDD.n463 VDD.t130 63.1425
R3956 VDD.n465 VDD.t177 63.1425
R3957 VDD.n742 VDD.t72 63.1021
R3958 VDD.n743 VDD.t106 63.1021
R3959 VDD.n927 VDD.t112 63.1021
R3960 VDD.n928 VDD.t78 63.1021
R3961 VDD.n262 VDD.t118 63.1021
R3962 VDD.n263 VDD.t97 63.1021
R3963 VDD.n114 VDD.t116 63.1021
R3964 VDD.n115 VDD.t87 63.1021
R3965 VDD.n734 VDD.t35 61.7074
R3966 VDD.n243 VDD.t127 61.7074
R3967 VDD.n259 VDD.t49 61.7074
R3968 VDD.n736 VDD.t207 58.8374
R3969 VDD.n107 VDD.t168 58.8374
R3970 VDD.n728 VDD.t208 58.4849
R3971 VDD.n727 VDD.t229 58.4849
R3972 VDD.n914 VDD.t16 58.4849
R3973 VDD.n913 VDD.t146 58.4849
R3974 VDD.n94 VDD.t225 58.4849
R3975 VDD.n93 VDD.t169 58.4849
R3976 VDD.n252 VDD.t158 58.4849
R3977 VDD.n251 VDD.t160 58.4849
R3978 VDD.n1225 VDD.t53 57.4023
R3979 VDD.n924 VDD.t15 57.4023
R3980 VDD.t23 VDD.n1147 57.4023
R3981 VDD.t27 VDD.n629 57.4023
R3982 VDD.n579 VDD.t157 57.4023
R3983 VDD.n503 VDD.t124 57.4023
R3984 VDD.n465 VDD.t7 57.4023
R3985 VDD.t134 VDD.n1202 55.9673
R3986 VDD.t138 VDD.n1122 55.9673
R3987 VDD.n589 VDD.t218 55.9673
R3988 VDD.n2967 VDD.t236 55.4067
R3989 VDD.t55 VDD.n1243 54.5322
R3990 VDD.t11 VDD.n1161 54.5322
R3991 VDD.n111 VDD.t164 54.5322
R3992 VDD.t153 VDD.n577 54.5322
R3993 VDD.n359 VDD.t147 54.5322
R3994 VDD.n748 VDD.t205 53.0972
R3995 VDD.t133 VDD.n1212 53.0972
R3996 VDD.t17 VDD.n1177 53.0972
R3997 VDD.n128 VDD.t12 53.0972
R3998 VDD.n980 VDD.t140 51.6621
R3999 VDD.t217 VDD.n606 51.6621
R4000 VDD.t5 VDD.n488 51.6621
R4001 VDD.n846 VDD 50.8144
R4002 VDD.n1050 VDD 50.8144
R4003 VDD.n647 VDD 50.8144
R4004 VDD.n539 VDD 50.8144
R4005 VDD.t83 VDD.n1160 50.2271
R4006 VDD.n761 VDD.t65 48.792
R4007 VDD.n362 VDD.t62 48.792
R4008 VDD.n129 VDD.t74 47.357
R4009 VDD.n2904 VDD.t237 47.1434
R4010 VDD.n2904 VDD.t234 47.1434
R4011 VDD.n749 VDD.t71 45.9219
R4012 VDD.t77 VDD.n1176 45.9219
R4013 VDD.t86 VDD.n110 45.9219
R4014 VDD.n351 VDD.t96 44.4869
R4015 VDD.n35 VDD.n34 41.7728
R4016 VDD.n986 VDD.t220 41.5552
R4017 VDD.n986 VDD.t186 41.5552
R4018 VDD.n985 VDD.t139 41.5552
R4019 VDD.n985 VDD.t184 41.5552
R4020 VDD.n793 VDD.t135 41.5552
R4021 VDD.n793 VDD.t176 41.5552
R4022 VDD.n792 VDD.t200 41.5552
R4023 VDD.n792 VDD.t185 41.5552
R4024 VDD.n247 VDD.t238 41.5552
R4025 VDD.n247 VDD.t182 41.5552
R4026 VDD.n246 VDD.t219 41.5552
R4027 VDD.n246 VDD.t180 41.5552
R4028 VDD.n449 VDD.t8 41.5552
R4029 VDD.n449 VDD.t181 41.5552
R4030 VDD.n448 VDD.t162 41.5552
R4031 VDD.n448 VDD.t178 41.5552
R4032 VDD.n490 VDD.t122 40.1818
R4033 VDD.n3015 VDD.n2 39.0005
R4034 VDD.n1214 VDD.t51 38.7467
R4035 VDD.n1136 VDD.t25 38.7467
R4036 VDD.n958 VDD.t60 38.6969
R4037 VDD.n957 VDD.t41 38.6969
R4038 VDD.n768 VDD.t204 38.6969
R4039 VDD.n767 VDD.t223 38.6969
R4040 VDD.n138 VDD.t48 38.6969
R4041 VDD.n137 VDD.t171 38.6969
R4042 VDD.n337 VDD.t33 38.6969
R4043 VDD.n336 VDD.t4 38.6969
R4044 VDD.t29 VDD.n211 37.3117
R4045 VDD.n2967 VDD.t189 34.0906
R4046 VDD.n2089 VDD.n2088 33.746
R4047 VDD.n2315 VDD.n2314 33.746
R4048 VDD.n2541 VDD.n2540 33.746
R4049 VDD.n3017 VDD.n3016 33.6517
R4050 VDD.n1826 VDD.n1819 32.9702
R4051 VDD.n1692 VDD.n1685 32.9702
R4052 VDD.n1558 VDD.n1551 32.9702
R4053 VDD.n1424 VDD.n1417 32.9702
R4054 VDD.n728 VDD.t152 31.831
R4055 VDD.n727 VDD.t36 31.831
R4056 VDD.n914 VDD.t44 31.831
R4057 VDD.n913 VDD.t58 31.831
R4058 VDD.n94 VDD.t149 31.831
R4059 VDD.n93 VDD.t163 31.831
R4060 VDD.n252 VDD.t192 31.831
R4061 VDD.n251 VDD.t50 31.831
R4062 VDD.t37 VDD.n2992 30.5388
R4063 VDD.n2953 VDD.n2893 29.4128
R4064 VDD.n2676 VDD.n2675 28.2358
R4065 VDD.n2714 VDD.n2712 28.2358
R4066 VDD.n2768 VDD.n1356 28.2358
R4067 VDD.n2658 VDD.n2657 28.2358
R4068 VDD.n2450 VDD.n2449 28.2358
R4069 VDD.n2488 VDD.n2486 28.2358
R4070 VDD.n2537 VDD.n1491 28.2358
R4071 VDD.n2432 VDD.n2431 28.2358
R4072 VDD.n2224 VDD.n2223 28.2358
R4073 VDD.n2262 VDD.n2260 28.2358
R4074 VDD.n2311 VDD.n1625 28.2358
R4075 VDD.n2206 VDD.n2205 28.2358
R4076 VDD.n1998 VDD.n1997 28.2358
R4077 VDD.n2036 VDD.n2034 28.2358
R4078 VDD.n2085 VDD.n1759 28.2358
R4079 VDD.n1892 VDD.n1891 28.2358
R4080 VDD.n1980 VDD.n1979 28.2358
R4081 VDD.n2814 VDD.n1333 28.2358
R4082 VDD.n2833 VDD.n1322 28.2358
R4083 VDD.n2852 VDD.n1311 28.2358
R4084 VDD.n2872 VDD.n1299 28.2358
R4085 VDD.n742 VDD.t206 28.0332
R4086 VDD.n743 VDD.t227 28.0332
R4087 VDD.n927 VDD.t18 28.0332
R4088 VDD.n928 VDD.t145 28.0332
R4089 VDD.n262 VDD.t154 28.0332
R4090 VDD.n263 VDD.t161 28.0332
R4091 VDD.n114 VDD.t165 28.0332
R4092 VDD.n115 VDD.t224 28.0332
R4093 VDD.n2999 VDD.n2998 27.3454
R4094 VDD.t201 VDD.n1244 25.8313
R4095 VDD.n1234 VDD.t209 25.8313
R4096 VDD.n953 VDD.t13 25.8313
R4097 VDD.n127 VDD.t45 25.8313
R4098 VDD.n132 VDD.t166 25.8313
R4099 VDD.n358 VDD.t1 25.8313
R4100 VDD.t155 VDD.n361 25.8313
R4101 VDD.n1162 VDD.t38 24.3963
R4102 VDD VDD.n911 22.9612
R4103 VDD.n3013 VDD.n1 22.8875
R4104 VDD.n2956 VDD.n2954 20.7428
R4105 VDD.n2951 VDD.n2895 20.7428
R4106 VDD.n2952 VDD.n2894 20.7428
R4107 VDD.n2950 VDD.n2949 20.7428
R4108 VDD.n2924 VDD.n29 20.7428
R4109 VDD.n1079 VDD.n1078 19.7005
R4110 VDD.n819 VDD.n818 19.7005
R4111 VDD.n161 VDD.n160 19.7005
R4112 VDD.n520 VDD.n519 19.7005
R4113 VDD.t99 VDD.n771 18.6561
R4114 VDD.n1137 VDD.t68 18.6561
R4115 VDD.t80 VDD.n210 18.6561
R4116 VDD.t89 VDD.n375 18.6561
R4117 VDD.n2952 VDD.t126 17.4304
R4118 VDD.n2989 VDD.n36 17.0672
R4119 VDD VDD.t215 15.5577
R4120 VDD.n3022 VDD.n3021 15.4666
R4121 VDD.n2951 VDD.t121 15.4137
R4122 VDD.n28 VDD 15.1421
R4123 VDD.n2974 VDD.n2965 14.0991
R4124 VDD.n1078 VDD 13.6005
R4125 VDD.n818 VDD 13.6005
R4126 VDD.n160 VDD 13.6005
R4127 VDD.n519 VDD 13.6005
R4128 VDD.n2893 VDD.n2892 13.3673
R4129 VDD.n2679 VDD.n2678 13.1177
R4130 VDD.n2743 VDD.n2742 13.1177
R4131 VDD.n2569 VDD.n1463 13.1177
R4132 VDD.n2590 VDD.n1448 13.1177
R4133 VDD.n2619 VDD.n2618 13.1177
R4134 VDD.n2639 VDD.n2638 13.1177
R4135 VDD.n2453 VDD.n2452 13.1177
R4136 VDD.n2517 VDD.n2516 13.1177
R4137 VDD.n2543 VDD.n2542 13.1177
R4138 VDD.n2343 VDD.n1597 13.1177
R4139 VDD.n2364 VDD.n1582 13.1177
R4140 VDD.n2393 VDD.n2392 13.1177
R4141 VDD.n2413 VDD.n2412 13.1177
R4142 VDD.n2227 VDD.n2226 13.1177
R4143 VDD.n2291 VDD.n2290 13.1177
R4144 VDD.n2317 VDD.n2316 13.1177
R4145 VDD.n2117 VDD.n1731 13.1177
R4146 VDD.n2138 VDD.n1716 13.1177
R4147 VDD.n2167 VDD.n2166 13.1177
R4148 VDD.n2187 VDD.n2186 13.1177
R4149 VDD.n2001 VDD.n2000 13.1177
R4150 VDD.n2065 VDD.n2064 13.1177
R4151 VDD.n2091 VDD.n2090 13.1177
R4152 VDD.n1912 VDD.n1850 13.1177
R4153 VDD.n1941 VDD.n1940 13.1177
R4154 VDD.n1961 VDD.n1960 13.1177
R4155 VDD.n2795 VDD.n1344 13.1177
R4156 VDD.n1297 VDD.n1296 13.1177
R4157 VDD.n2776 VDD.n1344 13.1177
R4158 VDD.n2000 VDD.n1789 13.1177
R4159 VDD.n2066 VDD.n2065 13.1177
R4160 VDD.n2226 VDD.n1655 13.1177
R4161 VDD.n2292 VDD.n2291 13.1177
R4162 VDD.n2452 VDD.n1521 13.1177
R4163 VDD.n2518 VDD.n2517 13.1177
R4164 VDD.n2678 VDD.n1387 13.1177
R4165 VDD.n2744 VDD.n2743 13.1177
R4166 VDD.n2638 VDD.n2637 13.1177
R4167 VDD.n2618 VDD.n2617 13.1177
R4168 VDD.n2591 VDD.n2590 13.1177
R4169 VDD.n2570 VDD.n2569 13.1177
R4170 VDD.n2539 VDD.n1474 13.1177
R4171 VDD.n2412 VDD.n2411 13.1177
R4172 VDD.n2392 VDD.n2391 13.1177
R4173 VDD.n2365 VDD.n2364 13.1177
R4174 VDD.n2344 VDD.n2343 13.1177
R4175 VDD.n2313 VDD.n1608 13.1177
R4176 VDD.n2186 VDD.n2185 13.1177
R4177 VDD.n2166 VDD.n2165 13.1177
R4178 VDD.n2139 VDD.n2138 13.1177
R4179 VDD.n2118 VDD.n2117 13.1177
R4180 VDD.n2087 VDD.n1742 13.1177
R4181 VDD.n1960 VDD.n1959 13.1177
R4182 VDD.n1940 VDD.n1939 13.1177
R4183 VDD.n1913 VDD.n1912 13.1177
R4184 VDD.t9 VDD.n954 12.9159
R4185 VDD.n2969 VDD.n2968 12.4295
R4186 VDD.n3015 VDD.n4 12.0005
R4187 VDD.n3020 VDD.n1 11.9758
R4188 VDD.t42 VDD.n29 11.8125
R4189 VDD.n2770 VDD.n2769 11.5452
R4190 VDD.n1890 VDD.n1889 11.5452
R4191 VDD.n1233 VDD.t56 11.4809
R4192 VDD.n360 VDD.t198 11.4809
R4193 VDD.n2999 VDD.n2996 11.2229
R4194 VDD.n2950 VDD.t42 10.8041
R4195 VDD.n3016 VDD.n3 10.3547
R4196 VDD.t19 VDD.n133 10.0458
R4197 VDD.n858 VDD.n855 9.49444
R4198 VDD.n1044 VDD.n1041 9.49444
R4199 VDD.n659 VDD.n656 9.49444
R4200 VDD.n552 VDD.n548 9.49444
R4201 VDD.n2674 VDD.n2673 9.38471
R4202 VDD.n2660 VDD.n2659 9.38471
R4203 VDD.n2448 VDD.n2447 9.38471
R4204 VDD.n2434 VDD.n2433 9.38471
R4205 VDD.n2222 VDD.n2221 9.38471
R4206 VDD.n2208 VDD.n2207 9.38471
R4207 VDD.n1996 VDD.n1995 9.38471
R4208 VDD.n1982 VDD.n1981 9.38471
R4209 VDD.n86 VDD 9.37843
R4210 VDD.n715 VDD 9.37838
R4211 VDD.n1826 VDD.n1825 9.3005
R4212 VDD.n2083 VDD.n2082 9.3005
R4213 VDD.n2039 VDD.n2038 9.3005
R4214 VDD.n2006 VDD.n2005 9.3005
R4215 VDD.n1820 VDD.n1819 9.3005
R4216 VDD.n1791 VDD.n1790 9.3005
R4217 VDD.n1776 VDD.n1775 9.3005
R4218 VDD.n1692 VDD.n1691 9.3005
R4219 VDD.n2309 VDD.n2308 9.3005
R4220 VDD.n2265 VDD.n2264 9.3005
R4221 VDD.n2232 VDD.n2231 9.3005
R4222 VDD.n1686 VDD.n1685 9.3005
R4223 VDD.n1657 VDD.n1656 9.3005
R4224 VDD.n1642 VDD.n1641 9.3005
R4225 VDD.n1558 VDD.n1557 9.3005
R4226 VDD.n2535 VDD.n2534 9.3005
R4227 VDD.n2491 VDD.n2490 9.3005
R4228 VDD.n2458 VDD.n2457 9.3005
R4229 VDD.n1552 VDD.n1551 9.3005
R4230 VDD.n1523 VDD.n1522 9.3005
R4231 VDD.n1508 VDD.n1507 9.3005
R4232 VDD.n1424 VDD.n1423 9.3005
R4233 VDD.n2766 VDD.n2765 9.3005
R4234 VDD.n2717 VDD.n2716 9.3005
R4235 VDD.n2684 VDD.n2683 9.3005
R4236 VDD.n1418 VDD.n1417 9.3005
R4237 VDD.n1389 VDD.n1388 9.3005
R4238 VDD.n1374 VDD.n1373 9.3005
R4239 VDD.n2655 VDD.n2654 9.3005
R4240 VDD.n2635 VDD.n2634 9.3005
R4241 VDD.n1454 VDD.n1453 9.3005
R4242 VDD.n2594 VDD.n2593 9.3005
R4243 VDD.n2573 VDD.n2572 9.3005
R4244 VDD.n2429 VDD.n2428 9.3005
R4245 VDD.n2409 VDD.n2408 9.3005
R4246 VDD.n1588 VDD.n1587 9.3005
R4247 VDD.n2368 VDD.n2367 9.3005
R4248 VDD.n2347 VDD.n2346 9.3005
R4249 VDD.n2203 VDD.n2202 9.3005
R4250 VDD.n2183 VDD.n2182 9.3005
R4251 VDD.n1722 VDD.n1721 9.3005
R4252 VDD.n2142 VDD.n2141 9.3005
R4253 VDD.n2121 VDD.n2120 9.3005
R4254 VDD.n1977 VDD.n1976 9.3005
R4255 VDD.n1957 VDD.n1956 9.3005
R4256 VDD.n1856 VDD.n1855 9.3005
R4257 VDD.n1895 VDD.n1894 9.3005
R4258 VDD.n1916 VDD.n1915 9.3005
R4259 VDD.n2975 VDD.n2974 9.3005
R4260 VDD.n1076 VDD.n1075 9.3005
R4261 VDD.n816 VDD.n815 9.3005
R4262 VDD.n830 VDD.n719 9.3005
R4263 VDD.n977 VDD.n976 9.3005
R4264 VDD.n921 VDD.n920 9.3005
R4265 VDD.n931 VDD.n908 9.3005
R4266 VDD.n1018 VDD.n1017 9.3005
R4267 VDD.n1017 VDD.n1016 9.3005
R4268 VDD.n1259 VDD.n1258 9.3005
R4269 VDD.n851 VDD.n850 9.3005
R4270 VDD.n848 VDD.n845 9.3005
R4271 VDD.n848 VDD.n847 9.3005
R4272 VDD.n860 VDD.n843 9.3005
R4273 VDD.n1055 VDD.n1054 9.3005
R4274 VDD.n1052 VDD.n1049 9.3005
R4275 VDD.n1052 VDD.n1051 9.3005
R4276 VDD.n1047 VDD.n1046 9.3005
R4277 VDD.n272 VDD.n268 9.3005
R4278 VDD.n275 VDD.n274 9.3005
R4279 VDD.n158 VDD.n157 9.3005
R4280 VDD.n379 VDD.n377 9.3005
R4281 VDD.n497 VDD.n378 9.3005
R4282 VDD.n175 VDD.n172 9.3005
R4283 VDD.n77 VDD.n74 9.3005
R4284 VDD.n121 VDD.n120 9.3005
R4285 VDD.n239 VDD.n238 9.3005
R4286 VDD.n223 VDD.n205 9.3005
R4287 VDD.n201 VDD.n200 9.3005
R4288 VDD.n370 VDD.n342 9.3005
R4289 VDD.n483 VDD.n387 9.3005
R4290 VDD.n452 VDD.n451 9.3005
R4291 VDD.n456 VDD.n455 9.3005
R4292 VDD.n517 VDD.n516 9.3005
R4293 VDD.n686 VDD.n682 9.3005
R4294 VDD.n686 VDD.n685 9.3005
R4295 VDD.n652 VDD.n651 9.3005
R4296 VDD.n649 VDD.n646 9.3005
R4297 VDD.n649 VDD.n648 9.3005
R4298 VDD.n662 VDD.n661 9.3005
R4299 VDD.n316 VDD.n315 9.3005
R4300 VDD.n313 VDD.n312 9.3005
R4301 VDD.n541 VDD.n538 9.3005
R4302 VDD.n541 VDD.n540 9.3005
R4303 VDD.n544 VDD.n543 9.3005
R4304 VDD.n554 VDD.n549 9.3005
R4305 VDD.n2793 VDD.n2792 9.3005
R4306 VDD.n2812 VDD.n2811 9.3005
R4307 VDD.n2831 VDD.n2830 9.3005
R4308 VDD.n2850 VDD.n2849 9.3005
R4309 VDD.n2870 VDD.n2869 9.3005
R4310 VDD.n2799 VDD.n2798 9.3005
R4311 VDD.n2798 VDD.n2797 9.3005
R4312 VDD.n2818 VDD.n2817 9.3005
R4313 VDD.n2817 VDD.n2816 9.3005
R4314 VDD.n2837 VDD.n2836 9.3005
R4315 VDD.n2836 VDD.n2835 9.3005
R4316 VDD.n2856 VDD.n2855 9.3005
R4317 VDD.n2855 VDD.n2854 9.3005
R4318 VDD.n2876 VDD.n2875 9.3005
R4319 VDD.n2875 VDD.n2874 9.3005
R4320 VDD.n2778 VDD.n2777 9.3005
R4321 VDD.n2777 VDD.n1298 9.3005
R4322 VDD.n2094 VDD.n2093 9.3005
R4323 VDD.n2093 VDD.n2092 9.3005
R4324 VDD.n2062 VDD.n2061 9.3005
R4325 VDD.n2062 VDD.n1771 9.3005
R4326 VDD.n2003 VDD.n1793 9.3005
R4327 VDD.n2003 VDD.n2002 9.3005
R4328 VDD.n1995 VDD.n1994 9.3005
R4329 VDD.n2031 VDD.n1787 9.3005
R4330 VDD.n2032 VDD.n2031 9.3005
R4331 VDD.n2070 VDD.n2069 9.3005
R4332 VDD.n2069 VDD.n2068 9.3005
R4333 VDD.n2320 VDD.n2319 9.3005
R4334 VDD.n2319 VDD.n2318 9.3005
R4335 VDD.n2288 VDD.n2287 9.3005
R4336 VDD.n2288 VDD.n1637 9.3005
R4337 VDD.n2229 VDD.n1659 9.3005
R4338 VDD.n2229 VDD.n2228 9.3005
R4339 VDD.n2221 VDD.n2220 9.3005
R4340 VDD.n2257 VDD.n1653 9.3005
R4341 VDD.n2258 VDD.n2257 9.3005
R4342 VDD.n2296 VDD.n2295 9.3005
R4343 VDD.n2295 VDD.n2294 9.3005
R4344 VDD.n2546 VDD.n2545 9.3005
R4345 VDD.n2545 VDD.n2544 9.3005
R4346 VDD.n2514 VDD.n2513 9.3005
R4347 VDD.n2514 VDD.n1503 9.3005
R4348 VDD.n2455 VDD.n1525 9.3005
R4349 VDD.n2455 VDD.n2454 9.3005
R4350 VDD.n2447 VDD.n2446 9.3005
R4351 VDD.n2483 VDD.n1519 9.3005
R4352 VDD.n2484 VDD.n2483 9.3005
R4353 VDD.n2522 VDD.n2521 9.3005
R4354 VDD.n2521 VDD.n2520 9.3005
R4355 VDD.n2740 VDD.n2739 9.3005
R4356 VDD.n2740 VDD.n1369 9.3005
R4357 VDD.n2681 VDD.n1391 9.3005
R4358 VDD.n2681 VDD.n2680 9.3005
R4359 VDD.n2673 VDD.n2672 9.3005
R4360 VDD.n2709 VDD.n1385 9.3005
R4361 VDD.n2710 VDD.n2709 9.3005
R4362 VDD.n2748 VDD.n2747 9.3005
R4363 VDD.n2747 VDD.n2746 9.3005
R4364 VDD.n2771 VDD.n2770 9.3005
R4365 VDD.n2642 VDD.n2641 9.3005
R4366 VDD.n2641 VDD.n2640 9.3005
R4367 VDD.n2622 VDD.n2621 9.3005
R4368 VDD.n2621 VDD.n1437 9.3005
R4369 VDD.n1437 VDD.n1355 9.3005
R4370 VDD.n2615 VDD.n2614 9.3005
R4371 VDD.n2616 VDD.n2615 9.3005
R4372 VDD.n2616 VDD.n1355 9.3005
R4373 VDD.n2588 VDD.n2587 9.3005
R4374 VDD.n2589 VDD.n2588 9.3005
R4375 VDD.n2589 VDD.n1355 9.3005
R4376 VDD.n2661 VDD.n2660 9.3005
R4377 VDD.n2567 VDD.n2566 9.3005
R4378 VDD.n2568 VDD.n2567 9.3005
R4379 VDD.n2568 VDD.n1355 9.3005
R4380 VDD.n2416 VDD.n2415 9.3005
R4381 VDD.n2415 VDD.n2414 9.3005
R4382 VDD.n2396 VDD.n2395 9.3005
R4383 VDD.n2395 VDD.n1571 9.3005
R4384 VDD.n1571 VDD.n1355 9.3005
R4385 VDD.n2389 VDD.n2388 9.3005
R4386 VDD.n2390 VDD.n2389 9.3005
R4387 VDD.n2390 VDD.n1355 9.3005
R4388 VDD.n2362 VDD.n2361 9.3005
R4389 VDD.n2363 VDD.n2362 9.3005
R4390 VDD.n2363 VDD.n1355 9.3005
R4391 VDD.n2435 VDD.n2434 9.3005
R4392 VDD.n2341 VDD.n2340 9.3005
R4393 VDD.n2342 VDD.n2341 9.3005
R4394 VDD.n2342 VDD.n1355 9.3005
R4395 VDD.n2190 VDD.n2189 9.3005
R4396 VDD.n2189 VDD.n2188 9.3005
R4397 VDD.n2170 VDD.n2169 9.3005
R4398 VDD.n2169 VDD.n1705 9.3005
R4399 VDD.n1705 VDD.n1355 9.3005
R4400 VDD.n2163 VDD.n2162 9.3005
R4401 VDD.n2164 VDD.n2163 9.3005
R4402 VDD.n2164 VDD.n1355 9.3005
R4403 VDD.n2136 VDD.n2135 9.3005
R4404 VDD.n2137 VDD.n2136 9.3005
R4405 VDD.n2137 VDD.n1355 9.3005
R4406 VDD.n2209 VDD.n2208 9.3005
R4407 VDD.n2115 VDD.n2114 9.3005
R4408 VDD.n2116 VDD.n2115 9.3005
R4409 VDD.n2116 VDD.n1355 9.3005
R4410 VDD.n1964 VDD.n1963 9.3005
R4411 VDD.n1963 VDD.n1962 9.3005
R4412 VDD.n1944 VDD.n1943 9.3005
R4413 VDD.n1943 VDD.n1839 9.3005
R4414 VDD.n1839 VDD.n1355 9.3005
R4415 VDD.n1937 VDD.n1936 9.3005
R4416 VDD.n1938 VDD.n1937 9.3005
R4417 VDD.n1938 VDD.n1355 9.3005
R4418 VDD.n1983 VDD.n1982 9.3005
R4419 VDD.n1889 VDD.n1888 9.3005
R4420 VDD.n1910 VDD.n1909 9.3005
R4421 VDD.n1911 VDD.n1910 9.3005
R4422 VDD.n2972 VDD.n2971 9.3005
R4423 VDD.n2998 VDD.n2997 9.3005
R4424 VDD.n3012 VDD.n3011 9.3005
R4425 VDD.n3012 VDD.n4 9.3005
R4426 VDD.n4 VDD.n3 9.3005
R4427 VDD.n936 VDD 9.2607
R4428 VDD.n936 VDD.n935 9.14483
R4429 VDD.t121 VDD.n2950 9.07556
R4430 VDD.n1028 VDD.n941 9.05896
R4431 VDD.n1028 VDD.n944 9.05896
R4432 VDD.n1152 VDD.n1151 9.05896
R4433 VDD.n1151 VDD.n951 9.05896
R4434 VDD.n961 VDD.n951 9.05896
R4435 VDD.n1140 VDD.n1139 9.05896
R4436 VDD.n1133 VDD.n971 9.05896
R4437 VDD.n1130 VDD.n1129 9.05896
R4438 VDD.n738 VDD.n725 9.05896
R4439 VDD.n741 VDD.n738 9.05896
R4440 VDD.n1241 VDD.n752 9.05896
R4441 VDD.n1236 VDD.n759 9.05896
R4442 VDD.n1231 VDD.n759 9.05896
R4443 VDD.n1231 VDD.n764 9.05896
R4444 VDD.n1227 VDD.n764 9.05896
R4445 VDD.n1221 VDD.n773 9.05896
R4446 VDD.n1221 VDD.n774 9.05896
R4447 VDD.n1216 VDD.n781 9.05896
R4448 VDD.n1210 VDD.n781 9.05896
R4449 VDD.n1210 VDD.n784 9.05896
R4450 VDD.n1206 VDD.n784 9.05896
R4451 VDD.n1196 VDD.n1195 9.05896
R4452 VDD.n105 VDD.n100 9.05896
R4453 VDD.n105 VDD.n102 9.05896
R4454 VDD.n586 VDD.n250 9.05896
R4455 VDD.n301 VDD.n257 9.05896
R4456 VDD.n356 VDD.n349 9.05896
R4457 VDD.n364 VDD.n349 9.05896
R4458 VDD.n368 VDD.n367 9.05896
R4459 VDD.n506 VDD.n505 9.05896
R4460 VDD.n429 VDD.n383 9.05896
R4461 VDD.n1156 VDD.n947 8.9605
R4462 VDD.n1144 VDD.n960 8.9605
R4463 VDD.n1133 VDD.n972 8.9605
R4464 VDD.n1126 VDD.n975 8.9605
R4465 VDD.n1200 VDD.n791 8.9605
R4466 VDD.n1181 VDD.n907 8.9605
R4467 VDD.n125 VDD.n83 8.9605
R4468 VDD.n82 VDD.n71 8.9605
R4469 VDD.n633 VDD.n65 8.9605
R4470 VDD.n625 VDD.n140 8.9605
R4471 VDD.n603 VDD.n214 8.9605
R4472 VDD.n602 VDD.n215 8.9605
R4473 VDD.n582 VDD.n581 8.9605
R4474 VDD.n1894 VDD.n1893 8.92171
R4475 VDD.n1915 VDD.n1914 8.92171
R4476 VDD.n1855 VDD.n1849 8.92171
R4477 VDD.n1958 VDD.n1957 8.92171
R4478 VDD.n1978 VDD.n1977 8.92171
R4479 VDD.n2005 VDD.n1803 8.92171
R4480 VDD.n1804 VDD.n1790 8.92171
R4481 VDD.n2038 VDD.n2037 8.92171
R4482 VDD.n1775 VDD.n1770 8.92171
R4483 VDD.n2084 VDD.n2083 8.92171
R4484 VDD.n2120 VDD.n2119 8.92171
R4485 VDD.n2141 VDD.n2140 8.92171
R4486 VDD.n1721 VDD.n1715 8.92171
R4487 VDD.n2184 VDD.n2183 8.92171
R4488 VDD.n2204 VDD.n2203 8.92171
R4489 VDD.n2231 VDD.n1669 8.92171
R4490 VDD.n1670 VDD.n1656 8.92171
R4491 VDD.n2264 VDD.n2263 8.92171
R4492 VDD.n1641 VDD.n1636 8.92171
R4493 VDD.n2310 VDD.n2309 8.92171
R4494 VDD.n2346 VDD.n2345 8.92171
R4495 VDD.n2367 VDD.n2366 8.92171
R4496 VDD.n1587 VDD.n1581 8.92171
R4497 VDD.n2410 VDD.n2409 8.92171
R4498 VDD.n2430 VDD.n2429 8.92171
R4499 VDD.n2457 VDD.n1535 8.92171
R4500 VDD.n1536 VDD.n1522 8.92171
R4501 VDD.n2490 VDD.n2489 8.92171
R4502 VDD.n1507 VDD.n1502 8.92171
R4503 VDD.n2536 VDD.n2535 8.92171
R4504 VDD.n2572 VDD.n2571 8.92171
R4505 VDD.n2593 VDD.n2592 8.92171
R4506 VDD.n1453 VDD.n1447 8.92171
R4507 VDD.n2636 VDD.n2635 8.92171
R4508 VDD.n2656 VDD.n2655 8.92171
R4509 VDD.n2683 VDD.n1401 8.92171
R4510 VDD.n1402 VDD.n1388 8.92171
R4511 VDD.n2716 VDD.n2715 8.92171
R4512 VDD.n1373 VDD.n1368 8.92171
R4513 VDD.n2767 VDD.n2766 8.92171
R4514 VDD.n2794 VDD.n2793 8.92171
R4515 VDD.n2813 VDD.n2812 8.92171
R4516 VDD.n2832 VDD.n2831 8.92171
R4517 VDD.n2851 VDD.n2850 8.92171
R4518 VDD.n2871 VDD.n2870 8.92171
R4519 VDD.n1196 VDD.n794 8.86204
R4520 VDD.n921 VDD.n917 8.86204
R4521 VDD.n2796 VDD.n1298 8.77616
R4522 VDD.n2815 VDD.n1298 8.77616
R4523 VDD.n2834 VDD.n1298 8.77616
R4524 VDD.n2853 VDD.n1298 8.77616
R4525 VDD.n1996 VDD.n1355 8.77616
R4526 VDD.n2033 VDD.n1355 8.77616
R4527 VDD.n2067 VDD.n1355 8.77616
R4528 VDD.n2222 VDD.n1355 8.77616
R4529 VDD.n2259 VDD.n1355 8.77616
R4530 VDD.n2293 VDD.n1355 8.77616
R4531 VDD.n2448 VDD.n1355 8.77616
R4532 VDD.n2485 VDD.n1355 8.77616
R4533 VDD.n2519 VDD.n1355 8.77616
R4534 VDD.n2674 VDD.n1355 8.77616
R4535 VDD.n2711 VDD.n1355 8.77616
R4536 VDD.n2745 VDD.n1355 8.77616
R4537 VDD.n2659 VDD.n1355 8.77616
R4538 VDD.n2433 VDD.n1355 8.77616
R4539 VDD.n2207 VDD.n1355 8.77616
R4540 VDD.n1981 VDD.n1355 8.77616
R4541 VDD.n1865 VDD.n1355 8.77616
R4542 VDD.n860 VDD.n855 8.76429
R4543 VDD.n1046 VDD.n1041 8.76429
R4544 VDD.n661 VDD.n656 8.76429
R4545 VDD.n554 VDD.n548 8.76429
R4546 VDD.n1120 VDD.n984 8.76358
R4547 VDD.n1206 VDD.n787 8.76358
R4548 VDD.n592 VDD.n591 8.76358
R4549 VDD.n249 VDD.n248 8.76358
R4550 VDD.n622 VDD.n621 8.66512
R4551 VDD.n628 VDD.t47 8.61077
R4552 VDD.n1116 VDD.n987 8.56665
R4553 VDD.n732 VDD.n730 8.56665
R4554 VDD.n1241 VDD.n751 8.56665
R4555 VDD.n98 VDD.n95 8.56665
R4556 VDD.n637 VDD.n636 8.56665
R4557 VDD.n586 VDD.n253 8.56665
R4558 VDD.n480 VDD.n479 8.56665
R4559 VDD.n368 VDD.n342 8.46819
R4560 VDD.n481 VDD.n387 8.46819
R4561 VDD.n2972 VDD.n30 8.45089
R4562 VDD.n2990 VDD.n2989 8.45089
R4563 VDD.n610 VDD.n204 8.36973
R4564 VDD.n1257 VDD.n1256 8.30364
R4565 VDD.n272 VDD.n271 8.30364
R4566 VDD.n633 VDD.n68 8.27127
R4567 VDD.n499 VDD.n378 8.27127
R4568 VDD.n2991 VDD.n2990 8.25289
R4569 VDD.n175 VDD.n174 8.17281
R4570 VDD.n468 VDD.n447 8.17281
R4571 VDD.n459 VDD.n455 8.17281
R4572 VDD.n811 VDD.n810 8.00414
R4573 VDD.n512 VDD.n511 8.00414
R4574 VDD.n1071 VDD.n1070 8.00389
R4575 VDD.n153 VDD.n152 8.00389
R4576 VDD.n499 VDD.n377 7.97588
R4577 VDD.n429 VDD.n386 7.97588
R4578 VDD.n86 VDD.n85 7.96107
R4579 VDD.n715 VDD.n714 7.96106
R4580 VDD.n213 VDD.n205 7.87742
R4581 VDD.n343 VDD.n335 7.87742
R4582 VDD.n1015 VDD 7.7918
R4583 VDD.n453 VDD.n452 7.6805
R4584 VDD.t173 VDD.t235 7.63507
R4585 VDD.n1157 VDD.n1156 7.58204
R4586 VDD.n1126 VDD.n977 7.58204
R4587 VDD.n1236 VDD.n758 7.58204
R4588 VDD.n239 VDD.n237 7.58204
R4589 VDD.n367 VDD.n346 7.58204
R4590 VDD.n746 VDD.n741 7.57296
R4591 VDD.n301 VDD.n261 7.57296
R4592 VDD.n684 VDD 7.51354
R4593 VDD.n1195 VDD.n796 7.48358
R4594 VDD.n101 VDD.n89 7.4745
R4595 VDD.n847 VDD.n846 7.34676
R4596 VDD.n1051 VDD.n1050 7.34676
R4597 VDD.n648 VDD.n647 7.34676
R4598 VDD.n540 VDD.n539 7.34676
R4599 VDD.n313 VDD.n284 7.21714
R4600 VDD.n1224 VDD.t203 7.17573
R4601 VDD.n1146 VDD.t40 7.17573
R4602 VDD VDD.t173 7.05888
R4603 VDD.n1076 VDD.n1074 6.95412
R4604 VDD.n816 VDD.n814 6.95412
R4605 VDD.n158 VDD.n156 6.95412
R4606 VDD.n517 VDD.n515 6.95412
R4607 VDD.n34 VDD.n33 6.85649
R4608 VDD.n1258 VDD 6.67876
R4609 VDD.n274 VDD 6.67876
R4610 VDD.n1016 VDD.n1014 6.54941
R4611 VDD.n685 VDD.n683 6.54941
R4612 VDD.n78 VDD.n77 6.4005
R4613 VDD.n315 VDD 6.4005
R4614 VDD.n1139 VDD.n967 6.10512
R4615 VDD.n780 VDD.n774 6.10512
R4616 VDD.n932 VDD.n908 5.99758
R4617 VDD.n502 VDD.t3 5.74068
R4618 VDD.n2873 VDD.n1298 5.63319
R4619 VDD.n1828 VDD.n1355 5.63319
R4620 VDD.n2086 VDD.n1355 5.63319
R4621 VDD.n2035 VDD.n1355 5.63319
R4622 VDD.n1999 VDD.n1355 5.63319
R4623 VDD.n1694 VDD.n1355 5.63319
R4624 VDD.n2312 VDD.n1355 5.63319
R4625 VDD.n2261 VDD.n1355 5.63319
R4626 VDD.n2225 VDD.n1355 5.63319
R4627 VDD.n1560 VDD.n1355 5.63319
R4628 VDD.n2538 VDD.n1355 5.63319
R4629 VDD.n2487 VDD.n1355 5.63319
R4630 VDD.n2451 VDD.n1355 5.63319
R4631 VDD.n1426 VDD.n1355 5.63319
R4632 VDD.n2713 VDD.n1355 5.63319
R4633 VDD.n2677 VDD.n1355 5.63319
R4634 VDD.t187 VDD.n32 5.23391
R4635 VDD.n494 VDD.n493 5.21896
R4636 VDD.n1890 VDD.n1355 5.1329
R4637 VDD.n2769 VDD.n1355 5.1329
R4638 VDD.n850 VDD 5.0092
R4639 VDD.n1054 VDD 5.0092
R4640 VDD.n651 VDD 5.0092
R4641 VDD.n543 VDD 5.0092
R4642 VDD.n961 VDD.n959 4.82512
R4643 VDD.n1227 VDD.n769 4.82512
R4644 VDD.n174 VDD.n139 4.82512
R4645 VDD.n202 VDD.n201 4.82512
R4646 VDD.n505 VDD.n338 4.82512
R4647 VDD.n2993 VDD.t37 4.7541
R4648 VDD.n33 VDD 4.7541
R4649 VDD.n1258 VDD.n1257 4.73093
R4650 VDD.n2977 VDD.n2965 4.6505
R4651 VDD.n2973 VDD.n2966 4.6505
R4652 VDD.n37 VDD.n36 4.6505
R4653 VDD.n849 VDD.n844 4.6505
R4654 VDD.n1053 VDD.n1048 4.6505
R4655 VDD.n650 VDD.n645 4.6505
R4656 VDD.n542 VDD.n537 4.6505
R4657 VDD.n7 VDD.n1 4.6505
R4658 VDD.n3000 VDD.n2999 4.6505
R4659 VDD.n811 VDD 4.55532
R4660 VDD.n512 VDD 4.55532
R4661 VDD.n1071 VDD 4.55472
R4662 VDD.n153 VDD 4.55472
R4663 VDD.n682 VDD.n681 4.54858
R4664 VDD.n1019 VDD.n1018 4.54617
R4665 VDD.n688 VDD.n687 4.54479
R4666 VDD.n1012 VDD.n1009 4.54309
R4667 VDD.n1888 VDD.n1876 4.54027
R4668 VDD.n2772 VDD.n2771 4.54027
R4669 VDD.n549 VDD.n534 4.53929
R4670 VDD.n2906 VDD.n2905 4.52882
R4671 VDD.n1259 VDD.n1255 4.51252
R4672 VDD.n276 VDD.n275 4.51252
R4673 VDD.n317 VDD.n316 4.51012
R4674 VDD.n1874 VDD.n1873 4.5005
R4675 VDD.n1875 VDD.n1874 4.5005
R4676 VDD.n1897 VDD.n1896 4.5005
R4677 VDD.n1918 VDD.n1917 4.5005
R4678 VDD.n1824 VDD.n1823 4.5005
R4679 VDD.n1832 VDD.n1816 4.5005
R4680 VDD.n2104 VDD.n1744 4.5005
R4681 VDD.n1756 VDD.n1749 4.5005
R4682 VDD.n2081 VDD.n2080 4.5005
R4683 VDD.n1755 VDD.n1753 4.5005
R4684 VDD.n1757 VDD.n1755 4.5005
R4685 VDD.n2060 VDD.n2059 4.5005
R4686 VDD.n2042 VDD.n2041 4.5005
R4687 VDD.n2040 VDD.n1773 4.5005
R4688 VDD.n1773 VDD.n1772 4.5005
R4689 VDD.n2025 VDD.n2024 4.5005
R4690 VDD.n2008 VDD.n2007 4.5005
R4691 VDD.n1802 VDD.n1800 4.5005
R4692 VDD.n2004 VDD.n1802 4.5005
R4693 VDD.n1801 VDD.n1799 4.5005
R4694 VDD.n1822 VDD.n1821 4.5005
R4695 VDD.n1809 VDD.n1808 4.5005
R4696 VDD.n1808 VDD.n1807 4.5005
R4697 VDD.n2044 VDD.n2043 4.5005
R4698 VDD.n2027 VDD.n2026 4.5005
R4699 VDD.n2029 VDD.n2028 4.5005
R4700 VDD.n2030 VDD.n2029 4.5005
R4701 VDD.n1762 VDD.n1761 4.5005
R4702 VDD.n1779 VDD.n1777 4.5005
R4703 VDD.n1768 VDD.n1766 4.5005
R4704 VDD.n1769 VDD.n1768 4.5005
R4705 VDD.n1690 VDD.n1689 4.5005
R4706 VDD.n1698 VDD.n1682 4.5005
R4707 VDD.n2330 VDD.n1610 4.5005
R4708 VDD.n1622 VDD.n1615 4.5005
R4709 VDD.n2307 VDD.n2306 4.5005
R4710 VDD.n1621 VDD.n1619 4.5005
R4711 VDD.n1623 VDD.n1621 4.5005
R4712 VDD.n2286 VDD.n2285 4.5005
R4713 VDD.n2268 VDD.n2267 4.5005
R4714 VDD.n2266 VDD.n1639 4.5005
R4715 VDD.n1639 VDD.n1638 4.5005
R4716 VDD.n2251 VDD.n2250 4.5005
R4717 VDD.n2234 VDD.n2233 4.5005
R4718 VDD.n1668 VDD.n1666 4.5005
R4719 VDD.n2230 VDD.n1668 4.5005
R4720 VDD.n1667 VDD.n1665 4.5005
R4721 VDD.n1688 VDD.n1687 4.5005
R4722 VDD.n1675 VDD.n1674 4.5005
R4723 VDD.n1674 VDD.n1673 4.5005
R4724 VDD.n2270 VDD.n2269 4.5005
R4725 VDD.n2253 VDD.n2252 4.5005
R4726 VDD.n2255 VDD.n2254 4.5005
R4727 VDD.n2256 VDD.n2255 4.5005
R4728 VDD.n1628 VDD.n1627 4.5005
R4729 VDD.n1645 VDD.n1643 4.5005
R4730 VDD.n1634 VDD.n1632 4.5005
R4731 VDD.n1635 VDD.n1634 4.5005
R4732 VDD.n1556 VDD.n1555 4.5005
R4733 VDD.n1564 VDD.n1548 4.5005
R4734 VDD.n2556 VDD.n1476 4.5005
R4735 VDD.n1488 VDD.n1481 4.5005
R4736 VDD.n2533 VDD.n2532 4.5005
R4737 VDD.n1487 VDD.n1485 4.5005
R4738 VDD.n1489 VDD.n1487 4.5005
R4739 VDD.n2512 VDD.n2511 4.5005
R4740 VDD.n2494 VDD.n2493 4.5005
R4741 VDD.n2492 VDD.n1505 4.5005
R4742 VDD.n1505 VDD.n1504 4.5005
R4743 VDD.n2477 VDD.n2476 4.5005
R4744 VDD.n2460 VDD.n2459 4.5005
R4745 VDD.n1534 VDD.n1532 4.5005
R4746 VDD.n2456 VDD.n1534 4.5005
R4747 VDD.n1533 VDD.n1531 4.5005
R4748 VDD.n1554 VDD.n1553 4.5005
R4749 VDD.n1541 VDD.n1540 4.5005
R4750 VDD.n1540 VDD.n1539 4.5005
R4751 VDD.n2496 VDD.n2495 4.5005
R4752 VDD.n2479 VDD.n2478 4.5005
R4753 VDD.n2481 VDD.n2480 4.5005
R4754 VDD.n2482 VDD.n2481 4.5005
R4755 VDD.n1494 VDD.n1493 4.5005
R4756 VDD.n1511 VDD.n1509 4.5005
R4757 VDD.n1500 VDD.n1498 4.5005
R4758 VDD.n1501 VDD.n1500 4.5005
R4759 VDD.n1422 VDD.n1421 4.5005
R4760 VDD.n1430 VDD.n1414 4.5005
R4761 VDD.n2764 VDD.n2763 4.5005
R4762 VDD.n2738 VDD.n2737 4.5005
R4763 VDD.n2720 VDD.n2719 4.5005
R4764 VDD.n2718 VDD.n1371 4.5005
R4765 VDD.n1371 VDD.n1370 4.5005
R4766 VDD.n2703 VDD.n2702 4.5005
R4767 VDD.n2686 VDD.n2685 4.5005
R4768 VDD.n1400 VDD.n1398 4.5005
R4769 VDD.n2682 VDD.n1400 4.5005
R4770 VDD.n1399 VDD.n1397 4.5005
R4771 VDD.n1420 VDD.n1419 4.5005
R4772 VDD.n1407 VDD.n1406 4.5005
R4773 VDD.n1406 VDD.n1405 4.5005
R4774 VDD.n2722 VDD.n2721 4.5005
R4775 VDD.n2705 VDD.n2704 4.5005
R4776 VDD.n2707 VDD.n2706 4.5005
R4777 VDD.n2708 VDD.n2707 4.5005
R4778 VDD.n1359 VDD.n1358 4.5005
R4779 VDD.n1377 VDD.n1375 4.5005
R4780 VDD.n1366 VDD.n1364 4.5005
R4781 VDD.n1367 VDD.n1366 4.5005
R4782 VDD.n2762 VDD.n1352 4.5005
R4783 VDD.n1354 VDD.n1352 4.5005
R4784 VDD.n2576 VDD.n1465 4.5005
R4785 VDD.n2653 VDD.n2652 4.5005
R4786 VDD.n1441 VDD.n1435 4.5005
R4787 VDD.n1429 VDD.n1428 4.5005
R4788 VDD.n1428 VDD.n1427 4.5005
R4789 VDD.n2633 VDD.n2632 4.5005
R4790 VDD.n1455 VDD.n1446 4.5005
R4791 VDD.n1440 VDD.n1439 4.5005
R4792 VDD.n1439 VDD.n1438 4.5005
R4793 VDD.n2611 VDD.n2610 4.5005
R4794 VDD.n2598 VDD.n1451 4.5005
R4795 VDD.n2613 VDD.n2612 4.5005
R4796 VDD.n2613 VDD.n1450 4.5005
R4797 VDD.n1461 VDD.n1460 4.5005
R4798 VDD.n1462 VDD.n1461 4.5005
R4799 VDD.n2596 VDD.n2595 4.5005
R4800 VDD.n1415 VDD.n1413 4.5005
R4801 VDD.n1425 VDD.n1415 4.5005
R4802 VDD.n1472 VDD.n1471 4.5005
R4803 VDD.n1473 VDD.n1472 4.5005
R4804 VDD.n2575 VDD.n2574 4.5005
R4805 VDD.n2350 VDD.n1599 4.5005
R4806 VDD.n2427 VDD.n2426 4.5005
R4807 VDD.n1575 VDD.n1569 4.5005
R4808 VDD.n1563 VDD.n1562 4.5005
R4809 VDD.n1562 VDD.n1561 4.5005
R4810 VDD.n2407 VDD.n2406 4.5005
R4811 VDD.n1589 VDD.n1580 4.5005
R4812 VDD.n1574 VDD.n1573 4.5005
R4813 VDD.n1573 VDD.n1572 4.5005
R4814 VDD.n2385 VDD.n2384 4.5005
R4815 VDD.n2372 VDD.n1585 4.5005
R4816 VDD.n2387 VDD.n2386 4.5005
R4817 VDD.n2387 VDD.n1584 4.5005
R4818 VDD.n1595 VDD.n1594 4.5005
R4819 VDD.n1596 VDD.n1595 4.5005
R4820 VDD.n2370 VDD.n2369 4.5005
R4821 VDD.n1549 VDD.n1547 4.5005
R4822 VDD.n1559 VDD.n1549 4.5005
R4823 VDD.n1606 VDD.n1605 4.5005
R4824 VDD.n1607 VDD.n1606 4.5005
R4825 VDD.n2349 VDD.n2348 4.5005
R4826 VDD.n2124 VDD.n1733 4.5005
R4827 VDD.n2201 VDD.n2200 4.5005
R4828 VDD.n1709 VDD.n1703 4.5005
R4829 VDD.n1697 VDD.n1696 4.5005
R4830 VDD.n1696 VDD.n1695 4.5005
R4831 VDD.n2181 VDD.n2180 4.5005
R4832 VDD.n1723 VDD.n1714 4.5005
R4833 VDD.n1708 VDD.n1707 4.5005
R4834 VDD.n1707 VDD.n1706 4.5005
R4835 VDD.n2159 VDD.n2158 4.5005
R4836 VDD.n2146 VDD.n1719 4.5005
R4837 VDD.n2161 VDD.n2160 4.5005
R4838 VDD.n2161 VDD.n1718 4.5005
R4839 VDD.n1729 VDD.n1728 4.5005
R4840 VDD.n1730 VDD.n1729 4.5005
R4841 VDD.n2144 VDD.n2143 4.5005
R4842 VDD.n1683 VDD.n1681 4.5005
R4843 VDD.n1693 VDD.n1683 4.5005
R4844 VDD.n1740 VDD.n1739 4.5005
R4845 VDD.n1741 VDD.n1740 4.5005
R4846 VDD.n2123 VDD.n2122 4.5005
R4847 VDD.n1920 VDD.n1853 4.5005
R4848 VDD.n1975 VDD.n1974 4.5005
R4849 VDD.n1843 VDD.n1837 4.5005
R4850 VDD.n1831 VDD.n1830 4.5005
R4851 VDD.n1830 VDD.n1829 4.5005
R4852 VDD.n1955 VDD.n1954 4.5005
R4853 VDD.n1857 VDD.n1848 4.5005
R4854 VDD.n1842 VDD.n1841 4.5005
R4855 VDD.n1841 VDD.n1840 4.5005
R4856 VDD.n1935 VDD.n1934 4.5005
R4857 VDD.n1935 VDD.n1852 4.5005
R4858 VDD.n1933 VDD.n1932 4.5005
R4859 VDD.n1817 VDD.n1815 4.5005
R4860 VDD.n1827 VDD.n1817 4.5005
R4861 VDD.n1863 VDD.n1862 4.5005
R4862 VDD.n1864 VDD.n1863 4.5005
R4863 VDD.n1898 VDD.n1867 4.5005
R4864 VDD.n836 VDD.n753 4.5005
R4865 VDD.n833 VDD.n829 4.5005
R4866 VDD.n833 VDD.n751 4.5005
R4867 VDD.n1115 VDD.n1114 4.5005
R4868 VDD.n1185 VDD.n1184 4.5005
R4869 VDD.n1182 VDD.n906 4.5005
R4870 VDD.n1182 VDD.n1181 4.5005
R4871 VDD.n1172 VDD.n1171 4.5005
R4872 VDD.n1172 VDD.n930 4.5005
R4873 VDD.n1169 VDD.n1168 4.5005
R4874 VDD.n1110 VDD.n1109 4.5005
R4875 VDD.n1109 VDD.n984 4.5005
R4876 VDD.n1193 VDD.n1192 4.5005
R4877 VDD.n918 VDD.n800 4.5005
R4878 VDD.n918 VDD.n796 4.5005
R4879 VDD.n1011 VDD.n1010 4.5005
R4880 VDD.n854 VDD.n842 4.5005
R4881 VDD.n863 VDD.n862 4.5005
R4882 VDD.n1038 VDD.n1037 4.5005
R4883 VDD.n1059 VDD.n1058 4.5005
R4884 VDD.n273 VDD.n270 4.5005
R4885 VDD.n418 VDD.n380 4.5005
R4886 VDD.n494 VDD.n380 4.5005
R4887 VDD.n427 VDD.n426 4.5005
R4888 VDD.n408 VDD.n407 4.5005
R4889 VDD.n415 VDD.n414 4.5005
R4890 VDD.n414 VDD.n413 4.5005
R4891 VDD.n166 VDD.n67 4.5005
R4892 VDD.n639 VDD.n638 4.5005
R4893 VDD.n638 VDD.n637 4.5005
R4894 VDD.n118 VDD.n117 4.5005
R4895 VDD.n291 VDD.n290 4.5005
R4896 VDD.n594 VDD.n593 4.5005
R4897 VDD.n593 VDD.n592 4.5005
R4898 VDD.n600 VDD.n599 4.5005
R4899 VDD.n601 VDD.n217 4.5005
R4900 VDD.n226 VDD.n225 4.5005
R4901 VDD.n611 VDD.n197 4.5005
R4902 VDD.n611 VDD.n610 4.5005
R4903 VDD.n614 VDD.n613 4.5005
R4904 VDD.n620 VDD.n619 4.5005
R4905 VDD.n621 VDD.n620 4.5005
R4906 VDD.n188 VDD.n142 4.5005
R4907 VDD.n167 VDD.n66 4.5005
R4908 VDD.n431 VDD.n397 4.5005
R4909 VDD.n434 VDD.n388 4.5005
R4910 VDD.n388 VDD.n386 4.5005
R4911 VDD.n437 VDD.n389 4.5005
R4912 VDD.n478 VDD.n477 4.5005
R4913 VDD.n479 VDD.n478 4.5005
R4914 VDD.n472 VDD.n471 4.5005
R4915 VDD.n469 VDD.n446 4.5005
R4916 VDD.n469 VDD.n468 4.5005
R4917 VDD.n178 VDD.n166 4.5005
R4918 VDD.n178 VDD.n68 4.5005
R4919 VDD.n508 VDD.n333 4.5005
R4920 VDD.n343 VDD.n333 4.5005
R4921 VDD.n509 VDD.n508 4.5005
R4922 VDD.n664 VDD.n663 4.5005
R4923 VDD.n655 VDD.n643 4.5005
R4924 VDD.n283 VDD.n282 4.5005
R4925 VDD.n557 VDD.n556 4.5005
R4926 VDD.n547 VDD.n536 4.5005
R4927 VDD.n2868 VDD.n2867 4.5005
R4928 VDD.n2879 VDD.n1283 4.5005
R4929 VDD.n1347 VDD.n1346 4.5005
R4930 VDD.n1336 VDD.n1335 4.5005
R4931 VDD.n2791 VDD.n2790 4.5005
R4932 VDD.n1325 VDD.n1324 4.5005
R4933 VDD.n2810 VDD.n2809 4.5005
R4934 VDD.n1314 VDD.n1313 4.5005
R4935 VDD.n2829 VDD.n2828 4.5005
R4936 VDD.n1302 VDD.n1301 4.5005
R4937 VDD.n2848 VDD.n2847 4.5005
R4938 VDD.n1293 VDD.n1291 4.5005
R4939 VDD.n1294 VDD.n1293 4.5005
R4940 VDD.n1342 VDD.n1340 4.5005
R4941 VDD.n1343 VDD.n1342 4.5005
R4942 VDD.n1331 VDD.n1329 4.5005
R4943 VDD.n1332 VDD.n1331 4.5005
R4944 VDD.n1320 VDD.n1318 4.5005
R4945 VDD.n1321 VDD.n1320 4.5005
R4946 VDD.n1309 VDD.n1307 4.5005
R4947 VDD.n1310 VDD.n1309 4.5005
R4948 VDD.n27 VDD.n26 4.5005
R4949 VDD.n9 VDD.n6 4.5005
R4950 VDD.n10 VDD.n8 4.5005
R4951 VDD.t126 VDD.n2951 4.466
R4952 VDD.n1077 VDD.n1073 4.46483
R4953 VDD.n817 VDD.n813 4.46483
R4954 VDD.n159 VDD.n155 4.46483
R4955 VDD.n518 VDD.n514 4.46483
R4956 VDD.n274 VDD.n273 4.45267
R4957 VDD.n315 VDD.n314 4.45267
R4958 VDD.t136 VDD.n1223 4.30564
R4959 VDD.t34 VDD.n501 4.30564
R4960 VDD.n1144 VDD.n959 4.23435
R4961 VDD.n773 VDD.n769 4.23435
R4962 VDD.n1247 VDD.n720 4.17639
R4963 VDD.n572 VDD.n264 4.17639
R4964 VDD.n684 VDD.n50 4.17441
R4965 VDD.n125 VDD.n73 4.15683
R4966 VDD.n356 VDD.n354 4.15683
R4967 VDD.n626 VDD.n139 4.13588
R4968 VDD.n1165 VDD.n1164 4.05837
R4969 VDD.n1298 VDD 4.03386
R4970 VDD.t235 VDD.t187 4.03386
R4971 VDD.n87 VDD.n86 3.97836
R4972 VDD.n1174 VDD.n929 3.94944
R4973 VDD.n744 VDD.n720 3.94944
R4974 VDD.n122 VDD.n121 3.94944
R4975 VDD.n574 VDD.n573 3.90405
R4976 VDD.n1015 VDD.n1013 3.89615
R4977 VDD.n413 VDD.n338 3.64358
R4978 VDD.n2928 VDD.n2909 3.62088
R4979 VDD.n1017 VDD.n1012 3.56525
R4980 VDD.n1083 VDD.n1082 3.52848
R4981 VDD.n2927 VDD.n2926 3.47503
R4982 VDD.n1169 VDD.n939 3.47069
R4983 VDD.n1104 VDD.n1103 3.46971
R4984 VDD.n1098 VDD.n1096 3.46971
R4985 VDD.n886 VDD.n776 3.46971
R4986 VDD.n869 VDD.n754 3.46971
R4987 VDD.n1273 VDD.n1272 3.46971
R4988 VDD.n892 VDD.n891 3.46971
R4989 VDD.n1064 VDD.n949 3.46971
R4990 VDD.n1268 VDD.n1267 3.46971
R4991 VDD.n1032 VDD.n1031 3.46971
R4992 VDD.n898 VDD.n897 3.46971
R4993 VDD.n1091 VDD.n963 3.46971
R4994 VDD.n694 VDD.n693 3.46971
R4995 VDD.n699 VDD.n698 3.46971
R4996 VDD.n532 VDD.n531 3.46971
R4997 VDD.n565 VDD.n564 3.46971
R4998 VDD.n304 VDD.n300 3.46971
R4999 VDD.n295 VDD.n254 3.46971
R5000 VDD.n185 VDD.n184 3.46971
R5001 VDD.n677 VDD.n676 3.46971
R5002 VDD.n672 VDD.n671 3.46971
R5003 VDD.n3002 VDD.n25 3.46788
R5004 VDD.n1192 VDD.n799 3.46752
R5005 VDD.n20 VDD.n19 3.46651
R5006 VDD.n1084 VDD.n1069 3.46532
R5007 VDD.n2979 VDD.n2978 3.46323
R5008 VDD.n2985 VDD.n38 3.46323
R5009 VDD.n2907 VDD.n2901 3.46321
R5010 VDD.n311 VDD.n309 3.46041
R5011 VDD.n841 VDD.n839 3.45822
R5012 VDD.n1039 VDD.n1035 3.45822
R5013 VDD.n642 VDD.n57 3.45754
R5014 VDD.n422 VDD.n397 3.45655
R5015 VDD.n2917 VDD.n2916 3.45407
R5016 VDD.n2958 VDD.n2957 3.45407
R5017 VDD.n2933 VDD.n2932 3.45407
R5018 VDD.n2948 VDD.n2897 3.45407
R5019 VDD.n2942 VDD.n2940 3.45407
R5020 VDD.n473 VDD.n472 3.45217
R5021 VDD.n2914 VDD.n2913 3.45149
R5022 VDD.n2955 VDD.n1279 3.45149
R5023 VDD.n426 VDD.n425 3.44997
R5024 VDD.n1111 VDD.n1110 3.44778
R5025 VDD.n615 VDD.n614 3.44778
R5026 VDD.n407 VDD.n406 3.44778
R5027 VDD.n1114 VDD.n1113 3.44676
R5028 VDD.n1005 VDD.n906 3.44559
R5029 VDD.n595 VDD.n594 3.44559
R5030 VDD.n1263 VDD.n1262 3.445
R5031 VDD.n438 VDD.n437 3.44339
R5032 VDD.n446 VDD.n441 3.44237
R5033 VDD.n829 VDD.n828 3.4412
R5034 VDD.n837 VDD.n836 3.4412
R5035 VDD.n189 VDD.n188 3.4412
R5036 VDD.n619 VDD.n618 3.4412
R5037 VDD.n640 VDD.n639 3.4412
R5038 VDD.n168 VDD.n167 3.4412
R5039 VDD.n2936 VDD.n2935 3.44028
R5040 VDD.n2898 VDD.n2896 3.44028
R5041 VDD.n2941 VDD.n2911 3.44028
R5042 VDD.n477 VDD.n476 3.43901
R5043 VDD.n1186 VDD.n1185 3.43682
R5044 VDD.n292 VDD.n291 3.43682
R5045 VDD.n220 VDD.n197 3.43462
R5046 VDD.n416 VDD.n415 3.43462
R5047 VDD.n419 VDD.n418 3.43243
R5048 VDD.n668 VDD.n57 3.43119
R5049 VDD.n561 VDD.n324 3.43092
R5050 VDD.n536 VDD.n325 3.43069
R5051 VDD.n1035 VDD.n1034 3.43066
R5052 VDD.n867 VDD.n839 3.43015
R5053 VDD.n643 VDD.n58 3.42988
R5054 VDD.n2782 VDD.n2775 3.42985
R5055 VDD.n227 VDD.n226 3.42804
R5056 VDD.n1060 VDD.n1059 3.42768
R5057 VDD.n2964 VDD.n2963 3.4267
R5058 VDD.n842 VDD.n840 3.42631
R5059 VDD.n1020 VDD.n1019 3.42585
R5060 VDD.n435 VDD.n434 3.42585
R5061 VDD.n534 VDD.n324 3.42585
R5062 VDD.n13 VDD.n10 3.4257
R5063 VDD.n568 VDD.n567 3.42489
R5064 VDD.n1089 VDD.n1088 3.42488
R5065 VDD.n2984 VDD.n39 3.42476
R5066 VDD.n2930 VDD.n2929 3.42476
R5067 VDD.n2889 VDD.n1285 3.42443
R5068 VDD.n1252 VDD.n1251 3.42429
R5069 VDD.n1102 VDD.n1101 3.42429
R5070 VDD.n1100 VDD.n1099 3.42429
R5071 VDD.n889 VDD.n888 3.42429
R5072 VDD.n872 VDD.n871 3.42429
R5073 VDD.n1271 VDD.n1270 3.42429
R5074 VDD.n894 VDD.n893 3.42429
R5075 VDD.n1067 VDD.n1066 3.42429
R5076 VDD.n1266 VDD.n1265 3.42429
R5077 VDD.n1027 VDD.n1026 3.42429
R5078 VDD.n896 VDD.n895 3.42429
R5079 VDD.n1094 VDD.n1093 3.42429
R5080 VDD.n692 VDD.n691 3.42429
R5081 VDD.n697 VDD.n696 3.42429
R5082 VDD.n530 VDD.n529 3.42429
R5083 VDD.n563 VDD.n562 3.42429
R5084 VDD.n306 VDD.n305 3.42429
R5085 VDD.n298 VDD.n297 3.42429
R5086 VDD.n187 VDD.n186 3.42429
R5087 VDD.n675 VDD.n674 3.42429
R5088 VDD.n670 VDD.n669 3.42429
R5089 VDD.n884 VDD.n883 3.42428
R5090 VDD.n874 VDD.n873 3.42428
R5091 VDD.n1880 VDD.n1876 3.42376
R5092 VDD.n2773 VDD.n2772 3.42376
R5093 VDD.n1255 VDD.n1254 3.42366
R5094 VDD.n689 VDD.n688 3.42366
R5095 VDD.n182 VDD.n181 3.42296
R5096 VDD.n681 VDD.n680 3.42146
R5097 VDD.n171 VDD.n170 3.4199
R5098 VDD.n528 VDD.n527 3.4199
R5099 VDD.n1009 VDD.n1008 3.41927
R5100 VDD.n2903 VDD.n2900 3.41853
R5101 VDD.n599 VDD.n598 3.41708
R5102 VDD.n318 VDD.n317 3.41708
R5103 VDD.n801 VDD.n800 3.41489
R5104 VDD.n26 VDD.n11 3.41388
R5105 VDD.n2774 VDD.n2773 3.41326
R5106 VDD.n1880 VDD.n1879 3.41257
R5107 VDD.n2917 VDD.n2912 3.41218
R5108 VDD.n2958 VDD.n1278 3.41218
R5109 VDD.n2980 VDD.n2979 3.41218
R5110 VDD.n2981 VDD.n38 3.41218
R5111 VDD.n2937 VDD.n2936 3.41218
R5112 VDD.n2932 VDD.n2931 3.41218
R5113 VDD.n2922 VDD.n2898 3.41218
R5114 VDD.n2925 VDD.n2897 3.41218
R5115 VDD.n2939 VDD.n2911 3.41218
R5116 VDD.n2940 VDD.n2939 3.41218
R5117 VDD.n1105 VDD.n1104 3.41212
R5118 VDD.n1096 VDD.n1095 3.41212
R5119 VDD.n1069 VDD.n1068 3.41212
R5120 VDD.n886 VDD.n885 3.41212
R5121 VDD.n869 VDD.n868 3.41212
R5122 VDD.n716 VDD.n707 3.41212
R5123 VDD.n1274 VDD.n1273 3.41212
R5124 VDD.n891 VDD.n890 3.41212
R5125 VDD.n1064 VDD.n1063 3.41212
R5126 VDD.n1187 VDD.n1186 3.41212
R5127 VDD.n1006 VDD.n1005 3.41212
R5128 VDD.n1023 VDD.n1022 3.41212
R5129 VDD.n1025 VDD.n939 3.41212
R5130 VDD.n1112 VDD.n1111 3.41212
R5131 VDD.n1269 VDD.n1268 3.41212
R5132 VDD.n828 VDD.n712 3.41212
R5133 VDD.n838 VDD.n837 3.41212
R5134 VDD.n877 VDD.n876 3.41212
R5135 VDD.n881 VDD.n809 3.41212
R5136 VDD.n1033 VDD.n1032 3.41212
R5137 VDD.n899 VDD.n898 3.41212
R5138 VDD.n1091 VDD.n1090 3.41212
R5139 VDD.n900 VDD.n799 3.41212
R5140 VDD.n1188 VDD.n801 3.41212
R5141 VDD.n1008 VDD.n1007 3.41212
R5142 VDD.n1021 VDD.n1020 3.41212
R5143 VDD.n1264 VDD.n1263 3.41212
R5144 VDD.n1254 VDD.n1253 3.41212
R5145 VDD.n695 VDD.n694 3.41212
R5146 VDD.n700 VDD.n699 3.41212
R5147 VDD.n423 VDD.n422 3.41212
R5148 VDD.n436 VDD.n435 3.41212
R5149 VDD.n439 VDD.n438 3.41212
R5150 VDD.n476 VDD.n475 3.41212
R5151 VDD.n533 VDD.n532 3.41212
R5152 VDD.n566 VDD.n565 3.41212
R5153 VDD.n280 VDD.n267 3.41212
R5154 VDD.n300 VDD.n299 3.41212
R5155 VDD.n295 VDD.n294 3.41212
R5156 VDD.n184 VDD.n183 3.41212
R5157 VDD.n678 VDD.n677 3.41212
R5158 VDD.n190 VDD.n189 3.41212
R5159 VDD.n618 VDD.n617 3.41212
R5160 VDD.n616 VDD.n615 3.41212
R5161 VDD.n221 VDD.n220 3.41212
R5162 VDD.n228 VDD.n227 3.41212
R5163 VDD.n598 VDD.n597 3.41212
R5164 VDD.n596 VDD.n595 3.41212
R5165 VDD.n293 VDD.n292 3.41212
R5166 VDD.n474 VDD.n473 3.41212
R5167 VDD.n673 VDD.n672 3.41212
R5168 VDD.n641 VDD.n640 3.41212
R5169 VDD.n169 VDD.n168 3.41212
R5170 VDD.n406 VDD.n405 3.41212
R5171 VDD.n417 VDD.n416 3.41212
R5172 VDD.n420 VDD.n419 3.41212
R5173 VDD.n425 VDD.n424 3.41212
R5174 VDD.n404 VDD.n332 3.41212
R5175 VDD.n690 VDD.n689 3.41212
R5176 VDD.n680 VDD.n679 3.41212
R5177 VDD.n309 VDD.n308 3.41212
R5178 VDD.n319 VDD.n318 3.41212
R5179 VDD.n2902 VDD.n2899 3.41162
R5180 VDD.n1900 VDD.n1899 3.4105
R5181 VDD.n1908 VDD.n1907 3.4105
R5182 VDD.n1993 VDD.n1992 3.4105
R5183 VDD.n2012 VDD.n1794 3.4105
R5184 VDD.n2017 VDD.n1785 3.4105
R5185 VDD.n2051 VDD.n1774 3.4105
R5186 VDD.n2072 VDD.n2071 3.4105
R5187 VDD.n2096 VDD.n2095 3.4105
R5188 VDD.n2106 VDD.n2105 3.4105
R5189 VDD.n2219 VDD.n2218 3.4105
R5190 VDD.n2238 VDD.n1660 3.4105
R5191 VDD.n2243 VDD.n1651 3.4105
R5192 VDD.n2277 VDD.n1640 3.4105
R5193 VDD.n2298 VDD.n2297 3.4105
R5194 VDD.n2322 VDD.n2321 3.4105
R5195 VDD.n2332 VDD.n2331 3.4105
R5196 VDD.n2445 VDD.n2444 3.4105
R5197 VDD.n2464 VDD.n1526 3.4105
R5198 VDD.n2469 VDD.n1517 3.4105
R5199 VDD.n2503 VDD.n1506 3.4105
R5200 VDD.n2524 VDD.n2523 3.4105
R5201 VDD.n2548 VDD.n2547 3.4105
R5202 VDD.n2558 VDD.n2557 3.4105
R5203 VDD.n2671 VDD.n2670 3.4105
R5204 VDD.n2690 VDD.n1392 3.4105
R5205 VDD.n2695 VDD.n1383 3.4105
R5206 VDD.n2729 VDD.n1372 3.4105
R5207 VDD.n2750 VDD.n2749 3.4105
R5208 VDD.n2754 VDD.n1353 3.4105
R5209 VDD.n2761 VDD.n2760 3.4105
R5210 VDD.n2736 VDD.n2735 3.4105
R5211 VDD.n1384 VDD.n1380 3.4105
R5212 VDD.n1394 VDD.n1390 3.4105
R5213 VDD.n2688 VDD.n2687 3.4105
R5214 VDD.n2644 VDD.n2643 3.4105
R5215 VDD.n2631 VDD.n2630 3.4105
R5216 VDD.n2624 VDD.n2623 3.4105
R5217 VDD.n2609 VDD.n2608 3.4105
R5218 VDD.n2602 VDD.n1452 3.4105
R5219 VDD.n2597 VDD.n1458 3.4105
R5220 VDD.n2586 VDD.n2585 3.4105
R5221 VDD.n2578 VDD.n2577 3.4105
R5222 VDD.n2651 VDD.n2650 3.4105
R5223 VDD.n2663 VDD.n2662 3.4105
R5224 VDD.n2565 VDD.n2564 3.4105
R5225 VDD.n2555 VDD.n2554 3.4105
R5226 VDD.n2531 VDD.n2530 3.4105
R5227 VDD.n2510 VDD.n2509 3.4105
R5228 VDD.n1518 VDD.n1514 3.4105
R5229 VDD.n1528 VDD.n1524 3.4105
R5230 VDD.n2462 VDD.n2461 3.4105
R5231 VDD.n2418 VDD.n2417 3.4105
R5232 VDD.n2405 VDD.n2404 3.4105
R5233 VDD.n2398 VDD.n2397 3.4105
R5234 VDD.n2383 VDD.n2382 3.4105
R5235 VDD.n2376 VDD.n1586 3.4105
R5236 VDD.n2371 VDD.n1592 3.4105
R5237 VDD.n2360 VDD.n2359 3.4105
R5238 VDD.n2352 VDD.n2351 3.4105
R5239 VDD.n2425 VDD.n2424 3.4105
R5240 VDD.n2437 VDD.n2436 3.4105
R5241 VDD.n2339 VDD.n2338 3.4105
R5242 VDD.n2329 VDD.n2328 3.4105
R5243 VDD.n2305 VDD.n2304 3.4105
R5244 VDD.n2284 VDD.n2283 3.4105
R5245 VDD.n1652 VDD.n1648 3.4105
R5246 VDD.n1662 VDD.n1658 3.4105
R5247 VDD.n2236 VDD.n2235 3.4105
R5248 VDD.n2192 VDD.n2191 3.4105
R5249 VDD.n2179 VDD.n2178 3.4105
R5250 VDD.n2172 VDD.n2171 3.4105
R5251 VDD.n2157 VDD.n2156 3.4105
R5252 VDD.n2150 VDD.n1720 3.4105
R5253 VDD.n2145 VDD.n1726 3.4105
R5254 VDD.n2134 VDD.n2133 3.4105
R5255 VDD.n2126 VDD.n2125 3.4105
R5256 VDD.n2199 VDD.n2198 3.4105
R5257 VDD.n2211 VDD.n2210 3.4105
R5258 VDD.n2113 VDD.n2112 3.4105
R5259 VDD.n2103 VDD.n2102 3.4105
R5260 VDD.n2079 VDD.n2078 3.4105
R5261 VDD.n2058 VDD.n2057 3.4105
R5262 VDD.n1786 VDD.n1782 3.4105
R5263 VDD.n1796 VDD.n1792 3.4105
R5264 VDD.n2010 VDD.n2009 3.4105
R5265 VDD.n1966 VDD.n1965 3.4105
R5266 VDD.n1953 VDD.n1952 3.4105
R5267 VDD.n1946 VDD.n1945 3.4105
R5268 VDD.n1931 VDD.n1930 3.4105
R5269 VDD.n1924 VDD.n1854 3.4105
R5270 VDD.n1919 VDD.n1860 3.4105
R5271 VDD.n1973 VDD.n1972 3.4105
R5272 VDD.n1985 VDD.n1984 3.4105
R5273 VDD.n1887 VDD.n1886 3.4105
R5274 VDD.n2903 VDD.n2902 3.4105
R5275 VDD.n2908 VDD.n2907 3.4105
R5276 VDD.n1083 VDD.n997 3.4105
R5277 VDD.n717 VDD.n716 3.4105
R5278 VDD.n1022 VDD.n937 3.4105
R5279 VDD.n878 VDD.n877 3.4105
R5280 VDD.n881 VDD.n880 3.4105
R5281 VDD.n866 VDD.n865 3.4105
R5282 VDD.n1062 VDD.n1061 3.4105
R5283 VDD.n279 VDD.n278 3.4105
R5284 VDD.n569 VDD.n267 3.4105
R5285 VDD.n165 VDD.n151 3.4105
R5286 VDD.n524 VDD.n330 3.4105
R5287 VDD.n526 VDD.n332 3.4105
R5288 VDD.n560 VDD.n559 3.4105
R5289 VDD.n667 VDD.n666 3.4105
R5290 VDD.n2945 VDD.n2944 3.4105
R5291 VDD.n2960 VDD.n2959 3.4105
R5292 VDD.n2959 VDD.n1280 3.4105
R5293 VDD.n2919 VDD.n2918 3.4105
R5294 VDD.n2920 VDD.n2919 3.4105
R5295 VDD.n1882 VDD.n1881 3.4105
R5296 VDD.n1885 VDD.n1884 3.4105
R5297 VDD.n1906 VDD.n1905 3.4105
R5298 VDD.n2757 VDD.n1361 3.4105
R5299 VDD.n1350 VDD.n1349 3.4105
R5300 VDD.n2759 VDD.n2758 3.4105
R5301 VDD.n1363 VDD.n1362 3.4105
R5302 VDD.n2753 VDD.n1360 3.4105
R5303 VDD.n2734 VDD.n2733 3.4105
R5304 VDD.n2728 VDD.n1379 3.4105
R5305 VDD.n2732 VDD.n1378 3.4105
R5306 VDD.n2727 VDD.n2726 3.4105
R5307 VDD.n2696 VDD.n2694 3.4105
R5308 VDD.n2725 VDD.n2724 3.4105
R5309 VDD.n2698 VDD.n2697 3.4105
R5310 VDD.n2692 VDD.n2691 3.4105
R5311 VDD.n2700 VDD.n2699 3.4105
R5312 VDD.n2689 VDD.n1395 3.4105
R5313 VDD.n2666 VDD.n1409 3.4105
R5314 VDD.n2667 VDD.n1396 3.4105
R5315 VDD.n2584 VDD.n2583 3.4105
R5316 VDD.n1470 VDD.n1469 3.4105
R5317 VDD.n2580 VDD.n2579 3.4105
R5318 VDD.n2604 VDD.n2603 3.4105
R5319 VDD.n2582 VDD.n1468 3.4105
R5320 VDD.n2600 VDD.n1459 3.4105
R5321 VDD.n2626 VDD.n2625 3.4105
R5322 VDD.n2605 VDD.n1456 3.4105
R5323 VDD.n2607 VDD.n2606 3.4105
R5324 VDD.n2646 VDD.n2645 3.4105
R5325 VDD.n2627 VDD.n1442 3.4105
R5326 VDD.n2629 VDD.n2628 3.4105
R5327 VDD.n2665 VDD.n2664 3.4105
R5328 VDD.n2647 VDD.n1431 3.4105
R5329 VDD.n2649 VDD.n2648 3.4105
R5330 VDD.n2563 VDD.n2562 3.4105
R5331 VDD.n1480 VDD.n1479 3.4105
R5332 VDD.n2560 VDD.n2559 3.4105
R5333 VDD.n2553 VDD.n2552 3.4105
R5334 VDD.n1484 VDD.n1483 3.4105
R5335 VDD.n2551 VDD.n1482 3.4105
R5336 VDD.n2529 VDD.n2528 3.4105
R5337 VDD.n1497 VDD.n1496 3.4105
R5338 VDD.n2527 VDD.n1495 3.4105
R5339 VDD.n2508 VDD.n2507 3.4105
R5340 VDD.n2502 VDD.n1513 3.4105
R5341 VDD.n2506 VDD.n1512 3.4105
R5342 VDD.n2501 VDD.n2500 3.4105
R5343 VDD.n2470 VDD.n2468 3.4105
R5344 VDD.n2499 VDD.n2498 3.4105
R5345 VDD.n2472 VDD.n2471 3.4105
R5346 VDD.n2466 VDD.n2465 3.4105
R5347 VDD.n2474 VDD.n2473 3.4105
R5348 VDD.n2463 VDD.n1529 3.4105
R5349 VDD.n2440 VDD.n1543 3.4105
R5350 VDD.n2441 VDD.n1530 3.4105
R5351 VDD.n2358 VDD.n2357 3.4105
R5352 VDD.n1604 VDD.n1603 3.4105
R5353 VDD.n2354 VDD.n2353 3.4105
R5354 VDD.n2378 VDD.n2377 3.4105
R5355 VDD.n2356 VDD.n1602 3.4105
R5356 VDD.n2374 VDD.n1593 3.4105
R5357 VDD.n2400 VDD.n2399 3.4105
R5358 VDD.n2379 VDD.n1590 3.4105
R5359 VDD.n2381 VDD.n2380 3.4105
R5360 VDD.n2420 VDD.n2419 3.4105
R5361 VDD.n2401 VDD.n1576 3.4105
R5362 VDD.n2403 VDD.n2402 3.4105
R5363 VDD.n2439 VDD.n2438 3.4105
R5364 VDD.n2421 VDD.n1565 3.4105
R5365 VDD.n2423 VDD.n2422 3.4105
R5366 VDD.n2337 VDD.n2336 3.4105
R5367 VDD.n1614 VDD.n1613 3.4105
R5368 VDD.n2334 VDD.n2333 3.4105
R5369 VDD.n2327 VDD.n2326 3.4105
R5370 VDD.n1618 VDD.n1617 3.4105
R5371 VDD.n2325 VDD.n1616 3.4105
R5372 VDD.n2303 VDD.n2302 3.4105
R5373 VDD.n1631 VDD.n1630 3.4105
R5374 VDD.n2301 VDD.n1629 3.4105
R5375 VDD.n2282 VDD.n2281 3.4105
R5376 VDD.n2276 VDD.n1647 3.4105
R5377 VDD.n2280 VDD.n1646 3.4105
R5378 VDD.n2275 VDD.n2274 3.4105
R5379 VDD.n2244 VDD.n2242 3.4105
R5380 VDD.n2273 VDD.n2272 3.4105
R5381 VDD.n2246 VDD.n2245 3.4105
R5382 VDD.n2240 VDD.n2239 3.4105
R5383 VDD.n2248 VDD.n2247 3.4105
R5384 VDD.n2237 VDD.n1663 3.4105
R5385 VDD.n2214 VDD.n1677 3.4105
R5386 VDD.n2215 VDD.n1664 3.4105
R5387 VDD.n2132 VDD.n2131 3.4105
R5388 VDD.n1738 VDD.n1737 3.4105
R5389 VDD.n2128 VDD.n2127 3.4105
R5390 VDD.n2152 VDD.n2151 3.4105
R5391 VDD.n2130 VDD.n1736 3.4105
R5392 VDD.n2148 VDD.n1727 3.4105
R5393 VDD.n2174 VDD.n2173 3.4105
R5394 VDD.n2153 VDD.n1724 3.4105
R5395 VDD.n2155 VDD.n2154 3.4105
R5396 VDD.n2194 VDD.n2193 3.4105
R5397 VDD.n2175 VDD.n1710 3.4105
R5398 VDD.n2177 VDD.n2176 3.4105
R5399 VDD.n2213 VDD.n2212 3.4105
R5400 VDD.n2195 VDD.n1699 3.4105
R5401 VDD.n2197 VDD.n2196 3.4105
R5402 VDD.n2111 VDD.n2110 3.4105
R5403 VDD.n1748 VDD.n1747 3.4105
R5404 VDD.n2108 VDD.n2107 3.4105
R5405 VDD.n2101 VDD.n2100 3.4105
R5406 VDD.n1752 VDD.n1751 3.4105
R5407 VDD.n2099 VDD.n1750 3.4105
R5408 VDD.n2077 VDD.n2076 3.4105
R5409 VDD.n1765 VDD.n1764 3.4105
R5410 VDD.n2075 VDD.n1763 3.4105
R5411 VDD.n2056 VDD.n2055 3.4105
R5412 VDD.n2050 VDD.n1781 3.4105
R5413 VDD.n2054 VDD.n1780 3.4105
R5414 VDD.n2049 VDD.n2048 3.4105
R5415 VDD.n2018 VDD.n2016 3.4105
R5416 VDD.n2047 VDD.n2046 3.4105
R5417 VDD.n2020 VDD.n2019 3.4105
R5418 VDD.n2014 VDD.n2013 3.4105
R5419 VDD.n2022 VDD.n2021 3.4105
R5420 VDD.n2011 VDD.n1797 3.4105
R5421 VDD.n1988 VDD.n1811 3.4105
R5422 VDD.n1989 VDD.n1798 3.4105
R5423 VDD.n1926 VDD.n1925 3.4105
R5424 VDD.n1904 VDD.n1870 3.4105
R5425 VDD.n1922 VDD.n1861 3.4105
R5426 VDD.n1948 VDD.n1947 3.4105
R5427 VDD.n1927 VDD.n1858 3.4105
R5428 VDD.n1929 VDD.n1928 3.4105
R5429 VDD.n1968 VDD.n1967 3.4105
R5430 VDD.n1949 VDD.n1844 3.4105
R5431 VDD.n1951 VDD.n1950 3.4105
R5432 VDD.n1987 VDD.n1986 3.4105
R5433 VDD.n1969 VDD.n1833 3.4105
R5434 VDD.n1971 VDD.n1970 3.4105
R5435 VDD.n1902 VDD.n1901 3.4105
R5436 VDD.n1872 VDD.n1871 3.4105
R5437 VDD.n2884 VDD.n2883 3.4105
R5438 VDD.n2862 VDD.n1304 3.4105
R5439 VDD.n1306 VDD.n1305 3.4105
R5440 VDD.n2864 VDD.n2863 3.4105
R5441 VDD.n2844 VDD.n2843 3.4105
R5442 VDD.n1317 VDD.n1316 3.4105
R5443 VDD.n1328 VDD.n1327 3.4105
R5444 VDD.n2825 VDD.n2824 3.4105
R5445 VDD.n2806 VDD.n2805 3.4105
R5446 VDD.n1339 VDD.n1338 3.4105
R5447 VDD.n2787 VDD.n2786 3.4105
R5448 VDD.n2886 VDD.n2885 3.4105
R5449 VDD.n1286 VDD.n1284 3.4105
R5450 VDD.n2878 VDD.n1288 3.4105
R5451 VDD.n2861 VDD.n1303 3.4105
R5452 VDD.n2842 VDD.n1315 3.4105
R5453 VDD.n2823 VDD.n1326 3.4105
R5454 VDD.n2804 VDD.n1337 3.4105
R5455 VDD.n2782 VDD.n2781 3.4105
R5456 VDD.n2789 VDD.n2788 3.4105
R5457 VDD.n2866 VDD.n2865 3.4105
R5458 VDD.n2858 VDD.n2857 3.4105
R5459 VDD.n2846 VDD.n2845 3.4105
R5460 VDD.n2839 VDD.n2838 3.4105
R5461 VDD.n2827 VDD.n2826 3.4105
R5462 VDD.n2820 VDD.n2819 3.4105
R5463 VDD.n2808 VDD.n2807 3.4105
R5464 VDD.n2801 VDD.n2800 3.4105
R5465 VDD.n2785 VDD.n1348 3.4105
R5466 VDD.n2882 VDD.n2881 3.4105
R5467 VDD.n2877 VDD.n1292 3.4105
R5468 VDD.n3006 VDD.n3005 3.4105
R5469 VDD.n16 VDD.n15 3.4105
R5470 VDD.n18 VDD.n17 3.4105
R5471 VDD.n3004 VDD.n23 3.4105
R5472 VDD.n22 VDD.n21 3.4105
R5473 VDD.n3008 VDD.n3007 3.4105
R5474 VDD.n24 VDD.n22 3.4105
R5475 VDD.n1166 VDD.n930 3.40476
R5476 VDD.n117 VDD.n116 3.40476
R5477 VDD.n2680 VDD.n2677 3.38568
R5478 VDD.n2713 VDD.n1369 3.38568
R5479 VDD.n2454 VDD.n2451 3.38568
R5480 VDD.n2487 VDD.n1503 3.38568
R5481 VDD.n2544 VDD.n2538 3.38568
R5482 VDD.n2228 VDD.n2225 3.38568
R5483 VDD.n2261 VDD.n1637 3.38568
R5484 VDD.n2318 VDD.n2312 3.38568
R5485 VDD.n2002 VDD.n1999 3.38568
R5486 VDD.n2035 VDD.n1771 3.38568
R5487 VDD.n2092 VDD.n2086 3.38568
R5488 VDD.n2874 VDD.n2873 3.38568
R5489 VDD.n2640 VDD.n1426 3.38568
R5490 VDD.n2414 VDD.n1560 3.38568
R5491 VDD.n2188 VDD.n1694 3.38568
R5492 VDD.n1962 VDD.n1828 3.38568
R5493 VDD.n937 VDD.n936 3.36713
R5494 VDD.n2993 VDD.n29 3.31362
R5495 VDD.n165 VDD.n164 3.3098
R5496 VDD.n524 VDD.n523 3.29413
R5497 VDD.n2972 VDD.n2969 3.15412
R5498 VDD.n2989 VDD 3.15412
R5499 VDD.n717 VDD.n715 3.10575
R5500 VDD.n1894 VDD.n1875 3.10353
R5501 VDD.n1893 VDD.n1866 3.10353
R5502 VDD.n1915 VDD.n1864 3.10353
R5503 VDD.n1914 VDD.n1851 3.10353
R5504 VDD.n1855 VDD.n1852 3.10353
R5505 VDD.n1942 VDD.n1849 3.10353
R5506 VDD.n1957 VDD.n1840 3.10353
R5507 VDD.n1958 VDD.n1838 3.10353
R5508 VDD.n1977 VDD.n1829 3.10353
R5509 VDD.n1978 VDD.n1818 3.10353
R5510 VDD.n1827 VDD.n1826 3.10353
R5511 VDD.n1819 VDD.n1807 3.10353
R5512 VDD.n1806 VDD.n1803 3.10353
R5513 VDD.n2005 VDD.n2004 3.10353
R5514 VDD.n1805 VDD.n1804 3.10353
R5515 VDD.n2030 VDD.n1790 3.10353
R5516 VDD.n2037 VDD.n1788 3.10353
R5517 VDD.n2038 VDD.n1772 3.10353
R5518 VDD.n2063 VDD.n1770 3.10353
R5519 VDD.n1775 VDD.n1769 3.10353
R5520 VDD.n2084 VDD.n1760 3.10353
R5521 VDD.n2083 VDD.n1757 3.10353
R5522 VDD.n2089 VDD.n1758 3.10353
R5523 VDD.n2088 VDD.n1743 3.10353
R5524 VDD.n2120 VDD.n1741 3.10353
R5525 VDD.n2119 VDD.n1732 3.10353
R5526 VDD.n2141 VDD.n1730 3.10353
R5527 VDD.n2140 VDD.n1717 3.10353
R5528 VDD.n1721 VDD.n1718 3.10353
R5529 VDD.n2168 VDD.n1715 3.10353
R5530 VDD.n2183 VDD.n1706 3.10353
R5531 VDD.n2184 VDD.n1704 3.10353
R5532 VDD.n2203 VDD.n1695 3.10353
R5533 VDD.n2204 VDD.n1684 3.10353
R5534 VDD.n1693 VDD.n1692 3.10353
R5535 VDD.n1685 VDD.n1673 3.10353
R5536 VDD.n1672 VDD.n1669 3.10353
R5537 VDD.n2231 VDD.n2230 3.10353
R5538 VDD.n1671 VDD.n1670 3.10353
R5539 VDD.n2256 VDD.n1656 3.10353
R5540 VDD.n2263 VDD.n1654 3.10353
R5541 VDD.n2264 VDD.n1638 3.10353
R5542 VDD.n2289 VDD.n1636 3.10353
R5543 VDD.n1641 VDD.n1635 3.10353
R5544 VDD.n2310 VDD.n1626 3.10353
R5545 VDD.n2309 VDD.n1623 3.10353
R5546 VDD.n2315 VDD.n1624 3.10353
R5547 VDD.n2314 VDD.n1609 3.10353
R5548 VDD.n2346 VDD.n1607 3.10353
R5549 VDD.n2345 VDD.n1598 3.10353
R5550 VDD.n2367 VDD.n1596 3.10353
R5551 VDD.n2366 VDD.n1583 3.10353
R5552 VDD.n1587 VDD.n1584 3.10353
R5553 VDD.n2394 VDD.n1581 3.10353
R5554 VDD.n2409 VDD.n1572 3.10353
R5555 VDD.n2410 VDD.n1570 3.10353
R5556 VDD.n2429 VDD.n1561 3.10353
R5557 VDD.n2430 VDD.n1550 3.10353
R5558 VDD.n1559 VDD.n1558 3.10353
R5559 VDD.n1551 VDD.n1539 3.10353
R5560 VDD.n1538 VDD.n1535 3.10353
R5561 VDD.n2457 VDD.n2456 3.10353
R5562 VDD.n1537 VDD.n1536 3.10353
R5563 VDD.n2482 VDD.n1522 3.10353
R5564 VDD.n2489 VDD.n1520 3.10353
R5565 VDD.n2490 VDD.n1504 3.10353
R5566 VDD.n2515 VDD.n1502 3.10353
R5567 VDD.n1507 VDD.n1501 3.10353
R5568 VDD.n2536 VDD.n1492 3.10353
R5569 VDD.n2535 VDD.n1489 3.10353
R5570 VDD.n2541 VDD.n1490 3.10353
R5571 VDD.n2540 VDD.n1475 3.10353
R5572 VDD.n2572 VDD.n1473 3.10353
R5573 VDD.n2571 VDD.n1464 3.10353
R5574 VDD.n2593 VDD.n1462 3.10353
R5575 VDD.n2592 VDD.n1449 3.10353
R5576 VDD.n1453 VDD.n1450 3.10353
R5577 VDD.n2620 VDD.n1447 3.10353
R5578 VDD.n2635 VDD.n1438 3.10353
R5579 VDD.n2636 VDD.n1436 3.10353
R5580 VDD.n2655 VDD.n1427 3.10353
R5581 VDD.n2656 VDD.n1416 3.10353
R5582 VDD.n1425 VDD.n1424 3.10353
R5583 VDD.n1417 VDD.n1405 3.10353
R5584 VDD.n1404 VDD.n1401 3.10353
R5585 VDD.n2683 VDD.n2682 3.10353
R5586 VDD.n1403 VDD.n1402 3.10353
R5587 VDD.n2708 VDD.n1388 3.10353
R5588 VDD.n2715 VDD.n1386 3.10353
R5589 VDD.n2716 VDD.n1370 3.10353
R5590 VDD.n2741 VDD.n1368 3.10353
R5591 VDD.n1373 VDD.n1367 3.10353
R5592 VDD.n2767 VDD.n1357 3.10353
R5593 VDD.n2766 VDD.n1354 3.10353
R5594 VDD.n849 VDD.n848 3.10353
R5595 VDD.n1053 VDD.n1052 3.10353
R5596 VDD.n650 VDD.n649 3.10353
R5597 VDD.n542 VDD.n541 3.10353
R5598 VDD.n2794 VDD.n1345 3.10353
R5599 VDD.n2793 VDD.n1343 3.10353
R5600 VDD.n2813 VDD.n1334 3.10353
R5601 VDD.n2812 VDD.n1332 3.10353
R5602 VDD.n2832 VDD.n1323 3.10353
R5603 VDD.n2831 VDD.n1321 3.10353
R5604 VDD.n2851 VDD.n1312 3.10353
R5605 VDD.n2850 VDD.n1310 3.10353
R5606 VDD.n2871 VDD.n1300 3.10353
R5607 VDD.n2870 VDD.n1294 3.10353
R5608 VDD.n2989 VDD.n2988 3.1005
R5609 VDD.n861 VDD.n860 3.07837
R5610 VDD.n1257 VDD.n709 3.03311
R5611 VDD.n314 VDD.n283 3.03311
R5612 VDD.n6 VDD.n5 3.03311
R5613 VDD.n687 VDD.n686 3.02758
R5614 VDD VDD.n852 3.02729
R5615 VDD VDD.n1056 3.02729
R5616 VDD VDD.n653 3.02729
R5617 VDD.n546 VDD.n545 3.01836
R5618 VDD.n1046 VDD.n1040 3.01733
R5619 VDD.n830 VDD.n721 2.9753
R5620 VDD.n2974 VDD.n2973 2.96862
R5621 VDD.n32 VDD.t172 2.96725
R5622 VDD.n971 VDD.n967 2.95435
R5623 VDD.n1216 VDD.n780 2.95435
R5624 VDD.n203 VDD.n202 2.95435
R5625 VDD.n858 VDD.n857 2.92171
R5626 VDD.n1044 VDD.n1043 2.92171
R5627 VDD.n659 VDD.n658 2.92171
R5628 VDD.n552 VDD.n551 2.92171
R5629 VDD.n1077 VDD 2.89456
R5630 VDD.n817 VDD 2.89456
R5631 VDD.n159 VDD 2.89456
R5632 VDD.n518 VDD 2.89456
R5633 VDD.n969 VDD.t31 2.87059
R5634 VDD.n982 VDD 2.87059
R5635 VDD.n208 VDD.t213 2.87059
R5636 VDD.n493 VDD.n492 2.85588
R5637 VDD.n661 VDD.n644 2.80926
R5638 VDD.n555 VDD.n554 2.80434
R5639 VDD.n2954 VDD 2.73742
R5640 VDD.n3014 VDD.n3013 2.64177
R5641 VDD.n1117 VDD.n1116 2.62088
R5642 VDD.n2779 VDD.n2778 2.5429
R5643 VDD.n1078 VDD.n1076 2.52171
R5644 VDD.n818 VDD.n816 2.52171
R5645 VDD.n160 VDD.n158 2.52171
R5646 VDD.n519 VDD.n517 2.52171
R5647 VDD.n2998 VDD.n5 2.4386
R5648 VDD.n732 VDD.n731 2.3854
R5649 VDD.n99 VDD.n98 2.3854
R5650 VDD.n1119 VDD.n1118 2.3255
R5651 VDD.n731 VDD.n725 2.3255
R5652 VDD.n739 VDD.n738 2.3255
R5653 VDD.n741 VDD.n740 2.3255
R5654 VDD.n746 VDD.n745 2.3255
R5655 VDD.n720 VDD.n718 2.3255
R5656 VDD.n1248 VDD.n1247 2.3255
R5657 VDD.n832 VDD.n831 2.3255
R5658 VDD.n1241 VDD.n1240 2.3255
R5659 VDD.n1239 VDD.n752 2.3255
R5660 VDD.n1237 VDD.n1236 2.3255
R5661 VDD.n759 VDD.n755 2.3255
R5662 VDD.n1231 VDD.n1230 2.3255
R5663 VDD.n1229 VDD.n764 2.3255
R5664 VDD.n1228 VDD.n1227 2.3255
R5665 VDD.n775 VDD.n773 2.3255
R5666 VDD.n1221 VDD.n1220 2.3255
R5667 VDD.n1218 VDD.n774 2.3255
R5668 VDD.n1217 VDD.n1216 2.3255
R5669 VDD.n785 VDD.n781 2.3255
R5670 VDD.n1210 VDD.n1209 2.3255
R5671 VDD.n1208 VDD.n784 2.3255
R5672 VDD.n1207 VDD.n1206 2.3255
R5673 VDD.n795 VDD.n791 2.3255
R5674 VDD.n1199 VDD.n1198 2.3255
R5675 VDD.n1197 VDD.n1196 2.3255
R5676 VDD.n1195 VDD.n1194 2.3255
R5677 VDD.n919 VDD.n916 2.3255
R5678 VDD.n907 VDD.n904 2.3255
R5679 VDD.n1180 VDD.n905 2.3255
R5680 VDD.n933 VDD.n932 2.3255
R5681 VDD.n1167 VDD.n1166 2.3255
R5682 VDD.n941 VDD.n940 2.3255
R5683 VDD.n1029 VDD.n1028 2.3255
R5684 VDD.n948 VDD.n944 2.3255
R5685 VDD.n1156 VDD.n1155 2.3255
R5686 VDD.n1153 VDD.n1152 2.3255
R5687 VDD.n1151 VDD.n950 2.3255
R5688 VDD.n1085 VDD.n951 2.3255
R5689 VDD.n962 VDD.n961 2.3255
R5690 VDD.n1144 VDD.n1143 2.3255
R5691 VDD.n1141 VDD.n1140 2.3255
R5692 VDD.n1139 VDD.n964 2.3255
R5693 VDD.n973 VDD.n971 2.3255
R5694 VDD.n1133 VDD.n1132 2.3255
R5695 VDD.n1131 VDD.n1130 2.3255
R5696 VDD.n1129 VDD.n1128 2.3255
R5697 VDD.n1127 VDD.n1126 2.3255
R5698 VDD.n1108 VDD.n1107 2.3255
R5699 VDD.n467 VDD.n445 2.3255
R5700 VDD.n392 VDD.n390 2.3255
R5701 VDD.n499 VDD.n498 2.3255
R5702 VDD.n237 VDD.n218 2.3255
R5703 VDD.n289 VDD.n236 2.3255
R5704 VDD.n583 VDD.n582 2.3255
R5705 VDD.n265 VDD.n261 2.3255
R5706 VDD.n572 VDD.n571 2.3255
R5707 VDD.n365 VDD.n364 2.3255
R5708 VDD.n367 VDD.n366 2.3255
R5709 VDD.n369 VDD.n368 2.3255
R5710 VDD.n372 VDD.n371 2.3255
R5711 VDD.n412 VDD.n410 2.3255
R5712 VDD.n505 VDD.n334 2.3255
R5713 VDD.n507 VDD.n506 2.3255
R5714 VDD.n349 VDD.n348 2.3255
R5715 VDD.n266 VDD.n264 2.3255
R5716 VDD.n356 VDD.n355 2.3255
R5717 VDD.n302 VDD.n301 2.3255
R5718 VDD.n257 VDD.n255 2.3255
R5719 VDD.n586 VDD.n585 2.3255
R5720 VDD.n288 VDD.n250 2.3255
R5721 VDD.n235 VDD.n233 2.3255
R5722 VDD.n224 VDD.n214 2.3255
R5723 VDD.n609 VDD.n196 2.3255
R5724 VDD.n203 VDD.n195 2.3255
R5725 VDD.n145 VDD.n143 2.3255
R5726 VDD.n623 VDD.n622 2.3255
R5727 VDD.n625 VDD.n624 2.3255
R5728 VDD.n174 VDD.n173 2.3255
R5729 VDD.n485 VDD.n484 2.3255
R5730 VDD.n496 VDD.n495 2.3255
R5731 VDD.n428 VDD.n383 2.3255
R5732 VDD.n430 VDD.n429 2.3255
R5733 VDD.n482 VDD.n481 2.3255
R5734 VDD.n447 VDD.n444 2.3255
R5735 VDD.n458 VDD.n457 2.3255
R5736 VDD.n100 VDD.n99 2.3255
R5737 VDD.n105 VDD.n104 2.3255
R5738 VDD.n103 VDD.n102 2.3255
R5739 VDD.n89 VDD.n88 2.3255
R5740 VDD.n119 VDD.n84 2.3255
R5741 VDD.n123 VDD.n122 2.3255
R5742 VDD.n125 VDD.n124 2.3255
R5743 VDD.n82 VDD.n81 2.3255
R5744 VDD.n80 VDD.n79 2.3255
R5745 VDD.n64 VDD.n62 2.3255
R5746 VDD.n636 VDD.n635 2.3255
R5747 VDD.n634 VDD.n633 2.3255
R5748 VDD.n177 VDD.n176 2.3255
R5749 VDD.n1295 VDD.n1282 2.28608
R5750 VDD.n276 VDD.n269 2.26295
R5751 VDD.n1262 VDD.n709 2.2521
R5752 VDD.n2914 VDD.n2894 2.24869
R5753 VDD.n2956 VDD.n2955 2.24869
R5754 VDD.n2935 VDD.n2924 2.24869
R5755 VDD.n2949 VDD.n2896 2.24869
R5756 VDD.n2941 VDD.n2895 2.24869
R5757 VDD.n860 VDD.n859 2.21917
R5758 VDD.n856 VDD 2.21917
R5759 VDD.n1046 VDD.n1045 2.21917
R5760 VDD.n1042 VDD 2.21917
R5761 VDD.n661 VDD.n660 2.21917
R5762 VDD.n657 VDD 2.21917
R5763 VDD.n554 VDD.n553 2.21917
R5764 VDD.n550 VDD 2.21917
R5765 VDD.n2992 VDD.n2991 2.17384
R5766 VDD.n2893 VDD.n1282 2.15377
R5767 VDD.n34 VDD.n30 2.10088
R5768 VDD.n2978 VDD.n2977 1.95502
R5769 VDD.n2986 VDD.n2985 1.94045
R5770 VDD.n1142 VDD.n963 1.94045
R5771 VDD.n897 VDD.n786 1.94045
R5772 VDD.n1031 VDD.n1030 1.94045
R5773 VDD.n808 VDD.n766 1.94045
R5774 VDD.n1267 VDD.n706 1.94045
R5775 VDD.n1170 VDD.n934 1.94045
R5776 VDD.n1154 VDD.n949 1.94045
R5777 VDD.n892 VDD.n777 1.94045
R5778 VDD.n1183 VDD.n903 1.94045
R5779 VDD.n989 VDD.n988 1.94045
R5780 VDD.n1272 VDD.n703 1.94045
R5781 VDD.n1250 VDD.n1249 1.94045
R5782 VDD.n835 VDD.n834 1.94045
R5783 VDD.n1238 VDD.n754 1.94045
R5784 VDD.n823 VDD.n765 1.94045
R5785 VDD.n1219 VDD.n776 1.94045
R5786 VDD.n1087 VDD.n1086 1.94045
R5787 VDD.n1098 VDD.n1097 1.94045
R5788 VDD.n1103 VDD.n974 1.94045
R5789 VDD.n1191 VDD.n798 1.94045
R5790 VDD.n180 VDD.n179 1.94045
R5791 VDD.n671 VDD.n56 1.94045
R5792 VDD.n470 VDD.n443 1.94045
R5793 VDD.n676 VDD.n53 1.94045
R5794 VDD.n63 VDD.n61 1.94045
R5795 VDD.n185 VDD.n141 1.94045
R5796 VDD.n146 VDD.n144 1.94045
R5797 VDD.n612 VDD.n194 1.94045
R5798 VDD.n222 VDD.n216 1.94045
R5799 VDD.n234 VDD.n232 1.94045
R5800 VDD.n584 VDD.n254 1.94045
R5801 VDD.n304 VDD.n303 1.94045
R5802 VDD.n570 VDD.n569 1.94045
R5803 VDD.n564 VDD.n323 1.94045
R5804 VDD.n531 VDD.n328 1.94045
R5805 VDD.n393 VDD.n391 1.94045
R5806 VDD.n433 VDD.n432 1.94045
R5807 VDD.n698 VDD.n42 1.94045
R5808 VDD.n693 VDD.n45 1.94045
R5809 VDD.n409 VDD.n403 1.94045
R5810 VDD.n399 VDD.n398 1.94045
R5811 VDD.n558 VDD.n535 1.94045
R5812 VDD.n2891 VDD.n2890 1.94045
R5813 VDD.n19 VDD.n0 1.94045
R5814 VDD.n3002 VDD.n3001 1.94045
R5815 VDD.n525 VDD.n510 1.93962
R5816 VDD.n1072 VDD 1.93354
R5817 VDD.n812 VDD 1.93354
R5818 VDD.n154 VDD 1.90675
R5819 VDD.n513 VDD 1.89336
R5820 VDD.n2953 VDD.n2952 1.87313
R5821 VDD.n1174 VDD.n1173 1.8605
R5822 VDD VDD.n1071 1.85098
R5823 VDD VDD.n153 1.85098
R5824 VDD VDD.n811 1.85046
R5825 VDD VDD.n512 1.85046
R5826 VDD.n2680 VDD.n2679 1.76521
R5827 VDD.n2742 VDD.n1369 1.76521
R5828 VDD.n2568 VDD.n1474 1.76521
R5829 VDD.n2589 VDD.n1463 1.76521
R5830 VDD.n2616 VDD.n1448 1.76521
R5831 VDD.n2619 VDD.n1437 1.76521
R5832 VDD.n2640 VDD.n2639 1.76521
R5833 VDD.n2454 VDD.n2453 1.76521
R5834 VDD.n2516 VDD.n1503 1.76521
R5835 VDD.n2544 VDD.n2543 1.76521
R5836 VDD.n2342 VDD.n1608 1.76521
R5837 VDD.n2363 VDD.n1597 1.76521
R5838 VDD.n2390 VDD.n1582 1.76521
R5839 VDD.n2393 VDD.n1571 1.76521
R5840 VDD.n2414 VDD.n2413 1.76521
R5841 VDD.n2228 VDD.n2227 1.76521
R5842 VDD.n2290 VDD.n1637 1.76521
R5843 VDD.n2318 VDD.n2317 1.76521
R5844 VDD.n2116 VDD.n1742 1.76521
R5845 VDD.n2137 VDD.n1731 1.76521
R5846 VDD.n2164 VDD.n1716 1.76521
R5847 VDD.n2167 VDD.n1705 1.76521
R5848 VDD.n2188 VDD.n2187 1.76521
R5849 VDD.n2002 VDD.n2001 1.76521
R5850 VDD.n2064 VDD.n1771 1.76521
R5851 VDD.n2092 VDD.n2091 1.76521
R5852 VDD.n1938 VDD.n1850 1.76521
R5853 VDD.n1941 VDD.n1839 1.76521
R5854 VDD.n1962 VDD.n1961 1.76521
R5855 VDD.n2777 VDD.n2776 1.76521
R5856 VDD.n2874 VDD.n1296 1.76521
R5857 VDD.n180 VDD.n171 1.70236
R5858 VDD.n527 VDD.n526 1.70236
R5859 VDD.n331 VDD.n330 1.70194
R5860 VDD.n2796 VDD.n1333 1.66612
R5861 VDD.n2815 VDD.n1322 1.66612
R5862 VDD.n2834 VDD.n1311 1.66612
R5863 VDD.n2853 VDD.n1299 1.66612
R5864 VDD.n1997 VDD.n1996 1.66612
R5865 VDD.n2034 VDD.n2033 1.66612
R5866 VDD.n2067 VDD.n1759 1.66612
R5867 VDD.n2223 VDD.n2222 1.66612
R5868 VDD.n2260 VDD.n2259 1.66612
R5869 VDD.n2293 VDD.n1625 1.66612
R5870 VDD.n2449 VDD.n2448 1.66612
R5871 VDD.n2486 VDD.n2485 1.66612
R5872 VDD.n2519 VDD.n1491 1.66612
R5873 VDD.n2675 VDD.n2674 1.66612
R5874 VDD.n2712 VDD.n2711 1.66612
R5875 VDD.n2745 VDD.n1356 1.66612
R5876 VDD.n2659 VDD.n2658 1.66612
R5877 VDD.n2433 VDD.n2432 1.66612
R5878 VDD.n2207 VDD.n2206 1.66612
R5879 VDD.n1981 VDD.n1980 1.66612
R5880 VDD.n1891 VDD.n1865 1.66612
R5881 VDD.n2954 VDD.t142 1.58503
R5882 VDD.n546 VDD 1.5824
R5883 VDD.n1180 VDD.n908 1.57588
R5884 VDD.n458 VDD 1.57588
R5885 VDD.n602 VDD.n601 1.53347
R5886 VDD.n277 VDD.n268 1.49861
R5887 VDD.n758 VDD.n752 1.47742
R5888 VDD.n79 VDD.n78 1.47742
R5889 VDD.n364 VDD.n346 1.47742
R5890 VDD.n1166 VDD.n1165 1.45298
R5891 VDD.n1247 VDD.n721 1.45298
R5892 VDD.n122 VDD.n73 1.45298
R5893 VDD.n354 VDD.n264 1.45298
R5894 VDD.n911 VDD 1.43555
R5895 VDD.n513 VDD 1.39336
R5896 VDD.n1081 VDD.n1080 1.37996
R5897 VDD.n154 VDD 1.37996
R5898 VDD.n1158 VDD.n1157 1.37896
R5899 VDD.n240 VDD.n239 1.37896
R5900 VDD.n821 VDD.n820 1.3755
R5901 VDD.n879 VDD.n822 1.37165
R5902 VDD.n1040 VDD.n1039 1.36384
R5903 VDD.n163 VDD.n162 1.36211
R5904 VDD.n644 VDD.n642 1.3585
R5905 VDD.n843 VDD.n841 1.35813
R5906 VDD.n1004 VDD.n1003 1.35607
R5907 VDD.n1261 VDD.n1260 1.35607
R5908 VDD.n2877 VDD.n2876 1.35607
R5909 VDD.n1909 VDD.n1908 1.35607
R5910 VDD.n1994 VDD.n1993 1.35607
R5911 VDD.n1794 VDD.n1793 1.35607
R5912 VDD.n1787 VDD.n1785 1.35607
R5913 VDD.n2061 VDD.n1774 1.35607
R5914 VDD.n2071 VDD.n2070 1.35607
R5915 VDD.n2095 VDD.n2094 1.35607
R5916 VDD.n2220 VDD.n2219 1.35607
R5917 VDD.n1660 VDD.n1659 1.35607
R5918 VDD.n1653 VDD.n1651 1.35607
R5919 VDD.n2287 VDD.n1640 1.35607
R5920 VDD.n2297 VDD.n2296 1.35607
R5921 VDD.n2321 VDD.n2320 1.35607
R5922 VDD.n2446 VDD.n2445 1.35607
R5923 VDD.n1526 VDD.n1525 1.35607
R5924 VDD.n1519 VDD.n1517 1.35607
R5925 VDD.n2513 VDD.n1506 1.35607
R5926 VDD.n2523 VDD.n2522 1.35607
R5927 VDD.n2547 VDD.n2546 1.35607
R5928 VDD.n2672 VDD.n2671 1.35607
R5929 VDD.n1392 VDD.n1391 1.35607
R5930 VDD.n1385 VDD.n1383 1.35607
R5931 VDD.n2739 VDD.n1372 1.35607
R5932 VDD.n2749 VDD.n2748 1.35607
R5933 VDD.n2771 VDD.n1353 1.35607
R5934 VDD.n2643 VDD.n2642 1.35607
R5935 VDD.n2623 VDD.n2622 1.35607
R5936 VDD.n2614 VDD.n1452 1.35607
R5937 VDD.n2587 VDD.n2586 1.35607
R5938 VDD.n2662 VDD.n2661 1.35607
R5939 VDD.n2566 VDD.n2565 1.35607
R5940 VDD.n2417 VDD.n2416 1.35607
R5941 VDD.n2397 VDD.n2396 1.35607
R5942 VDD.n2388 VDD.n1586 1.35607
R5943 VDD.n2361 VDD.n2360 1.35607
R5944 VDD.n2436 VDD.n2435 1.35607
R5945 VDD.n2340 VDD.n2339 1.35607
R5946 VDD.n2191 VDD.n2190 1.35607
R5947 VDD.n2171 VDD.n2170 1.35607
R5948 VDD.n2162 VDD.n1720 1.35607
R5949 VDD.n2135 VDD.n2134 1.35607
R5950 VDD.n2210 VDD.n2209 1.35607
R5951 VDD.n2114 VDD.n2113 1.35607
R5952 VDD.n1965 VDD.n1964 1.35607
R5953 VDD.n1945 VDD.n1944 1.35607
R5954 VDD.n1936 VDD.n1854 1.35607
R5955 VDD.n1984 VDD.n1983 1.35607
R5956 VDD.n1888 VDD.n1887 1.35607
R5957 VDD.n2857 VDD.n2856 1.35607
R5958 VDD.n2838 VDD.n2837 1.35607
R5959 VDD.n2819 VDD.n2818 1.35607
R5960 VDD.n2800 VDD.n2799 1.35607
R5961 VDD.n3010 VDD.n3009 1.35607
R5962 VDD.n1072 VDD 1.35318
R5963 VDD.n812 VDD 1.35318
R5964 VDD.n522 VDD.n521 1.34871
R5965 VDD.n2968 VDD.n36 1.29905
R5966 VDD.n1106 VDD.n977 1.2805
R5967 VDD.n201 VDD.n143 1.2805
R5968 VDD.n452 VDD.n390 1.2805
R5969 VDD.n831 VDD.n830 1.18204
R5970 VDD.n77 VDD.n64 1.18204
R5971 VDD.n181 VDD.n180 1.13877
R5972 VDD.n2756 VDD.n2755 1.13717
R5973 VDD.n1881 VDD.n1877 1.13717
R5974 VDD.n1351 VDD.n1350 1.13717
R5975 VDD.n2752 VDD.n2751 1.13717
R5976 VDD.n1365 VDD.n1360 1.13717
R5977 VDD.n2731 VDD.n2730 1.13717
R5978 VDD.n1378 VDD.n1376 1.13717
R5979 VDD.n1382 VDD.n1381 1.13717
R5980 VDD.n2724 VDD.n2723 1.13717
R5981 VDD.n2693 VDD.n1393 1.13717
R5982 VDD.n2701 VDD.n2700 1.13717
R5983 VDD.n2669 VDD.n2668 1.13717
R5984 VDD.n1408 VDD.n1396 1.13717
R5985 VDD.n2581 VDD.n1467 1.13717
R5986 VDD.n2579 VDD.n1466 1.13717
R5987 VDD.n2601 VDD.n1457 1.13717
R5988 VDD.n2600 VDD.n2599 1.13717
R5989 VDD.n1444 VDD.n1443 1.13717
R5990 VDD.n2607 VDD.n1445 1.13717
R5991 VDD.n1433 VDD.n1432 1.13717
R5992 VDD.n2629 VDD.n1434 1.13717
R5993 VDD.n1411 VDD.n1410 1.13717
R5994 VDD.n2649 VDD.n1412 1.13717
R5995 VDD.n2561 VDD.n1478 1.13717
R5996 VDD.n2559 VDD.n1477 1.13717
R5997 VDD.n2550 VDD.n2549 1.13717
R5998 VDD.n1486 VDD.n1482 1.13717
R5999 VDD.n2526 VDD.n2525 1.13717
R6000 VDD.n1499 VDD.n1495 1.13717
R6001 VDD.n2505 VDD.n2504 1.13717
R6002 VDD.n1512 VDD.n1510 1.13717
R6003 VDD.n1516 VDD.n1515 1.13717
R6004 VDD.n2498 VDD.n2497 1.13717
R6005 VDD.n2467 VDD.n1527 1.13717
R6006 VDD.n2475 VDD.n2474 1.13717
R6007 VDD.n2443 VDD.n2442 1.13717
R6008 VDD.n1542 VDD.n1530 1.13717
R6009 VDD.n2355 VDD.n1601 1.13717
R6010 VDD.n2353 VDD.n1600 1.13717
R6011 VDD.n2375 VDD.n1591 1.13717
R6012 VDD.n2374 VDD.n2373 1.13717
R6013 VDD.n1578 VDD.n1577 1.13717
R6014 VDD.n2381 VDD.n1579 1.13717
R6015 VDD.n1567 VDD.n1566 1.13717
R6016 VDD.n2403 VDD.n1568 1.13717
R6017 VDD.n1545 VDD.n1544 1.13717
R6018 VDD.n2423 VDD.n1546 1.13717
R6019 VDD.n2335 VDD.n1612 1.13717
R6020 VDD.n2333 VDD.n1611 1.13717
R6021 VDD.n2324 VDD.n2323 1.13717
R6022 VDD.n1620 VDD.n1616 1.13717
R6023 VDD.n2300 VDD.n2299 1.13717
R6024 VDD.n1633 VDD.n1629 1.13717
R6025 VDD.n2279 VDD.n2278 1.13717
R6026 VDD.n1646 VDD.n1644 1.13717
R6027 VDD.n1650 VDD.n1649 1.13717
R6028 VDD.n2272 VDD.n2271 1.13717
R6029 VDD.n2241 VDD.n1661 1.13717
R6030 VDD.n2249 VDD.n2248 1.13717
R6031 VDD.n2217 VDD.n2216 1.13717
R6032 VDD.n1676 VDD.n1664 1.13717
R6033 VDD.n2129 VDD.n1735 1.13717
R6034 VDD.n2127 VDD.n1734 1.13717
R6035 VDD.n2149 VDD.n1725 1.13717
R6036 VDD.n2148 VDD.n2147 1.13717
R6037 VDD.n1712 VDD.n1711 1.13717
R6038 VDD.n2155 VDD.n1713 1.13717
R6039 VDD.n1701 VDD.n1700 1.13717
R6040 VDD.n2177 VDD.n1702 1.13717
R6041 VDD.n1679 VDD.n1678 1.13717
R6042 VDD.n2197 VDD.n1680 1.13717
R6043 VDD.n2109 VDD.n1746 1.13717
R6044 VDD.n2107 VDD.n1745 1.13717
R6045 VDD.n2098 VDD.n2097 1.13717
R6046 VDD.n1754 VDD.n1750 1.13717
R6047 VDD.n2074 VDD.n2073 1.13717
R6048 VDD.n1767 VDD.n1763 1.13717
R6049 VDD.n2053 VDD.n2052 1.13717
R6050 VDD.n1780 VDD.n1778 1.13717
R6051 VDD.n1784 VDD.n1783 1.13717
R6052 VDD.n2046 VDD.n2045 1.13717
R6053 VDD.n2015 VDD.n1795 1.13717
R6054 VDD.n2023 VDD.n2022 1.13717
R6055 VDD.n1991 VDD.n1990 1.13717
R6056 VDD.n1810 VDD.n1798 1.13717
R6057 VDD.n1923 VDD.n1859 1.13717
R6058 VDD.n1922 VDD.n1921 1.13717
R6059 VDD.n1846 VDD.n1845 1.13717
R6060 VDD.n1929 VDD.n1847 1.13717
R6061 VDD.n1835 VDD.n1834 1.13717
R6062 VDD.n1951 VDD.n1836 1.13717
R6063 VDD.n1813 VDD.n1812 1.13717
R6064 VDD.n1971 VDD.n1814 1.13717
R6065 VDD.n1901 VDD.n1868 1.13717
R6066 VDD.n1903 VDD.n1869 1.13717
R6067 VDD.n1883 VDD.n1878 1.13717
R6068 VDD.n1290 VDD.n1289 1.13717
R6069 VDD.n2784 VDD.n2783 1.13717
R6070 VDD.n2803 VDD.n2802 1.13717
R6071 VDD.n2822 VDD.n2821 1.13717
R6072 VDD.n2841 VDD.n2840 1.13717
R6073 VDD.n2860 VDD.n2859 1.13717
R6074 VDD.n1308 VDD.n1303 1.13717
R6075 VDD.n1319 VDD.n1315 1.13717
R6076 VDD.n1330 VDD.n1326 1.13717
R6077 VDD.n1341 VDD.n1337 1.13717
R6078 VDD.n2780 VDD.n1348 1.13717
R6079 VDD.n2881 VDD.n2880 1.13717
R6080 VDD.n3008 VDD.n12 1.13717
R6081 VDD.n2944 VDD.n2921 1.13671
R6082 VDD.n1279 VDD.n1278 1.13462
R6083 VDD.n2913 VDD.n2912 1.13462
R6084 VDD.n2907 VDD.n2906 1.13005
R6085 VDD.n915 VDD.n796 1.08358
R6086 VDD.n609 VDD.n205 1.08358
R6087 VDD.n372 VDD.n343 1.08358
R6088 VDD.n312 VDD.n311 1.04507
R6089 VDD.n49 VDD.n48 1.04225
R6090 VDD.n2916 VDD.n2894 1.04017
R6091 VDD.n2957 VDD.n2956 1.04017
R6092 VDD.n2933 VDD.n2924 1.04017
R6093 VDD.n2949 VDD.n2948 1.04017
R6094 VDD.n2942 VDD.n2895 1.04017
R6095 VDD.n278 VDD.n277 1.03323
R6096 VDD.n3012 VDD.n5 1.01637
R6097 VDD.n411 VDD.n377 0.985115
R6098 VDD.n486 VDD.n386 0.985115
R6099 VDD.n176 VDD.n175 0.886654
R6100 VDD.n495 VDD.n494 0.886654
R6101 VDD.n468 VDD.n467 0.886654
R6102 VDD.n1081 VDD 0.882712
R6103 VDD.n821 VDD 0.880308
R6104 VDD.n163 VDD 0.873096
R6105 VDD.n25 VDD.n23 0.870766
R6106 VDD.n20 VDD.n18 0.870578
R6107 VDD VDD.t142 0.864791
R6108 VDD.n1170 VDD.n938 0.854208
R6109 VDD.n1088 VDD.n1087 0.854028
R6110 VDD.n668 VDD.n58 0.853705
R6111 VDD.n1060 VDD.n1034 0.853631
R6112 VDD.n47 VDD.n46 0.853592
R6113 VDD.n710 VDD.n708 0.853567
R6114 VDD.n307 VDD.n281 0.853567
R6115 VDD.n561 VDD.n325 0.853479
R6116 VDD.n867 VDD.n840 0.853372
R6117 VDD.n2930 VDD.n2926 0.853362
R6118 VDD.n569 VDD.n568 0.853335
R6119 VDD.n2900 VDD.n2899 0.853291
R6120 VDD.n2944 VDD.n2943 0.853
R6121 VDD.n990 VDD.n989 0.853
R6122 VDD.n835 VDD.n827 0.853
R6123 VDD.n1191 VDD.n1190 0.853
R6124 VDD.n1003 VDD.n1002 0.853
R6125 VDD.n1261 VDD.n708 0.853
R6126 VDD.n865 VDD.n864 0.853
R6127 VDD.n1061 VDD.n1036 0.853
R6128 VDD.n1002 VDD.n1001 0.853
R6129 VDD.n1190 VDD.n1189 0.853
R6130 VDD.n805 VDD.n804 0.853
R6131 VDD.n875 VDD.n824 0.853
R6132 VDD.n705 VDD.n704 0.853
R6133 VDD.n702 VDD.n701 0.853
R6134 VDD.n713 VDD.n711 0.853
R6135 VDD.n827 VDD.n826 0.853
R6136 VDD.n994 VDD.n993 0.853
R6137 VDD.n1092 VDD.n995 0.853
R6138 VDD.n887 VDD.n806 0.853
R6139 VDD.n1024 VDD.n938 0.853
R6140 VDD.n1065 VDD.n998 0.853
R6141 VDD.n1000 VDD.n999 0.853
R6142 VDD.n903 VDD.n902 0.853
R6143 VDD.n902 VDD.n901 0.853
R6144 VDD.n803 VDD.n802 0.853
R6145 VDD.n870 VDD.n825 0.853
R6146 VDD.n882 VDD.n807 0.853
R6147 VDD.n997 VDD.n996 0.853
R6148 VDD.n992 VDD.n991 0.853
R6149 VDD.n433 VDD.n396 0.853
R6150 VDD.n394 VDD.n393 0.853
R6151 VDD.n147 VDD.n146 0.853
R6152 VDD.n194 VDD.n193 0.853
R6153 VDD.n222 VDD.n219 0.853
R6154 VDD.n232 VDD.n231 0.853
R6155 VDD.n443 VDD.n442 0.853
R6156 VDD.n61 VDD.n60 0.853
R6157 VDD.n403 VDD.n402 0.853
R6158 VDD.n48 VDD.n47 0.853
R6159 VDD.n666 VDD.n665 0.853
R6160 VDD.n310 VDD.n281 0.853
R6161 VDD.n559 VDD.n558 0.853
R6162 VDD.n330 VDD.n329 0.853
R6163 VDD.n41 VDD.n40 0.853
R6164 VDD.n44 VDD.n43 0.853
R6165 VDD.n52 VDD.n51 0.853
R6166 VDD.n55 VDD.n54 0.853
R6167 VDD.n60 VDD.n59 0.853
R6168 VDD.n191 VDD.n147 0.853
R6169 VDD.n193 VDD.n192 0.853
R6170 VDD.n229 VDD.n219 0.853
R6171 VDD.n231 VDD.n230 0.853
R6172 VDD.n296 VDD.n287 0.853
R6173 VDD.n286 VDD.n285 0.853
R6174 VDD.n320 VDD.n279 0.853
R6175 VDD.n322 VDD.n321 0.853
R6176 VDD.n327 VDD.n326 0.853
R6177 VDD.n440 VDD.n394 0.853
R6178 VDD.n396 VDD.n395 0.853
R6179 VDD.n402 VDD.n401 0.853
R6180 VDD.n149 VDD.n148 0.853
R6181 VDD.n151 VDD.n150 0.853
R6182 VDD.n400 VDD.n399 0.853
R6183 VDD.n421 VDD.n400 0.853
R6184 VDD.n2947 VDD.n2946 0.853
R6185 VDD.n2946 VDD.n2945 0.853
R6186 VDD.n2934 VDD.n2923 0.853
R6187 VDD.n2923 VDD.n2910 0.853
R6188 VDD.n2983 VDD.n2982 0.853
R6189 VDD.n2962 VDD.n1277 0.853
R6190 VDD.n2959 VDD.n1281 0.853
R6191 VDD.n2919 VDD.n2915 0.853
R6192 VDD.n2888 VDD.n2887 0.853
R6193 VDD.n3009 VDD.n3008 0.853
R6194 VDD.n522 VDD 0.849557
R6195 VDD.n2781 VDD.n2779 0.849366
R6196 VDD.n1017 VDD.n1013 0.835283
R6197 VDD.n2996 VDD.n28 0.813198
R6198 VDD.n3014 VDD.n3012 0.813198
R6199 VDD.n495 VDD.n378 0.788192
R6200 VDD.n1174 VDD.n930 0.772131
R6201 VDD.n1113 VDD.n1112 0.683764
R6202 VDD.n474 VDD.n441 0.683764
R6203 VDD.n1251 VDD.n1250 0.683297
R6204 VDD.n859 VDD.n856 0.683167
R6205 VDD.n1045 VDD.n1042 0.683167
R6206 VDD.n660 VDD.n657 0.683167
R6207 VDD.n553 VDD.n550 0.683167
R6208 VDD.n1103 VDD.n1102 0.683034
R6209 VDD.n1099 VDD.n1098 0.683034
R6210 VDD.n888 VDD.n776 0.683034
R6211 VDD.n871 VDD.n754 0.683034
R6212 VDD.n1272 VDD.n1271 0.683034
R6213 VDD.n893 VDD.n892 0.683034
R6214 VDD.n1066 VDD.n949 0.683034
R6215 VDD.n1267 VDD.n1266 0.683034
R6216 VDD.n1031 VDD.n1027 0.683034
R6217 VDD.n897 VDD.n896 0.683034
R6218 VDD.n1093 VDD.n963 0.683034
R6219 VDD.n693 VDD.n692 0.683034
R6220 VDD.n698 VDD.n697 0.683034
R6221 VDD.n531 VDD.n530 0.683034
R6222 VDD.n564 VDD.n563 0.683034
R6223 VDD.n305 VDD.n304 0.683034
R6224 VDD.n297 VDD.n254 0.683034
R6225 VDD.n186 VDD.n185 0.683034
R6226 VDD.n676 VDD.n675 0.683034
R6227 VDD.n671 VDD.n670 0.683034
R6228 VDD.n19 VDD.n14 0.682713
R6229 VDD.n3003 VDD.n3002 0.682713
R6230 VDD.n2978 VDD.n2964 0.682697
R6231 VDD.n2985 VDD.n2984 0.682697
R6232 VDD.n2929 VDD.n2927 0.682697
R6233 VDD.n873 VDD.n823 0.682474
R6234 VDD.n883 VDD.n808 0.682474
R6235 VDD.n2890 VDD.n2889 0.682447
R6236 VDD.n2909 VDD.n2908 0.644064
R6237 VDD.n135 VDD.n68 0.591269
R6238 VDD.n610 VDD.n609 0.591269
R6239 VDD.n372 VDD.n342 0.591269
R6240 VDD.n413 VDD.n412 0.591269
R6241 VDD.n485 VDD.n387 0.591269
R6242 VDD.n455 VDD.n450 0.591269
R6243 VDD.t215 VDD.n2953 0.576694
R6244 VDD.n686 VDD.n50 0.557022
R6245 VDD.n117 VDD.n84 0.545181
R6246 VDD.n831 VDD.n751 0.492808
R6247 VDD.n916 VDD.n915 0.492808
R6248 VDD.n100 VDD.n95 0.492808
R6249 VDD.n637 VDD.n64 0.492808
R6250 VDD.n1355 VDD.n1298 0.432646
R6251 VDD.t0 VDD.t172 0.432646
R6252 VDD.n31 VDD.t0 0.419342
R6253 VDD.n3021 VDD.n3020 0.406849
R6254 VDD.n556 VDD 0.403278
R6255 VDD.n730 VDD.n729 0.394346
R6256 VDD.n621 VDD.n143 0.394346
R6257 VDD.n256 VDD.n253 0.394346
R6258 VDD.n479 VDD.n390 0.394346
R6259 VDD.n1078 VDD.n1077 0.373349
R6260 VDD.n818 VDD.n817 0.373349
R6261 VDD.n160 VDD.n159 0.373349
R6262 VDD.n519 VDD.n518 0.373349
R6263 VDD.n1756 VDD.n1744 0.314894
R6264 VDD.n1622 VDD.n1610 0.314894
R6265 VDD.n1488 VDD.n1476 0.314894
R6266 VDD.n1824 VDD.n1821 0.30353
R6267 VDD.n1690 VDD.n1687 0.30353
R6268 VDD.n1556 VDD.n1553 0.30353
R6269 VDD.n1422 VDD.n1419 0.30353
R6270 VDD.n1823 VDD.n1822 0.30353
R6271 VDD.n1689 VDD.n1688 0.30353
R6272 VDD.n1555 VDD.n1554 0.30353
R6273 VDD.n1421 VDD.n1420 0.30353
R6274 VDD.n791 VDD.n787 0.295885
R6275 VDD.n2105 VDD.n2103 0.288379
R6276 VDD.n2331 VDD.n2329 0.288379
R6277 VDD.n2557 VDD.n2555 0.288379
R6278 VDD.n273 VDD.n272 0.278761
R6279 VDD.n314 VDD.n313 0.278761
R6280 VDD.n2976 VDD 0.267102
R6281 VDD.n1080 VDD 0.259429
R6282 VDD.n820 VDD 0.259429
R6283 VDD.n852 VDD 0.259429
R6284 VDD.n1056 VDD 0.259429
R6285 VDD.n162 VDD 0.259429
R6286 VDD.n521 VDD 0.259429
R6287 VDD.n653 VDD 0.259429
R6288 VDD.n545 VDD 0.259429
R6289 VDD.n1276 VDD.n1275 0.240048
R6290 VDD.n2970 VDD 0.237479
R6291 VDD.n932 VDD.n929 0.22745
R6292 VDD.n746 VDD.n744 0.22745
R6293 VDD.n121 VDD.n84 0.22745
R6294 VDD.n2991 VDD.n33 0.219459
R6295 VDD.n1107 VDD.n1106 0.197423
R6296 VDD.n1107 VDD.n984 0.197423
R6297 VDD.n1119 VDD.n987 0.197423
R6298 VDD.n1199 VDD.n794 0.197423
R6299 VDD.n176 VDD.n135 0.197423
R6300 VDD.n592 VDD.n235 0.197423
R6301 VDD.n248 VDD.n236 0.197423
R6302 VDD.n467 VDD.n450 0.197423
R6303 VDD.n1889 VDD.n1875 0.194439
R6304 VDD.n1910 VDD.n1866 0.194439
R6305 VDD.n1910 VDD.n1864 0.194439
R6306 VDD.n1937 VDD.n1851 0.194439
R6307 VDD.n1937 VDD.n1852 0.194439
R6308 VDD.n1943 VDD.n1942 0.194439
R6309 VDD.n1943 VDD.n1840 0.194439
R6310 VDD.n1963 VDD.n1838 0.194439
R6311 VDD.n1963 VDD.n1829 0.194439
R6312 VDD.n1982 VDD.n1818 0.194439
R6313 VDD.n1982 VDD.n1827 0.194439
R6314 VDD.n1995 VDD.n1807 0.194439
R6315 VDD.n1995 VDD.n1806 0.194439
R6316 VDD.n2004 VDD.n2003 0.194439
R6317 VDD.n2003 VDD.n1805 0.194439
R6318 VDD.n2031 VDD.n2030 0.194439
R6319 VDD.n2031 VDD.n1788 0.194439
R6320 VDD.n2062 VDD.n1772 0.194439
R6321 VDD.n2063 VDD.n2062 0.194439
R6322 VDD.n2069 VDD.n1769 0.194439
R6323 VDD.n2069 VDD.n1760 0.194439
R6324 VDD.n2093 VDD.n1757 0.194439
R6325 VDD.n2093 VDD.n1758 0.194439
R6326 VDD.n2115 VDD.n1743 0.194439
R6327 VDD.n2115 VDD.n1741 0.194439
R6328 VDD.n2136 VDD.n1732 0.194439
R6329 VDD.n2136 VDD.n1730 0.194439
R6330 VDD.n2163 VDD.n1717 0.194439
R6331 VDD.n2163 VDD.n1718 0.194439
R6332 VDD.n2169 VDD.n2168 0.194439
R6333 VDD.n2169 VDD.n1706 0.194439
R6334 VDD.n2189 VDD.n1704 0.194439
R6335 VDD.n2189 VDD.n1695 0.194439
R6336 VDD.n2208 VDD.n1684 0.194439
R6337 VDD.n2208 VDD.n1693 0.194439
R6338 VDD.n2221 VDD.n1673 0.194439
R6339 VDD.n2221 VDD.n1672 0.194439
R6340 VDD.n2230 VDD.n2229 0.194439
R6341 VDD.n2229 VDD.n1671 0.194439
R6342 VDD.n2257 VDD.n2256 0.194439
R6343 VDD.n2257 VDD.n1654 0.194439
R6344 VDD.n2288 VDD.n1638 0.194439
R6345 VDD.n2289 VDD.n2288 0.194439
R6346 VDD.n2295 VDD.n1635 0.194439
R6347 VDD.n2295 VDD.n1626 0.194439
R6348 VDD.n2319 VDD.n1623 0.194439
R6349 VDD.n2319 VDD.n1624 0.194439
R6350 VDD.n2341 VDD.n1609 0.194439
R6351 VDD.n2341 VDD.n1607 0.194439
R6352 VDD.n2362 VDD.n1598 0.194439
R6353 VDD.n2362 VDD.n1596 0.194439
R6354 VDD.n2389 VDD.n1583 0.194439
R6355 VDD.n2389 VDD.n1584 0.194439
R6356 VDD.n2395 VDD.n2394 0.194439
R6357 VDD.n2395 VDD.n1572 0.194439
R6358 VDD.n2415 VDD.n1570 0.194439
R6359 VDD.n2415 VDD.n1561 0.194439
R6360 VDD.n2434 VDD.n1550 0.194439
R6361 VDD.n2434 VDD.n1559 0.194439
R6362 VDD.n2447 VDD.n1539 0.194439
R6363 VDD.n2447 VDD.n1538 0.194439
R6364 VDD.n2456 VDD.n2455 0.194439
R6365 VDD.n2455 VDD.n1537 0.194439
R6366 VDD.n2483 VDD.n2482 0.194439
R6367 VDD.n2483 VDD.n1520 0.194439
R6368 VDD.n2514 VDD.n1504 0.194439
R6369 VDD.n2515 VDD.n2514 0.194439
R6370 VDD.n2521 VDD.n1501 0.194439
R6371 VDD.n2521 VDD.n1492 0.194439
R6372 VDD.n2545 VDD.n1489 0.194439
R6373 VDD.n2545 VDD.n1490 0.194439
R6374 VDD.n2567 VDD.n1475 0.194439
R6375 VDD.n2567 VDD.n1473 0.194439
R6376 VDD.n2588 VDD.n1464 0.194439
R6377 VDD.n2588 VDD.n1462 0.194439
R6378 VDD.n2615 VDD.n1449 0.194439
R6379 VDD.n2615 VDD.n1450 0.194439
R6380 VDD.n2621 VDD.n2620 0.194439
R6381 VDD.n2621 VDD.n1438 0.194439
R6382 VDD.n2641 VDD.n1436 0.194439
R6383 VDD.n2641 VDD.n1427 0.194439
R6384 VDD.n2660 VDD.n1416 0.194439
R6385 VDD.n2660 VDD.n1425 0.194439
R6386 VDD.n2673 VDD.n1405 0.194439
R6387 VDD.n2673 VDD.n1404 0.194439
R6388 VDD.n2682 VDD.n2681 0.194439
R6389 VDD.n2681 VDD.n1403 0.194439
R6390 VDD.n2709 VDD.n2708 0.194439
R6391 VDD.n2709 VDD.n1386 0.194439
R6392 VDD.n2740 VDD.n1370 0.194439
R6393 VDD.n2741 VDD.n2740 0.194439
R6394 VDD.n2747 VDD.n1367 0.194439
R6395 VDD.n2747 VDD.n1357 0.194439
R6396 VDD.n2770 VDD.n1354 0.194439
R6397 VDD.n850 VDD.n849 0.194439
R6398 VDD.n848 VDD 0.194439
R6399 VDD.n1054 VDD.n1053 0.194439
R6400 VDD.n1052 VDD 0.194439
R6401 VDD.n651 VDD.n650 0.194439
R6402 VDD.n649 VDD 0.194439
R6403 VDD.n543 VDD.n542 0.194439
R6404 VDD.n541 VDD 0.194439
R6405 VDD.n2778 VDD.n1345 0.194439
R6406 VDD.n2798 VDD.n1343 0.194439
R6407 VDD.n2798 VDD.n1334 0.194439
R6408 VDD.n2817 VDD.n1332 0.194439
R6409 VDD.n2817 VDD.n1323 0.194439
R6410 VDD.n2836 VDD.n1321 0.194439
R6411 VDD.n2836 VDD.n1312 0.194439
R6412 VDD.n2855 VDD.n1310 0.194439
R6413 VDD.n2855 VDD.n1300 0.194439
R6414 VDD.n2875 VDD.n1294 0.194439
R6415 VDD.n2875 VDD.n1295 0.194439
R6416 VDD.n879 VDD.n878 0.188833
R6417 VDD.n2973 VDD.n2972 0.186007
R6418 VDD.n116 VDD.n113 0.18206
R6419 VDD.n575 VDD.n574 0.18206
R6420 VDD.n1275 VDD.n1274 0.169867
R6421 VDD.n2892 VDD.n2891 0.132407
R6422 VDD.n2891 VDD.n1283 0.127283
R6423 VDD.n880 VDD.n879 0.1205
R6424 VDD.n2961 VDD 0.103213
R6425 VDD.n1986 VDD.n1811 0.102103
R6426 VDD.n2212 VDD.n1677 0.102103
R6427 VDD.n2438 VDD.n1543 0.102103
R6428 VDD.n2664 VDD.n1409 0.102103
R6429 VDD.n2101 VDD.n1748 0.100721
R6430 VDD.n2327 VDD.n1614 0.100721
R6431 VDD.n2553 VDD.n1480 0.100721
R6432 VDD.n2775 VDD 0.100533
R6433 VDD.n1164 VDD.n941 0.0989615
R6434 VDD.n1158 VDD.n944 0.0989615
R6435 VDD.n1152 VDD.n947 0.0989615
R6436 VDD.n1140 VDD.n960 0.0989615
R6437 VDD.n1130 VDD.n972 0.0989615
R6438 VDD.n1129 VDD.n975 0.0989615
R6439 VDD.n1120 VDD.n1119 0.0989615
R6440 VDD.n729 VDD.n725 0.0989615
R6441 VDD.n1200 VDD.n1199 0.0989615
R6442 VDD.n921 VDD.n916 0.0989615
R6443 VDD.n917 VDD.n907 0.0989615
R6444 VDD.n1181 VDD.n1180 0.0989615
R6445 VDD.n102 VDD.n101 0.0989615
R6446 VDD.n83 VDD.n82 0.0989615
R6447 VDD.n79 VDD.n71 0.0989615
R6448 VDD.n636 VDD.n65 0.0989615
R6449 VDD.n626 VDD.n625 0.0989615
R6450 VDD.n622 VDD.n140 0.0989615
R6451 VDD.n204 VDD.n203 0.0989615
R6452 VDD.n214 VDD.n213 0.0989615
R6453 VDD.n603 VDD.n602 0.0989615
R6454 VDD.n237 VDD.n215 0.0989615
R6455 VDD.n240 VDD.n235 0.0989615
R6456 VDD.n591 VDD.n236 0.0989615
R6457 VDD.n250 VDD.n249 0.0989615
R6458 VDD.n582 VDD.n256 0.0989615
R6459 VDD.n581 VDD.n257 0.0989615
R6460 VDD.n506 VDD.n335 0.0989615
R6461 VDD.n412 VDD.n411 0.0989615
R6462 VDD.n492 VDD.n383 0.0989615
R6463 VDD.n486 VDD.n485 0.0989615
R6464 VDD.n481 VDD.n480 0.0989615
R6465 VDD.n453 VDD.n447 0.0989615
R6466 VDD.n459 VDD.n458 0.0989615
R6467 VDD.n3000 VDD.n27 0.0981562
R6468 VDD.n1988 VDD.n1987 0.0890769
R6469 VDD.n2214 VDD.n2213 0.0890769
R6470 VDD.n2440 VDD.n2439 0.0890769
R6471 VDD.n2666 VDD.n2665 0.0890769
R6472 VDD.n2711 VDD.n2710 0.0847059
R6473 VDD.n2746 VDD.n2745 0.0847059
R6474 VDD.n2485 VDD.n2484 0.0847059
R6475 VDD.n2520 VDD.n2519 0.0847059
R6476 VDD.n2259 VDD.n2258 0.0847059
R6477 VDD.n2294 VDD.n2293 0.0847059
R6478 VDD.n2033 VDD.n2032 0.0847059
R6479 VDD.n2068 VDD.n2067 0.0847059
R6480 VDD.n1911 VDD.n1865 0.0847059
R6481 VDD.n2797 VDD.n2796 0.0847059
R6482 VDD.n2816 VDD.n2815 0.0847059
R6483 VDD.n2835 VDD.n2834 0.0847059
R6484 VDD.n2854 VDD.n2853 0.0847059
R6485 VDD.n1082 VDD.n1081 0.0822308
R6486 VDD.n822 VDD.n812 0.0822308
R6487 VDD.n822 VDD.n821 0.0798269
R6488 VDD.n2878 VDD.n1284 0.0796667
R6489 VDD.n1082 VDD.n1072 0.0774231
R6490 VDD.n164 VDD.n154 0.0774231
R6491 VDD.n164 VDD.n163 0.0774231
R6492 VDD.n1080 VDD.n1079 0.076587
R6493 VDD.n820 VDD.n819 0.076587
R6494 VDD.n852 VDD.n851 0.076587
R6495 VDD.n1056 VDD.n1055 0.076587
R6496 VDD.n162 VDD.n161 0.076587
R6497 VDD.n521 VDD.n520 0.076587
R6498 VDD.n653 VDD.n652 0.076587
R6499 VDD.n545 VDD.n544 0.076587
R6500 VDD.n523 VDD.n513 0.0759717
R6501 VDD.n523 VDD.n522 0.0759717
R6502 VDD.n2987 VDD 0.0717891
R6503 VDD.n2963 VDD.n2961 0.0707339
R6504 VDD.n2791 VDD.n1346 0.0705758
R6505 VDD.n2810 VDD.n1335 0.0705758
R6506 VDD.n2829 VDD.n1324 0.0705758
R6507 VDD.n2848 VDD.n1313 0.0705758
R6508 VDD.n2868 VDD.n1301 0.0705758
R6509 VDD.n1896 VDD.n1867 0.0705758
R6510 VDD.n1917 VDD.n1853 0.0705758
R6511 VDD.n1932 VDD.n1848 0.0705758
R6512 VDD.n1955 VDD.n1837 0.0705758
R6513 VDD.n1975 VDD.n1816 0.0705758
R6514 VDD.n2007 VDD.n1801 0.0705758
R6515 VDD.n2026 VDD.n2025 0.0705758
R6516 VDD.n2043 VDD.n2042 0.0705758
R6517 VDD.n2060 VDD.n1777 0.0705758
R6518 VDD.n2081 VDD.n1761 0.0705758
R6519 VDD.n2122 VDD.n1733 0.0705758
R6520 VDD.n2143 VDD.n1719 0.0705758
R6521 VDD.n2158 VDD.n1714 0.0705758
R6522 VDD.n2181 VDD.n1703 0.0705758
R6523 VDD.n2201 VDD.n1682 0.0705758
R6524 VDD.n2233 VDD.n1667 0.0705758
R6525 VDD.n2252 VDD.n2251 0.0705758
R6526 VDD.n2269 VDD.n2268 0.0705758
R6527 VDD.n2286 VDD.n1643 0.0705758
R6528 VDD.n2307 VDD.n1627 0.0705758
R6529 VDD.n2348 VDD.n1599 0.0705758
R6530 VDD.n2369 VDD.n1585 0.0705758
R6531 VDD.n2384 VDD.n1580 0.0705758
R6532 VDD.n2407 VDD.n1569 0.0705758
R6533 VDD.n2427 VDD.n1548 0.0705758
R6534 VDD.n2459 VDD.n1533 0.0705758
R6535 VDD.n2478 VDD.n2477 0.0705758
R6536 VDD.n2495 VDD.n2494 0.0705758
R6537 VDD.n2512 VDD.n1509 0.0705758
R6538 VDD.n2533 VDD.n1493 0.0705758
R6539 VDD.n2574 VDD.n1465 0.0705758
R6540 VDD.n2595 VDD.n1451 0.0705758
R6541 VDD.n2610 VDD.n1446 0.0705758
R6542 VDD.n2633 VDD.n1435 0.0705758
R6543 VDD.n2653 VDD.n1414 0.0705758
R6544 VDD.n2685 VDD.n1399 0.0705758
R6545 VDD.n2704 VDD.n2703 0.0705758
R6546 VDD.n2721 VDD.n2720 0.0705758
R6547 VDD.n2738 VDD.n1375 0.0705758
R6548 VDD.n2764 VDD.n1358 0.0705758
R6549 VDD.n2987 VDD.n2986 0.063
R6550 VDD.n1250 VDD.n717 0.063
R6551 VDD.n2100 VDD 0.0619615
R6552 VDD.n2326 VDD 0.0619615
R6553 VDD.n2552 VDD 0.0619615
R6554 VDD VDD.n2774 0.0619615
R6555 VDD.n2971 VDD.n2970 0.0616979
R6556 VDD.n7 VDD.n0 0.0616979
R6557 VDD.n2988 VDD 0.0603958
R6558 VDD.n740 VDD.n739 0.0603958
R6559 VDD.n745 VDD.n718 0.0603958
R6560 VDD.n1240 VDD.n1239 0.0603958
R6561 VDD.n1237 VDD.n755 0.0603958
R6562 VDD.n1230 VDD.n1229 0.0603958
R6563 VDD.n1229 VDD.n1228 0.0603958
R6564 VDD.n1220 VDD.n775 0.0603958
R6565 VDD.n1218 VDD.n1217 0.0603958
R6566 VDD.n1209 VDD.n785 0.0603958
R6567 VDD.n1209 VDD.n1208 0.0603958
R6568 VDD.n1208 VDD.n1207 0.0603958
R6569 VDD.n1198 VDD.n795 0.0603958
R6570 VDD.n1198 VDD.n1197 0.0603958
R6571 VDD.n1173 VDD.n933 0.0603958
R6572 VDD.n1167 VDD.n940 0.0603958
R6573 VDD.n1029 VDD.n948 0.0603958
R6574 VDD.n1155 VDD.n948 0.0603958
R6575 VDD.n1153 VDD.n950 0.0603958
R6576 VDD.n1085 VDD.n962 0.0603958
R6577 VDD.n1143 VDD.n962 0.0603958
R6578 VDD.n1141 VDD.n964 0.0603958
R6579 VDD.n1132 VDD.n973 0.0603958
R6580 VDD.n1132 VDD.n1131 0.0603958
R6581 VDD.n1128 VDD.n1127 0.0603958
R6582 VDD.n1118 VDD.n1117 0.0603958
R6583 VDD.n104 VDD.n103 0.0603958
R6584 VDD.n124 VDD.n123 0.0603958
R6585 VDD.n81 VDD.n80 0.0603958
R6586 VDD.n635 VDD.n634 0.0603958
R6587 VDD.n624 VDD.n623 0.0603958
R6588 VDD.n289 VDD.n288 0.0603958
R6589 VDD.n583 VDD.n255 0.0603958
R6590 VDD.n302 VDD.n265 0.0603958
R6591 VDD.n571 VDD.n265 0.0603958
R6592 VDD.n355 VDD.n266 0.0603958
R6593 VDD.n365 VDD.n348 0.0603958
R6594 VDD.n366 VDD.n365 0.0603958
R6595 VDD.n507 VDD.n334 0.0603958
R6596 VDD.n430 VDD.n428 0.0603958
R6597 VDD VDD.n7 0.0603958
R6598 VDD.n775 VDD.n766 0.0597448
R6599 VDD.n1219 VDD.n1218 0.0597448
R6600 VDD.n920 VDD.n904 0.0597448
R6601 VDD.n739 VDD.n703 0.0590938
R6602 VDD.n369 VDD.n328 0.0590938
R6603 VDD.n3022 VDD.n0 0.0590938
R6604 VDD.n124 VDD.n56 0.0584427
R6605 VDD.n1171 VDD.n1170 0.0583704
R6606 VDD.n1287 VDD 0.0579444
R6607 VDD.n745 VDD.n706 0.0577917
R6608 VDD.n3001 VDD.n3000 0.0577917
R6609 VDD.n1899 VDD.n1897 0.0573182
R6610 VDD.n1919 VDD.n1918 0.0573182
R6611 VDD.n1933 VDD.n1931 0.0573182
R6612 VDD.n1954 VDD.n1953 0.0573182
R6613 VDD.n1974 VDD.n1973 0.0573182
R6614 VDD.n2009 VDD.n2008 0.0573182
R6615 VDD.n2027 VDD.n1792 0.0573182
R6616 VDD.n2041 VDD.n1786 0.0573182
R6617 VDD.n2058 VDD.n1779 0.0573182
R6618 VDD.n2080 VDD.n2079 0.0573182
R6619 VDD.n2125 VDD.n2123 0.0573182
R6620 VDD.n2145 VDD.n2144 0.0573182
R6621 VDD.n2159 VDD.n2157 0.0573182
R6622 VDD.n2180 VDD.n2179 0.0573182
R6623 VDD.n2200 VDD.n2199 0.0573182
R6624 VDD.n2235 VDD.n2234 0.0573182
R6625 VDD.n2253 VDD.n1658 0.0573182
R6626 VDD.n2267 VDD.n1652 0.0573182
R6627 VDD.n2284 VDD.n1645 0.0573182
R6628 VDD.n2306 VDD.n2305 0.0573182
R6629 VDD.n2351 VDD.n2349 0.0573182
R6630 VDD.n2371 VDD.n2370 0.0573182
R6631 VDD.n2385 VDD.n2383 0.0573182
R6632 VDD.n2406 VDD.n2405 0.0573182
R6633 VDD.n2426 VDD.n2425 0.0573182
R6634 VDD.n2461 VDD.n2460 0.0573182
R6635 VDD.n2479 VDD.n1524 0.0573182
R6636 VDD.n2493 VDD.n1518 0.0573182
R6637 VDD.n2510 VDD.n1511 0.0573182
R6638 VDD.n2532 VDD.n2531 0.0573182
R6639 VDD.n2577 VDD.n2575 0.0573182
R6640 VDD.n2597 VDD.n2596 0.0573182
R6641 VDD.n2611 VDD.n2609 0.0573182
R6642 VDD.n2632 VDD.n2631 0.0573182
R6643 VDD.n2652 VDD.n2651 0.0573182
R6644 VDD.n2687 VDD.n2686 0.0573182
R6645 VDD.n2705 VDD.n1390 0.0573182
R6646 VDD.n2719 VDD.n1384 0.0573182
R6647 VDD.n2736 VDD.n1377 0.0573182
R6648 VDD.n2763 VDD.n2761 0.0573182
R6649 VDD.n2790 VDD.n2789 0.0573182
R6650 VDD.n2809 VDD.n2808 0.0573182
R6651 VDD.n2828 VDD.n2827 0.0573182
R6652 VDD.n2847 VDD.n2846 0.0573182
R6653 VDD.n2867 VDD.n2866 0.0573182
R6654 VDD.n104 VDD.n42 0.0571406
R6655 VDD.n370 VDD.n369 0.0564896
R6656 VDD.n483 VDD.n482 0.0564896
R6657 VDD.n1191 VDD.n800 0.0553246
R6658 VDD.n498 VDD.n497 0.0551875
R6659 VDD.n457 VDD.n456 0.0551875
R6660 VDD.n173 VDD.n172 0.0545365
R6661 VDD.n303 VDD.n255 0.0545365
R6662 VDD.n1249 VDD.n1248 0.0532344
R6663 VDD.n224 VDD.n223 0.0532344
R6664 VDD.n498 VDD.n379 0.0532344
R6665 VDD.n1248 VDD.n719 0.0525833
R6666 VDD.n80 VDD.n74 0.0525833
R6667 VDD.n200 VDD.n195 0.0519323
R6668 VDD.n451 VDD.n444 0.0519323
R6669 VDD.n3006 VDD.n23 0.0517727
R6670 VDD.n1030 VDD.n940 0.0512812
R6671 VDD.n1154 VDD.n1153 0.0512812
R6672 VDD.n1127 VDD.n976 0.0506302
R6673 VDD.n238 VDD.n218 0.0506302
R6674 VDD.n933 VDD.n931 0.0499792
R6675 VDD.n1275 VDD.n700 0.0493412
R6676 VDD.n570 VDD.n266 0.0493281
R6677 VDD.n681 VDD.n48 0.0487456
R6678 VDD.n2977 VDD.n2976 0.0483516
R6679 VDD.n1084 VDD.n1083 0.0482941
R6680 VDD.n1238 VDD.n1237 0.048026
R6681 VDD.n600 VDD.n218 0.048026
R6682 VDD.n1261 VDD.n1255 0.0465526
R6683 VDD.n688 VDD.n48 0.0465526
R6684 VDD.n557 VDD.n536 0.0465526
R6685 VDD.n113 VDD.n89 0.0458901
R6686 VDD.n575 VDD.n261 0.0458901
R6687 VDD.n573 VDD.n572 0.0458901
R6688 VDD.n878 VDD.n823 0.0455
R6689 VDD.n880 VDD.n808 0.0455
R6690 VDD.n2890 VDD.n1284 0.0455
R6691 VDD.n225 VDD.n224 0.0447708
R6692 VDD.n1010 VDD.n1009 0.0443596
R6693 VDD.n1019 VDD.n1003 0.0443596
R6694 VDD.n434 VDD.n433 0.0443596
R6695 VDD.n317 VDD.n282 0.0443596
R6696 VDD.n558 VDD.n534 0.0443596
R6697 VDD.n1142 VDD.n1141 0.0441198
R6698 VDD.n173 VDD.n141 0.0441198
R6699 VDD.n1075 VDD.n1073 0.0439783
R6700 VDD.n815 VDD.n813 0.0439783
R6701 VDD.n845 VDD.n844 0.0439783
R6702 VDD.n1049 VDD.n1048 0.0439783
R6703 VDD.n157 VDD.n155 0.0439783
R6704 VDD.n516 VDD.n514 0.0439783
R6705 VDD.n646 VDD.n645 0.0439783
R6706 VDD.n538 VDD.n537 0.0439783
R6707 VDD.n18 VDD.n15 0.0438377
R6708 VDD.n2970 VDD.n37 0.0434688
R6709 VDD.n2779 VDD.n1346 0.0429036
R6710 VDD.n1184 VDD.n904 0.0428177
R6711 VDD.n88 VDD.n87 0.042644
R6712 VDD.n1118 VDD.n1115 0.0421667
R6713 VDD.n226 VDD.n222 0.0421667
R6714 VDD.n599 VDD.n217 0.0421667
R6715 VDD.n290 VDD.n289 0.0421667
R6716 VDD.n664 VDD.n643 0.0421667
R6717 VDD.n3005 VDD.n3004 0.041625
R6718 VDD.n1131 VDD.n974 0.0415156
R6719 VDD.n1097 VDD.n964 0.0408646
R6720 VDD.n120 VDD.n53 0.0408646
R6721 VDD.n623 VDD.n142 0.0408646
R6722 VDD.n482 VDD.n389 0.0408646
R6723 VDD.n3001 VDD 0.0408646
R6724 VDD.n2799 VDD.n1335 0.0402727
R6725 VDD.n2818 VDD.n1324 0.0402727
R6726 VDD.n2837 VDD.n1313 0.0402727
R6727 VDD.n2856 VDD.n1301 0.0402727
R6728 VDD.n2876 VDD.n1283 0.0402727
R6729 VDD.n1909 VDD.n1867 0.0402727
R6730 VDD.n1936 VDD.n1853 0.0402727
R6731 VDD.n1944 VDD.n1848 0.0402727
R6732 VDD.n1964 VDD.n1837 0.0402727
R6733 VDD.n1983 VDD.n1816 0.0402727
R6734 VDD.n1994 VDD.n1801 0.0402727
R6735 VDD.n2025 VDD.n1793 0.0402727
R6736 VDD.n2043 VDD.n1787 0.0402727
R6737 VDD.n2061 VDD.n2060 0.0402727
R6738 VDD.n2070 VDD.n1761 0.0402727
R6739 VDD.n2094 VDD.n1756 0.0402727
R6740 VDD.n2114 VDD.n1744 0.0402727
R6741 VDD.n2135 VDD.n1733 0.0402727
R6742 VDD.n2162 VDD.n1719 0.0402727
R6743 VDD.n2170 VDD.n1714 0.0402727
R6744 VDD.n2190 VDD.n1703 0.0402727
R6745 VDD.n2209 VDD.n1682 0.0402727
R6746 VDD.n2220 VDD.n1667 0.0402727
R6747 VDD.n2251 VDD.n1659 0.0402727
R6748 VDD.n2269 VDD.n1653 0.0402727
R6749 VDD.n2287 VDD.n2286 0.0402727
R6750 VDD.n2296 VDD.n1627 0.0402727
R6751 VDD.n2320 VDD.n1622 0.0402727
R6752 VDD.n2340 VDD.n1610 0.0402727
R6753 VDD.n2361 VDD.n1599 0.0402727
R6754 VDD.n2388 VDD.n1585 0.0402727
R6755 VDD.n2396 VDD.n1580 0.0402727
R6756 VDD.n2416 VDD.n1569 0.0402727
R6757 VDD.n2435 VDD.n1548 0.0402727
R6758 VDD.n2446 VDD.n1533 0.0402727
R6759 VDD.n2477 VDD.n1525 0.0402727
R6760 VDD.n2495 VDD.n1519 0.0402727
R6761 VDD.n2513 VDD.n2512 0.0402727
R6762 VDD.n2522 VDD.n1493 0.0402727
R6763 VDD.n2546 VDD.n1488 0.0402727
R6764 VDD.n2566 VDD.n1476 0.0402727
R6765 VDD.n2587 VDD.n1465 0.0402727
R6766 VDD.n2614 VDD.n1451 0.0402727
R6767 VDD.n2622 VDD.n1446 0.0402727
R6768 VDD.n2642 VDD.n1435 0.0402727
R6769 VDD.n2661 VDD.n1414 0.0402727
R6770 VDD.n2672 VDD.n1399 0.0402727
R6771 VDD.n2703 VDD.n1391 0.0402727
R6772 VDD.n2721 VDD.n1385 0.0402727
R6773 VDD.n2739 VDD.n2738 0.0402727
R6774 VDD.n2748 VDD.n1358 0.0402727
R6775 VDD.n1897 VDD.n1873 0.0402727
R6776 VDD.n1918 VDD.n1862 0.0402727
R6777 VDD.n1934 VDD.n1933 0.0402727
R6778 VDD.n1954 VDD.n1842 0.0402727
R6779 VDD.n1974 VDD.n1831 0.0402727
R6780 VDD.n1823 VDD.n1815 0.0402727
R6781 VDD.n1822 VDD.n1809 0.0402727
R6782 VDD.n2008 VDD.n1800 0.0402727
R6783 VDD.n2028 VDD.n2027 0.0402727
R6784 VDD.n2041 VDD.n2040 0.0402727
R6785 VDD.n1779 VDD.n1766 0.0402727
R6786 VDD.n2080 VDD.n1753 0.0402727
R6787 VDD.n2123 VDD.n1739 0.0402727
R6788 VDD.n2144 VDD.n1728 0.0402727
R6789 VDD.n2160 VDD.n2159 0.0402727
R6790 VDD.n2180 VDD.n1708 0.0402727
R6791 VDD.n2200 VDD.n1697 0.0402727
R6792 VDD.n1689 VDD.n1681 0.0402727
R6793 VDD.n1688 VDD.n1675 0.0402727
R6794 VDD.n2234 VDD.n1666 0.0402727
R6795 VDD.n2254 VDD.n2253 0.0402727
R6796 VDD.n2267 VDD.n2266 0.0402727
R6797 VDD.n1645 VDD.n1632 0.0402727
R6798 VDD.n2306 VDD.n1619 0.0402727
R6799 VDD.n2349 VDD.n1605 0.0402727
R6800 VDD.n2370 VDD.n1594 0.0402727
R6801 VDD.n2386 VDD.n2385 0.0402727
R6802 VDD.n2406 VDD.n1574 0.0402727
R6803 VDD.n2426 VDD.n1563 0.0402727
R6804 VDD.n1555 VDD.n1547 0.0402727
R6805 VDD.n1554 VDD.n1541 0.0402727
R6806 VDD.n2460 VDD.n1532 0.0402727
R6807 VDD.n2480 VDD.n2479 0.0402727
R6808 VDD.n2493 VDD.n2492 0.0402727
R6809 VDD.n1511 VDD.n1498 0.0402727
R6810 VDD.n2532 VDD.n1485 0.0402727
R6811 VDD.n2575 VDD.n1471 0.0402727
R6812 VDD.n2596 VDD.n1460 0.0402727
R6813 VDD.n2612 VDD.n2611 0.0402727
R6814 VDD.n2632 VDD.n1440 0.0402727
R6815 VDD.n2652 VDD.n1429 0.0402727
R6816 VDD.n1421 VDD.n1413 0.0402727
R6817 VDD.n1420 VDD.n1407 0.0402727
R6818 VDD.n2686 VDD.n1398 0.0402727
R6819 VDD.n2706 VDD.n2705 0.0402727
R6820 VDD.n2719 VDD.n2718 0.0402727
R6821 VDD.n1377 VDD.n1364 0.0402727
R6822 VDD.n2763 VDD.n2762 0.0402727
R6823 VDD.n2790 VDD.n1340 0.0402727
R6824 VDD.n2809 VDD.n1329 0.0402727
R6825 VDD.n2828 VDD.n1318 0.0402727
R6826 VDD.n2847 VDD.n1307 0.0402727
R6827 VDD.n2867 VDD.n1291 0.0402727
R6828 VDD.n1240 VDD.n753 0.0402135
R6829 VDD.n635 VDD.n66 0.0402135
R6830 VDD.n863 VDD.n842 0.0399737
R6831 VDD.n1059 VDD.n1037 0.0399737
R6832 VDD.n446 VDD.n443 0.0399737
R6833 VDD.n795 VDD.n786 0.0395625
R6834 VDD.n613 VDD.n195 0.0395625
R6835 VDD.n408 VDD.n334 0.0395625
R6836 VDD.n1260 VDD.n1259 0.0389615
R6837 VDD.n275 VDD.n270 0.0389615
R6838 VDD.n316 VDD.n283 0.0389615
R6839 VDD.n569 VDD.n278 0.0388523
R6840 VDD.n634 VDD.n67 0.0382604
R6841 VDD.n418 VDD.n399 0.0377807
R6842 VDD.n555 VDD.n547 0.0377545
R6843 VDD.n428 VDD.n427 0.0376094
R6844 VDD.n471 VDD.n444 0.0376094
R6845 VDD.n180 VDD.n166 0.0374318
R6846 VDD.n1086 VDD.n950 0.0369583
R6847 VDD.n355 VDD.n323 0.0369583
R6848 VDD.n1877 VDD.n1876 0.0364848
R6849 VDD.n1898 VDD.n1868 0.0364848
R6850 VDD.n1921 VDD.n1920 0.0364848
R6851 VDD.n1857 VDD.n1847 0.0364848
R6852 VDD.n1843 VDD.n1836 0.0364848
R6853 VDD.n1832 VDD.n1814 0.0364848
R6854 VDD.n1810 VDD.n1799 0.0364848
R6855 VDD.n2024 VDD.n2023 0.0364848
R6856 VDD.n2045 VDD.n2044 0.0364848
R6857 VDD.n2059 VDD.n1778 0.0364848
R6858 VDD.n1767 VDD.n1762 0.0364848
R6859 VDD.n1754 VDD.n1749 0.0364848
R6860 VDD.n2104 VDD.n1745 0.0364848
R6861 VDD.n2124 VDD.n1734 0.0364848
R6862 VDD.n2147 VDD.n2146 0.0364848
R6863 VDD.n1723 VDD.n1713 0.0364848
R6864 VDD.n1709 VDD.n1702 0.0364848
R6865 VDD.n1698 VDD.n1680 0.0364848
R6866 VDD.n1676 VDD.n1665 0.0364848
R6867 VDD.n2250 VDD.n2249 0.0364848
R6868 VDD.n2271 VDD.n2270 0.0364848
R6869 VDD.n2285 VDD.n1644 0.0364848
R6870 VDD.n1633 VDD.n1628 0.0364848
R6871 VDD.n1620 VDD.n1615 0.0364848
R6872 VDD.n2330 VDD.n1611 0.0364848
R6873 VDD.n2350 VDD.n1600 0.0364848
R6874 VDD.n2373 VDD.n2372 0.0364848
R6875 VDD.n1589 VDD.n1579 0.0364848
R6876 VDD.n1575 VDD.n1568 0.0364848
R6877 VDD.n1564 VDD.n1546 0.0364848
R6878 VDD.n1542 VDD.n1531 0.0364848
R6879 VDD.n2476 VDD.n2475 0.0364848
R6880 VDD.n2497 VDD.n2496 0.0364848
R6881 VDD.n2511 VDD.n1510 0.0364848
R6882 VDD.n1499 VDD.n1494 0.0364848
R6883 VDD.n1486 VDD.n1481 0.0364848
R6884 VDD.n2556 VDD.n1477 0.0364848
R6885 VDD.n2576 VDD.n1466 0.0364848
R6886 VDD.n2599 VDD.n2598 0.0364848
R6887 VDD.n1455 VDD.n1445 0.0364848
R6888 VDD.n1441 VDD.n1434 0.0364848
R6889 VDD.n1430 VDD.n1412 0.0364848
R6890 VDD.n1408 VDD.n1397 0.0364848
R6891 VDD.n2702 VDD.n2701 0.0364848
R6892 VDD.n2723 VDD.n2722 0.0364848
R6893 VDD.n2737 VDD.n1376 0.0364848
R6894 VDD.n1365 VDD.n1359 0.0364848
R6895 VDD.n2772 VDD.n1351 0.0364848
R6896 VDD.n2780 VDD.n1347 0.0364848
R6897 VDD.n1341 VDD.n1336 0.0364848
R6898 VDD.n1330 VDD.n1325 0.0364848
R6899 VDD.n1319 VDD.n1314 0.0364848
R6900 VDD.n1308 VDD.n1302 0.0364848
R6901 VDD.n2880 VDD.n2879 0.0364848
R6902 VDD.n509 VDD.n507 0.0363073
R6903 VDD.n431 VDD.n430 0.0363073
R6904 VDD.n1075 VDD 0.0358261
R6905 VDD.n815 VDD 0.0358261
R6906 VDD.n845 VDD 0.0358261
R6907 VDD.n1049 VDD 0.0358261
R6908 VDD.n157 VDD 0.0358261
R6909 VDD.n516 VDD 0.0358261
R6910 VDD.n646 VDD 0.0358261
R6911 VDD.n538 VDD 0.0358261
R6912 VDD.n2988 VDD.n2987 0.0356562
R6913 VDD.n2976 VDD.n2975 0.0356562
R6914 VDD.n1230 VDD.n765 0.0356562
R6915 VDD.n585 VDD.n584 0.0356562
R6916 VDD.n1114 VDD.n989 0.0355877
R6917 VDD.n197 VDD.n194 0.0355877
R6918 VDD.n415 VDD.n403 0.0355877
R6919 VDD.n17 VDD.n16 0.0351948
R6920 VDD.n1217 VDD.n777 0.0350052
R6921 VDD.n1185 VDD.n903 0.0333947
R6922 VDD.n291 VDD.n232 0.0333947
R6923 VDD.n1194 VDD.n1193 0.0330521
R6924 VDD.n1168 VDD.n1167 0.032401
R6925 VDD.n88 VDD.n45 0.032401
R6926 VDD.n900 VDD.n899 0.0321887
R6927 VDD.n477 VDD.n393 0.0312018
R6928 VDD.n3009 VDD.n10 0.0309054
R6929 VDD.n2792 VDD.n1342 0.030803
R6930 VDD.n2811 VDD.n1331 0.030803
R6931 VDD.n2830 VDD.n1320 0.030803
R6932 VDD.n2849 VDD.n1309 0.030803
R6933 VDD.n2869 VDD.n1293 0.030803
R6934 VDD.n1895 VDD.n1874 0.030803
R6935 VDD.n1916 VDD.n1863 0.030803
R6936 VDD.n1935 VDD.n1856 0.030803
R6937 VDD.n1956 VDD.n1841 0.030803
R6938 VDD.n1976 VDD.n1830 0.030803
R6939 VDD.n1825 VDD.n1817 0.030803
R6940 VDD.n1820 VDD.n1808 0.030803
R6941 VDD.n2006 VDD.n1802 0.030803
R6942 VDD.n2029 VDD.n1791 0.030803
R6943 VDD.n2039 VDD.n1773 0.030803
R6944 VDD.n1776 VDD.n1768 0.030803
R6945 VDD.n2082 VDD.n1755 0.030803
R6946 VDD.n2121 VDD.n1740 0.030803
R6947 VDD.n2142 VDD.n1729 0.030803
R6948 VDD.n2161 VDD.n1722 0.030803
R6949 VDD.n2182 VDD.n1707 0.030803
R6950 VDD.n2202 VDD.n1696 0.030803
R6951 VDD.n1691 VDD.n1683 0.030803
R6952 VDD.n1686 VDD.n1674 0.030803
R6953 VDD.n2232 VDD.n1668 0.030803
R6954 VDD.n2255 VDD.n1657 0.030803
R6955 VDD.n2265 VDD.n1639 0.030803
R6956 VDD.n1642 VDD.n1634 0.030803
R6957 VDD.n2308 VDD.n1621 0.030803
R6958 VDD.n2347 VDD.n1606 0.030803
R6959 VDD.n2368 VDD.n1595 0.030803
R6960 VDD.n2387 VDD.n1588 0.030803
R6961 VDD.n2408 VDD.n1573 0.030803
R6962 VDD.n2428 VDD.n1562 0.030803
R6963 VDD.n1557 VDD.n1549 0.030803
R6964 VDD.n1552 VDD.n1540 0.030803
R6965 VDD.n2458 VDD.n1534 0.030803
R6966 VDD.n2481 VDD.n1523 0.030803
R6967 VDD.n2491 VDD.n1505 0.030803
R6968 VDD.n1508 VDD.n1500 0.030803
R6969 VDD.n2534 VDD.n1487 0.030803
R6970 VDD.n2573 VDD.n1472 0.030803
R6971 VDD.n2594 VDD.n1461 0.030803
R6972 VDD.n2613 VDD.n1454 0.030803
R6973 VDD.n2634 VDD.n1439 0.030803
R6974 VDD.n2654 VDD.n1428 0.030803
R6975 VDD.n1423 VDD.n1415 0.030803
R6976 VDD.n1418 VDD.n1406 0.030803
R6977 VDD.n2684 VDD.n1400 0.030803
R6978 VDD.n2707 VDD.n1389 0.030803
R6979 VDD.n2717 VDD.n1371 0.030803
R6980 VDD.n1374 VDD.n1366 0.030803
R6981 VDD.n2765 VDD.n1352 0.030803
R6982 VDD.n1194 VDD 0.0304479
R6983 VDD.n585 VDD 0.0304479
R6984 VDD.n861 VDD.n854 0.0299674
R6985 VDD.n26 VDD.n9 0.0292162
R6986 VDD.n835 VDD.n829 0.0290088
R6987 VDD.n836 VDD.n835 0.0290088
R6988 VDD.n188 VDD.n146 0.0290088
R6989 VDD.n619 VDD.n146 0.0290088
R6990 VDD.n639 VDD.n61 0.0290088
R6991 VDD.n167 VDD.n61 0.0290088
R6992 VDD.n103 VDD.n45 0.0284948
R6993 VDD.n895 VDD.n894 0.0283124
R6994 VDD.n525 VDD.n524 0.0280028
R6995 VDD.n1047 VDD.n1038 0.0271393
R6996 VDD.n437 VDD.n393 0.0268158
R6997 VDD.n8 VDD 0.0265417
R6998 VDD.n1262 VDD.n1261 0.0259749
R6999 VDD.n785 VDD.n777 0.0258906
R7000 VDD.n294 VDD.n293 0.0254052
R7001 VDD.n765 VDD.n755 0.0252396
R7002 VDD.n584 VDD.n583 0.0252396
R7003 VDD.n906 VDD.n903 0.0246228
R7004 VDD.n594 VDD.n232 0.0246228
R7005 VDD.n663 VDD.n662 0.0243971
R7006 VDD.n2915 VDD.n2914 0.0242893
R7007 VDD.n2955 VDD.n1281 0.0242893
R7008 VDD.n2935 VDD.n2934 0.0242893
R7009 VDD.n2947 VDD.n2896 0.0242893
R7010 VDD.n2943 VDD.n2941 0.0242893
R7011 VDD.n1086 VDD.n1085 0.0239375
R7012 VDD.n348 VDD.n323 0.0239375
R7013 VDD.n3010 VDD.n8 0.0239375
R7014 VDD.n2905 VDD.n2904 0.0234759
R7015 VDD VDD.n3022 0.0226354
R7016 VDD.n1110 VDD.n989 0.0224298
R7017 VDD.n614 VDD.n194 0.0224298
R7018 VDD.n407 VDD.n403 0.0224298
R7019 VDD.n1101 VDD.n1100 0.0215289
R7020 VDD.n2975 VDD.n2966 0.0213333
R7021 VDD.n1207 VDD.n786 0.0213333
R7022 VDD.n2885 VDD.n2884 0.0206084
R7023 VDD.n1886 VDD.n1885 0.0205441
R7024 VDD.n1907 VDD.n1906 0.0205441
R7025 VDD.n1925 VDD.n1924 0.0205441
R7026 VDD.n1947 VDD.n1946 0.0205441
R7027 VDD.n1967 VDD.n1966 0.0205441
R7028 VDD.n1986 VDD.n1985 0.0205441
R7029 VDD.n2112 VDD.n2111 0.0205441
R7030 VDD.n2133 VDD.n2132 0.0205441
R7031 VDD.n2151 VDD.n2150 0.0205441
R7032 VDD.n2173 VDD.n2172 0.0205441
R7033 VDD.n2193 VDD.n2192 0.0205441
R7034 VDD.n2212 VDD.n2211 0.0205441
R7035 VDD.n2338 VDD.n2337 0.0205441
R7036 VDD.n2359 VDD.n2358 0.0205441
R7037 VDD.n2377 VDD.n2376 0.0205441
R7038 VDD.n2399 VDD.n2398 0.0205441
R7039 VDD.n2419 VDD.n2418 0.0205441
R7040 VDD.n2438 VDD.n2437 0.0205441
R7041 VDD.n2564 VDD.n2563 0.0205441
R7042 VDD.n2585 VDD.n2584 0.0205441
R7043 VDD.n2603 VDD.n2602 0.0205441
R7044 VDD.n2625 VDD.n2624 0.0205441
R7045 VDD.n2645 VDD.n2644 0.0205441
R7046 VDD.n2664 VDD.n2663 0.0205441
R7047 VDD.n426 VDD.n399 0.0202368
R7048 VDD.n1097 VDD.n973 0.0200312
R7049 VDD.n1992 VDD.n1811 0.0198529
R7050 VDD.n2013 VDD.n2012 0.0198529
R7051 VDD.n2018 VDD.n2017 0.0198529
R7052 VDD.n2051 VDD.n2050 0.0198529
R7053 VDD.n2072 VDD.n1765 0.0198529
R7054 VDD.n2096 VDD.n1752 0.0198529
R7055 VDD.n2218 VDD.n1677 0.0198529
R7056 VDD.n2239 VDD.n2238 0.0198529
R7057 VDD.n2244 VDD.n2243 0.0198529
R7058 VDD.n2277 VDD.n2276 0.0198529
R7059 VDD.n2298 VDD.n1631 0.0198529
R7060 VDD.n2322 VDD.n1618 0.0198529
R7061 VDD.n2444 VDD.n1543 0.0198529
R7062 VDD.n2465 VDD.n2464 0.0198529
R7063 VDD.n2470 VDD.n2469 0.0198529
R7064 VDD.n2503 VDD.n2502 0.0198529
R7065 VDD.n2524 VDD.n1497 0.0198529
R7066 VDD.n2548 VDD.n1484 0.0198529
R7067 VDD.n2670 VDD.n1409 0.0198529
R7068 VDD.n2691 VDD.n2690 0.0198529
R7069 VDD.n2696 VDD.n2695 0.0198529
R7070 VDD.n2729 VDD.n2728 0.0198529
R7071 VDD.n2750 VDD.n1363 0.0198529
R7072 VDD.n2754 VDD.n1361 0.0198529
R7073 VDD.n2801 VDD.n1339 0.0198529
R7074 VDD.n2820 VDD.n1328 0.0198529
R7075 VDD.n2839 VDD.n1317 0.0198529
R7076 VDD.n2858 VDD.n1306 0.0198529
R7077 VDD.n1304 VDD.n1292 0.0198529
R7078 VDD.n2922 VDD.n39 0.0194294
R7079 VDD.n1128 VDD.n974 0.0193802
R7080 VDD.n3006 VDD.n12 0.0188117
R7081 VDD.n15 VDD.n12 0.0188117
R7082 VDD.n1884 VDD.n1883 0.0185769
R7083 VDD.n1905 VDD.n1903 0.0185769
R7084 VDD.n1926 VDD.n1859 0.0185769
R7085 VDD.n1948 VDD.n1845 0.0185769
R7086 VDD.n1968 VDD.n1834 0.0185769
R7087 VDD.n1987 VDD.n1812 0.0185769
R7088 VDD.n1989 VDD.n1797 0.0185769
R7089 VDD.n2021 VDD.n2020 0.0185769
R7090 VDD.n2048 VDD.n2047 0.0185769
R7091 VDD.n2055 VDD.n2054 0.0185769
R7092 VDD.n2076 VDD.n2075 0.0185769
R7093 VDD.n2100 VDD.n2099 0.0185769
R7094 VDD.n2110 VDD.n2109 0.0185769
R7095 VDD.n2131 VDD.n2129 0.0185769
R7096 VDD.n2152 VDD.n1725 0.0185769
R7097 VDD.n2174 VDD.n1711 0.0185769
R7098 VDD.n2194 VDD.n1700 0.0185769
R7099 VDD.n2213 VDD.n1678 0.0185769
R7100 VDD.n2215 VDD.n1663 0.0185769
R7101 VDD.n2247 VDD.n2246 0.0185769
R7102 VDD.n2274 VDD.n2273 0.0185769
R7103 VDD.n2281 VDD.n2280 0.0185769
R7104 VDD.n2302 VDD.n2301 0.0185769
R7105 VDD.n2326 VDD.n2325 0.0185769
R7106 VDD.n2336 VDD.n2335 0.0185769
R7107 VDD.n2357 VDD.n2355 0.0185769
R7108 VDD.n2378 VDD.n1591 0.0185769
R7109 VDD.n2400 VDD.n1577 0.0185769
R7110 VDD.n2420 VDD.n1566 0.0185769
R7111 VDD.n2439 VDD.n1544 0.0185769
R7112 VDD.n2441 VDD.n1529 0.0185769
R7113 VDD.n2473 VDD.n2472 0.0185769
R7114 VDD.n2500 VDD.n2499 0.0185769
R7115 VDD.n2507 VDD.n2506 0.0185769
R7116 VDD.n2528 VDD.n2527 0.0185769
R7117 VDD.n2552 VDD.n2551 0.0185769
R7118 VDD.n2562 VDD.n2561 0.0185769
R7119 VDD.n2583 VDD.n2581 0.0185769
R7120 VDD.n2604 VDD.n1457 0.0185769
R7121 VDD.n2626 VDD.n1443 0.0185769
R7122 VDD.n2646 VDD.n1432 0.0185769
R7123 VDD.n2665 VDD.n1410 0.0185769
R7124 VDD.n2667 VDD.n1395 0.0185769
R7125 VDD.n2699 VDD.n2698 0.0185769
R7126 VDD.n2726 VDD.n2725 0.0185769
R7127 VDD.n2733 VDD.n2732 0.0185769
R7128 VDD.n2758 VDD.n2753 0.0185769
R7129 VDD.n2774 VDD.n1349 0.0185769
R7130 VDD.n2886 VDD.n1287 0.0185349
R7131 VDD.n1881 VDD.n1880 0.0184706
R7132 VDD.n1901 VDD.n1900 0.0184706
R7133 VDD.n1922 VDD.n1860 0.0184706
R7134 VDD.n1930 VDD.n1929 0.0184706
R7135 VDD.n1952 VDD.n1951 0.0184706
R7136 VDD.n1972 VDD.n1971 0.0184706
R7137 VDD.n2010 VDD.n1798 0.0184706
R7138 VDD.n2022 VDD.n1796 0.0184706
R7139 VDD.n2046 VDD.n1782 0.0184706
R7140 VDD.n2057 VDD.n1780 0.0184706
R7141 VDD.n2078 VDD.n1763 0.0184706
R7142 VDD.n2102 VDD.n1750 0.0184706
R7143 VDD.n2107 VDD.n2106 0.0184706
R7144 VDD.n2127 VDD.n2126 0.0184706
R7145 VDD.n2148 VDD.n1726 0.0184706
R7146 VDD.n2156 VDD.n2155 0.0184706
R7147 VDD.n2178 VDD.n2177 0.0184706
R7148 VDD.n2198 VDD.n2197 0.0184706
R7149 VDD.n2236 VDD.n1664 0.0184706
R7150 VDD.n2248 VDD.n1662 0.0184706
R7151 VDD.n2272 VDD.n1648 0.0184706
R7152 VDD.n2283 VDD.n1646 0.0184706
R7153 VDD.n2304 VDD.n1629 0.0184706
R7154 VDD.n2328 VDD.n1616 0.0184706
R7155 VDD.n2333 VDD.n2332 0.0184706
R7156 VDD.n2353 VDD.n2352 0.0184706
R7157 VDD.n2374 VDD.n1592 0.0184706
R7158 VDD.n2382 VDD.n2381 0.0184706
R7159 VDD.n2404 VDD.n2403 0.0184706
R7160 VDD.n2424 VDD.n2423 0.0184706
R7161 VDD.n2462 VDD.n1530 0.0184706
R7162 VDD.n2474 VDD.n1528 0.0184706
R7163 VDD.n2498 VDD.n1514 0.0184706
R7164 VDD.n2509 VDD.n1512 0.0184706
R7165 VDD.n2530 VDD.n1495 0.0184706
R7166 VDD.n2554 VDD.n1482 0.0184706
R7167 VDD.n2559 VDD.n2558 0.0184706
R7168 VDD.n2579 VDD.n2578 0.0184706
R7169 VDD.n2600 VDD.n1458 0.0184706
R7170 VDD.n2608 VDD.n2607 0.0184706
R7171 VDD.n2630 VDD.n2629 0.0184706
R7172 VDD.n2650 VDD.n2649 0.0184706
R7173 VDD.n2688 VDD.n1396 0.0184706
R7174 VDD.n2700 VDD.n1394 0.0184706
R7175 VDD.n2724 VDD.n1380 0.0184706
R7176 VDD.n2735 VDD.n1378 0.0184706
R7177 VDD.n2760 VDD.n1360 0.0184706
R7178 VDD.n2773 VDD.n1350 0.0184706
R7179 VDD.n2788 VDD.n1348 0.0184706
R7180 VDD.n2807 VDD.n1337 0.0184706
R7181 VDD.n2826 VDD.n1326 0.0184706
R7182 VDD.n2845 VDD.n1315 0.0184706
R7183 VDD.n2865 VDD.n1303 0.0184706
R7184 VDD.n2881 VDD.n1288 0.0184706
R7185 VDD.n1090 VDD.n1089 0.0184278
R7186 VDD.n472 VDD.n443 0.0180439
R7187 VDD.n1882 VDD.n1879 0.0179744
R7188 VDD.n1902 VDD.n1871 0.0179744
R7189 VDD.n1904 VDD.n1861 0.0179744
R7190 VDD.n1928 VDD.n1927 0.0179744
R7191 VDD.n1950 VDD.n1949 0.0179744
R7192 VDD.n1970 VDD.n1969 0.0179744
R7193 VDD.n1990 VDD.n1988 0.0179744
R7194 VDD.n2015 VDD.n2014 0.0179744
R7195 VDD.n2016 VDD.n1783 0.0179744
R7196 VDD.n2053 VDD.n1781 0.0179744
R7197 VDD.n2074 VDD.n1764 0.0179744
R7198 VDD.n2098 VDD.n1751 0.0179744
R7199 VDD.n2108 VDD.n1747 0.0179744
R7200 VDD.n2128 VDD.n1737 0.0179744
R7201 VDD.n2130 VDD.n1727 0.0179744
R7202 VDD.n2154 VDD.n2153 0.0179744
R7203 VDD.n2176 VDD.n2175 0.0179744
R7204 VDD.n2196 VDD.n2195 0.0179744
R7205 VDD.n2216 VDD.n2214 0.0179744
R7206 VDD.n2241 VDD.n2240 0.0179744
R7207 VDD.n2242 VDD.n1649 0.0179744
R7208 VDD.n2279 VDD.n1647 0.0179744
R7209 VDD.n2300 VDD.n1630 0.0179744
R7210 VDD.n2324 VDD.n1617 0.0179744
R7211 VDD.n2334 VDD.n1613 0.0179744
R7212 VDD.n2354 VDD.n1603 0.0179744
R7213 VDD.n2356 VDD.n1593 0.0179744
R7214 VDD.n2380 VDD.n2379 0.0179744
R7215 VDD.n2402 VDD.n2401 0.0179744
R7216 VDD.n2422 VDD.n2421 0.0179744
R7217 VDD.n2442 VDD.n2440 0.0179744
R7218 VDD.n2467 VDD.n2466 0.0179744
R7219 VDD.n2468 VDD.n1515 0.0179744
R7220 VDD.n2505 VDD.n1513 0.0179744
R7221 VDD.n2526 VDD.n1496 0.0179744
R7222 VDD.n2550 VDD.n1483 0.0179744
R7223 VDD.n2560 VDD.n1479 0.0179744
R7224 VDD.n2580 VDD.n1469 0.0179744
R7225 VDD.n2582 VDD.n1459 0.0179744
R7226 VDD.n2606 VDD.n2605 0.0179744
R7227 VDD.n2628 VDD.n2627 0.0179744
R7228 VDD.n2648 VDD.n2647 0.0179744
R7229 VDD.n2668 VDD.n2666 0.0179744
R7230 VDD.n2693 VDD.n2692 0.0179744
R7231 VDD.n2694 VDD.n1381 0.0179744
R7232 VDD.n2731 VDD.n1379 0.0179744
R7233 VDD.n2752 VDD.n1362 0.0179744
R7234 VDD.n2757 VDD.n2756 0.0179744
R7235 VDD.n2786 VDD.n2785 0.0179074
R7236 VDD.n2805 VDD.n2804 0.0179074
R7237 VDD.n2824 VDD.n2823 0.0179074
R7238 VDD.n2843 VDD.n2842 0.0179074
R7239 VDD.n2863 VDD.n2861 0.0179074
R7240 VDD.n2883 VDD.n2882 0.0179074
R7241 VDD.n876 VDD.n809 0.0178464
R7242 VDD.n547 VDD 0.0177414
R7243 VDD.n890 VDD.n889 0.0175557
R7244 VDD.n854 VDD.n853 0.0174492
R7245 VDD.n2784 VDD.n2775 0.0173272
R7246 VDD.n2803 VDD.n1338 0.0173272
R7247 VDD.n2822 VDD.n1327 0.0173272
R7248 VDD.n2841 VDD.n1316 0.0173272
R7249 VDD.n2860 VDD.n1305 0.0173272
R7250 VDD.n2862 VDD.n1289 0.0173272
R7251 VDD.n2908 VDD.n2899 0.0172857
R7252 VDD.n170 VDD.n169 0.017168
R7253 VDD.n420 VDD.n417 0.017168
R7254 VDD.n2921 VDD.n2920 0.0171448
R7255 VDD.n655 VDD.n654 0.0170441
R7256 VDD.n2887 VDD.n2886 0.0168953
R7257 VDD.n2887 VDD.n1285 0.0168953
R7258 VDD.n1058 VDD.n1057 0.0168934
R7259 VDD.n918 VDD.n798 0.016776
R7260 VDD.n1172 VDD.n934 0.016776
R7261 VDD.n1143 VDD.n1142 0.016776
R7262 VDD.n123 VDD.n53 0.016776
R7263 VDD.n624 VDD.n141 0.016776
R7264 VDD.n1068 VDD.n1067 0.0165866
R7265 VDD.n1112 VDD.n1105 0.0164897
R7266 VDD.n405 VDD.n404 0.0163928
R7267 VDD.n567 VDD.n566 0.0162959
R7268 VDD.n696 VDD.n695 0.016199
R7269 VDD.n2997 VDD.n6 0.016125
R7270 VDD.n1095 VDD.n1094 0.0161021
R7271 VDD.n1026 VDD.n1025 0.0160052
R7272 VDD.n424 VDD.n423 0.0159082
R7273 VDD.n864 VDD.n863 0.0158509
R7274 VDD.n1037 VDD.n1036 0.0158509
R7275 VDD.n2919 VDD.n2917 0.0156071
R7276 VDD.n2959 VDD.n2958 0.0156071
R7277 VDD.n2979 VDD.n1277 0.0156071
R7278 VDD.n2983 VDD.n38 0.0156071
R7279 VDD.n2936 VDD.n2923 0.0156071
R7280 VDD.n2932 VDD.n2923 0.0156071
R7281 VDD.n2946 VDD.n2898 0.0156071
R7282 VDD.n2946 VDD.n2897 0.0156071
R7283 VDD.n2944 VDD.n2911 0.0156071
R7284 VDD.n2944 VDD.n2940 0.0156071
R7285 VDD.n1188 VDD.n1187 0.0153268
R7286 VDD.n299 VDD.n298 0.0153268
R7287 VDD.n2888 VDD.n1286 0.0152558
R7288 VDD.n529 VDD.n528 0.0152299
R7289 VDD.n1104 VDD.n992 0.0150862
R7290 VDD.n1096 VDD.n994 0.0150862
R7291 VDD.n1069 VDD.n997 0.0150862
R7292 VDD.n887 VDD.n886 0.0150862
R7293 VDD.n870 VDD.n869 0.0150862
R7294 VDD.n716 VDD.n713 0.0150862
R7295 VDD.n1273 VDD.n702 0.0150862
R7296 VDD.n891 VDD.n805 0.0150862
R7297 VDD.n1065 VDD.n1064 0.0150862
R7298 VDD.n1186 VDD.n902 0.0150862
R7299 VDD.n1005 VDD.n902 0.0150862
R7300 VDD.n1022 VDD.n938 0.0150862
R7301 VDD.n939 VDD.n938 0.0150862
R7302 VDD.n1111 VDD.n990 0.0150862
R7303 VDD.n1268 VDD.n705 0.0150862
R7304 VDD.n828 VDD.n827 0.0150862
R7305 VDD.n837 VDD.n827 0.0150862
R7306 VDD.n877 VDD.n824 0.0150862
R7307 VDD.n882 VDD.n881 0.0150862
R7308 VDD.n1032 VDD.n1000 0.0150862
R7309 VDD.n898 VDD.n803 0.0150862
R7310 VDD.n1092 VDD.n1091 0.0150862
R7311 VDD.n1190 VDD.n799 0.0150862
R7312 VDD.n1190 VDD.n801 0.0150862
R7313 VDD.n1008 VDD.n1002 0.0150862
R7314 VDD.n1020 VDD.n1002 0.0150862
R7315 VDD.n1263 VDD.n708 0.0150862
R7316 VDD.n1254 VDD.n708 0.0150862
R7317 VDD.n865 VDD.n839 0.0150862
R7318 VDD.n1061 VDD.n1035 0.0150862
R7319 VDD.n694 VDD.n44 0.0150862
R7320 VDD.n699 VDD.n41 0.0150862
R7321 VDD.n422 VDD.n396 0.0150862
R7322 VDD.n435 VDD.n396 0.0150862
R7323 VDD.n438 VDD.n394 0.0150862
R7324 VDD.n476 VDD.n394 0.0150862
R7325 VDD.n532 VDD.n327 0.0150862
R7326 VDD.n565 VDD.n322 0.0150862
R7327 VDD.n279 VDD.n267 0.0150862
R7328 VDD.n300 VDD.n286 0.0150862
R7329 VDD.n296 VDD.n295 0.0150862
R7330 VDD.n184 VDD.n149 0.0150862
R7331 VDD.n677 VDD.n52 0.0150862
R7332 VDD.n189 VDD.n147 0.0150862
R7333 VDD.n618 VDD.n147 0.0150862
R7334 VDD.n615 VDD.n193 0.0150862
R7335 VDD.n220 VDD.n193 0.0150862
R7336 VDD.n227 VDD.n219 0.0150862
R7337 VDD.n598 VDD.n219 0.0150862
R7338 VDD.n595 VDD.n231 0.0150862
R7339 VDD.n292 VDD.n231 0.0150862
R7340 VDD.n473 VDD.n442 0.0150862
R7341 VDD.n672 VDD.n55 0.0150862
R7342 VDD.n640 VDD.n60 0.0150862
R7343 VDD.n168 VDD.n60 0.0150862
R7344 VDD.n406 VDD.n402 0.0150862
R7345 VDD.n416 VDD.n402 0.0150862
R7346 VDD.n419 VDD.n400 0.0150862
R7347 VDD.n425 VDD.n400 0.0150862
R7348 VDD.n332 VDD.n330 0.0150862
R7349 VDD.n689 VDD.n47 0.0150862
R7350 VDD.n680 VDD.n47 0.0150862
R7351 VDD.n666 VDD.n57 0.0150862
R7352 VDD.n309 VDD.n281 0.0150862
R7353 VDD.n318 VDD.n281 0.0150862
R7354 VDD.n559 VDD.n324 0.0150862
R7355 VDD.n2906 VDD.n2903 0.0148621
R7356 VDD.n674 VDD.n673 0.0146485
R7357 VDD.n874 VDD.n872 0.0143577
R7358 VDD.n1885 VDD.n1872 0.0143235
R7359 VDD.n1906 VDD.n1870 0.0143235
R7360 VDD.n1925 VDD.n1858 0.0143235
R7361 VDD.n1947 VDD.n1844 0.0143235
R7362 VDD.n1967 VDD.n1833 0.0143235
R7363 VDD.n2013 VDD.n2011 0.0143235
R7364 VDD.n2019 VDD.n2018 0.0143235
R7365 VDD.n2050 VDD.n2049 0.0143235
R7366 VDD.n2056 VDD.n1765 0.0143235
R7367 VDD.n2077 VDD.n1752 0.0143235
R7368 VDD.n2111 VDD.n1738 0.0143235
R7369 VDD.n2132 VDD.n1736 0.0143235
R7370 VDD.n2151 VDD.n1724 0.0143235
R7371 VDD.n2173 VDD.n1710 0.0143235
R7372 VDD.n2193 VDD.n1699 0.0143235
R7373 VDD.n2239 VDD.n2237 0.0143235
R7374 VDD.n2245 VDD.n2244 0.0143235
R7375 VDD.n2276 VDD.n2275 0.0143235
R7376 VDD.n2282 VDD.n1631 0.0143235
R7377 VDD.n2303 VDD.n1618 0.0143235
R7378 VDD.n2337 VDD.n1604 0.0143235
R7379 VDD.n2358 VDD.n1602 0.0143235
R7380 VDD.n2377 VDD.n1590 0.0143235
R7381 VDD.n2399 VDD.n1576 0.0143235
R7382 VDD.n2419 VDD.n1565 0.0143235
R7383 VDD.n2465 VDD.n2463 0.0143235
R7384 VDD.n2471 VDD.n2470 0.0143235
R7385 VDD.n2502 VDD.n2501 0.0143235
R7386 VDD.n2508 VDD.n1497 0.0143235
R7387 VDD.n2529 VDD.n1484 0.0143235
R7388 VDD.n2563 VDD.n1470 0.0143235
R7389 VDD.n2584 VDD.n1468 0.0143235
R7390 VDD.n2603 VDD.n1456 0.0143235
R7391 VDD.n2625 VDD.n1442 0.0143235
R7392 VDD.n2645 VDD.n1431 0.0143235
R7393 VDD.n2691 VDD.n2689 0.0143235
R7394 VDD.n2697 VDD.n2696 0.0143235
R7395 VDD.n2728 VDD.n2727 0.0143235
R7396 VDD.n2734 VDD.n1363 0.0143235
R7397 VDD.n2759 VDD.n1361 0.0143235
R7398 VDD.n2787 VDD.n1339 0.0143235
R7399 VDD.n2806 VDD.n1328 0.0143235
R7400 VDD.n2825 VDD.n1317 0.0143235
R7401 VDD.n2844 VDD.n1306 0.0143235
R7402 VDD.n2864 VDD.n1304 0.0143235
R7403 VDD.n597 VDD.n596 0.0142608
R7404 VDD.n228 VDD.n221 0.0141639
R7405 VDD.n3009 VDD.n9 0.0140135
R7406 VDD.n277 VDD.n276 0.0140001
R7407 VDD.n439 VDD.n436 0.0137763
R7408 VDD.n1899 VDD.n1898 0.0137576
R7409 VDD.n1920 VDD.n1919 0.0137576
R7410 VDD.n1931 VDD.n1857 0.0137576
R7411 VDD.n1953 VDD.n1843 0.0137576
R7412 VDD.n1973 VDD.n1832 0.0137576
R7413 VDD.n2009 VDD.n1799 0.0137576
R7414 VDD.n2024 VDD.n1792 0.0137576
R7415 VDD.n2044 VDD.n1786 0.0137576
R7416 VDD.n2059 VDD.n2058 0.0137576
R7417 VDD.n2079 VDD.n1762 0.0137576
R7418 VDD.n2103 VDD.n1749 0.0137576
R7419 VDD.n2105 VDD.n2104 0.0137576
R7420 VDD.n2125 VDD.n2124 0.0137576
R7421 VDD.n2146 VDD.n2145 0.0137576
R7422 VDD.n2157 VDD.n1723 0.0137576
R7423 VDD.n2179 VDD.n1709 0.0137576
R7424 VDD.n2199 VDD.n1698 0.0137576
R7425 VDD.n2235 VDD.n1665 0.0137576
R7426 VDD.n2250 VDD.n1658 0.0137576
R7427 VDD.n2270 VDD.n1652 0.0137576
R7428 VDD.n2285 VDD.n2284 0.0137576
R7429 VDD.n2305 VDD.n1628 0.0137576
R7430 VDD.n2329 VDD.n1615 0.0137576
R7431 VDD.n2331 VDD.n2330 0.0137576
R7432 VDD.n2351 VDD.n2350 0.0137576
R7433 VDD.n2372 VDD.n2371 0.0137576
R7434 VDD.n2383 VDD.n1589 0.0137576
R7435 VDD.n2405 VDD.n1575 0.0137576
R7436 VDD.n2425 VDD.n1564 0.0137576
R7437 VDD.n2461 VDD.n1531 0.0137576
R7438 VDD.n2476 VDD.n1524 0.0137576
R7439 VDD.n2496 VDD.n1518 0.0137576
R7440 VDD.n2511 VDD.n2510 0.0137576
R7441 VDD.n2531 VDD.n1494 0.0137576
R7442 VDD.n2555 VDD.n1481 0.0137576
R7443 VDD.n2557 VDD.n2556 0.0137576
R7444 VDD.n2577 VDD.n2576 0.0137576
R7445 VDD.n2598 VDD.n2597 0.0137576
R7446 VDD.n2609 VDD.n1455 0.0137576
R7447 VDD.n2631 VDD.n1441 0.0137576
R7448 VDD.n2651 VDD.n1430 0.0137576
R7449 VDD.n2687 VDD.n1397 0.0137576
R7450 VDD.n2702 VDD.n1390 0.0137576
R7451 VDD.n2722 VDD.n1384 0.0137576
R7452 VDD.n2737 VDD.n2736 0.0137576
R7453 VDD.n2761 VDD.n1359 0.0137576
R7454 VDD.n2789 VDD.n1347 0.0137576
R7455 VDD.n2808 VDD.n1336 0.0137576
R7456 VDD.n2827 VDD.n1325 0.0137576
R7457 VDD.n2846 VDD.n1314 0.0137576
R7458 VDD.n2866 VDD.n1302 0.0137576
R7459 VDD.n2879 VDD.n2878 0.0137576
R7460 VDD.n2905 VDD.n2901 0.0137243
R7461 VDD.n3008 VDD.n11 0.0137188
R7462 VDD.n3008 VDD.n13 0.0137188
R7463 VDD.n433 VDD.n397 0.0136579
R7464 VDD.n432 VDD.n388 0.0135208
R7465 VDD.n665 VDD.n642 0.013404
R7466 VDD.n190 VDD.n187 0.0132918
R7467 VDD.n31 VDD.t129 0.0132807
R7468 VDD.n1252 VDD.n712 0.0131948
R7469 VDD.n3004 VDD.n3003 0.0130393
R7470 VDD.n17 VDD.n14 0.0130393
R7471 VDD.n1239 VDD.n1238 0.0128698
R7472 VDD.n225 VDD.n216 0.0128698
R7473 VDD.n601 VDD.n600 0.0128698
R7474 VDD.n510 VDD.n333 0.0128698
R7475 VDD.n1039 VDD.n1036 0.0127516
R7476 VDD.n864 VDD.n841 0.0127493
R7477 VDD.n1270 VDD.n1269 0.0127103
R7478 VDD.n868 VDD.n838 0.0126134
R7479 VDD.n183 VDD.n182 0.0126134
R7480 VDD.n2918 VDD.n1280 0.0126104
R7481 VDD.n1884 VDD.n1871 0.0125513
R7482 VDD.n1905 VDD.n1904 0.0125513
R7483 VDD.n1927 VDD.n1926 0.0125513
R7484 VDD.n1949 VDD.n1948 0.0125513
R7485 VDD.n1969 VDD.n1968 0.0125513
R7486 VDD.n2014 VDD.n1797 0.0125513
R7487 VDD.n2020 VDD.n2016 0.0125513
R7488 VDD.n2048 VDD.n1781 0.0125513
R7489 VDD.n2055 VDD.n1764 0.0125513
R7490 VDD.n2076 VDD.n1751 0.0125513
R7491 VDD.n2110 VDD.n1737 0.0125513
R7492 VDD.n2131 VDD.n2130 0.0125513
R7493 VDD.n2153 VDD.n2152 0.0125513
R7494 VDD.n2175 VDD.n2174 0.0125513
R7495 VDD.n2195 VDD.n2194 0.0125513
R7496 VDD.n2240 VDD.n1663 0.0125513
R7497 VDD.n2246 VDD.n2242 0.0125513
R7498 VDD.n2274 VDD.n1647 0.0125513
R7499 VDD.n2281 VDD.n1630 0.0125513
R7500 VDD.n2302 VDD.n1617 0.0125513
R7501 VDD.n2336 VDD.n1603 0.0125513
R7502 VDD.n2357 VDD.n2356 0.0125513
R7503 VDD.n2379 VDD.n2378 0.0125513
R7504 VDD.n2401 VDD.n2400 0.0125513
R7505 VDD.n2421 VDD.n2420 0.0125513
R7506 VDD.n2466 VDD.n1529 0.0125513
R7507 VDD.n2472 VDD.n2468 0.0125513
R7508 VDD.n2500 VDD.n1513 0.0125513
R7509 VDD.n2507 VDD.n1496 0.0125513
R7510 VDD.n2528 VDD.n1483 0.0125513
R7511 VDD.n2562 VDD.n1469 0.0125513
R7512 VDD.n2583 VDD.n2582 0.0125513
R7513 VDD.n2605 VDD.n2604 0.0125513
R7514 VDD.n2627 VDD.n2626 0.0125513
R7515 VDD.n2647 VDD.n2646 0.0125513
R7516 VDD.n2692 VDD.n1395 0.0125513
R7517 VDD.n2698 VDD.n2694 0.0125513
R7518 VDD.n2726 VDD.n1379 0.0125513
R7519 VDD.n2733 VDD.n1362 0.0125513
R7520 VDD.n2758 VDD.n2757 0.0125513
R7521 VDD.n885 VDD.n884 0.0125165
R7522 VDD.n118 VDD.n87 0.0123994
R7523 VDD.n508 VDD.n331 0.0123859
R7524 VDD.n526 VDD.n331 0.0123641
R7525 VDD.n179 VDD.n178 0.0122188
R7526 VDD.n470 VDD.n469 0.0122188
R7527 VDD.n2786 VDD.n1338 0.0121049
R7528 VDD.n2805 VDD.n1327 0.0121049
R7529 VDD.n2824 VDD.n1316 0.0121049
R7530 VDD.n2843 VDD.n1305 0.0121049
R7531 VDD.n2863 VDD.n2862 0.0121049
R7532 VDD.n617 VDD.n616 0.012032
R7533 VDD.n2981 VDD.n2980 0.0118253
R7534 VDD.n475 VDD.n474 0.0116443
R7535 VDD.n1173 VDD.n1172 0.0115677
R7536 VDD.n571 VDD.n570 0.0115677
R7537 VDD.n398 VDD.n380 0.0115677
R7538 VDD.n662 VDD.n655 0.0115294
R7539 VDD.n222 VDD.n217 0.0114649
R7540 VDD.n665 VDD.n664 0.0114649
R7541 VDD.n1007 VDD.n1006 0.0114505
R7542 VDD.n308 VDD.n306 0.0114505
R7543 VDD.n1197 VDD 0.0109167
R7544 VDD.n919 VDD.n918 0.0109167
R7545 VDD.n931 VDD.n905 0.0109167
R7546 VDD.n1115 VDD.n988 0.0109167
R7547 VDD.n1117 VDD 0.0109167
R7548 VDD.n612 VDD.n611 0.0109167
R7549 VDD.n288 VDD 0.0109167
R7550 VDD.n414 VDD.n409 0.0109167
R7551 VDD.n457 VDD 0.0109167
R7552 VDD.n1058 VDD.n1047 0.0107459
R7553 VDD.n2907 VDD.n2902 0.0105714
R7554 VDD.n311 VDD.n310 0.0105041
R7555 VDD.n1265 VDD.n1264 0.0104814
R7556 VDD.n2916 VDD.n2915 0.0103794
R7557 VDD.n2957 VDD.n1281 0.0103794
R7558 VDD.n2934 VDD.n2933 0.0103794
R7559 VDD.n2948 VDD.n2947 0.0103794
R7560 VDD.n2943 VDD.n2942 0.0103794
R7561 VDD.n1184 VDD.n1183 0.0102656
R7562 VDD.n1108 VDD.n976 0.0102656
R7563 VDD.n238 VDD.n233 0.0102656
R7564 VDD.n290 VDD.n234 0.0102656
R7565 VDD.n862 VDD.n861 0.0101138
R7566 VDD.n2792 VDD.n2791 0.0099697
R7567 VDD.n2811 VDD.n2810 0.0099697
R7568 VDD.n2830 VDD.n2829 0.0099697
R7569 VDD.n2849 VDD.n2848 0.0099697
R7570 VDD.n2869 VDD.n2868 0.0099697
R7571 VDD.n1896 VDD.n1895 0.0099697
R7572 VDD.n1917 VDD.n1916 0.0099697
R7573 VDD.n1932 VDD.n1856 0.0099697
R7574 VDD.n1956 VDD.n1955 0.0099697
R7575 VDD.n1976 VDD.n1975 0.0099697
R7576 VDD.n1825 VDD.n1824 0.0099697
R7577 VDD.n1821 VDD.n1820 0.0099697
R7578 VDD.n2007 VDD.n2006 0.0099697
R7579 VDD.n2026 VDD.n1791 0.0099697
R7580 VDD.n2042 VDD.n2039 0.0099697
R7581 VDD.n1777 VDD.n1776 0.0099697
R7582 VDD.n2082 VDD.n2081 0.0099697
R7583 VDD.n2122 VDD.n2121 0.0099697
R7584 VDD.n2143 VDD.n2142 0.0099697
R7585 VDD.n2158 VDD.n1722 0.0099697
R7586 VDD.n2182 VDD.n2181 0.0099697
R7587 VDD.n2202 VDD.n2201 0.0099697
R7588 VDD.n1691 VDD.n1690 0.0099697
R7589 VDD.n1687 VDD.n1686 0.0099697
R7590 VDD.n2233 VDD.n2232 0.0099697
R7591 VDD.n2252 VDD.n1657 0.0099697
R7592 VDD.n2268 VDD.n2265 0.0099697
R7593 VDD.n1643 VDD.n1642 0.0099697
R7594 VDD.n2308 VDD.n2307 0.0099697
R7595 VDD.n2348 VDD.n2347 0.0099697
R7596 VDD.n2369 VDD.n2368 0.0099697
R7597 VDD.n2384 VDD.n1588 0.0099697
R7598 VDD.n2408 VDD.n2407 0.0099697
R7599 VDD.n2428 VDD.n2427 0.0099697
R7600 VDD.n1557 VDD.n1556 0.0099697
R7601 VDD.n1553 VDD.n1552 0.0099697
R7602 VDD.n2459 VDD.n2458 0.0099697
R7603 VDD.n2478 VDD.n1523 0.0099697
R7604 VDD.n2494 VDD.n2491 0.0099697
R7605 VDD.n1509 VDD.n1508 0.0099697
R7606 VDD.n2534 VDD.n2533 0.0099697
R7607 VDD.n2574 VDD.n2573 0.0099697
R7608 VDD.n2595 VDD.n2594 0.0099697
R7609 VDD.n2610 VDD.n1454 0.0099697
R7610 VDD.n2634 VDD.n2633 0.0099697
R7611 VDD.n2654 VDD.n2653 0.0099697
R7612 VDD.n1423 VDD.n1422 0.0099697
R7613 VDD.n1419 VDD.n1418 0.0099697
R7614 VDD.n2685 VDD.n2684 0.0099697
R7615 VDD.n2704 VDD.n1389 0.0099697
R7616 VDD.n2720 VDD.n2717 0.0099697
R7617 VDD.n1375 VDD.n1374 0.0099697
R7618 VDD.n2765 VDD.n2764 0.0099697
R7619 VDD.n1030 VDD.n1029 0.00961458
R7620 VDD.n1155 VDD.n1154 0.00961458
R7621 VDD.n478 VDD.n391 0.00961458
R7622 VDD.n562 VDD.n561 0.00951237
R7623 VDD.n556 VDD.n555 0.00944537
R7624 VDD.n310 VDD.n282 0.00927193
R7625 VDD.n862 VDD.n843 0.00897458
R7626 VDD.n834 VDD.n833 0.00896354
R7627 VDD.n834 VDD.n753 0.00896354
R7628 VDD.n638 VDD.n63 0.00896354
R7629 VDD.n66 VDD.n63 0.00896354
R7630 VDD.n144 VDD.n142 0.00896354
R7631 VDD.n620 VDD.n144 0.00896354
R7632 VDD.n200 VDD.n145 0.00896354
R7633 VDD.n451 VDD.n392 0.00896354
R7634 VDD.n667 VDD.n641 0.00883402
R7635 VDD.n853 VDD 0.00865217
R7636 VDD.n1057 VDD 0.00865217
R7637 VDD.n1063 VDD.n1062 0.00864021
R7638 VDD.n832 VDD.n719 0.0083125
R7639 VDD.n119 VDD.n118 0.0083125
R7640 VDD.n74 VDD.n62 0.0083125
R7641 VDD.n391 VDD.n389 0.0083125
R7642 VDD.n527 VDD.n330 0.00827754
R7643 VDD.n171 VDD.n151 0.00827754
R7644 VDD.n1011 VDD.n1004 0.00771154
R7645 VDD.n1249 VDD.n718 0.00766146
R7646 VDD.n1183 VDD.n1182 0.00766146
R7647 VDD.n223 VDD.n196 0.00766146
R7648 VDD.n593 VDD.n234 0.00766146
R7649 VDD.n371 VDD.n333 0.00766146
R7650 VDD.n410 VDD.n379 0.00766146
R7651 VDD.n484 VDD.n388 0.00766146
R7652 VDD.n687 VDD.n49 0.00761015
R7653 VDD.n1010 VDD.n1003 0.00707895
R7654 VDD.n1109 VDD.n988 0.00701042
R7655 VDD.n613 VDD.n612 0.00701042
R7656 VDD.n409 VDD.n408 0.00701042
R7657 VDD.n2997 VDD.n27 0.00701042
R7658 VDD.n3011 VDD.n6 0.00701042
R7659 VDD.n560 VDD.n533 0.00699278
R7660 VDD.n1012 VDD.n1011 0.00693001
R7661 VDD.n1034 VDD.n1033 0.00689588
R7662 VDD.n853 VDD 0.00685593
R7663 VDD.n1057 VDD 0.00664754
R7664 VDD.n177 VDD.n172 0.00635938
R7665 VDD.n303 VDD.n302 0.00635938
R7666 VDD.n496 VDD.n380 0.00635938
R7667 VDD.n427 VDD.n398 0.00635938
R7668 VDD.n469 VDD.n445 0.00635938
R7669 VDD.n2919 VDD.n2913 0.00635126
R7670 VDD.n2959 VDD.n1279 0.00635126
R7671 VDD.n181 VDD.n151 0.00619964
R7672 VDD.n691 VDD.n690 0.00612062
R7673 VDD.n669 VDD.n668 0.00602371
R7674 VDD.n179 VDD.n67 0.00570833
R7675 VDD.n178 VDD.n177 0.00570833
R7676 VDD.n497 VDD.n496 0.00570833
R7677 VDD.n471 VDD.n470 0.00570833
R7678 VDD.n456 VDD.n445 0.00570833
R7679 VDD.n682 VDD.n49 0.00530769
R7680 VDD.n1088 VDD.n997 0.00527274
R7681 VDD.n568 VDD.n279 0.00526787
R7682 VDD.n1061 VDD.n1060 0.00523977
R7683 VDD.n666 VDD.n58 0.0052393
R7684 VDD.n1171 VDD.n937 0.00512963
R7685 VDD.n510 VDD.n509 0.00505729
R7686 VDD.n25 VDD.n24 0.00490305
R7687 VDD.n558 VDD.n557 0.00488596
R7688 VDD.n2960 VDD.n1278 0.00482515
R7689 VDD.n1280 VDD.n1278 0.00482515
R7690 VDD.n2918 VDD.n2912 0.00482515
R7691 VDD.n2920 VDD.n2912 0.00482515
R7692 VDD.n549 VDD.n535 0.00481034
R7693 VDD.n556 VDD.n535 0.00481034
R7694 VDD VDD.n546 0.00481034
R7695 VDD.n2928 VDD.n2926 0.00476089
R7696 VDD.n865 VDD.n840 0.00461828
R7697 VDD.n559 VDD.n325 0.00461763
R7698 VDD.n611 VDD.n196 0.00440625
R7699 VDD.n371 VDD.n370 0.00440625
R7700 VDD.n414 VDD.n410 0.00440625
R7701 VDD.n432 VDD.n431 0.00440625
R7702 VDD.n484 VDD.n483 0.00440625
R7703 VDD.n3011 VDD.n3010 0.00440625
R7704 VDD.n1887 VDD.n1877 0.00428788
R7705 VDD.n1908 VDD.n1868 0.00428788
R7706 VDD.n1921 VDD.n1854 0.00428788
R7707 VDD.n1945 VDD.n1847 0.00428788
R7708 VDD.n1965 VDD.n1836 0.00428788
R7709 VDD.n1984 VDD.n1814 0.00428788
R7710 VDD.n1993 VDD.n1810 0.00428788
R7711 VDD.n2023 VDD.n1794 0.00428788
R7712 VDD.n2045 VDD.n1785 0.00428788
R7713 VDD.n1778 VDD.n1774 0.00428788
R7714 VDD.n2071 VDD.n1767 0.00428788
R7715 VDD.n2095 VDD.n1754 0.00428788
R7716 VDD.n2113 VDD.n1745 0.00428788
R7717 VDD.n2134 VDD.n1734 0.00428788
R7718 VDD.n2147 VDD.n1720 0.00428788
R7719 VDD.n2171 VDD.n1713 0.00428788
R7720 VDD.n2191 VDD.n1702 0.00428788
R7721 VDD.n2210 VDD.n1680 0.00428788
R7722 VDD.n2219 VDD.n1676 0.00428788
R7723 VDD.n2249 VDD.n1660 0.00428788
R7724 VDD.n2271 VDD.n1651 0.00428788
R7725 VDD.n1644 VDD.n1640 0.00428788
R7726 VDD.n2297 VDD.n1633 0.00428788
R7727 VDD.n2321 VDD.n1620 0.00428788
R7728 VDD.n2339 VDD.n1611 0.00428788
R7729 VDD.n2360 VDD.n1600 0.00428788
R7730 VDD.n2373 VDD.n1586 0.00428788
R7731 VDD.n2397 VDD.n1579 0.00428788
R7732 VDD.n2417 VDD.n1568 0.00428788
R7733 VDD.n2436 VDD.n1546 0.00428788
R7734 VDD.n2445 VDD.n1542 0.00428788
R7735 VDD.n2475 VDD.n1526 0.00428788
R7736 VDD.n2497 VDD.n1517 0.00428788
R7737 VDD.n1510 VDD.n1506 0.00428788
R7738 VDD.n2523 VDD.n1499 0.00428788
R7739 VDD.n2547 VDD.n1486 0.00428788
R7740 VDD.n2565 VDD.n1477 0.00428788
R7741 VDD.n2586 VDD.n1466 0.00428788
R7742 VDD.n2599 VDD.n1452 0.00428788
R7743 VDD.n2623 VDD.n1445 0.00428788
R7744 VDD.n2643 VDD.n1434 0.00428788
R7745 VDD.n2662 VDD.n1412 0.00428788
R7746 VDD.n2671 VDD.n1408 0.00428788
R7747 VDD.n2701 VDD.n1392 0.00428788
R7748 VDD.n2723 VDD.n1383 0.00428788
R7749 VDD.n1376 VDD.n1372 0.00428788
R7750 VDD.n2749 VDD.n1365 0.00428788
R7751 VDD.n1353 VDD.n1351 0.00428788
R7752 VDD.n2781 VDD.n2780 0.00428788
R7753 VDD.n2800 VDD.n1341 0.00428788
R7754 VDD.n2819 VDD.n1330 0.00428788
R7755 VDD.n2838 VDD.n1319 0.00428788
R7756 VDD.n2857 VDD.n1308 0.00428788
R7757 VDD.n2880 VDD.n2877 0.00428788
R7758 VDD.n21 VDD.n20 0.00428087
R7759 VDD.n2964 VDD.n1277 0.00397409
R7760 VDD.n2984 VDD.n2983 0.00397409
R7761 VDD.n2929 VDD.n2928 0.00397409
R7762 VDD.n679 VDD.n46 0.00395565
R7763 VDD.n2889 VDD.n2888 0.00391036
R7764 VDD.n1113 VDD.n990 0.00390422
R7765 VDD.n442 VDD.n441 0.00390422
R7766 VDD.n873 VDD.n824 0.00387702
R7767 VDD.n883 VDD.n882 0.00387702
R7768 VDD.n1102 VDD.n992 0.00386759
R7769 VDD.n1099 VDD.n994 0.00386759
R7770 VDD.n888 VDD.n887 0.00386759
R7771 VDD.n871 VDD.n870 0.00386759
R7772 VDD.n1271 VDD.n702 0.00386759
R7773 VDD.n893 VDD.n805 0.00386759
R7774 VDD.n1066 VDD.n1065 0.00386759
R7775 VDD.n1266 VDD.n705 0.00386759
R7776 VDD.n1027 VDD.n1000 0.00386759
R7777 VDD.n896 VDD.n803 0.00386759
R7778 VDD.n1093 VDD.n1092 0.00386759
R7779 VDD.n692 VDD.n44 0.00386759
R7780 VDD.n697 VDD.n41 0.00386759
R7781 VDD.n530 VDD.n327 0.00386759
R7782 VDD.n563 VDD.n322 0.00386759
R7783 VDD.n305 VDD.n286 0.00386759
R7784 VDD.n297 VDD.n296 0.00386759
R7785 VDD.n186 VDD.n149 0.00386759
R7786 VDD.n675 VDD.n52 0.00386759
R7787 VDD.n670 VDD.n55 0.00386759
R7788 VDD.n1251 VDD.n713 0.00386598
R7789 VDD.n690 VDD.n46 0.00385878
R7790 VDD.n308 VDD.n307 0.00385877
R7791 VDD.n1285 VDD 0.00377907
R7792 VDD.n711 VDD.n710 0.00376184
R7793 VDD.n833 VDD.n832 0.00375521
R7794 VDD.n99 VDD.n42 0.00375521
R7795 VDD.n120 VDD.n119 0.00375521
R7796 VDD.n638 VDD.n62 0.00375521
R7797 VDD.n601 VDD.n216 0.00375521
R7798 VDD.n1040 VDD.n1038 0.0036585
R7799 VDD.n3003 VDD.n24 0.00360776
R7800 VDD.n21 VDD.n14 0.00360776
R7801 VDD.n2907 VDD.n2900 0.00351641
R7802 VDD.n1274 VDD.n701 0.00340722
R7803 VDD.n1270 VDD.n701 0.00340722
R7804 VDD.n1269 VDD.n704 0.00340722
R7805 VDD.n1265 VDD.n704 0.00340722
R7806 VDD.n826 VDD.n712 0.00340722
R7807 VDD.n838 VDD.n826 0.00340722
R7808 VDD.n872 VDD.n825 0.00340722
R7809 VDD.n875 VDD.n874 0.00340722
R7810 VDD.n876 VDD.n875 0.00340722
R7811 VDD.n809 VDD.n807 0.00340722
R7812 VDD.n884 VDD.n807 0.00340722
R7813 VDD.n885 VDD.n806 0.00340722
R7814 VDD.n889 VDD.n806 0.00340722
R7815 VDD.n890 VDD.n804 0.00340722
R7816 VDD.n894 VDD.n804 0.00340722
R7817 VDD.n895 VDD.n802 0.00340722
R7818 VDD.n899 VDD.n802 0.00340722
R7819 VDD.n1189 VDD.n900 0.00340722
R7820 VDD.n1189 VDD.n1188 0.00340722
R7821 VDD.n1187 VDD.n901 0.00340722
R7822 VDD.n1006 VDD.n901 0.00340722
R7823 VDD.n1007 VDD.n1001 0.00340722
R7824 VDD.n1021 VDD.n1001 0.00340722
R7825 VDD.n1024 VDD.n1023 0.00340722
R7826 VDD.n1025 VDD.n1024 0.00340722
R7827 VDD.n1026 VDD.n999 0.00340722
R7828 VDD.n1033 VDD.n999 0.00340722
R7829 VDD.n1063 VDD.n998 0.00340722
R7830 VDD.n1067 VDD.n998 0.00340722
R7831 VDD.n1068 VDD.n996 0.00340722
R7832 VDD.n1089 VDD.n996 0.00340722
R7833 VDD.n1090 VDD.n995 0.00340722
R7834 VDD.n1094 VDD.n995 0.00340722
R7835 VDD.n1095 VDD.n993 0.00340722
R7836 VDD.n1100 VDD.n993 0.00340722
R7837 VDD.n1101 VDD.n991 0.00340722
R7838 VDD.n1105 VDD.n991 0.00340722
R7839 VDD.n700 VDD.n40 0.00340722
R7840 VDD.n696 VDD.n40 0.00340722
R7841 VDD.n695 VDD.n43 0.00340722
R7842 VDD.n691 VDD.n43 0.00340722
R7843 VDD.n679 VDD.n678 0.00340722
R7844 VDD.n678 VDD.n51 0.00340722
R7845 VDD.n674 VDD.n51 0.00340722
R7846 VDD.n673 VDD.n54 0.00340722
R7847 VDD.n669 VDD.n54 0.00340722
R7848 VDD.n641 VDD.n59 0.00340722
R7849 VDD.n169 VDD.n59 0.00340722
R7850 VDD.n170 VDD.n150 0.00340722
R7851 VDD.n182 VDD.n150 0.00340722
R7852 VDD.n183 VDD.n148 0.00340722
R7853 VDD.n187 VDD.n148 0.00340722
R7854 VDD.n191 VDD.n190 0.00340722
R7855 VDD.n617 VDD.n191 0.00340722
R7856 VDD.n616 VDD.n192 0.00340722
R7857 VDD.n221 VDD.n192 0.00340722
R7858 VDD.n229 VDD.n228 0.00340722
R7859 VDD.n597 VDD.n229 0.00340722
R7860 VDD.n596 VDD.n230 0.00340722
R7861 VDD.n293 VDD.n230 0.00340722
R7862 VDD.n294 VDD.n287 0.00340722
R7863 VDD.n298 VDD.n287 0.00340722
R7864 VDD.n299 VDD.n285 0.00340722
R7865 VDD.n306 VDD.n285 0.00340722
R7866 VDD.n567 VDD.n320 0.00340722
R7867 VDD.n566 VDD.n321 0.00340722
R7868 VDD.n562 VDD.n321 0.00340722
R7869 VDD.n533 VDD.n326 0.00340722
R7870 VDD.n529 VDD.n326 0.00340722
R7871 VDD.n528 VDD.n329 0.00340722
R7872 VDD.n404 VDD.n329 0.00340722
R7873 VDD.n405 VDD.n401 0.00340722
R7874 VDD.n417 VDD.n401 0.00340722
R7875 VDD.n421 VDD.n420 0.00340722
R7876 VDD.n424 VDD.n421 0.00340722
R7877 VDD.n423 VDD.n395 0.00340722
R7878 VDD.n436 VDD.n395 0.00340722
R7879 VDD.n440 VDD.n439 0.00340722
R7880 VDD.n475 VDD.n440 0.00340722
R7881 VDD.n526 VDD.n525 0.00334133
R7882 VDD.n2011 VDD.n2010 0.00326471
R7883 VDD.n2019 VDD.n1796 0.00326471
R7884 VDD.n2049 VDD.n1782 0.00326471
R7885 VDD.n2057 VDD.n2056 0.00326471
R7886 VDD.n2078 VDD.n2077 0.00326471
R7887 VDD.n2102 VDD.n2101 0.00326471
R7888 VDD.n2237 VDD.n2236 0.00326471
R7889 VDD.n2245 VDD.n1662 0.00326471
R7890 VDD.n2275 VDD.n1648 0.00326471
R7891 VDD.n2283 VDD.n2282 0.00326471
R7892 VDD.n2304 VDD.n2303 0.00326471
R7893 VDD.n2328 VDD.n2327 0.00326471
R7894 VDD.n2463 VDD.n2462 0.00326471
R7895 VDD.n2471 VDD.n1528 0.00326471
R7896 VDD.n2501 VDD.n1514 0.00326471
R7897 VDD.n2509 VDD.n2508 0.00326471
R7898 VDD.n2530 VDD.n2529 0.00326471
R7899 VDD.n2554 VDD.n2553 0.00326471
R7900 VDD.n2689 VDD.n2688 0.00326471
R7901 VDD.n2697 VDD.n1394 0.00326471
R7902 VDD.n2727 VDD.n1380 0.00326471
R7903 VDD.n2735 VDD.n2734 0.00326471
R7904 VDD.n2760 VDD.n2759 0.00326471
R7905 VDD.n2788 VDD.n2787 0.00326471
R7906 VDD.n2807 VDD.n2806 0.00326471
R7907 VDD.n2826 VDD.n2825 0.00326471
R7908 VDD.n2845 VDD.n2844 0.00326471
R7909 VDD.n2865 VDD.n2864 0.00326471
R7910 VDD.n2884 VDD.n1288 0.00326471
R7911 VDD.n663 VDD.n644 0.00322032
R7912 VDD.n1079 VDD.n1073 0.00321739
R7913 VDD.n819 VDD.n813 0.00321739
R7914 VDD.n851 VDD.n844 0.00321739
R7915 VDD.n1055 VDD.n1048 0.00321739
R7916 VDD.n161 VDD.n155 0.00321739
R7917 VDD.n520 VDD.n514 0.00321739
R7918 VDD.n652 VDD.n645 0.00321739
R7919 VDD.n654 VDD 0.00321739
R7920 VDD.n544 VDD.n537 0.00321739
R7921 VDD.n1264 VDD.n707 0.0032134
R7922 VDD.n1253 VDD.n1252 0.0032134
R7923 VDD.n866 VDD.n825 0.00311649
R7924 VDD.n740 VDD.n706 0.00310417
R7925 VDD.n620 VDD.n145 0.00310417
R7926 VDD.n478 VDD.n392 0.00310417
R7927 VDD.n2982 VDD.n2981 0.00292685
R7928 VDD.n2982 VDD.n39 0.00292685
R7929 VDD.n1018 VDD.n1004 0.00290385
R7930 VDD.n1260 VDD.n709 0.00290385
R7931 VDD.n312 VDD.n283 0.00290385
R7932 VDD.n2925 VDD.n2910 0.00284596
R7933 VDD.n1170 VDD.n1169 0.00281481
R7934 VDD.n319 VDD.n280 0.00272887
R7935 VDD.n1192 VDD.n1191 0.00269298
R7936 VDD.n1900 VDD.n1872 0.00257353
R7937 VDD.n1870 VDD.n1860 0.00257353
R7938 VDD.n1930 VDD.n1858 0.00257353
R7939 VDD.n1952 VDD.n1844 0.00257353
R7940 VDD.n1972 VDD.n1833 0.00257353
R7941 VDD.n2106 VDD.n1748 0.00257353
R7942 VDD.n2126 VDD.n1738 0.00257353
R7943 VDD.n1736 VDD.n1726 0.00257353
R7944 VDD.n2156 VDD.n1724 0.00257353
R7945 VDD.n2178 VDD.n1710 0.00257353
R7946 VDD.n2198 VDD.n1699 0.00257353
R7947 VDD.n2332 VDD.n1614 0.00257353
R7948 VDD.n2352 VDD.n1604 0.00257353
R7949 VDD.n1602 VDD.n1592 0.00257353
R7950 VDD.n2382 VDD.n1590 0.00257353
R7951 VDD.n2404 VDD.n1576 0.00257353
R7952 VDD.n2424 VDD.n1565 0.00257353
R7953 VDD.n2558 VDD.n1480 0.00257353
R7954 VDD.n2578 VDD.n1470 0.00257353
R7955 VDD.n1468 VDD.n1458 0.00257353
R7956 VDD.n2608 VDD.n1456 0.00257353
R7957 VDD.n2630 VDD.n1442 0.00257353
R7958 VDD.n2650 VDD.n1431 0.00257353
R7959 VDD.n81 VDD.n56 0.00245312
R7960 VDD.n2939 VDD.n2921 0.0024405
R7961 VDD.n2799 VDD.n1342 0.00239394
R7962 VDD.n2818 VDD.n1331 0.00239394
R7963 VDD.n2837 VDD.n1320 0.00239394
R7964 VDD.n2856 VDD.n1309 0.00239394
R7965 VDD.n2876 VDD.n1293 0.00239394
R7966 VDD.n1888 VDD.n1874 0.00239394
R7967 VDD.n1909 VDD.n1863 0.00239394
R7968 VDD.n1936 VDD.n1935 0.00239394
R7969 VDD.n1944 VDD.n1841 0.00239394
R7970 VDD.n1964 VDD.n1830 0.00239394
R7971 VDD.n1983 VDD.n1817 0.00239394
R7972 VDD.n1994 VDD.n1808 0.00239394
R7973 VDD.n1802 VDD.n1793 0.00239394
R7974 VDD.n2029 VDD.n1787 0.00239394
R7975 VDD.n2061 VDD.n1773 0.00239394
R7976 VDD.n2070 VDD.n1768 0.00239394
R7977 VDD.n2094 VDD.n1755 0.00239394
R7978 VDD.n2114 VDD.n1740 0.00239394
R7979 VDD.n2135 VDD.n1729 0.00239394
R7980 VDD.n2162 VDD.n2161 0.00239394
R7981 VDD.n2170 VDD.n1707 0.00239394
R7982 VDD.n2190 VDD.n1696 0.00239394
R7983 VDD.n2209 VDD.n1683 0.00239394
R7984 VDD.n2220 VDD.n1674 0.00239394
R7985 VDD.n1668 VDD.n1659 0.00239394
R7986 VDD.n2255 VDD.n1653 0.00239394
R7987 VDD.n2287 VDD.n1639 0.00239394
R7988 VDD.n2296 VDD.n1634 0.00239394
R7989 VDD.n2320 VDD.n1621 0.00239394
R7990 VDD.n2340 VDD.n1606 0.00239394
R7991 VDD.n2361 VDD.n1595 0.00239394
R7992 VDD.n2388 VDD.n2387 0.00239394
R7993 VDD.n2396 VDD.n1573 0.00239394
R7994 VDD.n2416 VDD.n1562 0.00239394
R7995 VDD.n2435 VDD.n1549 0.00239394
R7996 VDD.n2446 VDD.n1540 0.00239394
R7997 VDD.n1534 VDD.n1525 0.00239394
R7998 VDD.n2481 VDD.n1519 0.00239394
R7999 VDD.n2513 VDD.n1505 0.00239394
R8000 VDD.n2522 VDD.n1500 0.00239394
R8001 VDD.n2546 VDD.n1487 0.00239394
R8002 VDD.n2566 VDD.n1472 0.00239394
R8003 VDD.n2587 VDD.n1461 0.00239394
R8004 VDD.n2614 VDD.n2613 0.00239394
R8005 VDD.n2622 VDD.n1439 0.00239394
R8006 VDD.n2642 VDD.n1428 0.00239394
R8007 VDD.n2661 VDD.n1415 0.00239394
R8008 VDD.n2672 VDD.n1406 0.00239394
R8009 VDD.n1400 VDD.n1391 0.00239394
R8010 VDD.n2707 VDD.n1385 0.00239394
R8011 VDD.n2739 VDD.n1371 0.00239394
R8012 VDD.n2748 VDD.n1366 0.00239394
R8013 VDD.n2771 VDD.n1352 0.00239394
R8014 VDD.n1887 VDD.n1873 0.00239394
R8015 VDD.n1908 VDD.n1862 0.00239394
R8016 VDD.n1934 VDD.n1854 0.00239394
R8017 VDD.n1945 VDD.n1842 0.00239394
R8018 VDD.n1965 VDD.n1831 0.00239394
R8019 VDD.n1984 VDD.n1815 0.00239394
R8020 VDD.n1993 VDD.n1809 0.00239394
R8021 VDD.n1800 VDD.n1794 0.00239394
R8022 VDD.n2028 VDD.n1785 0.00239394
R8023 VDD.n2040 VDD.n1774 0.00239394
R8024 VDD.n2071 VDD.n1766 0.00239394
R8025 VDD.n2095 VDD.n1753 0.00239394
R8026 VDD.n2113 VDD.n1739 0.00239394
R8027 VDD.n2134 VDD.n1728 0.00239394
R8028 VDD.n2160 VDD.n1720 0.00239394
R8029 VDD.n2171 VDD.n1708 0.00239394
R8030 VDD.n2191 VDD.n1697 0.00239394
R8031 VDD.n2210 VDD.n1681 0.00239394
R8032 VDD.n2219 VDD.n1675 0.00239394
R8033 VDD.n1666 VDD.n1660 0.00239394
R8034 VDD.n2254 VDD.n1651 0.00239394
R8035 VDD.n2266 VDD.n1640 0.00239394
R8036 VDD.n2297 VDD.n1632 0.00239394
R8037 VDD.n2321 VDD.n1619 0.00239394
R8038 VDD.n2339 VDD.n1605 0.00239394
R8039 VDD.n2360 VDD.n1594 0.00239394
R8040 VDD.n2386 VDD.n1586 0.00239394
R8041 VDD.n2397 VDD.n1574 0.00239394
R8042 VDD.n2417 VDD.n1563 0.00239394
R8043 VDD.n2436 VDD.n1547 0.00239394
R8044 VDD.n2445 VDD.n1541 0.00239394
R8045 VDD.n1532 VDD.n1526 0.00239394
R8046 VDD.n2480 VDD.n1517 0.00239394
R8047 VDD.n2492 VDD.n1506 0.00239394
R8048 VDD.n2523 VDD.n1498 0.00239394
R8049 VDD.n2547 VDD.n1485 0.00239394
R8050 VDD.n2565 VDD.n1471 0.00239394
R8051 VDD.n2586 VDD.n1460 0.00239394
R8052 VDD.n2612 VDD.n1452 0.00239394
R8053 VDD.n2623 VDD.n1440 0.00239394
R8054 VDD.n2643 VDD.n1429 0.00239394
R8055 VDD.n2662 VDD.n1413 0.00239394
R8056 VDD.n2671 VDD.n1407 0.00239394
R8057 VDD.n1398 VDD.n1392 0.00239394
R8058 VDD.n2706 VDD.n1383 0.00239394
R8059 VDD.n2718 VDD.n1372 0.00239394
R8060 VDD.n2749 VDD.n1364 0.00239394
R8061 VDD.n2762 VDD.n1353 0.00239394
R8062 VDD.n2800 VDD.n1340 0.00239394
R8063 VDD.n2819 VDD.n1329 0.00239394
R8064 VDD.n2838 VDD.n1318 0.00239394
R8065 VDD.n2857 VDD.n1307 0.00239394
R8066 VDD.n2877 VDD.n1291 0.00239394
R8067 VDD.n1087 VDD.n1084 0.00233824
R8068 VDD.n654 VDD 0.00233824
R8069 VDD.n2931 VDD.n2930 0.00227969
R8070 VDD.n2883 VDD.n1287 0.00224074
R8071 VDD.n269 VDD.n268 0.00220831
R8072 VDD.n270 VDD.n269 0.0021949
R8073 VDD.n2885 VDD.n1286 0.00213953
R8074 VDD.n2939 VDD.n2938 0.00208589
R8075 VDD.n3005 VDD.n11 0.00196875
R8076 VDD.n16 VDD.n13 0.00196875
R8077 VDD.n166 VDD.n165 0.00192045
R8078 VDD.n2971 VDD.n2966 0.00180208
R8079 VDD.n731 VDD.n703 0.00180208
R8080 VDD.n1109 VDD.n1108 0.00180208
R8081 VDD.n593 VDD.n233 0.00180208
R8082 VDD.n366 VDD.n328 0.00180208
R8083 VDD.n2962 VDD.n1276 0.00179432
R8084 VDD.n307 VDD.n280 0.00172678
R8085 VDD.n1879 VDD 0.00170513
R8086 VDD VDD.n1747 0.00170513
R8087 VDD VDD.n1613 0.00170513
R8088 VDD VDD.n1479 0.00170513
R8089 VDD.n2980 VDD.n1276 0.00163253
R8090 VDD.n2938 VDD.n2937 0.00163253
R8091 VDD.n2986 VDD.n37 0.00147656
R8092 VDD.n2945 VDD.n2909 0.00138985
R8093 VDD.n1881 VDD.n1878 0.00119118
R8094 VDD.n1886 VDD.n1878 0.00119118
R8095 VDD.n1901 VDD.n1869 0.00119118
R8096 VDD.n1907 VDD.n1869 0.00119118
R8097 VDD.n1923 VDD.n1922 0.00119118
R8098 VDD.n1924 VDD.n1923 0.00119118
R8099 VDD.n1929 VDD.n1846 0.00119118
R8100 VDD.n1946 VDD.n1846 0.00119118
R8101 VDD.n1951 VDD.n1835 0.00119118
R8102 VDD.n1966 VDD.n1835 0.00119118
R8103 VDD.n1971 VDD.n1813 0.00119118
R8104 VDD.n1985 VDD.n1813 0.00119118
R8105 VDD.n1992 VDD.n1991 0.00119118
R8106 VDD.n1991 VDD.n1798 0.00119118
R8107 VDD.n2012 VDD.n1795 0.00119118
R8108 VDD.n2022 VDD.n1795 0.00119118
R8109 VDD.n2017 VDD.n1784 0.00119118
R8110 VDD.n2046 VDD.n1784 0.00119118
R8111 VDD.n2052 VDD.n2051 0.00119118
R8112 VDD.n2052 VDD.n1780 0.00119118
R8113 VDD.n2073 VDD.n2072 0.00119118
R8114 VDD.n2073 VDD.n1763 0.00119118
R8115 VDD.n2097 VDD.n2096 0.00119118
R8116 VDD.n2097 VDD.n1750 0.00119118
R8117 VDD.n2107 VDD.n1746 0.00119118
R8118 VDD.n2112 VDD.n1746 0.00119118
R8119 VDD.n2127 VDD.n1735 0.00119118
R8120 VDD.n2133 VDD.n1735 0.00119118
R8121 VDD.n2149 VDD.n2148 0.00119118
R8122 VDD.n2150 VDD.n2149 0.00119118
R8123 VDD.n2155 VDD.n1712 0.00119118
R8124 VDD.n2172 VDD.n1712 0.00119118
R8125 VDD.n2177 VDD.n1701 0.00119118
R8126 VDD.n2192 VDD.n1701 0.00119118
R8127 VDD.n2197 VDD.n1679 0.00119118
R8128 VDD.n2211 VDD.n1679 0.00119118
R8129 VDD.n2218 VDD.n2217 0.00119118
R8130 VDD.n2217 VDD.n1664 0.00119118
R8131 VDD.n2238 VDD.n1661 0.00119118
R8132 VDD.n2248 VDD.n1661 0.00119118
R8133 VDD.n2243 VDD.n1650 0.00119118
R8134 VDD.n2272 VDD.n1650 0.00119118
R8135 VDD.n2278 VDD.n2277 0.00119118
R8136 VDD.n2278 VDD.n1646 0.00119118
R8137 VDD.n2299 VDD.n2298 0.00119118
R8138 VDD.n2299 VDD.n1629 0.00119118
R8139 VDD.n2323 VDD.n2322 0.00119118
R8140 VDD.n2323 VDD.n1616 0.00119118
R8141 VDD.n2333 VDD.n1612 0.00119118
R8142 VDD.n2338 VDD.n1612 0.00119118
R8143 VDD.n2353 VDD.n1601 0.00119118
R8144 VDD.n2359 VDD.n1601 0.00119118
R8145 VDD.n2375 VDD.n2374 0.00119118
R8146 VDD.n2376 VDD.n2375 0.00119118
R8147 VDD.n2381 VDD.n1578 0.00119118
R8148 VDD.n2398 VDD.n1578 0.00119118
R8149 VDD.n2403 VDD.n1567 0.00119118
R8150 VDD.n2418 VDD.n1567 0.00119118
R8151 VDD.n2423 VDD.n1545 0.00119118
R8152 VDD.n2437 VDD.n1545 0.00119118
R8153 VDD.n2444 VDD.n2443 0.00119118
R8154 VDD.n2443 VDD.n1530 0.00119118
R8155 VDD.n2464 VDD.n1527 0.00119118
R8156 VDD.n2474 VDD.n1527 0.00119118
R8157 VDD.n2469 VDD.n1516 0.00119118
R8158 VDD.n2498 VDD.n1516 0.00119118
R8159 VDD.n2504 VDD.n2503 0.00119118
R8160 VDD.n2504 VDD.n1512 0.00119118
R8161 VDD.n2525 VDD.n2524 0.00119118
R8162 VDD.n2525 VDD.n1495 0.00119118
R8163 VDD.n2549 VDD.n2548 0.00119118
R8164 VDD.n2549 VDD.n1482 0.00119118
R8165 VDD.n2559 VDD.n1478 0.00119118
R8166 VDD.n2564 VDD.n1478 0.00119118
R8167 VDD.n2579 VDD.n1467 0.00119118
R8168 VDD.n2585 VDD.n1467 0.00119118
R8169 VDD.n2601 VDD.n2600 0.00119118
R8170 VDD.n2602 VDD.n2601 0.00119118
R8171 VDD.n2607 VDD.n1444 0.00119118
R8172 VDD.n2624 VDD.n1444 0.00119118
R8173 VDD.n2629 VDD.n1433 0.00119118
R8174 VDD.n2644 VDD.n1433 0.00119118
R8175 VDD.n2649 VDD.n1411 0.00119118
R8176 VDD.n2663 VDD.n1411 0.00119118
R8177 VDD.n2670 VDD.n2669 0.00119118
R8178 VDD.n2669 VDD.n1396 0.00119118
R8179 VDD.n2690 VDD.n1393 0.00119118
R8180 VDD.n2700 VDD.n1393 0.00119118
R8181 VDD.n2695 VDD.n1382 0.00119118
R8182 VDD.n2724 VDD.n1382 0.00119118
R8183 VDD.n2730 VDD.n2729 0.00119118
R8184 VDD.n2730 VDD.n1378 0.00119118
R8185 VDD.n2751 VDD.n2750 0.00119118
R8186 VDD.n2751 VDD.n1360 0.00119118
R8187 VDD.n2755 VDD.n2754 0.00119118
R8188 VDD.n2755 VDD.n1350 0.00119118
R8189 VDD.n2783 VDD.n2782 0.00119118
R8190 VDD.n2783 VDD.n1348 0.00119118
R8191 VDD.n2802 VDD.n2801 0.00119118
R8192 VDD.n2802 VDD.n1337 0.00119118
R8193 VDD.n2821 VDD.n2820 0.00119118
R8194 VDD.n2821 VDD.n1326 0.00119118
R8195 VDD.n2840 VDD.n2839 0.00119118
R8196 VDD.n2840 VDD.n1315 0.00119118
R8197 VDD.n2859 VDD.n2858 0.00119118
R8198 VDD.n2859 VDD.n1303 0.00119118
R8199 VDD.n1292 VDD.n1290 0.00119118
R8200 VDD.n2881 VDD.n1290 0.00119118
R8201 VDD.n320 VDD.n319 0.00117835
R8202 VDD.n1228 VDD.n766 0.00115104
R8203 VDD.n1220 VDD.n1219 0.00115104
R8204 VDD.n1193 VDD.n798 0.00115104
R8205 VDD.n920 VDD.n919 0.00115104
R8206 VDD.n1182 VDD.n905 0.00115104
R8207 VDD.n1168 VDD.n934 0.00115104
R8208 VDD.n710 VDD.n707 0.00114537
R8209 VDD.n2903 VDD.n2901 0.0011215
R8210 VDD.n1883 VDD.n1882 0.00110256
R8211 VDD.n1903 VDD.n1902 0.00110256
R8212 VDD.n1861 VDD.n1859 0.00110256
R8213 VDD.n1928 VDD.n1845 0.00110256
R8214 VDD.n1950 VDD.n1834 0.00110256
R8215 VDD.n1970 VDD.n1812 0.00110256
R8216 VDD.n1990 VDD.n1989 0.00110256
R8217 VDD.n2021 VDD.n2015 0.00110256
R8218 VDD.n2047 VDD.n1783 0.00110256
R8219 VDD.n2054 VDD.n2053 0.00110256
R8220 VDD.n2075 VDD.n2074 0.00110256
R8221 VDD.n2099 VDD.n2098 0.00110256
R8222 VDD.n2109 VDD.n2108 0.00110256
R8223 VDD.n2129 VDD.n2128 0.00110256
R8224 VDD.n1727 VDD.n1725 0.00110256
R8225 VDD.n2154 VDD.n1711 0.00110256
R8226 VDD.n2176 VDD.n1700 0.00110256
R8227 VDD.n2196 VDD.n1678 0.00110256
R8228 VDD.n2216 VDD.n2215 0.00110256
R8229 VDD.n2247 VDD.n2241 0.00110256
R8230 VDD.n2273 VDD.n1649 0.00110256
R8231 VDD.n2280 VDD.n2279 0.00110256
R8232 VDD.n2301 VDD.n2300 0.00110256
R8233 VDD.n2325 VDD.n2324 0.00110256
R8234 VDD.n2335 VDD.n2334 0.00110256
R8235 VDD.n2355 VDD.n2354 0.00110256
R8236 VDD.n1593 VDD.n1591 0.00110256
R8237 VDD.n2380 VDD.n1577 0.00110256
R8238 VDD.n2402 VDD.n1566 0.00110256
R8239 VDD.n2422 VDD.n1544 0.00110256
R8240 VDD.n2442 VDD.n2441 0.00110256
R8241 VDD.n2473 VDD.n2467 0.00110256
R8242 VDD.n2499 VDD.n1515 0.00110256
R8243 VDD.n2506 VDD.n2505 0.00110256
R8244 VDD.n2527 VDD.n2526 0.00110256
R8245 VDD.n2551 VDD.n2550 0.00110256
R8246 VDD.n2561 VDD.n2560 0.00110256
R8247 VDD.n2581 VDD.n2580 0.00110256
R8248 VDD.n1459 VDD.n1457 0.00110256
R8249 VDD.n2606 VDD.n1443 0.00110256
R8250 VDD.n2628 VDD.n1432 0.00110256
R8251 VDD.n2648 VDD.n1410 0.00110256
R8252 VDD.n2668 VDD.n2667 0.00110256
R8253 VDD.n2699 VDD.n2693 0.00110256
R8254 VDD.n2725 VDD.n1381 0.00110256
R8255 VDD.n2732 VDD.n2731 0.00110256
R8256 VDD.n2753 VDD.n2752 0.00110256
R8257 VDD.n2756 VDD.n1349 0.00110256
R8258 VDD.n2785 VDD.n2784 0.00108025
R8259 VDD.n2804 VDD.n2803 0.00108025
R8260 VDD.n2823 VDD.n2822 0.00108025
R8261 VDD.n2842 VDD.n2841 0.00108025
R8262 VDD.n2861 VDD.n2860 0.00108025
R8263 VDD.n2882 VDD.n1289 0.00108025
R8264 VDD.n2963 VDD.n2962 0.00098537
R8265 VDD.n1023 VDD.n1021 0.000984536
R8266 VDD.n2961 VDD.n2960 0.000932515
R8267 VDD.n3007 VDD.n3006 0.000837321
R8268 VDD.n2938 VDD.n2909 0.00082358
R8269 VDD VDD.n22 0.00072488
R8270 VDD.n1253 VDD.n711 0.000693814
R8271 VDD.n867 VDD.n866 0.000693814
R8272 VDD.n1062 VDD.n1034 0.000693814
R8273 VDD.n668 VDD.n667 0.000693814
R8274 VDD.n561 VDD.n560 0.000693814
R8275 VDD.n3007 VDD.n22 0.00061244
R8276 VDD.n868 VDD.n867 0.000596907
R8277 VDD.n2937 VDD.n2922 0.000580895
R8278 VDD.n2945 VDD.n2910 0.000580895
R8279 VDD.n2931 VDD.n2925 0.000580895
R8280 sar_retimer[3].n0 sar_retimer[3].t1 207.373
R8281 sar_retimer[3].n1 sar_retimer[3] 67.3346
R8282 sar_retimer[3].n1 sar_retimer[3].t0 32.6903
R8283 sar_retimer[3] sar_retimer[3].n0 9.01934
R8284 sar_retimer[3].n0 sar_retimer[3] 7.45876
R8285 sar_retimer[3] sar_retimer[3].n2 3.7337
R8286 sar_retimer[3].n2 sar_retimer[3] 2.09635
R8287 sar_retimer[3].n2 sar_retimer[3].n1 1.20577
R8288 sar_logic[6].n0 sar_logic[6].t1 331.51
R8289 sar_logic[6].n0 sar_logic[6].t0 209.403
R8290 sar_logic[6].n1 sar_logic[6].n0 76.0005
R8291 sar_logic[6] sar_logic[6].n1 8.58587
R8292 sar_logic[6].n1 sar_logic[6] 2.02977
R8293 eob.t11 eob.t5 221.72
R8294 eob.t16 eob.t11 221.72
R8295 eob.t10 eob.t16 221.72
R8296 eob.t7 eob.t10 221.72
R8297 eob.t13 eob.t7 221.72
R8298 eob.t14 eob.t20 221.72
R8299 eob.t1 eob.t14 221.72
R8300 eob.t15 eob.t1 221.72
R8301 eob.t9 eob.t15 221.72
R8302 eob.t2 eob.t9 221.72
R8303 eob.t17 eob.t2 221.72
R8304 eob.t3 eob.t17 221.72
R8305 eob.t18 eob.t0 221.72
R8306 eob.t4 eob.t18 221.72
R8307 eob.t19 eob.t4 221.72
R8308 eob.t12 eob.t19 221.72
R8309 eob.t6 eob.t12 221.72
R8310 eob.t21 eob.t6 221.72
R8311 eob.t8 eob.t21 221.72
R8312 eob.n5 eob.t13 154.8
R8313 eob.n0 eob 89.9738
R8314 eob.n1 eob.t3 78.7272
R8315 eob.n0 eob.t8 74.6592
R8316 eob.n2 eob 40.1672
R8317 eob.n3 eob.n1 32.1338
R8318 eob eob.n1 21.4227
R8319 eob.n4 eob.n0 21.3547
R8320 eob.n4 eob.n3 17.8279
R8321 eob.n5 eob.n4 13.4163
R8322 eob.n2 eob 11.8854
R8323 eob.n3 eob.n2 3.96214
R8324 eob.n6 eob 1.64944
R8325 eob.n6 eob 0.10169
R8326 eob eob.n6 0.00215441
R8327 eob.n6 eob.n5 0.00197059
R8328 sar_retimer[2].n2 sar_retimer[2].t0 117.424
R8329 sar_retimer[2].n1 sar_retimer[2].n0 73.2739
R8330 sar_retimer[2].n0 sar_retimer[2].t1 71.9813
R8331 sar_retimer[2] sar_retimer[2].n2 66.6967
R8332 sar_retimer[2].n1 sar_retimer[2] 13.6746
R8333 sar_retimer[2].n4 sar_retimer[2].n3 12.8005
R8334 sar_retimer[2].n2 sar_retimer[2] 6.64665
R8335 sar_retimer[2] sar_retimer[2].n4 2.21588
R8336 sar_retimer[2] sar_retimer[2].n1 1.9648
R8337 sar_retimer[2].n3 sar_retimer[2] 1.72358
R8338 delay_code[1] delay_code[1].t0 140.387
R8339 delay_code[1].n0 delay_code[1].t1 140.34
R8340 delay_code[1].n0 delay_code[1] 0.204667
R8341 delay_code[1] delay_code[1].n0 0.00218919
R8342 sar_logic[3].n2 sar_logic[3].t0 330.616
R8343 sar_logic[3].n0 sar_logic[3].t1 195.121
R8344 sar_logic[3].n3 sar_logic[3] 14.9071
R8345 sar_logic[3].n1 sar_logic[3].n0 14.282
R8346 sar_logic[3].n4 sar_logic[3].n2 8.76429
R8347 sar_logic[3].n3 sar_logic[3] 7.37062
R8348 sar_logic[3] sar_logic[3].n5 2.02977
R8349 sar_logic[3].n2 sar_logic[3].n1 0.893093
R8350 sar_logic[3].n4 sar_logic[3].n3 0.620445
R8351 sar_logic[3].n5 sar_logic[3].n4 0.156598
R8352 sar_logic[2].n2 sar_logic[2].t0 329.724
R8353 sar_logic[2].n0 sar_logic[2].t1 196.013
R8354 sar_logic[2].n1 sar_logic[2].n0 13.3894
R8355 sar_logic[2].n4 sar_logic[2].n2 8.76429
R8356 sar_logic[2].n3 sar_logic[2] 7.21403
R8357 sar_logic[2].n3 sar_logic[2] 3.7454
R8358 sar_logic[2] sar_logic[2].n5 2.02977
R8359 sar_logic[2].n2 sar_logic[2].n1 1.78569
R8360 sar_logic[2].n4 sar_logic[2].n3 0.620934
R8361 sar_logic[2].n5 sar_logic[2].n4 0.312695
R8362 sar_retimer[1].n2 sar_retimer[1].t1 425.096
R8363 sar_retimer[1].n3 sar_retimer[1].t1 417.519
R8364 sar_retimer[1].n4 sar_retimer[1].n3 64.3701
R8365 sar_retimer[1].n1 sar_retimer[1].t0 32.9519
R8366 sar_retimer[1] sar_retimer[1].n2 10.0928
R8367 sar_retimer[1].n3 sar_retimer[1] 6.64665
R8368 sar_retimer[1].n2 sar_retimer[1] 6.64665
R8369 sar_retimer[1].n1 sar_retimer[1].n0 4.64355
R8370 sar_retimer[1] sar_retimer[1].n4 1.85845
R8371 sar_retimer[1] sar_retimer[1].n1 0.492808
R8372 sar_retimer[1].n0 sar_retimer[1] 0.426349
R8373 sar_retimer[0].n0 sar_retimer[0].t1 417.519
R8374 sar_retimer[0].n1 sar_retimer[0].t1 143.925
R8375 sar_retimer[0] sar_retimer[0].t0 119.147
R8376 sar_retimer[0].n0 sar_retimer[0] 66.6967
R8377 sar_retimer[0].n2 sar_retimer[0] 12.7994
R8378 sar_retimer[0].n1 sar_retimer[0] 10.3226
R8379 sar_retimer[0] sar_retimer[0].n0 6.64665
R8380 sar_retimer[0] sar_retimer[0].n2 3.97979
R8381 sar_retimer[0].n2 sar_retimer[0].n1 1.42978
R8382 x2.x10.Y x2.x10.Y.t5 154.847
R8383 x2.x10.Y x2.x10.Y.t2 154.8
R8384 x2.x10.Y x2.x10.Y.t9 154.8
R8385 x2.x10.Y x2.x10.Y.t3 154.8
R8386 x2.x10.Y x2.x10.Y.t6 154.8
R8387 x2.x10.Y x2.x10.Y.t4 154.8
R8388 x2.x10.Y x2.x10.Y.t7 154.8
R8389 x2.x10.Y x2.x10.Y.t8 154.8
R8390 x2.x10.Y.n0 x2.x10.Y 134.239
R8391 x2.x10.Y x2.x10.Y.t0 106.635
R8392 x2.x10.Y.n2 x2.x10.Y.t1 24.6567
R8393 x2.x10.Y.n5 x2.x10.Y.n4 12.4089
R8394 x2.x10.Y.n3 x2.x10.Y.n2 9.12522
R8395 x2.x10.Y.n4 x2.x10.Y.n3 7.34048
R8396 x2.x10.Y.n5 x2.x10.Y 2.22659
R8397 x2.x10.Y.n2 x2.x10.Y.n1 1.93377
R8398 x2.x10.Y x2.x10.Y.n5 1.55202
R8399 x2.x10.Y.n3 x2.x10.Y.n0 0.69928
R8400 x2.x5[7].floating.n154 x2.x5[7].floating.t1 68.0345
R8401 x2.x5[7].floating.n142 x2.x5[7].floating.t2 68.0345
R8402 x2.x5[7].floating.n12 x2.x5[7].floating.t5 68.0345
R8403 x2.x5[7].floating.n24 x2.x5[7].floating.t3 68.0345
R8404 x2.x5[7].floating.n54 x2.x5[7].floating.t0 68.0345
R8405 x2.x5[7].floating.n72 x2.x5[7].floating.t7 68.0345
R8406 x2.x5[7].floating.n84 x2.x5[7].floating.t4 68.0345
R8407 x2.x5[7].floating.n42 x2.x5[7].floating.t6 68.0345
R8408 x2.x5[7].floating.n103 x2.x5[7].floating.n65 0.660401
R8409 x2.x5[7].floating.n112 x2.x5[7].floating.n50 0.660401
R8410 x2.x5[7].floating.n121 x2.x5[7].floating.n35 0.660401
R8411 x2.x5[7].floating.n130 x2.x5[7].floating.n20 0.660401
R8412 x2.x5[7].floating.n139 x2.x5[7].floating.n5 0.660401
R8413 x2.x5[7].floating.n90 x2.x5[7].floating.n89 0.320345
R8414 x2.x5[7].floating.n160 x2.x5[7].floating.n159 0.308269
R8415 x2.x5[7].floating.n161 x2.x5[7].floating.n160 0.173084
R8416 x2.x5[7].floating.n91 x2.x5[7].floating.n90 0.162103
R8417 x2.x5[7].floating.n160 x2.x5[7].floating 0.100688
R8418 x2.x5[7].floating.n90 x2.x5[7].floating 0.0755007
R8419 x2.x5[7].floating.n66 x2.x5[7].floating.n65 0.0716912
R8420 x2.x5[7].floating.n65 x2.x5[7].floating.n64 0.0716912
R8421 x2.x5[7].floating.n36 x2.x5[7].floating.n35 0.0716912
R8422 x2.x5[7].floating.n35 x2.x5[7].floating.n34 0.0716912
R8423 x2.x5[7].floating.n6 x2.x5[7].floating.n5 0.0716912
R8424 x2.x5[7].floating.n5 x2.x5[7].floating.n4 0.0716912
R8425 x2.x5[7].floating.n104 x2.x5[7].floating.n103 0.0716912
R8426 x2.x5[7].floating.n122 x2.x5[7].floating.n121 0.0716912
R8427 x2.x5[7].floating.n140 x2.x5[7].floating.n139 0.0716912
R8428 x2.x5[7].floating.n70 x2.x5[7].floating.n69 0.0557941
R8429 x2.x5[7].floating.n69 x2.x5[7].floating.n68 0.0557941
R8430 x2.x5[7].floating.n68 x2.x5[7].floating.n67 0.0557941
R8431 x2.x5[7].floating.n67 x2.x5[7].floating.n66 0.0557941
R8432 x2.x5[7].floating.n64 x2.x5[7].floating.n63 0.0557941
R8433 x2.x5[7].floating.n63 x2.x5[7].floating.n62 0.0557941
R8434 x2.x5[7].floating.n62 x2.x5[7].floating.n61 0.0557941
R8435 x2.x5[7].floating.n61 x2.x5[7].floating.n60 0.0557941
R8436 x2.x5[7].floating.n40 x2.x5[7].floating.n39 0.0557941
R8437 x2.x5[7].floating.n39 x2.x5[7].floating.n38 0.0557941
R8438 x2.x5[7].floating.n38 x2.x5[7].floating.n37 0.0557941
R8439 x2.x5[7].floating.n37 x2.x5[7].floating.n36 0.0557941
R8440 x2.x5[7].floating.n34 x2.x5[7].floating.n33 0.0557941
R8441 x2.x5[7].floating.n33 x2.x5[7].floating.n32 0.0557941
R8442 x2.x5[7].floating.n32 x2.x5[7].floating.n31 0.0557941
R8443 x2.x5[7].floating.n31 x2.x5[7].floating.n30 0.0557941
R8444 x2.x5[7].floating.n10 x2.x5[7].floating.n9 0.0557941
R8445 x2.x5[7].floating.n9 x2.x5[7].floating.n8 0.0557941
R8446 x2.x5[7].floating.n8 x2.x5[7].floating.n7 0.0557941
R8447 x2.x5[7].floating.n7 x2.x5[7].floating.n6 0.0557941
R8448 x2.x5[7].floating.n4 x2.x5[7].floating.n3 0.0557941
R8449 x2.x5[7].floating.n3 x2.x5[7].floating.n2 0.0557941
R8450 x2.x5[7].floating.n2 x2.x5[7].floating.n1 0.0557941
R8451 x2.x5[7].floating.n1 x2.x5[7].floating.n0 0.0557941
R8452 x2.x5[7].floating.n99 x2.x5[7].floating.n98 0.0557941
R8453 x2.x5[7].floating.n100 x2.x5[7].floating.n99 0.0557941
R8454 x2.x5[7].floating.n101 x2.x5[7].floating.n100 0.0557941
R8455 x2.x5[7].floating.n102 x2.x5[7].floating.n101 0.0557941
R8456 x2.x5[7].floating.n106 x2.x5[7].floating.n105 0.0557941
R8457 x2.x5[7].floating.n107 x2.x5[7].floating.n106 0.0557941
R8458 x2.x5[7].floating.n108 x2.x5[7].floating.n107 0.0557941
R8459 x2.x5[7].floating.n117 x2.x5[7].floating.n116 0.0557941
R8460 x2.x5[7].floating.n118 x2.x5[7].floating.n117 0.0557941
R8461 x2.x5[7].floating.n119 x2.x5[7].floating.n118 0.0557941
R8462 x2.x5[7].floating.n120 x2.x5[7].floating.n119 0.0557941
R8463 x2.x5[7].floating.n124 x2.x5[7].floating.n123 0.0557941
R8464 x2.x5[7].floating.n125 x2.x5[7].floating.n124 0.0557941
R8465 x2.x5[7].floating.n126 x2.x5[7].floating.n125 0.0557941
R8466 x2.x5[7].floating.n135 x2.x5[7].floating.n134 0.0557941
R8467 x2.x5[7].floating.n136 x2.x5[7].floating.n135 0.0557941
R8468 x2.x5[7].floating.n137 x2.x5[7].floating.n136 0.0557941
R8469 x2.x5[7].floating.n138 x2.x5[7].floating.n137 0.0557941
R8470 x2.x5[7].floating.n171 x2.x5[7].floating.n170 0.0557941
R8471 x2.x5[7].floating.n170 x2.x5[7].floating.n169 0.0557941
R8472 x2.x5[7].floating.n169 x2.x5[7].floating.n168 0.0557941
R8473 x2.x5[7].floating.n95 x2.x5[7].floating.n94 0.0537206
R8474 x2.x5[7].floating.n113 x2.x5[7].floating.n112 0.0537206
R8475 x2.x5[7].floating.n131 x2.x5[7].floating.n130 0.0537206
R8476 x2.x5[7].floating.n164 x2.x5[7].floating.n163 0.0537206
R8477 x2.x5[7].floating.n94 x2.x5[7].floating.n93 0.0530294
R8478 x2.x5[7].floating.n112 x2.x5[7].floating.n111 0.0530294
R8479 x2.x5[7].floating.n130 x2.x5[7].floating.n129 0.0530294
R8480 x2.x5[7].floating.n165 x2.x5[7].floating.n164 0.0530294
R8481 x2.x5[7].floating.n80 x2.x5[7].floating.n79 0.0529559
R8482 x2.x5[7].floating.n50 x2.x5[7].floating.n49 0.0529559
R8483 x2.x5[7].floating.n20 x2.x5[7].floating.n19 0.0529559
R8484 x2.x5[7].floating.n151 x2.x5[7].floating.n150 0.0529559
R8485 x2.x5[7].floating.n81 x2.x5[7].floating.n80 0.0524559
R8486 x2.x5[7].floating.n51 x2.x5[7].floating.n50 0.0524559
R8487 x2.x5[7].floating.n21 x2.x5[7].floating.n20 0.0524559
R8488 x2.x5[7].floating.n150 x2.x5[7].floating.n149 0.0524559
R8489 x2.x5[7].floating.n109 x2.x5[7].floating.n108 0.0523382
R8490 x2.x5[7].floating.n127 x2.x5[7].floating.n126 0.0523382
R8491 x2.x5[7].floating.n168 x2.x5[7].floating.n167 0.0523382
R8492 x2.x5[7].floating.n98 x2.x5[7].floating.n97 0.0516471
R8493 x2.x5[7].floating.n116 x2.x5[7].floating.n115 0.0516471
R8494 x2.x5[7].floating.n134 x2.x5[7].floating.n133 0.0516471
R8495 x2.x5[7].floating.n103 x2.x5[7].floating 0.0495735
R8496 x2.x5[7].floating.n121 x2.x5[7].floating 0.0495735
R8497 x2.x5[7].floating.n139 x2.x5[7].floating 0.0495735
R8498 x2.x5[7].floating.n157 x2.x5[7].floating.n156 0.0408846
R8499 x2.x5[7].floating.n15 x2.x5[7].floating.n14 0.0408846
R8500 x2.x5[7].floating.n75 x2.x5[7].floating.n74 0.0408846
R8501 x2.x5[7].floating.n45 x2.x5[7].floating.n44 0.0408846
R8502 x2.x5[7].floating.n105 x2.x5[7].floating 0.0336765
R8503 x2.x5[7].floating.n123 x2.x5[7].floating 0.0336765
R8504 x2.x5[7].floating x2.x5[7].floating.n171 0.0336765
R8505 x2.x5[7].floating.n60 x2.x5[7].floating.n59 0.0271618
R8506 x2.x5[7].floating.n30 x2.x5[7].floating.n29 0.0271618
R8507 x2.x5[7].floating.n71 x2.x5[7].floating.n70 0.0266618
R8508 x2.x5[7].floating.n41 x2.x5[7].floating.n40 0.0266618
R8509 x2.x5[7].floating.n11 x2.x5[7].floating.n10 0.0266618
R8510 x2.x5[7].floating x2.x5[7].floating.n102 0.0226176
R8511 x2.x5[7].floating x2.x5[7].floating.n104 0.0226176
R8512 x2.x5[7].floating x2.x5[7].floating.n120 0.0226176
R8513 x2.x5[7].floating x2.x5[7].floating.n122 0.0226176
R8514 x2.x5[7].floating x2.x5[7].floating.n138 0.0226176
R8515 x2.x5[7].floating x2.x5[7].floating.n140 0.0226176
R8516 x2.x5[7].floating.n93 x2.x5[7].floating.n92 0.0191618
R8517 x2.x5[7].floating.n111 x2.x5[7].floating.n110 0.0191618
R8518 x2.x5[7].floating.n129 x2.x5[7].floating.n128 0.0191618
R8519 x2.x5[7].floating.n166 x2.x5[7].floating.n165 0.0191618
R8520 x2.x5[7].floating.n96 x2.x5[7].floating.n95 0.0184706
R8521 x2.x5[7].floating.n114 x2.x5[7].floating.n113 0.0184706
R8522 x2.x5[7].floating.n132 x2.x5[7].floating.n131 0.0184706
R8523 x2.x5[7].floating.n163 x2.x5[7].floating.n162 0.0184706
R8524 x2.x5[7].floating.n82 x2.x5[7].floating.n81 0.014
R8525 x2.x5[7].floating.n76 x2.x5[7].floating.n71 0.014
R8526 x2.x5[7].floating.n52 x2.x5[7].floating.n51 0.014
R8527 x2.x5[7].floating.n46 x2.x5[7].floating.n41 0.014
R8528 x2.x5[7].floating.n22 x2.x5[7].floating.n21 0.014
R8529 x2.x5[7].floating.n16 x2.x5[7].floating.n11 0.014
R8530 x2.x5[7].floating.n149 x2.x5[7].floating.n148 0.014
R8531 x2.x5[7].floating.n159 x2.x5[7].floating.n158 0.014
R8532 x2.x5[7].floating.n89 x2.x5[7].floating.n88 0.0135
R8533 x2.x5[7].floating.n79 x2.x5[7].floating.n78 0.0135
R8534 x2.x5[7].floating.n59 x2.x5[7].floating.n58 0.0135
R8535 x2.x5[7].floating.n49 x2.x5[7].floating.n48 0.0135
R8536 x2.x5[7].floating.n29 x2.x5[7].floating.n28 0.0135
R8537 x2.x5[7].floating.n19 x2.x5[7].floating.n18 0.0135
R8538 x2.x5[7].floating.n146 x2.x5[7].floating.n141 0.0135
R8539 x2.x5[7].floating.n152 x2.x5[7].floating.n151 0.0135
R8540 x2.x5[7].floating.n145 x2.x5[7].floating.n144 0.0120385
R8541 x2.x5[7].floating.n27 x2.x5[7].floating.n26 0.0120385
R8542 x2.x5[7].floating.n57 x2.x5[7].floating.n56 0.0120385
R8543 x2.x5[7].floating.n87 x2.x5[7].floating.n86 0.0120385
R8544 x2.x5[7].floating.n97 x2.x5[7].floating.n96 0.00464706
R8545 x2.x5[7].floating.n115 x2.x5[7].floating.n114 0.00464706
R8546 x2.x5[7].floating.n133 x2.x5[7].floating.n132 0.00464706
R8547 x2.x5[7].floating.n162 x2.x5[7].floating.n161 0.00464706
R8548 x2.x5[7].floating.n92 x2.x5[7].floating.n91 0.00395588
R8549 x2.x5[7].floating.n110 x2.x5[7].floating.n109 0.00395588
R8550 x2.x5[7].floating.n128 x2.x5[7].floating.n127 0.00395588
R8551 x2.x5[7].floating.n167 x2.x5[7].floating.n166 0.00395588
R8552 x2.x5[7].floating.n143 x2.x5[7].floating.n142 0.00359614
R8553 x2.x5[7].floating.n25 x2.x5[7].floating.n24 0.00359614
R8554 x2.x5[7].floating.n55 x2.x5[7].floating.n54 0.00359614
R8555 x2.x5[7].floating.n85 x2.x5[7].floating.n84 0.00359614
R8556 x2.x5[7].floating.n88 x2.x5[7].floating.n83 0.0035
R8557 x2.x5[7].floating.n78 x2.x5[7].floating.n77 0.0035
R8558 x2.x5[7].floating.n58 x2.x5[7].floating.n53 0.0035
R8559 x2.x5[7].floating.n48 x2.x5[7].floating.n47 0.0035
R8560 x2.x5[7].floating.n28 x2.x5[7].floating.n23 0.0035
R8561 x2.x5[7].floating.n18 x2.x5[7].floating.n17 0.0035
R8562 x2.x5[7].floating.n147 x2.x5[7].floating.n146 0.0035
R8563 x2.x5[7].floating.n153 x2.x5[7].floating.n152 0.0035
R8564 x2.x5[7].floating.n83 x2.x5[7].floating.n82 0.003
R8565 x2.x5[7].floating.n77 x2.x5[7].floating.n76 0.003
R8566 x2.x5[7].floating.n53 x2.x5[7].floating.n52 0.003
R8567 x2.x5[7].floating.n47 x2.x5[7].floating.n46 0.003
R8568 x2.x5[7].floating.n23 x2.x5[7].floating.n22 0.003
R8569 x2.x5[7].floating.n17 x2.x5[7].floating.n16 0.003
R8570 x2.x5[7].floating.n148 x2.x5[7].floating.n147 0.003
R8571 x2.x5[7].floating.n158 x2.x5[7].floating.n153 0.003
R8572 x2.x5[7].floating.n155 x2.x5[7].floating.n154 0.00277942
R8573 x2.x5[7].floating.n43 x2.x5[7].floating.n42 0.0023396
R8574 x2.x5[7].floating.n13 x2.x5[7].floating.n12 0.0023396
R8575 x2.x5[7].floating.n73 x2.x5[7].floating.n72 0.0023396
R8576 x2.x5[7].floating.n157 x2.x5[7].floating.n155 0.00233747
R8577 x2.x5[7].floating.n15 x2.x5[7].floating.n13 0.00200689
R8578 x2.x5[7].floating.n75 x2.x5[7].floating.n73 0.00200689
R8579 x2.x5[7].floating.n45 x2.x5[7].floating.n43 0.00200689
R8580 x2.x5[7].floating.n145 x2.x5[7].floating.n143 0.0010233
R8581 x2.x5[7].floating.n27 x2.x5[7].floating.n25 0.0010233
R8582 x2.x5[7].floating.n57 x2.x5[7].floating.n55 0.0010233
R8583 x2.x5[7].floating.n87 x2.x5[7].floating.n85 0.0010233
R8584 x2.x5[7].floating.n88 x2.x5[7].floating.n87 0.00053972
R8585 x2.x5[7].floating.n76 x2.x5[7].floating.n75 0.00053972
R8586 x2.x5[7].floating.n58 x2.x5[7].floating.n57 0.00053972
R8587 x2.x5[7].floating.n28 x2.x5[7].floating.n27 0.00053972
R8588 x2.x5[7].floating.n16 x2.x5[7].floating.n15 0.00053972
R8589 x2.x5[7].floating.n146 x2.x5[7].floating.n145 0.00053972
R8590 x2.x5[7].floating.n158 x2.x5[7].floating.n157 0.00053972
R8591 x2.x5[7].floating.n46 x2.x5[7].floating.n45 0.00053972
R8592 sar_logic[7].n2 sar_logic[7].t0 330.616
R8593 sar_logic[7].n0 sar_logic[7].t1 195.121
R8594 sar_logic[7].n3 sar_logic[7] 15.0398
R8595 sar_logic[7].n1 sar_logic[7].n0 14.282
R8596 sar_logic[7].n4 sar_logic[7].n2 8.76429
R8597 sar_logic[7].n3 sar_logic[7] 7.37078
R8598 sar_logic[7] sar_logic[7].n5 2.02977
R8599 sar_logic[7].n2 sar_logic[7].n1 0.893093
R8600 sar_logic[7].n4 sar_logic[7].n3 0.620283
R8601 sar_logic[7].n5 sar_logic[7].n4 0.156598
R8602 delay_code[3].n0 delay_code[3].t0 229.971
R8603 delay_code[3].n0 delay_code[3].t1 158.35
R8604 delay_code[3].n1 delay_code[3].n0 8.50845
R8605 delay_code[3].n1 delay_code[3] 3.95275
R8606 delay_code[3].n2 delay_code[3].n1 1.73287
R8607 delay_code[3].n3 delay_code[3] 0.474765
R8608 delay_code[3] delay_code[3].n3 0.366977
R8609 delay_code[3].n2 delay_code[3] 0.339042
R8610 delay_code[3].n3 delay_code[3].n2 0.00334091
R8611 sar_logic[5].n0 sar_logic[5].t1 329.661
R8612 sar_logic[5].n0 sar_logic[5].t0 209.947
R8613 sar_logic[5].n1 sar_logic[5] 14.9701
R8614 sar_logic[5].n1 sar_logic[5].n0 7.71604
R8615 sar_logic[5] sar_logic[5].n1 1.75049
R8616 delay_code[2] delay_code[2].t1 140.387
R8617 delay_code[2].n1 delay_code[2].t2 140.34
R8618 delay_code[2].n0 delay_code[2].t0 140.34
R8619 delay_code[2].n2 delay_code[2].t3 140.34
R8620 delay_code[2].n3 delay_code[2] 3.93354
R8621 delay_code[2].n2 delay_code[2] 2.82659
R8622 delay_code[2].n1 delay_code[2] 0.285826
R8623 delay_code[2].n2 delay_code[2].n0 0.264087
R8624 delay_code[2].n0 delay_code[2] 0.0466957
R8625 delay_code[2] delay_code[2].n1 0.0466957
R8626 delay_code[2] delay_code[2].n2 0.0371379
R8627 delay_code[2] delay_code[2].n3 0.0306724
R8628 delay_code[2].n3 delay_code[2] 0.0242069
R8629 sar_logic[4].n0 sar_logic[4].t1 331.51
R8630 sar_logic[4].n0 sar_logic[4].t0 209.403
R8631 sar_logic[4] sar_logic[4].n0 79.2785
R8632 sar_logic[4].n1 sar_logic[4] 6.57147
R8633 sar_logic[4].n1 sar_logic[4] 6.4005
R8634 sar_logic[4] sar_logic[4].n1 4.21513
R8635 delay_offset.n2 delay_offset.t1 230.016
R8636 delay_offset.n1 delay_offset.t2 153.665
R8637 delay_offset.n2 delay_offset 153.601
R8638 delay_offset delay_offset.t0 140.379
R8639 delay_offset.n1 delay_offset.n0 73.8234
R8640 delay_offset.n3 delay_offset.n2 9.3005
R8641 delay_offset.n2 delay_offset.n1 4.91671
R8642 delay_offset.n5 delay_offset.n3 4.9013
R8643 delay_offset.n4 delay_offset 4.22092
R8644 delay_offset delay_offset.n0 2.4005
R8645 delay_offset.n7 delay_offset 2.38729
R8646 delay_offset.n4 delay_offset 1.01229
R8647 delay_offset.n5 delay_offset.n4 0.726043
R8648 delay_offset.n3 delay_offset.n0 0.533833
R8649 delay_offset.n6 delay_offset.n5 0.421696
R8650 delay_offset.n7 delay_offset 0.276542
R8651 delay_offset delay_offset.n7 0.2505
R8652 delay_offset.n6 delay_offset 0.0195217
R8653 delay_offset delay_offset.n6 0.0170094
R8654 sar_retimer[7].n0 sar_retimer[7].t1 207.373
R8655 sar_retimer[7].n1 sar_retimer[7] 67.6033
R8656 sar_retimer[7].n1 sar_retimer[7].t0 31.1614
R8657 sar_retimer[7] sar_retimer[7].n0 9.01934
R8658 sar_retimer[7].n0 sar_retimer[7] 7.45876
R8659 sar_retimer[7] sar_retimer[7].n2 3.45135
R8660 sar_retimer[7].n2 sar_retimer[7] 2.07756
R8661 sar_retimer[7].n2 sar_retimer[7].n1 1.22829
R8662 sar_retimer[6].n2 sar_retimer[6].t0 117.424
R8663 sar_retimer[6].n0 sar_retimer[6].t1 75.7697
R8664 sar_retimer[6].n1 sar_retimer[6].n0 73.0808
R8665 sar_retimer[6] sar_retimer[6].n2 66.6967
R8666 sar_retimer[6].n1 sar_retimer[6] 13.7503
R8667 sar_retimer[6].n4 sar_retimer[6].n3 13.0467
R8668 sar_retimer[6].n2 sar_retimer[6] 6.64665
R8669 sar_retimer[6] sar_retimer[6].n1 2.2023
R8670 sar_retimer[6] sar_retimer[6].n4 1.96973
R8671 sar_retimer[6].n3 sar_retimer[6] 1.72358
R8672 sar_retimer[5].n2 sar_retimer[5].t1 425.096
R8673 sar_retimer[5].n3 sar_retimer[5].t1 417.519
R8674 sar_retimer[5].n4 sar_retimer[5].n3 64.2795
R8675 sar_retimer[5].n1 sar_retimer[5].t0 30.6015
R8676 sar_retimer[5] sar_retimer[5].n2 10.0928
R8677 sar_retimer[5].n3 sar_retimer[5] 6.64665
R8678 sar_retimer[5].n2 sar_retimer[5] 6.64665
R8679 sar_retimer[5].n1 sar_retimer[5].n0 4.64234
R8680 sar_retimer[5] sar_retimer[5].n4 2.01398
R8681 sar_retimer[5] sar_retimer[5].n1 0.492808
R8682 sar_retimer[5].n0 sar_retimer[5] 0.373238
R8683 sar_retimer[4].n0 sar_retimer[4].t1 417.519
R8684 sar_retimer[4].n1 sar_retimer[4].t1 136.689
R8685 sar_retimer[4] sar_retimer[4].t0 119.147
R8686 sar_retimer[4].n0 sar_retimer[4] 66.6967
R8687 sar_retimer[4].n2 sar_retimer[4] 12.8551
R8688 sar_retimer[4].n1 sar_retimer[4] 9.84585
R8689 sar_retimer[4] sar_retimer[4].n0 6.64665
R8690 sar_retimer[4] sar_retimer[4].n2 4.56529
R8691 sar_retimer[4].n2 sar_retimer[4].n1 1.2499
R8692 sar_logic[1].n0 sar_logic[1].t0 330.514
R8693 sar_logic[1].n0 sar_logic[1].t1 209.107
R8694 sar_logic[1].n1 sar_logic[1] 14.9981
R8695 sar_logic[1].n1 sar_logic[1].n0 7.74846
R8696 sar_logic[1] sar_logic[1].n1 1.90643
R8697 sar_logic[0].n0 sar_logic[0].t0 331.51
R8698 sar_logic[0].n0 sar_logic[0].t1 209.403
R8699 sar_logic[0] sar_logic[0].n0 79.2785
R8700 sar_logic[0].n1 sar_logic[0] 7.02489
R8701 sar_logic[0].n1 sar_logic[0] 6.54661
R8702 sar_logic[0] sar_logic[0].n1 3.59074
R8703 delay_code[0] delay_code[0].t0 140.343
C0 delay_code[1] a_14312_7267# 2.44e-19
C1 a_16236_5787# sar_retimer[4] 0.0297f
C2 x2.x4[3].floating x3.X 5.28e-19
C3 delay_offset sar_logic[1] 1.65e-21
C4 a_17126_6165# sar_logic[5] 2.69e-20
C5 a_13844_7067# sar_logic[1] 0.0391f
C6 x1[6].Q_N a_16704_5121# 2.97e-20
C7 a_14799_7041# a_15506_7083# 0.0968f
C8 a_14312_7267# a_15789_7073# 2.82e-19
C9 a_13397_5793# a_15789_5793# 0.00176f
C10 a_17017_7445# a_17307_7433# 0.0282f
C11 delay_code[2] a_14625_7445# 6.64e-21
C12 a_15955_6427# a_16875_6709# 1.09e-19
C13 a_16410_6401# a_16654_6709# 0.0104f
C14 sar_retimer[0] sar_retimer[2] 0.0138f
C15 a_14625_6427# a_14711_6793# 0.00976f
C16 a_14312_5121# a_14483_5429# 0.00652f
C17 a_16704_7267# sar_retimer[0] 0.168f
C18 a_13563_5147# a_13952_5147# 0.00116f
C19 a_14018_5121# a_14158_5147# 0.07f
C20 a_16875_7067# a_16410_7041# 9.46e-19
C21 a_14262_6709# a_13563_6427# 2.46e-19
C22 a_13928_6793# a_14018_6401# 6.69e-20
C23 delay_offset a_12385_8002# 1.6e-19
C24 a_14625_5147# a_13397_5793# 5.98e-20
C25 a_17307_5147# sar_logic[7] 7.45e-20
C26 sar_retimer[7] a_15955_5147# 4.16e-20
C27 a_13397_7073# a_14018_7041# 0.117f
C28 sar_logic[0] a_13563_7073# 0.16f
C29 sar_retimer[4] a_14799_5761# 0.00452f
C30 a_16236_5787# x3.X 0.00441f
C31 x2.x3[1].floating x2.x9.output_stack 0.341f
C32 a_13563_6427# a_14018_6401# 0.152f
C33 sar_retimer[6] a_17017_5147# 0.0348f
C34 sar_logic[3] a_16410_6401# 2.88e-19
C35 a_17191_7041# a_16704_6401# 7.68e-20
C36 sar_logic[6] a_13844_5513# 0.0014f
C37 a_12385_8830# x2.x7.floating 8.52e-19
C38 sar_logic[3] sar_logic[2] 0.0778f
C39 sar_retimer[4] a_14711_5787# 8.82e-20
C40 a_13563_5147# a_15506_5147# 7.7e-21
C41 x2.x5[7].floating delay_offset 0.00308f
C42 a_12297_8278# delay_offset 5.57e-19
C43 x2.x5[7].floating a_12410_10219# 0.00154f
C44 x2.x4[3].floating sar_logic[0] 2.28e-19
C45 a_15789_6427# a_13563_6427# 4e-20
C46 a_13397_5147# a_13928_5513# 0.0018f
C47 delay_offset x2.x6.SW 0.19f
C48 x3.A x3.X 0.018f
C49 a_14799_5761# a_14625_6427# 2.23e-20
C50 a_17126_6427# a_16550_6427# 2.46e-21
C51 a_14625_6165# a_14799_6401# 2.23e-20
C52 a_14799_5761# x3.X 0.0152f
C53 a_13397_5147# a_13397_5793# 0.015f
C54 a_14018_5761# a_14018_6401# 0.00923f
C55 a_13844_5787# a_13563_6427# 1.56e-19
C56 sar_logic[3] a_15506_6427# 0.0433f
C57 x2.x4[3].floating x2.x10.Y 0.00668f
C58 a_17017_7445# sar_retimer[2] 1.27e-20
C59 sar_retimer[0] x3.X 0.117f
C60 a_16704_7267# a_17017_7445# 0.119f
C61 a_13844_5513# x3.X 0.00281f
C62 a_17017_6165# a_15955_5147# 8.13e-20
C63 sar_retimer[3] a_17191_6401# 0.00445f
C64 a_15955_7073# a_16410_7041# 0.153f
C65 a_14711_5787# x3.X 2.62e-19
C66 a_17425_5429# sar_retimer[6] 0.00258f
C67 x1[3].Q_N sar_retimer[3] 8.75e-19
C68 a_12297_8830# x2.x10.Y 1.69e-19
C69 a_12457_8692# a_12457_8416# 0.0316f
C70 a_12297_8554# a_12385_8554# 0.00227f
C71 a_12457_8692# x2.x6.floating 0.00278f
C72 a_17191_7041# x2.x3[1].floating 5.96e-19
C73 a_14018_5761# a_13844_5787# 0.205f
C74 a_13563_5793# a_14312_5987# 0.139f
C75 a_15789_5793# a_15955_5147# 1.39e-19
C76 a_14734_6427# a_14625_6427# 0.00707f
C77 a_16410_5121# a_16654_5429# 0.0104f
C78 a_15955_5147# a_16875_5429# 1.09e-19
C79 sar_retimer[7] a_17126_5147# 5e-20
C80 a_14734_6427# x3.X 8.02e-20
C81 a_15033_6709# a_13397_6427# 1.25e-19
C82 a_14312_5121# a_16236_5513# 4.38e-20
C83 a_15033_5429# sar_retimer[6] 1.51e-19
C84 x1[6].Q_N a_15506_5147# 0.178f
C85 a_15955_5793# a_16704_5987# 0.139f
C86 a_16704_5987# a_16704_6401# 0.0107f
C87 x3.A x2.x10.Y 1.17e-19
C88 sar_logic[3] a_14799_6401# 0.0312f
C89 sar_logic[7] a_16410_5121# 2.89e-19
C90 a_15789_5147# a_16236_5513# 0.14f
C91 a_17017_7445# x3.X 9.16e-19
C92 sar_retimer[0] a_16654_7067# 0.00292f
C93 a_12457_8140# x2.x9.output_stack 8.05e-20
C94 a_16143_6427# a_15789_6427# 0.0658f
C95 a_14915_6153# a_14799_5761# 0.0397f
C96 a_13952_6165# sar_logic[5] 0.00178f
C97 x1[4].Q_N a_13563_5793# 2.25e-21
C98 a_14483_5787# a_14018_5761# 9.46e-19
C99 a_14734_6165# a_14625_6165# 0.00707f
C100 sar_logic[5] a_15955_6427# 1.99e-20
C101 x1[7].Q_N a_17017_5147# 9.58e-21
C102 a_13397_5147# a_15955_5147# 2.9e-21
C103 sar_logic[5] a_13397_6427# 1.81e-19
C104 x3.X delay_offset 1.22e-20
C105 a_14530_7389# a_14625_7445# 0.00276f
C106 a_13751_7067# sar_logic[1] 0.0198f
C107 a_14915_7433# a_14312_7267# 0.051f
C108 a_14483_7067# a_13563_7073# 1.09e-19
C109 a_14312_6401# a_14799_7041# 7.68e-20
C110 a_14799_6401# a_14312_7267# 7.68e-20
C111 a_13928_7067# a_13844_7067# 0.00972f
C112 a_14734_7445# a_14799_7041# 4.2e-20
C113 a_14262_7067# a_14018_7041# 0.0104f
C114 sar_retimer[0] a_17191_6401# 1.29e-19
C115 x3.X a_13844_7067# 0.00457f
C116 a_13751_5787# a_13397_5793# 0.0663f
C117 a_16704_5987# x1[5].Q_N 0.00553f
C118 a_13563_6427# a_13563_7073# 0.0099f
C119 a_16550_6153# a_16236_6793# 8.58e-20
C120 a_15955_5793# a_15789_5147# 1.39e-19
C121 a_18195_9356# x3.A 0.148f
C122 a_15789_6427# a_16410_7041# 4.47e-20
C123 a_16550_5147# a_15789_5147# 6.04e-20
C124 delay_code[0] a_13397_7073# 4.1e-19
C125 delay_code[1] a_14625_7445# 8.64e-20
C126 a_17191_5761# sar_retimer[4] 0.0849f
C127 delay_code[2] delay_code[1] 0.553f
C128 a_14625_7445# a_15789_7073# 6.38e-20
C129 a_14799_7041# sar_logic[1] 0.0313f
C130 a_14158_5147# a_14734_5147# 2.46e-21
C131 a_16654_5787# a_15789_5793# 0.00119f
C132 a_16410_5761# sar_retimer[6] 8.16e-20
C133 sar_logic[4] sar_logic[5] 0.0459f
C134 a_16143_7067# a_15789_7073# 0.0657f
C135 a_16704_6401# a_16654_6709# 1.21e-20
C136 a_16143_6427# a_16320_6793# 8.94e-19
C137 a_15955_6427# a_16550_6427# 0.00118f
C138 a_13952_6427# x3.X 1.35e-19
C139 a_15955_5793# a_17103_5787# 2.13e-19
C140 a_14312_6401# a_15033_6709# 0.00185f
C141 a_14625_5147# a_14483_5429# 0.00412f
C142 a_14018_5121# a_14530_5147# 9.75e-19
C143 a_13844_5513# a_13952_5147# 0.00812f
C144 a_14312_5121# a_14158_5147# 0.00943f
C145 a_14799_5121# a_14711_5513# 7.71e-20
C146 a_17425_5429# x1[7].Q_N 2.02e-20
C147 a_17898_6427# a_15789_6427# 1.03e-19
C148 a_13751_5147# sar_logic[4] 3.37e-20
C149 a_14711_6793# a_13563_6427# 2.13e-19
C150 a_14483_6709# a_14018_6401# 9.46e-19
C151 a_17898_5147# a_16704_5121# 6.04e-19
C152 sar_logic[0] a_13844_7067# 0.00105f
C153 x2.x2.floating a_18195_9015# 0.0104f
C154 a_13397_7073# a_14312_7267# 0.125f
C155 sar_retimer[7] a_16236_5513# 1.89e-20
C156 a_16550_7433# delay_code[1] 9.16e-21
C157 sar_retimer[4] a_15506_5803# 0.0744f
C158 a_17191_5761# x3.X 6.15e-19
C159 a_15955_5793# sar_logic[3] 1.99e-20
C160 a_14799_5761# a_15506_5147# 3.56e-19
C161 sar_logic[3] a_16704_6401# 2.8e-19
C162 sar_retimer[6] a_16320_5513# 0.0022f
C163 a_17017_7445# a_17191_6401# 5.77e-20
C164 a_16410_5761# sar_retimer[5] 8.72e-20
C165 a_17191_7041# a_17017_6427# 5.77e-20
C166 a_12410_10219# x2.x10.Y 1.49e-19
C167 delay_offset x2.x10.Y 0.0402f
C168 a_12297_8554# x2.x7.floating 0.00409f
C169 sar_logic[6] a_14799_5121# 1.14e-20
C170 a_16550_7433# a_15789_7073# 6.04e-20
C171 a_14018_5121# sar_retimer[6] 7.99e-20
C172 a_16875_6709# sar_retimer[2] 0.00626f
C173 sar_logic[6] sar_logic[7] 0.05f
C174 a_12385_8278# delay_offset 2.7e-19
C175 sar_retimer[4] sar_logic[7] 1.21e-20
C176 a_13397_5147# a_14483_5429# 0.00907f
C177 sar_logic[5] a_14312_6401# 8.03e-20
C178 a_15506_5803# x3.X 0.0327f
C179 a_16654_5429# x3.X 2.64e-19
C180 a_14312_5987# a_14018_6401# 6.09e-20
C181 x2.x2.floating x2.x9.output_stack 0.193f
C182 a_17191_7041# a_15955_7073# 0.0264f
C183 a_14483_7067# sar_retimer[0] 1.58e-19
C184 a_16550_5147# sar_retimer[7] 8.53e-20
C185 sar_retimer[1] a_15955_7073# 4.55e-20
C186 a_16550_7433# a_17126_7445# 2.46e-21
C187 a_14799_5121# x3.X 0.0111f
C188 a_17425_7067# a_15789_7073# 1.25e-19
C189 a_16704_5987# a_17191_5121# 7.68e-20
C190 a_17191_5761# a_16704_5121# 7.68e-20
C191 a_16410_7041# a_16236_7067# 0.205f
C192 a_16550_6153# x3.X 9.96e-19
C193 a_13397_5793# a_13844_6793# 9.21e-20
C194 sar_logic[7] x3.X 0.0828f
C195 sar_retimer[4] a_17425_5787# 0.00258f
C196 a_16550_6427# a_16922_6427# 3.34e-19
C197 a_15033_5429# x1[6].Q_N 2.02e-20
C198 a_12457_8140# a_12297_8002# 0.0388f
C199 a_16410_5761# a_16143_5787# 6.99e-20
C200 a_12297_8554# a_12297_8278# 0.0316f
C201 x2.x3[1].floating delay_code[0] 0.0429f
C202 a_13563_5793# a_14625_6165# 0.137f
C203 a_13844_5787# a_14312_5987# 0.0633f
C204 a_12297_8554# x2.x6.SW 8.11e-20
C205 a_15789_5793# a_16236_5513# 8.13e-20
C206 a_16875_6709# x3.X 7.12e-20
C207 a_16704_7267# a_14799_7041# 2.71e-20
C208 a_16704_5121# a_16654_5429# 1.21e-20
C209 a_16143_5147# a_16320_5513# 8.94e-19
C210 a_17425_5787# x3.X 5.66e-20
C211 a_14018_5121# a_13844_5787# 1.29e-19
C212 a_13844_5513# a_14018_5761# 1.29e-19
C213 a_14799_5121# a_16704_5121# 3.71e-20
C214 a_15955_5793# a_17017_6165# 0.137f
C215 a_16143_5787# a_14312_5987# 3.27e-20
C216 a_17191_5761# a_17191_6401# 0.0172f
C217 sar_logic[7] a_16704_5121# 2.81e-19
C218 a_15789_5147# a_17191_5121# 0.0492f
C219 sar_logic[3] a_13751_6427# 0.0194f
C220 a_13751_7067# x3.X 0.00446f
C221 a_14158_7433# a_14734_7445# 2.46e-21
C222 a_13751_7067# a_13928_7067# 8.94e-19
C223 a_13563_5147# a_14018_5121# 0.152f
C224 a_17191_5761# x1[3].Q_N 3.57e-19
C225 a_13751_5787# sar_logic[2] 4.77e-20
C226 a_17191_7041# x2.x2.floating 7.24e-19
C227 sar_retimer[0] x1[1].Q_N 0.0258f
C228 a_15955_6427# a_13397_6427# 2.9e-21
C229 a_17898_6427# sar_retimer[3] 0.0749f
C230 x1[2].Q_N a_15506_6427# 0.178f
C231 a_15033_6709# sar_retimer[2] 1.4e-19
C232 a_16143_5787# a_16344_6165# 3.67e-19
C233 a_14483_5787# a_14312_5987# 0.00652f
C234 a_14530_6109# sar_logic[5] 0.00372f
C235 a_15955_5793# a_15789_5793# 0.74f
C236 a_15789_5793# a_16704_6401# 1.07e-20
C237 a_14158_7433# sar_logic[1] 0.0375f
C238 a_14915_7433# a_14625_7445# 0.0282f
C239 a_14799_6401# a_14625_7445# 5.77e-20
C240 a_14262_7067# a_14312_7267# 1.21e-20
C241 a_14625_6427# a_14799_7041# 5.77e-20
C242 x2.x6.floating a_12322_10081# 0.00996f
C243 x3.X a_14799_7041# 0.0162f
C244 a_17017_6165# x1[5].Q_N 9.58e-21
C245 a_14158_6153# a_13397_5793# 6.04e-20
C246 a_14018_6401# a_14018_7041# 0.00947f
C247 a_15955_5793# a_16922_6109# 0.00126f
C248 a_13563_6427# a_13844_7067# 1.14e-19
C249 a_13563_5793# sar_logic[3] 1.45e-19
C250 a_17307_6427# a_16704_6401# 0.0552f
C251 a_16704_7267# a_17103_7067# 3.35e-19
C252 a_16922_5147# a_15789_5147# 2.56e-19
C253 a_16344_5147# sar_logic[7] 3e-19
C254 delay_code[1] a_15789_7073# 2.13e-19
C255 a_13751_7067# sar_logic[0] 0.163f
C256 a_17898_5803# sar_retimer[4] 0.0353f
C257 x1[5].Q_N a_15789_5793# 1.07e-19
C258 a_16704_5987# sar_retimer[6] 6.53e-20
C259 a_15506_7083# sar_logic[1] 0.0438f
C260 a_16344_7445# sar_logic[1] 2.92e-19
C261 a_15033_7067# x3.X 4.06e-19
C262 sar_retimer[0] a_16410_7041# 0.0295f
C263 a_17017_7445# x1[1].Q_N 9.58e-21
C264 a_15955_6427# a_16922_6427# 0.00126f
C265 a_16236_6793# a_16550_6427# 0.0258f
C266 a_16704_6401# a_17103_6793# 3.57e-19
C267 a_15033_6709# x3.X 1.87e-21
C268 a_14799_6401# x1[2].Q_N 0.124f
C269 a_14625_5147# a_14158_5147# 0.00316f
C270 a_14312_5121# a_14530_5147# 3.73e-19
C271 sar_logic[6] sar_logic[5] 5.62e-20
C272 a_13952_6427# a_13563_6427# 0.00116f
C273 a_14158_6427# a_14018_6401# 0.07f
C274 sar_retimer[4] sar_logic[5] 0.044f
C275 a_13952_5147# sar_logic[7] 0.00175f
C276 sar_logic[0] a_14799_7041# 7.83e-21
C277 sar_retimer[7] a_17191_5121# 0.00433f
C278 a_13397_7073# a_14625_7445# 0.0334f
C279 a_14158_6153# a_13844_6793# 8.58e-20
C280 a_16143_7067# a_13397_7073# 3.65e-21
C281 a_15506_5803# a_15506_5147# 0.00419f
C282 delay_code[2] a_13397_7073# 1.8e-19
C283 sar_logic[3] a_17017_6427# 1.22e-19
C284 a_16704_5987# sar_retimer[5] 6.31e-19
C285 a_15955_6427# a_14312_6401# 5.51e-20
C286 sar_logic[6] a_13751_5147# 0.164f
C287 a_12385_8554# x2.x7.floating 8.52e-19
C288 a_16922_7389# sar_logic[1] 1.18e-19
C289 a_12322_10081# a_12322_9805# 0.0316f
C290 a_17103_7067# x3.X 6.95e-20
C291 a_14312_6401# a_13397_6427# 0.126f
C292 a_16143_7067# a_16320_7067# 8.94e-19
C293 a_13844_6793# sar_logic[2] 7.67e-19
C294 a_14799_5121# a_15506_5147# 0.0968f
C295 a_16410_5761# a_16236_5787# 0.205f
C296 a_14312_5121# sar_retimer[6] 3.93e-19
C297 x2.x4[3].floating x2.x9.output_stack 0.636f
C298 a_15506_5147# sar_logic[7] 0.0425f
C299 sar_retimer[6] a_15789_5147# 0.689f
C300 a_13397_5147# a_14158_5147# 6.04e-20
C301 a_13844_5787# a_14158_6427# 8.58e-20
C302 sar_logic[5] a_14625_6427# 2.01e-20
C303 sar_logic[5] x3.X 0.129f
C304 a_18195_9015# x3.A 0.152f
C305 a_16704_5987# a_15789_6427# 1.07e-20
C306 a_16410_6401# a_15789_7073# 4.47e-20
C307 delay_code[0] a_15955_7073# 3.02e-19
C308 a_17017_7445# a_16410_7041# 0.00187f
C309 a_17191_7041# a_16236_7067# 4.7e-22
C310 a_12297_8830# x2.x9.output_stack 0.0388f
C311 a_16236_5787# a_14312_5987# 4.15e-20
C312 sar_retimer[1] a_16236_7067# 2.31e-20
C313 a_13751_5147# x3.X 0.0026f
C314 a_16922_5147# sar_retimer[7] 9.55e-20
C315 a_17017_6165# a_17191_5121# 5.77e-20
C316 a_17191_5761# a_17017_5147# 5.77e-20
C317 a_17126_6165# x3.X 5.56e-20
C318 a_17126_6427# x3.X 5.56e-20
C319 a_12297_8554# x2.x10.Y 6.65e-20
C320 a_16704_5987# a_16143_5787# 3.79e-20
C321 a_16236_5787# a_16344_6165# 0.00812f
C322 a_18499_9105# x2.x5[7].floating 0.00264f
C323 a_14312_7267# a_15955_7073# 5.33e-20
C324 a_12457_8416# x2.x6.floating 0.00167f
C325 a_13563_5793# a_15789_5793# 4e-20
C326 a_14312_5987# a_14799_5761# 0.272f
C327 a_16704_6401# x1[2].Q_N 2.35e-20
C328 a_16704_7267# a_15506_7083# 3.54e-20
C329 x3.A x2.x9.output_stack 0.128f
C330 a_16704_5121# a_17103_5513# 4.23e-19
C331 a_16550_6427# x3.X 9.96e-19
C332 sar_logic[5] sar_logic[0] 4.09e-19
C333 a_14625_5147# a_13563_5793# 8.13e-20
C334 a_13563_5147# a_14625_6165# 8.13e-20
C335 a_14312_5121# a_16143_5147# 3.42e-20
C336 a_14799_5121# a_17017_5147# 1.86e-21
C337 a_17017_6165# a_17017_6427# 0.00421f
C338 a_13563_7073# a_14018_7041# 0.153f
C339 a_17898_5803# a_17191_6401# 3.81e-19
C340 a_14711_5787# a_14312_5987# 0.00133f
C341 a_15955_6427# a_16236_6793# 0.155f
C342 a_15789_5147# a_16143_5147# 0.066f
C343 sar_logic[7] a_17017_5147# 1.22e-19
C344 a_13844_6793# a_14799_6401# 4.7e-22
C345 a_14158_7433# x3.X 9.37e-19
C346 a_14018_5121# a_13844_5513# 0.205f
C347 a_13563_5147# a_14312_5121# 0.139f
C348 a_17898_7083# x2.x2.floating 4.52e-19
C349 x2.x2.floating delay_code[0] 0.164f
C350 x2.x3[1].floating delay_code[2] 0.00115f
C351 sar_logic[3] a_14018_6401# 0.0134f
C352 sar_retimer[7] sar_retimer[6] 0.0478f
C353 a_13563_5147# a_15789_5147# 4e-20
C354 a_16654_6709# a_15789_6427# 0.00119f
C355 a_16704_7267# a_16922_7389# 3.73e-19
C356 x1[4].Q_N a_14799_5761# 0.124f
C357 a_14483_5787# a_14625_6165# 0.00412f
C358 a_14915_6153# sar_logic[5] 0.0397f
C359 x2.x4[3].floating a_14018_7041# 3.7e-20
C360 a_15789_5793# a_17017_6427# 7.69e-20
C361 a_13397_5147# a_13563_5793# 1.39e-19
C362 x3.X a_15506_7083# 0.0333f
C363 x1[0].Q_N a_14312_7267# 0.00553f
C364 a_14734_7445# sar_logic[1] 0.00114f
C365 x2.x6.floating a_12322_9805# 0.00996f
C366 x2.x5[7].floating a_12410_9943# 0.00169f
C367 sar_logic[3] a_15789_6427# 0.269f
C368 a_15955_6427# sar_retimer[2] 0.0229f
C369 a_16344_7445# x3.X 3.03e-19
C370 a_15955_5793# a_13397_5793# 2.9e-21
C371 a_17307_6153# a_16704_6401# 1.41e-19
C372 a_14018_6401# a_14312_7267# 4.94e-20
C373 a_13844_5787# sar_logic[3] 2.64e-20
C374 sar_retimer[2] a_13397_6427# 9.28e-20
C375 a_17307_6427# a_17017_6427# 0.0282f
C376 a_17126_6427# a_17191_6401# 4.2e-20
C377 x1[7].Q_N a_15789_5147# 1.07e-19
C378 a_14530_7389# a_13397_7073# 2.56e-19
C379 a_13844_6793# a_13397_7073# 8.13e-20
C380 x2.x4[3].floating a_12297_8002# 7.17e-20
C381 a_17191_7041# sar_retimer[0] 0.0858f
C382 a_17191_5761# a_17898_6427# 3.81e-19
C383 a_16143_5787# sar_logic[3] 4.77e-20
C384 a_17017_6165# sar_retimer[6] 1.28e-20
C385 sar_retimer[0] sar_retimer[1] 0.0487f
C386 a_14915_6427# a_14734_6427# 4.11e-20
C387 a_17017_6427# a_17103_6793# 0.00976f
C388 a_16922_7389# x3.X 2.71e-19
C389 a_14799_5121# a_15033_5429# 0.00945f
C390 a_13751_5147# a_13952_5147# 3.67e-19
C391 delay_code[1] a_13397_7073# 3.3e-19
C392 a_14625_5147# a_14530_5147# 0.00276f
C393 a_14312_5121# x1[6].Q_N 0.00553f
C394 delay_offset x2.x9.output_stack 0.255f
C395 a_18499_9105# x3.X 0.167f
C396 a_12410_10219# x2.x9.output_stack 1.5e-19
C397 a_14530_6427# a_14018_6401# 9.75e-19
C398 a_12297_8830# a_12385_8968# 0.00227f
C399 a_13397_7073# a_15789_7073# 0.00176f
C400 x1[6].Q_N a_15789_5147# 2.94e-19
C401 a_15789_5793# sar_retimer[6] 1.2e-19
C402 a_13952_6165# x3.X 1.27e-19
C403 sar_retimer[0] a_14018_7041# 7.97e-20
C404 a_17017_6165# sar_retimer[5] 2.27e-19
C405 sar_retimer[6] a_16875_5429# 0.00627f
C406 a_16236_6793# a_14312_6401# 2.6e-20
C407 a_15955_5147# a_16236_5513# 0.155f
C408 a_15955_6427# x3.X 0.013f
C409 a_12297_8278# x2.x7.floating 0.00409f
C410 x2.x5[7].floating x2.x7.floating 0.182f
C411 a_16320_7067# a_15789_7073# 6.02e-19
C412 a_17307_7433# sar_logic[1] 7.07e-20
C413 sar_logic[6] sar_logic[4] 0.00949f
C414 a_14799_6401# sar_logic[2] 2.04e-21
C415 a_13397_6427# x3.X 0.276f
C416 a_14625_6427# a_13397_6427# 0.0334f
C417 x2.x7.floating x2.x6.SW 9.72e-19
C418 a_16236_5787# a_16704_5987# 0.0633f
C419 a_14625_5147# sar_retimer[6] 2.1e-19
C420 sar_retimer[4] a_16320_5787# 0.00223f
C421 a_17191_7041# a_17017_7445# 0.197f
C422 a_13397_5147# a_14530_5147# 2.56e-19
C423 sar_retimer[5] a_15789_5793# 1.24e-19
C424 a_17017_6165# a_15789_6427# 7.69e-20
C425 sar_logic[5] a_13563_6427# 1.51e-19
C426 a_17017_7445# sar_retimer[1] 2.13e-19
C427 delay_code[0] a_16236_7067# 1.2e-19
C428 a_16704_6401# a_15789_7073# 8.63e-20
C429 a_14312_6401# sar_retimer[2] 3.85e-19
C430 a_14799_6401# a_15506_6427# 0.0968f
C431 a_16704_5987# a_14799_5761# 3.59e-20
C432 a_13751_5787# a_13563_5793# 0.158f
C433 x1[7].Q_N sar_retimer[7] 8.13e-19
C434 a_14262_5429# x3.X 3.62e-19
C435 a_16320_5787# x3.X 2.86e-19
C436 a_15955_5793# a_15955_5147# 0.0099f
C437 sar_logic[4] x3.X 0.0765f
C438 a_16922_6109# sar_retimer[5] 9.99e-20
C439 a_16550_5147# a_15955_5147# 0.00118f
C440 a_13397_5147# sar_retimer[6] 9.32e-20
C441 a_18499_9105# x2.x10.Y 2.48e-19
C442 delay_code[0] a_13563_7073# 3.02e-19
C443 a_15789_5793# a_15789_6427# 0.0151f
C444 a_16410_5761# a_16550_6153# 0.07f
C445 a_13397_6427# sar_logic[0] 3.23e-21
C446 a_12457_8416# a_12385_8416# 0.00227f
C447 a_16236_5787# a_15789_5147# 8.13e-20
C448 a_14312_7267# a_16236_7067# 2.51e-20
C449 a_14312_5987# a_15506_5803# 6.04e-19
C450 a_14018_5761# sar_logic[5] 0.0137f
C451 sar_retimer[2] sar_logic[1] 1.21e-20
C452 a_14799_5761# a_14625_6165# 0.197f
C453 delay_offset a_12322_10357# 3.28e-19
C454 a_12297_8278# x2.x6.SW 4.74e-20
C455 a_16143_7067# a_15955_7073# 0.158f
C456 a_12410_10219# a_12322_10357# 0.0704f
C457 a_14915_5147# a_14734_5147# 4.11e-20
C458 a_16704_7267# sar_logic[1] 2.76e-19
C459 a_17017_5147# a_17103_5513# 0.00976f
C460 a_16922_6427# x3.X 2.45e-19
C461 a_14734_6427# a_14158_6427# 2.46e-21
C462 x2.x5[7].floating x2.x6.SW 0.00138f
C463 a_14799_5121# a_14312_5987# 7.68e-20
C464 a_13751_5787# a_13928_5787# 8.94e-19
C465 x2.x4[3].floating delay_code[0] 8.57e-20
C466 a_14158_6153# a_14734_6165# 2.46e-21
C467 x2.x3[1].floating delay_code[1] 0.227f
C468 a_14312_5121# a_14799_5761# 7.68e-20
C469 a_14312_5121# a_14915_5147# 0.0511f
C470 a_17307_5147# a_16704_5121# 0.0552f
C471 a_13563_7073# a_14312_7267# 0.139f
C472 a_15033_5787# a_14799_5761# 0.00945f
C473 a_14711_5787# a_14625_6165# 0.00976f
C474 a_13397_5793# a_13563_5793# 0.744f
C475 a_14018_7041# a_13844_7067# 0.205f
C476 a_16143_5787# a_15789_5793# 0.0658f
C477 a_15955_5793# a_16410_6401# 2.37e-20
C478 a_15955_6427# a_17191_6401# 0.0264f
C479 a_16410_6401# a_16704_6401# 0.199f
C480 a_14312_6401# x3.X 0.00505f
C481 a_14734_7445# x3.X 7.88e-20
C482 a_13844_6793# a_13751_6427# 0.0367f
C483 a_14312_6401# a_14625_6427# 0.124f
C484 x2.x3[1].floating a_15789_7073# 7.89e-19
C485 a_13844_5513# a_14312_5121# 0.0633f
C486 a_13563_5147# a_14625_5147# 0.137f
C487 a_16550_7433# a_15955_7073# 0.00118f
C488 x1[3].Q_N a_15955_6427# 4.18e-21
C489 a_18195_9356# a_18499_9105# 0.0406f
C490 a_14018_5121# sar_logic[7] 0.0134f
C491 a_16704_7267# a_17307_7433# 0.055f
C492 sar_retimer[4] a_16410_5121# 8.65e-20
C493 x1[4].Q_N a_15506_5803# 0.178f
C494 x2.x4[3].floating a_14312_7267# 4.99e-19
C495 x3.X x2.x7.floating 9.09e-19
C496 sar_logic[5] a_16143_6427# 4.77e-20
C497 a_12410_9943# x2.x10.Y 4.2e-19
C498 a_14711_7067# a_13563_7073# 2.13e-19
C499 a_13397_5147# a_13844_5787# 8.13e-20
C500 delay_offset a_12297_8002# 2.98e-19
C501 a_13397_5147# a_16143_5147# 3.65e-21
C502 x3.X sar_logic[1] 0.125f
C503 x1[0].Q_N a_14625_7445# 9.58e-21
C504 x1[4].Q_N a_14799_5121# 3.56e-19
C505 a_12385_8968# delay_offset 9.08e-19
C506 a_16236_6793# sar_retimer[2] 0.0297f
C507 a_16704_6401# a_15506_6427# 3.66e-20
C508 a_13928_5787# a_13397_5793# 0.0018f
C509 a_17307_6153# a_17017_6427# 6.09e-20
C510 a_16550_5147# a_17126_5147# 2.46e-21
C511 x1[0].Q_N delay_code[2] 7.35e-21
C512 a_15955_5793# a_16654_5787# 2.46e-19
C513 a_14799_5761# sar_logic[3] 8.24e-20
C514 x3.A delay_code[0] 4.31e-19
C515 a_13397_5147# a_13563_5147# 0.746f
C516 a_13563_5793# a_13844_6793# 1.56e-19
C517 a_16410_5121# x3.X 0.00214f
C518 sar_retimer[0] sar_logic[3] 1.21e-20
C519 a_17898_5803# a_17898_6427# 0.00442f
C520 a_17898_7083# sar_retimer[0] 0.0356f
C521 x2.x4[3].floating a_12457_8692# 8.29e-19
C522 a_17307_7433# x3.X 2.12e-19
C523 a_16704_7267# sar_retimer[2] 7.44e-20
C524 a_14625_5147# x1[6].Q_N 9.58e-21
C525 x2.x5[7].floating x3.X 8.06e-19
C526 sar_logic[0] sar_logic[1] 0.0457f
C527 a_12297_8830# a_12457_8692# 0.0388f
C528 x2.x7.floating x2.x10.Y 0.00345f
C529 sar_retimer[0] a_14312_7267# 3.94e-19
C530 a_14530_6109# x3.X 3.45e-19
C531 a_14915_6153# a_14312_6401# 1.41e-19
C532 a_16704_6401# a_14799_6401# 2.76e-20
C533 a_16410_5121# a_16704_5121# 0.199f
C534 sar_logic[3] a_14734_6427# 0.00113f
C535 a_15955_5147# a_17191_5121# 0.0264f
C536 a_16236_6793# x3.X 0.0044f
C537 a_16875_7067# a_15789_7073# 0.00571f
C538 a_12385_8278# x2.x7.floating 8.52e-19
C539 a_13928_6793# a_13397_6427# 0.0018f
C540 a_13751_6427# sar_logic[2] 0.163f
C541 a_17898_5147# a_15789_5147# 1.03e-19
C542 sar_retimer[4] a_16875_5787# 0.00626f
C543 a_16704_5987# a_17191_5761# 0.27f
C544 x1[2].Q_N a_15789_6427# 2.94e-19
C545 sar_retimer[3] a_17307_6427# 5.08e-19
C546 a_13397_6427# a_13563_6427# 0.749f
C547 a_17017_7445# delay_code[0] 1.08e-19
C548 a_13397_5147# x1[6].Q_N 1.07e-19
C549 sar_retimer[0] a_14711_7067# 8.75e-20
C550 a_17017_6427# a_15789_7073# 5.98e-20
C551 a_14625_6427# sar_retimer[2] 1.96e-19
C552 a_17017_6165# a_14799_5761# 1.86e-21
C553 a_12457_8140# a_12385_8140# 0.00227f
C554 a_16410_5761# sar_logic[5] 2.98e-19
C555 a_16236_5787# a_15789_5793# 0.14f
C556 sar_retimer[2] x3.X 0.117f
C557 a_14158_6153# a_13563_5793# 0.00118f
C558 a_16704_5987# a_15506_5803# 5.37e-20
C559 a_13751_5787# a_13844_5787# 0.0367f
C560 a_15955_5793# a_16236_5513# 1.14e-19
C561 a_16704_7267# x3.X 0.00204f
C562 a_16875_5787# x3.X 3.98e-19
C563 a_17307_6153# sar_retimer[5] 5.43e-19
C564 a_16550_5147# a_16236_5513# 0.0258f
C565 a_16922_5147# a_15955_5147# 0.00126f
C566 delay_code[0] delay_offset 1.92e-20
C567 a_12297_8278# x2.x10.Y 4.07e-20
C568 a_13952_7445# a_13563_7073# 0.00114f
C569 delay_code[0] a_13844_7067# 1.2e-19
C570 x2.x5[7].floating x2.x10.Y 1.01f
C571 a_13563_5793# sar_logic[2] 1.99e-20
C572 sar_logic[4] a_13563_6427# 1.99e-20
C573 a_13751_7067# a_14018_7041# 6.99e-20
C574 delay_code[1] a_15955_7073# 1.32e-19
C575 a_16704_5987# a_16550_6153# 0.00943f
C576 x2.x10.Y x2.x6.SW 0.788f
C577 a_12457_8140# x2.x6.floating 0.00109f
C578 sar_logic[6] x3.X 0.0799f
C579 a_12297_8278# a_12385_8278# 0.00227f
C580 a_12457_8416# a_12457_8140# 0.0316f
C581 a_15789_7073# a_15955_7073# 0.742f
C582 sar_retimer[4] x3.X 0.117f
C583 a_14799_5761# a_15789_5793# 0.00116f
C584 a_14312_5987# sar_logic[5] 0.0863f
C585 a_16143_7067# a_16236_7067# 0.0367f
C586 a_14799_5121# a_14625_6165# 5.77e-20
C587 a_14625_5147# a_14799_5761# 5.77e-20
C588 a_17126_5147# a_17191_5121# 4.2e-20
C589 a_17307_5147# a_17017_5147# 0.0282f
C590 a_14625_5147# a_14915_5147# 0.0282f
C591 a_14799_5121# a_14734_5147# 4.2e-20
C592 a_16344_6165# sar_logic[5] 3.12e-19
C593 sar_logic[4] a_14018_5761# 6.04e-19
C594 a_13397_5793# a_13844_5787# 0.15f
C595 a_13563_7073# a_14625_7445# 0.137f
C596 a_13844_7067# a_14312_7267# 0.0633f
C597 a_15955_5793# a_16704_6401# 1.45e-20
C598 a_15789_5147# a_16654_5429# 0.00126f
C599 a_16410_6401# a_17017_6427# 0.00187f
C600 a_15955_6427# a_16143_6427# 0.158f
C601 delay_code[2] a_13563_7073# 1.15e-19
C602 a_16236_6793# a_17191_6401# 4.7e-22
C603 sar_logic[7] a_14734_5147# 0.00113f
C604 sar_logic[3] a_13952_6427# 0.00175f
C605 a_17191_5761# a_17103_5787# 7.71e-20
C606 a_14625_6427# x3.X 6.62e-19
C607 a_17898_5147# sar_retimer[7] 0.0747f
C608 a_13928_7067# x3.X 4.41e-19
C609 a_16704_5987# a_17425_5787# 7.95e-19
C610 a_14018_5121# a_13751_5147# 6.99e-20
C611 a_14312_5121# a_14799_5121# 0.272f
C612 a_13563_5147# a_13928_5513# 4.45e-20
C613 a_16922_7389# a_16410_7041# 9.75e-19
C614 a_16550_7433# a_16236_7067# 0.0258f
C615 a_17425_6709# a_16704_6401# 7.95e-19
C616 a_16143_6427# a_13397_6427# 3.65e-21
C617 a_18195_9356# x2.x5[7].floating 0.0132f
C618 a_13563_5147# a_13397_5793# 1.39e-19
C619 a_13844_6793# a_14018_6401# 0.205f
C620 a_14312_6401# a_13563_6427# 0.139f
C621 a_14799_5121# a_15789_5147# 0.00116f
C622 a_14312_5121# sar_logic[7] 0.0879f
C623 a_16143_5787# a_13397_5793# 3.65e-21
C624 a_16704_7267# a_16654_7067# 1.21e-20
C625 sar_retimer[4] a_16704_5121# 7.44e-20
C626 x1[4].Q_N sar_logic[5] 0.0243f
C627 sar_retimer[6] a_15955_5147# 0.0224f
C628 a_15789_5147# sar_logic[7] 0.27f
C629 x2.x4[3].floating a_14625_7445# 4.05e-21
C630 x2.x4[3].floating delay_code[2] 0.532f
C631 x2.x2.floating delay_code[1] 0.0027f
C632 a_17191_7041# a_17103_7067# 7.71e-20
C633 x1[0].Q_N a_15789_7073# 2.94e-19
C634 a_12457_8692# delay_offset 0.00297f
C635 a_17191_6401# sar_retimer[2] 0.0849f
C636 a_14483_5787# a_13397_5793# 0.00907f
C637 a_14262_5787# sar_logic[4] 8.37e-22
C638 a_16704_7267# a_17191_6401# 7.68e-20
C639 a_15955_5793# x1[5].Q_N 1.68e-21
C640 x1[3].Q_N sar_retimer[2] 0.0257f
C641 a_13397_5147# a_13844_5513# 0.15f
C642 a_15506_5803# sar_logic[3] 9.57e-21
C643 a_13844_5787# a_13844_6793# 0.00451f
C644 a_14018_5761# a_14312_6401# 6.09e-20
C645 a_16704_5121# x3.X 8.07e-19
C646 a_14262_7067# a_13397_7073# 0.00276f
C647 x3.X sar_logic[0] 0.0782f
C648 a_17898_6427# a_15955_6427# 7.7e-21
C649 a_15789_6427# a_15789_7073# 0.015f
C650 a_16654_7067# x3.X 2.64e-19
C651 x3.X x2.x10.Y 1.41e-20
C652 a_18195_9015# a_18499_9105# 0.0314f
C653 a_12385_8830# a_12457_8692# 0.00227f
C654 sar_retimer[0] a_14625_7445# 2.15e-19
C655 a_14915_6153# x3.X 0.00113f
C656 a_14915_6153# a_14625_6427# 6.09e-20
C657 a_16143_6427# a_14312_6401# 2.23e-20
C658 a_17017_6427# a_14799_6401# 1.86e-21
C659 a_16236_5513# a_17191_5121# 4.7e-22
C660 a_15955_5147# a_16143_5147# 0.158f
C661 a_16410_5121# a_17017_5147# 0.00187f
C662 sar_retimer[0] a_16143_7067# 0.0142f
C663 a_17191_6401# x3.X 1e-19
C664 a_14483_6709# a_13397_6427# 0.00907f
C665 a_17191_5761# a_17017_6165# 0.197f
C666 a_14483_5429# sar_retimer[6] 1.58e-19
C667 a_16704_5987# a_17898_5803# 6.04e-19
C668 sar_logic[2] a_14018_6401# 8.01e-20
C669 a_16410_5761# a_15955_6427# 2.37e-20
C670 a_14799_5761# x1[2].Q_N 3.57e-19
C671 a_18195_9356# x3.X 0.0021f
C672 a_16143_6427# sar_logic[1] 3.37e-20
C673 a_18499_9105# x2.x9.output_stack 5.27e-19
C674 a_16410_6401# a_15789_6427# 0.111f
C675 a_14530_6109# a_14018_5761# 9.75e-19
C676 a_14158_6153# a_13844_5787# 0.0258f
C677 a_16704_5987# sar_logic[5] 2.9e-19
C678 a_17191_5761# a_15789_5793# 0.0492f
C679 sar_retimer[2] a_13563_6427# 3.91e-20
C680 x1[7].Q_N a_15955_5147# 4.5e-21
C681 a_13952_7445# a_13844_7067# 0.00812f
C682 a_13751_7067# a_14312_7267# 4.94e-21
C683 delay_code[0] a_14799_7041# 5.05e-19
C684 a_14530_7389# a_13563_7073# 0.00126f
C685 a_13844_6793# a_13563_7073# 1.14e-19
C686 delay_code[1] a_16236_7067# 3.77e-19
C687 a_14312_5987# a_13397_6427# 1.07e-20
C688 a_14158_7433# a_14018_7041# 0.07f
C689 a_16704_5987# a_17126_6165# 2.87e-21
C690 a_17017_6165# a_16550_6153# 0.00316f
C691 a_16410_5761# a_16320_5787# 6.69e-20
C692 a_15789_7073# a_16236_7067# 0.14f
C693 sar_logic[1] a_16410_7041# 2.83e-19
C694 a_14625_6165# sar_logic[5] 0.0363f
C695 a_15506_5803# a_15789_5793# 8.18e-19
C696 sar_retimer[0] a_17425_7067# 0.00259f
C697 a_15506_5147# x3.X 0.0296f
C698 a_15506_6427# a_15789_6427# 8.18e-19
C699 delay_code[1] a_13563_7073# 2.43e-19
C700 a_13563_7073# a_15789_7073# 4e-20
C701 a_14312_7267# a_14799_7041# 0.272f
C702 a_13397_7073# a_15955_7073# 2.9e-21
C703 a_16550_6153# a_15789_5793# 6.04e-20
C704 a_13397_5793# a_14799_5761# 0.0492f
C705 a_16704_5987# a_16550_6427# 1.58e-19
C706 sar_logic[4] a_14312_5987# 0.00305f
C707 a_17017_7445# a_16550_7433# 0.00316f
C708 delay_code[2] delay_offset 0.0105f
C709 a_15955_5793# a_17017_6427# 9.03e-20
C710 x1[5].Q_N a_17191_5121# 3.56e-19
C711 a_16704_6401# a_17017_6427# 0.12f
C712 a_18195_9356# x2.x10.Y 0.00127f
C713 a_16410_6401# a_16320_6793# 6.69e-20
C714 a_16236_6793# a_16143_6427# 0.0367f
C715 delay_code[2] a_13844_7067# 0.00111f
C716 x1[0].Q_N a_14799_6401# 3.56e-19
C717 a_13928_6793# x3.X 4.41e-19
C718 a_14312_6401# a_14483_6709# 0.00652f
C719 a_14483_7067# x3.X 9.28e-19
C720 a_14312_5121# a_13751_5147# 5.76e-21
C721 a_16550_5147# a_16922_5147# 3.34e-19
C722 a_13844_5513# a_13928_5513# 0.00972f
C723 a_13563_5147# a_14483_5429# 1.09e-19
C724 a_12410_9943# x2.x9.output_stack 0.032f
C725 a_14799_5121# a_14625_5147# 0.197f
C726 a_16922_7389# sar_retimer[1] 9.46e-20
C727 a_14018_5121# a_14262_5429# 0.0104f
C728 a_16320_7067# a_15955_7073# 4.45e-20
C729 x1[3].Q_N a_17191_6401# 0.124f
C730 a_13563_6427# x3.X 0.0148f
C731 x2.x4[3].floating delay_code[1] 0.0307f
C732 a_14625_6427# a_13563_6427# 0.137f
C733 a_13844_5513# a_13397_5793# 8.13e-20
C734 a_16550_6153# a_16922_6109# 3.34e-19
C735 a_14625_5147# sar_logic[7] 0.0362f
C736 sar_retimer[4] a_14018_5761# 7.8e-20
C737 a_16704_7267# x1[1].Q_N 0.00553f
C738 sar_retimer[4] a_17017_5147# 1.27e-20
C739 x2.x4[3].floating a_15789_7073# 2.59e-19
C740 sar_retimer[6] a_16236_5513# 0.0292f
C741 a_15506_5147# a_16704_5121# 5.62e-20
C742 a_17425_5787# a_15789_5793# 1.25e-19
C743 a_15033_7067# a_14312_7267# 0.00185f
C744 a_14711_7067# a_14799_7041# 7.71e-20
C745 a_16236_6793# a_16410_7041# 1.29e-19
C746 a_16410_6401# a_16236_7067# 1.29e-19
C747 a_14799_6401# a_15789_6427# 0.00116f
C748 a_16143_6427# sar_retimer[2] 0.0139f
C749 a_12385_8692# delay_offset 6.22e-19
C750 a_13397_5147# a_14799_5121# 0.0492f
C751 a_14312_5987# a_14312_6401# 0.0107f
C752 sar_logic[5] sar_logic[3] 0.0128f
C753 a_14018_5761# x3.X 0.0028f
C754 a_17017_5147# x3.X 1.4e-20
C755 a_13397_5147# sar_logic[7] 0.0426f
C756 x1[0].Q_N a_13397_7073# 1.07e-19
C757 a_14483_7067# sar_logic[0] 1.46e-21
C758 a_14262_5787# sar_retimer[4] 5.09e-20
C759 a_13397_6427# a_14018_7041# 4.47e-20
C760 a_14018_6401# a_13397_7073# 4.47e-20
C761 a_15955_5793# sar_retimer[6] 8.71e-20
C762 a_16410_5761# a_16410_5121# 0.00947f
C763 x3.A delay_code[1] 5.47e-22
C764 sar_retimer[3] a_16410_6401# 8.19e-20
C765 a_16236_5787# a_15955_5147# 1.14e-19
C766 a_17126_6427# sar_logic[3] 2.66e-20
C767 sar_retimer[2] a_16410_7041# 8.65e-20
C768 x2.x4[3].floating a_12457_8416# 8.29e-19
C769 x2.x7.floating x2.x9.output_stack 0.185f
C770 a_16704_7267# a_16410_7041# 0.199f
C771 a_14158_5147# a_14530_5147# 3.34e-19
C772 a_12457_8692# a_12297_8554# 0.0388f
C773 a_14262_5787# x3.X 4.92e-19
C774 sar_retimer[0] a_15789_7073# 0.715f
C775 a_16704_5121# a_17017_5147# 0.12f
C776 a_14915_6427# a_14312_6401# 0.0511f
C777 a_16236_5513# a_16143_5147# 0.0367f
C778 sar_logic[3] a_16550_6427# 3.51e-19
C779 a_16410_5121# a_16320_5513# 6.69e-20
C780 a_16143_6427# x3.X 0.00503f
C781 x2.x3[1].floating a_15955_7073# 3.31e-19
C782 a_15955_5793# sar_retimer[5] 5e-20
C783 a_12322_10081# delay_offset 6.38e-19
C784 a_17898_6427# sar_retimer[2] 0.0354f
C785 a_12410_10219# a_12322_10081# 0.0704f
C786 a_14158_6427# a_13397_6427# 6.04e-20
C787 a_16704_5987# a_15955_6427# 1.45e-20
C788 a_16236_5787# a_16410_6401# 3.66e-20
C789 a_16410_5761# a_16236_6793# 3.66e-20
C790 a_13751_7067# a_13952_7445# 3.67e-19
C791 x2.x5[7].floating x2.x9.output_stack 1.19f
C792 x3.X a_16410_7041# 0.00295f
C793 a_15955_5793# a_15789_6427# 4.5e-20
C794 a_16704_6401# a_15789_6427# 0.124f
C795 a_14483_6709# sar_retimer[2] 1.5e-19
C796 a_17898_5803# a_15789_5793# 1.03e-19
C797 a_14530_6109# a_14312_5987# 3.73e-19
C798 a_13928_5787# a_13563_5793# 4.45e-20
C799 a_17017_6165# sar_logic[5] 1.28e-19
C800 x2.x6.SW x2.x9.output_stack 0.164f
C801 a_17425_6709# a_15789_6427# 1.25e-19
C802 x1[5].Q_N sar_retimer[5] 9.81e-19
C803 a_17425_5429# a_16704_5121# 8.46e-19
C804 a_14625_6165# a_13397_6427# 7.69e-20
C805 a_17191_7041# sar_logic[1] 7.3e-20
C806 a_14312_6401# a_14018_7041# 4.94e-20
C807 a_14158_7433# a_14312_7267# 0.00943f
C808 a_17017_7445# a_15789_7073# 0.0322f
C809 delay_code[0] a_15506_7083# 1.16e-19
C810 a_13844_6793# a_13844_7067# 0.00445f
C811 sar_retimer[0] a_16410_6401# 8.82e-20
C812 a_17191_5761# a_17307_6153# 0.0397f
C813 a_16410_5761# a_16875_5787# 9.46e-19
C814 a_17017_6165# a_17126_6165# 0.00707f
C815 a_15955_5793# a_16143_5787# 0.158f
C816 a_15789_5793# sar_logic[5] 0.266f
C817 a_17191_6401# x1[1].Q_N 3.56e-19
C818 x2.x3[1].floating x2.x2.floating 1.17f
C819 delay_code[1] delay_offset 2.09e-20
C820 delay_code[1] a_13844_7067# 9.67e-20
C821 a_16410_5761# sar_retimer[4] 0.0293f
C822 a_14799_5761# a_15506_6427# 3.81e-19
C823 a_14312_7267# a_15506_7083# 6.04e-19
C824 a_14018_7041# sar_logic[1] 0.0137f
C825 a_16922_6109# sar_logic[5] 1.23e-19
C826 a_14799_7041# a_14625_7445# 0.197f
C827 sar_logic[4] a_14625_6165# 4.67e-20
C828 a_13397_5793# a_15506_5803# 1.03e-19
C829 a_16143_7067# a_14799_7041# 8.26e-21
C830 a_17017_7445# a_17126_7445# 0.00707f
C831 a_17191_7041# a_17307_7433# 0.0397f
C832 a_15955_6427# a_16654_6709# 2.46e-19
C833 delay_code[2] a_14799_7041# 1.33e-20
C834 a_14483_6709# x3.X 1.5e-19
C835 a_13844_6793# a_13952_6427# 0.00812f
C836 a_17307_7433# sar_retimer[1] 4.85e-19
C837 a_14799_6401# a_14711_6793# 7.71e-20
C838 a_14625_6427# a_14483_6709# 0.00412f
C839 a_14312_6401# a_14158_6427# 0.00943f
C840 a_14312_5121# a_14262_5429# 1.21e-20
C841 a_13563_5147# a_14158_5147# 0.00118f
C842 a_18195_9015# x3.X 0.0163f
C843 a_16320_7067# a_16236_7067# 0.00972f
C844 a_18499_9105# delay_code[0] 1.68e-19
C845 a_16654_7067# a_16410_7041# 0.0104f
C846 a_16875_7067# a_15955_7073# 1.09e-19
C847 a_13751_6427# a_14018_6401# 6.99e-20
C848 delay_offset a_12385_8140# 2.1e-19
C849 a_13928_6793# a_13563_6427# 4.45e-20
C850 a_17898_5147# a_15955_5147# 8.33e-21
C851 a_13397_7073# a_13563_7073# 0.747f
C852 sar_retimer[4] a_14312_5987# 3.88e-19
C853 a_17307_6427# a_17126_6427# 4.11e-20
C854 a_16410_5761# x3.X 0.0027f
C855 x2.x7.floating a_12297_8002# 0.00218f
C856 sar_logic[3] a_15955_6427# 0.249f
C857 sar_retimer[6] a_17191_5121# 0.0824f
C858 x2.x5[7].floating a_12322_10357# 2.14e-19
C859 sar_logic[6] a_14018_5121# 5.73e-19
C860 a_12385_8968# x2.x7.floating 8.52e-19
C861 sar_logic[3] a_13397_6427# 0.04f
C862 x2.x6.SW a_12322_10357# 5.11e-20
C863 a_17017_6427# a_15955_7073# 8.13e-20
C864 x1[2].Q_N a_14799_7041# 3.56e-19
C865 x2.x6.floating delay_offset 0.0624f
C866 a_12457_8416# delay_offset 8.34e-19
C867 x2.x6.floating a_12410_10219# 0.0191f
C868 x2.x4[3].floating a_13397_7073# 5.64e-19
C869 a_13397_5147# a_13751_5147# 0.0669f
C870 a_14799_5761# a_14799_6401# 0.0172f
C871 a_14312_5987# x3.X 0.00416f
C872 a_16320_5513# x3.X 3.02e-19
C873 x3.X x2.x9.output_stack 0.00468f
C874 a_12297_8002# a_12385_8002# 0.0022f
C875 a_14018_5761# a_13563_6427# 2.37e-20
C876 a_13563_5793# a_14018_6401# 2.37e-20
C877 a_17191_7041# sar_retimer[2] 1.27e-19
C878 x1[4].Q_N sar_retimer[4] 7.76e-19
C879 a_14018_5121# x3.X 0.00223f
C880 a_16704_7267# a_17191_7041# 0.27f
C881 a_13397_6427# a_14312_7267# 8.63e-20
C882 a_16236_5787# a_16236_5513# 0.00445f
C883 a_16410_5761# a_16704_5121# 4.94e-20
C884 sar_retimer[3] a_16704_6401# 6.06e-19
C885 sar_logic[4] sar_logic[3] 2.96e-20
C886 a_16704_5987# a_16410_5121# 4.94e-20
C887 a_17898_6427# a_17191_6401# 0.0968f
C888 a_16344_6165# x3.X 3.03e-19
C889 a_16704_7267# sar_retimer[1] 5.85e-19
C890 x1[3].Q_N a_17898_6427# 0.178f
C891 a_15033_6709# x1[2].Q_N 2.02e-20
C892 a_12297_8278# a_12297_8002# 0.0316f
C893 a_12297_8554# a_12385_8692# 0.00227f
C894 x2.x6.SW a_12297_8002# 3.1e-20
C895 a_13563_5793# a_13844_5787# 0.146f
C896 sar_logic[3] a_16922_6427# 1.17e-19
C897 x1[4].Q_N x3.X 0.00411f
C898 a_15955_5147# a_16654_5429# 2.46e-19
C899 a_14734_6427# a_14799_6401# 4.2e-20
C900 a_14915_6427# a_14625_6427# 0.0282f
C901 a_14915_6427# x3.X 0.00112f
C902 x2.x3[1].floating a_16236_7067# 7.62e-21
C903 sar_retimer[7] a_17307_5147# 4.56e-19
C904 a_12322_9805# delay_offset 0.00273f
C905 a_14530_6427# a_13397_6427# 2.56e-19
C906 a_13563_5147# a_13563_5793# 0.0099f
C907 a_14312_5121# a_16410_5121# 4.53e-20
C908 a_14799_5121# a_15955_5147# 2.24e-20
C909 a_15955_5793# a_16236_5787# 0.155f
C910 a_17017_6165# a_15955_6427# 9.03e-20
C911 sar_retimer[0] a_13397_7073# 9.26e-20
C912 sar_logic[3] a_14312_6401# 0.0879f
C913 a_15789_5147# a_16410_5121# 0.111f
C914 sar_logic[7] a_15955_5147# 0.25f
C915 x2.x10.Y x2.x9.output_stack 1.01f
C916 a_17191_7041# x3.X 0.0015f
C917 sar_retimer[0] a_16320_7067# 0.00224f
C918 a_18195_9015# a_18195_9356# 0.0121f
C919 sar_retimer[1] x3.X 0.0175f
C920 a_17017_6427# a_15789_6427# 0.0322f
C921 a_14262_5787# a_14018_5761# 0.0104f
C922 a_13928_5787# a_13844_5787# 0.00972f
C923 a_14734_6165# a_14799_5761# 4.2e-20
C924 a_13751_5787# sar_logic[5] 0.0198f
C925 a_14483_5787# a_13563_5793# 1.09e-19
C926 a_14915_6153# a_14312_5987# 0.051f
C927 a_14530_6109# a_14625_6165# 0.00276f
C928 a_15955_5793# a_14799_5761# 2.24e-20
C929 delay_code[0] x2.x7.floating 1.4e-20
C930 a_15789_5793# a_15955_6427# 4.5e-20
C931 x1[7].Q_N a_17191_5121# 0.124f
C932 x2.x4[3].floating x2.x3[1].floating 1.19f
C933 sar_logic[3] sar_logic[1] 0.0041f
C934 a_13928_7067# a_14018_7041# 6.69e-20
C935 a_14262_7067# a_13563_7073# 2.46e-19
C936 a_14312_6401# a_14312_7267# 0.0106f
C937 a_14734_7445# a_14312_7267# 2.87e-21
C938 a_14158_7433# a_14625_7445# 0.00316f
C939 delay_code[0] sar_logic[1] 1.1e-19
C940 sar_retimer[0] a_16704_6401# 7.74e-20
C941 x3.X a_14018_7041# 0.0034f
C942 a_16704_5987# a_16875_5787# 0.00652f
C943 a_14158_7433# delay_code[2] 4.56e-21
C944 a_15789_6427# a_15955_7073# 1.39e-19
C945 a_18195_9356# x2.x9.output_stack 0.00887f
C946 delay_code[1] a_14799_7041# 4.08e-19
C947 a_15506_5803# a_15506_6427# 0.00442f
C948 a_16704_5987# sar_retimer[4] 0.167f
C949 a_14799_7041# a_15789_7073# 0.00116f
C950 a_14312_7267# sar_logic[1] 0.0872f
C951 a_16320_5787# a_15789_5793# 6.27e-19
C952 a_17307_6153# sar_logic[5] 8.74e-20
C953 a_13397_5793# sar_logic[5] 0.0433f
C954 a_17307_7433# delay_code[0] 6.85e-21
C955 a_16143_7067# a_16344_7445# 3.67e-19
C956 a_16410_6401# a_16875_6709# 9.46e-19
C957 a_15955_6427# a_17103_6793# 2.13e-19
C958 a_14158_6427# x3.X 9.18e-19
C959 a_14625_6427# a_14158_6427# 0.00316f
C960 a_14312_6401# a_14530_6427# 3.73e-19
C961 a_13751_5147# a_13928_5513# 8.94e-19
C962 a_13563_5147# a_14530_5147# 0.00126f
C963 a_13844_5513# a_14158_5147# 0.0258f
C964 a_14312_5121# a_14711_5513# 0.00133f
C965 x2.x5[7].floating delay_code[0] 0.00132f
C966 delay_offset a_13397_7073# 3.76e-21
C967 a_14483_6709# a_13563_6427# 1.09e-19
C968 a_14262_6709# a_14018_6401# 0.0104f
C969 a_17126_6165# a_17307_6153# 4.11e-20
C970 a_17126_5147# sar_logic[7] 2.67e-20
C971 x2.x10.Y a_12322_10357# 1.02e-19
C972 sar_retimer[7] a_16410_5121# 7.43e-20
C973 x2.x3[1].floating x3.A 5.37e-20
C974 sar_retimer[4] a_14625_6165# 1.99e-19
C975 a_13397_7073# a_13844_7067# 0.15f
C976 sar_logic[0] a_14018_7041# 5.76e-19
C977 a_16704_5987# x3.X 0.00116f
C978 sar_logic[3] a_16236_6793# 0.00143f
C979 sar_retimer[6] a_16143_5147# 0.0134f
C980 a_17017_7445# a_16704_6401# 1.96e-20
C981 a_17191_7041# a_17191_6401# 0.016f
C982 a_12457_8692# x2.x7.floating 0.00959f
C983 sar_logic[6] a_14312_5121# 0.00283f
C984 a_15033_7067# a_15789_7073# 4.06e-20
C985 a_17191_7041# x1[3].Q_N 3.56e-19
C986 a_13751_7067# sar_logic[2] 3.37e-20
C987 sar_retimer[4] a_15033_5787# 1.41e-19
C988 a_16654_6709# sar_retimer[2] 0.00291f
C989 a_13563_5147# sar_retimer[6] 3.67e-20
C990 a_12385_8416# delay_offset 3.54e-19
C991 sar_retimer[4] a_15789_5147# 1.32e-19
C992 a_15506_5803# a_14799_6401# 3.81e-19
C993 a_14625_6165# a_14625_6427# 0.00421f
C994 sar_logic[5] a_13844_6793# 2.74e-20
C995 a_13397_5147# a_14262_5429# 0.00276f
C996 a_14625_6165# x3.X 0.00205f
C997 a_13397_5147# sar_logic[4] 3.22e-21
C998 a_13844_5787# a_14018_6401# 3.66e-20
C999 a_14312_5987# a_13563_6427# 1.45e-20
C1000 a_14262_7067# sar_retimer[0] 5.15e-20
C1001 sar_logic[3] sar_retimer[2] 0.044f
C1002 a_16704_7267# a_17898_7083# 6.04e-19
C1003 a_16704_7267# delay_code[0] 0.00142f
C1004 a_16550_7433# a_16922_7389# 3.34e-19
C1005 a_13397_6427# a_14625_7445# 5.98e-20
C1006 a_14312_5121# x3.X 0.00108f
C1007 sar_retimer[3] a_17017_6427# 2.37e-19
C1008 a_16704_5987# a_16704_5121# 0.0106f
C1009 a_15955_7073# a_16236_7067# 0.155f
C1010 a_15033_5787# x3.X 4.06e-19
C1011 x2.x10.Y a_12297_8002# 2.2e-20
C1012 x2.x4[3].floating a_12457_8140# 7.47e-19
C1013 sar_retimer[4] a_17103_5787# 0.00209f
C1014 a_15789_5147# x3.X 0.262f
C1015 x1[7].Q_N sar_retimer[6] 0.0256f
C1016 a_12297_8554# a_12457_8416# 0.0388f
C1017 a_17017_7445# x2.x3[1].floating 9.21e-21
C1018 a_14018_5761# a_14312_5987# 0.199f
C1019 a_13563_5793# a_14799_5761# 0.0264f
C1020 a_15506_6427# a_14799_7041# 3.56e-19
C1021 a_15789_5793# a_16410_5121# 4.47e-20
C1022 a_12457_8692# x2.x6.SW 2.44e-19
C1023 a_15955_5147# a_17103_5513# 2.13e-19
C1024 a_16410_5121# a_16875_5429# 9.46e-19
C1025 a_16704_7267# a_14312_7267# 2.22e-20
C1026 a_16654_6709# x3.X 2.64e-19
C1027 a_17103_5787# x3.X 7.09e-20
C1028 a_13563_5147# a_13844_5787# 1.14e-19
C1029 a_13844_5513# a_13563_5793# 1.14e-19
C1030 x1[2].Q_N a_13397_6427# 1.07e-19
C1031 a_14018_5121# a_14018_5761# 0.00947f
C1032 a_14312_5121# a_16704_5121# 3.6e-20
C1033 a_13751_5787# a_13952_6165# 3.67e-19
C1034 x1[6].Q_N sar_retimer[6] 7.77e-19
C1035 a_14799_5121# a_16236_5513# 7.98e-21
C1036 a_16704_5987# a_17191_6401# 6.54e-20
C1037 a_14711_5787# a_13563_5793# 2.13e-19
C1038 a_17191_5761# a_16704_6401# 6.54e-20
C1039 a_15955_5793# a_17191_5761# 0.0264f
C1040 sar_logic[7] a_16236_5513# 0.00144f
C1041 a_15789_5147# a_16704_5121# 0.124f
C1042 sar_logic[3] a_14625_6427# 0.0362f
C1043 a_14158_7433# a_14530_7389# 3.34e-19
C1044 delay_code[0] x3.X 0.0284f
C1045 sar_logic[3] x3.X 0.108f
C1046 a_17898_7083# x3.X 2.09e-19
C1047 sar_retimer[0] a_16875_7067# 0.00627f
C1048 a_16320_6793# a_15789_6427# 6.27e-19
C1049 a_14915_6153# a_14625_6165# 0.0282f
C1050 a_14158_6153# sar_logic[5] 0.0375f
C1051 sar_retimer[3] sar_retimer[6] 1.41e-19
C1052 a_14262_5787# a_14312_5987# 1.21e-20
C1053 a_15789_5793# a_16236_6793# 9.21e-20
C1054 sar_logic[5] sar_logic[2] 3.33e-19
C1055 a_14483_7067# a_14018_7041# 9.46e-19
C1056 a_13952_7445# sar_logic[1] 0.00177f
C1057 a_14312_6401# a_14625_7445# 1.96e-20
C1058 a_14915_7433# a_14799_7041# 0.0397f
C1059 a_14734_7445# a_14625_7445# 0.00707f
C1060 a_14799_6401# a_14799_7041# 0.016f
C1061 a_14625_6427# a_14312_7267# 1.96e-20
C1062 x3.X a_14312_7267# 0.00549f
C1063 sar_retimer[0] a_17017_6427# 1.27e-20
C1064 a_13751_5787# sar_logic[4] 0.164f
C1065 a_17017_6165# a_16875_5787# 0.00412f
C1066 a_17191_5761# x1[5].Q_N 0.124f
C1067 a_15955_5793# a_16550_6153# 0.00118f
C1068 a_16550_6153# a_16704_6401# 1.58e-19
C1069 a_15789_6427# a_16236_7067# 8.13e-20
C1070 sar_retimer[5] sar_retimer[3] 0.0129f
C1071 a_16550_5147# sar_logic[7] 3.52e-19
C1072 delay_code[0] sar_logic[0] 1.1e-19
C1073 delay_code[1] a_15506_7083# 9.3e-20
C1074 a_13397_5793# a_13397_6427# 0.0151f
C1075 a_13751_7067# a_13397_7073# 0.0662f
C1076 a_17017_6165# sar_retimer[4] 0.0352f
C1077 delay_code[2] x2.x7.floating 0.0102f
C1078 sar_logic[5] a_15506_6427# 1.11e-20
C1079 a_16875_5787# a_15789_5793# 0.00576f
C1080 a_14625_7445# sar_logic[1] 0.0363f
C1081 a_15506_7083# a_15789_7073# 8.18e-19
C1082 a_16236_5787# sar_retimer[6] 1.36e-20
C1083 a_17191_7041# x1[1].Q_N 0.124f
C1084 delay_code[0] x2.x10.Y 0.0125f
C1085 a_17017_7445# a_16875_7067# 0.00412f
C1086 a_14711_7067# x3.X 2.62e-19
C1087 sar_retimer[0] a_15955_7073# 0.0231f
C1088 a_16143_7067# sar_logic[1] 0.165f
C1089 a_16410_6401# a_16550_6427# 0.07f
C1090 a_16704_6401# a_16875_6709# 0.00652f
C1091 a_15955_6427# a_16344_6427# 0.0019f
C1092 delay_code[2] sar_logic[1] 3.62e-21
C1093 a_14625_6427# a_14530_6427# 0.00276f
C1094 a_14799_6401# a_15033_6709# 0.00945f
C1095 a_13563_5147# x1[6].Q_N 4.18e-21
C1096 x1[1].Q_N sar_retimer[1] 8.3e-19
C1097 a_13751_6427# a_13952_6427# 3.67e-19
C1098 a_14530_6427# x3.X 3.13e-19
C1099 a_14625_5147# a_14711_5513# 0.00976f
C1100 a_14312_6401# x1[2].Q_N 0.00553f
C1101 sar_retimer[3] a_15789_6427# 9.98e-20
C1102 a_14158_6427# a_13563_6427# 0.00118f
C1103 sar_logic[0] a_14312_7267# 0.00299f
C1104 a_14158_5147# sar_logic[7] 0.0379f
C1105 a_17898_5147# a_17191_5121# 0.0968f
C1106 sar_retimer[7] a_16704_5121# 5.71e-19
C1107 a_13397_7073# a_14799_7041# 0.0492f
C1108 a_13397_5793# sar_logic[4] 0.313f
C1109 sar_retimer[4] a_15789_5793# 0.708f
C1110 a_17017_6165# x3.X 9.29e-19
C1111 sar_logic[3] a_17191_6401# 7.27e-20
C1112 a_16236_5787# sar_retimer[5] 2.42e-20
C1113 a_17898_7083# a_17191_6401# 3.56e-19
C1114 a_17017_7445# a_17017_6427# 0.0041f
C1115 a_12385_8692# x2.x7.floating 8.52e-19
C1116 sar_logic[6] a_14625_5147# 4.22e-20
C1117 a_16922_7389# a_15789_7073# 2.56e-19
C1118 a_12322_10081# a_12410_9943# 0.0704f
C1119 a_16550_7433# sar_logic[1] 3.4e-19
C1120 a_13844_6793# a_13397_6427# 0.15f
C1121 a_17103_6793# sar_retimer[2] 0.00209f
C1122 a_13844_5513# sar_retimer[6] 2.25e-20
C1123 a_14312_5121# a_15506_5147# 6.04e-19
C1124 a_12457_8140# delay_offset 3.98e-19
C1125 a_15506_5147# a_15789_5147# 8.18e-19
C1126 sar_logic[5] a_14799_6401# 8.35e-20
C1127 a_15789_5793# x3.X 0.27f
C1128 x2.x5[7].floating delay_code[2] 0.00564f
C1129 a_16875_5429# x3.X 1.26e-19
C1130 x2.x2.floating x3.A 0.0198f
C1131 a_15033_7067# a_13397_7073# 1.25e-19
C1132 x1[5].Q_N a_17425_5787# 2.02e-20
C1133 a_16236_5787# a_15789_6427# 9.21e-20
C1134 a_14625_6165# a_13563_6427# 9.03e-20
C1135 a_18195_9015# x2.x9.output_stack 0.00892f
C1136 a_17017_7445# a_15955_7073# 0.137f
C1137 a_15955_6427# a_15789_7073# 1.39e-19
C1138 x1[0].Q_N sar_retimer[0] 7.57e-19
C1139 sar_retimer[1] a_16410_7041# 8.29e-20
C1140 a_16410_5761# a_14312_5987# 4.35e-20
C1141 a_14625_5147# x3.X 8.27e-20
C1142 a_16922_6109# x3.X 2.71e-19
C1143 a_17017_6165# a_16704_5121# 1.96e-20
C1144 a_13397_5147# sar_logic[6] 0.298f
C1145 a_17191_5761# a_17191_5121# 0.016f
C1146 a_16704_5987# a_17017_5147# 1.96e-20
C1147 a_13397_5793# a_14312_6401# 1.07e-20
C1148 a_17307_6427# x3.X 1.91e-19
C1149 a_16236_5787# a_16143_5787# 0.0367f
C1150 a_12385_8554# a_12457_8416# 0.00227f
C1151 a_13844_5787# a_14799_5761# 4.7e-22
C1152 a_17191_7041# a_17898_6427# 3.56e-19
C1153 a_13563_5793# a_15506_5803# 4.46e-21
C1154 a_15506_6427# a_15506_7083# 0.00419f
C1155 a_14018_5761# a_14625_6165# 0.00187f
C1156 a_15789_5793# a_16704_5121# 8.63e-20
C1157 a_16704_5121# a_16875_5429# 0.00652f
C1158 sar_retimer[0] a_15789_6427# 1.36e-19
C1159 a_16704_7267# a_16143_7067# 3.79e-20
C1160 a_13397_5147# x3.X 0.263f
C1161 a_14018_5121# a_14312_5987# 4.94e-20
C1162 a_14312_5121# a_14018_5761# 4.94e-20
C1163 a_13844_5513# a_13844_5787# 0.00445f
C1164 a_17017_6165# a_17191_6401# 2.23e-20
C1165 a_16143_5787# a_14799_5761# 8.26e-21
C1166 a_17191_5761# a_17017_6427# 2.23e-20
C1167 a_15955_5793# a_17898_5803# 4.84e-21
C1168 sar_logic[7] a_17191_5121# 7.2e-20
C1169 a_15789_5147# a_17017_5147# 0.0322f
C1170 a_15955_6427# a_16410_6401# 0.152f
C1171 a_13952_7445# x3.X 1.27e-19
C1172 a_13844_6793# a_14312_6401# 0.0633f
C1173 a_13563_5147# a_13844_5513# 0.146f
C1174 sar_logic[3] a_13563_6427# 0.271f
C1175 a_17898_5147# sar_retimer[6] 0.035f
C1176 a_16704_7267# a_16550_7433# 0.00943f
C1177 x1[2].Q_N sar_retimer[2] 7.51e-19
C1178 sar_retimer[1] a_18195_9015# 6.48e-21
C1179 a_13397_6427# sar_logic[2] 0.243f
C1180 x1[4].Q_N a_14312_5987# 0.00553f
C1181 a_14734_6165# sar_logic[5] 0.00114f
C1182 x2.x4[3].floating a_13563_7073# 9.83e-19
C1183 a_15955_5793# sar_logic[5] 0.252f
C1184 a_14312_5987# a_14915_6427# 1.41e-19
C1185 a_14799_6401# a_15506_7083# 3.56e-19
C1186 a_14530_7389# sar_logic[1] 0.00372f
C1187 a_14483_7067# a_14312_7267# 0.00652f
C1188 a_14625_6427# a_14625_7445# 0.0041f
C1189 x2.x6.floating a_12410_9943# 0.0194f
C1190 x3.X a_14625_7445# 0.00213f
C1191 x2.x5[7].floating a_12322_10081# 2.76e-19
C1192 a_16143_7067# x3.X 0.00452f
C1193 a_14530_6109# a_13397_5793# 2.56e-19
C1194 a_17898_5803# x1[5].Q_N 0.178f
C1195 a_17017_7445# a_15789_6427# 5.98e-20
C1196 a_14018_6401# a_13844_7067# 1.29e-19
C1197 delay_code[2] x3.X 2.69e-19
C1198 delay_code[1] x2.x7.floating 1.53e-20
C1199 a_12322_10081# x2.x6.SW 9.98e-20
C1200 a_17126_6427# a_16704_6401# 2.87e-21
C1201 a_17307_6427# a_17191_6401# 0.0397f
C1202 a_14018_5761# sar_logic[3] 8.96e-20
C1203 a_15506_6427# a_13397_6427# 1.03e-19
C1204 a_16922_5147# sar_logic[7] 1.17e-19
C1205 a_16704_7267# a_17425_7067# 7.78e-19
C1206 a_17425_5429# a_15789_5147# 1.25e-19
C1207 sar_logic[4] sar_logic[2] 0.00425f
C1208 delay_code[1] sar_logic[1] 8.75e-20
C1209 a_13751_5787# sar_logic[6] 3.37e-20
C1210 a_14158_7433# a_13397_7073# 6.04e-20
C1211 sar_retimer[1] x2.x9.output_stack 4.28e-21
C1212 x1[6].Q_N a_14799_5761# 3.56e-19
C1213 a_17191_5761# sar_retimer[6] 1.19e-19
C1214 a_15789_7073# sar_logic[1] 0.273f
C1215 x2.x4[3].floating a_12297_8830# 1.17e-19
C1216 a_17898_7083# x1[1].Q_N 0.178f
C1217 a_16550_7433# x3.X 9.96e-19
C1218 sar_retimer[0] a_16236_7067# 0.0299f
C1219 x2.x7.floating a_12385_8140# 8.52e-19
C1220 a_17191_6401# a_17103_6793# 7.71e-20
C1221 a_16410_6401# a_16922_6427# 9.75e-19
C1222 a_16236_6793# a_16344_6427# 0.00812f
C1223 a_17017_6427# a_16875_6709# 0.00412f
C1224 a_16704_6401# a_16550_6427# 0.00943f
C1225 x1[2].Q_N x3.X 0.00412f
C1226 a_14625_6427# x1[2].Q_N 9.58e-21
C1227 a_14312_5121# a_15033_5429# 0.00185f
C1228 a_17307_5147# a_17126_5147# 4.11e-20
C1229 a_14530_6427# a_13563_6427# 0.00126f
C1230 a_14530_5147# sar_logic[7] 0.00358f
C1231 a_15033_5429# a_15789_5147# 4.06e-20
C1232 a_13397_7073# a_15506_7083# 1.03e-19
C1233 sar_logic[0] a_14625_7445# 1.88e-20
C1234 sar_retimer[7] a_17017_5147# 2.27e-19
C1235 a_13751_5787# x3.X 0.0044f
C1236 a_14158_6153# a_14312_6401# 1.58e-19
C1237 sar_retimer[0] a_13563_7073# 3.45e-20
C1238 sar_logic[3] a_16143_6427# 0.165f
C1239 sar_retimer[6] a_16654_5429# 0.00292f
C1240 delay_code[2] sar_logic[0] 7.09e-20
C1241 a_17191_5761# sar_retimer[5] 0.00464f
C1242 a_15955_5147# a_16410_5121# 0.152f
C1243 a_16410_6401# a_14312_6401# 3.1e-20
C1244 a_15955_6427# a_14799_6401# 2.24e-20
C1245 x2.x6.floating x2.x7.floating 0.202f
C1246 a_12457_8416# x2.x7.floating 0.00959f
C1247 a_17126_7445# sar_logic[1] 2.61e-20
C1248 x2.x5[7].floating delay_code[1] 0.00228f
C1249 a_12410_9943# a_12322_9805# 0.0704f
C1250 a_17425_7067# x3.X 5.66e-20
C1251 a_14799_6401# a_13397_6427# 0.0492f
C1252 sar_logic[6] a_13397_5793# 3.13e-21
C1253 a_14312_6401# sar_logic[2] 1.88e-19
C1254 a_14799_5121# sar_retimer[6] 0.00447f
C1255 a_16410_5761# a_16704_5987# 0.199f
C1256 sar_retimer[4] a_13397_5793# 9.31e-20
C1257 delay_code[2] x2.x10.Y 0.00203f
C1258 sar_retimer[6] sar_logic[7] 0.0435f
C1259 a_14312_5987# a_14158_6427# 1.58e-19
C1260 a_17191_7041# sar_retimer[1] 0.00444f
C1261 a_16236_6793# a_15789_7073# 8.13e-20
C1262 a_12385_8968# x2.x9.output_stack 0.00227f
C1263 delay_code[0] a_16410_7041# 2.45e-19
C1264 a_13844_6793# sar_retimer[2] 2.2e-20
C1265 a_14312_6401# a_15506_6427# 6.04e-19
C1266 a_16236_5787# a_14799_5761# 7.98e-21
C1267 a_16704_5987# a_14312_5987# 3.43e-20
C1268 x1[7].Q_N a_17898_5147# 0.178f
C1269 a_17126_7445# a_17307_7433# 4.11e-20
C1270 a_13928_5513# x3.X 4.41e-19
C1271 a_17017_6165# a_17017_5147# 0.0041f
C1272 a_17307_6153# x3.X 2.01e-19
C1273 a_13397_5793# a_14625_6427# 7.69e-20
C1274 a_17898_5803# a_17191_5121# 3.56e-19
C1275 a_13397_5793# x3.X 0.271f
C1276 a_16550_6153# sar_retimer[5] 9.61e-20
C1277 a_13397_5147# a_15506_5147# 1.03e-19
C1278 a_16704_7267# delay_code[1] 1.69e-20
C1279 a_12457_8416# a_12297_8278# 0.0388f
C1280 a_13397_6427# a_13397_7073# 0.015f
C1281 x2.x6.floating x2.x5[7].floating 1.18f
C1282 a_16410_5761# a_15789_5147# 4.47e-20
C1283 a_14312_7267# a_16410_7041# 3.01e-20
C1284 a_14799_7041# a_15955_7073# 2.24e-20
C1285 a_13563_5793# sar_logic[5] 0.274f
C1286 a_14312_5987# a_14625_6165# 0.124f
C1287 sar_retimer[2] a_15789_7073# 1.32e-19
C1288 a_17898_7083# a_17898_6427# 0.00419f
C1289 a_15789_5793# a_17017_5147# 5.98e-20
C1290 a_12457_8416# x2.x6.SW 1.28e-19
C1291 a_16344_6427# x3.X 3.03e-19
C1292 a_17191_5121# a_17103_5513# 7.71e-20
C1293 x2.x6.floating x2.x6.SW 0.13f
C1294 a_17017_5147# a_16875_5429# 0.00412f
C1295 a_16704_7267# a_15789_7073# 0.124f
C1296 a_16704_5987# x1[4].Q_N 2.9e-20
C1297 a_14312_5121# a_14312_5987# 0.0106f
C1298 a_14158_6153# a_14530_6109# 3.34e-19
C1299 a_14799_5121# a_16143_5147# 8.26e-21
C1300 a_14711_5787# a_14799_5761# 7.71e-20
C1301 a_15033_5787# a_14312_5987# 0.00185f
C1302 a_13563_7073# a_13844_7067# 0.146f
C1303 a_17191_5761# x1[7].Q_N 3.56e-19
C1304 a_15955_5793# a_15955_6427# 0.0109f
C1305 a_16410_6401# a_16236_6793# 0.205f
C1306 a_15955_6427# a_16704_6401# 0.139f
C1307 sar_logic[7] a_16143_5147# 0.165f
C1308 a_15789_5147# a_16320_5513# 7.03e-19
C1309 a_14734_7445# a_14915_7433# 4.11e-20
C1310 a_14312_6401# a_14799_6401# 0.272f
C1311 a_14530_7389# x3.X 3.48e-19
C1312 a_13844_6793# x3.X 0.00438f
C1313 a_13563_5147# a_14799_5121# 0.0264f
C1314 a_14018_5121# a_14312_5121# 0.199f
C1315 a_18195_9015# delay_code[0] 0.00169f
C1316 a_13563_5147# sar_logic[7] 0.271f
C1317 a_16875_6709# a_15789_6427# 0.00576f
C1318 a_16704_7267# a_17126_7445# 2.87e-21
C1319 x2.x4[3].floating delay_offset 0.00402f
C1320 a_16143_5787# sar_logic[7] 3.37e-20
C1321 sar_retimer[4] a_15955_5147# 1.01e-19
C1322 x1[4].Q_N a_14625_6165# 9.58e-21
C1323 x2.x4[3].floating a_13844_7067# 1.78e-19
C1324 a_14625_6165# a_14915_6427# 6.09e-20
C1325 delay_code[1] x3.X 6.2e-19
C1326 a_12322_10081# x2.x10.Y 2.35e-19
C1327 a_13397_5147# a_14018_5761# 4.47e-20
C1328 x1[0].Q_N a_14799_7041# 0.124f
C1329 x3.X a_15789_7073# 0.268f
C1330 a_14483_7067# a_14625_7445# 0.00412f
C1331 a_14915_7433# sar_logic[1] 0.0397f
C1332 a_16410_6401# sar_retimer[2] 0.0293f
C1333 a_12297_8830# delay_offset 0.0165f
C1334 x2.x5[7].floating a_12322_9805# 2.76e-19
C1335 x1[4].Q_N a_15033_5787# 2.02e-20
C1336 a_17103_7067# a_15955_7073# 2.13e-19
C1337 a_15955_5793# a_16320_5787# 4.45e-20
C1338 a_13563_6427# a_14625_7445# 8.13e-20
C1339 a_16704_7267# a_16410_6401# 4.94e-20
C1340 a_12322_9805# x2.x6.SW 0.00707f
C1341 a_14312_5987# sar_logic[3] 8.06e-20
C1342 a_17126_6427# a_17017_6427# 0.00707f
C1343 x2.x3[1].floating a_18499_9105# 4.53e-20
C1344 a_15955_5147# x3.X 0.00724f
C1345 delay_code[0] x2.x9.output_stack 0.0322f
C1346 a_14312_6401# a_13397_7073# 8.63e-20
C1347 a_17017_7445# sar_retimer[0] 0.0354f
C1348 x1[0].Q_N a_15033_7067# 2.02e-20
C1349 a_15506_6427# sar_retimer[2] 0.0744f
C1350 a_16704_6401# a_16922_6427# 3.73e-19
C1351 a_17126_7445# x3.X 5.56e-20
C1352 a_17017_6427# a_16550_6427# 0.00316f
C1353 delay_code[1] sar_logic[0] 8.75e-20
C1354 a_14799_5121# x1[6].Q_N 0.124f
C1355 x1[2].Q_N a_13563_6427# 4.89e-21
C1356 x1[6].Q_N sar_logic[7] 0.0243f
C1357 a_12297_8830# a_12385_8830# 0.00227f
C1358 a_13397_7073# sar_logic[1] 0.0432f
C1359 sar_retimer[0] a_13844_7067# 2.24e-20
C1360 a_14158_6153# x3.X 9.34e-19
C1361 delay_code[1] x2.x10.Y 7.14e-19
C1362 sar_logic[5] sar_retimer[6] 1.22e-20
C1363 a_16704_6401# a_14312_6401# 2.29e-20
C1364 sar_logic[3] a_14915_6427# 0.0398f
C1365 a_16410_5121# a_16236_5513# 0.205f
C1366 sar_retimer[6] a_17103_5513# 0.00205f
C1367 a_17898_5803# sar_retimer[5] 0.0764f
C1368 a_16236_6793# a_14799_6401# 7.98e-21
C1369 a_15955_5147# a_16704_5121# 0.139f
C1370 a_16410_6401# x3.X 0.00261f
C1371 a_12385_8416# x2.x7.floating 8.52e-19
C1372 a_16654_7067# a_15789_7073# 0.00117f
C1373 sar_logic[2] x3.X 0.084f
C1374 a_13751_6427# a_13397_6427# 0.0695f
C1375 a_14625_6427# sar_logic[2] 1.19e-20
C1376 a_16410_5761# a_17017_6165# 0.00187f
C1377 sar_retimer[4] a_16654_5787# 0.00291f
C1378 a_16236_5787# a_17191_5761# 4.7e-22
C1379 a_15033_6709# a_15789_6427# 4.06e-20
C1380 a_17191_7041# a_17898_7083# 0.0968f
C1381 a_17191_7041# delay_code[0] 1.11e-19
C1382 a_13397_5147# a_15033_5429# 1.25e-19
C1383 sar_logic[5] a_14018_6401# 9.19e-20
C1384 a_17898_7083# sar_retimer[1] 0.0748f
C1385 a_12457_8692# x2.x9.output_stack 0.032f
C1386 a_14799_6401# sar_retimer[2] 0.00449f
C1387 a_15506_6427# x3.X 0.0331f
C1388 a_13952_6165# a_13563_5793# 0.00114f
C1389 a_13751_5787# a_14018_5761# 6.99e-20
C1390 a_16410_5761# a_15789_5793# 0.111f
C1391 a_14483_5429# x3.X 1.52e-19
C1392 sar_logic[4] a_13751_6427# 4.77e-20
C1393 a_16654_5787# x3.X 2.64e-19
C1394 a_16344_5147# a_15955_5147# 0.0019f
C1395 a_17126_6165# sar_retimer[5] 4.55e-20
C1396 a_16550_5147# a_16410_5121# 0.07f
C1397 a_13751_7067# a_13563_7073# 0.158f
C1398 a_13563_5793# a_13397_6427# 4.5e-20
C1399 x2.x6.floating x2.x10.Y 0.0881f
C1400 a_13397_5793# a_13563_6427# 4.5e-20
C1401 delay_code[0] a_14018_7041# 2.45e-19
C1402 sar_logic[5] a_15789_6427# 6.82e-20
C1403 a_16410_5761# a_16922_6109# 9.75e-19
C1404 a_16236_5787# a_16550_6153# 0.0258f
C1405 sar_logic[2] sar_logic[0] 0.00838f
C1406 a_12297_8278# a_12385_8416# 0.00227f
C1407 a_16704_5987# a_15789_5147# 8.63e-20
C1408 a_14799_7041# a_16236_7067# 7.98e-21
C1409 a_14312_5987# a_15789_5793# 3.34e-19
C1410 a_13844_5787# sar_logic[5] 0.0391f
C1411 a_14799_5761# a_15506_5803# 0.0968f
C1412 a_16143_7067# a_16410_7041# 6.99e-20
C1413 a_16344_7445# a_15955_7073# 0.0019f
C1414 sar_logic[5] a_16143_5147# 3.37e-20
C1415 x1[1].Q_N a_17425_7067# 2.02e-20
C1416 a_14625_5147# a_14312_5987# 1.96e-20
C1417 a_14312_5121# a_14625_6165# 1.96e-20
C1418 a_12410_10219# delay_offset 1.9e-19
C1419 a_14799_5121# a_14799_5761# 0.016f
C1420 a_17307_5147# a_17191_5121# 0.0397f
C1421 a_17126_5147# a_16704_5121# 2.87e-21
C1422 a_14312_5121# a_14734_5147# 2.87e-21
C1423 a_14799_5121# a_14915_5147# 0.0397f
C1424 a_13563_7073# a_14799_7041# 0.0264f
C1425 a_16143_5787# sar_logic[5] 0.166f
C1426 a_14018_7041# a_14312_7267# 0.199f
C1427 a_13397_5793# a_14018_5761# 0.117f
C1428 sar_logic[4] a_13563_5793# 0.165f
C1429 a_15955_5793# a_16236_6793# 1.56e-19
C1430 a_15955_6427# a_17017_6427# 0.137f
C1431 sar_logic[7] a_14915_5147# 0.0398f
C1432 a_16236_6793# a_16704_6401# 0.0633f
C1433 sar_logic[3] a_14158_6427# 0.0379f
C1434 a_14915_7433# x3.X 0.00114f
C1435 x2.x3[1].floating sar_logic[1] 6.32e-19
C1436 a_16704_5987# a_17103_5787# 3.57e-19
C1437 a_14799_6401# x3.X 0.0128f
C1438 a_14312_6401# a_13751_6427# 3.79e-20
C1439 a_14799_6401# a_14625_6427# 0.197f
C1440 a_13844_6793# a_13928_6793# 0.00972f
C1441 a_13844_5513# a_14799_5121# 4.7e-22
C1442 a_13563_5147# a_13751_5147# 0.158f
C1443 a_14018_5121# a_14625_5147# 0.00187f
C1444 a_16922_7389# a_15955_7073# 0.00126f
C1445 a_16550_7433# a_16410_7041# 0.07f
C1446 a_13844_6793# a_13563_6427# 0.146f
C1447 a_14312_5121# a_15789_5147# 3.41e-19
C1448 a_16550_6427# a_15789_6427# 6.04e-20
C1449 a_13844_5513# sar_logic[7] 0.0388f
C1450 sar_retimer[4] a_16236_5513# 1.35e-20
C1451 x1[4].Q_N a_15789_5793# 2.94e-19
C1452 x2.x4[3].floating a_14799_7041# 0.00104f
C1453 a_12322_9805# x2.x10.Y 0.039f
C1454 a_13397_5147# a_14312_5987# 8.63e-20
C1455 x1[0].Q_N a_15506_7083# 0.178f
C1456 a_15955_6427# a_15955_7073# 0.0099f
C1457 a_12385_8830# delay_offset 7.9e-19
C1458 a_16704_6401# sar_retimer[2] 0.167f
C1459 a_14262_5787# a_13397_5793# 0.00276f
C1460 a_15955_5793# a_16875_5787# 1.09e-19
C1461 a_16704_7267# a_16704_6401# 0.0106f
C1462 a_14625_6165# sar_logic[3] 1.95e-20
C1463 a_13397_5147# a_14018_5121# 0.117f
C1464 a_17425_6709# sar_retimer[2] 0.00258f
C1465 x2.x3[1].floating x2.x5[7].floating 0.8f
C1466 a_14018_5761# a_13844_6793# 3.66e-20
C1467 a_13563_5793# a_14312_6401# 1.45e-20
C1468 a_16236_5513# x3.X 0.00252f
C1469 a_17191_5761# a_17898_5147# 3.56e-19
C1470 a_14625_6427# a_13397_7073# 5.98e-20
C1471 a_13928_7067# a_13397_7073# 0.0018f
C1472 x3.X a_13397_7073# 0.269f
C1473 a_15955_5793# sar_retimer[4] 0.0229f
C1474 x2.x4[3].floating a_12297_8554# 1.17e-19
C1475 a_16320_7067# x3.X 2.8e-19
C1476 a_17017_6427# a_16922_6427# 0.00276f
C1477 a_16143_6427# a_16344_6427# 3.67e-19
C1478 a_14158_6427# a_14530_6427# 3.34e-19
C1479 x2.x2.floating a_18499_9105# 0.00119f
C1480 a_12297_8830# a_12297_8554# 0.0316f
C1481 delay_code[2] x2.x9.output_stack 0.332f
C1482 a_14734_6165# x3.X 7.88e-20
C1483 sar_retimer[0] a_14799_7041# 0.00439f
C1484 a_15955_5793# x3.X 0.0134f
C1485 a_16236_5513# a_16704_5121# 0.0633f
C1486 a_15955_5147# a_17017_5147# 0.137f
C1487 a_16704_6401# x3.X 0.00155f
C1488 x1[1].Q_N a_15789_7073# 1.07e-19
C1489 a_12457_8140# x2.x7.floating 0.00925f
C1490 a_16704_7267# x2.x3[1].floating 6.81e-19
C1491 a_14262_6709# a_13397_6427# 0.00276f
C1492 a_14262_5429# sar_retimer[6] 5.18e-20
C1493 sar_retimer[7] a_15789_5147# 9.3e-20
C1494 a_16704_5987# a_17017_6165# 0.12f
C1495 a_13397_7073# sar_logic[0] 0.309f
C1496 sar_retimer[4] x1[5].Q_N 0.0257f
C1497 sar_retimer[3] a_17126_6427# 5.17e-20
C1498 a_13397_6427# a_14018_6401# 0.117f
C1499 sar_logic[2] a_13563_6427# 0.217f
C1500 sar_retimer[0] a_15033_7067# 1.56e-19
C1501 a_15955_6427# a_15789_6427# 0.741f
C1502 a_14158_6153# a_14018_5761# 0.07f
C1503 a_13952_6165# a_13844_5787# 0.00812f
C1504 a_13751_5787# a_14312_5987# 5.76e-21
C1505 a_16236_5787# sar_logic[5] 0.0015f
C1506 a_16704_5987# a_15789_5793# 0.124f
C1507 a_14530_6109# a_13563_5793# 0.00126f
C1508 a_15789_6427# a_13397_6427# 0.00176f
C1509 a_15506_6427# a_13563_6427# 1.06e-20
C1510 sar_retimer[3] a_16550_6427# 9.43e-20
C1511 a_16922_5147# a_16410_5121# 9.75e-19
C1512 a_16550_5147# a_16704_5121# 0.00943f
C1513 a_16344_5147# a_16236_5513# 0.00812f
C1514 a_14158_7433# a_13563_7073# 0.00118f
C1515 delay_code[0] a_14312_7267# 3.02e-19
C1516 a_13751_7067# a_13844_7067# 0.0367f
C1517 a_13844_5787# a_13397_6427# 9.21e-20
C1518 a_17017_7445# a_14799_7041# 1.86e-21
C1519 delay_code[1] a_16410_7041# 8.75e-20
C1520 a_16704_5987# a_16922_6109# 3.73e-19
C1521 a_12297_8278# a_12457_8140# 0.0388f
C1522 a_16704_5987# a_17307_6427# 1.41e-19
C1523 a_15789_7073# a_16410_7041# 0.111f
C1524 sar_logic[1] a_15955_7073# 0.246f
C1525 x2.x3[1].floating x3.X 3.43e-20
C1526 a_17017_6165# a_15789_5147# 5.98e-20
C1527 sar_retimer[0] a_17103_7067# 0.00211f
C1528 a_14625_6165# a_15789_5793# 6.38e-20
C1529 a_14799_5761# sar_logic[5] 0.0311f
C1530 a_12457_8140# x2.x6.SW 7.9e-20
C1531 a_16344_7445# a_16236_7067# 0.00812f
C1532 a_14799_5121# a_15506_5803# 3.56e-19
C1533 a_14625_5147# a_14625_6165# 0.0041f
C1534 a_14734_6165# a_14915_6153# 4.11e-20
C1535 a_14625_5147# a_14734_5147# 0.00707f
C1536 a_13844_7067# a_14799_7041# 4.7e-22
C1537 a_14018_7041# a_14625_7445# 0.00187f
C1538 a_17126_5147# a_17017_5147# 0.00707f
C1539 sar_logic[4] a_13844_5787# 0.00149f
C1540 a_13397_5793# a_14312_5987# 0.125f
C1541 a_15033_5787# a_15789_5793# 4.06e-20
C1542 a_16236_5787# a_16550_6427# 8.58e-20
C1543 a_15789_5793# a_15789_5147# 0.015f
C1544 a_16704_6401# a_17191_6401# 0.27f
C1545 a_15789_5147# a_16875_5429# 0.00592f
C1546 delay_code[2] a_14018_7041# 7.81e-20
C1547 a_15955_6427# a_16320_6793# 4.45e-20
C1548 a_16410_6401# a_16143_6427# 6.99e-20
C1549 sar_logic[3] a_14530_6427# 0.00362f
C1550 a_14312_6401# a_14262_6709# 1.21e-20
C1551 a_17017_6165# a_17103_5787# 0.00976f
C1552 a_14262_7067# x3.X 4.92e-19
C1553 a_17191_5761# a_17425_5787# 0.00945f
C1554 a_13751_6427# x3.X 0.00505f
C1555 a_13844_5513# a_13751_5147# 0.0367f
C1556 a_14018_5121# a_13928_5513# 6.69e-20
C1557 a_14312_5121# a_14625_5147# 0.124f
C1558 a_13563_5147# a_14262_5429# 2.46e-19
C1559 a_16550_7433# sar_retimer[1] 8.77e-20
C1560 a_17425_6709# a_17191_6401# 0.00945f
C1561 x1[3].Q_N a_16704_6401# 0.00553f
C1562 a_14018_5121# a_13397_5793# 4.47e-20
C1563 a_14312_6401# a_14018_6401# 0.199f
C1564 a_14799_6401# a_13563_6427# 0.0264f
C1565 a_14625_5147# a_15789_5147# 6.38e-20
C1566 a_14799_5121# sar_logic[7] 0.0309f
C1567 a_16143_5787# a_16320_5787# 8.94e-19
C1568 a_16922_6427# a_15789_6427# 2.56e-19
C1569 sar_retimer[4] a_13563_5793# 3.88e-20
C1570 a_16704_7267# a_16875_7067# 0.00652f
C1571 sar_retimer[4] a_17191_5121# 1.27e-19
C1572 a_17425_6709# x1[3].Q_N 2.02e-20
C1573 x2.x4[3].floating a_15506_7083# 4.83e-19
C1574 sar_retimer[6] a_16410_5121# 0.0289f
C1575 a_18195_9015# delay_code[1] 3.4e-20
C1576 a_13397_5147# a_14625_6165# 5.98e-20
C1577 a_14711_7067# a_14312_7267# 0.00133f
C1578 a_17017_7445# a_17103_7067# 0.00976f
C1579 a_17191_7041# a_17425_7067# 0.00945f
C1580 a_16236_6793# a_15955_7073# 1.14e-19
C1581 x1[0].Q_N sar_logic[1] 0.0244f
C1582 a_15955_6427# a_16236_7067# 1.14e-19
C1583 a_16410_6401# a_16410_7041# 0.00947f
C1584 a_17017_6427# sar_retimer[2] 0.0352f
C1585 x2.x3[1].floating x2.x10.Y 0.00302f
C1586 a_12297_8554# delay_offset 0.0014f
C1587 a_14312_6401# a_15789_6427# 2.85e-19
C1588 x1[4].Q_N a_13397_5793# 1.07e-19
C1589 a_16704_7267# a_17017_6427# 1.96e-20
C1590 x1[5].Q_N a_17191_6401# 3.57e-19
C1591 a_13397_5147# a_14312_5121# 0.125f
C1592 a_15789_5793# sar_logic[3] 5.58e-20
C1593 a_13563_5793# a_14625_6427# 9.03e-20
C1594 a_13563_5793# x3.X 0.021f
C1595 a_13397_5147# a_15789_5147# 0.00176f
C1596 a_14262_7067# sar_logic[0] 2.51e-21
C1597 a_13751_6427# sar_logic[0] 3.37e-20
C1598 a_17898_5803# a_17898_5147# 0.00419f
C1599 a_14483_7067# a_13397_7073# 0.00907f
C1600 a_13397_6427# a_13563_7073# 1.39e-19
C1601 a_13563_6427# a_13397_7073# 1.39e-19
C1602 sar_retimer[3] a_15955_6427# 4.6e-20
C1603 a_17307_6427# sar_logic[3] 7.35e-20
C1604 sar_retimer[2] a_15955_7073# 1.01e-19
C1605 a_16875_7067# x3.X 3.98e-19
C1606 delay_code[1] x2.x9.output_stack 0.0746f
C1607 a_16704_7267# a_15955_7073# 0.139f
C1608 x2.x2.floating x2.x5[7].floating 0.441f
C1609 a_12322_10081# a_12322_10357# 0.0316f
C1610 sar_retimer[0] a_15506_7083# 0.0744f
C1611 a_13928_5787# x3.X 4.41e-19
C1612 a_16704_5121# a_17191_5121# 0.27f
C1613 a_15955_5147# a_16320_5513# 4.45e-20
C1614 a_16143_6427# a_14799_6401# 8.26e-21
C1615 a_16410_5121# a_16143_5147# 6.99e-20
C1616 a_17017_6427# x3.X 3.22e-19
C1617 a_14711_5513# sar_retimer[6] 8.94e-20
C1618 a_17191_5761# a_17898_5803# 0.0968f
C1619 a_16236_5787# a_15955_6427# 1.56e-19
C1620 a_16410_5761# a_16410_6401# 0.00923f
C1621 x3.A a_18499_9105# 0.171f
C1622 x2.x6.floating x2.x9.output_stack 0.229f
C1623 a_12457_8416# x2.x9.output_stack 1.74e-19
C1624 x3.X a_15955_7073# 0.0123f
C1625 a_16236_6793# a_15789_6427# 0.14f
C1626 a_14262_6709# sar_retimer[2] 5.06e-20
C1627 a_17191_5761# sar_logic[5] 7.67e-20
C1628 sar_retimer[4] sar_retimer[6] 0.0139f
C1629 a_14158_6153# a_14312_5987# 0.00943f
C1630 a_17017_6165# a_15789_5793# 0.0322f
C1631 a_16704_7267# x1[0].Q_N 2.27e-20
C1632 sar_retimer[3] a_16922_6427# 1.03e-19
C1633 sar_retimer[2] a_14018_6401# 7.75e-20
C1634 a_15955_5793# a_17017_5147# 8.13e-20
C1635 a_16704_7267# x2.x2.floating 3.8e-19
C1636 a_16922_5147# a_16704_5121# 3.73e-19
C1637 a_16550_5147# a_17017_5147# 0.00316f
C1638 a_17191_7041# a_15789_7073# 0.0492f
C1639 a_14530_7389# a_14018_7041# 9.75e-19
C1640 a_13844_6793# a_14018_7041# 1.29e-19
C1641 delay_code[0] a_14625_7445# 1.08e-19
C1642 a_14158_7433# a_13844_7067# 0.0258f
C1643 sar_retimer[0] a_15955_6427# 1.06e-19
C1644 a_16143_7067# sar_logic[3] 3.37e-20
C1645 a_16410_5761# a_16654_5787# 0.0104f
C1646 a_17017_6165# a_16922_6109# 0.00276f
C1647 a_16704_5987# a_17307_6153# 0.0549f
C1648 a_17191_5761# a_17126_6165# 4.2e-20
C1649 a_16236_5787# a_16320_5787# 0.00972f
C1650 a_17017_6165# a_17307_6427# 6.09e-20
C1651 a_12385_8278# a_12457_8140# 0.00227f
C1652 sar_retimer[1] a_15789_7073# 1.18e-19
C1653 delay_code[2] delay_code[0] 7.66e-20
C1654 sar_logic[1] a_16236_7067# 0.00139f
C1655 a_15506_5803# sar_logic[5] 0.043f
C1656 sar_retimer[6] x3.X 0.112f
C1657 sar_retimer[4] sar_retimer[5] 0.0492f
C1658 sar_retimer[2] a_15789_6427# 0.708f
C1659 a_16704_7267# a_15789_6427# 8.63e-20
C1660 delay_code[1] a_14018_7041# 1.97e-19
C1661 a_14312_7267# a_14625_7445# 0.124f
C1662 a_16922_6109# a_15789_5793# 2.56e-19
C1663 a_13563_7073# sar_logic[1] 0.274f
C1664 a_16550_6153# sar_logic[5] 3.58e-19
C1665 sar_logic[4] a_14799_5761# 1.34e-20
C1666 a_13397_5793# a_14625_6165# 0.0334f
C1667 a_16143_7067# a_14312_7267# 2.15e-20
C1668 sar_logic[5] sar_logic[7] 0.0041f
C1669 a_17017_7445# a_16922_7389# 0.00276f
C1670 a_17191_7041# a_17126_7445# 4.2e-20
C1671 a_16236_6793# a_16320_6793# 0.00972f
C1672 sar_logic[3] x1[2].Q_N 0.0243f
C1673 delay_code[2] a_14312_7267# 1.33e-20
C1674 a_16704_6401# a_16143_6427# 3.79e-20
C1675 a_17191_6401# a_17017_6427# 0.197f
C1676 a_14262_6709# x3.X 3.69e-19
C1677 a_14312_6401# a_14711_6793# 0.00133f
C1678 a_13844_6793# a_14158_6427# 0.0258f
C1679 a_13751_6427# a_13928_6793# 8.94e-19
C1680 x1[0].Q_N x3.X 0.00412f
C1681 a_17126_7445# sar_retimer[1] 4.44e-20
C1682 a_13563_5147# a_14711_5513# 2.13e-19
C1683 a_14018_5121# a_14483_5429# 9.46e-19
C1684 a_12322_9805# x2.x9.output_stack 0.0702f
C1685 x2.x2.floating x3.X 0.01f
C1686 a_16320_7067# a_16410_7041# 6.69e-20
C1687 x1[3].Q_N a_17017_6427# 9.58e-21
C1688 a_16654_7067# a_15955_7073# 2.46e-19
C1689 x2.x4[3].floating x2.x7.floating 1.18f
C1690 a_14625_6427# a_14018_6401# 0.00187f
C1691 a_13751_6427# a_13563_6427# 0.155f
C1692 a_14018_6401# x3.X 0.0029f
C1693 a_14312_5121# a_13397_5793# 8.63e-20
C1694 a_16550_6153# a_17126_6165# 2.46e-21
C1695 a_13751_5147# sar_logic[7] 0.0194f
C1696 a_15033_5787# a_13397_5793# 1.25e-19
C1697 sar_retimer[4] a_13844_5787# 2.21e-20
C1698 sar_retimer[6] a_16704_5121# 0.164f
C1699 a_17017_7445# a_15955_6427# 8.13e-20
C1700 x2.x6.floating a_12322_10357# 0.00578f
C1701 a_12297_8830# x2.x7.floating 0.00409f
C1702 sar_logic[6] a_13563_5147# 0.167f
C1703 a_15033_7067# a_14799_7041# 0.00945f
C1704 a_14711_7067# a_14625_7445# 0.00976f
C1705 sar_retimer[4] a_16143_5787# 0.0139f
C1706 a_16236_6793# a_16236_7067# 0.00445f
C1707 a_16704_6401# a_16410_7041# 4.94e-20
C1708 a_16320_6793# sar_retimer[2] 0.00223f
C1709 a_14625_6427# a_15789_6427# 6.38e-20
C1710 a_12385_8554# delay_offset 4.7e-19
C1711 a_15789_6427# x3.X 0.27f
C1712 a_14799_5761# a_14312_6401# 6.54e-20
C1713 a_13397_5147# a_14625_5147# 0.0334f
C1714 a_14312_5987# a_14799_6401# 6.54e-20
C1715 a_13844_5787# x3.X 0.00421f
C1716 a_16143_5147# x3.X 0.00275f
C1717 a_12297_8002# a_12385_8140# 0.00227f
C1718 a_13563_5793# a_13563_6427# 0.0109f
C1719 a_14483_5787# sar_retimer[4] 1.51e-19
C1720 a_13563_5147# x3.X 0.0147f
C1721 a_13397_6427# a_13844_7067# 8.13e-20
C1722 a_13397_5793# sar_logic[3] 1.75e-19
C1723 a_16410_5761# a_16236_5513# 1.29e-19
C1724 a_16236_5787# a_16410_5121# 1.29e-19
C1725 sar_retimer[3] a_16236_6793# 2.14e-20
C1726 a_17898_6427# a_16704_6401# 6.04e-19
C1727 sar_retimer[2] a_16236_7067# 1.35e-20
C1728 x2.x4[3].floating a_12297_8278# 1.17e-19
C1729 a_16143_5787# x3.X 0.00503f
C1730 x2.x4[3].floating x2.x5[7].floating 1.55f
C1731 a_16704_7267# a_16236_7067# 0.0633f
C1732 x2.x2.floating x2.x10.Y 0.00202f
C1733 a_12457_8692# a_12385_8692# 0.00227f
C1734 a_13563_5793# a_14018_5761# 0.153f
C1735 x1[4].Q_N a_14799_6401# 3.57e-19
C1736 sar_retimer[0] sar_logic[1] 0.0441f
C1737 a_14483_5787# x3.X 9.28e-19
C1738 sar_logic[3] a_16344_6427# 2.99e-19
C1739 a_12297_8830# x2.x6.SW 0.00179f
C1740 a_16704_5121# a_16143_5147# 3.79e-20
C1741 a_16236_5513# a_16320_5513# 0.00972f
C1742 a_14734_6427# a_14312_6401# 2.87e-21
C1743 a_14915_6427# a_14799_6401# 0.0397f
C1744 a_17191_5121# a_17017_5147# 0.197f
C1745 a_16320_6793# x3.X 2.86e-19
C1746 x2.x3[1].floating a_16410_7041# 1.08e-19
C1747 a_12410_9943# delay_offset 3.64e-19
C1748 sar_retimer[3] sar_retimer[2] 0.0479f
C1749 a_12410_10219# a_12410_9943# 0.0316f
C1750 a_14312_5121# a_15955_5147# 8.45e-20
C1751 a_15955_5793# a_16410_5761# 0.153f
C1752 a_16410_5761# a_16704_6401# 6.09e-20
C1753 a_16704_5987# a_16410_6401# 6.09e-20
C1754 a_16236_5787# a_16236_6793# 0.00451f
C1755 sar_logic[3] a_13844_6793# 0.0388f
C1756 a_15789_5147# a_15955_5147# 0.741f
C1757 x3.A x2.x5[7].floating 0.0216f
C1758 x3.X a_16236_7067# 0.00382f
C1759 sar_retimer[4] sar_retimer[3] 2.05e-19
C1760 a_14711_6793# sar_retimer[2] 8.74e-20
C1761 a_17191_6401# a_15789_6427# 0.0492f
C1762 x1[6].Q_N x3.X 0.00281f
C1763 a_14734_6165# a_14312_5987# 2.87e-21
C1764 a_14158_6153# a_14625_6165# 0.00316f
C1765 a_14262_5787# a_13563_5793# 2.46e-19
C1766 a_13928_5787# a_14018_5761# 6.69e-20
C1767 a_15506_5147# sar_retimer[6] 0.0744f
C1768 a_15955_5793# a_14312_5987# 8.09e-20
C1769 x1[3].Q_N a_15789_6427# 1.07e-19
C1770 delay_code[1] delay_code[0] 1.97f
C1771 x1[7].Q_N a_16704_5121# 0.00553f
C1772 a_17425_5429# a_17191_5121# 0.00945f
C1773 a_16344_5147# a_16143_5147# 3.67e-19
C1774 a_16922_5147# a_17017_5147# 0.00276f
C1775 a_14625_6427# a_13563_7073# 8.13e-20
C1776 a_13928_7067# a_13563_7073# 4.45e-20
C1777 a_17898_7083# a_15789_7073# 1.03e-19
C1778 delay_code[0] a_15789_7073# 4.1e-19
C1779 a_17017_7445# sar_logic[1] 1.2e-19
C1780 a_14530_7389# a_14312_7267# 3.73e-19
C1781 sar_retimer[0] a_16236_6793# 1.34e-20
C1782 x3.X a_13563_7073# 0.0188f
C1783 a_16704_5987# a_16654_5787# 1.21e-20
C1784 a_17017_6165# a_17307_6153# 0.0282f
C1785 a_15955_5793# a_16344_6165# 0.0019f
C1786 x2.x3[1].floating a_18195_9015# 3.09e-19
C1787 sar_retimer[3] x3.X 1.82e-19
C1788 x2.x7.floating delay_offset 0.17f
C1789 a_17126_5147# 0 0.00271f
C1790 a_17307_5147# 0 0.167f
C1791 sar_retimer[7] 0 0.257f
C1792 a_17898_5147# 0 0.26f
C1793 x1[7].Q_N 0 0.114f
C1794 a_17425_5429# 0 0.00115f
C1795 a_16922_5147# 0 0.012f
C1796 a_16344_5147# 0 0.00291f
C1797 a_16550_5147# 0 0.191f
C1798 a_17103_5513# 0 7.41e-19
C1799 a_16875_5429# 0 0.00209f
C1800 a_16654_5429# 0 9.29e-19
C1801 a_14734_5147# 0 0.00178f
C1802 a_14915_5147# 0 0.157f
C1803 a_16320_5513# 0 7.05e-19
C1804 a_16143_5147# 0 0.109f
C1805 a_17017_5147# 0 0.272f
C1806 a_17191_5121# 0 0.487f
C1807 a_16704_5121# 0 0.433f
C1808 a_16236_5513# 0 0.281f
C1809 a_16410_5121# 0 0.296f
C1810 a_15955_5147# 0 0.585f
C1811 sar_logic[7] 0 1.71f
C1812 a_15789_5147# 0 0.544f
C1813 sar_retimer[6] 0 0.216f
C1814 a_15506_5147# 0 0.227f
C1815 x1[6].Q_N 0 0.101f
C1816 a_15033_5429# 0 0.00121f
C1817 a_14530_5147# 0 0.00861f
C1818 a_13952_5147# 0 0.00124f
C1819 a_14158_5147# 0 0.18f
C1820 a_14711_5513# 0 8.96e-19
C1821 a_14483_5429# 0 0.00223f
C1822 a_14262_5429# 0 0.00195f
C1823 a_13928_5513# 0 0.00146f
C1824 a_13751_5147# 0 0.102f
C1825 a_14625_5147# 0 0.257f
C1826 a_14799_5121# 0 0.453f
C1827 a_14312_5121# 0 0.368f
C1828 a_13844_5513# 0 0.275f
C1829 a_14018_5121# 0 0.299f
C1830 a_13563_5147# 0 0.425f
C1831 sar_logic[6] 0 0.186f
C1832 a_13397_5147# 0 0.597f
C1833 a_17425_5787# 0 1.82e-20
C1834 a_17103_5787# 0 5.79e-19
C1835 sar_retimer[5] 0 0.228f
C1836 x1[5].Q_N 0 0.107f
C1837 a_16875_5787# 0 0.00266f
C1838 a_16654_5787# 0 0.0011f
C1839 a_16320_5787# 0 7.93e-20
C1840 a_17307_6153# 0 0.168f
C1841 a_17126_6165# 0 0.00272f
C1842 a_16922_6109# 0 0.0118f
C1843 a_16550_6153# 0 0.186f
C1844 a_15033_5787# 0 0.0013f
C1845 a_14711_5787# 0 4.17e-19
C1846 a_16344_6165# 0 0.002f
C1847 a_16143_5787# 0 0.104f
C1848 sar_retimer[4] 0 0.17f
C1849 x1[4].Q_N 0 0.0929f
C1850 a_14483_5787# 0 0.00143f
C1851 a_13928_5787# 0 0.00102f
C1852 a_14915_6153# 0 0.156f
C1853 a_14734_6165# 0 0.00196f
C1854 a_14530_6109# 0 0.00926f
C1855 a_14158_6153# 0 0.183f
C1856 a_13952_6165# 0 0.00142f
C1857 a_13751_5787# 0 0.0996f
C1858 a_17898_5803# 0 0.245f
C1859 a_17017_6165# 0 0.256f
C1860 a_17191_5761# 0 0.452f
C1861 a_16704_5987# 0 0.386f
C1862 a_16236_5787# 0 0.266f
C1863 a_16410_5761# 0 0.286f
C1864 a_15955_5793# 0 0.532f
C1865 sar_logic[5] 0 1.62f
C1866 a_15789_5793# 0 0.483f
C1867 a_15506_5803# 0 0.219f
C1868 a_14625_6165# 0 0.244f
C1869 a_14799_5761# 0 0.426f
C1870 a_14312_5987# 0 0.327f
C1871 a_13844_5787# 0 0.261f
C1872 a_14018_5761# 0 0.276f
C1873 a_13563_5793# 0 0.386f
C1874 sar_logic[4] 0 0.164f
C1875 a_13397_5793# 0 0.542f
C1876 a_17126_6427# 0 0.00266f
C1877 a_17307_6427# 0 0.168f
C1878 sar_retimer[3] 0 0.242f
C1879 a_17898_6427# 0 0.256f
C1880 x1[3].Q_N 0 0.112f
C1881 a_17425_6709# 0 6.16e-19
C1882 a_16922_6427# 0 0.0117f
C1883 a_16344_6427# 0 0.00228f
C1884 a_16550_6427# 0 0.188f
C1885 a_17103_6793# 0 4.96e-19
C1886 a_16875_6709# 0 0.00146f
C1887 a_16654_6709# 0 0.0015f
C1888 a_14734_6427# 0 0.00193f
C1889 a_14915_6427# 0 0.157f
C1890 a_16320_6793# 0 1.99e-19
C1891 a_16143_6427# 0 0.107f
C1892 a_17017_6427# 0 0.265f
C1893 a_17191_6401# 0 0.463f
C1894 a_16704_6401# 0 0.416f
C1895 a_16236_6793# 0 0.277f
C1896 a_16410_6401# 0 0.291f
C1897 a_15955_6427# 0 0.565f
C1898 sar_logic[3] 0 1.67f
C1899 a_15789_6427# 0 0.505f
C1900 sar_retimer[2] 0 0.196f
C1901 a_15506_6427# 0 0.225f
C1902 x1[2].Q_N 0 0.0981f
C1903 a_15033_6709# 0 0.00118f
C1904 a_14530_6427# 0 0.00927f
C1905 a_13952_6427# 0 0.00129f
C1906 a_14158_6427# 0 0.181f
C1907 a_14711_6793# 0 7.03e-19
C1908 a_14483_6709# 0 0.00226f
C1909 a_14262_6709# 0 0.00106f
C1910 a_13928_6793# 0 0.00141f
C1911 a_13751_6427# 0 0.102f
C1912 a_14625_6427# 0 0.254f
C1913 a_14799_6401# 0 0.441f
C1914 a_14312_6401# 0 0.356f
C1915 a_13844_6793# 0 0.268f
C1916 a_14018_6401# 0 0.284f
C1917 a_13563_6427# 0 0.418f
C1918 sar_logic[2] 0 0.18f
C1919 a_13397_6427# 0 0.567f
C1920 a_17425_7067# 0 6.19e-19
C1921 a_17103_7067# 0 5.37e-19
C1922 sar_retimer[1] 0 0.226f
C1923 x1[1].Q_N 0 0.114f
C1924 a_16875_7067# 0 0.0029f
C1925 a_16654_7067# 0 0.00134f
C1926 a_16320_7067# 0 3.15e-19
C1927 a_17307_7433# 0 0.167f
C1928 a_17126_7445# 0 0.00295f
C1929 a_16922_7389# 0 0.0129f
C1930 a_16550_7433# 0 0.189f
C1931 a_15033_7067# 0 7.46e-19
C1932 a_14711_7067# 0 6.03e-19
C1933 a_16344_7445# 0 0.00263f
C1934 a_16143_7067# 0 0.104f
C1935 sar_retimer[0] 0 0.168f
C1936 x1[0].Q_N 0 0.0979f
C1937 a_14483_7067# 0 0.00321f
C1938 a_14262_7067# 0 5.48e-19
C1939 a_13928_7067# 0 0.00107f
C1940 a_14915_7433# 0 0.161f
C1941 a_14734_7445# 0 0.00207f
C1942 a_14530_7389# 0 0.0105f
C1943 a_14158_7433# 0 0.183f
C1944 a_13952_7445# 0 0.0013f
C1945 a_13751_7067# 0 0.101f
C1946 a_17898_7083# 0 0.256f
C1947 a_17017_7445# 0 0.266f
C1948 a_17191_7041# 0 0.47f
C1949 a_16704_7267# 0 0.401f
C1950 a_16236_7067# 0 0.275f
C1951 a_16410_7041# 0 0.297f
C1952 a_15955_7073# 0 0.55f
C1953 sar_logic[1] 0 1.68f
C1954 a_15789_7073# 0 0.504f
C1955 a_15506_7083# 0 0.219f
C1956 a_14625_7445# 0 0.255f
C1957 a_14799_7041# 0 0.453f
C1958 a_14312_7267# 0 0.346f
C1959 a_13844_7067# 0 0.266f
C1960 a_14018_7041# 0 0.288f
C1961 a_13563_7073# 0 0.4f
C1962 sar_logic[0] 0 0.169f
C1963 a_13397_7073# 0 0.565f
C1964 a_12385_8002# 0 0.00426f
C1965 a_12385_8140# 0 9.21e-19
C1966 a_12297_8002# 0 0.179f
C1967 a_12457_8140# 0 0.164f
C1968 a_12385_8278# 0 8.65e-19
C1969 a_12385_8416# 0 8.09e-19
C1970 a_12297_8278# 0 0.114f
C1971 a_12457_8416# 0 0.114f
C1972 a_12385_8554# 0 7.57e-19
C1973 a_12385_8692# 0 7.1e-19
C1974 a_12297_8554# 0 0.114f
C1975 a_12457_8692# 0 0.111f
C1976 a_12385_8830# 0 6.69e-19
C1977 a_12385_8968# 0 6.32e-19
C1978 a_12297_8830# 0 0.119f
C1979 a_18195_9015# 0 0.308f
C1980 x2.x2.floating 0 6.43f
C1981 x2.x3[1].floating 0 10.9f
C1982 x2.x4[3].floating 0 21.7f
C1983 x2.x7.floating 0 5.91f
C1984 x3.X 0 8.92f
C1985 delay_code[0] 0 3.75f
C1986 delay_code[1] 0 1.92f
C1987 delay_code[2] 0 1.96f
C1988 x2.x5[7].floating 0 0.107p
C1989 x2.x6.floating 0 0.412f
C1990 a_18499_9105# 0 0.359f
C1991 x3.A 0 0.587f
C1992 a_18195_9356# 0 0.275f
C1993 x2.x9.output_stack 0 1.52f
C1994 x2.x6.SW 0 0.299f
C1995 x2.x10.Y 0 2.76f
C1996 delay_offset 0 1.12f
C1997 a_12322_9805# 0 0.0147f
C1998 a_12410_9943# 0 0.0402f
C1999 a_12322_10081# 0 0.0815f
C2000 a_12410_10219# 0 0.032f
C2001 a_12322_10357# 0 0.0953f
C2002 x2.x5[7].floating.n0 0 -7.99f
C2003 x2.x5[7].floating.n1 0 -28.9f
C2004 x2.x5[7].floating.n2 0 3.83f
C2005 x2.x5[7].floating.n3 0 -7.07f
C2006 x2.x5[7].floating.n4 0 -28.3f
C2007 x2.x5[7].floating.n5 0 52.7f
C2008 x2.x5[7].floating.n6 0 -28.3f
C2009 x2.x5[7].floating.n7 0 -7.07f
C2010 x2.x5[7].floating.n8 0 3.83f
C2011 x2.x5[7].floating.n9 0 -28.9f
C2012 x2.x5[7].floating.n10 0 -8.01f
C2013 x2.x5[7].floating.n11 0 2.21f
C2014 x2.x5[7].floating.t5 0 0.859f
C2015 x2.x5[7].floating.n12 0 6.65f
C2016 x2.x5[7].floating.n13 0 1.21f
C2017 x2.x5[7].floating.n14 0 1.17f
C2018 x2.x5[7].floating.n15 0 2.18f
C2019 x2.x5[7].floating.n16 0 1.06f
C2020 x2.x5[7].floating.n17 0 0.366f
C2021 x2.x5[7].floating.n18 0 1.06f
C2022 x2.x5[7].floating.n19 0 2.8f
C2023 x2.x5[7].floating.n20 0 51.4f
C2024 x2.x5[7].floating.n21 0 2.79f
C2025 x2.x5[7].floating.n22 0 1.06f
C2026 x2.x5[7].floating.n23 0 0.364f
C2027 x2.x5[7].floating.t3 0 0.859f
C2028 x2.x5[7].floating.n24 0 6.48f
C2029 x2.x5[7].floating.n25 0 1.15f
C2030 x2.x5[7].floating.n26 0 1.36f
C2031 x2.x5[7].floating.n27 0 2.2f
C2032 x2.x5[7].floating.n28 0 1.06f
C2033 x2.x5[7].floating.n29 0 2.23f
C2034 x2.x5[7].floating.n30 0 -7.99f
C2035 x2.x5[7].floating.n31 0 -28.9f
C2036 x2.x5[7].floating.n32 0 3.83f
C2037 x2.x5[7].floating.n33 0 -7.07f
C2038 x2.x5[7].floating.n34 0 -28.3f
C2039 x2.x5[7].floating.n35 0 52.7f
C2040 x2.x5[7].floating.n36 0 -28.3f
C2041 x2.x5[7].floating.n37 0 -7.07f
C2042 x2.x5[7].floating.n38 0 3.83f
C2043 x2.x5[7].floating.n39 0 -28.9f
C2044 x2.x5[7].floating.n40 0 -8.01f
C2045 x2.x5[7].floating.n41 0 2.21f
C2046 x2.x5[7].floating.t6 0 0.859f
C2047 x2.x5[7].floating.n42 0 6.65f
C2048 x2.x5[7].floating.n43 0 1.21f
C2049 x2.x5[7].floating.n44 0 1.17f
C2050 x2.x5[7].floating.n45 0 2.18f
C2051 x2.x5[7].floating.n46 0 1.06f
C2052 x2.x5[7].floating.n47 0 0.366f
C2053 x2.x5[7].floating.n48 0 1.06f
C2054 x2.x5[7].floating.n49 0 2.8f
C2055 x2.x5[7].floating.n50 0 51.4f
C2056 x2.x5[7].floating.n51 0 2.79f
C2057 x2.x5[7].floating.n52 0 1.06f
C2058 x2.x5[7].floating.n53 0 0.364f
C2059 x2.x5[7].floating.t0 0 0.859f
C2060 x2.x5[7].floating.n54 0 6.48f
C2061 x2.x5[7].floating.n55 0 1.15f
C2062 x2.x5[7].floating.n56 0 1.36f
C2063 x2.x5[7].floating.n57 0 2.2f
C2064 x2.x5[7].floating.n58 0 1.06f
C2065 x2.x5[7].floating.n59 0 2.23f
C2066 x2.x5[7].floating.n60 0 -7.99f
C2067 x2.x5[7].floating.n61 0 -28.9f
C2068 x2.x5[7].floating.n62 0 3.83f
C2069 x2.x5[7].floating.n63 0 -7.07f
C2070 x2.x5[7].floating.n64 0 -28.3f
C2071 x2.x5[7].floating.n65 0 52.7f
C2072 x2.x5[7].floating.n66 0 -28.3f
C2073 x2.x5[7].floating.n67 0 -7.07f
C2074 x2.x5[7].floating.n68 0 3.83f
C2075 x2.x5[7].floating.n69 0 -28.9f
C2076 x2.x5[7].floating.n70 0 -8.01f
C2077 x2.x5[7].floating.n71 0 2.21f
C2078 x2.x5[7].floating.t7 0 0.859f
C2079 x2.x5[7].floating.n72 0 6.65f
C2080 x2.x5[7].floating.n73 0 1.21f
C2081 x2.x5[7].floating.n74 0 1.17f
C2082 x2.x5[7].floating.n75 0 2.18f
C2083 x2.x5[7].floating.n76 0 1.06f
C2084 x2.x5[7].floating.n77 0 0.366f
C2085 x2.x5[7].floating.n78 0 1.06f
C2086 x2.x5[7].floating.n79 0 2.8f
C2087 x2.x5[7].floating.n80 0 51.4f
C2088 x2.x5[7].floating.n81 0 2.79f
C2089 x2.x5[7].floating.n82 0 1.06f
C2090 x2.x5[7].floating.n83 0 0.364f
C2091 x2.x5[7].floating.t4 0 0.859f
C2092 x2.x5[7].floating.n84 0 6.48f
C2093 x2.x5[7].floating.n85 0 1.15f
C2094 x2.x5[7].floating.n86 0 1.36f
C2095 x2.x5[7].floating.n87 0 2.2f
C2096 x2.x5[7].floating.n88 0 1.06f
C2097 x2.x5[7].floating.n89 0 -15.2f
C2098 x2.x5[7].floating.n90 0 -15.2f
C2099 x2.x5[7].floating.n91 0 -41.6f
C2100 x2.x5[7].floating.n92 0 0.766f
C2101 x2.x5[7].floating.n93 0 2.47f
C2102 x2.x5[7].floating.n94 0 51.5f
C2103 x2.x5[7].floating.n95 0 2.47f
C2104 x2.x5[7].floating.n96 0 0.766f
C2105 x2.x5[7].floating.n97 0 -33.5f
C2106 x2.x5[7].floating.n98 0 -4.56f
C2107 x2.x5[7].floating.n99 0 3.83f
C2108 x2.x5[7].floating.n100 0 -28.9f
C2109 x2.x5[7].floating.n101 0 -7.07f
C2110 x2.x5[7].floating.n102 0 2.68f
C2111 x2.x5[7].floating.n103 0 52f
C2112 x2.x5[7].floating.n104 0 3.23f
C2113 x2.x5[7].floating.n105 0 -7.84f
C2114 x2.x5[7].floating.n106 0 -28.9f
C2115 x2.x5[7].floating.n107 0 3.83f
C2116 x2.x5[7].floating.n108 0 -5.01f
C2117 x2.x5[7].floating.n109 0 -33f
C2118 x2.x5[7].floating.n110 0 0.766f
C2119 x2.x5[7].floating.n111 0 2.47f
C2120 x2.x5[7].floating.n112 0 51.5f
C2121 x2.x5[7].floating.n113 0 2.47f
C2122 x2.x5[7].floating.n114 0 0.766f
C2123 x2.x5[7].floating.n115 0 -33.5f
C2124 x2.x5[7].floating.n116 0 -4.56f
C2125 x2.x5[7].floating.n117 0 3.83f
C2126 x2.x5[7].floating.n118 0 -28.9f
C2127 x2.x5[7].floating.n119 0 -7.07f
C2128 x2.x5[7].floating.n120 0 2.68f
C2129 x2.x5[7].floating.n121 0 52f
C2130 x2.x5[7].floating.n122 0 3.23f
C2131 x2.x5[7].floating.n123 0 -7.84f
C2132 x2.x5[7].floating.n124 0 -28.9f
C2133 x2.x5[7].floating.n125 0 3.83f
C2134 x2.x5[7].floating.n126 0 -5.01f
C2135 x2.x5[7].floating.n127 0 -33f
C2136 x2.x5[7].floating.n128 0 0.766f
C2137 x2.x5[7].floating.n129 0 2.47f
C2138 x2.x5[7].floating.n130 0 51.5f
C2139 x2.x5[7].floating.n131 0 2.47f
C2140 x2.x5[7].floating.n132 0 0.766f
C2141 x2.x5[7].floating.n133 0 -33.5f
C2142 x2.x5[7].floating.n134 0 -4.56f
C2143 x2.x5[7].floating.n135 0 3.83f
C2144 x2.x5[7].floating.n136 0 -28.9f
C2145 x2.x5[7].floating.n137 0 -7.07f
C2146 x2.x5[7].floating.n138 0 2.68f
C2147 x2.x5[7].floating.n139 0 52f
C2148 x2.x5[7].floating.n140 0 3.23f
C2149 x2.x5[7].floating.n141 0 2.23f
C2150 x2.x5[7].floating.t2 0 0.859f
C2151 x2.x5[7].floating.n142 0 6.48f
C2152 x2.x5[7].floating.n143 0 1.15f
C2153 x2.x5[7].floating.n144 0 1.36f
C2154 x2.x5[7].floating.n145 0 2.2f
C2155 x2.x5[7].floating.n146 0 1.06f
C2156 x2.x5[7].floating.n147 0 0.364f
C2157 x2.x5[7].floating.n148 0 1.06f
C2158 x2.x5[7].floating.n149 0 2.79f
C2159 x2.x5[7].floating.n150 0 51.4f
C2160 x2.x5[7].floating.n151 0 2.8f
C2161 x2.x5[7].floating.n152 0 1.06f
C2162 x2.x5[7].floating.n153 0 0.366f
C2163 x2.x5[7].floating.t1 0 0.859f
C2164 x2.x5[7].floating.n154 0 7.16f
C2165 x2.x5[7].floating.n155 0 1.21f
C2166 x2.x5[7].floating.n156 0 1.17f
C2167 x2.x5[7].floating.n157 0 1.67f
C2168 x2.x5[7].floating.n158 0 1.06f
C2169 x2.x5[7].floating.n159 0 -17.4f
C2170 x2.x5[7].floating.n160 0 -17.2f
C2171 x2.x5[7].floating.n161 0 -43.6f
C2172 x2.x5[7].floating.n162 0 0.766f
C2173 x2.x5[7].floating.n163 0 2.47f
C2174 x2.x5[7].floating.n164 0 51.5f
C2175 x2.x5[7].floating.n165 0 2.47f
C2176 x2.x5[7].floating.n166 0 0.766f
C2177 x2.x5[7].floating.n167 0 -33f
C2178 x2.x5[7].floating.n168 0 -5.01f
C2179 x2.x5[7].floating.n169 0 3.83f
C2180 x2.x5[7].floating.n170 0 -28.9f
C2181 x2.x5[7].floating.n171 0 -7.84f
C2182 x2.x10.Y.t0 0 0.0462f
C2183 x2.x10.Y.t5 0 0.0167f
C2184 x2.x10.Y.t2 0 0.0167f
C2185 x2.x10.Y.t9 0 0.0167f
C2186 x2.x10.Y.t3 0 0.0167f
C2187 x2.x10.Y.t6 0 0.0167f
C2188 x2.x10.Y.t4 0 0.0167f
C2189 x2.x10.Y.t7 0 0.0167f
C2190 x2.x10.Y.t8 0 0.0167f
C2191 x2.x10.Y.n0 0 0.222f
C2192 x2.x10.Y.n1 0 0.0366f
C2193 x2.x10.Y.t1 0 0.0174f
C2194 x2.x10.Y.n2 0 0.0188f
C2195 x2.x10.Y.n3 0 0.0186f
C2196 x2.x10.Y.n4 0 0.0151f
C2197 x2.x10.Y.n5 0 0.0211f
C2198 VDD.n0 0 0.00798f
C2199 VDD.t231 0 0.0192f
C2200 VDD.n1 0 0.00373f
C2201 VDD.n2 0 0.0047f
C2202 VDD.n3 0 0.0345f
C2203 VDD.n4 0 0.00527f
C2204 VDD.n5 0 9.66e-19
C2205 VDD.n6 0 0.00147f
C2206 VDD.n7 0 0.00806f
C2207 VDD.n8 0 0.0033f
C2208 VDD.n9 0 0.00167f
C2209 VDD.n10 0 0.00254f
C2210 VDD.n11 0 0.0026f
C2211 VDD.n12 0 0.00417f
C2212 VDD.n13 0 0.0026f
C2213 VDD.n14 0 3.08e-19
C2214 VDD.n15 0 0.00702f
C2215 VDD.n16 0 0.00643f
C2216 VDD.n17 0 0.00875f
C2217 VDD.n18 0 0.0154f
C2218 VDD.n19 0 0.00745f
C2219 VDD.n20 0 0.00602f
C2220 VDD.n21 0 0.00468f
C2221 VDD.n22 0 0.00113f
C2222 VDD.n23 0 0.0229f
C2223 VDD.n24 0 0.00468f
C2224 VDD.n25 0 0.0103f
C2225 VDD.n26 0 0.00154f
C2226 VDD.n27 0 0.00694f
C2227 VDD.t233 0 0.0192f
C2228 VDD.n28 0 0.0212f
C2229 VDD.n29 0 0.635f
C2230 VDD.n30 0 0.00966f
C2231 VDD.t172 0 0.387f
C2232 VDD.t0 0 0.164f
C2233 VDD.t129 0 0.162f
C2234 VDD.n31 0 0.221f
C2235 VDD.n32 0 5.57e-19
C2236 VDD.t187 0 0.533f
C2237 VDD.t235 0 0.483f
C2238 VDD.t173 0 0.608f
C2239 VDD.n33 0 0.298f
C2240 VDD.n35 0 0.00595f
C2241 VDD.n36 0 0.00617f
C2242 VDD.n37 0 0.0052f
C2243 VDD.n38 0 0.00755f
C2244 VDD.n39 0 0.139f
C2245 VDD.n40 0 0.0263f
C2246 VDD.n41 0 0.00424f
C2247 VDD.n42 0 0.016f
C2248 VDD.n43 0 0.0263f
C2249 VDD.n44 0 0.00424f
C2250 VDD.n45 0 0.016f
C2251 VDD.n46 0 0.0257f
C2252 VDD.n47 0 0.00424f
C2253 VDD.n48 0 0.00221f
C2254 VDD.n49 0 7.98e-19
C2255 VDD.n50 0 7.06e-19
C2256 VDD.n51 0 0.0263f
C2257 VDD.n52 0 0.00424f
C2258 VDD.n53 0 0.0151f
C2259 VDD.n54 0 0.0263f
C2260 VDD.n55 0 0.00424f
C2261 VDD.n56 0 0.016f
C2262 VDD.n57 0 0.00721f
C2263 VDD.n58 0 0.00654f
C2264 VDD.n59 0 0.0263f
C2265 VDD.n60 0 0.00424f
C2266 VDD.n61 0 0.00134f
C2267 VDD.n62 0 0.00295f
C2268 VDD.n63 0 0.00451f
C2269 VDD.n64 0 0.002f
C2270 VDD.n65 0 0.0108f
C2271 VDD.n66 0 0.0128f
C2272 VDD.n67 0 0.0114f
C2273 VDD.n68 0 0.0106f
C2274 VDD.n69 0 0.00565f
C2275 VDD.t166 0 0.0556f
C2276 VDD.n70 0 0.00562f
C2277 VDD.n71 0 0.0108f
C2278 VDD.t45 0 0.055f
C2279 VDD.n72 0 0.00565f
C2280 VDD.t170 0 0.0136f
C2281 VDD.t46 0 0.0136f
C2282 VDD.n73 0 0.0284f
C2283 VDD.n74 0 0.016f
C2284 VDD.t102 0 0.00296f
C2285 VDD.t167 0 0.00296f
C2286 VDD.n75 0 0.00613f
C2287 VDD.t75 0 0.00296f
C2288 VDD.t226 0 0.00296f
C2289 VDD.n76 0 0.00613f
C2290 VDD.n77 0 0.00904f
C2291 VDD.n78 0 0.0298f
C2292 VDD.n79 0 0.00188f
C2293 VDD.n80 0 0.0298f
C2294 VDD.n81 0 0.0165f
C2295 VDD.n82 0 0.0108f
C2296 VDD.n83 0 0.0108f
C2297 VDD.n84 0 0.00433f
C2298 VDD.t85 0 0.00531f
C2299 VDD.t258 0 0.00451f
C2300 VDD.n85 0 0.0125f
C2301 VDD.n86 0 0.0232f
C2302 VDD.n87 0 0.0383f
C2303 VDD.n88 0 0.02f
C2304 VDD.n89 0 0.0194f
C2305 VDD.n90 0 0.00568f
C2306 VDD.n91 0 0.00562f
C2307 VDD.t168 0 0.055f
C2308 VDD.n92 0 0.00565f
C2309 VDD.t163 0 -0.0014f
C2310 VDD.t169 0 0.00439f
C2311 VDD.n93 0 0.0202f
C2312 VDD.t149 0 -0.0014f
C2313 VDD.t225 0 0.00439f
C2314 VDD.n94 0 0.0202f
C2315 VDD.n95 0 0.0445f
C2316 VDD.n96 0 0.0568f
C2317 VDD.t148 0 0.129f
C2318 VDD.n97 0 0.0608f
C2319 VDD.n98 0 0.0218f
C2320 VDD.n99 0 0.0479f
C2321 VDD.n100 0 0.0114f
C2322 VDD.n101 0 0.00999f
C2323 VDD.n102 0 0.0109f
C2324 VDD.n103 0 0.0234f
C2325 VDD.n104 0 0.031f
C2326 VDD.n105 0 0.0216f
C2327 VDD.n106 0 0.00568f
C2328 VDD.n107 0 0.0801f
C2329 VDD.n108 0 0.0879f
C2330 VDD.t164 0 0.055f
C2331 VDD.n109 0 0.0993f
C2332 VDD.n110 0 0.0741f
C2333 VDD.t86 0 0.0544f
C2334 VDD.n111 0 0.058f
C2335 VDD.n112 0 0.00562f
C2336 VDD.n113 0 0.00127f
C2337 VDD.t165 0 -0.00262f
C2338 VDD.t116 0 0.00474f
C2339 VDD.n114 0 0.0186f
C2340 VDD.t224 0 -0.00262f
C2341 VDD.t87 0 0.00474f
C2342 VDD.n115 0 0.0186f
C2343 VDD.n116 0 0.0232f
C2344 VDD.n117 0 0.0222f
C2345 VDD.n118 0 0.0062f
C2346 VDD.n119 0 0.00295f
C2347 VDD.n120 0 0.0116f
C2348 VDD.n121 0 0.0234f
C2349 VDD.n122 0 0.0303f
C2350 VDD.n123 0 0.0203f
C2351 VDD.n124 0 0.0314f
C2352 VDD.n125 0 0.018f
C2353 VDD.n126 0 0.00562f
C2354 VDD.n127 0 0.0431f
C2355 VDD.t12 0 0.0544f
C2356 VDD.n128 0 0.0574f
C2357 VDD.t74 0 0.055f
C2358 VDD.n129 0 0.0646f
C2359 VDD.n130 0 0.00568f
C2360 VDD.n131 0 0.00571f
C2361 VDD.n132 0 0.0664f
C2362 VDD.n133 0 0.0598f
C2363 VDD.t19 0 0.0544f
C2364 VDD.t216 0 0.104f
C2365 VDD.n134 0 0.00568f
C2366 VDD.n135 0 9.39e-19
C2367 VDD.t47 0 0.0538f
C2368 VDD.n136 0 0.00568f
C2369 VDD.t212 0 0.0112f
C2370 VDD.t171 0 0.00501f
C2371 VDD.n137 0 0.0175f
C2372 VDD.t28 0 0.0112f
C2373 VDD.t48 0 0.00501f
C2374 VDD.n138 0 0.0175f
C2375 VDD.n139 0 0.0426f
C2376 VDD.n140 0 0.0108f
C2377 VDD.n141 0 0.016f
C2378 VDD.n142 0 0.013f
C2379 VDD.n143 0 0.002f
C2380 VDD.n144 0 0.00451f
C2381 VDD.n145 0 0.00295f
C2382 VDD.n146 0 0.00134f
C2383 VDD.n147 0 0.00424f
C2384 VDD.n148 0 0.0263f
C2385 VDD.n149 0 0.00424f
C2386 VDD.n150 0 0.0263f
C2387 VDD.n151 0 0.00427f
C2388 VDD.t73 0 0.00769f
C2389 VDD.t250 0 0.00326f
C2390 VDD.n152 0 0.0156f
C2391 VDD.n153 0 0.00639f
C2392 VDD.n154 0 0.0201f
C2393 VDD.n155 0 7.06e-19
C2394 VDD.t107 0 0.00772f
C2395 VDD.t241 0 0.00326f
C2396 VDD.n156 0 0.0145f
C2397 VDD.n157 0 0.0012f
C2398 VDD.n158 0 0.00425f
C2399 VDD.n159 0 8.83e-19
C2400 VDD.n160 0 0.00167f
C2401 VDD.n161 0 0.00146f
C2402 VDD.n162 0 0.0103f
C2403 VDD.n163 0 0.0263f
C2404 VDD.n164 0 0.00921f
C2405 VDD.n165 0 0.03f
C2406 VDD.n166 0 0.00215f
C2407 VDD.n167 0 0.00312f
C2408 VDD.n168 0 0.00653f
C2409 VDD.n169 0 0.0885f
C2410 VDD.n170 0 0.0885f
C2411 VDD.n171 0 0.00713f
C2412 VDD.n172 0 0.016f
C2413 VDD.n173 0 0.026f
C2414 VDD.n174 0 0.0155f
C2415 VDD.n175 0 0.0108f
C2416 VDD.n176 0 0.00129f
C2417 VDD.n177 0 0.00295f
C2418 VDD.n178 0 0.00451f
C2419 VDD.n179 0 0.00451f
C2420 VDD.n180 0 0.00712f
C2421 VDD.n181 0 0.0065f
C2422 VDD.n182 0 0.0679f
C2423 VDD.n183 0 0.0679f
C2424 VDD.n184 0 0.00719f
C2425 VDD.n185 0 0.00763f
C2426 VDD.n186 0 0.00654f
C2427 VDD.n187 0 0.071f
C2428 VDD.n188 0 0.00323f
C2429 VDD.n189 0 0.00716f
C2430 VDD.n190 0 0.071f
C2431 VDD.n191 0 0.0263f
C2432 VDD.n192 0 0.0263f
C2433 VDD.n193 0 0.00424f
C2434 VDD.n194 0 0.00134f
C2435 VDD.n195 0 0.0241f
C2436 VDD.n196 0 0.00295f
C2437 VDD.n197 0 0.00297f
C2438 VDD.t81 0 0.00296f
C2439 VDD.t211 0 0.00281f
C2440 VDD.n198 0 0.00604f
C2441 VDD.t108 0 0.00296f
C2442 VDD.t30 0 0.00281f
C2443 VDD.n199 0 0.00604f
C2444 VDD.n200 0 0.016f
C2445 VDD.n201 0 0.00728f
C2446 VDD.n202 0 0.0323f
C2447 VDD.n203 0 0.00364f
C2448 VDD.n204 0 0.0101f
C2449 VDD.n205 0 0.0107f
C2450 VDD.n206 0 0.00565f
C2451 VDD.n207 0 0.00562f
C2452 VDD.t213 0 0.0514f
C2453 VDD.n208 0 0.0568f
C2454 VDD.n209 0 0.00571f
C2455 VDD.n210 0 0.0634f
C2456 VDD.t80 0 0.0556f
C2457 VDD.n211 0 0.0634f
C2458 VDD.t29 0 0.0544f
C2459 VDD.t127 0 0.055f
C2460 VDD.n212 0 0.00565f
C2461 VDD.n213 0 0.00951f
C2462 VDD.n214 0 0.0108f
C2463 VDD.n215 0 0.0108f
C2464 VDD.n216 0 0.00416f
C2465 VDD.n217 0 0.00123f
C2466 VDD.n218 0 0.026f
C2467 VDD.n219 0 0.00424f
C2468 VDD.n220 0 0.00653f
C2469 VDD.n221 0 0.0749f
C2470 VDD.n222 0 0.00123f
C2471 VDD.n223 0 0.016f
C2472 VDD.n224 0 0.0258f
C2473 VDD.n225 0 0.0151f
C2474 VDD.n226 0 0.00293f
C2475 VDD.n227 0 0.00715f
C2476 VDD.n228 0 0.0749f
C2477 VDD.n229 0 0.0263f
C2478 VDD.n230 0 0.0263f
C2479 VDD.n231 0 0.00424f
C2480 VDD.n232 0 0.00134f
C2481 VDD.n233 0 0.00295f
C2482 VDD.n234 0 0.00451f
C2483 VDD.n235 0 3.52e-19
C2484 VDD.n236 0 3.52e-19
C2485 VDD.t128 0 0.0072f
C2486 VDD.t197 0 0.0072f
C2487 VDD.n237 0 0.0358f
C2488 VDD.n238 0 0.016f
C2489 VDD.n239 0 0.0107f
C2490 VDD.n240 0 0.00176f
C2491 VDD.n241 0 0.00565f
C2492 VDD.n242 0 0.00568f
C2493 VDD.n243 0 0.0807f
C2494 VDD.n244 0 0.0867f
C2495 VDD.t218 0 0.055f
C2496 VDD.t49 0 0.0544f
C2497 VDD.n245 0 0.00562f
C2498 VDD.t219 0 0.00312f
C2499 VDD.t180 0 0.00312f
C2500 VDD.n246 0 0.00661f
C2501 VDD.t238 0 0.00312f
C2502 VDD.t182 0 0.00312f
C2503 VDD.n247 0 0.00661f
C2504 VDD.n248 0 0.0338f
C2505 VDD.n249 0 0.0106f
C2506 VDD.n250 0 0.0109f
C2507 VDD.t50 0 -0.0014f
C2508 VDD.t160 0 0.00439f
C2509 VDD.n251 0 0.0202f
C2510 VDD.t192 0 -0.0014f
C2511 VDD.t158 0 0.00439f
C2512 VDD.n252 0 0.0202f
C2513 VDD.n253 0 0.0444f
C2514 VDD.n254 0 0.00763f
C2515 VDD.n255 0 0.0303f
C2516 VDD.n256 0 5.87e-19
C2517 VDD.n257 0 0.0109f
C2518 VDD.n258 0 0.00571f
C2519 VDD.n259 0 0.0568f
C2520 VDD.t157 0 0.055f
C2521 VDD.t96 0 0.0538f
C2522 VDD.n260 0 0.00562f
C2523 VDD.n261 0 0.0196f
C2524 VDD.t154 0 -0.00262f
C2525 VDD.t118 0 0.00474f
C2526 VDD.n262 0 0.0186f
C2527 VDD.t161 0 -0.00262f
C2528 VDD.t97 0 0.00474f
C2529 VDD.n263 0 0.0186f
C2530 VDD.n264 0 0.0316f
C2531 VDD.n265 0 0.0319f
C2532 VDD.n266 0 0.029f
C2533 VDD.n267 0 0.00715f
C2534 VDD.n268 0 0.00305f
C2535 VDD.n270 0 7.98e-19
C2536 VDD.t117 0 0.00529f
C2537 VDD.t244 0 0.00455f
C2538 VDD.n271 0 0.0122f
C2539 VDD.n272 0 0.0028f
C2540 VDD.n273 0 7.06e-19
C2541 VDD.n274 0 0.00166f
C2542 VDD.n275 0 0.00216f
C2543 VDD.n276 0 0.0044f
C2544 VDD.n277 0 0.0107f
C2545 VDD.n278 0 0.0146f
C2546 VDD.n279 0 0.00428f
C2547 VDD.n280 0 0.0149f
C2548 VDD.n281 0 0.00424f
C2549 VDD.n282 0 0.00124f
C2550 VDD.n283 0 7.98e-19
C2551 VDD.t248 0 0.00458f
C2552 VDD.t95 0 0.00524f
C2553 VDD.n284 0 0.0122f
C2554 VDD.n285 0 0.0263f
C2555 VDD.n286 0 0.00424f
C2556 VDD.n287 0 0.0263f
C2557 VDD.n288 0 0.0187f
C2558 VDD.n289 0 0.0271f
C2559 VDD.n290 0 0.0137f
C2560 VDD.n291 0 0.00302f
C2561 VDD.n292 0 0.00653f
C2562 VDD.n293 0 0.126f
C2563 VDD.n294 0 0.126f
C2564 VDD.n295 0 0.00719f
C2565 VDD.n296 0 0.00424f
C2566 VDD.n297 0 0.00654f
C2567 VDD.n298 0 0.0802f
C2568 VDD.n299 0 0.0802f
C2569 VDD.n300 0 0.00719f
C2570 VDD.n301 0 0.0208f
C2571 VDD.n302 0 0.0175f
C2572 VDD.n303 0 0.016f
C2573 VDD.n304 0 0.00763f
C2574 VDD.n305 0 0.00654f
C2575 VDD.n306 0 0.0627f
C2576 VDD.n307 0 0.016f
C2577 VDD.n308 0 0.065f
C2578 VDD.n309 0 0.00718f
C2579 VDD.n310 0 0.00118f
C2580 VDD.n311 0 0.00294f
C2581 VDD.n312 0 0.00338f
C2582 VDD.n313 0 0.00286f
C2583 VDD.n314 0 7.06e-19
C2584 VDD.n315 0 0.00162f
C2585 VDD.n316 0 0.00197f
C2586 VDD.n317 0 0.00237f
C2587 VDD.n318 0 0.00652f
C2588 VDD.n319 0 0.0131f
C2589 VDD.n320 0 0.0162f
C2590 VDD.n321 0 0.0263f
C2591 VDD.n322 0 0.00424f
C2592 VDD.n323 0 0.016f
C2593 VDD.n324 0 0.00718f
C2594 VDD.n325 0 0.00654f
C2595 VDD.n326 0 0.0263f
C2596 VDD.n327 0 0.00424f
C2597 VDD.n328 0 0.016f
C2598 VDD.n329 0 0.0263f
C2599 VDD.n330 0 0.00424f
C2600 VDD.n332 0 0.00652f
C2601 VDD.n333 0 0.0052f
C2602 VDD.n334 0 0.0264f
C2603 VDD.n335 0 0.00951f
C2604 VDD.t193 0 0.0112f
C2605 VDD.t4 0 0.00501f
C2606 VDD.n336 0 0.0175f
C2607 VDD.t125 0 0.0112f
C2608 VDD.t33 0 0.00501f
C2609 VDD.n337 0 0.0175f
C2610 VDD.n338 0 0.042f
C2611 VDD.n339 0 0.00565f
C2612 VDD.n340 0 0.00565f
C2613 VDD.t198 0 0.055f
C2614 VDD.n341 0 0.00565f
C2615 VDD.n342 0 0.0108f
C2616 VDD.n343 0 0.0107f
C2617 VDD.t63 0 0.00296f
C2618 VDD.t159 0 0.00296f
C2619 VDD.n344 0 0.00613f
C2620 VDD.t92 0 0.00296f
C2621 VDD.t156 0 0.00296f
C2622 VDD.n345 0 0.00613f
C2623 VDD.n346 0 0.0313f
C2624 VDD.n347 0 0.00565f
C2625 VDD.n348 0 0.0222f
C2626 VDD.n349 0 0.0216f
C2627 VDD.n350 0 0.00565f
C2628 VDD.t1 0 0.055f
C2629 VDD.n351 0 0.0741f
C2630 VDD.n352 0 0.0999f
C2631 VDD.n353 0 0.00568f
C2632 VDD.t32 0 0.0136f
C2633 VDD.t2 0 0.0136f
C2634 VDD.n354 0 0.0284f
C2635 VDD.n355 0 0.0257f
C2636 VDD.n356 0 0.0181f
C2637 VDD.n357 0 0.00565f
C2638 VDD.n358 0 0.0431f
C2639 VDD.t147 0 0.055f
C2640 VDD.n359 0 0.0574f
C2641 VDD.t62 0 0.055f
C2642 VDD.n360 0 0.0598f
C2643 VDD.n361 0 0.0658f
C2644 VDD.t155 0 0.055f
C2645 VDD.n362 0 0.0646f
C2646 VDD.n363 0 0.00565f
C2647 VDD.n364 0 0.0126f
C2648 VDD.n365 0 0.0319f
C2649 VDD.n366 0 0.0163f
C2650 VDD.n367 0 0.0198f
C2651 VDD.n368 0 0.0209f
C2652 VDD.n369 0 0.0305f
C2653 VDD.n370 0 0.016f
C2654 VDD.n371 0 0.00295f
C2655 VDD.n372 0 0.002f
C2656 VDD.n373 0 0.00562f
C2657 VDD.t6 0 0.105f
C2658 VDD.n374 0 0.0861f
C2659 VDD.t124 0 0.0556f
C2660 VDD.n375 0 0.0628f
C2661 VDD.n376 0 0.00562f
C2662 VDD.n377 0 0.0107f
C2663 VDD.n378 0 0.0108f
C2664 VDD.n379 0 0.016f
C2665 VDD.n380 0 0.00451f
C2666 VDD.t114 0 0.00296f
C2667 VDD.t194 0 0.00281f
C2668 VDD.n381 0 0.00604f
C2669 VDD.t90 0 0.00296f
C2670 VDD.t123 0 0.00281f
C2671 VDD.n382 0 0.00604f
C2672 VDD.n383 0 0.0109f
C2673 VDD.n384 0 0.00565f
C2674 VDD.t89 0 0.0544f
C2675 VDD.t199 0 0.0562f
C2676 VDD.n385 0 0.00568f
C2677 VDD.n386 0 0.0107f
C2678 VDD.n387 0 0.0108f
C2679 VDD.n388 0 0.00538f
C2680 VDD.n389 0 0.0128f
C2681 VDD.t137 0 0.0072f
C2682 VDD.t131 0 0.0072f
C2683 VDD.n390 0 0.0287f
C2684 VDD.n391 0 0.00451f
C2685 VDD.n392 0 0.00295f
C2686 VDD.n393 0 0.00134f
C2687 VDD.n394 0 0.00424f
C2688 VDD.n395 0 0.0263f
C2689 VDD.n396 0 0.00424f
C2690 VDD.n397 0 0.00357f
C2691 VDD.n398 0 0.00451f
C2692 VDD.n399 0 0.00134f
C2693 VDD.n400 0 0.00424f
C2694 VDD.n401 0 0.0263f
C2695 VDD.n402 0 0.00424f
C2696 VDD.n403 0 0.00134f
C2697 VDD.n404 0 0.085f
C2698 VDD.n405 0 0.085f
C2699 VDD.n406 0 0.00717f
C2700 VDD.n407 0 0.00337f
C2701 VDD.n408 0 0.0121f
C2702 VDD.n409 0 0.00451f
C2703 VDD.n410 0 0.00295f
C2704 VDD.n411 0 0.00129f
C2705 VDD.n412 0 8.22e-19
C2706 VDD.n413 0 0.00505f
C2707 VDD.n414 0 0.00382f
C2708 VDD.n415 0 0.00297f
C2709 VDD.n416 0 0.00653f
C2710 VDD.n417 0 0.0885f
C2711 VDD.n418 0 0.00303f
C2712 VDD.n419 0 0.00716f
C2713 VDD.n420 0 0.0885f
C2714 VDD.n421 0 0.0263f
C2715 VDD.n422 0 0.00718f
C2716 VDD.n423 0 0.0828f
C2717 VDD.n424 0 0.0828f
C2718 VDD.n425 0 0.00654f
C2719 VDD.n426 0 0.00332f
C2720 VDD.n427 0 0.0114f
C2721 VDD.n428 0 0.0258f
C2722 VDD.n429 0 0.0203f
C2723 VDD.n430 0 0.0255f
C2724 VDD.n431 0 0.0106f
C2725 VDD.n432 0 0.00451f
C2726 VDD.n433 0 0.00134f
C2727 VDD.n434 0 0.00277f
C2728 VDD.n435 0 0.00652f
C2729 VDD.n436 0 0.0732f
C2730 VDD.n437 0 0.00328f
C2731 VDD.n438 0 0.00716f
C2732 VDD.n439 0 0.0732f
C2733 VDD.n440 0 0.0263f
C2734 VDD.n441 0 0.00746f
C2735 VDD.n442 0 0.00424f
C2736 VDD.n443 0 0.00134f
C2737 VDD.n444 0 0.0236f
C2738 VDD.n445 0 0.00295f
C2739 VDD.n446 0 0.0029f
C2740 VDD.n447 0 0.00986f
C2741 VDD.t162 0 0.00312f
C2742 VDD.t178 0 0.00312f
C2743 VDD.n448 0 0.00661f
C2744 VDD.t8 0 0.00312f
C2745 VDD.t181 0 0.00312f
C2746 VDD.n449 0 0.00661f
C2747 VDD.n450 0 0.0241f
C2748 VDD.n451 0 0.016f
C2749 VDD.n452 0 0.0107f
C2750 VDD.n453 0 0.00928f
C2751 VDD.n454 0 0.00565f
C2752 VDD.n455 0 0.0105f
C2753 VDD.n456 0 0.016f
C2754 VDD.n457 0 0.0173f
C2755 VDD.n458 0 0.002f
C2756 VDD.n459 0 0.00986f
C2757 VDD.n460 0 0.00568f
C2758 VDD.n461 0 0.0556f
C2759 VDD.t130 0 0.0544f
C2760 VDD.n462 0 0.00559f
C2761 VDD.n463 0 0.0807f
C2762 VDD.n464 0 0.0861f
C2763 VDD.t7 0 0.0556f
C2764 VDD.t177 0 0.0544f
C2765 VDD.n465 0 0.0502f
C2766 VDD.n466 0 0.00565f
C2767 VDD.n467 0 0.00129f
C2768 VDD.n468 0 0.0108f
C2769 VDD.n469 0 0.00468f
C2770 VDD.n470 0 0.00451f
C2771 VDD.n471 0 0.0113f
C2772 VDD.n472 0 0.00347f
C2773 VDD.n473 0 0.00717f
C2774 VDD.n474 0 0.255f
C2775 VDD.n475 0 0.0635f
C2776 VDD.n476 0 0.00653f
C2777 VDD.n477 0 0.00307f
C2778 VDD.n478 0 0.00312f
C2779 VDD.n479 0 0.0107f
C2780 VDD.n480 0 0.0103f
C2781 VDD.n481 0 0.0102f
C2782 VDD.n482 0 0.0257f
C2783 VDD.n483 0 0.016f
C2784 VDD.n484 0 0.00295f
C2785 VDD.n485 0 8.22e-19
C2786 VDD.n486 0 0.00129f
C2787 VDD.n487 0 0.00568f
C2788 VDD.n488 0 0.0502f
C2789 VDD.t5 0 0.0544f
C2790 VDD.n489 0 0.0718f
C2791 VDD.t122 0 0.0556f
C2792 VDD.n490 0 0.0634f
C2793 VDD.n491 0 0.00565f
C2794 VDD.n492 0 0.00352f
C2795 VDD.n493 0 0.0327f
C2796 VDD.n494 0 0.00728f
C2797 VDD.n495 0 0.002f
C2798 VDD.n496 0 0.00295f
C2799 VDD.n497 0 0.016f
C2800 VDD.n498 0 0.0286f
C2801 VDD.n499 0 0.0194f
C2802 VDD.n500 0 0.00562f
C2803 VDD.n501 0 0.0568f
C2804 VDD.t34 0 0.052f
C2805 VDD.t3 0 0.0526f
C2806 VDD.n502 0 0.058f
C2807 VDD.n503 0 0.0795f
C2808 VDD.n504 0 0.00571f
C2809 VDD.n505 0 0.0166f
C2810 VDD.n506 0 0.0109f
C2811 VDD.n507 0 0.0255f
C2812 VDD.n508 0 0.00363f
C2813 VDD.n509 0 0.0108f
C2814 VDD.n510 0 0.00451f
C2815 VDD.t91 0 0.00769f
C2816 VDD.t251 0 0.00326f
C2817 VDD.n511 0 0.0156f
C2818 VDD.n512 0 0.00639f
C2819 VDD.n513 0 0.0201f
C2820 VDD.n514 0 7.06e-19
C2821 VDD.t88 0 0.00772f
C2822 VDD.t245 0 0.00326f
C2823 VDD.n515 0 0.0145f
C2824 VDD.n516 0 0.0012f
C2825 VDD.n517 0 0.00425f
C2826 VDD.n518 0 8.83e-19
C2827 VDD.n519 0 0.00167f
C2828 VDD.n520 0 0.00146f
C2829 VDD.n521 0 0.0103f
C2830 VDD.n522 0 0.0264f
C2831 VDD.n523 0 0.00927f
C2832 VDD.n524 0 0.04f
C2833 VDD.n525 0 0.00244f
C2834 VDD.n526 0 0.0027f
C2835 VDD.n527 0 0.00713f
C2836 VDD.n528 0 0.0797f
C2837 VDD.n529 0 0.0798f
C2838 VDD.n530 0 0.00654f
C2839 VDD.n531 0 0.00763f
C2840 VDD.n532 0 0.00719f
C2841 VDD.n533 0 0.0425f
C2842 VDD.n534 0 0.00288f
C2843 VDD.n535 0 2.1e-19
C2844 VDD.n536 0 0.00254f
C2845 VDD.n537 0 7.06e-19
C2846 VDD.n538 0 0.0012f
C2847 VDD.t253 0 0.00323f
C2848 VDD.t113 0 0.00758f
C2849 VDD.n539 0 0.00998f
C2850 VDD.n540 0 0.00485f
C2851 VDD.n541 0 0.00101f
C2852 VDD.n542 0 0.00101f
C2853 VDD.n543 0 0.00214f
C2854 VDD.n544 0 0.0012f
C2855 VDD.n545 0 0.0197f
C2856 VDD.n546 0 0.0557f
C2857 VDD.n547 0 0.00143f
C2858 VDD.t257 0 0.00322f
C2859 VDD.n548 0 0.00481f
C2860 VDD.n549 0 0.00215f
C2861 VDD.n550 0 0.00115f
C2862 VDD.t61 0 0.00742f
C2863 VDD.n551 0 0.00939f
C2864 VDD.n552 0 0.00101f
C2865 VDD.n553 0 0.00115f
C2866 VDD.n554 0 0.00366f
C2867 VDD.n555 0 5.09e-19
C2868 VDD.n556 0 0.00359f
C2869 VDD.n557 0 0.00118f
C2870 VDD.n558 0 0.00113f
C2871 VDD.n559 0 0.00424f
C2872 VDD.n560 0 0.0302f
C2873 VDD.n561 0 0.056f
C2874 VDD.n562 0 0.0539f
C2875 VDD.n563 0 0.00654f
C2876 VDD.n564 0 0.00763f
C2877 VDD.n565 0 0.00719f
C2878 VDD.n566 0 0.0845f
C2879 VDD.n567 0 0.0846f
C2880 VDD.n568 0 0.00649f
C2881 VDD.n569 0 0.00736f
C2882 VDD.n570 0 0.016f
C2883 VDD.n571 0 0.0189f
C2884 VDD.n572 0 0.0237f
C2885 VDD.n573 0 0.0222f
C2886 VDD.n574 0 0.026f
C2887 VDD.n575 0 0.00127f
C2888 VDD.n576 0 0.00562f
C2889 VDD.n577 0 0.058f
C2890 VDD.t153 0 0.0556f
C2891 VDD.n578 0 0.0885f
C2892 VDD.n579 0 0.0795f
C2893 VDD.n580 0 0.00568f
C2894 VDD.n581 0 0.0108f
C2895 VDD.n582 0 0.0108f
C2896 VDD.n583 0 0.0225f
C2897 VDD.n584 0 0.016f
C2898 VDD.n585 0 0.0173f
C2899 VDD.n586 0 0.021f
C2900 VDD.n587 0 0.00565f
C2901 VDD.n588 0 0.0741f
C2902 VDD.t179 0 0.055f
C2903 VDD.n589 0 0.0502f
C2904 VDD.n590 0 0.00565f
C2905 VDD.n591 0 0.0106f
C2906 VDD.n592 0 0.0107f
C2907 VDD.n593 0 0.00225f
C2908 VDD.n594 0 0.00333f
C2909 VDD.n595 0 0.00717f
C2910 VDD.n596 0 0.0754f
C2911 VDD.n597 0 0.0753f
C2912 VDD.n598 0 0.00652f
C2913 VDD.n599 0 0.00231f
C2914 VDD.n600 0 0.016f
C2915 VDD.n601 0 0.00416f
C2916 VDD.n602 0 0.0108f
C2917 VDD.n603 0 0.0108f
C2918 VDD.n604 0 0.00565f
C2919 VDD.n605 0 0.0556f
C2920 VDD.t20 0 0.055f
C2921 VDD.n606 0 0.0502f
C2922 VDD.t217 0 0.0544f
C2923 VDD.n607 0 0.0718f
C2924 VDD.n608 0 0.00559f
C2925 VDD.n609 0 0.002f
C2926 VDD.n610 0 0.0107f
C2927 VDD.n611 0 0.00382f
C2928 VDD.n612 0 0.00451f
C2929 VDD.n613 0 0.0121f
C2930 VDD.n614 0 0.00337f
C2931 VDD.n615 0 0.00717f
C2932 VDD.n616 0 0.0653f
C2933 VDD.n617 0 0.0653f
C2934 VDD.n618 0 0.00653f
C2935 VDD.n619 0 0.00312f
C2936 VDD.n620 0 0.00295f
C2937 VDD.n621 0 0.0108f
C2938 VDD.n622 0 0.0105f
C2939 VDD.n623 0 0.0267f
C2940 VDD.n624 0 0.0203f
C2941 VDD.n625 0 0.0108f
C2942 VDD.n626 0 0.00505f
C2943 VDD.n627 0 0.00562f
C2944 VDD.n628 0 0.058f
C2945 VDD.n629 0 0.0783f
C2946 VDD.t27 0 0.0562f
C2947 VDD.n630 0 0.0861f
C2948 VDD.n631 0 0.00565f
C2949 VDD.n632 0 0.00556f
C2950 VDD.n633 0 0.0205f
C2951 VDD.n634 0 0.026f
C2952 VDD.n635 0 0.0265f
C2953 VDD.n636 0 0.0103f
C2954 VDD.n637 0 0.0108f
C2955 VDD.n638 0 0.00312f
C2956 VDD.n639 0 0.00323f
C2957 VDD.n640 0 0.00716f
C2958 VDD.n641 0 0.0508f
C2959 VDD.n642 0 0.00292f
C2960 VDD.n643 0 0.00234f
C2961 VDD.n644 0 0.00245f
C2962 VDD.n645 0 7.06e-19
C2963 VDD.n646 0 0.0012f
C2964 VDD.t246 0 0.00323f
C2965 VDD.t79 0 0.00758f
C2966 VDD.n647 0 0.00998f
C2967 VDD.n648 0 0.00485f
C2968 VDD.n649 0 0.00101f
C2969 VDD.n650 0 0.00101f
C2970 VDD.n651 0 0.00214f
C2971 VDD.n652 0 0.0012f
C2972 VDD.n653 0 0.0198f
C2973 VDD.n654 0 6.56e-19
C2974 VDD.n655 0 9.21e-19
C2975 VDD.t256 0 0.00322f
C2976 VDD.n656 0 0.00481f
C2977 VDD.n657 0 0.00115f
C2978 VDD.t101 0 0.00742f
C2979 VDD.n658 0 0.00939f
C2980 VDD.n659 0 0.00101f
C2981 VDD.n660 0 0.00115f
C2982 VDD.n661 0 0.00366f
C2983 VDD.n662 0 0.00117f
C2984 VDD.n663 0 0.00314f
C2985 VDD.n664 0 0.00123f
C2986 VDD.n665 0 0.00123f
C2987 VDD.n666 0 0.00424f
C2988 VDD.n667 0 0.0386f
C2989 VDD.n668 0 0.04f
C2990 VDD.n669 0 0.0381f
C2991 VDD.n670 0 0.00654f
C2992 VDD.n671 0 0.00763f
C2993 VDD.n672 0 0.00719f
C2994 VDD.n673 0 0.0771f
C2995 VDD.n674 0 0.0771f
C2996 VDD.n675 0 0.00654f
C2997 VDD.n676 0 0.00763f
C2998 VDD.n677 0 0.00719f
C2999 VDD.n678 0 0.0263f
C3000 VDD.n679 0 0.0285f
C3001 VDD.n680 0 0.00652f
C3002 VDD.n681 0 0.00269f
C3003 VDD.n682 0 0.00299f
C3004 VDD.t239 0 0.00439f
C3005 VDD.n683 0 0.00566f
C3006 VDD.n684 0 0.00175f
C3007 VDD.t115 0 0.00526f
C3008 VDD.n685 0 0.00663f
C3009 VDD.n686 0 0.00175f
C3010 VDD.n687 0 0.00328f
C3011 VDD.n688 0 0.00285f
C3012 VDD.n689 0 0.00715f
C3013 VDD.n690 0 0.041f
C3014 VDD.n691 0 0.0386f
C3015 VDD.n692 0 0.00654f
C3016 VDD.n693 0 0.00763f
C3017 VDD.n694 0 0.00719f
C3018 VDD.n695 0 0.0841f
C3019 VDD.n696 0 0.0841f
C3020 VDD.n697 0 0.00654f
C3021 VDD.n698 0 0.00763f
C3022 VDD.n699 0 0.00719f
C3023 VDD.n700 0 0.234f
C3024 VDD.n701 0 0.0263f
C3025 VDD.n702 0 0.00424f
C3026 VDD.n703 0 0.016f
C3027 VDD.n704 0 0.0263f
C3028 VDD.n705 0 0.00424f
C3029 VDD.n706 0 0.016f
C3030 VDD.n707 0 0.0171f
C3031 VDD.n708 0 0.00424f
C3032 VDD.n709 0 0.00303f
C3033 VDD.n710 0 0.0109f
C3034 VDD.n711 0 0.0154f
C3035 VDD.n712 0 0.0705f
C3036 VDD.n713 0 0.00424f
C3037 VDD.t70 0 0.00531f
C3038 VDD.t243 0 0.00451f
C3039 VDD.n714 0 0.0125f
C3040 VDD.n715 0 0.0132f
C3041 VDD.n716 0 0.00715f
C3042 VDD.n717 0 0.0268f
C3043 VDD.n718 0 0.0179f
C3044 VDD.n719 0 0.016f
C3045 VDD.n720 0 0.0456f
C3046 VDD.t202 0 0.0136f
C3047 VDD.t222 0 0.0136f
C3048 VDD.n721 0 0.026f
C3049 VDD.n722 0 0.00565f
C3050 VDD.n723 0 0.00565f
C3051 VDD.t205 0 0.055f
C3052 VDD.n724 0 0.00565f
C3053 VDD.n725 0 0.0109f
C3054 VDD.n726 0 0.00565f
C3055 VDD.t36 0 -0.0014f
C3056 VDD.t229 0 0.00439f
C3057 VDD.n727 0 0.0202f
C3058 VDD.t152 0 -0.0014f
C3059 VDD.t208 0 0.00439f
C3060 VDD.n728 0 0.0202f
C3061 VDD.n729 0 5.87e-19
C3062 VDD.n730 0 0.0444f
C3063 VDD.n731 0 0.0474f
C3064 VDD.n732 0 0.0218f
C3065 VDD.n733 0 0.0607f
C3066 VDD.t35 0 0.128f
C3067 VDD.n734 0 0.0568f
C3068 VDD.t207 0 0.0556f
C3069 VDD.n735 0 0.0879f
C3070 VDD.n736 0 0.0795f
C3071 VDD.n737 0 0.00568f
C3072 VDD.n738 0 0.0216f
C3073 VDD.n739 0 0.0316f
C3074 VDD.n740 0 0.0166f
C3075 VDD.n741 0 0.0208f
C3076 VDD.t206 0 -0.00262f
C3077 VDD.t72 0 0.00474f
C3078 VDD.n742 0 0.0186f
C3079 VDD.t227 0 -0.00262f
C3080 VDD.t106 0 0.00474f
C3081 VDD.n743 0 0.0186f
C3082 VDD.n744 0 0.0265f
C3083 VDD.n745 0 0.0312f
C3084 VDD.n746 0 0.0206f
C3085 VDD.n747 0 0.00565f
C3086 VDD.n748 0 0.058f
C3087 VDD.t71 0 0.055f
C3088 VDD.n749 0 0.0741f
C3089 VDD.t65 0 0.055f
C3090 VDD.n750 0 0.00565f
C3091 VDD.n751 0 0.0108f
C3092 VDD.n752 0 0.0126f
C3093 VDD.n753 0 0.0128f
C3094 VDD.n754 0 0.00763f
C3095 VDD.n755 0 0.0225f
C3096 VDD.t94 0 0.00296f
C3097 VDD.t228 0 0.00296f
C3098 VDD.n756 0 0.00613f
C3099 VDD.t66 0 0.00296f
C3100 VDD.t210 0 0.00296f
C3101 VDD.n757 0 0.00613f
C3102 VDD.n758 0 0.0313f
C3103 VDD.n759 0 0.0216f
C3104 VDD.n760 0 0.00565f
C3105 VDD.n761 0 0.0646f
C3106 VDD.t209 0 0.055f
C3107 VDD.n762 0 0.0861f
C3108 VDD.n763 0 0.00565f
C3109 VDD.n764 0 0.0216f
C3110 VDD.n765 0 0.016f
C3111 VDD.n766 0 0.016f
C3112 VDD.t54 0 0.0112f
C3113 VDD.t223 0 0.00501f
C3114 VDD.n767 0 0.0175f
C3115 VDD.t196 0 0.0112f
C3116 VDD.t204 0 0.00501f
C3117 VDD.n768 0 0.0175f
C3118 VDD.n769 0 0.0427f
C3119 VDD.n770 0 0.00565f
C3120 VDD.t53 0 0.055f
C3121 VDD.n771 0 0.0628f
C3122 VDD.n772 0 0.00565f
C3123 VDD.n773 0 0.0159f
C3124 VDD.n774 0 0.0181f
C3125 VDD.n775 0 0.0317f
C3126 VDD.n776 0 0.00763f
C3127 VDD.n777 0 0.016f
C3128 VDD.t120 0 0.00296f
C3129 VDD.t52 0 0.00281f
C3130 VDD.n778 0 0.00604f
C3131 VDD.t100 0 0.00296f
C3132 VDD.t195 0 0.00281f
C3133 VDD.n779 0 0.00604f
C3134 VDD.n780 0 0.0339f
C3135 VDD.n781 0 0.0216f
C3136 VDD.n782 0 0.00565f
C3137 VDD.t99 0 0.055f
C3138 VDD.t57 0 0.055f
C3139 VDD.n783 0 0.00565f
C3140 VDD.n784 0 0.0216f
C3141 VDD.n785 0 0.0227f
C3142 VDD.n786 0 0.016f
C3143 VDD.t22 0 0.0072f
C3144 VDD.t221 0 0.0072f
C3145 VDD.n787 0 0.0108f
C3146 VDD.n788 0 0.00562f
C3147 VDD.n789 0 0.0556f
C3148 VDD.t21 0 0.055f
C3149 VDD.t175 0 0.055f
C3150 VDD.n790 0 0.00568f
C3151 VDD.n791 0 0.011f
C3152 VDD.t200 0 0.00312f
C3153 VDD.t185 0 0.00312f
C3154 VDD.n792 0 0.00661f
C3155 VDD.t135 0 0.00312f
C3156 VDD.t176 0 0.00312f
C3157 VDD.n793 0 0.00661f
C3158 VDD.n794 0 0.0339f
C3159 VDD.n795 0 0.0264f
C3160 VDD.n796 0 0.0102f
C3161 VDD.n797 0 0.00568f
C3162 VDD.n798 0 0.00451f
C3163 VDD.n799 0 0.00719f
C3164 VDD.n800 0 0.00252f
C3165 VDD.n801 0 0.00652f
C3166 VDD.n802 0 0.0263f
C3167 VDD.n803 0 0.00424f
C3168 VDD.n804 0 0.0263f
C3169 VDD.n805 0 0.00424f
C3170 VDD.n806 0 0.0263f
C3171 VDD.n807 0 0.0263f
C3172 VDD.n808 0 0.0072f
C3173 VDD.n809 0 0.0916f
C3174 VDD.t64 0 0.00769f
C3175 VDD.t260 0 0.00326f
C3176 VDD.n810 0 0.0156f
C3177 VDD.n811 0 0.00639f
C3178 VDD.n812 0 0.0202f
C3179 VDD.n813 0 7.06e-19
C3180 VDD.t98 0 0.00772f
C3181 VDD.t249 0 0.00326f
C3182 VDD.n814 0 0.0145f
C3183 VDD.n815 0 0.0012f
C3184 VDD.n816 0 0.00425f
C3185 VDD.n817 0 8.83e-19
C3186 VDD.n818 0 0.00167f
C3187 VDD.n819 0 0.00146f
C3188 VDD.n820 0 0.0104f
C3189 VDD.n821 0 0.0265f
C3190 VDD.n822 0 0.0193f
C3191 VDD.n823 0 0.00693f
C3192 VDD.n824 0 0.00424f
C3193 VDD.n825 0 0.025f
C3194 VDD.n826 0 0.0263f
C3195 VDD.n827 0 0.00424f
C3196 VDD.n828 0 0.00716f
C3197 VDD.n829 0 0.00323f
C3198 VDD.n830 0 0.00829f
C3199 VDD.n831 0 0.002f
C3200 VDD.n832 0 0.00295f
C3201 VDD.n833 0 0.00312f
C3202 VDD.n834 0 0.00451f
C3203 VDD.n835 0 0.00134f
C3204 VDD.n836 0 0.00312f
C3205 VDD.n837 0 0.00653f
C3206 VDD.n838 0 0.0679f
C3207 VDD.n839 0 0.00721f
C3208 VDD.n840 0 0.00654f
C3209 VDD.n841 0 0.00296f
C3210 VDD.n842 0 0.00218f
C3211 VDD.n843 0 0.00183f
C3212 VDD.n844 0 7.06e-19
C3213 VDD.n845 0 0.0012f
C3214 VDD.t255 0 0.00323f
C3215 VDD.t119 0 0.00758f
C3216 VDD.n846 0 0.00998f
C3217 VDD.n847 0 0.00485f
C3218 VDD.n848 0 0.00101f
C3219 VDD.n849 0 0.00101f
C3220 VDD.n850 0 0.00214f
C3221 VDD.n851 0 0.0012f
C3222 VDD.n852 0 0.0198f
C3223 VDD.n853 0 7.1e-19
C3224 VDD.n854 0 0.00131f
C3225 VDD.t240 0 0.00322f
C3226 VDD.n855 0 0.00481f
C3227 VDD.n856 0 0.00115f
C3228 VDD.t93 0 0.00742f
C3229 VDD.n857 0 0.00939f
C3230 VDD.n858 0 0.00101f
C3231 VDD.n859 0 0.00115f
C3232 VDD.n860 0 0.00357f
C3233 VDD.n861 0 3.44e-19
C3234 VDD.n862 0 0.00309f
C3235 VDD.n863 0 0.00129f
C3236 VDD.n864 0 0.00129f
C3237 VDD.n865 0 0.00424f
C3238 VDD.n866 0 0.0127f
C3239 VDD.n867 0 0.0163f
C3240 VDD.n868 0 0.0552f
C3241 VDD.n869 0 0.00719f
C3242 VDD.n870 0 0.00424f
C3243 VDD.n871 0 0.00654f
C3244 VDD.n872 0 0.0758f
C3245 VDD.n873 0 0.00716f
C3246 VDD.n874 0 0.0758f
C3247 VDD.n875 0 0.0263f
C3248 VDD.n876 0 0.0916f
C3249 VDD.n877 0 0.00652f
C3250 VDD.n878 0 0.00948f
C3251 VDD.n879 0 0.0257f
C3252 VDD.n880 0 0.00671f
C3253 VDD.n881 0 0.00715f
C3254 VDD.n882 0 0.00424f
C3255 VDD.n883 0 0.00654f
C3256 VDD.n884 0 0.0675f
C3257 VDD.n885 0 0.0675f
C3258 VDD.n886 0 0.00719f
C3259 VDD.n887 0 0.00424f
C3260 VDD.n888 0 0.00654f
C3261 VDD.n889 0 0.0903f
C3262 VDD.n890 0 0.0902f
C3263 VDD.n891 0 0.00719f
C3264 VDD.n892 0 0.00763f
C3265 VDD.n893 0 0.00654f
C3266 VDD.n894 0 0.139f
C3267 VDD.n895 0 0.139f
C3268 VDD.n896 0 0.00716f
C3269 VDD.n897 0 0.00763f
C3270 VDD.n898 0 0.00656f
C3271 VDD.n899 0 0.156f
C3272 VDD.n900 0 0.156f
C3273 VDD.n901 0 0.0263f
C3274 VDD.n902 0 0.00424f
C3275 VDD.n903 0 0.00134f
C3276 VDD.n904 0 0.0271f
C3277 VDD.n905 0 0.00295f
C3278 VDD.n906 0 0.00322f
C3279 VDD.n907 0 0.0108f
C3280 VDD.n908 0 0.0102f
C3281 VDD.n909 0 0.00562f
C3282 VDD.n910 0 0.00565f
C3283 VDD.n911 0 0.0102f
C3284 VDD.n912 0 0.0741f
C3285 VDD.t43 0 0.0556f
C3286 VDD.t58 0 -0.0014f
C3287 VDD.t146 0 0.00439f
C3288 VDD.n913 0 0.0202f
C3289 VDD.t44 0 -0.0014f
C3290 VDD.t16 0 0.00439f
C3291 VDD.n914 0 0.0202f
C3292 VDD.n915 0 0.0356f
C3293 VDD.n916 0 7.05e-19
C3294 VDD.n917 0 0.0107f
C3295 VDD.n918 0 0.00711f
C3296 VDD.n919 0 0.00295f
C3297 VDD.n920 0 0.016f
C3298 VDD.n921 0 0.0107f
C3299 VDD.n922 0 0.00562f
C3300 VDD.n923 0 0.0568f
C3301 VDD.t15 0 0.0538f
C3302 VDD.n924 0 0.0795f
C3303 VDD.n925 0 0.0993f
C3304 VDD.n926 0 0.00562f
C3305 VDD.t18 0 -0.00262f
C3306 VDD.t112 0 0.00474f
C3307 VDD.n927 0 0.0186f
C3308 VDD.t145 0 -0.00262f
C3309 VDD.t78 0 0.00474f
C3310 VDD.n928 0 0.0186f
C3311 VDD.n929 0 0.0265f
C3312 VDD.n930 0 0.0234f
C3313 VDD.n931 0 0.016f
C3314 VDD.n932 0 0.0185f
C3315 VDD.n933 0 0.0291f
C3316 VDD.n934 0 0.00451f
C3317 VDD.t111 0 0.00529f
C3318 VDD.t252 0 0.00455f
C3319 VDD.n935 0 0.0125f
C3320 VDD.n936 0 0.013f
C3321 VDD.n937 0 0.0339f
C3322 VDD.n938 0 0.00424f
C3323 VDD.n939 0 0.00656f
C3324 VDD.n940 0 0.0295f
C3325 VDD.t39 0 0.0136f
C3326 VDD.t59 0 0.0136f
C3327 VDD.n941 0 0.0109f
C3328 VDD.n942 0 0.00571f
C3329 VDD.t38 0 0.0544f
C3330 VDD.t13 0 0.0544f
C3331 VDD.n943 0 0.00559f
C3332 VDD.n944 0 0.0109f
C3333 VDD.t110 0 0.00296f
C3334 VDD.t144 0 0.00296f
C3335 VDD.n945 0 0.00613f
C3336 VDD.t84 0 0.00296f
C3337 VDD.t14 0 0.00296f
C3338 VDD.n946 0 0.00613f
C3339 VDD.n947 0 0.0108f
C3340 VDD.n948 0 0.0319f
C3341 VDD.n949 0 0.00763f
C3342 VDD.n950 0 0.0257f
C3343 VDD.n951 0 0.0216f
C3344 VDD.n952 0 0.00565f
C3345 VDD.n953 0 0.0652f
C3346 VDD.n954 0 0.0598f
C3347 VDD.t9 0 0.0556f
C3348 VDD.t141 0 0.105f
C3349 VDD.n955 0 0.00565f
C3350 VDD.t40 0 0.0532f
C3351 VDD.n956 0 0.00565f
C3352 VDD.t191 0 0.0112f
C3353 VDD.t41 0 0.00501f
C3354 VDD.n957 0 0.0175f
C3355 VDD.t24 0 0.0112f
C3356 VDD.t60 0 0.00501f
C3357 VDD.n958 0 0.0175f
C3358 VDD.n959 0 0.0427f
C3359 VDD.n960 0 0.0108f
C3360 VDD.n961 0 0.0166f
C3361 VDD.n962 0 0.0319f
C3362 VDD.n963 0 0.00763f
C3363 VDD.n964 0 0.0267f
C3364 VDD.t104 0 0.00296f
C3365 VDD.t190 0 0.00281f
C3366 VDD.n965 0 0.00604f
C3367 VDD.t69 0 0.00296f
C3368 VDD.t26 0 0.00281f
C3369 VDD.n966 0 0.00604f
C3370 VDD.n967 0 0.0339f
C3371 VDD.n968 0 0.00565f
C3372 VDD.t31 0 0.0514f
C3373 VDD.n969 0 0.0568f
C3374 VDD.t140 0 0.0544f
C3375 VDD.n970 0 0.00568f
C3376 VDD.n971 0 0.0143f
C3377 VDD.n972 0 0.0108f
C3378 VDD.n973 0 0.0212f
C3379 VDD.n974 0 0.016f
C3380 VDD.n975 0 0.0108f
C3381 VDD.n976 0 0.016f
C3382 VDD.t151 0 0.0072f
C3383 VDD.t214 0 0.0072f
C3384 VDD.n977 0 0.0106f
C3385 VDD.n978 0 0.00568f
C3386 VDD.n979 0 0.00562f
C3387 VDD.n980 0 0.0502f
C3388 VDD.t10 0 0.0562f
C3389 VDD.n981 0 0.0556f
C3390 VDD.t150 0 0.0544f
C3391 VDD.t183 0 0.0538f
C3392 VDD.n982 0 0.0281f
C3393 VDD.n983 0 0.00577f
C3394 VDD.n984 0 0.0107f
C3395 VDD.t139 0 0.00312f
C3396 VDD.t184 0 0.00312f
C3397 VDD.n985 0 0.00661f
C3398 VDD.t220 0 0.00312f
C3399 VDD.t186 0 0.00312f
C3400 VDD.n986 0 0.00661f
C3401 VDD.n987 0 0.0336f
C3402 VDD.n988 0 0.00451f
C3403 VDD.n989 0 0.00134f
C3404 VDD.n990 0 0.00424f
C3405 VDD.n991 0 0.0263f
C3406 VDD.n992 0 0.00424f
C3407 VDD.n993 0 0.0263f
C3408 VDD.n994 0 0.00424f
C3409 VDD.n995 0 0.0263f
C3410 VDD.n996 0 0.0263f
C3411 VDD.n997 0 0.00427f
C3412 VDD.n998 0 0.0263f
C3413 VDD.n999 0 0.0263f
C3414 VDD.n1000 0 0.00424f
C3415 VDD.n1001 0 0.024f
C3416 VDD.n1002 0 0.00424f
C3417 VDD.n1003 0 0.00118f
C3418 VDD.n1004 0 1.88e-19
C3419 VDD.n1005 0 0.00654f
C3420 VDD.n1006 0 0.0626f
C3421 VDD.n1007 0 0.0625f
C3422 VDD.n1008 0 0.00715f
C3423 VDD.n1009 0 0.00259f
C3424 VDD.n1010 0 0.00118f
C3425 VDD.n1011 0 7.51e-19
C3426 VDD.n1012 0 0.00323f
C3427 VDD.n1013 0 7.06e-19
C3428 VDD.t259 0 0.00439f
C3429 VDD.n1014 0 0.00566f
C3430 VDD.n1015 0 0.00175f
C3431 VDD.t76 0 0.00526f
C3432 VDD.n1016 0 0.00663f
C3433 VDD.n1017 0 0.00158f
C3434 VDD.n1018 0 0.00303f
C3435 VDD.n1019 0 0.00279f
C3436 VDD.n1020 0 0.00652f
C3437 VDD.n1021 0 0.0153f
C3438 VDD.n1022 0 0.00715f
C3439 VDD.n1023 0 0.0153f
C3440 VDD.n1024 0 0.0263f
C3441 VDD.n1025 0 0.0832f
C3442 VDD.n1026 0 0.0833f
C3443 VDD.n1027 0 0.00716f
C3444 VDD.n1028 0 0.0216f
C3445 VDD.n1029 0 0.0184f
C3446 VDD.n1030 0 0.016f
C3447 VDD.n1031 0 0.00763f
C3448 VDD.n1032 0 0.00656f
C3449 VDD.n1033 0 0.0421f
C3450 VDD.n1034 0 0.0443f
C3451 VDD.n1035 0 0.00721f
C3452 VDD.n1036 0 0.00129f
C3453 VDD.n1037 0 0.00129f
C3454 VDD.n1038 0 0.00311f
C3455 VDD.n1039 0 0.00297f
C3456 VDD.n1040 0 0.00192f
C3457 VDD.t242 0 0.00322f
C3458 VDD.n1041 0 0.00481f
C3459 VDD.n1042 0 0.00115f
C3460 VDD.t109 0 0.00742f
C3461 VDD.n1043 0 0.00939f
C3462 VDD.n1044 0 0.00101f
C3463 VDD.n1045 0 0.00115f
C3464 VDD.n1046 0 0.00358f
C3465 VDD.n1047 0 9.9e-19
C3466 VDD.n1048 0 7.06e-19
C3467 VDD.n1049 0 0.0012f
C3468 VDD.t262 0 0.00323f
C3469 VDD.t103 0 0.00758f
C3470 VDD.n1050 0 0.00998f
C3471 VDD.n1051 0 0.00485f
C3472 VDD.n1052 0 0.00101f
C3473 VDD.n1053 0 0.00101f
C3474 VDD.n1054 0 0.00214f
C3475 VDD.n1055 0 0.0012f
C3476 VDD.n1056 0 0.0198f
C3477 VDD.n1057 0 7.3e-19
C3478 VDD.n1058 0 7.15e-19
C3479 VDD.n1059 0 0.00219f
C3480 VDD.n1060 0 0.00654f
C3481 VDD.n1061 0 0.00424f
C3482 VDD.n1062 0 0.0377f
C3483 VDD.n1063 0 0.0499f
C3484 VDD.n1064 0 0.00719f
C3485 VDD.n1065 0 0.00424f
C3486 VDD.n1066 0 0.00654f
C3487 VDD.n1067 0 0.0859f
C3488 VDD.n1068 0 0.0859f
C3489 VDD.n1069 0 0.00718f
C3490 VDD.t82 0 0.00769f
C3491 VDD.t261 0 0.00326f
C3492 VDD.n1070 0 0.0156f
C3493 VDD.n1071 0 0.00639f
C3494 VDD.n1072 0 0.0201f
C3495 VDD.n1073 0 7.06e-19
C3496 VDD.t67 0 0.00772f
C3497 VDD.t254 0 0.00326f
C3498 VDD.n1074 0 0.0145f
C3499 VDD.n1075 0 0.0012f
C3500 VDD.n1076 0 0.00425f
C3501 VDD.n1077 0 8.83e-19
C3502 VDD.n1078 0 0.00167f
C3503 VDD.n1079 0 0.00146f
C3504 VDD.n1080 0 0.0104f
C3505 VDD.n1081 0 0.0266f
C3506 VDD.n1082 0 0.00963f
C3507 VDD.n1083 0 0.0252f
C3508 VDD.n1084 0 0.00533f
C3509 VDD.n1085 0 0.0222f
C3510 VDD.n1086 0 0.016f
C3511 VDD.n1087 0 0.00372f
C3512 VDD.n1088 0 0.00649f
C3513 VDD.n1089 0 0.0942f
C3514 VDD.n1090 0 0.0942f
C3515 VDD.n1091 0 0.00719f
C3516 VDD.n1092 0 0.00424f
C3517 VDD.n1093 0 0.00654f
C3518 VDD.n1094 0 0.0837f
C3519 VDD.n1095 0 0.0837f
C3520 VDD.n1096 0 0.00719f
C3521 VDD.n1097 0 0.016f
C3522 VDD.n1098 0 0.00763f
C3523 VDD.n1099 0 0.00654f
C3524 VDD.n1100 0 0.108f
C3525 VDD.n1101 0 0.108f
C3526 VDD.n1102 0 0.00716f
C3527 VDD.n1103 0 0.00763f
C3528 VDD.n1104 0 0.00656f
C3529 VDD.n1105 0 0.0854f
C3530 VDD.n1106 0 0.00176f
C3531 VDD.n1107 0 4.7e-19
C3532 VDD.n1108 0 0.00295f
C3533 VDD.n1109 0 0.00208f
C3534 VDD.n1110 0 0.00337f
C3535 VDD.n1111 0 0.00717f
C3536 VDD.n1112 0 0.326f
C3537 VDD.n1113 0 0.00772f
C3538 VDD.n1114 0 0.003f
C3539 VDD.n1115 0 0.0139f
C3540 VDD.n1116 0 0.0205f
C3541 VDD.n1117 0 0.02f
C3542 VDD.n1118 0 0.0271f
C3543 VDD.n1119 0 3.52e-19
C3544 VDD.n1120 0 0.0106f
C3545 VDD.n1121 0 0.00562f
C3546 VDD.n1122 0 0.0502f
C3547 VDD.t138 0 0.0556f
C3548 VDD.n1123 0 0.0861f
C3549 VDD.n1124 0 0.0801f
C3550 VDD.n1125 0 0.00556f
C3551 VDD.n1126 0 0.0464f
C3552 VDD.n1127 0 0.0293f
C3553 VDD.n1128 0 0.021f
C3554 VDD.n1129 0 0.0109f
C3555 VDD.n1130 0 0.0109f
C3556 VDD.n1131 0 0.0269f
C3557 VDD.n1132 0 0.0319f
C3558 VDD.n1133 0 0.0215f
C3559 VDD.n1134 0 0.00562f
C3560 VDD.n1135 0 0.0718f
C3561 VDD.t25 0 0.055f
C3562 VDD.n1136 0 0.0634f
C3563 VDD.t68 0 0.055f
C3564 VDD.n1137 0 0.0634f
C3565 VDD.n1138 0 0.00568f
C3566 VDD.n1139 0 0.0181f
C3567 VDD.n1140 0 0.0109f
C3568 VDD.n1141 0 0.0276f
C3569 VDD.n1142 0 0.016f
C3570 VDD.n1143 0 0.0203f
C3571 VDD.n1144 0 0.0157f
C3572 VDD.n1145 0 0.00562f
C3573 VDD.n1146 0 0.058f
C3574 VDD.n1147 0 0.0789f
C3575 VDD.t23 0 0.055f
C3576 VDD.n1148 0 0.0861f
C3577 VDD.n1149 0 0.00565f
C3578 VDD.n1150 0 0.00568f
C3579 VDD.n1151 0 0.0216f
C3580 VDD.n1152 0 0.0109f
C3581 VDD.n1153 0 0.0295f
C3582 VDD.n1154 0 0.016f
C3583 VDD.n1155 0 0.0184f
C3584 VDD.n1156 0 0.0197f
C3585 VDD.n1157 0 0.0311f
C3586 VDD.n1158 0 0.00176f
C3587 VDD.n1159 0 0.00565f
C3588 VDD.n1160 0 0.0646f
C3589 VDD.t83 0 0.0556f
C3590 VDD.n1161 0 0.0574f
C3591 VDD.t11 0 0.0556f
C3592 VDD.n1162 0 0.0431f
C3593 VDD.n1163 0 0.00565f
C3594 VDD.n1164 0 0.0074f
C3595 VDD.n1165 0 0.0282f
C3596 VDD.n1166 0 0.0273f
C3597 VDD.n1167 0 0.0245f
C3598 VDD.n1168 0 0.00867f
C3599 VDD.n1169 0 0.00352f
C3600 VDD.n1170 0 0.00167f
C3601 VDD.n1171 0 0.00132f
C3602 VDD.n1172 0 0.00728f
C3603 VDD.n1173 0 0.0189f
C3604 VDD.n1174 0 0.0265f
C3605 VDD.n1175 0 0.00565f
C3606 VDD.n1176 0 0.0741f
C3607 VDD.t77 0 0.055f
C3608 VDD.n1177 0 0.058f
C3609 VDD.t17 0 0.055f
C3610 VDD.n1178 0 0.0885f
C3611 VDD.n1179 0 0.00568f
C3612 VDD.n1180 0 0.002f
C3613 VDD.n1181 0 0.0108f
C3614 VDD.n1182 0 0.00208f
C3615 VDD.n1183 0 0.00451f
C3616 VDD.n1184 0 0.0139f
C3617 VDD.n1185 0 0.00313f
C3618 VDD.n1186 0 0.00716f
C3619 VDD.n1187 0 0.0802f
C3620 VDD.n1188 0 0.0802f
C3621 VDD.n1189 0 0.0263f
C3622 VDD.n1190 0 0.00424f
C3623 VDD.n1191 0 0.00134f
C3624 VDD.n1192 0 0.00382f
C3625 VDD.n1193 0 0.00884f
C3626 VDD.n1194 0 0.0166f
C3627 VDD.n1195 0 0.0197f
C3628 VDD.n1196 0 0.0214f
C3629 VDD.n1197 0 0.0187f
C3630 VDD.n1198 0 0.0319f
C3631 VDD.n1199 0 3.52e-19
C3632 VDD.n1200 0 0.0108f
C3633 VDD.n1201 0 0.00574f
C3634 VDD.n1202 0 0.0502f
C3635 VDD.t134 0 0.0562f
C3636 VDD.n1203 0 0.0861f
C3637 VDD.n1204 0 0.0795f
C3638 VDD.n1205 0 0.00556f
C3639 VDD.n1206 0 0.0479f
C3640 VDD.n1207 0 0.0215f
C3641 VDD.n1208 0 0.0319f
C3642 VDD.n1209 0 0.0319f
C3643 VDD.n1210 0 0.0216f
C3644 VDD.n1211 0 0.00565f
C3645 VDD.n1212 0 0.0502f
C3646 VDD.t133 0 0.055f
C3647 VDD.n1213 0 0.0718f
C3648 VDD.t51 0 0.055f
C3649 VDD.n1214 0 0.0634f
C3650 VDD.n1215 0 0.00565f
C3651 VDD.n1216 0 0.0143f
C3652 VDD.n1217 0 0.0251f
C3653 VDD.n1218 0 0.0317f
C3654 VDD.n1219 0 0.016f
C3655 VDD.n1220 0 0.0161f
C3656 VDD.n1221 0 0.0216f
C3657 VDD.n1222 0 0.00565f
C3658 VDD.n1223 0 0.0568f
C3659 VDD.t136 0 0.052f
C3660 VDD.t203 0 0.0532f
C3661 VDD.n1224 0 0.058f
C3662 VDD.n1225 0 0.0789f
C3663 VDD.n1226 0 0.00565f
C3664 VDD.n1227 0 0.0166f
C3665 VDD.n1228 0 0.0161f
C3666 VDD.n1229 0 0.0319f
C3667 VDD.n1230 0 0.0253f
C3668 VDD.n1231 0 0.0216f
C3669 VDD.n1232 0 0.00565f
C3670 VDD.t132 0 0.105f
C3671 VDD.t56 0 0.055f
C3672 VDD.n1233 0 0.0598f
C3673 VDD.n1234 0 0.0658f
C3674 VDD.n1235 0 0.00565f
C3675 VDD.n1236 0 0.0198f
C3676 VDD.n1237 0 0.0286f
C3677 VDD.n1238 0 0.016f
C3678 VDD.n1239 0 0.0192f
C3679 VDD.n1240 0 0.0265f
C3680 VDD.n1241 0 0.021f
C3681 VDD.n1242 0 0.00565f
C3682 VDD.n1243 0 0.0574f
C3683 VDD.t55 0 0.055f
C3684 VDD.n1244 0 0.0431f
C3685 VDD.t201 0 0.055f
C3686 VDD.n1245 0 0.0993f
C3687 VDD.n1246 0 0.00565f
C3688 VDD.n1247 0 0.0316f
C3689 VDD.n1248 0 0.0279f
C3690 VDD.n1249 0 0.016f
C3691 VDD.n1250 0 0.00529f
C3692 VDD.n1251 0 0.00654f
C3693 VDD.n1252 0 0.0697f
C3694 VDD.n1253 0 0.0131f
C3695 VDD.n1254 0 0.00652f
C3696 VDD.n1255 0 0.00273f
C3697 VDD.t247 0 0.00455f
C3698 VDD.t105 0 0.00529f
C3699 VDD.n1256 0 0.0122f
C3700 VDD.n1257 0 0.00346f
C3701 VDD.n1258 0 0.0017f
C3702 VDD.n1259 0 0.00234f
C3703 VDD.n1260 0 7.98e-19
C3704 VDD.n1261 0 0.00216f
C3705 VDD.n1262 0 0.00282f
C3706 VDD.n1263 0 0.00717f
C3707 VDD.n1264 0 0.0574f
C3708 VDD.n1265 0 0.0583f
C3709 VDD.n1266 0 0.00654f
C3710 VDD.n1267 0 0.00763f
C3711 VDD.n1268 0 0.00719f
C3712 VDD.n1269 0 0.0683f
C3713 VDD.n1270 0 0.0684f
C3714 VDD.n1271 0 0.00654f
C3715 VDD.n1272 0 0.00763f
C3716 VDD.n1273 0 0.00719f
C3717 VDD.n1274 0 0.951f
C3718 VDD.n1275 0 2.21f
C3719 VDD.n1276 0 1.15f
C3720 VDD.n1277 0 0.0041f
C3721 VDD.n1278 0 0.0177f
C3722 VDD.n1279 0 0.00751f
C3723 VDD.n1280 0 0.0336f
C3724 VDD.n1281 0 0.00239f
C3725 VDD.t142 0 0.101f
C3726 VDD.n1282 0 0.00384f
C3727 VDD.t143 0 0.0022f
C3728 VDD.n1283 0 0.00596f
C3729 VDD.n1284 0 0.00459f
C3730 VDD.n1285 0 0.0028f
C3731 VDD.n1286 0 0.00233f
C3732 VDD.n1287 0 0.01f
C3733 VDD.n1288 0 0.00184f
C3734 VDD.n1289 0 -0.0325f
C3735 VDD.n1290 0 1.23e-19
C3736 VDD.n1291 0 0.00131f
C3737 VDD.n1292 0 0.00178f
C3738 VDD.n1293 0 0.00101f
C3739 VDD.n1294 0 0.00101f
C3740 VDD.n1295 0 0.00114f
C3741 VDD.n1296 0 0.00104f
C3742 VDD.n1297 0 0.00654f
C3743 VDD.n1298 0 0.185f
C3744 VDD.n1299 0 0.00104f
C3745 VDD.n1300 0 0.00101f
C3746 VDD.n1301 0 0.00346f
C3747 VDD.n1302 0 0.00155f
C3748 VDD.n1303 0 0.00166f
C3749 VDD.n1304 0 0.00295f
C3750 VDD.n1305 0 0.00358f
C3751 VDD.n1306 0 0.00295f
C3752 VDD.n1307 0 0.00131f
C3753 VDD.n1308 0 0.00125f
C3754 VDD.n1309 0 0.00101f
C3755 VDD.n1310 0 0.00101f
C3756 VDD.n1311 0 0.00104f
C3757 VDD.n1312 0 0.00101f
C3758 VDD.n1313 0 0.00346f
C3759 VDD.n1314 0 0.00155f
C3760 VDD.n1315 0 -0.0284f
C3761 VDD.n1316 0 0.00358f
C3762 VDD.n1317 0 0.00295f
C3763 VDD.n1318 0 0.00131f
C3764 VDD.n1319 0 0.00125f
C3765 VDD.n1320 0 0.00101f
C3766 VDD.n1321 0 0.00101f
C3767 VDD.n1322 0 0.00104f
C3768 VDD.n1323 0 0.00101f
C3769 VDD.n1324 0 0.00346f
C3770 VDD.n1325 0 0.00155f
C3771 VDD.n1326 0 0.00166f
C3772 VDD.n1327 0 -0.0734f
C3773 VDD.n1328 0 0.00295f
C3774 VDD.n1329 0 0.00131f
C3775 VDD.n1330 0 0.00125f
C3776 VDD.n1331 0 0.00101f
C3777 VDD.n1332 0 0.00101f
C3778 VDD.n1333 0 0.00104f
C3779 VDD.n1334 0 0.00101f
C3780 VDD.n1335 0 0.00346f
C3781 VDD.n1336 0 0.00155f
C3782 VDD.n1337 0 0.00166f
C3783 VDD.n1338 0 0.00358f
C3784 VDD.n1339 0 0.00295f
C3785 VDD.n1340 0 0.00131f
C3786 VDD.n1341 0 0.00125f
C3787 VDD.n1342 0 0.00101f
C3788 VDD.n1343 0 0.00101f
C3789 VDD.n1345 0 0.00101f
C3790 VDD.n1346 0 0.00358f
C3791 VDD.n1347 0 0.00155f
C3792 VDD.n1348 0 -0.0284f
C3793 VDD.n1349 0 0.00218f
C3794 VDD.n1350 0 0.00166f
C3795 VDD.n1351 0 0.00125f
C3796 VDD.n1352 0 0.00101f
C3797 VDD.n1353 0 1.79e-19
C3798 VDD.n1354 0 0.00101f
C3799 VDD.n1355 0 1.02f
C3800 VDD.n1356 0 0.00104f
C3801 VDD.n1357 0 0.00101f
C3802 VDD.n1358 0 0.00346f
C3803 VDD.n1359 0 0.00155f
C3804 VDD.n1360 0 0.00166f
C3805 VDD.n1361 0 0.00295f
C3806 VDD.n1362 0 0.00345f
C3807 VDD.n1363 0 0.00295f
C3808 VDD.n1364 0 0.00131f
C3809 VDD.n1365 0 0.00125f
C3810 VDD.n1366 0 0.00101f
C3811 VDD.n1367 0 0.00101f
C3812 VDD.n1368 0 0.0037f
C3813 VDD.n1369 0 0.00393f
C3814 VDD.n1370 0 0.00101f
C3815 VDD.n1371 0 0.00101f
C3816 VDD.n1372 0 1.79e-19
C3817 VDD.n1373 0 0.0037f
C3818 VDD.n1374 0 0.00125f
C3819 VDD.n1375 0 0.0025f
C3820 VDD.n1376 0 0.00125f
C3821 VDD.n1377 0 0.00304f
C3822 VDD.n1378 0 -0.0284f
C3823 VDD.n1379 0 0.00345f
C3824 VDD.n1380 0 0.00184f
C3825 VDD.n1381 0 -0.0325f
C3826 VDD.n1382 0 1.23e-19
C3827 VDD.n1383 0 1.79e-19
C3828 VDD.n1384 0 0.00221f
C3829 VDD.n1385 0 0.00131f
C3830 VDD.n1386 0 0.00101f
C3831 VDD.n1387 0 0.00485f
C3832 VDD.n1388 0 0.0037f
C3833 VDD.n1389 0 0.00125f
C3834 VDD.n1390 0 0.00221f
C3835 VDD.n1391 0 0.00131f
C3836 VDD.n1392 0 1.79e-19
C3837 VDD.n1393 0 1.23e-19
C3838 VDD.n1394 0 0.00184f
C3839 VDD.n1395 0 0.00352f
C3840 VDD.n1396 0 -0.0284f
C3841 VDD.n1397 0 0.00155f
C3842 VDD.n1398 0 0.00131f
C3843 VDD.n1399 0 0.00346f
C3844 VDD.n1400 0 0.00101f
C3845 VDD.n1401 0 0.0037f
C3846 VDD.n1402 0 0.0037f
C3847 VDD.n1403 0 0.00101f
C3848 VDD.n1404 0 0.00101f
C3849 VDD.n1405 0 0.00101f
C3850 VDD.n1406 0 0.00101f
C3851 VDD.n1407 0 0.00131f
C3852 VDD.n1408 0 0.00125f
C3853 VDD.n1409 0 0.0107f
C3854 VDD.n1410 0 0.00218f
C3855 VDD.n1411 0 1.23e-19
C3856 VDD.n1412 0 0.00125f
C3857 VDD.n1413 0 0.00131f
C3858 VDD.n1414 0 0.00346f
C3859 VDD.n1415 0 0.00101f
C3860 VDD.n1416 0 0.00101f
C3861 VDD.n1417 0 0.0111f
C3862 VDD.n1418 0 0.00125f
C3863 VDD.n1419 0 0.00984f
C3864 VDD.n1420 0 0.0108f
C3865 VDD.n1421 0 0.0108f
C3866 VDD.n1422 0 0.00984f
C3867 VDD.n1423 0 0.00125f
C3868 VDD.n1424 0 0.0111f
C3869 VDD.n1425 0 0.00101f
C3870 VDD.n1427 0 0.00101f
C3871 VDD.n1428 0 0.00101f
C3872 VDD.n1429 0 0.00131f
C3873 VDD.n1430 0 0.00155f
C3874 VDD.n1431 0 0.00141f
C3875 VDD.n1432 0 0.00218f
C3876 VDD.n1433 0 1.23e-19
C3877 VDD.n1434 0 0.00125f
C3878 VDD.n1435 0 0.00346f
C3879 VDD.n1436 0 0.00101f
C3880 VDD.n1437 0 0.00393f
C3881 VDD.n1438 0 0.00101f
C3882 VDD.n1439 0 0.00101f
C3883 VDD.n1440 0 0.00131f
C3884 VDD.n1441 0 0.00155f
C3885 VDD.n1442 0 0.00141f
C3886 VDD.n1443 0 -0.035f
C3887 VDD.n1444 0 1.23e-19
C3888 VDD.n1445 0 0.00125f
C3889 VDD.n1446 0 0.00346f
C3890 VDD.n1447 0 0.0037f
C3891 VDD.n1448 0 0.00104f
C3892 VDD.n1449 0 0.00101f
C3893 VDD.n1450 0 0.00101f
C3894 VDD.n1451 0 0.00346f
C3895 VDD.n1452 0 1.79e-19
C3896 VDD.n1453 0 0.0037f
C3897 VDD.n1454 0 0.00125f
C3898 VDD.n1455 0 0.00155f
C3899 VDD.n1456 0 0.00141f
C3900 VDD.n1457 0 0.00218f
C3901 VDD.n1458 0 -0.0798f
C3902 VDD.n1459 0 0.00211f
C3903 VDD.n1460 0 0.00131f
C3904 VDD.n1461 0 0.00101f
C3905 VDD.n1462 0 0.00101f
C3906 VDD.n1463 0 0.00104f
C3907 VDD.n1464 0 0.00101f
C3908 VDD.n1465 0 0.00346f
C3909 VDD.n1466 0 0.00125f
C3910 VDD.n1467 0 1.23e-19
C3911 VDD.n1468 0 0.00141f
C3912 VDD.n1469 0 0.00345f
C3913 VDD.n1470 0 0.00141f
C3914 VDD.n1471 0 0.00131f
C3915 VDD.n1472 0 0.00101f
C3916 VDD.n1473 0 0.00101f
C3917 VDD.n1474 0 0.00104f
C3918 VDD.n1475 0 0.00101f
C3919 VDD.n1476 0 0.0111f
C3920 VDD.n1477 0 0.00125f
C3921 VDD.n1478 0 1.23e-19
C3922 VDD.n1479 0 0.00218f
C3923 VDD.n1480 0 0.00909f
C3924 VDD.n1481 0 0.00155f
C3925 VDD.n1482 0 0.00166f
C3926 VDD.n1483 0 -0.0735f
C3927 VDD.n1484 0 0.00295f
C3928 VDD.n1485 0 0.00131f
C3929 VDD.n1486 0 0.00125f
C3930 VDD.n1487 0 0.00101f
C3931 VDD.n1488 0 0.0111f
C3932 VDD.n1489 0 0.00101f
C3933 VDD.n1490 0 0.00101f
C3934 VDD.n1491 0 0.00104f
C3935 VDD.n1492 0 0.00101f
C3936 VDD.n1493 0 0.00346f
C3937 VDD.n1494 0 0.00155f
C3938 VDD.n1495 0 0.00166f
C3939 VDD.n1496 0 0.00345f
C3940 VDD.n1497 0 0.00295f
C3941 VDD.n1498 0 0.00131f
C3942 VDD.n1499 0 0.00125f
C3943 VDD.n1500 0 0.00101f
C3944 VDD.n1501 0 0.00101f
C3945 VDD.n1502 0 0.0037f
C3946 VDD.n1503 0 0.00393f
C3947 VDD.n1504 0 0.00101f
C3948 VDD.n1505 0 0.00101f
C3949 VDD.n1506 0 1.79e-19
C3950 VDD.n1507 0 0.0037f
C3951 VDD.n1508 0 0.00125f
C3952 VDD.n1509 0 0.0025f
C3953 VDD.n1510 0 0.00125f
C3954 VDD.n1511 0 0.00304f
C3955 VDD.n1512 0 -0.0284f
C3956 VDD.n1513 0 0.00345f
C3957 VDD.n1514 0 0.00184f
C3958 VDD.n1515 0 -0.0325f
C3959 VDD.n1516 0 1.23e-19
C3960 VDD.n1517 0 1.79e-19
C3961 VDD.n1518 0 0.00221f
C3962 VDD.n1519 0 0.00131f
C3963 VDD.n1520 0 0.00101f
C3964 VDD.n1521 0 0.00485f
C3965 VDD.n1522 0 0.0037f
C3966 VDD.n1523 0 0.00125f
C3967 VDD.n1524 0 0.00221f
C3968 VDD.n1525 0 0.00131f
C3969 VDD.n1526 0 1.79e-19
C3970 VDD.n1527 0 1.23e-19
C3971 VDD.n1528 0 0.00184f
C3972 VDD.n1529 0 0.00352f
C3973 VDD.n1530 0 -0.0284f
C3974 VDD.n1531 0 0.00155f
C3975 VDD.n1532 0 0.00131f
C3976 VDD.n1533 0 0.00346f
C3977 VDD.n1534 0 0.00101f
C3978 VDD.n1535 0 0.0037f
C3979 VDD.n1536 0 0.0037f
C3980 VDD.n1537 0 0.00101f
C3981 VDD.n1538 0 0.00101f
C3982 VDD.n1539 0 0.00101f
C3983 VDD.n1540 0 0.00101f
C3984 VDD.n1541 0 0.00131f
C3985 VDD.n1542 0 0.00125f
C3986 VDD.n1543 0 0.0107f
C3987 VDD.n1544 0 0.00218f
C3988 VDD.n1545 0 1.23e-19
C3989 VDD.n1546 0 0.00125f
C3990 VDD.n1547 0 0.00131f
C3991 VDD.n1548 0 0.00346f
C3992 VDD.n1549 0 0.00101f
C3993 VDD.n1550 0 0.00101f
C3994 VDD.n1551 0 0.0111f
C3995 VDD.n1552 0 0.00125f
C3996 VDD.n1553 0 0.00984f
C3997 VDD.n1554 0 0.0108f
C3998 VDD.n1555 0 0.0108f
C3999 VDD.n1556 0 0.00984f
C4000 VDD.n1557 0 0.00125f
C4001 VDD.n1558 0 0.0111f
C4002 VDD.n1559 0 0.00101f
C4003 VDD.n1561 0 0.00101f
C4004 VDD.n1562 0 0.00101f
C4005 VDD.n1563 0 0.00131f
C4006 VDD.n1564 0 0.00155f
C4007 VDD.n1565 0 0.00141f
C4008 VDD.n1566 0 0.00218f
C4009 VDD.n1567 0 1.23e-19
C4010 VDD.n1568 0 0.00125f
C4011 VDD.n1569 0 0.00346f
C4012 VDD.n1570 0 0.00101f
C4013 VDD.n1571 0 0.00393f
C4014 VDD.n1572 0 0.00101f
C4015 VDD.n1573 0 0.00101f
C4016 VDD.n1574 0 0.00131f
C4017 VDD.n1575 0 0.00155f
C4018 VDD.n1576 0 0.00141f
C4019 VDD.n1577 0 -0.035f
C4020 VDD.n1578 0 1.23e-19
C4021 VDD.n1579 0 0.00125f
C4022 VDD.n1580 0 0.00346f
C4023 VDD.n1581 0 0.0037f
C4024 VDD.n1582 0 0.00104f
C4025 VDD.n1583 0 0.00101f
C4026 VDD.n1584 0 0.00101f
C4027 VDD.n1585 0 0.00346f
C4028 VDD.n1586 0 1.79e-19
C4029 VDD.n1587 0 0.0037f
C4030 VDD.n1588 0 0.00125f
C4031 VDD.n1589 0 0.00155f
C4032 VDD.n1590 0 0.00141f
C4033 VDD.n1591 0 0.00218f
C4034 VDD.n1592 0 -0.0798f
C4035 VDD.n1593 0 0.00211f
C4036 VDD.n1594 0 0.00131f
C4037 VDD.n1595 0 0.00101f
C4038 VDD.n1596 0 0.00101f
C4039 VDD.n1597 0 0.00104f
C4040 VDD.n1598 0 0.00101f
C4041 VDD.n1599 0 0.00346f
C4042 VDD.n1600 0 0.00125f
C4043 VDD.n1601 0 1.23e-19
C4044 VDD.n1602 0 0.00141f
C4045 VDD.n1603 0 0.00345f
C4046 VDD.n1604 0 0.00141f
C4047 VDD.n1605 0 0.00131f
C4048 VDD.n1606 0 0.00101f
C4049 VDD.n1607 0 0.00101f
C4050 VDD.n1608 0 0.00104f
C4051 VDD.n1609 0 0.00101f
C4052 VDD.n1610 0 0.0111f
C4053 VDD.n1611 0 0.00125f
C4054 VDD.n1612 0 1.23e-19
C4055 VDD.n1613 0 0.00218f
C4056 VDD.n1614 0 0.00909f
C4057 VDD.n1615 0 0.00155f
C4058 VDD.n1616 0 0.00166f
C4059 VDD.n1617 0 -0.0735f
C4060 VDD.n1618 0 0.00295f
C4061 VDD.n1619 0 0.00131f
C4062 VDD.n1620 0 0.00125f
C4063 VDD.n1621 0 0.00101f
C4064 VDD.n1622 0 0.0111f
C4065 VDD.n1623 0 0.00101f
C4066 VDD.n1624 0 0.00101f
C4067 VDD.n1625 0 0.00104f
C4068 VDD.n1626 0 0.00101f
C4069 VDD.n1627 0 0.00346f
C4070 VDD.n1628 0 0.00155f
C4071 VDD.n1629 0 0.00166f
C4072 VDD.n1630 0 0.00345f
C4073 VDD.n1631 0 0.00295f
C4074 VDD.n1632 0 0.00131f
C4075 VDD.n1633 0 0.00125f
C4076 VDD.n1634 0 0.00101f
C4077 VDD.n1635 0 0.00101f
C4078 VDD.n1636 0 0.0037f
C4079 VDD.n1637 0 0.00393f
C4080 VDD.n1638 0 0.00101f
C4081 VDD.n1639 0 0.00101f
C4082 VDD.n1640 0 1.79e-19
C4083 VDD.n1641 0 0.0037f
C4084 VDD.n1642 0 0.00125f
C4085 VDD.n1643 0 0.0025f
C4086 VDD.n1644 0 0.00125f
C4087 VDD.n1645 0 0.00304f
C4088 VDD.n1646 0 -0.0284f
C4089 VDD.n1647 0 0.00345f
C4090 VDD.n1648 0 0.00184f
C4091 VDD.n1649 0 -0.0325f
C4092 VDD.n1650 0 1.23e-19
C4093 VDD.n1651 0 1.79e-19
C4094 VDD.n1652 0 0.00221f
C4095 VDD.n1653 0 0.00131f
C4096 VDD.n1654 0 0.00101f
C4097 VDD.n1655 0 0.00485f
C4098 VDD.n1656 0 0.0037f
C4099 VDD.n1657 0 0.00125f
C4100 VDD.n1658 0 0.00221f
C4101 VDD.n1659 0 0.00131f
C4102 VDD.n1660 0 1.79e-19
C4103 VDD.n1661 0 1.23e-19
C4104 VDD.n1662 0 0.00184f
C4105 VDD.n1663 0 0.00352f
C4106 VDD.n1664 0 -0.0284f
C4107 VDD.n1665 0 0.00155f
C4108 VDD.n1666 0 0.00131f
C4109 VDD.n1667 0 0.00346f
C4110 VDD.n1668 0 0.00101f
C4111 VDD.n1669 0 0.0037f
C4112 VDD.n1670 0 0.0037f
C4113 VDD.n1671 0 0.00101f
C4114 VDD.n1672 0 0.00101f
C4115 VDD.n1673 0 0.00101f
C4116 VDD.n1674 0 0.00101f
C4117 VDD.n1675 0 0.00131f
C4118 VDD.n1676 0 0.00125f
C4119 VDD.n1677 0 0.0107f
C4120 VDD.n1678 0 0.00218f
C4121 VDD.n1679 0 1.23e-19
C4122 VDD.n1680 0 0.00125f
C4123 VDD.n1681 0 0.00131f
C4124 VDD.n1682 0 0.00346f
C4125 VDD.n1683 0 0.00101f
C4126 VDD.n1684 0 0.00101f
C4127 VDD.n1685 0 0.0111f
C4128 VDD.n1686 0 0.00125f
C4129 VDD.n1687 0 0.00984f
C4130 VDD.n1688 0 0.0108f
C4131 VDD.n1689 0 0.0108f
C4132 VDD.n1690 0 0.00984f
C4133 VDD.n1691 0 0.00125f
C4134 VDD.n1692 0 0.0111f
C4135 VDD.n1693 0 0.00101f
C4136 VDD.n1695 0 0.00101f
C4137 VDD.n1696 0 0.00101f
C4138 VDD.n1697 0 0.00131f
C4139 VDD.n1698 0 0.00155f
C4140 VDD.n1699 0 0.00141f
C4141 VDD.n1700 0 0.00218f
C4142 VDD.n1701 0 1.23e-19
C4143 VDD.n1702 0 0.00125f
C4144 VDD.n1703 0 0.00346f
C4145 VDD.n1704 0 0.00101f
C4146 VDD.n1705 0 0.00393f
C4147 VDD.n1706 0 0.00101f
C4148 VDD.n1707 0 0.00101f
C4149 VDD.n1708 0 0.00131f
C4150 VDD.n1709 0 0.00155f
C4151 VDD.n1710 0 0.00141f
C4152 VDD.n1711 0 -0.035f
C4153 VDD.n1712 0 1.23e-19
C4154 VDD.n1713 0 0.00125f
C4155 VDD.n1714 0 0.00346f
C4156 VDD.n1715 0 0.0037f
C4157 VDD.n1716 0 0.00104f
C4158 VDD.n1717 0 0.00101f
C4159 VDD.n1718 0 0.00101f
C4160 VDD.n1719 0 0.00346f
C4161 VDD.n1720 0 1.79e-19
C4162 VDD.n1721 0 0.0037f
C4163 VDD.n1722 0 0.00125f
C4164 VDD.n1723 0 0.00155f
C4165 VDD.n1724 0 0.00141f
C4166 VDD.n1725 0 0.00218f
C4167 VDD.n1726 0 -0.0798f
C4168 VDD.n1727 0 0.00211f
C4169 VDD.n1728 0 0.00131f
C4170 VDD.n1729 0 0.00101f
C4171 VDD.n1730 0 0.00101f
C4172 VDD.n1731 0 0.00104f
C4173 VDD.n1732 0 0.00101f
C4174 VDD.n1733 0 0.00346f
C4175 VDD.n1734 0 0.00125f
C4176 VDD.n1735 0 1.23e-19
C4177 VDD.n1736 0 0.00141f
C4178 VDD.n1737 0 0.00345f
C4179 VDD.n1738 0 0.00141f
C4180 VDD.n1739 0 0.00131f
C4181 VDD.n1740 0 0.00101f
C4182 VDD.n1741 0 0.00101f
C4183 VDD.n1742 0 0.00104f
C4184 VDD.n1743 0 0.00101f
C4185 VDD.n1744 0 0.0111f
C4186 VDD.n1745 0 0.00125f
C4187 VDD.n1746 0 1.23e-19
C4188 VDD.n1747 0 0.00218f
C4189 VDD.n1748 0 0.00909f
C4190 VDD.n1749 0 0.00155f
C4191 VDD.n1750 0 0.00166f
C4192 VDD.n1751 0 -0.0735f
C4193 VDD.n1752 0 0.00295f
C4194 VDD.n1753 0 0.00131f
C4195 VDD.n1754 0 0.00125f
C4196 VDD.n1755 0 0.00101f
C4197 VDD.n1756 0 0.0111f
C4198 VDD.n1757 0 0.00101f
C4199 VDD.n1758 0 0.00101f
C4200 VDD.n1759 0 0.00104f
C4201 VDD.n1760 0 0.00101f
C4202 VDD.n1761 0 0.00346f
C4203 VDD.n1762 0 0.00155f
C4204 VDD.n1763 0 0.00166f
C4205 VDD.n1764 0 0.00345f
C4206 VDD.n1765 0 0.00295f
C4207 VDD.n1766 0 0.00131f
C4208 VDD.n1767 0 0.00125f
C4209 VDD.n1768 0 0.00101f
C4210 VDD.n1769 0 0.00101f
C4211 VDD.n1770 0 0.0037f
C4212 VDD.n1771 0 0.00393f
C4213 VDD.n1772 0 0.00101f
C4214 VDD.n1773 0 0.00101f
C4215 VDD.n1774 0 1.79e-19
C4216 VDD.n1775 0 0.0037f
C4217 VDD.n1776 0 0.00125f
C4218 VDD.n1777 0 0.0025f
C4219 VDD.n1778 0 0.00125f
C4220 VDD.n1779 0 0.00304f
C4221 VDD.n1780 0 -0.0284f
C4222 VDD.n1781 0 0.00345f
C4223 VDD.n1782 0 0.00184f
C4224 VDD.n1783 0 -0.0325f
C4225 VDD.n1784 0 1.23e-19
C4226 VDD.n1785 0 1.79e-19
C4227 VDD.n1786 0 0.00221f
C4228 VDD.n1787 0 0.00131f
C4229 VDD.n1788 0 0.00101f
C4230 VDD.n1789 0 0.00485f
C4231 VDD.n1790 0 0.0037f
C4232 VDD.n1791 0 0.00125f
C4233 VDD.n1792 0 0.00221f
C4234 VDD.n1793 0 0.00131f
C4235 VDD.n1794 0 1.79e-19
C4236 VDD.n1795 0 1.23e-19
C4237 VDD.n1796 0 0.00184f
C4238 VDD.n1797 0 0.00352f
C4239 VDD.n1798 0 -0.0284f
C4240 VDD.n1799 0 0.00155f
C4241 VDD.n1800 0 0.00131f
C4242 VDD.n1801 0 0.00346f
C4243 VDD.n1802 0 0.00101f
C4244 VDD.n1803 0 0.0037f
C4245 VDD.n1804 0 0.0037f
C4246 VDD.n1805 0 0.00101f
C4247 VDD.n1806 0 0.00101f
C4248 VDD.n1807 0 0.00101f
C4249 VDD.n1808 0 0.00101f
C4250 VDD.n1809 0 0.00131f
C4251 VDD.n1810 0 0.00125f
C4252 VDD.n1811 0 0.0107f
C4253 VDD.n1812 0 0.00218f
C4254 VDD.n1813 0 1.23e-19
C4255 VDD.n1814 0 0.00125f
C4256 VDD.n1815 0 0.00131f
C4257 VDD.n1816 0 0.00346f
C4258 VDD.n1817 0 0.00101f
C4259 VDD.n1818 0 0.00101f
C4260 VDD.n1819 0 0.0111f
C4261 VDD.n1820 0 0.00125f
C4262 VDD.n1821 0 0.00984f
C4263 VDD.n1822 0 0.0108f
C4264 VDD.n1823 0 0.0108f
C4265 VDD.n1824 0 0.00984f
C4266 VDD.n1825 0 0.00125f
C4267 VDD.n1826 0 0.0111f
C4268 VDD.n1827 0 0.00101f
C4269 VDD.n1829 0 0.00101f
C4270 VDD.n1830 0 0.00101f
C4271 VDD.n1831 0 0.00131f
C4272 VDD.n1832 0 0.00155f
C4273 VDD.n1833 0 0.00141f
C4274 VDD.n1834 0 0.00218f
C4275 VDD.n1835 0 1.23e-19
C4276 VDD.n1836 0 0.00125f
C4277 VDD.n1837 0 0.00346f
C4278 VDD.n1838 0 0.00101f
C4279 VDD.n1839 0 0.00393f
C4280 VDD.n1840 0 0.00101f
C4281 VDD.n1841 0 0.00101f
C4282 VDD.n1842 0 0.00131f
C4283 VDD.n1843 0 0.00155f
C4284 VDD.n1844 0 0.00141f
C4285 VDD.n1845 0 -0.035f
C4286 VDD.n1846 0 1.23e-19
C4287 VDD.n1847 0 0.00125f
C4288 VDD.n1848 0 0.00346f
C4289 VDD.n1849 0 0.0037f
C4290 VDD.n1850 0 0.00104f
C4291 VDD.n1851 0 0.00101f
C4292 VDD.n1852 0 0.00101f
C4293 VDD.n1853 0 0.00346f
C4294 VDD.n1854 0 1.79e-19
C4295 VDD.n1855 0 0.0037f
C4296 VDD.n1856 0 0.00125f
C4297 VDD.n1857 0 0.00155f
C4298 VDD.n1858 0 0.00141f
C4299 VDD.n1859 0 0.00218f
C4300 VDD.n1860 0 -0.0798f
C4301 VDD.n1861 0 0.00211f
C4302 VDD.n1862 0 0.00131f
C4303 VDD.n1863 0 0.00101f
C4304 VDD.n1864 0 0.00101f
C4305 VDD.n1866 0 0.00101f
C4306 VDD.n1867 0 0.00346f
C4307 VDD.n1868 0 0.00125f
C4308 VDD.n1869 0 1.23e-19
C4309 VDD.n1870 0 0.00141f
C4310 VDD.n1871 0 0.00345f
C4311 VDD.n1872 0 0.00141f
C4312 VDD.n1873 0 0.00131f
C4313 VDD.n1874 0 0.00101f
C4314 VDD.n1875 0 0.00101f
C4315 VDD.n1876 0 0.0147f
C4316 VDD.n1877 0 0.00125f
C4317 VDD.n1878 0 1.23e-19
C4318 VDD.n1879 0 0.00219f
C4319 VDD.n1880 0 0.015f
C4320 VDD.n1881 0 0.00166f
C4321 VDD.n1882 0 0.00211f
C4322 VDD.n1883 0 -0.035f
C4323 VDD.n1884 0 -0.0709f
C4324 VDD.n1885 0 0.00301f
C4325 VDD.n1886 0 0.00184f
C4326 VDD.n1887 0 1.79e-19
C4327 VDD.n1888 0 0.0159f
C4328 VDD.n1889 0 0.0195f
C4329 VDD.n1890 0 0.00764f
C4330 VDD.n1891 0 0.00104f
C4331 VDD.n1892 0 0.00485f
C4332 VDD.n1893 0 0.0037f
C4333 VDD.n1894 0 0.0037f
C4334 VDD.n1895 0 0.00125f
C4335 VDD.n1896 0 0.0025f
C4336 VDD.n1897 0 0.00304f
C4337 VDD.n1898 0 0.00155f
C4338 VDD.n1899 0 0.00221f
C4339 VDD.n1900 0 0.00178f
C4340 VDD.n1901 0 0.00166f
C4341 VDD.n1902 0 0.00211f
C4342 VDD.n1903 0 0.00218f
C4343 VDD.n1904 0 0.00345f
C4344 VDD.n1905 0 0.00352f
C4345 VDD.n1906 0 0.00301f
C4346 VDD.n1907 0 0.00184f
C4347 VDD.n1908 0 1.79e-19
C4348 VDD.n1909 0 0.00131f
C4349 VDD.n1910 0 1.19e-19
C4350 VDD.n1911 0 0.00393f
C4351 VDD.n1913 0 0.00485f
C4352 VDD.n1914 0 0.0037f
C4353 VDD.n1915 0 0.0037f
C4354 VDD.n1916 0 0.00125f
C4355 VDD.n1917 0 0.0025f
C4356 VDD.n1918 0 0.00304f
C4357 VDD.n1919 0 0.00221f
C4358 VDD.n1920 0 0.00155f
C4359 VDD.n1921 0 0.00125f
C4360 VDD.n1922 0 -0.0284f
C4361 VDD.n1923 0 1.23e-19
C4362 VDD.n1924 0 0.00184f
C4363 VDD.n1925 0 0.00301f
C4364 VDD.n1926 0 0.00352f
C4365 VDD.n1927 0 0.00345f
C4366 VDD.n1928 0 0.00211f
C4367 VDD.n1929 0 0.00166f
C4368 VDD.n1930 0 0.00178f
C4369 VDD.n1931 0 0.00221f
C4370 VDD.n1932 0 0.0025f
C4371 VDD.n1933 0 0.00304f
C4372 VDD.n1934 0 0.00131f
C4373 VDD.n1935 0 0.00101f
C4374 VDD.n1936 0 0.00131f
C4375 VDD.n1937 0 1.19e-19
C4376 VDD.n1938 0 0.00393f
C4377 VDD.n1939 0 0.00485f
C4378 VDD.n1941 0 0.00104f
C4379 VDD.n1942 0 0.00101f
C4380 VDD.n1943 0 1.19e-19
C4381 VDD.n1944 0 0.00131f
C4382 VDD.n1945 0 1.79e-19
C4383 VDD.n1946 0 0.00184f
C4384 VDD.n1947 0 0.00301f
C4385 VDD.n1948 0 -0.0709f
C4386 VDD.n1949 0 0.00345f
C4387 VDD.n1950 0 0.00211f
C4388 VDD.n1951 0 0.00166f
C4389 VDD.n1952 0 0.00178f
C4390 VDD.n1953 0 0.00221f
C4391 VDD.n1954 0 0.00304f
C4392 VDD.n1955 0 0.0025f
C4393 VDD.n1956 0 0.00125f
C4394 VDD.n1957 0 0.0037f
C4395 VDD.n1958 0 0.0037f
C4396 VDD.n1959 0 0.00485f
C4397 VDD.n1961 0 0.00104f
C4398 VDD.n1962 0 0.00393f
C4399 VDD.n1963 0 1.19e-19
C4400 VDD.n1964 0 0.00131f
C4401 VDD.n1965 0 1.79e-19
C4402 VDD.n1966 0 0.00184f
C4403 VDD.n1967 0 0.00301f
C4404 VDD.n1968 0 0.00352f
C4405 VDD.n1969 0 0.00345f
C4406 VDD.n1970 0 0.00211f
C4407 VDD.n1971 0 -0.0284f
C4408 VDD.n1972 0 -0.0798f
C4409 VDD.n1973 0 0.00221f
C4410 VDD.n1974 0 0.00304f
C4411 VDD.n1975 0 0.0025f
C4412 VDD.n1976 0 0.00125f
C4413 VDD.n1977 0 0.0037f
C4414 VDD.n1978 0 0.0037f
C4415 VDD.n1979 0 0.00485f
C4416 VDD.n1980 0 0.00104f
C4417 VDD.n1981 0 0.00883f
C4418 VDD.n1982 0 1.99e-19
C4419 VDD.n1983 0 0.00131f
C4420 VDD.n1984 0 1.79e-19
C4421 VDD.n1985 0 0.00184f
C4422 VDD.n1986 0 0.0108f
C4423 VDD.n1987 0 0.0125f
C4424 VDD.n1988 0 0.0124f
C4425 VDD.n1989 0 0.00218f
C4426 VDD.n1990 0 0.00211f
C4427 VDD.n1991 0 1.23e-19
C4428 VDD.n1992 0 0.00178f
C4429 VDD.n1993 0 1.79e-19
C4430 VDD.n1994 0 0.00131f
C4431 VDD.n1995 0 1.99e-19
C4432 VDD.n1996 0 0.00883f
C4433 VDD.n1997 0 0.00104f
C4434 VDD.n1998 0 0.00485f
C4435 VDD.n2001 0 0.00104f
C4436 VDD.n2002 0 0.00393f
C4437 VDD.n2003 0 1.19e-19
C4438 VDD.n2004 0 0.00101f
C4439 VDD.n2005 0 0.0037f
C4440 VDD.n2006 0 0.00125f
C4441 VDD.n2007 0 0.0025f
C4442 VDD.n2008 0 0.00304f
C4443 VDD.n2009 0 0.00221f
C4444 VDD.n2010 0 -0.0797f
C4445 VDD.n2011 0 0.00147f
C4446 VDD.n2012 0 0.00178f
C4447 VDD.n2013 0 0.00295f
C4448 VDD.n2014 0 0.00345f
C4449 VDD.n2015 0 0.00211f
C4450 VDD.n2016 0 -0.0735f
C4451 VDD.n2017 0 0.00178f
C4452 VDD.n2018 0 0.00295f
C4453 VDD.n2019 0 0.00147f
C4454 VDD.n2020 0 0.00352f
C4455 VDD.n2021 0 0.00218f
C4456 VDD.n2022 0 0.00166f
C4457 VDD.n2023 0 0.00125f
C4458 VDD.n2024 0 0.00155f
C4459 VDD.n2025 0 0.00346f
C4460 VDD.n2026 0 0.0025f
C4461 VDD.n2027 0 0.00304f
C4462 VDD.n2028 0 0.00131f
C4463 VDD.n2029 0 0.00101f
C4464 VDD.n2030 0 0.00101f
C4465 VDD.n2031 0 1.19e-19
C4466 VDD.n2032 0 0.00393f
C4467 VDD.n2034 0 0.00104f
C4468 VDD.n2036 0 0.00485f
C4469 VDD.n2037 0 0.0037f
C4470 VDD.n2038 0 0.0037f
C4471 VDD.n2039 0 0.00125f
C4472 VDD.n2040 0 0.00131f
C4473 VDD.n2041 0 0.00304f
C4474 VDD.n2042 0 0.0025f
C4475 VDD.n2043 0 0.00346f
C4476 VDD.n2044 0 0.00155f
C4477 VDD.n2045 0 0.00125f
C4478 VDD.n2046 0 0.00166f
C4479 VDD.n2047 0 0.00218f
C4480 VDD.n2048 0 0.00352f
C4481 VDD.n2049 0 0.00147f
C4482 VDD.n2050 0 0.00295f
C4483 VDD.n2051 0 0.00178f
C4484 VDD.n2052 0 1.23e-19
C4485 VDD.n2053 0 0.00211f
C4486 VDD.n2054 0 0.00218f
C4487 VDD.n2055 0 0.00352f
C4488 VDD.n2056 0 0.00147f
C4489 VDD.n2057 0 -0.0797f
C4490 VDD.n2058 0 0.00221f
C4491 VDD.n2059 0 0.00155f
C4492 VDD.n2060 0 0.00346f
C4493 VDD.n2061 0 0.00131f
C4494 VDD.n2062 0 1.19e-19
C4495 VDD.n2063 0 0.00101f
C4496 VDD.n2064 0 0.00104f
C4497 VDD.n2066 0 0.00485f
C4498 VDD.n2068 0 0.00393f
C4499 VDD.n2069 0 1.19e-19
C4500 VDD.n2070 0 0.00131f
C4501 VDD.n2071 0 1.79e-19
C4502 VDD.n2072 0 0.00178f
C4503 VDD.n2073 0 1.23e-19
C4504 VDD.n2074 0 0.00211f
C4505 VDD.n2075 0 0.00218f
C4506 VDD.n2076 0 0.00352f
C4507 VDD.n2077 0 0.00147f
C4508 VDD.n2078 0 0.00184f
C4509 VDD.n2079 0 0.00221f
C4510 VDD.n2080 0 0.00304f
C4511 VDD.n2081 0 0.0025f
C4512 VDD.n2082 0 0.00125f
C4513 VDD.n2083 0 0.0037f
C4514 VDD.n2084 0 0.0037f
C4515 VDD.n2085 0 0.00485f
C4516 VDD.n2087 0 0.00654f
C4517 VDD.n2088 0 0.0118f
C4518 VDD.n2089 0 0.0118f
C4519 VDD.n2090 0 0.00654f
C4520 VDD.n2091 0 0.00104f
C4521 VDD.n2092 0 0.00393f
C4522 VDD.n2093 0 1.19e-19
C4523 VDD.n2094 0 0.00131f
C4524 VDD.n2095 0 1.79e-19
C4525 VDD.n2096 0 0.00178f
C4526 VDD.n2097 0 1.23e-19
C4527 VDD.n2098 0 -0.0325f
C4528 VDD.n2099 0 0.00218f
C4529 VDD.n2100 0 0.0093f
C4530 VDD.n2101 0 0.00915f
C4531 VDD.n2102 0 0.00184f
C4532 VDD.n2103 0 0.00948f
C4533 VDD.n2104 0 0.00155f
C4534 VDD.n2105 0 0.00948f
C4535 VDD.n2106 0 0.00178f
C4536 VDD.n2107 0 0.00166f
C4537 VDD.n2108 0 0.00211f
C4538 VDD.n2109 0 -0.035f
C4539 VDD.n2110 0 -0.0709f
C4540 VDD.n2111 0 0.00301f
C4541 VDD.n2112 0 0.00184f
C4542 VDD.n2113 0 1.79e-19
C4543 VDD.n2114 0 0.00131f
C4544 VDD.n2115 0 1.19e-19
C4545 VDD.n2116 0 0.00393f
C4546 VDD.n2118 0 0.00485f
C4547 VDD.n2119 0 0.0037f
C4548 VDD.n2120 0 0.0037f
C4549 VDD.n2121 0 0.00125f
C4550 VDD.n2122 0 0.0025f
C4551 VDD.n2123 0 0.00304f
C4552 VDD.n2124 0 0.00155f
C4553 VDD.n2125 0 0.00221f
C4554 VDD.n2126 0 0.00178f
C4555 VDD.n2127 0 0.00166f
C4556 VDD.n2128 0 0.00211f
C4557 VDD.n2129 0 0.00218f
C4558 VDD.n2130 0 0.00345f
C4559 VDD.n2131 0 0.00352f
C4560 VDD.n2132 0 0.00301f
C4561 VDD.n2133 0 0.00184f
C4562 VDD.n2134 0 1.79e-19
C4563 VDD.n2135 0 0.00131f
C4564 VDD.n2136 0 1.19e-19
C4565 VDD.n2137 0 0.00393f
C4566 VDD.n2139 0 0.00485f
C4567 VDD.n2140 0 0.0037f
C4568 VDD.n2141 0 0.0037f
C4569 VDD.n2142 0 0.00125f
C4570 VDD.n2143 0 0.0025f
C4571 VDD.n2144 0 0.00304f
C4572 VDD.n2145 0 0.00221f
C4573 VDD.n2146 0 0.00155f
C4574 VDD.n2147 0 0.00125f
C4575 VDD.n2148 0 -0.0284f
C4576 VDD.n2149 0 1.23e-19
C4577 VDD.n2150 0 0.00184f
C4578 VDD.n2151 0 0.00301f
C4579 VDD.n2152 0 0.00352f
C4580 VDD.n2153 0 0.00345f
C4581 VDD.n2154 0 0.00211f
C4582 VDD.n2155 0 0.00166f
C4583 VDD.n2156 0 0.00178f
C4584 VDD.n2157 0 0.00221f
C4585 VDD.n2158 0 0.0025f
C4586 VDD.n2159 0 0.00304f
C4587 VDD.n2160 0 0.00131f
C4588 VDD.n2161 0 0.00101f
C4589 VDD.n2162 0 0.00131f
C4590 VDD.n2163 0 1.19e-19
C4591 VDD.n2164 0 0.00393f
C4592 VDD.n2165 0 0.00485f
C4593 VDD.n2167 0 0.00104f
C4594 VDD.n2168 0 0.00101f
C4595 VDD.n2169 0 1.19e-19
C4596 VDD.n2170 0 0.00131f
C4597 VDD.n2171 0 1.79e-19
C4598 VDD.n2172 0 0.00184f
C4599 VDD.n2173 0 0.00301f
C4600 VDD.n2174 0 -0.0709f
C4601 VDD.n2175 0 0.00345f
C4602 VDD.n2176 0 0.00211f
C4603 VDD.n2177 0 0.00166f
C4604 VDD.n2178 0 0.00178f
C4605 VDD.n2179 0 0.00221f
C4606 VDD.n2180 0 0.00304f
C4607 VDD.n2181 0 0.0025f
C4608 VDD.n2182 0 0.00125f
C4609 VDD.n2183 0 0.0037f
C4610 VDD.n2184 0 0.0037f
C4611 VDD.n2185 0 0.00485f
C4612 VDD.n2187 0 0.00104f
C4613 VDD.n2188 0 0.00393f
C4614 VDD.n2189 0 1.19e-19
C4615 VDD.n2190 0 0.00131f
C4616 VDD.n2191 0 1.79e-19
C4617 VDD.n2192 0 0.00184f
C4618 VDD.n2193 0 0.00301f
C4619 VDD.n2194 0 0.00352f
C4620 VDD.n2195 0 0.00345f
C4621 VDD.n2196 0 0.00211f
C4622 VDD.n2197 0 -0.0284f
C4623 VDD.n2198 0 -0.0798f
C4624 VDD.n2199 0 0.00221f
C4625 VDD.n2200 0 0.00304f
C4626 VDD.n2201 0 0.0025f
C4627 VDD.n2202 0 0.00125f
C4628 VDD.n2203 0 0.0037f
C4629 VDD.n2204 0 0.0037f
C4630 VDD.n2205 0 0.00485f
C4631 VDD.n2206 0 0.00104f
C4632 VDD.n2207 0 0.00883f
C4633 VDD.n2208 0 1.99e-19
C4634 VDD.n2209 0 0.00131f
C4635 VDD.n2210 0 1.79e-19
C4636 VDD.n2211 0 0.00184f
C4637 VDD.n2212 0 0.0108f
C4638 VDD.n2213 0 0.0125f
C4639 VDD.n2214 0 0.0124f
C4640 VDD.n2215 0 0.00218f
C4641 VDD.n2216 0 0.00211f
C4642 VDD.n2217 0 1.23e-19
C4643 VDD.n2218 0 0.00178f
C4644 VDD.n2219 0 1.79e-19
C4645 VDD.n2220 0 0.00131f
C4646 VDD.n2221 0 1.99e-19
C4647 VDD.n2222 0 0.00883f
C4648 VDD.n2223 0 0.00104f
C4649 VDD.n2224 0 0.00485f
C4650 VDD.n2227 0 0.00104f
C4651 VDD.n2228 0 0.00393f
C4652 VDD.n2229 0 1.19e-19
C4653 VDD.n2230 0 0.00101f
C4654 VDD.n2231 0 0.0037f
C4655 VDD.n2232 0 0.00125f
C4656 VDD.n2233 0 0.0025f
C4657 VDD.n2234 0 0.00304f
C4658 VDD.n2235 0 0.00221f
C4659 VDD.n2236 0 -0.0797f
C4660 VDD.n2237 0 0.00147f
C4661 VDD.n2238 0 0.00178f
C4662 VDD.n2239 0 0.00295f
C4663 VDD.n2240 0 0.00345f
C4664 VDD.n2241 0 0.00211f
C4665 VDD.n2242 0 -0.0735f
C4666 VDD.n2243 0 0.00178f
C4667 VDD.n2244 0 0.00295f
C4668 VDD.n2245 0 0.00147f
C4669 VDD.n2246 0 0.00352f
C4670 VDD.n2247 0 0.00218f
C4671 VDD.n2248 0 0.00166f
C4672 VDD.n2249 0 0.00125f
C4673 VDD.n2250 0 0.00155f
C4674 VDD.n2251 0 0.00346f
C4675 VDD.n2252 0 0.0025f
C4676 VDD.n2253 0 0.00304f
C4677 VDD.n2254 0 0.00131f
C4678 VDD.n2255 0 0.00101f
C4679 VDD.n2256 0 0.00101f
C4680 VDD.n2257 0 1.19e-19
C4681 VDD.n2258 0 0.00393f
C4682 VDD.n2260 0 0.00104f
C4683 VDD.n2262 0 0.00485f
C4684 VDD.n2263 0 0.0037f
C4685 VDD.n2264 0 0.0037f
C4686 VDD.n2265 0 0.00125f
C4687 VDD.n2266 0 0.00131f
C4688 VDD.n2267 0 0.00304f
C4689 VDD.n2268 0 0.0025f
C4690 VDD.n2269 0 0.00346f
C4691 VDD.n2270 0 0.00155f
C4692 VDD.n2271 0 0.00125f
C4693 VDD.n2272 0 0.00166f
C4694 VDD.n2273 0 0.00218f
C4695 VDD.n2274 0 0.00352f
C4696 VDD.n2275 0 0.00147f
C4697 VDD.n2276 0 0.00295f
C4698 VDD.n2277 0 0.00178f
C4699 VDD.n2278 0 1.23e-19
C4700 VDD.n2279 0 0.00211f
C4701 VDD.n2280 0 0.00218f
C4702 VDD.n2281 0 0.00352f
C4703 VDD.n2282 0 0.00147f
C4704 VDD.n2283 0 -0.0797f
C4705 VDD.n2284 0 0.00221f
C4706 VDD.n2285 0 0.00155f
C4707 VDD.n2286 0 0.00346f
C4708 VDD.n2287 0 0.00131f
C4709 VDD.n2288 0 1.19e-19
C4710 VDD.n2289 0 0.00101f
C4711 VDD.n2290 0 0.00104f
C4712 VDD.n2292 0 0.00485f
C4713 VDD.n2294 0 0.00393f
C4714 VDD.n2295 0 1.19e-19
C4715 VDD.n2296 0 0.00131f
C4716 VDD.n2297 0 1.79e-19
C4717 VDD.n2298 0 0.00178f
C4718 VDD.n2299 0 1.23e-19
C4719 VDD.n2300 0 0.00211f
C4720 VDD.n2301 0 0.00218f
C4721 VDD.n2302 0 0.00352f
C4722 VDD.n2303 0 0.00147f
C4723 VDD.n2304 0 0.00184f
C4724 VDD.n2305 0 0.00221f
C4725 VDD.n2306 0 0.00304f
C4726 VDD.n2307 0 0.0025f
C4727 VDD.n2308 0 0.00125f
C4728 VDD.n2309 0 0.0037f
C4729 VDD.n2310 0 0.0037f
C4730 VDD.n2311 0 0.00485f
C4731 VDD.n2313 0 0.00654f
C4732 VDD.n2314 0 0.0118f
C4733 VDD.n2315 0 0.0118f
C4734 VDD.n2316 0 0.00654f
C4735 VDD.n2317 0 0.00104f
C4736 VDD.n2318 0 0.00393f
C4737 VDD.n2319 0 1.19e-19
C4738 VDD.n2320 0 0.00131f
C4739 VDD.n2321 0 1.79e-19
C4740 VDD.n2322 0 0.00178f
C4741 VDD.n2323 0 1.23e-19
C4742 VDD.n2324 0 -0.0325f
C4743 VDD.n2325 0 0.00218f
C4744 VDD.n2326 0 0.0093f
C4745 VDD.n2327 0 0.00915f
C4746 VDD.n2328 0 0.00184f
C4747 VDD.n2329 0 0.00948f
C4748 VDD.n2330 0 0.00155f
C4749 VDD.n2331 0 0.00948f
C4750 VDD.n2332 0 0.00178f
C4751 VDD.n2333 0 0.00166f
C4752 VDD.n2334 0 0.00211f
C4753 VDD.n2335 0 -0.035f
C4754 VDD.n2336 0 -0.0709f
C4755 VDD.n2337 0 0.00301f
C4756 VDD.n2338 0 0.00184f
C4757 VDD.n2339 0 1.79e-19
C4758 VDD.n2340 0 0.00131f
C4759 VDD.n2341 0 1.19e-19
C4760 VDD.n2342 0 0.00393f
C4761 VDD.n2344 0 0.00485f
C4762 VDD.n2345 0 0.0037f
C4763 VDD.n2346 0 0.0037f
C4764 VDD.n2347 0 0.00125f
C4765 VDD.n2348 0 0.0025f
C4766 VDD.n2349 0 0.00304f
C4767 VDD.n2350 0 0.00155f
C4768 VDD.n2351 0 0.00221f
C4769 VDD.n2352 0 0.00178f
C4770 VDD.n2353 0 0.00166f
C4771 VDD.n2354 0 0.00211f
C4772 VDD.n2355 0 0.00218f
C4773 VDD.n2356 0 0.00345f
C4774 VDD.n2357 0 0.00352f
C4775 VDD.n2358 0 0.00301f
C4776 VDD.n2359 0 0.00184f
C4777 VDD.n2360 0 1.79e-19
C4778 VDD.n2361 0 0.00131f
C4779 VDD.n2362 0 1.19e-19
C4780 VDD.n2363 0 0.00393f
C4781 VDD.n2365 0 0.00485f
C4782 VDD.n2366 0 0.0037f
C4783 VDD.n2367 0 0.0037f
C4784 VDD.n2368 0 0.00125f
C4785 VDD.n2369 0 0.0025f
C4786 VDD.n2370 0 0.00304f
C4787 VDD.n2371 0 0.00221f
C4788 VDD.n2372 0 0.00155f
C4789 VDD.n2373 0 0.00125f
C4790 VDD.n2374 0 -0.0284f
C4791 VDD.n2375 0 1.23e-19
C4792 VDD.n2376 0 0.00184f
C4793 VDD.n2377 0 0.00301f
C4794 VDD.n2378 0 0.00352f
C4795 VDD.n2379 0 0.00345f
C4796 VDD.n2380 0 0.00211f
C4797 VDD.n2381 0 0.00166f
C4798 VDD.n2382 0 0.00178f
C4799 VDD.n2383 0 0.00221f
C4800 VDD.n2384 0 0.0025f
C4801 VDD.n2385 0 0.00304f
C4802 VDD.n2386 0 0.00131f
C4803 VDD.n2387 0 0.00101f
C4804 VDD.n2388 0 0.00131f
C4805 VDD.n2389 0 1.19e-19
C4806 VDD.n2390 0 0.00393f
C4807 VDD.n2391 0 0.00485f
C4808 VDD.n2393 0 0.00104f
C4809 VDD.n2394 0 0.00101f
C4810 VDD.n2395 0 1.19e-19
C4811 VDD.n2396 0 0.00131f
C4812 VDD.n2397 0 1.79e-19
C4813 VDD.n2398 0 0.00184f
C4814 VDD.n2399 0 0.00301f
C4815 VDD.n2400 0 -0.0709f
C4816 VDD.n2401 0 0.00345f
C4817 VDD.n2402 0 0.00211f
C4818 VDD.n2403 0 0.00166f
C4819 VDD.n2404 0 0.00178f
C4820 VDD.n2405 0 0.00221f
C4821 VDD.n2406 0 0.00304f
C4822 VDD.n2407 0 0.0025f
C4823 VDD.n2408 0 0.00125f
C4824 VDD.n2409 0 0.0037f
C4825 VDD.n2410 0 0.0037f
C4826 VDD.n2411 0 0.00485f
C4827 VDD.n2413 0 0.00104f
C4828 VDD.n2414 0 0.00393f
C4829 VDD.n2415 0 1.19e-19
C4830 VDD.n2416 0 0.00131f
C4831 VDD.n2417 0 1.79e-19
C4832 VDD.n2418 0 0.00184f
C4833 VDD.n2419 0 0.00301f
C4834 VDD.n2420 0 0.00352f
C4835 VDD.n2421 0 0.00345f
C4836 VDD.n2422 0 0.00211f
C4837 VDD.n2423 0 -0.0284f
C4838 VDD.n2424 0 -0.0798f
C4839 VDD.n2425 0 0.00221f
C4840 VDD.n2426 0 0.00304f
C4841 VDD.n2427 0 0.0025f
C4842 VDD.n2428 0 0.00125f
C4843 VDD.n2429 0 0.0037f
C4844 VDD.n2430 0 0.0037f
C4845 VDD.n2431 0 0.00485f
C4846 VDD.n2432 0 0.00104f
C4847 VDD.n2433 0 0.00883f
C4848 VDD.n2434 0 1.99e-19
C4849 VDD.n2435 0 0.00131f
C4850 VDD.n2436 0 1.79e-19
C4851 VDD.n2437 0 0.00184f
C4852 VDD.n2438 0 0.0108f
C4853 VDD.n2439 0 0.0125f
C4854 VDD.n2440 0 0.0124f
C4855 VDD.n2441 0 0.00218f
C4856 VDD.n2442 0 0.00211f
C4857 VDD.n2443 0 1.23e-19
C4858 VDD.n2444 0 0.00178f
C4859 VDD.n2445 0 1.79e-19
C4860 VDD.n2446 0 0.00131f
C4861 VDD.n2447 0 1.99e-19
C4862 VDD.n2448 0 0.00883f
C4863 VDD.n2449 0 0.00104f
C4864 VDD.n2450 0 0.00485f
C4865 VDD.n2453 0 0.00104f
C4866 VDD.n2454 0 0.00393f
C4867 VDD.n2455 0 1.19e-19
C4868 VDD.n2456 0 0.00101f
C4869 VDD.n2457 0 0.0037f
C4870 VDD.n2458 0 0.00125f
C4871 VDD.n2459 0 0.0025f
C4872 VDD.n2460 0 0.00304f
C4873 VDD.n2461 0 0.00221f
C4874 VDD.n2462 0 -0.0797f
C4875 VDD.n2463 0 0.00147f
C4876 VDD.n2464 0 0.00178f
C4877 VDD.n2465 0 0.00295f
C4878 VDD.n2466 0 0.00345f
C4879 VDD.n2467 0 0.00211f
C4880 VDD.n2468 0 -0.0735f
C4881 VDD.n2469 0 0.00178f
C4882 VDD.n2470 0 0.00295f
C4883 VDD.n2471 0 0.00147f
C4884 VDD.n2472 0 0.00352f
C4885 VDD.n2473 0 0.00218f
C4886 VDD.n2474 0 0.00166f
C4887 VDD.n2475 0 0.00125f
C4888 VDD.n2476 0 0.00155f
C4889 VDD.n2477 0 0.00346f
C4890 VDD.n2478 0 0.0025f
C4891 VDD.n2479 0 0.00304f
C4892 VDD.n2480 0 0.00131f
C4893 VDD.n2481 0 0.00101f
C4894 VDD.n2482 0 0.00101f
C4895 VDD.n2483 0 1.19e-19
C4896 VDD.n2484 0 0.00393f
C4897 VDD.n2486 0 0.00104f
C4898 VDD.n2488 0 0.00485f
C4899 VDD.n2489 0 0.0037f
C4900 VDD.n2490 0 0.0037f
C4901 VDD.n2491 0 0.00125f
C4902 VDD.n2492 0 0.00131f
C4903 VDD.n2493 0 0.00304f
C4904 VDD.n2494 0 0.0025f
C4905 VDD.n2495 0 0.00346f
C4906 VDD.n2496 0 0.00155f
C4907 VDD.n2497 0 0.00125f
C4908 VDD.n2498 0 0.00166f
C4909 VDD.n2499 0 0.00218f
C4910 VDD.n2500 0 0.00352f
C4911 VDD.n2501 0 0.00147f
C4912 VDD.n2502 0 0.00295f
C4913 VDD.n2503 0 0.00178f
C4914 VDD.n2504 0 1.23e-19
C4915 VDD.n2505 0 0.00211f
C4916 VDD.n2506 0 0.00218f
C4917 VDD.n2507 0 0.00352f
C4918 VDD.n2508 0 0.00147f
C4919 VDD.n2509 0 -0.0797f
C4920 VDD.n2510 0 0.00221f
C4921 VDD.n2511 0 0.00155f
C4922 VDD.n2512 0 0.00346f
C4923 VDD.n2513 0 0.00131f
C4924 VDD.n2514 0 1.19e-19
C4925 VDD.n2515 0 0.00101f
C4926 VDD.n2516 0 0.00104f
C4927 VDD.n2518 0 0.00485f
C4928 VDD.n2520 0 0.00393f
C4929 VDD.n2521 0 1.19e-19
C4930 VDD.n2522 0 0.00131f
C4931 VDD.n2523 0 1.79e-19
C4932 VDD.n2524 0 0.00178f
C4933 VDD.n2525 0 1.23e-19
C4934 VDD.n2526 0 0.00211f
C4935 VDD.n2527 0 0.00218f
C4936 VDD.n2528 0 0.00352f
C4937 VDD.n2529 0 0.00147f
C4938 VDD.n2530 0 0.00184f
C4939 VDD.n2531 0 0.00221f
C4940 VDD.n2532 0 0.00304f
C4941 VDD.n2533 0 0.0025f
C4942 VDD.n2534 0 0.00125f
C4943 VDD.n2535 0 0.0037f
C4944 VDD.n2536 0 0.0037f
C4945 VDD.n2537 0 0.00485f
C4946 VDD.n2539 0 0.00654f
C4947 VDD.n2540 0 0.0118f
C4948 VDD.n2541 0 0.0118f
C4949 VDD.n2542 0 0.00654f
C4950 VDD.n2543 0 0.00104f
C4951 VDD.n2544 0 0.00393f
C4952 VDD.n2545 0 1.19e-19
C4953 VDD.n2546 0 0.00131f
C4954 VDD.n2547 0 1.79e-19
C4955 VDD.n2548 0 0.00178f
C4956 VDD.n2549 0 1.23e-19
C4957 VDD.n2550 0 -0.0325f
C4958 VDD.n2551 0 0.00218f
C4959 VDD.n2552 0 0.0093f
C4960 VDD.n2553 0 0.00915f
C4961 VDD.n2554 0 0.00184f
C4962 VDD.n2555 0 0.00948f
C4963 VDD.n2556 0 0.00155f
C4964 VDD.n2557 0 0.00948f
C4965 VDD.n2558 0 0.00178f
C4966 VDD.n2559 0 0.00166f
C4967 VDD.n2560 0 0.00211f
C4968 VDD.n2561 0 -0.035f
C4969 VDD.n2562 0 -0.0709f
C4970 VDD.n2563 0 0.00301f
C4971 VDD.n2564 0 0.00184f
C4972 VDD.n2565 0 1.79e-19
C4973 VDD.n2566 0 0.00131f
C4974 VDD.n2567 0 1.19e-19
C4975 VDD.n2568 0 0.00393f
C4976 VDD.n2570 0 0.00485f
C4977 VDD.n2571 0 0.0037f
C4978 VDD.n2572 0 0.0037f
C4979 VDD.n2573 0 0.00125f
C4980 VDD.n2574 0 0.0025f
C4981 VDD.n2575 0 0.00304f
C4982 VDD.n2576 0 0.00155f
C4983 VDD.n2577 0 0.00221f
C4984 VDD.n2578 0 0.00178f
C4985 VDD.n2579 0 0.00166f
C4986 VDD.n2580 0 0.00211f
C4987 VDD.n2581 0 0.00218f
C4988 VDD.n2582 0 0.00345f
C4989 VDD.n2583 0 0.00352f
C4990 VDD.n2584 0 0.00301f
C4991 VDD.n2585 0 0.00184f
C4992 VDD.n2586 0 1.79e-19
C4993 VDD.n2587 0 0.00131f
C4994 VDD.n2588 0 1.19e-19
C4995 VDD.n2589 0 0.00393f
C4996 VDD.n2591 0 0.00485f
C4997 VDD.n2592 0 0.0037f
C4998 VDD.n2593 0 0.0037f
C4999 VDD.n2594 0 0.00125f
C5000 VDD.n2595 0 0.0025f
C5001 VDD.n2596 0 0.00304f
C5002 VDD.n2597 0 0.00221f
C5003 VDD.n2598 0 0.00155f
C5004 VDD.n2599 0 0.00125f
C5005 VDD.n2600 0 -0.0284f
C5006 VDD.n2601 0 1.23e-19
C5007 VDD.n2602 0 0.00184f
C5008 VDD.n2603 0 0.00301f
C5009 VDD.n2604 0 0.00352f
C5010 VDD.n2605 0 0.00345f
C5011 VDD.n2606 0 0.00211f
C5012 VDD.n2607 0 0.00166f
C5013 VDD.n2608 0 0.00178f
C5014 VDD.n2609 0 0.00221f
C5015 VDD.n2610 0 0.0025f
C5016 VDD.n2611 0 0.00304f
C5017 VDD.n2612 0 0.00131f
C5018 VDD.n2613 0 0.00101f
C5019 VDD.n2614 0 0.00131f
C5020 VDD.n2615 0 1.19e-19
C5021 VDD.n2616 0 0.00393f
C5022 VDD.n2617 0 0.00485f
C5023 VDD.n2619 0 0.00104f
C5024 VDD.n2620 0 0.00101f
C5025 VDD.n2621 0 1.19e-19
C5026 VDD.n2622 0 0.00131f
C5027 VDD.n2623 0 1.79e-19
C5028 VDD.n2624 0 0.00184f
C5029 VDD.n2625 0 0.00301f
C5030 VDD.n2626 0 -0.0709f
C5031 VDD.n2627 0 0.00345f
C5032 VDD.n2628 0 0.00211f
C5033 VDD.n2629 0 0.00166f
C5034 VDD.n2630 0 0.00178f
C5035 VDD.n2631 0 0.00221f
C5036 VDD.n2632 0 0.00304f
C5037 VDD.n2633 0 0.0025f
C5038 VDD.n2634 0 0.00125f
C5039 VDD.n2635 0 0.0037f
C5040 VDD.n2636 0 0.0037f
C5041 VDD.n2637 0 0.00485f
C5042 VDD.n2639 0 0.00104f
C5043 VDD.n2640 0 0.00393f
C5044 VDD.n2641 0 1.19e-19
C5045 VDD.n2642 0 0.00131f
C5046 VDD.n2643 0 1.79e-19
C5047 VDD.n2644 0 0.00184f
C5048 VDD.n2645 0 0.00301f
C5049 VDD.n2646 0 0.00352f
C5050 VDD.n2647 0 0.00345f
C5051 VDD.n2648 0 0.00211f
C5052 VDD.n2649 0 -0.0284f
C5053 VDD.n2650 0 -0.0798f
C5054 VDD.n2651 0 0.00221f
C5055 VDD.n2652 0 0.00304f
C5056 VDD.n2653 0 0.0025f
C5057 VDD.n2654 0 0.00125f
C5058 VDD.n2655 0 0.0037f
C5059 VDD.n2656 0 0.0037f
C5060 VDD.n2657 0 0.00485f
C5061 VDD.n2658 0 0.00104f
C5062 VDD.n2659 0 0.00883f
C5063 VDD.n2660 0 1.99e-19
C5064 VDD.n2661 0 0.00131f
C5065 VDD.n2662 0 1.79e-19
C5066 VDD.n2663 0 0.00184f
C5067 VDD.n2664 0 0.0108f
C5068 VDD.n2665 0 0.0125f
C5069 VDD.n2666 0 0.0124f
C5070 VDD.n2667 0 0.00218f
C5071 VDD.n2668 0 0.00211f
C5072 VDD.n2669 0 1.23e-19
C5073 VDD.n2670 0 0.00178f
C5074 VDD.n2671 0 1.79e-19
C5075 VDD.n2672 0 0.00131f
C5076 VDD.n2673 0 1.99e-19
C5077 VDD.n2674 0 0.00883f
C5078 VDD.n2675 0 0.00104f
C5079 VDD.n2676 0 0.00485f
C5080 VDD.n2679 0 0.00104f
C5081 VDD.n2680 0 0.00393f
C5082 VDD.n2681 0 1.19e-19
C5083 VDD.n2682 0 0.00101f
C5084 VDD.n2683 0 0.0037f
C5085 VDD.n2684 0 0.00125f
C5086 VDD.n2685 0 0.0025f
C5087 VDD.n2686 0 0.00304f
C5088 VDD.n2687 0 0.00221f
C5089 VDD.n2688 0 -0.0797f
C5090 VDD.n2689 0 0.00147f
C5091 VDD.n2690 0 0.00178f
C5092 VDD.n2691 0 0.00295f
C5093 VDD.n2692 0 0.00345f
C5094 VDD.n2693 0 0.00211f
C5095 VDD.n2694 0 -0.0735f
C5096 VDD.n2695 0 0.00178f
C5097 VDD.n2696 0 0.00295f
C5098 VDD.n2697 0 0.00147f
C5099 VDD.n2698 0 0.00352f
C5100 VDD.n2699 0 0.00218f
C5101 VDD.n2700 0 0.00166f
C5102 VDD.n2701 0 0.00125f
C5103 VDD.n2702 0 0.00155f
C5104 VDD.n2703 0 0.00346f
C5105 VDD.n2704 0 0.0025f
C5106 VDD.n2705 0 0.00304f
C5107 VDD.n2706 0 0.00131f
C5108 VDD.n2707 0 0.00101f
C5109 VDD.n2708 0 0.00101f
C5110 VDD.n2709 0 1.19e-19
C5111 VDD.n2710 0 0.00393f
C5112 VDD.n2712 0 0.00104f
C5113 VDD.n2714 0 0.00485f
C5114 VDD.n2715 0 0.0037f
C5115 VDD.n2716 0 0.0037f
C5116 VDD.n2717 0 0.00125f
C5117 VDD.n2718 0 0.00131f
C5118 VDD.n2719 0 0.00304f
C5119 VDD.n2720 0 0.0025f
C5120 VDD.n2721 0 0.00346f
C5121 VDD.n2722 0 0.00155f
C5122 VDD.n2723 0 0.00125f
C5123 VDD.n2724 0 0.00166f
C5124 VDD.n2725 0 0.00218f
C5125 VDD.n2726 0 0.00352f
C5126 VDD.n2727 0 0.00147f
C5127 VDD.n2728 0 0.00295f
C5128 VDD.n2729 0 0.00178f
C5129 VDD.n2730 0 1.23e-19
C5130 VDD.n2731 0 0.00211f
C5131 VDD.n2732 0 0.00218f
C5132 VDD.n2733 0 0.00352f
C5133 VDD.n2734 0 0.00147f
C5134 VDD.n2735 0 -0.0797f
C5135 VDD.n2736 0 0.00221f
C5136 VDD.n2737 0 0.00155f
C5137 VDD.n2738 0 0.00346f
C5138 VDD.n2739 0 0.00131f
C5139 VDD.n2740 0 1.19e-19
C5140 VDD.n2741 0 0.00101f
C5141 VDD.n2742 0 0.00104f
C5142 VDD.n2744 0 0.00485f
C5143 VDD.n2746 0 0.00393f
C5144 VDD.n2747 0 1.19e-19
C5145 VDD.n2748 0 0.00131f
C5146 VDD.n2749 0 1.79e-19
C5147 VDD.n2750 0 0.00178f
C5148 VDD.n2751 0 1.23e-19
C5149 VDD.n2752 0 0.00211f
C5150 VDD.n2753 0 0.00218f
C5151 VDD.n2754 0 0.00178f
C5152 VDD.n2755 0 1.23e-19
C5153 VDD.n2756 0 -0.0325f
C5154 VDD.n2757 0 -0.0735f
C5155 VDD.n2758 0 0.00352f
C5156 VDD.n2759 0 0.00147f
C5157 VDD.n2760 0 0.00184f
C5158 VDD.n2761 0 0.00221f
C5159 VDD.n2762 0 0.00131f
C5160 VDD.n2763 0 0.00304f
C5161 VDD.n2764 0 0.0025f
C5162 VDD.n2765 0 0.00125f
C5163 VDD.n2766 0 0.0037f
C5164 VDD.n2767 0 0.0037f
C5165 VDD.n2768 0 0.00485f
C5166 VDD.n2769 0 0.00764f
C5167 VDD.n2770 0 0.0195f
C5168 VDD.n2771 0 0.0159f
C5169 VDD.n2772 0 0.0147f
C5170 VDD.n2773 0 0.015f
C5171 VDD.n2774 0 0.00931f
C5172 VDD.n2775 0 0.0147f
C5173 VDD.n2776 0 0.00104f
C5174 VDD.n2777 0 0.00891f
C5175 VDD.n2778 0 0.0118f
C5176 VDD.n2779 0 0.0218f
C5177 VDD.n2780 0 0.00125f
C5178 VDD.n2781 0 0.0163f
C5179 VDD.n2782 0 0.0166f
C5180 VDD.n2783 0 1.23e-19
C5181 VDD.n2784 0 0.00219f
C5182 VDD.n2785 0 0.00227f
C5183 VDD.n2786 0 0.00366f
C5184 VDD.n2787 0 0.00147f
C5185 VDD.n2788 0 -0.0797f
C5186 VDD.n2789 0 0.00221f
C5187 VDD.n2790 0 0.00304f
C5188 VDD.n2791 0 0.0025f
C5189 VDD.n2792 0 0.00125f
C5190 VDD.n2793 0 0.0037f
C5191 VDD.n2794 0 0.0037f
C5192 VDD.n2795 0 0.00485f
C5193 VDD.n2797 0 0.00393f
C5194 VDD.n2798 0 1.19e-19
C5195 VDD.n2799 0 0.00131f
C5196 VDD.n2800 0 1.79e-19
C5197 VDD.n2801 0 0.00178f
C5198 VDD.n2802 0 1.23e-19
C5199 VDD.n2803 0 0.00219f
C5200 VDD.n2804 0 0.00227f
C5201 VDD.n2805 0 0.00366f
C5202 VDD.n2806 0 0.00147f
C5203 VDD.n2807 0 0.00184f
C5204 VDD.n2808 0 0.00221f
C5205 VDD.n2809 0 0.00304f
C5206 VDD.n2810 0 0.0025f
C5207 VDD.n2811 0 0.00125f
C5208 VDD.n2812 0 0.0037f
C5209 VDD.n2813 0 0.0037f
C5210 VDD.n2814 0 0.00485f
C5211 VDD.n2816 0 0.00393f
C5212 VDD.n2817 0 1.19e-19
C5213 VDD.n2818 0 0.00131f
C5214 VDD.n2819 0 1.79e-19
C5215 VDD.n2820 0 0.00178f
C5216 VDD.n2821 0 1.23e-19
C5217 VDD.n2822 0 -0.0325f
C5218 VDD.n2823 0 0.00227f
C5219 VDD.n2824 0 0.00366f
C5220 VDD.n2825 0 0.00147f
C5221 VDD.n2826 0 0.00184f
C5222 VDD.n2827 0 0.00221f
C5223 VDD.n2828 0 0.00304f
C5224 VDD.n2829 0 0.0025f
C5225 VDD.n2830 0 0.00125f
C5226 VDD.n2831 0 0.0037f
C5227 VDD.n2832 0 0.0037f
C5228 VDD.n2833 0 0.00485f
C5229 VDD.n2835 0 0.00393f
C5230 VDD.n2836 0 1.19e-19
C5231 VDD.n2837 0 0.00131f
C5232 VDD.n2838 0 1.79e-19
C5233 VDD.n2839 0 0.00178f
C5234 VDD.n2840 0 1.23e-19
C5235 VDD.n2841 0 0.00219f
C5236 VDD.n2842 0 0.00227f
C5237 VDD.n2843 0 0.00366f
C5238 VDD.n2844 0 0.00147f
C5239 VDD.n2845 0 -0.0797f
C5240 VDD.n2846 0 0.00221f
C5241 VDD.n2847 0 0.00304f
C5242 VDD.n2848 0 0.0025f
C5243 VDD.n2849 0 0.00125f
C5244 VDD.n2850 0 0.0037f
C5245 VDD.n2851 0 0.0037f
C5246 VDD.n2852 0 0.00485f
C5247 VDD.n2854 0 0.00393f
C5248 VDD.n2855 0 1.19e-19
C5249 VDD.n2856 0 0.00131f
C5250 VDD.n2857 0 1.79e-19
C5251 VDD.n2858 0 0.00178f
C5252 VDD.n2859 0 1.23e-19
C5253 VDD.n2860 0 0.00219f
C5254 VDD.n2861 0 0.00227f
C5255 VDD.n2862 0 -0.0734f
C5256 VDD.n2863 0 0.00366f
C5257 VDD.n2864 0 0.00147f
C5258 VDD.n2865 0 0.00184f
C5259 VDD.n2866 0 0.00221f
C5260 VDD.n2867 0 0.00304f
C5261 VDD.n2868 0 0.0025f
C5262 VDD.n2869 0 0.00125f
C5263 VDD.n2870 0 0.0037f
C5264 VDD.n2871 0 0.0037f
C5265 VDD.n2872 0 0.00485f
C5266 VDD.n2874 0 0.00393f
C5267 VDD.n2875 0 1.19e-19
C5268 VDD.n2876 0 0.00131f
C5269 VDD.n2877 0 1.79e-19
C5270 VDD.n2878 0 0.00294f
C5271 VDD.n2879 0 0.00155f
C5272 VDD.n2880 0 0.00125f
C5273 VDD.n2881 0 0.00166f
C5274 VDD.n2882 0 0.00227f
C5275 VDD.n2883 0 0.00241f
C5276 VDD.n2884 0 0.00289f
C5277 VDD.n2885 0 0.00308f
C5278 VDD.n2886 0 0.00489f
C5279 VDD.n2887 0 0.00466f
C5280 VDD.n2888 0 0.00419f
C5281 VDD.n2889 0 4.01e-19
C5282 VDD.n2890 0 0.00655f
C5283 VDD.n2891 0 0.0136f
C5284 VDD.n2892 0 0.0219f
C5285 VDD.n2893 0 0.0239f
C5286 VDD.n2894 0 0.0307f
C5287 VDD.n2895 0 0.0307f
C5288 VDD.n2896 0 0.00311f
C5289 VDD.n2897 0 0.00754f
C5290 VDD.n2898 0 0.00753f
C5291 VDD.n2899 0 0.00727f
C5292 VDD.n2900 0 0.00647f
C5293 VDD.n2901 0 0.00296f
C5294 VDD.n2902 0 0.00635f
C5295 VDD.n2903 0 0.0025f
C5296 VDD.t237 0 0.0025f
C5297 VDD.t234 0 0.0025f
C5298 VDD.n2904 0 0.00614f
C5299 VDD.n2905 0 0.0182f
C5300 VDD.n2906 0 0.00304f
C5301 VDD.n2907 0 0.00621f
C5302 VDD.n2908 0 0.051f
C5303 VDD.n2909 0 0.0324f
C5304 VDD.n2910 0 0.0157f
C5305 VDD.n2911 0 0.00753f
C5306 VDD.n2912 0 0.0177f
C5307 VDD.n2913 0 0.00751f
C5308 VDD.n2914 0 0.00314f
C5309 VDD.n2915 0 0.00239f
C5310 VDD.n2916 0 0.00309f
C5311 VDD.n2917 0 0.00754f
C5312 VDD.n2918 0 0.0336f
C5313 VDD.n2919 0 0.0041f
C5314 VDD.n2920 0 0.0432f
C5315 VDD.n2921 0 0.0286f
C5316 VDD.n2922 0 0.123f
C5317 VDD.n2923 0 0.0041f
C5318 VDD.n2924 0 0.0307f
C5319 VDD.n2925 0 0.0157f
C5320 VDD.n2926 0 0.0078f
C5321 VDD.t174 0 0.00356f
C5322 VDD.n2927 0 0.0515f
C5323 VDD.n2928 0 0.00434f
C5324 VDD.n2929 0 0.00752f
C5325 VDD.n2930 0 0.111f
C5326 VDD.n2931 0 0.0121f
C5327 VDD.n2932 0 0.00754f
C5328 VDD.n2933 0 0.00309f
C5329 VDD.n2934 0 0.00239f
C5330 VDD.n2935 0 0.00311f
C5331 VDD.n2936 0 0.00753f
C5332 VDD.n2937 0 0.00787f
C5333 VDD.n2938 0 0.0127f
C5334 VDD.n2939 0 0.0121f
C5335 VDD.n2940 0 0.00754f
C5336 VDD.n2941 0 0.00311f
C5337 VDD.n2942 0 0.00309f
C5338 VDD.n2943 0 0.00239f
C5339 VDD.n2944 0 0.0041f
C5340 VDD.n2945 0 0.0063f
C5341 VDD.n2946 0 0.0041f
C5342 VDD.n2947 0 0.00239f
C5343 VDD.n2948 0 0.00309f
C5344 VDD.n2949 0 0.0307f
C5345 VDD.t42 0 0.935f
C5346 VDD.n2950 0 0.832f
C5347 VDD.t121 0 1.01f
C5348 VDD.n2951 0 0.831f
C5349 VDD.t126 0 0.905f
C5350 VDD.n2952 0 0.808f
C5351 VDD.n2953 0 0.122f
C5352 VDD.t215 0 0.667f
C5353 VDD.n2954 0 0.188f
C5354 VDD.n2955 0 0.00314f
C5355 VDD.n2956 0 0.0307f
C5356 VDD.n2957 0 0.00309f
C5357 VDD.n2958 0 0.00754f
C5358 VDD.n2959 0 0.0041f
C5359 VDD.n2960 0 0.00972f
C5360 VDD.n2961 0 0.164f
C5361 VDD.n2962 0 0.0115f
C5362 VDD.n2963 0 0.48f
C5363 VDD.n2964 0 0.00765f
C5364 VDD.t188 0 0.0197f
C5365 VDD.n2965 0 0.0315f
C5366 VDD.n2966 0 0.00147f
C5367 VDD.t189 0 -6.65e-20
C5368 VDD.t236 0 0.00416f
C5369 VDD.n2967 0 0.0188f
C5370 VDD.n2968 0 0.0214f
C5371 VDD.n2969 0 0.00523f
C5372 VDD.n2970 0 0.0249f
C5373 VDD.n2971 0 0.00416f
C5374 VDD.n2972 0 0.00112f
C5375 VDD.n2973 0 0.00106f
C5376 VDD.n2974 0 0.00573f
C5377 VDD.n2975 0 0.00373f
C5378 VDD.n2976 0 0.0396f
C5379 VDD.n2977 0 0.0221f
C5380 VDD.n2978 0 0.00857f
C5381 VDD.n2979 0 0.00755f
C5382 VDD.n2980 0 0.0808f
C5383 VDD.n2981 0 0.0892f
C5384 VDD.n2982 0 0.0315f
C5385 VDD.n2983 0 0.0041f
C5386 VDD.n2984 0 0.00752f
C5387 VDD.n2985 0 0.00847f
C5388 VDD.n2986 0 0.00313f
C5389 VDD.n2987 0 0.0182f
C5390 VDD.n2988 0 0.00633f
C5391 VDD.n2989 0 0.00679f
C5392 VDD.n2990 0 0.00839f
C5393 VDD.n2992 0 1.36f
C5394 VDD.t37 0 1.46f
C5395 VDD.n2993 0 0.365f
C5396 VDD.t232 0 0.0471f
C5397 VDD.n2994 0 0.0239f
C5398 VDD.n2995 0 0.0119f
C5399 VDD.n2996 0 0.00301f
C5400 VDD.n2997 0 0.00147f
C5401 VDD.n2998 0 0.00413f
C5402 VDD.n2999 0 0.00402f
C5403 VDD.n3000 0 0.0103f
C5404 VDD.n3001 0 0.0065f
C5405 VDD.n3002 0 0.00747f
C5406 VDD.n3003 0 3.08e-19
C5407 VDD.n3004 0 0.00986f
C5408 VDD.n3005 0 0.00754f
C5409 VDD.n3006 0 0.00906f
C5410 VDD.n3007 0 0.00151f
C5411 VDD.n3008 0 0.00468f
C5412 VDD.n3009 0 0.00174f
C5413 VDD.n3010 0 0.00182f
C5414 VDD.n3011 0 6.94e-19
C5415 VDD.n3012 0 5.11e-19
C5416 VDD.n3013 0 0.00408f
C5417 VDD.n3014 0 9.66e-19
C5418 VDD.n3015 0 6.14e-19
C5419 VDD.n3016 0 0.00563f
C5420 VDD.n3017 0 0.0285f
C5421 VDD.t230 0 0.0388f
C5422 VDD.n3018 0 0.0351f
C5423 VDD.n3019 0 0.00762f
C5424 VDD.n3020 0 0.00301f
C5425 VDD.n3021 0 0.021f
C5426 VDD.n3022 0 0.00848f
.ends

