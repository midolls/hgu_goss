* NGSPICE file created from hgu_cdac_cap_4.ext - technology: sky130A


* Top level circuit hgu_cdac_cap_4

C0 hgu_cdac_unit_3.CTOP hgu_cdac_unit_3.SUB 4.58f $ **FLOATING
.end

