magic
tech sky130A
magscale 1 2
timestamp 1698575955
<< pwell >>
rect 484 1736 906 2240
rect 689 963 715 995
<< nmos >>
rect 680 1946 710 2030
<< ndiff >>
rect 622 2018 680 2030
rect 622 1958 634 2018
rect 668 1958 680 2018
rect 622 1946 680 1958
rect 710 2018 768 2030
rect 710 1958 722 2018
rect 756 1958 768 2018
rect 710 1946 768 1958
<< ndiffc >>
rect 634 1958 668 2018
rect 722 1958 756 2018
<< psubdiff >>
rect 520 2170 616 2204
rect 774 2170 870 2204
rect 520 2108 554 2170
rect 836 2108 870 2170
rect 520 1806 554 1868
rect 836 1806 870 1868
rect 520 1772 616 1806
rect 774 1772 870 1806
<< psubdiffcont >>
rect 616 2170 774 2204
rect 520 1868 554 2108
rect 836 1868 870 2108
rect 616 1772 774 1806
<< poly >>
rect 662 2102 728 2118
rect 662 2068 678 2102
rect 712 2068 728 2102
rect 662 2052 728 2068
rect 680 2030 710 2052
rect 680 1924 710 1946
rect 662 1908 728 1924
rect 662 1874 678 1908
rect 712 1874 728 1908
rect 662 1858 728 1874
<< polycont >>
rect 678 2068 712 2102
rect 678 1874 712 1908
<< locali >>
rect 520 2170 616 2204
rect 774 2170 870 2204
rect 520 2108 554 2170
rect 836 2108 870 2170
rect 662 2068 678 2102
rect 712 2068 728 2102
rect 634 2018 668 2034
rect 634 1942 668 1958
rect 722 2018 756 2034
rect 722 1942 756 1958
rect 662 1874 678 1908
rect 712 1874 728 1908
rect 520 1806 554 1868
rect 836 1806 870 1868
rect 520 1772 616 1806
rect 774 1772 870 1806
<< viali >>
rect 678 2068 712 2102
rect 634 1958 668 2018
rect 722 1958 756 2018
rect 678 1874 712 1908
<< metal1 >>
rect 666 2102 724 2108
rect 666 2068 678 2102
rect 712 2068 724 2102
rect 666 2062 724 2068
rect 628 2018 674 2030
rect 628 1958 634 2018
rect 668 1958 674 2018
rect 628 1946 674 1958
rect 716 2018 762 2030
rect 716 1958 722 2018
rect 756 1958 762 2018
rect 716 1946 762 1958
rect 666 1908 724 1914
rect 666 1874 678 1908
rect 712 1874 724 1908
rect 666 1868 724 1874
<< metal3 >>
rect 369 1773 1041 1775
rect 369 1709 473 1773
rect 537 1709 553 1773
rect 617 1709 633 1773
rect 697 1709 713 1773
rect 777 1709 793 1773
rect 857 1709 873 1773
rect 937 1709 1041 1773
rect 369 1707 1041 1709
rect 369 1553 435 1707
rect 369 1489 370 1553
rect 434 1489 435 1553
rect 369 1473 435 1489
rect 369 1409 370 1473
rect 434 1409 435 1473
rect 369 1393 435 1409
rect 369 1329 370 1393
rect 434 1329 435 1393
rect 369 1313 435 1329
rect 369 1249 370 1313
rect 434 1249 435 1313
rect 369 1233 435 1249
rect 369 1169 370 1233
rect 434 1169 435 1233
rect 369 1153 435 1169
rect 369 1089 370 1153
rect 434 1089 435 1153
rect 369 1073 435 1089
rect 369 1009 370 1073
rect 434 1009 435 1073
rect 369 993 435 1009
rect 369 929 370 993
rect 434 929 435 993
rect 369 913 435 929
rect 369 849 370 913
rect 434 849 435 913
rect 369 833 435 849
rect 369 769 370 833
rect 434 769 435 833
rect 369 679 435 769
rect 495 675 555 1707
rect 615 615 675 1645
rect 735 675 795 1707
rect 855 615 915 1645
rect 975 1553 1041 1707
rect 975 1489 976 1553
rect 1040 1489 1041 1553
rect 975 1473 1041 1489
rect 975 1409 976 1473
rect 1040 1409 1041 1473
rect 975 1393 1041 1409
rect 975 1329 976 1393
rect 1040 1329 1041 1393
rect 975 1313 1041 1329
rect 975 1249 976 1313
rect 1040 1249 1041 1313
rect 975 1233 1041 1249
rect 975 1169 976 1233
rect 1040 1169 1041 1233
rect 975 1153 1041 1169
rect 975 1089 976 1153
rect 1040 1089 1041 1153
rect 975 1073 1041 1089
rect 975 1009 976 1073
rect 1040 1009 1041 1073
rect 975 993 1041 1009
rect 975 929 976 993
rect 1040 929 1041 993
rect 975 913 1041 929
rect 975 849 976 913
rect 1040 849 1041 913
rect 975 833 1041 849
rect 975 769 976 833
rect 1040 769 1041 833
rect 975 679 1041 769
rect 369 613 1041 615
rect 369 549 473 613
rect 537 549 553 613
rect 617 549 633 613
rect 697 549 713 613
rect 777 549 793 613
rect 857 549 873 613
rect 937 549 1041 613
rect 369 547 1041 549
<< via3 >>
rect 473 1709 537 1773
rect 553 1709 617 1773
rect 633 1709 697 1773
rect 713 1709 777 1773
rect 793 1709 857 1773
rect 873 1709 937 1773
rect 370 1489 434 1553
rect 370 1409 434 1473
rect 370 1329 434 1393
rect 370 1249 434 1313
rect 370 1169 434 1233
rect 370 1089 434 1153
rect 370 1009 434 1073
rect 370 929 434 993
rect 370 849 434 913
rect 370 769 434 833
rect 976 1489 1040 1553
rect 976 1409 1040 1473
rect 976 1329 1040 1393
rect 976 1249 1040 1313
rect 976 1169 1040 1233
rect 976 1089 1040 1153
rect 976 1009 1040 1073
rect 976 929 1040 993
rect 976 849 1040 913
rect 976 769 1040 833
rect 473 549 537 613
rect 553 549 617 613
rect 633 549 697 613
rect 713 549 777 613
rect 793 549 857 613
rect 873 549 937 613
<< metal4 >>
rect 369 1773 1041 1775
rect 369 1709 473 1773
rect 537 1709 553 1773
rect 617 1709 633 1773
rect 697 1709 713 1773
rect 777 1709 793 1773
rect 857 1709 873 1773
rect 937 1709 1041 1773
rect 369 1707 1041 1709
rect 369 1553 435 1707
rect 369 1489 370 1553
rect 434 1489 435 1553
rect 369 1473 435 1489
rect 369 1409 370 1473
rect 434 1409 435 1473
rect 369 1393 435 1409
rect 369 1329 370 1393
rect 434 1329 435 1393
rect 369 1313 435 1329
rect 369 1249 370 1313
rect 434 1249 435 1313
rect 369 1233 435 1249
rect 369 1169 370 1233
rect 434 1169 435 1233
rect 369 1153 435 1169
rect 369 1089 370 1153
rect 434 1089 435 1153
rect 369 1073 435 1089
rect 369 1009 370 1073
rect 434 1009 435 1073
rect 369 993 435 1009
rect 369 929 370 993
rect 434 929 435 993
rect 369 913 435 929
rect 369 849 370 913
rect 434 849 435 913
rect 369 833 435 849
rect 369 769 370 833
rect 434 769 435 833
rect 369 679 435 769
rect 495 615 555 1645
rect 615 675 675 1707
rect 735 615 795 1645
rect 855 675 915 1707
rect 975 1553 1041 1707
rect 975 1489 976 1553
rect 1040 1489 1041 1553
rect 975 1473 1041 1489
rect 975 1409 976 1473
rect 1040 1409 1041 1473
rect 975 1393 1041 1409
rect 975 1329 976 1393
rect 1040 1329 1041 1393
rect 975 1313 1041 1329
rect 975 1249 976 1313
rect 1040 1249 1041 1313
rect 975 1233 1041 1249
rect 975 1169 976 1233
rect 1040 1169 1041 1233
rect 975 1153 1041 1169
rect 975 1089 976 1153
rect 1040 1089 1041 1153
rect 975 1073 1041 1089
rect 975 1009 976 1073
rect 1040 1009 1041 1073
rect 975 993 1041 1009
rect 975 929 976 993
rect 1040 929 1041 993
rect 975 913 1041 929
rect 975 849 976 913
rect 1040 849 1041 913
rect 975 833 1041 849
rect 975 769 976 833
rect 1040 769 1041 833
rect 975 679 1041 769
rect 369 613 1041 615
rect 369 549 473 613
rect 537 549 553 613
rect 617 549 633 613
rect 697 549 713 613
rect 777 549 793 613
rect 857 549 873 613
rect 937 549 1041 613
rect 369 547 1041 549
<< labels >>
flabel pwell 689 963 715 995 0 FreeSans 160 0 0 0 x2.SUB
flabel metal4 631 1297 657 1329 0 FreeSans 320 0 0 0 x2.CBOT
flabel metal4 749 707 775 739 0 FreeSans 320 0 0 0 x2.CTOP
<< end >>
