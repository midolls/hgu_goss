magic
tech sky130A
magscale 1 2
timestamp 1699484509
<< error_p >>
rect -41 855 324 905
rect -127 769 324 855
rect 41 754 156 769
rect 41 737 190 754
rect 41 733 359 737
rect 41 723 127 733
rect 5 720 127 723
rect 156 720 359 733
rect 5 699 359 720
rect 41 687 359 699
rect 41 674 295 687
rect 79 -521 113 -351
rect 43 -550 149 -521
rect 195 -548 359 -452
rect 79 -557 113 -550
rect 195 -557 551 -548
rect 79 -605 551 -557
rect -323 -705 157 -680
rect 195 -706 551 -605
rect -359 -741 193 -716
<< nwell >>
rect -359 737 359 769
rect -359 687 127 737
rect -359 674 41 687
rect 156 674 359 737
rect -359 -557 359 674
rect -359 -605 79 -557
rect 113 -605 359 -557
rect -359 -694 359 -605
rect -359 -706 195 -694
rect -359 -716 551 -706
<< pmos >>
rect -159 -550 -129 550
rect -63 -550 -33 550
rect 33 -550 63 550
rect 129 -550 159 550
<< pdiff >>
rect -221 538 -159 550
rect -221 -538 -209 538
rect -175 -538 -159 538
rect -221 -550 -159 -538
rect -129 538 -63 550
rect -129 -538 -113 538
rect -79 -538 -63 538
rect -129 -550 -63 -538
rect -33 538 33 550
rect -33 -538 -17 538
rect 17 -538 33 538
rect -33 -550 33 -538
rect 63 538 129 550
rect 63 -538 79 538
rect 113 -538 129 538
rect 63 -550 129 -538
rect 159 538 221 550
rect 159 -538 175 538
rect 209 -538 221 538
rect 159 -550 221 -538
<< pdiffc >>
rect -209 -538 -175 538
rect -113 -538 -79 538
rect -17 -538 17 538
rect 79 -538 113 538
rect 175 -538 209 538
<< nsubdiff >>
rect -323 699 -217 733
rect -167 699 -121 733
rect -71 699 -25 733
rect 25 699 71 733
rect 121 720 166 733
rect 121 699 127 720
rect 156 699 166 720
rect -323 637 -289 699
rect -323 -671 -289 -594
rect -323 -705 -217 -671
rect -167 -705 -121 -671
rect -71 -705 -25 -671
rect 25 -705 71 -671
rect 121 -705 157 -671
<< nsubdiffcont >>
rect -217 699 -167 733
rect -121 699 -71 733
rect -25 699 25 733
rect 71 699 121 733
rect -323 -594 -289 637
rect -217 -705 -167 -671
rect -121 -705 -71 -671
rect -25 -705 25 -671
rect 71 -705 121 -671
<< poly >>
rect -159 550 -129 576
rect -63 550 -33 576
rect 33 550 63 576
rect 129 550 159 576
rect -159 -576 -129 -550
rect -63 -576 -33 -550
rect 33 -576 63 -550
rect 129 -576 159 -550
<< locali >>
rect -323 699 -217 733
rect -167 699 -121 733
rect -71 699 -25 733
rect 25 699 71 733
rect 121 720 166 733
rect 121 699 127 720
rect 156 699 166 720
rect -323 637 -289 699
rect -209 538 -175 554
rect -209 -554 -175 -538
rect -113 538 -79 554
rect -113 -554 -79 -538
rect -17 538 17 554
rect -17 -554 17 -538
rect 79 538 113 554
rect 79 -554 113 -538
rect 175 538 209 589
rect 175 -554 209 -538
rect -323 -671 -289 -594
rect -323 -705 -217 -671
rect -167 -705 -121 -671
rect -71 -705 -25 -671
rect 25 -705 71 -671
rect 121 -705 157 -671
<< viali >>
rect -209 -538 -175 538
rect -113 -538 -79 538
rect -17 -538 17 538
rect 79 -538 113 538
rect 175 -538 209 538
<< metal1 >>
rect -215 538 -169 550
rect -215 -538 -209 538
rect -175 -538 -169 538
rect -215 -550 -169 -538
rect -119 538 -73 550
rect -119 -538 -113 538
rect -79 -538 -73 538
rect -119 -550 -73 -538
rect -23 538 23 550
rect -23 -538 -17 538
rect 17 -538 23 538
rect -23 -550 23 -538
rect 73 538 119 550
rect 73 -538 79 538
rect 113 -538 119 538
rect 73 -550 119 -538
rect 169 538 215 550
rect 169 -538 175 538
rect 209 -538 215 538
rect 169 -550 215 -538
rect -113 -588 -79 -550
rect 79 -588 113 -550
rect -113 -622 113 -588
<< properties >>
string FIXED_BBOX -306 -716 306 716
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 5.5 l 0.15 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
