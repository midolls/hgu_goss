magic
tech sky130A
magscale 1 2
timestamp 1699479866
<< error_p >>
rect -121 449 -97 473
rect -95 449 -71 473
rect -25 449 -1 473
rect -145 415 -17 449
rect -121 391 -97 415
rect -95 391 -71 415
rect -25 391 -1 415
rect -120 -415 -96 -391
rect -144 -449 -133 -415
rect -120 -473 -96 -449
<< nmos >>
rect -63 -275 -33 275
rect 33 -275 63 275
<< ndiff >>
rect -125 263 -63 275
rect -125 -263 -113 263
rect -79 -263 -63 263
rect -125 -275 -63 -263
rect -33 263 33 275
rect -33 -263 -17 263
rect 17 -263 33 263
rect -33 -275 33 -263
rect 63 263 125 275
rect 63 -263 79 263
rect 113 -263 125 263
rect 63 -275 125 -263
<< ndiffc >>
rect -113 -263 -79 263
rect -17 -263 17 263
rect 79 -263 113 263
<< psubdiff >>
rect 25 415 71 449
rect 121 415 227 449
rect 193 353 227 415
rect 193 -415 227 -353
rect -133 -449 -120 -415
rect -70 -449 -24 -415
rect 26 -449 72 -415
rect 122 -449 227 -415
<< psubdiffcont >>
rect -121 415 -71 449
rect -25 415 25 449
rect 71 415 121 449
rect 193 -353 227 353
rect -120 -449 -70 -415
rect -24 -449 26 -415
rect 72 -449 122 -415
<< poly >>
rect -63 275 -33 301
rect 33 275 63 301
rect -63 -301 -33 -275
rect 33 -301 63 -275
<< locali >>
rect 25 415 71 449
rect 121 415 227 449
rect 193 353 227 415
rect -113 263 -79 279
rect -113 -279 -79 -263
rect -17 263 17 279
rect -17 -314 17 -263
rect 79 263 113 279
rect 79 -314 113 -263
rect -78 -348 113 -314
rect 193 -415 227 -353
rect -133 -449 -120 -415
rect -70 -449 -24 -415
rect 26 -449 72 -415
rect 122 -449 227 -415
<< viali >>
rect -113 -263 -79 263
rect -17 -263 17 263
rect 79 -263 113 263
<< metal1 >>
rect 79 275 113 633
rect -119 263 -73 275
rect -119 -263 -113 263
rect -79 -263 -73 263
rect -119 -275 -73 -263
rect -23 263 23 275
rect -23 -263 -17 263
rect 17 -263 23 263
rect -23 -275 23 -263
rect 73 263 119 275
rect 73 -263 79 263
rect 113 -263 119 263
rect 73 -275 119 -263
<< labels >>
flabel metal1 86 454 109 490 0 FreeSans 320 0 0 0 tah_vp
flabel space -204 1779 -175 1797 0 FreeSans 320 0 0 0 vip
<< properties >>
string FIXED_BBOX -210 -432 210 432
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2.75 l 0.15 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
