** sch_path: /foss/designs/hgu_goss/hgu/tutorial_jh/ring.sch
*.PININFO EN:I OSIL:O GND:I VDD:I
x1 net1 GND GND VDD VDD net2 sky130_fd_sc_hd__inv_1
x5 EN OSIL GND GND VDD VDD net1 sky130_fd_sc_hd__nand2_1
x2 net2 GND GND VDD VDD net3 sky130_fd_sc_hd__inv_1
x3 net3 GND GND VDD VDD net4 sky130_fd_sc_hd__inv_1
x4 net4 GND GND VDD VDD OSIL sky130_fd_sc_hd__inv_1
.end
