magic
tech sky130A
magscale 1 2
timestamp 1698655018
<< checkpaint >>
rect -1260 -2889 1460 1460
rect -1260 -8060 94878 -2889
<< error_s >>
rect 182 3113 240 3119
rect 925 3113 983 3119
rect 1668 3113 1726 3119
rect 2411 3113 2469 3119
rect 3154 3113 3212 3119
rect 3897 3113 3955 3119
rect 4640 3113 4698 3119
rect 5383 3113 5441 3119
rect 6126 3113 6184 3119
rect 6869 3113 6927 3119
rect 7612 3113 7670 3119
rect 8355 3113 8413 3119
rect 9098 3113 9156 3119
rect 9841 3113 9899 3119
rect 10584 3113 10642 3119
rect 11327 3113 11385 3119
rect 12070 3113 12128 3119
rect 12813 3113 12871 3119
rect 13556 3113 13614 3119
rect 14299 3113 14357 3119
rect 15042 3113 15100 3119
rect 15785 3113 15843 3119
rect 16528 3113 16586 3119
rect 17271 3113 17329 3119
rect 18014 3113 18072 3119
rect 18757 3113 18815 3119
rect 19500 3113 19558 3119
rect 20243 3113 20301 3119
rect 20986 3113 21044 3119
rect 21729 3113 21787 3119
rect 22472 3113 22530 3119
rect 23215 3113 23273 3119
rect 23958 3113 24016 3119
rect 24701 3113 24759 3119
rect 25444 3113 25502 3119
rect 26187 3113 26245 3119
rect 26930 3113 26988 3119
rect 27673 3113 27731 3119
rect 28416 3113 28474 3119
rect 29159 3113 29217 3119
rect 29902 3113 29960 3119
rect 30645 3113 30703 3119
rect 31388 3113 31446 3119
rect 32131 3113 32189 3119
rect 32874 3113 32932 3119
rect 33617 3113 33675 3119
rect 34360 3113 34418 3119
rect 35103 3113 35161 3119
rect 35846 3113 35904 3119
rect 36589 3113 36647 3119
rect 37332 3113 37390 3119
rect 38075 3113 38133 3119
rect 38818 3113 38876 3119
rect 39561 3113 39619 3119
rect 40304 3113 40362 3119
rect 41047 3113 41105 3119
rect 41790 3113 41848 3119
rect 42533 3113 42591 3119
rect 43276 3113 43334 3119
rect 44019 3113 44077 3119
rect 44762 3113 44820 3119
rect 45505 3113 45563 3119
rect 46248 3113 46306 3119
rect 46991 3113 47049 3119
rect 47734 3113 47792 3119
rect 48477 3113 48535 3119
rect 49220 3113 49278 3119
rect 49963 3113 50021 3119
rect 50706 3113 50764 3119
rect 51449 3113 51507 3119
rect 52192 3113 52250 3119
rect 52935 3113 52993 3119
rect 53678 3113 53736 3119
rect 54421 3113 54479 3119
rect 55164 3113 55222 3119
rect 55907 3113 55965 3119
rect 56650 3113 56708 3119
rect 57393 3113 57451 3119
rect 58136 3113 58194 3119
rect 58879 3113 58937 3119
rect 59622 3113 59680 3119
rect 60365 3113 60423 3119
rect 61108 3113 61166 3119
rect 61851 3113 61909 3119
rect 62594 3113 62652 3119
rect 63337 3113 63395 3119
rect 64080 3113 64138 3119
rect 64823 3113 64881 3119
rect 65566 3113 65624 3119
rect 66309 3113 66367 3119
rect 67052 3113 67110 3119
rect 67795 3113 67853 3119
rect 68538 3113 68596 3119
rect 69281 3113 69339 3119
rect 70024 3113 70082 3119
rect 70767 3113 70825 3119
rect 71510 3113 71568 3119
rect 72253 3113 72311 3119
rect 72996 3113 73054 3119
rect 73739 3113 73797 3119
rect 74482 3113 74540 3119
rect 75225 3113 75283 3119
rect 75968 3113 76026 3119
rect 76711 3113 76769 3119
rect 77454 3113 77512 3119
rect 78197 3113 78255 3119
rect 78940 3113 78998 3119
rect 79683 3113 79741 3119
rect 80426 3113 80484 3119
rect 81169 3113 81227 3119
rect 81912 3113 81970 3119
rect 82655 3113 82713 3119
rect 83398 3113 83456 3119
rect 84141 3113 84199 3119
rect 84884 3113 84942 3119
rect 85627 3113 85685 3119
rect 86370 3113 86428 3119
rect 87113 3113 87171 3119
rect 87856 3113 87914 3119
rect 88599 3113 88657 3119
rect 89342 3113 89400 3119
rect 90085 3113 90143 3119
rect 90828 3113 90886 3119
rect 91571 3113 91629 3119
rect 92314 3113 92372 3119
rect 93057 3113 93115 3119
rect 93800 3113 93858 3119
rect 182 3079 194 3113
rect 925 3079 937 3113
rect 1668 3079 1680 3113
rect 2411 3079 2423 3113
rect 3154 3079 3166 3113
rect 3897 3079 3909 3113
rect 4640 3079 4652 3113
rect 5383 3079 5395 3113
rect 6126 3079 6138 3113
rect 6869 3079 6881 3113
rect 7612 3079 7624 3113
rect 8355 3079 8367 3113
rect 9098 3079 9110 3113
rect 9841 3079 9853 3113
rect 10584 3079 10596 3113
rect 11327 3079 11339 3113
rect 12070 3079 12082 3113
rect 12813 3079 12825 3113
rect 13556 3079 13568 3113
rect 14299 3079 14311 3113
rect 15042 3079 15054 3113
rect 15785 3079 15797 3113
rect 16528 3079 16540 3113
rect 17271 3079 17283 3113
rect 18014 3079 18026 3113
rect 18757 3079 18769 3113
rect 19500 3079 19512 3113
rect 20243 3079 20255 3113
rect 20986 3079 20998 3113
rect 21729 3079 21741 3113
rect 22472 3079 22484 3113
rect 23215 3079 23227 3113
rect 23958 3079 23970 3113
rect 24701 3079 24713 3113
rect 25444 3079 25456 3113
rect 26187 3079 26199 3113
rect 26930 3079 26942 3113
rect 27673 3079 27685 3113
rect 28416 3079 28428 3113
rect 29159 3079 29171 3113
rect 29902 3079 29914 3113
rect 30645 3079 30657 3113
rect 31388 3079 31400 3113
rect 32131 3079 32143 3113
rect 32874 3079 32886 3113
rect 33617 3079 33629 3113
rect 34360 3079 34372 3113
rect 35103 3079 35115 3113
rect 35846 3079 35858 3113
rect 36589 3079 36601 3113
rect 37332 3079 37344 3113
rect 38075 3079 38087 3113
rect 38818 3079 38830 3113
rect 39561 3079 39573 3113
rect 40304 3079 40316 3113
rect 41047 3079 41059 3113
rect 41790 3079 41802 3113
rect 42533 3079 42545 3113
rect 43276 3079 43288 3113
rect 44019 3079 44031 3113
rect 44762 3079 44774 3113
rect 45505 3079 45517 3113
rect 46248 3079 46260 3113
rect 46991 3079 47003 3113
rect 47734 3079 47746 3113
rect 48477 3079 48489 3113
rect 49220 3079 49232 3113
rect 49963 3079 49975 3113
rect 50706 3079 50718 3113
rect 51449 3079 51461 3113
rect 52192 3079 52204 3113
rect 52935 3079 52947 3113
rect 53678 3079 53690 3113
rect 54421 3079 54433 3113
rect 55164 3079 55176 3113
rect 55907 3079 55919 3113
rect 56650 3079 56662 3113
rect 57393 3079 57405 3113
rect 58136 3079 58148 3113
rect 58879 3079 58891 3113
rect 59622 3079 59634 3113
rect 60365 3079 60377 3113
rect 61108 3079 61120 3113
rect 61851 3079 61863 3113
rect 62594 3079 62606 3113
rect 63337 3079 63349 3113
rect 64080 3079 64092 3113
rect 64823 3079 64835 3113
rect 65566 3079 65578 3113
rect 66309 3079 66321 3113
rect 67052 3079 67064 3113
rect 67795 3079 67807 3113
rect 68538 3079 68550 3113
rect 69281 3079 69293 3113
rect 70024 3079 70036 3113
rect 70767 3079 70779 3113
rect 71510 3079 71522 3113
rect 72253 3079 72265 3113
rect 72996 3079 73008 3113
rect 73739 3079 73751 3113
rect 74482 3079 74494 3113
rect 75225 3079 75237 3113
rect 75968 3079 75980 3113
rect 76711 3079 76723 3113
rect 77454 3079 77466 3113
rect 78197 3079 78209 3113
rect 78940 3079 78952 3113
rect 79683 3079 79695 3113
rect 80426 3079 80438 3113
rect 81169 3079 81181 3113
rect 81912 3079 81924 3113
rect 82655 3079 82667 3113
rect 83398 3079 83410 3113
rect 84141 3079 84153 3113
rect 84884 3079 84896 3113
rect 85627 3079 85639 3113
rect 86370 3079 86382 3113
rect 87113 3079 87125 3113
rect 87856 3079 87868 3113
rect 88599 3079 88611 3113
rect 89342 3079 89354 3113
rect 90085 3079 90097 3113
rect 90828 3079 90840 3113
rect 91571 3079 91583 3113
rect 92314 3079 92326 3113
rect 93057 3079 93069 3113
rect 93800 3079 93812 3113
rect 182 3073 240 3079
rect 925 3073 983 3079
rect 1668 3073 1726 3079
rect 2411 3073 2469 3079
rect 3154 3073 3212 3079
rect 3897 3073 3955 3079
rect 4640 3073 4698 3079
rect 5383 3073 5441 3079
rect 6126 3073 6184 3079
rect 6869 3073 6927 3079
rect 7612 3073 7670 3079
rect 8355 3073 8413 3079
rect 9098 3073 9156 3079
rect 9841 3073 9899 3079
rect 10584 3073 10642 3079
rect 11327 3073 11385 3079
rect 12070 3073 12128 3079
rect 12813 3073 12871 3079
rect 13556 3073 13614 3079
rect 14299 3073 14357 3079
rect 15042 3073 15100 3079
rect 15785 3073 15843 3079
rect 16528 3073 16586 3079
rect 17271 3073 17329 3079
rect 18014 3073 18072 3079
rect 18757 3073 18815 3079
rect 19500 3073 19558 3079
rect 20243 3073 20301 3079
rect 20986 3073 21044 3079
rect 21729 3073 21787 3079
rect 22472 3073 22530 3079
rect 23215 3073 23273 3079
rect 23958 3073 24016 3079
rect 24701 3073 24759 3079
rect 25444 3073 25502 3079
rect 26187 3073 26245 3079
rect 26930 3073 26988 3079
rect 27673 3073 27731 3079
rect 28416 3073 28474 3079
rect 29159 3073 29217 3079
rect 29902 3073 29960 3079
rect 30645 3073 30703 3079
rect 31388 3073 31446 3079
rect 32131 3073 32189 3079
rect 32874 3073 32932 3079
rect 33617 3073 33675 3079
rect 34360 3073 34418 3079
rect 35103 3073 35161 3079
rect 35846 3073 35904 3079
rect 36589 3073 36647 3079
rect 37332 3073 37390 3079
rect 38075 3073 38133 3079
rect 38818 3073 38876 3079
rect 39561 3073 39619 3079
rect 40304 3073 40362 3079
rect 41047 3073 41105 3079
rect 41790 3073 41848 3079
rect 42533 3073 42591 3079
rect 43276 3073 43334 3079
rect 44019 3073 44077 3079
rect 44762 3073 44820 3079
rect 45505 3073 45563 3079
rect 46248 3073 46306 3079
rect 46991 3073 47049 3079
rect 47734 3073 47792 3079
rect 48477 3073 48535 3079
rect 49220 3073 49278 3079
rect 49963 3073 50021 3079
rect 50706 3073 50764 3079
rect 51449 3073 51507 3079
rect 52192 3073 52250 3079
rect 52935 3073 52993 3079
rect 53678 3073 53736 3079
rect 54421 3073 54479 3079
rect 55164 3073 55222 3079
rect 55907 3073 55965 3079
rect 56650 3073 56708 3079
rect 57393 3073 57451 3079
rect 58136 3073 58194 3079
rect 58879 3073 58937 3079
rect 59622 3073 59680 3079
rect 60365 3073 60423 3079
rect 61108 3073 61166 3079
rect 61851 3073 61909 3079
rect 62594 3073 62652 3079
rect 63337 3073 63395 3079
rect 64080 3073 64138 3079
rect 64823 3073 64881 3079
rect 65566 3073 65624 3079
rect 66309 3073 66367 3079
rect 67052 3073 67110 3079
rect 67795 3073 67853 3079
rect 68538 3073 68596 3079
rect 69281 3073 69339 3079
rect 70024 3073 70082 3079
rect 70767 3073 70825 3079
rect 71510 3073 71568 3079
rect 72253 3073 72311 3079
rect 72996 3073 73054 3079
rect 73739 3073 73797 3079
rect 74482 3073 74540 3079
rect 75225 3073 75283 3079
rect 75968 3073 76026 3079
rect 76711 3073 76769 3079
rect 77454 3073 77512 3079
rect 78197 3073 78255 3079
rect 78940 3073 78998 3079
rect 79683 3073 79741 3079
rect 80426 3073 80484 3079
rect 81169 3073 81227 3079
rect 81912 3073 81970 3079
rect 82655 3073 82713 3079
rect 83398 3073 83456 3079
rect 84141 3073 84199 3079
rect 84884 3073 84942 3079
rect 85627 3073 85685 3079
rect 86370 3073 86428 3079
rect 87113 3073 87171 3079
rect 87856 3073 87914 3079
rect 88599 3073 88657 3079
rect 89342 3073 89400 3079
rect 90085 3073 90143 3079
rect 90828 3073 90886 3079
rect 91571 3073 91629 3079
rect 92314 3073 92372 3079
rect 93057 3073 93115 3079
rect 93800 3073 93858 3079
rect 182 2919 240 2925
rect 925 2919 983 2925
rect 1668 2919 1726 2925
rect 2411 2919 2469 2925
rect 3154 2919 3212 2925
rect 3897 2919 3955 2925
rect 4640 2919 4698 2925
rect 5383 2919 5441 2925
rect 6126 2919 6184 2925
rect 6869 2919 6927 2925
rect 7612 2919 7670 2925
rect 8355 2919 8413 2925
rect 9098 2919 9156 2925
rect 9841 2919 9899 2925
rect 10584 2919 10642 2925
rect 11327 2919 11385 2925
rect 12070 2919 12128 2925
rect 12813 2919 12871 2925
rect 13556 2919 13614 2925
rect 14299 2919 14357 2925
rect 15042 2919 15100 2925
rect 15785 2919 15843 2925
rect 16528 2919 16586 2925
rect 17271 2919 17329 2925
rect 18014 2919 18072 2925
rect 18757 2919 18815 2925
rect 19500 2919 19558 2925
rect 20243 2919 20301 2925
rect 20986 2919 21044 2925
rect 21729 2919 21787 2925
rect 22472 2919 22530 2925
rect 23215 2919 23273 2925
rect 23958 2919 24016 2925
rect 24701 2919 24759 2925
rect 25444 2919 25502 2925
rect 26187 2919 26245 2925
rect 26930 2919 26988 2925
rect 27673 2919 27731 2925
rect 28416 2919 28474 2925
rect 29159 2919 29217 2925
rect 29902 2919 29960 2925
rect 30645 2919 30703 2925
rect 31388 2919 31446 2925
rect 32131 2919 32189 2925
rect 32874 2919 32932 2925
rect 33617 2919 33675 2925
rect 34360 2919 34418 2925
rect 35103 2919 35161 2925
rect 35846 2919 35904 2925
rect 36589 2919 36647 2925
rect 37332 2919 37390 2925
rect 38075 2919 38133 2925
rect 38818 2919 38876 2925
rect 39561 2919 39619 2925
rect 40304 2919 40362 2925
rect 41047 2919 41105 2925
rect 41790 2919 41848 2925
rect 42533 2919 42591 2925
rect 43276 2919 43334 2925
rect 44019 2919 44077 2925
rect 44762 2919 44820 2925
rect 45505 2919 45563 2925
rect 46248 2919 46306 2925
rect 46991 2919 47049 2925
rect 47734 2919 47792 2925
rect 48477 2919 48535 2925
rect 49220 2919 49278 2925
rect 49963 2919 50021 2925
rect 50706 2919 50764 2925
rect 51449 2919 51507 2925
rect 52192 2919 52250 2925
rect 52935 2919 52993 2925
rect 53678 2919 53736 2925
rect 54421 2919 54479 2925
rect 55164 2919 55222 2925
rect 55907 2919 55965 2925
rect 56650 2919 56708 2925
rect 57393 2919 57451 2925
rect 58136 2919 58194 2925
rect 58879 2919 58937 2925
rect 59622 2919 59680 2925
rect 60365 2919 60423 2925
rect 61108 2919 61166 2925
rect 61851 2919 61909 2925
rect 62594 2919 62652 2925
rect 63337 2919 63395 2925
rect 64080 2919 64138 2925
rect 64823 2919 64881 2925
rect 65566 2919 65624 2925
rect 66309 2919 66367 2925
rect 67052 2919 67110 2925
rect 67795 2919 67853 2925
rect 68538 2919 68596 2925
rect 69281 2919 69339 2925
rect 70024 2919 70082 2925
rect 70767 2919 70825 2925
rect 71510 2919 71568 2925
rect 72253 2919 72311 2925
rect 72996 2919 73054 2925
rect 73739 2919 73797 2925
rect 74482 2919 74540 2925
rect 75225 2919 75283 2925
rect 75968 2919 76026 2925
rect 76711 2919 76769 2925
rect 77454 2919 77512 2925
rect 78197 2919 78255 2925
rect 78940 2919 78998 2925
rect 79683 2919 79741 2925
rect 80426 2919 80484 2925
rect 81169 2919 81227 2925
rect 81912 2919 81970 2925
rect 82655 2919 82713 2925
rect 83398 2919 83456 2925
rect 84141 2919 84199 2925
rect 84884 2919 84942 2925
rect 85627 2919 85685 2925
rect 86370 2919 86428 2925
rect 87113 2919 87171 2925
rect 87856 2919 87914 2925
rect 88599 2919 88657 2925
rect 89342 2919 89400 2925
rect 90085 2919 90143 2925
rect 90828 2919 90886 2925
rect 91571 2919 91629 2925
rect 92314 2919 92372 2925
rect 93057 2919 93115 2925
rect 93800 2919 93858 2925
rect 182 2885 194 2919
rect 925 2885 937 2919
rect 1668 2885 1680 2919
rect 2411 2885 2423 2919
rect 3154 2885 3166 2919
rect 3897 2885 3909 2919
rect 4640 2885 4652 2919
rect 5383 2885 5395 2919
rect 6126 2885 6138 2919
rect 6869 2885 6881 2919
rect 7612 2885 7624 2919
rect 8355 2885 8367 2919
rect 9098 2885 9110 2919
rect 9841 2885 9853 2919
rect 10584 2885 10596 2919
rect 11327 2885 11339 2919
rect 12070 2885 12082 2919
rect 12813 2885 12825 2919
rect 13556 2885 13568 2919
rect 14299 2885 14311 2919
rect 15042 2885 15054 2919
rect 15785 2885 15797 2919
rect 16528 2885 16540 2919
rect 17271 2885 17283 2919
rect 18014 2885 18026 2919
rect 18757 2885 18769 2919
rect 19500 2885 19512 2919
rect 20243 2885 20255 2919
rect 20986 2885 20998 2919
rect 21729 2885 21741 2919
rect 22472 2885 22484 2919
rect 23215 2885 23227 2919
rect 23958 2885 23970 2919
rect 24701 2885 24713 2919
rect 25444 2885 25456 2919
rect 26187 2885 26199 2919
rect 26930 2885 26942 2919
rect 27673 2885 27685 2919
rect 28416 2885 28428 2919
rect 29159 2885 29171 2919
rect 29902 2885 29914 2919
rect 30645 2885 30657 2919
rect 31388 2885 31400 2919
rect 32131 2885 32143 2919
rect 32874 2885 32886 2919
rect 33617 2885 33629 2919
rect 34360 2885 34372 2919
rect 35103 2885 35115 2919
rect 35846 2885 35858 2919
rect 36589 2885 36601 2919
rect 37332 2885 37344 2919
rect 38075 2885 38087 2919
rect 38818 2885 38830 2919
rect 39561 2885 39573 2919
rect 40304 2885 40316 2919
rect 41047 2885 41059 2919
rect 41790 2885 41802 2919
rect 42533 2885 42545 2919
rect 43276 2885 43288 2919
rect 44019 2885 44031 2919
rect 44762 2885 44774 2919
rect 45505 2885 45517 2919
rect 46248 2885 46260 2919
rect 46991 2885 47003 2919
rect 47734 2885 47746 2919
rect 48477 2885 48489 2919
rect 49220 2885 49232 2919
rect 49963 2885 49975 2919
rect 50706 2885 50718 2919
rect 51449 2885 51461 2919
rect 52192 2885 52204 2919
rect 52935 2885 52947 2919
rect 53678 2885 53690 2919
rect 54421 2885 54433 2919
rect 55164 2885 55176 2919
rect 55907 2885 55919 2919
rect 56650 2885 56662 2919
rect 57393 2885 57405 2919
rect 58136 2885 58148 2919
rect 58879 2885 58891 2919
rect 59622 2885 59634 2919
rect 60365 2885 60377 2919
rect 61108 2885 61120 2919
rect 61851 2885 61863 2919
rect 62594 2885 62606 2919
rect 63337 2885 63349 2919
rect 64080 2885 64092 2919
rect 64823 2885 64835 2919
rect 65566 2885 65578 2919
rect 66309 2885 66321 2919
rect 67052 2885 67064 2919
rect 67795 2885 67807 2919
rect 68538 2885 68550 2919
rect 69281 2885 69293 2919
rect 70024 2885 70036 2919
rect 70767 2885 70779 2919
rect 71510 2885 71522 2919
rect 72253 2885 72265 2919
rect 72996 2885 73008 2919
rect 73739 2885 73751 2919
rect 74482 2885 74494 2919
rect 75225 2885 75237 2919
rect 75968 2885 75980 2919
rect 76711 2885 76723 2919
rect 77454 2885 77466 2919
rect 78197 2885 78209 2919
rect 78940 2885 78952 2919
rect 79683 2885 79695 2919
rect 80426 2885 80438 2919
rect 81169 2885 81181 2919
rect 81912 2885 81924 2919
rect 82655 2885 82667 2919
rect 83398 2885 83410 2919
rect 84141 2885 84153 2919
rect 84884 2885 84896 2919
rect 85627 2885 85639 2919
rect 86370 2885 86382 2919
rect 87113 2885 87125 2919
rect 87856 2885 87868 2919
rect 88599 2885 88611 2919
rect 89342 2885 89354 2919
rect 90085 2885 90097 2919
rect 90828 2885 90840 2919
rect 91571 2885 91583 2919
rect 92314 2885 92326 2919
rect 93057 2885 93069 2919
rect 93800 2885 93812 2919
rect 182 2879 240 2885
rect 925 2879 983 2885
rect 1668 2879 1726 2885
rect 2411 2879 2469 2885
rect 3154 2879 3212 2885
rect 3897 2879 3955 2885
rect 4640 2879 4698 2885
rect 5383 2879 5441 2885
rect 6126 2879 6184 2885
rect 6869 2879 6927 2885
rect 7612 2879 7670 2885
rect 8355 2879 8413 2885
rect 9098 2879 9156 2885
rect 9841 2879 9899 2885
rect 10584 2879 10642 2885
rect 11327 2879 11385 2885
rect 12070 2879 12128 2885
rect 12813 2879 12871 2885
rect 13556 2879 13614 2885
rect 14299 2879 14357 2885
rect 15042 2879 15100 2885
rect 15785 2879 15843 2885
rect 16528 2879 16586 2885
rect 17271 2879 17329 2885
rect 18014 2879 18072 2885
rect 18757 2879 18815 2885
rect 19500 2879 19558 2885
rect 20243 2879 20301 2885
rect 20986 2879 21044 2885
rect 21729 2879 21787 2885
rect 22472 2879 22530 2885
rect 23215 2879 23273 2885
rect 23958 2879 24016 2885
rect 24701 2879 24759 2885
rect 25444 2879 25502 2885
rect 26187 2879 26245 2885
rect 26930 2879 26988 2885
rect 27673 2879 27731 2885
rect 28416 2879 28474 2885
rect 29159 2879 29217 2885
rect 29902 2879 29960 2885
rect 30645 2879 30703 2885
rect 31388 2879 31446 2885
rect 32131 2879 32189 2885
rect 32874 2879 32932 2885
rect 33617 2879 33675 2885
rect 34360 2879 34418 2885
rect 35103 2879 35161 2885
rect 35846 2879 35904 2885
rect 36589 2879 36647 2885
rect 37332 2879 37390 2885
rect 38075 2879 38133 2885
rect 38818 2879 38876 2885
rect 39561 2879 39619 2885
rect 40304 2879 40362 2885
rect 41047 2879 41105 2885
rect 41790 2879 41848 2885
rect 42533 2879 42591 2885
rect 43276 2879 43334 2885
rect 44019 2879 44077 2885
rect 44762 2879 44820 2885
rect 45505 2879 45563 2885
rect 46248 2879 46306 2885
rect 46991 2879 47049 2885
rect 47734 2879 47792 2885
rect 48477 2879 48535 2885
rect 49220 2879 49278 2885
rect 49963 2879 50021 2885
rect 50706 2879 50764 2885
rect 51449 2879 51507 2885
rect 52192 2879 52250 2885
rect 52935 2879 52993 2885
rect 53678 2879 53736 2885
rect 54421 2879 54479 2885
rect 55164 2879 55222 2885
rect 55907 2879 55965 2885
rect 56650 2879 56708 2885
rect 57393 2879 57451 2885
rect 58136 2879 58194 2885
rect 58879 2879 58937 2885
rect 59622 2879 59680 2885
rect 60365 2879 60423 2885
rect 61108 2879 61166 2885
rect 61851 2879 61909 2885
rect 62594 2879 62652 2885
rect 63337 2879 63395 2885
rect 64080 2879 64138 2885
rect 64823 2879 64881 2885
rect 65566 2879 65624 2885
rect 66309 2879 66367 2885
rect 67052 2879 67110 2885
rect 67795 2879 67853 2885
rect 68538 2879 68596 2885
rect 69281 2879 69339 2885
rect 70024 2879 70082 2885
rect 70767 2879 70825 2885
rect 71510 2879 71568 2885
rect 72253 2879 72311 2885
rect 72996 2879 73054 2885
rect 73739 2879 73797 2885
rect 74482 2879 74540 2885
rect 75225 2879 75283 2885
rect 75968 2879 76026 2885
rect 76711 2879 76769 2885
rect 77454 2879 77512 2885
rect 78197 2879 78255 2885
rect 78940 2879 78998 2885
rect 79683 2879 79741 2885
rect 80426 2879 80484 2885
rect 81169 2879 81227 2885
rect 81912 2879 81970 2885
rect 82655 2879 82713 2885
rect 83398 2879 83456 2885
rect 84141 2879 84199 2885
rect 84884 2879 84942 2885
rect 85627 2879 85685 2885
rect 86370 2879 86428 2885
rect 87113 2879 87171 2885
rect 87856 2879 87914 2885
rect 88599 2879 88657 2885
rect 89342 2879 89400 2885
rect 90085 2879 90143 2885
rect 90828 2879 90886 2885
rect 91571 2879 91629 2885
rect 92314 2879 92372 2885
rect 93057 2879 93115 2885
rect 93800 2879 93858 2885
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
rect 0 -2400 200 -2200
rect 0 -2800 200 -2600
rect 0 -3200 200 -3000
rect 0 -3600 200 -3400
rect 0 -4000 200 -3800
rect 0 -4400 200 -4200
rect 0 -4800 200 -4600
rect 0 -5200 200 -5000
rect 0 -5600 200 -5400
rect 0 -6000 200 -5800
rect 0 -6400 200 -6200
rect 0 -6800 200 -6600
use hgu_inverter  hgu_inverter_0
timestamp 1698632956
transform 1 0 46862 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x1
timestamp 1698632956
transform 1 0 47605 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x2[0]
timestamp 1698632956
transform 1 0 48348 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x2[0]
timestamp 1698632956
transform 1 0 49091 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x2[1]
timestamp 1698632956
transform 1 0 47605 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x2[1]
timestamp 1698632956
transform 1 0 48348 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x3[0]
timestamp 1698632956
transform 1 0 51320 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x3[0]
timestamp 1698632956
transform 1 0 52063 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x3[1]
timestamp 1698632956
transform 1 0 50577 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x3[1]
timestamp 1698632956
transform 1 0 51320 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x3[2]
timestamp 1698632956
transform 1 0 49834 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x3[2]
timestamp 1698632956
transform 1 0 50577 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x3[3]
timestamp 1698632956
transform 1 0 49091 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x3[3]
timestamp 1698632956
transform 1 0 49834 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x4[0]
timestamp 1698632956
transform 1 0 57264 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x4[0]
timestamp 1698632956
transform 1 0 58007 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x4[1]
timestamp 1698632956
transform 1 0 56521 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x4[1]
timestamp 1698632956
transform 1 0 57264 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x4[2]
timestamp 1698632956
transform 1 0 55778 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x4[2]
timestamp 1698632956
transform 1 0 56521 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x4[3]
timestamp 1698632956
transform 1 0 55035 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x4[3]
timestamp 1698632956
transform 1 0 55778 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x4[4]
timestamp 1698632956
transform 1 0 54292 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x4[4]
timestamp 1698632956
transform 1 0 55035 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x4[5]
timestamp 1698632956
transform 1 0 53549 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x4[5]
timestamp 1698632956
transform 1 0 54292 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x4[6]
timestamp 1698632956
transform 1 0 52806 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x4[6]
timestamp 1698632956
transform 1 0 53549 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x4[7]
timestamp 1698632956
transform 1 0 52063 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x4[7]
timestamp 1698632956
transform 1 0 52806 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x5[0]
timestamp 1698632956
transform 1 0 69152 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x5[0]
timestamp 1698632956
transform 1 0 69895 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x5[1]
timestamp 1698632956
transform 1 0 68409 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x5[1]
timestamp 1698632956
transform 1 0 69152 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x5[2]
timestamp 1698632956
transform 1 0 67666 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x5[2]
timestamp 1698632956
transform 1 0 68409 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x5[3]
timestamp 1698632956
transform 1 0 66923 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x5[3]
timestamp 1698632956
transform 1 0 67666 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x5[4]
timestamp 1698632956
transform 1 0 66180 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x5[4]
timestamp 1698632956
transform 1 0 66923 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x5[5]
timestamp 1698632956
transform 1 0 65437 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x5[5]
timestamp 1698632956
transform 1 0 66180 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x5[6]
timestamp 1698632956
transform 1 0 64694 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x5[6]
timestamp 1698632956
transform 1 0 65437 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x5[7]
timestamp 1698632956
transform 1 0 63951 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x5[7]
timestamp 1698632956
transform 1 0 64694 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x5[8]
timestamp 1698632956
transform 1 0 63208 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x5[8]
timestamp 1698632956
transform 1 0 63951 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x5[9]
timestamp 1698632956
transform 1 0 62465 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x5[9]
timestamp 1698632956
transform 1 0 63208 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x5[10]
timestamp 1698632956
transform 1 0 61722 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x5[10]
timestamp 1698632956
transform 1 0 62465 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x5[11]
timestamp 1698632956
transform 1 0 60979 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x5[11]
timestamp 1698632956
transform 1 0 61722 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x5[12]
timestamp 1698632956
transform 1 0 60236 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x5[12]
timestamp 1698632956
transform 1 0 60979 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x5[13]
timestamp 1698632956
transform 1 0 59493 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x5[13]
timestamp 1698632956
transform 1 0 60236 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x5[14]
timestamp 1698632956
transform 1 0 58750 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x5[14]
timestamp 1698632956
transform 1 0 59493 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x5[15]
timestamp 1698632956
transform 1 0 58007 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x5[15]
timestamp 1698632956
transform 1 0 58750 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x6[0]
timestamp 1698632956
transform 1 0 92928 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x6[0]
timestamp 1698632956
transform 1 0 93671 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x6[1]
timestamp 1698632956
transform 1 0 92185 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x6[1]
timestamp 1698632956
transform 1 0 92928 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x6[2]
timestamp 1698632956
transform 1 0 91442 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x6[2]
timestamp 1698632956
transform 1 0 92185 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x6[3]
timestamp 1698632956
transform 1 0 90699 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x6[3]
timestamp 1698632956
transform 1 0 91442 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x6[4]
timestamp 1698632956
transform 1 0 89956 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x6[4]
timestamp 1698632956
transform 1 0 90699 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x6[5]
timestamp 1698632956
transform 1 0 89213 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x6[5]
timestamp 1698632956
transform 1 0 89956 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x6[6]
timestamp 1698632956
transform 1 0 88470 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x6[6]
timestamp 1698632956
transform 1 0 89213 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x6[7]
timestamp 1698632956
transform 1 0 87727 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x6[7]
timestamp 1698632956
transform 1 0 88470 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x6[8]
timestamp 1698632956
transform 1 0 86984 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x6[8]
timestamp 1698632956
transform 1 0 87727 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x6[9]
timestamp 1698632956
transform 1 0 86241 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x6[9]
timestamp 1698632956
transform 1 0 86984 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x6[10]
timestamp 1698632956
transform 1 0 85498 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x6[10]
timestamp 1698632956
transform 1 0 86241 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x6[11]
timestamp 1698632956
transform 1 0 84755 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x6[11]
timestamp 1698632956
transform 1 0 85498 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x6[12]
timestamp 1698632956
transform 1 0 84012 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x6[12]
timestamp 1698632956
transform 1 0 84755 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x6[13]
timestamp 1698632956
transform 1 0 83269 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x6[13]
timestamp 1698632956
transform 1 0 84012 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x6[14]
timestamp 1698632956
transform 1 0 82526 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x6[14]
timestamp 1698632956
transform 1 0 83269 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x6[15]
timestamp 1698632956
transform 1 0 81783 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x6[15]
timestamp 1698632956
transform 1 0 82526 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x6[16]
timestamp 1698632956
transform 1 0 81040 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x6[16]
timestamp 1698632956
transform 1 0 81783 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x6[17]
timestamp 1698632956
transform 1 0 80297 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x6[17]
timestamp 1698632956
transform 1 0 81040 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x6[18]
timestamp 1698632956
transform 1 0 79554 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x6[18]
timestamp 1698632956
transform 1 0 80297 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x6[19]
timestamp 1698632956
transform 1 0 78811 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x6[19]
timestamp 1698632956
transform 1 0 79554 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x6[20]
timestamp 1698632956
transform 1 0 78068 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x6[20]
timestamp 1698632956
transform 1 0 78811 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x6[21]
timestamp 1698632956
transform 1 0 77325 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x6[21]
timestamp 1698632956
transform 1 0 78068 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x6[22]
timestamp 1698632956
transform 1 0 76582 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x6[22]
timestamp 1698632956
transform 1 0 77325 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x6[23]
timestamp 1698632956
transform 1 0 75839 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x6[23]
timestamp 1698632956
transform 1 0 76582 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x6[24]
timestamp 1698632956
transform 1 0 75096 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x6[24]
timestamp 1698632956
transform 1 0 75839 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x6[25]
timestamp 1698632956
transform 1 0 74353 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x6[25]
timestamp 1698632956
transform 1 0 75096 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x6[26]
timestamp 1698632956
transform 1 0 73610 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x6[26]
timestamp 1698632956
transform 1 0 74353 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x6[27]
timestamp 1698632956
transform 1 0 72867 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x6[27]
timestamp 1698632956
transform 1 0 73610 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x6[28]
timestamp 1698632956
transform 1 0 72124 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x6[28]
timestamp 1698632956
transform 1 0 72867 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x6[29]
timestamp 1698632956
transform 1 0 71381 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x6[29]
timestamp 1698632956
transform 1 0 72124 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x6[30]
timestamp 1698632956
transform 1 0 70638 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x6[30]
timestamp 1698632956
transform 1 0 71381 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x6[31]
timestamp 1698632956
transform 1 0 69895 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x6[31]
timestamp 1698632956
transform 1 0 70638 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x7[0]
timestamp 1698632956
transform 1 0 46119 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x7[0]
timestamp 1698632956
transform 1 0 46862 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x7[1]
timestamp 1698632956
transform 1 0 45376 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x7[1]
timestamp 1698632956
transform 1 0 46119 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x7[2]
timestamp 1698632956
transform 1 0 44633 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x7[2]
timestamp 1698632956
transform 1 0 45376 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x7[3]
timestamp 1698632956
transform 1 0 43890 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x7[3]
timestamp 1698632956
transform 1 0 44633 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x7[4]
timestamp 1698632956
transform 1 0 43147 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x7[4]
timestamp 1698632956
transform 1 0 43890 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x7[5]
timestamp 1698632956
transform 1 0 42404 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x7[5]
timestamp 1698632956
transform 1 0 43147 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x7[6]
timestamp 1698632956
transform 1 0 41661 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x7[6]
timestamp 1698632956
transform 1 0 42404 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x7[7]
timestamp 1698632956
transform 1 0 40918 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x7[7]
timestamp 1698632956
transform 1 0 41661 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x7[8]
timestamp 1698632956
transform 1 0 40175 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x7[8]
timestamp 1698632956
transform 1 0 40918 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x7[9]
timestamp 1698632956
transform 1 0 39432 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x7[9]
timestamp 1698632956
transform 1 0 40175 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x7[10]
timestamp 1698632956
transform 1 0 38689 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x7[10]
timestamp 1698632956
transform 1 0 39432 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x7[11]
timestamp 1698632956
transform 1 0 37946 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x7[11]
timestamp 1698632956
transform 1 0 38689 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x7[12]
timestamp 1698632956
transform 1 0 37203 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x7[12]
timestamp 1698632956
transform 1 0 37946 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x7[13]
timestamp 1698632956
transform 1 0 36460 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x7[13]
timestamp 1698632956
transform 1 0 37203 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x7[14]
timestamp 1698632956
transform 1 0 35717 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x7[14]
timestamp 1698632956
transform 1 0 36460 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x7[15]
timestamp 1698632956
transform 1 0 34974 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x7[15]
timestamp 1698632956
transform 1 0 35717 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x7[16]
timestamp 1698632956
transform 1 0 34231 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x7[16]
timestamp 1698632956
transform 1 0 34974 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x7[17]
timestamp 1698632956
transform 1 0 33488 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x7[17]
timestamp 1698632956
transform 1 0 34231 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x7[18]
timestamp 1698632956
transform 1 0 32745 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x7[18]
timestamp 1698632956
transform 1 0 33488 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x7[19]
timestamp 1698632956
transform 1 0 32002 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x7[19]
timestamp 1698632956
transform 1 0 32745 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x7[20]
timestamp 1698632956
transform 1 0 31259 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x7[20]
timestamp 1698632956
transform 1 0 32002 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x7[21]
timestamp 1698632956
transform 1 0 30516 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x7[21]
timestamp 1698632956
transform 1 0 31259 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x7[22]
timestamp 1698632956
transform 1 0 29773 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x7[22]
timestamp 1698632956
transform 1 0 30516 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x7[23]
timestamp 1698632956
transform 1 0 29030 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x7[23]
timestamp 1698632956
transform 1 0 29773 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x7[24]
timestamp 1698632956
transform 1 0 28287 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x7[24]
timestamp 1698632956
transform 1 0 29030 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x7[25]
timestamp 1698632956
transform 1 0 27544 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x7[25]
timestamp 1698632956
transform 1 0 28287 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x7[26]
timestamp 1698632956
transform 1 0 26801 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x7[26]
timestamp 1698632956
transform 1 0 27544 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x7[27]
timestamp 1698632956
transform 1 0 26058 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x7[27]
timestamp 1698632956
transform 1 0 26801 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x7[28]
timestamp 1698632956
transform 1 0 25315 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x7[28]
timestamp 1698632956
transform 1 0 26058 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x7[29]
timestamp 1698632956
transform 1 0 24572 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x7[29]
timestamp 1698632956
transform 1 0 25315 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x7[30]
timestamp 1698632956
transform 1 0 23829 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x7[30]
timestamp 1698632956
transform 1 0 24572 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x7[31]
timestamp 1698632956
transform 1 0 23086 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x7[31]
timestamp 1698632956
transform 1 0 23829 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x7[32]
timestamp 1698632956
transform 1 0 22343 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x7[32]
timestamp 1698632956
transform 1 0 23086 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x7[33]
timestamp 1698632956
transform 1 0 21600 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x7[33]
timestamp 1698632956
transform 1 0 22343 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x7[34]
timestamp 1698632956
transform 1 0 20857 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x7[34]
timestamp 1698632956
transform 1 0 21600 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x7[35]
timestamp 1698632956
transform 1 0 20114 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x7[35]
timestamp 1698632956
transform 1 0 20857 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x7[36]
timestamp 1698632956
transform 1 0 19371 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x7[36]
timestamp 1698632956
transform 1 0 20114 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x7[37]
timestamp 1698632956
transform 1 0 18628 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x7[37]
timestamp 1698632956
transform 1 0 19371 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x7[38]
timestamp 1698632956
transform 1 0 17885 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x7[38]
timestamp 1698632956
transform 1 0 18628 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x7[39]
timestamp 1698632956
transform 1 0 17142 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x7[39]
timestamp 1698632956
transform 1 0 17885 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x7[40]
timestamp 1698632956
transform 1 0 16399 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x7[40]
timestamp 1698632956
transform 1 0 17142 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x7[41]
timestamp 1698632956
transform 1 0 15656 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x7[41]
timestamp 1698632956
transform 1 0 16399 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x7[42]
timestamp 1698632956
transform 1 0 14913 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x7[42]
timestamp 1698632956
transform 1 0 15656 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x7[43]
timestamp 1698632956
transform 1 0 14170 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x7[43]
timestamp 1698632956
transform 1 0 14913 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x7[44]
timestamp 1698632956
transform 1 0 13427 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x7[44]
timestamp 1698632956
transform 1 0 14170 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x7[45]
timestamp 1698632956
transform 1 0 12684 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x7[45]
timestamp 1698632956
transform 1 0 13427 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x7[46]
timestamp 1698632956
transform 1 0 11941 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x7[46]
timestamp 1698632956
transform 1 0 12684 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x7[47]
timestamp 1698632956
transform 1 0 11198 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x7[47]
timestamp 1698632956
transform 1 0 11941 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x7[48]
timestamp 1698632956
transform 1 0 10455 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x7[48]
timestamp 1698632956
transform 1 0 11198 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x7[49]
timestamp 1698632956
transform 1 0 9712 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x7[49]
timestamp 1698632956
transform 1 0 10455 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x7[50]
timestamp 1698632956
transform 1 0 8969 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x7[50]
timestamp 1698632956
transform 1 0 9712 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x7[51]
timestamp 1698632956
transform 1 0 8226 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x7[51]
timestamp 1698632956
transform 1 0 8969 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x7[52]
timestamp 1698632956
transform 1 0 7483 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x7[52]
timestamp 1698632956
transform 1 0 8226 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x7[53]
timestamp 1698632956
transform 1 0 6740 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x7[53]
timestamp 1698632956
transform 1 0 7483 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x7[54]
timestamp 1698632956
transform 1 0 5997 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x7[54]
timestamp 1698632956
transform 1 0 6740 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x7[55]
timestamp 1698632956
transform 1 0 5254 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x7[55]
timestamp 1698632956
transform 1 0 5997 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x7[56]
timestamp 1698632956
transform 1 0 4511 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x7[56]
timestamp 1698632956
transform 1 0 5254 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x7[57]
timestamp 1698632956
transform 1 0 3768 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x7[57]
timestamp 1698632956
transform 1 0 4511 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x7[58]
timestamp 1698632956
transform 1 0 3025 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x7[58]
timestamp 1698632956
transform 1 0 3768 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x7[59]
timestamp 1698632956
transform 1 0 2282 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x7[59]
timestamp 1698632956
transform 1 0 3025 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x7[60]
timestamp 1698632956
transform 1 0 1539 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x7[60]
timestamp 1698632956
transform 1 0 2282 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x7[61]
timestamp 1698632956
transform 1 0 796 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x7[61]
timestamp 1698632956
transform 1 0 1539 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x7[62]
timestamp 1698632956
transform 1 0 53 0 1 -5200
box -53 -1600 690 1051
use hgu_inverter  x7[62]
timestamp 1698632956
transform 1 0 796 0 1 2200
box -53 -1600 690 1051
use hgu_inverter  x7[63]
timestamp 1698632956
transform 1 0 53 0 1 2200
box -53 -1600 690 1051
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 VREF
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 SAR<4>
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 SAR<1>
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 SAR<2>
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 SAR<3>
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 SAR<5>
port 5 nsew
flabel metal1 0 -2400 200 -2200 0 FreeSans 256 0 0 0 SAR<6>
port 6 nsew
flabel metal1 0 -2800 200 -2600 0 FreeSans 256 0 0 0 SAR<0>
port 7 nsew
flabel metal1 0 -3200 200 -3000 0 FreeSans 256 0 0 0 C<3:0>
port 8 nsew
flabel metal1 0 -3600 200 -3400 0 FreeSans 256 0 0 0 C<7:0>
port 9 nsew
flabel metal1 0 -4000 200 -3800 0 FreeSans 256 0 0 0 C<15:0>
port 10 nsew
flabel metal1 0 -4400 200 -4200 0 FreeSans 256 0 0 0 {}
port 11 nsew
flabel metal1 0 -4800 200 -4600 0 FreeSans 256 0 0 0 C<31:0>
port 12 nsew
flabel metal1 0 -5200 200 -5000 0 FreeSans 256 0 0 0 C<0>
port 13 nsew
flabel metal1 0 -5600 200 -5400 0 FreeSans 256 0 0 0 C<1:0>
port 14 nsew
flabel metal1 0 -6000 200 -5800 0 FreeSans 256 0 0 0 C<63:0>
port 15 nsew
flabel metal1 0 -6400 200 -6200 0 FreeSans 256 0 0 0 VSS
port 16 nsew
flabel metal1 0 -6800 200 -6600 0 FreeSans 256 0 0 0 VDD
port 17 nsew
<< end >>
