magic
tech sky130A
timestamp 1697298256
<< checkpaint >>
rect -630 -330 1016 1170
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  XC2
timestamp 0
transform 1 0 193 0 1 420
box -193 -120 193 120
<< end >>
