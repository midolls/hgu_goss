* NGSPICE file created from hgu_cdac_cap_8.ext - technology: sky130A


* Top level circuit hgu_cdac_cap_8

C0 hgu_cdac_cap_4_1.hgu_cdac_cap_2_1.hgu_cdac_unit_1.C1 hgu_cdac_cap_4_0.hgu_cdac_cap_2_1.hgu_cdac_unit_1.C0 4.31f
C1 hgu_cdac_cap_4_1.hgu_cdac_cap_2_1.hgu_cdac_unit_1.C1 hgu_cdac_cap_4_1.hgu_cdac_cap_2_0.hgu_cdac_unit_1.C0 4.31f
C2 hgu_cdac_cap_4_1.hgu_cdac_cap_2_1.hgu_cdac_unit_1.C0 hgu_cdac_cap_4_1.hgu_cdac_cap_2_1.hgu_cdac_unit_1.C1 4.31f
C3 hgu_cdac_cap_4_1.hgu_cdac_cap_2_1.hgu_cdac_unit_1.C1 hgu_cdac_cap_4_1.hgu_cdac_cap_2_1.hgu_cdac_unit_0.C1 17.7f
C4 hgu_cdac_cap_4_1.hgu_cdac_cap_2_1.hgu_cdac_unit_1.C1 hgu_cdac_cap_4_0.hgu_cdac_cap_2_0.hgu_cdac_unit_1.C0 4.31f
C5 hgu_cdac_cap_4_1.hgu_cdac_cap_2_1.hgu_cdac_unit_1.C1 VSUBS 2.53f $ **FLOATING
C6 hgu_cdac_cap_4_1.hgu_cdac_cap_2_1.hgu_cdac_unit_0.C1 VSUBS 2.6f $ **FLOATING
.end

