magic
tech sky130A
magscale 1 2
timestamp 1697717772
<< error_p >>
rect 73 34 119 49
rect -23 5 23 18
rect -23 -30 -17 5
rect 73 0 79 34
rect 73 -12 119 0
rect -23 -42 23 -30
rect -17 -44 17 -42
<< nmos >>
rect -63 -42 -33 42
rect 33 -42 63 42
<< ndiff >>
rect -125 30 -63 42
rect -125 -30 -113 30
rect -79 -30 -63 30
rect -125 -42 -63 -30
rect -33 5 33 42
rect -33 -30 -17 5
rect 17 -30 33 5
rect -33 -42 33 -30
rect 63 34 125 42
rect 63 0 79 34
rect 113 0 125 34
rect 63 -42 125 0
rect -17 -44 17 -42
<< ndiffc >>
rect -113 -30 -79 30
rect -17 -30 17 5
rect 79 0 113 34
<< poly >>
rect -63 42 -33 68
rect 33 42 63 68
rect -63 -64 -33 -42
rect -81 -80 -15 -64
rect 33 -68 63 -42
rect -81 -114 -65 -80
rect -31 -114 -15 -80
rect -81 -130 -15 -114
<< polycont >>
rect -65 -114 -31 -80
<< locali >>
rect -113 30 -79 46
rect -113 -46 -79 -30
rect -17 5 17 46
rect -17 -46 17 -30
rect 79 34 113 52
rect 79 -45 113 0
rect -81 -114 -65 -80
rect -31 -114 -15 -80
<< viali >>
rect -113 -30 -79 30
rect -17 -30 17 5
rect 79 0 113 34
<< metal1 >>
rect -119 30 -73 46
rect -119 -30 -113 30
rect -79 -30 -73 30
rect 73 34 119 49
rect -119 -42 -73 -30
rect -23 5 23 18
rect -23 -30 -17 5
rect 17 -30 23 5
rect 73 0 79 34
rect 113 0 119 34
rect 73 -12 119 0
rect -23 -42 23 -30
rect -17 -44 17 -42
<< properties >>
string FIXED_BBOX -210 -199 210 199
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.42 l 0.15 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
