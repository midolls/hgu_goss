magic
tech sky130A
magscale 1 2
timestamp 1701186871
<< nwell >>
rect 11513 8777 11713 8794
rect 11513 8765 11968 8777
rect 11513 8048 11815 8765
rect 24490 7367 26123 7481
<< metal1 >>
rect 13198 12668 13224 12702
rect 19914 12668 19940 12702
rect 2324 12193 2356 12227
rect 10869 12169 10912 12233
rect 2330 11810 2393 11857
rect 10914 11288 11232 11530
rect 13479 10913 13504 10941
rect 13481 10857 13506 10885
rect 13483 10801 13508 10829
rect 13484 10745 13509 10773
rect 13486 10689 13511 10717
rect 13485 10633 13510 10661
rect 13473 10493 13506 10605
rect 2930 10449 4871 10477
rect 13482 10438 13506 10464
rect 2931 10393 7297 10421
rect 13484 10382 13510 10408
rect 2929 10337 8154 10365
rect 13486 10326 13512 10352
rect 2928 10281 8154 10309
rect 13482 10270 13508 10296
rect 2932 10225 7297 10253
rect 13486 10214 13512 10240
rect 2930 10169 4871 10197
rect 13484 10158 13510 10184
rect 11827 8983 11873 9018
rect 2324 8419 2366 8453
rect 11771 8426 11874 8460
rect 11771 8122 11799 8426
rect 19956 8407 19982 8441
rect 26659 8407 26685 8441
rect 11563 8066 11799 8122
rect 11750 7849 11836 7855
rect 11802 7834 11836 7849
rect 11802 7806 11830 7834
rect 11859 7831 11887 7839
rect 11750 7790 11802 7797
rect 10305 7481 10311 7533
rect 10363 7522 10369 7533
rect 11743 7522 11749 7532
rect 10363 7494 11749 7522
rect 10363 7481 10369 7494
rect 11743 7480 11749 7494
rect 11801 7480 11807 7532
rect 9945 7358 9951 7410
rect 10003 7358 10009 7410
rect 10623 7282 10629 7334
rect 10681 7323 10687 7334
rect 23915 7323 23921 7333
rect 10681 7295 23921 7323
rect 10681 7282 10687 7295
rect 10623 7281 10687 7282
rect 23915 7281 23921 7295
rect 23973 7281 23979 7333
rect 23915 7280 23979 7281
rect 10922 6824 10956 6858
rect 9982 6744 9988 6796
rect 10040 6788 10046 6796
rect 10040 6754 10952 6788
rect 10040 6744 10046 6754
rect 10927 6687 10962 6722
rect 23937 6371 24075 6405
rect 23914 5985 23921 6037
rect 23973 6035 23979 6037
rect 23973 5988 23980 6035
rect 23973 5985 23979 5988
rect 23914 5984 23979 5985
rect 24237 5786 24349 5834
rect 10311 5240 10363 5246
rect 10363 5197 10949 5231
rect 10311 5182 10363 5188
rect 25545 4635 26484 4663
rect 25545 4579 28910 4607
rect 25545 4523 29767 4551
rect 10623 4311 10630 4363
rect 10682 4354 10688 4363
rect 10682 4320 10949 4354
rect 10682 4311 10688 4320
rect 25226 4155 25511 4203
rect 10933 3942 10967 3977
rect 14907 3096 14914 3148
rect 14966 3143 14972 3148
rect 20834 3143 20840 3149
rect 14966 3115 20840 3143
rect 14966 3096 14972 3115
rect 20834 3097 20840 3115
rect 20892 3097 20898 3149
rect 20996 3097 21002 3149
rect 21054 3142 21060 3149
rect 24881 3142 24887 3155
rect 21054 3114 24887 3142
rect 21054 3097 21060 3114
rect 24881 3103 24887 3114
rect 24940 3142 24946 3155
rect 25226 3142 25254 4155
rect 30445 4145 30754 4193
rect 24940 3114 25254 3142
rect 25282 3951 25525 3999
rect 24940 3103 24946 3114
rect 18599 3018 18605 3086
rect 18657 3069 18663 3086
rect 25282 3069 25310 3951
rect 30455 3815 30764 3863
rect 30447 3516 30756 3564
rect 18657 3041 25310 3069
rect 25338 3308 25528 3356
rect 18657 3018 18663 3041
rect 9983 2924 9989 2976
rect 10041 2965 10047 2976
rect 11905 2965 11911 2978
rect 10041 2937 11911 2965
rect 10041 2924 10047 2937
rect 11905 2926 11911 2937
rect 11963 2926 11969 2978
rect 19695 2961 19701 3013
rect 19753 3003 19759 3013
rect 21245 3003 21251 3013
rect 19753 2975 21251 3003
rect 19753 2961 19759 2975
rect 21245 2961 21251 2975
rect 21303 2961 21309 3013
rect 22486 2961 22493 3013
rect 22545 3003 22551 3013
rect 23380 3003 23386 3013
rect 22545 2975 23386 3003
rect 22545 2961 22551 2975
rect 23380 2961 23386 2975
rect 23438 3003 23444 3013
rect 25338 3003 25366 3308
rect 23438 2975 25366 3003
rect 25394 3174 25529 3222
rect 30461 3174 30770 3222
rect 23438 2961 23444 2975
rect 12518 2904 12524 2956
rect 12576 2949 12583 2956
rect 18429 2949 18435 2954
rect 12576 2907 18435 2949
rect 12576 2904 12583 2907
rect 18429 2902 18435 2907
rect 18487 2902 18494 2954
rect 20092 2892 20099 2944
rect 20151 2933 20157 2944
rect 21076 2933 21082 2944
rect 20151 2905 21082 2933
rect 20151 2892 20157 2905
rect 21076 2892 21082 2905
rect 21134 2933 21140 2944
rect 25394 2933 25422 3174
rect 21134 2905 25422 2933
rect 21134 2892 21140 2905
rect 15309 2824 15316 2876
rect 15368 2864 15374 2876
rect 16296 2864 16302 2877
rect 15368 2836 16302 2864
rect 15368 2824 15374 2836
rect 16296 2825 16302 2836
rect 16354 2864 16360 2877
rect 25504 2864 25549 2886
rect 30450 2864 30759 2912
rect 16354 2836 25549 2864
rect 16354 2825 16360 2836
rect 8498 2735 8505 2787
rect 8557 2773 8563 2787
rect 10303 2773 10310 2783
rect 8557 2745 10310 2773
rect 8557 2735 8563 2745
rect 8498 2734 8563 2735
rect 10303 2731 10310 2745
rect 10362 2731 10368 2783
rect 17701 2756 17708 2808
rect 17760 2797 17766 2808
rect 18685 2797 18691 2808
rect 17760 2769 18691 2797
rect 17760 2756 17766 2769
rect 18685 2756 18691 2769
rect 18743 2797 18750 2808
rect 18743 2769 25550 2797
rect 18743 2756 18750 2769
rect 10303 2730 10368 2731
rect 12922 2700 12928 2752
rect 12980 2728 12987 2752
rect 13898 2728 13904 2752
rect 12980 2700 13904 2728
rect 13956 2728 13963 2752
rect 13956 2700 25477 2728
rect 25505 2711 25550 2769
rect 10529 2637 10535 2689
rect 10587 2672 10594 2689
rect 11509 2672 11515 2686
rect 10587 2644 11515 2672
rect 10587 2637 10594 2644
rect 11509 2634 11515 2644
rect 11567 2672 11574 2686
rect 11567 2644 25420 2672
rect 11567 2634 11574 2644
rect 10126 2568 10132 2620
rect 10184 2605 10191 2620
rect 16033 2605 16039 2614
rect 10184 2577 16039 2605
rect 10184 2568 10191 2577
rect 16033 2562 16039 2577
rect 16091 2562 16097 2614
rect 16434 2561 16440 2613
rect 16492 2605 16498 2613
rect 24475 2605 24482 2616
rect 16492 2577 24482 2605
rect 16492 2561 16498 2577
rect 24475 2564 24482 2577
rect 24534 2564 24540 2616
rect 17301 2496 17307 2548
rect 17359 2537 17366 2548
rect 23224 2537 23230 2549
rect 17359 2509 23230 2537
rect 17359 2496 17366 2509
rect 23224 2497 23230 2509
rect 23282 2497 23288 2549
rect 18857 2429 18863 2481
rect 18915 2469 18922 2481
rect 22083 2469 22089 2481
rect 18915 2441 22089 2469
rect 18915 2429 18922 2441
rect 22083 2429 22089 2441
rect 22141 2429 22147 2481
rect 9823 2360 9829 2412
rect 9881 2401 9887 2412
rect 25247 2401 25253 2413
rect 9881 2371 25253 2401
rect 9881 2360 9887 2371
rect 25247 2361 25253 2371
rect 25305 2361 25312 2413
rect 9736 2291 9742 2343
rect 9794 2332 9800 2343
rect 22853 2332 22859 2342
rect 9794 2302 22859 2332
rect 9794 2291 9800 2302
rect 22853 2290 22859 2302
rect 22911 2290 22918 2342
rect 9649 2222 9655 2274
rect 9707 2262 9713 2274
rect 20462 2262 20468 2271
rect 9707 2232 20468 2262
rect 9707 2222 9713 2232
rect 20462 2219 20468 2232
rect 20520 2219 20527 2271
rect 9563 2152 9569 2204
rect 9621 2192 9627 2204
rect 18070 2192 18076 2203
rect 9621 2162 18076 2192
rect 9621 2152 9627 2162
rect 18070 2151 18076 2162
rect 18128 2151 18135 2203
rect 9477 2082 9483 2134
rect 9535 2123 9541 2134
rect 15679 2123 15685 2133
rect 9535 2093 15685 2123
rect 9535 2082 9541 2093
rect 15679 2081 15685 2093
rect 15737 2081 15744 2133
rect 9390 2013 9396 2065
rect 9448 2053 9454 2065
rect 13285 2053 13291 2064
rect 9448 2023 13291 2053
rect 9448 2013 9454 2023
rect 13285 2012 13291 2023
rect 13343 2012 13350 2064
rect 9304 1943 9310 1995
rect 9362 1983 9368 1995
rect 10893 1983 10899 1994
rect 9362 1953 10899 1983
rect 9362 1943 9368 1953
rect 10893 1942 10899 1953
rect 10951 1942 10958 1994
rect 25391 1942 25420 2644
rect 25448 2141 25477 2700
rect 30456 2533 30765 2581
rect 30453 2237 30762 2285
rect 25448 2093 25551 2141
rect 9218 1873 9224 1925
rect 9276 1913 9282 1925
rect 23055 1913 23061 1924
rect 9276 1883 23061 1913
rect 9276 1873 9282 1883
rect 23055 1872 23061 1883
rect 23113 1872 23120 1924
rect 25391 1894 25509 1942
rect 30451 1893 30760 1941
rect 9132 1803 9138 1855
rect 9190 1844 9196 1855
rect 20666 1844 20672 1854
rect 9190 1814 20672 1844
rect 9190 1803 9196 1814
rect 20666 1802 20672 1814
rect 20724 1802 20731 1854
rect 9045 1734 9051 1786
rect 9103 1774 9109 1786
rect 18273 1774 18279 1785
rect 9103 1744 18279 1774
rect 9103 1734 9109 1744
rect 18273 1733 18279 1744
rect 18331 1733 18338 1785
rect 8959 1664 8965 1716
rect 9017 1705 9023 1716
rect 15880 1705 15886 1715
rect 9017 1675 15886 1705
rect 9017 1664 9023 1675
rect 15880 1663 15886 1675
rect 15938 1663 15945 1715
rect 8872 1595 8878 1647
rect 8930 1635 8936 1647
rect 13488 1635 13494 1646
rect 8930 1605 13494 1635
rect 8930 1595 8936 1605
rect 13488 1594 13494 1605
rect 13546 1594 13553 1646
rect 8786 1525 8792 1577
rect 8844 1565 8850 1577
rect 11098 1565 11104 1575
rect 8844 1535 11104 1565
rect 8844 1525 8850 1535
rect 11098 1523 11104 1535
rect 11156 1523 11163 1575
rect 8489 1164 8497 1216
rect 8549 1164 8555 1216
rect 11910 967 11916 1019
rect 11968 967 11974 1019
<< via1 >>
rect 11750 7797 11802 7849
rect 10311 7481 10363 7533
rect 11749 7480 11801 7532
rect 9951 7358 10003 7410
rect 10629 7282 10681 7334
rect 23921 7281 23973 7333
rect 9988 6744 10040 6796
rect 23921 5985 23973 6037
rect 10311 5188 10363 5240
rect 10630 4311 10682 4363
rect 14914 3096 14966 3148
rect 20840 3097 20892 3149
rect 21002 3097 21054 3149
rect 24887 3103 24940 3155
rect 18605 3018 18657 3086
rect 9989 2924 10041 2976
rect 11911 2926 11963 2978
rect 19701 2961 19753 3013
rect 21251 2961 21303 3013
rect 22493 2961 22545 3013
rect 23386 2961 23438 3013
rect 12524 2904 12576 2956
rect 18435 2902 18487 2954
rect 20099 2892 20151 2944
rect 21082 2892 21134 2944
rect 15316 2824 15368 2876
rect 16302 2825 16354 2877
rect 8505 2735 8557 2787
rect 10310 2731 10362 2783
rect 17708 2756 17760 2808
rect 18691 2756 18743 2808
rect 12928 2700 12980 2752
rect 13904 2700 13956 2752
rect 10535 2637 10587 2689
rect 11515 2634 11567 2686
rect 10132 2568 10184 2620
rect 16039 2562 16091 2614
rect 16440 2561 16492 2613
rect 24482 2564 24534 2616
rect 17307 2496 17359 2548
rect 23230 2497 23282 2549
rect 18863 2429 18915 2481
rect 22089 2429 22141 2481
rect 9829 2360 9881 2412
rect 25253 2361 25305 2413
rect 9742 2291 9794 2343
rect 22859 2290 22911 2342
rect 9655 2222 9707 2274
rect 20468 2219 20520 2271
rect 9569 2152 9621 2204
rect 18076 2151 18128 2203
rect 9483 2082 9535 2134
rect 15685 2081 15737 2133
rect 9396 2013 9448 2065
rect 13291 2012 13343 2064
rect 9310 1943 9362 1995
rect 10899 1942 10951 1994
rect 9224 1873 9276 1925
rect 23061 1872 23113 1924
rect 9138 1803 9190 1855
rect 20672 1802 20724 1854
rect 9051 1734 9103 1786
rect 18279 1733 18331 1785
rect 8965 1664 9017 1716
rect 15886 1663 15938 1715
rect 8878 1595 8930 1647
rect 13494 1594 13546 1646
rect 8792 1525 8844 1577
rect 11104 1523 11156 1575
rect 8497 1164 8549 1216
rect 11916 967 11968 1019
<< metal2 >>
rect 2737 9041 2790 11605
rect 10624 8067 10765 8124
rect 10305 7481 10311 7533
rect 10363 7481 10369 7533
rect 9945 7358 9951 7410
rect 10003 7358 10029 7410
rect 10001 6796 10029 7358
rect 9982 6744 9988 6796
rect 10040 6744 10046 6796
rect 10001 2976 10029 6744
rect 10323 5246 10351 7481
rect 10624 7334 10652 8067
rect 11750 7849 11802 7855
rect 11750 7790 11802 7797
rect 11762 7532 11790 7790
rect 11743 7480 11749 7532
rect 11801 7480 11807 7532
rect 10623 7282 10629 7334
rect 10681 7282 10687 7334
rect 10623 7281 10687 7282
rect 23915 7281 23921 7333
rect 23973 7281 23979 7333
rect 10311 5240 10363 5246
rect 10311 5182 10363 5188
rect 8498 2735 8505 2787
rect 8557 2735 8563 2787
rect 8498 2734 8563 2735
rect 8506 1216 8543 2734
rect 8489 1164 8497 1216
rect 8549 1164 8555 1216
rect 8716 -1261 8758 2925
rect 8798 1577 8840 2925
rect 8882 1647 8924 2925
rect 8970 1716 9012 2925
rect 9057 1786 9099 2925
rect 9143 1855 9185 2925
rect 9229 1925 9271 2925
rect 9316 1995 9358 2925
rect 9402 2065 9444 2925
rect 9488 2134 9530 2925
rect 9575 2204 9617 2925
rect 9660 2274 9702 2925
rect 9747 2343 9789 2925
rect 9834 2412 9876 2925
rect 9983 2924 9989 2976
rect 10041 2924 10047 2976
rect 10323 2783 10351 5182
rect 10642 4363 10670 7281
rect 23915 7280 23979 7281
rect 23933 6037 23963 7280
rect 23914 5985 23921 6037
rect 23973 5985 23979 6037
rect 23914 5984 23979 5985
rect 10623 4311 10630 4363
rect 10682 4311 10688 4363
rect 14907 3096 14914 3148
rect 14966 3096 14972 3148
rect 20834 3097 20840 3149
rect 20892 3097 20898 3149
rect 20996 3097 21002 3149
rect 21054 3097 21060 3149
rect 24881 3103 24887 3155
rect 24940 3103 24946 3155
rect 11905 2926 11911 2978
rect 11963 2926 11969 2978
rect 10303 2731 10310 2783
rect 10362 2731 10368 2783
rect 10303 2730 10368 2731
rect 10529 2637 10535 2689
rect 10587 2637 10594 2689
rect 10126 2568 10132 2620
rect 10184 2568 10191 2620
rect 9823 2360 9829 2412
rect 9881 2360 9887 2412
rect 9736 2291 9742 2343
rect 9794 2291 9800 2343
rect 9649 2222 9655 2274
rect 9707 2222 9713 2274
rect 9563 2152 9569 2204
rect 9621 2152 9627 2204
rect 9477 2082 9483 2134
rect 9535 2082 9541 2134
rect 9390 2013 9396 2065
rect 9448 2013 9454 2065
rect 9304 1943 9310 1995
rect 9362 1943 9368 1995
rect 9218 1873 9224 1925
rect 9276 1873 9282 1925
rect 9132 1803 9138 1855
rect 9190 1803 9196 1855
rect 9045 1734 9051 1786
rect 9103 1734 9109 1786
rect 8959 1664 8965 1716
rect 9017 1664 9023 1716
rect 8872 1595 8878 1647
rect 8930 1595 8936 1647
rect 10137 1602 10179 2568
rect 10539 1676 10581 2637
rect 11509 2634 11515 2686
rect 11567 2634 11574 2686
rect 10893 1942 10899 1994
rect 10951 1942 10958 1994
rect 10905 1728 10947 1942
rect 8786 1525 8792 1577
rect 8844 1525 8850 1577
rect 11098 1523 11104 1575
rect 11156 1523 11163 1575
rect 11922 1019 11950 2926
rect 12518 2904 12524 2956
rect 12576 2904 12583 2956
rect 12529 2703 12571 2904
rect 12528 1703 12571 2703
rect 12922 2700 12928 2752
rect 12980 2700 12987 2752
rect 13898 2700 13904 2752
rect 13956 2700 13963 2752
rect 12931 1714 12973 2700
rect 13913 2676 13947 2700
rect 13285 2012 13291 2064
rect 13343 2012 13350 2064
rect 13297 1727 13339 2012
rect 14919 1716 14961 3096
rect 18599 3018 18605 3086
rect 18657 3018 18663 3086
rect 19695 2961 19701 3013
rect 19753 2961 19759 3013
rect 21245 2961 21251 3013
rect 21303 2961 21309 3013
rect 22486 2961 22493 3013
rect 22545 2961 22551 3013
rect 23380 2961 23386 3013
rect 23438 2961 23444 3013
rect 18429 2902 18435 2954
rect 18487 2902 18494 2954
rect 15309 2824 15316 2876
rect 15368 2824 15374 2876
rect 16296 2825 16302 2877
rect 16354 2825 16360 2877
rect 15322 1724 15364 2824
rect 17701 2756 17708 2808
rect 17760 2756 17766 2808
rect 18685 2756 18691 2808
rect 18743 2756 18750 2808
rect 16049 2614 16083 2662
rect 16033 2562 16039 2614
rect 16091 2562 16097 2614
rect 16449 2613 16483 2660
rect 16434 2561 16440 2613
rect 16492 2561 16498 2613
rect 17301 2496 17307 2548
rect 17359 2496 17366 2548
rect 15679 2081 15685 2133
rect 15737 2081 15744 2133
rect 15689 1727 15731 2081
rect 15880 1663 15886 1715
rect 15938 1663 15945 1715
rect 13488 1594 13494 1646
rect 13546 1594 13553 1646
rect 17313 1522 17355 2496
rect 17715 1703 17757 2756
rect 18701 2733 18735 2756
rect 18869 2481 18903 2661
rect 18857 2429 18863 2481
rect 18915 2429 18922 2481
rect 18070 2151 18076 2203
rect 18128 2151 18135 2203
rect 18081 1728 18123 2151
rect 18273 1733 18279 1785
rect 18331 1733 18338 1785
rect 19705 1704 19747 2961
rect 20092 2892 20099 2944
rect 20151 2892 20157 2944
rect 21076 2892 21082 2944
rect 21134 2892 21140 2944
rect 20106 1704 20148 2892
rect 21092 2891 21120 2892
rect 22083 2429 22089 2481
rect 22141 2429 22147 2481
rect 20462 2219 20468 2271
rect 20520 2219 20527 2271
rect 20473 1728 20515 2219
rect 20666 1802 20672 1854
rect 20724 1802 20731 1854
rect 20677 1730 20719 1802
rect 22094 1464 22136 2429
rect 22499 1722 22541 2961
rect 23239 2549 23273 2657
rect 24475 2564 24482 2616
rect 24534 2564 24540 2616
rect 23224 2497 23230 2549
rect 23282 2497 23288 2549
rect 22853 2290 22859 2342
rect 22911 2290 22918 2342
rect 22865 1731 22907 2290
rect 23055 1872 23061 1924
rect 23113 1872 23120 1924
rect 23068 1730 23110 1872
rect 24489 1726 24531 2564
rect 24892 1721 24934 3103
rect 25247 2361 25253 2413
rect 25305 2361 25312 2413
rect 25257 1729 25299 2361
rect 11910 967 11916 1019
rect 11968 967 11974 1019
rect 8876 -1908 8918 -1331
rect 10621 -1908 10663 -652
rect 11268 -1908 11310 -1331
rect 13013 -1908 13055 -651
rect 13659 -1908 13701 -1331
rect 15404 -1908 15446 -651
rect 16052 -1908 16094 -1331
rect 17797 -1908 17839 -650
rect 18444 -1908 18486 -1331
rect 20188 -1908 20230 -651
rect 20835 -1908 20877 -1330
rect 22581 -1908 22623 -652
rect 23228 -1908 23270 -1331
rect 24974 -1908 25016 -650
<< metal4 >>
rect 9023 12571 10729 13159
rect 10055 2874 10580 7673
rect 12824 7444 13488 7540
rect 12826 7376 13488 7444
rect 12826 7292 13822 7376
rect 24043 7336 27157 7437
rect 24043 7330 24460 7336
rect 12826 7212 13488 7292
rect 13654 7212 13822 7292
rect 12826 3212 13822 7212
rect 8122 2660 10580 2874
rect 8122 2503 10581 2660
rect 8122 -1451 8351 2503
rect 10751 2451 13822 3212
rect 23794 4382 25158 4546
rect 23794 3834 24814 4382
rect 25024 3834 25158 4382
rect 23794 3643 25158 3834
rect 23794 3431 24798 3643
rect 25030 3431 25158 3643
rect 23794 3120 25158 3431
rect 25369 2465 25451 2471
rect 25338 2459 25451 2465
rect 10751 1359 13823 2451
rect 24345 2367 25451 2459
rect 24345 2207 24914 2367
rect 25004 2207 25451 2367
rect 24345 2044 25451 2207
rect 24342 1532 25452 2044
rect 24346 1446 25452 1532
rect 24346 1138 24410 1446
rect 24500 1138 25452 1446
rect 24346 902 25452 1138
rect 8122 -1771 9605 -1451
use hgu_clk_async  x1
timestamp 1699633333
transform 1 0 9186 0 -1 9828
box -7122 -3534 2561 2470
use hgu_clk_sample  x2
timestamp 1699539229
transform 1 0 9205 0 1 5836
box 1440 1522 17950 7913
use hgu_sarlogic_8bit_logic  x3
timestamp 1699717961
transform 1 0 10463 0 1 906
box 290 1745 13444 6250
use hgu_sarlogic_sw_ctrl  x4
timestamp 1699632744
transform 1 0 8575 0 1 -1565
box -144 -343 16876 3300
use hgu_sarlogic_retimer  x5
timestamp 1699720582
transform 1 0 12207 0 1 -3283
box 11730 5040 19043 10661
<< labels >>
flabel metal1 10933 3942 10967 3977 0 FreeSans 320 0 0 0 comp_result
port 55 nsew
flabel metal2 10001 2976 10029 6744 0 FreeSans 320 0 0 0 sar_clk
port 8 nsew
flabel metal2 11750 7806 11802 7855 0 FreeSans 320 0 0 0 sample_clk_b
port 7 nsew
flabel metal1 11827 8983 11873 9018 0 FreeSans 320 0 0 0 sample_clk
port 6 nsew
flabel metal1 10869 12169 10912 12233 0 FreeSans 320 0 0 0 ext_clk
port 4 nsew
flabel metal1 2330 11810 2393 11857 0 FreeSans 320 0 0 0 ready
port 1 nsew
flabel metal4 12826 2361 13488 7539 0 FreeSans 1600 0 0 0 VDD
port 10 nsew
flabel metal4 10055 2503 10580 7673 0 FreeSans 1600 0 0 0 VSS
port 9 nsew
flabel metal1 10922 6824 10956 6858 0 FreeSans 320 0 0 0 sel_bit[0]
port 11 nsew
flabel metal1 10927 6687 10962 6722 0 FreeSans 320 0 0 0 sel_bit[1]
port 12 nsew
flabel metal1 30455 3815 30764 3863 0 FreeSans 320 0 0 0 sar_result[0]
port 20 nsew
flabel metal1 30445 4145 30754 4193 0 FreeSans 320 0 0 0 sar_result[1]
port 13 nsew
flabel metal1 30447 3516 30756 3564 0 FreeSans 320 0 0 0 sar_result[2]
port 14 nsew
flabel metal1 30461 3174 30770 3222 0 FreeSans 320 0 0 0 sar_result[3]
port 15 nsew
flabel metal1 30450 2864 30759 2912 0 FreeSans 320 0 0 0 sar_result[5]
port 16 nsew
flabel metal1 30456 2533 30765 2581 0 FreeSans 320 0 0 0 sar_result[4]
port 17 nsew
flabel metal1 30453 2237 30762 2285 0 FreeSans 320 0 0 0 sar_result[6]
port 18 nsew
flabel metal1 30451 1893 30760 1941 0 FreeSans 320 0 0 0 sar_result[7]
port 19 nsew
flabel metal1 13479 10913 13504 10941 0 FreeSans 320 0 0 0 sample_delay_cap_ctrl_code[2]
port 21 nsew
flabel metal1 13481 10857 13506 10885 0 FreeSans 320 0 0 0 sample_delay_cap_ctrl_code[1]
port 22 nsew
flabel metal1 13483 10801 13508 10829 0 FreeSans 320 0 0 0 sample_delay_cap_ctrl_code[0]
port 23 nsew
flabel metal1 13484 10745 13509 10773 0 FreeSans 320 0 0 0 sample_delay_cap_ctrl_code[6]
port 24 nsew
flabel metal1 13486 10689 13511 10717 0 FreeSans 320 0 0 0 sample_delay_cap_ctrl_code[5]
port 25 nsew
flabel metal1 13485 10633 13510 10661 0 FreeSans 320 0 0 0 sample_delay_cap_ctrl_code[4]
port 26 nsew
flabel metal1 13473 10493 13505 10605 0 FreeSans 320 0 0 0 sample_delay_offset
port 35 nsew
flabel metal1 13198 12668 13224 12702 0 FreeSans 320 0 0 0 sample_delay_cap_ctrl_code[3]
port 36 nsew
flabel metal1 19914 12668 19940 12702 0 FreeSans 320 0 0 0 sample_delay_cap_ctrl_code[7]
port 37 nsew
flabel metal1 26659 8407 26685 8441 0 FreeSans 320 0 0 0 sample_delay_cap_ctrl_code[11]
port 38 nsew
flabel metal1 19956 8407 19982 8441 0 FreeSans 320 0 0 0 sample_delay_cap_ctrl_code[15]
port 39 nsew
flabel metal1 2930 10449 4871 10477 0 FreeSans 320 0 0 0 async_setb_delay_cap_ctrl_code[2]
port 40 nsew
flabel metal1 2931 10393 7297 10421 0 FreeSans 320 0 0 0 async_setb_delay_cap_ctrl_code[1]
port 41 nsew
flabel metal1 2929 10337 8154 10365 0 FreeSans 320 0 0 0 async_setb_delay_cap_ctrl_code[0]
port 42 nsew
flabel metal1 2928 10281 8154 10309 0 FreeSans 320 0 0 0 async_resetb_delay_cap_ctrl_code[0]
port 43 nsew
flabel metal1 2932 10225 7297 10253 0 FreeSans 320 0 0 0 async_resetb_delay_cap_ctrl_code[1]
port 44 nsew
flabel metal1 2930 10169 4871 10197 0 FreeSans 320 0 0 0 async_resetb_delay_cap_ctrl_code[2]
port 45 nsew
flabel metal1 2324 12193 2356 12227 0 FreeSans 320 0 0 0 async_setb_delay_cap_ctrl_code[3]
port 46 nsew
flabel metal1 2324 8419 2366 8453 0 FreeSans 320 0 0 0 async_resetb_delay_cap_ctrl_code[3]
port 47 nsew
flabel metal2 2737 9041 2790 11605 0 FreeSans 320 0 0 0 async_delay_offset
port 48 nsew
flabel metal1 23937 6371 24075 6405 0 FreeSans 320 0 0 0 retimer_delay_code[3]
port 50 nsew
flabel metal1 25545 4635 26484 4663 0 FreeSans 320 0 0 0 retimer_delay_code[2]
port 51 nsew
flabel metal1 25545 4579 28910 4607 0 FreeSans 320 0 0 0 retimer_delay_code[1]
port 52 nsew
flabel metal1 25545 4523 29767 4551 0 FreeSans 320 0 0 0 retimer_delay_code[0]
port 54 nsew
flabel metal2 8716 -1261 8758 2925 0 FreeSans 320 0 0 0 vss_sw[7]
port 56 nsew
flabel metal2 8798 1577 8840 2925 0 FreeSans 320 0 0 0 vss_sw[6]
port 57 nsew
flabel metal2 8882 1647 8924 2925 0 FreeSans 320 0 0 0 vss_sw[5]
port 58 nsew
flabel metal2 8970 1716 9012 2925 0 FreeSans 320 0 0 0 vss_sw[4]
port 59 nsew
flabel metal2 9057 1786 9099 2925 0 FreeSans 320 0 0 0 vss_sw[3]
port 60 nsew
flabel metal2 9143 1855 9185 2925 0 FreeSans 320 0 0 0 vss_sw[2]
port 61 nsew
flabel metal2 9229 1925 9271 2925 0 FreeSans 320 0 0 0 vss_sw[1]
port 62 nsew
flabel metal2 9316 1995 9358 2925 0 FreeSans 320 0 0 0 vdd_sw[7]
port 63 nsew
flabel metal2 9402 2065 9444 2925 0 FreeSans 320 0 0 0 vdd_sw[6]
port 64 nsew
flabel metal2 9488 2134 9530 2925 0 FreeSans 320 0 0 0 vdd_sw[5]
port 65 nsew
flabel metal2 9575 2204 9617 2925 0 FreeSans 320 0 0 0 vdd_sw[4]
port 66 nsew
flabel metal2 9660 2274 9702 2925 0 FreeSans 320 0 0 0 vdd_sw[3]
port 67 nsew
flabel metal2 9747 2343 9789 2925 0 FreeSans 320 0 0 0 vdd_sw[2]
port 68 nsew
flabel metal2 9834 2412 9876 2925 0 FreeSans 320 0 0 0 vdd_sw[1]
port 69 nsew
flabel metal2 8876 -1908 8918 -1331 0 FreeSans 320 0 0 0 vss_sw_b[7]
port 70 nsew
flabel metal2 11268 -1908 11310 -1331 0 FreeSans 320 0 0 0 vss_sw_b[6]
port 71 nsew
flabel metal2 13659 -1908 13701 -1331 0 FreeSans 320 0 0 0 vss_sw_b[5]
port 72 nsew
flabel metal2 16052 -1908 16094 -1331 0 FreeSans 320 0 0 0 vss_sw_b[4]
port 73 nsew
flabel metal2 18444 -1908 18486 -1331 0 FreeSans 320 0 0 0 vss_sw_b[3]
port 74 nsew
flabel metal2 20835 -1908 20877 -1330 0 FreeSans 320 0 0 0 vss_sw_b[2]
port 75 nsew
flabel metal2 23228 -1908 23270 -1331 0 FreeSans 320 0 0 0 vss_sw_b[1]
port 76 nsew
flabel metal2 24974 -1908 25016 -650 0 FreeSans 320 0 0 0 vdd_sw_b[1]
port 77 nsew
flabel metal2 22581 -1908 22623 -652 0 FreeSans 320 0 0 0 vdd_sw_b[2]
port 78 nsew
flabel metal2 20188 -1908 20230 -651 0 FreeSans 320 0 0 0 vdd_sw_b[3]
port 79 nsew
flabel metal2 17797 -1908 17839 -650 0 FreeSans 320 0 0 0 vdd_sw_b[4]
port 80 nsew
flabel metal2 15404 -1908 15446 -651 0 FreeSans 320 0 0 0 vdd_sw_b[5]
port 81 nsew
flabel metal2 13013 -1908 13055 -651 0 FreeSans 320 0 0 0 vdd_sw_b[6]
port 82 nsew
flabel metal2 10621 -1908 10663 -652 0 FreeSans 320 0 0 0 vdd_sw_b[7]
port 83 nsew
flabel metal1 13484 10382 13510 10408 0 FreeSans 320 0 0 0 sample_delay_cap_ctrl_code[9]
port 88 nsew
flabel metal1 13486 10326 13512 10352 0 FreeSans 320 0 0 0 sample_delay_cap_ctrl_code[8]
port 89 nsew
flabel metal1 13482 10270 13508 10296 0 FreeSans 320 0 0 0 sample_delay_cap_ctrl_code[14]
port 90 nsew
flabel metal1 13486 10214 13512 10240 0 FreeSans 320 0 0 0 sample_delay_cap_ctrl_code[13]
port 91 nsew
flabel metal1 13484 10158 13510 10184 0 FreeSans 320 0 0 0 sample_delay_cap_ctrl_code[12]
port 92 nsew
flabel metal1 13482 10438 13506 10464 0 FreeSans 320 0 0 0 sample_delay_cap_ctrl_code[10]
port 93 nsew
flabel metal1 24237 5786 24349 5834 0 FreeSans 320 0 0 0 retimer_eob_delay_offset
port 49 nsew
<< end >>
