* NGSPICE file created from hgu_top_block_flat.ext - technology: sky130A

.subckt hgu_top_block_flat sel_bit[0] sel_bit[1] EXT_CLK sample_delay_cap_ctrl_code[11]
+ sample_delay_cap_ctrl_code[3] sample_delay_cap_ctrl_code[2] sample_delay_cap_ctrl_code[1]
+ sample_delay_cap_ctrl_code[0] sample_delay_cap_ctrl_code[6] sample_delay_cap_ctrl_code[5]
+ sample_delay_cap_ctrl_code[4] sample_delay_cap_ctrl_code[10] sample_delay_cap_ctrl_code[9]
+ sample_delay_cap_ctrl_code[8] sample_delay_cap_ctrl_code[14] sample_delay_cap_ctrl_code[13]
+ sample_delay_offset async_resetb_delay_cap_ctrl_code[2] async_resetb_delay_cap_ctrl_code[1]
+ async_setb_delay_cap_ctrl_code[1] async_setb_delay_cap_ctrl_code[2] async_setb_delay_cap_ctrl_code[3]
+ retimer_delay_code[2] retimer_delay_code[1] retimer_delay_offset async_delay_offset
+ vip vin result[2] result[5] async_resetb_delay_cap_ctrl_code[0] result[0] async_resetb_delay_cap_ctrl_code[3]
+ result[1] retimer_delay_code[0] result[3] result[4] retimer_delay_code[3] result[6]
+ sample_delay_cap_ctrl_code[12] result[7] async_setb_delay_cap_ctrl_code[0] sample_delay_cap_ctrl_code[15]
+ sample_delay_cap_ctrl_code[7] VDD VSS
X0 a_n982_1868# hgu_sarlogic_flat_0.x4.x5.D VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X1 hgu_cdac_half_1.VREF hgu_cdac_half_1.d<5> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2 hgu_sarlogic_flat_0.x2.x2.x3.x5[7].floating hgu_sarlogic_flat_0.x2.x2.x3.x10.Y hgu_sarlogic_flat_0.x2.x2.x3.x9.output_stack VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X3 VSS a_n607_7947# hgu_cdac_sw_buffer_2.x7.X VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X4 VSS a_12012_2136# a_12733_1868# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X5 hgu_sarlogic_flat_0.x4.x19.Q_N a_2444_2136# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X6 hgu_cdac_half_1.VREF hgu_cdac_half_1.d<6> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X7 VSS hgu_cdac_half_1.db<3> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<7:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X8 VDD a_2036_7824# hgu_sarlogic_flat_0.x3.x4.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9 a_10681_7824# a_9763_7798# a_10235_8008# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X10 a_7071_6052# a_7369_6352# a_7305_6444# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0924 ps=0.86 w=0.42 l=0.15
X11 VDD a_12069_8487# a_12790_8795# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X12 VDD a_n871_7253# hgu_cdac_half_1.d<3> VDD sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X13 a_12494_6078# a_12626_6262# a_12358_6052# VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0864 ps=0.91 w=0.64 l=0.15
X14 VSS a_1196_n1740# hgu_cdac_half_0.d<6> VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X15 a_2975_1179# a_2058_1153# a_2530_1363# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0675 ps=0.735 w=0.36 l=0.15
X16 hgu_cdac_half_1.VREF hgu_cdac_half_1.d<6> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X17 hgu_cdac_half_1.VREF hgu_cdac_half_1.db<6> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X18 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<15:0> hgu_cdac_half_1.d<4> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X19 a_n7766_6446# a_n7390_7871# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.139 pd=1.17 as=0.139 ps=1.17 w=0.84 l=0.15
X20 VSS a_n148_n1104# hgu_cdac_half_0.db<4> VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X21 hgu_cdac_half_1.d<6> a_n2219_8368# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X22 a_7371_7798# hgu_sarlogic_flat_0.x3.x5.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X23 a_n6887_13761# hgu_comp_flat_0.ready a_n6959_13899# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X24 a_9523_8513# a_9677_8487# a_9383_8487# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X25 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<7:0> hgu_cdac_half_1.d<3> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X26 VDD hgu_comp_flat_0.RS_p a_n7216_6420# VDD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0.244 ps=2.26 w=0.84 l=0.15
X27 hgu_cdac_sw_buffer_0.VDD a_n1158_n1744# hgu_cdac_half_0.db<6> hgu_cdac_sw_buffer_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X28 a_1993_1179# a_1203_1153# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0703 ps=0.755 w=0.42 l=0.15
X29 VSS a_10164_8487# a_10099_8513# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X30 hgu_sarlogic_flat_0.x4.x25.Q_N a_7228_2136# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X31 VSS a_8909_7798# hgu_sarlogic_flat_0.x3.x42.Q_N VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X32 a_4532_6951# a_4143_6951# a_4424_7317# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X33 hgu_cdac_half_0.VREF hgu_cdac_half_0.d<2> hgu_cdac_half_0.hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.35
X34 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.db<6> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X35 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X36 a_18224_5950# a_18058_5950# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X37 a_14490_1363# a_14018_1153# a_14734_1545# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X38 hgu_cdac_sw_buffer_3.x11.X a_n4397_8367# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X39 VSS hgu_comp_flat_0.clk a_n7660_7467# VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X40 hgu_cdac_half_1.d<0> a_15125_1868# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X41 hgu_vgen_vref_0.vcm hgu_vgen_vref_0.phi1 hgu_vgen_vref_0.mimtop2 VSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=0.5
X42 hgu_sarlogic_flat_0.x4.x2.X a_n424_3698# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X43 a_18224_6596# a_18058_6596# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X44 a_12291_6444# a_12154_6052# a_11855_6052# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X45 hgu_cdac_sw_buffer_0.VDD hgu_cdac_sw_buffer_0.x11.A a_n1158_n1744# hgu_cdac_sw_buffer_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X46 hgu_cdac_half_1.d<6> a_n2219_8368# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X47 VSS hgu_sarlogic_flat_0.x4.D[5] a_5367_1179# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X48 a_11856_7798# a_12155_7798# a_12090_7824# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.066 ps=0.745 w=0.36 l=0.15
X49 a_8798_1179# a_8925_1347# a_8379_1153# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.03 as=0.0864 ps=0.91 w=0.64 l=0.15
X50 VDD a_8281_2708# hgu_sarlogic_flat_0.x4.x14.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X51 VSS hgu_cdac_half_1.d<6> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X52 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X53 a_4976_1868# a_4362_1842# a_4836_2136# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X54 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<15:0> hgu_cdac_half_1.d<4> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X55 hgu_cdac_half_1.VREF hgu_cdac_half_1.d<6> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X56 a_n4397_8367# hgu_cdac_sw_buffer_3.x11.A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X57 hgu_cdac_half_0.d<6> a_1196_n1740# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X58 VDD VDD a_16581_5924# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X59 VSS VDD a_9146_1842# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X60 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_1.d<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X61 a_10279_6951# hgu_sarlogic_flat_0.x3.x42.Q_N VSS VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X62 a_14654_8353# hgu_sarlogic_flat_0.x5.eob a_14566_8353# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X63 VSS a_1454_6950# hgu_sarlogic_flat_0.x3.x7.X VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X64 VSS hgu_cdac_half_0.db<5> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X65 a_4141_1347# a_4450_1153# a_4385_1179# VSS sky130_fd_pr__nfet_01v8 ad=0.0486 pd=0.63 as=0.066 ps=0.745 w=0.36 l=0.15
X66 hgu_sarlogic_flat_0.x5.x2.x10.Y retimer_delay_code[3] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X67 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X68 hgu_cdac_half_0.VREF hgu_cdac_half_0.d<6> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X69 VSS hgu_cdac_half_0.db<6> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X70 a_611_11594# a_n134_11726# a_747_11682# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X71 hgu_vgen_vref_0.mimtop1 hgu_vgen_vref_0.mimbot1 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X72 hgu_cdac_half_0.VREF hgu_cdac_half_0.d<4> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<15:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X73 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_0.d<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X74 a_6829_6078# hgu_sarlogic_flat_0.x3.x4.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.154 ps=1.34 w=0.64 l=0.15
X75 hgu_sarlogic_flat_0.x4.x13.X a_7570_2883# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.113 ps=1.04 w=0.65 l=0.15
X76 a_17068_6564# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X77 VDD a_9620_2136# a_9545_2234# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0956 pd=0.875 as=0.0787 ps=0.795 w=0.42 l=0.15
X78 VSS hgu_sarlogic_flat_0.x2.x3.Y a_2323_11578# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X79 a_3314_11664# hgu_sarlogic_flat_0.x2.x7.A VDD VSS sky130_fd_pr__nfet_01v8 ad=0.0651 pd=0.73 as=0.0693 ps=0.75 w=0.42 l=0.15
X80 a_555_10641# hgu_sarlogic_flat_0.x1.x3.X a_192_10793# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X81 VDD hgu_cdac_sw_buffer_3.x9.X a_n4479_7727# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X82 a_5891_1331# a_5987_1153# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X83 a_12152_1868# hgu_sarlogic_flat_0.x4.x2.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.03 as=0.0703 ps=0.755 w=0.42 l=0.15
X84 VDD a_18973_5924# a_19694_6232# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X85 VSS VSS a_1390_n460# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X86 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<15:0> hgu_cdac_half_0.db<4> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X87 hgu_comp_flat_0.RS_n a_n6526_6819# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.15
X88 a_18224_4670# a_18058_4670# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X89 a_20464_8538# hgu_sarlogic_flat_0.x5.x2.x9.output_stack hgu_sarlogic_flat_0.x5.x3.A VSS sky130_fd_pr__nfet_01v8 ad=0.0651 pd=0.73 as=0.122 ps=1.42 w=0.42 l=0.15
X90 VSS hgu_sarlogic_flat_0.x3.x4.A a_2036_7824# VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X91 hgu_cdac_half_0.VREF hgu_cdac_half_0.db<3> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<7:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X92 VDD a_3960_3698# hgu_sarlogic_flat_0.x4.x9.A1 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X93 hgu_sarlogic_flat_0.x4.x9.A1 a_3960_3698# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X94 vin hgu_tah_0.sw hgu_tah_0.tah_vn VSS sky130_fd_pr__nfet_01v8 ad=0.454 pd=3.08 as=0.853 ps=6.12 w=2.75 l=0.15
X95 VSS hgu_sarlogic_flat_0.x4.x14.X a_8232_1868# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X96 VDD VDD a_4362_1842# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.17 ps=1.81 w=0.64 l=0.15
X97 VDD sample_delay_offset hgu_sarlogic_flat_0.x2.x2.x4.x6.SW VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X98 VSS a_4979_7798# a_4978_8098# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X99 a_2725_6078# a_2585_6352# a_2287_6052# VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.0711 ps=0.755 w=0.36 l=0.15
X100 hgu_vgen_vref_0.mimtop2 VSS sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X101 a_5205_6951# a_4143_6951# a_5110_6951# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X102 a_12342_1179# a_11830_1153# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0882 ps=0.84 w=0.42 l=0.15
X103 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.d<6> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X104 a_n2219_8368# hgu_cdac_sw_buffer_2.x11.A VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X105 VSS VDD a_n770_1179# VSS sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.109 ps=1.03 w=0.42 l=0.15
X106 VSS hgu_cdac_half_0.db<6> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X107 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X108 hgu_vgen_vref_0.phi1 a_n55304_8227# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X109 VSS hgu_cdac_half_0.d<4> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<15:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X110 a_9574_1179# a_9706_1363# a_9438_1153# VSS sky130_fd_pr__nfet_01v8 ad=0.0974 pd=0.97 as=0.0864 ps=0.91 w=0.64 l=0.15
X111 a_14674_2883# a_14492_2883# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X112 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_1.db<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X113 VSS hgu_cdac_half_0.db<6> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X114 hgu_cdac_half_1.VREF hgu_cdac_half_1.d<6> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X115 VSS hgu_cdac_half_1.db<2> hgu_cdac_half_1.hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT VSS sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.35
X116 hgu_tah_0.tah_vn hgu_tah_0.sw hgu_tah_0.tah_vn hgu_tah_0.VDD sky130_fd_pr__pfet_01v8 ad=8.85 pd=58.2 as=0.908 ps=5.83 w=5.5 l=0.15
X117 a_7228_2136# hgu_sarlogic_flat_0.x4.x2.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.132 pd=1.22 as=0.0956 ps=0.875 w=0.42 l=0.15
X118 hgu_cdac_half_1.VREF hgu_cdac_half_1.db<5> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X119 hgu_cdac_sw_buffer_3.x11.X a_n4397_8367# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X120 hgu_cdac_half_1.VREF hgu_cdac_half_1.db<6> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X121 VSS a_n3387_7727# hgu_cdac_half_1.db<4> VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X122 a_n7760_6349# a_n6526_6819# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0759 pd=0.79 as=0.143 ps=1.54 w=0.46 l=0.15
X123 VSS hgu_cdac_half_0.d<5> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X124 a_6252_2556# VSS a_5889_2708# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X125 VSS a_2268_n241# hgu_cdac_sw_buffer_1.x4.X VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X126 hgu_sarlogic_flat_0.x2.x3.A a_3080_14774# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X127 VDD a_11774_6925# a_11684_7317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X128 VDD hgu_sarlogic_flat_0.x2.x2.x1.IN a_10575_16177# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X129 hgu_sarlogic_flat_0.x1.x2.x4[3].floating async_setb_delay_cap_ctrl_code[2] hgu_sarlogic_flat_0.x1.x2.x9.output_stack VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X130 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.d<6> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X131 a_7131_8513# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X132 hgu_vgen_vref_0.phi2_n a_n54752_6595# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X133 VSS hgu_cdac_half_0.db<5> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X134 a_13182_1868# a_13016_1868# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X135 a_13494_2530# hgu_sarlogic_flat_0.x4.x20.S VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X136 a_n134_11726# hgu_sarlogic_flat_0.x1.x10.Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.154 ps=1.34 w=0.64 l=0.15
X137 hgu_sarlogic_flat_0.x2.x7.A hgu_sarlogic_flat_0.x2.x2.x3.x9.output_stack a_3314_11461# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.0651 ps=0.73 w=0.42 l=0.15
X138 a_14654_7525# hgu_sarlogic_flat_0.x5.eob a_14566_7525# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X139 a_n472_2150# a_n890_2234# a_n716_1842# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X140 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.db<6> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X141 hgu_cdac_half_0.db<5> a_n688_n1104# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X142 VDD hgu_sarlogic_flat_0.x4.x9.S a_3000_2883# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.0767 ps=0.785 w=0.42 l=0.15
X143 hgu_cdac_half_1.hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT hgu_cdac_half_1.d<2> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X144 a_2057_1453# hgu_sarlogic_flat_0.x4.x9.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X145 hgu_sarlogic_flat_0.x3.D[0] a_8478_6951# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X146 VSS a_5182_6052# a_5117_6078# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0935 ps=0.965 w=0.64 l=0.15
X147 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_0.db<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X148 VDD a_11775_8487# a_11685_8879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X149 a_n3049_7252# hgu_cdac_sw_buffer_3.x6.A VSS VSS sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X150 a_13494_2530# hgu_sarlogic_flat_0.x4.x20.S VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X151 VSS a_11300_6052# hgu_sarlogic_flat_0.x3.x63.Q_N VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X152 a_9371_1545# a_9234_1153# a_8925_1347# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X153 hgu_cdac_half_1.d<1> a_12733_1868# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X154 hgu_sarlogic_flat_0.x1.x2.x2.floating async_setb_delay_cap_ctrl_code[0] hgu_sarlogic_flat_0.x1.x2.x9.output_stack VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.124 ps=1.43 w=0.42 l=0.15
X155 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X156 hgu_sarlogic_flat_0.x2.x2.x2.x9.output_stack hgu_sarlogic_flat_0.x2.x2.x2.x10.Y hgu_sarlogic_flat_0.x2.x2.x2.x5[7].floating VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X157 a_7306_8190# a_6517_7798# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0819 ps=0.81 w=0.42 l=0.15
X158 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.db<6> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.35
X159 VSS hgu_sarlogic_flat_0.x4.x9.S a_3007_2556# VSS sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.0693 ps=0.75 w=0.42 l=0.15
X160 VDD hgu_sarlogic_flat_0.x4.x14.X a_8232_1868# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X161 hgu_tah_0.VDD a_n54567_7371# a_n54754_7113# hgu_tah_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X162 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X163 a_13709_1347# a_14018_1153# a_13953_1179# VSS sky130_fd_pr__nfet_01v8 ad=0.0486 pd=0.63 as=0.066 ps=0.745 w=0.36 l=0.15
X164 VDD a_5889_2708# hgu_sarlogic_flat_0.x4.x12.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X165 a_2786_2883# VSS a_2786_2556# VSS sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X166 VDD a_4979_7798# a_4978_8098# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X167 a_n7660_7467# hgu_tah_0.tah_vn hgu_comp_flat_0.Q VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X168 hgu_sarlogic_flat_0.x5.x1[3].Q_N a_19460_5924# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X169 hgu_sarlogic_flat_0.x4.x2.X a_n424_3698# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X170 a_7508_8190# a_7371_7798# a_7072_7798# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X171 a_2584_1868# a_1970_1842# a_2444_2136# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X172 VSS hgu_cdac_half_0.d<6> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X173 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<7:0> hgu_cdac_half_1.d<3> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X174 hgu_tah_0.VDD hgu_vgen_vref_0.clk hgu_vgen_vref_0.sky130_fd_sc_hd__nand2_1_0.Y hgu_tah_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X175 a_16287_4644# a_16113_5036# a_16427_4670# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X176 VDD a_n6292_6446# hgu_comp_flat_0.comp_outn VDD sky130_fd_pr__pfet_01v8 ad=0.139 pd=1.17 as=0.139 ps=1.17 w=0.84 l=0.15
X177 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_0.d<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X178 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.d<6> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X179 hgu_cdac_half_1.VREF hgu_cdac_half_1.d<4> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<15:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X180 hgu_cdac_half_0.VREF hgu_cdac_half_0.db<2> hgu_cdac_half_0.hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X181 a_7176_1868# a_6006_1868# a_7069_2234# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0486 ps=0.63 w=0.36 l=0.15
X182 a_6421_6052# a_6516_6052# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X183 VSS a_2036_7824# hgu_sarlogic_flat_0.x3.x4.X VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X184 a_7575_7798# a_7843_8008# a_7789_8106# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X185 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X186 VDD a_n2219_8368# hgu_cdac_half_1.d<6> VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X187 VDD a_7772_8487# a_8479_8513# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X188 a_7888_8513# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X189 a_9222_7824# hgu_sarlogic_flat_0.x3.x4.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X190 a_n3877_7252# hgu_cdac_sw_buffer_3.x3.A VSS VSS sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X191 VSS hgu_tah_0.sw_n a_n1334_3698# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X192 hgu_cdac_half_0.d<6> a_1196_n1740# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X193 VSS hgu_cdac_half_0.db<6> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X194 VSS async_delay_offset hgu_sarlogic_flat_0.x1.x4.x6.SW VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X195 a_13966_1545# a_13163_1153# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0787 pd=0.795 as=0.0956 ps=0.875 w=0.42 l=0.15
X196 a_4001_13960# hgu_sarlogic_flat_0.x2.x3.A a_3929_14098# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X197 hgu_sarlogic_flat_0.x2.x2.x3.x5[7].floating hgu_sarlogic_flat_0.x2.x2.x3.x10.Y hgu_sarlogic_flat_0.x2.x2.x3.x9.output_stack VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X198 VDD a_n4397_8367# hgu_cdac_sw_buffer_3.x11.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X199 VDD a_17068_4644# a_17775_4670# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X200 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.db<6> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X201 a_13182_1868# a_13016_1868# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X202 a_n806_2234# a_n1170_1868# a_n890_2234# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X203 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_1.d<5> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X204 hgu_sarlogic_flat_0.x4.x9.A1 a_3960_3698# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X205 a_6194_1868# hgu_sarlogic_flat_0.x4.D[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X206 a_5291_7317# a_4143_6951# a_5205_6951# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X207 VDD a_17068_6564# a_17775_6606# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X208 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_0.d<5> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X209 hgu_cdac_half_1.VREF hgu_cdac_half_1.db<5> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X210 VSS a_4030_7798# hgu_sarlogic_flat_0.x3.x48.Q VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X211 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X212 a_n28_11682# a_108_11334# a_n447_11350# VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0864 ps=0.91 w=0.64 l=0.15
X213 a_12352_2883# hgu_sarlogic_flat_0.x4.x9.A1 a_12280_2883# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X214 VDD a_17068_6564# a_16980_6590# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X215 VDD a_16581_5510# a_17302_5310# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X216 VDD a_19460_5284# a_19372_5310# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X217 VDD a_n424_3698# hgu_sarlogic_flat_0.x4.x2.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X218 a_3378_9360# sel_bit[0] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X219 a_12490_6951# a_11153_6951# a_12381_6951# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X220 VSS a_1196_n1740# hgu_cdac_half_0.d<6> VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X221 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X222 a_11507_6951# hgu_sarlogic_flat_0.x3.x7.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X223 VSS hgu_sarlogic_flat_0.x4.x12.X a_5840_1868# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X224 a_5292_8879# a_4144_8513# a_5206_8513# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X225 hgu_sarlogic_flat_0.x5.x2.x9.output_stack hgu_sarlogic_flat_0.x5.x2.x10.Y hgu_sarlogic_flat_0.x5.x2.x5[7].floating VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X226 VDD a_19460_5924# a_19372_6316# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X227 VDD VDD a_1970_1842# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.17 ps=1.81 w=0.64 l=0.15
X228 VDD hgu_cdac_sw_buffer_2.x3.X a_n1749_7728# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X229 VSS a_1422_7824# hgu_sarlogic_flat_0.x3.x4.A VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X230 VSS hgu_sarlogic_flat_0.x3.x7.X a_3504_6078# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X231 VDD a_4654_1153# a_4587_1545# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X232 a_12352_2556# a_12098_2883# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.145 ps=1.11 w=0.42 l=0.15
X233 VDD a_18679_5284# a_18589_5310# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X234 hgu_cdac_half_0.VREF hgu_cdac_half_0.db<5> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X235 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X236 a_n53014_7459# hgu_vgen_vref_0.sky130_fd_sc_hd__inv_1_2.Y hgu_vgen_vref_0.sky130_fd_sc_hd__nand2_1_1.Y VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X237 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X238 a_9404_12677# hgu_sarlogic_flat_0.x2.x2.x3.IN a_9332_12677# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X239 hgu_cdac_sw_buffer_2.x8.X a_n2025_7088# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X240 VDD a_18679_5924# a_18589_6316# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X241 VSS hgu_cdac_half_0.db<6> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X242 VSS a_n447_11350# hgu_sarlogic_flat_0.x1.x27.Q_N VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X243 a_n1190_n245# hgu_cdac_sw_buffer_0.x9.A VSS VSS sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X244 hgu_cdac_half_0.db<4> a_n148_n1104# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X245 a_8762_2234# a_8398_1868# a_8678_2234# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X246 hgu_cdac_half_1.VREF hgu_cdac_half_1.d<6> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X247 VSS hgu_cdac_half_1.db<4> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<15:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X248 a_4836_2136# hgu_sarlogic_flat_0.x4.x2.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.132 pd=1.22 as=0.0956 ps=0.875 w=0.42 l=0.15
X249 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<15:0> hgu_cdac_half_1.d<4> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X250 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_1.d<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X251 a_7069_2234# a_6006_1868# a_6925_2150# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X252 VDD a_n3927_7727# hgu_cdac_half_1.db<5> VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X253 hgu_cdac_sw_buffer_2.x12.X a_n1473_7088# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X254 VDD a_2036_7824# hgu_sarlogic_flat_0.x3.x4.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X255 a_6535_6951# a_6369_6951# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X256 a_3860_2556# VSS a_3497_2708# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X257 a_2926_6078# a_3058_6262# a_2790_6052# VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0864 ps=0.91 w=0.64 l=0.15
X258 hgu_sarlogic_flat_0.x4.x3.X a_n1058_3698# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X259 hgu_vgen_vref_0.mimtop1 hgu_vgen_vref_0.mimbot1 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X260 hgu_cdac_half_0.VREF hgu_cdac_half_0.d<4> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<15:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X261 VDD a_2501_8487# a_3222_8795# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X262 hgu_sarlogic_flat_0.x5.x1[5].Q_N a_19460_5284# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X263 hgu_cdac_sw_buffer_0.VDD a_n688_n1104# hgu_cdac_half_0.db<5> hgu_cdac_sw_buffer_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X264 VSS hgu_cdac_half_0.db<4> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<15:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X265 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<1:0> hgu_cdac_half_1.db<1> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.35
X266 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_0.d<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X267 hgu_sarlogic_flat_0.x2.x2.x4.x5[7].floating hgu_sarlogic_flat_0.x2.x2.x4.x10.Y hgu_sarlogic_flat_0.x2.x2.x4.x9.output_stack VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X268 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.d<6> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X269 a_10790_1868# a_10624_1868# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X270 VSS a_3326_3698# hgu_sarlogic_flat_0.x4.x30.A VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X271 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.db<6> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X272 hgu_cdac_half_0.VREF hgu_cdac_half_0.d<5> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X273 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_0.db<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X274 a_2489_15124# hgu_sarlogic_flat_0.x2.x1.x3.Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X275 VDD a_8908_6052# hgu_sarlogic_flat_0.x3.x60.Q_N VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X276 a_n607_7947# VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X277 VSS hgu_sarlogic_flat_0.x4.D[2] a_12543_1179# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X278 VDD hgu_sarlogic_flat_0.x5.eob a_14591_9880# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X279 a_7771_6925# hgu_sarlogic_flat_0.x3.x45.Q_N VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X280 VSS a_2790_6052# a_2725_6078# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0935 ps=0.965 w=0.64 l=0.15
X281 VSS hgu_sarlogic_flat_0.x3.x30.Q_N a_6935_6078# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.12 ps=1.08 w=0.42 l=0.15
X282 VSS a_n54567_7835# a_n54754_7657# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X283 a_n1158_n1744# hgu_cdac_sw_buffer_0.x11.A hgu_cdac_sw_buffer_0.VDD hgu_cdac_sw_buffer_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X284 a_n6959_12137# hgu_comp_flat_0.clk a_n7047_12137# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X285 a_5111_8513# a_4599_8487# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X286 VDD hgu_sarlogic_flat_0.x4.x30.A a_3960_3698# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X287 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.db<6> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X288 VDD a_n2219_8368# hgu_cdac_half_1.d<6> VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X289 VDD hgu_sarlogic_flat_0.x5.x3.X a_15666_6596# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X290 a_n1285_1331# a_n1189_1153# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X291 VDD hgu_sarlogic_flat_0.x4.x7.S a_140_2883# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.118 ps=1.4 w=0.42 l=0.15
X292 hgu_cdac_half_0.d<5> a_1666_n1100# hgu_cdac_sw_buffer_1.VDD hgu_cdac_sw_buffer_1.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X293 VDD VDD a_8379_1153# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0956 pd=0.875 as=0.132 ps=1.22 w=0.42 l=0.15
X294 a_4922_1363# a_4450_1153# a_5166_1545# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X295 VDD a_n2219_8368# hgu_cdac_half_1.d<6> VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X296 a_4914_8190# a_4125_7798# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0819 ps=0.81 w=0.42 l=0.15
X297 VDD hgu_sarlogic_flat_0.x4.x12.X a_5840_1868# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X298 VSS hgu_cdac_half_1.d<6> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X299 a_11317_1347# a_11626_1153# a_11561_1179# VSS sky130_fd_pr__nfet_01v8 ad=0.0486 pd=0.63 as=0.066 ps=0.745 w=0.36 l=0.15
X300 a_n2251_7253# hgu_cdac_sw_buffer_2.x9.A VSS VSS sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X301 VSS hgu_cdac_half_0.d<6> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X302 hgu_cdac_half_0.VREF hgu_cdac_half_0.db<6> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X303 a_6936_7824# a_7072_7798# a_6517_7798# VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0864 ps=0.91 w=0.64 l=0.15
X304 VSS hgu_cdac_half_1.db<6> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X305 vip hgu_tah_0.sw_n hgu_tah_0.tah_vp hgu_tah_0.VDD sky130_fd_pr__pfet_01v8 ad=0.908 pd=5.83 as=0.908 ps=5.83 w=5.5 l=0.15
X306 VSS a_2036_7824# hgu_sarlogic_flat_0.x3.x4.X VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X307 VSS hgu_sarlogic_flat_0.x4.x7.S a_140_2883# VSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.109 ps=1.36 w=0.42 l=0.15
X308 VDD VDD a_6517_7798# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.123 ps=1.17 w=0.42 l=0.15
X309 hgu_sarlogic_flat_0.x4.x9.A1 a_3960_3698# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X310 VDD a_n858_2530# a_n828_2883# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X311 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.d<6> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X312 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X313 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<7:0> hgu_cdac_half_0.db<3> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X314 VSS hgu_cdac_half_1.db<6> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X315 a_8086_6444# a_7574_6052# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X316 VDD a_n4397_8367# hgu_cdac_sw_buffer_3.x11.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X317 VSS a_190_n245# hgu_cdac_half_0.db<3> VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X318 a_4784_1868# a_3614_1868# a_4677_2234# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0486 ps=0.63 w=0.36 l=0.15
X319 hgu_sarlogic_flat_0.x2.x2.x4.x9.output_stack sample_delay_cap_ctrl_code[1] hgu_sarlogic_flat_0.x2.x2.x4.x3[1].floating VSS sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X320 hgu_sarlogic_flat_0.x4.x27.A a_3050_3698# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X321 VSS a_n1158_n1744# hgu_cdac_half_0.db<6> VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X322 hgu_cdac_half_0.VREF hgu_cdac_half_0.d<6> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X323 VSS a_7772_8487# a_8479_8513# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X324 a_n1149_11676# hgu_sarlogic_flat_0.x1.x4.x9.output_stack hgu_sarlogic_flat_0.x1.x10.A VSS sky130_fd_pr__nfet_01v8 ad=0.0651 pd=0.73 as=0.122 ps=1.42 w=0.42 l=0.15
X325 a_9404_11849# hgu_sarlogic_flat_0.x2.x2.x3.IN a_9332_11849# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X326 a_1123_11360# a_611_11594# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X327 VSS a_n2785_7946# hgu_cdac_sw_buffer_3.x7.X VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X328 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_0.d<5> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X329 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.db<6> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X330 a_11613_6078# hgu_sarlogic_flat_0.x3.x4.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X331 VSS a_17068_4644# a_17775_4670# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X332 a_10151_1179# a_9233_1453# a_9706_1363# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.0567 ps=0.69 w=0.42 l=0.15
X333 hgu_sarlogic_flat_0.x5.x3.X a_20768_8628# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X334 a_19395_5950# a_18058_5950# a_19286_5950# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X335 a_10790_1868# a_10624_1868# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X336 a_10710_14512# hgu_sarlogic_flat_0.x2.x2.x1.IN a_10638_14650# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X337 hgu_vgen_vref_0.mimtop2 VSS sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X338 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X339 VSS a_17068_5284# a_17775_5326# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X340 a_3802_1868# hgu_sarlogic_flat_0.x4.D[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X341 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.d<6> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X342 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.db<6> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.35
X343 VDD a_8814_7798# hgu_sarlogic_flat_0.x4.x17.S VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X344 a_7843_8008# a_7370_8098# a_8087_7824# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0671 ps=0.75 w=0.36 l=0.15
X345 VSS a_12155_7798# a_12154_8098# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X346 VDD hgu_sarlogic_flat_0.x3.D[0] a_8761_6951# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X347 hgu_vgen_vref_0.sky130_fd_sc_hd__inv_1_3.Y hgu_vgen_vref_0.sky130_fd_sc_hd__inv_1_3.A VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X348 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.db<6> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X349 hgu_sarlogic_flat_0.x5.eob a_2914_9360# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.175 ps=1.35 w=1 l=0.15
X350 hgu_cdac_half_1.VREF hgu_cdac_half_1.d<5> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X351 VSS a_1203_1153# hgu_sarlogic_flat_0.x4.x21.Q_N VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X352 hgu_sarlogic_flat_0.x3.x5.X a_1863_9386# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X353 a_14726_7939# hgu_sarlogic_flat_0.x5.eob a_14654_8077# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X354 hgu_vgen_vref_0.mimtop2 VSS sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X355 a_2262_1153# a_2530_1363# a_2476_1461# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X356 hgu_cdac_half_0.VREF hgu_cdac_half_0.db<5> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X357 a_2900_8879# a_1752_8513# a_2814_8513# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X358 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X359 VSS a_7228_2136# a_7176_1868# VSS sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.066 ps=0.745 w=0.42 l=0.15
X360 a_n1149_14701# hgu_sarlogic_flat_0.x1.x9.A VSS VDD sky130_fd_pr__pfet_01v8_hvt ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X361 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X362 a_9332_12401# hgu_sarlogic_flat_0.x2.x2.x3.IN a_9244_12263# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X363 a_5380_8487# a_5206_8513# a_5496_8513# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X364 hgu_tah_0.VDD a_n53930_7835# hgu_vgen_vref_0.sky130_fd_sc_hd__dlymetal6s6s_1_2.A hgu_tah_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X365 VSS hgu_cdac_half_1.d<3> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<7:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.35
X366 a_19286_5688# a_18224_5316# a_19191_5632# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X367 hgu_cdac_sw_buffer_3.x12.X a_n3651_7087# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X368 VSS hgu_cdac_half_0.d<6> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X369 a_1203_1153# a_1749_1347# a_1707_1461# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.132 pd=1.22 as=0.0882 ps=1.05 w=0.84 l=0.15
X370 a_9096_2150# a_8678_2234# a_8852_1842# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X371 VSS hgu_cdac_half_1.d<6> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X372 VSS a_n4479_7727# hgu_cdac_sw_buffer_3.x11.A VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X373 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<15:0> hgu_cdac_half_1.d<4> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X374 VSS hgu_sarlogic_flat_0.x3.x30.Q_N a_7710_6078# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.101 ps=0.99 w=0.42 l=0.15
X375 hgu_sarlogic_flat_0.x2.x2.x2.x9.output_stack hgu_sarlogic_flat_0.x2.x2.x2.x10.Y hgu_sarlogic_flat_0.x2.x2.x2.x5[7].floating VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X376 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_0.d<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X377 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.d<6> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X378 VSS a_n53647_7371# a_n53834_7113# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X379 a_4677_2234# a_3614_1868# a_4533_2150# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X380 VSS a_7575_7798# a_7510_7824# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0935 ps=0.965 w=0.64 l=0.15
X381 VDD a_1534_2530# a_1564_2883# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X382 VSS hgu_cdac_half_0.db<4> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<15:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X383 VDD hgu_sarlogic_flat_0.x4.x15.S a_10176_2883# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.0767 ps=0.785 w=0.42 l=0.15
X384 hgu_tah_0.VDD hgu_vgen_vref_0.sky130_fd_sc_hd__inv_1_3.Y a_n54752_6595# hgu_tah_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X385 VSS a_n86_n245# hgu_cdac_sw_buffer_0.x4.X VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X386 a_2268_n241# hgu_cdac_sw_buffer_1.x4.A hgu_cdac_sw_buffer_1.VDD hgu_cdac_sw_buffer_1.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X387 a_n6959_14175# hgu_comp_flat_0.ready a_n7047_14175# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X388 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<15:0> hgu_cdac_half_1.db<4> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X389 VSS a_12358_6052# a_12293_6078# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0935 ps=0.965 w=0.64 l=0.15
X390 hgu_tah_0.VDD a_n55487_7835# a_n55674_7657# hgu_tah_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X391 VSS a_n688_n1104# hgu_cdac_half_0.db<5> VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X392 a_13780_1868# hgu_sarlogic_flat_0.x4.x2.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0974 pd=0.97 as=0.0882 ps=0.84 w=0.42 l=0.15
X393 a_10280_8513# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X394 VSS hgu_cdac_sw_buffer_0.x9.X a_n1240_n1104# VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X395 hgu_cdac_half_1.d<6> a_n2219_8368# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X396 a_11600_7317# a_11153_6951# a_11507_6951# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X397 a_4124_6052# a_4437_6078# a_4543_6078# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X398 hgu_vgen_vref_0.mimtop2 VSS sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X399 VSS hgu_sarlogic_flat_0.x4.x15.S a_10183_2556# VSS sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.0693 ps=0.75 w=0.42 l=0.15
X400 a_3926_2530# hgu_sarlogic_flat_0.x4.x11.S VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X401 a_10280_8513# a_9677_8487# a_10164_8487# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X402 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_0.d<5> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X403 VSS a_11774_6925# a_11708_6951# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X404 VSS hgu_sarlogic_flat_0.x3.x27.Q_N a_4543_6078# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.12 ps=1.08 w=0.42 l=0.15
X405 VDD a_12155_7798# a_12154_8098# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X406 a_7597_6951# a_6369_6951# a_7455_7233# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X407 hgu_sarlogic_flat_0.x1.x2.x9.output_stack hgu_sarlogic_flat_0.x1.x2.x10.Y hgu_sarlogic_flat_0.x1.x2.x5[7].floating VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X408 hgu_cdac_half_1.VREF hgu_cdac_half_1.db<5> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X409 hgu_sarlogic_flat_0.x2.x2.x3.x6.SW sample_delay_offset VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X410 VSS a_1454_6950# hgu_sarlogic_flat_0.x3.x7.X VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X411 hgu_cdac_half_0.VREF hgu_cdac_half_0.db<6> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X412 VSS hgu_sarlogic_flat_0.x2.x2.x1.IN a_10638_13822# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X413 hgu_sarlogic_flat_0.x2.x2.x3.x5[7].floating hgu_sarlogic_flat_0.x2.x2.x3.x10.Y hgu_sarlogic_flat_0.x2.x2.x3.x9.output_stack VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X414 hgu_comp_flat_0.ready a_n7678_6446# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X415 a_2530_1363# a_2058_1153# a_2774_1545# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X416 a_3926_2530# hgu_sarlogic_flat_0.x4.x11.S VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X417 a_192_10793# VSS a_334_10641# VSS sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X418 a_8814_7798# a_8909_7798# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X419 VSS hgu_cdac_half_0.d<3> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<7:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.35
X420 VDD hgu_sarlogic_flat_0.x1.x9.A a_n1149_14360# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0651 ps=0.73 w=0.42 l=0.15
X421 a_4544_7824# a_4680_7798# a_4125_7798# VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0864 ps=0.91 w=0.64 l=0.15
X422 VDD a_16581_6790# a_16531_6590# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X423 a_11614_7824# hgu_sarlogic_flat_0.x3.x4.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.154 ps=1.34 w=0.64 l=0.15
X424 VDD VDD a_4125_7798# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.123 ps=1.17 w=0.42 l=0.15
X425 a_10176_2883# VSS a_9962_2883# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.193 ps=1.34 w=0.42 l=0.15
X426 hgu_vgen_vref_0.mimtop1 hgu_vgen_vref_0.mimbot1 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X427 hgu_sarlogic_flat_0.x2.x2.x1.x9.output_stack hgu_sarlogic_flat_0.x2.x2.x1.x10.Y hgu_sarlogic_flat_0.x2.x2.x1.x5[7].floating VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X428 a_5694_6444# a_5182_6052# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X429 a_13163_1153# a_13476_1179# a_13582_1179# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X430 a_66_11360# a_n134_11726# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X431 hgu_sarlogic_flat_0.x2.x2.x2.x9.output_stack sample_delay_cap_ctrl_code[10] hgu_sarlogic_flat_0.x2.x2.x2.x4[3].floating VSS sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X432 VDD a_n4479_7727# hgu_cdac_sw_buffer_3.x11.A VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X433 hgu_cdac_half_0.VREF hgu_cdac_half_0.d<6> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X434 VDD hgu_comp_flat_0.clk a_n6994_7879# VDD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X435 VSS VDD a_n422_1842# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X436 hgu_vgen_vref_0.mimtop1 hgu_vgen_vref_0.mimbot1 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X437 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<15:0> hgu_cdac_half_0.db<4> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X438 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X439 VSS hgu_sarlogic_flat_0.x2.x7.Y a_2820_11667# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X440 hgu_cdac_half_1.VREF hgu_cdac_half_1.d<2> hgu_cdac_half_1.hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.35
X441 a_12467_7317# a_11319_6951# a_12381_6951# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X442 hgu_sarlogic_flat_0.x1.x9.Y hgu_sarlogic_flat_0.x1.x9.A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X443 hgu_cdac_half_1.VREF hgu_cdac_half_1.d<6> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X444 VSS hgu_sarlogic_flat_0.x3.x4.A a_2036_7824# VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X445 VSS a_11206_7798# hgu_sarlogic_flat_0.x4.x15.S VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X446 a_n1190_n245# hgu_cdac_sw_buffer_0.x9.A hgu_cdac_sw_buffer_0.VDD hgu_cdac_sw_buffer_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X447 a_3960_3698# hgu_sarlogic_flat_0.x4.x30.A VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X448 VSS a_n1285_1331# hgu_cdac_sw_buffer_3.x9.A VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X449 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X450 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_1.d<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X451 hgu_cdac_half_1.VREF hgu_cdac_half_1.db<6> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X452 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_0.d<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X453 VDD a_611_11594# a_544_11360# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X454 hgu_vgen_vref_0.mimtop1 hgu_vgen_vref_0.phi2 hgu_tah_0.VDD VSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=0.5
X455 a_17003_5950# a_15666_5950# a_16894_5950# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X456 a_n572_1868# a_n422_1842# a_n716_1842# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X457 VSS hgu_cdac_half_1.db<5> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X458 a_4398_1545# a_3595_1153# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0787 pd=0.795 as=0.0956 ps=0.875 w=0.42 l=0.15
X459 a_12468_8879# a_11320_8513# a_12382_8513# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X460 hgu_vgen_vref_0.mimtop2 VSS sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X461 a_9522_6951# hgu_sarlogic_flat_0.x3.x42.Q_N VSS VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X462 VSS hgu_cdac_half_1.db<5> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X463 a_5451_8008# a_4978_8098# a_5695_7824# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0671 ps=0.75 w=0.36 l=0.15
X464 VDD a_13067_1331# hgu_cdac_half_1.db<0> VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X465 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.d<6> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X466 a_n6959_13347# hgu_comp_flat_0.ready a_n7047_13347# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X467 VSS a_9763_7798# a_9762_8098# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X468 hgu_comp_flat_0.comp_outn a_n6292_6446# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.54 as=0.0759 ps=0.79 w=0.46 l=0.15
X469 hgu_cdac_half_0.VREF hgu_cdac_half_0.db<3> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<7:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X470 VSS VDD a_2501_8487# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X471 a_10234_6262# a_9761_6352# a_10478_6078# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0671 ps=0.75 w=0.36 l=0.15
X472 hgu_cdac_sw_buffer_0.x11.A a_n1240_n1104# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X473 a_10163_6925# hgu_sarlogic_flat_0.x3.x42.Q_N VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X474 hgu_sarlogic_flat_0.x2.x2.x4.x5[7].floating hgu_sarlogic_flat_0.x2.x2.x4.x10.Y hgu_sarlogic_flat_0.x2.x2.x4.x9.output_stack VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X475 VDD a_9676_6925# a_10397_7233# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X476 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X477 hgu_cdac_sw_buffer_3.x11.X a_n4397_8367# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X478 hgu_cdac_half_1.VREF hgu_cdac_half_1.db<6> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X479 hgu_sarlogic_flat_0.x1.x4.x10.Y async_resetb_delay_cap_ctrl_code[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X480 VDD hgu_sarlogic_flat_0.x3.x7.X a_8288_6078# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0662 ps=0.735 w=0.42 l=0.15
X481 VSS hgu_cdac_half_0.d<6> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X482 hgu_sarlogic_flat_0.x2.x2.x2.x6.SW sample_delay_offset VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X483 a_5319_7824# a_5451_8008# a_5183_7798# VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0864 ps=0.91 w=0.64 l=0.15
X484 a_10164_8487# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X485 hgu_vgen_vref_0.phi2_n a_n54752_6595# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X486 a_16894_5688# a_15832_5316# a_16799_5632# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X487 a_10102_6078# a_10234_6262# a_9966_6052# VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0864 ps=0.91 w=0.64 l=0.15
X488 result[6] a_17775_4670# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X489 a_19460_4644# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X490 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.d<6> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X491 a_6704_2150# a_6286_2234# a_6460_1842# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X492 a_13524_2883# hgu_sarlogic_flat_0.x4.x9.A1 a_13065_2708# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X493 VSS a_19460_5924# a_19395_5950# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X494 VSS a_n7390_7871# a_n7766_6446# VSS sky130_fd_pr__nfet_01v8 ad=0.0759 pd=0.79 as=0.143 ps=1.54 w=0.46 l=0.15
X495 VSS hgu_cdac_half_0.d<3> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<7:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X496 a_18505_6316# a_18058_5950# a_18412_5950# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X497 hgu_sarlogic_flat_0.x2.x1.x3.Y VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X498 VSS hgu_cdac_half_1.db<6> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X499 hgu_tah_0.tah_vn hgu_tah_0.sw_n vin hgu_tah_0.VDD sky130_fd_pr__pfet_01v8 ad=0.908 pd=5.83 as=0.908 ps=5.83 w=5.5 l=0.15
X500 VSS a_19460_6564# a_19395_6968# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X501 a_10638_14788# hgu_sarlogic_flat_0.x2.x2.x1.IN a_10550_14650# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X502 VSS hgu_cdac_half_0.d<5> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X503 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X504 hgu_vgen_vref_0.sky130_fd_sc_hd__inv_1_2.A hgu_vgen_vref_0.sky130_fd_sc_hd__inv_1_0.A VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X505 a_2714_2883# a_2532_2883# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X506 hgu_cdac_half_0.VREF hgu_cdac_half_0.d<6> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X507 VSS a_9438_1153# a_9348_1179# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.116 ps=1.09 w=0.64 l=0.15
X508 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.db<6> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X509 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X510 a_12871_8190# a_12359_7798# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X511 a_11813_6360# a_11613_6078# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X512 VSS a_18679_5924# a_18613_5950# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X513 VSS a_13494_2530# a_13428_2556# VSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X514 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X515 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_0.d<5> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X516 a_13636_1842# hgu_sarlogic_flat_0.x4.x2.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X517 hgu_vgen_vref_0.vcm hgu_vgen_vref_0.phi1_n hgu_vgen_vref_0.mimtop2 hgu_tah_0.VDD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=0.5
X518 VSS hgu_cdac_sw_buffer_2.x4.X a_n1209_7728# VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X519 hgu_cdac_sw_buffer_0.VDD a_190_n245# hgu_cdac_half_0.db<3> hgu_cdac_sw_buffer_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X520 a_14222_1153# a_13476_1179# a_14358_1179# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X521 a_12287_8513# a_11775_8487# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X522 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X523 VSS a_18679_6564# a_18613_6968# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X524 hgu_cdac_sw_buffer_0.x8.X a_n964_n464# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X525 VSS a_1592_14732# a_1526_15136# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X526 a_9626_7233# a_9208_7317# a_9382_6925# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X527 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_1.db<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X528 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X529 hgu_sarlogic_flat_0.x4.x2.X a_n424_3698# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X530 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_0.db<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X531 a_1222_1868# a_1056_1868# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X532 VDD a_n422_1842# a_309_2150# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X533 VDD a_1448_10615# a_1478_10968# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X534 a_4679_6052# a_4977_6352# a_4913_6444# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0924 ps=0.86 w=0.42 l=0.15
X535 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_1.d<5> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X536 VDD a_9763_7798# a_9762_8098# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X537 VDD a_11538_1842# a_11488_2150# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X538 VSS hgu_sarlogic_flat_0.x2.x2.x3.x9.output_stack a_3314_11664# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X539 a_11775_8487# a_11601_8879# a_11915_8513# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X540 hgu_vgen_vref_0.mimtop1 hgu_vgen_vref_0.mimbot1 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X541 a_16041_12125# hgu_sarlogic_flat_0.x2.x2.x2.IN a_15953_11987# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X542 VSS retimer_delay_offset hgu_sarlogic_flat_0.x5.x2.x6.SW VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X543 a_9627_8795# a_9209_8879# a_9383_8487# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X544 hgu_cdac_half_1.d<5> a_n1749_7728# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X545 VSS hgu_cdac_half_0.db<2> hgu_cdac_half_0.hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT VSS sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.35
X546 a_3954_16039# hgu_sarlogic_flat_0.x2.x3.A a_3866_16177# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X547 VSS a_n542_11334# hgu_sarlogic_flat_0.x1.x3.A0 VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X548 VSS hgu_cdac_half_0.db<6> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X549 a_1732_15124# hgu_sarlogic_flat_0.x2.x1.x3.Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X550 VSS a_2036_7824# hgu_sarlogic_flat_0.x3.x4.X VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X551 a_7570_2883# hgu_sarlogic_flat_0.x4.x9.A1 a_7498_2883# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X552 hgu_cdac_half_1.VREF hgu_cdac_half_1.d<4> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<15:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X553 VDD a_3960_3698# hgu_sarlogic_flat_0.x4.x9.A1 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X554 hgu_sarlogic_flat_0.x4.x9.A1 a_3960_3698# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X555 hgu_sarlogic_flat_0.x4.x30.A a_3326_3698# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X556 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<7:0> hgu_cdac_half_0.d<3> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X557 a_13709_1347# a_14017_1453# a_13966_1545# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0787 ps=0.795 w=0.42 l=0.15
X558 a_4868_1461# a_3908_1179# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X559 hgu_cdac_half_1.VREF hgu_cdac_half_1.d<5> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X560 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X561 a_1749_1347# a_2058_1153# a_1993_1179# VSS sky130_fd_pr__nfet_01v8 ad=0.0486 pd=0.63 as=0.066 ps=0.745 w=0.36 l=0.15
X562 a_16448_14835# hgu_sarlogic_flat_0.x2.x2.x1.x9.output_stack VSS VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X563 VDD a_n4397_8367# hgu_cdac_sw_buffer_3.x11.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X564 a_11709_8513# a_11320_8513# a_11601_8879# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X565 VSS hgu_cdac_half_0.d<6> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X566 hgu_cdac_half_0.d<5> a_1666_n1100# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X567 VSS hgu_vgen_vref_0.sky130_fd_sc_hd__inv_1_4.Y a_n53014_7459# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X568 hgu_cdac_half_0.VREF hgu_cdac_half_0.d<3> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<7:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.35
X569 hgu_cdac_half_0.db<6> a_n1158_n1744# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X570 a_7570_2556# a_7316_2883# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.145 ps=1.11 w=0.42 l=0.15
X571 a_11856_7798# a_12154_8098# a_12090_8190# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0924 ps=0.86 w=0.42 l=0.15
X572 a_2820_n241# hgu_cdac_sw_buffer_1.x5.A VSS VSS sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X573 hgu_vgen_vref_0.mimtop2 VSS sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X574 a_10978_1868# hgu_sarlogic_flat_0.x4.D[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X575 VSS a_621_10615# a_555_10641# VSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X576 a_4437_6078# hgu_sarlogic_flat_0.x3.x4.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.154 ps=1.34 w=0.64 l=0.15
X577 VDD hgu_sarlogic_flat_0.x4.x17.S a_12098_2883# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.118 ps=1.4 w=0.42 l=0.15
X578 a_17068_5284# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X579 VDD a_7228_2136# a_7153_2234# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0956 pd=0.875 as=0.0787 ps=0.795 w=0.42 l=0.15
X580 VDD a_2444_2136# a_3165_1868# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X581 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_0.db<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X582 a_n6934_10472# hgu_comp_flat_0.clk a_n7022_10334# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X583 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_1.d<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X584 a_2790_6052# a_2045_6078# a_2926_6078# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X585 a_17068_5924# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X586 a_12573_8106# a_11614_7824# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X587 hgu_cdac_sw_buffer_0.VDD a_n86_n245# hgu_cdac_sw_buffer_0.x4.X hgu_cdac_sw_buffer_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X588 VSS hgu_sarlogic_flat_0.x3.x3.A a_1422_7824# VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X589 VSS a_1164_n241# hgu_cdac_sw_buffer_1.x9.X VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X590 a_2006_1545# a_1203_1153# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0787 pd=0.795 as=0.0956 ps=0.875 w=0.42 l=0.15
X591 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X592 VSS hgu_sarlogic_flat_0.x4.x17.S a_12098_2883# VSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.109 ps=1.36 w=0.42 l=0.15
X593 a_n4397_8367# hgu_cdac_sw_buffer_3.x11.A VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X594 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_0.d<5> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X595 VSS a_14404_2136# a_14352_1868# VSS sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.066 ps=0.745 w=0.42 l=0.15
X596 a_1222_1868# a_1056_1868# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X597 a_7314_1363# a_6841_1453# a_7558_1179# VSS sky130_fd_pr__nfet_01v8 ad=0.0675 pd=0.735 as=0.0671 ps=0.75 w=0.36 l=0.15
X598 VSS hgu_cdac_half_1.d<5> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X599 VSS hgu_cdac_half_0.d<2> hgu_cdac_half_0.hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X600 VDD a_10675_1331# hgu_cdac_half_1.db<1> VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X601 a_1196_n1740# hgu_cdac_sw_buffer_1.x11.A hgu_cdac_sw_buffer_1.VDD hgu_cdac_sw_buffer_1.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X602 a_3929_14512# hgu_sarlogic_flat_0.x2.x3.A a_3841_14374# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X603 hgu_cdac_half_1.d<4> a_n1209_7728# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X604 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_1.db<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X605 a_15832_4670# a_15666_4670# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X606 VSS a_n1209_7728# hgu_cdac_half_1.d<4> VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X607 a_611_11594# a_879_11334# a_825_11360# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X608 a_n2785_7946# VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X609 a_15832_5316# a_15666_5316# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X610 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X611 a_13462_2234# a_13182_1868# a_13370_1868# VSS sky130_fd_pr__nfet_01v8 ad=0.0675 pd=0.735 as=0.066 ps=0.745 w=0.36 l=0.15
X612 a_16088_10322# hgu_sarlogic_flat_0.x2.x2.x2.IN a_16000_10460# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X613 a_n220_1179# a_n335_1453# a_n643_1347# VSS sky130_fd_pr__nfet_01v8 ad=0.116 pd=1.09 as=0.0486 ps=0.63 w=0.36 l=0.15
X614 hgu_cdac_half_1.VREF hgu_cdac_half_1.db<5> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X615 hgu_sarlogic_flat_0.x1.x4.x4[3].floating async_resetb_delay_cap_ctrl_code[2] hgu_sarlogic_flat_0.x1.x4.x9.output_stack VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X616 VDD hgu_sarlogic_flat_0.x3.x7.X a_5896_6078# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0662 ps=0.735 w=0.42 l=0.15
X617 hgu_cdac_half_1.hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT hgu_cdac_half_1.db<2> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X618 a_11206_7798# a_11301_7798# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X619 VDD a_10163_6925# a_10075_7317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X620 hgu_vgen_vref_0.mimtop2 VSS sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X621 a_7182_1179# a_7314_1363# a_7046_1153# VSS sky130_fd_pr__nfet_01v8 ad=0.0974 pd=0.97 as=0.0864 ps=0.91 w=0.64 l=0.15
X622 a_3639_2883# hgu_sarlogic_flat_0.x4.x11.S VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X623 hgu_cdac_sw_buffer_1.VDD a_1196_n1740# hgu_cdac_half_0.d<6> hgu_cdac_sw_buffer_1.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X624 a_6517_7798# a_6830_7824# a_6936_7824# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X625 VSS hgu_sarlogic_flat_0.x4.x27.A a_3326_3698# VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X626 hgu_comp_flat_0.P hgu_tah_0.tah_vp a_n7660_7467# VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X627 a_18819_5676# a_18973_5510# a_18679_5284# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X628 a_19286_4670# a_18058_4670# a_19144_4952# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X629 hgu_sarlogic_flat_0.x4.x20.X a_14746_2883# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.158 ps=1.39 w=1 l=0.15
X630 hgu_cdac_half_0.VREF hgu_cdac_half_0.d<6> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X631 a_11084_1179# hgu_sarlogic_flat_0.x4.x2.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X632 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.db<6> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X633 a_1592_14732# a_1418_14758# a_1732_15124# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X634 a_3639_2556# hgu_sarlogic_flat_0.x4.x11.S VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X635 a_2489_15124# a_1886_14958# a_2373_14732# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X636 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X637 VDD a_10164_8487# a_10076_8879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X638 a_18923_4952# a_18505_5036# a_18679_4644# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X639 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X640 hgu_vgen_vref_0.mimtop2 VSS sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X641 hgu_sarlogic_flat_0.x1.x4.x2.floating async_resetb_delay_cap_ctrl_code[0] hgu_sarlogic_flat_0.x1.x4.x9.output_stack VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.124 ps=1.43 w=0.42 l=0.15
X642 hgu_tah_0.VDD a_n54850_7371# hgu_vgen_vref_0.sky130_fd_sc_hd__dlymetal6s6s_1_5.A hgu_tah_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X643 a_4143_6951# a_3977_6951# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X644 hgu_cdac_half_0.VREF hgu_cdac_half_0.d<3> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<7:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X645 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X646 a_342_11360# a_n447_11350# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0819 ps=0.81 w=0.42 l=0.15
X647 result[3] a_20167_5950# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X648 a_13462_2234# a_13016_1868# a_13370_1868# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0651 ps=0.73 w=0.42 l=0.15
X649 VSS hgu_cdac_half_1.db<4> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<15:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X650 VDD a_n2219_8368# hgu_cdac_half_1.d<6> VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X651 hgu_comp_flat_0.comp_outp a_n7216_6420# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0759 pd=0.79 as=0.0759 ps=0.79 w=0.46 l=0.15
X652 a_7305_6078# a_6516_6052# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0588 ps=0.7 w=0.42 l=0.15
X653 VDD hgu_sarlogic_flat_0.x5.x3.X a_18058_5950# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X654 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X655 hgu_cdac_half_0.VREF hgu_cdac_half_0.d<5> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X656 hgu_sarlogic_flat_0.x2.x2.x1.x9.output_stack hgu_sarlogic_flat_0.x2.x2.x1.x10.Y hgu_sarlogic_flat_0.x2.x2.x1.x5[7].floating VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X657 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X658 a_4212_1868# hgu_sarlogic_flat_0.x4.x2.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0974 pd=0.97 as=0.0882 ps=0.84 w=0.42 l=0.15
X659 hgu_cdac_half_0.d<6> a_1196_n1740# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X660 VDD VDD a_13163_1153# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0956 pd=0.875 as=0.132 ps=1.22 w=0.42 l=0.15
X661 a_5889_2708# hgu_sarlogic_flat_0.x4.x9.A1 a_6031_2556# VSS sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X662 a_n7760_6349# a_n6526_6819# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.3 as=0.139 ps=1.17 w=0.84 l=0.15
X663 VSS hgu_sarlogic_flat_0.x4.D[1] a_11153_6951# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X664 hgu_cdac_sw_buffer_2.x5.A a_10341_1868# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X665 a_19144_6590# a_18679_6564# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X666 VSS a_2036_7824# hgu_sarlogic_flat_0.x3.x4.X VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X667 VSS hgu_cdac_half_1.db<5> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X668 hgu_sarlogic_flat_0.x3.x4.A a_1422_7824# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X669 hgu_sarlogic_flat_0.x4.x9.A1 a_3960_3698# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X670 hgu_sarlogic_flat_0.x4.x7.X a_394_2883# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.113 ps=1.04 w=0.65 l=0.15
X671 VSS hgu_cdac_half_1.db<6> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X672 a_11720_7824# a_11856_7798# a_11301_7798# VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0864 ps=0.91 w=0.64 l=0.15
X673 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<1:0> hgu_cdac_half_1.d<1> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.122 ps=1.42 w=0.42 l=0.35
X674 a_4030_7798# a_4125_7798# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X675 hgu_cdac_half_1.VREF hgu_cdac_half_1.d<4> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<15:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.35
X676 VDD a_n4397_8367# hgu_cdac_sw_buffer_3.x11.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X677 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_1.db<5> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X678 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.db<6> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X679 a_n6887_12275# hgu_comp_flat_0.clk a_n6959_12275# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X680 VSS a_1196_n1740# hgu_cdac_half_0.d<6> VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X681 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<0> hgu_cdac_half_1.d<0> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.244 ps=2.26 w=0.84 l=0.35
X682 hgu_tah_0.tah_vp hgu_tah_0.sw_n hgu_tah_0.tah_vp VSS sky130_fd_pr__nfet_01v8 ad=4.43 pd=30.7 as=0.454 ps=3.08 w=2.75 l=0.15
X683 VSS hgu_cdac_half_0.d<4> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<15:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X684 VDD a_n2219_8368# hgu_cdac_half_1.d<6> VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X685 hgu_vgen_vref_0.phi2 a_n55304_6595# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X686 VSS hgu_cdac_half_0.d<6> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.35
X687 VSS a_n595_7253# hgu_cdac_half_1.d<2> VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X688 a_16113_12401# hgu_sarlogic_flat_0.x2.x2.x2.IN a_16041_12401# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X689 a_12382_8513# a_11320_8513# a_12287_8513# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X690 VSS a_4125_7798# hgu_sarlogic_flat_0.x3.x48.Q_N VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X691 a_19576_5676# a_18973_5510# a_19460_5284# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X692 hgu_sarlogic_flat_0.x2.x2.x4.x5[7].floating hgu_sarlogic_flat_0.x2.x2.x4.x10.Y hgu_sarlogic_flat_0.x2.x2.x4.x9.output_stack VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X693 VDD a_5380_8487# a_6087_8513# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X694 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<7:0> hgu_cdac_half_0.d<3> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X695 VDD sample_delay_cap_ctrl_code[15] hgu_sarlogic_flat_0.x2.x2.x3.x10.Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X696 VSS hgu_cdac_half_0.d<5> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.35
X697 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_0.db<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X698 a_16197_6590# a_15666_6596# a_16113_6590# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X699 VDD a_11205_6052# hgu_sarlogic_flat_0.x4.D[3] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X700 hgu_cdac_half_0.VREF hgu_cdac_half_0.d<6> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X701 a_3595_1153# a_3908_1179# a_4014_1179# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X702 VDD a_4836_2136# a_4761_2234# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0956 pd=0.875 as=0.0787 ps=0.795 w=0.42 l=0.15
X703 a_12627_8008# a_12154_8098# a_12871_7824# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0671 ps=0.75 w=0.36 l=0.15
X704 VDD a_5987_1153# hgu_sarlogic_flat_0.x4.x26.Q_N VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X705 hgu_cdac_half_0.hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT hgu_cdac_half_0.db<2> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.35
X706 VDD a_3497_2708# hgu_sarlogic_flat_0.x4.x10.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X707 VDD hgu_cdac_sw_buffer_3.x3.X a_n3927_7727# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X708 a_52_2136# hgu_sarlogic_flat_0.x4.x2.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.132 pd=1.22 as=0.0956 ps=0.875 w=0.42 l=0.15
X709 VSS hgu_sarlogic_flat_0.x2.x2.x1.IN a_9739_15176# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0651 ps=0.73 w=0.42 l=0.15
X710 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X711 a_9332_11987# hgu_sarlogic_flat_0.x2.x2.x3.IN a_9244_11987# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X712 a_16427_6956# a_16581_6790# a_16287_6564# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X713 a_583_1179# a_n335_1453# a_138_1363# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.0567 ps=0.69 w=0.42 l=0.15
X714 VDD a_17068_5284# a_16980_5310# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X715 hgu_cdac_sw_buffer_0.x11.A a_n1240_n1104# hgu_cdac_sw_buffer_0.VDD hgu_cdac_sw_buffer_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X716 a_14661_2150# a_14245_2234# a_14404_2136# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.132 ps=1.22 w=0.84 l=0.15
X717 VSS hgu_cdac_half_1.d<5> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X718 a_10098_6951# a_8761_6951# a_9989_6951# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X719 hgu_tah_0.VDD hgu_vgen_vref_0.sky130_fd_sc_hd__inv_1_2.Y a_n54752_8227# hgu_tah_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X720 hgu_cdac_sw_buffer_0.x8.X a_n964_n464# hgu_cdac_sw_buffer_0.VDD hgu_cdac_sw_buffer_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X721 VDD a_17068_5924# a_16980_6316# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X722 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X723 VSS hgu_cdac_half_1.d<6> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X724 hgu_sarlogic_flat_0.x2.x2.x2.x3[1].floating sample_delay_cap_ctrl_code[9] hgu_sarlogic_flat_0.x2.x2.x2.x9.output_stack VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X725 a_n6934_10748# hgu_comp_flat_0.clk a_n7022_10610# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X726 VSS hgu_sarlogic_flat_0.x4.x17.S a_3518_9386# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0786 ps=0.805 w=0.42 l=0.15
X727 VDD a_2262_1153# a_2195_1545# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X728 VSS hgu_cdac_half_1.d<6> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X729 a_n1149_14360# hgu_sarlogic_flat_0.x1.x2.x9.output_stack VSS VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X730 VSS hgu_cdac_half_1.db<4> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<15:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X731 hgu_cdac_sw_buffer_3.x12.X a_n3651_7087# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X732 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<15:0> hgu_cdac_half_1.d<4> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X733 result[5] a_20167_5326# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X734 VDD hgu_sarlogic_flat_0.x4.x30.A a_3960_3698# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X735 VSS a_n424_3698# hgu_sarlogic_flat_0.x4.x2.X VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X736 hgu_cdac_half_0.VREF hgu_cdac_half_0.d<2> hgu_cdac_half_0.hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X737 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_1.d<5> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X738 VSS hgu_cdac_half_1.db<6> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X739 a_108_11334# a_406_11482# a_342_11360# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0924 ps=0.86 w=0.42 l=0.15
X740 hgu_tah_0.sw_n a_1945_10648# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X741 a_4790_1179# a_4922_1363# a_4654_1153# VSS sky130_fd_pr__nfet_01v8 ad=0.0974 pd=0.97 as=0.0864 ps=0.91 w=0.64 l=0.15
X742 hgu_sarlogic_flat_0.x3.x36.Q_N a_12556_8487# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X743 hgu_cdac_half_1.VREF hgu_cdac_half_1.d<5> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X744 hgu_cdac_half_1.d<6> a_n2219_8368# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X745 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.d<6> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X746 VSS a_n54850_7835# hgu_vgen_vref_0.sky130_fd_sc_hd__dlymetal6s6s_1_3.A VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X747 a_n1147_7253# hgu_cdac_sw_buffer_2.x4.A VSS VSS sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X748 a_16894_4670# a_15666_4670# a_16752_4952# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X749 a_1468_2556# VSS a_1105_2708# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X750 a_10663_15763# hgu_sarlogic_flat_0.x2.x2.x1.IN a_10575_15901# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X751 hgu_cdac_half_1.d<6> a_n2219_8368# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X752 a_14017_1453# hgu_sarlogic_flat_0.x4.x20.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X753 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X754 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_1.db<5> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X755 VDD hgu_cdac_sw_buffer_2.x11.A a_n2219_8368# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X756 a_2347_8513# hgu_sarlogic_flat_0.x3.x4.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X757 a_18412_6590# hgu_sarlogic_flat_0.x4.D[1] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X758 a_16088_10598# hgu_sarlogic_flat_0.x2.x2.x2.IN a_16000_10736# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X759 VSS hgu_sarlogic_flat_0.x4.x10.X a_3448_1868# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X760 VDD a_9967_7798# a_9900_8190# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X761 VSS a_n424_3698# hgu_sarlogic_flat_0.x4.x2.X VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X762 VSS sample_delay_cap_ctrl_code[11] hgu_sarlogic_flat_0.x2.x2.x2.x10.Y VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X763 a_n55204_7835# hgu_vgen_vref_0.sky130_fd_sc_hd__dlymetal6s6s_1_3.A hgu_tah_0.VDD hgu_tah_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.141 ps=1.33 w=0.42 l=0.15
X764 a_4913_6078# a_4124_6052# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0588 ps=0.7 w=0.42 l=0.15
X765 a_4068_1842# hgu_sarlogic_flat_0.x4.x2.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X766 VSS a_1945_10648# hgu_tah_0.sw_n VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X767 a_17184_6956# a_16581_6790# a_17068_6564# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X768 a_1820_1868# hgu_sarlogic_flat_0.x4.x2.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0974 pd=0.97 as=0.0882 ps=0.84 w=0.42 l=0.15
X769 a_1137_14764# a_971_14764# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X770 VSS hgu_cdac_half_1.d<6> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X771 hgu_tah_0.VDD a_n54752_6595# hgu_vgen_vref_0.phi2_n hgu_tah_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X772 hgu_cdac_half_0.VREF hgu_cdac_half_0.db<5> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X773 VDD hgu_cdac_sw_buffer_3.x11.A a_n4397_8367# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X774 a_4587_1545# a_4450_1153# a_4141_1347# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X775 a_n6934_15564# hgu_comp_flat_0.ready a_n7022_15702# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X776 a_16752_6590# a_16287_6564# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X777 VDD hgu_sarlogic_flat_0.x5.x3.X a_15666_5316# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X778 a_14746_2883# hgu_sarlogic_flat_0.x4.x9.A1 a_14674_2883# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X779 a_9739_15176# hgu_sarlogic_flat_0.x2.x2.x1.IN VSS VDD sky130_fd_pr__pfet_01v8_hvt ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X780 VSS hgu_cdac_half_1.db<6> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X781 VSS hgu_sarlogic_flat_0.x3.x5.X a_8762_8513# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X782 hgu_sarlogic_flat_0.x5.x2.x2.floating retimer_delay_code[0] hgu_sarlogic_flat_0.x5.x2.x9.output_stack VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.124 ps=1.43 w=0.42 l=0.15
X783 hgu_vgen_vref_0.mimtop2 VSS sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X784 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.d<6> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X785 hgu_vgen_vref_0.phi1_n a_n54752_8227# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X786 VDD a_18973_5924# a_18923_6232# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X787 hgu_cdac_half_0.d<6> a_1196_n1740# hgu_cdac_sw_buffer_1.VDD hgu_cdac_sw_buffer_1.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X788 a_n53647_7371# a_n53551_7113# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X789 a_14746_2556# a_14492_2883# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.145 ps=1.11 w=0.42 l=0.15
X790 VSS VDD a_12495_7824# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.101 ps=0.99 w=0.42 l=0.15
X791 a_6990_6925# hgu_sarlogic_flat_0.x3.x45.Q_N VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X792 a_1502_14758# a_971_14764# a_1418_14758# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X793 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X794 VSS a_1666_n1100# hgu_cdac_half_0.d<5> VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X795 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_1.db<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X796 a_19694_4952# a_19286_4670# a_19460_4644# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X797 a_3960_3698# hgu_sarlogic_flat_0.x4.x30.A VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X798 hgu_cdac_sw_buffer_0.x11.A a_n1240_n1104# hgu_cdac_sw_buffer_0.VDD hgu_cdac_sw_buffer_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X799 hgu_cdac_half_1.VREF hgu_cdac_half_1.db<6> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X800 a_6516_6052# a_7071_6052# a_7029_6360# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0882 ps=1.05 w=0.84 l=0.15
X801 a_n6959_12551# hgu_comp_flat_0.clk a_n7047_12413# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X802 a_7071_6052# a_7370_6052# a_7305_6078# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.066 ps=0.745 w=0.36 l=0.15
X803 a_9379_10874# hgu_sarlogic_flat_0.x2.x2.x3.IN hgu_sarlogic_flat_0.x2.x2.x3.x9.output_stack VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X804 VSS a_5380_8487# a_6087_8513# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X805 hgu_cdac_half_0.VREF hgu_cdac_half_0.d<4> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<15:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X806 VDD a_2988_8487# a_3695_8513# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X807 a_6991_8487# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X808 a_8005_7233# a_7597_6951# a_7771_6925# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X809 a_608_2883# VSS a_394_2883# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.193 ps=1.34 w=0.42 l=0.15
X810 hgu_cdac_sw_buffer_0.VDD a_454_n939# hgu_cdac_sw_buffer_0.x7.X hgu_cdac_sw_buffer_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X811 hgu_cdac_half_0.db<5> a_n688_n1104# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X812 hgu_cdac_half_0.VREF hgu_cdac_half_0.d<6> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.35
X813 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X814 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_0.d<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X815 VDD hgu_sarlogic_flat_0.x4.x11.S a_5390_2883# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.0767 ps=0.785 w=0.42 l=0.15
X816 VDD hgu_sarlogic_flat_0.x4.x3.X a_n424_3698# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X817 a_1203_1153# a_1516_1179# a_1622_1179# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X818 VSS hgu_cdac_half_0.db<3> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<7:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X819 VDD hgu_sarlogic_flat_0.x4.x10.X a_3448_1868# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X820 hgu_vgen_vref_0.mimtop1 hgu_vgen_vref_0.mimbot1 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X821 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_0.d<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X822 hgu_cdac_half_1.VREF hgu_cdac_half_1.db<3> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<7:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.35
X823 hgu_cdac_sw_buffer_0.VDD a_n1158_n1744# hgu_cdac_half_0.db<6> hgu_cdac_sw_buffer_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X824 VDD a_3595_1153# hgu_sarlogic_flat_0.x4.x24.Q_N VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X825 a_8006_8795# a_7598_8513# a_7772_8487# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X826 hgu_cdac_sw_buffer_3.x11.X a_n4397_8367# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X827 hgu_vgen_vref_0.mimtop2 VSS sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X828 hgu_cdac_half_0.VREF hgu_cdac_half_0.d<5> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.35
X829 VSS hgu_sarlogic_flat_0.x4.x11.S a_5397_2556# VSS sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.0693 ps=0.75 w=0.42 l=0.15
X830 a_621_10615# hgu_sarlogic_flat_0.x5.eob VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X831 hgu_cdac_half_0.VREF hgu_cdac_half_0.db<6> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X832 a_n1149_11676# hgu_sarlogic_flat_0.x1.x10.A VDD VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X833 hgu_cdac_half_0.VREF hgu_cdac_half_0.db<6> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X834 a_17068_5284# a_16894_5688# a_17184_5676# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X835 VDD a_3960_3698# hgu_sarlogic_flat_0.x4.x9.A1 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X836 hgu_cdac_sw_buffer_1.VDD hgu_cdac_sw_buffer_1.x11.A a_1196_n1740# hgu_cdac_sw_buffer_1.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X837 VDD VDD a_n130_1153# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X838 hgu_cdac_half_0.VREF hgu_cdac_half_0.db<4> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<15:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X839 VSS a_n53930_7371# hgu_vgen_vref_0.sky130_fd_sc_hd__dlymetal6s6s_1_4.A VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X840 a_9364_1868# a_8852_1842# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.116 pd=1.09 as=0.166 ps=1.8 w=0.64 l=0.15
X841 VSS hgu_cdac_half_1.d<6> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X842 hgu_sarlogic_flat_0.x1.x2.x9.output_stack async_setb_delay_cap_ctrl_code[1] hgu_sarlogic_flat_0.x1.x2.x3[1].floating VSS sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X843 a_11709_2150# a_11244_1842# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X844 a_7707_8513# a_6370_8513# a_7598_8513# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X845 VSS hgu_cdac_half_1.db<6> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X846 a_2141_8513# a_1752_8513# a_2033_8879# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X847 a_n6887_13485# hgu_comp_flat_0.ready a_n6959_13485# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X848 hgu_tah_0.VDD a_n55770_7835# hgu_vgen_vref_0.sky130_fd_sc_hd__inv_1_0.A hgu_tah_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X849 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<7:0> hgu_cdac_half_1.d<3> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.35
X850 VSS hgu_cdac_half_1.db<6> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X851 a_n3325_7252# hgu_cdac_sw_buffer_3.x4.A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X852 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X853 a_5390_2883# VSS a_5176_2883# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.193 ps=1.34 w=0.42 l=0.15
X854 hgu_cdac_half_1.VREF hgu_cdac_half_1.d<4> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<15:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X855 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_0.db<5> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X856 a_3978_2234# a_3614_1868# a_3894_2234# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X857 hgu_sarlogic_flat_0.x3.x33.Q_N a_10164_8487# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X858 VSS a_n55487_7371# a_n55674_7113# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X859 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X860 a_9698_7824# a_8909_7798# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0588 ps=0.7 w=0.42 l=0.15
X861 a_2373_14732# a_2199_15136# a_2489_15124# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X862 hgu_cdac_half_1.VREF hgu_cdac_half_1.d<5> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.35
X863 hgu_cdac_half_1.VREF hgu_cdac_half_1.db<4> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<15:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X864 a_9522_6951# a_9676_6925# a_9382_6925# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X865 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<15:0> hgu_cdac_half_0.d<4> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X866 a_11625_1453# hgu_sarlogic_flat_0.x4.x17.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X867 hgu_sarlogic_flat_0.x2.x2.x4.x9.output_stack hgu_sarlogic_flat_0.x2.x3.A a_3929_14788# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X868 a_9967_7798# a_9222_7824# a_10103_7824# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X869 a_11388_1868# hgu_sarlogic_flat_0.x4.x2.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0974 pd=0.97 as=0.0882 ps=0.84 w=0.42 l=0.15
X870 VSS a_10163_6925# a_10098_6951# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X871 a_16020_6590# hgu_sarlogic_flat_0.x3.D[0] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X872 VSS hgu_sarlogic_flat_0.x5.x3.X a_15666_5950# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X873 hgu_sarlogic_flat_0.x5.x2.x9.output_stack hgu_sarlogic_flat_0.x5.eob a_14654_8491# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X874 a_8786_1868# a_8232_1868# a_8678_2234# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0675 ps=0.735 w=0.36 l=0.15
X875 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.122 ps=1.42 w=0.42 l=0.35
X876 hgu_sarlogic_flat_0.x4.x31.Q_N a_12012_2136# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X877 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X878 hgu_cdac_half_1.d<5> a_n1749_7728# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X879 VDD hgu_sarlogic_flat_0.x3.x4.A a_2036_7824# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X880 VSS hgu_sarlogic_flat_0.x5.x3.X a_15666_6596# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X881 VSS a_1196_n1740# hgu_cdac_half_0.d<6> VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X882 VDD hgu_sarlogic_flat_0.x4.x3.X a_n424_3698# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X883 hgu_cdac_half_0.VREF hgu_cdac_half_0.db<6> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X884 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<15:0> hgu_cdac_half_1.db<4> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.35
X885 a_1676_1842# hgu_sarlogic_flat_0.x4.x2.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X886 VSS a_2036_7824# hgu_sarlogic_flat_0.x3.x4.X VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X887 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X888 a_2262_1153# a_1516_1179# a_2398_1179# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X889 VDD hgu_sarlogic_flat_0.x4.x13.S a_7316_2883# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.118 ps=1.4 w=0.42 l=0.15
X890 hgu_cdac_sw_buffer_3.x8.X a_n4203_7087# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X891 hgu_sarlogic_flat_0.x4.x30.A a_3326_3698# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X892 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<7:0> hgu_cdac_half_1.d<3> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X893 hgu_sarlogic_flat_0.x1.x10.Y hgu_sarlogic_flat_0.x1.x10.A VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X894 VSS a_2914_9360# hgu_sarlogic_flat_0.x5.eob VSS sky130_fd_pr__nfet_01v8 ad=0.107 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X895 a_18679_6564# a_18505_6590# a_18819_6956# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X896 a_16113_5310# a_15666_5316# a_16020_5310# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X897 a_13780_1868# a_13930_1842# a_13636_1842# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X898 hgu_vgen_vref_0.mimtop1 hgu_vgen_vref_0.mimbot1 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X899 VDD VDD a_3595_1153# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0956 pd=0.875 as=0.132 ps=1.22 w=0.42 l=0.15
X900 VSS a_52_2136# a_773_1868# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X901 VSS a_1863_9386# hgu_sarlogic_flat_0.x3.x5.X VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X902 VSS hgu_cdac_half_0.db<2> hgu_cdac_half_0.hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X903 VSS hgu_cdac_half_1.d<4> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<15:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X904 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.d<6> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X905 hgu_cdac_half_0.d<6> a_1196_n1740# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X906 VDD hgu_sarlogic_flat_0.x4.D[5] a_5367_1179# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X907 VSS hgu_sarlogic_flat_0.x4.x13.S a_7316_2883# VSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.109 ps=1.36 w=0.42 l=0.15
X908 hgu_comp_flat_0.Q hgu_tah_0.tah_vn a_n7660_7467# VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X909 a_14017_1453# hgu_sarlogic_flat_0.x4.x20.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X910 VDD a_6318_2530# a_6348_2883# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X911 VDD a_16581_5510# a_16531_5310# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X912 VSS hgu_cdac_half_0.d<6> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X913 hgu_cdac_sw_buffer_1.x11.A a_1114_n1100# hgu_cdac_sw_buffer_1.VDD hgu_cdac_sw_buffer_1.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X914 a_n55204_7371# hgu_vgen_vref_0.sky130_fd_sc_hd__dlymetal6s6s_1_5.A hgu_tah_0.VDD hgu_tah_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.141 ps=1.33 w=0.42 l=0.15
X915 a_1732_6052# a_2045_6078# a_2151_6078# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X916 hgu_cdac_half_1.VREF hgu_cdac_half_1.d<6> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X917 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.db<6> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X918 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X919 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_1.d<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X920 VDD a_4124_6052# hgu_sarlogic_flat_0.x3.x54.Q_N VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X921 hgu_cdac_half_1.VREF hgu_cdac_half_1.d<6> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X922 hgu_cdac_half_1.VREF hgu_cdac_half_1.db<6> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X923 VSS hgu_sarlogic_flat_0.x3.x20.Q_N a_2151_6078# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.12 ps=1.08 w=0.42 l=0.15
X924 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.d<6> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X925 a_1749_1347# a_2057_1453# a_2006_1545# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0787 ps=0.795 w=0.42 l=0.15
X926 VSS a_2988_8487# a_3695_8513# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X927 VDD hgu_sarlogic_flat_0.x3.x5.X a_6370_8513# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X928 a_n4397_8367# hgu_cdac_sw_buffer_3.x11.A VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X929 VDD a_7370_6052# a_7369_6352# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X930 VSS hgu_cdac_half_1.db<5> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X931 VDD hgu_sarlogic_flat_0.x5.x3.X a_15666_4670# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X932 VSS a_n1158_n1744# hgu_cdac_half_0.db<6> VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X933 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_1.db<5> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X934 VDD hgu_tah_0.sw_n a_1146_7824# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X935 VSS a_1666_n1100# hgu_cdac_half_0.d<5> VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X936 a_2373_14732# hgu_sarlogic_flat_0.x2.x1.x3.Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X937 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_0.d<5> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X938 hgu_tah_0.VDD hgu_vgen_vref_0.sky130_fd_sc_hd__inv_1_3.A a_n55304_6595# hgu_tah_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X939 hgu_cdac_half_1.VREF hgu_cdac_half_1.d<1> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<1:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.35
X940 a_n6959_12827# hgu_comp_flat_0.clk a_n7047_12689# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X941 hgu_tah_0.VDD hgu_vgen_vref_0.clk hgu_vgen_vref_0.sky130_fd_sc_hd__inv_1_4.Y hgu_tah_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X942 VSS hgu_cdac_half_0.db<5> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X943 VDD hgu_sarlogic_flat_0.x2.x2.x2.IN a_16448_14835# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0651 ps=0.73 w=0.42 l=0.15
X944 a_n828_2883# hgu_sarlogic_flat_0.x4.x9.A1 a_n1287_2708# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X945 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_0.d<5> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X946 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_0.db<5> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X947 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X948 VDD a_11301_7798# hgu_sarlogic_flat_0.x3.x39.Q_N VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X949 a_14726_7663# hgu_sarlogic_flat_0.x5.eob a_14654_7663# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X950 hgu_cdac_half_1.VREF hgu_cdac_half_1.db<5> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X951 hgu_sarlogic_flat_0.x3.x4.X a_2036_7824# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X952 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X953 hgu_sarlogic_flat_0.x1.x2.x5[7].floating hgu_sarlogic_flat_0.x1.x2.x10.Y hgu_sarlogic_flat_0.x1.x2.x9.output_stack VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X954 a_6972_1868# a_6460_1842# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.116 pd=1.09 as=0.166 ps=1.8 w=0.64 l=0.15
X955 a_5093_2150# a_4677_2234# a_4836_2136# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.132 ps=1.22 w=0.84 l=0.15
X956 VSS a_2444_2136# a_2392_1868# VSS sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.066 ps=0.745 w=0.42 l=0.15
X957 a_n572_1868# hgu_sarlogic_flat_0.x4.x2.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0974 pd=0.97 as=0.0882 ps=0.84 w=0.42 l=0.15
X958 VSS hgu_cdac_half_1.d<6> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X959 hgu_sarlogic_flat_0.x1.x4.x5[7].floating hgu_sarlogic_flat_0.x1.x4.x10.Y hgu_sarlogic_flat_0.x1.x4.x9.output_stack VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X960 VDD a_n1749_7728# hgu_cdac_half_1.d<5> VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X961 VDD VDD a_7575_7798# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X962 VSS a_n858_2530# a_n924_2556# VSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X963 hgu_sarlogic_flat_0.x4.x7.S a_6087_8513# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X964 VDD a_8852_1842# a_8762_2234# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X965 hgu_sarlogic_flat_0.x5.x2.x9.output_stack hgu_sarlogic_flat_0.x5.x2.x10.Y hgu_sarlogic_flat_0.x5.x2.x5[7].floating VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X966 hgu_vgen_vref_0.mimtop2 hgu_vgen_vref_0.phi2_n hgu_vgen_vref_0.mimbot1 hgu_tah_0.VDD sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=0.5
X967 VDD a_7574_6052# a_7507_6444# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X968 VSS hgu_cdac_sw_buffer_3.x4.X a_n3387_7727# VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X969 a_12342_1545# a_11830_1153# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X970 VSS a_17068_5924# a_17003_5950# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X971 VSS a_n1158_n1744# hgu_cdac_half_0.db<6> VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X972 VSS a_8283_1331# hgu_cdac_sw_buffer_3.x5.A VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X973 a_n447_11350# a_n134_11726# a_n28_11682# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X974 a_12870_6078# a_12358_6052# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.084 ps=0.82 w=0.42 l=0.15
X975 VDD a_n1189_1153# hgu_cdac_sw_buffer_0.x9.A VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X976 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X977 VSS a_n1209_7728# hgu_cdac_half_1.d<4> VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X978 hgu_sarlogic_flat_0.x5.x1[6].Q_N a_17068_4644# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X979 a_1502_2234# a_1222_1868# a_1410_1868# VSS sky130_fd_pr__nfet_01v8 ad=0.0675 pd=0.735 as=0.066 ps=0.745 w=0.36 l=0.15
X980 a_n6959_13761# hgu_comp_flat_0.ready a_n7047_13623# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X981 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X982 hgu_sarlogic_flat_0.x5.x2.x9.output_stack hgu_sarlogic_flat_0.x5.x2.x6.SW hgu_sarlogic_flat_0.x5.x2.x6.floating VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X983 a_7130_6951# hgu_sarlogic_flat_0.x3.x45.Q_N VSS VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X984 VSS a_17068_6564# a_17003_6968# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X985 hgu_vgen_vref_0.sky130_fd_sc_hd__inv_1_2.Y hgu_vgen_vref_0.sky130_fd_sc_hd__inv_1_2.A VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X986 a_n7660_7467# hgu_tah_0.tah_vp hgu_comp_flat_0.P VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X987 hgu_vgen_vref_0.mimtop1 hgu_vgen_vref_0.mimbot1 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X988 hgu_cdac_sw_buffer_2.x6.A a_7949_1868# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X989 hgu_cdac_half_1.VREF hgu_cdac_half_1.d<6> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X990 a_n424_3698# hgu_sarlogic_flat_0.x4.x3.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X991 VDD VDD a_13930_1842# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.17 ps=1.81 w=0.64 l=0.15
X992 a_10479_8190# a_9967_7798# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X993 hgu_sarlogic_flat_0.x2.x2.x4.x2.floating sample_delay_cap_ctrl_code[0] hgu_sarlogic_flat_0.x2.x2.x4.x9.output_stack VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.124 ps=1.43 w=0.42 l=0.15
X994 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_0.d<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X995 a_11830_1153# a_11084_1179# a_11966_1179# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X996 a_16448_15176# hgu_sarlogic_flat_0.x2.x2.x1.x9.output_stack hgu_sarlogic_flat_0.x2.x2.x2.IN VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.122 ps=1.42 w=0.42 l=0.15
X997 hgu_cdac_half_1.VREF hgu_cdac_half_1.db<6> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X998 VSS a_2036_7824# hgu_sarlogic_flat_0.x3.x4.X VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X999 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1000 hgu_sarlogic_flat_0.x4.x9.X a_2786_2883# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.158 ps=1.39 w=1 l=0.15
X1001 hgu_sarlogic_flat_0.x3.x4.A a_1422_7824# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1002 hgu_sarlogic_flat_0.x4.x9.A1 a_3960_3698# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1003 a_n638_n245# hgu_cdac_sw_buffer_0.x3.A VSS VSS sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1004 hgu_cdac_half_0.db<6> a_n1158_n1744# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1005 hgu_vgen_vref_0.vcm hgu_vgen_vref_0.phi1_n hgu_vgen_vref_0.mimtop1 hgu_tah_0.VDD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=0.5
X1006 a_16799_6912# a_16287_6564# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X1007 a_11275_1461# a_11084_1179# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X1008 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<15:0> hgu_cdac_half_0.d<4> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1009 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.d<6> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1010 hgu_sarlogic_flat_0.x2.x3.Y VSS a_2323_10792# VDD sky130_fd_pr__pfet_01v8 ad=0.551 pd=4.38 as=0.551 ps=4.38 w=1.9 l=0.15
X1011 VDD a_n7390_7871# a_n7766_6446# VDD sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.3 as=0.139 ps=1.17 w=0.84 l=0.15
X1012 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X1013 VDD a_n4397_8367# hgu_cdac_sw_buffer_3.x11.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1014 VSS a_n6292_6446# hgu_comp_flat_0.comp_outn VSS sky130_fd_pr__nfet_01v8 ad=0.0759 pd=0.79 as=0.0759 ps=0.79 w=0.46 l=0.15
X1015 a_1716_n241# hgu_cdac_sw_buffer_1.x3.A VSS VSS sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1016 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.db<6> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1017 VSS a_7772_8487# a_7707_8513# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X1018 VSS a_n148_n1104# hgu_cdac_half_0.db<4> VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1019 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<7:0> hgu_cdac_half_0.db<3> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1020 VSS hgu_cdac_half_0.db<6> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1021 a_6817_8879# a_6370_8513# a_6724_8513# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X1022 a_16113_11849# hgu_sarlogic_flat_0.x2.x2.x2.IN a_16041_11987# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X1023 a_3309_9708# hgu_sarlogic_flat_0.x4.x15.S VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=0.995 as=0.154 ps=1.34 w=0.64 l=0.15
X1024 a_1502_2234# a_1056_1868# a_1410_1868# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0651 ps=0.73 w=0.42 l=0.15
X1025 a_11132_2883# hgu_sarlogic_flat_0.x4.x9.A1 a_10673_2708# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X1026 hgu_sarlogic_flat_0.x2.x2.x3.x7.floating sample_delay_offset hgu_sarlogic_flat_0.x2.x2.x3.x9.output_stack VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X1027 VDD a_n2219_8368# hgu_cdac_half_1.d<6> VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1028 hgu_vgen_vref_0.mimtop2 VSS sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X1029 VDD VDD a_1203_1153# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0956 pd=0.875 as=0.132 ps=1.22 w=0.42 l=0.15
X1030 a_n54567_7835# a_n54471_7657# hgu_tah_0.VDD hgu_tah_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.141 ps=1.33 w=0.42 l=0.15
X1031 a_n55204_7835# hgu_vgen_vref_0.sky130_fd_sc_hd__dlymetal6s6s_1_3.A VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1032 a_7842_6262# a_7370_6052# a_8086_6444# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X1033 hgu_cdac_sw_buffer_0.x11.A a_n1240_n1104# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1034 a_9464_7798# a_9763_7798# a_9698_7824# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.066 ps=0.745 w=0.36 l=0.15
X1035 a_1418_14758# a_1137_14764# a_1325_14758# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X1036 VSS a_11102_2530# a_11036_2556# VSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X1037 a_n7660_7467# hgu_comp_flat_0.clk VSS VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.165 ps=1.33 w=1 l=0.15
X1038 a_11625_1453# hgu_sarlogic_flat_0.x4.x17.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1039 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.db<6> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1040 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1041 hgu_tah_0.tah_vp hgu_tah_0.sw vip VSS sky130_fd_pr__nfet_01v8 ad=0.454 pd=3.08 as=0.454 ps=3.08 w=2.75 l=0.15
X1042 a_14654_8215# hgu_sarlogic_flat_0.x5.eob a_14566_8077# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X1043 a_7234_7233# a_6816_7317# a_6990_6925# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X1044 a_7887_6951# hgu_sarlogic_flat_0.x3.x45.Q_N VSS VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X1045 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1046 VDD hgu_sarlogic_flat_0.x4.x17.S a_12566_2883# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.0767 ps=0.785 w=0.42 l=0.15
X1047 VDD hgu_sarlogic_flat_0.x4.x13.S a_13073_7824# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0662 ps=0.735 w=0.42 l=0.15
X1048 a_4424_7317# a_4143_6951# a_4331_6951# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X1049 VDD a_1732_6052# hgu_sarlogic_flat_0.x3.x51.Q_N VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X1050 VSS a_n688_n1104# hgu_cdac_half_0.db<5> VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1051 hgu_vgen_vref_0.mimtop2 hgu_vgen_vref_0.phi1 hgu_vgen_vref_0.vcm VSS sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=0.5
X1052 a_2544_n241# hgu_cdac_sw_buffer_1.x6.A VSS VSS sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1053 hgu_cdac_half_0.VREF hgu_cdac_half_0.d<6> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1054 VDD a_10771_1153# hgu_sarlogic_flat_0.x4.x32.Q_N VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X1055 VDD hgu_sarlogic_flat_0.x3.x5.A a_1863_9386# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1056 hgu_sarlogic_flat_0.x5.x1[0].Q_N a_17068_6564# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X1057 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1058 VSS hgu_sarlogic_flat_0.x4.x17.S a_12573_2556# VSS sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.0693 ps=0.75 w=0.42 l=0.15
X1059 a_7235_8795# a_6817_8879# a_6991_8487# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X1060 a_12090_7824# a_11301_7798# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0588 ps=0.7 w=0.42 l=0.15
X1061 a_4425_8879# a_4144_8513# a_4332_8513# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X1062 hgu_sarlogic_flat_0.x4.x13.S a_13263_8513# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X1063 hgu_cdac_sw_buffer_2.x11.A a_n2301_7728# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1064 hgu_cdac_half_1.db<4> a_n3387_7727# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1065 hgu_cdac_sw_buffer_2.x9.A a_773_1868# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X1066 a_2057_14758# a_1592_14732# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X1067 VSS hgu_cdac_half_1.d<5> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1068 hgu_cdac_half_0.VREF hgu_cdac_half_0.db<4> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<15:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1069 a_13072_6078# a_12153_6352# a_12626_6262# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X1070 VSS hgu_cdac_half_0.db<5> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1071 a_9404_12125# hgu_sarlogic_flat_0.x2.x2.x3.IN a_9332_12263# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X1072 hgu_sarlogic_flat_0.x3.x4.X a_2036_7824# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1073 VSS hgu_tah_0.sw_n a_1146_7824# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1074 VDD VDD a_18973_6790# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X1075 a_9760_1868# hgu_sarlogic_flat_0.x4.x2.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.03 as=0.0703 ps=0.755 w=0.42 l=0.15
X1076 a_20464_8538# hgu_sarlogic_flat_0.x5.x2.x9.output_stack VSS VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X1077 VDD hgu_sarlogic_flat_0.x4.x30.A a_3960_3698# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1078 VSS a_n424_3698# hgu_sarlogic_flat_0.x4.x2.X VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1079 a_4144_8513# a_3978_8513# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1080 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_1.d<5> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1081 hgu_cdac_half_1.VREF hgu_cdac_half_1.db<5> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1082 a_1161_10641# hgu_tah_0.sw VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X1083 hgu_tah_0.VDD a_n55204_7371# a_n55391_7113# hgu_tah_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X1084 hgu_cdac_half_0.d<5> a_1666_n1100# hgu_cdac_sw_buffer_1.VDD hgu_cdac_sw_buffer_1.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1085 a_n982_1868# hgu_sarlogic_flat_0.x4.x5.D VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X1086 hgu_tah_0.VDD VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X1087 hgu_cdac_half_1.VREF hgu_cdac_half_1.db<5> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1088 hgu_vgen_vref_0.mimbot1 hgu_vgen_vref_0.phi1_n VSS hgu_tah_0.VDD sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=0.5
X1089 a_2701_2150# a_2285_2234# a_2444_2136# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.132 ps=1.22 w=0.84 l=0.15
X1090 a_12566_2883# VSS a_12352_2883# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.193 ps=1.34 w=0.42 l=0.15
X1091 a_1123_11726# a_611_11594# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.084 ps=0.82 w=0.42 l=0.15
X1092 hgu_sarlogic_flat_0.x2.x2.x2.x9.output_stack hgu_sarlogic_flat_0.x2.x2.x2.x10.Y hgu_sarlogic_flat_0.x2.x2.x2.x5[7].floating VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X1093 a_5182_6052# a_5450_6262# a_5396_6360# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X1094 a_8281_2708# VSS a_8423_2883# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X1095 hgu_sarlogic_flat_0.x3.x27.D a_3695_8513# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X1096 hgu_cdac_half_1.d<6> a_n2219_8368# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1097 VSS a_2036_7824# hgu_sarlogic_flat_0.x3.x4.X VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1098 VDD hgu_sarlogic_flat_0.x3.x7.X a_3504_6078# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0662 ps=0.735 w=0.42 l=0.15
X1099 a_9221_6078# hgu_sarlogic_flat_0.x3.x4.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.154 ps=1.34 w=0.64 l=0.15
X1100 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.db<6> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1101 hgu_tah_0.VDD a_n54752_8227# hgu_vgen_vref_0.phi1_n hgu_tah_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1102 a_n53010_7683# hgu_vgen_vref_0.sky130_fd_sc_hd__inv_1_3.Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1103 VSS a_7370_6052# a_7369_6352# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1104 VSS hgu_cdac_half_0.d<6> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1105 a_9950_1179# a_9438_1153# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0882 ps=0.84 w=0.42 l=0.15
X1106 a_18589_5036# a_18058_4670# a_18505_5036# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X1107 VSS hgu_vgen_vref_0.phi1 hgu_vgen_vref_0.mimbot1 VSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=0.5
X1108 a_14726_7939# hgu_sarlogic_flat_0.x5.eob a_14654_7939# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X1109 VSS a_n424_3698# hgu_sarlogic_flat_0.x4.x2.X VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1110 VSS a_5891_1331# hgu_cdac_sw_buffer_3.x6.A VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X1111 VDD a_n4397_8367# hgu_cdac_sw_buffer_3.x11.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1112 a_17302_6232# a_16894_5950# a_17068_5924# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X1113 VSS hgu_cdac_half_1.db<4> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<15:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1114 hgu_cdac_sw_buffer_1.x11.A a_1114_n1100# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1115 a_14222_1153# a_14490_1363# a_14436_1461# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X1116 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1117 hgu_tah_0.VDD a_n54752_6595# hgu_vgen_vref_0.phi2_n hgu_tah_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1118 hgu_cdac_half_1.VREF hgu_cdac_half_1.d<6> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1119 VDD hgu_sarlogic_flat_0.x2.x2.x3.x9.output_stack a_3314_11461# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X1120 VDD hgu_sarlogic_flat_0.x4.x20.S a_14492_2883# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.118 ps=1.4 w=0.42 l=0.15
X1121 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<15:0> hgu_cdac_half_1.db<4> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1122 hgu_cdac_half_1.VREF hgu_cdac_half_1.db<6> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1123 hgu_tah_0.tah_vn hgu_tah_0.sw hgu_tah_0.tah_vn hgu_tah_0.VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.908 ps=5.83 w=5.5 l=0.15
X1124 VSS hgu_cdac_half_0.d<5> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1125 VSS hgu_cdac_half_0.db<6> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1126 a_5110_6951# a_4598_6925# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X1127 a_16287_4644# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X1128 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_0.d<5> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1129 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.d<6> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1130 hgu_vgen_vref_0.phi1_n a_n54752_8227# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1131 a_2141_2150# a_1676_1842# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X1132 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_1.db<5> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1133 a_19144_5310# a_18679_5284# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X1134 VDD hgu_sarlogic_flat_0.x4.D[2] a_12543_1179# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X1135 VSS hgu_sarlogic_flat_0.x4.x20.S a_14492_2883# VSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.109 ps=1.36 w=0.42 l=0.15
X1136 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.db<6> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1137 a_8423_2883# hgu_sarlogic_flat_0.x4.x15.S VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X1138 a_3954_15763# hgu_sarlogic_flat_0.x2.x3.A a_3866_15625# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X1139 VSS hgu_comp_flat_0.clk a_3050_3698# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1140 VDD a_13494_2530# a_13524_2883# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1141 a_9379_10598# hgu_sarlogic_flat_0.x2.x2.x3.IN a_9291_10460# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X1142 VDD a_n2301_7728# hgu_cdac_sw_buffer_2.x11.A VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1143 hgu_sarlogic_flat_0.x2.x2.x4.x10.Y sample_delay_cap_ctrl_code[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1144 hgu_sarlogic_flat_0.x4.x9.A1 a_3960_3698# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1145 a_4212_1868# a_4362_1842# a_4068_1842# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1146 hgu_cdac_half_1.VREF hgu_cdac_half_1.db<6> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1147 a_5450_6262# a_4978_6052# a_5694_6444# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X1148 a_16531_4952# a_16113_5036# a_16287_4644# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X1149 a_2786_2883# hgu_sarlogic_flat_0.x4.x9.A1 a_2714_2883# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X1150 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<15:0> hgu_cdac_half_0.db<4> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1151 a_8423_2556# hgu_sarlogic_flat_0.x4.x15.S VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X1152 hgu_sarlogic_flat_0.x2.x2.x1.x9.output_stack sample_delay_offset hgu_sarlogic_flat_0.x2.x2.x1.x7.floating VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X1153 VDD hgu_comp_flat_0.comp_outp a_1178_6950# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1154 a_11300_6052# a_11855_6052# a_11813_6360# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0882 ps=1.05 w=0.84 l=0.15
X1155 VDD a_19460_5284# a_20167_5326# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X1156 VSS hgu_cdac_half_1.d<2> hgu_cdac_half_1.hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT VSS sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.35
X1157 a_5063_7233# a_4598_6925# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X1158 VSS hgu_cdac_half_1.d<6> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1159 VSS VDD a_18973_5924# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1160 a_3929_14098# hgu_sarlogic_flat_0.x2.x3.A a_3841_14098# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X1161 a_4842_7233# a_4424_7317# a_4598_6925# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X1162 VSS a_7771_6925# a_8478_6951# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1163 hgu_sarlogic_flat_0.x1.x2.x5[7].floating hgu_sarlogic_flat_0.x1.x2.x10.Y hgu_sarlogic_flat_0.x1.x2.x9.output_stack VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X1164 VDD hgu_sarlogic_flat_0.x4.x15.S a_10681_7824# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0662 ps=0.735 w=0.42 l=0.15
X1165 hgu_comp_flat_0.Q hgu_tah_0.tah_vn a_n7660_7467# VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1166 a_2786_2556# a_2532_2883# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.145 ps=1.11 w=0.42 l=0.15
X1167 VSS hgu_cdac_sw_buffer_2.x11.A a_n2219_8368# VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1168 VSS VDD a_18973_6790# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1169 hgu_vgen_vref_0.mimtop1 hgu_vgen_vref_0.mimbot1 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X1170 hgu_sarlogic_flat_0.x2.x2.x2.x9.output_stack sample_delay_cap_ctrl_code[8] hgu_sarlogic_flat_0.x2.x2.x2.x2.floating VSS sky130_fd_pr__nfet_01v8 ad=0.124 pd=1.43 as=0.122 ps=1.42 w=0.42 l=0.15
X1171 a_5064_8795# a_4599_8487# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X1172 a_16197_5310# a_15666_5316# a_16113_5310# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X1173 VSS hgu_cdac_half_0.d<6> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1174 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.d<6> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1175 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1176 a_4843_8795# a_4425_8879# a_4599_8487# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X1177 a_n54567_7371# a_n54471_7113# hgu_tah_0.VDD hgu_tah_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.141 ps=1.33 w=0.42 l=0.15
X1178 VDD a_1105_2708# hgu_sarlogic_flat_0.x4.x8.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X1179 hgu_cdac_half_0.VREF hgu_cdac_half_0.db<4> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<15:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.35
X1180 VSS hgu_cdac_half_0.db<3> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<7:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1181 VSS a_2323_10792# a_1945_10648# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X1182 a_6_1179# a_138_1363# a_n130_1153# VSS sky130_fd_pr__nfet_01v8 ad=0.0974 pd=0.97 as=0.0864 ps=0.91 w=0.64 l=0.15
X1183 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1184 a_16197_6316# a_15666_5950# a_16113_6316# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X1185 VSS a_n55204_7835# a_n55391_7657# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X1186 a_10680_6078# a_9761_6352# a_10234_6262# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X1187 hgu_sarlogic_flat_0.x2.x2.x1.x3[1].floating sample_delay_cap_ctrl_code[5] hgu_sarlogic_flat_0.x2.x2.x1.x9.output_stack VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X1188 VDD hgu_tah_0.sw_n a_n1334_3698# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1189 a_8283_1331# a_8379_1153# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X1190 a_12269_2150# a_11853_2234# a_12012_2136# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.132 ps=1.22 w=0.84 l=0.15
X1191 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X1192 a_n638_n245# hgu_cdac_sw_buffer_0.x3.A hgu_cdac_sw_buffer_0.VDD hgu_cdac_sw_buffer_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1193 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_1.d<5> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1194 a_1752_8513# a_1586_8513# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1195 VSS hgu_cdac_half_1.db<6> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1196 a_16041_12815# hgu_sarlogic_flat_0.x2.x2.x2.IN VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X1197 VSS a_6421_6052# hgu_sarlogic_flat_0.x4.D[5] VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X1198 a_18819_4670# a_18973_4644# a_18679_4644# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1199 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<15:0> hgu_cdac_half_1.db<4> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1200 a_5379_6925# a_5205_6951# a_5495_6951# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X1201 a_n3325_7252# hgu_cdac_sw_buffer_3.x4.A VSS VSS sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1202 a_1418_14758# a_971_14764# a_1325_14758# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X1203 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.db<6> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1204 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.db<6> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1205 VDD hgu_cdac_sw_buffer_3.x11.A a_n4397_8367# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1206 hgu_cdac_half_1.VREF hgu_cdac_half_1.d<5> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1207 a_9404_12401# hgu_sarlogic_flat_0.x2.x2.x3.IN a_9332_12539# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X1208 hgu_cdac_half_0.db<6> a_n1158_n1744# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1209 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_1.db<5> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1210 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1211 a_12627_8008# a_12155_7798# a_12871_8190# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X1212 a_1382_10641# hgu_sarlogic_flat_0.x1.x3.A0 a_1019_10793# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X1213 a_19372_6590# a_18224_6596# a_19286_6968# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X1214 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1215 a_466_n245# hgu_cdac_sw_buffer_0.x5.A VSS VSS sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1216 hgu_sarlogic_flat_0.x4.x15.X a_9962_2883# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.158 ps=1.39 w=1 l=0.15
X1217 VDD a_6841_1453# a_6842_1153# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1218 a_3302_6078# a_2790_6052# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.084 ps=0.82 w=0.42 l=0.15
X1219 hgu_cdac_half_0.VREF hgu_cdac_half_0.d<6> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1220 VSS a_1019_10793# hgu_sarlogic_flat_0.x1.x3.X VSS sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X1221 a_18412_5310# hgu_sarlogic_flat_0.x4.D[5] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X1222 VSS hgu_sarlogic_flat_0.x4.x8.X a_1056_1868# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1223 VSS a_n1158_n1744# hgu_cdac_half_0.db<6> VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1224 hgu_vgen_vref_0.mimtop2 VSS sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X1225 hgu_cdac_half_0.VREF hgu_cdac_half_0.db<5> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1226 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_1.d<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1227 a_18412_5950# hgu_sarlogic_flat_0.x4.D[3] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X1228 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<1:0> hgu_cdac_half_0.d<1> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.122 ps=1.42 w=0.42 l=0.35
X1229 a_10279_6951# a_9676_6925# a_10163_6925# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1230 a_3504_6078# a_2586_6052# a_3058_6262# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1231 VDD a_7046_1153# a_6979_1545# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X1232 VSS a_1863_9386# hgu_sarlogic_flat_0.x3.x5.X VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1233 a_n53930_7371# a_n53834_7113# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1234 hgu_cdac_sw_buffer_3.x8.X a_n4203_7087# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1235 hgu_cdac_sw_buffer_2.x12.X a_n1473_7088# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1236 a_19576_4670# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X1237 VSS hgu_cdac_half_1.d<4> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<15:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1238 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.d<6> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1239 a_16113_5036# a_15832_4670# a_16020_4670# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X1240 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.db<6> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1241 a_16752_5310# a_16287_5284# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X1242 VSS hgu_cdac_half_1.d<5> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1243 a_19576_5676# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X1244 hgu_cdac_half_0.VREF hgu_cdac_half_0.d<5> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1245 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.db<6> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1246 hgu_sarlogic_flat_0.x3.x7.X a_1454_6950# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1247 a_19576_4670# a_18973_4644# a_19460_4644# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1248 VSS a_n1240_n1104# hgu_cdac_sw_buffer_0.x11.A VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1249 hgu_sarlogic_flat_0.x1.x4.x9.output_stack hgu_comp_flat_0.clk a_n6959_11861# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X1250 VDD a_7771_6925# a_8478_6951# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X1251 hgu_cdac_half_1.VREF hgu_cdac_half_1.db<1> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<1:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.35
X1252 hgu_sarlogic_flat_0.x2.x2.x3.x6.floating hgu_sarlogic_flat_0.x2.x2.x3.x6.SW hgu_sarlogic_flat_0.x2.x2.x3.x9.output_stack VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X1253 a_11814_8106# a_11614_7824# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X1254 VDD hgu_sarlogic_flat_0.x4.x3.X a_n424_3698# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1255 VDD hgu_sarlogic_flat_0.x2.x2.x3.IN a_10023_11664# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1256 result[2] a_17775_5950# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X1257 a_n643_1347# a_n335_1453# a_n386_1545# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0787 ps=0.795 w=0.42 l=0.15
X1258 a_n55487_7371# a_n55391_7113# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1259 hgu_cdac_sw_buffer_1.VDD a_1196_n1740# hgu_cdac_half_0.d<6> hgu_cdac_sw_buffer_1.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1260 hgu_vgen_vref_0.mimtop1 hgu_vgen_vref_0.mimbot1 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X1261 VSS VDD a_4790_1179# VSS sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0974 ps=0.97 w=0.42 l=0.15
X1262 a_9545_2234# a_8232_1868# a_9461_2234# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0787 pd=0.795 as=0.0567 ps=0.69 w=0.42 l=0.15
X1263 a_1820_1868# a_1970_1842# a_1676_1842# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1264 hgu_tah_0.VDD hgu_vgen_vref_0.sky130_fd_sc_hd__inv_1_2.A a_n55304_8227# hgu_tah_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1265 VSS VDD a_10103_7824# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.101 ps=0.99 w=0.42 l=0.15
X1266 hgu_sarlogic_flat_0.x4.x2.X a_n424_3698# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1267 a_n542_11334# a_n447_11350# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1268 VSS hgu_comp_flat_0.comp_outp a_1178_6950# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1269 a_7788_6360# a_6829_6078# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X1270 hgu_sarlogic_flat_0.x4.x2.X a_n424_3698# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1271 hgu_vgen_vref_0.mimtop1 hgu_vgen_vref_0.mimbot1 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X1272 a_16427_4670# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X1273 a_9327_6078# a_9463_6052# a_8908_6052# VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0864 ps=0.91 w=0.64 l=0.15
X1274 a_12543_1179# a_11626_1153# a_12098_1363# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0675 ps=0.735 w=0.36 l=0.15
X1275 a_20464_8879# hgu_sarlogic_flat_0.x5.x2.x9.output_stack hgu_sarlogic_flat_0.x5.x3.A VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.122 ps=1.42 w=0.42 l=0.15
X1276 a_16427_5950# a_16581_5924# a_16287_5924# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1277 a_1105_2708# hgu_sarlogic_flat_0.x4.x9.A1 a_1247_2556# VSS sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X1278 a_n54567_7835# a_n54471_7657# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1279 a_n2251_7253# hgu_cdac_sw_buffer_2.x9.A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1280 hgu_tah_0.VDD a_n55304_6595# hgu_vgen_vref_0.phi2 hgu_tah_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1281 VDD hgu_sarlogic_flat_0.x3.x4.X a_7284_6925# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X1282 a_16427_5676# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X1283 a_6194_1868# hgu_sarlogic_flat_0.x4.D[4] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X1284 hgu_tah_0.tah_vp hgu_tah_0.sw_n vip hgu_tah_0.VDD sky130_fd_pr__pfet_01v8 ad=0.908 pd=5.83 as=0.908 ps=5.83 w=5.5 l=0.15
X1285 a_n858_2530# hgu_sarlogic_flat_0.x4.x7.S VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X1286 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1287 hgu_cdac_half_0.VREF hgu_cdac_half_0.db<6> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1288 a_2672_8795# a_2207_8487# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X1289 VDD hgu_sarlogic_flat_0.x4.x8.X a_1056_1868# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1290 a_10710_14512# hgu_sarlogic_flat_0.x2.x2.x1.IN a_10638_14512# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X1291 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1292 a_3378_9360# sel_bit[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1293 hgu_sarlogic_flat_0.x3.x4.X a_2036_7824# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1294 a_11561_1179# a_10771_1153# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0703 ps=0.755 w=0.42 l=0.15
X1295 hgu_sarlogic_flat_0.x1.x4.x9.output_stack async_resetb_delay_cap_ctrl_code[1] hgu_sarlogic_flat_0.x1.x4.x3[1].floating VSS sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X1296 a_7759_1179# a_6841_1453# a_7314_1363# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.0567 ps=0.69 w=0.42 l=0.15
X1297 VDD hgu_sarlogic_flat_0.x3.x4.X a_7285_8487# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X1298 hgu_vgen_vref_0.phi1 a_n55304_8227# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1299 hgu_sarlogic_flat_0.x4.x27.A a_3050_3698# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1300 hgu_cdac_half_0.VREF hgu_cdac_half_0.d<6> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1301 a_n858_2530# hgu_sarlogic_flat_0.x4.x7.S VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X1302 a_n876_1179# hgu_sarlogic_flat_0.x4.x2.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.17 pd=1.81 as=0.154 ps=1.34 w=0.64 l=0.15
X1303 VDD hgu_sarlogic_flat_0.x3.x33.Q_N a_9966_6052# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X1304 a_5891_1331# a_5987_1153# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X1305 a_12358_6052# a_12626_6262# a_12572_6360# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X1306 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.d<6> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1307 VSS a_n3387_7727# hgu_cdac_half_1.db<4> VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1308 VSS a_1196_n1740# hgu_cdac_half_0.d<6> VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1309 VSS a_n55770_7371# hgu_vgen_vref_0.sky130_fd_sc_hd__inv_1_1.A VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X1310 a_5897_7824# a_4978_8098# a_5451_8008# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X1311 VDD a_14404_2136# a_15125_1868# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X1312 a_9989_6951# a_8927_6951# a_9894_6951# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X1313 VSS hgu_sarlogic_flat_0.x4.D[1] a_14935_1179# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1314 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.d<6> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1315 a_10638_14374# hgu_sarlogic_flat_0.x2.x2.x1.IN a_10550_14374# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X1316 VSS hgu_cdac_half_1.db<5> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1317 a_2808_n935# VSS hgu_cdac_sw_buffer_1.VDD hgu_cdac_sw_buffer_1.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1318 a_8087_7824# a_7575_7798# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.084 ps=0.82 w=0.42 l=0.15
X1319 VDD hgu_sarlogic_flat_0.x5.x3.X a_18058_6596# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1320 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1321 a_17184_5950# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X1322 a_n6934_15288# hgu_comp_flat_0.ready a_n7022_15150# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X1323 hgu_cdac_half_1.VREF hgu_cdac_half_1.db<6> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1324 hgu_cdac_half_1.VREF hgu_cdac_half_1.d<6> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1325 VSS a_2036_7824# hgu_sarlogic_flat_0.x3.x4.X VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1326 a_8289_7824# a_7371_7798# a_7843_8008# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1327 hgu_cdac_half_1.db<5> a_n3927_7727# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1328 a_17184_6956# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X1329 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<15:0> hgu_cdac_half_0.db<4> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1330 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X1331 hgu_cdac_half_1.VREF hgu_cdac_half_1.db<6> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1332 a_17184_5950# a_16581_5924# a_17068_5924# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1333 VSS hgu_cdac_sw_buffer_1.x9.X a_1114_n1100# VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1334 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<7:0> hgu_cdac_half_1.db<3> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1335 hgu_cdac_half_1.d<6> a_n2219_8368# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1336 a_16980_6590# a_15832_6596# a_16894_6968# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X1337 VDD a_4449_1453# a_4450_1153# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1338 VDD a_13930_1842# a_14661_2150# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X1339 a_9233_1453# hgu_sarlogic_flat_0.x4.x15.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1340 hgu_cdac_half_0.VREF hgu_cdac_half_0.db<5> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1341 a_n6959_14037# hgu_comp_flat_0.ready a_n7047_13899# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X1342 a_12286_6951# a_11774_6925# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X1343 hgu_sarlogic_flat_0.x2.x3.Y hgu_sarlogic_flat_0.x2.x3.A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1344 a_16020_5310# hgu_sarlogic_flat_0.x4.D[4] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X1345 result[4] a_17775_5326# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X1346 VSS hgu_cdac_half_0.d<4> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<15:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1347 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X1348 VDD hgu_sarlogic_flat_0.x4.x13.S a_7784_2883# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.0767 ps=0.785 w=0.42 l=0.15
X1349 VDD a_n2219_8368# hgu_cdac_half_1.d<6> VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1350 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.d<6> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1351 hgu_sarlogic_flat_0.x2.x2.x3.x4[3].floating sample_delay_cap_ctrl_code[14] hgu_sarlogic_flat_0.x2.x2.x3.x9.output_stack VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X1352 VSS a_9966_6052# a_9901_6078# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0935 ps=0.965 w=0.64 l=0.15
X1353 a_16020_5950# hgu_sarlogic_flat_0.x4.D[2] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X1354 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X1355 VSS a_n55304_6595# hgu_vgen_vref_0.phi2 VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1356 hgu_cdac_sw_buffer_1.VDD a_2820_n241# hgu_cdac_half_0.d<2> hgu_cdac_sw_buffer_1.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1357 a_546_11738# a_406_11482# a_108_11334# VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.0711 ps=0.755 w=0.36 l=0.15
X1358 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X1359 VSS hgu_cdac_half_1.d<4> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<15:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.35
X1360 a_11774_6925# a_11600_7317# a_11914_6951# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X1361 hgu_sarlogic_flat_0.x4.x2.X a_n424_3698# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1362 VSS hgu_sarlogic_flat_0.x4.x13.S a_7791_2556# VSS sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.0693 ps=0.75 w=0.42 l=0.15
X1363 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<0> hgu_cdac_half_1.d<0> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.35
X1364 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1365 a_4173_9684# hgu_sarlogic_flat_0.x3.x48.Q VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.164 pd=1.33 as=0.0864 ps=0.91 w=0.64 l=0.15
X1366 a_16221_4670# a_15832_4670# a_16113_5036# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X1367 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<1:0> hgu_cdac_half_0.d<1> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.35
X1368 a_11388_1868# a_11538_1842# a_11244_1842# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1369 hgu_sarlogic_flat_0.x5.x2.x10.Y retimer_delay_code[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1370 hgu_sarlogic_flat_0.x5.x2.x9.output_stack retimer_delay_code[2] hgu_sarlogic_flat_0.x5.x2.x4[3].floating VSS sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X1371 a_12239_7233# a_11774_6925# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X1372 a_7510_7824# a_7370_8098# a_7072_7798# VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.0711 ps=0.755 w=0.36 l=0.15
X1373 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<15:0> hgu_cdac_half_1.d<4> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1374 VSS a_6841_1453# a_6842_1153# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1375 a_12293_6078# a_12153_6352# a_11855_6052# VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.0711 ps=0.755 w=0.36 l=0.15
X1376 hgu_sarlogic_flat_0.x4.x34.Q_N a_14404_2136# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X1377 a_11708_6951# a_11319_6951# a_11600_7317# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X1378 a_342_11726# a_n447_11350# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0588 ps=0.7 w=0.42 l=0.15
X1379 VSS VDD a_2398_1179# VSS sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0974 ps=0.97 w=0.42 l=0.15
X1380 hgu_sarlogic_flat_0.x4.x28.Q_N a_9620_2136# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X1381 VSS hgu_comp_flat_0.clk a_n7660_7467# VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.31 ps=2.62 w=1 l=0.15
X1382 VDD VDD a_16581_4644# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X1383 hgu_cdac_half_1.db<4> a_n3387_7727# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1384 VDD a_16287_6564# a_16197_6590# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X1385 a_1732_6052# a_2287_6052# a_2245_6360# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0882 ps=1.05 w=0.84 l=0.15
X1386 a_2808_n935# VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1387 a_7784_2883# VSS a_7570_2883# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.193 ps=1.34 w=0.42 l=0.15
X1388 hgu_cdac_half_1.VREF hgu_cdac_half_1.d<5> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1389 hgu_vgen_vref_0.mimtop2 VSS sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X1390 hgu_cdac_half_0.hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT hgu_cdac_half_0.db<2> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.122 ps=1.42 w=0.42 l=0.35
X1391 a_n53364_7835# hgu_vgen_vref_0.sky130_fd_sc_hd__nand2_1_0.Y hgu_tah_0.VDD hgu_tah_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.141 ps=1.33 w=0.42 l=0.15
X1392 a_2287_6052# a_2586_6052# a_2521_6078# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.066 ps=0.745 w=0.36 l=0.15
X1393 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<15:0> hgu_cdac_half_0.d<4> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1394 a_n6292_6446# hgu_comp_flat_0.RS_n VDD VDD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0.244 ps=2.26 w=0.84 l=0.15
X1395 a_18613_5688# a_18224_5316# a_18505_5310# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X1396 hgu_cdac_half_0.VREF hgu_cdac_half_0.db<6> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1397 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_1.db<5> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1398 VDD hgu_sarlogic_flat_0.x3.x4.X a_4892_6925# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X1399 a_n7678_6446# a_n7760_6349# a_n7766_6446# VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.15
X1400 VDD a_4978_6052# a_4977_6352# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1401 a_6421_6052# a_6516_6052# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X1402 a_3595_1153# a_4141_1347# a_4099_1461# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.132 pd=1.22 as=0.0882 ps=1.05 w=0.84 l=0.15
X1403 a_7228_2136# a_7069_2234# a_7368_1868# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.109 ps=1.03 w=0.64 l=0.15
X1404 a_17068_4644# a_16894_4670# a_17184_4670# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X1405 a_3802_1868# hgu_sarlogic_flat_0.x4.D[5] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X1406 a_466_n245# hgu_cdac_sw_buffer_0.x5.A hgu_cdac_sw_buffer_0.VDD hgu_cdac_sw_buffer_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1407 VSS sample_delay_offset hgu_sarlogic_flat_0.x2.x2.x4.x6.SW VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1408 a_1836_14758# a_1418_14758# a_1592_14732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X1409 VSS a_8814_7798# hgu_sarlogic_flat_0.x4.x17.S VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X1410 VSS hgu_cdac_half_0.d<6> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1411 hgu_cdac_half_0.d<5> a_1666_n1100# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1412 a_n1170_1868# a_n1336_1868# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1413 a_n424_3698# hgu_sarlogic_flat_0.x4.x3.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1414 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.d<6> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1415 VDD hgu_sarlogic_flat_0.x3.x4.X a_4893_8487# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X1416 VDD VDD a_7046_1153# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X1417 a_12555_6925# a_12381_6951# a_12671_6951# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X1418 VSS a_8379_1153# hgu_sarlogic_flat_0.x4.x29.Q_N VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X1419 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_1.d<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1420 a_9438_1153# a_9706_1363# a_9652_1461# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X1421 VDD a_18973_4644# a_19694_4952# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X1422 hgu_tah_0.VDD a_n54752_8227# hgu_vgen_vref_0.phi1_n hgu_tah_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1423 hgu_cdac_half_0.d<6> a_1196_n1740# hgu_cdac_sw_buffer_1.VDD hgu_cdac_sw_buffer_1.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1424 a_n2219_8368# hgu_cdac_sw_buffer_2.x11.A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1425 VSS VDD a_8798_1179# VSS sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.109 ps=1.03 w=0.42 l=0.15
X1426 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X1427 hgu_vgen_vref_0.mimtop1 hgu_vgen_vref_0.mimbot1 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X1428 VDD a_12012_2136# a_12733_1868# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X1429 VDD VDD a_5183_7798# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X1430 VSS hgu_cdac_half_1.d<5> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1431 a_2207_8487# hgu_sarlogic_flat_0.x3.x4.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X1432 hgu_sarlogic_flat_0.x5.x2.x5[7].floating hgu_sarlogic_flat_0.x5.x2.x10.Y hgu_sarlogic_flat_0.x5.x2.x9.output_stack VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X1433 VDD a_5182_6052# a_5115_6444# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X1434 a_9762_6052# hgu_sarlogic_flat_0.x4.D[3] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1435 a_12152_1868# a_11538_1842# a_12012_2136# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1436 a_5695_7824# a_5183_7798# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.084 ps=0.82 w=0.42 l=0.15
X1437 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_1.db<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1438 hgu_tah_0.VDD hgu_vgen_vref_0.phi2 hgu_vgen_vref_0.mimtop1 VSS sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=0.5
X1439 hgu_cdac_sw_buffer_2.x11.A a_n2301_7728# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1440 a_n2773_7252# hgu_cdac_sw_buffer_3.x5.A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1441 hgu_cdac_half_1.VREF hgu_cdac_half_1.d<6> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1442 a_10478_6078# a_9966_6052# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.084 ps=0.82 w=0.42 l=0.15
X1443 hgu_cdac_sw_buffer_1.VDD a_2206_n1100# hgu_cdac_half_0.d<4> hgu_cdac_sw_buffer_1.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1444 hgu_cdac_sw_buffer_1.VDD a_1196_n1740# hgu_cdac_half_0.d<6> hgu_cdac_sw_buffer_1.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1445 hgu_cdac_half_1.VREF hgu_cdac_half_1.db<6> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1446 a_7772_8487# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X1447 a_5897_7824# a_4979_7798# a_5451_8008# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1448 a_7710_6078# a_7842_6262# a_7574_6052# VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0864 ps=0.91 w=0.64 l=0.15
X1449 hgu_cdac_half_1.VREF hgu_cdac_half_1.db<5> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.35
X1450 a_10180_6360# a_9221_6078# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X1451 VDD a_14222_1153# a_14155_1545# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X1452 a_1478_10968# VSS a_1019_10793# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X1453 a_18679_5924# a_18505_6316# a_18819_5950# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X1454 VSS hgu_cdac_half_0.db<5> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1455 hgu_cdac_half_1.VREF hgu_cdac_half_1.db<3> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<7:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1456 a_n1189_1153# a_n876_1179# a_n770_1179# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1457 a_n54850_7835# a_n54754_7657# hgu_tah_0.VDD hgu_tah_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.141 ps=1.33 w=0.42 l=0.15
X1458 a_n1170_1868# a_n1336_1868# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1459 a_9895_8513# a_9383_8487# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X1460 a_n595_7253# hgu_cdac_sw_buffer_2.x5.A VSS VSS sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1461 vin hgu_tah_0.sw_n hgu_tah_0.tah_vn hgu_tah_0.VDD sky130_fd_pr__pfet_01v8 ad=0.908 pd=5.83 as=0.908 ps=5.83 w=5.5 l=0.15
X1462 a_7305_6444# a_6516_6052# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0819 ps=0.81 w=0.42 l=0.15
X1463 hgu_cdac_half_0.VREF hgu_cdac_half_0.d<4> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<15:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1464 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1465 a_16221_6968# a_15832_6596# a_16113_6590# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X1466 VDD hgu_sarlogic_flat_0.x4.x9.S a_2532_2883# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.118 ps=1.4 w=0.42 l=0.15
X1467 hgu_sarlogic_flat_0.x2.x2.x1.x10.Y sample_delay_cap_ctrl_code[7] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1468 a_13428_2556# VSS a_13065_2708# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X1469 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1470 hgu_cdac_half_0.hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT hgu_cdac_half_0.db<2> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1471 a_18412_5950# hgu_sarlogic_flat_0.x4.D[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X1472 a_7507_6444# a_7370_6052# a_7071_6052# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X1473 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.db<6> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1474 a_3954_16039# hgu_sarlogic_flat_0.x2.x3.A a_3866_15901# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X1475 VSS hgu_sarlogic_flat_0.x4.x17.S a_8289_7824# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1476 hgu_sarlogic_flat_0.x3.x77.Y hgu_sarlogic_flat_0.x5.eob VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1477 a_n130_1153# a_n876_1179# a_6_1179# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1478 hgu_cdac_half_0.d<6> a_1196_n1740# hgu_cdac_sw_buffer_1.VDD hgu_cdac_sw_buffer_1.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1479 a_n1285_1331# a_n1189_1153# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X1480 VDD VDD a_11538_1842# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.17 ps=1.81 w=0.64 l=0.15
X1481 a_18412_6590# hgu_sarlogic_flat_0.x4.D[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X1482 VSS hgu_sarlogic_flat_0.x3.x7.X a_13072_6078# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1483 hgu_cdac_sw_buffer_1.x8.X a_1390_n460# hgu_cdac_sw_buffer_1.VDD hgu_cdac_sw_buffer_1.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1484 a_6300_1179# hgu_sarlogic_flat_0.x4.x2.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.17 pd=1.81 as=0.154 ps=1.34 w=0.64 l=0.15
X1485 VSS hgu_sarlogic_flat_0.x4.x9.S a_2532_2883# VSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.109 ps=1.36 w=0.42 l=0.15
X1486 hgu_vgen_vref_0.mimtop2 hgu_vgen_vref_0.phi1_n hgu_vgen_vref_0.vcm hgu_tah_0.VDD sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=0.5
X1487 VSS a_4449_1453# a_4450_1153# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1488 a_9233_1453# hgu_sarlogic_flat_0.x4.x15.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1489 a_12381_6951# a_11319_6951# a_12286_6951# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X1490 hgu_sarlogic_flat_0.x5.x1[7].Q_N a_19460_4644# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X1491 VSS VDD a_4362_1842# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1492 hgu_cdac_half_1.VREF hgu_cdac_half_1.d<4> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<15:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1493 hgu_cdac_sw_buffer_3.x11.A a_n4479_7727# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1494 a_108_11334# a_407_11578# a_342_11726# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.066 ps=0.745 w=0.36 l=0.15
X1495 hgu_sarlogic_flat_0.x4.D[1] a_10870_6951# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X1496 hgu_sarlogic_flat_0.x2.x2.x4.x4[3].floating sample_delay_cap_ctrl_code[2] hgu_sarlogic_flat_0.x2.x2.x4.x9.output_stack VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X1497 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X1498 a_14404_2136# hgu_sarlogic_flat_0.x4.x2.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.132 pd=1.22 as=0.0956 ps=0.875 w=0.42 l=0.15
X1499 VSS hgu_cdac_half_0.d<6> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1500 a_2268_n241# hgu_cdac_sw_buffer_1.x4.A VSS VSS sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1501 hgu_cdac_half_0.VREF hgu_cdac_half_0.db<5> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1502 VDD hgu_sarlogic_flat_0.x3.x5.X a_1586_8513# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1503 a_n7660_7467# hgu_tah_0.tah_vn hgu_comp_flat_0.Q VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1504 hgu_sarlogic_flat_0.x5.x1[4].Q_N a_17068_5284# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X1505 a_14935_1179# a_14017_1453# a_14490_1363# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.0567 ps=0.69 w=0.42 l=0.15
X1506 VSS hgu_cdac_half_1.db<3> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<7:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1507 hgu_sarlogic_flat_0.x5.x2.x4[3].floating retimer_delay_code[2] hgu_sarlogic_flat_0.x5.x2.x9.output_stack VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X1508 VSS hgu_sarlogic_flat_0.x3.x4.X a_9676_6925# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1509 VDD a_2586_6052# a_2585_6352# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1510 VSS hgu_cdac_half_0.db<6> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1511 a_9464_7798# a_9762_8098# a_9698_8190# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0924 ps=0.86 w=0.42 l=0.15
X1512 VSS a_n424_3698# hgu_sarlogic_flat_0.x4.x2.X VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1513 VSS hgu_cdac_half_0.d<6> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1514 VSS hgu_cdac_half_0.db<6> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1515 VSS a_6460_1842# a_6394_1868# VSS sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0671 ps=0.75 w=0.42 l=0.15
X1516 VDD hgu_comp_flat_0.clk a_n7022_10334# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X1517 hgu_sarlogic_flat_0.x4.x11.S a_10871_8513# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X1518 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<15:0> hgu_cdac_half_0.d<4> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1519 VSS hgu_cdac_half_0.db<4> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<15:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1520 a_9461_2234# a_8232_1868# a_9364_1868# VSS sky130_fd_pr__nfet_01v8 ad=0.0486 pd=0.63 as=0.116 ps=1.09 w=0.36 l=0.15
X1521 a_7368_1868# hgu_sarlogic_flat_0.x4.x2.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.03 as=0.0703 ps=0.755 w=0.42 l=0.15
X1522 VDD hgu_cdac_sw_buffer_3.x11.A a_n4397_8367# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1523 hgu_cdac_sw_buffer_3.x11.X a_n4397_8367# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1524 hgu_cdac_half_0.d<6> a_1196_n1740# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1525 VSS hgu_cdac_half_0.d<5> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1526 a_6517_7798# a_7072_7798# a_7030_8106# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0882 ps=1.05 w=0.84 l=0.15
X1527 hgu_cdac_half_0.VREF hgu_cdac_half_0.d<6> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1528 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<7:0> hgu_cdac_half_1.d<3> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.122 ps=1.42 w=0.42 l=0.35
X1529 hgu_sarlogic_flat_0.x3.x5.X a_1863_9386# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1530 a_n53364_7371# hgu_vgen_vref_0.sky130_fd_sc_hd__nand2_1_1.Y hgu_tah_0.VDD hgu_tah_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.141 ps=1.33 w=0.42 l=0.15
X1531 a_20464_8538# hgu_sarlogic_flat_0.x5.x3.A VDD VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1532 VSS VDD a_6406_1179# VSS sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.109 ps=1.03 w=0.42 l=0.15
X1533 a_4564_1179# a_4449_1453# a_4141_1347# VSS sky130_fd_pr__nfet_01v8 ad=0.116 pd=1.09 as=0.0486 ps=0.63 w=0.36 l=0.15
X1534 hgu_sarlogic_flat_0.x2.x2.x3.x4[3].floating sample_delay_cap_ctrl_code[14] hgu_sarlogic_flat_0.x2.x2.x3.x9.output_stack VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X1535 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_0.db<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1536 VSS hgu_cdac_half_1.d<4> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<15:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1537 hgu_cdac_half_0.db<6> a_n1158_n1744# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1538 a_2790_6052# a_3058_6262# a_3004_6360# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X1539 a_16088_10322# hgu_sarlogic_flat_0.x2.x2.x2.IN VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X1540 VSS hgu_cdac_half_1.d<5> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.35
X1541 a_2033_8879# a_1752_8513# a_1940_8513# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X1542 hgu_sarlogic_flat_0.x3.x66.Q_N a_12555_6925# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X1543 VDD a_2790_6052# a_2723_6444# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X1544 VSS a_4978_6052# a_4977_6352# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1545 a_7558_1179# a_7046_1153# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0882 ps=0.84 w=0.42 l=0.15
X1546 a_16799_5950# a_16287_5924# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X1547 VDD a_7771_6925# a_7683_7317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X1548 hgu_sarlogic_flat_0.x5.x1[1].Q_N a_19460_6564# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X1549 a_7260_1461# a_6300_1179# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X1550 a_14352_1868# a_13182_1868# a_14245_2234# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0486 ps=0.63 w=0.36 l=0.15
X1551 a_9332_12677# hgu_sarlogic_flat_0.x2.x2.x3.IN a_9244_12539# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X1552 a_7598_8513# a_6370_8513# a_7456_8795# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X1553 a_2036_7824# hgu_sarlogic_flat_0.x3.x4.A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1554 a_11830_1153# a_12098_1363# a_12044_1461# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X1555 VSS hgu_cdac_half_0.db<6> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1556 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<15:0> hgu_cdac_half_0.d<4> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1557 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X1558 VDD a_11830_1153# a_11763_1545# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X1559 VSS hgu_cdac_half_0.d<6> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1560 a_8692_1179# hgu_sarlogic_flat_0.x4.x2.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1561 VSS a_3960_3698# hgu_sarlogic_flat_0.x4.x9.A1 VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1562 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X1563 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.db<6> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1564 VDD a_7772_8487# a_7684_8879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X1565 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<15:0> hgu_cdac_half_0.db<4> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1566 a_8398_1868# a_8232_1868# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1567 hgu_vgen_vref_0.phi2 a_n55304_6595# hgu_tah_0.VDD hgu_tah_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1568 a_18224_4670# a_18058_4670# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1569 VDD a_4362_1842# a_5093_2150# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X1570 a_8710_2530# hgu_sarlogic_flat_0.x4.x15.S VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X1571 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_1.db<5> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1572 a_n7660_7467# hgu_tah_0.tah_vp hgu_comp_flat_0.P VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1573 VSS hgu_cdac_half_0.d<6> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1574 a_5889_2708# VSS a_6031_2883# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X1575 hgu_cdac_half_1.VREF hgu_cdac_half_1.db<2> hgu_cdac_half_1.hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.35
X1576 a_4979_7798# hgu_sarlogic_flat_0.x3.x5.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1577 a_13370_1868# hgu_sarlogic_flat_0.x4.D[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X1578 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1579 a_18224_5316# a_18058_5316# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1580 VSS a_2988_8487# a_2923_8513# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X1581 a_4913_6444# a_4124_6052# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0819 ps=0.81 w=0.42 l=0.15
X1582 a_9762_6052# hgu_sarlogic_flat_0.x4.D[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1583 hgu_tah_0.VDD a_n55304_8227# hgu_vgen_vref_0.phi1 hgu_tah_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1584 VDD a_3960_3698# hgu_sarlogic_flat_0.x4.x9.A1 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1585 VSS a_3499_1331# hgu_cdac_sw_buffer_3.x4.A VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X1586 VSS hgu_sarlogic_flat_0.x3.D[0] a_8761_6951# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1587 a_19286_5950# a_18224_5950# a_19191_5950# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X1588 hgu_cdac_half_0.db<4> a_n148_n1104# hgu_cdac_sw_buffer_0.VDD hgu_cdac_sw_buffer_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1589 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.db<6> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1590 a_8710_2530# hgu_sarlogic_flat_0.x4.x15.S VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X1591 hgu_sarlogic_flat_0.x3.x5.A a_1587_9386# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1592 a_5182_6052# a_4437_6078# a_5318_6078# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1593 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<15:0> hgu_cdac_half_0.db<4> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.35
X1594 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1595 a_544_11360# a_407_11578# a_108_11334# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X1596 VDD hgu_comp_flat_0.clk hgu_comp_flat_0.P VDD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X1597 hgu_vgen_vref_0.mimtop2 VSS sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X1598 VSS hgu_cdac_half_1.d<6> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1599 a_11915_8513# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X1600 a_16020_5950# hgu_sarlogic_flat_0.x4.D[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X1601 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1602 hgu_sarlogic_flat_0.x1.x2.x3[1].floating async_setb_delay_cap_ctrl_code[1] hgu_sarlogic_flat_0.x1.x2.x9.output_stack VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X1603 VSS hgu_sarlogic_flat_0.x4.x20.S a_5897_7824# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1604 VDD hgu_sarlogic_flat_0.x3.x30.Q_N a_6516_6052# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.123 ps=1.17 w=0.42 l=0.15
X1605 hgu_cdac_sw_buffer_2.x3.A a_3165_1868# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X1606 a_4680_7798# a_4979_7798# a_4914_7824# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.066 ps=0.745 w=0.36 l=0.15
X1607 hgu_cdac_half_0.VREF hgu_cdac_half_0.db<6> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1608 VSS hgu_cdac_half_1.d<6> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1609 a_n6887_11999# hgu_comp_flat_0.clk a_n6959_12137# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X1610 a_16020_6590# hgu_sarlogic_flat_0.x3.D[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X1611 VSS hgu_sarlogic_flat_0.x3.x7.X a_10680_6078# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1612 a_3908_1179# hgu_sarlogic_flat_0.x4.x2.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.17 pd=1.81 as=0.154 ps=1.34 w=0.64 l=0.15
X1613 a_14654_7801# hgu_sarlogic_flat_0.x5.eob a_14566_7801# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X1614 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<15:0> hgu_cdac_half_1.db<4> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1615 VSS hgu_cdac_half_1.db<6> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1616 hgu_sarlogic_flat_0.x5.x3.X a_20768_8628# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X1617 a_n54850_7371# a_n54754_7113# hgu_tah_0.VDD hgu_tah_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.141 ps=1.33 w=0.42 l=0.15
X1618 a_n2219_8368# hgu_cdac_sw_buffer_2.x11.A VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1619 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.d<6> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1620 a_10771_1153# a_11317_1347# a_11275_1461# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.132 pd=1.22 as=0.0882 ps=1.05 w=0.84 l=0.15
X1621 VSS VDD a_1970_1842# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1622 VSS a_5379_6925# a_6086_6951# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1623 hgu_vgen_vref_0.mimtop2 VSS sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X1624 a_10978_1868# hgu_sarlogic_flat_0.x4.D[2] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X1625 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X1626 a_4401_9752# sel_bit[0] a_3898_9386# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0974 pd=0.97 as=0.0567 ps=0.69 w=0.42 l=0.15
X1627 hgu_cdac_half_0.VREF hgu_cdac_half_0.db<5> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1628 a_14679_9466# hgu_sarlogic_flat_0.x5.eob a_14591_9328# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X1629 a_9990_8513# a_8928_8513# a_9895_8513# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X1630 VSS a_9620_2136# a_10341_1868# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1631 hgu_sarlogic_flat_0.x4.x11.X a_5176_2883# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.158 ps=1.39 w=1 l=0.15
X1632 a_n54284_7371# hgu_vgen_vref_0.sky130_fd_sc_hd__dlymetal6s6s_1_4.A VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1633 a_n1158_n1744# hgu_cdac_sw_buffer_0.x11.A VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1634 a_14245_2234# a_13182_1868# a_14101_2150# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X1635 VSS hgu_cdac_half_1.d<1> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<1:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.35
X1636 hgu_cdac_half_0.d<6> a_1196_n1740# hgu_cdac_sw_buffer_1.VDD hgu_cdac_sw_buffer_1.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1637 a_6031_2883# hgu_sarlogic_flat_0.x4.x13.S VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X1638 hgu_tah_0.tah_vp hgu_tah_0.sw_n hgu_tah_0.tah_vp VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.454 ps=3.08 w=2.75 l=0.15
X1639 VSS a_6516_6052# hgu_sarlogic_flat_0.x3.x57.Q_N VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X1640 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1641 hgu_sarlogic_flat_0.x2.x2.x2.x5[7].floating hgu_sarlogic_flat_0.x2.x2.x2.x10.Y hgu_sarlogic_flat_0.x2.x2.x2.x9.output_stack VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X1642 VDD a_n595_7253# hgu_cdac_half_1.d<2> VDD sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1643 vip hgu_tah_0.sw_n hgu_tah_0.tah_vp hgu_tah_0.VDD sky130_fd_pr__pfet_01v8 ad=0.908 pd=5.83 as=1.71 ps=11.6 w=5.5 l=0.15
X1644 VDD a_9677_8487# a_10398_8795# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X1645 a_8909_7798# a_9222_7824# a_9328_7824# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1646 hgu_vgen_vref_0.mimtop2 VSS sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X1647 VSS hgu_cdac_sw_buffer_1.x3.X a_1666_n1100# VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1648 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_0.db<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1649 VDD a_8813_6052# hgu_sarlogic_flat_0.x4.D[4] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X1650 hgu_cdac_half_0.VREF hgu_cdac_half_0.d<6> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1651 a_8398_1868# a_8232_1868# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1652 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<7:0> hgu_cdac_half_1.db<3> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.122 ps=1.42 w=0.42 l=0.35
X1653 a_n53364_7835# hgu_vgen_vref_0.sky130_fd_sc_hd__nand2_1_0.Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1654 VDD hgu_sarlogic_flat_0.x4.x3.A a_n1058_3698# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1655 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<15:0> hgu_cdac_half_0.d<4> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1656 a_6031_2556# hgu_sarlogic_flat_0.x4.x13.S VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X1657 a_9332_11849# hgu_sarlogic_flat_0.x2.x2.x3.IN hgu_sarlogic_flat_0.x2.x2.x3.x9.output_stack VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X1658 a_4979_7798# hgu_sarlogic_flat_0.x3.x5.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1659 VSS VDD a_9328_7824# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.12 ps=1.08 w=0.42 l=0.15
X1660 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.db<6> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1661 a_7131_8513# a_7285_8487# a_6991_8487# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1662 VDD hgu_comp_flat_0.RS_n hgu_comp_flat_0.RS_p VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.15
X1663 hgu_cdac_half_0.VREF hgu_cdac_half_0.d<6> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1664 a_4976_1868# hgu_sarlogic_flat_0.x4.x2.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.03 as=0.0703 ps=0.755 w=0.42 l=0.15
X1665 hgu_sarlogic_flat_0.x1.x4.x5[7].floating hgu_sarlogic_flat_0.x1.x4.x10.Y hgu_sarlogic_flat_0.x1.x4.x9.output_stack VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X1666 hgu_cdac_sw_buffer_1.VDD a_1196_n1740# hgu_cdac_half_0.d<6> hgu_cdac_sw_buffer_1.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1667 a_4125_7798# a_4680_7798# a_4638_8106# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0882 ps=1.05 w=0.84 l=0.15
X1668 VSS a_4029_6052# hgu_sarlogic_flat_0.x4.D[6] VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X1669 hgu_sarlogic_flat_0.x4.x23.Q_N a_4836_2136# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X1670 VSS hgu_sarlogic_flat_0.x2.x7.A a_3314_11461# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1671 a_7706_6951# a_6369_6951# a_7597_6951# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X1672 hgu_sarlogic_flat_0.x3.x4.X a_2036_7824# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1673 a_12098_1363# a_11626_1153# a_12342_1545# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X1674 VSS a_n2251_7253# hgu_cdac_sw_buffer_2.x9.X VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1675 a_4001_14236# hgu_sarlogic_flat_0.x2.x3.A a_3929_14374# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X1676 hgu_cdac_half_0.VREF hgu_cdac_half_0.d<5> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1677 VSS hgu_cdac_half_1.d<6> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1678 hgu_sarlogic_flat_0.x3.x69.Q_N a_10163_6925# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X1679 VSS a_2586_6052# a_2585_6352# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1680 VSS hgu_cdac_sw_buffer_0.x3.X a_n688_n1104# VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1681 VSS hgu_sarlogic_flat_0.x4.D[6] a_2975_1179# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1682 a_6406_1179# a_6533_1347# a_5987_1153# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.03 as=0.0864 ps=0.91 w=0.64 l=0.15
X1683 hgu_cdac_sw_buffer_3.x11.X a_n4397_8367# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1684 a_10235_8008# a_9763_7798# a_10479_8190# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X1685 a_n890_2234# a_n1336_1868# a_n982_1868# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0651 ps=0.73 w=0.42 l=0.15
X1686 a_19372_5310# a_18224_5316# a_19286_5688# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X1687 hgu_cdac_half_0.VREF hgu_cdac_half_0.db<6> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1688 VSS hgu_cdac_half_1.db<6> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1689 hgu_tah_0.sw_n a_1945_10648# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X1690 a_11960_1868# a_10790_1868# a_11853_2234# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0486 ps=0.63 w=0.36 l=0.15
X1691 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1692 VSS hgu_cdac_half_0.d<6> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1693 VDD a_n3387_7727# hgu_cdac_half_1.db<4> VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1694 a_19372_6316# a_18224_5950# a_19286_5950# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X1695 a_1526_15136# a_1137_14764# a_1418_14758# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X1696 hgu_sarlogic_flat_0.x4.x2.X a_n424_3698# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1697 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<15:0> hgu_cdac_half_0.db<4> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1698 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<7:0> hgu_cdac_half_0.db<3> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1699 hgu_sarlogic_flat_0.x2.x2.x1.x5[7].floating hgu_sarlogic_flat_0.x2.x2.x1.x10.Y hgu_sarlogic_flat_0.x2.x2.x1.x9.output_stack VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X1700 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<15:0> hgu_cdac_half_1.db<4> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1701 VSS hgu_cdac_half_0.d<4> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<15:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1702 hgu_cdac_half_1.VREF hgu_cdac_half_1.d<5> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1703 hgu_tah_0.VDD a_n53364_7371# a_n53551_7113# hgu_tah_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X1704 a_6006_1868# a_5840_1868# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1705 a_n55770_7371# a_n55674_7113# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1706 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.122 ps=1.42 w=0.42 l=0.35
X1707 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<15:0> hgu_cdac_half_0.d<4> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1708 VDD a_1970_1842# a_2701_2150# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X1709 hgu_sarlogic_flat_0.x2.x2.x4.x4[3].floating sample_delay_cap_ctrl_code[2] hgu_sarlogic_flat_0.x2.x2.x4.x9.output_stack VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X1710 hgu_cdac_half_1.VREF hgu_cdac_half_1.db<4> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<15:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1711 VDD a_7575_7798# a_7508_8190# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X1712 a_n1147_7253# hgu_cdac_sw_buffer_2.x4.A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1713 hgu_vgen_vref_0.mimtop1 hgu_vgen_vref_0.mimbot1 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X1714 a_3497_2708# VSS a_3639_2883# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X1715 hgu_sarlogic_flat_0.x3.x4.A a_1422_7824# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1716 hgu_vgen_vref_0.mimtop1 hgu_vgen_vref_0.mimbot1 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X1717 VSS hgu_cdac_half_0.d<5> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1718 a_n6887_14037# hgu_comp_flat_0.ready a_n6959_14175# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X1719 hgu_cdac_half_0.VREF hgu_cdac_half_0.d<6> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1720 hgu_sarlogic_flat_0.x2.x2.x4.x9.output_stack hgu_sarlogic_flat_0.x2.x2.x4.x10.Y hgu_sarlogic_flat_0.x2.x2.x4.x5[7].floating VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X1721 a_13476_1179# hgu_sarlogic_flat_0.x4.x2.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.17 pd=1.81 as=0.154 ps=1.34 w=0.64 l=0.15
X1722 VDD a_1945_10648# hgu_tah_0.sw_n VDD sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.391 ps=3.14 w=1.26 l=0.15
X1723 VSS hgu_sarlogic_flat_0.x3.x4.X a_12069_8487# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1724 a_16894_5950# a_15832_5950# a_16799_5950# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X1725 hgu_cdac_half_0.VREF hgu_cdac_half_0.d<6> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1726 a_3499_1331# a_3595_1153# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1727 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1728 a_10023_11664# hgu_sarlogic_flat_0.x2.x2.x3.IN VDD VSS sky130_fd_pr__nfet_01v8 ad=0.0651 pd=0.73 as=0.0693 ps=0.75 w=0.42 l=0.15
X1729 a_n54850_7835# a_n54754_7657# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1730 VDD a_5379_6925# a_6086_6951# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X1731 VDD a_16581_5924# a_17302_6232# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X1732 hgu_cdac_half_0.VREF hgu_cdac_half_0.db<6> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1733 hgu_sarlogic_flat_0.x2.x2.x3.x5[7].floating hgu_sarlogic_flat_0.x2.x2.x3.x10.Y hgu_sarlogic_flat_0.x2.x2.x3.x9.output_stack VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X1734 VDD hgu_sarlogic_flat_0.x3.x27.Q_N a_4124_6052# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.123 ps=1.17 w=0.42 l=0.15
X1735 VSS hgu_cdac_half_1.db<6> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1736 VSS a_n2301_7728# hgu_cdac_sw_buffer_2.x11.A VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1737 VDD a_n1058_3698# hgu_sarlogic_flat_0.x4.x3.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1738 hgu_cdac_sw_buffer_0.VDD hgu_cdac_sw_buffer_0.x4.X a_n148_n1104# hgu_cdac_sw_buffer_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1739 a_12556_8487# a_12382_8513# a_12672_8513# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X1740 a_n335_1453# hgu_sarlogic_flat_0.x4.x7.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1741 a_3960_3698# hgu_sarlogic_flat_0.x4.x30.A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1742 VSS a_13636_1842# a_13570_1868# VSS sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0671 ps=0.75 w=0.42 l=0.15
X1743 VDD a_192_10793# hgu_comp_flat_0.clk VDD sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X1744 VSS hgu_cdac_half_0.db<4> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<15:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1745 VDD sample_delay_offset hgu_sarlogic_flat_0.x2.x2.x1.x6.SW VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1746 a_n6959_12413# hgu_comp_flat_0.clk a_n7047_12413# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X1747 VDD a_n6994_7879# a_n7390_7871# VDD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0.244 ps=2.26 w=0.84 l=0.15
X1748 hgu_cdac_sw_buffer_0.VDD a_n1158_n1744# hgu_cdac_half_0.db<6> hgu_cdac_sw_buffer_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1749 a_n424_3698# hgu_sarlogic_flat_0.x4.x3.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1750 hgu_cdac_half_1.VREF hgu_cdac_half_1.d<6> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1751 a_11853_2234# a_10790_1868# a_11709_2150# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X1752 hgu_sarlogic_flat_0.vdd_sw_b[7] a_52_2136# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X1753 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_1.db<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1754 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1755 hgu_cdac_half_1.VREF hgu_cdac_half_1.db<6> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1756 a_6829_6078# hgu_sarlogic_flat_0.x3.x4.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1757 VDD a_17068_5284# a_17775_5326# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X1758 a_18923_6590# a_18505_6590# a_18679_6564# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X1759 hgu_cdac_half_0.VREF hgu_cdac_half_0.db<1> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<1:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.35
X1760 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_1.d<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1761 hgu_cdac_half_1.VREF hgu_cdac_half_1.db<6> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1762 hgu_cdac_half_1.d<6> a_n2219_8368# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1763 a_11300_6052# a_11613_6078# a_11719_6078# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1764 a_6006_1868# a_5840_1868# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1765 a_9739_15176# hgu_sarlogic_flat_0.x2.x2.x4.x9.output_stack VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X1766 VSS hgu_cdac_half_1.db<5> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1767 VDD hgu_sarlogic_flat_0.x1.x9.Y a_611_11594# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X1768 hgu_sarlogic_flat_0.x5.eob a_2914_9360# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.335 ps=2.67 w=1 l=0.15
X1769 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.d<6> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1770 VSS VDD a_13582_1179# VSS sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.109 ps=1.03 w=0.42 l=0.15
X1771 a_11102_2530# hgu_sarlogic_flat_0.x4.x17.S VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X1772 VDD hgu_sarlogic_flat_0.x2.x3.Y a_2323_11578# VDD sky130_fd_pr__pfet_01v8 ad=0.406 pd=3.38 as=0.406 ps=3.38 w=1.4 l=0.15
X1773 a_4739_8513# a_4893_8487# a_4599_8487# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1774 VDD a_19460_4644# a_19372_5036# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X1775 VDD a_n4429_7252# hgu_cdac_sw_buffer_3.x9.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1776 VSS hgu_sarlogic_flat_0.x3.x36.Q_N a_11719_6078# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.12 ps=1.08 w=0.42 l=0.15
X1777 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1778 VSS a_1637_6052# hgu_sarlogic_flat_0.x4.x5.D VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X1779 hgu_sarlogic_flat_0.x5.x1[2].Q_N a_17068_5924# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X1780 hgu_cdac_sw_buffer_1.VDD hgu_cdac_sw_buffer_1.x4.X a_2206_n1100# hgu_cdac_sw_buffer_1.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1781 hgu_sarlogic_flat_0.x2.x1.x3.Y VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1782 hgu_sarlogic_flat_0.x2.x2.x3.IN hgu_sarlogic_flat_0.x2.x2.x2.x9.output_stack a_10023_11461# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.0651 ps=0.73 w=0.42 l=0.15
X1783 hgu_sarlogic_flat_0.x3.x75.Q a_6086_6951# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X1784 hgu_cdac_sw_buffer_1.VDD a_1716_n241# hgu_cdac_sw_buffer_1.x3.X hgu_cdac_sw_buffer_1.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1785 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<15:0> hgu_cdac_half_0.d<4> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1786 VSS hgu_cdac_half_0.d<5> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1787 a_n2773_7252# hgu_cdac_sw_buffer_3.x5.A VSS VSS sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1788 VDD a_18679_4644# a_18589_5036# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X1789 a_11102_2530# hgu_sarlogic_flat_0.x4.x17.S VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X1790 VSS VSS a_n2025_7088# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1791 a_5397_2556# hgu_sarlogic_flat_0.x4.x9.A1 a_5176_2883# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X1792 VSS hgu_comp_flat_0.ready a_n6959_13347# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X1793 VDD hgu_sarlogic_flat_0.x5.x3.X a_18058_5316# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1794 VDD a_2373_14732# a_3080_14774# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X1795 a_14436_1461# a_13476_1179# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X1796 a_3929_14788# hgu_sarlogic_flat_0.x2.x3.A a_3841_14650# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X1797 hgu_vgen_vref_0.mimtop1 hgu_vgen_vref_0.mimbot1 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X1798 VSS hgu_cdac_half_1.d<6> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1799 hgu_cdac_half_0.VREF hgu_cdac_half_0.db<6> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1800 VDD VDD a_11301_7798# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.123 ps=1.17 w=0.42 l=0.15
X1801 VSS a_n424_3698# hgu_sarlogic_flat_0.x4.x2.X VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1802 VSS hgu_cdac_half_1.db<6> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1803 a_n6994_7879# a_n6676_7789# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X1804 hgu_vgen_vref_0.mimtop2 VSS sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X1805 a_5116_8190# a_4979_7798# a_4680_7798# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X1806 a_12870_6444# a_12358_6052# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X1807 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X1808 a_n716_1842# hgu_sarlogic_flat_0.x4.x2.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X1809 a_16980_5310# a_15832_5316# a_16894_5688# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X1810 VDD a_2057_1453# a_2058_1153# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1811 VSS a_n53364_7835# a_n53551_7657# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X1812 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1813 a_16980_6316# a_15832_5950# a_16894_5950# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X1814 a_14726_8215# hgu_sarlogic_flat_0.x5.eob a_14654_8353# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X1815 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1816 a_4029_6052# a_4124_6052# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1817 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1818 a_8996_1868# hgu_sarlogic_flat_0.x4.x2.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0974 pd=0.97 as=0.0882 ps=0.84 w=0.42 l=0.15
X1819 a_5183_7798# a_5451_8008# a_5397_8106# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X1820 a_7575_7798# a_6830_7824# a_7711_7824# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1821 VSS a_7771_6925# a_7706_6951# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X1822 hgu_cdac_sw_buffer_1.VDD a_2544_n241# hgu_cdac_half_0.d<3> hgu_cdac_sw_buffer_1.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1823 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X1824 a_5496_8513# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X1825 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1826 hgu_sarlogic_flat_0.x3.x4.X a_2036_7824# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1827 a_6816_7317# a_6369_6951# a_6723_6951# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X1828 a_12358_6052# a_11613_6078# a_12494_6078# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1829 hgu_cdac_half_0.VREF hgu_cdac_half_0.d<6> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1830 a_11574_1545# a_10771_1153# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0787 pd=0.795 as=0.0956 ps=0.875 w=0.42 l=0.15
X1831 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_0.db<5> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1832 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<15:0> hgu_cdac_half_1.d<4> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1833 hgu_cdac_half_0.VREF hgu_cdac_half_0.d<4> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<15:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1834 a_5496_8513# a_4893_8487# a_5380_8487# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1835 a_8814_7798# a_8909_7798# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X1836 hgu_vgen_vref_0.mimtop2 VSS sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X1837 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_0.d<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1838 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.d<6> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.35
X1839 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<15:0> hgu_cdac_half_1.db<4> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1840 a_3408_9386# sel_bit[0] a_3309_9708# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.105 ps=0.995 w=0.42 l=0.15
X1841 VSS hgu_sarlogic_flat_0.x1.x9.A a_n1149_14701# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0651 ps=0.73 w=0.42 l=0.15
X1842 a_10710_13960# hgu_sarlogic_flat_0.x2.x2.x1.IN a_10638_14098# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X1843 hgu_sarlogic_flat_0.x2.x2.x2.x5[7].floating hgu_sarlogic_flat_0.x2.x2.x2.x10.Y hgu_sarlogic_flat_0.x2.x2.x2.x9.output_stack VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X1844 VSS hgu_sarlogic_flat_0.x3.x4.X a_9677_8487# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1845 hgu_cdac_sw_buffer_3.x11.A a_n4479_7727# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1846 a_5118_7824# a_4978_8098# a_4680_7798# VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.0711 ps=0.755 w=0.36 l=0.15
X1847 hgu_cdac_half_0.db<6> a_n1158_n1744# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1848 hgu_cdac_half_0.VREF hgu_cdac_half_0.d<5> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1849 hgu_sarlogic_flat_0.x4.x9.A1 a_3960_3698# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1850 hgu_cdac_half_0.VREF hgu_cdac_half_0.db<6> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1851 hgu_sarlogic_flat_0.x4.x17.X a_12352_2883# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.158 ps=1.39 w=1 l=0.15
X1852 a_14101_2150# a_13636_1842# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X1853 a_12495_7824# a_12627_8008# a_12359_7798# VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0864 ps=0.91 w=0.64 l=0.15
X1854 hgu_cdac_half_0.VREF hgu_cdac_half_0.db<4> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<15:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1855 a_11855_6052# a_12153_6352# a_12089_6444# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0924 ps=0.86 w=0.42 l=0.15
X1856 VSS hgu_cdac_half_0.db<4> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<15:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.35
X1857 a_4543_6078# a_4679_6052# a_4124_6052# VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0864 ps=0.91 w=0.64 l=0.15
X1858 VDD a_16287_5284# a_16197_5310# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X1859 a_13880_2150# a_13462_2234# a_13636_1842# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X1860 VSS hgu_cdac_sw_buffer_0.x11.A a_n1158_n1744# VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1861 a_9116_8513# hgu_sarlogic_flat_0.x4.x9.S VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X1862 hgu_tah_0.tah_vn hgu_tah_0.sw_n hgu_tah_0.tah_vn VSS sky130_fd_pr__nfet_01v8 ad=4.43 pd=30.7 as=0.454 ps=3.08 w=2.75 l=0.15
X1863 VDD a_16287_5924# a_16197_6316# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X1864 a_19395_4670# a_18058_4670# a_19286_4670# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X1865 hgu_cdac_half_1.VREF hgu_cdac_half_1.d<6> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1866 a_16113_12677# hgu_sarlogic_flat_0.x2.x2.x2.IN a_16041_12677# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X1867 hgu_cdac_sw_buffer_3.x11.X a_n4397_8367# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1868 hgu_vgen_vref_0.mimtop1 hgu_vgen_vref_0.mimbot1 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X1869 a_8928_8513# a_8762_8513# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1870 a_6370_2234# a_6006_1868# a_6286_2234# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X1871 a_2444_2136# hgu_sarlogic_flat_0.x4.x2.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.132 pd=1.22 as=0.0956 ps=0.875 w=0.42 l=0.15
X1872 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_1.d<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1873 hgu_sarlogic_flat_0.x3.x7.X a_1454_6950# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1874 a_11301_7798# a_11856_7798# a_11814_8106# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0882 ps=1.05 w=0.84 l=0.15
X1875 a_2975_1179# a_2057_1453# a_2530_1363# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.0567 ps=0.69 w=0.42 l=0.15
X1876 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_0.db<5> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1877 a_4143_6951# a_3977_6951# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1878 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1879 VSS a_n1287_2708# hgu_sarlogic_flat_0.x4.x6.X VSS sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X1880 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.db<6> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1881 VSS hgu_sarlogic_flat_0.x5.x3.X a_18058_5950# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1882 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1883 VSS hgu_cdac_half_1.d<5> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1884 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.db<6> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1885 a_18679_6564# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X1886 a_10638_13960# hgu_sarlogic_flat_0.x2.x2.x1.IN a_10550_13822# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X1887 a_6830_7824# hgu_sarlogic_flat_0.x3.x4.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.154 ps=1.34 w=0.64 l=0.15
X1888 VSS hgu_sarlogic_flat_0.x5.eob a_14654_7525# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X1889 VSS hgu_sarlogic_flat_0.x5.x3.X a_18058_6596# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1890 VDD hgu_sarlogic_flat_0.x4.x7.S a_608_2883# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.0767 ps=0.785 w=0.42 l=0.15
X1891 hgu_sarlogic_flat_0.x2.x2.x1.x5[7].floating hgu_sarlogic_flat_0.x2.x2.x1.x10.Y hgu_sarlogic_flat_0.x2.x2.x1.x9.output_stack VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X1892 a_9292_7317# a_8761_6951# a_9208_7317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X1893 VSS hgu_sarlogic_flat_0.x4.D[3] a_10151_1179# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1894 a_n335_1453# hgu_sarlogic_flat_0.x4.x7.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1895 a_2308_15136# a_971_14764# a_2199_15136# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X1896 a_5379_6925# hgu_sarlogic_flat_0.x3.x77.Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X1897 a_13582_1179# a_13709_1347# a_13163_1153# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.03 as=0.0864 ps=0.91 w=0.64 l=0.15
X1898 a_n782_1868# a_n1336_1868# a_n890_2234# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0675 ps=0.735 w=0.36 l=0.15
X1899 a_9962_2883# VSS a_9962_2556# VSS sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X1900 hgu_vgen_vref_0.phi1 a_n55304_8227# hgu_tah_0.VDD hgu_tah_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1901 VDD a_13065_2708# hgu_sarlogic_flat_0.x4.x18.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X1902 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_1.d<5> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.35
X1903 hgu_cdac_half_1.VREF hgu_cdac_half_1.db<5> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1904 hgu_tah_0.VDD a_n54284_7835# a_n54471_7657# hgu_tah_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X1905 VSS hgu_sarlogic_flat_0.x4.x7.S a_615_2556# VSS sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.0693 ps=0.75 w=0.42 l=0.15
X1906 hgu_cdac_half_1.VREF hgu_cdac_half_1.db<5> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1907 hgu_sarlogic_flat_0.x2.x2.x4.x9.output_stack hgu_sarlogic_flat_0.x2.x2.x4.x10.Y hgu_sarlogic_flat_0.x2.x2.x4.x5[7].floating VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X1908 a_9293_8879# a_8762_8513# a_9209_8879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X1909 hgu_cdac_half_0.VREF hgu_cdac_half_0.d<5> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1910 VSS hgu_cdac_half_0.db<5> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1911 a_5380_8487# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X1912 a_n607_7947# VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1913 a_9950_1545# a_9438_1153# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X1914 VDD a_n4479_7727# hgu_cdac_sw_buffer_3.x11.A VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1915 a_19694_6590# a_19286_6968# a_19460_6564# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X1916 a_n6959_13623# hgu_comp_flat_0.ready a_n7047_13623# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X1917 VSS hgu_cdac_sw_buffer_2.x11.A a_n2219_8368# VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1918 a_n716_1842# a_n890_2234# a_n572_1868# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.0974 ps=0.97 w=0.64 l=0.15
X1919 hgu_sarlogic_flat_0.x2.x2.x4.x9.output_stack hgu_sarlogic_flat_0.x2.x2.x4.x10.Y hgu_sarlogic_flat_0.x2.x2.x4.x5[7].floating VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X1920 hgu_sarlogic_flat_0.x2.x2.x3.x9.output_stack sample_delay_cap_ctrl_code[14] hgu_sarlogic_flat_0.x2.x2.x3.x4[3].floating VSS sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X1921 VSS hgu_sarlogic_flat_0.x3.x4.A a_2036_7824# VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1922 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1923 VSS hgu_cdac_half_0.d<6> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1924 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<7:0> hgu_cdac_half_0.d<3> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.122 ps=1.42 w=0.42 l=0.35
X1925 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1926 a_7029_6360# a_6829_6078# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X1927 VDD a_14404_2136# a_14329_2234# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0956 pd=0.875 as=0.0787 ps=0.795 w=0.42 l=0.15
X1928 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1929 a_1637_6052# a_1732_6052# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1930 a_9438_1153# a_8692_1179# a_9574_1179# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1931 a_8852_1842# hgu_sarlogic_flat_0.x4.x2.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X1932 a_2392_1868# a_1222_1868# a_2285_2234# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0486 ps=0.63 w=0.36 l=0.15
X1933 VDD hgu_sarlogic_flat_0.x3.x7.A a_1454_6950# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1934 VSS hgu_cdac_half_1.db<4> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<15:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1935 VSS hgu_cdac_half_0.d<6> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1936 hgu_cdac_half_1.VREF hgu_cdac_half_1.d<6> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1937 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1938 VSS a_n4397_8367# hgu_cdac_sw_buffer_3.x11.X VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1939 a_8883_1461# a_8692_1179# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X1940 hgu_sarlogic_flat_0.x3.x5.A a_1587_9386# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1941 hgu_comp_flat_0.P hgu_tah_0.tah_vp a_n7660_7467# VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1942 result[7] a_20167_4670# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X1943 hgu_cdac_half_1.VREF hgu_cdac_half_1.db<6> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1944 hgu_sarlogic_flat_0.x5.x2.x9.output_stack hgu_sarlogic_flat_0.x5.x2.x10.Y hgu_sarlogic_flat_0.x5.x2.x5[7].floating VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X1945 VDD hgu_sarlogic_flat_0.x5.x3.X a_18058_4670# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1946 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.d<6> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1947 VSS a_4836_2136# a_5557_1868# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1948 a_16113_11849# hgu_sarlogic_flat_0.x2.x2.x2.IN a_16041_11849# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X1949 hgu_vgen_vref_0.sky130_fd_sc_hd__inv_1_3.A hgu_vgen_vref_0.sky130_fd_sc_hd__inv_1_1.A hgu_tah_0.VDD hgu_tah_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1950 VDD a_n7216_6420# hgu_comp_flat_0.comp_outp VDD sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.3 as=0.139 ps=1.17 w=0.84 l=0.15
X1951 a_52_2136# a_n107_2234# a_192_1868# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.109 ps=1.03 w=0.64 l=0.15
X1952 a_14490_1363# a_14017_1453# a_14734_1179# VSS sky130_fd_pr__nfet_01v8 ad=0.0675 pd=0.735 as=0.0671 ps=0.75 w=0.36 l=0.15
X1953 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.d<6> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1954 VSS hgu_sarlogic_flat_0.x4.x18.X a_13016_1868# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1955 VDD a_6754_1842# a_6704_2150# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X1956 a_1410_1868# hgu_sarlogic_flat_0.x4.D[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X1957 a_8740_2883# hgu_sarlogic_flat_0.x4.x9.A1 a_8281_2708# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X1958 VDD VDD a_9146_1842# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.17 ps=1.81 w=0.64 l=0.15
X1959 VDD a_n422_1842# a_n472_2150# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X1960 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.db<6> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1961 VDD a_6422_7798# hgu_sarlogic_flat_0.x4.x20.S VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X1962 VDD hgu_sarlogic_flat_0.x3.x75.Q a_6369_6951# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1963 a_11319_6951# a_11153_6951# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1964 a_1164_n241# hgu_cdac_sw_buffer_1.x9.A hgu_cdac_sw_buffer_1.VDD hgu_cdac_sw_buffer_1.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1965 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_1.db<5> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1966 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_0.d<5> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1967 VSS a_2057_1453# a_2058_1153# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1968 VSS a_1114_n1100# hgu_cdac_sw_buffer_1.x11.A VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1969 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X1970 hgu_vgen_vref_0.mimtop1 hgu_vgen_vref_0.phi1_n hgu_vgen_vref_0.vcm hgu_tah_0.VDD sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=0.5
X1971 VSS a_8710_2530# a_8644_2556# VSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X1972 VSS hgu_cdac_half_1.db<3> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<7:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1973 VSS a_n55304_8227# hgu_vgen_vref_0.phi1 VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1974 a_n7760_6349# a_n6526_6819# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.139 pd=1.17 as=0.26 ps=2.3 w=0.84 l=0.15
X1975 a_8925_1347# a_9233_1453# a_9182_1545# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0787 ps=0.795 w=0.42 l=0.15
X1976 VSS hgu_cdac_half_0.db<6> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1977 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X1978 VSS a_611_11594# a_546_11738# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0935 ps=0.965 w=0.64 l=0.15
X1979 hgu_cdac_half_0.db<6> a_n1158_n1744# hgu_cdac_sw_buffer_0.VDD hgu_cdac_sw_buffer_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1980 hgu_vgen_vref_0.mimtop1 hgu_vgen_vref_0.mimbot1 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X1981 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X1982 a_2988_8487# a_2814_8513# a_3104_8513# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X1983 a_19395_6968# a_18058_6596# a_19286_6968# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X1984 a_6724_8513# hgu_sarlogic_flat_0.x4.x7.S VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X1985 a_11036_2556# VSS a_10673_2708# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X1986 a_17003_4670# a_15666_4670# a_16894_4670# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X1987 VSS a_4068_1842# a_4002_1868# VSS sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0671 ps=0.75 w=0.42 l=0.15
X1988 a_16041_12401# hgu_sarlogic_flat_0.x2.x2.x2.IN a_15953_12263# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X1989 VSS hgu_sarlogic_flat_0.x3.x27.Q_N a_5318_6078# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.101 ps=0.99 w=0.42 l=0.15
X1990 vip hgu_tah_0.sw hgu_tah_0.tah_vp VSS sky130_fd_pr__nfet_01v8 ad=0.454 pd=3.08 as=0.454 ps=3.08 w=2.75 l=0.15
X1991 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1992 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1993 a_2036_7824# hgu_sarlogic_flat_0.x3.x4.A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1994 VSS a_5183_7798# a_5118_7824# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0935 ps=0.965 w=0.64 l=0.15
X1995 a_2285_2234# a_1222_1868# a_2141_2150# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X1996 a_9404_12125# hgu_sarlogic_flat_0.x2.x2.x3.IN a_9332_12125# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X1997 hgu_cdac_sw_buffer_1.x12.X a_1942_n460# hgu_cdac_sw_buffer_1.VDD hgu_cdac_sw_buffer_1.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1998 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1999 hgu_sarlogic_flat_0.x4.D[2] a_13262_6951# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X2000 hgu_sarlogic_flat_0.x3.x4.X a_2036_7824# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2001 a_7789_8106# a_6830_7824# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X2002 VSS a_11301_7798# hgu_sarlogic_flat_0.x3.x39.Q_N VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X2003 VDD VDD a_2262_1153# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X2004 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2005 hgu_sarlogic_flat_0.x3.x72.Q_N a_7771_6925# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X2006 VSS a_3960_3698# hgu_sarlogic_flat_0.x4.x9.A1 VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2007 a_13065_2708# hgu_sarlogic_flat_0.x4.x9.A1 a_13207_2556# VSS sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X2008 a_19191_6912# a_18679_6564# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X2009 VDD a_3326_3698# hgu_sarlogic_flat_0.x4.x30.A VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2010 a_14155_1545# a_14018_1153# a_13709_1347# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X2011 hgu_cdac_half_0.VREF hgu_cdac_half_0.db<6> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2012 hgu_vgen_vref_0.sky130_fd_sc_hd__nand2_1_1.Y hgu_vgen_vref_0.sky130_fd_sc_hd__inv_1_2.Y hgu_tah_0.VDD hgu_tah_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2013 result[1] a_20167_6606# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X2014 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_0.d<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2015 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.d<6> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2016 VSS VDD a_4014_1179# VSS sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.109 ps=1.03 w=0.42 l=0.15
X2017 VSS hgu_cdac_half_1.d<6> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2018 hgu_cdac_sw_buffer_3.x11.X a_n4397_8367# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2019 a_18505_6590# a_18224_6596# a_18412_6590# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X2020 VDD hgu_sarlogic_flat_0.x4.x18.X a_13016_1868# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2021 a_n1149_14701# hgu_sarlogic_flat_0.x1.x2.x9.output_stack VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X2022 VDD a_n447_11350# hgu_sarlogic_flat_0.x1.x27.Q_N VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X2023 a_6900_7317# a_6369_6951# a_6816_7317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X2024 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<15:0> hgu_cdac_half_0.db<4> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2025 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_1.d<5> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2026 a_9209_8879# a_8762_8513# a_9116_8513# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X2027 a_11206_7798# a_11301_7798# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X2028 VDD a_10673_2708# hgu_sarlogic_flat_0.x4.x16.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X2029 hgu_sarlogic_flat_0.x3.x30.Q_N a_7772_8487# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X2030 a_5205_6951# a_3977_6951# a_5063_7233# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X2031 hgu_vgen_vref_0.vcm hgu_vgen_vref_0.phi1 hgu_vgen_vref_0.mimtop1 VSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=0.5
X2032 VSS a_19460_4644# a_19395_4670# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X2033 VSS hgu_cdac_half_0.db<5> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2034 a_18505_5036# a_18058_4670# a_18412_4670# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X2035 hgu_sarlogic_flat_0.x4.x2.X a_n424_3698# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2036 VDD hgu_sarlogic_flat_0.x4.x20.S a_4401_9752# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.0974 ps=0.97 w=0.64 l=0.15
X2037 VSS a_9383_8487# a_9317_8513# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X2038 VDD a_5379_6925# a_5291_7317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X2039 VSS a_19460_5284# a_19395_5688# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X2040 hgu_sarlogic_flat_0.x2.x2.x2.x6.SW sample_delay_offset VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2041 a_6901_8879# a_6370_8513# a_6817_8879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X2042 a_6422_7798# a_6517_7798# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2043 hgu_sarlogic_flat_0.x5.x1[5].Q_N a_19460_5284# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X2044 hgu_sarlogic_flat_0.x2.x2.x2.x5[7].floating hgu_sarlogic_flat_0.x2.x2.x2.x10.Y hgu_sarlogic_flat_0.x2.x2.x2.x9.output_stack VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X2045 VSS a_18679_4644# a_18613_4670# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X2046 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_1.db<5> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2047 a_5206_8513# a_3978_8513# a_5064_8795# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X2048 a_12359_7798# a_12627_8008# a_12573_8106# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X2049 hgu_sarlogic_flat_0.x3.x4.A a_1422_7824# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2050 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X2051 VSS a_2373_14732# a_2308_15136# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X2052 VDD a_12556_8487# a_13263_8513# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X2053 VSS hgu_cdac_half_0.d<6> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2054 hgu_vgen_vref_0.mimtop2 VSS sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X2055 VSS a_18679_5284# a_18613_5688# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X2056 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X2057 a_3302_6444# a_2790_6052# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X2058 a_3898_9386# sel_bit[0] a_4196_9386# VSS sky130_fd_pr__nfet_01v8 ad=0.072 pd=0.76 as=0.0671 ps=0.75 w=0.36 l=0.15
X2059 a_10771_1153# a_11084_1179# a_11190_1179# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2060 a_2199_15136# a_1137_14764# a_2104_15080# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X2061 VSS a_n1158_n1744# hgu_cdac_half_0.db<6> VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2062 VDD hgu_cdac_sw_buffer_2.x4.X a_n1209_7728# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2063 hgu_cdac_half_0.d<6> a_1196_n1740# hgu_cdac_sw_buffer_1.VDD hgu_cdac_sw_buffer_1.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2064 VDD a_13163_1153# hgu_sarlogic_flat_0.x4.x35.Q_N VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X2065 a_8678_2234# a_8232_1868# a_8586_1868# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0651 ps=0.73 w=0.42 l=0.15
X2066 hgu_sarlogic_flat_0.x1.x4.x3[1].floating async_resetb_delay_cap_ctrl_code[1] hgu_sarlogic_flat_0.x1.x4.x9.output_stack VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X2067 a_11320_8513# a_11154_8513# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2068 a_10075_7317# a_8927_6951# a_9989_6951# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X2069 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<15:0> hgu_cdac_half_1.d<4> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2070 hgu_cdac_half_1.VREF hgu_cdac_half_1.d<6> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2071 hgu_sarlogic_flat_0.x5.x2.x9.output_stack retimer_delay_offset hgu_sarlogic_flat_0.x5.x2.x7.floating VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X2072 VSS hgu_cdac_half_0.d<5> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2073 VSS hgu_cdac_sw_buffer_1.x11.A a_1196_n1740# VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2074 hgu_vgen_vref_0.mimtop2 VSS sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X2075 hgu_cdac_half_0.VREF hgu_cdac_half_0.d<6> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2076 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<7:0> hgu_cdac_half_0.d<3> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.35
X2077 VSS a_1107_1331# hgu_cdac_sw_buffer_3.x3.A VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X2078 hgu_sarlogic_flat_0.x2.x2.x4.x9.output_stack hgu_sarlogic_flat_0.x2.x3.A a_3866_15625# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X2079 VDD a_n1058_3698# hgu_sarlogic_flat_0.x4.x3.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2080 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<15:0> hgu_cdac_half_1.db<4> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2081 VSS hgu_cdac_half_1.db<6> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2082 hgu_cdac_half_0.VREF hgu_cdac_half_0.d<6> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2083 a_n6959_11999# hgu_comp_flat_0.clk a_n7047_11861# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X2084 hgu_cdac_half_0.db<6> a_n1158_n1744# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2085 VSS hgu_sarlogic_flat_0.x4.x16.X a_10624_1868# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2086 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.d<6> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2087 a_10076_8879# a_8928_8513# a_9990_8513# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X2088 hgu_vgen_vref_0.mimtop2 VSS sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X2089 hgu_cdac_half_1.VREF hgu_cdac_half_1.db<4> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<15:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2090 VDD a_2323_10792# a_1945_10648# VDD sky130_fd_pr__pfet_01v8 ad=0.365 pd=3.1 as=0.365 ps=3.1 w=1.26 l=0.15
X2091 hgu_cdac_half_1.d<5> a_n1749_7728# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2092 hgu_cdac_sw_buffer_1.VDD a_1196_n1740# hgu_cdac_half_0.d<6> hgu_cdac_sw_buffer_1.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2093 a_1516_1179# hgu_sarlogic_flat_0.x4.x2.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.17 pd=1.81 as=0.154 ps=1.34 w=0.64 l=0.15
X2094 VSS hgu_cdac_half_1.d<5> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2095 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.db<6> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2096 VSS hgu_sarlogic_flat_0.x2.x7.A hgu_sarlogic_flat_0.x2.x7.Y VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2097 a_19460_6564# a_19286_6968# a_19576_6956# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X2098 VSS hgu_cdac_half_0.db<6> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2099 a_192_1868# hgu_sarlogic_flat_0.x4.x2.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.03 as=0.0703 ps=0.755 w=0.42 l=0.15
X2100 VDD a_18973_4644# a_18923_4952# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X2101 hgu_cdac_half_1.VREF hgu_cdac_half_1.d<6> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2102 VDD hgu_comp_flat_0.clk a_3050_3698# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X2103 hgu_cdac_half_1.db<5> a_n3927_7727# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2104 a_6533_1347# a_6841_1453# a_6790_1545# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0787 ps=0.795 w=0.42 l=0.15
X2105 hgu_cdac_half_1.VREF hgu_cdac_half_1.db<5> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2106 a_1448_10615# hgu_tah_0.sw VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X2107 hgu_sarlogic_flat_0.x2.x2.x1.x5[7].floating hgu_sarlogic_flat_0.x2.x2.x1.x10.Y hgu_sarlogic_flat_0.x2.x2.x1.x9.output_stack VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X2108 hgu_cdac_half_1.VREF hgu_cdac_half_1.db<6> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2109 VSS hgu_cdac_half_1.db<2> hgu_cdac_half_1.hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2110 hgu_cdac_sw_buffer_1.VDD hgu_cdac_sw_buffer_1.x3.X a_1666_n1100# hgu_cdac_sw_buffer_1.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2111 a_13546_2234# a_13182_1868# a_13462_2234# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X2112 hgu_cdac_half_1.d<6> a_n2219_8368# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2113 a_7598_8513# a_6536_8513# a_7503_8513# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X2114 a_n871_7253# hgu_cdac_sw_buffer_2.x6.A VSS VSS sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2115 hgu_sarlogic_flat_0.x3.x4.X a_2036_7824# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2116 a_17003_6968# a_15666_6596# a_16894_6968# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X2117 a_17068_4644# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X2118 hgu_cdac_sw_buffer_2.x4.A a_5557_1868# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X2119 a_4312_2150# a_3894_2234# a_4068_1842# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X2120 hgu_sarlogic_flat_0.x3.x4.X a_2036_7824# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2121 VSS a_1676_1842# a_1610_1868# VSS sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0671 ps=0.75 w=0.42 l=0.15
X2122 a_3408_9386# a_3378_9360# a_3313_9386# VSS sky130_fd_pr__nfet_01v8 ad=0.072 pd=0.76 as=0.066 ps=0.745 w=0.36 l=0.15
X2123 a_16113_6316# a_15666_5950# a_16020_5950# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X2124 hgu_sarlogic_flat_0.x4.x3.A a_n1334_3698# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2125 VSS a_3960_3698# hgu_sarlogic_flat_0.x4.x9.A1 VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2126 VSS hgu_cdac_half_0.d<6> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2127 VSS VDD a_14358_1179# VSS sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0974 ps=0.97 w=0.42 l=0.15
X2128 a_382_1179# a_n130_1153# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0882 ps=0.84 w=0.42 l=0.15
X2129 VDD hgu_sarlogic_flat_0.x4.x11.S a_4922_2883# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.118 ps=1.4 w=0.42 l=0.15
X2130 a_n6887_12551# hgu_comp_flat_0.clk a_n6959_12551# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X2131 hgu_sarlogic_flat_0.x2.x1.x2.D a_2373_14732# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X2132 hgu_sarlogic_flat_0.x2.x2.x4.x9.output_stack hgu_sarlogic_flat_0.x2.x2.x4.x10.Y hgu_sarlogic_flat_0.x2.x2.x4.x5[7].floating VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X2133 hgu_sarlogic_flat_0.x2.x2.x3.x9.output_stack sample_delay_cap_ctrl_code[14] hgu_sarlogic_flat_0.x2.x2.x3.x4[3].floating VSS sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X2134 VSS a_n4429_7252# hgu_cdac_sw_buffer_3.x9.X VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X2135 a_n7660_7467# hgu_tah_0.tah_vn hgu_comp_flat_0.Q VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.165 ps=1.33 w=1 l=0.15
X2136 VSS a_7046_1153# a_6956_1179# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.116 ps=1.09 w=0.64 l=0.15
X2137 hgu_cdac_sw_buffer_3.x11.X a_n4397_8367# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2138 VSS hgu_cdac_half_0.d<6> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2139 a_3314_11461# hgu_sarlogic_flat_0.x2.x7.A VSS VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.0693 ps=0.75 w=0.42 l=0.15
X2140 VSS a_16287_5924# a_16221_5950# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X2141 hgu_sarlogic_flat_0.x4.x2.X a_n424_3698# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2142 a_11244_1842# hgu_sarlogic_flat_0.x4.x2.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X2143 a_n1189_1153# a_n643_1347# a_n685_1461# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.132 pd=1.22 as=0.0882 ps=1.05 w=0.84 l=0.15
X2144 hgu_sarlogic_flat_0.x3.x75.Q_N a_5379_6925# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X2145 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.d<6> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2146 a_9877_2150# a_9461_2234# a_9620_2136# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.132 ps=1.22 w=0.84 l=0.15
X2147 a_10673_2708# hgu_sarlogic_flat_0.x4.x9.A1 a_10815_2556# VSS sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X2148 VSS hgu_sarlogic_flat_0.x4.x11.S a_4922_2883# VSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.109 ps=1.36 w=0.42 l=0.15
X2149 hgu_cdac_half_1.d<6> a_n2219_8368# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2150 VSS a_16287_6564# a_16221_6968# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X2151 a_11763_1545# a_11626_1153# a_11317_1347# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X2152 hgu_sarlogic_flat_0.x4.x19.Q_N a_2444_2136# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X2153 VSS hgu_cdac_half_1.d<6> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2154 a_14679_9742# hgu_sarlogic_flat_0.x5.eob a_14591_9880# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X2155 VSS VDD a_1622_1179# VSS sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.109 ps=1.03 w=0.42 l=0.15
X2156 VSS a_n424_3698# hgu_sarlogic_flat_0.x4.x2.X VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2157 VDD hgu_sarlogic_flat_0.x4.x16.X a_10624_1868# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2158 VSS hgu_cdac_half_0.d<5> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2159 hgu_vgen_vref_0.mimtop1 hgu_vgen_vref_0.mimbot1 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X2160 VDD hgu_sarlogic_flat_0.x4.D[1] a_14935_1179# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X2161 hgu_cdac_half_0.VREF hgu_cdac_half_0.db<6> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2162 VDD a_n1209_7728# hgu_cdac_half_1.d<4> VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2163 VSS hgu_cdac_half_1.db<6> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2164 hgu_sarlogic_flat_0.x3.x27.Q_N a_5380_8487# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X2165 hgu_vgen_vref_0.mimbot1 hgu_vgen_vref_0.phi2 hgu_vgen_vref_0.mimtop2 VSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=0.5
X2166 a_18505_6590# a_18058_6596# a_18412_6590# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X2167 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_0.d<5> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2168 a_2914_9360# a_3783_9360# a_3408_9386# VSS sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2169 hgu_tah_0.VDD a_n53647_7371# a_n53834_7113# hgu_tah_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X2170 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.d<6> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2171 hgu_tah_0.sw a_1945_11268# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2172 hgu_vgen_vref_0.mimtop1 hgu_vgen_vref_0.mimbot1 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X2173 VSS hgu_sarlogic_flat_0.x2.x2.x2.x9.output_stack a_10023_11664# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X2174 VSS a_6991_8487# a_6925_8513# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X2175 a_10663_16039# hgu_sarlogic_flat_0.x2.x2.x1.IN a_10575_16177# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X2176 hgu_cdac_half_1.VREF hgu_cdac_half_1.d<4> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<15:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2177 hgu_cdac_half_1.VREF hgu_cdac_half_1.d<5> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2178 a_2476_1461# a_1516_1179# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X2179 a_2814_8513# a_1586_8513# a_2672_8795# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X2180 hgu_sarlogic_flat_0.x4.x13.X a_7570_2883# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.158 ps=1.39 w=1 l=0.15
X2181 hgu_cdac_half_1.VREF hgu_cdac_half_1.db<4> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<15:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2182 VSS a_12556_8487# a_13263_8513# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X2183 a_11614_7824# hgu_sarlogic_flat_0.x3.x4.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2184 VDD a_10164_8487# a_10871_8513# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X2185 a_3908_1179# hgu_sarlogic_flat_0.x4.x2.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2186 hgu_cdac_half_1.VREF hgu_cdac_half_1.db<6> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2187 VDD a_2988_8487# a_2900_8879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X2188 VDD a_12068_6925# a_12018_7233# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X2189 hgu_cdac_half_0.hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT hgu_cdac_half_0.db<2> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2190 a_1325_14758# hgu_sarlogic_flat_0.x2.x1.x2.D VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X2191 VSS a_n4397_8367# hgu_cdac_sw_buffer_3.x11.X VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2192 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2193 a_n107_2234# a_n1170_1868# a_n251_2150# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X2194 a_2045_6078# hgu_sarlogic_flat_0.x3.x4.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.154 ps=1.34 w=0.64 l=0.15
X2195 hgu_cdac_half_0.VREF hgu_cdac_half_0.d<6> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2196 VSS a_1945_11268# hgu_tah_0.sw VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2197 hgu_sarlogic_flat_0.x4.x9.A1 a_3960_3698# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2198 VDD a_12069_8487# a_12019_8795# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X2199 hgu_sarlogic_flat_0.x2.x2.x4.x9.output_stack hgu_sarlogic_flat_0.x2.x2.x4.x6.SW hgu_sarlogic_flat_0.x2.x2.x4.x6.floating VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X2200 a_n6292_6446# hgu_comp_flat_0.RS_n VSS VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X2201 a_10181_8106# a_9222_7824# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X2202 a_n7678_6901# a_n7760_6349# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.15
X2203 VSS hgu_cdac_half_1.d<4> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<15:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2204 hgu_comp_flat_0.Q a_n6676_7789# a_n6994_7879# VSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X2205 hgu_cdac_half_0.VREF hgu_cdac_half_0.d<5> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2206 VSS a_12012_2136# a_11960_1868# VSS sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.066 ps=0.745 w=0.42 l=0.15
X2207 a_4922_1363# a_4449_1453# a_5166_1179# VSS sky130_fd_pr__nfet_01v8 ad=0.0675 pd=0.735 as=0.0671 ps=0.75 w=0.36 l=0.15
X2208 VSS a_n2219_8368# hgu_cdac_half_1.d<6> VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2209 a_n2219_8368# hgu_cdac_sw_buffer_2.x11.A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2210 a_10164_8487# a_9990_8513# a_10280_8513# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X2211 VSS hgu_cdac_half_0.db<5> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2212 hgu_cdac_sw_buffer_1.VDD a_2206_n1100# hgu_cdac_half_0.d<4> hgu_cdac_sw_buffer_1.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2213 VSS VDD a_7711_7824# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.101 ps=0.99 w=0.42 l=0.15
X2214 hgu_sarlogic_flat_0.x1.x4.x9.output_stack hgu_sarlogic_flat_0.x1.x4.x10.Y hgu_sarlogic_flat_0.x1.x4.x5[7].floating VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X2215 VDD hgu_sarlogic_flat_0.x2.x7.Y hgu_sarlogic_flat_0.x2.x3.Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2216 hgu_cdac_half_1.VREF hgu_cdac_half_1.d<6> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2217 hgu_cdac_sw_buffer_3.x11.X a_n4397_8367# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2218 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.db<6> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2219 hgu_cdac_half_1.VREF hgu_cdac_half_1.db<6> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2220 a_11070_2234# a_10790_1868# a_10978_1868# VSS sky130_fd_pr__nfet_01v8 ad=0.0675 pd=0.735 as=0.066 ps=0.745 w=0.36 l=0.15
X2221 a_15832_5950# a_15666_5950# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2222 a_1247_2883# hgu_sarlogic_flat_0.x4.x9.S VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X2223 VSS hgu_cdac_half_1.db<5> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2224 hgu_vgen_vref_0.phi2_n a_n54752_6595# hgu_tah_0.VDD hgu_tah_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2225 hgu_tah_0.tah_vn hgu_tah_0.sw vin VSS sky130_fd_pr__nfet_01v8 ad=0.454 pd=3.08 as=0.454 ps=3.08 w=2.75 l=0.15
X2226 VSS a_12359_7798# a_12294_7824# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0935 ps=0.965 w=0.64 l=0.15
X2227 hgu_cdac_half_1.hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT hgu_cdac_half_1.db<2> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.122 ps=1.42 w=0.42 l=0.35
X2228 VSS hgu_cdac_half_0.d<6> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2229 a_1107_1331# a_1203_1153# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2230 a_n399_1179# a_n1189_1153# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0703 ps=0.755 w=0.42 l=0.15
X2231 a_4125_7798# a_4438_7824# a_4544_7824# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2232 a_1920_2150# a_1502_2234# a_1676_1842# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X2233 a_16427_5676# a_16581_5510# a_16287_5284# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2234 a_18923_5310# a_18505_5310# a_18679_5284# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X2235 a_n2785_7946# VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2236 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_1.db<5> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2237 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2238 VSS hgu_cdac_half_0.d<3> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<7:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2239 a_1247_2556# hgu_sarlogic_flat_0.x4.x9.S VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X2240 VSS VDD a_4544_7824# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.12 ps=1.08 w=0.42 l=0.15
X2241 hgu_vgen_vref_0.mimtop1 hgu_vgen_vref_0.mimbot1 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X2242 VDD a_11300_6052# hgu_sarlogic_flat_0.x3.x63.Q_N VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X2243 VDD a_17068_4644# a_16980_5036# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X2244 VSS a_4654_1153# a_4564_1179# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.116 ps=1.09 w=0.64 l=0.15
X2245 hgu_cdac_half_0.VREF hgu_cdac_half_0.db<5> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2246 VSS hgu_cdac_half_0.d<5> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2247 hgu_vgen_vref_0.mimtop1 hgu_vgen_vref_0.mimbot1 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X2248 hgu_cdac_half_0.VREF hgu_cdac_half_0.d<6> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2249 a_11070_2234# a_10624_1868# a_10978_1868# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0651 ps=0.73 w=0.42 l=0.15
X2250 VDD hgu_sarlogic_flat_0.x3.x30.Q_N a_7574_6052# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X2251 a_4001_13960# hgu_sarlogic_flat_0.x2.x3.A a_3929_13960# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X2252 VSS a_n53647_7835# a_n53834_7657# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X2253 hgu_cdac_half_0.VREF hgu_cdac_half_0.d<6> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2254 VDD VDD a_10771_1153# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0956 pd=0.875 as=0.132 ps=1.22 w=0.42 l=0.15
X2255 hgu_cdac_half_0.VREF hgu_cdac_half_0.db<6> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2256 a_10638_14236# hgu_sarlogic_flat_0.x2.x2.x1.IN a_10550_14098# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X2257 VSS hgu_comp_flat_0.clk a_n6959_12827# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X2258 VSS a_n6526_6819# a_n7760_6349# VSS sky130_fd_pr__nfet_01v8 ad=0.0759 pd=0.79 as=0.0759 ps=0.79 w=0.46 l=0.15
X2259 VSS a_n1699_7253# hgu_cdac_sw_buffer_2.x3.X VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X2260 VSS hgu_cdac_half_1.db<6> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2261 VSS a_2914_9360# hgu_sarlogic_flat_0.x5.eob VSS sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X2262 a_16531_6590# a_16113_6590# a_16287_6564# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X2263 a_4437_6078# hgu_sarlogic_flat_0.x3.x4.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2264 hgu_sarlogic_flat_0.x4.x3.X a_n1058_3698# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2265 VSS hgu_sarlogic_flat_0.x4.x5.D a_583_1179# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2266 hgu_vgen_vref_0.sky130_fd_sc_hd__inv_1_2.A hgu_vgen_vref_0.sky130_fd_sc_hd__inv_1_0.A hgu_tah_0.VDD hgu_tah_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2267 a_11774_6925# hgu_sarlogic_flat_0.x3.x39.Q_N VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X2268 a_1622_1179# a_1749_1347# a_1203_1153# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.03 as=0.0864 ps=0.91 w=0.64 l=0.15
X2269 hgu_cdac_half_0.VREF hgu_cdac_half_0.d<5> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2270 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<15:0> hgu_cdac_half_0.db<4> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2271 a_10478_6444# a_9966_6052# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X2272 hgu_sarlogic_flat_0.x2.x2.x4.x9.output_stack sample_delay_cap_ctrl_code[2] hgu_sarlogic_flat_0.x2.x2.x4.x4[3].floating VSS sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X2273 hgu_cdac_half_1.VREF hgu_cdac_half_1.d<6> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2274 a_2347_8513# a_2501_8487# a_2207_8487# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2275 hgu_cdac_half_1.VREF hgu_cdac_half_1.d<6> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2276 hgu_cdac_half_1.VREF hgu_cdac_half_1.db<6> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2277 VSS a_10164_8487# a_10871_8513# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X2278 a_11775_8487# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X2279 hgu_cdac_half_0.db<6> a_n1158_n1744# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2280 hgu_cdac_half_1.VREF hgu_cdac_half_1.db<6> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2281 a_9894_6951# a_9382_6925# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X2282 a_17184_5676# a_16581_5510# a_17068_5284# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2283 hgu_sarlogic_flat_0.x4.x9.A1 a_3960_3698# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2284 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2285 VSS a_5379_6925# a_5314_6951# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X2286 hgu_cdac_sw_buffer_1.VDD a_1196_n1740# hgu_cdac_half_0.d<6> hgu_cdac_sw_buffer_1.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2287 a_n6887_13761# hgu_comp_flat_0.ready a_n6959_13761# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X2288 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<15:0> hgu_cdac_half_0.db<4> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.122 ps=1.42 w=0.42 l=0.35
X2289 VDD hgu_sarlogic_flat_0.x1.x10.A a_n1149_11676# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0651 ps=0.73 w=0.42 l=0.15
X2290 a_1196_n1740# hgu_cdac_sw_buffer_1.x11.A VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2291 hgu_sarlogic_flat_0.x2.x2.x1.x5[7].floating hgu_sarlogic_flat_0.x2.x2.x1.x10.Y hgu_sarlogic_flat_0.x2.x2.x1.x9.output_stack VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X2292 a_n86_n245# hgu_cdac_sw_buffer_0.x4.A VSS VSS sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2293 VSS a_1945_10648# hgu_tah_0.sw_n VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2294 hgu_sarlogic_flat_0.x5.x1[3].Q_N a_19460_5924# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X2295 VSS hgu_cdac_half_0.db<6> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2296 VDD a_2444_2136# a_2369_2234# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0956 pd=0.875 as=0.0787 ps=0.795 w=0.42 l=0.15
X2297 VDD a_52_2136# a_773_1868# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X2298 VDD a_n542_11334# hgu_sarlogic_flat_0.x1.x3.A0 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X2299 VDD sample_delay_cap_ctrl_code[11] hgu_sarlogic_flat_0.x2.x2.x2.x10.Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2300 a_10235_8008# a_9762_8098# a_10479_7824# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0671 ps=0.75 w=0.36 l=0.15
X2301 hgu_sarlogic_flat_0.x2.x1.x4.Y VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2302 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2303 hgu_cdac_half_0.d<6> a_1196_n1740# hgu_cdac_sw_buffer_1.VDD hgu_cdac_sw_buffer_1.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2304 VSS hgu_sarlogic_flat_0.x2.x2.x2.IN a_16448_15176# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0651 ps=0.73 w=0.42 l=0.15
X2305 hgu_cdac_half_1.VREF hgu_cdac_half_1.d<3> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<7:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2306 a_5176_2883# VSS a_5176_2556# VSS sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X2307 a_9847_7233# a_9382_6925# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X2308 VSS hgu_cdac_half_0.d<5> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2309 VSS hgu_cdac_half_0.db<5> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2310 a_16041_11987# hgu_sarlogic_flat_0.x2.x2.x2.IN a_15953_11987# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X2311 hgu_tah_0.VDD hgu_vgen_vref_0.sky130_fd_sc_hd__inv_1_4.Y hgu_vgen_vref_0.sky130_fd_sc_hd__nand2_1_1.Y hgu_tah_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2312 VDD a_n7390_7871# a_n7766_6446# VDD sky130_fd_pr__pfet_01v8 ad=0.139 pd=1.17 as=0.26 ps=2.3 w=0.84 l=0.15
X2313 hgu_sarlogic_flat_0.x4.x13.S a_13263_8513# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X2314 VDD hgu_sarlogic_flat_0.x3.x7.X a_13072_6078# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0662 ps=0.735 w=0.42 l=0.15
X2315 a_2530_1363# a_2057_1453# a_2774_1179# VSS sky130_fd_pr__nfet_01v8 ad=0.0675 pd=0.735 as=0.0671 ps=0.75 w=0.36 l=0.15
X2316 VDD a_621_10615# a_651_10968# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X2317 a_8289_7824# a_7370_8098# a_7843_8008# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X2318 a_10103_7824# a_10235_8008# a_9967_7798# VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0864 ps=0.91 w=0.64 l=0.15
X2319 a_9901_6078# a_9761_6352# a_9463_6052# VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.0711 ps=0.755 w=0.36 l=0.15
X2320 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.db<6> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2321 a_11488_2150# a_11070_2234# a_11244_1842# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X2322 hgu_sarlogic_flat_0.x4.x25.Q_N a_7228_2136# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X2323 a_9848_8795# a_9383_8487# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X2324 VSS a_n1749_7728# hgu_cdac_half_1.d<5> VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2325 a_2036_7824# hgu_sarlogic_flat_0.x3.x4.A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2326 hgu_sarlogic_flat_0.x1.x4.x9.output_stack hgu_sarlogic_flat_0.x1.x4.x6.SW hgu_sarlogic_flat_0.x1.x4.x6.floating VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X2327 hgu_sarlogic_flat_0.x3.x4.X a_2036_7824# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2328 a_2398_1179# a_2530_1363# a_2262_1153# VSS sky130_fd_pr__nfet_01v8 ad=0.0974 pd=0.97 as=0.0864 ps=0.91 w=0.64 l=0.15
X2329 hgu_cdac_half_1.d<0> a_15125_1868# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X2330 a_8852_1842# a_8678_2234# a_8996_1868# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.0974 ps=0.97 w=0.64 l=0.15
X2331 hgu_comp_flat_0.Q hgu_comp_flat_0.clk VDD VDD sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X2332 VSS a_3960_3698# hgu_sarlogic_flat_0.x4.x9.A1 VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2333 hgu_cdac_sw_buffer_0.VDD a_n1158_n1744# hgu_cdac_half_0.db<6> hgu_cdac_sw_buffer_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2334 VDD a_3326_3698# hgu_sarlogic_flat_0.x4.x30.A VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2335 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<15:0> hgu_cdac_half_0.db<4> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2336 hgu_cdac_half_1.VREF hgu_cdac_half_1.d<5> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2337 VSS hgu_comp_flat_0.RS_p a_n7216_6420# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X2338 a_n1149_11335# hgu_sarlogic_flat_0.x1.x4.x9.output_stack hgu_sarlogic_flat_0.x1.x10.A VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.122 ps=1.42 w=0.42 l=0.15
X2339 VSS VDD a_13930_1842# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X2340 hgu_tah_0.VDD a_n54567_7835# a_n54754_7657# hgu_tah_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X2341 hgu_cdac_half_0.VREF hgu_cdac_half_0.d<6> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2342 a_454_n939# VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2343 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<0> hgu_cdac_half_0.db<0> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.244 ps=2.26 w=0.84 l=0.35
X2344 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_1.d<5> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2345 a_n6526_6819# a_n6676_7789# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0.244 ps=2.26 w=0.84 l=0.15
X2346 a_18679_5284# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X2347 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<7:0> hgu_cdac_half_0.d<3> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2348 VDD a_n3877_7252# hgu_cdac_sw_buffer_3.x3.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X2349 VDD a_1454_6950# hgu_sarlogic_flat_0.x3.x7.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2350 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_0.d<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2351 VSS hgu_cdac_half_0.d<4> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<15:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2352 hgu_cdac_half_1.VREF hgu_cdac_half_1.db<5> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2353 a_2521_6078# a_1732_6052# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0588 ps=0.7 w=0.42 l=0.15
X2354 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X2355 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.d<6> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2356 hgu_cdac_half_0.VREF hgu_cdac_half_0.d<3> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<7:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2357 a_9332_12263# hgu_sarlogic_flat_0.x2.x2.x3.IN a_9244_12263# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X2358 hgu_sarlogic_flat_0.x5.x2.x3[1].floating retimer_delay_code[1] hgu_sarlogic_flat_0.x5.x2.x9.output_stack VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X2359 VSS a_n54284_7371# a_n54471_7113# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X2360 a_18679_5924# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X2361 VSS hgu_cdac_half_0.db<6> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2362 hgu_cdac_half_0.VREF hgu_cdac_half_0.d<5> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2363 a_2195_1545# a_2058_1153# a_1749_1347# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X2364 a_6536_8513# a_6370_8513# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2365 hgu_sarlogic_flat_0.x4.x9.A1 a_3960_3698# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2366 hgu_cdac_sw_buffer_1.x11.A a_1114_n1100# hgu_cdac_sw_buffer_1.VDD hgu_cdac_sw_buffer_1.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2367 hgu_sarlogic_flat_0.x1.x4.x9.output_stack hgu_comp_flat_0.clk a_n7022_10886# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X2368 a_7370_6052# hgu_sarlogic_flat_0.x4.D[4] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2369 hgu_cdac_sw_buffer_0.VDD a_n1158_n1744# hgu_cdac_half_0.db<6> hgu_cdac_sw_buffer_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2370 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<15:0> hgu_cdac_half_0.db<4> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2371 a_9760_1868# a_9146_1842# a_9620_2136# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2372 a_9739_14835# hgu_sarlogic_flat_0.x2.x2.x4.x9.output_stack hgu_sarlogic_flat_0.x2.x2.x1.IN VSS sky130_fd_pr__nfet_01v8 ad=0.0651 pd=0.73 as=0.122 ps=1.42 w=0.42 l=0.15
X2373 VSS hgu_sarlogic_flat_0.x3.x5.X a_6370_8513# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2374 a_7558_1545# a_7046_1153# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X2375 VSS hgu_cdac_half_1.d<5> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2376 VDD a_16581_5924# a_16531_6232# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X2377 a_19694_5310# a_19286_5688# a_19460_5284# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X2378 a_11600_7317# a_11319_6951# a_11507_6951# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X2379 VSS hgu_sarlogic_flat_0.x5.x3.X a_15666_4670# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2380 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_0.db<5> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.35
X2381 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_1.db<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2382 a_n6676_7789# hgu_comp_flat_0.clk VDD VDD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X2383 VSS a_8281_2708# hgu_sarlogic_flat_0.x4.x14.X VSS sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X2384 hgu_cdac_half_1.VREF hgu_cdac_half_1.d<6> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2385 VSS hgu_cdac_half_1.db<4> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<15:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.35
X2386 VSS hgu_sarlogic_flat_0.x5.x3.X a_15666_5316# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2387 a_17302_4952# a_16894_4670# a_17068_4644# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X2388 a_n4397_8367# hgu_cdac_sw_buffer_3.x11.A VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2389 hgu_cdac_half_0.db<6> a_n1158_n1744# hgu_cdac_sw_buffer_0.VDD hgu_cdac_sw_buffer_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2390 hgu_cdac_half_1.VREF hgu_cdac_half_1.d<6> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2391 VDD a_6517_7798# hgu_sarlogic_flat_0.x3.x45.Q_N VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X2392 a_2104_15080# a_1592_14732# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X2393 a_11601_8879# a_11320_8513# a_11508_8513# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X2394 hgu_cdac_sw_buffer_1.VDD VSS a_1942_n460# hgu_cdac_sw_buffer_1.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X2395 hgu_sarlogic_flat_0.x1.x4.x9.output_stack hgu_sarlogic_flat_0.x1.x4.x10.Y hgu_sarlogic_flat_0.x1.x4.x5[7].floating VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X2396 a_5613_7233# a_5205_6951# a_5379_6925# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X2397 VSS hgu_cdac_half_0.db<6> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2398 hgu_cdac_half_1.d<5> a_n1749_7728# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2399 a_18679_5284# a_18505_5310# a_18819_5676# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X2400 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.db<6> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2401 a_16088_10874# hgu_sarlogic_flat_0.x2.x2.x2.IN hgu_sarlogic_flat_0.x2.x2.x2.x9.output_stack VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X2402 hgu_vgen_vref_0.sky130_fd_sc_hd__inv_1_3.Y hgu_vgen_vref_0.sky130_fd_sc_hd__inv_1_3.A hgu_tah_0.VDD hgu_tah_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2403 a_n1158_n1744# hgu_cdac_sw_buffer_0.x11.A VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2404 a_11914_6951# hgu_sarlogic_flat_0.x3.x39.Q_N VSS VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X2405 a_12098_1363# a_11625_1453# a_12342_1179# VSS sky130_fd_pr__nfet_01v8 ad=0.0675 pd=0.735 as=0.0671 ps=0.75 w=0.36 l=0.15
X2406 a_9115_6951# hgu_sarlogic_flat_0.x3.x7.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X2407 a_6348_2883# hgu_sarlogic_flat_0.x4.x9.A1 a_5889_2708# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X2408 VDD a_1203_1153# hgu_sarlogic_flat_0.x4.x21.Q_N VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X2409 VDD VSS a_3977_6951# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2410 a_5614_8795# a_5206_8513# a_5380_8487# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X2411 a_n595_7253# hgu_cdac_sw_buffer_2.x5.A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X2412 VSS VDD a_9574_1179# VSS sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0974 ps=0.97 w=0.42 l=0.15
X2413 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X2414 hgu_sarlogic_flat_0.x5.x2.x9.output_stack retimer_delay_code[1] hgu_sarlogic_flat_0.x5.x2.x3[1].floating VSS sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X2415 hgu_cdac_half_1.d<4> a_n1209_7728# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2416 hgu_tah_0.tah_vn hgu_tah_0.sw_n vin hgu_tah_0.VDD sky130_fd_pr__pfet_01v8 ad=0.908 pd=5.83 as=0.908 ps=5.83 w=5.5 l=0.15
X2417 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X2418 VSS hgu_cdac_half_1.d<6> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2419 a_4637_6360# a_4437_6078# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X2420 VSS a_6318_2530# a_6252_2556# VSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X2421 hgu_sarlogic_flat_0.x2.x2.x1.x9.output_stack sample_delay_cap_ctrl_code[5] hgu_sarlogic_flat_0.x2.x2.x1.x3[1].floating VSS sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X2422 a_9116_8513# hgu_sarlogic_flat_0.x4.x9.S VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X2423 VDD hgu_sarlogic_flat_0.x3.x7.X a_10680_6078# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0662 ps=0.735 w=0.42 l=0.15
X2424 a_n130_1153# a_138_1363# a_84_1461# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X2425 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X2426 hgu_vgen_vref_0.mimtop2 VSS sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X2427 hgu_tah_0.sw a_1945_11268# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X2428 VSS a_3960_3698# hgu_sarlogic_flat_0.x4.x9.A1 VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2429 VSS hgu_cdac_half_0.db<1> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<1:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.35
X2430 a_5315_8513# a_3978_8513# a_5206_8513# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X2431 hgu_cdac_half_0.VREF hgu_cdac_half_0.d<5> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2432 VSS hgu_cdac_half_1.db<6> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2433 hgu_sarlogic_flat_0.x3.D[0] a_8478_6951# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X2434 hgu_cdac_half_0.hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT hgu_cdac_half_0.d<2> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2435 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.db<6> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2436 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.db<6> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2437 hgu_sarlogic_flat_0.x1.x2.x5[7].floating hgu_sarlogic_flat_0.x1.x2.x10.Y hgu_sarlogic_flat_0.x1.x2.x9.output_stack VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X2438 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<15:0> hgu_cdac_half_0.db<4> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2439 hgu_cdac_half_1.d<1> a_12733_1868# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X2440 a_6460_1842# a_6286_2234# a_6604_1868# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.0974 ps=0.97 w=0.64 l=0.15
X2441 a_4599_8487# a_4425_8879# a_4739_8513# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X2442 a_1586_2234# a_1222_1868# a_1502_2234# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X2443 hgu_cdac_half_1.d<6> a_n2219_8368# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2444 VSS a_2820_n241# hgu_cdac_half_0.d<2> VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X2445 a_7306_7824# a_6517_7798# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0588 ps=0.7 w=0.42 l=0.15
X2446 VSS hgu_cdac_half_0.d<6> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2447 hgu_sarlogic_flat_0.x4.x9.S a_8479_8513# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X2448 a_7130_6951# a_7284_6925# a_6990_6925# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2449 a_13072_6078# a_12154_6052# a_12626_6262# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2450 a_12089_6078# a_11300_6052# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0588 ps=0.7 w=0.42 l=0.15
X2451 hgu_sarlogic_flat_0.x2.x2.x4.x9.output_stack sample_delay_cap_ctrl_code[2] hgu_sarlogic_flat_0.x2.x2.x4.x4[3].floating VSS sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X2452 a_12018_7233# a_11600_7317# a_11774_6925# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X2453 hgu_comp_flat_0.Q hgu_tah_0.tah_vn a_n7660_7467# VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X2454 VDD a_1945_11268# hgu_tah_0.sw VDD sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.391 ps=3.14 w=1.26 l=0.15
X2455 a_3898_9386# sel_bit[1] a_2914_9360# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X2456 hgu_sarlogic_flat_0.x2.x2.x1.x9.output_stack hgu_sarlogic_flat_0.x2.x2.x1.IN a_10638_14788# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X2457 a_6394_1868# a_5840_1868# a_6286_2234# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0675 ps=0.735 w=0.36 l=0.15
X2458 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_1.d<5> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2459 result[5] a_20167_5326# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X2460 hgu_cdac_half_0.VREF hgu_cdac_half_0.db<5> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2461 a_18505_5310# a_18224_5316# a_18412_5310# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X2462 VSS hgu_cdac_half_0.db<6> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2463 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<7:0> hgu_cdac_half_1.db<3> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2464 a_4332_8513# hgu_sarlogic_flat_0.x3.x27.D VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X2465 a_4508_7317# a_3977_6951# a_4424_7317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X2466 a_n86_n245# hgu_cdac_sw_buffer_0.x4.A hgu_cdac_sw_buffer_0.VDD hgu_cdac_sw_buffer_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X2467 a_12019_8795# a_11601_8879# a_11775_8487# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X2468 hgu_comp_flat_0.comp_outn a_n6292_6446# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.139 pd=1.17 as=0.26 ps=2.3 w=0.84 l=0.15
X2469 VDD a_n130_1153# a_n197_1545# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X2470 a_18505_6316# a_18224_5950# a_18412_5950# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X2471 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X2472 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<7:0> hgu_cdac_half_0.d<3> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2473 hgu_sarlogic_flat_0.x3.x7.A a_1178_6950# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X2474 VSS a_17068_4644# a_17003_4670# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X2475 a_16287_6564# a_16113_6590# a_16427_6956# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X2476 VSS hgu_cdac_sw_buffer_0.x11.A a_n1158_n1744# VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2477 a_12626_6262# a_12154_6052# a_12870_6444# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X2478 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_0.d<5> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2479 hgu_cdac_half_0.VREF hgu_cdac_half_0.d<4> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<15:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2480 hgu_cdac_sw_buffer_0.VDD a_n1240_n1104# hgu_cdac_sw_buffer_0.x11.A hgu_cdac_sw_buffer_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2481 a_2607_14758# a_2199_15136# a_2373_14732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X2482 VSS a_17068_5284# a_17003_5688# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X2483 a_4509_8879# a_3978_8513# a_4425_8879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X2484 VDD hgu_cdac_sw_buffer_3.x4.X a_n3387_7727# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2485 a_16448_14835# hgu_sarlogic_flat_0.x2.x2.x2.IN VDD VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2486 VDD hgu_sarlogic_flat_0.x5.x3.A a_20464_8538# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0651 ps=0.73 w=0.42 l=0.15
X2487 VSS hgu_cdac_sw_buffer_2.x9.X a_n2301_7728# VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2488 VDD hgu_sarlogic_flat_0.x4.D[6] a_2975_1179# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X2489 a_10183_2556# hgu_sarlogic_flat_0.x4.x9.A1 a_9962_2883# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X2490 a_9332_12539# hgu_sarlogic_flat_0.x2.x2.x3.IN a_9244_12539# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X2491 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X2492 VDD a_n1209_7728# hgu_cdac_half_1.d<4> VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2493 a_16799_5632# a_16287_5284# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X2494 VSS a_5889_2708# hgu_sarlogic_flat_0.x4.x12.X VSS sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X2495 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<15:0> hgu_cdac_half_1.d<4> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2496 a_3898_9386# a_3783_9360# a_2914_9360# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.6 as=0.0729 ps=0.81 w=0.54 l=0.15
X2497 a_3960_3698# hgu_sarlogic_flat_0.x4.x30.A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2498 hgu_sarlogic_flat_0.x4.x2.X a_n424_3698# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2499 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_0.db<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2500 hgu_vgen_vref_0.mimtop1 hgu_vgen_vref_0.mimbot1 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X2501 VDD a_n1285_1331# hgu_cdac_sw_buffer_3.x9.A VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X2502 VSS hgu_cdac_half_1.db<6> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2503 a_12240_8795# a_11775_8487# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X2504 a_18819_5950# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X2505 a_7887_6951# a_7284_6925# a_7771_6925# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2506 VDD hgu_sarlogic_flat_0.x3.x5.X a_3978_8513# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2507 hgu_vgen_vref_0.sky130_fd_sc_hd__nand2_1_0.Y hgu_vgen_vref_0.clk a_n53010_7683# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2508 a_18819_6956# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X2509 hgu_sarlogic_flat_0.x3.x4.X a_2036_7824# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2510 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.d<6> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2511 hgu_sarlogic_flat_0.x2.x7.A hgu_sarlogic_flat_0.x2.x2.x3.x9.output_stack a_3314_11664# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0651 ps=0.73 w=0.42 l=0.15
X2512 VSS hgu_sarlogic_flat_0.x3.x4.X a_12068_6925# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X2513 hgu_cdac_half_1.VREF hgu_cdac_half_1.db<4> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<15:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2514 hgu_cdac_half_0.db<5> a_n688_n1104# hgu_cdac_sw_buffer_0.VDD hgu_cdac_sw_buffer_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2515 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.db<6> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2516 VSS a_n2219_8368# hgu_cdac_half_1.d<6> VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2517 VDD a_14017_1453# a_14018_1153# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2518 a_12352_2883# VSS a_12352_2556# VSS sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X2519 hgu_cdac_half_0.VREF hgu_cdac_half_0.db<6> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2520 hgu_vgen_vref_0.phi1_n a_n54752_8227# hgu_tah_0.VDD hgu_tah_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2521 a_7370_6052# hgu_sarlogic_flat_0.x4.D[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2522 VSS hgu_cdac_half_0.db<6> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2523 a_3956_2883# hgu_sarlogic_flat_0.x4.x9.A1 a_3497_2708# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X2524 VSS a_n4397_8367# hgu_cdac_sw_buffer_3.x11.X VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2525 a_6723_6951# hgu_sarlogic_flat_0.x3.x7.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X2526 VDD a_18973_6790# a_19694_6590# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X2527 VSS hgu_cdac_half_0.db<4> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<15:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2528 hgu_cdac_sw_buffer_3.x11.X a_n4397_8367# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2529 hgu_vgen_vref_0.phi2_n a_n54752_6595# hgu_tah_0.VDD hgu_tah_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2530 VSS a_3926_2530# a_3860_2556# VSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X2531 VSS hgu_cdac_half_1.d<6> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2532 a_6724_8513# hgu_sarlogic_flat_0.x4.x7.S VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X2533 result[6] a_17775_4670# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X2534 VDD async_delay_offset hgu_sarlogic_flat_0.x1.x2.x6.SW VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2535 VSS a_n424_3698# hgu_sarlogic_flat_0.x4.x2.X VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2536 a_4580_1868# a_4068_1842# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.116 pd=1.09 as=0.166 ps=1.8 w=0.64 l=0.15
X2537 a_8379_1153# a_8925_1347# a_8883_1461# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.132 pd=1.22 as=0.0882 ps=1.05 w=0.84 l=0.15
X2538 VDD a_6460_1842# a_6370_2234# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X2539 hgu_sarlogic_flat_0.x5.x2.x9.output_stack hgu_sarlogic_flat_0.x5.eob a_14591_9328# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X2540 a_2923_8513# a_1586_8513# a_2814_8513# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X2541 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_0.db<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2542 VSS hgu_cdac_half_1.db<6> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.35
X2543 a_19191_5950# a_18679_5924# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X2544 hgu_cdac_half_0.VREF hgu_cdac_half_0.db<5> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2545 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2546 a_9379_10874# hgu_sarlogic_flat_0.x2.x2.x3.IN a_9291_10736# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X2547 VSS VDD a_11966_1179# VSS sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0974 ps=0.97 w=0.42 l=0.15
X2548 hgu_cdac_half_0.VREF hgu_cdac_half_0.db<6> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.35
X2549 VDD VDD a_18973_5510# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X2550 hgu_cdac_half_0.hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT hgu_cdac_half_0.d<2> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2551 hgu_sarlogic_flat_0.x2.x2.x2.x9.output_stack sample_delay_cap_ctrl_code[9] hgu_sarlogic_flat_0.x2.x2.x2.x3[1].floating VSS sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X2552 a_4914_7824# a_4125_7798# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0588 ps=0.7 w=0.42 l=0.15
X2553 VSS a_19460_5924# a_20167_5950# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X2554 a_9169_1179# a_8379_1153# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0703 ps=0.755 w=0.42 l=0.15
X2555 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_1.db<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2556 hgu_cdac_sw_buffer_2.x11.A a_n2301_7728# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2557 a_4738_6951# a_4892_6925# a_4598_6925# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2558 a_10680_6078# a_9762_6052# a_10234_6262# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2559 VSS hgu_sarlogic_flat_0.x5.x3.A a_20768_8628# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X2560 hgu_vgen_vref_0.mimtop1 hgu_vgen_vref_0.mimbot1 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X2561 hgu_tah_0.VDD a_n53930_7371# hgu_vgen_vref_0.sky130_fd_sc_hd__dlymetal6s6s_1_4.A hgu_tah_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X2562 VDD a_9382_6925# a_9292_7317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X2563 VSS a_19460_6564# a_20167_6606# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X2564 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_1.d<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.122 ps=1.42 w=0.42 l=0.35
X2565 a_3929_14374# hgu_sarlogic_flat_0.x2.x3.A a_3841_14374# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X2566 a_5896_6078# a_4977_6352# a_5450_6262# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X2567 hgu_cdac_half_0.VREF hgu_cdac_half_0.db<5> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2568 hgu_sarlogic_flat_0.x4.x3.X a_n1058_3698# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2569 hgu_cdac_sw_buffer_0.x12.X a_n412_n464# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2570 hgu_cdac_half_0.VREF hgu_cdac_half_0.d<6> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2571 a_n7766_6446# a_n7390_7871# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0759 pd=0.79 as=0.0759 ps=0.79 w=0.46 l=0.15
X2572 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X2573 a_4002_1868# a_3448_1868# a_3894_2234# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0675 ps=0.735 w=0.36 l=0.15
X2574 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.d<6> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2575 VSS a_1114_n1100# hgu_cdac_sw_buffer_1.x11.A VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2576 a_19144_6232# a_18679_5924# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X2577 hgu_cdac_sw_buffer_1.x8.X a_1390_n460# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2578 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.db<6> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2579 VSS a_5380_8487# a_5315_8513# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X2580 VSS a_n7390_7871# hgu_comp_flat_0.RS_p VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.15
X2581 hgu_sarlogic_flat_0.x1.x4.x9.output_stack hgu_sarlogic_flat_0.x1.x4.x10.Y hgu_sarlogic_flat_0.x1.x4.x5[7].floating VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X2582 a_1940_8513# hgu_sarlogic_flat_0.x5.eob VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X2583 VDD a_9383_8487# a_9293_8879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X2584 hgu_sarlogic_flat_0.x4.x9.A1 a_3960_3698# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2585 a_4001_14236# hgu_sarlogic_flat_0.x2.x3.A a_3929_14236# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X2586 hgu_sarlogic_flat_0.x3.x20.Q_N a_2988_8487# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X2587 a_4425_8879# a_3978_8513# a_4332_8513# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X2588 a_407_11578# hgu_tah_0.sw VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2589 VSS a_8908_6052# hgu_sarlogic_flat_0.x3.x60.Q_N VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X2590 a_18613_5950# a_18224_5950# a_18505_6316# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X2591 hgu_cdac_half_0.db<6> a_n1158_n1744# hgu_cdac_sw_buffer_0.VDD hgu_cdac_sw_buffer_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2592 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_0.d<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.122 ps=1.42 w=0.42 l=0.35
X2593 hgu_tah_0.VDD a_n55487_7371# a_n55674_7113# hgu_tah_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X2594 hgu_sarlogic_flat_0.x5.x1[0].Q_N a_17068_6564# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X2595 hgu_vgen_vref_0.mimtop2 VSS sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X2596 hgu_sarlogic_flat_0.x3.x7.A a_1178_6950# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2597 VSS a_4599_8487# a_4533_8513# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X2598 a_2036_7824# hgu_sarlogic_flat_0.x3.x4.A VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2599 hgu_cdac_half_1.VREF hgu_cdac_half_1.db<6> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2600 hgu_sarlogic_flat_0.x2.x2.x2.x7.floating sample_delay_offset hgu_sarlogic_flat_0.x2.x2.x2.x9.output_stack VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X2601 VSS a_n2219_8368# hgu_cdac_half_1.d<6> VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2602 VSS hgu_sarlogic_flat_0.x4.x30.A a_3960_3698# VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2603 a_7072_7798# a_7371_7798# a_7306_7824# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.066 ps=0.745 w=0.36 l=0.15
X2604 VDD a_n2251_7253# hgu_cdac_sw_buffer_2.x9.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X2605 result[0] a_17775_6606# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X2606 VSS a_n2219_8368# hgu_cdac_half_1.d<6> VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2607 a_11855_6052# a_12154_6052# a_12089_6078# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.066 ps=0.745 w=0.36 l=0.15
X2608 hgu_cdac_half_0.VREF hgu_cdac_half_0.db<3> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<7:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2609 VSS hgu_cdac_half_1.d<6> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2610 a_1019_10793# VSS a_1161_10641# VSS sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X2611 hgu_cdac_sw_buffer_0.VDD a_n1158_n1744# hgu_cdac_half_0.db<6> hgu_cdac_sw_buffer_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2612 a_12789_7233# a_12381_6951# a_12555_6925# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X2613 a_13370_1868# hgu_sarlogic_flat_0.x4.D[1] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X2614 a_5104_2883# a_4922_2883# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X2615 a_5495_6951# hgu_sarlogic_flat_0.x3.x77.Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X2616 VDD a_1592_14732# a_1502_14758# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X2617 a_9404_12677# hgu_sarlogic_flat_0.x2.x2.x3.IN a_9332_12815# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X2618 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2619 a_5495_6951# a_4892_6925# a_5379_6925# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2620 hgu_vgen_vref_0.mimtop2 VSS sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X2621 hgu_sarlogic_flat_0.x1.x10.Y hgu_sarlogic_flat_0.x1.x10.A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2622 a_n6887_14037# hgu_comp_flat_0.ready a_n6959_14037# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X2623 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2624 VSS a_n4397_8367# hgu_cdac_sw_buffer_3.x11.X VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2625 a_n4397_8367# hgu_cdac_sw_buffer_3.x11.A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2626 a_19460_5924# a_19286_5950# a_19576_5950# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X2627 hgu_vgen_vref_0.mimtop2 VSS sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X2628 hgu_cdac_half_0.VREF hgu_cdac_half_0.db<6> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2629 VDD a_11625_1453# a_11626_1153# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2630 VSS hgu_cdac_half_0.d<5> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2631 VDD VDD a_16581_6790# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X2632 a_14148_1868# a_13636_1842# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.116 pd=1.09 as=0.166 ps=1.8 w=0.64 l=0.15
X2633 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X2634 VSS hgu_cdac_half_1.db<4> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<15:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2635 hgu_tah_0.VDD VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X2636 a_16113_12125# hgu_sarlogic_flat_0.x2.x2.x2.IN a_16041_12263# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X2637 VSS VDD a_18973_4644# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X2638 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X2639 VDD a_1886_14958# a_2607_14758# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X2640 VSS VDD a_18973_5510# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X2641 a_9115_6951# hgu_sarlogic_flat_0.x3.x7.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X2642 VDD hgu_sarlogic_flat_0.x4.x27.A a_3326_3698# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2643 hgu_sarlogic_flat_0.x5.eob a_2914_9360# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X2644 a_13636_1842# a_13462_2234# a_13780_1868# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.0974 ps=0.97 w=0.64 l=0.15
X2645 hgu_vgen_vref_0.mimtop1 hgu_vgen_vref_0.mimbot1 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X2646 VDD a_19460_5924# a_20167_5950# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X2647 hgu_vgen_vref_0.mimtop1 hgu_vgen_vref_0.mimbot1 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X2648 a_7759_1179# a_6842_1153# a_7314_1363# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0675 ps=0.735 w=0.36 l=0.15
X2649 hgu_sarlogic_flat_0.x3.x5.X a_1863_9386# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2650 hgu_cdac_half_0.VREF hgu_cdac_half_0.db<5> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.35
X2651 hgu_vgen_vref_0.mimtop1 hgu_vgen_vref_0.phi2_n hgu_tah_0.VDD hgu_tah_0.VDD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=0.5
X2652 a_20464_8879# hgu_sarlogic_flat_0.x5.x3.A VSS VDD sky130_fd_pr__pfet_01v8_hvt ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2653 a_16197_5036# a_15666_4670# a_16113_5036# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X2654 VSS a_14017_1453# a_14018_1153# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2655 VSS a_52_2136# a_0_1868# VSS sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.066 ps=0.745 w=0.42 l=0.15
X2656 VSS a_n53930_7835# hgu_vgen_vref_0.sky130_fd_sc_hd__dlymetal6s6s_1_2.A VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X2657 VSS hgu_cdac_half_0.db<6> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2658 a_9890_2883# a_9708_2883# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X2659 VDD a_1454_6950# hgu_sarlogic_flat_0.x3.x7.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2660 VSS a_n3877_7252# hgu_cdac_sw_buffer_3.x3.X VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X2661 a_6777_1179# a_5987_1153# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0703 ps=0.755 w=0.42 l=0.15
X2662 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_1.d<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2663 hgu_vgen_vref_0.mimtop2 VSS sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X2664 hgu_cdac_half_1.VREF hgu_cdac_half_1.d<6> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.35
X2665 hgu_sarlogic_flat_0.x3.x4.X a_2036_7824# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2666 VDD a_6990_6925# a_6900_7317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X2667 hgu_sarlogic_flat_0.x4.x9.A1 a_3960_3698# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2668 hgu_sarlogic_flat_0.x4.x7.X a_394_2883# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.158 ps=1.39 w=1 l=0.15
X2669 VSS hgu_cdac_half_0.d<6> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2670 VSS hgu_vgen_vref_0.sky130_fd_sc_hd__inv_1_3.Y a_n54752_6595# VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2671 VDD hgu_sarlogic_flat_0.x3.x27.Q_N a_5182_6052# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X2672 hgu_cdac_sw_buffer_1.VDD a_1196_n1740# hgu_cdac_half_0.d<6> hgu_cdac_sw_buffer_1.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2673 VDD hgu_sarlogic_flat_0.x2.x2.x2.x9.output_stack a_10023_11461# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X2674 VSS hgu_cdac_half_0.d<4> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<15:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.35
X2675 VSS hgu_cdac_half_1.db<5> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2676 VSS a_n55487_7835# a_n55674_7657# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X2677 hgu_cdac_half_0.d<6> a_1196_n1740# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2678 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.db<6> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2679 a_n1149_11676# hgu_sarlogic_flat_0.x1.x4.x9.output_stack VSS VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X2680 a_16752_6232# a_16287_5924# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X2681 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2682 a_n107_2234# a_n1336_1868# a_n204_1868# VSS sky130_fd_pr__nfet_01v8 ad=0.0486 pd=0.63 as=0.116 ps=1.09 w=0.36 l=0.15
X2683 VDD a_6991_8487# a_6901_8879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X2684 VDD hgu_sarlogic_flat_0.x4.D[3] a_10151_1179# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X2685 hgu_vgen_vref_0.phi2 a_n55304_6595# hgu_tah_0.VDD hgu_tah_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2686 VDD a_11102_2530# a_11132_2883# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X2687 a_16531_5310# a_16113_5310# a_16287_5284# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X2688 VDD VDD a_14222_1153# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X2689 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_1.db<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2690 hgu_vgen_vref_0.sky130_fd_sc_hd__inv_1_2.Y hgu_vgen_vref_0.sky130_fd_sc_hd__inv_1_2.A hgu_tah_0.VDD hgu_tah_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2691 a_10663_15763# hgu_sarlogic_flat_0.x2.x2.x1.IN a_10575_15625# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X2692 VDD a_2323_11578# a_1945_11268# VDD sky130_fd_pr__pfet_01v8 ad=0.365 pd=3.1 as=0.365 ps=3.1 w=1.26 l=0.15
X2693 VSS a_n7216_6420# hgu_comp_flat_0.comp_outp VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.54 as=0.0759 ps=0.79 w=0.46 l=0.15
X2694 a_3058_6262# a_2586_6052# a_3302_6444# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X2695 result[3] a_20167_5950# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X2696 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_0.d<5> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.35
X2697 a_8925_1347# a_9234_1153# a_9169_1179# VSS sky130_fd_pr__nfet_01v8 ad=0.0486 pd=0.63 as=0.066 ps=0.745 w=0.36 l=0.15
X2698 hgu_sarlogic_flat_0.x2.x2.x1.x10.Y sample_delay_cap_ctrl_code[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2699 hgu_cdac_half_1.VREF hgu_cdac_half_1.db<5> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2700 a_16088_10598# hgu_sarlogic_flat_0.x2.x2.x2.IN a_16000_10460# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X2701 a_14960_2883# VSS a_14746_2883# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.193 ps=1.34 w=0.42 l=0.15
X2702 VDD VSS a_n2025_7088# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X2703 VDD hgu_sarlogic_flat_0.x3.x5.X a_11154_8513# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2704 a_18412_4670# hgu_sarlogic_flat_0.x4.x5.D VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X2705 a_n685_1461# a_n876_1179# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X2706 VSS hgu_cdac_half_1.d<6> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2707 VSS VDD a_16581_5924# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X2708 VDD a_9146_1842# a_9877_2150# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X2709 hgu_sarlogic_flat_0.x2.x2.x3.x9.output_stack hgu_sarlogic_flat_0.x2.x2.x3.x10.Y hgu_sarlogic_flat_0.x2.x2.x3.x5[7].floating VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X2710 a_14726_8215# hgu_sarlogic_flat_0.x5.eob a_14654_8215# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X2711 VDD a_12154_6052# a_12153_6352# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2712 VSS a_n1190_n245# hgu_cdac_sw_buffer_0.x9.X VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X2713 a_14404_2136# a_14245_2234# a_14544_1868# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.109 ps=1.03 w=0.64 l=0.15
X2714 a_n251_2150# a_n716_1842# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X2715 a_10638_14650# hgu_sarlogic_flat_0.x2.x2.x1.IN a_10550_14650# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X2716 VSS VSS a_n1473_7088# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X2717 VSS VDD a_16581_6790# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X2718 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X2719 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2720 a_n6934_15564# hgu_comp_flat_0.ready a_n7022_15426# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X2721 hgu_cdac_half_1.VREF hgu_cdac_half_1.d<3> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<7:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2722 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2723 a_9221_6078# hgu_sarlogic_flat_0.x3.x4.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2724 a_2451_8795# a_2033_8879# a_2207_8487# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X2725 VSS a_1448_10615# a_1382_10641# VSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X2726 hgu_sarlogic_flat_0.x1.x9.Y hgu_sarlogic_flat_0.x1.x9.A VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2727 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2728 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.db<6> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2729 VSS hgu_cdac_half_1.d<6> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2730 VDD a_n607_7947# hgu_cdac_sw_buffer_2.x7.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X2731 VSS a_n3927_7727# hgu_cdac_half_1.db<5> VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2732 a_14132_1179# a_14017_1453# a_13709_1347# VSS sky130_fd_pr__nfet_01v8 ad=0.116 pd=1.09 as=0.0486 ps=0.63 w=0.36 l=0.15
X2733 a_n6959_14313# hgu_comp_flat_0.ready a_n7047_14175# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X2734 VDD a_n424_3698# hgu_sarlogic_flat_0.x4.x2.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2735 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<0> hgu_cdac_half_0.d<0> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.35
X2736 a_11756_1868# a_11244_1842# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.116 pd=1.09 as=0.166 ps=1.8 w=0.64 l=0.15
X2737 VDD VDD a_12359_7798# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X2738 hgu_cdac_sw_buffer_0.x12.X a_n412_n464# hgu_cdac_sw_buffer_0.VDD hgu_cdac_sw_buffer_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X2739 a_4449_1453# hgu_sarlogic_flat_0.x4.x11.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2740 VDD a_13636_1842# a_13546_2234# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X2741 hgu_sarlogic_flat_0.x4.x11.S a_10871_8513# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X2742 vin hgu_tah_0.sw_n hgu_tah_0.tah_vn hgu_tah_0.VDD sky130_fd_pr__pfet_01v8 ad=0.908 pd=5.83 as=1.71 ps=11.6 w=5.5 l=0.15
X2743 a_7509_6078# a_7369_6352# a_7071_6052# VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.0711 ps=0.755 w=0.36 l=0.15
X2744 VDD a_12358_6052# a_12291_6444# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X2745 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.db<6> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2746 a_12871_7824# a_12359_7798# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.084 ps=0.82 w=0.42 l=0.15
X2747 a_16427_4670# a_16581_4644# a_16287_4644# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2748 hgu_cdac_half_0.VREF hgu_cdac_half_0.d<5> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2749 VSS a_13067_1331# hgu_cdac_half_1.db<0> VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X2750 hgu_cdac_half_1.VREF hgu_cdac_half_1.d<4> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<15:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2751 hgu_cdac_half_1.d<6> a_n2219_8368# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2752 a_6723_6951# hgu_sarlogic_flat_0.x3.x7.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X2753 hgu_tah_0.VDD a_n54850_7835# hgu_vgen_vref_0.sky130_fd_sc_hd__dlymetal6s6s_1_3.A hgu_tah_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X2754 a_9463_6052# a_9761_6352# a_9697_6444# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0924 ps=0.86 w=0.42 l=0.15
X2755 hgu_cdac_half_1.d<6> a_n2219_8368# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2756 VDD async_delay_offset hgu_sarlogic_flat_0.x1.x4.x6.SW VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2757 a_16113_12401# hgu_sarlogic_flat_0.x2.x2.x2.IN a_16041_12539# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X2758 VDD a_n424_3698# hgu_sarlogic_flat_0.x4.x2.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2759 VSS a_n54567_7371# a_n54754_7113# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X2760 a_190_n245# hgu_cdac_sw_buffer_0.x6.A VSS VSS sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2761 VSS a_11625_1453# a_11626_1153# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2762 hgu_tah_0.tah_vn hgu_tah_0.sw_n hgu_tah_0.tah_vn VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.454 ps=3.08 w=2.75 l=0.15
X2763 hgu_sarlogic_flat_0.x1.x2.x10.Y async_setb_delay_cap_ctrl_code[3] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2764 VSS a_12556_8487# a_12491_8513# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X2765 VSS hgu_cdac_half_0.db<6> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2766 VDD VSS a_n3651_7087# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X2767 hgu_cdac_sw_buffer_1.x11.A a_1114_n1100# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2768 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2769 a_10638_13822# hgu_sarlogic_flat_0.x2.x2.x1.IN a_10550_13822# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X2770 a_9208_7317# a_8761_6951# a_9115_6951# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X2771 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2772 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.d<6> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2773 a_n1149_11335# hgu_sarlogic_flat_0.x1.x10.A VSS VDD sky130_fd_pr__pfet_01v8_hvt ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2774 VDD a_n3387_7727# hgu_cdac_half_1.db<4> VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2775 a_17184_4670# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X2776 VSS hgu_cdac_half_1.d<4> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<15:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2777 VSS hgu_cdac_half_1.d<5> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2778 VDD a_407_11578# a_406_11482# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2779 a_7888_8513# a_7285_8487# a_7772_8487# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2780 hgu_cdac_half_0.VREF hgu_cdac_half_0.d<6> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2781 VSS hgu_sarlogic_flat_0.x4.D[4] a_7759_1179# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2782 a_7570_2883# VSS a_7570_2556# VSS sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X2783 VSS a_9382_6925# a_9316_6951# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X2784 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_0.db<5> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2785 a_17184_5676# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X2786 a_17184_4670# a_16581_4644# a_17068_4644# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2787 a_3960_3698# hgu_sarlogic_flat_0.x4.x30.A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2788 hgu_sarlogic_flat_0.x4.x2.X a_n424_3698# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2789 hgu_cdac_half_0.VREF hgu_cdac_half_0.d<4> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<15:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.35
X2790 VDD VDD a_18973_5924# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X2791 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.db<6> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2792 hgu_vgen_vref_0.mimtop2 VSS sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X2793 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.d<6> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2794 VSS VDD a_11538_1842# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X2795 a_n1149_14360# hgu_sarlogic_flat_0.x1.x2.x9.output_stack hgu_sarlogic_flat_0.x1.x9.A VSS sky130_fd_pr__nfet_01v8 ad=0.0651 pd=0.73 as=0.122 ps=1.42 w=0.42 l=0.15
X2796 hgu_cdac_sw_buffer_1.VDD a_1666_n1100# hgu_cdac_half_0.d<5> hgu_cdac_sw_buffer_1.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2797 a_7153_2234# a_5840_1868# a_7069_2234# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0787 pd=0.795 as=0.0567 ps=0.69 w=0.42 l=0.15
X2798 VSS a_n716_1842# a_n782_1868# VSS sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0671 ps=0.75 w=0.42 l=0.15
X2799 hgu_cdac_half_1.db<5> a_n3927_7727# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2800 a_6533_1347# a_6842_1153# a_6777_1179# VSS sky130_fd_pr__nfet_01v8 ad=0.0486 pd=0.63 as=0.066 ps=0.745 w=0.36 l=0.15
X2801 hgu_sarlogic_flat_0.x2.x2.x2.x6.floating hgu_sarlogic_flat_0.x2.x2.x2.x6.SW hgu_sarlogic_flat_0.x2.x2.x2.x9.output_stack VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X2802 hgu_sarlogic_flat_0.x3.x4.X a_2036_7824# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2803 VSS a_2808_n935# hgu_cdac_sw_buffer_1.x7.X VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X2804 hgu_cdac_half_0.VREF hgu_cdac_half_0.db<6> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2805 hgu_sarlogic_flat_0.x2.x2.x4.x5[7].floating hgu_sarlogic_flat_0.x2.x2.x4.x10.Y hgu_sarlogic_flat_0.x2.x2.x4.x9.output_stack VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X2806 a_5396_6360# a_4437_6078# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X2807 a_16020_4670# hgu_sarlogic_flat_0.x4.D[6] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X2808 hgu_cdac_half_0.db<5> a_n688_n1104# hgu_cdac_sw_buffer_0.VDD hgu_cdac_sw_buffer_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2809 hgu_sarlogic_flat_0.x3.x4.X a_2036_7824# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2810 a_9222_7824# hgu_sarlogic_flat_0.x3.x4.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.154 ps=1.34 w=0.64 l=0.15
X2811 a_615_2556# hgu_sarlogic_flat_0.x4.x9.A1 a_394_2883# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X2812 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_1.db<5> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2813 a_6935_6078# a_7071_6052# a_6516_6052# VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0864 ps=0.91 w=0.64 l=0.15
X2814 VDD a_9762_6052# a_9761_6352# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2815 VSS a_3960_3698# hgu_sarlogic_flat_0.x4.x9.A1 VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2816 a_10151_1179# a_9234_1153# a_9706_1363# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0675 ps=0.735 w=0.36 l=0.15
X2817 hgu_vgen_vref_0.phi1_n a_n54752_8227# hgu_tah_0.VDD hgu_tah_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2818 hgu_sarlogic_flat_0.x4.x30.A a_3326_3698# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2819 hgu_vgen_vref_0.mimtop2 VSS sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X2820 a_19460_6564# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X2821 hgu_cdac_sw_buffer_3.x11.X a_n4397_8367# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2822 VSS a_n4397_8367# hgu_cdac_sw_buffer_3.x11.X VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2823 VSS a_1196_n1740# hgu_cdac_half_0.d<6> VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2824 a_n876_1179# hgu_sarlogic_flat_0.x4.x2.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2825 a_14544_1868# hgu_sarlogic_flat_0.x4.x2.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.03 as=0.0703 ps=0.755 w=0.42 l=0.15
X2826 a_15832_6596# a_15666_6596# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2827 hgu_vgen_vref_0.mimtop2 VSS sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X2828 hgu_cdac_half_1.VREF hgu_cdac_half_1.d<2> hgu_cdac_half_1.hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2829 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2830 VSS a_1716_n241# hgu_cdac_sw_buffer_1.x3.X VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X2831 a_5367_1179# a_4449_1453# a_4922_1363# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.0567 ps=0.69 w=0.42 l=0.15
X2832 VDD a_20768_8628# hgu_sarlogic_flat_0.x5.x3.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X2833 VSS hgu_cdac_half_1.d<6> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2834 a_11740_1179# a_11625_1453# a_11317_1347# VSS sky130_fd_pr__nfet_01v8 ad=0.116 pd=1.09 as=0.0486 ps=0.63 w=0.36 l=0.15
X2835 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2836 a_3499_1331# a_3595_1153# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X2837 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X2838 VSS hgu_cdac_half_1.db<6> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2839 a_n7660_7467# hgu_tah_0.tah_vp hgu_comp_flat_0.P VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X2840 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2841 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.db<6> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2842 VDD VDD a_6754_1842# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.17 ps=1.81 w=0.64 l=0.15
X2843 VSS a_7371_7798# a_7370_8098# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2844 a_8927_6951# a_8761_6951# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2845 a_9966_6052# a_10234_6262# a_10180_6360# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X2846 hgu_tah_0.VDD VSS sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X2847 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.d<6> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2848 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<15:0> hgu_cdac_half_1.db<4> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2849 a_7842_6262# a_7369_6352# a_8086_6078# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0671 ps=0.75 w=0.36 l=0.15
X2850 VSS a_12154_6052# a_12153_6352# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2851 a_7597_6951# a_6535_6951# a_7502_6951# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X2852 a_14734_1179# a_14222_1153# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0882 ps=0.84 w=0.42 l=0.15
X2853 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.db<6> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2854 VDD a_7284_6925# a_8005_7233# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X2855 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<0> hgu_cdac_half_0.d<0> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.244 ps=2.26 w=0.84 l=0.35
X2856 VSS a_10675_1331# hgu_cdac_half_1.db<1> VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X2857 hgu_cdac_half_0.db<6> a_n1158_n1744# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2858 hgu_vgen_vref_0.mimtop2 VSS sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X2859 VDD VDD a_n1189_1153# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0956 pd=0.875 as=0.132 ps=1.22 w=0.42 l=0.15
X2860 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_1.db<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.122 ps=1.42 w=0.42 l=0.35
X2861 hgu_cdac_sw_buffer_2.x5.A a_10341_1868# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X2862 a_4068_1842# a_3894_2234# a_4212_1868# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.0974 ps=0.97 w=0.64 l=0.15
X2863 VSS hgu_cdac_half_0.db<5> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2864 VDD hgu_sarlogic_flat_0.x2.x3.A a_3866_16177# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X2865 VSS a_2544_n241# hgu_cdac_half_0.d<3> VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X2866 a_1196_n1740# hgu_cdac_sw_buffer_1.x11.A VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2867 a_8644_2556# VSS a_8281_2708# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X2868 VDD a_7285_8487# a_8006_8795# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X2869 a_n6959_12689# hgu_comp_flat_0.clk a_n7047_12689# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X2870 a_382_1545# a_n130_1153# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X2871 hgu_cdac_half_0.VREF hgu_cdac_half_0.db<6> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2872 VDD a_11538_1842# a_12269_2150# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X2873 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<7:0> hgu_cdac_half_1.db<3> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2874 VSS a_n1158_n1744# hgu_cdac_half_0.db<6> VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2875 VSS hgu_cdac_half_0.db<6> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2876 a_12155_7798# hgu_sarlogic_flat_0.x3.x5.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2877 hgu_cdac_sw_buffer_0.VDD a_n1190_n245# hgu_cdac_sw_buffer_0.x9.X hgu_cdac_sw_buffer_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X2878 hgu_sarlogic_flat_0.x4.x20.X a_14746_2883# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.113 ps=1.04 w=0.65 l=0.15
X2879 hgu_cdac_half_0.d<6> a_1196_n1740# hgu_cdac_sw_buffer_1.VDD hgu_cdac_sw_buffer_1.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2880 a_4449_1453# hgu_sarlogic_flat_0.x4.x11.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2881 a_9421_6360# a_9221_6078# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X2882 hgu_cdac_half_1.VREF hgu_cdac_half_1.db<3> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<7:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2883 VDD a_2914_9360# hgu_sarlogic_flat_0.x5.eob VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.135 ps=1.27 w=1 l=0.15
X2884 VSS a_7574_6052# a_7509_6078# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0935 ps=0.965 w=0.64 l=0.15
X2885 hgu_sarlogic_flat_0.x2.x2.x3.x9.output_stack hgu_sarlogic_flat_0.x2.x2.x3.x10.Y hgu_sarlogic_flat_0.x2.x2.x3.x5[7].floating VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X2886 hgu_tah_0.tah_vp hgu_tah_0.sw vip VSS sky130_fd_pr__nfet_01v8 ad=0.454 pd=3.08 as=0.454 ps=3.08 w=2.75 l=0.15
X2887 VSS hgu_cdac_sw_buffer_1.x11.A a_1196_n1740# VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2888 hgu_vgen_vref_0.mimtop1 hgu_vgen_vref_0.mimbot1 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X2889 a_13207_2883# hgu_sarlogic_flat_0.x4.x20.S VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X2890 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<0> hgu_cdac_half_1.db<0> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.35
X2891 a_n55204_7371# hgu_vgen_vref_0.sky130_fd_sc_hd__dlymetal6s6s_1_5.A VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2892 VSS hgu_cdac_sw_buffer_3.x9.X a_n4479_7727# VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2893 VSS hgu_cdac_half_0.d<6> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2894 a_13067_1331# a_13163_1153# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2895 VDD a_1863_9386# hgu_sarlogic_flat_0.x3.x5.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2896 hgu_cdac_half_0.db<6> a_n1158_n1744# hgu_cdac_sw_buffer_0.VDD hgu_cdac_sw_buffer_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2897 hgu_sarlogic_flat_0.x2.x2.x2.x4[3].floating sample_delay_cap_ctrl_code[10] hgu_sarlogic_flat_0.x2.x2.x2.x9.output_stack VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X2898 a_9698_8190# a_8909_7798# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0819 ps=0.81 w=0.42 l=0.15
X2899 hgu_vgen_vref_0.mimtop1 hgu_vgen_vref_0.mimbot1 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X2900 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X2901 VSS a_7228_2136# a_7949_1868# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X2902 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2903 VSS a_n2219_8368# hgu_cdac_half_1.d<6> VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2904 VSS hgu_cdac_half_1.d<6> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2905 a_n6934_10472# hgu_comp_flat_0.clk a_n7022_10610# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X2906 a_10234_6262# a_9762_6052# a_10478_6444# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X2907 VDD a_7371_7798# a_7370_8098# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2908 VSS a_6990_6925# a_6924_6951# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X2909 a_13207_2556# hgu_sarlogic_flat_0.x4.x20.S VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X2910 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.d<6> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2911 VDD a_9146_1842# a_9096_2150# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X2912 VSS hgu_cdac_half_1.d<6> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2913 a_9383_8487# a_9209_8879# a_9523_8513# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X2914 VSS hgu_sarlogic_flat_0.x3.x5.X a_1586_8513# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2915 a_n53647_7835# a_n53551_7657# hgu_tah_0.VDD hgu_tah_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.141 ps=1.33 w=0.42 l=0.15
X2916 VSS hgu_cdac_half_1.db<6> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2917 VSS a_12555_6925# a_13262_6951# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X2918 a_18679_4644# a_18505_5036# a_18819_4670# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X2919 hgu_cdac_half_0.VREF hgu_cdac_half_0.db<6> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2920 hgu_sarlogic_flat_0.x4.x31.Q_N a_12012_2136# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X2921 a_4761_2234# a_3448_1868# a_4677_2234# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0787 pd=0.795 as=0.0567 ps=0.69 w=0.42 l=0.15
X2922 a_8813_6052# a_8908_6052# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2923 a_9568_1868# a_8398_1868# a_9461_2234# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0486 ps=0.63 w=0.36 l=0.15
X2924 a_n4397_8367# hgu_cdac_sw_buffer_3.x11.A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2925 VSS a_n4397_8367# hgu_cdac_sw_buffer_3.x11.X VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2926 hgu_cdac_half_1.VREF hgu_cdac_half_1.d<4> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<15:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2927 hgu_cdac_half_1.VREF hgu_cdac_half_1.d<5> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2928 a_3004_6360# a_2045_6078# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X2929 hgu_sarlogic_flat_0.x2.x2.x3.x3[1].floating sample_delay_cap_ctrl_code[13] hgu_sarlogic_flat_0.x2.x2.x3.x9.output_stack VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X2930 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X2931 a_9317_8513# a_8928_8513# a_9209_8879# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X2932 VSS a_n2219_8368# hgu_cdac_half_1.d<6> VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2933 hgu_cdac_half_1.VREF hgu_cdac_half_1.d<5> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2934 a_16221_5688# a_15832_5316# a_16113_5310# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X2935 a_8379_1153# a_8692_1179# a_8798_1179# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2936 hgu_vgen_vref_0.mimtop1 hgu_vgen_vref_0.phi1 hgu_vgen_vref_0.vcm VSS sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=0.5
X2937 a_4029_6052# a_4124_6052# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X2938 a_4836_2136# a_4677_2234# a_4976_1868# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.109 ps=1.03 w=0.64 l=0.15
X2939 a_1410_1868# hgu_sarlogic_flat_0.x4.D[6] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X2940 hgu_sarlogic_flat_0.x2.x3.A a_3080_14774# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X2941 VSS hgu_cdac_half_1.d<3> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<7:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2942 a_19286_6968# a_18058_6596# a_19144_6590# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X2943 a_18412_4670# hgu_sarlogic_flat_0.x4.x5.D VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X2944 a_8586_1868# hgu_sarlogic_flat_0.x4.D[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X2945 a_12155_7798# hgu_sarlogic_flat_0.x3.x5.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2946 a_7683_7317# a_6535_6951# a_7597_6951# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X2947 a_190_n245# hgu_cdac_sw_buffer_0.x6.A hgu_cdac_sw_buffer_0.VDD hgu_cdac_sw_buffer_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X2948 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_0.db<5> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2949 VSS a_6422_7798# hgu_sarlogic_flat_0.x4.x20.S VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X2950 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2951 VSS VSS a_n964_n464# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X2952 VSS sample_delay_offset hgu_sarlogic_flat_0.x2.x2.x1.x6.SW VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2953 VSS a_192_10793# hgu_comp_flat_0.clk VSS sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X2954 a_4196_9386# hgu_sarlogic_flat_0.x3.x48.Q VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0819 ps=0.81 w=0.42 l=0.15
X2955 a_18412_5310# hgu_sarlogic_flat_0.x4.D[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X2956 VSS a_11205_6052# hgu_sarlogic_flat_0.x4.D[3] VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X2957 VDD a_18973_5510# a_19694_5310# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X2958 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2959 VDD VDD a_2501_8487# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X2960 a_10163_6925# a_9989_6951# a_10279_6951# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X2961 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2962 VSS a_n1158_n1744# hgu_cdac_half_0.db<6> VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2963 VDD VDD a_4654_1153# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X2964 VSS a_3497_2708# hgu_sarlogic_flat_0.x4.x10.X VSS sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X2965 a_7046_1153# a_7314_1363# a_7260_1461# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X2966 VSS a_5987_1153# hgu_sarlogic_flat_0.x4.x26.Q_N VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X2967 a_7684_8879# a_6536_8513# a_7598_8513# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X2968 a_14654_8077# hgu_sarlogic_flat_0.x5.eob a_14566_8077# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X2969 a_334_10968# hgu_sarlogic_flat_0.x5.eob VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X2970 VDD a_16581_4644# a_17302_4952# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X2971 a_10673_2708# VSS a_10815_2883# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X2972 VDD a_8283_1331# hgu_cdac_sw_buffer_3.x5.A VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X2973 a_11613_6078# hgu_sarlogic_flat_0.x3.x4.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.154 ps=1.34 w=0.64 l=0.15
X2974 a_2188_1868# a_1676_1842# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.116 pd=1.09 as=0.166 ps=1.8 w=0.64 l=0.15
X2975 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.d<6> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2976 VSS hgu_vgen_vref_0.phi1_n hgu_vgen_vref_0.mimbot1 hgu_tah_0.VDD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=0.5
X2977 a_5450_6262# a_4977_6352# a_5694_6078# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0671 ps=0.75 w=0.36 l=0.15
X2978 VSS a_9762_6052# a_9761_6352# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2979 VDD a_9620_2136# a_10341_1868# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X2980 VSS hgu_cdac_sw_buffer_0.x11.A a_n1158_n1744# VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2981 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<15:0> hgu_cdac_half_0.db<4> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2982 VSS hgu_cdac_half_1.d<5> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2983 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.db<6> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2984 hgu_cdac_sw_buffer_3.x11.A a_n4479_7727# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2985 VDD a_4892_6925# a_5613_7233# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X2986 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_0.d<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X2987 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.d<6> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2988 VDD a_4068_1842# a_3978_2234# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X2989 a_n1158_n1744# hgu_cdac_sw_buffer_0.x11.A hgu_cdac_sw_buffer_0.VDD hgu_cdac_sw_buffer_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2990 a_n424_3698# hgu_sarlogic_flat_0.x4.x3.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2991 hgu_cdac_half_1.VREF hgu_cdac_half_1.d<6> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2992 a_n197_1545# a_n334_1153# a_n643_1347# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X2993 a_2036_7824# hgu_sarlogic_flat_0.x3.x4.A VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2994 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<0> hgu_cdac_half_0.db<0> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.35
X2995 a_1676_1842# a_1502_2234# a_1820_1868# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.0974 ps=0.97 w=0.64 l=0.15
X2996 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<15:0> hgu_cdac_half_1.db<4> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X2997 hgu_vgen_vref_0.phi1 a_n55304_8227# hgu_tah_0.VDD hgu_tah_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2998 a_n1699_7253# hgu_cdac_sw_buffer_2.x3.A VSS VSS sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2999 a_4331_6951# VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X3000 hgu_sarlogic_flat_0.x4.x9.A1 a_3960_3698# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3001 VSS hgu_sarlogic_flat_0.x4.x30.A a_3960_3698# VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3002 hgu_cdac_sw_buffer_0.VDD a_n148_n1104# hgu_cdac_half_0.db<4> hgu_cdac_sw_buffer_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3003 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_1.d<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3004 hgu_cdac_half_1.VREF hgu_cdac_half_1.db<6> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3005 VDD a_4893_8487# a_5614_8795# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X3006 a_5318_6078# a_5450_6262# a_5182_6052# VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0864 ps=0.91 w=0.64 l=0.15
X3007 hgu_cdac_half_0.VREF hgu_cdac_half_0.db<6> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3008 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X3009 a_n6887_12275# hgu_comp_flat_0.clk a_n6959_12413# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X3010 hgu_vgen_vref_0.mimtop2 VSS sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X3011 a_1325_11738# a_406_11482# a_879_11334# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X3012 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X3013 a_n871_7253# hgu_cdac_sw_buffer_2.x6.A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3014 a_8908_6052# a_9221_6078# a_9327_6078# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3015 hgu_sarlogic_flat_0.x5.x2.x9.output_stack retimer_delay_code[2] hgu_sarlogic_flat_0.x5.x2.x4[3].floating VSS sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X3016 hgu_tah_0.VDD a_n55770_7371# hgu_vgen_vref_0.sky130_fd_sc_hd__inv_1_1.A hgu_tah_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X3017 a_16287_5924# a_16113_6316# a_16427_5950# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X3018 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.db<6> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3019 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X3020 a_4332_8513# hgu_sarlogic_flat_0.x3.x27.D VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X3021 VSS hgu_cdac_sw_buffer_2.x11.A a_n2219_8368# VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3022 VSS hgu_cdac_half_0.d<6> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3023 a_14679_9742# hgu_sarlogic_flat_0.x5.eob a_14591_9604# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X3024 hgu_sarlogic_flat_0.x4.x3.A a_n1334_3698# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3025 VDD VDD a_1325_11738# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0662 ps=0.735 w=0.42 l=0.15
X3026 a_14358_1179# a_14490_1363# a_14222_1153# VSS sky130_fd_pr__nfet_01v8 ad=0.0974 pd=0.97 as=0.0864 ps=0.91 w=0.64 l=0.15
X3027 a_10815_2883# hgu_sarlogic_flat_0.x4.x17.S VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X3028 a_7503_8513# a_6991_8487# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X3029 a_1164_n241# hgu_cdac_sw_buffer_1.x9.A VSS VSS sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3030 a_10675_1331# a_10771_1153# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3031 hgu_sarlogic_flat_0.x1.x4.x10.Y async_resetb_delay_cap_ctrl_code[3] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3032 a_192_10793# hgu_sarlogic_flat_0.x1.x3.X a_334_10968# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X3033 hgu_sarlogic_flat_0.x1.x2.x9.output_stack async_setb_delay_cap_ctrl_code[2] hgu_sarlogic_flat_0.x1.x2.x4[3].floating VSS sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X3034 VSS hgu_sarlogic_flat_0.x4.x20.S a_4402_9386# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.066 ps=0.745 w=0.42 l=0.15
X3035 VDD a_12555_6925# a_13262_6951# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X3036 VSS hgu_cdac_half_0.d<3> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<7:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3037 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<7:0> hgu_cdac_half_1.db<3> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.35
X3038 a_16799_4670# a_16287_4644# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X3039 a_7314_1363# a_6842_1153# a_7558_1545# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X3040 VSS hgu_cdac_half_0.d<1> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<1:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.35
X3041 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_0.db<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.122 ps=1.42 w=0.42 l=0.35
X3042 hgu_cdac_sw_buffer_2.x6.A a_7949_1868# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X3043 VSS hgu_cdac_half_1.d<6> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3044 VDD hgu_sarlogic_flat_0.x3.x36.Q_N a_11300_6052# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.123 ps=1.17 w=0.42 l=0.15
X3045 hgu_vgen_vref_0.mimtop2 VSS sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X3046 a_3313_9386# hgu_sarlogic_flat_0.x4.x15.S VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.107 ps=1 w=0.42 l=0.15
X3047 VSS a_n54752_6595# hgu_vgen_vref_0.phi2_n VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3048 a_5115_6444# a_4978_6052# a_4679_6052# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X3049 hgu_cdac_half_0.VREF hgu_cdac_half_0.d<6> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3050 a_10815_2556# hgu_sarlogic_flat_0.x4.x17.S VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X3051 VSS hgu_cdac_half_1.d<6> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3052 VSS hgu_cdac_sw_buffer_3.x11.A a_n4397_8367# VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3053 a_9328_7824# a_9464_7798# a_8909_7798# VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0864 ps=0.91 w=0.64 l=0.15
X3054 hgu_sarlogic_flat_0.x2.x2.x1.x2.floating sample_delay_cap_ctrl_code[4] hgu_sarlogic_flat_0.x2.x2.x1.x9.output_stack VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.124 ps=1.43 w=0.42 l=0.15
X3055 VDD a_n2785_7946# hgu_cdac_sw_buffer_3.x7.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3056 VDD hgu_sarlogic_flat_0.x4.x5.D a_583_1179# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X3057 VSS hgu_cdac_half_1.db<5> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3058 VSS hgu_cdac_sw_buffer_2.x3.X a_n1749_7728# VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3059 result[4] a_17775_5326# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X3060 a_10663_16039# hgu_sarlogic_flat_0.x2.x2.x1.IN a_10575_15901# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X3061 VSS hgu_cdac_half_1.db<6> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3062 VSS a_10163_6925# a_10870_6951# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X3063 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_0.db<5> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3064 VDD hgu_sarlogic_flat_0.x3.x4.X a_12068_6925# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X3065 VSS a_466_n245# hgu_cdac_half_0.db<2> VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X3066 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3067 a_12012_2136# hgu_sarlogic_flat_0.x4.x2.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.132 pd=1.22 as=0.0956 ps=0.875 w=0.42 l=0.15
X3068 a_4001_14512# hgu_sarlogic_flat_0.x2.x3.A a_3929_14650# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X3069 a_n6959_13899# hgu_comp_flat_0.ready a_n7047_13899# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X3070 a_6925_8513# a_6536_8513# a_6817_8879# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X3071 a_3000_2883# VSS a_2786_2883# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.193 ps=1.34 w=0.42 l=0.15
X3072 hgu_cdac_sw_buffer_1.x12.X a_1942_n460# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3073 hgu_sarlogic_flat_0.x2.x2.x1.x4[3].floating sample_delay_cap_ctrl_code[6] hgu_sarlogic_flat_0.x2.x2.x1.x9.output_stack VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X3074 a_2033_8879# a_1586_8513# a_1940_8513# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X3075 VDD a_9676_6925# a_9626_7233# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X3076 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X3077 hgu_cdac_half_1.VREF hgu_cdac_half_1.d<6> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3078 hgu_vgen_vref_0.mimtop2 hgu_vgen_vref_0.phi2 hgu_vgen_vref_0.mimbot1 VSS sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=0.5
X3079 VSS a_n3927_7727# hgu_cdac_half_1.db<5> VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3080 a_12543_1179# a_11625_1453# a_12098_1363# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.0567 ps=0.69 w=0.42 l=0.15
X3081 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<7:0> hgu_cdac_half_0.db<3> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.35
X3082 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<15:0> hgu_cdac_half_1.d<4> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.35
X3083 a_19286_4670# a_18224_4670# a_19191_4670# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X3084 VDD a_n424_3698# hgu_sarlogic_flat_0.x4.x2.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3085 hgu_cdac_half_1.VREF hgu_cdac_half_1.db<6> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3086 a_n53647_7371# a_n53551_7113# hgu_tah_0.VDD hgu_tah_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.141 ps=1.33 w=0.42 l=0.15
X3087 a_7072_7798# a_7370_8098# a_7306_8190# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0924 ps=0.86 w=0.42 l=0.15
X3088 a_1637_6052# a_1732_6052# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X3089 a_2444_2136# a_2285_2234# a_2584_1868# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.109 ps=1.03 w=0.64 l=0.15
X3090 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_1.d<5> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3091 a_16894_6968# a_15666_6596# a_16752_6590# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X3092 a_16020_4670# hgu_sarlogic_flat_0.x4.D[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X3093 a_n1145_2883# hgu_sarlogic_flat_0.x4.x7.S VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X3094 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<15:0> hgu_cdac_half_1.d<4> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3095 VSS a_2207_8487# a_2141_8513# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X3096 hgu_vgen_vref_0.mimtop1 hgu_vgen_vref_0.mimbot1 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X3097 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<15:0> hgu_cdac_half_1.db<4> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3098 hgu_sarlogic_flat_0.x5.x2.x5[7].floating hgu_sarlogic_flat_0.x5.x2.x10.Y hgu_sarlogic_flat_0.x5.x2.x9.output_stack VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X3099 VSS hgu_sarlogic_flat_0.x4.x3.X a_n424_3698# VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3100 VSS hgu_sarlogic_flat_0.x3.x4.X a_7285_8487# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X3101 VDD a_9677_8487# a_9627_8795# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X3102 a_16020_5310# hgu_sarlogic_flat_0.x4.D[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X3103 VSS hgu_cdac_half_0.d<6> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3104 a_7069_2234# a_5840_1868# a_6972_1868# VSS sky130_fd_pr__nfet_01v8 ad=0.0486 pd=0.63 as=0.116 ps=1.09 w=0.36 l=0.15
X3105 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X3106 hgu_sarlogic_flat_0.x5.x1[1].Q_N a_19460_6564# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X3107 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_0.db<5> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3108 a_n1145_2556# hgu_sarlogic_flat_0.x4.x7.S VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X3109 a_1592_14732# hgu_sarlogic_flat_0.x2.x1.x3.Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X3110 hgu_cdac_half_1.d<6> a_n2219_8368# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3111 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.d<6> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3112 VSS a_3595_1153# hgu_sarlogic_flat_0.x4.x24.Q_N VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X3113 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3114 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X3115 hgu_vgen_vref_0.sky130_fd_sc_hd__nand2_1_0.Y hgu_vgen_vref_0.sky130_fd_sc_hd__inv_1_3.Y hgu_tah_0.VDD hgu_tah_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3116 a_4654_1153# a_4922_1363# a_4868_1461# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X3117 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3118 VSS a_9620_2136# a_9568_1868# VSS sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.066 ps=0.745 w=0.42 l=0.15
X3119 a_12573_2556# hgu_sarlogic_flat_0.x4.x9.A1 a_12352_2883# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X3120 VSS sel_bit[1] a_3783_9360# VSS sky130_fd_pr__nfet_01v8 ad=0.0819 pd=0.81 as=0.113 ps=1.38 w=0.42 l=0.15
X3121 VDD a_n424_3698# hgu_sarlogic_flat_0.x4.x2.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3122 VDD a_5891_1331# hgu_cdac_sw_buffer_3.x6.A VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X3123 a_2172_1179# a_2057_1453# a_1749_1347# VSS sky130_fd_pr__nfet_01v8 ad=0.116 pd=1.09 as=0.0486 ps=0.63 w=0.36 l=0.15
X3124 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<15:0> hgu_cdac_half_0.db<4> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3125 a_309_2150# a_n107_2234# a_52_2136# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.132 ps=1.22 w=0.84 l=0.15
X3126 hgu_sarlogic_flat_0.x1.x2.x5[7].floating hgu_sarlogic_flat_0.x1.x2.x10.Y hgu_sarlogic_flat_0.x1.x2.x9.output_stack VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X3127 VDD sel_bit[1] a_3783_9360# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3128 a_7772_8487# a_7598_8513# a_7888_8513# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X3129 a_12090_8190# a_11301_7798# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0819 ps=0.81 w=0.42 l=0.15
X3130 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.d<6> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3131 hgu_sarlogic_flat_0.x3.x4.X a_2036_7824# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3132 hgu_sarlogic_flat_0.x2.x2.x3.x9.output_stack hgu_sarlogic_flat_0.x2.x2.x3.x10.Y hgu_sarlogic_flat_0.x2.x2.x3.x5[7].floating VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X3133 VSS a_3960_3698# hgu_sarlogic_flat_0.x4.x9.A1 VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3134 VDD a_1676_1842# a_1586_2234# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X3135 a_n7660_7467# hgu_tah_0.tah_vp hgu_comp_flat_0.P VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.165 ps=1.33 w=1 l=0.15
X3136 a_12292_8190# a_12155_7798# a_11856_7798# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X3137 a_5166_1179# a_4654_1153# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0882 ps=0.84 w=0.42 l=0.15
X3138 VDD a_9233_1453# a_9234_1153# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3139 a_8678_2234# a_8398_1868# a_8586_1868# VSS sky130_fd_pr__nfet_01v8 ad=0.0675 pd=0.735 as=0.066 ps=0.745 w=0.36 l=0.15
X3140 hgu_cdac_half_1.VREF hgu_cdac_half_1.db<6> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3141 VSS a_n55770_7835# hgu_vgen_vref_0.sky130_fd_sc_hd__inv_1_0.A VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X3142 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_0.d<5> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3143 a_7498_2883# a_7316_2883# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X3144 VSS a_9967_7798# a_9902_7824# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0935 ps=0.965 w=0.64 l=0.15
X3145 a_n1287_2708# VSS a_n1145_2883# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X3146 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_1.d<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3147 VSS hgu_cdac_half_0.db<5> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3148 a_11205_6052# a_11300_6052# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3149 a_4638_8106# a_4438_7824# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X3150 VSS VSS a_n3651_7087# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X3151 a_3929_13960# hgu_sarlogic_flat_0.x2.x3.A a_3841_13822# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X3152 VSS hgu_cdac_half_1.db<5> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3153 a_12672_8513# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X3154 a_16041_12677# hgu_sarlogic_flat_0.x2.x2.x2.IN a_15953_12539# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X3155 a_6516_6052# a_6829_6078# a_6935_6078# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3156 a_6300_1179# hgu_sarlogic_flat_0.x4.x2.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3157 hgu_cdac_half_1.VREF hgu_cdac_half_1.d<5> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3158 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.d<6> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3159 VDD a_4598_6925# a_4508_7317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X3160 VDD a_5380_8487# a_5292_8879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X3161 vin hgu_tah_0.sw hgu_tah_0.tah_vn VSS sky130_fd_pr__nfet_01v8 ad=0.454 pd=3.08 as=0.454 ps=3.08 w=2.75 l=0.15
X3162 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.db<6> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3163 a_1940_8513# hgu_sarlogic_flat_0.x5.eob VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X3164 a_6318_2530# hgu_sarlogic_flat_0.x4.x13.S VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X3165 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_1.db<5> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3166 a_12672_8513# a_12069_8487# a_12556_8487# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3167 a_407_11578# hgu_tah_0.sw VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3168 VSS hgu_sarlogic_flat_0.x2.x3.A a_3929_13822# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X3169 a_2199_15136# a_971_14764# a_2057_14758# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X3170 a_12294_7824# a_12154_8098# a_11856_7798# VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.0711 ps=0.755 w=0.36 l=0.15
X3171 a_18224_5950# a_18058_5950# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3172 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<15:0> hgu_cdac_half_0.d<4> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3173 VDD a_4599_8487# a_4509_8879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X3174 VDD a_10163_6925# a_10870_6951# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X3175 a_2521_6444# a_1732_6052# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0819 ps=0.81 w=0.42 l=0.15
X3176 VSS a_17068_5924# a_17775_5950# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X3177 hgu_cdac_half_1.VREF hgu_cdac_half_1.db<5> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3178 VSS hgu_sarlogic_flat_0.x3.x75.Q a_6369_6951# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3179 VSS hgu_sarlogic_flat_0.x4.x3.X a_n424_3698# VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3180 hgu_cdac_sw_buffer_0.VDD VSS a_n964_n464# hgu_cdac_sw_buffer_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3181 hgu_cdac_half_0.VREF hgu_cdac_half_0.d<6> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3182 a_n643_1347# a_n334_1153# a_n399_1179# VSS sky130_fd_pr__nfet_01v8 ad=0.0486 pd=0.63 as=0.066 ps=0.745 w=0.36 l=0.15
X3183 a_6318_2530# hgu_sarlogic_flat_0.x4.x13.S VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X3184 a_11319_6951# a_11153_6951# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3185 a_11937_2234# a_10624_1868# a_11853_2234# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0787 pd=0.795 as=0.0567 ps=0.69 w=0.42 l=0.15
X3186 hgu_cdac_half_0.VREF hgu_cdac_half_0.db<4> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<15:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3187 VSS a_17068_6564# a_17775_6606# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X3188 a_2723_6444# a_2586_6052# a_2287_6052# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X3189 a_n54567_7371# a_n54471_7113# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3190 VDD a_18973_6790# a_18923_6590# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X3191 hgu_sarlogic_flat_0.x4.x30.A a_3326_3698# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3192 hgu_cdac_half_0.VREF hgu_cdac_half_0.d<3> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<7:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3193 a_19372_5036# a_18224_4670# a_19286_4670# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X3194 hgu_cdac_half_0.VREF hgu_cdac_half_0.d<1> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<1:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.35
X3195 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_0.db<5> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3196 VDD hgu_cdac_sw_buffer_2.x11.A a_n2219_8368# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3197 a_n7760_6349# a_n6526_6819# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.54 as=0.0759 ps=0.79 w=0.46 l=0.15
X3198 VDD a_n1699_7253# hgu_cdac_sw_buffer_2.x3.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3199 a_11719_6078# a_11855_6052# a_11300_6052# VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0864 ps=0.91 w=0.64 l=0.15
X3200 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_0.d<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3201 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3202 VDD hgu_sarlogic_flat_0.x3.x4.X a_9676_6925# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X3203 hgu_vgen_vref_0.mimtop1 hgu_vgen_vref_0.mimbot1 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X3204 hgu_cdac_half_0.VREF hgu_cdac_half_0.db<6> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3205 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<1:0> hgu_cdac_half_1.db<1> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.122 ps=1.42 w=0.42 l=0.35
X3206 a_n53647_7835# a_n53551_7657# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3207 VSS hgu_cdac_half_0.db<6> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3208 hgu_cdac_half_1.VREF hgu_cdac_half_1.d<6> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3209 a_n6887_13485# hgu_comp_flat_0.ready a_n6959_13623# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X3210 VSS a_n1147_7253# hgu_cdac_sw_buffer_2.x4.X VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X3211 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<7:0> hgu_cdac_half_0.db<3> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3212 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3213 hgu_sarlogic_flat_0.x1.x2.x9.output_stack async_delay_offset hgu_sarlogic_flat_0.x1.x2.x7.floating VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X3214 hgu_tah_0.VDD a_n55204_7835# a_n55391_7657# hgu_tah_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X3215 a_19286_6968# a_18224_6596# a_19191_6912# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X3216 hgu_cdac_half_1.VREF hgu_cdac_half_1.d<6> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3217 hgu_cdac_half_1.VREF hgu_cdac_half_1.db<6> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3218 VDD hgu_sarlogic_flat_0.x3.x4.X a_9677_8487# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X3219 VSS a_4124_6052# hgu_sarlogic_flat_0.x3.x54.Q_N VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X3220 a_16894_4670# a_15832_4670# a_16799_4670# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X3221 hgu_cdac_sw_buffer_1.VDD a_2808_n935# hgu_cdac_sw_buffer_1.x7.X hgu_cdac_sw_buffer_1.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3222 a_583_1179# a_n334_1153# a_138_1363# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0675 ps=0.735 w=0.36 l=0.15
X3223 VDD VDD a_11830_1153# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X3224 VDD a_1422_7824# hgu_sarlogic_flat_0.x3.x4.A VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3225 VDD a_6421_6052# hgu_sarlogic_flat_0.x4.D[5] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X3226 VDD a_1945_10648# hgu_tah_0.sw_n VDD sky130_fd_pr__pfet_01v8 ad=0.391 pd=3.14 as=0.208 ps=1.59 w=1.26 l=0.15
X3227 hgu_cdac_half_0.db<6> a_n1158_n1744# hgu_cdac_sw_buffer_0.VDD hgu_cdac_sw_buffer_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3228 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.db<6> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3229 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_0.db<5> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3230 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.d<6> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3231 VSS hgu_sarlogic_flat_0.x3.x4.X a_4893_8487# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X3232 VSS VDD a_6936_7824# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.12 ps=1.08 w=0.42 l=0.15
X3233 a_12626_6262# a_12153_6352# a_12870_6078# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0671 ps=0.75 w=0.36 l=0.15
X3234 a_4677_2234# a_3448_1868# a_4580_1868# VSS sky130_fd_pr__nfet_01v8 ad=0.0486 pd=0.63 as=0.116 ps=1.09 w=0.36 l=0.15
X3235 a_2584_1868# hgu_sarlogic_flat_0.x4.x2.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.03 as=0.0703 ps=0.755 w=0.42 l=0.15
X3236 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.db<6> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3237 a_12555_6925# hgu_sarlogic_flat_0.x3.x39.Q_N VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X3238 a_16041_11849# hgu_sarlogic_flat_0.x2.x2.x2.IN hgu_sarlogic_flat_0.x2.x2.x2.x9.output_stack VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X3239 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3240 a_5176_2883# hgu_sarlogic_flat_0.x4.x9.A1 a_5104_2883# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X3241 VSS a_n54850_7371# hgu_vgen_vref_0.sky130_fd_sc_hd__dlymetal6s6s_1_5.A VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X3242 VSS hgu_vgen_vref_0.sky130_fd_sc_hd__inv_1_3.A a_n55304_6595# VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3243 a_10479_7824# a_9967_7798# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.084 ps=0.82 w=0.42 l=0.15
X3244 a_5314_6951# a_3977_6951# a_5205_6951# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X3245 hgu_cdac_sw_buffer_0.VDD hgu_cdac_sw_buffer_0.x9.X a_n1240_n1104# hgu_cdac_sw_buffer_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3246 hgu_sarlogic_flat_0.x2.x2.x3.x6.SW sample_delay_offset VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3247 VDD a_n2301_7728# hgu_cdac_sw_buffer_2.x11.A VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3248 VSS hgu_cdac_half_0.db<5> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3249 VDD a_n7216_6420# hgu_comp_flat_0.comp_outp VDD sky130_fd_pr__pfet_01v8 ad=0.139 pd=1.17 as=0.26 ps=2.3 w=0.84 l=0.15
X3250 a_n1158_n1744# hgu_cdac_sw_buffer_0.x11.A VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3251 hgu_cdac_half_0.VREF hgu_cdac_half_0.d<6> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3252 a_9706_1363# a_9234_1153# a_9950_1545# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X3253 hgu_cdac_half_0.VREF hgu_cdac_half_0.db<6> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3254 VSS hgu_cdac_half_0.db<6> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.35
X3255 VSS hgu_sarlogic_flat_0.x2.x2.x3.IN a_10023_11461# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3256 hgu_cdac_sw_buffer_0.VDD hgu_cdac_sw_buffer_0.x11.A a_n1158_n1744# hgu_cdac_sw_buffer_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3257 a_9317_2150# a_8852_1842# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X3258 a_7711_7824# a_7843_8008# a_7575_7798# VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0864 ps=0.91 w=0.64 l=0.15
X3259 a_12556_8487# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X3260 a_5176_2556# a_4922_2883# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.145 ps=1.11 w=0.42 l=0.15
X3261 hgu_sarlogic_flat_0.x1.x2.x9.output_stack async_setb_delay_cap_ctrl_code[2] hgu_sarlogic_flat_0.x1.x2.x4[3].floating VSS sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X3262 a_4598_6925# a_4424_7317# a_4738_6951# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X3263 a_10710_14236# hgu_sarlogic_flat_0.x2.x2.x1.IN a_10638_14374# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X3264 a_2774_1179# a_2262_1153# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0882 ps=0.84 w=0.42 l=0.15
X3265 hgu_comp_flat_0.comp_outn a_n6292_6446# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0759 pd=0.79 as=0.143 ps=1.54 w=0.46 l=0.15
X3266 a_4014_1179# a_4141_1347# a_3595_1153# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.03 as=0.0864 ps=0.91 w=0.64 l=0.15
X3267 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<7:0> hgu_cdac_half_1.d<3> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3268 VSS hgu_cdac_half_0.db<5> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3269 a_3494_9752# a_3378_9360# a_3408_9386# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.16 as=0.0567 ps=0.69 w=0.42 l=0.15
X3270 a_n7760_6349# a_n7766_6446# a_n7678_6446# VDD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.15
X3271 hgu_sarlogic_flat_0.x3.x30.Q_N a_7772_8487# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X3272 VSS a_n4479_7727# hgu_cdac_sw_buffer_3.x11.A VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3273 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3274 a_n1149_11335# hgu_sarlogic_flat_0.x1.x4.x9.output_stack VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X3275 VDD a_1863_9386# hgu_sarlogic_flat_0.x3.x5.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3276 hgu_cdac_sw_buffer_0.VDD a_466_n245# hgu_cdac_half_0.db<2> hgu_cdac_sw_buffer_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3277 a_454_n939# VSS hgu_cdac_sw_buffer_0.VDD hgu_cdac_sw_buffer_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3278 VSS hgu_cdac_sw_buffer_0.x4.X a_n148_n1104# VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3279 VSS a_n1189_1153# hgu_cdac_sw_buffer_0.x9.A VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X3280 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.122 ps=1.42 w=0.42 l=0.35
X3281 hgu_vgen_vref_0.mimtop2 VSS sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X3282 a_12089_6444# a_11300_6052# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0819 ps=0.81 w=0.42 l=0.15
X3283 VDD a_17068_5924# a_17775_5950# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X3284 hgu_sarlogic_flat_0.x5.x1[6].Q_N a_17068_4644# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X3285 hgu_tah_0.VDD VSS sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X3286 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3287 hgu_sarlogic_flat_0.x1.x4.x9.output_stack hgu_sarlogic_flat_0.x1.x4.x10.Y hgu_sarlogic_flat_0.x1.x4.x5[7].floating VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X3288 a_4331_6951# VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X3289 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X3290 a_3614_1868# a_3448_1868# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3291 VDD a_5183_7798# a_5116_8190# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X3292 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.db<6> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3293 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_1.d<5> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3294 a_1105_2708# VSS a_1247_2883# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X3295 a_9332_12125# hgu_sarlogic_flat_0.x2.x2.x3.IN a_9244_11987# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X3296 vip hgu_tah_0.sw hgu_tah_0.tah_vp VSS sky130_fd_pr__nfet_01v8 ad=0.454 pd=3.08 as=0.853 ps=6.12 w=2.75 l=0.15
X3297 VSS hgu_sarlogic_flat_0.x4.x13.S a_13073_7824# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3298 VDD a_13930_1842# a_13880_2150# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X3299 hgu_sarlogic_flat_0.x4.x9.X a_2786_2883# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.113 ps=1.04 w=0.65 l=0.15
X3300 VSS hgu_cdac_half_0.d<6> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3301 hgu_sarlogic_flat_0.x2.x2.x1.x4[3].floating sample_delay_cap_ctrl_code[6] hgu_sarlogic_flat_0.x2.x2.x1.x9.output_stack VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X3302 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_1.d<5> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3303 hgu_vgen_vref_0.mimtop2 VSS sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X3304 a_11084_1179# hgu_sarlogic_flat_0.x4.x2.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.17 pd=1.81 as=0.154 ps=1.34 w=0.64 l=0.15
X3305 VSS a_n6994_7879# a_n7390_7871# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X3306 hgu_cdac_half_0.VREF hgu_cdac_half_0.db<4> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<15:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3307 VSS hgu_cdac_half_0.db<3> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<7:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3308 VSS a_9233_1453# a_9234_1153# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3309 VSS a_n4397_8367# hgu_cdac_sw_buffer_3.x11.X VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3310 hgu_sarlogic_flat_0.x2.x2.x1.x9.output_stack hgu_sarlogic_flat_0.x2.x2.x1.x10.Y hgu_sarlogic_flat_0.x2.x2.x1.x5[7].floating VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X3311 a_9962_2883# hgu_sarlogic_flat_0.x4.x9.A1 a_9890_2883# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X3312 a_9739_14835# hgu_sarlogic_flat_0.x2.x2.x4.x9.output_stack VSS VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X3313 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<15:0> hgu_cdac_half_0.d<4> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3314 VSS a_n2219_8368# hgu_cdac_half_1.d<6> VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3315 hgu_cdac_sw_buffer_2.x9.A a_773_1868# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X3316 hgu_cdac_half_1.VREF hgu_cdac_half_1.d<5> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3317 VDD hgu_sarlogic_flat_0.x3.x20.Q_N a_1732_6052# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.123 ps=1.17 w=0.42 l=0.15
X3318 VSS hgu_cdac_half_0.d<5> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3319 a_8928_8513# a_8762_8513# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3320 a_16980_5036# a_15832_4670# a_16894_4670# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X3321 hgu_sarlogic_flat_0.x2.x2.x2.x5[7].floating hgu_sarlogic_flat_0.x2.x2.x2.x10.Y hgu_sarlogic_flat_0.x2.x2.x2.x9.output_stack VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X3322 VSS hgu_vgen_vref_0.sky130_fd_sc_hd__inv_1_2.Y a_n54752_8227# VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3323 a_14726_7663# hgu_sarlogic_flat_0.x5.eob a_14654_7801# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X3324 VDD a_n3325_7252# hgu_cdac_sw_buffer_3.x4.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3325 a_9962_2556# a_9708_2883# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.145 ps=1.11 w=0.42 l=0.15
X3326 VSS hgu_cdac_half_0.db<6> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3327 VSS a_11244_1842# a_11178_1868# VSS sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0671 ps=0.75 w=0.42 l=0.15
X3328 VSS hgu_sarlogic_flat_0.x3.x36.Q_N a_12494_6078# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.101 ps=0.99 w=0.42 l=0.15
X3329 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_0.d<5> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3330 a_n386_1545# a_n1189_1153# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0787 pd=0.795 as=0.0956 ps=0.875 w=0.42 l=0.15
X3331 a_n1149_14360# hgu_sarlogic_flat_0.x1.x9.A VDD VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3332 hgu_sarlogic_flat_0.x3.x7.X a_1454_6950# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3333 a_19460_5284# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X3334 VDD a_4836_2136# a_5557_1868# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X3335 hgu_sarlogic_flat_0.x2.x2.x3.x9.output_stack hgu_sarlogic_flat_0.x2.x2.x3.x10.Y hgu_sarlogic_flat_0.x2.x2.x3.x5[7].floating VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X3336 a_16894_6968# a_15832_6596# a_16799_6912# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X3337 hgu_comp_flat_0.Q hgu_tah_0.tah_vn a_n7660_7467# VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.31 ps=2.62 w=1 l=0.15
X3338 result[2] a_17775_5950# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X3339 a_19460_5924# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X3340 a_14245_2234# a_13016_1868# a_14148_1868# VSS sky130_fd_pr__nfet_01v8 ad=0.0486 pd=0.63 as=0.116 ps=1.09 w=0.36 l=0.15
X3341 VSS a_1732_6052# hgu_sarlogic_flat_0.x3.x51.Q_N VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X3342 a_15832_5316# a_15666_5316# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3343 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3344 VSS a_10771_1153# hgu_sarlogic_flat_0.x4.x32.Q_N VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X3345 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.d<6> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3346 VSS hgu_cdac_half_1.db<5> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3347 VSS hgu_sarlogic_flat_0.x3.x5.A a_1863_9386# VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3348 hgu_tah_0.VDD VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X3349 a_3614_1868# a_3448_1868# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3350 VSS hgu_sarlogic_flat_0.x1.x9.Y a_747_11682# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.101 ps=0.99 w=0.42 l=0.15
X3351 VSS VDD a_11190_1179# VSS sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.109 ps=1.03 w=0.42 l=0.15
X3352 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.d<6> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3353 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.db<6> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3354 hgu_cdac_sw_buffer_3.x11.A a_n4479_7727# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3355 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3356 a_16448_15176# hgu_sarlogic_flat_0.x2.x2.x1.x9.output_stack VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X3357 hgu_cdac_half_1.VREF hgu_cdac_half_1.db<4> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<15:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3358 hgu_tah_0.tah_vp hgu_tah_0.sw hgu_tah_0.tah_vp hgu_tah_0.VDD sky130_fd_pr__pfet_01v8 ad=8.85 pd=58.2 as=0.908 ps=5.83 w=5.5 l=0.15
X3359 VDD VSS a_n4203_7087# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3360 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.db<6> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3361 a_9379_10322# hgu_sarlogic_flat_0.x2.x2.x3.IN a_9291_10460# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X3362 VSS hgu_cdac_half_0.db<5> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.35
X3363 a_12381_6951# a_11153_6951# a_12239_7233# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X3364 hgu_cdac_half_0.VREF hgu_cdac_half_0.db<6> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3365 a_2036_7824# hgu_sarlogic_flat_0.x3.x4.A VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3366 hgu_cdac_sw_buffer_1.VDD VSS a_1390_n460# hgu_cdac_sw_buffer_1.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3367 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<1:0> hgu_cdac_half_0.db<1> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.35
X3368 a_n6887_11999# hgu_comp_flat_0.clk a_n6959_11999# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X3369 VDD a_8909_7798# hgu_sarlogic_flat_0.x3.x42.Q_N VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X3370 VSS hgu_sarlogic_flat_0.x4.x30.A a_3960_3698# VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3371 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X3372 VDD a_16287_4644# a_16197_5036# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X3373 VDD a_12555_6925# a_12467_7317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X3374 a_6925_2150# a_6460_1842# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X3375 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.d<6> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3376 a_n447_11350# a_108_11334# a_66_11360# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0882 ps=1.05 w=0.84 l=0.15
X3377 a_12044_1461# a_11084_1179# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X3378 a_12382_8513# a_11154_8513# a_12240_8795# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X3379 VSS hgu_cdac_half_1.d<6> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.35
X3380 a_394_2883# VSS a_394_2556# VSS sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X3381 hgu_vgen_vref_0.mimtop1 hgu_vgen_vref_0.mimbot1 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X3382 a_13476_1179# hgu_sarlogic_flat_0.x4.x2.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3383 hgu_vgen_vref_0.mimtop1 hgu_vgen_vref_0.mimbot1 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X3384 a_192_1868# a_n422_1842# a_52_2136# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3385 VSS hgu_cdac_half_1.db<6> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3386 VDD a_12556_8487# a_12468_8879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X3387 hgu_cdac_half_1.hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT hgu_cdac_half_1.d<2> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.35
X3388 hgu_cdac_half_1.VREF hgu_cdac_half_1.db<3> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<7:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3389 hgu_tah_0.VDD a_n55304_6595# hgu_vgen_vref_0.phi2 hgu_tah_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3390 VSS hgu_sarlogic_flat_0.x5.x3.X a_18058_4670# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3391 a_1107_1331# a_1203_1153# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X3392 hgu_sarlogic_flat_0.x3.x27.Q_N a_5380_8487# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X3393 a_1448_10615# hgu_tah_0.sw VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X3394 VSS a_n4397_8367# hgu_cdac_sw_buffer_3.x11.X VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3395 a_6535_6951# a_6369_6951# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3396 a_9763_7798# hgu_sarlogic_flat_0.x3.x5.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3397 VSS hgu_sarlogic_flat_0.x5.x3.X a_18058_5316# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3398 a_3898_9386# a_3378_9360# a_4173_9684# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.164 ps=1.33 w=0.42 l=0.15
X3399 a_8087_8190# a_7575_7798# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X3400 a_n53930_7835# a_n53834_7657# hgu_tah_0.VDD hgu_tah_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.141 ps=1.33 w=0.42 l=0.15
X3401 a_9697_6078# a_8908_6052# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0588 ps=0.7 w=0.42 l=0.15
X3402 VSS a_407_11578# a_406_11482# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3403 hgu_sarlogic_flat_0.x3.x3.A a_1146_7824# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3404 a_5183_7798# a_4438_7824# a_5319_7824# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3405 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.db<6> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3406 a_6604_1868# hgu_sarlogic_flat_0.x4.x2.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0974 pd=0.97 as=0.0882 ps=0.84 w=0.42 l=0.15
X3407 a_n204_1868# a_n716_1842# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.116 pd=1.09 as=0.166 ps=1.8 w=0.64 l=0.15
X3408 a_3104_8513# hgu_sarlogic_flat_0.x3.x4.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X3409 VSS a_n54752_6595# hgu_vgen_vref_0.phi2_n VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3410 hgu_cdac_sw_buffer_1.VDD a_2268_n241# hgu_cdac_sw_buffer_1.x4.X hgu_cdac_sw_buffer_1.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3411 hgu_cdac_half_0.d<4> a_2206_n1100# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3412 a_8281_2708# hgu_sarlogic_flat_0.x4.x9.A1 a_8423_2556# VSS sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X3413 a_4424_7317# a_3977_6951# a_4331_6951# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X3414 a_9966_6052# a_9221_6078# a_10102_6078# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3415 VSS hgu_cdac_half_1.db<6> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3416 VSS hgu_sarlogic_flat_0.x4.x15.S a_10681_7824# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3417 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3418 a_3104_8513# a_2501_8487# a_2988_8487# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3419 hgu_sarlogic_flat_0.x2.x2.x3.x9.output_stack sample_delay_cap_ctrl_code[12] hgu_sarlogic_flat_0.x2.x2.x3.x2.floating VSS sky130_fd_pr__nfet_01v8 ad=0.124 pd=1.43 as=0.122 ps=1.42 w=0.42 l=0.15
X3420 VSS a_4598_6925# a_4532_6951# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X3421 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.d<6> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.35
X3422 a_6422_7798# a_6517_7798# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X3423 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3424 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.db<6> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3425 a_n55487_7835# a_n55391_7657# hgu_tah_0.VDD hgu_tah_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.141 ps=1.33 w=0.42 l=0.15
X3426 a_9404_12401# hgu_sarlogic_flat_0.x2.x2.x3.IN a_9332_12401# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X3427 hgu_cdac_half_1.d<4> a_n1209_7728# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3428 VSS a_2206_n1100# hgu_cdac_half_0.d<4> VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3429 hgu_cdac_half_0.VREF hgu_cdac_half_0.d<6> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3430 VSS a_n871_7253# hgu_cdac_half_1.d<3> VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X3431 hgu_cdac_half_1.VREF hgu_cdac_half_1.d<5> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3432 VDD hgu_sarlogic_flat_0.x3.x4.A a_2036_7824# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3433 VSS a_454_n939# hgu_cdac_sw_buffer_0.x7.X VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X3434 VSS VDD a_6_1179# VSS sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0974 ps=0.97 w=0.42 l=0.15
X3435 hgu_cdac_half_0.VREF hgu_cdac_half_0.db<5> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3436 a_2369_2234# a_1056_1868# a_2285_2234# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0787 pd=0.795 as=0.0567 ps=0.69 w=0.42 l=0.15
X3437 a_7791_2556# hgu_sarlogic_flat_0.x4.x9.A1 a_7570_2883# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X3438 VSS a_6517_7798# hgu_sarlogic_flat_0.x3.x45.Q_N VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X3439 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X3440 VSS hgu_cdac_half_1.d<3> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<7:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3441 a_15832_5950# a_15666_5950# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3442 hgu_sarlogic_flat_0.x4.x9.A1 a_3960_3698# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3443 VDD VDD a_n422_1842# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.17 ps=1.81 w=0.64 l=0.15
X3444 a_2151_6078# a_2287_6052# a_1732_6052# VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0864 ps=0.91 w=0.64 l=0.15
X3445 hgu_cdac_sw_buffer_0.VDD a_n1158_n1744# hgu_cdac_half_0.db<6> hgu_cdac_sw_buffer_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3446 hgu_cdac_half_0.VREF hgu_cdac_half_0.d<5> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3447 a_5987_1153# a_6300_1179# a_6406_1179# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3448 a_15832_6596# a_15666_6596# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3449 a_18589_6590# a_18058_6596# a_18505_6590# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X3450 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3451 a_n424_3698# hgu_sarlogic_flat_0.x4.x3.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3452 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X3453 a_9763_7798# hgu_sarlogic_flat_0.x3.x5.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3454 a_19286_5688# a_18058_5316# a_19144_5310# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X3455 hgu_cdac_sw_buffer_1.VDD hgu_cdac_sw_buffer_1.x11.A a_1196_n1740# hgu_cdac_sw_buffer_1.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3456 VSS a_14222_1153# a_14132_1179# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.116 ps=1.09 w=0.64 l=0.15
X3457 VDD a_8379_1153# hgu_sarlogic_flat_0.x4.x29.Q_N VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X3458 a_6991_8487# a_6817_8879# a_7131_8513# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X3459 a_11915_8513# a_12069_8487# a_11775_8487# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3460 VSS a_n638_n245# hgu_cdac_sw_buffer_0.x3.X VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X3461 a_11853_2234# a_10624_1868# a_11756_1868# VSS sky130_fd_pr__nfet_01v8 ad=0.0486 pd=0.63 as=0.116 ps=1.09 w=0.36 l=0.15
X3462 VDD EXT_CLK a_971_14764# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3463 a_n7660_7467# hgu_comp_flat_0.clk VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X3464 a_18819_6956# a_18973_6790# a_18679_6564# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3465 a_19286_5950# a_18058_5950# a_19144_6232# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X3466 hgu_cdac_half_0.db<6> a_n1158_n1744# hgu_cdac_sw_buffer_0.VDD hgu_cdac_sw_buffer_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3467 hgu_cdac_half_0.VREF hgu_cdac_half_0.db<3> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<7:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.35
X3468 hgu_sarlogic_flat_0.x4.x28.Q_N a_9620_2136# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X3469 VSS hgu_cdac_half_1.d<4> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<15:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3470 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.d<6> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3471 VSS a_1105_2708# hgu_sarlogic_flat_0.x4.x8.X VSS sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X3472 VDD hgu_comp_flat_0.clk a_1587_9386# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3473 a_4438_7824# hgu_sarlogic_flat_0.x3.x4.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.154 ps=1.34 w=0.64 l=0.15
X3474 a_16287_6564# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X3475 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.d<6> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3476 hgu_cdac_sw_buffer_1.VDD a_1114_n1100# hgu_cdac_sw_buffer_1.x11.A hgu_cdac_sw_buffer_1.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3477 hgu_vgen_vref_0.mimtop1 hgu_vgen_vref_0.mimbot1 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X3478 a_3058_6262# a_2585_6352# a_3302_6078# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0671 ps=0.75 w=0.36 l=0.15
X3479 a_19395_5688# a_18058_5316# a_19286_5688# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X3480 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<15:0> hgu_cdac_half_1.db<4> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3481 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.d<6> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3482 a_11190_1179# a_11317_1347# a_10771_1153# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.03 as=0.0864 ps=0.91 w=0.64 l=0.15
X3483 hgu_cdac_half_1.VREF hgu_cdac_half_1.db<6> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3484 hgu_cdac_half_0.VREF hgu_cdac_half_0.db<6> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3485 a_3954_15763# hgu_sarlogic_flat_0.x2.x3.A a_3866_15901# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X3486 hgu_vgen_vref_0.mimbot1 hgu_vgen_vref_0.phi1 VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=0.5
X3487 VSS hgu_cdac_sw_buffer_3.x11.A a_n4397_8367# VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3488 a_9379_10598# hgu_sarlogic_flat_0.x2.x2.x3.IN a_9291_10736# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X3489 a_2988_8487# hgu_sarlogic_flat_0.x3.x4.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X3490 a_15832_4670# a_15666_4670# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3491 a_11320_8513# a_11154_8513# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3492 a_17302_6590# a_16894_6968# a_17068_6564# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X3493 VSS VSS a_1942_n460# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X3494 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X3495 hgu_sarlogic_flat_0.x2.x2.x1.x9.output_stack hgu_sarlogic_flat_0.x2.x2.x1.x10.Y hgu_sarlogic_flat_0.x2.x2.x1.x5[7].floating VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X3496 a_4739_8513# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X3497 a_14654_8491# hgu_sarlogic_flat_0.x5.eob a_14566_8353# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X3498 VDD a_n335_1453# a_n334_1153# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3499 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X3500 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3501 hgu_cdac_half_1.VREF hgu_cdac_half_1.db<2> hgu_cdac_half_1.hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3502 hgu_sarlogic_flat_0.x1.x4.x9.output_stack async_resetb_delay_cap_ctrl_code[2] hgu_sarlogic_flat_0.x1.x4.x4[3].floating VSS sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X3503 VDD a_12359_7798# a_12292_8190# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X3504 a_19191_5632# a_18679_5284# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X3505 VSS sample_delay_cap_ctrl_code[15] hgu_sarlogic_flat_0.x2.x2.x3.x10.Y VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3506 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X3507 hgu_sarlogic_flat_0.x4.x15.X a_9962_2883# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.113 ps=1.04 w=0.65 l=0.15
X3508 a_3929_14236# hgu_sarlogic_flat_0.x2.x3.A a_3841_14098# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X3509 a_5695_8190# a_5183_7798# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X3510 VDD a_12012_2136# a_11937_2234# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0956 pd=0.875 as=0.0787 ps=0.795 w=0.42 l=0.15
X3511 a_19576_6956# a_18973_6790# a_19460_6564# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3512 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_0.db<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3513 a_6460_1842# hgu_sarlogic_flat_0.x4.x2.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X3514 a_7046_1153# a_6300_1179# a_7182_1179# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3515 VDD a_2036_7824# hgu_sarlogic_flat_0.x3.x4.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3516 hgu_comp_flat_0.RS_n hgu_comp_flat_0.RS_p VDD VDD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.15
X3517 VSS hgu_cdac_sw_buffer_3.x3.X a_n3927_7727# VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3518 hgu_sarlogic_flat_0.x3.x3.A a_1146_7824# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3519 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3520 a_6979_1545# a_6842_1153# a_6533_1347# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X3521 a_6491_1461# a_6300_1179# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X3522 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3523 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<15:0> hgu_cdac_half_0.d<4> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3524 VSS a_2444_2136# a_3165_1868# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X3525 VSS hgu_cdac_half_1.db<5> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3526 VSS hgu_cdac_half_0.d<6> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3527 VSS hgu_cdac_half_0.db<6> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3528 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.d<6> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3529 hgu_cdac_half_1.hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT hgu_cdac_half_1.db<2> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3530 hgu_cdac_half_0.db<4> a_n148_n1104# hgu_cdac_sw_buffer_0.VDD hgu_cdac_sw_buffer_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3531 VDD a_4362_1842# a_4312_2150# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X3532 VSS a_n7390_7871# a_n7766_6446# VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.54 as=0.0759 ps=0.79 w=0.46 l=0.15
X3533 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.d<6> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3534 VDD a_4030_7798# hgu_sarlogic_flat_0.x3.x48.Q VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X3535 a_9382_6925# hgu_sarlogic_flat_0.x3.x42.Q_N VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X3536 hgu_sarlogic_flat_0.x1.x2.x9.output_stack hgu_comp_flat_0.ready a_n7022_15150# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X3537 VSS hgu_vgen_vref_0.clk hgu_vgen_vref_0.sky130_fd_sc_hd__inv_1_4.Y VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3538 a_n53930_7371# a_n53834_7113# hgu_tah_0.VDD hgu_tah_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.141 ps=1.33 w=0.42 l=0.15
X3539 a_1196_n1740# hgu_cdac_sw_buffer_1.x11.A VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3540 hgu_vgen_vref_0.mimtop1 hgu_vgen_vref_0.mimbot1 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X3541 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.d<6> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3542 hgu_cdac_half_1.VREF hgu_cdac_half_1.d<6> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3543 a_8908_6052# a_9463_6052# a_9421_6360# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0882 ps=1.05 w=0.84 l=0.15
X3544 VSS hgu_sarlogic_flat_0.x4.x3.X a_n424_3698# VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3545 hgu_sarlogic_flat_0.x2.x1.x4.Y VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3546 VDD a_n424_3698# hgu_sarlogic_flat_0.x4.x2.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3547 hgu_cdac_half_1.VREF hgu_cdac_half_1.db<6> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3548 a_9463_6052# a_9762_6052# a_9697_6078# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.066 ps=0.745 w=0.36 l=0.15
X3549 a_11966_1179# a_12098_1363# a_11830_1153# VSS sky130_fd_pr__nfet_01v8 ad=0.0974 pd=0.97 as=0.0864 ps=0.91 w=0.64 l=0.15
X3550 hgu_sarlogic_flat_0.x3.x4.X a_2036_7824# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3551 a_9383_8487# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X3552 VDD a_1422_7824# hgu_sarlogic_flat_0.x3.x4.A VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3553 VSS hgu_cdac_half_1.d<2> hgu_cdac_half_1.hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3554 a_n53364_7371# hgu_vgen_vref_0.sky130_fd_sc_hd__nand2_1_1.Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3555 a_11301_7798# a_11614_7824# a_11720_7824# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3556 VDD a_7284_6925# a_7234_7233# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X3557 result[1] a_20167_6606# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X3558 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X3559 VDD hgu_sarlogic_flat_0.x4.x17.S a_8289_7824# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0662 ps=0.735 w=0.42 l=0.15
X3560 hgu_sarlogic_flat_0.x4.x2.X a_n424_3698# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3561 hgu_sarlogic_flat_0.x3.x77.Y hgu_sarlogic_flat_0.x5.eob VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3562 hgu_sarlogic_flat_0.x4.x2.X a_n424_3698# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3563 hgu_cdac_sw_buffer_3.x11.X a_n4397_8367# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3564 VSS a_1196_n1740# hgu_cdac_half_0.d<6> VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3565 a_n55487_7371# a_n55391_7113# hgu_tah_0.VDD hgu_tah_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.141 ps=1.33 w=0.42 l=0.15
X3566 VSS hgu_sarlogic_flat_0.x3.x20.Q_N a_2926_6078# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.101 ps=0.99 w=0.42 l=0.15
X3567 VSS VDD a_11720_7824# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.12 ps=1.08 w=0.42 l=0.15
X3568 a_16894_5688# a_15666_5316# a_16752_5310# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X3569 hgu_vgen_vref_0.mimtop2 VSS sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X3570 hgu_sarlogic_flat_0.x3.x5.X a_1863_9386# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3571 VSS a_11830_1153# a_11740_1179# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.116 ps=1.09 w=0.64 l=0.15
X3572 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3573 VSS a_n55304_6595# hgu_vgen_vref_0.phi2 VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3574 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3575 VDD a_7285_8487# a_7235_8795# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X3576 a_16894_5950# a_15666_5950# a_16752_6232# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X3577 a_14654_7663# hgu_sarlogic_flat_0.x5.eob a_14566_7525# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X3578 hgu_sarlogic_flat_0.x4.D[1] a_10870_6951# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X3579 a_5397_8106# a_4438_7824# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X3580 a_8288_6078# a_7369_6352# a_7842_6262# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X3581 a_19460_5284# a_19286_5688# a_19576_5676# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X3582 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_1.db<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3583 VSS async_delay_offset hgu_sarlogic_flat_0.x1.x2.x6.SW VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3584 hgu_cdac_half_1.VREF hgu_cdac_half_1.d<3> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<7:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3585 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3586 a_16113_12125# hgu_sarlogic_flat_0.x2.x2.x2.IN a_16041_12125# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X3587 a_6830_7824# hgu_sarlogic_flat_0.x3.x4.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3588 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X3589 a_4533_8513# a_4144_8513# a_4425_8879# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X3590 a_16113_6590# a_15832_6596# a_16020_6590# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X3591 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3592 a_17003_5688# a_15666_5316# a_16894_5688# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X3593 hgu_cdac_half_1.db<5> a_n3927_7727# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3594 a_4680_7798# a_4978_8098# a_4914_8190# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0924 ps=0.86 w=0.42 l=0.15
X3595 VSS hgu_cdac_half_0.db<6> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3596 a_6286_2234# a_6006_1868# a_6194_1868# VSS sky130_fd_pr__nfet_01v8 ad=0.0675 pd=0.735 as=0.066 ps=0.745 w=0.36 l=0.15
X3597 a_651_10968# VSS a_192_10793# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X3598 a_16113_5036# a_15666_4670# a_16020_4670# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X3599 VDD a_3960_3698# hgu_sarlogic_flat_0.x4.x9.A1 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3600 a_138_1363# a_n334_1153# a_382_1545# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X3601 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.db<6> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3602 a_4030_7798# a_4125_7798# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3603 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_0.d<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3604 a_9967_7798# a_10235_8008# a_10181_8106# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X3605 a_12359_7798# a_11614_7824# a_12495_7824# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3606 VSS a_16287_4644# a_16221_4670# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X3607 hgu_sarlogic_flat_0.x5.x2.x9.output_stack hgu_sarlogic_flat_0.x5.x2.x10.Y hgu_sarlogic_flat_0.x5.x2.x5[7].floating VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X3608 VSS a_12555_6925# a_12490_6951# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X3609 VDD a_2036_7824# hgu_sarlogic_flat_0.x3.x4.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3610 VSS a_16287_5284# a_16221_5688# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X3611 hgu_sarlogic_flat_0.x2.x1.x2.D a_2373_14732# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X3612 VDD retimer_delay_offset hgu_sarlogic_flat_0.x5.x2.x6.SW VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3613 hgu_sarlogic_flat_0.x4.x34.Q_N a_14404_2136# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X3614 hgu_cdac_half_1.d<6> a_n2219_8368# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3615 VSS hgu_cdac_sw_buffer_1.x4.X a_2206_n1100# VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3616 VDD a_3499_1331# hgu_cdac_sw_buffer_3.x4.A VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X3617 VSS hgu_sarlogic_flat_0.x5.x3.A a_20464_8879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0651 ps=0.73 w=0.42 l=0.15
X3618 a_n54850_7371# a_n54754_7113# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3619 hgu_cdac_half_1.hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT hgu_cdac_half_1.db<2> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.35
X3620 hgu_cdac_half_1.VREF hgu_cdac_half_1.db<5> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3621 a_4654_1153# a_3908_1179# a_4790_1179# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3622 VDD hgu_sarlogic_flat_0.x4.x15.S a_9708_2883# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.118 ps=1.4 w=0.42 l=0.15
X3623 a_2719_8513# a_2207_8487# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X3624 hgu_tah_0.VDD hgu_vgen_vref_0.phi2_n hgu_vgen_vref_0.mimtop1 hgu_tah_0.VDD sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=0.5
X3625 a_6286_2234# a_5840_1868# a_6194_1868# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0651 ps=0.73 w=0.42 l=0.15
X3626 a_n4429_7252# hgu_cdac_sw_buffer_3.x9.A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3627 a_18505_5310# a_18058_5316# a_18412_5310# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X3628 hgu_vgen_vref_0.mimtop1 hgu_vgen_vref_0.mimbot1 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X3629 VSS a_n2219_8368# hgu_cdac_half_1.d<6> VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3630 a_1325_11738# a_407_11578# a_879_11334# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3631 VSS hgu_cdac_half_0.d<6> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3632 hgu_cdac_sw_buffer_0.VDD a_n638_n245# hgu_cdac_sw_buffer_0.x3.X hgu_cdac_sw_buffer_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3633 VDD VDD a_5987_1153# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0956 pd=0.875 as=0.132 ps=1.22 w=0.42 l=0.15
X3634 VSS hgu_cdac_half_0.db<6> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3635 hgu_sarlogic_flat_0.x1.x2.x9.output_stack hgu_sarlogic_flat_0.x1.x2.x6.SW hgu_sarlogic_flat_0.x1.x2.x6.floating VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X3636 VSS VSS a_3977_6951# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3637 a_879_11334# a_407_11578# a_1123_11360# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X3638 a_n2219_8368# hgu_cdac_sw_buffer_2.x11.A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3639 a_n53930_7835# a_n53834_7657# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3640 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.d<6> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3641 VDD hgu_sarlogic_flat_0.x4.D[4] a_7759_1179# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X3642 a_14967_2556# hgu_sarlogic_flat_0.x4.x9.A1 a_14746_2883# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X3643 VSS hgu_sarlogic_flat_0.x4.x15.S a_9708_2883# VSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.109 ps=1.36 w=0.42 l=0.15
X3644 hgu_cdac_sw_buffer_2.x8.X a_n2025_7088# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3645 VDD a_8710_2530# a_8740_2883# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3646 hgu_sarlogic_flat_0.x2.x2.x1.x9.output_stack hgu_sarlogic_flat_0.x2.x2.x1.IN a_10575_15625# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X3647 VSS hgu_cdac_half_1.d<4> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<15:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3648 VSS hgu_cdac_half_1.d<5> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3649 VSS a_n3325_7252# hgu_cdac_sw_buffer_3.x4.X VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X3650 hgu_sarlogic_flat_0.x4.x2.X a_n424_3698# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3651 VDD a_1970_1842# a_1920_2150# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X3652 hgu_comp_flat_0.P hgu_tah_0.tah_vp a_n7660_7467# VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X3653 VDD a_18973_5510# a_18923_5310# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X3654 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<15:0> hgu_cdac_half_0.d<4> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3655 VSS hgu_cdac_half_1.d<5> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3656 a_9422_8106# a_9222_7824# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X3657 VSS hgu_cdac_half_0.d<5> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3658 VSS a_n335_1453# a_n334_1153# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3659 hgu_sarlogic_flat_0.x1.x4.x9.output_stack async_delay_offset hgu_sarlogic_flat_0.x1.x4.x7.floating VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X3660 a_9208_7317# a_8927_6951# a_9115_6951# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X3661 hgu_cdac_half_0.VREF hgu_cdac_half_0.d<6> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3662 a_17068_6564# a_16894_6968# a_17184_6956# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X3663 hgu_cdac_half_1.VREF hgu_cdac_half_1.d<6> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3664 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_1.db<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3665 VDD a_6516_6052# hgu_sarlogic_flat_0.x3.x57.Q_N VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X3666 VDD a_16581_4644# a_16531_4952# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X3667 hgu_sarlogic_flat_0.x5.x2.x5[7].floating hgu_sarlogic_flat_0.x5.x2.x10.Y hgu_sarlogic_flat_0.x5.x2.x9.output_stack VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X3668 VSS a_n55204_7371# a_n55391_7113# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X3669 hgu_cdac_half_0.db<6> a_n1158_n1744# hgu_cdac_sw_buffer_0.VDD hgu_cdac_sw_buffer_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3670 hgu_vgen_vref_0.mimtop2 VSS sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X3671 a_4141_1347# a_4449_1453# a_4398_1545# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0787 ps=0.795 w=0.42 l=0.15
X3672 a_10638_14512# hgu_sarlogic_flat_0.x2.x2.x1.IN a_10550_14374# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X3673 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_0.db<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3674 hgu_cdac_half_1.VREF hgu_cdac_half_1.db<6> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3675 VDD hgu_sarlogic_flat_0.x3.x5.X a_8762_8513# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3676 a_n55487_7835# a_n55391_7657# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3677 a_11154_2234# a_10790_1868# a_11070_2234# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X3678 VSS a_2323_11578# a_1945_11268# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X3679 a_5206_8513# a_4144_8513# a_5111_8513# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X3680 hgu_sarlogic_flat_0.x1.x2.x9.output_stack hgu_sarlogic_flat_0.x1.x2.x10.Y hgu_sarlogic_flat_0.x1.x2.x5[7].floating VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X3681 VDD a_2207_8487# a_2117_8879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X3682 a_9209_8879# a_8928_8513# a_9116_8513# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X3683 VDD a_4892_6925# a_4842_7233# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X3684 hgu_cdac_half_0.VREF hgu_cdac_half_0.db<5> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3685 VDD hgu_sarlogic_flat_0.x4.x20.S a_5897_7824# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0662 ps=0.735 w=0.42 l=0.15
X3686 a_1196_n1740# hgu_cdac_sw_buffer_1.x11.A hgu_cdac_sw_buffer_1.VDD hgu_cdac_sw_buffer_1.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3687 a_n6934_15288# hgu_comp_flat_0.ready a_n7022_15426# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X3688 hgu_cdac_sw_buffer_2.x3.A a_3165_1868# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X3689 VSS a_1945_11268# hgu_tah_0.sw VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3690 VSS a_n54752_8227# hgu_vgen_vref_0.phi1_n VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3691 a_18923_6232# a_18505_6316# a_18679_5924# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X3692 VDD hgu_sarlogic_flat_0.x2.x2.x1.IN a_9739_14835# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0651 ps=0.73 w=0.42 l=0.15
X3693 VDD a_4029_6052# hgu_sarlogic_flat_0.x4.D[6] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X3694 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3695 VDD a_4893_8487# a_4843_8795# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X3696 VSS VSS a_n4203_7087# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X3697 a_322_2883# a_140_2883# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X3698 hgu_cdac_sw_buffer_0.VDD a_n1240_n1104# hgu_cdac_sw_buffer_0.x11.A hgu_cdac_sw_buffer_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3699 VDD VSS a_n1473_7088# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3700 a_n542_11334# a_n447_11350# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X3701 a_2285_2234# a_1056_1868# a_2188_1868# VSS sky130_fd_pr__nfet_01v8 ad=0.0486 pd=0.63 as=0.116 ps=1.09 w=0.36 l=0.15
X3702 hgu_sarlogic_flat_0.x2.x3.Y VDD a_2323_10792# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X3703 hgu_tah_0.VDD a_n55304_8227# hgu_vgen_vref_0.phi1 hgu_tah_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3704 hgu_sarlogic_flat_0.x1.x4.x9.output_stack async_resetb_delay_cap_ctrl_code[2] hgu_sarlogic_flat_0.x1.x4.x4[3].floating VSS sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X3705 a_7485_2150# a_7069_2234# a_7228_2136# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.132 ps=1.22 w=0.84 l=0.15
X3706 a_10023_11461# hgu_sarlogic_flat_0.x2.x2.x3.IN VSS VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.0693 ps=0.75 w=0.42 l=0.15
X3707 VSS a_4836_2136# a_4784_1868# VSS sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.066 ps=0.745 w=0.42 l=0.15
X3708 VSS hgu_cdac_half_1.d<6> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3709 hgu_tah_0.tah_vp hgu_tah_0.sw_n vip hgu_tah_0.VDD sky130_fd_pr__pfet_01v8 ad=0.908 pd=5.83 as=0.908 ps=5.83 w=5.5 l=0.15
X3710 VSS hgu_cdac_half_0.d<6> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3711 a_n6959_12275# hgu_comp_flat_0.clk a_n7047_12137# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X3712 hgu_sarlogic_flat_0.x4.x9.S a_8479_8513# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X3713 a_0_1868# a_n1170_1868# a_n107_2234# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0486 ps=0.63 w=0.36 l=0.15
X3714 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<7:0> hgu_cdac_half_1.d<3> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3715 VSS hgu_cdac_half_1.db<6> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3716 a_14734_1545# a_14222_1153# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X3717 VSS hgu_cdac_half_0.db<6> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3718 a_n2219_8368# hgu_cdac_sw_buffer_2.x11.A VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3719 a_14654_7939# hgu_sarlogic_flat_0.x5.eob a_14566_7801# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X3720 a_16113_6590# a_15666_6596# a_16020_6590# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X3721 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.db<6> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3722 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.d<6> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3723 a_3894_2234# a_3614_1868# a_3802_1868# VSS sky130_fd_pr__nfet_01v8 ad=0.0675 pd=0.735 as=0.066 ps=0.745 w=0.36 l=0.15
X3724 hgu_cdac_half_0.d<6> a_1196_n1740# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3725 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3726 a_9739_15176# hgu_sarlogic_flat_0.x2.x2.x4.x9.output_stack hgu_sarlogic_flat_0.x2.x2.x1.IN VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.122 ps=1.42 w=0.42 l=0.15
X3727 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X3728 hgu_cdac_half_1.VREF hgu_cdac_half_1.d<6> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3729 VSS hgu_cdac_half_1.db<3> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<7:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.35
X3730 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<15:0> hgu_cdac_half_1.d<4> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3731 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_0.d<5> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3732 a_13667_1461# a_13476_1179# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X3733 a_6841_1453# hgu_sarlogic_flat_0.x4.x13.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3734 a_1516_1179# hgu_sarlogic_flat_0.x4.x2.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3735 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_1.d<5> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3736 a_9404_11849# hgu_sarlogic_flat_0.x2.x2.x3.IN a_9332_11987# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X3737 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X3738 hgu_cdac_half_0.VREF hgu_cdac_half_0.db<5> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3739 hgu_cdac_half_0.VREF hgu_cdac_half_0.db<6> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3740 a_3894_2234# a_3448_1868# a_3802_1868# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0651 ps=0.73 w=0.42 l=0.15
X3741 VDD hgu_sarlogic_flat_0.x4.D[1] a_11153_6951# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3742 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3743 a_12790_8795# a_12382_8513# a_12556_8487# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X3744 VDD hgu_sarlogic_flat_0.x3.x4.A a_2036_7824# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3745 VDD a_11206_7798# hgu_sarlogic_flat_0.x4.x15.S VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X3746 a_9739_14835# hgu_sarlogic_flat_0.x2.x2.x1.IN VDD VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3747 a_9382_6925# a_9208_7317# a_9522_6951# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X3748 VSS a_n1158_n1744# hgu_cdac_half_0.db<6> VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3749 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_0.db<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3750 a_8996_1868# a_9146_1842# a_8852_1842# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3751 hgu_sarlogic_flat_0.x2.x2.x1.x9.output_stack hgu_sarlogic_flat_0.x2.x2.x1.x6.SW hgu_sarlogic_flat_0.x2.x2.x1.x6.floating VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X3752 VSS hgu_cdac_sw_buffer_1.x11.A a_1196_n1740# VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3753 hgu_cdac_half_0.VREF hgu_cdac_half_0.d<6> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3754 VSS a_n1749_7728# hgu_cdac_half_1.d<5> VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3755 VSS hgu_cdac_half_1.d<6> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3756 a_12491_8513# a_11154_8513# a_12382_8513# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X3757 VDD a_n3049_7252# hgu_cdac_half_1.db<3> VDD sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3758 a_n424_3698# hgu_sarlogic_flat_0.x4.x3.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3759 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<15:0> hgu_cdac_half_1.d<4> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.122 ps=1.42 w=0.42 l=0.35
X3760 VSS hgu_cdac_half_1.db<4> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<15:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3761 a_11508_8513# hgu_sarlogic_flat_0.x4.x11.S VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X3762 a_6816_7317# a_6535_6951# a_6723_6951# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X3763 a_9316_6951# a_8927_6951# a_9208_7317# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X3764 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<15:0> hgu_cdac_half_0.db<4> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3765 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<7:0> hgu_cdac_half_0.db<3> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.122 ps=1.42 w=0.42 l=0.35
X3766 VSS VDD a_5319_7824# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.101 ps=0.99 w=0.42 l=0.15
X3767 VSS VDD a_1325_11738# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3768 a_1534_2530# hgu_sarlogic_flat_0.x4.x9.S VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X3769 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<15:0> hgu_cdac_half_1.d<4> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3770 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_1.d<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3771 VSS hgu_sarlogic_flat_0.x3.x33.Q_N a_10102_6078# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.101 ps=0.99 w=0.42 l=0.15
X3772 a_n54284_7835# hgu_vgen_vref_0.sky130_fd_sc_hd__dlymetal6s6s_1_2.A hgu_tah_0.VDD hgu_tah_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.141 ps=1.33 w=0.42 l=0.15
X3773 hgu_sarlogic_flat_0.x5.x1[7].Q_N a_19460_4644# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X3774 hgu_cdac_half_0.VREF hgu_cdac_half_0.d<5> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3775 a_2814_8513# a_1752_8513# a_2719_8513# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X3776 a_6817_8879# a_6536_8513# a_6724_8513# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X3777 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<15:0> hgu_cdac_half_1.db<4> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.122 ps=1.42 w=0.42 l=0.35
X3778 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_0.db<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3779 a_1534_2530# hgu_sarlogic_flat_0.x4.x9.S VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X3780 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_1.db<5> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3781 a_n1158_n1744# hgu_cdac_sw_buffer_0.x11.A hgu_cdac_sw_buffer_0.VDD hgu_cdac_sw_buffer_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3782 hgu_cdac_half_1.VREF hgu_cdac_half_1.db<4> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<15:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.35
X3783 hgu_sarlogic_flat_0.x3.x66.Q_N a_12555_6925# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X3784 VDD hgu_sarlogic_flat_0.x2.x7.A hgu_sarlogic_flat_0.x2.x7.Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3785 hgu_cdac_sw_buffer_1.VDD a_1114_n1100# hgu_cdac_sw_buffer_1.x11.A hgu_cdac_sw_buffer_1.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3786 hgu_cdac_half_0.VREF hgu_cdac_half_0.db<6> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3787 VSS hgu_comp_flat_0.clk a_1587_9386# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X3788 VDD a_1637_6052# hgu_sarlogic_flat_0.x4.x5.D VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X3789 a_2820_n241# hgu_cdac_sw_buffer_1.x5.A hgu_cdac_sw_buffer_1.VDD hgu_cdac_sw_buffer_1.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3790 hgu_cdac_half_0.VREF hgu_cdac_half_0.db<6> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3791 hgu_sarlogic_flat_0.x1.x4.x5[7].floating hgu_sarlogic_flat_0.x1.x4.x10.Y hgu_sarlogic_flat_0.x1.x4.x9.output_stack VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X3792 VDD hgu_sarlogic_flat_0.x5.x3.A a_20768_8628# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X3793 a_13570_1868# a_13016_1868# a_13462_2234# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0675 ps=0.735 w=0.36 l=0.15
X3794 a_6536_8513# a_6370_8513# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3795 hgu_vgen_vref_0.mimtop1 hgu_vgen_vref_0.mimbot1 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X3796 VSS a_2262_1153# a_2172_1179# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.116 ps=1.09 w=0.64 l=0.15
X3797 a_11684_7317# a_11153_6951# a_11600_7317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X3798 hgu_sarlogic_flat_0.x1.x2.x4[3].floating async_setb_delay_cap_ctrl_code[2] hgu_sarlogic_flat_0.x1.x2.x9.output_stack VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X3799 hgu_sarlogic_flat_0.x3.x36.Q_N a_12556_8487# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X3800 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X3801 hgu_sarlogic_flat_0.vdd_sw_b[7] a_52_2136# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X3802 hgu_cdac_sw_buffer_1.VDD a_1164_n241# hgu_cdac_sw_buffer_1.x9.X hgu_cdac_sw_buffer_1.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3803 hgu_cdac_half_0.VREF hgu_cdac_half_0.db<5> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3804 VSS hgu_cdac_sw_buffer_3.x11.A a_n4397_8367# VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3805 a_7574_6052# a_7842_6262# a_7788_6360# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X3806 VDD a_n424_3698# hgu_sarlogic_flat_0.x4.x2.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3807 VDD hgu_sarlogic_flat_0.x1.x9.Y a_n447_11350# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.123 ps=1.17 w=0.42 l=0.15
X3808 a_10710_13960# hgu_sarlogic_flat_0.x2.x2.x1.IN a_10638_13960# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X3809 VSS hgu_cdac_half_1.db<6> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3810 a_11685_8879# a_11154_8513# a_11601_8879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X3811 hgu_cdac_half_1.hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT hgu_cdac_half_1.d<2> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3812 hgu_tah_0.VDD a_n53364_7835# a_n53551_7657# hgu_tah_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X3813 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_0.db<5> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3814 a_2045_6078# hgu_sarlogic_flat_0.x3.x4.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3815 VSS hgu_cdac_half_0.d<5> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3816 VDD a_n1749_7728# hgu_cdac_half_1.d<5> VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3817 hgu_cdac_half_0.VREF hgu_cdac_half_0.d<6> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3818 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3819 a_18224_6596# a_18058_6596# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3820 a_19694_6232# a_19286_5950# a_19460_5924# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X3821 hgu_vgen_vref_0.mimtop2 VSS sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X3822 VSS hgu_cdac_half_1.d<5> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3823 a_8086_6078# a_7574_6052# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.084 ps=0.82 w=0.42 l=0.15
X3824 a_16448_15176# hgu_sarlogic_flat_0.x2.x2.x2.IN VSS VDD sky130_fd_pr__pfet_01v8_hvt ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3825 a_20464_8879# hgu_sarlogic_flat_0.x5.x2.x9.output_stack VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X3826 hgu_sarlogic_flat_0.x1.x2.x10.Y async_setb_delay_cap_ctrl_code[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3827 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_1.db<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3828 VDD a_2036_7824# hgu_sarlogic_flat_0.x3.x4.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3829 hgu_sarlogic_flat_0.x3.x20.Q_N a_2988_8487# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X3830 a_8288_6078# a_7370_6052# a_7842_6262# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3831 hgu_sarlogic_flat_0.x2.x2.x1.x9.output_stack sample_delay_cap_ctrl_code[6] hgu_sarlogic_flat_0.x2.x2.x1.x4[3].floating VSS sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X3832 hgu_cdac_half_1.VREF hgu_cdac_half_1.db<6> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3833 a_621_10615# hgu_sarlogic_flat_0.x5.eob VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X3834 VSS hgu_vgen_vref_0.sky130_fd_sc_hd__inv_1_2.A a_n55304_8227# VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3835 a_n55770_7835# a_n55674_7657# hgu_tah_0.VDD hgu_tah_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.141 ps=1.33 w=0.42 l=0.15
X3836 a_7502_6951# a_6990_6925# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X3837 a_18679_4644# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X3838 a_84_1461# a_n876_1179# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X3839 hgu_cdac_half_1.db<4> a_n3387_7727# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3840 VSS hgu_cdac_half_0.db<4> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<15:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3841 a_4533_2150# a_4068_1842# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X3842 VSS hgu_cdac_half_1.db<5> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3843 a_2287_6052# a_2585_6352# a_2521_6444# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0924 ps=0.86 w=0.42 l=0.15
X3844 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3845 hgu_vgen_vref_0.phi2 a_n55304_6595# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3846 hgu_sarlogic_flat_0.x1.x2.x9.output_stack hgu_sarlogic_flat_0.x1.x2.x10.Y hgu_sarlogic_flat_0.x1.x2.x5[7].floating VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X3847 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_0.db<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3848 hgu_cdac_sw_buffer_0.VDD hgu_cdac_sw_buffer_0.x11.A a_n1158_n1744# hgu_cdac_sw_buffer_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3849 hgu_vgen_vref_0.mimtop2 VSS sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X3850 hgu_sarlogic_flat_0.x2.x2.x4.x9.output_stack sample_delay_offset hgu_sarlogic_flat_0.x2.x2.x4.x7.floating VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X3851 a_19144_4952# a_18679_4644# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X3852 hgu_cdac_half_0.db<4> a_n148_n1104# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3853 VDD a_n716_1842# a_n806_2234# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X3854 hgu_comp_flat_0.ready a_n7678_6446# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0.244 ps=2.26 w=0.84 l=0.15
X3855 hgu_cdac_half_0.VREF hgu_cdac_half_0.db<6> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3856 VSS hgu_cdac_half_0.db<6> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3857 a_6604_1868# a_6754_1842# a_6460_1842# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3858 a_n6959_13485# hgu_comp_flat_0.ready a_n7047_13347# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X3859 hgu_sarlogic_flat_0.x3.x4.X a_2036_7824# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3860 VDD hgu_sarlogic_flat_0.x3.x3.A a_1422_7824# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3861 VSS a_3960_3698# hgu_sarlogic_flat_0.x4.x9.A1 VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3862 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.d<6> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3863 a_11317_1347# a_11625_1453# a_11574_1545# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0787 ps=0.795 w=0.42 l=0.15
X3864 a_7455_7233# a_6990_6925# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X3865 VSS hgu_cdac_half_1.d<6> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3866 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<7:0> hgu_cdac_half_1.db<3> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3867 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<7:0> hgu_cdac_half_0.db<3> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3868 hgu_cdac_sw_buffer_3.x11.X a_n4397_8367# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3869 VDD a_n2773_7252# hgu_cdac_half_1.db<2> VDD sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3870 a_6841_1453# hgu_sarlogic_flat_0.x4.x13.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3871 VSS hgu_cdac_half_1.d<6> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3872 VSS a_2373_14732# a_3080_14774# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X3873 a_6924_6951# a_6535_6951# a_6816_7317# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X3874 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X3875 VSS hgu_cdac_half_1.db<6> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3876 hgu_vgen_vref_0.mimtop1 hgu_vgen_vref_0.mimbot1 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X3877 a_n6526_6819# a_n6676_7789# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X3878 hgu_sarlogic_flat_0.x4.x23.Q_N a_4836_2136# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X3879 a_7456_8795# a_6991_8487# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X3880 a_18589_5310# a_18058_5316# a_18505_5310# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X3881 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3882 hgu_vgen_vref_0.mimtop1 hgu_vgen_vref_0.mimbot1 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X3883 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X3884 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_0.db<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3885 VDD a_n1287_2708# hgu_sarlogic_flat_0.x4.x6.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X3886 hgu_sarlogic_flat_0.x2.x2.x4.x3[1].floating sample_delay_cap_ctrl_code[1] hgu_sarlogic_flat_0.x2.x2.x4.x9.output_stack VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X3887 a_18589_6316# a_18058_5950# a_18505_6316# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X3888 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3889 hgu_sarlogic_flat_0.x4.x11.X a_5176_2883# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.113 ps=1.04 w=0.65 l=0.15
X3890 VSS hgu_sarlogic_flat_0.x3.x4.X a_7284_6925# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X3891 VSS VSS a_n412_n464# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X3892 hgu_cdac_half_0.VREF hgu_cdac_half_0.db<6> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3893 VDD hgu_sarlogic_flat_0.x4.x17.S a_3494_9752# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.138 ps=1.16 w=0.64 l=0.15
X3894 hgu_sarlogic_flat_0.x3.x69.Q_N a_10163_6925# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X3895 a_9332_12815# hgu_sarlogic_flat_0.x2.x2.x3.IN VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X3896 hgu_cdac_half_1.VREF hgu_cdac_half_1.db<6> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3897 VSS hgu_cdac_half_0.db<6> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3898 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<15:0> hgu_cdac_half_1.d<4> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3899 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_1.d<5> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3900 VSS a_8813_6052# hgu_sarlogic_flat_0.x4.D[4] VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X3901 a_2820_11667# hgu_sarlogic_flat_0.x2.x3.A hgu_sarlogic_flat_0.x2.x3.Y VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3902 a_n54284_7371# hgu_vgen_vref_0.sky130_fd_sc_hd__dlymetal6s6s_1_4.A hgu_tah_0.VDD hgu_tah_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.141 ps=1.33 w=0.42 l=0.15
X3903 hgu_cdac_half_1.d<4> a_n1209_7728# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3904 a_7771_6925# a_7597_6951# a_7887_6951# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X3905 a_16287_5284# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X3906 VSS hgu_sarlogic_flat_0.x4.x3.A a_n1058_3698# VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3907 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3908 hgu_sarlogic_flat_0.x3.x33.Q_N a_10164_8487# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X3909 a_11601_8879# a_11154_8513# a_11508_8513# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X3910 hgu_cdac_half_0.VREF hgu_cdac_half_0.db<4> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<15:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3911 a_16287_5924# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X3912 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<7:0> hgu_cdac_half_1.d<3> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3913 VDD hgu_cdac_sw_buffer_2.x11.A a_n2219_8368# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3914 VSS a_11775_8487# a_11709_8513# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X3915 VSS a_n2301_7728# hgu_cdac_sw_buffer_2.x11.A VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3916 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_0.db<5> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3917 a_16041_12263# hgu_sarlogic_flat_0.x2.x2.x2.IN a_15953_12263# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X3918 a_4144_8513# a_3978_8513# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3919 VDD a_2036_7824# hgu_sarlogic_flat_0.x3.x4.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3920 a_4978_6052# hgu_sarlogic_flat_0.x4.D[5] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3921 a_7368_1868# a_6754_1842# a_7228_2136# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3922 VDD a_19460_4644# a_20167_4670# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X3923 hgu_cdac_sw_buffer_0.VDD hgu_cdac_sw_buffer_0.x3.X a_n688_n1104# hgu_cdac_sw_buffer_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3924 VSS hgu_sarlogic_flat_0.x3.x5.X a_3978_8513# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3925 VSS a_n1240_n1104# hgu_cdac_sw_buffer_0.x11.A VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3926 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_0.d<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3927 a_5166_1545# a_4654_1153# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X3928 a_n890_2234# a_n1170_1868# a_n982_1868# VSS sky130_fd_pr__nfet_01v8 ad=0.0675 pd=0.735 as=0.066 ps=0.745 w=0.36 l=0.15
X3929 a_17302_5310# a_16894_5688# a_17068_5284# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X3930 a_12280_2883# a_12098_2883# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X3931 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X3932 a_12671_6951# hgu_sarlogic_flat_0.x3.x39.Q_N VSS VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X3933 a_5694_6078# a_5182_6052# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.084 ps=0.82 w=0.42 l=0.15
X3934 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3935 VSS hgu_sarlogic_flat_0.x4.x6.X a_n1336_1868# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3936 a_16448_14835# hgu_sarlogic_flat_0.x2.x2.x1.x9.output_stack hgu_sarlogic_flat_0.x2.x2.x2.IN VSS sky130_fd_pr__nfet_01v8 ad=0.0651 pd=0.73 as=0.122 ps=1.42 w=0.42 l=0.15
X3937 hgu_cdac_sw_buffer_3.x11.X a_n4397_8367# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3938 VDD a_19460_6564# a_20167_6606# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X3939 hgu_cdac_half_0.VREF hgu_cdac_half_0.d<5> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3940 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_1.d<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3941 VDD a_n4397_8367# hgu_cdac_sw_buffer_3.x11.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3942 hgu_cdac_half_1.VREF hgu_cdac_half_1.d<6> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3943 a_12671_6951# a_12068_6925# a_12555_6925# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3944 a_5896_6078# a_4978_6052# a_5450_6262# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3945 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_1.d<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3946 hgu_cdac_half_1.VREF hgu_cdac_half_1.db<6> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.35
X3947 a_n4429_7252# hgu_cdac_sw_buffer_3.x9.A VSS VSS sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3948 VDD hgu_sarlogic_flat_0.x5.x3.X a_15666_5950# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3949 hgu_cdac_sw_buffer_1.VDD a_1666_n1100# hgu_cdac_half_0.d<5> hgu_cdac_sw_buffer_1.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3950 VDD a_9438_1153# a_9371_1545# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X3951 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X3952 VSS hgu_cdac_half_0.db<4> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<15:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3953 VDD a_1945_11268# hgu_tah_0.sw VDD sky130_fd_pr__pfet_01v8 ad=0.391 pd=3.14 as=0.208 ps=1.59 w=1.26 l=0.15
X3954 VDD a_4125_7798# hgu_sarlogic_flat_0.x3.x48.Q_N VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X3955 a_n1699_7253# hgu_cdac_sw_buffer_2.x3.A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3956 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<7:0> hgu_cdac_half_0.db<3> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3957 VSS hgu_cdac_half_1.db<5> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3958 a_14679_9466# hgu_sarlogic_flat_0.x5.eob a_14591_9604# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X3959 a_18505_5036# a_18224_4670# a_18412_4670# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X3960 hgu_sarlogic_flat_0.x4.x2.X a_n424_3698# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3961 a_4099_1461# a_3908_1179# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X3962 a_16287_5284# a_16113_5310# a_16427_5676# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X3963 VSS hgu_cdac_half_1.d<5> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3964 VSS hgu_cdac_half_1.db<5> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3965 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_1.db<5> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3966 VDD hgu_sarlogic_flat_0.x2.x7.A a_3314_11664# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3967 a_9706_1363# a_9233_1453# a_9950_1179# VSS sky130_fd_pr__nfet_01v8 ad=0.0675 pd=0.735 as=0.0671 ps=0.75 w=0.36 l=0.15
X3968 a_16752_4952# a_16287_4644# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X3969 hgu_cdac_half_0.d<4> a_2206_n1100# hgu_cdac_sw_buffer_1.VDD hgu_cdac_sw_buffer_1.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3970 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.d<6> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3971 a_3222_8795# a_2814_8513# a_2988_8487# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X3972 VSS VDD a_7182_1179# VSS sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0974 ps=0.97 w=0.42 l=0.15
X3973 hgu_sarlogic_flat_0.x2.x2.x2.x9.output_stack sample_delay_cap_ctrl_code[10] hgu_sarlogic_flat_0.x2.x2.x2.x4[3].floating VSS sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X3974 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.db<6> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3975 VDD a_52_2136# a_n23_2234# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0956 pd=0.875 as=0.0787 ps=0.795 w=0.42 l=0.15
X3976 a_9523_8513# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X3977 a_n55770_7371# a_n55674_7113# hgu_tah_0.VDD hgu_tah_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.141 ps=1.33 w=0.42 l=0.15
X3978 a_3929_14650# hgu_sarlogic_flat_0.x2.x3.A a_3841_14650# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X3979 hgu_sarlogic_flat_0.x1.x4.x5[7].floating hgu_sarlogic_flat_0.x1.x4.x10.Y hgu_sarlogic_flat_0.x1.x4.x9.output_stack VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X3980 VSS hgu_sarlogic_flat_0.x3.x7.A a_1454_6950# VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3981 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<15:0> hgu_cdac_half_0.d<4> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.122 ps=1.42 w=0.42 l=0.35
X3982 VDD hgu_cdac_sw_buffer_2.x9.X a_n2301_7728# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3983 VSS hgu_sarlogic_flat_0.x3.x7.X a_8288_6078# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3984 a_13065_2708# VSS a_13207_2883# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X3985 a_2245_6360# a_2045_6078# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X3986 a_18819_4670# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X3987 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3988 a_14935_1179# a_14018_1153# a_14490_1363# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0675 ps=0.735 w=0.36 l=0.15
X3989 a_3007_2556# hgu_sarlogic_flat_0.x4.x9.A1 a_2786_2883# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X3990 VSS a_n54752_8227# hgu_vgen_vref_0.phi1_n VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3991 a_18819_5950# a_18973_5924# a_18679_5924# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3992 VSS hgu_cdac_half_0.d<5> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3993 a_3497_2708# hgu_sarlogic_flat_0.x4.x9.A1 a_3639_2556# VSS sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X3994 a_18819_5676# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X3995 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<15:0> hgu_cdac_half_1.db<4> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X3996 hgu_sarlogic_flat_0.x5.x1[2].Q_N a_17068_5924# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X3997 VSS a_n1058_3698# hgu_sarlogic_flat_0.x4.x3.X VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3998 a_8586_1868# hgu_sarlogic_flat_0.x4.D[3] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X3999 a_4001_14512# hgu_sarlogic_flat_0.x2.x3.A a_3929_14512# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X4000 VSS hgu_cdac_half_1.db<6> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X4001 a_4402_9386# a_3378_9360# a_3898_9386# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.072 ps=0.76 w=0.36 l=0.15
X4002 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X4003 hgu_sarlogic_flat_0.x3.x75.Q a_6086_6951# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X4004 VDD hgu_sarlogic_flat_0.x4.x6.X a_n1336_1868# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4005 a_9620_2136# hgu_sarlogic_flat_0.x4.x2.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.132 pd=1.22 as=0.0956 ps=0.875 w=0.42 l=0.15
X4006 VSS a_n7216_6420# hgu_comp_flat_0.comp_outp VSS sky130_fd_pr__nfet_01v8 ad=0.0759 pd=0.79 as=0.143 ps=1.54 w=0.46 l=0.15
X4007 hgu_cdac_half_0.d<4> a_2206_n1100# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4008 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X4009 VDD a_3960_3698# hgu_sarlogic_flat_0.x4.x9.A1 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4010 a_3960_3698# hgu_sarlogic_flat_0.x4.x30.A VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4011 a_13953_1179# a_13163_1153# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0703 ps=0.755 w=0.42 l=0.15
X4012 a_2285_14758# a_1137_14764# a_2199_15136# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X4013 hgu_comp_flat_0.comp_outn a_n6292_6446# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.3 as=0.139 ps=1.17 w=0.84 l=0.15
X4014 hgu_cdac_half_1.VREF hgu_cdac_half_1.d<3> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<7:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.35
X4015 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_1.db<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X4016 a_2207_8487# a_2033_8879# a_2347_8513# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X4017 VDD a_1886_14958# a_1836_14758# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X4018 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X4019 VDD a_n6526_6819# a_n7760_6349# VDD sky130_fd_pr__pfet_01v8 ad=0.139 pd=1.17 as=0.139 ps=1.17 w=0.84 l=0.15
X4020 VSS hgu_sarlogic_flat_0.x3.x4.X a_4892_6925# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X4021 VSS hgu_cdac_half_0.db<6> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X4022 a_n54284_7835# hgu_vgen_vref_0.sky130_fd_sc_hd__dlymetal6s6s_1_2.A VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X4023 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<1:0> hgu_cdac_half_0.db<1> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.122 ps=1.42 w=0.42 l=0.35
X4024 hgu_cdac_half_1.VREF hgu_cdac_half_1.d<6> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X4025 hgu_sarlogic_flat_0.x4.x7.S a_6087_8513# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X4026 VDD hgu_sarlogic_flat_0.x3.x36.Q_N a_12358_6052# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X4027 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<15:0> hgu_cdac_half_1.d<4> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X4028 a_n7678_6446# a_n7766_6446# a_n7678_6901# VSS sky130_fd_pr__nfet_01v8 ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.15
X4029 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X4030 VSS hgu_cdac_half_1.db<6> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X4031 hgu_cdac_half_1.d<6> a_n2219_8368# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4032 hgu_cdac_half_0.VREF hgu_cdac_half_0.db<4> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<15:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X4033 hgu_sarlogic_flat_0.x2.x2.x1.x9.output_stack sample_delay_cap_ctrl_code[6] hgu_sarlogic_flat_0.x2.x2.x1.x4[3].floating VSS sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X4034 a_4438_7824# hgu_sarlogic_flat_0.x3.x4.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X4035 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.db<6> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X4036 hgu_sarlogic_flat_0.x5.eob a_2914_9360# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.218 ps=1.97 w=0.65 l=0.15
X4037 a_16113_5310# a_15832_5316# a_16020_5310# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X4038 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<7:0> hgu_cdac_half_0.d<3> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X4039 hgu_sarlogic_flat_0.x1.x2.x9.output_stack hgu_comp_flat_0.ready a_n6959_14313# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X4040 a_19576_5950# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X4041 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X4042 VSS hgu_cdac_half_0.d<4> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<15:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X4043 hgu_cdac_half_1.hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT hgu_cdac_half_1.d<2> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.122 ps=1.42 w=0.42 l=0.35
X4044 a_16113_6316# a_15832_5950# a_16020_5950# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X4045 a_19191_4670# a_18679_4644# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X4046 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.d<6> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X4047 hgu_cdac_half_1.VREF hgu_cdac_half_1.db<4> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<15:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X4048 a_1752_8513# a_1586_8513# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4049 a_19576_6956# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X4050 a_n1287_2708# hgu_sarlogic_flat_0.x4.x9.A1 a_n1145_2556# VSS sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X4051 hgu_sarlogic_flat_0.x1.x2.x9.output_stack hgu_sarlogic_flat_0.x1.x2.x10.Y hgu_sarlogic_flat_0.x1.x2.x5[7].floating VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X4052 a_2586_6052# hgu_sarlogic_flat_0.x4.D[6] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4053 a_19576_5950# a_18973_5924# a_19460_5924# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4054 a_2117_8879# a_1586_8513# a_2033_8879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X4055 a_9900_8190# a_9763_7798# a_9464_7798# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X4056 hgu_sarlogic_flat_0.x3.x72.Q_N a_7771_6925# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X4057 VSS a_19460_4644# a_20167_4670# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X4058 a_2774_1545# a_2262_1153# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X4059 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X4060 a_7843_8008# a_7371_7798# a_8087_8190# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X4061 a_3518_9386# sel_bit[0] a_3408_9386# VSS sky130_fd_pr__nfet_01v8 ad=0.0786 pd=0.805 as=0.072 ps=0.76 w=0.36 l=0.15
X4062 hgu_sarlogic_flat_0.x5.x2.x5[7].floating hgu_sarlogic_flat_0.x5.x2.x10.Y hgu_sarlogic_flat_0.x5.x2.x9.output_stack VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X4063 VSS a_19460_5284# a_20167_5326# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X4064 a_3929_13822# hgu_sarlogic_flat_0.x2.x3.A a_3841_13822# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X4065 a_825_11360# a_n134_11726# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X4066 a_16041_12539# hgu_sarlogic_flat_0.x2.x2.x2.IN a_15953_12539# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X4067 hgu_tah_0.VDD a_n54284_7371# a_n54471_7113# hgu_tah_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X4068 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_0.d<5> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X4069 VDD a_1107_1331# hgu_cdac_sw_buffer_3.x3.A VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X4070 a_16427_5950# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X4071 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.122 ps=1.42 w=0.42 l=0.35
X4072 a_1161_10968# hgu_tah_0.sw VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X4073 hgu_cdac_half_0.d<6> a_1196_n1740# hgu_cdac_sw_buffer_1.VDD hgu_cdac_sw_buffer_1.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4074 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<15:0> hgu_cdac_half_1.db<4> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X4075 a_16427_6956# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X4076 a_18613_4670# a_18224_4670# a_18505_5036# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X4077 a_1707_1461# a_1516_1179# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X4078 hgu_sarlogic_flat_0.x5.x1[4].Q_N a_17068_5284# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X4079 hgu_vgen_vref_0.mimtop2 VSS sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X4080 VSS hgu_sarlogic_flat_0.x2.x1.x4.Y a_1886_14958# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X4081 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X4082 hgu_cdac_sw_buffer_0.VDD VSS a_n412_n464# hgu_cdac_sw_buffer_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X4083 VSS hgu_cdac_half_1.d<5> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X4084 a_n6676_7789# a_n6994_7879# hgu_comp_flat_0.P VSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X4085 a_13067_1331# a_13163_1153# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X4086 VSS hgu_cdac_half_0.db<5> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X4087 hgu_sarlogic_flat_0.x2.x2.x3.IN hgu_sarlogic_flat_0.x2.x2.x2.x9.output_stack a_10023_11664# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0651 ps=0.73 w=0.42 l=0.15
X4088 a_n55770_7835# a_n55674_7657# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X4089 a_4978_6052# hgu_sarlogic_flat_0.x4.D[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4090 hgu_tah_0.tah_vn hgu_tah_0.sw vin VSS sky130_fd_pr__nfet_01v8 ad=0.454 pd=3.08 as=0.454 ps=3.08 w=2.75 l=0.15
X4091 a_9902_7824# a_9762_8098# a_9464_7798# VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.0711 ps=0.755 w=0.36 l=0.15
X4092 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X4093 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_1.db<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X4094 a_13073_7824# a_12154_8098# a_12627_8008# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X4095 VDD a_16581_6790# a_17302_6590# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X4096 VDD a_19460_6564# a_19372_6590# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X4097 a_1564_2883# hgu_sarlogic_flat_0.x4.x9.A1 a_1105_2708# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X4098 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.db<6> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X4099 VSS a_n3049_7252# hgu_cdac_half_1.db<3> VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X4100 a_8927_6951# a_8761_6951# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4101 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X4102 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_1.d<5> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X4103 hgu_sarlogic_flat_0.x3.x7.X a_1454_6950# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4104 hgu_cdac_half_1.VREF hgu_cdac_half_1.db<5> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X4105 a_n6934_10748# hgu_comp_flat_0.clk a_n7022_10886# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X4106 VDD a_2373_14732# a_2285_14758# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X4107 VDD VDD a_18973_4644# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X4108 VSS hgu_cdac_half_0.d<6> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X4109 VDD a_18679_6564# a_18589_6590# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X4110 a_4124_6052# a_4679_6052# a_4637_6360# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0882 ps=1.05 w=0.84 l=0.15
X4111 VSS hgu_sarlogic_flat_0.x3.x7.X a_5896_6078# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4112 VSS a_1534_2530# a_1468_2556# VSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X4113 a_4679_6052# a_4978_6052# a_4913_6078# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.066 ps=0.745 w=0.36 l=0.15
X4114 VSS a_20768_8628# hgu_sarlogic_flat_0.x5.x3.X VSS sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X4115 VDD a_3960_3698# hgu_sarlogic_flat_0.x4.x9.A1 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4116 hgu_sarlogic_flat_0.x4.x9.A1 a_3960_3698# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4117 hgu_cdac_sw_buffer_1.VDD hgu_cdac_sw_buffer_1.x9.X a_1114_n1100# hgu_cdac_sw_buffer_1.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4118 hgu_sarlogic_flat_0.x4.x17.X a_12352_2883# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.113 ps=1.04 w=0.65 l=0.15
X4119 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_1.db<5> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X4120 a_8813_6052# a_8908_6052# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X4121 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<15:0> hgu_cdac_half_0.d<4> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.35
X4122 a_5987_1153# a_6533_1347# a_6491_1461# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.132 pd=1.22 as=0.0882 ps=1.05 w=0.84 l=0.15
X4123 a_9620_2136# a_9461_2234# a_9760_1868# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.109 ps=1.03 w=0.64 l=0.15
X4124 a_19460_4644# a_19286_4670# a_19576_4670# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X4125 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.d<6> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X4126 VSS hgu_cdac_half_0.db<3> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<7:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.35
X4127 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X4128 hgu_cdac_half_0.VREF hgu_cdac_half_0.d<5> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X4129 a_1019_10793# hgu_sarlogic_flat_0.x1.x3.A0 a_1161_10968# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X4130 a_14329_2234# a_13016_1868# a_14245_2234# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0787 pd=0.795 as=0.0567 ps=0.69 w=0.42 l=0.15
X4131 a_9461_2234# a_8398_1868# a_9317_2150# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X4132 VDD VDD a_16581_5510# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X4133 VDD hgu_sarlogic_flat_0.x4.x20.S a_14960_2883# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.0767 ps=0.785 w=0.42 l=0.15
X4134 hgu_cdac_sw_buffer_0.VDD a_n148_n1104# hgu_cdac_half_0.db<4> hgu_cdac_sw_buffer_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4135 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X4136 a_16088_10874# hgu_sarlogic_flat_0.x2.x2.x2.IN a_16000_10736# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X4137 a_4598_6925# hgu_sarlogic_flat_0.x3.x77.Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X4138 VDD VDD a_9438_1153# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X4139 a_7030_8106# a_6830_7824# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X4140 VDD a_n1147_7253# hgu_cdac_sw_buffer_2.x4.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X4141 VDD a_n424_3698# hgu_sarlogic_flat_0.x4.x2.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4142 hgu_sarlogic_flat_0.x3.x27.D a_3695_8513# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X4143 VSS hgu_cdac_half_1.db<1> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<1:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.35
X4144 result[0] a_17775_6606# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X4145 a_3504_6078# a_2585_6352# a_3058_6262# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X4146 a_9348_1179# a_9233_1453# a_8925_1347# VSS sky130_fd_pr__nfet_01v8 ad=0.116 pd=1.09 as=0.0486 ps=0.63 w=0.36 l=0.15
X4147 VSS hgu_cdac_half_0.db<6> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X4148 VSS hgu_sarlogic_flat_0.x4.x20.S a_14967_2556# VSS sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.0693 ps=0.75 w=0.42 l=0.15
X4149 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.d<6> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X4150 VDD hgu_sarlogic_flat_0.x2.x1.x4.Y a_1886_14958# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X4151 VSS hgu_sarlogic_flat_0.x3.x33.Q_N a_9327_6078# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.12 ps=1.08 w=0.42 l=0.15
X4152 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.db<6> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X4153 a_1610_1868# a_1056_1868# a_1502_2234# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0675 ps=0.735 w=0.36 l=0.15
X4154 a_14746_2883# VSS a_14746_2556# VSS sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X4155 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.db<6> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X4156 a_4599_8487# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X4157 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.d<6> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X4158 a_12154_6052# hgu_sarlogic_flat_0.x4.D[2] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4159 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X4160 a_14544_1868# a_13930_1842# a_14404_2136# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4161 VDD hgu_comp_flat_0.ready a_n7022_15702# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X4162 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.db<6> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X4163 VSS hgu_sarlogic_flat_0.x3.x5.X a_11154_8513# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4164 VDD a_2036_7824# hgu_sarlogic_flat_0.x3.x4.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4165 a_n3049_7252# hgu_cdac_sw_buffer_3.x6.A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X4166 a_16531_6232# a_16113_6316# a_16287_5924# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X4167 a_16221_5950# a_15832_5950# a_16113_6316# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X4168 hgu_vgen_vref_0.mimtop1 hgu_vgen_vref_0.mimbot1 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X4169 a_10710_14236# hgu_sarlogic_flat_0.x2.x2.x1.IN a_10638_14236# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X4170 VSS a_n55304_8227# hgu_vgen_vref_0.phi1 VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4171 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<15:0> hgu_cdac_half_0.d<4> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X4172 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<7:0> hgu_cdac_half_0.d<3> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X4173 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_0.db<5> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X4174 VSS a_13065_2708# hgu_sarlogic_flat_0.x4.x18.X VSS sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X4175 VSS a_1196_n1740# hgu_cdac_half_0.d<6> VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4176 VDD a_2501_8487# a_2451_8795# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X4177 hgu_sarlogic_flat_0.x3.x75.Q_N a_5379_6925# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X4178 a_12572_6360# a_11613_6078# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X4179 hgu_cdac_half_0.VREF hgu_cdac_half_0.d<4> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<15:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X4180 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X4181 VSS a_n54284_7835# a_n54471_7657# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X4182 hgu_cdac_half_1.db<4> a_n3387_7727# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4183 hgu_comp_flat_0.comp_outp a_n7216_6420# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.139 pd=1.17 as=0.139 ps=1.17 w=0.84 l=0.15
X4184 VSS hgu_sarlogic_flat_0.x1.x9.Y a_n28_11682# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.12 ps=1.08 w=0.42 l=0.15
X4185 VDD a_n4397_8367# hgu_cdac_sw_buffer_3.x11.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4186 a_5451_8008# a_4979_7798# a_5695_8190# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X4187 VDD VDD a_8909_7798# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.123 ps=1.17 w=0.42 l=0.15
X4188 hgu_sarlogic_flat_0.x5.x2.x4[3].floating retimer_delay_code[2] hgu_sarlogic_flat_0.x5.x2.x9.output_stack VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X4189 hgu_cdac_half_0.VREF hgu_cdac_half_0.db<2> hgu_cdac_half_0.hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.35
X4190 a_10397_7233# a_9989_6951# a_10163_6925# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X4191 hgu_cdac_half_0.VREF hgu_cdac_half_0.db<6> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X4192 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X4193 hgu_sarlogic_flat_0.x2.x2.x4.x10.Y sample_delay_cap_ctrl_code[3] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X4194 a_747_11682# a_879_11334# a_611_11594# VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0864 ps=0.91 w=0.64 l=0.15
X4195 a_10638_14098# hgu_sarlogic_flat_0.x2.x2.x1.IN a_10550_14098# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X4196 a_n6887_12551# hgu_comp_flat_0.clk a_n6959_12689# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X4197 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X4198 a_9697_6444# a_8908_6052# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0819 ps=0.81 w=0.42 l=0.15
X4199 a_18613_6968# a_18224_6596# a_18505_6590# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X4200 hgu_sarlogic_flat_0.x2.x2.x3.x9.output_stack sample_delay_cap_ctrl_code[13] hgu_sarlogic_flat_0.x2.x2.x3.x3[1].floating VSS sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X4201 a_16113_12677# hgu_sarlogic_flat_0.x2.x2.x2.IN a_16041_12815# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X4202 a_10398_8795# a_9990_8513# a_10164_8487# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X4203 VDD hgu_sarlogic_flat_0.x3.x4.X a_12069_8487# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X4204 a_n3877_7252# hgu_cdac_sw_buffer_3.x3.A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X4205 a_17068_5924# a_16894_5950# a_17184_5950# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X4206 hgu_cdac_half_0.hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT hgu_cdac_half_0.d<2> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.122 ps=1.42 w=0.42 l=0.35
X4207 hgu_sarlogic_flat_0.x2.x2.x2.x4[3].floating sample_delay_cap_ctrl_code[10] hgu_sarlogic_flat_0.x2.x2.x2.x9.output_stack VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X4208 a_9899_6444# a_9762_6052# a_9463_6052# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X4209 a_9182_1545# a_8379_1153# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0787 pd=0.795 as=0.0956 ps=0.875 w=0.42 l=0.15
X4210 VDD a_n2219_8368# hgu_cdac_half_1.d<6> VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4211 a_n1149_14701# hgu_sarlogic_flat_0.x1.x2.x9.output_stack hgu_sarlogic_flat_0.x1.x9.A VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.122 ps=1.42 w=0.42 l=0.15
X4212 VSS hgu_cdac_half_1.d<6> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X4213 a_10675_1331# a_10771_1153# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X4214 a_n134_11726# hgu_sarlogic_flat_0.x1.x10.Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X4215 a_2586_6052# hgu_sarlogic_flat_0.x4.D[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4216 a_8692_1179# hgu_sarlogic_flat_0.x4.x2.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.17 pd=1.81 as=0.154 ps=1.34 w=0.64 l=0.15
X4217 result[7] a_20167_4670# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X4218 a_1716_n241# hgu_cdac_sw_buffer_1.x3.A hgu_cdac_sw_buffer_1.VDD hgu_cdac_sw_buffer_1.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X4219 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_0.db<5> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X4220 VSS hgu_cdac_half_1.db<6> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X4221 a_10681_7824# a_9762_8098# a_10235_8008# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X4222 VDD a_3926_2530# a_3956_2883# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X4223 a_879_11334# a_406_11482# a_1123_11726# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0671 ps=0.75 w=0.36 l=0.15
X4224 hgu_vgen_vref_0.sky130_fd_sc_hd__inv_1_3.A hgu_vgen_vref_0.sky130_fd_sc_hd__inv_1_1.A VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X4225 VSS a_n2773_7252# hgu_cdac_half_1.db<2> VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X4226 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_1.d<5> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X4227 VSS hgu_cdac_half_1.db<6> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X4228 a_10099_8513# a_8762_8513# a_9990_8513# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X4229 VSS VDD a_16581_4644# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X4230 VSS VDD a_6754_1842# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X4231 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<7:0> hgu_cdac_half_1.db<3> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X4232 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.db<6> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X4233 VSS EXT_CLK a_971_14764# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4234 hgu_sarlogic_flat_0.x4.D[2] a_13262_6951# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X4235 hgu_cdac_sw_buffer_2.x11.A a_n2301_7728# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4236 VSS VDD a_16581_5510# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X4237 VSS a_14404_2136# a_15125_1868# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X4238 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X4239 a_11244_1842# a_11070_2234# a_11388_1868# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.0974 ps=0.97 w=0.64 l=0.15
X4240 a_1325_14758# hgu_sarlogic_flat_0.x2.x1.x2.D VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X4241 hgu_cdac_half_1.VREF hgu_cdac_half_1.d<5> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X4242 VDD a_n6994_7879# a_n6676_7789# VDD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X4243 a_13073_7824# a_12155_7798# a_12627_8008# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4244 VSS a_2206_n1100# hgu_cdac_half_0.d<4> VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4245 hgu_cdac_half_0.VREF hgu_cdac_half_0.d<6> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X4246 a_5367_1179# a_4450_1153# a_4922_1363# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0675 ps=0.735 w=0.36 l=0.15
X4247 a_6990_6925# a_6816_7317# a_7130_6951# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X4248 a_11914_6951# a_12068_6925# a_11774_6925# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4249 VSS a_8852_1842# a_8786_1868# VSS sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0671 ps=0.75 w=0.42 l=0.15
X4250 VSS a_1422_7824# hgu_sarlogic_flat_0.x3.x4.A VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4251 hgu_cdac_sw_buffer_1.VDD a_1196_n1740# hgu_cdac_half_0.d<6> hgu_cdac_sw_buffer_1.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4252 VSS a_n130_1153# a_n220_1179# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.116 ps=1.09 w=0.64 l=0.15
X4253 hgu_sarlogic_flat_0.x1.x4.x4[3].floating async_resetb_delay_cap_ctrl_code[2] hgu_sarlogic_flat_0.x1.x4.x9.output_stack VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X4254 VSS hgu_cdac_half_1.d<3> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<7:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X4255 a_2544_n241# hgu_cdac_sw_buffer_1.x6.A hgu_cdac_sw_buffer_1.VDD hgu_cdac_sw_buffer_1.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X4256 VSS hgu_sarlogic_flat_0.x1.x10.A a_n1149_11335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0651 ps=0.73 w=0.42 l=0.15
X4257 a_2914_9360# sel_bit[1] a_3408_9386# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0729 pd=0.81 as=0.14 ps=1.6 w=0.54 l=0.15
X4258 VSS hgu_cdac_half_0.d<2> hgu_cdac_half_0.hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT VSS sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.35
X4259 a_11178_1868# a_10624_1868# a_11070_2234# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0675 ps=0.735 w=0.36 l=0.15
X4260 hgu_tah_0.VDD a_n53647_7835# a_n53834_7657# hgu_tah_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X4261 a_8909_7798# a_9464_7798# a_9422_8106# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0882 ps=1.05 w=0.84 l=0.15
X4262 a_4385_1179# a_3595_1153# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0703 ps=0.755 w=0.42 l=0.15
X4263 VDD a_n3927_7727# hgu_cdac_half_1.db<5> VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4264 a_6956_1179# a_6841_1453# a_6533_1347# VSS sky130_fd_pr__nfet_01v8 ad=0.116 pd=1.09 as=0.0486 ps=0.63 w=0.36 l=0.15
X4265 a_n6959_11861# hgu_comp_flat_0.clk a_n7047_11861# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X4266 a_9379_10322# hgu_sarlogic_flat_0.x2.x2.x3.IN VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X4267 VDD a_2914_9360# hgu_sarlogic_flat_0.x5.eob VDD sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X4268 VDD a_2036_7824# hgu_sarlogic_flat_0.x3.x4.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4269 a_n7660_7467# hgu_tah_0.tah_vn hgu_comp_flat_0.Q VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X4270 a_n23_2234# a_n1336_1868# a_n107_2234# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0787 pd=0.795 as=0.0567 ps=0.69 w=0.42 l=0.15
X4271 VDD hgu_sarlogic_flat_0.x3.x20.Q_N a_2790_6052# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X4272 hgu_sarlogic_flat_0.x4.x3.X a_n1058_3698# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4273 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.d<6> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X4274 VSS a_n53364_7371# a_n53551_7113# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X4275 hgu_cdac_sw_buffer_0.VDD a_n688_n1104# hgu_cdac_half_0.db<5> hgu_cdac_sw_buffer_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4276 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.db<6> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X4277 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_0.db<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X4278 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.d<6> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X4279 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.db<6> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X4280 a_9989_6951# a_8761_6951# a_9847_7233# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X4281 VSS a_3326_3698# hgu_sarlogic_flat_0.x4.x30.A VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4282 hgu_cdac_half_0.db<6> a_n1158_n1744# hgu_cdac_sw_buffer_0.VDD hgu_cdac_sw_buffer_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4283 VDD a_1019_10793# hgu_sarlogic_flat_0.x1.x3.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X4284 hgu_cdac_sw_buffer_3.x11.X a_n4397_8367# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4285 hgu_tah_0.tah_vp hgu_tah_0.sw hgu_tah_0.tah_vp hgu_tah_0.VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.908 ps=5.83 w=5.5 l=0.15
X4286 VSS hgu_cdac_half_0.d<6> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X4287 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_1.db<5> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X4288 a_18224_5316# a_18058_5316# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4289 VSS a_10673_2708# hgu_sarlogic_flat_0.x4.x16.X VSS sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X4290 hgu_cdac_half_1.VREF hgu_cdac_half_1.db<6> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X4291 a_4738_6951# hgu_sarlogic_flat_0.x3.x77.Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X4292 a_1196_n1740# hgu_cdac_sw_buffer_1.x11.A hgu_cdac_sw_buffer_1.VDD hgu_cdac_sw_buffer_1.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4293 a_9652_1461# a_8692_1179# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X4294 a_334_10641# hgu_sarlogic_flat_0.x5.eob VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X4295 a_9990_8513# a_8762_8513# a_9848_8795# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X4296 VSS hgu_cdac_half_0.d<4> hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<15:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X4297 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<15:0> hgu_cdac_half_1.db<4> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X4298 a_394_2883# hgu_sarlogic_flat_0.x4.x9.A1 a_322_2883# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X4299 a_1137_14764# a_971_14764# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4300 hgu_vgen_vref_0.mimtop2 VSS sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X4301 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<1:0> hgu_cdac_half_1.d<1> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.35
X4302 hgu_sarlogic_flat_0.x4.x2.X a_n424_3698# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4303 hgu_cdac_sw_buffer_0.VDD a_n1158_n1744# hgu_cdac_half_0.db<6> hgu_cdac_sw_buffer_0.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4304 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<15:0> hgu_cdac_half_0.d<4> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X4305 VDD a_6754_1842# a_7485_2150# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X4306 a_11205_6052# a_11300_6052# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X4307 a_12012_2136# a_11853_2234# a_12152_1868# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.109 ps=1.03 w=0.64 l=0.15
X4308 a_7371_7798# hgu_sarlogic_flat_0.x3.x5.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4309 a_394_2556# a_140_2883# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.145 ps=1.11 w=0.42 l=0.15
X4310 hgu_cdac_sw_buffer_1.VDD hgu_cdac_sw_buffer_1.x11.A a_1196_n1740# hgu_cdac_sw_buffer_1.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4311 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_1.db<5> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.35
X4312 hgu_sarlogic_flat_0.x2.x2.x2.x9.output_stack hgu_sarlogic_flat_0.x2.x2.x2.x10.Y hgu_sarlogic_flat_0.x2.x2.x2.x5[7].floating VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X4313 hgu_comp_flat_0.P hgu_tah_0.tah_vp a_n7660_7467# VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.31 ps=2.62 w=1 l=0.15
X4314 VDD a_7228_2136# a_7949_1868# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X4315 a_12154_6052# hgu_sarlogic_flat_0.x4.D[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4316 hgu_cdac_half_0.d<4> a_2206_n1100# hgu_cdac_sw_buffer_1.VDD hgu_cdac_sw_buffer_1.VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4317 hgu_vgen_vref_0.mimbot1 hgu_vgen_vref_0.phi2_n hgu_vgen_vref_0.mimtop2 hgu_tah_0.VDD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=0.5
X4318 a_11507_6951# hgu_sarlogic_flat_0.x3.x7.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X4319 a_7574_6052# a_6829_6078# a_7710_6078# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4320 a_8283_1331# a_8379_1153# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X4321 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<7:0> hgu_cdac_half_1.db<3> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X4322 a_n924_2556# VSS a_n1287_2708# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X4323 hgu_vgen_vref_0.mimtop1 hgu_vgen_vref_0.mimbot1 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X4324 VSS a_13163_1153# hgu_sarlogic_flat_0.x4.x35.Q_N VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X4325 a_6790_1545# a_5987_1153# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0787 pd=0.795 as=0.0956 ps=0.875 w=0.42 l=0.15
X4326 hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_half_0.db<5> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X4327 VDD hgu_sarlogic_flat_0.x3.x33.Q_N a_8908_6052# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.123 ps=1.17 w=0.42 l=0.15
X4328 hgu_vgen_vref_0.mimtop1 hgu_vgen_vref_0.mimbot1 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X4329 hgu_cdac_sw_buffer_2.x4.A a_5557_1868# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X4330 VSS hgu_cdac_half_1.d<6> hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X4331 a_11508_8513# hgu_sarlogic_flat_0.x4.x11.S VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X4332 VSS a_n1058_3698# hgu_sarlogic_flat_0.x4.x3.X VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4333 hgu_cdac_half_0.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_0.d<6> VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X4334 hgu_tah_0.VDD VSS sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X4335 hgu_cdac_half_0.hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT hgu_cdac_half_0.d<2> hgu_cdac_half_0.VREF hgu_cdac_half_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.35
X4336 a_n770_1179# a_n643_1347# a_n1189_1153# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.03 as=0.0864 ps=0.91 w=0.64 l=0.15
X4337 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<0> hgu_cdac_half_1.db<0> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.244 ps=2.26 w=0.84 l=0.35
X4338 VSS hgu_cdac_half_1.db<6> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X4339 hgu_cdac_half_0.d<6> a_1196_n1740# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4340 a_1732_15124# a_1886_14958# a_1592_14732# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4341 VDD VDD a_9967_7798# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X4342 a_138_1363# a_n335_1453# a_382_1179# VSS sky130_fd_pr__nfet_01v8 ad=0.0675 pd=0.735 as=0.0671 ps=0.75 w=0.36 l=0.15
X4343 hgu_cdac_half_1.hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_half_1.d<6> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X4344 VSS hgu_cdac_half_1.db<5> hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.35
X4345 VDD a_12068_6925# a_12789_7233# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X4346 a_13163_1153# a_13709_1347# a_13667_1461# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.132 pd=1.22 as=0.0882 ps=1.05 w=0.84 l=0.15
X4347 a_2057_1453# hgu_sarlogic_flat_0.x4.x9.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4348 VSS hgu_cdac_half_0.db<5> hgu_cdac_half_0.hgu_cdac_8bit_array_2.drv<31:0> VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X4349 VDD a_11244_1842# a_11154_2234# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X4350 a_5117_6078# a_4977_6352# a_4679_6052# VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.0711 ps=0.755 w=0.36 l=0.15
X4351 VDD a_9966_6052# a_9899_6444# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X4352 hgu_cdac_half_1.hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_half_1.db<6> hgu_cdac_half_1.VREF hgu_cdac_half_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X4353 VDD a_3960_3698# hgu_sarlogic_flat_0.x4.x9.A1 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4354 hgu_vgen_vref_0.vcm VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
.ends

