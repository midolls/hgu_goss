* NGSPICE file created from hgu_comp_flat.ext - technology: sky130A

.subckt hgu_comp_flat cdac_vn cdac_vp clk comp_outp comp_outn ready VDD VSS
X0 Q cdac_vn a_582_n702# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1 ready a_564_n1721# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0.244 ps=2.26 w=0.84 l=0.15
X2 a_564_n1721# a_476_n1721# a_564_n1266# VSS sky130_fd_pr__nfet_01v8 ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.15
X3 comp_outn a_1950_n1721# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.3 as=0.139 ps=1.17 w=0.84 l=0.15
X4 a_582_n702# cdac_vn Q VSS sky130_fd_pr__nfet_01v8_lvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X5 a_1950_n1721# RS_n VDD VDD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0.244 ps=2.26 w=0.84 l=0.15
X6 a_482_n1818# a_1716_n1348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0759 pd=0.79 as=0.143 ps=1.54 w=0.46 l=0.15
X7 a_564_n1721# a_482_n1818# a_476_n1721# VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.15
X8 VDD a_1026_n1747# comp_outp VDD sky130_fd_pr__pfet_01v8 ad=0.139 pd=1.17 as=0.26 ps=2.3 w=0.84 l=0.15
X9 VSS RS_p a_1026_n1747# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X10 VDD clk a_1248_n288# VDD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X11 a_674_n702# cdac_vp a_582_n702# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.165 pd=1.33 as=0.31 ps=2.62 w=1 l=0.15
X12 VDD a_852_n296# a_476_n1721# VDD sky130_fd_pr__pfet_01v8 ad=0.139 pd=1.17 as=0.26 ps=2.3 w=0.84 l=0.15
X13 comp_outp a_1026_n1747# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.139 pd=1.17 as=0.139 ps=1.17 w=0.84 l=0.15
X14 a_476_n1721# a_852_n296# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.139 pd=1.17 as=0.139 ps=1.17 w=0.84 l=0.15
X15 a_582_n702# cdac_vn Q VSS sky130_fd_pr__nfet_01v8_lvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X16 a_582_n702# cdac_vp a_674_n702# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X17 comp_outn a_1950_n1721# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.54 as=0.0759 ps=0.79 w=0.46 l=0.15
X18 VDD RS_p a_1026_n1747# VDD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0.244 ps=2.26 w=0.84 l=0.15
X19 VDD a_852_n296# a_476_n1721# VDD sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.3 as=0.139 ps=1.17 w=0.84 l=0.15
X20 a_674_n702# cdac_vp a_582_n702# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X21 Q cdac_vn a_582_n702# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X22 a_564_n1266# a_482_n1818# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.15
X23 VSS a_1026_n1747# comp_outp VSS sky130_fd_pr__nfet_01v8 ad=0.0759 pd=0.79 as=0.143 ps=1.54 w=0.46 l=0.15
X24 a_1950_n1721# RS_n VSS VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X25 a_1566_n378# clk VDD VDD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X26 VSS a_852_n296# a_476_n1721# VSS sky130_fd_pr__nfet_01v8 ad=0.0759 pd=0.79 as=0.143 ps=1.54 w=0.46 l=0.15
X27 VDD a_1248_n288# a_852_n296# VDD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0.244 ps=2.26 w=0.84 l=0.15
X28 a_482_n1818# a_1716_n1348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.54 as=0.0759 ps=0.79 w=0.46 l=0.15
X29 a_582_n702# clk VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X30 comp_outp a_1026_n1747# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0759 pd=0.79 as=0.0759 ps=0.79 w=0.46 l=0.15
X31 VSS a_1248_n288# a_852_n296# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X32 a_674_n702# cdac_vp a_582_n702# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X33 a_582_n702# cdac_vn Q VSS sky130_fd_pr__nfet_01v8_lvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X34 a_1248_n288# a_1566_n378# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X35 Q clk VDD VDD sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X36 a_582_n702# cdac_vp a_674_n702# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X37 VDD a_1026_n1747# comp_outp VDD sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.3 as=0.139 ps=1.17 w=0.84 l=0.15
X38 RS_n a_1716_n1348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.15
X39 comp_outn a_1950_n1721# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.139 pd=1.17 as=0.26 ps=2.3 w=0.84 l=0.15
X40 a_1716_n1348# a_1566_n378# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X41 VSS a_1716_n1348# a_482_n1818# VSS sky130_fd_pr__nfet_01v8 ad=0.0759 pd=0.79 as=0.0759 ps=0.79 w=0.46 l=0.15
X42 VSS clk a_582_n702# VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.31 ps=2.62 w=1 l=0.15
X43 a_582_n702# cdac_vn Q VSS sky130_fd_pr__nfet_01v8_lvt ad=0.31 pd=2.62 as=0.165 ps=1.33 w=1 l=0.15
X44 VSS a_852_n296# a_476_n1721# VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.54 as=0.0759 ps=0.79 w=0.46 l=0.15
X45 Q a_1566_n378# a_1248_n288# VSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X46 Q cdac_vn a_582_n702# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.165 pd=1.33 as=0.31 ps=2.62 w=1 l=0.15
X47 RS_n RS_p VDD VDD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.15
X48 VDD a_1950_n1721# comp_outn VDD sky130_fd_pr__pfet_01v8 ad=0.139 pd=1.17 as=0.139 ps=1.17 w=0.84 l=0.15
X49 a_1716_n1348# a_1566_n378# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0.244 ps=2.26 w=0.84 l=0.15
X50 a_582_n702# clk VSS VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.165 ps=1.33 w=1 l=0.15
X51 VDD clk a_674_n702# VDD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X52 a_674_n702# cdac_vp a_582_n702# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X53 VSS a_1026_n1747# comp_outp VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.54 as=0.0759 ps=0.79 w=0.46 l=0.15
X54 comp_outn a_1950_n1721# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0759 pd=0.79 as=0.143 ps=1.54 w=0.46 l=0.15
X55 a_482_n1818# a_1716_n1348# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.139 pd=1.17 as=0.26 ps=2.3 w=0.84 l=0.15
X56 a_482_n1818# a_1716_n1348# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.3 as=0.139 ps=1.17 w=0.84 l=0.15
X57 a_582_n702# cdac_vp a_674_n702# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.31 pd=2.62 as=0.165 ps=1.33 w=1 l=0.15
X58 VSS a_852_n296# RS_p VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.15
X59 VDD a_1716_n1348# a_482_n1818# VDD sky130_fd_pr__pfet_01v8 ad=0.139 pd=1.17 as=0.139 ps=1.17 w=0.84 l=0.15
X60 Q cdac_vn a_582_n702# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X61 ready a_564_n1721# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X62 a_482_n1818# a_476_n1721# a_564_n1721# VDD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.15
X63 VSS a_1950_n1721# comp_outn VSS sky130_fd_pr__nfet_01v8 ad=0.0759 pd=0.79 as=0.0759 ps=0.79 w=0.46 l=0.15
X64 a_476_n1721# a_852_n296# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0759 pd=0.79 as=0.0759 ps=0.79 w=0.46 l=0.15
X65 VDD a_1248_n288# a_1566_n378# VDD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X66 a_1566_n378# a_1248_n288# a_674_n702# VSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X67 a_582_n702# cdac_vp a_674_n702# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X68 VSS clk a_582_n702# VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X69 VDD RS_n RS_p VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.15
.ends

