magic
tech sky130A
magscale 1 2
timestamp 1697713470
<< nwell >>
rect -489 -128 490 124
<< pmos >>
rect -395 -88 395 88
<< pdiff >>
rect -453 76 -395 88
rect -453 -76 -441 76
rect -407 -76 -395 76
rect -453 -88 -395 -76
rect 395 76 453 88
rect 395 -76 407 76
rect 441 -76 453 76
rect 395 -88 453 -76
<< pdiffc >>
rect -441 -76 -407 76
rect 407 -76 441 76
<< poly >>
rect -395 169 395 185
rect -395 135 -379 169
rect 379 135 395 169
rect -395 88 395 135
rect -395 -135 395 -88
rect -395 -169 -379 -135
rect 379 -169 395 -135
rect -395 -185 395 -169
<< polycont >>
rect -379 135 379 169
rect -379 -169 379 -135
<< locali >>
rect -395 135 -379 169
rect 379 135 395 169
rect -441 76 -407 92
rect -441 -92 -407 -76
rect 407 76 441 92
rect 407 -92 441 -76
rect -395 -169 -379 -135
rect 379 -169 395 -135
<< viali >>
rect -379 135 379 169
rect -441 -76 -407 76
rect 407 -76 441 76
<< metal1 >>
rect -391 169 391 175
rect -391 135 -379 169
rect 379 135 391 169
rect -391 129 391 135
rect -447 76 -401 88
rect -447 -76 -441 76
rect -407 -76 -401 76
rect -447 -88 -401 -76
rect 401 76 447 88
rect 401 -76 407 76
rect 441 -76 447 76
rect 401 -88 447 -76
<< properties >>
string FIXED_BBOX -538 -254 538 254
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.875 l 3.95 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
