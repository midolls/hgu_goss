magic
tech sky130A
magscale 1 2
timestamp 1700415065
<< psubdiff >>
rect -87 5794 436 5840
rect 818 5794 1345 5840
rect 1983 5794 2878 5840
rect 4028 5794 5429 5840
rect 14738 5794 20301 5840
rect -109 5106 565 5152
rect 4598 5106 8013 5152
rect 10187 5106 15171 5152
rect 19393 5106 20225 5152
rect 20308 5106 20314 5152
<< poly >>
rect -249 5978 -179 6110
rect 656 5978 726 6110
rect 1437 6023 1891 6093
rect 2970 6023 3936 6093
rect 5521 6023 7511 6093
rect 10608 6023 14646 6093
rect 20393 6023 28527 6093
rect -271 5290 -201 5422
rect 657 5290 727 5422
rect 1921 5335 2375 5405
rect 3540 5335 4506 5405
rect 8105 5335 10095 5405
rect 15263 5335 19301 5405
rect 20317 5335 28451 5405
<< locali >>
rect -87 6374 436 6420
rect 818 6374 1345 6420
rect 1983 6374 2878 6420
rect 4028 6374 5429 6420
rect 7603 6374 10516 6420
rect 14738 6374 20301 6420
rect -87 5794 436 5840
rect 818 5794 1345 5840
rect 1983 5794 2878 5840
rect 4028 5794 5429 5840
rect 7603 5794 10516 5840
rect 14738 5794 20301 5840
rect -109 5686 565 5732
rect 947 5686 1829 5732
rect 2467 5686 3448 5732
rect 4598 5686 8013 5732
rect 10187 5686 15171 5732
rect 19393 5686 20264 5732
rect -109 5106 565 5152
rect 947 5106 1829 5152
rect 2467 5106 3448 5152
rect 4598 5106 8013 5152
rect 10187 5106 15171 5152
rect 19393 5106 20225 5152
rect 20308 5106 20314 5152
<< metal1 >>
rect 29502 6422 29566 6426
rect -95 6372 440 6422
rect 818 6372 1345 6422
rect 1983 6372 2878 6422
rect 4028 6372 5429 6422
rect 7603 6372 10516 6422
rect 14738 6372 20301 6422
rect 28616 6420 29566 6422
rect 28616 6372 29508 6420
rect 29502 6368 29508 6372
rect 29560 6368 29566 6420
rect 29502 6362 29566 6368
rect -87 6311 436 6343
rect 818 6311 1345 6343
rect 1983 6311 2878 6343
rect 4028 6311 5429 6343
rect 7603 6311 10516 6343
rect 14738 6311 20301 6343
rect 28619 6337 28783 6343
rect 28619 6311 28725 6337
rect 28719 6285 28725 6311
rect 28777 6285 28783 6337
rect 28719 6279 28783 6285
rect -95 6083 -31 6089
rect -95 6073 -89 6083
rect -133 6040 -89 6073
rect -95 6031 -89 6040
rect -37 6031 -31 6083
rect -95 6025 -31 6031
rect 357 6061 421 6067
rect 357 6009 363 6061
rect 415 6053 421 6061
rect 1268 6061 1332 6067
rect 415 6017 643 6053
rect 415 6009 421 6017
rect 357 6003 421 6009
rect 1268 6009 1274 6061
rect 1326 6050 1332 6061
rect 1326 6019 1553 6050
rect 2803 6049 2867 6055
rect 1326 6009 1332 6019
rect 1268 6003 1332 6009
rect 2803 5997 2809 6049
rect 2861 6038 2867 6049
rect 5353 6047 5417 6053
rect 2861 6009 3052 6038
rect 2861 5997 2867 6009
rect 2803 5991 2867 5997
rect 5353 5995 5359 6047
rect 5411 6036 5417 6047
rect 10326 6047 10390 6053
rect 5411 6007 5603 6036
rect 5411 5995 5417 6007
rect 5353 5989 5417 5995
rect 10326 5995 10332 6047
rect 10384 6036 10390 6047
rect 28631 6047 28695 6053
rect 28631 6036 28637 6047
rect 10384 6006 10690 6036
rect 28445 6007 28637 6036
rect 10384 5995 10390 6006
rect 10326 5989 10390 5995
rect 28631 5995 28637 6007
rect 28689 5995 28695 6047
rect 28631 5989 28695 5995
rect 28824 5843 28888 5849
rect 28824 5842 28830 5843
rect -87 5792 436 5842
rect 818 5792 1345 5842
rect 1983 5792 2878 5842
rect 4028 5792 5429 5842
rect 7603 5792 10516 5842
rect 14738 5792 20301 5842
rect 28619 5792 28830 5842
rect 28824 5791 28830 5792
rect 28882 5791 28888 5843
rect 28824 5785 28888 5791
rect 29504 5736 29568 5742
rect 29504 5734 29510 5736
rect -109 5684 565 5734
rect 947 5684 1829 5734
rect 2467 5684 3448 5734
rect 4598 5684 8013 5734
rect 10187 5684 15171 5734
rect 19393 5684 20264 5734
rect 28543 5684 29510 5734
rect 29562 5684 29568 5736
rect 29504 5678 29568 5684
rect -109 5623 565 5655
rect 947 5623 1829 5655
rect 2467 5623 3448 5655
rect 4598 5623 8013 5655
rect 10187 5623 15171 5655
rect 19393 5623 20264 5655
rect 28543 5649 28783 5655
rect 28543 5623 28725 5649
rect 28719 5597 28725 5623
rect 28777 5597 28783 5649
rect 28719 5591 28783 5597
rect 962 5401 1026 5407
rect 962 5394 968 5401
rect -95 5363 -31 5369
rect -95 5356 -89 5363
rect -173 5322 -89 5356
rect -95 5311 -89 5322
rect -37 5311 -31 5363
rect 773 5358 968 5394
rect 962 5349 968 5358
rect 1020 5349 1026 5401
rect 2480 5364 2544 5370
rect 2480 5354 2486 5364
rect 962 5343 1026 5349
rect 2293 5323 2486 5354
rect -95 5305 -31 5311
rect 2480 5312 2486 5323
rect 2538 5312 2544 5364
rect 4620 5359 4684 5365
rect 4620 5348 4626 5359
rect 4424 5319 4626 5348
rect 2480 5306 2544 5312
rect 4620 5307 4626 5319
rect 4678 5307 4684 5359
rect 10200 5362 10264 5368
rect 10200 5353 10206 5362
rect 10013 5324 10206 5353
rect 4620 5301 4684 5307
rect 10200 5310 10206 5324
rect 10258 5310 10264 5362
rect 19416 5358 19480 5364
rect 19416 5347 19422 5358
rect 19219 5318 19422 5347
rect 10200 5304 10264 5310
rect 19416 5306 19422 5318
rect 19474 5306 19480 5358
rect 19416 5300 19480 5306
rect 20149 5358 20213 5364
rect 20149 5306 20155 5358
rect 20207 5348 20213 5358
rect 20207 5319 20399 5348
rect 20207 5306 20213 5319
rect 20149 5300 20213 5306
rect 28825 5158 28889 5164
rect 28825 5154 28831 5158
rect -109 5104 565 5154
rect 947 5104 1829 5154
rect 2467 5104 3448 5154
rect 4598 5104 8013 5154
rect 10187 5104 15171 5154
rect 19393 5104 20225 5154
rect 28543 5106 28831 5154
rect 28883 5106 28889 5158
rect 28543 5104 28889 5106
rect 28825 5100 28889 5104
rect 150 4070 210 4078
rect 150 4018 154 4070
rect 206 4018 210 4070
rect 150 4007 210 4018
rect 162 3998 196 4007
rect 10327 3271 10391 3282
rect 10327 3219 10332 3271
rect 10384 3219 10391 3271
rect 10327 3208 10391 3219
rect 10341 3204 10375 3208
rect 28633 3177 28697 3183
rect 5352 3163 5418 3174
rect 1270 3143 1330 3149
rect 1270 3091 1274 3143
rect 1326 3091 1330 3143
rect 1270 3082 1330 3091
rect 2804 3131 2864 3137
rect 358 3074 418 3080
rect 358 3022 362 3074
rect 414 3022 418 3074
rect 1282 3071 1316 3082
rect 2804 3079 2808 3131
rect 2860 3079 2864 3131
rect 5352 3111 5358 3163
rect 5410 3111 5418 3163
rect 28633 3125 28639 3177
rect 28691 3125 28697 3177
rect 28633 3119 28697 3125
rect 28647 3114 28681 3119
rect 5352 3100 5418 3111
rect 5367 3096 5401 3100
rect 2804 3070 2864 3079
rect 2816 3059 2850 3070
rect 358 3013 418 3022
rect 370 3002 404 3013
rect -93 2598 -33 2604
rect -93 2546 -89 2598
rect -37 2546 -33 2598
rect -93 2540 -33 2546
rect -81 2526 -47 2540
rect 964 2459 1024 2465
rect 964 2407 968 2459
rect 1020 2407 1024 2459
rect 964 2398 1024 2407
rect 2482 2459 2542 2465
rect 2482 2407 2486 2459
rect 2538 2407 2542 2459
rect 2482 2398 2542 2407
rect 4620 2449 4684 2455
rect 976 2387 1010 2398
rect 2494 2387 2528 2398
rect 4620 2397 4626 2449
rect 4678 2397 4684 2449
rect 4620 2391 4684 2397
rect 10200 2451 10266 2462
rect 10200 2399 10206 2451
rect 10258 2399 10266 2451
rect 19417 2459 19481 2465
rect 19417 2407 19423 2459
rect 19475 2407 19481 2459
rect 19417 2401 19481 2407
rect 20149 2460 20213 2466
rect 20149 2408 20155 2460
rect 20207 2408 20213 2460
rect 20149 2402 20213 2408
rect 4634 2377 4668 2391
rect 10200 2388 10266 2399
rect 19431 2396 19465 2401
rect 20163 2397 20197 2402
rect 10215 2379 10249 2388
<< via1 >>
rect 29508 6368 29560 6420
rect 28725 6285 28777 6337
rect -89 6031 -37 6083
rect 363 6009 415 6061
rect 1274 6009 1326 6061
rect 2809 5997 2861 6049
rect 5359 5995 5411 6047
rect 10332 5995 10384 6047
rect 28637 5995 28689 6047
rect 28830 5791 28882 5843
rect 29510 5684 29562 5736
rect 28725 5597 28777 5649
rect -89 5311 -37 5363
rect 968 5349 1020 5401
rect 2486 5312 2538 5364
rect 4626 5307 4678 5359
rect 10206 5310 10258 5362
rect 19422 5306 19474 5358
rect 20155 5306 20207 5358
rect 28831 5106 28883 5158
rect 154 4018 206 4070
rect 10332 3219 10384 3271
rect 1274 3091 1326 3143
rect 362 3022 414 3074
rect 2808 3079 2860 3131
rect 5358 3111 5410 3163
rect 28639 3125 28691 3177
rect -89 2546 -37 2598
rect 968 2407 1020 2459
rect 2486 2407 2538 2459
rect 4626 2397 4678 2449
rect 10206 2399 10258 2451
rect 19423 2407 19475 2459
rect 20155 2408 20207 2460
<< metal2 >>
rect 29502 6420 29566 6426
rect 29502 6368 29508 6420
rect 29560 6368 29566 6420
rect 29502 6362 29566 6368
rect 28719 6337 28783 6343
rect 28719 6285 28725 6337
rect 28777 6285 28783 6337
rect 81 6248 196 6281
rect 28719 6279 28783 6285
rect -95 6083 -31 6089
rect -95 6031 -89 6083
rect -37 6073 -31 6083
rect 81 6073 114 6248
rect -37 6040 114 6073
rect -37 6031 -31 6040
rect -95 6025 -31 6031
rect -95 5363 -31 5369
rect -95 5311 -89 5363
rect -37 5311 -31 5363
rect -95 5305 -31 5311
rect -80 2609 -47 5305
rect 163 4081 196 6248
rect 357 6061 421 6067
rect 357 6009 363 6061
rect 415 6009 421 6061
rect 357 6003 421 6009
rect 1268 6061 1332 6067
rect 1268 6009 1274 6061
rect 1326 6009 1332 6061
rect 28734 6059 28768 6279
rect 29518 6078 29552 6362
rect 28734 6058 28928 6059
rect 1268 6003 1332 6009
rect 2803 6049 2867 6055
rect 150 4072 210 4081
rect 150 4016 152 4072
rect 208 4016 210 4072
rect 150 4007 210 4016
rect 371 3085 405 6003
rect 962 5401 1026 5407
rect 962 5349 968 5401
rect 1020 5349 1026 5401
rect 962 5343 1026 5349
rect 358 3076 418 3085
rect 358 3020 360 3076
rect 416 3020 418 3076
rect 358 3011 418 3020
rect -93 2600 -33 2609
rect -93 2544 -91 2600
rect -35 2544 -33 2600
rect -93 2535 -33 2544
rect 977 2470 1011 5343
rect 1283 3154 1317 6003
rect 2803 5997 2809 6049
rect 2861 5997 2867 6049
rect 2803 5991 2867 5997
rect 5353 6047 5417 6053
rect 5353 5995 5359 6047
rect 5411 5995 5417 6047
rect 2480 5364 2544 5370
rect 2480 5312 2486 5364
rect 2538 5312 2544 5364
rect 2480 5306 2544 5312
rect 1270 3145 1330 3154
rect 1270 3089 1272 3145
rect 1328 3089 1330 3145
rect 1270 3080 1330 3089
rect 2495 2470 2529 5306
rect 2817 3142 2850 5991
rect 5353 5989 5417 5995
rect 10326 6047 10390 6053
rect 10326 5995 10332 6047
rect 10384 5995 10390 6047
rect 10326 5989 10390 5995
rect 28631 6047 28695 6053
rect 28631 5995 28637 6047
rect 28689 5995 28695 6047
rect 28631 5989 28695 5995
rect 4620 5359 4684 5365
rect 4620 5307 4626 5359
rect 4678 5307 4684 5359
rect 4620 5301 4684 5307
rect 2804 3133 2864 3142
rect 2804 3077 2806 3133
rect 2862 3077 2864 3133
rect 2804 3068 2864 3077
rect 964 2461 1024 2470
rect 964 2405 966 2461
rect 1022 2405 1024 2461
rect 964 2396 1024 2405
rect 2482 2461 2542 2470
rect 2482 2405 2484 2461
rect 2540 2405 2542 2461
rect 4635 2460 4669 5301
rect 5367 3174 5401 5989
rect 10200 5362 10264 5368
rect 10200 5310 10206 5362
rect 10258 5310 10264 5362
rect 10200 5304 10264 5310
rect 5352 3165 5418 3174
rect 5352 3109 5357 3165
rect 5413 3109 5418 3165
rect 5352 3100 5418 3109
rect 10215 2462 10249 5304
rect 10341 3282 10375 5989
rect 19416 5358 19480 5364
rect 19416 5306 19422 5358
rect 19474 5306 19480 5358
rect 19416 5300 19480 5306
rect 20149 5358 20213 5364
rect 20149 5306 20155 5358
rect 20207 5306 20213 5358
rect 20149 5300 20213 5306
rect 10327 3273 10391 3282
rect 10327 3217 10331 3273
rect 10387 3217 10391 3273
rect 10327 3208 10391 3217
rect 19431 2470 19465 5300
rect 20163 2471 20197 5300
rect 28647 3188 28681 5989
rect 28734 5981 28941 6058
rect 28734 5655 28768 5981
rect 29518 5978 29744 6078
rect 28824 5843 28888 5849
rect 28824 5791 28830 5843
rect 28882 5791 28888 5843
rect 28824 5785 28888 5791
rect 28719 5649 28783 5655
rect 28719 5597 28725 5649
rect 28777 5597 28783 5649
rect 28719 5591 28783 5597
rect 28839 5429 28873 5785
rect 29518 5742 29552 5978
rect 29504 5736 29568 5742
rect 29504 5684 29510 5736
rect 29562 5684 29568 5736
rect 29504 5678 29568 5684
rect 28839 5352 29152 5429
rect 28839 5164 28873 5352
rect 28825 5158 28889 5164
rect 28825 5106 28831 5158
rect 28883 5106 28889 5158
rect 28825 5100 28889 5106
rect 28633 3179 28697 3188
rect 28633 3123 28637 3179
rect 28693 3123 28697 3179
rect 28633 3114 28697 3123
rect 2482 2396 2542 2405
rect 4620 2451 4684 2460
rect 4620 2395 4624 2451
rect 4680 2395 4684 2451
rect 4620 2386 4684 2395
rect 10200 2453 10266 2462
rect 10200 2397 10205 2453
rect 10261 2397 10266 2453
rect 10200 2388 10266 2397
rect 19417 2461 19481 2470
rect 19417 2405 19421 2461
rect 19477 2405 19481 2461
rect 19417 2396 19481 2405
rect 20149 2462 20213 2471
rect 20149 2406 20153 2462
rect 20209 2406 20213 2462
rect 20149 2397 20213 2406
<< via2 >>
rect 152 4070 208 4072
rect 152 4018 154 4070
rect 154 4018 206 4070
rect 206 4018 208 4070
rect 152 4016 208 4018
rect 360 3074 416 3076
rect 360 3022 362 3074
rect 362 3022 414 3074
rect 414 3022 416 3074
rect 360 3020 416 3022
rect -91 2598 -35 2600
rect -91 2546 -89 2598
rect -89 2546 -37 2598
rect -37 2546 -35 2598
rect -91 2544 -35 2546
rect 1272 3143 1328 3145
rect 1272 3091 1274 3143
rect 1274 3091 1326 3143
rect 1326 3091 1328 3143
rect 1272 3089 1328 3091
rect 2806 3131 2862 3133
rect 2806 3079 2808 3131
rect 2808 3079 2860 3131
rect 2860 3079 2862 3131
rect 2806 3077 2862 3079
rect 966 2459 1022 2461
rect 966 2407 968 2459
rect 968 2407 1020 2459
rect 1020 2407 1022 2459
rect 966 2405 1022 2407
rect 2484 2459 2540 2461
rect 2484 2407 2486 2459
rect 2486 2407 2538 2459
rect 2538 2407 2540 2459
rect 2484 2405 2540 2407
rect 5357 3163 5413 3165
rect 5357 3111 5358 3163
rect 5358 3111 5410 3163
rect 5410 3111 5413 3163
rect 5357 3109 5413 3111
rect 10331 3271 10387 3273
rect 10331 3219 10332 3271
rect 10332 3219 10384 3271
rect 10384 3219 10387 3271
rect 10331 3217 10387 3219
rect 28637 3177 28693 3179
rect 28637 3125 28639 3177
rect 28639 3125 28691 3177
rect 28691 3125 28693 3177
rect 28637 3123 28693 3125
rect 4624 2449 4680 2451
rect 4624 2397 4626 2449
rect 4626 2397 4678 2449
rect 4678 2397 4680 2449
rect 4624 2395 4680 2397
rect 10205 2451 10261 2453
rect 10205 2399 10206 2451
rect 10206 2399 10258 2451
rect 10258 2399 10261 2451
rect 10205 2397 10261 2399
rect 19421 2459 19477 2461
rect 19421 2407 19423 2459
rect 19423 2407 19475 2459
rect 19475 2407 19477 2459
rect 19421 2405 19477 2407
rect 20153 2460 20209 2462
rect 20153 2408 20155 2460
rect 20155 2408 20207 2460
rect 20207 2408 20209 2460
rect 20153 2406 20209 2408
<< metal3 >>
rect 150 4072 210 4087
rect 150 4016 152 4072
rect 208 4016 210 4072
rect 150 4007 210 4016
rect 10327 3203 10391 3213
rect 5352 3165 5367 3186
rect 5401 3165 5418 3186
rect 1267 3145 1333 3154
rect 358 3089 418 3091
rect 1267 3089 1272 3145
rect 1328 3089 1333 3145
rect 355 3076 421 3089
rect 1267 3079 1333 3089
rect 2804 3133 2864 3137
rect 355 3020 360 3076
rect 416 3020 421 3076
rect 1268 3074 1332 3079
rect 2804 3077 2806 3133
rect 2862 3077 2864 3133
rect 5352 3109 5357 3165
rect 5413 3109 5418 3165
rect 5352 3096 5418 3109
rect 28632 3183 28633 3192
rect 28697 3183 28698 3192
rect 28632 3179 28698 3183
rect 28632 3157 28637 3179
rect 28632 3156 28636 3157
rect 28632 3123 28637 3156
rect 28693 3158 28698 3179
rect 28694 3157 28698 3158
rect 28693 3123 28698 3157
rect 28632 3122 28642 3123
rect 28643 3122 28698 3123
rect 28632 3102 28698 3122
rect 2804 3071 2864 3077
rect 2866 3059 2867 3060
rect 1267 3040 1268 3042
rect 1332 3040 1333 3042
rect 355 3000 421 3020
rect 10205 2984 10261 2987
rect -93 2605 -33 2615
rect 2442 2538 2545 2548
rect 964 2465 1024 2476
rect 2482 2474 2542 2476
rect 2479 2465 2545 2474
rect 2479 2401 2480 2465
rect 2544 2401 2545 2465
rect 964 2396 1024 2401
rect 2479 2384 2545 2401
rect 4620 2456 4685 2472
rect 19416 2465 19482 2470
rect 4620 2392 4621 2456
rect 10200 2453 10266 2462
rect 10200 2397 10205 2453
rect 10261 2397 10266 2453
rect 4620 2377 4685 2392
rect 10200 2388 10266 2397
rect 19416 2401 19417 2465
rect 19481 2401 19482 2465
rect 19416 2384 19482 2401
<< via3 >>
rect 962 2461 1026 2465
rect 962 2405 966 2461
rect 966 2405 1022 2461
rect 1022 2405 1026 2461
rect 962 2401 1026 2405
rect 2480 2461 2544 2465
rect 2480 2405 2484 2461
rect 2484 2405 2540 2461
rect 2540 2405 2544 2461
rect 2480 2401 2544 2405
<< metal4 >>
rect 29171 6320 29404 6321
rect 28942 5756 29404 6320
rect 29749 5770 30141 6341
rect 29171 5755 29404 5756
rect 29146 5204 29501 5596
rect -209 4434 -158 4641
rect 150 3994 210 4087
rect -324 3245 -280 3393
rect 10327 3203 10391 3282
rect 5352 3163 5367 3186
rect 5401 3163 5418 3186
rect 355 3000 421 3089
rect 1267 3071 1333 3154
rect 5352 3096 5418 3163
rect 1267 3040 1268 3042
rect 1332 3040 1333 3042
rect 8383 2928 8447 2992
rect -93 2605 -33 2615
rect -93 2526 -33 2541
rect 964 2465 1024 2474
rect 2479 2465 2545 2474
rect 2479 2401 2480 2465
rect 2544 2401 2545 2465
rect 964 2384 1024 2401
rect 2479 2384 2545 2401
rect 4620 2456 4685 2472
rect 19417 2465 19481 2469
rect 4620 2392 4621 2456
rect 4620 2377 4685 2392
rect 10200 2388 10266 2462
rect 20148 2385 20214 2475
rect -205 2058 -161 2188
rect -329 832 -283 967
<< metal5 >>
rect 287 5026 524 5262
rect 1717 5026 1954 5262
rect 3301 5026 3538 5262
rect 5394 5026 5631 5262
rect 10368 5026 10605 5262
rect 39298 5026 39534 5262
rect 287 50 524 286
rect 1717 50 1954 286
rect 3301 50 3538 286
rect 5394 50 5631 286
rect 10368 50 10605 286
rect 39298 50 39534 286
use hgu_cdac_8bit_array  hgu_cdac_8bit_array_2
timestamp 1699890160
transform 1 0 4202 0 -1 -4800
box -4661 -7612 35404 -4800
use hgu_cdac_8bit_array  hgu_cdac_8bit_array_3
timestamp 1699890160
transform 1 0 4202 0 -1 -2312
box -4661 -7612 35404 -4800
use hgu_cdac_unit  hgu_cdac_unit_0
timestamp 1699890160
transform 1 0 -1145 0 -1 2044
box 686 598 1358 1826
use hgu_cdac_unit  hgu_cdac_unit_1
timestamp 1699890160
transform 1 0 -1145 0 -1 4532
box 686 598 1358 1826
use hgu_inverter  hgu_inverter_0
timestamp 1699345134
transform 1 0 -747 0 1 4944
box 347 160 675 824
use hgu_inverter  hgu_inverter_1
timestamp 1699345134
transform 1 0 -725 0 1 5632
box 347 160 675 824
use inv_2_test  inv_2_test_0
timestamp 1699782319
transform 1 0 128 0 1 2744
box 400 2360 856 3024
use inv_2_test  inv_2_test_1
timestamp 1699782319
transform 1 0 -1 0 1 3432
box 400 2360 856 3024
use inv_4_test  inv_4_test_1
timestamp 1699782319
transform 1 0 2239 0 1 3780
box -447 1324 265 1988
use inv_4_test  inv_4_test_2
timestamp 1699782319
transform 1 0 1755 0 1 4468
box -447 1324 265 1988
use inv_8_test  inv_8_test_0
timestamp 1699782319
transform 1 0 3315 0 1 2784
box 96 2320 1320 2984
use inv_8_test  inv_8_test_1
timestamp 1699782319
transform 1 0 2745 0 1 3472
box 96 2320 1320 2984
use inv_16_test  inv_16_test_0
timestamp 1699782319
transform 1 0 8625 0 1 5144
box -649 -40 1599 624
use inv_16_test  inv_16_test_1
timestamp 1699782319
transform 1 0 6041 0 1 5832
box -649 -40 1599 624
use inv_32_test  inv_32_test_0
timestamp 1699782319
transform 1 0 12782 0 1 8194
box -2303 -2402 1993 -1738
use inv_32_test  inv_32_test_1
timestamp 1699782319
transform 1 0 17437 0 1 7506
box -2303 -2402 1993 -1738
use inv_64_test  inv_64_test_0
timestamp 1699782319
transform 1 0 23771 0 1 7506
box -3583 -2402 4809 -1738
use inv_64_test  inv_64_test_1
timestamp 1699782319
transform 1 0 23847 0 1 8194
box -3583 -2402 4809 -1738
<< labels >>
flabel metal4 -209 4434 -158 4641 0 FreeSans 480 0 0 0 t<0>
port 27 nsew
flabel metal4 -205 2058 -161 2188 0 FreeSans 320 0 0 0 tb<0>
port 76 nsew
flabel metal4 -324 3245 -280 3393 0 FreeSans 320 0 0 0 tu
port 90 nsew
flabel poly 2970 6023 3936 6093 0 FreeSans 320 0 0 0 d<3>
port 102 nsew
flabel poly 1437 6023 1891 6093 0 FreeSans 320 0 0 0 d<2>
port 104 nsew
flabel poly 656 5978 726 6110 0 FreeSans 320 0 0 0 d<1>
port 106 nsew
flabel poly -249 5978 -179 6110 0 FreeSans 320 0 0 0 d<0>
port 109 nsew
flabel poly 5521 6023 7511 6093 0 FreeSans 320 0 0 0 d<4>
port 111 nsew
flabel poly 10608 6023 14646 6093 0 FreeSans 320 0 0 0 d<5>
port 113 nsew
flabel poly 20393 6023 28527 6093 0 FreeSans 320 0 0 0 d<6>
port 115 nsew
flabel poly -271 5290 -201 5422 0 FreeSans 320 0 0 0 db<0>
port 117 nsew
flabel poly 657 5290 727 5422 0 FreeSans 320 0 0 0 db<1>
port 119 nsew
flabel poly 1921 5335 2375 5405 0 FreeSans 320 0 0 0 db<2>
port 121 nsew
flabel poly 3540 5335 4506 5405 0 FreeSans 320 0 0 0 db<3>
port 123 nsew
flabel poly 8105 5335 10095 5405 0 FreeSans 320 0 0 0 db<4>
port 125 nsew
flabel poly 15263 5335 19301 5405 0 FreeSans 320 0 0 0 db<5>
port 127 nsew
flabel metal4 -329 832 -283 967 0 FreeSans 320 0 0 0 tub
port 131 nsew
flabel poly 20317 5335 28451 5405 0 FreeSans 320 0 0 0 db<6>
port 133 nsew
flabel metal5 287 5026 524 5262 0 FreeSans 320 0 0 0 t<1>
port 135 nsew
flabel metal5 1717 5026 1954 5262 0 FreeSans 320 0 0 0 t<2>
port 137 nsew
flabel metal5 3301 5026 3538 5262 0 FreeSans 320 0 0 0 t<3>
port 139 nsew
flabel metal5 5394 5026 5631 5262 0 FreeSans 320 0 0 0 t<4>
port 141 nsew
flabel metal5 10368 5026 10605 5262 0 FreeSans 480 0 0 0 t<5>
port 143 nsew
flabel metal5 39298 5026 39534 5262 0 FreeSans 480 0 0 0 t<6>
port 145 nsew
flabel metal5 287 50 524 286 0 FreeSans 480 0 0 0 tb<1>
port 147 nsew
flabel metal5 1717 50 1954 286 0 FreeSans 480 0 0 0 tb<2>
port 149 nsew
flabel metal5 3301 50 3538 286 0 FreeSans 480 0 0 0 tb<3>
port 151 nsew
flabel metal5 5394 50 5631 286 0 FreeSans 480 0 0 0 tb<4>
port 153 nsew
flabel metal5 10368 50 10605 286 0 FreeSans 480 0 0 0 tb<5>
port 155 nsew
flabel metal5 39298 50 39534 286 0 FreeSans 480 0 0 0 tb<6>
port 157 nsew
<< end >>
