* NGSPICE file created from hgu_sarlogic_sw_ctrl.ext - technology: sky130A

.subckt sky130_fd_sc_hd__buf_1 A VGND VPWR X VNB VPB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_4 A VGND VPWR X VNB VPB
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_16 A VGND VPWR X VNB VPB
X0 VGND A a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 a_109_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 VPWR A a_109_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 a_109_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X17 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X18 VPWR A a_109_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 VGND A a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X21 VGND A a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X22 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X23 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X24 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X25 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X26 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X27 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X28 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X29 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X30 a_109_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X31 a_109_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X32 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X33 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X34 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X35 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X36 VPWR A a_109_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X37 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X38 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X39 a_109_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X40 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X41 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X42 a_109_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X43 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfbbn_1 CLK_N D RESET_B SET_B VGND VPWR Q Q_N VNB VPB
X0 a_791_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0974 pd=0.97 as=0.0882 ps=0.84 w=0.42 l=0.15
X1 a_1555_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.03 as=0.0703 ps=0.755 w=0.42 l=0.15
X2 VPWR RESET_B a_941_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.17 ps=1.81 w=0.64 l=0.15
X3 a_1415_315# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.132 pd=1.22 as=0.0956 ps=0.875 w=0.42 l=0.15
X4 a_791_47# a_941_21# a_647_21# VNB sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5 VGND a_1415_315# a_1363_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.066 ps=0.745 w=0.42 l=0.15
X6 a_1340_413# a_27_47# a_1256_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0787 pd=0.795 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 VPWR CLK_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X8 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X9 a_473_413# a_193_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0675 pd=0.735 as=0.066 ps=0.745 w=0.36 l=0.15
X10 a_1555_47# a_941_21# a_1415_315# VNB sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X11 VPWR a_1415_315# a_2136_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X12 a_1256_413# a_193_47# a_1112_329# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X13 a_581_47# a_27_47# a_473_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0675 ps=0.735 w=0.36 l=0.15
X14 a_647_21# a_473_413# a_791_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.0974 ps=0.97 w=0.64 l=0.15
X15 a_647_21# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X16 VPWR a_941_21# a_891_329# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X17 a_557_413# a_193_47# a_473_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X18 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X19 Q a_2136_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X20 a_473_413# a_27_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0651 ps=0.73 w=0.42 l=0.15
X21 a_891_329# a_473_413# a_647_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X22 Q_N a_1415_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X23 VGND RESET_B a_941_21# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X24 Q a_2136_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X25 VPWR a_647_21# a_557_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X26 a_1112_329# a_647_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X27 VGND a_647_21# a_581_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0671 ps=0.75 w=0.42 l=0.15
X28 VGND a_1415_315# a_2136_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X29 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X30 VPWR a_941_21# a_1672_329# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X31 VPWR a_1415_315# a_1340_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0956 pd=0.875 as=0.0787 ps=0.795 w=0.42 l=0.15
X32 a_1363_47# a_193_47# a_1256_413# VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0486 ps=0.63 w=0.36 l=0.15
X33 Q_N a_1415_315# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X34 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X35 a_1159_47# a_647_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.116 pd=1.09 as=0.166 ps=1.8 w=0.64 l=0.15
X36 a_1672_329# a_1256_413# a_1415_315# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.132 ps=1.22 w=0.84 l=0.15
X37 VGND CLK_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X38 a_1256_413# a_27_47# a_1159_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0486 pd=0.63 as=0.116 ps=1.09 w=0.36 l=0.15
X39 a_1415_315# a_1256_413# a_1555_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.109 ps=1.03 w=0.64 l=0.15
.ends

.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VPWR X VNB VPB
X0 VPWR a_505_21# a_535_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1 a_505_21# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_218_374# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X3 VGND a_505_21# a_439_47# VNB sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_76_199# A0 a_218_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X5 a_505_21# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X6 a_439_47# A0 a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X7 a_535_374# A1 a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X8 a_76_199# A1 a_218_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X9 a_218_47# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X10 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt hgu_sarlogic_sw_ctrl VSS_SW[1] VSS_SW[2] VSS_SW[3] VSS_SW[4] VSS_SW[5] VSS_SW[6]
+ VSS_SW[7] VDD_SW[2] VDD_SW[3] VDD_SW[4] VDD_SW[5] VDD_SW[6] VDD_SW[7] D[2] D[3]
+ D[4] D[5] D[6] D[7] check[0] check[1] check[2] check[3] check[4] check[5] check[6]
+ VDD_SW_b[1] VDD_SW_b[2] VDD_SW_b[3] VDD_SW_b[4] VDD_SW_b[5] VDD_SW_b[6] VDD_SW_b[7]
+ VSS_SW_b[1] VSS_SW_b[2] VSS_SW_b[3] VSS_SW_b[4] VSS_SW_b[5] VSS_SW_b[6] VSS_SW_b[7]
+ D[1] VDD_SW[1] ready reset VDD VSS
Xx1 reset VSS VDD x3/A VSS VDD sky130_fd_sc_hd__buf_1
Xx3 x3/A VSS VDD x3/X VSS VDD sky130_fd_sc_hd__buf_4
Xx2 x3/X VSS VDD x2/X VSS VDD sky130_fd_sc_hd__buf_16
Xx5 x7/X D[7] x2/X VDD VSS VDD VSS_SW[7] VSS_SW_b[7] VSS VDD sky130_fd_sc_hd__dfbbn_1
Xx6 VSS x9/A1 check[6] VSS VDD x6/X VSS VDD sky130_fd_sc_hd__mux2_1
Xx7 VSS x9/A1 check[6] VSS VDD x7/X VSS VDD sky130_fd_sc_hd__mux2_1
Xx8 VSS x9/A1 check[5] VSS VDD x8/X VSS VDD sky130_fd_sc_hd__mux2_1
Xx9 VSS x9/A1 check[5] VSS VDD x9/X VSS VDD sky130_fd_sc_hd__mux2_1
Xx30 x30/A VSS VDD x9/A1 VSS VDD sky130_fd_sc_hd__buf_16
Xx20 VSS x9/A1 check[0] VSS VDD x20/X VSS VDD sky130_fd_sc_hd__mux2_1
Xx31 x16/X D[2] VDD x2/X VSS VDD VDD_SW[2] VDD_SW_b[2] VSS VDD sky130_fd_sc_hd__dfbbn_1
Xx10 VSS x9/A1 check[4] VSS VDD x10/X VSS VDD sky130_fd_sc_hd__mux2_1
Xx32 x17/X D[2] x2/X VDD VSS VDD VSS_SW[2] VSS_SW_b[2] VSS VDD sky130_fd_sc_hd__dfbbn_1
Xx21 x9/X D[6] x2/X VDD VSS VDD VSS_SW[6] VSS_SW_b[6] VSS VDD sky130_fd_sc_hd__dfbbn_1
Xx22 ready VSS VDD x27/A VSS VDD sky130_fd_sc_hd__buf_1
Xx11 VSS x9/A1 check[4] VSS VDD x11/X VSS VDD sky130_fd_sc_hd__mux2_1
Xx12 VSS x9/A1 check[3] VSS VDD x12/X VSS VDD sky130_fd_sc_hd__mux2_1
Xx34 x18/X D[1] VDD x2/X VSS VDD VDD_SW[1] VDD_SW_b[1] VSS VDD sky130_fd_sc_hd__dfbbn_1
Xx23 x10/X D[5] VDD x2/X VSS VDD VDD_SW[5] VDD_SW_b[5] VSS VDD sky130_fd_sc_hd__dfbbn_1
Xx13 VSS x9/A1 check[3] VSS VDD x13/X VSS VDD sky130_fd_sc_hd__mux2_1
Xx35 x20/X D[1] x2/X VDD VSS VDD VSS_SW[1] VSS_SW_b[1] VSS VDD sky130_fd_sc_hd__dfbbn_1
Xx24 x11/X D[5] x2/X VDD VSS VDD VSS_SW[5] VSS_SW_b[5] VSS VDD sky130_fd_sc_hd__dfbbn_1
Xx15 VSS x9/A1 check[2] VSS VDD x15/X VSS VDD sky130_fd_sc_hd__mux2_1
Xx14 VSS x9/A1 check[2] VSS VDD x14/X VSS VDD sky130_fd_sc_hd__mux2_1
Xx26 x13/X D[4] x2/X VDD VSS VDD VSS_SW[4] VSS_SW_b[4] VSS VDD sky130_fd_sc_hd__dfbbn_1
Xx25 x12/X D[4] VDD x2/X VSS VDD VDD_SW[4] VDD_SW_b[4] VSS VDD sky130_fd_sc_hd__dfbbn_1
Xx27 x27/A VSS VDD x30/A VSS VDD sky130_fd_sc_hd__buf_4
Xx16 VSS x9/A1 check[1] VSS VDD x16/X VSS VDD sky130_fd_sc_hd__mux2_1
Xx17 VSS x9/A1 check[1] VSS VDD x17/X VSS VDD sky130_fd_sc_hd__mux2_1
Xx28 x14/X D[3] VDD x2/X VSS VDD VDD_SW[3] VDD_SW_b[3] VSS VDD sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__dfbbn_1_0 x6/X D[7] VDD x2/X VSS VDD VDD_SW[7] VDD_SW_b[7] VSS VDD
+ sky130_fd_sc_hd__dfbbn_1
Xx18 VSS x9/A1 check[0] VSS VDD x18/X VSS VDD sky130_fd_sc_hd__mux2_1
Xx29 x15/X D[3] x2/X VDD VSS VDD VSS_SW[3] VSS_SW_b[3] VSS VDD sky130_fd_sc_hd__dfbbn_1
Xx19 x8/X D[6] VDD x2/X VSS VDD VDD_SW[6] VDD_SW_b[6] VSS VDD sky130_fd_sc_hd__dfbbn_1
.ends

