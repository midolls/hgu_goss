magic
tech sky130A
magscale 1 2
timestamp 1699599968
<< checkpaint >>
rect -949 -4662 2097 -1638
<< error_s >>
rect 2102 977 2533 1041
rect 2149 973 2213 977
rect 2104 944 2213 973
rect 2229 944 2293 977
rect 2309 973 2373 977
rect 2389 973 2453 977
rect 2309 944 2453 973
rect 2469 944 2533 977
rect 2104 942 2171 944
rect 318 375 353 409
rect 319 356 353 375
rect 705 356 758 357
rect 149 307 207 313
rect 149 273 161 307
rect 149 267 207 273
rect 338 -23 353 356
rect 372 322 407 356
rect 687 322 758 356
rect 372 -23 406 322
rect 688 321 758 322
rect 705 287 776 321
rect 1056 287 1091 321
rect 518 254 576 260
rect 518 220 530 254
rect 518 214 576 220
rect 518 60 576 66
rect 518 26 530 60
rect 518 20 576 26
rect 372 -57 387 -23
rect 705 -76 775 287
rect 1057 268 1091 287
rect 887 219 945 225
rect 887 185 899 219
rect 887 179 945 185
rect 887 7 945 13
rect 887 -27 899 7
rect 887 -33 945 -27
rect 705 -112 758 -76
rect 1076 -129 1091 268
rect 1110 234 1145 268
rect 1110 -129 1144 234
rect 1678 181 1736 187
rect 1256 166 1314 172
rect 1256 132 1268 166
rect 1678 147 1690 181
rect 1678 141 1736 147
rect 1256 126 1314 132
rect 1678 -13 1736 -7
rect 1256 -46 1314 -40
rect 1256 -80 1268 -46
rect 1678 -47 1690 -13
rect 1678 -53 1736 -47
rect 2104 -57 2111 942
rect 1256 -86 1314 -80
rect 2045 -86 2111 -57
rect 2164 -117 2171 942
rect 1985 -119 2171 -117
rect 2224 942 2291 944
rect 2224 -117 2231 942
rect 2284 -117 2291 942
rect 2224 -119 2291 -117
rect 2344 942 2411 944
rect 2344 -117 2351 942
rect 2404 -117 2411 942
rect 2464 -113 2471 942
rect 2524 -53 2531 942
rect 2531 -90 2591 -57
rect 2344 -119 2411 -117
rect 2464 -119 2590 -117
rect 1110 -163 1125 -129
rect 1985 -146 2590 -119
rect 2102 -150 2590 -146
rect 2102 -183 2533 -150
rect 2149 -216 2213 -183
rect 2229 -216 2293 -183
rect 2309 -216 2373 -183
rect 2389 -216 2453 -183
rect 2469 -216 2533 -183
rect 573 -1974 877 -1941
rect 893 -1974 957 -1941
rect 573 -1989 1004 -1974
rect 1020 -1989 1084 -1974
rect 573 -2005 1318 -1989
rect 1794 -2005 2225 -1941
rect 3015 -2005 3446 -1941
rect 4236 -2005 4667 -1941
rect 5457 -2005 5888 -1941
rect 6678 -2005 7109 -1941
rect 620 -2009 684 -2005
rect 575 -2038 684 -2009
rect 700 -2038 764 -2005
rect 780 -2038 1318 -2005
rect 1841 -2009 1905 -2005
rect 575 -2040 642 -2038
rect -4 -2653 30 -2649
rect 88 -2653 122 -2649
rect 180 -2653 214 -2649
rect -33 -2663 35 -2653
rect 77 -2663 239 -2653
rect -33 -2687 281 -2663
rect -67 -2699 281 -2687
rect -67 -2707 319 -2699
rect -42 -2711 319 -2707
rect -33 -2733 319 -2711
rect -33 -2827 281 -2733
rect 317 -2767 319 -2747
rect 319 -2827 353 -2795
rect -33 -3145 364 -2827
rect 463 -2849 521 -2843
rect 463 -2883 475 -2849
rect 463 -2889 521 -2883
rect 463 -3039 521 -3037
rect 575 -3039 582 -2040
rect 463 -3043 582 -3039
rect 463 -3077 475 -3043
rect 516 -3068 582 -3043
rect 463 -3083 521 -3077
rect 635 -3099 642 -2040
rect 456 -3101 642 -3099
rect 643 -3099 702 -2040
rect 703 -3083 762 -2040
rect 807 -2053 871 -2038
rect 887 -2053 1318 -2038
rect 815 -2055 882 -2053
rect 755 -3099 762 -3083
rect 643 -3101 762 -3099
rect 769 -3099 822 -2055
rect 829 -3099 882 -2055
rect 934 -2057 1002 -2053
rect 769 -3101 882 -3099
rect 889 -2088 1002 -2057
rect 1014 -2057 1158 -2053
rect 1174 -2057 1238 -2053
rect 1014 -2086 1238 -2057
rect 1254 -2086 1318 -2053
rect 1796 -2038 1905 -2009
rect 1921 -2038 1985 -2005
rect 2001 -2009 2065 -2005
rect 2081 -2009 2145 -2005
rect 2001 -2038 2145 -2009
rect 2161 -2038 2225 -2005
rect 3062 -2009 3126 -2005
rect 3017 -2038 3126 -2009
rect 3142 -2038 3206 -2005
rect 3222 -2009 3286 -2005
rect 3302 -2009 3366 -2005
rect 3222 -2038 3366 -2009
rect 3382 -2038 3446 -2005
rect 4283 -2009 4347 -2005
rect 4238 -2038 4347 -2009
rect 4363 -2038 4427 -2005
rect 4443 -2009 4507 -2005
rect 4523 -2009 4587 -2005
rect 4443 -2038 4587 -2009
rect 4603 -2038 4667 -2005
rect 5504 -2009 5568 -2005
rect 5459 -2038 5568 -2009
rect 5584 -2038 5648 -2005
rect 5664 -2009 5728 -2005
rect 5744 -2009 5808 -2005
rect 5664 -2038 5808 -2009
rect 5824 -2038 5888 -2005
rect 6725 -2009 6789 -2005
rect 6680 -2038 6789 -2009
rect 6805 -2038 6869 -2005
rect 6885 -2009 6949 -2005
rect 6965 -2009 7029 -2005
rect 6885 -2038 7029 -2009
rect 7045 -2038 7109 -2005
rect 1796 -2040 1863 -2038
rect 889 -3099 942 -2088
rect 949 -3099 1002 -2088
rect 456 -3128 877 -3101
rect 573 -3134 877 -3128
rect 889 -3132 1002 -3099
rect 1009 -2088 1122 -2086
rect 1009 -3132 1062 -2088
rect 1069 -3132 1122 -2088
rect 1129 -2088 1196 -2086
rect 1129 -3068 1188 -2088
rect 1129 -3132 1136 -3068
rect 889 -3134 957 -3132
rect 1009 -3134 1076 -3132
rect -33 -3165 387 -3145
rect 573 -3149 1004 -3134
rect 1020 -3149 1084 -3134
rect 1129 -3147 1188 -3132
rect 1189 -3147 1248 -2088
rect 1249 -3143 1256 -2088
rect 1309 -3083 1316 -2088
rect 1370 -2801 1428 -2795
rect 1370 -2835 1382 -2801
rect 1370 -2841 1428 -2835
rect 1370 -2995 1428 -2989
rect 1370 -3029 1382 -2995
rect 1370 -3035 1428 -3029
rect 1796 -3039 1803 -2040
rect 1737 -3068 1803 -3039
rect 1316 -3120 1376 -3087
rect 1856 -3099 1863 -2040
rect 1677 -3101 1863 -3099
rect 1916 -2040 1983 -2038
rect 1916 -3099 1923 -2040
rect 1976 -3099 1983 -2040
rect 1916 -3101 1983 -3099
rect 2036 -2040 2103 -2038
rect 3017 -2040 3084 -2038
rect 2036 -3099 2043 -2040
rect 2096 -3099 2103 -2040
rect 2156 -3095 2163 -2040
rect 2216 -3035 2223 -2040
rect 2591 -2801 2649 -2795
rect 2591 -2835 2603 -2801
rect 2591 -2841 2649 -2835
rect 2591 -2995 2649 -2989
rect 2591 -3029 2603 -2995
rect 2591 -3035 2649 -3029
rect 3017 -3039 3024 -2040
rect 2223 -3072 2283 -3039
rect 2958 -3068 3024 -3039
rect 3077 -3099 3084 -2040
rect 2036 -3101 2103 -3099
rect 2156 -3101 2282 -3099
rect 1677 -3128 2282 -3101
rect 2898 -3101 3084 -3099
rect 3137 -2040 3204 -2038
rect 3137 -3099 3144 -2040
rect 3197 -3099 3204 -2040
rect 3137 -3101 3204 -3099
rect 3257 -2040 3324 -2038
rect 4238 -2040 4305 -2038
rect 3257 -3099 3264 -2040
rect 3317 -3099 3324 -2040
rect 3377 -3095 3384 -2040
rect 3437 -3035 3444 -2040
rect 3812 -2801 3870 -2795
rect 3812 -2835 3824 -2801
rect 3812 -2841 3870 -2835
rect 3812 -2995 3870 -2989
rect 3812 -3029 3824 -2995
rect 3812 -3035 3870 -3029
rect 4238 -3039 4245 -2040
rect 3444 -3072 3504 -3039
rect 4179 -3068 4245 -3039
rect 4298 -3099 4305 -2040
rect 3257 -3101 3324 -3099
rect 3377 -3101 3503 -3099
rect 2898 -3128 3503 -3101
rect 4119 -3101 4305 -3099
rect 4358 -2040 4425 -2038
rect 4358 -3099 4365 -2040
rect 4418 -3099 4425 -2040
rect 4358 -3101 4425 -3099
rect 4478 -2040 4545 -2038
rect 5459 -2040 5526 -2038
rect 4478 -3099 4485 -2040
rect 4538 -3099 4545 -2040
rect 4598 -3095 4605 -2040
rect 4658 -3035 4665 -2040
rect 5033 -2801 5091 -2795
rect 5033 -2835 5045 -2801
rect 5033 -2841 5091 -2835
rect 5033 -2995 5091 -2989
rect 5033 -3029 5045 -2995
rect 5033 -3035 5091 -3029
rect 5459 -3039 5466 -2040
rect 4665 -3072 4725 -3039
rect 5400 -3068 5466 -3039
rect 5519 -3099 5526 -2040
rect 4478 -3101 4545 -3099
rect 4598 -3101 4724 -3099
rect 4119 -3128 4724 -3101
rect 5340 -3101 5526 -3099
rect 5579 -2040 5646 -2038
rect 5579 -3099 5586 -2040
rect 5639 -3099 5646 -2040
rect 5579 -3101 5646 -3099
rect 5699 -2040 5766 -2038
rect 6680 -2040 6747 -2038
rect 5699 -3099 5706 -2040
rect 5759 -3099 5766 -2040
rect 5819 -3095 5826 -2040
rect 5879 -3035 5886 -2040
rect 6254 -2801 6312 -2795
rect 6254 -2835 6266 -2801
rect 6254 -2841 6312 -2835
rect 6254 -2995 6312 -2989
rect 6254 -3029 6266 -2995
rect 6254 -3035 6312 -3029
rect 6680 -3039 6687 -2040
rect 5886 -3072 5946 -3039
rect 6621 -3068 6687 -3039
rect 6740 -3099 6747 -2040
rect 5699 -3101 5766 -3099
rect 5819 -3101 5945 -3099
rect 5340 -3128 5945 -3101
rect 6561 -3101 6747 -3099
rect 6800 -2040 6867 -2038
rect 6800 -3099 6807 -2040
rect 6860 -3099 6867 -2040
rect 6800 -3101 6867 -3099
rect 6920 -2040 6987 -2038
rect 6920 -3099 6927 -2040
rect 6980 -3099 6987 -2040
rect 7040 -3095 7047 -2040
rect 7100 -3035 7107 -2040
rect 7107 -3072 7167 -3039
rect 6920 -3101 6987 -3099
rect 7040 -3101 7166 -3099
rect 6561 -3128 7166 -3101
rect 1794 -3132 2282 -3128
rect 3015 -3132 3503 -3128
rect 4236 -3132 4724 -3128
rect 5457 -3132 5945 -3128
rect 6678 -3132 7166 -3128
rect 1129 -3149 1196 -3147
rect 1249 -3149 1375 -3147
rect 573 -3165 1375 -3149
rect 1794 -3165 2225 -3132
rect 3015 -3165 3446 -3132
rect 4236 -3165 4667 -3132
rect 5457 -3165 5888 -3132
rect 6678 -3165 7109 -3132
rect -33 -3167 364 -3165
rect -29 -3193 199 -3167
rect -29 -3197 214 -3193
rect -105 -3279 -92 -3197
rect -33 -3217 239 -3197
rect 281 -3215 364 -3167
rect 620 -3198 684 -3165
rect 700 -3198 764 -3165
rect 780 -3180 1375 -3165
rect 780 -3198 1318 -3180
rect 1841 -3198 1905 -3165
rect 1921 -3198 1985 -3165
rect 2001 -3198 2065 -3165
rect 2081 -3198 2145 -3165
rect 2161 -3198 2225 -3165
rect 3062 -3198 3126 -3165
rect 3142 -3198 3206 -3165
rect 3222 -3198 3286 -3165
rect 3302 -3198 3366 -3165
rect 3382 -3198 3446 -3165
rect 4283 -3198 4347 -3165
rect 4363 -3198 4427 -3165
rect 4443 -3198 4507 -3165
rect 4523 -3198 4587 -3165
rect 4603 -3198 4667 -3165
rect 5504 -3198 5568 -3165
rect 5584 -3198 5648 -3165
rect 5664 -3198 5728 -3165
rect 5744 -3198 5808 -3165
rect 5824 -3198 5888 -3165
rect 6725 -3198 6789 -3165
rect 6805 -3198 6869 -3165
rect 6885 -3198 6949 -3165
rect 6965 -3198 7029 -3165
rect 7045 -3198 7109 -3165
rect 807 -3213 871 -3198
rect 887 -3213 1318 -3198
rect -29 -3227 157 -3217
rect -29 -3231 -8 -3227
rect -71 -3245 -7 -3231
rect 39 -3245 205 -3231
rect -71 -3265 205 -3245
rect 934 -3246 998 -3213
rect 1014 -3246 1078 -3213
rect 1094 -3246 1158 -3213
rect 1174 -3246 1238 -3213
rect 1254 -3246 1318 -3213
rect -105 -3299 239 -3279
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
rect 0 -2400 200 -2200
rect 0 -2800 200 -2600
rect 0 -3200 200 -3000
use hgu_sw_cap  hgu_sw_cap_0
timestamp 1698477894
transform 1 0 1549 0 1 -732
box -53 514 1168 1775
use hgu_sw_cap  x3[0]
timestamp 1698477894
transform 1 0 1241 0 1 -3714
box -53 514 1168 1775
use hgu_sw_cap  x3[1]
timestamp 1698477894
transform 1 0 20 0 1 -3714
box -53 514 1168 1775
use hgu_sw_cap  x4[0]
timestamp 1698477894
transform 1 0 6125 0 1 -3714
box -53 514 1168 1775
use hgu_sw_cap  x4[1]
timestamp 1698477894
transform 1 0 4904 0 1 -3714
box -53 514 1168 1775
use hgu_sw_cap  x4[2]
timestamp 1698477894
transform 1 0 3683 0 1 -3714
box -53 514 1168 1775
use hgu_sw_cap  x4[3]
timestamp 1698477894
transform 1 0 2462 0 1 -3714
box -53 514 1168 1775
use hgu_sw_cap  x7
timestamp 1698477894
transform 1 0 334 0 1 -3762
box -53 514 1168 1775
use sky130_fd_sc_hd__inv_1  x10 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1697965495
transform 1 0 -33 0 1 -3200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x11
timestamp 1697965495
transform 1 0 -71 0 1 -3248
box -38 -48 314 592
use sky130_fd_pr__nfet_01v8_MVW3GX  XM1
timestamp 0
transform 1 0 574 0 1 -3150
box -263 -252 263 252
use sky130_fd_pr__nfet_01v8_L7T3GD  XM13
timestamp 0
transform 1 0 178 0 1 193
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_L7T3GD  XM15
timestamp 0
transform 1 0 547 0 1 140
box -211 -252 211 252
use sky130_fd_pr__pfet_01v8_hvt_M479BZ  XM46
timestamp 0
transform 1 0 916 0 1 96
box -211 -261 211 261
use sky130_fd_pr__pfet_01v8_hvt_M479BZ  XM47
timestamp 0
transform 1 0 1285 0 1 43
box -211 -261 211 261
use sky130_fd_pr__pfet_01v8_hvt_M433PY  XM48
timestamp 0
transform 1 0 101 0 1 -3088
box -263 -261 263 261
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 IN
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 OUT
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 VSS
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 {code\[0\]}
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 {code\[1\]}
port 5 nsew
flabel metal1 0 -2400 200 -2200 0 FreeSans 256 0 0 0 {code\[2\]}
port 6 nsew
flabel metal1 0 -2800 200 -2600 0 FreeSans 256 0 0 0 {code\[3\]}
port 7 nsew
flabel metal1 0 -3200 200 -3000 0 FreeSans 256 0 0 0 code_offset
port 8 nsew
<< end >>
