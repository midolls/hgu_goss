magic
tech sky130A
magscale 1 2
timestamp 1698469782
<< pwell >>
rect -2620 1602 -2594 1634
rect -2614 806 -2588 838
<< metal3 >>
rect -2940 2412 -2268 2414
rect -2940 2348 -2836 2412
rect -2772 2348 -2756 2412
rect -2692 2348 -2676 2412
rect -2612 2348 -2596 2412
rect -2532 2348 -2516 2412
rect -2452 2348 -2436 2412
rect -2372 2348 -2268 2412
rect -2940 2346 -2268 2348
rect -2940 2192 -2874 2346
rect -2940 2128 -2939 2192
rect -2875 2128 -2874 2192
rect -2940 2112 -2874 2128
rect -2940 2048 -2939 2112
rect -2875 2048 -2874 2112
rect -2940 2032 -2874 2048
rect -2940 1968 -2939 2032
rect -2875 1968 -2874 2032
rect -2940 1952 -2874 1968
rect -2940 1888 -2939 1952
rect -2875 1888 -2874 1952
rect -2940 1872 -2874 1888
rect -2940 1808 -2939 1872
rect -2875 1808 -2874 1872
rect -2940 1792 -2874 1808
rect -2940 1728 -2939 1792
rect -2875 1728 -2874 1792
rect -2940 1712 -2874 1728
rect -2940 1648 -2939 1712
rect -2875 1648 -2874 1712
rect -2940 1632 -2874 1648
rect -2940 1568 -2939 1632
rect -2875 1568 -2874 1632
rect -2940 1552 -2874 1568
rect -2940 1488 -2939 1552
rect -2875 1488 -2874 1552
rect -2940 1472 -2874 1488
rect -2940 1408 -2939 1472
rect -2875 1408 -2874 1472
rect -2940 1318 -2874 1408
rect -2814 1314 -2754 2346
rect -2694 1254 -2634 2284
rect -2574 1314 -2514 2346
rect -2454 1254 -2394 2284
rect -2334 2192 -2268 2346
rect -2334 2128 -2333 2192
rect -2269 2128 -2268 2192
rect -2334 2112 -2268 2128
rect -2334 2048 -2333 2112
rect -2269 2048 -2268 2112
rect -2334 2032 -2268 2048
rect -2334 1968 -2333 2032
rect -2269 1968 -2268 2032
rect -2334 1952 -2268 1968
rect -2334 1888 -2333 1952
rect -2269 1888 -2268 1952
rect -2334 1872 -2268 1888
rect -2334 1808 -2333 1872
rect -2269 1808 -2268 1872
rect -2334 1792 -2268 1808
rect -2334 1728 -2333 1792
rect -2269 1728 -2268 1792
rect -2334 1712 -2268 1728
rect -2334 1648 -2333 1712
rect -2269 1648 -2268 1712
rect -2334 1632 -2268 1648
rect -2334 1568 -2333 1632
rect -2269 1568 -2268 1632
rect -2334 1552 -2268 1568
rect -2334 1488 -2333 1552
rect -2269 1488 -2268 1552
rect -2334 1472 -2268 1488
rect -2334 1408 -2333 1472
rect -2269 1408 -2268 1472
rect -2334 1318 -2268 1408
rect -2940 1252 -2268 1254
rect -2940 1188 -2836 1252
rect -2772 1188 -2756 1252
rect -2692 1188 -2676 1252
rect -2612 1188 -2596 1252
rect -2532 1188 -2516 1252
rect -2452 1188 -2436 1252
rect -2372 1188 -2268 1252
rect -2940 1186 -2268 1188
rect -2940 1032 -2874 1122
rect -2940 968 -2939 1032
rect -2875 968 -2874 1032
rect -2940 952 -2874 968
rect -2940 888 -2939 952
rect -2875 888 -2874 952
rect -2940 872 -2874 888
rect -2940 808 -2939 872
rect -2875 808 -2874 872
rect -2940 792 -2874 808
rect -2940 728 -2939 792
rect -2875 728 -2874 792
rect -2940 712 -2874 728
rect -2940 648 -2939 712
rect -2875 648 -2874 712
rect -2940 632 -2874 648
rect -2940 568 -2939 632
rect -2875 568 -2874 632
rect -2940 552 -2874 568
rect -2940 488 -2939 552
rect -2875 488 -2874 552
rect -2940 472 -2874 488
rect -2940 408 -2939 472
rect -2875 408 -2874 472
rect -2940 392 -2874 408
rect -2940 328 -2939 392
rect -2875 328 -2874 392
rect -2940 312 -2874 328
rect -2940 248 -2939 312
rect -2875 248 -2874 312
rect -2940 94 -2874 248
rect -2814 156 -2754 1186
rect -2694 94 -2634 1126
rect -2574 156 -2514 1186
rect -2454 94 -2394 1126
rect -2334 1032 -2268 1122
rect -2334 968 -2333 1032
rect -2269 968 -2268 1032
rect -2334 952 -2268 968
rect -2334 888 -2333 952
rect -2269 888 -2268 952
rect -2334 872 -2268 888
rect -2334 808 -2333 872
rect -2269 808 -2268 872
rect -2334 792 -2268 808
rect -2334 728 -2333 792
rect -2269 728 -2268 792
rect -2334 712 -2268 728
rect -2334 648 -2333 712
rect -2269 648 -2268 712
rect -2334 632 -2268 648
rect -2334 568 -2333 632
rect -2269 568 -2268 632
rect -2334 552 -2268 568
rect -2334 488 -2333 552
rect -2269 488 -2268 552
rect -2334 472 -2268 488
rect -2334 408 -2333 472
rect -2269 408 -2268 472
rect -2334 392 -2268 408
rect -2334 328 -2333 392
rect -2269 328 -2268 392
rect -2334 312 -2268 328
rect -2334 248 -2333 312
rect -2269 248 -2268 312
rect -2334 94 -2268 248
rect -2940 92 -2268 94
rect -2940 28 -2836 92
rect -2772 28 -2756 92
rect -2692 28 -2676 92
rect -2612 28 -2596 92
rect -2532 28 -2516 92
rect -2452 28 -2436 92
rect -2372 28 -2268 92
rect -2940 26 -2268 28
<< via3 >>
rect -2836 2348 -2772 2412
rect -2756 2348 -2692 2412
rect -2676 2348 -2612 2412
rect -2596 2348 -2532 2412
rect -2516 2348 -2452 2412
rect -2436 2348 -2372 2412
rect -2939 2128 -2875 2192
rect -2939 2048 -2875 2112
rect -2939 1968 -2875 2032
rect -2939 1888 -2875 1952
rect -2939 1808 -2875 1872
rect -2939 1728 -2875 1792
rect -2939 1648 -2875 1712
rect -2939 1568 -2875 1632
rect -2939 1488 -2875 1552
rect -2939 1408 -2875 1472
rect -2333 2128 -2269 2192
rect -2333 2048 -2269 2112
rect -2333 1968 -2269 2032
rect -2333 1888 -2269 1952
rect -2333 1808 -2269 1872
rect -2333 1728 -2269 1792
rect -2333 1648 -2269 1712
rect -2333 1568 -2269 1632
rect -2333 1488 -2269 1552
rect -2333 1408 -2269 1472
rect -2836 1188 -2772 1252
rect -2756 1188 -2692 1252
rect -2676 1188 -2612 1252
rect -2596 1188 -2532 1252
rect -2516 1188 -2452 1252
rect -2436 1188 -2372 1252
rect -2939 968 -2875 1032
rect -2939 888 -2875 952
rect -2939 808 -2875 872
rect -2939 728 -2875 792
rect -2939 648 -2875 712
rect -2939 568 -2875 632
rect -2939 488 -2875 552
rect -2939 408 -2875 472
rect -2939 328 -2875 392
rect -2939 248 -2875 312
rect -2333 968 -2269 1032
rect -2333 888 -2269 952
rect -2333 808 -2269 872
rect -2333 728 -2269 792
rect -2333 648 -2269 712
rect -2333 568 -2269 632
rect -2333 488 -2269 552
rect -2333 408 -2269 472
rect -2333 328 -2269 392
rect -2333 248 -2269 312
rect -2836 28 -2772 92
rect -2756 28 -2692 92
rect -2676 28 -2612 92
rect -2596 28 -2532 92
rect -2516 28 -2452 92
rect -2436 28 -2372 92
<< metal4 >>
rect -2940 2412 -2268 2414
rect -2940 2348 -2836 2412
rect -2772 2348 -2756 2412
rect -2692 2348 -2676 2412
rect -2612 2348 -2596 2412
rect -2532 2348 -2516 2412
rect -2452 2348 -2436 2412
rect -2372 2348 -2268 2412
rect -2940 2346 -2268 2348
rect -2940 2192 -2874 2346
rect -2940 2128 -2939 2192
rect -2875 2128 -2874 2192
rect -2940 2112 -2874 2128
rect -2940 2048 -2939 2112
rect -2875 2048 -2874 2112
rect -2940 2032 -2874 2048
rect -2940 1968 -2939 2032
rect -2875 1968 -2874 2032
rect -2940 1952 -2874 1968
rect -2940 1888 -2939 1952
rect -2875 1888 -2874 1952
rect -2940 1872 -2874 1888
rect -2940 1808 -2939 1872
rect -2875 1808 -2874 1872
rect -2940 1792 -2874 1808
rect -2940 1728 -2939 1792
rect -2875 1728 -2874 1792
rect -2940 1712 -2874 1728
rect -2940 1648 -2939 1712
rect -2875 1648 -2874 1712
rect -2940 1632 -2874 1648
rect -2940 1568 -2939 1632
rect -2875 1568 -2874 1632
rect -2940 1552 -2874 1568
rect -2940 1488 -2939 1552
rect -2875 1488 -2874 1552
rect -2940 1472 -2874 1488
rect -2940 1408 -2939 1472
rect -2875 1408 -2874 1472
rect -2940 1318 -2874 1408
rect -2814 1254 -2754 2284
rect -2694 1314 -2634 2346
rect -2574 1254 -2514 2284
rect -2454 1314 -2394 2346
rect -2334 2192 -2268 2346
rect -2334 2128 -2333 2192
rect -2269 2128 -2268 2192
rect -2334 2112 -2268 2128
rect -2334 2048 -2333 2112
rect -2269 2048 -2268 2112
rect -2334 2032 -2268 2048
rect -2334 1968 -2333 2032
rect -2269 1968 -2268 2032
rect -2334 1952 -2268 1968
rect -2334 1888 -2333 1952
rect -2269 1888 -2268 1952
rect -2334 1872 -2268 1888
rect -2334 1808 -2333 1872
rect -2269 1808 -2268 1872
rect -2334 1792 -2268 1808
rect -2334 1728 -2333 1792
rect -2269 1728 -2268 1792
rect -2334 1712 -2268 1728
rect -2334 1648 -2333 1712
rect -2269 1648 -2268 1712
rect -2334 1632 -2268 1648
rect -2334 1568 -2333 1632
rect -2269 1568 -2268 1632
rect -2334 1552 -2268 1568
rect -2334 1488 -2333 1552
rect -2269 1488 -2268 1552
rect -2334 1472 -2268 1488
rect -2334 1408 -2333 1472
rect -2269 1408 -2268 1472
rect -2334 1318 -2268 1408
rect -2940 1252 -2268 1254
rect -2940 1188 -2836 1252
rect -2772 1188 -2756 1252
rect -2692 1188 -2676 1252
rect -2612 1188 -2596 1252
rect -2532 1188 -2516 1252
rect -2452 1188 -2436 1252
rect -2372 1188 -2268 1252
rect -2940 1186 -2268 1188
rect -2940 1032 -2874 1122
rect -2940 968 -2939 1032
rect -2875 968 -2874 1032
rect -2940 952 -2874 968
rect -2940 888 -2939 952
rect -2875 888 -2874 952
rect -2940 872 -2874 888
rect -2940 808 -2939 872
rect -2875 808 -2874 872
rect -2940 792 -2874 808
rect -2940 728 -2939 792
rect -2875 728 -2874 792
rect -2940 712 -2874 728
rect -2940 648 -2939 712
rect -2875 648 -2874 712
rect -2940 632 -2874 648
rect -2940 568 -2939 632
rect -2875 568 -2874 632
rect -2940 552 -2874 568
rect -2940 488 -2939 552
rect -2875 488 -2874 552
rect -2940 472 -2874 488
rect -2940 408 -2939 472
rect -2875 408 -2874 472
rect -2940 392 -2874 408
rect -2940 328 -2939 392
rect -2875 328 -2874 392
rect -2940 312 -2874 328
rect -2940 248 -2939 312
rect -2875 248 -2874 312
rect -2940 94 -2874 248
rect -2814 94 -2754 1126
rect -2694 156 -2634 1186
rect -2574 94 -2514 1126
rect -2454 156 -2394 1186
rect -2334 1032 -2268 1122
rect -2334 968 -2333 1032
rect -2269 968 -2268 1032
rect -2334 952 -2268 968
rect -2334 888 -2333 952
rect -2269 888 -2268 952
rect -2334 872 -2268 888
rect -2334 808 -2333 872
rect -2269 808 -2268 872
rect -2334 792 -2268 808
rect -2334 728 -2333 792
rect -2269 728 -2268 792
rect -2334 712 -2268 728
rect -2334 648 -2333 712
rect -2269 648 -2268 712
rect -2334 632 -2268 648
rect -2334 568 -2333 632
rect -2269 568 -2268 632
rect -2334 552 -2268 568
rect -2334 488 -2333 552
rect -2269 488 -2268 552
rect -2334 472 -2268 488
rect -2334 408 -2333 472
rect -2269 408 -2268 472
rect -2334 392 -2268 408
rect -2334 328 -2333 392
rect -2269 328 -2268 392
rect -2334 312 -2268 328
rect -2334 248 -2333 312
rect -2269 248 -2268 312
rect -2334 94 -2268 248
rect -2940 92 -2268 94
rect -2940 28 -2836 92
rect -2772 28 -2756 92
rect -2692 28 -2676 92
rect -2612 28 -2596 92
rect -2532 28 -2516 92
rect -2452 28 -2436 92
rect -2372 28 -2268 92
rect -2940 26 -2268 28
<< labels >>
flabel pwell -2614 806 -2588 838 0 FreeSans 160 0 0 0 x1.SUB
flabel metal4 -2556 472 -2530 504 0 FreeSans 320 0 0 0 x1.CBOT
flabel metal4 -2674 1062 -2648 1094 0 FreeSans 320 0 0 0 x1.CTOP
flabel pwell -2620 1602 -2594 1634 0 FreeSans 160 0 0 0 x2.SUB
flabel metal4 -2678 1936 -2652 1968 0 FreeSans 320 0 0 0 x2.CBOT
flabel metal4 -2560 1346 -2534 1378 0 FreeSans 320 0 0 0 x2.CTOP
<< end >>
