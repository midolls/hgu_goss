magic
tech sky130A
timestamp 1697681522
use hgu_cdac_unit  x1
timestamp 1697641878
transform 1 0 3429 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x2[0]
timestamp 1697641878
transform 1 0 3859 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x2[1]
timestamp 1697641878
transform 1 0 3644 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x3[0]
timestamp 1697641878
transform 1 0 4719 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x3[1]
timestamp 1697641878
transform 1 0 4504 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x3[2]
timestamp 1697641878
transform 1 0 4289 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x3[3]
timestamp 1697641878
transform 1 0 4074 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x4[0]
timestamp 1697641878
transform 1 0 6439 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x4[1]
timestamp 1697641878
transform 1 0 6224 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x4[2]
timestamp 1697641878
transform 1 0 6009 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x4[3]
timestamp 1697641878
transform 1 0 5794 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x4[4]
timestamp 1697641878
transform 1 0 5579 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x4[5]
timestamp 1697641878
transform 1 0 5364 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x4[6]
timestamp 1697641878
transform 1 0 5149 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x4[7]
timestamp 1697641878
transform 1 0 4934 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x5[0]
timestamp 1697641878
transform 1 0 9879 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x5[1]
timestamp 1697641878
transform 1 0 9664 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x5[2]
timestamp 1697641878
transform 1 0 9449 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x5[3]
timestamp 1697641878
transform 1 0 9234 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x5[4]
timestamp 1697641878
transform 1 0 9019 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x5[5]
timestamp 1697641878
transform 1 0 8804 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x5[6]
timestamp 1697641878
transform 1 0 8589 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x5[7]
timestamp 1697641878
transform 1 0 8374 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x5[8]
timestamp 1697641878
transform 1 0 8159 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x5[9]
timestamp 1697641878
transform 1 0 7944 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x5[10]
timestamp 1697641878
transform 1 0 7729 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x5[11]
timestamp 1697641878
transform 1 0 7514 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x5[12]
timestamp 1697641878
transform 1 0 7299 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x5[13]
timestamp 1697641878
transform 1 0 7084 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x5[14]
timestamp 1697641878
transform 1 0 6869 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x5[15]
timestamp 1697641878
transform 1 0 6654 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x6[0]
timestamp 1697641878
transform 1 0 16759 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x6[1]
timestamp 1697641878
transform 1 0 16544 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x6[2]
timestamp 1697641878
transform 1 0 16329 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x6[3]
timestamp 1697641878
transform 1 0 16114 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x6[4]
timestamp 1697641878
transform 1 0 15899 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x6[5]
timestamp 1697641878
transform 1 0 15684 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x6[6]
timestamp 1697641878
transform 1 0 15469 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x6[7]
timestamp 1697641878
transform 1 0 15254 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x6[8]
timestamp 1697641878
transform 1 0 15039 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x6[9]
timestamp 1697641878
transform 1 0 14824 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x6[10]
timestamp 1697641878
transform 1 0 14609 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x6[11]
timestamp 1697641878
transform 1 0 14394 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x6[12]
timestamp 1697641878
transform 1 0 14179 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x6[13]
timestamp 1697641878
transform 1 0 13964 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x6[14]
timestamp 1697641878
transform 1 0 13749 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x6[15]
timestamp 1697641878
transform 1 0 13534 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x6[16]
timestamp 1697641878
transform 1 0 13319 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x6[17]
timestamp 1697641878
transform 1 0 13104 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x6[18]
timestamp 1697641878
transform 1 0 12889 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x6[19]
timestamp 1697641878
transform 1 0 12674 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x6[20]
timestamp 1697641878
transform 1 0 12459 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x6[21]
timestamp 1697641878
transform 1 0 12244 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x6[22]
timestamp 1697641878
transform 1 0 12029 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x6[23]
timestamp 1697641878
transform 1 0 11814 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x6[24]
timestamp 1697641878
transform 1 0 11599 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x6[25]
timestamp 1697641878
transform 1 0 11384 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x6[26]
timestamp 1697641878
transform 1 0 11169 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x6[27]
timestamp 1697641878
transform 1 0 10954 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x6[28]
timestamp 1697641878
transform 1 0 10739 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x6[29]
timestamp 1697641878
transform 1 0 10524 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x6[30]
timestamp 1697641878
transform 1 0 10309 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x6[31]
timestamp 1697641878
transform 1 0 10094 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x7[0]
timestamp 1697641878
transform 1 0 30519 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x7[1]
timestamp 1697641878
transform 1 0 30304 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x7[2]
timestamp 1697641878
transform 1 0 30089 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x7[3]
timestamp 1697641878
transform 1 0 29874 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x7[4]
timestamp 1697641878
transform 1 0 29659 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x7[5]
timestamp 1697641878
transform 1 0 29444 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x7[6]
timestamp 1697641878
transform 1 0 29229 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x7[7]
timestamp 1697641878
transform 1 0 29014 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x7[8]
timestamp 1697641878
transform 1 0 28799 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x7[9]
timestamp 1697641878
transform 1 0 28584 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x7[10]
timestamp 1697641878
transform 1 0 28369 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x7[11]
timestamp 1697641878
transform 1 0 28154 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x7[12]
timestamp 1697641878
transform 1 0 27939 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x7[13]
timestamp 1697641878
transform 1 0 27724 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x7[14]
timestamp 1697641878
transform 1 0 27509 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x7[15]
timestamp 1697641878
transform 1 0 27294 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x7[16]
timestamp 1697641878
transform 1 0 27079 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x7[17]
timestamp 1697641878
transform 1 0 26864 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x7[18]
timestamp 1697641878
transform 1 0 26649 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x7[19]
timestamp 1697641878
transform 1 0 26434 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x7[20]
timestamp 1697641878
transform 1 0 26219 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x7[21]
timestamp 1697641878
transform 1 0 26004 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x7[22]
timestamp 1697641878
transform 1 0 25789 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x7[23]
timestamp 1697641878
transform 1 0 25574 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x7[24]
timestamp 1697641878
transform 1 0 25359 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x7[25]
timestamp 1697641878
transform 1 0 25144 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x7[26]
timestamp 1697641878
transform 1 0 24929 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x7[27]
timestamp 1697641878
transform 1 0 24714 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x7[28]
timestamp 1697641878
transform 1 0 24499 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x7[29]
timestamp 1697641878
transform 1 0 24284 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x7[30]
timestamp 1697641878
transform 1 0 24069 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x7[31]
timestamp 1697641878
transform 1 0 23854 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x7[32]
timestamp 1697641878
transform 1 0 23639 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x7[33]
timestamp 1697641878
transform 1 0 23424 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x7[34]
timestamp 1697641878
transform 1 0 23209 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x7[35]
timestamp 1697641878
transform 1 0 22994 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x7[36]
timestamp 1697641878
transform 1 0 22779 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x7[37]
timestamp 1697641878
transform 1 0 22564 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x7[38]
timestamp 1697641878
transform 1 0 22349 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x7[39]
timestamp 1697641878
transform 1 0 22134 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x7[40]
timestamp 1697641878
transform 1 0 21919 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x7[41]
timestamp 1697641878
transform 1 0 21704 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x7[42]
timestamp 1697641878
transform 1 0 21489 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x7[43]
timestamp 1697641878
transform 1 0 21274 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x7[44]
timestamp 1697641878
transform 1 0 21059 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x7[45]
timestamp 1697641878
transform 1 0 20844 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x7[46]
timestamp 1697641878
transform 1 0 20629 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x7[47]
timestamp 1697641878
transform 1 0 20414 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x7[48]
timestamp 1697641878
transform 1 0 20199 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x7[49]
timestamp 1697641878
transform 1 0 19984 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x7[50]
timestamp 1697641878
transform 1 0 19769 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x7[51]
timestamp 1697641878
transform 1 0 19554 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x7[52]
timestamp 1697641878
transform 1 0 19339 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x7[53]
timestamp 1697641878
transform 1 0 19124 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x7[54]
timestamp 1697641878
transform 1 0 18909 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x7[55]
timestamp 1697641878
transform 1 0 18694 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x7[56]
timestamp 1697641878
transform 1 0 18479 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x7[57]
timestamp 1697641878
transform 1 0 18264 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x7[58]
timestamp 1697641878
transform 1 0 18049 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x7[59]
timestamp 1697641878
transform 1 0 17834 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x7[60]
timestamp 1697641878
transform 1 0 17619 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x7[61]
timestamp 1697641878
transform 1 0 17404 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x7[62]
timestamp 1697641878
transform 1 0 17189 0 1 900
box 0 300 242 759
use hgu_cdac_unit  x7[63]
timestamp 1697641878
transform 1 0 16974 0 1 900
box 0 300 242 759
<< end >>
