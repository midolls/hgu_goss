* NGSPICE file created from hgu_cdac_cap_4.ext - technology: sky130A


* Top level circuit hgu_cdac_cap_4

C0 hgu_cdac_cap_2_1.hgu_cdac_unit_1.C1 hgu_cdac_cap_2_1.hgu_cdac_unit_1.C0 4.31f
C1 hgu_cdac_cap_2_1.hgu_cdac_unit_1.C1 hgu_cdac_cap_2_1.hgu_cdac_unit_0.C1 8.87f
C2 hgu_cdac_cap_2_1.hgu_cdac_unit_1.C1 hgu_cdac_cap_2_0.hgu_cdac_unit_1.C0 4.31f
C3 hgu_cdac_cap_2_1.hgu_cdac_unit_1.C1 VSUBS 1.68f $ **FLOATING
C4 hgu_cdac_cap_2_1.hgu_cdac_unit_0.C1 VSUBS 1.7f $ **FLOATING
.end

