* NGSPICE file created from hgu_vgen_vref_flat.ext - technology: sky130A

.subckt adc_vcm_generator VDD vcm clk VSS
X0 vcm.t8 VSS.t282 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X1 vcm.t9 VSS.t280 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X2 a_4324_38050# a_4147_38050# VSS.t87 VSS.t76 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X3 VDD.t57 a_3404_37506# a_3510_37506# VDD.t56 sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X4 mimtop2 VSS.t39 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X5 mimtop1.t7 phi1 vcm.t7 VSS.t329 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=0.5
X6 phi1_n a_3172_38568# VSS.t317 VSS.t316 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7 VDD.t113 sky130_fd_sc_hd__inv_1_3.Y sky130_fd_sc_hd__nand2_1_0.Y VDD.t112 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8 VDD.t99 sky130_fd_sc_hd__nand2_1_0.Y a_2024_38050# VDD.t98 sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X9 VSS.t46 a_3121_38050# a_3227_38050# VSS.t45 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X10 phi2_n a_3172_36936# VSS.t60 VSS.t59 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 vcm.t10 VSS.t278 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X12 VDD.t143 sky130_fd_sc_hd__inv_1_2.Y sky130_fd_sc_hd__nand2_1_1.Y VDD.t142 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X13 mimtop2 VSS.t38 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X14 a_4041_38050# a_3864_38050# VSS.t91 VSS.t90 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X15 a_3121_37506# a_2944_37506# VDD.t11 VDD.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X16 VDD.t144 VSS.t42 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X17 vcm.t11 VSS.t276 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X18 VDD.t121 sky130_fd_sc_hd__nand2_1_1.Y a_2024_37506# VDD.t120 sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X19 vcm.t12 VSS.t274 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X20 a_2201_37506# a_2024_37506# VSS.t319 VSS.t51 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X21 vcm.t13 VSS.t272 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X22 VSS.t75 a_2201_37506# a_2307_37506# VSS.t74 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X23 VSS.t58 a_3172_36936# phi2_n VSS.t57 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X24 vcm.t14 VSS.t270 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X25 sky130_fd_sc_hd__nand2_1_1.Y sky130_fd_sc_hd__inv_1_4.Y VDD.t97 VDD.t96 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X26 mimtop1.t8 mimbot1.t41 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X27 phi1 a_3724_38568# VSS.t303 VSS.t302 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X28 VSS.t301 a_3724_38568# phi1 VSS.t300 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X29 VSS.t119 a_3404_38050# a_3510_38050# VSS.t96 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X30 sky130_fd_sc_hd__dlymetal6s6s_1_4.A a_2590_37506# VDD.t35 VDD.t34 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X31 mimtop2 VSS.t37 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X32 mimtop1.t9 mimbot1.t40 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X33 vcm.t15 VSS.t268 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X34 mimtop2 VSS.t36 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X35 mimtop1.t10 mimbot1.t39 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X36 mimtop1.t11 mimbot1.t38 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X37 mimtop1.t12 mimbot1.t37 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X38 vcm.t16 VSS.t266 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X39 a_3121_38050# a_2944_38050# VSS.t295 VSS.t49 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X40 VSS.t294 sky130_fd_sc_hd__nand2_1_0.Y a_2024_38050# VSS.t293 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X41 mimtop2 VSS.t35 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X42 mimtop2 VSS.t34 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X43 vcm.t17 VSS.t264 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X44 VSS.t290 a_2484_37506# a_2590_37506# VSS.t288 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X45 mimtop2 VSS.t33 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X46 VSS.t118 a_3724_36936# phi2 VSS.t117 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X47 vcm.t18 VSS.t262 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X48 vcm.t19 VSS.t260 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X49 phi1_n a_3172_38568# VSS.t315 VSS.t314 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X50 VDD.t29 sky130_fd_sc_hd__inv_1_2.A sky130_fd_sc_hd__inv_1_2.Y VDD.t28 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X51 sky130_fd_sc_hd__dlymetal6s6s_1_2.A a_2590_38050# VSS.t109 VSS.t72 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X52 vcm.t20 VSS.t258 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X53 VSS.t328 phi1 mimbot1.t47 VSS.t327 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=0.5
X54 mimtop1.t13 mimbot1.t36 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X55 mimtop2 VSS.t32 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X56 vcm.t21 VSS.t256 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X57 VDD.t119 phi2_n mimtop1.t5 VDD.t118 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=0.5
X58 vcm.t22 VSS.t254 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X59 mimtop2 VSS.t31 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X60 mimtop1.t14 mimbot1.t35 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X61 a_3172_38568# sky130_fd_sc_hd__inv_1_2.Y VDD.t141 VDD.t140 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X62 vcm.t23 VSS.t252 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X63 vcm.t24 VSS.t250 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X64 mimtop1.t15 mimbot1.t34 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X65 mimtop1.t16 mimbot1.t33 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X66 VSS.t313 a_3172_38568# phi1_n VSS.t312 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X67 sky130_fd_sc_hd__dlymetal6s6s_1_3.A a_3510_38050# VDD.t133 VDD.t132 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X68 VSS.t56 a_3172_36936# phi2_n VSS.t55 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X69 mimtop2 VSS.t30 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X70 vcm.t25 VSS.t248 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X71 mimtop2 VSS.t29 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X72 VDD.t145 VSS.t43 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X73 VDD.t146 VSS.t105 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X74 mimtop2 VSS.t28 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X75 vcm.t26 VSS.t246 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X76 VSS.t86 a_4041_37506# a_4147_37506# VSS.t85 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X77 mimtop1.t4 phi2_n VDD.t117 VDD.t116 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=0.5
X78 VDD.t147 VSS.t107 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X79 sky130_fd_sc_hd__inv_1_1.A a_4430_37506# VDD.t65 VDD.t64 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X80 vcm.t27 VSS.t244 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X81 sky130_fd_sc_hd__dlymetal6s6s_1_5.A a_3510_37506# VSS.t99 VSS.t98 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X82 phi2 a_3724_36936# VDD.t77 VDD.t76 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X83 mimtop1.t17 mimbot1.t32 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X84 mimbot1.t45 phi2_n mimtop2 VDD.t115 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=0.5
X85 vcm.t28 VSS.t242 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X86 VSS.t299 a_3724_38568# phi1 VSS.t298 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X87 mimtop2 VSS.t27 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X88 vcm.t29 VSS.t240 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X89 vcm.t30 VSS.t238 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X90 vcm.t31 VSS.t236 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X91 mimtop1.t18 mimbot1.t31 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X92 mimtop1.t19 mimbot1.t30 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X93 VSS.t84 a_4324_37506# a_4430_37506# VSS.t83 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X94 a_3724_36936# sky130_fd_sc_hd__inv_1_3.A VDD.t33 VDD.t32 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X95 mimtop2 VSS.t26 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X96 vcm.t32 VSS.t234 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X97 VDD.t25 sky130_fd_sc_hd__inv_1_1.A sky130_fd_sc_hd__inv_1_3.A VDD.t24 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X98 vcm.t33 VSS.t232 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X99 mimtop1.t20 mimbot1.t29 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X100 a_2484_38050# a_2307_38050# VDD.t3 VDD.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X101 mimtop2 VSS.t25 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X102 mimtop2 VSS.t24 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X103 sky130_fd_sc_hd__inv_1_0.A a_4430_38050# VSS.t110 VSS.t103 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X104 mimtop2 phi2 mimbot1.t1 VSS.t82 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=0.5
X105 vcm.t34 VSS.t230 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X106 VDD.t91 a_2201_38050# a_2307_38050# VDD.t90 sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X107 VDD.t148 VSS.t92 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X108 vcm.t35 VSS.t228 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X109 mimtop2 VSS.t23 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X110 vcm.t36 VSS.t226 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X111 vcm.t37 VSS.t224 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X112 a_1794_38050# clk.t0 sky130_fd_sc_hd__nand2_1_0.Y VSS.t44 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X113 a_3404_37506# a_3227_37506# VDD.t7 VDD.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X114 VSS.t311 a_3172_38568# phi1_n VSS.t310 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X115 VDD.t37 a_2201_37506# a_2307_37506# VDD.t36 sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X116 a_2484_37506# a_2307_37506# VSS.t61 VSS.t40 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X117 VSS.t123 sky130_fd_sc_hd__dlymetal6s6s_1_5.A a_3864_37506# VSS.t122 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X118 vcm.t38 VSS.t222 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X119 mimtop2 VSS.t22 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X120 VSS.t71 sky130_fd_sc_hd__inv_1_3.A sky130_fd_sc_hd__inv_1_3.Y VSS.t70 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X121 vcm.t39 VSS.t220 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X122 vcm.t40 VSS.t218 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X123 mimtop2 VSS.t21 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X124 VDD.t93 a_2484_38050# a_2590_38050# VDD.t92 sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X125 phi2_n a_3172_36936# VDD.t21 VDD.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X126 mimtop1.t21 mimbot1.t28 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X127 mimtop1.t22 mimbot1.t27 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X128 vcm.t41 VSS.t216 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X129 vcm.t42 VSS.t214 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X130 vcm.t43 VSS.t212 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X131 mimtop1.t23 mimbot1.t26 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X132 vcm.t44 VSS.t210 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X133 a_3172_36936# sky130_fd_sc_hd__inv_1_3.Y VSS.t307 VSS.t306 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X134 vcm.t45 VSS.t208 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X135 mimtop2 VSS.t20 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X136 vcm.t3 phi1_n mimtop1.t3 VDD.t89 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=0.5
X137 a_3404_38050# a_3227_38050# VSS.t78 VSS.t47 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X138 VDD.t95 a_2484_37506# a_2590_37506# VDD.t94 sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X139 vcm.t46 VSS.t206 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X140 mimtop2 VSS.t19 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X141 mimtop1.t24 mimbot1.t25 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X142 VSS.t287 a_2201_38050# a_2307_38050# VSS.t74 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X143 vcm.t47 VSS.t204 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X144 VSS.t309 sky130_fd_sc_hd__dlymetal6s6s_1_4.A a_2944_37506# VSS.t101 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X145 a_2201_37506# a_2024_37506# VDD.t135 VDD.t134 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X146 vcm.t48 VSS.t202 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X147 phi2 a_3724_36936# VDD.t75 VDD.t74 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X148 mimtop2 VSS.t18 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X149 vcm.t49 VSS.t200 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X150 vcm.t50 VSS.t198 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X151 VDD.t73 a_3724_36936# phi2 VDD.t72 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X152 vcm.t51 VSS.t196 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X153 a_4324_38050# a_4147_38050# VDD.t49 VDD.t48 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X154 mimtop1.t25 mimbot1.t24 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X155 vcm.t52 VSS.t194 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X156 VDD.t83 a_4041_38050# a_4147_38050# VDD.t82 sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X157 mimtop1.t26 mimbot1.t23 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X158 mimtop1.t27 mimbot1.t22 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X159 vcm.t53 VSS.t192 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X160 a_4041_38050# a_3864_38050# VDD.t53 VDD.t52 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X161 VSS.t289 a_2484_38050# a_2590_38050# VSS.t288 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X162 mimtop2 VSS.t17 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X163 mimtop2 VSS.t16 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X164 vcm.t54 VSS.t190 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X165 VSS.t67 sky130_fd_sc_hd__inv_1_2.A sky130_fd_sc_hd__inv_1_2.Y VSS.t66 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X166 mimtop2 VSS.t15 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X167 mimtop2 VSS.t14 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X168 mimbot1.t46 phi1 VSS.t326 VSS.t325 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=0.5
X169 mimtop2 phi1 vcm.t5 VSS.t324 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=0.5
X170 a_2201_38050# a_2024_38050# VSS.t52 VSS.t51 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X171 VDD.t47 a_4041_37506# a_4147_37506# VDD.t46 sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X172 vcm.t55 VSS.t188 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X173 phi1 a_3724_38568# VDD.t109 VDD.t108 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X174 sky130_fd_sc_hd__inv_1_4.Y clk.t1 VSS.t121 VSS.t120 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X175 a_4324_37506# a_4147_37506# VSS.t77 VSS.t76 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X176 phi2_n a_3172_36936# VDD.t19 VDD.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X177 vcm.t56 VSS.t186 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X178 VSS.t305 sky130_fd_sc_hd__inv_1_3.Y a_1794_38050# VSS.t304 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X179 VDD.t149 VSS.t94 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X180 vcm.t57 VSS.t184 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X181 a_3172_38568# sky130_fd_sc_hd__inv_1_2.Y VSS.t332 VSS.t331 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X182 VDD.t55 a_4324_38050# a_4430_38050# VDD.t54 sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X183 a_4041_37506# a_3864_37506# VSS.t320 VSS.t90 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X184 a_3724_38568# sky130_fd_sc_hd__inv_1_2.A VDD.t27 VDD.t26 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X185 vcm.t4 phi1 mimtop2 VSS.t323 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=0.5
X186 VDD.t51 sky130_fd_sc_hd__inv_1_0.A sky130_fd_sc_hd__inv_1_2.A VDD.t50 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X187 vcm.t58 VSS.t182 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X188 a_3121_38050# a_2944_38050# VDD.t101 VDD.t100 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X189 vcm.t59 VSS.t180 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X190 mimtop1.t28 mimbot1.t21 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X191 VDD.t17 a_3172_36936# phi2_n VDD.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X192 mimtop2 VSS.t13 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X193 mimtop1.t29 mimbot1.t20 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X194 mimtop1.t30 mimbot1.t19 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X195 VDD.t45 a_4324_37506# a_4430_37506# VDD.t44 sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X196 vcm.t60 VSS.t178 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X197 mimtop1.t31 mimbot1.t18 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X198 VSS.t286 phi1_n mimbot1.t43 VDD.t88 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=0.5
X199 VSS.t284 a_4041_38050# a_4147_38050# VSS.t85 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X200 mimtop2 VSS.t12 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X201 mimtop2 VSS.t11 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X202 mimtop2 VSS.t10 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X203 vcm.t61 VSS.t176 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X204 vcm.t62 VSS.t174 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X205 mimtop1.t32 mimbot1.t17 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X206 mimtop2 phi1_n vcm.t1 VDD.t87 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=0.5
X207 sky130_fd_sc_hd__dlymetal6s6s_1_2.A a_2590_38050# VDD.t67 VDD.t66 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X208 sky130_fd_sc_hd__nand2_1_1.Y sky130_fd_sc_hd__inv_1_2.Y a_1798_37826# VSS.t330 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X209 VDD.t139 sky130_fd_sc_hd__dlymetal6s6s_1_3.A a_3864_38050# VDD.t138 sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X210 a_3121_37506# a_2944_37506# VSS.t50 VSS.t49 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X211 VDD.t43 phi2 mimtop1.t1 VSS.t81 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=0.5
X212 vcm.t63 VSS.t172 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X213 VSS.t100 a_3121_37506# a_3227_37506# VSS.t45 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X214 vcm.t6 phi1 mimtop1.t6 VSS.t322 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=0.5
X215 phi1_n a_3172_38568# VDD.t131 VDD.t130 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X216 VDD.t71 a_3724_36936# phi2 VDD.t70 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X217 vcm.t64 VSS.t170 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X218 VSS.t95 a_4324_38050# a_4430_38050# VSS.t83 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X219 sky130_fd_sc_hd__dlymetal6s6s_1_5.A a_3510_37506# VDD.t59 VDD.t58 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X220 VDD.t81 sky130_fd_sc_hd__dlymetal6s6s_1_5.A a_3864_37506# VDD.t80 sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X221 vcm.t65 VSS.t168 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X222 mimtop1.t33 mimbot1.t16 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X223 vcm.t0 phi1_n mimtop2 VDD.t86 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=0.5
X224 a_1798_37826# sky130_fd_sc_hd__inv_1_4.Y VSS.t292 VSS.t291 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X225 sky130_fd_sc_hd__dlymetal6s6s_1_4.A a_2590_37506# VSS.t73 VSS.t72 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X226 mimtop1.t0 phi2 VDD.t42 VSS.t80 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=0.5
X227 vcm.t66 VSS.t166 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X228 mimtop1.t34 mimbot1.t15 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X229 vcm.t67 VSS.t164 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X230 mimtop2 VSS.t9 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X231 VDD.t63 sky130_fd_sc_hd__dlymetal6s6s_1_2.A a_2944_38050# VDD.t62 sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X232 mimbot1.t0 phi2 mimtop2 VSS.t79 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=0.5
X233 mimtop2 VSS.t8 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X234 VSS.t97 a_3404_37506# a_3510_37506# VSS.t96 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X235 mimtop1.t35 mimbot1.t14 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X236 vcm.t68 VSS.t162 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X237 phi1 a_3724_38568# VDD.t107 VDD.t106 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X238 VDD.t105 a_3724_38568# phi1 VDD.t104 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X239 VSS.t321 sky130_fd_sc_hd__dlymetal6s6s_1_3.A a_3864_38050# VSS.t122 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X240 VDD.t15 a_3172_36936# phi2_n VDD.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X241 vcm.t69 VSS.t160 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X242 sky130_fd_sc_hd__dlymetal6s6s_1_3.A a_3510_38050# VSS.t318 VSS.t98 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X243 VDD.t123 sky130_fd_sc_hd__dlymetal6s6s_1_4.A a_2944_37506# VDD.t122 sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X244 VSS.t308 sky130_fd_sc_hd__nand2_1_1.Y a_2024_37506# VSS.t293 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X245 phi2 a_3724_36936# VSS.t116 VSS.t115 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X246 vcm.t70 VSS.t158 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X247 vcm.t71 VSS.t156 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X248 vcm.t72 VSS.t154 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X249 a_2484_37506# a_2307_37506# VDD.t23 VDD.t22 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X250 mimtop1.t36 mimbot1.t13 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X251 mimtop1.t37 mimbot1.t12 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X252 vcm.t73 VSS.t152 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X253 vcm.t74 VSS.t150 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X254 mimtop1.t2 phi1_n vcm.t2 VDD.t85 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=0.5
X255 a_3724_36936# sky130_fd_sc_hd__inv_1_3.A VSS.t69 VSS.t68 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X256 VSS.t63 sky130_fd_sc_hd__inv_1_1.A sky130_fd_sc_hd__inv_1_3.A VSS.t62 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X257 vcm.t75 VSS.t148 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X258 sky130_fd_sc_hd__inv_1_0.A a_4430_38050# VDD.t69 VDD.t68 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X259 phi1_n a_3172_38568# VDD.t129 VDD.t128 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X260 mimtop2 VSS.t7 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X261 mimtop1.t38 mimbot1.t11 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X262 vcm.t76 VSS.t146 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X263 vcm.t77 VSS.t144 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X264 VSS.t102 sky130_fd_sc_hd__dlymetal6s6s_1_2.A a_2944_38050# VSS.t101 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X265 mimtop1.t39 mimbot1.t10 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X266 sky130_fd_sc_hd__nand2_1_0.Y clk.t2 VDD.t1 VDD.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X267 vcm.t78 VSS.t142 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X268 vcm.t79 VSS.t140 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X269 mimtop2 VSS.t6 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X270 a_2484_38050# a_2307_38050# VSS.t41 VSS.t40 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X271 sky130_fd_sc_hd__inv_1_1.A a_4430_37506# VSS.t104 VSS.t103 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X272 VDD.t127 a_3172_38568# phi1_n VDD.t126 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X273 mimtop2 VSS.t5 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X274 mimtop1.t40 mimbot1.t9 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X275 phi2_n a_3172_36936# VSS.t54 VSS.t53 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X276 mimtop1.t41 mimbot1.t8 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X277 vcm.t80 VSS.t138 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X278 mimtop2 phi2_n mimbot1.t44 VDD.t114 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=0.5
X279 mimtop2 VSS.t4 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X280 phi1 a_3724_38568# VSS.t297 VSS.t296 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X281 a_3404_38050# a_3227_38050# VDD.t41 VDD.t40 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X282 VDD.t31 sky130_fd_sc_hd__inv_1_3.A sky130_fd_sc_hd__inv_1_3.Y VDD.t30 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X283 vcm.t81 VSS.t136 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X284 vcm.t82 VSS.t134 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X285 mimtop2 VSS.t3 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X286 mimtop1.t42 mimbot1.t7 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X287 vcm.t83 VSS.t132 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X288 VDD.t5 a_3121_38050# a_3227_38050# VDD.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X289 mimtop1.t43 mimbot1.t6 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X290 mimtop1.t44 mimbot1.t5 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X291 vcm.t84 VSS.t130 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X292 a_3724_38568# sky130_fd_sc_hd__inv_1_2.A VSS.t65 VSS.t64 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X293 VDD.t103 a_3724_38568# phi1 VDD.t102 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X294 VSS.t89 sky130_fd_sc_hd__inv_1_0.A sky130_fd_sc_hd__inv_1_2.A VSS.t88 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X295 sky130_fd_sc_hd__inv_1_4.Y clk.t3 VDD.t9 VDD.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X296 a_4324_37506# a_4147_37506# VDD.t39 VDD.t38 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X297 a_3172_36936# sky130_fd_sc_hd__inv_1_3.Y VDD.t111 VDD.t110 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X298 mimtop2 VSS.t2 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X299 a_3404_37506# a_3227_37506# VSS.t48 VSS.t47 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X300 VDD.t61 a_3121_37506# a_3227_37506# VDD.t60 sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X301 phi2 a_3724_36936# VSS.t114 VSS.t113 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X302 VSS.t112 a_3724_36936# phi2 VSS.t111 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X303 a_4041_37506# a_3864_37506# VDD.t137 VDD.t136 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X304 mimbot1.t42 phi1_n VSS.t285 VDD.t84 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=0.5
X305 mimtop1.t45 mimbot1.t4 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X306 vcm.t85 VSS.t128 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X307 vcm.t86 VSS.t126 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X308 VDD.t79 a_3404_38050# a_3510_38050# VDD.t78 sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X309 mimtop1.t46 mimbot1.t3 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X310 vcm.t87 VSS.t124 error sky130_fd_pr__cap_var_lvt w=16.4 l=16
X311 a_2201_38050# a_2024_38050# VDD.t13 VDD.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X312 mimtop2 VSS.t1 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X313 VDD.t125 a_3172_38568# phi1_n VDD.t124 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X314 mimtop2 VSS.t0 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X315 mimtop1.t47 mimbot1.t2 sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
R0 vcm.n752 vcm.t0 122.98
R1 vcm.n753 vcm.t1 122.98
R2 vcm.n755 vcm.t2 122.959
R3 vcm.n756 vcm.t3 122.959
R4 vcm.n755 vcm.t7 78.1964
R5 vcm.n752 vcm.t4 74.3032
R6 vcm.n754 vcm.t5 35.0208
R7 vcm.n757 vcm.t6 34.9023
R8 vcm.n759 vcm.n758 30.2261
R9 vcm.n387 vcm.t45 27.8779
R10 vcm.n75 vcm.t15 27.8779
R11 vcm.n62 vcm.t41 27.8779
R12 vcm.n106 vcm.t16 27.8779
R13 vcm.n120 vcm.t44 27.8779
R14 vcm.n28 vcm.t58 27.8779
R15 vcm.n919 vcm.t25 27.8779
R16 vcm.n501 vcm.t60 27.8779
R17 vcm.n297 vcm.t23 27.8779
R18 vcm.n373 vcm.t54 27.8779
R19 vcm.n488 vcm.t24 27.8779
R20 vcm.n267 vcm.t67 27.8779
R21 vcm.n187 vcm.t73 27.8779
R22 vcm.n178 vcm.t74 27.8779
R23 vcm.n169 vcm.t70 27.8779
R24 vcm.n160 vcm.t68 27.8779
R25 vcm.n243 vcm.t61 27.8779
R26 vcm.n232 vcm.t86 27.8779
R27 vcm.n221 vcm.t36 27.8779
R28 vcm.n341 vcm.t57 27.8779
R29 vcm.n415 vcm.t46 27.8779
R30 vcm.n472 vcm.t22 27.8779
R31 vcm.n538 vcm.t59 27.8779
R32 vcm.n527 vcm.t65 27.8779
R33 vcm.n516 vcm.t72 27.8779
R34 vcm.n715 vcm.t33 27.8779
R35 vcm.n644 vcm.t56 27.8779
R36 vcm.n698 vcm.t30 27.8779
R37 vcm.n622 vcm.t55 27.8779
R38 vcm.n681 vcm.t51 27.8779
R39 vcm.n907 vcm.t12 27.8779
R40 vcm.n738 vcm.t76 27.8779
R41 vcm.n813 vcm.t64 27.8779
R42 vcm.n963 vcm.t83 27.8779
R43 vcm.n1082 vcm.t42 27.8779
R44 vcm.n1071 vcm.t29 27.8779
R45 vcm.n1170 vcm.t20 27.8779
R46 vcm.n1157 vcm.t27 27.8779
R47 vcm.n1135 vcm.t26 27.8779
R48 vcm.n777 vcm.t80 27.8779
R49 vcm.n837 vcm.t78 27.8779
R50 vcm.n992 vcm.t87 27.8779
R51 vcm.n1052 vcm.t50 27.8779
R52 vcm.n39 vcm.t21 27.8779
R53 vcm.n652 vcm.t48 27.8769
R54 vcm.n464 vcm.t28 27.8769
R55 vcm.n480 vcm.t31 27.8769
R56 vcm.n423 vcm.t37 27.8769
R57 vcm.n308 vcm.t79 27.8769
R58 vcm.n330 vcm.t84 27.8769
R59 vcm.n401 vcm.t35 27.8769
R60 vcm.n549 vcm.t66 27.8769
R61 vcm.n706 vcm.t43 27.8769
R62 vcm.n630 vcm.t47 27.8769
R63 vcm.n689 vcm.t40 27.8769
R64 vcm.n608 vcm.t62 27.8769
R65 vcm.n785 vcm.t75 27.8769
R66 vcm.n1090 vcm.t32 27.8769
R67 vcm.n935 vcm.t11 27.8769
R68 vcm.n943 vcm.t19 27.8769
R69 vcm.n845 vcm.t69 27.8769
R70 vcm.n873 vcm.t71 27.8769
R71 vcm.n1000 vcm.t81 27.8769
R72 vcm.n1011 vcm.t9 27.8769
R73 vcm.n1060 vcm.t39 27.8769
R74 vcm.n1124 vcm.t34 27.8769
R75 vcm.n1146 vcm.t18 27.8769
R76 vcm.n768 vcm.t85 27.8769
R77 vcm.n1182 vcm.t10 27.8769
R78 vcm.n97 vcm.t53 27.8769
R79 vcm.n85 vcm.t8 27.8769
R80 vcm.n51 vcm.t52 27.8769
R81 vcm.n196 vcm.t77 27.8769
R82 vcm.n254 vcm.t13 27.8769
R83 vcm.n456 vcm.t38 27.8769
R84 vcm.n319 vcm.t49 27.8759
R85 vcm.n793 vcm.t82 27.8759
R86 vcm.n859 vcm.t63 27.8759
R87 vcm.n927 vcm.t17 27.8759
R88 vcm.n981 vcm.t14 27.8759
R89 vcm.n757 vcm.n756 22.9652
R90 vcm.n754 vcm.n753 21.2119
R91 vcm.n758 vcm.n754 8.17828
R92 vcm.n758 vcm.n757 6.99309
R93 vcm.n11 vcm 2.29217
R94 vcm.n915 vcm 2.29217
R95 vcm.n560 vcm 2.29217
R96 vcm.n290 vcm 2.29217
R97 vcm.n363 vcm 2.29217
R98 vcm.n426 vcm 2.29217
R99 vcm.n147 vcm 2.29217
R100 vcm.n265 vcm 2.29217
R101 vcm.n155 vcm 2.29217
R102 vcm.n214 vcm 2.29217
R103 vcm.n282 vcm 2.29217
R104 vcm.n452 vcm 2.29217
R105 vcm.n509 vcm 2.29217
R106 vcm.n598 vcm 2.29217
R107 vcm.n673 vcm 2.29217
R108 vcm.n887 vcm 2.29217
R109 vcm.n1117 vcm 2.29217
R110 vcm.n748 vcm 2.29217
R111 vcm.n827 vcm 2.29217
R112 vcm.n974 vcm 2.29217
R113 vcm.n1045 vcm 2.29217
R114 vcm.n17 vcm 2.29217
R115 vcm.n718 vcm.n717 1.63383
R116 vcm.n761 vcm.n759 1.59065
R117 vcm.n1024 vcm.n962 1.58855
R118 vcm.n118 vcm.n101 1.57342
R119 vcm.n93 vcm.n89 1.57342
R120 vcm.n60 vcm.n55 1.57342
R121 vcm.n26 vcm.n12 1.57342
R122 vcm.n925 vcm.n924 1.57342
R123 vcm.n917 vcm.n916 1.57342
R124 vcm.n651 vcm.n650 1.57342
R125 vcm.n547 vcm.n543 1.57342
R126 vcm.n295 vcm.n291 1.57342
R127 vcm.n385 vcm.n378 1.57342
R128 vcm.n371 vcm.n364 1.57342
R129 vcm.n372 vcm.n371 1.57342
R130 vcm.n471 vcm.n470 1.57342
R131 vcm.n489 vcm.n486 1.57342
R132 vcm.n486 vcm.n485 1.57342
R133 vcm.n479 vcm.n478 1.57342
R134 vcm.n422 vcm.n421 1.57342
R135 vcm.n266 vcm.n263 1.57342
R136 vcm.n263 vcm.n259 1.57342
R137 vcm.n185 vcm.n183 1.57342
R138 vcm.n158 vcm.n156 1.57342
R139 vcm.n231 vcm.n230 1.57342
R140 vcm.n241 vcm.n237 1.57342
R141 vcm.n230 vcm.n226 1.57342
R142 vcm.n219 vcm.n215 1.57342
R143 vcm.n220 vcm.n219 1.57342
R144 vcm.n159 vcm.n158 1.57342
R145 vcm.n167 vcm.n165 1.57342
R146 vcm.n168 vcm.n167 1.57342
R147 vcm.n176 vcm.n174 1.57342
R148 vcm.n177 vcm.n176 1.57342
R149 vcm.n242 vcm.n241 1.57342
R150 vcm.n252 vcm.n248 1.57342
R151 vcm.n253 vcm.n252 1.57342
R152 vcm.n186 vcm.n185 1.57342
R153 vcm.n194 vcm.n192 1.57342
R154 vcm.n195 vcm.n194 1.57342
R155 vcm.n328 vcm.n324 1.57342
R156 vcm.n317 vcm.n313 1.57342
R157 vcm.n318 vcm.n317 1.57342
R158 vcm.n329 vcm.n328 1.57342
R159 vcm.n339 vcm.n335 1.57342
R160 vcm.n340 vcm.n339 1.57342
R161 vcm.n421 vcm.n420 1.57342
R162 vcm.n413 vcm.n406 1.57342
R163 vcm.n414 vcm.n413 1.57342
R164 vcm.n478 vcm.n477 1.57342
R165 vcm.n470 vcm.n469 1.57342
R166 vcm.n463 vcm.n462 1.57342
R167 vcm.n462 vcm.n461 1.57342
R168 vcm.n454 vcm.n453 1.57342
R169 vcm.n455 vcm.n454 1.57342
R170 vcm.n526 vcm.n525 1.57342
R171 vcm.n536 vcm.n532 1.57342
R172 vcm.n525 vcm.n521 1.57342
R173 vcm.n514 vcm.n510 1.57342
R174 vcm.n515 vcm.n514 1.57342
R175 vcm.n296 vcm.n295 1.57342
R176 vcm.n306 vcm.n302 1.57342
R177 vcm.n307 vcm.n306 1.57342
R178 vcm.n386 vcm.n385 1.57342
R179 vcm.n399 vcm.n392 1.57342
R180 vcm.n400 vcm.n399 1.57342
R181 vcm.n537 vcm.n536 1.57342
R182 vcm.n548 vcm.n547 1.57342
R183 vcm.n558 vcm.n554 1.57342
R184 vcm.n559 vcm.n558 1.57342
R185 vcm.n705 vcm.n704 1.57342
R186 vcm.n713 vcm.n711 1.57342
R187 vcm.n714 vcm.n713 1.57342
R188 vcm.n650 vcm.n649 1.57342
R189 vcm.n629 vcm.n628 1.57342
R190 vcm.n642 vcm.n635 1.57342
R191 vcm.n643 vcm.n642 1.57342
R192 vcm.n704 vcm.n703 1.57342
R193 vcm.n688 vcm.n687 1.57342
R194 vcm.n696 vcm.n694 1.57342
R195 vcm.n697 vcm.n696 1.57342
R196 vcm.n628 vcm.n627 1.57342
R197 vcm.n606 vcm.n599 1.57342
R198 vcm.n607 vcm.n606 1.57342
R199 vcm.n620 vcm.n613 1.57342
R200 vcm.n621 vcm.n620 1.57342
R201 vcm.n687 vcm.n686 1.57342
R202 vcm.n679 vcm.n674 1.57342
R203 vcm.n680 vcm.n679 1.57342
R204 vcm.n1089 vcm.n1088 1.57342
R205 vcm.n941 vcm.n940 1.57342
R206 vcm.n942 vcm.n941 1.57342
R207 vcm.n949 vcm.n948 1.57342
R208 vcm.n950 vcm.n949 1.57342
R209 vcm.n792 vcm.n791 1.57342
R210 vcm.n800 vcm.n798 1.57342
R211 vcm.n801 vcm.n800 1.57342
R212 vcm.n871 vcm.n864 1.57342
R213 vcm.n857 vcm.n850 1.57342
R214 vcm.n844 vcm.n843 1.57342
R215 vcm.n858 vcm.n857 1.57342
R216 vcm.n872 vcm.n871 1.57342
R217 vcm.n885 vcm.n878 1.57342
R218 vcm.n886 vcm.n885 1.57342
R219 vcm.n1009 vcm.n1005 1.57342
R220 vcm.n999 vcm.n998 1.57342
R221 vcm.n1010 vcm.n1009 1.57342
R222 vcm.n1020 vcm.n1016 1.57342
R223 vcm.n1021 vcm.n1020 1.57342
R224 vcm.n1088 vcm.n1087 1.57342
R225 vcm.n1059 vcm.n1058 1.57342
R226 vcm.n1069 vcm.n1065 1.57342
R227 vcm.n1070 vcm.n1069 1.57342
R228 vcm.n1080 vcm.n1076 1.57342
R229 vcm.n1081 vcm.n1080 1.57342
R230 vcm.n1169 vcm.n1166 1.57342
R231 vcm.n1166 vcm.n1162 1.57342
R232 vcm.n1144 vcm.n1140 1.57342
R233 vcm.n1122 vcm.n1118 1.57342
R234 vcm.n1123 vcm.n1122 1.57342
R235 vcm.n1133 vcm.n1129 1.57342
R236 vcm.n1134 vcm.n1133 1.57342
R237 vcm.n1145 vcm.n1144 1.57342
R238 vcm.n1155 vcm.n1151 1.57342
R239 vcm.n1156 vcm.n1155 1.57342
R240 vcm.n791 vcm.n790 1.57342
R241 vcm.n784 vcm.n783 1.57342
R242 vcm.n783 vcm.n782 1.57342
R243 vcm.n766 vcm.n749 1.57342
R244 vcm.n767 vcm.n766 1.57342
R245 vcm.n775 vcm.n773 1.57342
R246 vcm.n776 vcm.n775 1.57342
R247 vcm.n843 vcm.n842 1.57342
R248 vcm.n835 vcm.n828 1.57342
R249 vcm.n836 vcm.n835 1.57342
R250 vcm.n918 vcm.n917 1.57342
R251 vcm.n926 vcm.n925 1.57342
R252 vcm.n933 vcm.n932 1.57342
R253 vcm.n934 vcm.n933 1.57342
R254 vcm.n998 vcm.n997 1.57342
R255 vcm.n979 vcm.n975 1.57342
R256 vcm.n980 vcm.n979 1.57342
R257 vcm.n990 vcm.n986 1.57342
R258 vcm.n991 vcm.n990 1.57342
R259 vcm.n1058 vcm.n1057 1.57342
R260 vcm.n1050 vcm.n1046 1.57342
R261 vcm.n1051 vcm.n1050 1.57342
R262 vcm.n47 vcm.n43 1.57342
R263 vcm.n22 vcm.n18 1.57342
R264 vcm.n27 vcm.n26 1.57342
R265 vcm.n49 vcm.n32 1.57342
R266 vcm.n50 vcm.n49 1.57342
R267 vcm.n83 vcm.n79 1.57342
R268 vcm.n84 vcm.n83 1.57342
R269 vcm.n61 vcm.n60 1.57342
R270 vcm.n95 vcm.n66 1.57342
R271 vcm.n96 vcm.n95 1.57342
R272 vcm.n114 vcm.n110 1.57342
R273 vcm.n121 vcm.n118 1.57342
R274 vcm.n1024 vcm.n1023 1.49217
R275 vcm.n718 vcm.n716 1.44689
R276 vcm.n953 vcm.n952 1.42133
R277 vcm.n492 vcm.n491 1.4005
R278 vcm.n1186 vcm.n1185 1.388
R279 vcm.n1197 vcm.n1196 1.388
R280 vcm.n1185 vcm 1.14633
R281 vcm.n655 vcm 1.14633
R282 vcm.n491 vcm 1.14633
R283 vcm.n717 vcm 1.14633
R284 vcm.n1030 vcm 1.14633
R285 vcm.n952 vcm 1.14633
R286 vcm.n803 vcm 1.14633
R287 vcm.n1023 vcm 1.14633
R288 vcm.n1167 vcm 1.14633
R289 vcm vcm.n1197 1.14633
R290 vcm.n158 vcm.n157 1.1065
R291 vcm.n167 vcm.n166 1.1065
R292 vcm.n176 vcm.n175 1.1065
R293 vcm.n185 vcm.n184 1.1065
R294 vcm.n194 vcm.n193 1.1065
R295 vcm.n800 vcm.n799 1.1065
R296 vcm.n791 vcm.n740 1.1065
R297 vcm.n783 vcm.n742 1.1065
R298 vcm.n775 vcm.n774 1.1065
R299 vcm.n713 vcm.n712 1.101
R300 vcm.n704 vcm.n665 1.101
R301 vcm.n696 vcm.n695 1.101
R302 vcm.n687 vcm.n668 1.101
R303 vcm.n26 vcm.n13 1.101
R304 vcm.n49 vcm.n33 1.101
R305 vcm.n60 vcm.n56 1.101
R306 vcm.n95 vcm.n67 1.101
R307 vcm.n118 vcm.n102 1.101
R308 vcm.n219 vcm.n218 1.1005
R309 vcm.n241 vcm.n240 1.1005
R310 vcm.n252 vcm.n251 1.1005
R311 vcm.n339 vcm.n338 1.1005
R312 vcm.n263 vcm.n262 1.1005
R313 vcm.n421 vcm.n352 1.1005
R314 vcm.n421 vcm.n355 1.1005
R315 vcm.n413 vcm.n409 1.1005
R316 vcm.n413 vcm.n412 1.1005
R317 vcm.n328 vcm.n327 1.1005
R318 vcm.n514 vcm.n513 1.1005
R319 vcm.n371 vcm.n367 1.1005
R320 vcm.n371 vcm.n370 1.1005
R321 vcm.n295 vcm.n294 1.1005
R322 vcm.n306 vcm.n305 1.1005
R323 vcm.n230 vcm.n229 1.1005
R324 vcm.n385 vcm.n381 1.1005
R325 vcm.n385 vcm.n384 1.1005
R326 vcm.n399 vcm.n395 1.1005
R327 vcm.n399 vcm.n398 1.1005
R328 vcm.n317 vcm.n316 1.1005
R329 vcm.n536 vcm.n535 1.1005
R330 vcm.n558 vcm.n557 1.1005
R331 vcm.n650 vcm.n581 1.1005
R332 vcm.n650 vcm.n584 1.1005
R333 vcm.n642 vcm.n638 1.1005
R334 vcm.n642 vcm.n641 1.1005
R335 vcm.n547 vcm.n546 1.1005
R336 vcm.n628 vcm.n589 1.1005
R337 vcm.n628 vcm.n592 1.1005
R338 vcm.n620 vcm.n616 1.1005
R339 vcm.n620 vcm.n619 1.1005
R340 vcm.n525 vcm.n524 1.1005
R341 vcm.n679 vcm.n678 1.1005
R342 vcm.n606 vcm.n602 1.1005
R343 vcm.n606 vcm.n605 1.1005
R344 vcm.n885 vcm.n881 1.1005
R345 vcm.n885 vcm.n884 1.1005
R346 vcm.n1020 vcm.n1019 1.1005
R347 vcm.n1088 vcm.n1034 1.1005
R348 vcm.n1069 vcm.n1068 1.1005
R349 vcm.n1133 vcm.n1132 1.1005
R350 vcm.n1155 vcm.n1154 1.1005
R351 vcm.n1080 vcm.n1079 1.1005
R352 vcm.n1009 vcm.n1008 1.1005
R353 vcm.n871 vcm.n867 1.1005
R354 vcm.n871 vcm.n870 1.1005
R355 vcm.n843 vcm.n819 1.1005
R356 vcm.n843 vcm.n822 1.1005
R357 vcm.n835 vcm.n831 1.1005
R358 vcm.n835 vcm.n834 1.1005
R359 vcm.n766 vcm.n765 1.1005
R360 vcm.n857 vcm.n853 1.1005
R361 vcm.n857 vcm.n856 1.1005
R362 vcm.n998 vcm.n968 1.1005
R363 vcm.n990 vcm.n989 1.1005
R364 vcm.n1058 vcm.n1040 1.1005
R365 vcm.n1050 vcm.n1049 1.1005
R366 vcm.n979 vcm.n978 1.1005
R367 vcm.n25 vcm.n22 1.1005
R368 vcm.n22 vcm.n21 1.1005
R369 vcm.n1122 vcm.n1121 1.1005
R370 vcm.n26 vcm.n25 1.1005
R371 vcm.n49 vcm.n48 1.1005
R372 vcm.n48 vcm.n47 1.1005
R373 vcm.n47 vcm.n46 1.1005
R374 vcm.n83 vcm.n82 1.1005
R375 vcm.n1144 vcm.n1143 1.1005
R376 vcm.n60 vcm.n59 1.1005
R377 vcm.n95 vcm.n94 1.1005
R378 vcm.n94 vcm.n93 1.1005
R379 vcm.n93 vcm.n92 1.1005
R380 vcm.n117 vcm.n114 1.1005
R381 vcm.n114 vcm.n113 1.1005
R382 vcm.n1166 vcm.n1165 1.1005
R383 vcm.n118 vcm.n117 1.1005
R384 vcm.n731 vcm.n730 1.05236
R385 vcm.n427 vcm.n426 1.013
R386 vcm.n656 vcm.n655 0.971333
R387 vcm.n656 vcm.n653 0.9255
R388 vcm.n427 vcm.n424 0.921888
R389 vcm.n198 vcm.n197 0.822638
R390 vcm.n269 vcm.n268 0.821888
R391 vcm.n730 vcm.n729 0.78775
R392 vcm.n343 vcm.n342 0.771888
R393 vcm.n561 vcm.n560 0.7005
R394 vcm.n804 vcm.n803 0.6755
R395 vcm.n888 vcm.n887 0.604667
R396 vcm.n756 vcm.n755 0.572017
R397 vcm.n1092 vcm.n1091 0.567167
R398 vcm.n1172 vcm.n1171 0.563
R399 vcm.n753 vcm.n752 0.562674
R400 vcm.n1187 vcm.n1186 0.539716
R401 vcm.n657 vcm.n656 0.539716
R402 vcm.n562 vcm.n561 0.539716
R403 vcm.n493 vcm.n492 0.539716
R404 vcm.n428 vcm.n427 0.539716
R405 vcm.n199 vcm.n198 0.539716
R406 vcm.n270 vcm.n269 0.539716
R407 vcm.n344 vcm.n343 0.539716
R408 vcm.n719 vcm.n718 0.539716
R409 vcm.n1093 vcm.n1092 0.539716
R410 vcm.n954 vcm.n953 0.539716
R411 vcm.n805 vcm.n804 0.539716
R412 vcm.n889 vcm.n888 0.539716
R413 vcm.n1025 vcm.n1024 0.539716
R414 vcm.n1173 vcm.n1172 0.539716
R415 vcm.n1196 vcm.n1195 0.539716
R416 vcm.n810 vcm.n809 0.48695
R417 vcm.n662 vcm.n661 0.475318
R418 vcm.n498 vcm.n497 0.469208
R419 vcm.n959 vcm.n958 0.458633
R420 vcm.n1178 vcm.n1177 0.458162
R421 vcm.n275 vcm.n274 0.458045
R422 vcm.n1104 vcm.n1103 0.456753
R423 vcm.n1192 vcm.n1191 0.456635
R424 vcm.n204 vcm.n203 0.456635
R425 vcm.n349 vcm.n348 0.452405
R426 vcm.n1096 vcm.n1029 0.452052
R427 vcm.n900 vcm.n899 0.447353
R428 vcm.n439 vcm.n438 0.43525
R429 vcm.n573 vcm.n572 0.43196
R430 vcm vcm.n98 0.3755
R431 vcm vcm.n86 0.3755
R432 vcm vcm.n52 0.3755
R433 vcm vcm.n374 0.3755
R434 vcm vcm.n481 0.3755
R435 vcm vcm.n255 0.3755
R436 vcm vcm.n179 0.3755
R437 vcm vcm.n233 0.3755
R438 vcm vcm.n222 0.3755
R439 vcm vcm.n161 0.3755
R440 vcm vcm.n170 0.3755
R441 vcm vcm.n244 0.3755
R442 vcm vcm.n188 0.3755
R443 vcm vcm.n309 0.3755
R444 vcm vcm.n320 0.3755
R445 vcm vcm.n331 0.3755
R446 vcm vcm.n416 0.3755
R447 vcm vcm.n402 0.3755
R448 vcm vcm.n473 0.3755
R449 vcm vcm.n465 0.3755
R450 vcm vcm.n457 0.3755
R451 vcm vcm.n528 0.3755
R452 vcm vcm.n517 0.3755
R453 vcm vcm.n298 0.3755
R454 vcm vcm.n388 0.3755
R455 vcm vcm.n539 0.3755
R456 vcm vcm.n550 0.3755
R457 vcm vcm.n707 0.3755
R458 vcm vcm.n645 0.3755
R459 vcm vcm.n631 0.3755
R460 vcm vcm.n699 0.3755
R461 vcm vcm.n690 0.3755
R462 vcm vcm.n623 0.3755
R463 vcm vcm.n609 0.3755
R464 vcm vcm.n682 0.3755
R465 vcm vcm.n936 0.3755
R466 vcm vcm.n944 0.3755
R467 vcm vcm.n794 0.3755
R468 vcm vcm.n846 0.3755
R469 vcm vcm.n860 0.3755
R470 vcm vcm.n874 0.3755
R471 vcm vcm.n1001 0.3755
R472 vcm vcm.n1012 0.3755
R473 vcm vcm.n1083 0.3755
R474 vcm vcm.n1061 0.3755
R475 vcm vcm.n1072 0.3755
R476 vcm vcm.n1158 0.3755
R477 vcm vcm.n1125 0.3755
R478 vcm vcm.n1136 0.3755
R479 vcm vcm.n1147 0.3755
R480 vcm vcm.n786 0.3755
R481 vcm vcm.n778 0.3755
R482 vcm vcm.n769 0.3755
R483 vcm vcm.n838 0.3755
R484 vcm vcm.n920 0.3755
R485 vcm vcm.n928 0.3755
R486 vcm vcm.n993 0.3755
R487 vcm vcm.n982 0.3755
R488 vcm vcm.n1053 0.3755
R489 vcm vcm.n40 0.3755
R490 vcm vcm.n29 0.3755
R491 vcm vcm.n76 0.3755
R492 vcm vcm.n63 0.3755
R493 vcm vcm.n107 0.3755
R494 vcm.n8 vcm 0.234474
R495 vcm.n912 vcm 0.234474
R496 vcm.n653 vcm 0.234474
R497 vcm.n287 vcm 0.234474
R498 vcm.n360 vcm 0.234474
R499 vcm.n152 vcm 0.234474
R500 vcm.n211 vcm 0.234474
R501 vcm.n449 vcm 0.234474
R502 vcm.n506 vcm 0.234474
R503 vcm.n595 vcm 0.234474
R504 vcm.n670 vcm 0.234474
R505 vcm.n1091 vcm 0.234474
R506 vcm.n737 vcm 0.234474
R507 vcm.n1171 vcm 0.234474
R508 vcm.n1114 vcm 0.234474
R509 vcm.n745 vcm 0.234474
R510 vcm.n824 vcm 0.234474
R511 vcm.n971 vcm 0.234474
R512 vcm.n1042 vcm 0.234474
R513 vcm.n14 vcm 0.234474
R514 vcm.n665 vcm 0.187646
R515 vcm.n668 vcm 0.187646
R516 vcm.n13 vcm 0.187646
R517 vcm.n56 vcm 0.187646
R518 vcm.n102 vcm 0.187646
R519 vcm.n712 vcm 0.186894
R520 vcm.n695 vcm 0.186894
R521 vcm.n33 vcm 0.186894
R522 vcm.n67 vcm 0.186894
R523 vcm.n157 vcm 0.185131
R524 vcm.n166 vcm 0.185131
R525 vcm.n184 vcm 0.185131
R526 vcm.n799 vcm 0.185131
R527 vcm.n740 vcm 0.185131
R528 vcm.n742 vcm 0.185131
R529 vcm.n175 vcm 0.185131
R530 vcm.n193 vcm 0.185131
R531 vcm.n774 vcm 0.185131
R532 vcm.n98 vcm 0.117487
R533 vcm.n86 vcm 0.117487
R534 vcm.n52 vcm 0.117487
R535 vcm.n374 vcm 0.117487
R536 vcm.n481 vcm 0.117487
R537 vcm.n255 vcm 0.117487
R538 vcm.n179 vcm 0.117487
R539 vcm.n233 vcm 0.117487
R540 vcm.n222 vcm 0.117487
R541 vcm.n161 vcm 0.117487
R542 vcm.n170 vcm 0.117487
R543 vcm.n244 vcm 0.117487
R544 vcm.n188 vcm 0.117487
R545 vcm.n309 vcm 0.117487
R546 vcm.n320 vcm 0.117487
R547 vcm.n331 vcm 0.117487
R548 vcm.n416 vcm 0.117487
R549 vcm.n402 vcm 0.117487
R550 vcm.n473 vcm 0.117487
R551 vcm.n465 vcm 0.117487
R552 vcm.n457 vcm 0.117487
R553 vcm.n528 vcm 0.117487
R554 vcm.n517 vcm 0.117487
R555 vcm.n298 vcm 0.117487
R556 vcm.n388 vcm 0.117487
R557 vcm.n539 vcm 0.117487
R558 vcm.n550 vcm 0.117487
R559 vcm.n707 vcm 0.117487
R560 vcm.n645 vcm 0.117487
R561 vcm.n631 vcm 0.117487
R562 vcm.n699 vcm 0.117487
R563 vcm.n690 vcm 0.117487
R564 vcm.n623 vcm 0.117487
R565 vcm.n609 vcm 0.117487
R566 vcm.n682 vcm 0.117487
R567 vcm.n936 vcm 0.117487
R568 vcm.n944 vcm 0.117487
R569 vcm.n794 vcm 0.117487
R570 vcm.n846 vcm 0.117487
R571 vcm.n860 vcm 0.117487
R572 vcm.n874 vcm 0.117487
R573 vcm.n1001 vcm 0.117487
R574 vcm.n1012 vcm 0.117487
R575 vcm.n1083 vcm 0.117487
R576 vcm.n1061 vcm 0.117487
R577 vcm.n1072 vcm 0.117487
R578 vcm.n1158 vcm 0.117487
R579 vcm.n1125 vcm 0.117487
R580 vcm.n1136 vcm 0.117487
R581 vcm.n1147 vcm 0.117487
R582 vcm.n786 vcm 0.117487
R583 vcm.n778 vcm 0.117487
R584 vcm.n769 vcm 0.117487
R585 vcm.n838 vcm 0.117487
R586 vcm.n920 vcm 0.117487
R587 vcm.n928 vcm 0.117487
R588 vcm.n993 vcm 0.117487
R589 vcm.n982 vcm 0.117487
R590 vcm.n1053 vcm 0.117487
R591 vcm.n40 vcm 0.117487
R592 vcm.n29 vcm 0.117487
R593 vcm.n76 vcm 0.117487
R594 vcm.n63 vcm 0.117487
R595 vcm.n107 vcm 0.117487
R596 vcm.n10 vcm 0.117222
R597 vcm.n914 vcm 0.117222
R598 vcm.n289 vcm 0.117222
R599 vcm.n362 vcm 0.117222
R600 vcm.n154 vcm 0.117222
R601 vcm.n213 vcm 0.117222
R602 vcm.n451 vcm 0.117222
R603 vcm.n508 vcm 0.117222
R604 vcm.n597 vcm 0.117222
R605 vcm.n672 vcm 0.117222
R606 vcm.n1116 vcm 0.117222
R607 vcm.n747 vcm 0.117222
R608 vcm.n826 vcm 0.117222
R609 vcm.n973 vcm 0.117222
R610 vcm.n1044 vcm 0.117222
R611 vcm.n16 vcm 0.117222
R612 vcm.n499 vcm 0.105191
R613 vcm.n425 vcm 0.105191
R614 vcm.n146 vcm 0.105191
R615 vcm.n264 vcm 0.105191
R616 vcm.n281 vcm 0.105191
R617 vcm.n811 vcm 0.105191
R618 vcm.n261 vcm 0.0970784
R619 vcm.n337 vcm 0.0970784
R620 vcm.n354 vcm 0.0970784
R621 vcm.n411 vcm 0.0970784
R622 vcm.n408 vcm 0.0970784
R623 vcm.n512 vcm 0.0970784
R624 vcm.n397 vcm 0.0970784
R625 vcm.n394 vcm 0.0970784
R626 vcm.n556 vcm 0.0970784
R627 vcm.n583 vcm 0.0970784
R628 vcm.n640 vcm 0.0970784
R629 vcm.n637 vcm 0.0970784
R630 vcm.n591 vcm 0.0970784
R631 vcm.n618 vcm 0.0970784
R632 vcm.n615 vcm 0.0970784
R633 vcm.n601 vcm 0.0970784
R634 vcm.n1078 vcm 0.0970784
R635 vcm.n1007 vcm 0.0970784
R636 vcm.n866 vcm 0.0970784
R637 vcm.n833 vcm 0.0970784
R638 vcm.n830 vcm 0.0970784
R639 vcm.n852 vcm 0.0970784
R640 vcm.n967 vcm 0.0970784
R641 vcm.n988 vcm 0.0970784
R642 vcm.n1039 vcm 0.0970784
R643 vcm.n35 vcm 0.0965779
R644 vcm.n69 vcm 0.0965779
R645 vcm.n326 vcm 0.0965766
R646 vcm.n351 vcm 0.0965766
R647 vcm.n545 vcm 0.0965766
R648 vcm.n604 vcm 0.0965766
R649 vcm.n523 vcm 0.0965766
R650 vcm.n380 vcm 0.0965766
R651 vcm.n534 vcm 0.0965766
R652 vcm.n580 vcm 0.0965766
R653 vcm.n588 vcm 0.0965766
R654 vcm.n1153 vcm 0.0965766
R655 vcm.n869 vcm 0.0965766
R656 vcm.n977 vcm 0.0965766
R657 vcm.n1142 vcm 0.0965766
R658 vcm.n1067 vcm 0.0965766
R659 vcm.n1131 vcm 0.0965766
R660 vcm.n217 vcm 0.0958266
R661 vcm.n228 vcm 0.0958266
R662 vcm.n315 vcm 0.0958266
R663 vcm.n250 vcm 0.0958266
R664 vcm.n366 vcm 0.0958266
R665 vcm.n369 vcm 0.0958266
R666 vcm.n304 vcm 0.0958266
R667 vcm.n883 vcm 0.0958266
R668 vcm.n1018 vcm 0.0958266
R669 vcm.n1164 vcm 0.0958266
R670 vcm.n855 vcm 0.0958266
R671 vcm.n818 vcm 0.0958266
R672 vcm.n1048 vcm 0.0958266
R673 vcm.n20 vcm 0.0958266
R674 vcm.n81 vcm 0.0958266
R675 vcm.n112 vcm 0.0958266
R676 vcm.n239 vcm 0.0956149
R677 vcm.n293 vcm 0.0956149
R678 vcm.n383 vcm 0.0956149
R679 vcm.n880 vcm 0.0956149
R680 vcm.n1033 vcm 0.0956149
R681 vcm.n821 vcm 0.0956149
R682 vcm.n1120 vcm 0.0956149
R683 vcm.n24 vcm 0.0956149
R684 vcm.n45 vcm 0.0956149
R685 vcm.n58 vcm 0.0956149
R686 vcm.n91 vcm 0.0956149
R687 vcm.n116 vcm 0.0956149
R688 vcm.n677 vcm.n676 0.0955985
R689 vcm.n1184 vcm.n1183 0.0915799
R690 vcm.n490 vcm.n489 0.0915799
R691 vcm.n714 vcm.n663 0.0915799
R692 vcm.n1089 vcm.n1031 0.0915799
R693 vcm.n951 vcm.n950 0.0915799
R694 vcm.n802 vcm.n801 0.0915799
R695 vcm.n1022 vcm.n1021 0.0915799
R696 vcm.n1169 vcm.n1168 0.0915799
R697 vcm.n122 vcm.n121 0.0915799
R698 vcm.n101 vcm.n100 0.0914585
R699 vcm.n89 vcm.n88 0.0914585
R700 vcm.n55 vcm.n54 0.0914585
R701 vcm.n378 vcm.n377 0.0914585
R702 vcm.n485 vcm.n484 0.0914585
R703 vcm.n259 vcm.n258 0.0914585
R704 vcm.n183 vcm.n182 0.0914585
R705 vcm.n237 vcm.n236 0.0914585
R706 vcm.n226 vcm.n225 0.0914585
R707 vcm.n165 vcm.n164 0.0914585
R708 vcm.n174 vcm.n173 0.0914585
R709 vcm.n248 vcm.n247 0.0914585
R710 vcm.n192 vcm.n191 0.0914585
R711 vcm.n313 vcm.n312 0.0914585
R712 vcm.n324 vcm.n323 0.0914585
R713 vcm.n335 vcm.n334 0.0914585
R714 vcm.n420 vcm.n419 0.0914585
R715 vcm.n406 vcm.n405 0.0914585
R716 vcm.n477 vcm.n476 0.0914585
R717 vcm.n469 vcm.n468 0.0914585
R718 vcm.n461 vcm.n460 0.0914585
R719 vcm.n532 vcm.n531 0.0914585
R720 vcm.n521 vcm.n520 0.0914585
R721 vcm.n302 vcm.n301 0.0914585
R722 vcm.n392 vcm.n391 0.0914585
R723 vcm.n543 vcm.n542 0.0914585
R724 vcm.n554 vcm.n553 0.0914585
R725 vcm.n711 vcm.n710 0.0914585
R726 vcm.n649 vcm.n648 0.0914585
R727 vcm.n635 vcm.n634 0.0914585
R728 vcm.n703 vcm.n702 0.0914585
R729 vcm.n694 vcm.n693 0.0914585
R730 vcm.n627 vcm.n626 0.0914585
R731 vcm.n613 vcm.n612 0.0914585
R732 vcm.n686 vcm.n685 0.0914585
R733 vcm.n940 vcm.n939 0.0914585
R734 vcm.n948 vcm.n947 0.0914585
R735 vcm.n798 vcm.n797 0.0914585
R736 vcm.n850 vcm.n849 0.0914585
R737 vcm.n864 vcm.n863 0.0914585
R738 vcm.n878 vcm.n877 0.0914585
R739 vcm.n1005 vcm.n1004 0.0914585
R740 vcm.n1016 vcm.n1015 0.0914585
R741 vcm.n1087 vcm.n1086 0.0914585
R742 vcm.n1065 vcm.n1064 0.0914585
R743 vcm.n1076 vcm.n1075 0.0914585
R744 vcm.n1162 vcm.n1161 0.0914585
R745 vcm.n1129 vcm.n1128 0.0914585
R746 vcm.n1140 vcm.n1139 0.0914585
R747 vcm.n1151 vcm.n1150 0.0914585
R748 vcm.n790 vcm.n789 0.0914585
R749 vcm.n782 vcm.n781 0.0914585
R750 vcm.n773 vcm.n772 0.0914585
R751 vcm.n842 vcm.n841 0.0914585
R752 vcm.n924 vcm.n923 0.0914585
R753 vcm.n932 vcm.n931 0.0914585
R754 vcm.n997 vcm.n996 0.0914585
R755 vcm.n986 vcm.n985 0.0914585
R756 vcm.n1057 vcm.n1056 0.0914585
R757 vcm.n43 vcm.n42 0.0914585
R758 vcm.n32 vcm.n31 0.0914585
R759 vcm.n79 vcm.n78 0.0914585
R760 vcm.n66 vcm.n65 0.0914585
R761 vcm.n110 vcm.n109 0.0914585
R762 vcm.n197 vcm.n196 0.0888628
R763 vcm.n1182 vcm.n1181 0.0888625
R764 vcm.n501 vcm.n500 0.0888625
R765 vcm.n488 vcm.n487 0.0888625
R766 vcm.n424 vcm.n423 0.0888625
R767 vcm.n268 vcm.n267 0.0888625
R768 vcm.n342 vcm.n341 0.0888625
R769 vcm.n716 vcm.n715 0.0888625
R770 vcm.n907 vcm.n906 0.0888625
R771 vcm.n813 vcm.n812 0.0888625
R772 vcm.n120 vcm.n119 0.0888625
R773 vcm.n675 vcm 0.0635002
R774 vcm.n751 vcm 0.063
R775 vcm.n730 vcm 0.0617502
R776 vcm.n12 vcm.n11 0.049413
R777 vcm.n916 vcm.n915 0.049413
R778 vcm.n560 vcm.n559 0.049413
R779 vcm.n291 vcm.n290 0.049413
R780 vcm.n364 vcm.n363 0.049413
R781 vcm.n195 vcm.n147 0.049413
R782 vcm.n266 vcm.n265 0.049413
R783 vcm.n156 vcm.n155 0.049413
R784 vcm.n215 vcm.n214 0.049413
R785 vcm.n340 vcm.n282 0.049413
R786 vcm.n453 vcm.n452 0.049413
R787 vcm.n510 vcm.n509 0.049413
R788 vcm.n599 vcm.n598 0.049413
R789 vcm.n674 vcm.n673 0.049413
R790 vcm.n887 vcm.n886 0.049413
R791 vcm.n1118 vcm.n1117 0.049413
R792 vcm.n749 vcm.n748 0.049413
R793 vcm.n828 vcm.n827 0.049413
R794 vcm.n975 vcm.n974 0.049413
R795 vcm.n1046 vcm.n1045 0.049413
R796 vcm.n18 vcm.n17 0.049413
R797 vcm.n98 vcm.n0 0.0466957
R798 vcm.n98 vcm.n97 0.0466957
R799 vcm.n86 vcm.n70 0.0466957
R800 vcm.n86 vcm.n85 0.0466957
R801 vcm.n52 vcm.n4 0.0466957
R802 vcm.n52 vcm.n51 0.0466957
R803 vcm.n9 vcm.n8 0.0466957
R804 vcm.n913 vcm.n912 0.0466957
R805 vcm.n653 vcm.n652 0.0466957
R806 vcm.n288 vcm.n287 0.0466957
R807 vcm.n374 vcm.n359 0.0466957
R808 vcm.n374 vcm.n373 0.0466957
R809 vcm.n361 vcm.n360 0.0466957
R810 vcm.n481 vcm.n445 0.0466957
R811 vcm.n481 vcm.n480 0.0466957
R812 vcm.n255 vcm.n207 0.0466957
R813 vcm.n255 vcm.n254 0.0466957
R814 vcm.n179 vcm.n149 0.0466957
R815 vcm.n179 vcm.n178 0.0466957
R816 vcm.n153 vcm.n152 0.0466957
R817 vcm.n233 vcm.n209 0.0466957
R818 vcm.n233 vcm.n232 0.0466957
R819 vcm.n222 vcm.n210 0.0466957
R820 vcm.n222 vcm.n221 0.0466957
R821 vcm.n212 vcm.n211 0.0466957
R822 vcm.n161 vcm.n160 0.0466957
R823 vcm.n161 vcm.n151 0.0466957
R824 vcm.n170 vcm.n169 0.0466957
R825 vcm.n170 vcm.n150 0.0466957
R826 vcm.n244 vcm.n243 0.0466957
R827 vcm.n244 vcm.n208 0.0466957
R828 vcm.n188 vcm.n187 0.0466957
R829 vcm.n188 vcm.n148 0.0466957
R830 vcm.n309 vcm.n308 0.0466957
R831 vcm.n309 vcm.n285 0.0466957
R832 vcm.n320 vcm.n319 0.0466957
R833 vcm.n320 vcm.n284 0.0466957
R834 vcm.n331 vcm.n330 0.0466957
R835 vcm.n331 vcm.n283 0.0466957
R836 vcm.n416 vcm.n356 0.0466957
R837 vcm.n416 vcm.n415 0.0466957
R838 vcm.n402 vcm.n401 0.0466957
R839 vcm.n402 vcm.n357 0.0466957
R840 vcm.n473 vcm.n446 0.0466957
R841 vcm.n473 vcm.n472 0.0466957
R842 vcm.n465 vcm.n447 0.0466957
R843 vcm.n465 vcm.n464 0.0466957
R844 vcm.n457 vcm.n448 0.0466957
R845 vcm.n457 vcm.n456 0.0466957
R846 vcm.n450 vcm.n449 0.0466957
R847 vcm.n528 vcm.n504 0.0466957
R848 vcm.n528 vcm.n527 0.0466957
R849 vcm.n517 vcm.n505 0.0466957
R850 vcm.n517 vcm.n516 0.0466957
R851 vcm.n507 vcm.n506 0.0466957
R852 vcm.n298 vcm.n297 0.0466957
R853 vcm.n298 vcm.n286 0.0466957
R854 vcm.n388 vcm.n387 0.0466957
R855 vcm.n388 vcm.n358 0.0466957
R856 vcm.n539 vcm.n538 0.0466957
R857 vcm.n539 vcm.n503 0.0466957
R858 vcm.n550 vcm.n549 0.0466957
R859 vcm.n550 vcm.n502 0.0466957
R860 vcm.n707 vcm.n706 0.0466957
R861 vcm.n707 vcm.n664 0.0466957
R862 vcm.n645 vcm.n585 0.0466957
R863 vcm.n645 vcm.n644 0.0466957
R864 vcm.n631 vcm.n630 0.0466957
R865 vcm.n631 vcm.n586 0.0466957
R866 vcm.n699 vcm.n666 0.0466957
R867 vcm.n699 vcm.n698 0.0466957
R868 vcm.n690 vcm.n689 0.0466957
R869 vcm.n690 vcm.n667 0.0466957
R870 vcm.n623 vcm.n593 0.0466957
R871 vcm.n623 vcm.n622 0.0466957
R872 vcm.n596 vcm.n595 0.0466957
R873 vcm.n609 vcm.n608 0.0466957
R874 vcm.n609 vcm.n594 0.0466957
R875 vcm.n682 vcm.n669 0.0466957
R876 vcm.n682 vcm.n681 0.0466957
R877 vcm.n671 vcm.n670 0.0466957
R878 vcm.n1091 vcm.n1090 0.0466957
R879 vcm.n936 vcm.n935 0.0466957
R880 vcm.n936 vcm.n909 0.0466957
R881 vcm.n944 vcm.n943 0.0466957
R882 vcm.n944 vcm.n908 0.0466957
R883 vcm.n738 vcm.n737 0.0466957
R884 vcm.n794 vcm.n793 0.0466957
R885 vcm.n794 vcm.n739 0.0466957
R886 vcm.n846 vcm.n845 0.0466957
R887 vcm.n846 vcm.n816 0.0466957
R888 vcm.n860 vcm.n859 0.0466957
R889 vcm.n860 vcm.n815 0.0466957
R890 vcm.n874 vcm.n873 0.0466957
R891 vcm.n874 vcm.n814 0.0466957
R892 vcm.n1001 vcm.n1000 0.0466957
R893 vcm.n1001 vcm.n965 0.0466957
R894 vcm.n1012 vcm.n1011 0.0466957
R895 vcm.n1012 vcm.n964 0.0466957
R896 vcm.n1083 vcm.n1035 0.0466957
R897 vcm.n1083 vcm.n1082 0.0466957
R898 vcm.n1061 vcm.n1060 0.0466957
R899 vcm.n1061 vcm.n1037 0.0466957
R900 vcm.n1072 vcm.n1071 0.0466957
R901 vcm.n1072 vcm.n1036 0.0466957
R902 vcm.n1171 vcm.n1170 0.0466957
R903 vcm.n1158 vcm.n1110 0.0466957
R904 vcm.n1158 vcm.n1157 0.0466957
R905 vcm.n1115 vcm.n1114 0.0466957
R906 vcm.n1125 vcm.n1124 0.0466957
R907 vcm.n1125 vcm.n1113 0.0466957
R908 vcm.n1136 vcm.n1135 0.0466957
R909 vcm.n1136 vcm.n1112 0.0466957
R910 vcm.n1147 vcm.n1146 0.0466957
R911 vcm.n1147 vcm.n1111 0.0466957
R912 vcm.n786 vcm.n741 0.0466957
R913 vcm.n786 vcm.n785 0.0466957
R914 vcm.n778 vcm.n743 0.0466957
R915 vcm.n778 vcm.n777 0.0466957
R916 vcm.n746 vcm.n745 0.0466957
R917 vcm.n769 vcm.n768 0.0466957
R918 vcm.n769 vcm.n744 0.0466957
R919 vcm.n838 vcm.n823 0.0466957
R920 vcm.n838 vcm.n837 0.0466957
R921 vcm.n825 vcm.n824 0.0466957
R922 vcm.n920 vcm.n919 0.0466957
R923 vcm.n920 vcm.n911 0.0466957
R924 vcm.n928 vcm.n927 0.0466957
R925 vcm.n928 vcm.n910 0.0466957
R926 vcm.n993 vcm.n969 0.0466957
R927 vcm.n993 vcm.n992 0.0466957
R928 vcm.n972 vcm.n971 0.0466957
R929 vcm.n982 vcm.n981 0.0466957
R930 vcm.n982 vcm.n970 0.0466957
R931 vcm.n1053 vcm.n1041 0.0466957
R932 vcm.n1053 vcm.n1052 0.0466957
R933 vcm.n1043 vcm.n1042 0.0466957
R934 vcm.n40 vcm.n36 0.0466957
R935 vcm.n40 vcm.n39 0.0466957
R936 vcm.n15 vcm.n14 0.0466957
R937 vcm.n29 vcm.n28 0.0466957
R938 vcm.n29 vcm.n6 0.0466957
R939 vcm.n76 vcm.n75 0.0466957
R940 vcm.n76 vcm.n72 0.0466957
R941 vcm.n63 vcm.n62 0.0466957
R942 vcm.n63 vcm.n2 0.0466957
R943 vcm.n107 vcm.n106 0.0466957
R944 vcm.n107 vcm.n103 0.0466957
R945 vcm.n560 vcm.n499 0.0394617
R946 vcm.n426 vcm.n425 0.0394617
R947 vcm.n147 vcm.n146 0.0394617
R948 vcm.n265 vcm.n264 0.0394617
R949 vcm.n282 vcm.n281 0.0394617
R950 vcm.n887 vcm.n811 0.0394617
R951 vcm.n1185 vcm.n1184 0.0385543
R952 vcm.n655 vcm.n654 0.0385543
R953 vcm.n491 vcm.n490 0.0385543
R954 vcm.n1031 vcm.n1030 0.0385543
R955 vcm.n952 vcm.n951 0.0385543
R956 vcm.n803 vcm.n802 0.0385543
R957 vcm.n1023 vcm.n1022 0.0385543
R958 vcm.n1168 vcm.n1167 0.0385543
R959 vcm.n1197 vcm.n122 0.0385543
R960 vcm.n763 vcm.n762 0.0302414
R961 vcm.n11 vcm.n10 0.0270767
R962 vcm.n915 vcm.n914 0.0270767
R963 vcm.n290 vcm.n289 0.0270767
R964 vcm.n363 vcm.n362 0.0270767
R965 vcm.n155 vcm.n154 0.0270767
R966 vcm.n214 vcm.n213 0.0270767
R967 vcm.n452 vcm.n451 0.0270767
R968 vcm.n509 vcm.n508 0.0270767
R969 vcm.n598 vcm.n597 0.0270767
R970 vcm.n673 vcm.n672 0.0270767
R971 vcm.n1117 vcm.n1116 0.0270767
R972 vcm.n748 vcm.n747 0.0270767
R973 vcm.n827 vcm.n826 0.0270767
R974 vcm.n974 vcm.n973 0.0270767
R975 vcm.n1045 vcm.n1044 0.0270767
R976 vcm.n17 vcm.n16 0.0270767
R977 vcm.n100 vcm 0.0209545
R978 vcm.n88 vcm 0.0209545
R979 vcm.n54 vcm 0.0209545
R980 vcm.n377 vcm 0.0209545
R981 vcm.n484 vcm 0.0209545
R982 vcm.n258 vcm 0.0209545
R983 vcm.n182 vcm 0.0209545
R984 vcm.n236 vcm 0.0209545
R985 vcm.n225 vcm 0.0209545
R986 vcm.n164 vcm 0.0209545
R987 vcm.n173 vcm 0.0209545
R988 vcm.n247 vcm 0.0209545
R989 vcm.n191 vcm 0.0209545
R990 vcm.n312 vcm 0.0209545
R991 vcm.n323 vcm 0.0209545
R992 vcm.n334 vcm 0.0209545
R993 vcm.n419 vcm 0.0209545
R994 vcm.n405 vcm 0.0209545
R995 vcm.n476 vcm 0.0209545
R996 vcm.n468 vcm 0.0209545
R997 vcm.n460 vcm 0.0209545
R998 vcm.n531 vcm 0.0209545
R999 vcm.n520 vcm 0.0209545
R1000 vcm.n301 vcm 0.0209545
R1001 vcm.n391 vcm 0.0209545
R1002 vcm.n542 vcm 0.0209545
R1003 vcm.n553 vcm 0.0209545
R1004 vcm.n710 vcm 0.0209545
R1005 vcm.n648 vcm 0.0209545
R1006 vcm.n634 vcm 0.0209545
R1007 vcm.n702 vcm 0.0209545
R1008 vcm.n693 vcm 0.0209545
R1009 vcm.n626 vcm 0.0209545
R1010 vcm.n612 vcm 0.0209545
R1011 vcm.n685 vcm 0.0209545
R1012 vcm.n939 vcm 0.0209545
R1013 vcm.n947 vcm 0.0209545
R1014 vcm.n797 vcm 0.0209545
R1015 vcm.n849 vcm 0.0209545
R1016 vcm.n863 vcm 0.0209545
R1017 vcm.n877 vcm 0.0209545
R1018 vcm.n1004 vcm 0.0209545
R1019 vcm.n1015 vcm 0.0209545
R1020 vcm.n1086 vcm 0.0209545
R1021 vcm.n1064 vcm 0.0209545
R1022 vcm.n1075 vcm 0.0209545
R1023 vcm.n1161 vcm 0.0209545
R1024 vcm.n1128 vcm 0.0209545
R1025 vcm.n1139 vcm 0.0209545
R1026 vcm.n1150 vcm 0.0209545
R1027 vcm.n789 vcm 0.0209545
R1028 vcm.n781 vcm 0.0209545
R1029 vcm.n772 vcm 0.0209545
R1030 vcm.n841 vcm 0.0209545
R1031 vcm.n923 vcm 0.0209545
R1032 vcm.n931 vcm 0.0209545
R1033 vcm.n996 vcm 0.0209545
R1034 vcm.n985 vcm 0.0209545
R1035 vcm.n1056 vcm 0.0209545
R1036 vcm.n42 vcm 0.0209545
R1037 vcm.n31 vcm 0.0209545
R1038 vcm.n78 vcm 0.0209545
R1039 vcm.n65 vcm 0.0209545
R1040 vcm.n109 vcm 0.0209545
R1041 vcm.n762 vcm.n751 0.0197903
R1042 vcm vcm.n99 0.0150455
R1043 vcm vcm.n87 0.0150455
R1044 vcm vcm.n53 0.0150455
R1045 vcm.n375 vcm 0.0150455
R1046 vcm.n482 vcm 0.0150455
R1047 vcm.n256 vcm 0.0150455
R1048 vcm.n180 vcm 0.0150455
R1049 vcm.n234 vcm 0.0150455
R1050 vcm.n223 vcm 0.0150455
R1051 vcm.n162 vcm 0.0150455
R1052 vcm.n171 vcm 0.0150455
R1053 vcm.n245 vcm 0.0150455
R1054 vcm.n189 vcm 0.0150455
R1055 vcm.n310 vcm 0.0150455
R1056 vcm.n321 vcm 0.0150455
R1057 vcm.n332 vcm 0.0150455
R1058 vcm.n417 vcm 0.0150455
R1059 vcm.n403 vcm 0.0150455
R1060 vcm.n474 vcm 0.0150455
R1061 vcm.n466 vcm 0.0150455
R1062 vcm.n458 vcm 0.0150455
R1063 vcm.n529 vcm 0.0150455
R1064 vcm.n518 vcm 0.0150455
R1065 vcm.n299 vcm 0.0150455
R1066 vcm.n389 vcm 0.0150455
R1067 vcm.n540 vcm 0.0150455
R1068 vcm.n551 vcm 0.0150455
R1069 vcm.n708 vcm 0.0150455
R1070 vcm.n646 vcm 0.0150455
R1071 vcm.n632 vcm 0.0150455
R1072 vcm.n700 vcm 0.0150455
R1073 vcm.n691 vcm 0.0150455
R1074 vcm.n624 vcm 0.0150455
R1075 vcm.n610 vcm 0.0150455
R1076 vcm.n683 vcm 0.0150455
R1077 vcm.n937 vcm 0.0150455
R1078 vcm.n945 vcm 0.0150455
R1079 vcm.n795 vcm 0.0150455
R1080 vcm.n847 vcm 0.0150455
R1081 vcm.n861 vcm 0.0150455
R1082 vcm.n875 vcm 0.0150455
R1083 vcm.n1002 vcm 0.0150455
R1084 vcm.n1013 vcm 0.0150455
R1085 vcm.n1084 vcm 0.0150455
R1086 vcm.n1062 vcm 0.0150455
R1087 vcm.n1073 vcm 0.0150455
R1088 vcm.n1159 vcm 0.0150455
R1089 vcm.n1126 vcm 0.0150455
R1090 vcm.n1137 vcm 0.0150455
R1091 vcm.n1148 vcm 0.0150455
R1092 vcm.n787 vcm 0.0150455
R1093 vcm.n779 vcm 0.0150455
R1094 vcm.n770 vcm 0.0150455
R1095 vcm.n839 vcm 0.0150455
R1096 vcm.n921 vcm 0.0150455
R1097 vcm.n929 vcm 0.0150455
R1098 vcm.n994 vcm 0.0150455
R1099 vcm.n983 vcm 0.0150455
R1100 vcm.n1054 vcm 0.0150455
R1101 vcm vcm.n41 0.0150455
R1102 vcm vcm.n30 0.0150455
R1103 vcm vcm.n77 0.0150455
R1104 vcm vcm.n64 0.0150455
R1105 vcm vcm.n108 0.0150455
R1106 vcm.n762 vcm.n761 0.00833208
R1107 vcm.n765 vcm.n764 0.00570833
R1108 vcm.n763 vcm.n750 0.00481034
R1109 vcm.n1183 vcm.n1182 0.00321739
R1110 vcm.n101 vcm.n0 0.00321739
R1111 vcm.n97 vcm.n96 0.00321739
R1112 vcm.n89 vcm.n70 0.00321739
R1113 vcm.n85 vcm.n84 0.00321739
R1114 vcm.n55 vcm.n4 0.00321739
R1115 vcm.n51 vcm.n50 0.00321739
R1116 vcm.n12 vcm.n9 0.00321739
R1117 vcm.n916 vcm.n913 0.00321739
R1118 vcm.n652 vcm.n651 0.00321739
R1119 vcm.n559 vcm.n501 0.00321739
R1120 vcm.n291 vcm.n288 0.00321739
R1121 vcm.n378 vcm.n359 0.00321739
R1122 vcm.n373 vcm.n372 0.00321739
R1123 vcm.n364 vcm.n361 0.00321739
R1124 vcm.n489 vcm.n488 0.00321739
R1125 vcm.n485 vcm.n445 0.00321739
R1126 vcm.n480 vcm.n479 0.00321739
R1127 vcm.n423 vcm.n422 0.00321739
R1128 vcm.n196 vcm.n195 0.00321739
R1129 vcm.n267 vcm.n266 0.00321739
R1130 vcm.n259 vcm.n207 0.00321739
R1131 vcm.n254 vcm.n253 0.00321739
R1132 vcm.n183 vcm.n149 0.00321739
R1133 vcm.n178 vcm.n177 0.00321739
R1134 vcm.n156 vcm.n153 0.00321739
R1135 vcm.n237 vcm.n209 0.00321739
R1136 vcm.n232 vcm.n231 0.00321739
R1137 vcm.n226 vcm.n210 0.00321739
R1138 vcm.n221 vcm.n220 0.00321739
R1139 vcm.n215 vcm.n212 0.00321739
R1140 vcm.n160 vcm.n159 0.00321739
R1141 vcm.n165 vcm.n151 0.00321739
R1142 vcm.n169 vcm.n168 0.00321739
R1143 vcm.n174 vcm.n150 0.00321739
R1144 vcm.n243 vcm.n242 0.00321739
R1145 vcm.n248 vcm.n208 0.00321739
R1146 vcm.n187 vcm.n186 0.00321739
R1147 vcm.n192 vcm.n148 0.00321739
R1148 vcm.n341 vcm.n340 0.00321739
R1149 vcm.n308 vcm.n307 0.00321739
R1150 vcm.n313 vcm.n285 0.00321739
R1151 vcm.n319 vcm.n318 0.00321739
R1152 vcm.n324 vcm.n284 0.00321739
R1153 vcm.n330 vcm.n329 0.00321739
R1154 vcm.n335 vcm.n283 0.00321739
R1155 vcm.n420 vcm.n356 0.00321739
R1156 vcm.n415 vcm.n414 0.00321739
R1157 vcm.n401 vcm.n400 0.00321739
R1158 vcm.n406 vcm.n357 0.00321739
R1159 vcm.n477 vcm.n446 0.00321739
R1160 vcm.n472 vcm.n471 0.00321739
R1161 vcm.n469 vcm.n447 0.00321739
R1162 vcm.n464 vcm.n463 0.00321739
R1163 vcm.n461 vcm.n448 0.00321739
R1164 vcm.n456 vcm.n455 0.00321739
R1165 vcm.n453 vcm.n450 0.00321739
R1166 vcm.n532 vcm.n504 0.00321739
R1167 vcm.n527 vcm.n526 0.00321739
R1168 vcm.n521 vcm.n505 0.00321739
R1169 vcm.n516 vcm.n515 0.00321739
R1170 vcm.n510 vcm.n507 0.00321739
R1171 vcm.n297 vcm.n296 0.00321739
R1172 vcm.n302 vcm.n286 0.00321739
R1173 vcm.n387 vcm.n386 0.00321739
R1174 vcm.n392 vcm.n358 0.00321739
R1175 vcm.n538 vcm.n537 0.00321739
R1176 vcm.n543 vcm.n503 0.00321739
R1177 vcm.n549 vcm.n548 0.00321739
R1178 vcm.n554 vcm.n502 0.00321739
R1179 vcm.n715 vcm.n714 0.00321739
R1180 vcm.n706 vcm.n705 0.00321739
R1181 vcm.n711 vcm.n664 0.00321739
R1182 vcm.n649 vcm.n585 0.00321739
R1183 vcm.n644 vcm.n643 0.00321739
R1184 vcm.n630 vcm.n629 0.00321739
R1185 vcm.n635 vcm.n586 0.00321739
R1186 vcm.n703 vcm.n666 0.00321739
R1187 vcm.n698 vcm.n697 0.00321739
R1188 vcm.n689 vcm.n688 0.00321739
R1189 vcm.n694 vcm.n667 0.00321739
R1190 vcm.n627 vcm.n593 0.00321739
R1191 vcm.n622 vcm.n621 0.00321739
R1192 vcm.n599 vcm.n596 0.00321739
R1193 vcm.n608 vcm.n607 0.00321739
R1194 vcm.n613 vcm.n594 0.00321739
R1195 vcm.n686 vcm.n669 0.00321739
R1196 vcm.n681 vcm.n680 0.00321739
R1197 vcm.n674 vcm.n671 0.00321739
R1198 vcm.n1090 vcm.n1089 0.00321739
R1199 vcm.n950 vcm.n907 0.00321739
R1200 vcm.n935 vcm.n934 0.00321739
R1201 vcm.n940 vcm.n909 0.00321739
R1202 vcm.n943 vcm.n942 0.00321739
R1203 vcm.n948 vcm.n908 0.00321739
R1204 vcm.n801 vcm.n738 0.00321739
R1205 vcm.n793 vcm.n792 0.00321739
R1206 vcm.n798 vcm.n739 0.00321739
R1207 vcm.n886 vcm.n813 0.00321739
R1208 vcm.n845 vcm.n844 0.00321739
R1209 vcm.n850 vcm.n816 0.00321739
R1210 vcm.n859 vcm.n858 0.00321739
R1211 vcm.n864 vcm.n815 0.00321739
R1212 vcm.n873 vcm.n872 0.00321739
R1213 vcm.n878 vcm.n814 0.00321739
R1214 vcm.n1021 vcm.n963 0.00321739
R1215 vcm.n1000 vcm.n999 0.00321739
R1216 vcm.n1005 vcm.n965 0.00321739
R1217 vcm.n1011 vcm.n1010 0.00321739
R1218 vcm.n1016 vcm.n964 0.00321739
R1219 vcm.n1087 vcm.n1035 0.00321739
R1220 vcm.n1082 vcm.n1081 0.00321739
R1221 vcm.n1060 vcm.n1059 0.00321739
R1222 vcm.n1065 vcm.n1037 0.00321739
R1223 vcm.n1071 vcm.n1070 0.00321739
R1224 vcm.n1076 vcm.n1036 0.00321739
R1225 vcm.n1170 vcm.n1169 0.00321739
R1226 vcm.n1162 vcm.n1110 0.00321739
R1227 vcm.n1157 vcm.n1156 0.00321739
R1228 vcm.n1118 vcm.n1115 0.00321739
R1229 vcm.n1124 vcm.n1123 0.00321739
R1230 vcm.n1129 vcm.n1113 0.00321739
R1231 vcm.n1135 vcm.n1134 0.00321739
R1232 vcm.n1140 vcm.n1112 0.00321739
R1233 vcm.n1146 vcm.n1145 0.00321739
R1234 vcm.n1151 vcm.n1111 0.00321739
R1235 vcm.n790 vcm.n741 0.00321739
R1236 vcm.n785 vcm.n784 0.00321739
R1237 vcm.n782 vcm.n743 0.00321739
R1238 vcm.n777 vcm.n776 0.00321739
R1239 vcm.n749 vcm.n746 0.00321739
R1240 vcm.n768 vcm.n767 0.00321739
R1241 vcm.n773 vcm.n744 0.00321739
R1242 vcm.n842 vcm.n823 0.00321739
R1243 vcm.n837 vcm.n836 0.00321739
R1244 vcm.n828 vcm.n825 0.00321739
R1245 vcm.n919 vcm.n918 0.00321739
R1246 vcm.n924 vcm.n911 0.00321739
R1247 vcm.n927 vcm.n926 0.00321739
R1248 vcm.n932 vcm.n910 0.00321739
R1249 vcm.n997 vcm.n969 0.00321739
R1250 vcm.n992 vcm.n991 0.00321739
R1251 vcm.n975 vcm.n972 0.00321739
R1252 vcm.n981 vcm.n980 0.00321739
R1253 vcm.n986 vcm.n970 0.00321739
R1254 vcm.n1057 vcm.n1041 0.00321739
R1255 vcm.n1052 vcm.n1051 0.00321739
R1256 vcm.n1046 vcm.n1043 0.00321739
R1257 vcm.n43 vcm.n36 0.00321739
R1258 vcm.n39 vcm.n38 0.00321739
R1259 vcm.n18 vcm.n15 0.00321739
R1260 vcm.n28 vcm.n27 0.00321739
R1261 vcm.n32 vcm.n6 0.00321739
R1262 vcm.n75 vcm.n74 0.00321739
R1263 vcm.n79 vcm.n72 0.00321739
R1264 vcm.n62 vcm.n61 0.00321739
R1265 vcm.n66 vcm.n2 0.00321739
R1266 vcm.n106 vcm.n105 0.00321739
R1267 vcm.n110 vcm.n103 0.00321739
R1268 vcm.n121 vcm.n120 0.00321739
R1269 vcm.n99 vcm.n1 0.00239652
R1270 vcm.n87 vcm.n71 0.00239652
R1271 vcm.n53 vcm.n5 0.00239652
R1272 vcm.n41 vcm.n37 0.00239652
R1273 vcm.n30 vcm.n7 0.00239652
R1274 vcm.n77 vcm.n73 0.00239652
R1275 vcm.n64 vcm.n3 0.00239652
R1276 vcm.n108 vcm.n104 0.00239652
R1277 vcm.n258 vcm.n257 0.00239442
R1278 vcm.n323 vcm.n322 0.00239442
R1279 vcm.n460 vcm.n459 0.00239442
R1280 vcm.n391 vcm.n390 0.00239442
R1281 vcm.n797 vcm.n796 0.00239442
R1282 vcm.n863 vcm.n862 0.00239442
R1283 vcm.n931 vcm.n930 0.00239442
R1284 vcm.n985 vcm.n984 0.00239442
R1285 vcm.n377 vcm.n376 0.00225049
R1286 vcm.n484 vcm.n483 0.00225049
R1287 vcm.n182 vcm.n181 0.00225049
R1288 vcm.n236 vcm.n235 0.00225049
R1289 vcm.n225 vcm.n224 0.00225049
R1290 vcm.n164 vcm.n163 0.00225049
R1291 vcm.n173 vcm.n172 0.00225049
R1292 vcm.n247 vcm.n246 0.00225049
R1293 vcm.n191 vcm.n190 0.00225049
R1294 vcm.n312 vcm.n311 0.00225049
R1295 vcm.n334 vcm.n333 0.00225049
R1296 vcm.n419 vcm.n418 0.00225049
R1297 vcm.n405 vcm.n404 0.00225049
R1298 vcm.n476 vcm.n475 0.00225049
R1299 vcm.n468 vcm.n467 0.00225049
R1300 vcm.n531 vcm.n530 0.00225049
R1301 vcm.n520 vcm.n519 0.00225049
R1302 vcm.n301 vcm.n300 0.00225049
R1303 vcm.n542 vcm.n541 0.00225049
R1304 vcm.n553 vcm.n552 0.00225049
R1305 vcm.n710 vcm.n709 0.00225049
R1306 vcm.n648 vcm.n647 0.00225049
R1307 vcm.n634 vcm.n633 0.00225049
R1308 vcm.n702 vcm.n701 0.00225049
R1309 vcm.n693 vcm.n692 0.00225049
R1310 vcm.n626 vcm.n625 0.00225049
R1311 vcm.n612 vcm.n611 0.00225049
R1312 vcm.n685 vcm.n684 0.00225049
R1313 vcm.n939 vcm.n938 0.00225049
R1314 vcm.n947 vcm.n946 0.00225049
R1315 vcm.n849 vcm.n848 0.00225049
R1316 vcm.n877 vcm.n876 0.00225049
R1317 vcm.n1004 vcm.n1003 0.00225049
R1318 vcm.n1015 vcm.n1014 0.00225049
R1319 vcm.n1086 vcm.n1085 0.00225049
R1320 vcm.n1064 vcm.n1063 0.00225049
R1321 vcm.n1075 vcm.n1074 0.00225049
R1322 vcm.n1161 vcm.n1160 0.00225049
R1323 vcm.n1128 vcm.n1127 0.00225049
R1324 vcm.n1139 vcm.n1138 0.00225049
R1325 vcm.n1150 vcm.n1149 0.00225049
R1326 vcm.n789 vcm.n788 0.00225049
R1327 vcm.n781 vcm.n780 0.00225049
R1328 vcm.n772 vcm.n771 0.00225049
R1329 vcm.n841 vcm.n840 0.00225049
R1330 vcm.n923 vcm.n922 0.00225049
R1331 vcm.n996 vcm.n995 0.00225049
R1332 vcm.n1056 vcm.n1055 0.00225049
R1333 vcm.n262 vcm.n261 0.00149648
R1334 vcm.n338 vcm.n337 0.00149648
R1335 vcm.n355 vcm.n354 0.00149648
R1336 vcm.n412 vcm.n411 0.00149648
R1337 vcm.n409 vcm.n408 0.00149648
R1338 vcm.n513 vcm.n512 0.00149648
R1339 vcm.n398 vcm.n397 0.00149648
R1340 vcm.n395 vcm.n394 0.00149648
R1341 vcm.n557 vcm.n556 0.00149648
R1342 vcm.n584 vcm.n583 0.00149648
R1343 vcm.n641 vcm.n640 0.00149648
R1344 vcm.n638 vcm.n637 0.00149648
R1345 vcm.n592 vcm.n591 0.00149648
R1346 vcm.n619 vcm.n618 0.00149648
R1347 vcm.n616 vcm.n615 0.00149648
R1348 vcm.n602 vcm.n601 0.00149648
R1349 vcm.n1079 vcm.n1078 0.00149648
R1350 vcm.n1008 vcm.n1007 0.00149648
R1351 vcm.n867 vcm.n866 0.00149648
R1352 vcm.n834 vcm.n833 0.00149648
R1353 vcm.n831 vcm.n830 0.00149648
R1354 vcm.n853 vcm.n852 0.00149648
R1355 vcm.n968 vcm.n967 0.00149648
R1356 vcm.n989 vcm.n988 0.00149648
R1357 vcm.n1040 vcm.n1039 0.00149648
R1358 vcm.n261 vcm.n260 0.00149647
R1359 vcm.n337 vcm.n336 0.00149647
R1360 vcm.n354 vcm.n353 0.00149647
R1361 vcm.n411 vcm.n410 0.00149647
R1362 vcm.n408 vcm.n407 0.00149647
R1363 vcm.n512 vcm.n511 0.00149647
R1364 vcm.n397 vcm.n396 0.00149647
R1365 vcm.n394 vcm.n393 0.00149647
R1366 vcm.n556 vcm.n555 0.00149647
R1367 vcm.n583 vcm.n582 0.00149647
R1368 vcm.n640 vcm.n639 0.00149647
R1369 vcm.n637 vcm.n636 0.00149647
R1370 vcm.n591 vcm.n590 0.00149647
R1371 vcm.n618 vcm.n617 0.00149647
R1372 vcm.n615 vcm.n614 0.00149647
R1373 vcm.n601 vcm.n600 0.00149647
R1374 vcm.n1078 vcm.n1077 0.00149647
R1375 vcm.n1007 vcm.n1006 0.00149647
R1376 vcm.n866 vcm.n865 0.00149647
R1377 vcm.n833 vcm.n832 0.00149647
R1378 vcm.n830 vcm.n829 0.00149647
R1379 vcm.n852 vcm.n851 0.00149647
R1380 vcm.n967 vcm.n966 0.00149647
R1381 vcm.n988 vcm.n987 0.00149647
R1382 vcm.n1039 vcm.n1038 0.00149647
R1383 vcm.n240 vcm.n239 0.00145928
R1384 vcm.n294 vcm.n293 0.00145928
R1385 vcm.n384 vcm.n383 0.00145928
R1386 vcm.n881 vcm.n880 0.00145928
R1387 vcm.n1034 vcm.n1033 0.00145928
R1388 vcm.n822 vcm.n821 0.00145928
R1389 vcm.n1121 vcm.n1120 0.00145928
R1390 vcm.n25 vcm.n24 0.00145928
R1391 vcm.n46 vcm.n45 0.00145928
R1392 vcm.n59 vcm.n58 0.00145928
R1393 vcm.n92 vcm.n91 0.00145928
R1394 vcm.n117 vcm.n116 0.00145928
R1395 vcm.n239 vcm.n238 0.00139285
R1396 vcm.n293 vcm.n292 0.00139285
R1397 vcm.n383 vcm.n382 0.00139285
R1398 vcm.n880 vcm.n879 0.00139285
R1399 vcm.n1033 vcm.n1032 0.00139285
R1400 vcm.n821 vcm.n820 0.00139285
R1401 vcm.n1120 vcm.n1119 0.00139285
R1402 vcm.n24 vcm.n23 0.00139285
R1403 vcm.n45 vcm.n44 0.00139285
R1404 vcm.n58 vcm.n57 0.00139285
R1405 vcm.n91 vcm.n90 0.00139285
R1406 vcm.n116 vcm.n115 0.00139285
R1407 vcm.n145 vcm.n143 0.00114214
R1408 vcm.n897 vcm.n896 0.00104325
R1409 vcm.n436 vcm.n435 0.00104325
R1410 vcm.n570 vcm.n569 0.00104325
R1411 vcm.n727 vcm.n726 0.00104325
R1412 vcm.n660 vcm.n578 0.00103325
R1413 vcm.n496 vcm.n444 0.00103325
R1414 vcm.n347 vcm.n280 0.00103325
R1415 vcm.n1102 vcm.n1101 0.00103325
R1416 vcm.n957 vcm.n905 0.00103325
R1417 vcm.n808 vcm.n736 0.00103325
R1418 vcm.n1176 vcm.n1109 0.00103325
R1419 vcm.n808 vcm.n807 0.00103325
R1420 vcm.n957 vcm.n956 0.00103325
R1421 vcm.n1028 vcm.n1027 0.00103325
R1422 vcm.n1176 vcm.n1175 0.00103325
R1423 vcm.n1190 vcm.n1189 0.00103325
R1424 vcm.n273 vcm.n272 0.00103325
R1425 vcm.n347 vcm.n346 0.00103325
R1426 vcm.n496 vcm.n495 0.00103325
R1427 vcm.n660 vcm.n659 0.00103325
R1428 vcm.n569 vcm.n568 0.00103323
R1429 vcm.n435 vcm.n434 0.00103323
R1430 vcm.n142 vcm.n141 0.00103323
R1431 vcm.n726 vcm.n725 0.00103323
R1432 vcm.n896 vcm.n895 0.00103323
R1433 vcm.n1180 vcm.n1178 0.00103319
R1434 vcm.n1106 vcm.n1104 0.00103319
R1435 vcm.n1098 vcm.n1096 0.00103319
R1436 vcm.n961 vcm.n959 0.00103319
R1437 vcm.n902 vcm.n900 0.00103319
R1438 vcm.n733 vcm.n731 0.00103319
R1439 vcm.n575 vcm.n573 0.00103319
R1440 vcm.n441 vcm.n439 0.00103319
R1441 vcm.n277 vcm.n275 0.00103319
R1442 vcm.n206 vcm.n204 0.00103319
R1443 vcm.n1191 vcm.n1180 0.00103319
R1444 vcm.n1177 vcm.n1106 0.00103319
R1445 vcm.n1103 vcm.n1098 0.00103319
R1446 vcm.n1029 vcm.n961 0.00103319
R1447 vcm.n958 vcm.n902 0.00103319
R1448 vcm.n809 vcm.n733 0.00103319
R1449 vcm.n661 vcm.n575 0.00103319
R1450 vcm.n497 vcm.n441 0.00103319
R1451 vcm.n348 vcm.n277 0.00103319
R1452 vcm.n274 vcm.n206 0.00103319
R1453 vcm.n128 vcm.n127 0.00103293
R1454 vcm.n203 vcm.n145 0.00103293
R1455 vcm.n202 vcm.n201 0.00102352
R1456 vcm.n892 vcm.n891 0.00102352
R1457 vcm.n431 vcm.n430 0.00102352
R1458 vcm.n565 vcm.n564 0.00102352
R1459 vcm.n722 vcm.n721 0.00102352
R1460 vcm.n899 vcm.n898 0.00102346
R1461 vcm.n438 vcm.n437 0.00102346
R1462 vcm.n572 vcm.n571 0.00102346
R1463 vcm.n729 vcm.n728 0.00102346
R1464 vcm.n898 vcm.n897 0.00101835
R1465 vcm.n728 vcm.n727 0.00101835
R1466 vcm.n571 vcm.n570 0.00101835
R1467 vcm.n437 vcm.n436 0.00101835
R1468 vcm.n899 vcm.n892 0.0010183
R1469 vcm.n729 vcm.n722 0.0010183
R1470 vcm.n572 vcm.n565 0.0010183
R1471 vcm.n438 vcm.n431 0.0010183
R1472 vcm.n203 vcm.n202 0.0010183
R1473 vcm.n125 vcm.n124 0.00100588
R1474 vcm.n131 vcm.n130 0.00100116
R1475 vcm.n577 vcm.n576 0.00100116
R1476 vcm.n567 vcm.n566 0.00100116
R1477 vcm.n443 vcm.n442 0.00100116
R1478 vcm.n433 vcm.n432 0.00100116
R1479 vcm.n140 vcm.n139 0.00100116
R1480 vcm.n137 vcm.n136 0.00100116
R1481 vcm.n279 vcm.n278 0.00100116
R1482 vcm.n724 vcm.n723 0.00100116
R1483 vcm.n1100 vcm.n1099 0.00100116
R1484 vcm.n904 vcm.n903 0.00100116
R1485 vcm.n735 vcm.n734 0.00100116
R1486 vcm.n894 vcm.n893 0.00100116
R1487 vcm.n134 vcm.n133 0.00100116
R1488 vcm.n1108 vcm.n1107 0.00100116
R1489 vcm.n127 vcm.n126 0.00100034
R1490 vcm.n145 vcm.n144 0.00100034
R1491 vcm.n257 vcm.n256 0.0010003
R1492 vcm.n322 vcm.n321 0.0010003
R1493 vcm.n459 vcm.n458 0.0010003
R1494 vcm.n390 vcm.n389 0.0010003
R1495 vcm.n796 vcm.n795 0.0010003
R1496 vcm.n862 vcm.n861 0.0010003
R1497 vcm.n930 vcm.n929 0.0010003
R1498 vcm.n984 vcm.n983 0.0010003
R1499 vcm.n376 vcm.n375 0.00100024
R1500 vcm.n483 vcm.n482 0.00100024
R1501 vcm.n181 vcm.n180 0.00100024
R1502 vcm.n235 vcm.n234 0.00100024
R1503 vcm.n224 vcm.n223 0.00100024
R1504 vcm.n163 vcm.n162 0.00100024
R1505 vcm.n172 vcm.n171 0.00100024
R1506 vcm.n246 vcm.n245 0.00100024
R1507 vcm.n190 vcm.n189 0.00100024
R1508 vcm.n311 vcm.n310 0.00100024
R1509 vcm.n333 vcm.n332 0.00100024
R1510 vcm.n418 vcm.n417 0.00100024
R1511 vcm.n404 vcm.n403 0.00100024
R1512 vcm.n475 vcm.n474 0.00100024
R1513 vcm.n467 vcm.n466 0.00100024
R1514 vcm.n530 vcm.n529 0.00100024
R1515 vcm.n519 vcm.n518 0.00100024
R1516 vcm.n300 vcm.n299 0.00100024
R1517 vcm.n541 vcm.n540 0.00100024
R1518 vcm.n552 vcm.n551 0.00100024
R1519 vcm.n709 vcm.n708 0.00100024
R1520 vcm.n647 vcm.n646 0.00100024
R1521 vcm.n633 vcm.n632 0.00100024
R1522 vcm.n701 vcm.n700 0.00100024
R1523 vcm.n692 vcm.n691 0.00100024
R1524 vcm.n625 vcm.n624 0.00100024
R1525 vcm.n611 vcm.n610 0.00100024
R1526 vcm.n684 vcm.n683 0.00100024
R1527 vcm.n938 vcm.n937 0.00100024
R1528 vcm.n946 vcm.n945 0.00100024
R1529 vcm.n848 vcm.n847 0.00100024
R1530 vcm.n876 vcm.n875 0.00100024
R1531 vcm.n1003 vcm.n1002 0.00100024
R1532 vcm.n1014 vcm.n1013 0.00100024
R1533 vcm.n1085 vcm.n1084 0.00100024
R1534 vcm.n1063 vcm.n1062 0.00100024
R1535 vcm.n1074 vcm.n1073 0.00100024
R1536 vcm.n1160 vcm.n1159 0.00100024
R1537 vcm.n1127 vcm.n1126 0.00100024
R1538 vcm.n1138 vcm.n1137 0.00100024
R1539 vcm.n1149 vcm.n1148 0.00100024
R1540 vcm.n788 vcm.n787 0.00100024
R1541 vcm.n780 vcm.n779 0.00100024
R1542 vcm.n771 vcm.n770 0.00100024
R1543 vcm.n840 vcm.n839 0.00100024
R1544 vcm.n922 vcm.n921 0.00100024
R1545 vcm.n995 vcm.n994 0.00100024
R1546 vcm.n1055 vcm.n1054 0.00100024
R1547 vcm.n100 vcm.n1 0.00100019
R1548 vcm.n88 vcm.n71 0.00100019
R1549 vcm.n54 vcm.n5 0.00100019
R1550 vcm.n42 vcm.n37 0.00100019
R1551 vcm.n31 vcm.n7 0.00100019
R1552 vcm.n78 vcm.n73 0.00100019
R1553 vcm.n65 vcm.n3 0.00100019
R1554 vcm.n109 vcm.n104 0.00100019
R1555 vcm.n676 vcm.n675 0.00100017
R1556 vcm.n1180 vcm.n1179 0.00100008
R1557 vcm.n1106 vcm.n1105 0.00100008
R1558 vcm.n1098 vcm.n1097 0.00100008
R1559 vcm.n961 vcm.n960 0.00100008
R1560 vcm.n902 vcm.n901 0.00100008
R1561 vcm.n733 vcm.n732 0.00100008
R1562 vcm.n575 vcm.n574 0.00100008
R1563 vcm.n441 vcm.n440 0.00100008
R1564 vcm.n277 vcm.n276 0.00100008
R1565 vcm.n206 vcm.n205 0.00100008
R1566 vcm.n143 vcm.n142 0.00100006
R1567 vcm.n1192 vcm.n129 0.00100006
R1568 vcm.n218 vcm.n217 0.00100005
R1569 vcm.n229 vcm.n228 0.00100005
R1570 vcm.n316 vcm.n315 0.00100005
R1571 vcm.n327 vcm.n326 0.00100005
R1572 vcm.n251 vcm.n250 0.00100005
R1573 vcm.n352 vcm.n351 0.00100005
R1574 vcm.n546 vcm.n545 0.00100005
R1575 vcm.n605 vcm.n604 0.00100005
R1576 vcm.n367 vcm.n366 0.00100005
R1577 vcm.n370 vcm.n369 0.00100005
R1578 vcm.n305 vcm.n304 0.00100005
R1579 vcm.n524 vcm.n523 0.00100005
R1580 vcm.n381 vcm.n380 0.00100005
R1581 vcm.n535 vcm.n534 0.00100005
R1582 vcm.n581 vcm.n580 0.00100005
R1583 vcm.n589 vcm.n588 0.00100005
R1584 vcm.n884 vcm.n883 0.00100005
R1585 vcm.n1019 vcm.n1018 0.00100005
R1586 vcm.n1165 vcm.n1164 0.00100005
R1587 vcm.n1154 vcm.n1153 0.00100005
R1588 vcm.n870 vcm.n869 0.00100005
R1589 vcm.n856 vcm.n855 0.00100005
R1590 vcm.n819 vcm.n818 0.00100005
R1591 vcm.n978 vcm.n977 0.00100005
R1592 vcm.n1143 vcm.n1142 0.00100005
R1593 vcm.n1068 vcm.n1067 0.00100005
R1594 vcm.n1132 vcm.n1131 0.00100005
R1595 vcm.n1049 vcm.n1048 0.00100005
R1596 vcm.n21 vcm.n20 0.00100005
R1597 vcm.n82 vcm.n81 0.00100005
R1598 vcm.n113 vcm.n112 0.00100005
R1599 vcm.n48 vcm.n35 0.00100005
R1600 vcm.n94 vcm.n69 0.00100005
R1601 vcm.n1191 vcm.n1190 0.00100005
R1602 vcm.n1177 vcm.n1176 0.00100005
R1603 vcm.n1103 vcm.n1102 0.00100005
R1604 vcm.n1029 vcm.n1028 0.00100005
R1605 vcm.n958 vcm.n957 0.00100005
R1606 vcm.n809 vcm.n808 0.00100005
R1607 vcm.n661 vcm.n660 0.00100005
R1608 vcm.n497 vcm.n496 0.00100005
R1609 vcm.n348 vcm.n347 0.00100005
R1610 vcm.n274 vcm.n273 0.00100005
R1611 vcm.n35 vcm.n34 0.00100004
R1612 vcm.n69 vcm.n68 0.00100004
R1613 vcm.n217 vcm.n216 0.00100004
R1614 vcm.n228 vcm.n227 0.00100004
R1615 vcm.n315 vcm.n314 0.00100004
R1616 vcm.n326 vcm.n325 0.00100004
R1617 vcm.n250 vcm.n249 0.00100004
R1618 vcm.n351 vcm.n350 0.00100004
R1619 vcm.n545 vcm.n544 0.00100004
R1620 vcm.n604 vcm.n603 0.00100004
R1621 vcm.n366 vcm.n365 0.00100004
R1622 vcm.n369 vcm.n368 0.00100004
R1623 vcm.n304 vcm.n303 0.00100004
R1624 vcm.n523 vcm.n522 0.00100004
R1625 vcm.n380 vcm.n379 0.00100004
R1626 vcm.n534 vcm.n533 0.00100004
R1627 vcm.n580 vcm.n579 0.00100004
R1628 vcm.n588 vcm.n587 0.00100004
R1629 vcm.n883 vcm.n882 0.00100004
R1630 vcm.n1018 vcm.n1017 0.00100004
R1631 vcm.n1164 vcm.n1163 0.00100004
R1632 vcm.n1153 vcm.n1152 0.00100004
R1633 vcm.n869 vcm.n868 0.00100004
R1634 vcm.n855 vcm.n854 0.00100004
R1635 vcm.n818 vcm.n817 0.00100004
R1636 vcm.n977 vcm.n976 0.00100004
R1637 vcm.n1142 vcm.n1141 0.00100004
R1638 vcm.n1067 vcm.n1066 0.00100004
R1639 vcm.n1131 vcm.n1130 0.00100004
R1640 vcm.n1048 vcm.n1047 0.00100004
R1641 vcm.n20 vcm.n19 0.00100004
R1642 vcm.n81 vcm.n80 0.00100004
R1643 vcm.n112 vcm.n111 0.00100004
R1644 vcm.n128 vcm.n123 0.000533349
R1645 vcm.n1193 vcm.n128 0.000533349
R1646 vcm.n891 vcm.n810 0.000533349
R1647 vcm.n959 vcm.n135 0.000533349
R1648 vcm.n1096 vcm.n1095 0.000533349
R1649 vcm.n1178 vcm.n132 0.000533349
R1650 vcm.n204 vcm.n138 0.000533349
R1651 vcm.n430 vcm.n349 0.000533349
R1652 vcm.n564 vcm.n498 0.000533349
R1653 vcm.n721 vcm.n662 0.000533349
R1654 vcm.n1193 vcm.n1192 0.000533349
R1655 vcm.n568 vcm.n567 0.00050467
R1656 vcm.n434 vcm.n433 0.00050467
R1657 vcm.n141 vcm.n140 0.00050467
R1658 vcm.n725 vcm.n724 0.00050467
R1659 vcm.n895 vcm.n894 0.00050467
R1660 vcm.n201 vcm.n200 0.00050467
R1661 vcm.n736 vcm.n735 0.00050467
R1662 vcm.n807 vcm.n806 0.00050467
R1663 vcm.n891 vcm.n890 0.00050467
R1664 vcm.n905 vcm.n904 0.00050467
R1665 vcm.n956 vcm.n955 0.00050467
R1666 vcm.n135 vcm.n134 0.00050467
R1667 vcm.n1027 vcm.n1026 0.00050467
R1668 vcm.n1101 vcm.n1100 0.00050467
R1669 vcm.n1095 vcm.n1094 0.00050467
R1670 vcm.n1109 vcm.n1108 0.00050467
R1671 vcm.n1175 vcm.n1174 0.00050467
R1672 vcm.n132 vcm.n131 0.00050467
R1673 vcm.n1189 vcm.n1188 0.00050467
R1674 vcm.n138 vcm.n137 0.00050467
R1675 vcm.n272 vcm.n271 0.00050467
R1676 vcm.n280 vcm.n279 0.00050467
R1677 vcm.n346 vcm.n345 0.00050467
R1678 vcm.n430 vcm.n429 0.00050467
R1679 vcm.n444 vcm.n443 0.00050467
R1680 vcm.n495 vcm.n494 0.00050467
R1681 vcm.n564 vcm.n563 0.00050467
R1682 vcm.n578 vcm.n577 0.00050467
R1683 vcm.n659 vcm.n658 0.00050467
R1684 vcm.n721 vcm.n720 0.00050467
R1685 vcm.n126 vcm.n125 0.00050467
R1686 vcm.n1194 vcm.n1193 0.00050467
R1687 vcm.n200 vcm.n199 0.000502311
R1688 vcm.n1195 vcm.n1194 0.000502311
R1689 vcm.n1188 vcm.n1187 0.000502311
R1690 vcm.n658 vcm.n657 0.000502311
R1691 vcm.n563 vcm.n562 0.000502311
R1692 vcm.n494 vcm.n493 0.000502311
R1693 vcm.n429 vcm.n428 0.000502311
R1694 vcm.n271 vcm.n270 0.000502311
R1695 vcm.n345 vcm.n344 0.000502311
R1696 vcm.n720 vcm.n719 0.000502311
R1697 vcm.n1094 vcm.n1093 0.000502311
R1698 vcm.n955 vcm.n954 0.000502311
R1699 vcm.n806 vcm.n805 0.000502311
R1700 vcm.n890 vcm.n889 0.000502311
R1701 vcm.n1026 vcm.n1025 0.000502311
R1702 vcm.n1174 vcm.n1173 0.000502311
R1703 vcm.n761 vcm.n760 0.000500172
R1704 vcm.n764 vcm.n763 0.000500095
R1705 vcm.n678 vcm.n677 0.000500095
R1706 VSS.n5935 VSS.n5934 34571.4
R1707 VSS.n2946 VSS.n2945 34571.4
R1708 VSS.n3070 VSS.n3069 34571.4
R1709 VSS.n3067 VSS.n3065 34571.4
R1710 VSS.n6054 VSS.n1943 34571.4
R1711 VSS.n6048 VSS.n1945 34571.4
R1712 VSS.n6042 VSS.n1948 34571.4
R1713 VSS.n2352 VSS.n2351 23783
R1714 VSS.n2947 VSS.n2946 22403.2
R1715 VSS.n6055 VSS.n6054 22403.2
R1716 VSS.n5882 VSS.n5881 21511.1
R1717 VSS.n6011 VSS.n6010 21511.1
R1718 VSS.n1900 VSS.n1899 21511.1
R1719 VSS.n6745 VSS.n1020 21511.1
R1720 VSS.n3256 VSS.n2961 21511.1
R1721 VSS.n3078 VSS.n2989 21511.1
R1722 VSS.n5504 VSS.n5501 21511.1
R1723 VSS.n5506 VSS.n2080 21511.1
R1724 VSS.n5555 VSS.n2076 21511.1
R1725 VSS.n3270 VSS.n3269 21511.1
R1726 VSS.n3126 VSS.n3125 21511.1
R1727 VSS.n3220 VSS.n3219 21511.1
R1728 VSS.n5520 VSS.n5493 21511.1
R1729 VSS.n5522 VSS.n2091 21511.1
R1730 VSS.n5490 VSS.n5489 21511.1
R1731 VSS.n6235 VSS.n1903 21511.1
R1732 VSS.n6038 VSS.n1949 21511.1
R1733 VSS.n6044 VSS.n1947 21511.1
R1734 VSS.n1931 VSS.n1930 21511.1
R1735 VSS.n1937 VSS.n1936 21511.1
R1736 VSS.n6050 VSS.n1944 21511.1
R1737 VSS.n6031 VSS.n1950 21511.1
R1738 VSS.n1908 VSS.n1021 21511.1
R1739 VSS.n6737 VSS.n6736 21511.1
R1740 VSS.n6758 VSS.n6757 21511.1
R1741 VSS.n2017 VSS.n2016 21511.1
R1742 VSS.n2083 VSS.n2082 21511.1
R1743 VSS.n5934 VSS.n5933 21229.4
R1744 VSS.n6033 VSS.n6032 18464.3
R1745 VSS.n6037 VSS.n6036 18464.3
R1746 VSS.n3067 VSS.n3066 18464.3
R1747 VSS.n3279 VSS.n3278 18464.3
R1748 VSS.n3272 VSS.n3271 18464.3
R1749 VSS.n6049 VSS.n6048 18464.3
R1750 VSS.n6043 VSS.n6042 18464.3
R1751 VSS.n2993 VSS.n2990 17285.7
R1752 VSS.n3084 VSS.n3083 17285.7
R1753 VSS.n3258 VSS.n2956 17285.7
R1754 VSS.n3267 VSS.n3266 17285.7
R1755 VSS.n3289 VSS.n3286 17285.7
R1756 VSS.n2999 VSS.n2987 17285.7
R1757 VSS.n3093 VSS.n3092 17285.7
R1758 VSS.n3160 VSS.n3157 17285.7
R1759 VSS.n3167 VSS.n3153 17285.7
R1760 VSS.n3170 VSS.n3169 17285.7
R1761 VSS.n3005 VSS.n2984 17285.7
R1762 VSS.n3102 VSS.n3101 17285.7
R1763 VSS.n3143 VSS.n3140 17285.7
R1764 VSS.n3187 VSS.n3186 17285.7
R1765 VSS.n3184 VSS.n3183 17285.7
R1766 VSS.n3048 VSS.n2981 17285.7
R1767 VSS.n3111 VSS.n3110 17285.7
R1768 VSS.n3198 VSS.n3195 17285.7
R1769 VSS.n3205 VSS.n3135 17285.7
R1770 VSS.n3208 VSS.n3207 17285.7
R1771 VSS.n3014 VSS.n3013 17285.7
R1772 VSS.n3121 VSS.n3119 17285.7
R1773 VSS.n3124 VSS.n3123 17285.7
R1774 VSS.n3229 VSS.n3228 17285.7
R1775 VSS.n3308 VSS.n2931 17285.7
R1776 VSS.n3020 VSS.n2786 17285.7
R1777 VSS.n5545 VSS.n5544 17285.7
R1778 VSS.n2792 VSS.n2791 17285.7
R1779 VSS.n2924 VSS.n2921 17285.7
R1780 VSS.n5552 VSS.n2783 17285.7
R1781 VSS.n5511 VSS.n5510 17285.7
R1782 VSS.n5517 VSS.n5516 17285.7
R1783 VSS.n5495 VSS.n5494 17285.7
R1784 VSS.n2041 VSS.n2040 17285.7
R1785 VSS.n2058 VSS.n2057 17285.7
R1786 VSS.n1986 VSS.n1980 17285.7
R1787 VSS.n6771 VSS.n1012 17285.7
R1788 VSS.n5953 VSS.n2007 17285.7
R1789 VSS.n5960 VSS.n2004 17285.7
R1790 VSS.n2002 VSS.n2001 17285.7
R1791 VSS.n1999 VSS.n1998 17285.7
R1792 VSS.n1996 VSS.n1995 17285.7
R1793 VSS.n5917 VSS.n1964 17285.7
R1794 VSS.n5982 VSS.n5981 17285.7
R1795 VSS.n5976 VSS.n5975 17285.7
R1796 VSS.n5973 VSS.n1004 17285.7
R1797 VSS.n6785 VSS.n6784 17285.7
R1798 VSS.n5991 VSS.n1960 17285.7
R1799 VSS.n6003 VSS.n6002 17285.7
R1800 VSS.n6000 VSS.n5999 17285.7
R1801 VSS.n6798 VSS.n6797 17285.7
R1802 VSS.n6026 VSS.n1951 17285.7
R1803 VSS.n6016 VSS.n6014 17285.7
R1804 VSS.n1934 VSS.n1933 17285.7
R1805 VSS.n1942 VSS.n1941 17285.7
R1806 VSS.n2030 VSS.n2029 17285.7
R1807 VSS.n2034 VSS.n2033 17285.7
R1808 VSS.n6764 VSS.n6762 17285.7
R1809 VSS.n2021 VSS.n2020 17285.7
R1810 VSS.n1866 VSS.n1028 17283.5
R1811 VSS.n2176 VSS.n2175 14040.1
R1812 VSS.n2961 VSS.n2960 12320
R1813 VSS.n3280 VSS.n3279 12320
R1814 VSS.n3271 VSS.n3270 12320
R1815 VSS.n6038 VSS.n6037 12320
R1816 VSS.n6044 VSS.n6043 12320
R1817 VSS.n6050 VSS.n6049 12320
R1818 VSS.n6032 VSS.n6031 12320
R1819 VSS.n5490 VSS.n2092 11061.4
R1820 VSS.n3085 VSS.n2990 11000
R1821 VSS.n3085 VSS.n3084 11000
R1822 VSS.n3258 VSS.n3257 11000
R1823 VSS.n3268 VSS.n2956 11000
R1824 VSS.n3268 VSS.n3267 11000
R1825 VSS.n3266 VSS.n2943 11000
R1826 VSS.n3286 VSS.n2943 11000
R1827 VSS.n3094 VSS.n2987 11000
R1828 VSS.n3094 VSS.n3093 11000
R1829 VSS.n3092 VSS.n3091 11000
R1830 VSS.n3161 VSS.n3160 11000
R1831 VSS.n3161 VSS.n3153 11000
R1832 VSS.n3171 VSS.n3167 11000
R1833 VSS.n3171 VSS.n3170 11000
R1834 VSS.n3103 VSS.n2984 11000
R1835 VSS.n3103 VSS.n3102 11000
R1836 VSS.n3101 VSS.n3100 11000
R1837 VSS.n3188 VSS.n3143 11000
R1838 VSS.n3188 VSS.n3187 11000
R1839 VSS.n3186 VSS.n3185 11000
R1840 VSS.n3185 VSS.n3184 11000
R1841 VSS.n3112 VSS.n2981 11000
R1842 VSS.n3112 VSS.n3111 11000
R1843 VSS.n3110 VSS.n3109 11000
R1844 VSS.n3199 VSS.n3198 11000
R1845 VSS.n3199 VSS.n3135 11000
R1846 VSS.n3209 VSS.n3205 11000
R1847 VSS.n3209 VSS.n3208 11000
R1848 VSS.n3014 VSS.n2978 11000
R1849 VSS.n3119 VSS.n2978 11000
R1850 VSS.n3121 VSS.n3120 11000
R1851 VSS.n3230 VSS.n3124 11000
R1852 VSS.n3230 VSS.n3229 11000
R1853 VSS.n3228 VSS.n3227 11000
R1854 VSS.n3227 VSS.n2931 11000
R1855 VSS.n5546 VSS.n2786 11000
R1856 VSS.n5546 VSS.n5545 11000
R1857 VSS.n2920 VSS.n2795 11000
R1858 VSS.n2921 VSS.n2920 11000
R1859 VSS.n5552 VSS.n5551 11000
R1860 VSS.n2059 VSS.n2041 11000
R1861 VSS.n2059 VSS.n2058 11000
R1862 VSS.n2057 VSS.n2056 11000
R1863 VSS.n2056 VSS.n2055 11000
R1864 VSS.n1978 VSS.n1977 11000
R1865 VSS.n1980 VSS.n1978 11000
R1866 VSS.n1986 VSS.n1985 11000
R1867 VSS.n1985 VSS.n1012 11000
R1868 VSS.n5954 VSS.n5953 11000
R1869 VSS.n5954 VSS.n2004 11000
R1870 VSS.n5961 VSS.n5960 11000
R1871 VSS.n2001 VSS.n2000 11000
R1872 VSS.n2000 VSS.n1999 11000
R1873 VSS.n1998 VSS.n1997 11000
R1874 VSS.n1997 VSS.n1996 11000
R1875 VSS.n5983 VSS.n1964 11000
R1876 VSS.n5983 VSS.n5982 11000
R1877 VSS.n5976 VSS.n5970 11000
R1878 VSS.n5975 VSS.n5974 11000
R1879 VSS.n5974 VSS.n5973 11000
R1880 VSS.n6786 VSS.n1004 11000
R1881 VSS.n6786 VSS.n6785 11000
R1882 VSS.n5992 VSS.n5991 11000
R1883 VSS.n5993 VSS.n5992 11000
R1884 VSS.n6004 VSS.n5996 11000
R1885 VSS.n6004 VSS.n6003 11000
R1886 VSS.n6002 VSS.n6001 11000
R1887 VSS.n6001 VSS.n6000 11000
R1888 VSS.n5999 VSS.n1001 11000
R1889 VSS.n6797 VSS.n1001 11000
R1890 VSS.n6026 VSS.n6025 11000
R1891 VSS.n6025 VSS.n6024 11000
R1892 VSS.n6013 VSS.n1954 11000
R1893 VSS.n6014 VSS.n6013 11000
R1894 VSS.n6016 VSS.n6015 11000
R1895 VSS.n6015 VSS.n1933 11000
R1896 VSS.n1940 VSS.n1934 11000
R1897 VSS.n1941 VSS.n1940 11000
R1898 VSS.n2035 VSS.n2030 11000
R1899 VSS.n2035 VSS.n2034 11000
R1900 VSS.n2049 VSS.n1904 11000
R1901 VSS.n1914 VSS.n1905 11000
R1902 VSS.n1914 VSS.n1913 11000
R1903 VSS.n1910 VSS.n1016 11000
R1904 VSS.n6762 VSS.n1016 11000
R1905 VSS.n2024 VSS.n2021 11000
R1906 VSS.n2024 VSS.n2023 11000
R1907 VSS.n6239 VSS.n6238 11000
R1908 VSS.n6238 VSS.n6237 11000
R1909 VSS.n6750 VSS.n6749 11000
R1910 VSS.n6751 VSS.n6750 11000
R1911 VSS.n6753 VSS.n1018 11000
R1912 VSS.n6597 VSS.n1018 11000
R1913 VSS.n2050 VSS.n2049 10951.1
R1914 VSS.n2056 VSS.n2044 10951.1
R1915 VSS.n2056 VSS.n2045 10951.1
R1916 VSS.n5962 VSS.n5961 10951.1
R1917 VSS.n5970 VSS.n5969 10951.1
R1918 VSS.n5984 VSS.n5983 10951.1
R1919 VSS.n5992 VSS.n1958 10951.1
R1920 VSS.n2060 VSS.n2059 10951.1
R1921 VSS.n5955 VSS.n5954 10951.1
R1922 VSS.n2036 VSS.n2035 10951.1
R1923 VSS.n2059 VSS.n2037 10951.1
R1924 VSS.n2025 VSS.n2024 10951.1
R1925 VSS.n2035 VSS.n2026 10951.1
R1926 VSS.n6238 VSS.n1900 10951.1
R1927 VSS.n6750 VSS.n1020 10951.1
R1928 VSS.n3120 VSS.n2977 10951.1
R1929 VSS.n3109 VSS.n2973 10951.1
R1930 VSS.n3100 VSS.n2969 10951.1
R1931 VSS.n3091 VSS.n2965 10951.1
R1932 VSS.n3086 VSS.n3085 10951.1
R1933 VSS.n3094 VSS.n2986 10951.1
R1934 VSS.n3095 VSS.n3094 10951.1
R1935 VSS.n3103 VSS.n2983 10951.1
R1936 VSS.n3104 VSS.n3103 10951.1
R1937 VSS.n3112 VSS.n2980 10951.1
R1938 VSS.n3257 VSS.n3256 10951.1
R1939 VSS.n3085 VSS.n2989 10951.1
R1940 VSS.n3113 VSS.n3112 10951.1
R1941 VSS.n3115 VSS.n2978 10951.1
R1942 VSS.n5500 VSS.n5499 10951.1
R1943 VSS.n3022 VSS.n2978 10951.1
R1944 VSS.n5546 VSS.n2785 10951.1
R1945 VSS.n5547 VSS.n5546 10951.1
R1946 VSS.n5551 VSS.n5550 10951.1
R1947 VSS.n5501 VSS.n5500 10951.1
R1948 VSS.n5505 VSS.n5504 10951.1
R1949 VSS.n5506 VSS.n5505 10951.1
R1950 VSS.n5870 VSS.n2080 10951.1
R1951 VSS.n5876 VSS.n2076 10951.1
R1952 VSS.n3282 VSS.n2943 10951.1
R1953 VSS.n3269 VSS.n3268 10951.1
R1954 VSS.n3162 VSS.n3161 10951.1
R1955 VSS.n3172 VSS.n3171 10951.1
R1956 VSS.n3185 VSS.n3145 10951.1
R1957 VSS.n3189 VSS.n3188 10951.1
R1958 VSS.n3200 VSS.n3199 10951.1
R1959 VSS.n3210 VSS.n3209 10951.1
R1960 VSS.n3227 VSS.n3226 10951.1
R1961 VSS.n3231 VSS.n3230 10951.1
R1962 VSS.n5488 VSS.n2798 10951.1
R1963 VSS.n5493 VSS.n5492 10951.1
R1964 VSS.n5521 VSS.n5520 10951.1
R1965 VSS.n5522 VSS.n5521 10951.1
R1966 VSS.n5864 VSS.n2091 10951.1
R1967 VSS.n5489 VSS.n5488 10951.1
R1968 VSS.n6238 VSS.n6235 10951.1
R1969 VSS.n2049 VSS.n1903 10951.1
R1970 VSS.n5954 VSS.n2006 10951.1
R1971 VSS.n5983 VSS.n1963 10951.1
R1972 VSS.n5992 VSS.n1959 10951.1
R1973 VSS.n6025 VSS.n1952 10951.1
R1974 VSS.n6005 VSS.n6004 10951.1
R1975 VSS.n1985 VSS.n1984 10951.1
R1976 VSS.n1997 VSS.n1971 10951.1
R1977 VSS.n2000 VSS.n1920 10951.1
R1978 VSS.n5974 VSS.n1924 10951.1
R1979 VSS.n6787 VSS.n6786 10951.1
R1980 VSS.n6793 VSS.n1001 10951.1
R1981 VSS.n6001 VSS.n1928 10951.1
R1982 VSS.n6025 VSS.n1950 10951.1
R1983 VSS.n6750 VSS.n1021 10951.1
R1984 VSS.n1914 VSS.n1908 10951.1
R1985 VSS.n1915 VSS.n1914 10951.1
R1986 VSS.n1978 VSS.n1916 10951.1
R1987 VSS.n6737 VSS.n1018 10951.1
R1988 VSS.n6757 VSS.n1018 10951.1
R1989 VSS.n3289 VSS.n3288 9232.14
R1990 VSS.n3169 VSS.n3168 9232.14
R1991 VSS.n3183 VSS.n3182 9232.14
R1992 VSS.n3207 VSS.n3206 9232.14
R1993 VSS.n3308 VSS.n3307 9232.14
R1994 VSS.n2928 VSS.n2924 9232.14
R1995 VSS.n2801 VSS.n2800 9232.14
R1996 VSS.n6771 VSS.n6770 9232.14
R1997 VSS.n1995 VSS.n1994 9232.14
R1998 VSS.n6784 VSS.n6783 9232.14
R1999 VSS.n6799 VSS.n6798 9232.14
R2000 VSS.n6198 VSS.n1942 9232.14
R2001 VSS.n6764 VSS.n6763 9232.14
R2002 VSS.n6603 VSS.n6602 9232.14
R2003 VSS.n2773 VSS.n2015 6020.82
R2004 VSS.n6247 VSS.n1897 6020.82
R2005 VSS.n2992 VSS.n2991 4827.93
R2006 VSS.n2998 VSS.n2997 4827.93
R2007 VSS.n3004 VSS.n3003 4827.93
R2008 VSS.n3010 VSS.n3009 4827.93
R2009 VSS.n3046 VSS.n3045 4827.93
R2010 VSS.n3043 VSS.n3042 4827.93
R2011 VSS.n3040 VSS.n3039 4827.93
R2012 VSS.n3037 VSS.n3036 4827.93
R2013 VSS.n5897 VSS.n5896 4827.93
R2014 VSS.n5902 VSS.n5901 4827.93
R2015 VSS.n5908 VSS.n5906 4827.93
R2016 VSS.n5913 VSS.n2008 4827.93
R2017 VSS.n5916 VSS.n5915 4827.93
R2018 VSS.n5926 VSS.n5925 4827.93
R2019 VSS.n5929 VSS.n5928 4827.93
R2020 VSS.n5933 VSS.n5932 4827.93
R2021 VSS.n1867 VSS.n1866 4810.3
R2022 VSS.n3288 VSS.n3287 4376.55
R2023 VSS.n3288 VSS.n2941 4376.55
R2024 VSS.n3168 VSS.n2940 4376.55
R2025 VSS.n3168 VSS.n2938 4376.55
R2026 VSS.n3182 VSS.n2937 4376.55
R2027 VSS.n3182 VSS.n2935 4376.55
R2028 VSS.n3206 VSS.n2934 4376.55
R2029 VSS.n3206 VSS.n2932 4376.55
R2030 VSS.n3307 VSS.n3306 4376.55
R2031 VSS.n3307 VSS.n2930 4376.55
R2032 VSS.n2929 VSS.n2928 4376.55
R2033 VSS.n2928 VSS.n2927 4376.55
R2034 VSS.n2802 VSS.n2801 4376.55
R2035 VSS.n6602 VSS.n6600 4376.55
R2036 VSS.n6602 VSS.n6601 4376.55
R2037 VSS.n6763 VSS.n1013 4376.55
R2038 VSS.n6770 VSS.n6769 4376.55
R2039 VSS.n6770 VSS.n1010 4376.55
R2040 VSS.n1994 VSS.n1009 4376.55
R2041 VSS.n1994 VSS.n1007 4376.55
R2042 VSS.n6783 VSS.n1006 4376.55
R2043 VSS.n6783 VSS.n6782 4376.55
R2044 VSS.n6800 VSS.n6799 4376.55
R2045 VSS.n6799 VSS.n960 4376.55
R2046 VSS.n6199 VSS.n6198 4376.55
R2047 VSS.n6198 VSS.n6197 4376.55
R2048 VSS.n2776 VSS.n2775 3147.35
R2049 VSS.n2774 VSS.n2073 3147.35
R2050 VSS.n5888 VSS.n5887 3147.35
R2051 VSS.n6246 VSS.n1898 3147.35
R2052 VSS.n6251 VSS.n6250 3147.35
R2053 VSS.n2996 VSS.n2992 3072.32
R2054 VSS.n2997 VSS.n2996 3072.32
R2055 VSS.n3002 VSS.n2998 3072.32
R2056 VSS.n3003 VSS.n3002 3072.32
R2057 VSS.n3008 VSS.n3004 3072.32
R2058 VSS.n3009 VSS.n3008 3072.32
R2059 VSS.n3011 VSS.n3010 3072.32
R2060 VSS.n3046 VSS.n3011 3072.32
R2061 VSS.n3045 VSS.n3044 3072.32
R2062 VSS.n3044 VSS.n3043 3072.32
R2063 VSS.n3042 VSS.n3041 3072.32
R2064 VSS.n3041 VSS.n3040 3072.32
R2065 VSS.n3039 VSS.n3038 3072.32
R2066 VSS.n3038 VSS.n3037 3072.32
R2067 VSS.n5897 VSS.n2012 3072.32
R2068 VSS.n5901 VSS.n2012 3072.32
R2069 VSS.n5902 VSS.n2010 3072.32
R2070 VSS.n5906 VSS.n2010 3072.32
R2071 VSS.n5908 VSS.n5907 3072.32
R2072 VSS.n5907 VSS.n2008 3072.32
R2073 VSS.n5914 VSS.n5913 3072.32
R2074 VSS.n5915 VSS.n5914 3072.32
R2075 VSS.n5924 VSS.n5916 3072.32
R2076 VSS.n5925 VSS.n5924 3072.32
R2077 VSS.n5927 VSS.n5926 3072.32
R2078 VSS.n5928 VSS.n5927 3072.32
R2079 VSS.n5931 VSS.n5929 3072.32
R2080 VSS.n5932 VSS.n5931 3072.32
R2081 VSS.n2780 VSS.n2779 3014.53
R2082 VSS.n5860 VSS.n2092 2895.44
R2083 VSS.n3036 VSS.n2781 2574.58
R2084 VSS.n2773 VSS.n2014 1881.22
R2085 VSS.n2776 VSS.n2015 1881.22
R2086 VSS.n2775 VSS.n2774 1881.22
R2087 VSS.n5884 VSS.n2073 1881.22
R2088 VSS.n5889 VSS.n5888 1881.22
R2089 VSS.n5887 VSS.n1898 1881.22
R2090 VSS.n6247 VSS.n6246 1881.22
R2091 VSS.n6250 VSS.n1897 1881.22
R2092 VSS.t83 VSS.t76 1584.67
R2093 VSS.t85 VSS.t90 1584.67
R2094 VSS.t96 VSS.t47 1584.67
R2095 VSS.t45 VSS.t49 1584.67
R2096 VSS.t288 VSS.t40 1584.67
R2097 VSS.t74 VSS.t51 1584.67
R2098 VSS.n6253 VSS.n6252 1544.68
R2099 VSS.n2247 VSS.t103 1475.1
R2100 VSS VSS.t98 1298.08
R2101 VSS VSS.t72 1298.08
R2102 VSS.n6714 VSS 1088
R2103 VSS.n5836 VSS 1088
R2104 VSS.n5485 VSS 1088
R2105 VSS.n3313 VSS 1088
R2106 VSS.n3302 VSS 1088
R2107 VSS.n3298 VSS 1088
R2108 VSS.n1011 VSS 1088
R2109 VSS.n6195 VSS 1088
R2110 VSS.n6804 VSS 1088
R2111 VSS.n1000 VSS 1088
R2112 VSS.n6252 VSS.n6251 1073.06
R2113 VSS.n6254 VSS.n1895 1043.16
R2114 VSS.n6304 VSS.n6302 922.486
R2115 VSS.n6254 VSS.n6253 918.338
R2116 VSS VSS.t120 893.487
R2117 VSS.t122 VSS 885.058
R2118 VSS.t101 VSS 885.058
R2119 VSS.t293 VSS 885.058
R2120 VSS.n4962 VSS.n4961 880.317
R2121 VSS.n4626 VSS.n4625 880.317
R2122 VSS.n4615 VSS.n4614 880.317
R2123 VSS.n5272 VSS.n5271 880.317
R2124 VSS.n4347 VSS.n4346 880.317
R2125 VSS.n4655 VSS.n4261 880.317
R2126 VSS.n4926 VSS.n4925 880.317
R2127 VSS.n5158 VSS.n5157 880.317
R2128 VSS.n5145 VSS.n5144 880.317
R2129 VSS.n4833 VSS.n4832 880.317
R2130 VSS.n4677 VSS.n4233 880.317
R2131 VSS.n4742 VSS.n4741 880.317
R2132 VSS.n4728 VSS.n4727 880.317
R2133 VSS.n5207 VSS.n5206 880.317
R2134 VSS.n4666 VSS.n4665 880.317
R2135 VSS.n4042 VSS.n4041 880.317
R2136 VSS.n4055 VSS.n4054 880.317
R2137 VSS.n4066 VSS.n3985 880.317
R2138 VSS.n4094 VSS.n4093 880.317
R2139 VSS.n3971 VSS.n3970 880.317
R2140 VSS.n5262 VSS.n5261 880.317
R2141 VSS.n5771 VSS.n5770 880.317
R2142 VSS.n5739 VSS.n5738 880.317
R2143 VSS.n5707 VSS.n5706 880.317
R2144 VSS.n2604 VSS.n2603 880.317
R2145 VSS.n2583 VSS.n2582 880.317
R2146 VSS.n2629 VSS.n2510 880.317
R2147 VSS.n7458 VSS.n7457 880.317
R2148 VSS.n533 VSS.n431 880.317
R2149 VSS.n661 VSS.n660 880.317
R2150 VSS.n7047 VSS.n7046 880.317
R2151 VSS.n7073 VSS.n758 880.317
R2152 VSS.n7194 VSS.n7193 880.317
R2153 VSS.n7414 VSS.n7413 880.317
R2154 VSS.n7361 VSS.n7255 880.317
R2155 VSS.n7619 VSS.n86 880.317
R2156 VSS.n687 VSS.n686 880.317
R2157 VSS.n7173 VSS.n7172 880.317
R2158 VSS.n7159 VSS.n7158 880.317
R2159 VSS.n7248 VSS.n7247 880.317
R2160 VSS.n6922 VSS.n6921 880.317
R2161 VSS.n7184 VSS.n7183 880.317
R2162 VSS.n7023 VSS.n7022 880.317
R2163 VSS.n903 VSS.n902 880.317
R2164 VSS.n6997 VSS.n6996 880.317
R2165 VSS.n6886 VSS.n6885 880.317
R2166 VSS.n6966 VSS.n6965 880.317
R2167 VSS.n838 VSS.n837 880.317
R2168 VSS.n7715 VSS.n7714 880.317
R2169 VSS.n7683 VSS.n7682 880.317
R2170 VSS.n7651 VSS.n7650 880.317
R2171 VSS.n5560 VSS.n2781 851.542
R2172 VSS.t103 VSS.t83 800.766
R2173 VSS.t76 VSS.t85 800.766
R2174 VSS.t90 VSS.t122 800.766
R2175 VSS.t98 VSS.t96 800.766
R2176 VSS.t47 VSS.t45 800.766
R2177 VSS.t49 VSS.t101 800.766
R2178 VSS.t72 VSS.t288 800.766
R2179 VSS.t40 VSS.t74 800.766
R2180 VSS.t51 VSS.t293 800.766
R2181 VSS.t120 VSS.n2350 800.766
R2182 VSS.n5561 VSS.n2075 745.378
R2183 VSS.n5873 VSS.n5872 745.378
R2184 VSS.n5867 VSS.n5866 745.378
R2185 VSS.n2353 VSS.n2352 708.047
R2186 VSS VSS.n5836 688
R2187 VSS VSS.n5485 688
R2188 VSS.n3313 VSS 688
R2189 VSS VSS.n3302 688
R2190 VSS VSS.n3298 688
R2191 VSS VSS.n1011 688
R2192 VSS.t304 VSS.t291 674.331
R2193 VSS.n6801 VSS.n1000 673.318
R2194 VSS.n6195 VSS.n6076 656.076
R2195 VSS.n6804 VSS.n959 656.076
R2196 VSS.n6714 VSS.n1029 656
R2197 VSS.n2353 VSS 632.184
R2198 VSS.n2350 VSS 623.755
R2199 VSS.n2182 VSS.n2181 617.899
R2200 VSS.n6306 VSS.n6305 617.899
R2201 VSS.n2354 VSS.n2353 613.249
R2202 VSS.n2350 VSS.n2349 613.249
R2203 VSS.t44 VSS 556.322
R2204 VSS.n6252 VSS.n1023 435.765
R2205 VSS.n2215 VSS.n2214 433.748
R2206 VSS.n5877 VSS.n5876 389.642
R2207 VSS.n5875 VSS.n5874 389.642
R2208 VSS.n5871 VSS.n5870 389.642
R2209 VSS.n5869 VSS.n5868 389.642
R2210 VSS.n5865 VSS.n5864 389.642
R2211 VSS.n2259 VSS.n2247 306.625
R2212 VSS.n5895 VSS.n5894 274.635
R2213 VSS.n3064 VSS.n3063 274.635
R2214 VSS VSS.t330 269.733
R2215 VSS.n5588 VSS.n2778 257.318
R2216 VSS.n5879 VSS.n2074 257.318
R2217 VSS.n5944 VSS.n5942 257.318
R2218 VSS.n6741 VSS.n6735 257.318
R2219 VSS.n5911 VSS.n5910 257.318
R2220 VSS.n5905 VSS.n5904 257.318
R2221 VSS.n5900 VSS.n5899 257.318
R2222 VSS.n5892 VSS.n5891 257.318
R2223 VSS.n6245 VSS.n6243 257.318
R2224 VSS.n6744 VSS.n6743 257.318
R2225 VSS.n2953 VSS.n2952 257.318
R2226 VSS.n3276 VSS.n3274 257.318
R2227 VSS.n3074 VSS.n3072 257.318
R2228 VSS.n3030 VSS.n3029 257.318
R2229 VSS.n3052 VSS.n3047 257.318
R2230 VSS.n3061 VSS.n3060 257.318
R2231 VSS.n3058 VSS.n3057 257.318
R2232 VSS.n3055 VSS.n3054 257.318
R2233 VSS.n3077 VSS.n3076 257.318
R2234 VSS.n3018 VSS.n3017 257.318
R2235 VSS.n3034 VSS.n3033 257.318
R2236 VSS.n5559 VSS 257.318
R2237 VSS VSS.n2077 257.318
R2238 VSS VSS.n2081 257.318
R2239 VSS.n5525 VSS 257.318
R2240 VSS VSS.n2097 257.318
R2241 VSS.n5950 VSS.n5949 257.318
R2242 VSS.n5947 VSS.n5946 257.318
R2243 VSS.n5940 VSS.n5939 257.318
R2244 VSS VSS.n5937 257.318
R2245 VSS.n6034 VSS 257.318
R2246 VSS.n6040 VSS 257.318
R2247 VSS.n6046 VSS 257.318
R2248 VSS.n6052 VSS 257.318
R2249 VSS.n2087 VSS.n2086 257.318
R2250 VSS VSS.n2089 257.318
R2251 VSS.n6248 VSS 257.318
R2252 VSS.n5885 VSS 257.318
R2253 VSS.n5587 VSS.n5562 257.318
R2254 VSS.n6605 VSS 240.076
R2255 VSS VSS.n2950 240.076
R2256 VSS VSS.n2804 240.076
R2257 VSS.n2925 VSS 240.076
R2258 VSS.n3310 VSS 240.076
R2259 VSS.n3303 VSS 240.076
R2260 VSS.n3299 VSS 240.076
R2261 VSS.n3295 VSS 240.076
R2262 VSS.n3291 VSS 240.076
R2263 VSS.n6766 VSS 240.076
R2264 VSS.n6777 VSS 240.076
R2265 VSS.n6773 VSS 240.076
R2266 VSS.n2086 VSS 240
R2267 VSS.n6208 VSS.n1932 240
R2268 VSS.n6008 VSS.n6007 240
R2269 VSS VSS.n5940 240
R2270 VSS.n6760 VSS.n1017 240
R2271 VSS.n5950 VSS 240
R2272 VSS.n5910 VSS 240
R2273 VSS.n5904 VSS 240
R2274 VSS.n5899 VSS 240
R2275 VSS VSS.n5892 240
R2276 VSS.n6243 VSS 240
R2277 VSS VSS.n1901 240
R2278 VSS.n6744 VSS 240
R2279 VSS VSS.n1019 240
R2280 VSS VSS.n6741 240
R2281 VSS.n6596 VSS 240
R2282 VSS VSS.n1015 240
R2283 VSS VSS.n1029 240
R2284 VSS VSS.n6715 240
R2285 VSS VSS.n2942 240
R2286 VSS.n3284 VSS.n2944 240
R2287 VSS.n3262 VSS.n3261 240
R2288 VSS VSS.n2953 240
R2289 VSS.n3274 VSS 240
R2290 VSS.n3033 VSS 240
R2291 VSS.n3017 VSS 240
R2292 VSS.n3077 VSS 240
R2293 VSS VSS.n3061 240
R2294 VSS VSS.n2988 240
R2295 VSS VSS.n3058 240
R2296 VSS VSS.n2985 240
R2297 VSS VSS.n3055 240
R2298 VSS VSS.n2982 240
R2299 VSS VSS.n3052 240
R2300 VSS VSS.n2979 240
R2301 VSS.n3117 VSS 240
R2302 VSS.n3107 VSS 240
R2303 VSS.n3098 VSS 240
R2304 VSS.n3089 VSS 240
R2305 VSS.n3081 VSS 240
R2306 VSS VSS.n3074 240
R2307 VSS.n3254 VSS.n2959 240
R2308 VSS VSS.n2959 240
R2309 VSS VSS.n3254 240
R2310 VSS.n3250 VSS.n2966 240
R2311 VSS VSS.n3156 240
R2312 VSS VSS.n2966 240
R2313 VSS VSS.n3250 240
R2314 VSS.n3246 VSS.n2970 240
R2315 VSS.n3192 VSS 240
R2316 VSS VSS.n2970 240
R2317 VSS VSS.n3246 240
R2318 VSS.n3242 VSS.n2974 240
R2319 VSS VSS.n3138 240
R2320 VSS VSS.n2974 240
R2321 VSS VSS.n3242 240
R2322 VSS VSS.n3238 240
R2323 VSS VSS.n3129 240
R2324 VSS.n3238 VSS.n3237 240
R2325 VSS.n3237 VSS 240
R2326 VSS.n3021 VSS 240
R2327 VSS.n3029 VSS 240
R2328 VSS VSS.n2782 240
R2329 VSS VSS.n2784 240
R2330 VSS VSS.n3025 240
R2331 VSS.n5542 VSS.n2789 240
R2332 VSS.n5514 VSS 240
R2333 VSS VSS.n2789 240
R2334 VSS VSS.n5542 240
R2335 VSS VSS.n5538 240
R2336 VSS VSS.n5498 240
R2337 VSS.n5538 VSS.n5537 240
R2338 VSS.n5537 VSS 240
R2339 VSS.n3130 VSS.n3129 240
R2340 VSS VSS.n3130 240
R2341 VSS.n3202 VSS.n3138 240
R2342 VSS.n3202 VSS 240
R2343 VSS.n3192 VSS.n3191 240
R2344 VSS.n3191 VSS 240
R2345 VSS.n3164 VSS.n3156 240
R2346 VSS.n3164 VSS 240
R2347 VSS.n3261 VSS 240
R2348 VSS.n3262 VSS 240
R2349 VSS VSS.n2944 240
R2350 VSS.n3175 VSS.n3174 240
R2351 VSS.n3174 VSS 240
R2352 VSS.n3175 VSS 240
R2353 VSS.n3180 VSS.n3148 240
R2354 VSS.n3180 VSS 240
R2355 VSS VSS.n3148 240
R2356 VSS.n3213 VSS.n3212 240
R2357 VSS.n3212 VSS 240
R2358 VSS.n3213 VSS 240
R2359 VSS.n3224 VSS.n3218 240
R2360 VSS VSS.n3218 240
R2361 VSS VSS.n3224 240
R2362 VSS.n5534 VSS.n2796 240
R2363 VSS.n2796 VSS 240
R2364 VSS VSS.n5534 240
R2365 VSS VSS.n5530 240
R2366 VSS.n5530 VSS.n5529 240
R2367 VSS.n5529 VSS 240
R2368 VSS.n5498 VSS.n5491 240
R2369 VSS VSS.n5491 240
R2370 VSS.n5514 VSS.n5513 240
R2371 VSS.n5513 VSS 240
R2372 VSS.n5554 VSS.n2782 240
R2373 VSS.n5554 VSS 240
R2374 VSS VSS.n3294 240
R2375 VSS.n3284 VSS 240
R2376 VSS.n6760 VSS 240
R2377 VSS.n6755 VSS 240
R2378 VSS VSS.n1022 240
R2379 VSS VSS.n1902 240
R2380 VSS VSS.n2018 240
R2381 VSS VSS.n2070 240
R2382 VSS VSS.n2027 240
R2383 VSS VSS.n2066 240
R2384 VSS VSS.n2047 240
R2385 VSS VSS.n2038 240
R2386 VSS VSS.n2062 240
R2387 VSS.n5957 VSS 240
R2388 VSS.n5965 VSS 240
R2389 VSS.n5918 VSS 240
R2390 VSS VSS.n5947 240
R2391 VSS VSS.n5944 240
R2392 VSS VSS.n5989 240
R2393 VSS.n1953 VSS 240
R2394 VSS VSS.n1957 240
R2395 VSS VSS.n1962 240
R2396 VSS VSS.n5921 240
R2397 VSS VSS.n5979 240
R2398 VSS.n5979 VSS.n5978 240
R2399 VSS.n5978 VSS 240
R2400 VSS.n5965 VSS.n5964 240
R2401 VSS.n5964 VSS 240
R2402 VSS.n2053 VSS 240
R2403 VSS.n2048 VSS 240
R2404 VSS VSS.n6232 240
R2405 VSS VSS.n6228 240
R2406 VSS.n6224 VSS.n1917 240
R2407 VSS.n1988 VSS.n1976 240
R2408 VSS.n1988 VSS 240
R2409 VSS VSS.n1917 240
R2410 VSS VSS.n6224 240
R2411 VSS.n6220 VSS.n1921 240
R2412 VSS VSS.n1974 240
R2413 VSS VSS.n1921 240
R2414 VSS VSS.n6220 240
R2415 VSS.n6216 VSS.n1925 240
R2416 VSS.n6790 VSS 240
R2417 VSS VSS.n1925 240
R2418 VSS VSS.n6216 240
R2419 VSS VSS.n6212 240
R2420 VSS VSS.n1002 240
R2421 VSS.n6212 VSS.n6211 240
R2422 VSS.n6211 VSS 240
R2423 VSS.n6007 VSS 240
R2424 VSS.n6008 VSS 240
R2425 VSS.n6021 VSS.n6019 240
R2426 VSS.n6019 VSS 240
R2427 VSS VSS.n6021 240
R2428 VSS.n1932 VSS 240
R2429 VSS VSS.n6208 240
R2430 VSS VSS.n6204 240
R2431 VSS.n6204 VSS.n6203 240
R2432 VSS.n6203 VSS 240
R2433 VSS.n6795 VSS.n1002 240
R2434 VSS.n6795 VSS 240
R2435 VSS.n6790 VSS.n6789 240
R2436 VSS.n6789 VSS 240
R2437 VSS.n1992 VSS.n1974 240
R2438 VSS.n1992 VSS 240
R2439 VSS.n6028 VSS 240
R2440 VSS.n6056 VSS 240
R2441 VSS VSS.n6196 240
R2442 VSS VSS.n6200 240
R2443 VSS.n6803 VSS 240
R2444 VSS.n6781 VSS 240
R2445 VSS VSS.n6780 240
R2446 VSS VSS.n6776 240
R2447 VSS VSS.n1976 240
R2448 VSS VSS.n1017 240
R2449 VSS.n1909 VSS 240
R2450 VSS.n5879 VSS 240
R2451 VSS.n4608 VSS.n4368 236.089
R2452 VSS.n3895 VSS.n3894 236.089
R2453 VSS.n4291 VSS.n4285 236.089
R2454 VSS.n4654 VSS.n4653 236.089
R2455 VSS.n4362 VSS.n4358 236.089
R2456 VSS.n4202 VSS.n4201 236.089
R2457 VSS.n4920 VSS.n4842 236.089
R2458 VSS.n5152 VSS.n4121 236.089
R2459 VSS.n5138 VSS.n5137 236.089
R2460 VSS.n4819 VSS.n4818 236.089
R2461 VSS.n4685 VSS.n4678 236.089
R2462 VSS.n4736 VSS.n4230 236.089
R2463 VSS.n4722 VSS.n4714 236.089
R2464 VSS.n5200 VSS.n5199 236.089
R2465 VSS.n4255 VSS.n4254 236.089
R2466 VSS.n4029 VSS.n4028 236.089
R2467 VSS.n4007 VSS.n4006 236.089
R2468 VSS.n4080 VSS.n4067 236.089
R2469 VSS.n3982 VSS.n3981 236.089
R2470 VSS.n3964 VSS.n3963 236.089
R2471 VSS.n5259 VSS.n3902 236.089
R2472 VSS.n5765 VSS.n2388 236.089
R2473 VSS.n5733 VSS.n2407 236.089
R2474 VSS.n5701 VSS.n2426 236.089
R2475 VSS.n2566 VSS.n2562 236.089
R2476 VSS.n2602 VSS.n2601 236.089
R2477 VSS.n5617 VSS.n5616 236.089
R2478 VSS.n673 VSS.n672 236.089
R2479 VSS.n6664 VSS.n792 236.089
R2480 VSS.n7067 VSS.n7066 236.089
R2481 VSS.n7084 VSS.n7083 236.089
R2482 VSS.n317 VSS.n314 236.089
R2483 VSS.n655 VSS.n642 236.089
R2484 VSS.n701 VSS.n696 236.089
R2485 VSS.n7369 VSS.n7362 236.089
R2486 VSS.n7613 VSS.n7612 236.089
R2487 VSS.n428 VSS.n427 236.089
R2488 VSS.n7167 VSS.n7112 236.089
R2489 VSS.n7153 VSS.n7140 236.089
R2490 VSS.n6891 VSS.n720 236.089
R2491 VSS.n6915 VSS.n6914 236.089
R2492 VSS.n7181 VSS.n7100 236.089
R2493 VSS.n852 VSS.n847 236.089
R2494 VSS.n896 VSS.n895 236.089
R2495 VSS.n918 VSS.n913 236.089
R2496 VSS.n6879 VSS.n6878 236.089
R2497 VSS.n6959 VSS.n6958 236.089
R2498 VSS.n831 VSS.n830 236.089
R2499 VSS.n7709 VSS.n31 236.089
R2500 VSS.n7677 VSS.n50 236.089
R2501 VSS.n7645 VSS.n69 236.089
R2502 VSS.n5561 VSS.n5560 232.895
R2503 VSS.n5877 VSS.n2075 232.895
R2504 VSS.n5876 VSS.n5875 232.895
R2505 VSS.n5874 VSS.n5873 232.895
R2506 VSS.n5872 VSS.n5871 232.895
R2507 VSS.n5870 VSS.n5869 232.895
R2508 VSS.n5868 VSS.n5867 232.895
R2509 VSS.n5866 VSS.n5865 232.895
R2510 VSS VSS.n2777 225.319
R2511 VSS.n2079 VSS 225.319
R2512 VSS VSS.n5941 225.319
R2513 VSS.n5912 VSS 225.319
R2514 VSS.n5909 VSS 225.319
R2515 VSS.n5903 VSS 225.319
R2516 VSS.n5898 VSS 225.319
R2517 VSS VSS.n5893 225.319
R2518 VSS VSS.n5890 225.319
R2519 VSS VSS.n6244 225.319
R2520 VSS VSS.n6742 225.319
R2521 VSS.n6716 VSS 225.319
R2522 VSS VSS.n2951 225.319
R2523 VSS.n3277 VSS 225.319
R2524 VSS.n3273 VSS 225.319
R2525 VSS.n3031 VSS 225.319
R2526 VSS.n3012 VSS 225.319
R2527 VSS.n3068 VSS 225.319
R2528 VSS VSS.n3062 225.319
R2529 VSS VSS.n3059 225.319
R2530 VSS VSS.n3056 225.319
R2531 VSS VSS.n3053 225.319
R2532 VSS VSS.n3075 225.319
R2533 VSS.n3019 VSS 225.319
R2534 VSS.n3035 VSS 225.319
R2535 VSS VSS.n5558 225.319
R2536 VSS.n2078 VSS 225.319
R2537 VSS.n2088 VSS 225.319
R2538 VSS.n5526 VSS 225.319
R2539 VSS.n5837 VSS 225.319
R2540 VSS.n3305 VSS.n3304 225.319
R2541 VSS VSS.n5948 225.319
R2542 VSS VSS.n5945 225.319
R2543 VSS VSS.n5938 225.319
R2544 VSS VSS.n5936 225.319
R2545 VSS.n6035 VSS 225.319
R2546 VSS.n6041 VSS 225.319
R2547 VSS.n6047 VSS 225.319
R2548 VSS.n6053 VSS 225.319
R2549 VSS.n2090 VSS 225.319
R2550 VSS VSS.n1896 225.319
R2551 VSS.n6249 VSS 225.319
R2552 VSS.n5886 VSS 225.319
R2553 VSS.n5878 VSS 225.319
R2554 VSS.n6595 VSS.n6594 208.076
R2555 VSS.n2949 VSS.n2948 208.076
R2556 VSS.n3293 VSS.n3292 208.076
R2557 VSS.n6779 VSS.n6778 208.076
R2558 VSS.n6775 VSS.n6774 208.076
R2559 VSS VSS.n6739 208
R2560 VSS VSS.n6739 208
R2561 VSS.n6599 VSS 208
R2562 VSS.n6599 VSS 208
R2563 VSS VSS.n3050 208
R2564 VSS VSS.n3050 208
R2565 VSS VSS.n2962 208
R2566 VSS VSS.n2962 208
R2567 VSS VSS.n3252 208
R2568 VSS VSS.n3252 208
R2569 VSS VSS.n3248 208
R2570 VSS VSS.n3248 208
R2571 VSS VSS.n3244 208
R2572 VSS VSS.n3244 208
R2573 VSS VSS.n3240 208
R2574 VSS VSS.n3240 208
R2575 VSS VSS.n3027 208
R2576 VSS VSS.n3027 208
R2577 VSS.n2788 VSS 208
R2578 VSS.n2788 VSS 208
R2579 VSS VSS.n5540 208
R2580 VSS VSS.n5540 208
R2581 VSS.n3264 VSS 208
R2582 VSS.n3264 VSS 208
R2583 VSS.n3152 VSS 208
R2584 VSS.n3152 VSS 208
R2585 VSS.n3178 VSS 208
R2586 VSS.n3178 VSS 208
R2587 VSS VSS.n3134 208
R2588 VSS VSS.n3134 208
R2589 VSS.n3216 VSS 208
R2590 VSS.n3216 VSS 208
R2591 VSS VSS.n3222 208
R2592 VSS VSS.n3222 208
R2593 VSS VSS.n5532 208
R2594 VSS VSS.n5532 208
R2595 VSS.n2803 VSS.n2101 208
R2596 VSS.n2926 VSS.n2806 208
R2597 VSS.n3312 VSS.n3311 208
R2598 VSS.n3301 VSS.n3300 208
R2599 VSS.n3297 VSS.n3296 208
R2600 VSS.n6768 VSS.n6767 208
R2601 VSS VSS.n2068 208
R2602 VSS VSS.n2068 208
R2603 VSS VSS.n2064 208
R2604 VSS VSS.n2064 208
R2605 VSS VSS.n2005 208
R2606 VSS VSS.n2005 208
R2607 VSS VSS.n1961 208
R2608 VSS VSS.n1961 208
R2609 VSS.n1966 VSS 208
R2610 VSS.n1966 VSS 208
R2611 VSS VSS.n6230 208
R2612 VSS VSS.n6230 208
R2613 VSS VSS.n6226 208
R2614 VSS VSS.n6226 208
R2615 VSS VSS.n6222 208
R2616 VSS VSS.n6222 208
R2617 VSS VSS.n6218 208
R2618 VSS VSS.n6218 208
R2619 VSS VSS.n6214 208
R2620 VSS VSS.n6214 208
R2621 VSS VSS.n1955 208
R2622 VSS VSS.n1955 208
R2623 VSS VSS.n6206 208
R2624 VSS VSS.n6206 208
R2625 VSS.n5588 VSS.n5587 208
R2626 VSS.n6317 VSS.n6316 203.197
R2627 VSS.n6721 VSS.t82 199.631
R2628 VSS.n5863 VSS.n5862 169.403
R2629 VSS.t88 VSS 166.407
R2630 VSS.t62 VSS 166.222
R2631 VSS.t302 VSS 151.725
R2632 VSS.t113 VSS 151.556
R2633 VSS.n6256 VSS 149.112
R2634 VSS.n2217 VSS.n2216 140.675
R2635 VSS.n5863 VSS.n5860 137.083
R2636 VSS.n5845 VSS.t316 137.042
R2637 VSS.n6718 VSS.t81 134.445
R2638 VSS.n5864 VSS.n5863 132.845
R2639 VSS.n2172 VSS.t285 122.206
R2640 VSS.n2171 VSS.t286 122.206
R2641 VSS.n5842 VSS.t323 120.749
R2642 VSS.n2180 VSS.n2177 120.749
R2643 VSS.n2156 VSS.n2119 113.834
R2644 VSS.n2144 VSS.n2122 113.834
R2645 VSS.n6289 VSS.n1887 113.834
R2646 VSS.n6277 VSS.n1890 113.834
R2647 VSS.n2039 VSS 112.659
R2648 VSS.n2028 VSS 112.659
R2649 VSS.n2019 VSS 112.659
R2650 VSS VSS.n2071 112.659
R2651 VSS VSS.n6241 112.659
R2652 VSS.n6747 VSS 112.659
R2653 VSS.n2955 VSS 112.659
R2654 VSS VSS.n2994 112.659
R2655 VSS VSS.n3000 112.659
R2656 VSS VSS.n3006 112.659
R2657 VSS.n3116 VSS 112.659
R2658 VSS VSS.n2975 112.659
R2659 VSS.n3106 VSS 112.659
R2660 VSS VSS.n2971 112.659
R2661 VSS.n3097 VSS 112.659
R2662 VSS VSS.n2967 112.659
R2663 VSS.n3088 VSS 112.659
R2664 VSS VSS.n2963 112.659
R2665 VSS.n3080 VSS 112.659
R2666 VSS.n3260 VSS 112.659
R2667 VSS.n3159 VSS 112.659
R2668 VSS.n3142 VSS 112.659
R2669 VSS.n3197 VSS 112.659
R2670 VSS VSS.n3233 112.659
R2671 VSS VSS.n2790 112.659
R2672 VSS.n3122 VSS 112.659
R2673 VSS.n3024 VSS 112.659
R2674 VSS VSS.n3015 112.659
R2675 VSS.n5549 VSS 112.659
R2676 VSS.n5503 VSS 112.659
R2677 VSS.n5519 VSS 112.659
R2678 VSS VSS.n5535 112.659
R2679 VSS VSS.n3127 112.659
R2680 VSS.n3132 VSS 112.659
R2681 VSS.n3232 VSS 112.659
R2682 VSS.n3204 VSS 112.659
R2683 VSS.n3201 VSS 112.659
R2684 VSS.n3144 VSS 112.659
R2685 VSS.n3190 VSS 112.659
R2686 VSS.n3166 VSS 112.659
R2687 VSS.n3163 VSS 112.659
R2688 VSS VSS.n2939 112.659
R2689 VSS VSS.n2936 112.659
R2690 VSS VSS.n2933 112.659
R2691 VSS.n3309 VSS 112.659
R2692 VSS.n2923 VSS 112.659
R2693 VSS VSS.n5486 112.659
R2694 VSS VSS.n5527 112.659
R2695 VSS VSS.n5496 112.659
R2696 VSS.n5524 VSS 112.659
R2697 VSS.n5518 VSS 112.659
R2698 VSS VSS.n5507 112.659
R2699 VSS.n5512 VSS 112.659
R2700 VSS.n5557 VSS 112.659
R2701 VSS.n5553 VSS 112.659
R2702 VSS.n3290 VSS 112.659
R2703 VSS.n3283 VSS 112.659
R2704 VSS.n6765 VSS 112.659
R2705 VSS.n6759 VSS 112.659
R2706 VSS.n6754 VSS 112.659
R2707 VSS.n1907 VSS 112.659
R2708 VSS.n6748 VSS 112.659
R2709 VSS VSS.n6233 112.659
R2710 VSS.n6240 VSS 112.659
R2711 VSS.n2032 VSS 112.659
R2712 VSS.n2043 VSS 112.659
R2713 VSS.n5959 VSS 112.659
R2714 VSS.n5920 VSS 112.659
R2715 VSS.n5952 VSS 112.659
R2716 VSS VSS.n5922 112.659
R2717 VSS VSS.n6022 112.659
R2718 VSS VSS.n5987 112.659
R2719 VSS.n5995 VSS 112.659
R2720 VSS.n5986 VSS 112.659
R2721 VSS.n6006 VSS 112.659
R2722 VSS VSS.n1926 112.659
R2723 VSS.n5968 VSS 112.659
R2724 VSS VSS.n1922 112.659
R2725 VSS.n5963 VSS 112.659
R2726 VSS VSS.n1918 112.659
R2727 VSS.n2052 VSS 112.659
R2728 VSS.n1991 VSS 112.659
R2729 VSS.n1987 VSS 112.659
R2730 VSS.n1970 VSS 112.659
R2731 VSS VSS.n5971 112.659
R2732 VSS.n5998 VSS 112.659
R2733 VSS VSS.n6209 112.659
R2734 VSS.n5997 VSS 112.659
R2735 VSS VSS.n6017 112.659
R2736 VSS.n6039 VSS 112.659
R2737 VSS.n6045 VSS 112.659
R2738 VSS.n6051 VSS 112.659
R2739 VSS VSS.n6201 112.659
R2740 VSS.n1938 VSS 112.659
R2741 VSS VSS.n961 112.659
R2742 VSS.n6794 VSS 112.659
R2743 VSS.n1005 VSS 112.659
R2744 VSS.n6788 VSS 112.659
R2745 VSS VSS.n1008 112.659
R2746 VSS.n6030 VSS 112.659
R2747 VSS.n6027 VSS 112.659
R2748 VSS.n6772 VSS 112.659
R2749 VSS.n1983 VSS 112.659
R2750 VSS VSS.n1911 112.659
R2751 VSS VSS.n2084 112.659
R2752 VSS.n5883 VSS 112.659
R2753 VSS.n6271 VSS.t71 111.925
R2754 VSS.n6265 VSS.t63 111.925
R2755 VSS.n2241 VSS.t121 111.924
R2756 VSS.n2138 VSS.t67 111.924
R2757 VSS.n2132 VSS.t89 111.924
R2758 VSS.n2161 VSS.n2160 108.016
R2759 VSS.n2149 VSS.n2148 108.016
R2760 VSS.n6294 VSS.n6293 108.016
R2761 VSS.n6282 VSS.n6281 108.016
R2762 VSS.n6724 VSS.t79 106.742
R2763 VSS.n6728 VSS.n6727 105.927
R2764 VSS.n2339 VSS.n2338 105.135
R2765 VSS.n2339 VSS.n2337 105.135
R2766 VSS.n2328 VSS.n2327 105.135
R2767 VSS.n2328 VSS.n2326 105.135
R2768 VSS.n2320 VSS.n2319 105.135
R2769 VSS.n2320 VSS.n2318 105.135
R2770 VSS.n2311 VSS.n2310 105.135
R2771 VSS.n2311 VSS.n2309 105.135
R2772 VSS.n2300 VSS.n2299 105.135
R2773 VSS.n2300 VSS.n2298 105.135
R2774 VSS.n2292 VSS.n2291 105.135
R2775 VSS.n2292 VSS.n2290 105.135
R2776 VSS.n2283 VSS.n2282 105.135
R2777 VSS.n2283 VSS.n2281 105.135
R2778 VSS.n2272 VSS.n2271 105.135
R2779 VSS.n2272 VSS.n2270 105.135
R2780 VSS.n2264 VSS.n2263 105.135
R2781 VSS.n2264 VSS.n2262 105.135
R2782 VSS.n2348 VSS.t292 104.666
R2783 VSS.n2344 VSS.t305 104.666
R2784 VSS.n2117 VSS.t317 103.507
R2785 VSS.n2120 VSS.t303 103.507
R2786 VSS.n1886 VSS.t54 103.507
R2787 VSS.n1888 VSS.t114 103.507
R2788 VSS.n5855 VSS.t66 101.15
R2789 VSS.n2177 VSS.n2176 91.3782
R2790 VSS.n2131 VSS.n2130 89.977
R2791 VSS.n6264 VSS.n6263 89.977
R2792 VSS.n7646 VSS.n7645 84.2672
R2793 VSS.n7678 VSS.n7677 84.2672
R2794 VSS.n7710 VSS.n7709 84.2672
R2795 VSS.n5702 VSS.n5701 84.2672
R2796 VSS.n5734 VSS.n5733 84.2672
R2797 VSS.n5766 VSS.n5765 84.2672
R2798 VSS.n4453 VSS.n4358 84.2672
R2799 VSS.n4408 VSS.n4368 84.2672
R2800 VSS.n4612 VSS.n4608 84.2672
R2801 VSS.n4608 VSS.n4607 84.2672
R2802 VSS.n4368 VSS.n4366 84.2672
R2803 VSS.n3894 VSS.n3888 84.2672
R2804 VSS.n5269 VSS.n3895 84.2672
R2805 VSS.n4299 VSS.n3895 84.2672
R2806 VSS.n4285 VSS.n4282 84.2672
R2807 VSS.n4344 VSS.n4291 84.2672
R2808 VSS.n4291 VSS.n4290 84.2672
R2809 VSS.n4316 VSS.n4285 84.2672
R2810 VSS.n4653 VSS.n4271 84.2672
R2811 VSS.n4654 VSS.n4259 84.2672
R2812 VSS.n4654 VSS.n4270 84.2672
R2813 VSS.n4623 VSS.n4362 84.2672
R2814 VSS.n4404 VSS.n4362 84.2672
R2815 VSS.n4358 VSS.n4356 84.2672
R2816 VSS.n4957 VSS.n4202 84.2672
R2817 VSS.n4372 VSS.n4202 84.2672
R2818 VSS.n4201 VSS.n4195 84.2672
R2819 VSS.n4842 VSS.n4747 84.2672
R2820 VSS.n4842 VSS.n4841 84.2672
R2821 VSS.n4920 VSS.n4919 84.2672
R2822 VSS.n5153 VSS.n5152 84.2672
R2823 VSS.n4121 VSS.n4118 84.2672
R2824 VSS.n4912 VSS.n4121 84.2672
R2825 VSS.n5137 VSS.n4127 84.2672
R2826 VSS.n5140 VSS.n5138 84.2672
R2827 VSS.n5138 VSS.n5136 84.2672
R2828 VSS.n4818 VSS.n4806 84.2672
R2829 VSS.n4828 VSS.n4819 84.2672
R2830 VSS.n4819 VSS.n4817 84.2672
R2831 VSS.n4686 VSS.n4685 84.2672
R2832 VSS.n4678 VSS.n4234 84.2672
R2833 VSS.n4678 VSS.n4235 84.2672
R2834 VSS.n4737 VSS.n4736 84.2672
R2835 VSS.n4694 VSS.n4230 84.2672
R2836 VSS.n4230 VSS.n4229 84.2672
R2837 VSS.n4723 VSS.n4722 84.2672
R2838 VSS.n4714 VSS.n4703 84.2672
R2839 VSS.n4714 VSS.n4713 84.2672
R2840 VSS.n5199 VSS.n4102 84.2672
R2841 VSS.n5202 VSS.n5200 84.2672
R2842 VSS.n5200 VSS.n5198 84.2672
R2843 VSS.n4254 VSS.n4253 84.2672
R2844 VSS.n4661 VSS.n4255 84.2672
R2845 VSS.n4263 VSS.n4255 84.2672
R2846 VSS.n4037 VSS.n4029 84.2672
R2847 VSS.n4029 VSS.n4018 84.2672
R2848 VSS.n4028 VSS.n4027 84.2672
R2849 VSS.n4050 VSS.n4007 84.2672
R2850 VSS.n4020 VSS.n4007 84.2672
R2851 VSS.n4006 VSS.n4005 84.2672
R2852 VSS.n4081 VSS.n4080 84.2672
R2853 VSS.n4067 VSS.n3986 84.2672
R2854 VSS.n4067 VSS.n3987 84.2672
R2855 VSS.n3981 VSS.n3980 84.2672
R2856 VSS.n4089 VSS.n3982 84.2672
R2857 VSS.n4070 VSS.n3982 84.2672
R2858 VSS.n3963 VSS.n3946 84.2672
R2859 VSS.n3966 VSS.n3964 84.2672
R2860 VSS.n3964 VSS.n3962 84.2672
R2861 VSS.n5259 VSS.n5258 84.2672
R2862 VSS.n3903 VSS.n3902 84.2672
R2863 VSS.n4295 VSS.n3902 84.2672
R2864 VSS.n2388 VSS.n2385 84.2672
R2865 VSS.n3955 VSS.n2388 84.2672
R2866 VSS.n2407 VSS.n2404 84.2672
R2867 VSS.n5191 VSS.n2407 84.2672
R2868 VSS.n2426 VSS.n2423 84.2672
R2869 VSS.n5129 VSS.n2426 84.2672
R2870 VSS.n5616 VSS.n2512 84.2672
R2871 VSS.n2601 VSS.n2600 84.2672
R2872 VSS.n2567 VSS.n2566 84.2672
R2873 VSS.n2578 VSS.n2562 84.2672
R2874 VSS.n2562 VSS.n2561 84.2672
R2875 VSS.n2602 VSS.n2532 84.2672
R2876 VSS.n2602 VSS.n2536 84.2672
R2877 VSS.n5617 VSS.n2511 84.2672
R2878 VSS.n5618 VSS.n5617 84.2672
R2879 VSS.n314 VSS.n311 84.2672
R2880 VSS.n672 VSS.n532 84.2672
R2881 VSS.n674 VSS.n673 84.2672
R2882 VSS.n673 VSS.n531 84.2672
R2883 VSS.n656 VSS.n655 84.2672
R2884 VSS.n6665 VSS.n6664 84.2672
R2885 VSS.n7042 VSS.n792 84.2672
R2886 VSS.n822 VSS.n792 84.2672
R2887 VSS.n7066 VSS.n781 84.2672
R2888 VSS.n7069 VSS.n7067 84.2672
R2889 VSS.n7067 VSS.n760 84.2672
R2890 VSS.n7066 VSS.n7065 84.2672
R2891 VSS.n7083 VSS.n753 84.2672
R2892 VSS.n7191 VSS.n7084 84.2672
R2893 VSS.n7091 VSS.n7084 84.2672
R2894 VSS.n7453 VSS.n317 84.2672
R2895 VSS.n645 VSS.n317 84.2672
R2896 VSS.n764 VSS.n314 84.2672
R2897 VSS.n642 VSS.n641 84.2672
R2898 VSS.n642 VSS.n628 84.2672
R2899 VSS.n696 VSS.n341 84.2672
R2900 VSS.n696 VSS.n695 84.2672
R2901 VSS.n7259 VSS.n701 84.2672
R2902 VSS.n7370 VSS.n7369 84.2672
R2903 VSS.n7362 VSS.n7256 84.2672
R2904 VSS.n7362 VSS.n7257 84.2672
R2905 VSS.n7612 VSS.n89 84.2672
R2906 VSS.n7615 VSS.n7613 84.2672
R2907 VSS.n7613 VSS.n88 84.2672
R2908 VSS.n427 VSS.n418 84.2672
R2909 VSS.n682 VSS.n428 84.2672
R2910 VSS.n433 VSS.n428 84.2672
R2911 VSS.n7168 VSS.n7167 84.2672
R2912 VSS.n7120 VSS.n7112 84.2672
R2913 VSS.n7112 VSS.n7111 84.2672
R2914 VSS.n7154 VSS.n7153 84.2672
R2915 VSS.n7140 VSS.n7133 84.2672
R2916 VSS.n7140 VSS.n7139 84.2672
R2917 VSS.n6892 VSS.n6891 84.2672
R2918 VSS.n7243 VSS.n720 84.2672
R2919 VSS.n7143 VSS.n720 84.2672
R2920 VSS.n6914 VSS.n6897 84.2672
R2921 VSS.n6917 VSS.n6915 84.2672
R2922 VSS.n6915 VSS.n6913 84.2672
R2923 VSS.n7181 VSS.n7180 84.2672
R2924 VSS.n7101 VSS.n7100 84.2672
R2925 VSS.n7100 VSS.n7099 84.2672
R2926 VSS.n847 VSS.n808 84.2672
R2927 VSS.n847 VSS.n846 84.2672
R2928 VSS.n886 VSS.n852 84.2672
R2929 VSS.n898 VSS.n896 84.2672
R2930 VSS.n896 VSS.n894 84.2672
R2931 VSS.n895 VSS.n877 84.2672
R2932 VSS.n913 VSS.n873 84.2672
R2933 VSS.n913 VSS.n912 84.2672
R2934 VSS.n6867 VSS.n918 84.2672
R2935 VSS.n6878 VSS.n6877 84.2672
R2936 VSS.n6881 VSS.n6879 84.2672
R2937 VSS.n6879 VSS.n6874 84.2672
R2938 VSS.n6958 VSS.n6857 84.2672
R2939 VSS.n6961 VSS.n6959 84.2672
R2940 VSS.n6959 VSS.n6957 84.2672
R2941 VSS.n830 VSS.n813 84.2672
R2942 VSS.n833 VSS.n831 84.2672
R2943 VSS.n831 VSS.n829 84.2672
R2944 VSS.n31 VSS.n28 84.2672
R2945 VSS.n6950 VSS.n31 84.2672
R2946 VSS.n50 VSS.n47 84.2672
R2947 VSS.n6906 VSS.n50 84.2672
R2948 VSS.n69 VSS.n66 84.2672
R2949 VSS.n80 VSS.n69 84.2672
R2950 VSS.n5839 VSS.t322 84.0354
R2951 VSS.n5860 VSS 82.3883
R2952 VSS.n2098 VSS.t325 70.1655
R2953 VSS.t64 VSS.t300 68.5211
R2954 VSS.t300 VSS.t296 68.5211
R2955 VSS.t331 VSS.t310 68.5211
R2956 VSS.t314 VSS.t312 68.5211
R2957 VSS.t68 VSS.t111 68.4449
R2958 VSS.t111 VSS.t115 68.4449
R2959 VSS.t117 VSS.t113 68.4449
R2960 VSS.t55 VSS.t59 68.4449
R2961 VSS.t53 VSS.t57 68.4449
R2962 VSS.n2227 VSS.n2226 66.4303
R2963 VSS.n5855 VSS 66.0739
R2964 VSS.t296 VSS.n5854 66.0739
R2965 VSS.n6721 VSS.t80 62.7412
R2966 VSS.n2098 VSS.t327 58.7433
R2967 VSS VSS.t88 58.7324
R2968 VSS.t66 VSS 58.7324
R2969 VSS VSS.t62 58.6672
R2970 VSS VSS.t70 58.6672
R2971 VSS.n6257 VSS.n6254 57.8524
R2972 VSS.t329 VSS.n5838 53.0322
R2973 VSS.n6734 VSS.n1024 50.519
R2974 VSS.n6305 VSS.n6304 48.0746
R2975 VSS.n2338 VSS.t308 45.7148
R2976 VSS.n2337 VSS.t294 45.7148
R2977 VSS.n2327 VSS.t75 45.7148
R2978 VSS.n2326 VSS.t287 45.7148
R2979 VSS.n2319 VSS.t290 45.7148
R2980 VSS.n2318 VSS.t289 45.7148
R2981 VSS.n2310 VSS.t309 45.7148
R2982 VSS.n2309 VSS.t102 45.7148
R2983 VSS.n2299 VSS.t100 45.7148
R2984 VSS.n2298 VSS.t46 45.7148
R2985 VSS.n2291 VSS.t97 45.7148
R2986 VSS.n2290 VSS.t119 45.7148
R2987 VSS.n2282 VSS.t123 45.7148
R2988 VSS.n2281 VSS.t321 45.7148
R2989 VSS.n2271 VSS.t86 45.7148
R2990 VSS.n2270 VSS.t284 45.7148
R2991 VSS.n2263 VSS.t84 45.7148
R2992 VSS.n2262 VSS.t95 45.7148
R2993 VSS.n5839 VSS.t329 44.8735
R2994 VSS.n2259 VSS.n2258 44.424
R2995 VSS.t310 VSS.n5851 43.2337
R2996 VSS.n2173 VSS.n2172 41.6396
R2997 VSS.n6733 VSS.t55 39.9264
R2998 VSS.n2181 VSS.n2180 39.1624
R2999 VSS.n6318 VSS.n6315 38.9511
R3000 VSS.n5853 VSS.t302 38.3394
R3001 VSS.n2169 VSS.t328 34.9023
R3002 VSS.n2173 VSS.t326 34.8109
R3003 VSS.n2316 VSS.n2315 34.6358
R3004 VSS.n2288 VSS.n2287 34.6358
R3005 VSS.n2155 VSS.n2154 34.6358
R3006 VSS.n2143 VSS.n2142 34.6358
R3007 VSS.n2137 VSS.n2123 34.6358
R3008 VSS.n6288 VSS.n1889 34.6358
R3009 VSS.n6276 VSS.n1891 34.6358
R3010 VSS.n6270 VSS.n1892 34.6358
R3011 VSS.n6594 VSS 34.5605
R3012 VSS.n6605 VSS 34.5605
R3013 VSS.n2950 VSS 34.5605
R3014 VSS.n2948 VSS 34.5605
R3015 VSS.n2804 VSS 34.5605
R3016 VSS.n2925 VSS 34.5605
R3017 VSS.n3310 VSS 34.5605
R3018 VSS.n3303 VSS 34.5605
R3019 VSS.n3299 VSS 34.5605
R3020 VSS.n3295 VSS 34.5605
R3021 VSS.n3293 VSS 34.5605
R3022 VSS.n3291 VSS 34.5605
R3023 VSS.n6766 VSS 34.5605
R3024 VSS.n6076 VSS 34.5605
R3025 VSS.n959 VSS 34.5605
R3026 VSS.n6779 VSS 34.5605
R3027 VSS.n6777 VSS 34.5605
R3028 VSS.n6775 VSS 34.5605
R3029 VSS.n6773 VSS 34.5605
R3030 VSS.n2338 VSS.t319 34.506
R3031 VSS.n2337 VSS.t52 34.506
R3032 VSS.n2327 VSS.t61 34.506
R3033 VSS.n2326 VSS.t41 34.506
R3034 VSS.n2319 VSS.t73 34.506
R3035 VSS.n2318 VSS.t109 34.506
R3036 VSS.n2310 VSS.t50 34.506
R3037 VSS.n2309 VSS.t295 34.506
R3038 VSS.n2299 VSS.t48 34.506
R3039 VSS.n2298 VSS.t78 34.506
R3040 VSS.n2291 VSS.t99 34.506
R3041 VSS.n2290 VSS.t318 34.506
R3042 VSS.n2282 VSS.t320 34.506
R3043 VSS.n2281 VSS.t91 34.506
R3044 VSS.n2271 VSS.t77 34.506
R3045 VSS.n2270 VSS.t87 34.506
R3046 VSS.n2263 VSS.t104 34.506
R3047 VSS.n2262 VSS.t110 34.506
R3048 VSS.t330 VSS.t304 33.717
R3049 VSS.t291 VSS.t44 33.717
R3050 VSS.n6728 VSS.t53 30.9635
R3051 VSS.t298 VSS.n5853 30.1822
R3052 VSS.n6726 VSS.n6723 28.5997
R3053 VSS.t306 VSS.n6733 28.519
R3054 VSS.n2218 VSS.n2213 26.9663
R3055 VSS.n5846 VSS.n5845 26.9193
R3056 VSS.n5851 VSS.t314 25.2879
R3057 VSS.n2160 VSS.t315 24.9236
R3058 VSS.n2160 VSS.t313 24.9236
R3059 VSS.n2119 VSS.t332 24.9236
R3060 VSS.n2119 VSS.t311 24.9236
R3061 VSS.n2148 VSS.t297 24.9236
R3062 VSS.n2148 VSS.t299 24.9236
R3063 VSS.n2122 VSS.t65 24.9236
R3064 VSS.n2122 VSS.t301 24.9236
R3065 VSS.n6293 VSS.t60 24.9236
R3066 VSS.n6293 VSS.t58 24.9236
R3067 VSS.n1887 VSS.t307 24.9236
R3068 VSS.n1887 VSS.t56 24.9236
R3069 VSS.n6281 VSS.t116 24.9236
R3070 VSS.n6281 VSS.t118 24.9236
R3071 VSS.n1890 VSS.t69 24.9236
R3072 VSS.n1890 VSS.t112 24.9236
R3073 VSS.n5858 VSS.n2095 24.921
R3074 VSS VSS.t64 24.4721
R3075 VSS VSS.t331 24.4721
R3076 VSS.n6257 VSS 24.4449
R3077 VSS VSS.t68 24.4449
R3078 VSS VSS.t306 24.4449
R3079 VSS.n2170 VSS.n2169 24.0738
R3080 VSS.n2354 VSS.n2240 23.7181
R3081 VSS.n2349 VSS.n2242 23.7181
R3082 VSS.n2344 VSS.n2343 23.7181
R3083 VSS.n2260 VSS.n2259 23.7181
R3084 VSS.n2167 VSS.n2166 23.7181
R3085 VSS.n6300 VSS.n6299 23.7181
R3086 VSS.n2187 VSS.n2186 23.4463
R3087 VSS.n2216 VSS.n2215 23.4463
R3088 VSS.n2345 VSS.n2344 22.2123
R3089 VSS.n6289 VSS.n6288 22.2123
R3090 VSS.n6277 VSS.n6276 22.2123
R3091 VSS.n6259 VSS.n1894 21.4231
R3092 VSS.n1894 VSS.n1026 21.4231
R3093 VSS.n6731 VSS.n1026 21.4231
R3094 VSS.n6723 VSS.n6720 21.4231
R3095 VSS.n6720 VSS.n1027 21.4231
R3096 VSS.n5858 VSS.n5857 20.3989
R3097 VSS.n5857 VSS.n2096 20.3989
R3098 VSS.n5849 VSS.n2096 20.3989
R3099 VSS.n5849 VSS.n5848 20.3989
R3100 VSS.n5848 VSS.n5844 20.3989
R3101 VSS.n5844 VSS.n5841 20.3989
R3102 VSS.n5841 VSS.n2100 20.3989
R3103 VSS.n2178 VSS.n2100 20.3989
R3104 VSS.n2207 VSS.n2204 19.3944
R3105 VSS.n1884 VSS.n1881 19.3944
R3106 VSS.n2178 VSS.n2116 19.0674
R3107 VSS.n5589 VSS 18.3101
R3108 VSS VSS.n5585 18.3101
R3109 VSS.n6731 VSS.n6730 18.1561
R3110 VSS.t70 VSS.n6256 17.9264
R3111 VSS.n2129 VSS.n2126 17.7168
R3112 VSS.n2257 VSS.n2251 17.7168
R3113 VSS.n2251 VSS.n1893 17.7168
R3114 VSS.n1870 VSS.n1869 17.649
R3115 VSS.n6730 VSS.n6726 17.5135
R3116 VSS.n2778 VSS 17.3181
R3117 VSS.n2777 VSS 17.3181
R3118 VSS VSS.n2079 17.3181
R3119 VSS VSS.n2074 17.3181
R3120 VSS.n5941 VSS 17.3181
R3121 VSS.n5942 VSS 17.3181
R3122 VSS.n5912 VSS 17.3181
R3123 VSS VSS.n5911 17.3181
R3124 VSS VSS.n5909 17.3181
R3125 VSS.n5905 VSS 17.3181
R3126 VSS VSS.n5903 17.3181
R3127 VSS.n5900 VSS 17.3181
R3128 VSS VSS.n5898 17.3181
R3129 VSS.n5895 VSS 17.3181
R3130 VSS.n5894 VSS 17.3181
R3131 VSS.n5893 VSS 17.3181
R3132 VSS.n5891 VSS 17.3181
R3133 VSS.n5890 VSS 17.3181
R3134 VSS.n6245 VSS 17.3181
R3135 VSS.n6244 VSS 17.3181
R3136 VSS.n6743 VSS 17.3181
R3137 VSS.n6742 VSS 17.3181
R3138 VSS.n6716 VSS 17.3181
R3139 VSS.n6735 VSS 17.3181
R3140 VSS.n2952 VSS 17.3181
R3141 VSS.n2951 VSS 17.3181
R3142 VSS.n3277 VSS 17.3181
R3143 VSS VSS.n3276 17.3181
R3144 VSS VSS.n3273 17.3181
R3145 VSS.n3072 VSS 17.3181
R3146 VSS VSS.n3031 17.3181
R3147 VSS VSS.n3030 17.3181
R3148 VSS VSS.n3012 17.3181
R3149 VSS.n3047 VSS 17.3181
R3150 VSS VSS.n3068 17.3181
R3151 VSS.n3064 VSS 17.3181
R3152 VSS.n3063 VSS 17.3181
R3153 VSS.n3062 VSS 17.3181
R3154 VSS.n3060 VSS 17.3181
R3155 VSS.n3059 VSS 17.3181
R3156 VSS.n3057 VSS 17.3181
R3157 VSS.n3056 VSS 17.3181
R3158 VSS.n3054 VSS 17.3181
R3159 VSS.n3053 VSS 17.3181
R3160 VSS.n3076 VSS 17.3181
R3161 VSS.n3075 VSS 17.3181
R3162 VSS VSS.n3018 17.3181
R3163 VSS VSS.n3019 17.3181
R3164 VSS VSS.n3034 17.3181
R3165 VSS.n3035 VSS 17.3181
R3166 VSS.n5559 VSS 17.3181
R3167 VSS.n5558 VSS 17.3181
R3168 VSS VSS.n2077 17.3181
R3169 VSS VSS.n2078 17.3181
R3170 VSS VSS.n2081 17.3181
R3171 VSS VSS.n2088 17.3181
R3172 VSS VSS.n5525 17.3181
R3173 VSS VSS.n5526 17.3181
R3174 VSS VSS.n2097 17.3181
R3175 VSS.n5837 VSS 17.3181
R3176 VSS.n5949 VSS 17.3181
R3177 VSS.n5948 VSS 17.3181
R3178 VSS.n5946 VSS 17.3181
R3179 VSS.n5945 VSS 17.3181
R3180 VSS.n5939 VSS 17.3181
R3181 VSS.n5938 VSS 17.3181
R3182 VSS.n5937 VSS 17.3181
R3183 VSS.n5936 VSS 17.3181
R3184 VSS VSS.n6034 17.3181
R3185 VSS.n6035 VSS 17.3181
R3186 VSS VSS.n6040 17.3181
R3187 VSS.n6041 VSS 17.3181
R3188 VSS VSS.n6046 17.3181
R3189 VSS.n6047 VSS 17.3181
R3190 VSS VSS.n6052 17.3181
R3191 VSS.n6053 VSS 17.3181
R3192 VSS VSS.n2087 17.3181
R3193 VSS.n2090 VSS 17.3181
R3194 VSS.n2089 VSS 17.3181
R3195 VSS VSS.n1896 17.3181
R3196 VSS.n6249 VSS 17.3181
R3197 VSS VSS.n6248 17.3181
R3198 VSS.n5886 VSS 17.3181
R3199 VSS VSS.n5885 17.3181
R3200 VSS VSS.n5878 17.3181
R3201 VSS.n5562 VSS 17.3181
R3202 VSS VSS.n2908 17.2429
R3203 VSS VSS.n6802 17.2429
R3204 VSS.n6263 VSS.n6262 16.8752
R3205 VSS.n1869 VSS.n1027 16.2614
R3206 VSS.n1885 VSS.n1884 15.952
R3207 VSS.n2208 VSS.n2207 15.7581
R3208 VSS.t115 VSS.n1024 15.482
R3209 VSS.n2156 VSS 15.4358
R3210 VSS.n2144 VSS 15.4358
R3211 VSS.n2196 VSS.n2116 14.4975
R3212 VSS.n2130 VSS.n2095 14.395
R3213 VSS.n2223 VSS.n2221 14.2324
R3214 VSS.n2349 VSS.n2348 12.8005
R3215 VSS.n6262 VSS.n6259 12.2814
R3216 VSS.t81 VSS.n6717 10.5931
R3217 VSS.n2242 VSS.n2241 10.5417
R3218 VSS.n2139 VSS.n2138 10.5417
R3219 VSS.n2133 VSS.n2132 10.5417
R3220 VSS.n6272 VSS.n6271 10.5417
R3221 VSS.n6266 VSS.n6265 10.5417
R3222 VSS.n2174 VSS.n2173 10.2904
R3223 VSS.n5910 VSS.n2009 8.65932
R3224 VSS VSS.n2009 8.65932
R3225 VSS.n5904 VSS.n2011 8.65932
R3226 VSS VSS.n2011 8.65932
R3227 VSS.n5899 VSS.n2013 8.65932
R3228 VSS VSS.n2013 8.65932
R3229 VSS.n5892 VSS.n2072 8.65932
R3230 VSS.n2072 VSS 8.65932
R3231 VSS.n6241 VSS 8.65932
R3232 VSS.n6243 VSS.n6242 8.65932
R3233 VSS.n6242 VSS 8.65932
R3234 VSS VSS.n6747 8.65932
R3235 VSS.n6746 VSS.n6744 8.65932
R3236 VSS VSS.n6746 8.65932
R3237 VSS.n6741 VSS.n6740 8.65932
R3238 VSS.n6740 VSS 8.65932
R3239 VSS.n6739 VSS.n6738 8.65932
R3240 VSS.n6738 VSS 8.65932
R3241 VSS.n6598 VSS.n6596 8.65932
R3242 VSS VSS.n6598 8.65932
R3243 VSS.n6604 VSS.n6599 8.65932
R3244 VSS VSS.n6604 8.65932
R3245 VSS.n3274 VSS.n2954 8.65932
R3246 VSS VSS.n2954 8.65932
R3247 VSS.n2994 VSS 8.65932
R3248 VSS.n3061 VSS.n2995 8.65932
R3249 VSS.n2995 VSS 8.65932
R3250 VSS.n3000 VSS 8.65932
R3251 VSS.n3058 VSS.n3001 8.65932
R3252 VSS.n3001 VSS 8.65932
R3253 VSS.n3006 VSS 8.65932
R3254 VSS.n3055 VSS.n3007 8.65932
R3255 VSS.n3007 VSS 8.65932
R3256 VSS.n3052 VSS.n3051 8.65932
R3257 VSS.n3051 VSS 8.65932
R3258 VSS.n3050 VSS.n3049 8.65932
R3259 VSS.n3049 VSS 8.65932
R3260 VSS VSS.n3116 8.65932
R3261 VSS.n3114 VSS.n2979 8.65932
R3262 VSS VSS.n3114 8.65932
R3263 VSS.n3108 VSS.n3107 8.65932
R3264 VSS.n3108 VSS 8.65932
R3265 VSS VSS.n3106 8.65932
R3266 VSS.n3105 VSS.n2982 8.65932
R3267 VSS VSS.n3105 8.65932
R3268 VSS.n3099 VSS.n3098 8.65932
R3269 VSS.n3099 VSS 8.65932
R3270 VSS VSS.n3097 8.65932
R3271 VSS.n3096 VSS.n2985 8.65932
R3272 VSS VSS.n3096 8.65932
R3273 VSS.n3090 VSS.n3089 8.65932
R3274 VSS.n3090 VSS 8.65932
R3275 VSS VSS.n3088 8.65932
R3276 VSS.n3087 VSS.n2988 8.65932
R3277 VSS VSS.n3087 8.65932
R3278 VSS.n3082 VSS.n3081 8.65932
R3279 VSS.n3082 VSS 8.65932
R3280 VSS VSS.n3080 8.65932
R3281 VSS.n3079 VSS.n3077 8.65932
R3282 VSS VSS.n3079 8.65932
R3283 VSS.n3074 VSS.n3073 8.65932
R3284 VSS.n3073 VSS 8.65932
R3285 VSS.n3259 VSS.n2959 8.65932
R3286 VSS VSS.n3259 8.65932
R3287 VSS.n3255 VSS.n2962 8.65932
R3288 VSS.n3255 VSS 8.65932
R3289 VSS VSS.n2963 8.65932
R3290 VSS.n3254 VSS.n3253 8.65932
R3291 VSS.n3253 VSS 8.65932
R3292 VSS.n3159 VSS 8.65932
R3293 VSS.n3158 VSS.n2966 8.65932
R3294 VSS VSS.n3158 8.65932
R3295 VSS.n3252 VSS.n3251 8.65932
R3296 VSS.n3251 VSS 8.65932
R3297 VSS VSS.n2967 8.65932
R3298 VSS.n3250 VSS.n3249 8.65932
R3299 VSS.n3249 VSS 8.65932
R3300 VSS.n3142 VSS 8.65932
R3301 VSS.n3141 VSS.n2970 8.65932
R3302 VSS VSS.n3141 8.65932
R3303 VSS.n3248 VSS.n3247 8.65932
R3304 VSS.n3247 VSS 8.65932
R3305 VSS VSS.n2971 8.65932
R3306 VSS.n3246 VSS.n3245 8.65932
R3307 VSS.n3245 VSS 8.65932
R3308 VSS.n3197 VSS 8.65932
R3309 VSS.n3196 VSS.n2974 8.65932
R3310 VSS VSS.n3196 8.65932
R3311 VSS.n3244 VSS.n3243 8.65932
R3312 VSS.n3243 VSS 8.65932
R3313 VSS VSS.n2975 8.65932
R3314 VSS.n3242 VSS.n3241 8.65932
R3315 VSS.n3241 VSS 8.65932
R3316 VSS.n3240 VSS.n3239 8.65932
R3317 VSS.n3239 VSS 8.65932
R3318 VSS.n3233 VSS 8.65932
R3319 VSS.n3238 VSS.n3234 8.65932
R3320 VSS.n3234 VSS 8.65932
R3321 VSS.n3237 VSS.n3236 8.65932
R3322 VSS.n3236 VSS 8.65932
R3323 VSS VSS.n3122 8.65932
R3324 VSS.n3118 VSS.n3117 8.65932
R3325 VSS.n3118 VSS 8.65932
R3326 VSS.n3023 VSS.n3021 8.65932
R3327 VSS VSS.n3023 8.65932
R3328 VSS.n3015 VSS 8.65932
R3329 VSS.n3017 VSS.n3016 8.65932
R3330 VSS.n3016 VSS 8.65932
R3331 VSS.n3029 VSS.n3028 8.65932
R3332 VSS.n3028 VSS 8.65932
R3333 VSS.n5549 VSS 8.65932
R3334 VSS.n5548 VSS.n2784 8.65932
R3335 VSS VSS.n5548 8.65932
R3336 VSS.n3027 VSS.n3026 8.65932
R3337 VSS.n3026 VSS 8.65932
R3338 VSS VSS.n3024 8.65932
R3339 VSS.n3025 VSS.n2787 8.65932
R3340 VSS VSS.n2787 8.65932
R3341 VSS.n5503 VSS 8.65932
R3342 VSS.n5502 VSS.n2789 8.65932
R3343 VSS VSS.n5502 8.65932
R3344 VSS.n5543 VSS.n2788 8.65932
R3345 VSS.n5543 VSS 8.65932
R3346 VSS VSS.n2790 8.65932
R3347 VSS.n5542 VSS.n5541 8.65932
R3348 VSS.n5541 VSS 8.65932
R3349 VSS.n5540 VSS.n5539 8.65932
R3350 VSS.n5539 VSS 8.65932
R3351 VSS.n5519 VSS 8.65932
R3352 VSS.n5538 VSS.n2793 8.65932
R3353 VSS VSS.n2793 8.65932
R3354 VSS.n5537 VSS.n5536 8.65932
R3355 VSS.n5536 VSS 8.65932
R3356 VSS.n3127 VSS 8.65932
R3357 VSS.n3129 VSS.n3128 8.65932
R3358 VSS.n3128 VSS 8.65932
R3359 VSS.n3131 VSS.n3130 8.65932
R3360 VSS VSS.n3131 8.65932
R3361 VSS VSS.n3232 8.65932
R3362 VSS.n3138 VSS.n3137 8.65932
R3363 VSS.n3137 VSS 8.65932
R3364 VSS.n3203 VSS.n3202 8.65932
R3365 VSS VSS.n3203 8.65932
R3366 VSS VSS.n3201 8.65932
R3367 VSS.n3194 VSS.n3192 8.65932
R3368 VSS VSS.n3194 8.65932
R3369 VSS.n3191 VSS.n3139 8.65932
R3370 VSS VSS.n3139 8.65932
R3371 VSS VSS.n3190 8.65932
R3372 VSS.n3156 VSS.n3155 8.65932
R3373 VSS.n3155 VSS 8.65932
R3374 VSS.n3165 VSS.n3164 8.65932
R3375 VSS VSS.n3165 8.65932
R3376 VSS VSS.n3163 8.65932
R3377 VSS.n3261 VSS.n2958 8.65932
R3378 VSS VSS.n2958 8.65932
R3379 VSS VSS.n3260 8.65932
R3380 VSS VSS.n2955 8.65932
R3381 VSS.n3263 VSS.n3262 8.65932
R3382 VSS VSS.n3263 8.65932
R3383 VSS.n3265 VSS.n3264 8.65932
R3384 VSS.n3265 VSS 8.65932
R3385 VSS.n3151 VSS.n2944 8.65932
R3386 VSS VSS.n3151 8.65932
R3387 VSS.n3174 VSS.n3149 8.65932
R3388 VSS.n3149 VSS 8.65932
R3389 VSS.n3173 VSS.n3152 8.65932
R3390 VSS VSS.n3173 8.65932
R3391 VSS.n3166 VSS 8.65932
R3392 VSS.n3177 VSS.n3175 8.65932
R3393 VSS VSS.n3177 8.65932
R3394 VSS.n3181 VSS.n3180 8.65932
R3395 VSS.n3181 VSS 8.65932
R3396 VSS.n3179 VSS.n3178 8.65932
R3397 VSS VSS.n3179 8.65932
R3398 VSS VSS.n3144 8.65932
R3399 VSS.n3148 VSS.n3147 8.65932
R3400 VSS.n3147 VSS 8.65932
R3401 VSS.n3212 VSS.n3133 8.65932
R3402 VSS.n3133 VSS 8.65932
R3403 VSS.n3211 VSS.n3134 8.65932
R3404 VSS VSS.n3211 8.65932
R3405 VSS.n3204 VSS 8.65932
R3406 VSS.n3215 VSS.n3213 8.65932
R3407 VSS VSS.n3215 8.65932
R3408 VSS.n3218 VSS.n3217 8.65932
R3409 VSS.n3217 VSS 8.65932
R3410 VSS.n3225 VSS.n3216 8.65932
R3411 VSS.n3225 VSS 8.65932
R3412 VSS VSS.n3132 8.65932
R3413 VSS.n3224 VSS.n3223 8.65932
R3414 VSS.n3223 VSS 8.65932
R3415 VSS.n2922 VSS.n2796 8.65932
R3416 VSS VSS.n2922 8.65932
R3417 VSS.n3222 VSS.n3221 8.65932
R3418 VSS.n3221 VSS 8.65932
R3419 VSS.n5535 VSS 8.65932
R3420 VSS.n5534 VSS.n5533 8.65932
R3421 VSS.n5533 VSS 8.65932
R3422 VSS.n5532 VSS.n5531 8.65932
R3423 VSS.n5531 VSS 8.65932
R3424 VSS.n5530 VSS.n5487 8.65932
R3425 VSS.n5487 VSS 8.65932
R3426 VSS.n5529 VSS.n5528 8.65932
R3427 VSS.n5528 VSS 8.65932
R3428 VSS.n5496 VSS 8.65932
R3429 VSS.n5498 VSS.n5497 8.65932
R3430 VSS.n5497 VSS 8.65932
R3431 VSS.n5523 VSS.n5491 8.65932
R3432 VSS VSS.n5523 8.65932
R3433 VSS VSS.n5518 8.65932
R3434 VSS.n5515 VSS.n5514 8.65932
R3435 VSS.n5515 VSS 8.65932
R3436 VSS.n5513 VSS.n5508 8.65932
R3437 VSS.n5508 VSS 8.65932
R3438 VSS VSS.n5512 8.65932
R3439 VSS.n5509 VSS.n2782 8.65932
R3440 VSS.n5509 VSS 8.65932
R3441 VSS.n5556 VSS.n5554 8.65932
R3442 VSS VSS.n5556 8.65932
R3443 VSS VSS.n5553 8.65932
R3444 VSS.n3033 VSS.n3032 8.65932
R3445 VSS.n3032 VSS 8.65932
R3446 VSS VSS.n5557 8.65932
R3447 VSS.n5507 VSS 8.65932
R3448 VSS VSS.n5524 8.65932
R3449 VSS.n5527 VSS 8.65932
R3450 VSS.n5486 VSS 8.65932
R3451 VSS.n2923 VSS 8.65932
R3452 VSS VSS.n3309 8.65932
R3453 VSS VSS.n2933 8.65932
R3454 VSS VSS.n2936 8.65932
R3455 VSS VSS.n2939 8.65932
R3456 VSS VSS.n3290 8.65932
R3457 VSS.n3285 VSS.n3284 8.65932
R3458 VSS.n3285 VSS 8.65932
R3459 VSS VSS.n3283 8.65932
R3460 VSS.n3281 VSS.n2953 8.65932
R3461 VSS VSS.n3281 8.65932
R3462 VSS VSS.n6765 8.65932
R3463 VSS.n6761 VSS.n6760 8.65932
R3464 VSS.n6761 VSS 8.65932
R3465 VSS VSS.n6759 8.65932
R3466 VSS.n6756 VSS.n6755 8.65932
R3467 VSS.n6756 VSS 8.65932
R3468 VSS VSS.n6754 8.65932
R3469 VSS.n6752 VSS.n1019 8.65932
R3470 VSS VSS.n6752 8.65932
R3471 VSS.n1906 VSS.n1022 8.65932
R3472 VSS VSS.n1906 8.65932
R3473 VSS.n6748 VSS 8.65932
R3474 VSS.n6236 VSS.n1901 8.65932
R3475 VSS.n6236 VSS 8.65932
R3476 VSS.n6234 VSS.n1902 8.65932
R3477 VSS.n6234 VSS 8.65932
R3478 VSS VSS.n6240 8.65932
R3479 VSS.n2022 VSS.n2018 8.65932
R3480 VSS.n2022 VSS 8.65932
R3481 VSS.n2071 VSS 8.65932
R3482 VSS VSS.n2019 8.65932
R3483 VSS.n2070 VSS.n2069 8.65932
R3484 VSS.n2069 VSS 8.65932
R3485 VSS.n2031 VSS.n2027 8.65932
R3486 VSS VSS.n2031 8.65932
R3487 VSS.n2068 VSS.n2067 8.65932
R3488 VSS.n2067 VSS 8.65932
R3489 VSS VSS.n2028 8.65932
R3490 VSS.n2066 VSS.n2065 8.65932
R3491 VSS.n2065 VSS 8.65932
R3492 VSS VSS.n2043 8.65932
R3493 VSS.n2042 VSS.n2038 8.65932
R3494 VSS VSS.n2042 8.65932
R3495 VSS.n2064 VSS.n2063 8.65932
R3496 VSS.n2063 VSS 8.65932
R3497 VSS VSS.n2039 8.65932
R3498 VSS.n2062 VSS.n2061 8.65932
R3499 VSS.n2061 VSS 8.65932
R3500 VSS.n5956 VSS.n2005 8.65932
R3501 VSS VSS.n5956 8.65932
R3502 VSS.n5959 VSS 8.65932
R3503 VSS.n5958 VSS.n5957 8.65932
R3504 VSS VSS.n5958 8.65932
R3505 VSS.n5919 VSS.n5918 8.65932
R3506 VSS VSS.n5919 8.65932
R3507 VSS.n5952 VSS 8.65932
R3508 VSS.n5951 VSS.n5950 8.65932
R3509 VSS VSS.n5951 8.65932
R3510 VSS.n5947 VSS.n5923 8.65932
R3511 VSS.n5923 VSS 8.65932
R3512 VSS.n5944 VSS.n5943 8.65932
R3513 VSS.n5943 VSS 8.65932
R3514 VSS.n5990 VSS.n1961 8.65932
R3515 VSS.n5990 VSS 8.65932
R3516 VSS.n6023 VSS.n1953 8.65932
R3517 VSS.n6023 VSS 8.65932
R3518 VSS.n5987 VSS 8.65932
R3519 VSS.n5989 VSS.n5988 8.65932
R3520 VSS.n5988 VSS 8.65932
R3521 VSS.n5994 VSS.n1957 8.65932
R3522 VSS VSS.n5994 8.65932
R3523 VSS VSS.n5986 8.65932
R3524 VSS.n5985 VSS.n1962 8.65932
R3525 VSS VSS.n5985 8.65932
R3526 VSS.n5922 VSS 8.65932
R3527 VSS VSS.n5920 8.65932
R3528 VSS.n5921 VSS.n1965 8.65932
R3529 VSS VSS.n1965 8.65932
R3530 VSS.n5980 VSS.n1966 8.65932
R3531 VSS.n5980 VSS 8.65932
R3532 VSS.n5979 VSS.n1968 8.65932
R3533 VSS.n1968 VSS 8.65932
R3534 VSS.n5978 VSS.n5977 8.65932
R3535 VSS.n5977 VSS 8.65932
R3536 VSS.n5968 VSS 8.65932
R3537 VSS.n5967 VSS.n5965 8.65932
R3538 VSS VSS.n5967 8.65932
R3539 VSS.n5964 VSS.n2003 8.65932
R3540 VSS.n2003 VSS 8.65932
R3541 VSS VSS.n5963 8.65932
R3542 VSS.n2047 VSS.n2046 8.65932
R3543 VSS.n2046 VSS 8.65932
R3544 VSS.n2054 VSS.n2053 8.65932
R3545 VSS.n2054 VSS 8.65932
R3546 VSS VSS.n2052 8.65932
R3547 VSS.n2051 VSS.n2048 8.65932
R3548 VSS VSS.n2051 8.65932
R3549 VSS.n2032 VSS 8.65932
R3550 VSS.n6233 VSS 8.65932
R3551 VSS.n6232 VSS.n6231 8.65932
R3552 VSS.n6231 VSS 8.65932
R3553 VSS.n6230 VSS.n6229 8.65932
R3554 VSS.n6229 VSS 8.65932
R3555 VSS.n6228 VSS.n6227 8.65932
R3556 VSS.n6227 VSS 8.65932
R3557 VSS.n1990 VSS.n1988 8.65932
R3558 VSS VSS.n1990 8.65932
R3559 VSS VSS.n1987 8.65932
R3560 VSS.n1979 VSS.n1917 8.65932
R3561 VSS.n1979 VSS 8.65932
R3562 VSS.n6226 VSS.n6225 8.65932
R3563 VSS.n6225 VSS 8.65932
R3564 VSS VSS.n1918 8.65932
R3565 VSS.n6224 VSS.n6223 8.65932
R3566 VSS.n6223 VSS 8.65932
R3567 VSS VSS.n1970 8.65932
R3568 VSS.n1969 VSS.n1921 8.65932
R3569 VSS VSS.n1969 8.65932
R3570 VSS.n6222 VSS.n6221 8.65932
R3571 VSS.n6221 VSS 8.65932
R3572 VSS VSS.n1922 8.65932
R3573 VSS.n6220 VSS.n6219 8.65932
R3574 VSS.n6219 VSS 8.65932
R3575 VSS.n5971 VSS 8.65932
R3576 VSS.n5972 VSS.n1925 8.65932
R3577 VSS.n5972 VSS 8.65932
R3578 VSS.n6218 VSS.n6217 8.65932
R3579 VSS.n6217 VSS 8.65932
R3580 VSS VSS.n1926 8.65932
R3581 VSS.n6216 VSS.n6215 8.65932
R3582 VSS.n6215 VSS 8.65932
R3583 VSS.n6214 VSS.n6213 8.65932
R3584 VSS.n6213 VSS 8.65932
R3585 VSS.n5998 VSS 8.65932
R3586 VSS.n6212 VSS.n1929 8.65932
R3587 VSS VSS.n1929 8.65932
R3588 VSS.n6211 VSS.n6210 8.65932
R3589 VSS.n6210 VSS 8.65932
R3590 VSS.n5997 VSS 8.65932
R3591 VSS.n6007 VSS.n1956 8.65932
R3592 VSS VSS.n1956 8.65932
R3593 VSS VSS.n6006 8.65932
R3594 VSS.n5995 VSS 8.65932
R3595 VSS.n6009 VSS.n6008 8.65932
R3596 VSS.n6009 VSS 8.65932
R3597 VSS.n6019 VSS.n6018 8.65932
R3598 VSS.n6018 VSS 8.65932
R3599 VSS.n6012 VSS.n1955 8.65932
R3600 VSS VSS.n6012 8.65932
R3601 VSS.n6022 VSS 8.65932
R3602 VSS.n6021 VSS.n6020 8.65932
R3603 VSS.n6020 VSS 8.65932
R3604 VSS.n1946 VSS.n1932 8.65932
R3605 VSS.n1946 VSS 8.65932
R3606 VSS.n6017 VSS 8.65932
R3607 VSS.n6209 VSS 8.65932
R3608 VSS.n6208 VSS.n6207 8.65932
R3609 VSS.n6207 VSS 8.65932
R3610 VSS.n6206 VSS.n6205 8.65932
R3611 VSS.n6205 VSS 8.65932
R3612 VSS.n6204 VSS.n1939 8.65932
R3613 VSS VSS.n1939 8.65932
R3614 VSS.n6203 VSS.n6202 8.65932
R3615 VSS.n6202 VSS 8.65932
R3616 VSS VSS.n1938 8.65932
R3617 VSS.n1935 VSS.n1002 8.65932
R3618 VSS.n1935 VSS 8.65932
R3619 VSS.n6796 VSS.n6795 8.65932
R3620 VSS.n6796 VSS 8.65932
R3621 VSS VSS.n6794 8.65932
R3622 VSS.n6792 VSS.n6790 8.65932
R3623 VSS VSS.n6792 8.65932
R3624 VSS.n6789 VSS.n1003 8.65932
R3625 VSS VSS.n1003 8.65932
R3626 VSS VSS.n6788 8.65932
R3627 VSS.n1974 VSS.n1973 8.65932
R3628 VSS.n1973 VSS 8.65932
R3629 VSS.n1993 VSS.n1992 8.65932
R3630 VSS.n1993 VSS 8.65932
R3631 VSS VSS.n1991 8.65932
R3632 VSS.n6029 VSS.n6028 8.65932
R3633 VSS VSS.n6029 8.65932
R3634 VSS VSS.n6027 8.65932
R3635 VSS.n5940 VSS.n5930 8.65932
R3636 VSS.n5930 VSS 8.65932
R3637 VSS.n6030 VSS 8.65932
R3638 VSS VSS.n6039 8.65932
R3639 VSS VSS.n6045 8.65932
R3640 VSS VSS.n6051 8.65932
R3641 VSS.n6201 VSS 8.65932
R3642 VSS VSS.n961 8.65932
R3643 VSS VSS.n1005 8.65932
R3644 VSS VSS.n1008 8.65932
R3645 VSS VSS.n6772 8.65932
R3646 VSS.n1976 VSS.n1975 8.65932
R3647 VSS.n1975 VSS 8.65932
R3648 VSS.n1983 VSS 8.65932
R3649 VSS.n1982 VSS.n1017 8.65932
R3650 VSS VSS.n1982 8.65932
R3651 VSS.n1911 VSS 8.65932
R3652 VSS.n1912 VSS.n1909 8.65932
R3653 VSS.n1912 VSS 8.65932
R3654 VSS.n1907 VSS 8.65932
R3655 VSS.n2086 VSS.n2085 8.65932
R3656 VSS.n2085 VSS 8.65932
R3657 VSS.n2084 VSS 8.65932
R3658 VSS VSS.n5883 8.65932
R3659 VSS.n5880 VSS.n5879 8.65932
R3660 VSS.n5880 VSS 8.65932
R3661 VSS.n4025 VSS.n4011 8.53683
R3662 VSS.n4003 VSS.n3993 8.53683
R3663 VSS.n5256 VSS.n3905 8.53683
R3664 VSS.n663 VSS.n627 8.53683
R3665 VSS.n7178 VSS.n7103 8.53683
R3666 VSS.n887 VSS.n848 8.53683
R3667 VSS.n905 VSS.n876 8.53683
R3668 VSS.n6868 VSS.n914 8.53683
R3669 VSS.n840 VSS.n812 8.53683
R3670 VSS.n6992 VSS.n917 8.53683
R3671 VSS.n880 VSS.n879 8.53683
R3672 VSS.n4057 VSS.n3991 8.53683
R3673 VSS.n4454 VSS.n4357 8.53683
R3674 VSS.n4409 VSS.n4367 8.53683
R3675 VSS.n4610 VSS.n4609 8.53683
R3676 VSS.n5274 VSS.n3887 8.53683
R3677 VSS.n3897 VSS.n3896 8.53683
R3678 VSS.n4310 VSS.n3889 8.53683
R3679 VSS.n4349 VSS.n4281 8.53683
R3680 VSS.n4293 VSS.n4292 8.53683
R3681 VSS.n4338 VSS.n4336 8.53683
R3682 VSS.n4657 VSS.n4258 8.53683
R3683 VSS.n4649 VSS.n4648 8.53683
R3684 VSS.n4364 VSS.n4363 8.53683
R3685 VSS.n4960 VSS.n4959 8.53683
R3686 VSS.n4373 VSS.n4199 8.53683
R3687 VSS.n4822 VSS.n4197 8.53683
R3688 VSS.n4964 VSS.n4194 8.53683
R3689 VSS.n4928 VSS.n4746 8.53683
R3690 VSS.n4839 VSS.n4748 8.53683
R3691 VSS.n4921 VSS.n4846 8.53683
R3692 VSS.n4917 VSS.n4843 8.53683
R3693 VSS.n5160 VSS.n4117 8.53683
R3694 VSS.n4913 VSS.n4119 8.53683
R3695 VSS.n4131 VSS.n4122 8.53683
R3696 VSS.n5147 VSS.n4126 8.53683
R3697 VSS.n5134 VSS.n5127 8.53683
R3698 VSS.n5123 VSS.n4128 8.53683
R3699 VSS.n4835 VSS.n4805 8.53683
R3700 VSS.n4831 VSS.n4830 8.53683
R3701 VSS.n4815 VSS.n4813 8.53683
R3702 VSS.n4809 VSS.n4808 8.53683
R3703 VSS.n4676 VSS.n4675 8.53683
R3704 VSS.n4246 VSS.n4236 8.53683
R3705 VSS.n4681 VSS.n4680 8.53683
R3706 VSS.n4697 VSS.n4696 8.53683
R3707 VSS.n4743 VSS.n4227 8.53683
R3708 VSS.n4707 VSS.n4698 8.53683
R3709 VSS.n4730 VSS.n4702 8.53683
R3710 VSS.n4711 VSS.n4704 8.53683
R3711 VSS.n4717 VSS.n4715 8.53683
R3712 VSS.n5209 VSS.n4101 8.53683
R3713 VSS.n5196 VSS.n5189 8.53683
R3714 VSS.n5185 VSS.n4103 8.53683
R3715 VSS.n4251 VSS.n4241 8.53683
R3716 VSS.n4664 VSS.n4257 8.53683
R3717 VSS.n4264 VSS.n4244 8.53683
R3718 VSS.n4668 VSS.n4239 8.53683
R3719 VSS.n4044 VSS.n4009 8.53683
R3720 VSS.n4040 VSS.n4039 8.53683
R3721 VSS.n4016 VSS.n4014 8.53683
R3722 VSS.n4053 VSS.n4052 8.53683
R3723 VSS.n4021 VSS.n3996 8.53683
R3724 VSS.n4065 VSS.n4064 8.53683
R3725 VSS.n3999 VSS.n3988 8.53683
R3726 VSS.n4076 VSS.n4075 8.53683
R3727 VSS.n4092 VSS.n4091 8.53683
R3728 VSS.n4071 VSS.n3943 8.53683
R3729 VSS.n4096 VSS.n3938 8.53683
R3730 VSS.n3973 VSS.n3945 8.53683
R3731 VSS.n3960 VSS.n3953 8.53683
R3732 VSS.n3949 VSS.n3947 8.53683
R3733 VSS.n5263 VSS.n3899 8.53683
R3734 VSS.n4296 VSS.n3900 8.53683
R3735 VSS.n4031 VSS.n3908 8.53683
R3736 VSS.n5773 VSS.n2384 8.53683
R3737 VSS.n3956 VSS.n2386 8.53683
R3738 VSS.n5759 VSS.n2389 8.53683
R3739 VSS.n5741 VSS.n2403 8.53683
R3740 VSS.n5192 VSS.n2405 8.53683
R3741 VSS.n5727 VSS.n2408 8.53683
R3742 VSS.n5709 VSS.n2422 8.53683
R3743 VSS.n5130 VSS.n2424 8.53683
R3744 VSS.n5695 VSS.n2427 8.53683
R3745 VSS.n2534 VSS.n2528 8.53683
R3746 VSS.n2581 VSS.n2580 8.53683
R3747 VSS.n2559 VSS.n2553 8.53683
R3748 VSS.n2585 VSS.n2548 8.53683
R3749 VSS.n2542 VSS.n2530 8.53683
R3750 VSS.n2606 VSS.n2523 8.53683
R3751 VSS.n2613 VSS.n2611 8.53683
R3752 VSS.n5621 VSS.n5620 8.53683
R3753 VSS.n5612 VSS.n5611 8.53683
R3754 VSS.n7460 VSS.n310 8.53683
R3755 VSS.n646 VSS.n315 8.53683
R3756 VSS.n633 VSS.n631 8.53683
R3757 VSS.n677 VSS.n676 8.53683
R3758 VSS.n668 VSS.n667 8.53683
R3759 VSS.n6666 VSS.n788 8.53683
R3760 VSS.n823 VSS.n790 8.53683
R3761 VSS.n7049 VSS.n785 8.53683
R3762 VSS.n779 VSS.n778 8.53683
R3763 VSS.n7074 VSS.n757 8.53683
R3764 VSS.n7196 VSS.n752 8.53683
R3765 VSS.n7086 VSS.n7085 8.53683
R3766 VSS.n7077 VSS.n754 8.53683
R3767 VSS.n639 VSS.n629 8.53683
R3768 VSS.n650 VSS.n643 8.53683
R3769 VSS.n7416 VSS.n340 8.53683
R3770 VSS.n693 VSS.n342 8.53683
R3771 VSS.n7409 VSS.n700 8.53683
R3772 VSS.n7260 VSS.n697 8.53683
R3773 VSS.n7360 VSS.n7359 8.53683
R3774 VSS.n7355 VSS.n7258 8.53683
R3775 VSS.n7365 VSS.n7364 8.53683
R3776 VSS.n7377 VSS.n7375 8.53683
R3777 VSS.n7620 VSS.n85 8.53683
R3778 VSS.n7608 VSS.n7607 8.53683
R3779 VSS.n689 VSS.n417 8.53683
R3780 VSS.n685 VSS.n684 8.53683
R3781 VSS.n434 VSS.n425 8.53683
R3782 VSS.n421 VSS.n420 8.53683
R3783 VSS.n7123 VSS.n7122 8.53683
R3784 VSS.n7174 VSS.n7109 8.53683
R3785 VSS.n7127 VSS.n7124 8.53683
R3786 VSS.n7161 VSS.n7132 8.53683
R3787 VSS.n7137 VSS.n7134 8.53683
R3788 VSS.n7148 VSS.n7141 8.53683
R3789 VSS.n7246 VSS.n7245 8.53683
R3790 VSS.n7144 VSS.n718 8.53683
R3791 VSS.n7250 VSS.n713 8.53683
R3792 VSS.n6924 VSS.n6896 8.53683
R3793 VSS.n6911 VSS.n6904 8.53683
R3794 VSS.n6900 VSS.n6898 8.53683
R3795 VSS.n7185 VSS.n7088 8.53683
R3796 VSS.n7097 VSS.n7089 8.53683
R3797 VSS.n7114 VSS.n7106 8.53683
R3798 VSS.n7018 VSS.n851 8.53683
R3799 VSS.n7025 VSS.n807 8.53683
R3800 VSS.n844 VSS.n809 8.53683
R3801 VSS.n901 VSS.n900 8.53683
R3802 VSS.n892 VSS.n884 8.53683
R3803 VSS.n6999 VSS.n872 8.53683
R3804 VSS.n910 VSS.n874 8.53683
R3805 VSS.n6884 VSS.n6883 8.53683
R3806 VSS.n6872 VSS.n6865 8.53683
R3807 VSS.n6888 VSS.n6860 8.53683
R3808 VSS.n6968 VSS.n6856 8.53683
R3809 VSS.n6955 VSS.n6948 8.53683
R3810 VSS.n6944 VSS.n6858 8.53683
R3811 VSS.n836 VSS.n835 8.53683
R3812 VSS.n827 VSS.n820 8.53683
R3813 VSS.n816 VSS.n815 8.53683
R3814 VSS.n7717 VSS.n27 8.53683
R3815 VSS.n6951 VSS.n29 8.53683
R3816 VSS.n7703 VSS.n32 8.53683
R3817 VSS.n7685 VSS.n46 8.53683
R3818 VSS.n6907 VSS.n48 8.53683
R3819 VSS.n7671 VSS.n51 8.53683
R3820 VSS.n7653 VSS.n65 8.53683
R3821 VSS.n81 VSS.n67 8.53683
R3822 VSS.n7639 VSS.n70 8.53683
R3823 VSS.n4923 VSS.n4845 8.53633
R3824 VSS.n7411 VSS.n699 8.53633
R3825 VSS.n7648 VSS.n7643 8.53632
R3826 VSS.n7680 VSS.n7675 8.53632
R3827 VSS.n7712 VSS.n7707 8.53632
R3828 VSS.n6994 VSS.n916 8.53632
R3829 VSS.n882 VSS.n878 8.53632
R3830 VSS.n5704 VSS.n5699 8.53632
R3831 VSS.n5736 VSS.n5731 8.53632
R3832 VSS.n5768 VSS.n5763 8.53632
R3833 VSS.n4056 VSS.n3992 8.53632
R3834 VSS.n4821 VSS.n4196 8.53632
R3835 VSS.n4405 VSS.n4360 8.53632
R3836 VSS.n4605 VSS.n4371 8.53632
R3837 VSS.n4617 VSS.n4616 8.53632
R3838 VSS.n4300 VSS.n3892 8.53632
R3839 VSS.n4309 VSS.n3890 8.53632
R3840 VSS.n4288 VSS.n4286 8.53632
R3841 VSS.n4317 VSS.n4283 8.53632
R3842 VSS.n4268 VSS.n4260 8.53632
R3843 VSS.n4651 VSS.n4272 8.53632
R3844 VSS.n4628 VSS.n4627 8.53632
R3845 VSS.n5155 VSS.n4125 8.53632
R3846 VSS.n4130 VSS.n4123 8.53632
R3847 VSS.n5142 VSS.n5139 8.53632
R3848 VSS.n5125 VSS.n4129 8.53632
R3849 VSS.n4811 VSS.n4807 8.53632
R3850 VSS.n4688 VSS.n4687 8.53632
R3851 VSS.n4683 VSS.n4679 8.53632
R3852 VSS.n4739 VSS.n4701 8.53632
R3853 VSS.n4706 VSS.n4699 8.53632
R3854 VSS.n4725 VSS.n4721 8.53632
R3855 VSS.n4719 VSS.n4716 8.53632
R3856 VSS.n5204 VSS.n5201 8.53632
R3857 VSS.n5187 VSS.n4104 8.53632
R3858 VSS.n4667 VSS.n4240 8.53632
R3859 VSS.n4043 VSS.n4010 8.53632
R3860 VSS.n4083 VSS.n4082 8.53632
R3861 VSS.n4078 VSS.n4068 8.53632
R3862 VSS.n3978 VSS.n3941 8.53632
R3863 VSS.n4095 VSS.n3939 8.53632
R3864 VSS.n3968 VSS.n3965 8.53632
R3865 VSS.n3951 VSS.n3948 8.53632
R3866 VSS.n3909 VSS.n3907 8.53632
R3867 VSS.n5761 VSS.n2390 8.53632
R3868 VSS.n5729 VSS.n2409 8.53632
R3869 VSS.n5697 VSS.n2428 8.53632
R3870 VSS.n2627 VSS.n2513 8.53632
R3871 VSS.n2598 VSS.n2526 8.53632
R3872 VSS.n2568 VSS.n2551 8.53632
R3873 VSS.n2584 VSS.n2549 8.53632
R3874 VSS.n2605 VSS.n2524 8.53632
R3875 VSS.n5614 VSS.n2630 8.53632
R3876 VSS.n530 VSS.n529 8.53632
R3877 VSS.n670 VSS.n534 8.53632
R3878 VSS.n658 VSS.n654 8.53632
R3879 VSS.n7044 VSS.n793 8.53632
R3880 VSS.n7048 VSS.n786 8.53632
R3881 VSS.n7071 VSS.n7068 8.53632
R3882 VSS.n7063 VSS.n782 8.53632
R3883 VSS.n7092 VSS.n7081 8.53632
R3884 VSS.n7079 VSS.n755 8.53632
R3885 VSS.n7455 VSS.n318 8.53632
R3886 VSS.n765 VSS.n312 8.53632
R3887 VSS.n652 VSS.n644 8.53632
R3888 VSS.n7372 VSS.n7371 8.53632
R3889 VSS.n7367 VSS.n7363 8.53632
R3890 VSS.n7617 VSS.n7614 8.53632
R3891 VSS.n7610 VSS.n90 8.53632
R3892 VSS.n423 VSS.n419 8.53632
R3893 VSS.n7170 VSS.n7131 8.53632
R3894 VSS.n7129 VSS.n7125 8.53632
R3895 VSS.n7156 VSS.n7152 8.53632
R3896 VSS.n7150 VSS.n7142 8.53632
R3897 VSS.n6893 VSS.n716 8.53632
R3898 VSS.n7249 VSS.n714 8.53632
R3899 VSS.n6919 VSS.n6916 8.53632
R3900 VSS.n6902 VSS.n6899 8.53632
R3901 VSS.n7107 VSS.n7105 8.53632
R3902 VSS.n7020 VSS.n850 8.53632
R3903 VSS.n6875 VSS.n6863 8.53632
R3904 VSS.n6887 VSS.n6861 8.53632
R3905 VSS.n6963 VSS.n6960 8.53632
R3906 VSS.n6946 VSS.n6859 8.53632
R3907 VSS.n818 VSS.n814 8.53632
R3908 VSS.n7705 VSS.n33 8.53632
R3909 VSS.n7673 VSS.n52 8.53632
R3910 VSS.n7641 VSS.n71 8.53632
R3911 VSS.n2258 VSS.n2257 8.28285
R3912 VSS.n5842 VSS.t324 8.15922
R3913 VSS VSS.n2155 6.77697
R3914 VSS VSS.n2143 6.77697
R3915 VSS.n2132 VSS.n2131 6.77697
R3916 VSS.n2138 VSS.n2137 6.77697
R3917 VSS.n6271 VSS.n6270 6.77697
R3918 VSS.n6265 VSS.n6264 6.77697
R3919 VSS.n2249 VSS.n2248 5.57294
R3920 VSS.n2259 VSS 4.68305
R3921 VSS.n2131 VSS 4.67264
R3922 VSS.n6264 VSS 4.67264
R3923 VSS.n2265 VSS.n2264 4.6505
R3924 VSS.n2293 VSS.n2292 4.6505
R3925 VSS.n2295 VSS.n2294 4.6505
R3926 VSS.n2321 VSS.n2320 4.6505
R3927 VSS.n2323 VSS.n2322 4.6505
R3928 VSS.n2344 VSS.n2246 4.6505
R3929 VSS.n2348 VSS.n2347 4.6505
R3930 VSS.n2349 VSS.n2245 4.6505
R3931 VSS.n2267 VSS.n2266 4.6505
R3932 VSS.n2269 VSS.n2268 4.6505
R3933 VSS.n2274 VSS.n2273 4.6505
R3934 VSS.n2276 VSS.n2275 4.6505
R3935 VSS.n2278 VSS.n2277 4.6505
R3936 VSS.n2280 VSS.n2279 4.6505
R3937 VSS.n2285 VSS.n2284 4.6505
R3938 VSS.n2287 VSS.n2286 4.6505
R3939 VSS.n2289 VSS.n2288 4.6505
R3940 VSS.n2297 VSS.n2296 4.6505
R3941 VSS.n2302 VSS.n2301 4.6505
R3942 VSS.n2304 VSS.n2303 4.6505
R3943 VSS.n2306 VSS.n2305 4.6505
R3944 VSS.n2308 VSS.n2307 4.6505
R3945 VSS.n2313 VSS.n2312 4.6505
R3946 VSS.n2315 VSS.n2314 4.6505
R3947 VSS.n2317 VSS.n2316 4.6505
R3948 VSS.n2325 VSS.n2324 4.6505
R3949 VSS.n2330 VSS.n2329 4.6505
R3950 VSS.n2332 VSS.n2331 4.6505
R3951 VSS.n2334 VSS.n2333 4.6505
R3952 VSS.n2336 VSS.n2335 4.6505
R3953 VSS.n2341 VSS.n2340 4.6505
R3954 VSS.n2343 VSS.n2342 4.6505
R3955 VSS.n2346 VSS.n2345 4.6505
R3956 VSS.n2244 VSS.n2242 4.6505
R3957 VSS.n2243 VSS.n2240 4.6505
R3958 VSS.n2261 VSS.n2260 4.6505
R3959 VSS.n2355 VSS.n2354 4.6505
R3960 VSS.n2134 VSS.n2133 4.6505
R3961 VSS.n2145 VSS.n2144 4.6505
R3962 VSS.n2150 VSS.n2149 4.6505
R3963 VSS.n2157 VSS.n2156 4.6505
R3964 VSS.n2162 VSS.n2161 4.6505
R3965 VSS.n2135 VSS.n2123 4.6505
R3966 VSS.n2137 VSS.n2136 4.6505
R3967 VSS.n2140 VSS.n2139 4.6505
R3968 VSS.n2142 VSS.n2141 4.6505
R3969 VSS.n2143 VSS.n2121 4.6505
R3970 VSS.n2147 VSS.n2146 4.6505
R3971 VSS.n2152 VSS.n2151 4.6505
R3972 VSS.n2154 VSS.n2153 4.6505
R3973 VSS.n2155 VSS.n2118 4.6505
R3974 VSS.n2159 VSS.n2158 4.6505
R3975 VSS.n2164 VSS.n2163 4.6505
R3976 VSS.n2166 VSS.n2165 4.6505
R3977 VSS.n2168 VSS.n2167 4.6505
R3978 VSS.n6278 VSS.n6277 4.6505
R3979 VSS.n6283 VSS.n6282 4.6505
R3980 VSS.n6290 VSS.n6289 4.6505
R3981 VSS.n6295 VSS.n6294 4.6505
R3982 VSS.n6267 VSS.n6266 4.6505
R3983 VSS.n6268 VSS.n1892 4.6505
R3984 VSS.n6270 VSS.n6269 4.6505
R3985 VSS.n6273 VSS.n6272 4.6505
R3986 VSS.n6274 VSS.n1891 4.6505
R3987 VSS.n6276 VSS.n6275 4.6505
R3988 VSS.n6280 VSS.n6279 4.6505
R3989 VSS.n6285 VSS.n6284 4.6505
R3990 VSS.n6286 VSS.n1889 4.6505
R3991 VSS.n6288 VSS.n6287 4.6505
R3992 VSS.n6292 VSS.n6291 4.6505
R3993 VSS.n6297 VSS.n6296 4.6505
R3994 VSS.n6299 VSS.n6298 4.6505
R3995 VSS.n6301 VSS.n6300 4.6505
R3996 VSS.n1876 VSS.n1875 4.61383
R3997 VSS.n1875 VSS.n1874 4.61383
R3998 VSS.n2229 VSS.n2228 4.61383
R3999 VSS.n2228 VSS.n2227 4.61383
R4000 VSS.n2188 VSS.n2185 4.4948
R4001 VSS.n2213 VSS.n2212 4.4948
R4002 VSS.n6263 VSS.n1893 4.47386
R4003 VSS.n6802 VSS.n999 4.4066
R4004 VSS VSS.n6593 4.4066
R4005 VSS.n6612 VSS 4.4066
R4006 VSS VSS.n6713 4.4066
R4007 VSS.n3849 VSS 4.4066
R4008 VSS.n3833 VSS 4.4066
R4009 VSS.n3444 VSS.n2908 4.4066
R4010 VSS VSS.n5835 4.4066
R4011 VSS.n5406 VSS 4.4066
R4012 VSS VSS.n5484 4.4066
R4013 VSS.n5371 VSS 4.4066
R4014 VSS.n3347 VSS 4.4066
R4015 VSS.n3363 VSS 4.4066
R4016 VSS.n3460 VSS 4.4066
R4017 VSS.n3541 VSS 4.4066
R4018 VSS.n3557 VSS 4.4066
R4019 VSS.n3638 VSS 4.4066
R4020 VSS.n3654 VSS 4.4066
R4021 VSS.n3736 VSS 4.4066
R4022 VSS.n3752 VSS 4.4066
R4023 VSS.n6516 VSS 4.4066
R4024 VSS.n6534 VSS 4.4066
R4025 VSS VSS.n6075 4.4066
R4026 VSS VSS.n6194 4.4066
R4027 VSS.n6116 VSS 4.4066
R4028 VSS.n6815 VSS 4.4066
R4029 VSS.n1311 VSS 4.4066
R4030 VSS.n1246 VSS 4.4066
R4031 VSS.n6385 VSS 4.4066
R4032 VSS.n6440 VSS 4.4066
R4033 VSS.n6456 VSS 4.4066
R4034 VSS.n1051 VSS 4.39702
R4035 VSS.n7665 VSS.n58 4.11196
R4036 VSS.n7697 VSS.n39 4.11196
R4037 VSS.n7729 VSS.n20 4.11196
R4038 VSS.n7035 VSS.n7034 4.11196
R4039 VSS.n863 VSS.n858 4.11196
R4040 VSS.n7008 VSS.n866 4.11196
R4041 VSS.n929 VSS.n924 4.11196
R4042 VSS.n6982 VSS.n932 4.11196
R4043 VSS.n7216 VSS.n740 4.11196
R4044 VSS.n7225 VSS.n736 4.11196
R4045 VSS.n7232 VSS.n730 4.11196
R4046 VSS.n7236 VSS.n728 4.11196
R4047 VSS.n7429 VSS.n7425 4.11196
R4048 VSS.n7398 VSS.n7393 4.11196
R4049 VSS.n7402 VSS.n7391 4.11196
R4050 VSS.n5721 VSS.n2415 4.11196
R4051 VSS.n5753 VSS.n2396 4.11196
R4052 VSS.n5785 VSS.n2377 4.11196
R4053 VSS.n5290 VSS.n2856 4.11196
R4054 VSS.n5299 VSS.n2852 4.11196
R4055 VSS.n5308 VSS.n2848 4.11196
R4056 VSS.n5317 VSS.n2844 4.11196
R4057 VSS.n5324 VSS.n2838 4.11196
R4058 VSS.n5247 VSS.n3917 4.11196
R4059 VSS.n5242 VSS.n5239 4.11196
R4060 VSS.n5234 VSS.n5231 4.11196
R4061 VSS.n5226 VSS.n5223 4.11196
R4062 VSS.n4941 VSS.n4937 4.11196
R4063 VSS.n4222 VSS.n4219 4.11196
R4064 VSS.n5172 VSS.n4110 4.11196
R4065 VSS.n2592 VSS.n2539 4.11196
R4066 VSS.n5281 VSS.n2860 4.11196
R4067 VSS.n4324 VSS.n4306 4.11196
R4068 VSS.n4329 VSS.n4328 4.11196
R4069 VSS.n4635 VSS.n4278 4.11196
R4070 VSS.n4640 VSS.n4639 4.11196
R4071 VSS.n4947 VSS.n4211 4.11196
R4072 VSS.n5178 VSS.n5176 4.11196
R4073 VSS.n5220 VSS.n5218 4.11196
R4074 VSS.n5330 VSS.n5328 4.11196
R4075 VSS.n2620 VSS.n2519 4.11196
R4076 VSS.n6676 VSS.n6675 4.11196
R4077 VSS.n7056 VSS.n7055 4.11196
R4078 VSS.n7207 VSS.n744 4.11196
R4079 VSS.n773 VSS.n772 4.11196
R4080 VSS.n7444 VSS.n7443 4.11196
R4081 VSS.n7438 VSS.n7435 4.11196
R4082 VSS.n7388 VSS.n7386 4.11196
R4083 VSS.n6937 VSS.n6935 4.11196
R4084 VSS.n6979 VSS.n6977 4.11196
R4085 VSS.n4463 VSS.n4462 3.89651
R4086 VSS.n5281 VSS.n5280 3.89651
R4087 VSS.n4324 VSS.n4323 3.89651
R4088 VSS.n4328 VSS.n4326 3.89651
R4089 VSS.n4635 VSS.n4634 3.89651
R4090 VSS.n4639 VSS.n4637 3.89651
R4091 VSS.n4949 VSS.n4947 3.89651
R4092 VSS.n5176 VSS.n5175 3.89651
R4093 VSS.n5172 VSS.n5171 3.89651
R4094 VSS.n4219 VSS.n4218 3.89651
R4095 VSS.n4937 VSS.n4214 3.89651
R4096 VSS.n5218 VSS.n5217 3.89651
R4097 VSS.n5223 VSS.n3932 3.89651
R4098 VSS.n5231 VSS.n3927 3.89651
R4099 VSS.n5239 VSS.n3922 3.89651
R4100 VSS.n5249 VSS.n5247 3.89651
R4101 VSS.n5328 VSS.n5327 3.89651
R4102 VSS.n5324 VSS.n5323 3.89651
R4103 VSS.n5317 VSS.n5316 3.89651
R4104 VSS.n5308 VSS.n5307 3.89651
R4105 VSS.n5299 VSS.n5298 3.89651
R4106 VSS.n5290 VSS.n5289 3.89651
R4107 VSS.n5785 VSS.n5784 3.89651
R4108 VSS.n5753 VSS.n5752 3.89651
R4109 VSS.n5721 VSS.n5720 3.89651
R4110 VSS.n5686 VSS.n5685 3.89651
R4111 VSS.n2593 VSS.n2592 3.89651
R4112 VSS.n2620 VSS.n2619 3.89651
R4113 VSS.n6675 VSS.n6672 3.89651
R4114 VSS.n7057 VSS.n7056 3.89651
R4115 VSS.n7207 VSS.n7206 3.89651
R4116 VSS.n772 VSS.n771 3.89651
R4117 VSS.n7443 VSS.n325 3.89651
R4118 VSS.n7435 VSS.n331 3.89651
R4119 VSS.n7470 VSS.n7469 3.89651
R4120 VSS.n7386 VSS.n7385 3.89651
R4121 VSS.n7391 VSS.n707 3.89651
R4122 VSS.n7398 VSS.n7397 3.89651
R4123 VSS.n7425 VSS.n334 3.89651
R4124 VSS.n6935 VSS.n6934 3.89651
R4125 VSS.n728 VSS.n727 3.89651
R4126 VSS.n7232 VSS.n7231 3.89651
R4127 VSS.n7225 VSS.n7224 3.89651
R4128 VSS.n7216 VSS.n7215 3.89651
R4129 VSS.n6977 VSS.n6976 3.89651
R4130 VSS.n6984 VSS.n6982 3.89651
R4131 VSS.n929 VSS.n928 3.89651
R4132 VSS.n7010 VSS.n7008 3.89651
R4133 VSS.n863 VSS.n862 3.89651
R4134 VSS.n7034 VSS.n799 3.89651
R4135 VSS.n7729 VSS.n7728 3.89651
R4136 VSS.n7697 VSS.n7696 3.89651
R4137 VSS.n7665 VSS.n7664 3.89651
R4138 VSS.n7630 VSS.n7629 3.89651
R4139 VSS.n2572 VSS.n2571 3.71869
R4140 VSS.n3815 VSS.n2865 3.59425
R4141 VSS.n6660 VSS.n6659 3.59425
R4142 VSS VSS.n1029 3.33963
R4143 VSS.n2130 VSS.n2129 3.3223
R4144 VSS.n7544 VSS 3.31776
R4145 VSS.n146 VSS.t145 3.18343
R4146 VSS.n7650 VSS.t153 3.18343
R4147 VSS.n7682 VSS.t151 3.18343
R4148 VSS.n7714 VSS.t159 3.18343
R4149 VSS.n838 VSS.t189 3.18343
R4150 VSS.n7183 VSS.t181 3.18343
R4151 VSS.n687 VSS.t237 3.18343
R4152 VSS.n7332 VSS.t225 3.18343
R4153 VSS.n7585 VSS.t185 3.18343
R4154 VSS.n197 VSS.t165 3.18343
R4155 VSS.n2486 VSS.t147 3.18343
R4156 VSS.n5706 VSS.t135 3.18343
R4157 VSS.n5738 VSS.t149 3.18343
R4158 VSS.n5770 VSS.t139 3.18343
R4159 VSS.n5261 VSS.t269 3.18343
R4160 VSS.n4666 VSS.t263 3.18343
R4161 VSS.n4833 VSS.t215 3.18343
R4162 VSS.n4891 VSS.t133 3.18343
R4163 VSS.n4783 VSS.t235 3.18343
R4164 VSS.n4482 VSS.t211 3.18343
R4165 VSS.n4625 VSS.t193 3.18343
R4166 VSS.n4987 VSS.t259 3.18343
R4167 VSS.n4583 VSS.t279 3.18343
R4168 VSS.n4614 VSS.t267 3.18343
R4169 VSS.n5271 VSS.t195 3.18343
R4170 VSS.n4346 VSS.t217 3.18343
R4171 VSS.n4655 VSS.t283 3.18343
R4172 VSS.n4962 VSS.t245 3.18343
R4173 VSS.n5101 VSS.t275 3.18343
R4174 VSS.n5672 VSS.t171 3.18343
R4175 VSS.n4925 VSS.t281 3.18343
R4176 VSS.n5157 VSS.t261 3.18343
R4177 VSS.n5144 VSS.t157 3.18343
R4178 VSS.n4233 VSS.t241 3.18343
R4179 VSS.n4741 VSS.t137 3.18343
R4180 VSS.n4727 VSS.t277 3.18343
R4181 VSS.n5206 VSS.t173 3.18343
R4182 VSS.n4042 VSS.t247 3.18343
R4183 VSS.n4055 VSS.t221 3.18343
R4184 VSS.n3985 VSS.t125 3.18343
R4185 VSS.n4094 VSS.t265 3.18343
R4186 VSS.n3970 VSS.t161 3.18343
R4187 VSS.n3699 VSS.t257 3.18343
R4188 VSS.n3601 VSS.t231 3.18343
R4189 VSS.n3504 VSS.t199 3.18343
R4190 VSS.n3407 VSS.t271 3.18343
R4191 VSS.n5345 VSS.t249 3.18343
R4192 VSS.n5447 VSS.t143 3.18343
R4193 VSS.n3795 VSS.t183 3.18343
R4194 VSS.n5799 VSS.t129 3.18343
R4195 VSS.n2603 VSS.t93 3.18343
R4196 VSS.n2629 VSS.t108 3.18343
R4197 VSS.n2583 VSS.t106 3.18343
R4198 VSS.n395 VSS.t251 3.18343
R4199 VSS.n7488 VSS.t233 3.18343
R4200 VSS.n7457 VSS.t213 3.18343
R4201 VSS.n661 VSS.t187 3.18343
R4202 VSS.n505 VSS.t179 3.18343
R4203 VSS.n606 VSS.t203 3.18343
R4204 VSS.n431 VSS.t167 3.18343
R4205 VSS.n7046 VSS.t219 3.18343
R4206 VSS.n7073 VSS.t239 3.18343
R4207 VSS.n7193 VSS.t205 3.18343
R4208 VSS.n7413 VSS.t207 3.18343
R4209 VSS.n7255 VSS.t131 3.18343
R4210 VSS.n7619 VSS.t273 3.18343
R4211 VSS.n7172 VSS.t255 3.18343
R4212 VSS.n7158 VSS.t229 3.18343
R4213 VSS.n7248 VSS.t201 3.18343
R4214 VSS.n6921 VSS.t177 3.18343
R4215 VSS.n7022 VSS.t169 3.18343
R4216 VSS.n903 VSS.t243 3.18343
R4217 VSS.n6996 VSS.t209 3.18343
R4218 VSS.n6886 VSS.t141 3.18343
R4219 VSS.n6965 VSS.t127 3.18343
R4220 VSS.n6564 VSS.t175 3.18343
R4221 VSS.n6497 VSS.t155 3.18343
R4222 VSS.n6411 VSS.t223 3.18343
R4223 VSS.n1287 VSS.t191 3.18343
R4224 VSS.n6849 VSS.t253 3.18343
R4225 VSS.n6154 VSS.t227 3.18343
R4226 VSS.n1069 VSS.t197 3.18343
R4227 VSS.n7743 VSS.t163 3.18343
R4228 VSS.n179 VSS.t144 3.14684
R4229 VSS.n7651 VSS.t152 3.14684
R4230 VSS.n7683 VSS.t150 3.14684
R4231 VSS.n7715 VSS.t158 3.14684
R4232 VSS.n6167 VSS.t162 3.14684
R4233 VSS.n7289 VSS.t184 3.14684
R4234 VSS.n102 VSS.t164 3.14684
R4235 VSS.n2462 VSS.t146 3.14684
R4236 VSS.n5707 VSS.t134 3.14684
R4237 VSS.n5739 VSS.t148 3.14684
R4238 VSS.n5771 VSS.t138 3.14684
R4239 VSS.n5435 VSS.t128 3.14684
R4240 VSS.n5002 VSS.t234 3.14684
R4241 VSS.n4961 VSS.t244 3.14684
R4242 VSS.n4626 VSS.t192 3.14684
R4243 VSS.n4445 VSS.t210 3.14684
R4244 VSS.n4615 VSS.t266 3.14684
R4245 VSS.n4543 VSS.t258 3.14684
R4246 VSS.n4496 VSS.t278 3.14684
R4247 VSS.n4261 VSS.t282 3.14684
R4248 VSS.n5272 VSS.t194 3.14684
R4249 VSS.n3879 VSS.t182 3.14684
R4250 VSS.n4347 VSS.t216 3.14684
R4251 VSS.n4866 VSS.t274 3.14684
R4252 VSS.n4145 VSS.t170 3.14684
R4253 VSS.n4763 VSS.t132 3.14684
R4254 VSS.n4926 VSS.t280 3.14684
R4255 VSS.n5158 VSS.t260 3.14684
R4256 VSS.n5145 VSS.t156 3.14684
R4257 VSS.n4832 VSS.t214 3.14684
R4258 VSS.n4677 VSS.t240 3.14684
R4259 VSS.n4742 VSS.t136 3.14684
R4260 VSS.n4728 VSS.t276 3.14684
R4261 VSS.n5207 VSS.t172 3.14684
R4262 VSS.n4665 VSS.t262 3.14684
R4263 VSS.n4041 VSS.t246 3.14684
R4264 VSS.n4054 VSS.t220 3.14684
R4265 VSS.n4066 VSS.t124 3.14684
R4266 VSS.n4093 VSS.t264 3.14684
R4267 VSS.n3971 VSS.t160 3.14684
R4268 VSS.n5262 VSS.t268 3.14684
R4269 VSS.n3782 VSS.t256 3.14684
R4270 VSS.n3684 VSS.t230 3.14684
R4271 VSS.n3586 VSS.t198 3.14684
R4272 VSS.n3489 VSS.t270 3.14684
R4273 VSS.n3392 VSS.t248 3.14684
R4274 VSS.n2829 VSS.t142 3.14684
R4275 VSS.n2510 VSS.t107 3.14684
R4276 VSS.n2604 VSS.t92 3.14684
R4277 VSS.n2582 VSS.t105 3.14684
R4278 VSS.n465 VSS.t250 3.14684
R4279 VSS.n2732 VSS.t232 3.14684
R4280 VSS.n7458 VSS.t212 3.14684
R4281 VSS.n563 VSS.t178 3.14684
R4282 VSS.n7501 VSS.t202 3.14684
R4283 VSS.n533 VSS.t166 3.14684
R4284 VSS.n660 VSS.t186 3.14684
R4285 VSS.n7194 VSS.t204 3.14684
R4286 VSS.n7047 VSS.t218 3.14684
R4287 VSS.n6689 VSS.t196 3.14684
R4288 VSS.n758 VSS.t238 3.14684
R4289 VSS.n375 VSS.t224 3.14684
R4290 VSS.n7414 VSS.t206 3.14684
R4291 VSS.n7361 VSS.t130 3.14684
R4292 VSS.n86 VSS.t272 3.14684
R4293 VSS.n686 VSS.t236 3.14684
R4294 VSS.n7173 VSS.t254 3.14684
R4295 VSS.n7159 VSS.t228 3.14684
R4296 VSS.n7247 VSS.t200 3.14684
R4297 VSS.n6922 VSS.t176 3.14684
R4298 VSS.n7184 VSS.t180 3.14684
R4299 VSS.n7023 VSS.t168 3.14684
R4300 VSS.n902 VSS.t242 3.14684
R4301 VSS.n6997 VSS.t208 3.14684
R4302 VSS.n6885 VSS.t140 3.14684
R4303 VSS.n6966 VSS.t126 3.14684
R4304 VSS.n837 VSS.t188 3.14684
R4305 VSS.n1082 VSS.t174 3.14684
R4306 VSS.n1116 VSS.t154 3.14684
R4307 VSS.n6482 VSS.t222 3.14684
R4308 VSS.n1167 VSS.t190 3.14684
R4309 VSS.n1272 VSS.t252 3.14684
R4310 VSS.n950 VSS.t226 3.14684
R4311 VSS.n538 VSS 2.84776
R4312 VSS.n2329 VSS.n2328 2.63579
R4313 VSS.n2301 VSS.n2300 2.63579
R4314 VSS.n2273 VSS.n2272 2.63579
R4315 VSS.n6319 VSS.n1885 2.52171
R4316 VSS.n5854 VSS.t298 2.44766
R4317 VSS.n6734 VSS.t117 2.44494
R4318 VSS.n440 VSS 2.37788
R4319 VSS.n6594 VSS 2.37087
R4320 VSS VSS.n6605 2.37087
R4321 VSS.n6714 VSS 2.37087
R4322 VSS.n2950 VSS 2.37087
R4323 VSS.n2948 VSS 2.37087
R4324 VSS.n5836 VSS 2.37087
R4325 VSS VSS.n2804 2.37087
R4326 VSS.n5485 VSS 2.37087
R4327 VSS.n2925 VSS 2.37087
R4328 VSS VSS.n3313 2.37087
R4329 VSS.n3310 VSS 2.37087
R4330 VSS.n3303 VSS 2.37087
R4331 VSS.n3302 VSS 2.37087
R4332 VSS.n3299 VSS 2.37087
R4333 VSS.n3298 VSS 2.37087
R4334 VSS.n3295 VSS 2.37087
R4335 VSS.n3293 VSS 2.37087
R4336 VSS.n3291 VSS 2.37087
R4337 VSS VSS.n1011 2.37087
R4338 VSS.n6766 VSS 2.37087
R4339 VSS.n6076 VSS 2.37087
R4340 VSS.n6195 VSS 2.37087
R4341 VSS VSS.n959 2.37087
R4342 VSS VSS.n6804 2.37087
R4343 VSS VSS.n1000 2.37087
R4344 VSS.n6779 VSS 2.37087
R4345 VSS.n6777 VSS 2.37087
R4346 VSS.n6775 VSS 2.37087
R4347 VSS.n6773 VSS 2.37087
R4348 VSS.n4783 VSS.n4781 1.9205
R4349 VSS.n4987 VSS.n4190 1.9205
R4350 VSS.n4614 VSS.n4608 1.9205
R4351 VSS.n5271 VSS.n3895 1.9205
R4352 VSS.n4346 VSS.n4291 1.9205
R4353 VSS.n4655 VSS.n4654 1.9205
R4354 VSS.n4625 VSS.n4362 1.9205
R4355 VSS.n4482 VSS.n4481 1.9205
R4356 VSS.n5144 VSS.n5138 1.9205
R4357 VSS.n5206 VSS.n5200 1.9205
R4358 VSS.n3970 VSS.n3964 1.9205
R4359 VSS.n5447 VSS.n5444 1.9205
R4360 VSS.n3795 VSS.n3793 1.9205
R4361 VSS.n2603 VSS.n2602 1.9205
R4362 VSS.n395 VSS.n393 1.9205
R4363 VSS.n673 VSS.n431 1.9205
R4364 VSS.n7046 VSS.n792 1.9205
R4365 VSS.n7073 VSS.n7067 1.9205
R4366 VSS.n7193 VSS.n7084 1.9205
R4367 VSS.n7457 VSS.n317 1.9205
R4368 VSS.n661 VSS.n642 1.9205
R4369 VSS.n7488 VSS.n303 1.9205
R4370 VSS.n505 VSS.n504 1.9205
R4371 VSS.n7619 VSS.n7613 1.9205
R4372 VSS.n6921 VSS.n6915 1.9205
R4373 VSS.n6965 VSS.n6959 1.9205
R4374 VSS.n6154 VSS.n6147 1.9205
R4375 VSS.n1069 VSS.n1063 1.9205
R4376 VSS.n358 VSS 1.90776
R4377 VSS.n7584 VSS.n7582 1.87823
R4378 VSS.n196 VSS.n194 1.87823
R4379 VSS.n4582 VSS.n4581 1.87823
R4380 VSS.n4201 VSS.n4198 1.87823
R4381 VSS.n5100 VSS.n5098 1.87823
R4382 VSS.n5671 VSS.n5669 1.87823
R4383 VSS.n4890 VSS.n4889 1.87823
R4384 VSS.n4924 VSS.n4920 1.87823
R4385 VSS.n5152 VSS.n4124 1.87823
R4386 VSS.n4818 VSS.n4812 1.87823
R4387 VSS.n4685 VSS.n4684 1.87823
R4388 VSS.n4736 VSS.n4700 1.87823
R4389 VSS.n4722 VSS.n4720 1.87823
R4390 VSS.n4254 VSS.n4243 1.87823
R4391 VSS.n4028 VSS.n4013 1.87823
R4392 VSS.n4006 VSS.n3995 1.87823
R4393 VSS.n4080 VSS.n4079 1.87823
R4394 VSS.n3981 VSS.n3940 1.87823
R4395 VSS.n5260 VSS.n5259 1.87823
R4396 VSS.n3698 VSS.n3696 1.87823
R4397 VSS.n3600 VSS.n3598 1.87823
R4398 VSS.n3503 VSS.n3501 1.87823
R4399 VSS.n3406 VSS.n3404 1.87823
R4400 VSS.n5344 VSS.n5342 1.87823
R4401 VSS.n5796 VSS.n5795 1.87823
R4402 VSS.n5765 VSS.n5762 1.87823
R4403 VSS.n5733 VSS.n5730 1.87823
R4404 VSS.n5701 VSS.n5698 1.87823
R4405 VSS.n2479 VSS.n2478 1.87823
R4406 VSS.n2566 VSS.n2550 1.87823
R4407 VSS.n5616 VSS.n5615 1.87823
R4408 VSS.n605 VSS.n604 1.87823
R4409 VSS.n7331 VSS.n7330 1.87823
R4410 VSS.n7412 VSS.n701 1.87823
R4411 VSS.n7369 VSS.n7368 1.87823
R4412 VSS.n427 VSS.n424 1.87823
R4413 VSS.n7167 VSS.n7130 1.87823
R4414 VSS.n7153 VSS.n7151 1.87823
R4415 VSS.n6891 VSS.n715 1.87823
R4416 VSS.n7182 VSS.n7181 1.87823
R4417 VSS.n7021 VSS.n852 1.87823
R4418 VSS.n895 VSS.n883 1.87823
R4419 VSS.n6995 VSS.n918 1.87823
R4420 VSS.n6878 VSS.n6862 1.87823
R4421 VSS.n830 VSS.n819 1.87823
R4422 VSS.n6563 VSS.n6561 1.87823
R4423 VSS.n6496 VSS.n6494 1.87823
R4424 VSS.n6410 VSS.n6408 1.87823
R4425 VSS.n1286 VSS.n1284 1.87823
R4426 VSS.n6848 VSS.n6846 1.87823
R4427 VSS.n7740 VSS.n7739 1.87823
R4428 VSS.n7709 VSS.n7706 1.87823
R4429 VSS.n7677 VSS.n7674 1.87823
R4430 VSS.n7645 VSS.n7642 1.87823
R4431 VSS.n139 VSS.n138 1.87823
R4432 VSS.n6306 VSS 1.85727
R4433 VSS.n7289 VSS.n7282 1.84939
R4434 VSS.n102 VSS.n95 1.84939
R4435 VSS.n5002 VSS.n5001 1.84939
R4436 VSS.n4543 VSS.n4542 1.84939
R4437 VSS.n4496 VSS.n4489 1.84939
R4438 VSS.n4615 VSS.n4368 1.84939
R4439 VSS.n4347 VSS.n4285 1.84939
R4440 VSS.n4626 VSS.n4358 1.84939
R4441 VSS.n4961 VSS.n4202 1.84939
R4442 VSS.n4866 VSS.n4859 1.84939
R4443 VSS.n4145 VSS.n4138 1.84939
R4444 VSS.n4763 VSS.n4756 1.84939
R4445 VSS.n4926 VSS.n4842 1.84939
R4446 VSS.n5158 VSS.n4121 1.84939
R4447 VSS.n4832 VSS.n4819 1.84939
R4448 VSS.n4678 VSS.n4677 1.84939
R4449 VSS.n4742 VSS.n4230 1.84939
R4450 VSS.n4728 VSS.n4714 1.84939
R4451 VSS.n4665 VSS.n4255 1.84939
R4452 VSS.n4041 VSS.n4029 1.84939
R4453 VSS.n4054 VSS.n4007 1.84939
R4454 VSS.n4067 VSS.n4066 1.84939
R4455 VSS.n4093 VSS.n3982 1.84939
R4456 VSS.n5262 VSS.n3902 1.84939
R4457 VSS.n3782 VSS.n3775 1.84939
R4458 VSS.n3684 VSS.n3677 1.84939
R4459 VSS.n3586 VSS.n3579 1.84939
R4460 VSS.n3489 VSS.n3482 1.84939
R4461 VSS.n3392 VSS.n3385 1.84939
R4462 VSS.n5435 VSS.n5428 1.84939
R4463 VSS.n5771 VSS.n2388 1.84939
R4464 VSS.n5739 VSS.n2407 1.84939
R4465 VSS.n5707 VSS.n2426 1.84939
R4466 VSS.n2462 VSS.n2455 1.84939
R4467 VSS.n2582 VSS.n2562 1.84939
R4468 VSS.n5617 VSS.n2510 1.84939
R4469 VSS.n465 VSS.n464 1.84939
R4470 VSS.n7501 VSS.n7494 1.84939
R4471 VSS.n7066 VSS.n758 1.84939
R4472 VSS.n7458 VSS.n314 1.84939
R4473 VSS.n2732 VSS.n2731 1.84939
R4474 VSS.n375 VSS.n368 1.84939
R4475 VSS.n7414 VSS.n696 1.84939
R4476 VSS.n7362 VSS.n7361 1.84939
R4477 VSS.n686 VSS.n428 1.84939
R4478 VSS.n7173 VSS.n7112 1.84939
R4479 VSS.n7159 VSS.n7140 1.84939
R4480 VSS.n7247 VSS.n720 1.84939
R4481 VSS.n7184 VSS.n7100 1.84939
R4482 VSS.n7023 VSS.n847 1.84939
R4483 VSS.n902 VSS.n896 1.84939
R4484 VSS.n6997 VSS.n913 1.84939
R4485 VSS.n6885 VSS.n6879 1.84939
R4486 VSS.n837 VSS.n831 1.84939
R4487 VSS.n1082 VSS.n1080 1.84939
R4488 VSS.n1116 VSS.n1114 1.84939
R4489 VSS.n6482 VSS.n6475 1.84939
R4490 VSS.n1167 VSS.n1165 1.84939
R4491 VSS.n1272 VSS.n1265 1.84939
R4492 VSS.n6689 VSS.n6688 1.84939
R4493 VSS.n6167 VSS.n6165 1.84939
R4494 VSS.n7715 VSS.n31 1.84939
R4495 VSS.n7683 VSS.n50 1.84939
R4496 VSS.n7651 VSS.n69 1.84939
R4497 VSS.n179 VSS.n172 1.84939
R4498 VSS.n3894 VSS.n3891 1.8102
R4499 VSS.n4653 VSS.n4652 1.8102
R4500 VSS.n4442 VSS.n4441 1.8102
R4501 VSS.n5137 VSS.n5126 1.8102
R4502 VSS.n5199 VSS.n5188 1.8102
R4503 VSS.n3963 VSS.n3952 1.8102
R4504 VSS.n2823 VSS.n2822 1.8102
R4505 VSS.n3878 VSS.n3877 1.8102
R4506 VSS.n2601 VSS.n2525 1.8102
R4507 VSS.n672 VSS.n671 1.8102
R4508 VSS.n6664 VSS.n787 1.8102
R4509 VSS.n7083 VSS.n7080 1.8102
R4510 VSS.n655 VSS.n653 1.8102
R4511 VSS.n556 VSS.n555 1.8102
R4512 VSS.n7612 VSS.n7611 1.8102
R4513 VSS.n6914 VSS.n6903 1.8102
R4514 VSS.n6958 VSS.n6947 1.8102
R4515 VSS.n948 VSS.n947 1.8102
R4516 VSS.n1877 VSS.n1876 1.79444
R4517 VSS.n2219 VSS.n2209 1.74595
R4518 VSS.n2193 VSS.n2189 1.45505
R4519 VSS.n7272 VSS 1.43788
R4520 VSS.n1876 VSS.n1873 1.35808
R4521 VSS.n2170 VSS 1.34946
R4522 VSS VSS.n5588 1.11354
R4523 VSS.n5587 VSS 1.11354
R4524 VSS.n6594 VSS.n1015 0.976535
R4525 VSS.n6605 VSS.n6595 0.976535
R4526 VSS.n6715 VSS.n6714 0.976535
R4527 VSS.n2950 VSS.n2949 0.976535
R4528 VSS.n2948 VSS.n2942 0.976535
R4529 VSS.n5836 VSS.n2101 0.976535
R4530 VSS.n2804 VSS.n2803 0.976535
R4531 VSS.n5485 VSS.n2806 0.976535
R4532 VSS.n2926 VSS.n2925 0.976535
R4533 VSS.n3313 VSS.n3312 0.976535
R4534 VSS.n3311 VSS.n3310 0.976535
R4535 VSS.n3304 VSS.n3303 0.976535
R4536 VSS.n3302 VSS.n3301 0.976535
R4537 VSS.n3300 VSS.n3299 0.976535
R4538 VSS.n3298 VSS.n3297 0.976535
R4539 VSS.n3296 VSS.n3295 0.976535
R4540 VSS.n3294 VSS.n3293 0.976535
R4541 VSS.n3292 VSS.n3291 0.976535
R4542 VSS.n6768 VSS.n1011 0.976535
R4543 VSS.n6767 VSS.n6766 0.976535
R4544 VSS.n6076 VSS.n6056 0.976535
R4545 VSS.n6196 VSS.n6195 0.976535
R4546 VSS.n6200 VSS.n959 0.976535
R4547 VSS.n6804 VSS.n6803 0.976535
R4548 VSS.n6781 VSS.n1000 0.976535
R4549 VSS.n6780 VSS.n6779 0.976535
R4550 VSS.n6778 VSS.n6777 0.976535
R4551 VSS.n6776 VSS.n6775 0.976535
R4552 VSS.n6774 VSS.n6773 0.976535
R4553 VSS.n256 VSS 0.967877
R4554 VSS.n5642 VSS.n5641 0.95507
R4555 VSS.n2225 VSS.n2224 0.921712
R4556 VSS.n6319 VSS.n6312 0.921712
R4557 VSS.n2229 VSS.n2225 0.824742
R4558 VSS.n2356 VSS 0.741385
R4559 VSS.n5814 VSS.n2369 0.614203
R4560 VSS.n2172 VSS.n2171 0.572017
R4561 VSS.n6333 VSS.n6332 0.542292
R4562 VSS.n211 VSS 0.497878
R4563 VSS.n3816 VSS 0.426857
R4564 VSS.n3719 VSS 0.426857
R4565 VSS.n6307 VSS 0.424356
R4566 VSS.n2174 VSS.n2170 0.411958
R4567 VSS.n3330 VSS 0.39425
R4568 VSS.n5467 VSS 0.389562
R4569 VSS.n3621 VSS 0.383312
R4570 VSS.n6129 VSS 0.380708
R4571 VSS.n4 VSS 0.380708
R4572 VSS.n3427 VSS 0.380187
R4573 VSS.n6423 VSS 0.379146
R4574 VSS.n2340 VSS.n2339 0.376971
R4575 VSS.n2312 VSS.n2311 0.376971
R4576 VSS.n2284 VSS.n2283 0.376971
R4577 VSS.n2166 VSS.n2117 0.376971
R4578 VSS.n2154 VSS.n2120 0.376971
R4579 VSS.n6299 VSS.n1886 0.376971
R4580 VSS.n1889 VSS.n1888 0.376971
R4581 VSS.n4397 VSS 0.3755
R4582 VSS.n4379 VSS 0.3755
R4583 VSS.n4185 VSS 0.3755
R4584 VSS.n5037 VSS 0.3755
R4585 VSS.n3524 VSS 0.369771
R4586 VSS.n2441 VSS 0.368208
R4587 VSS.n1132 VSS 0.361958
R4588 VSS.n5648 VSS.n5644 0.352765
R4589 VSS.n352 VSS 0.352583
R4590 VSS.n966 VSS 0.346333
R4591 VSS.n4849 VSS 0.341646
R4592 VSS.n5627 VSS.n5626 0.340206
R4593 VSS.n5606 VSS.n5604 0.339716
R4594 VSS.n1098 VSS 0.339563
R4595 VSS.n1217 VSS 0.336958
R4596 VSS.n2753 VSS.n2752 0.334553
R4597 VSS.n6658 VSS 0.330188
R4598 VSS.n5054 VSS.n5053 0.329265
R4599 VSS.n551 VSS 0.3255
R4600 VSS.n5070 VSS.n5069 0.324095
R4601 VSS.n155 VSS 0.322896
R4602 VSS.n251 VSS 0.322896
R4603 VSS.n216 VSS 0.322896
R4604 VSS.n7278 VSS 0.322896
R4605 VSS.n5606 VSS 0.318729
R4606 VSS.n454 VSS 0.317167
R4607 VSS.n4422 VSS.n4419 0.315283
R4608 VSS.n4527 VSS.n4526 0.315283
R4609 VSS.n4559 VSS.n4555 0.315283
R4610 VSS.n5032 VSS.n5031 0.315283
R4611 VSS.n4155 VSS 0.313
R4612 VSS.n5081 VSS.n5077 0.310818
R4613 VSS.n7539 VSS 0.304667
R4614 VSS.n2189 VSS.n2184 0.291409
R4615 VSS.n2209 VSS.n2208 0.291409
R4616 VSS.n5626 VSS 0.284875
R4617 VSS.n2183 VSS 0.278917
R4618 VSS.n5817 VSS 0.278625
R4619 VSS.n6636 VSS 0.265604
R4620 VSS.n2571 VSS.n2570 0.252499
R4621 VSS.n5804 VSS.n5803 0.25175
R4622 VSS.n7749 VSS.n7747 0.25175
R4623 VSS.n2231 VSS.n2230 0.247667
R4624 VSS.n5422 VSS 0.247375
R4625 VSS.n6322 VSS.n6321 0.24733
R4626 VSS.n6470 VSS 0.246854
R4627 VSS.n2182 VSS.n2174 0.24399
R4628 VSS.n491 VSS 0.242435
R4629 VSS.n4770 VSS 0.235396
R4630 VSS.n5354 VSS 0.234354
R4631 VSS.n6551 VSS 0.234354
R4632 VSS.n3871 VSS.n3870 0.232887
R4633 VSS.n2577 VSS.n2576 0.232887
R4634 VSS.n6694 VSS.n6693 0.232887
R4635 VSS.n3572 VSS 0.228104
R4636 VSS.n2471 VSS 0.226021
R4637 VSS.n6834 VSS 0.226021
R4638 VSS.n6178 VSS 0.226021
R4639 VSS.n6698 VSS 0.221854
R4640 VSS.n2743 VSS 0.221854
R4641 VSS.n1297 VSS 0.210917
R4642 VSS.n3378 VSS 0.209875
R4643 VSS.n4431 VSS 0.207271
R4644 VSS.n4506 VSS 0.207271
R4645 VSS.n4551 VSS 0.207271
R4646 VSS.n5011 VSS 0.207271
R4647 VSS.n6396 VSS 0.204146
R4648 VSS.n589 VSS 0.203203
R4649 VSS.n3475 VSS 0.201542
R4650 VSS.n3866 VSS 0.186437
R4651 VSS.n3768 VSS 0.186437
R4652 VSS.n3670 VSS 0.185396
R4653 VSS.n4875 VSS 0.183833
R4654 VSS.n7529 VSS 0.181229
R4655 VSS.n5086 VSS 0.180188
R4656 VSS.n261 VSS 0.178625
R4657 VSS.n225 VSS 0.178625
R4658 VSS.n7568 VSS 0.178625
R4659 VSS.n7316 VSS 0.178625
R4660 VSS.n3450 VSS.n3449 0.174048
R4661 VSS.n5569 VSS.n5568 0.17393
R4662 VSS.n3839 VSS.n3838 0.17393
R4663 VSS.n3742 VSS.n3741 0.17393
R4664 VSS.n5396 VSS.n5395 0.17393
R4665 VSS.n6446 VSS.n6445 0.17393
R4666 VSS.n3644 VSS.n3643 0.173813
R4667 VSS.n3547 VSS.n3546 0.173813
R4668 VSS.n3353 VSS.n3352 0.173813
R4669 VSS.n5377 VSS.n5376 0.173813
R4670 VSS.n6529 VSS.n6528 0.173813
R4671 VSS.n7316 VSS 0.172914
R4672 VSS.n7568 VSS 0.172914
R4673 VSS.n261 VSS 0.172914
R4674 VSS.n225 VSS 0.172914
R4675 VSS.n589 VSS 0.171854
R4676 VSS.n2491 VSS.n2475 0.169915
R4677 VSS.n4450 VSS.n4449 0.168417
R4678 VSS.n5277 VSS.n5276 0.168417
R4679 VSS.n4320 VSS.n4319 0.168417
R4680 VSS.n4631 VSS.n4630 0.168417
R4681 VSS.n2597 VSS.n2596 0.168417
R4682 VSS.n2616 VSS.n2615 0.168417
R4683 VSS.n6669 VSS.n6668 0.168417
R4684 VSS.n7061 VSS.n7060 0.168417
R4685 VSS.n768 VSS.n767 0.168417
R4686 VSS.n2727 VSS.n2726 0.168417
R4687 VSS.n4435 VSS.n4434 0.167667
R4688 VSS.n5623 VSS.n2508 0.167667
R4689 VSS.n5609 VSS.n5608 0.167667
R4690 VSS.n2740 VSS.n2738 0.167667
R4691 VSS.n152 VSS.n151 0.167667
R4692 VSS.n142 VSS.n72 0.167667
R4693 VSS.n7644 VSS.n53 0.167667
R4694 VSS.n7676 VSS.n34 0.167667
R4695 VSS.n7708 VSS.n15 0.167667
R4696 VSS.n2482 VSS.n2429 0.167667
R4697 VSS.n5700 VSS.n2410 0.167667
R4698 VSS.n5732 VSS.n2391 0.167667
R4699 VSS.n5764 VSS.n2372 0.167667
R4700 VSS.n2625 VSS.n2624 0.167667
R4701 VSS.n2547 VSS.n2544 0.167667
R4702 VSS.n5086 VSS 0.167167
R4703 VSS.n2574 VSS.n2573 0.167167
R4704 VSS.n491 VSS 0.165604
R4705 VSS.n2576 VSS.n2564 0.16503
R4706 VSS.n7529 VSS 0.163543
R4707 VSS.n4875 VSS 0.155139
R4708 VSS.n3670 VSS 0.1505
R4709 VSS.n3866 VSS 0.147559
R4710 VSS.n3768 VSS 0.147559
R4711 VSS.n4457 VSS 0.146833
R4712 VSS.n3884 VSS 0.146833
R4713 VSS.n4313 VSS 0.146833
R4714 VSS.n4352 VSS 0.146833
R4715 VSS VSS.n4435 0.146833
R4716 VSS VSS.n5789 0.146833
R4717 VSS VSS.n5757 0.146833
R4718 VSS VSS.n5725 0.146833
R4719 VSS VSS.n5693 0.146833
R4720 VSS.n2491 VSS 0.146833
R4721 VSS.n5623 VSS 0.146833
R4722 VSS VSS.n2515 0.146833
R4723 VSS VSS.n2557 0.146833
R4724 VSS.n2588 VSS 0.146833
R4725 VSS.n2609 VSS 0.146833
R4726 VSS VSS.n5609 0.146833
R4727 VSS.n2738 VSS 0.146833
R4728 VSS.n7463 VSS 0.146833
R4729 VSS VSS.n6679 0.146833
R4730 VSS.n7052 VSS 0.146833
R4731 VSS VSS.n776 0.146833
R4732 VSS VSS.n7733 0.146833
R4733 VSS VSS.n7701 0.146833
R4734 VSS VSS.n7669 0.146833
R4735 VSS VSS.n7637 0.146833
R4736 VSS.n151 VSS 0.146833
R4737 VSS.n3717 VSS.n2879 0.142792
R4738 VSS.n3814 VSS.n2870 0.142557
R4739 VSS.n2175 VSS.n2101 0.140147
R4740 VSS.n2803 VSS.n2802 0.140147
R4741 VSS.n2806 VSS.n2805 0.140147
R4742 VSS.n2927 VSS.n2926 0.140147
R4743 VSS.n3312 VSS.n2929 0.140147
R4744 VSS.n3311 VSS.n2930 0.140147
R4745 VSS.n3304 VSS.n2932 0.140147
R4746 VSS.n3301 VSS.n2934 0.140147
R4747 VSS.n3300 VSS.n2935 0.140147
R4748 VSS.n3297 VSS.n2937 0.140147
R4749 VSS.n3296 VSS.n2938 0.140147
R4750 VSS.n3294 VSS.n2940 0.140147
R4751 VSS.n3292 VSS.n2941 0.140147
R4752 VSS.n3287 VSS.n2942 0.140147
R4753 VSS.n2949 VSS.n2947 0.140147
R4754 VSS.n1015 VSS.n1014 0.140147
R4755 VSS.n6601 VSS.n6595 0.140147
R4756 VSS.n6715 VSS.n1028 0.140147
R4757 VSS.n6769 VSS.n6768 0.140147
R4758 VSS.n6767 VSS.n1013 0.140147
R4759 VSS.n6056 VSS.n6055 0.140147
R4760 VSS.n6197 VSS.n6196 0.140147
R4761 VSS.n6200 VSS.n6199 0.140147
R4762 VSS.n6803 VSS.n960 0.140147
R4763 VSS.n6782 VSS.n6781 0.140147
R4764 VSS.n6780 VSS.n1006 0.140147
R4765 VSS.n6778 VSS.n1007 0.140147
R4766 VSS.n6776 VSS.n1009 0.140147
R4767 VSS.n6774 VSS.n1010 0.140147
R4768 VSS.n4458 VSS.n4457 0.14005
R4769 VSS.n4314 VSS.n4313 0.14005
R4770 VSS.n3885 VSS.n3884 0.14005
R4771 VSS.n4353 VSS.n4352 0.14005
R4772 VSS.n2557 VSS.n2556 0.14005
R4773 VSS.n2609 VSS.n2522 0.14005
R4774 VSS.n7464 VSS.n7463 0.14005
R4775 VSS.n7053 VSS.n7052 0.14005
R4776 VSS.n6679 VSS.n6678 0.14005
R4777 VSS.n776 VSS.n775 0.14005
R4778 VSS.n5588 VSS.n2780 0.139843
R4779 VSS.n6600 VSS.n1029 0.139843
R4780 VSS.n5587 VSS.n5586 0.139843
R4781 VSS.n5278 VSS.n5277 0.13959
R4782 VSS.n4321 VSS.n4320 0.13959
R4783 VSS.n4632 VSS.n4631 0.13959
R4784 VSS.n2617 VSS.n2616 0.13959
R4785 VSS.n2596 VSS.n2595 0.13959
R4786 VSS.n6670 VSS.n6669 0.13959
R4787 VSS.n7060 VSS.n7059 0.13959
R4788 VSS.n769 VSS.n768 0.13959
R4789 VSS.n2708 VSS 0.137248
R4790 VSS.n4431 VSS.n4430 0.136775
R4791 VSS.n4506 VSS.n4505 0.136775
R4792 VSS.n4552 VSS.n4551 0.136775
R4793 VSS.n5011 VSS.n5010 0.136775
R4794 VSS.n4770 VSS.n4754 0.136775
R4795 VSS.n4156 VSS.n4155 0.136775
R4796 VSS.n2472 VSS.n2471 0.136775
R4797 VSS.n5086 VSS.n5084 0.136775
R4798 VSS.n4875 VSS.n4873 0.136775
R4799 VSS.n2744 VSS.n2743 0.136775
R4800 VSS.n551 VSS.n550 0.136775
R4801 VSS.n454 VSS.n452 0.136775
R4802 VSS.n589 VSS.n587 0.136775
R4803 VSS.n7529 VSS.n7527 0.136775
R4804 VSS.n7540 VSS.n7539 0.136775
R4805 VSS.n491 VSS.n489 0.136775
R4806 VSS.n262 VSS.n261 0.136775
R4807 VSS.n7278 VSS.n7276 0.136775
R4808 VSS.n252 VSS.n251 0.136775
R4809 VSS.n216 VSS.n215 0.136775
R4810 VSS.n226 VSS.n225 0.136775
R4811 VSS.n7568 VSS.n7566 0.136775
R4812 VSS.n7316 VSS.n7314 0.136775
R4813 VSS.n156 VSS.n155 0.136775
R4814 VSS.n2182 VSS 0.129576
R4815 VSS.n3425 VSS.n2911 0.128457
R4816 VSS.n4520 VSS.n4519 0.127988
R4817 VSS.n4563 VSS.n4562 0.127988
R4818 VSS.n5025 VSS.n5024 0.127988
R4819 VSS.n3522 VSS.n2899 0.127988
R4820 VSS.n3328 VSS.n3316 0.126108
R4821 VSS.n5063 VSS.n5062 0.125637
R4822 VSS.n153 VSS 0.1255
R4823 VSS.n73 VSS 0.1255
R4824 VSS.n55 VSS 0.1255
R4825 VSS.n36 VSS 0.1255
R4826 VSS.n17 VSS 0.1255
R4827 VSS.n93 VSS 0.1255
R4828 VSS.n7279 VSS 0.1255
R4829 VSS.n2430 VSS 0.1255
R4830 VSS.n2412 VSS 0.1255
R4831 VSS.n2393 VSS 0.1255
R4832 VSS.n2374 VSS 0.1255
R4833 VSS.n4853 VSS 0.1255
R4834 VSS.n4451 VSS 0.1255
R4835 VSS.n2862 VSS 0.1255
R4836 VSS.n4308 VSS 0.1255
R4837 VSS.n4280 VSS 0.1255
R4838 VSS.n4399 VSS 0.1255
R4839 VSS.n4568 VSS 0.1255
R4840 VSS.n4187 VSS 0.1255
R4841 VSS.n5039 VSS 0.1255
R4842 VSS.n4135 VSS 0.1255
R4843 VSS.n5657 VSS 0.1255
R4844 VSS.n2872 VSS 0.1255
R4845 VSS.n2881 VSS 0.1255
R4846 VSS.n2890 VSS 0.1255
R4847 VSS.n2901 VSS 0.1255
R4848 VSS.n2913 VSS 0.1255
R4849 VSS.n3318 VSS 0.1255
R4850 VSS.n5386 VSS 0.1255
R4851 VSS.n5805 VSS 0.1255
R4852 VSS.n5607 VSS 0.1255
R4853 VSS.n2514 VSS 0.1255
R4854 VSS.n2537 VSS 0.1255
R4855 VSS.n2565 VSS 0.1255
R4856 VSS.n2572 VSS.n2564 0.1255
R4857 VSS.n2546 VSS 0.1255
R4858 VSS.n2521 VSS 0.1255
R4859 VSS.n7537 VSS 0.1255
R4860 VSS.n6663 VSS 0.1255
R4861 VSS.n783 VSS 0.1255
R4862 VSS.n763 VSS 0.1255
R4863 VSS.n309 VSS 0.1255
R4864 VSS.n552 VSS 0.1255
R4865 VSS.n455 VSS 0.1255
R4866 VSS.n363 VSS 0.1255
R4867 VSS.n217 VSS 0.1255
R4868 VSS.n6641 VSS 0.1255
R4869 VSS.n1105 VSS 0.1255
R4870 VSS.n1139 VSS 0.1255
R4871 VSS.n1157 VSS 0.1255
R4872 VSS.n1257 VSS 0.1255
R4873 VSS.n976 VSS 0.1255
R4874 VSS.n6140 VSS 0.1255
R4875 VSS.n7748 VSS 0.1255
R4876 VSS.n3619 VSS.n2888 0.12505
R4877 VSS.n2699 VSS 0.1227
R4878 VSS.n5652 VSS.n5651 0.122113
R4879 VSS.n5465 VSS.n5384 0.122113
R4880 VSS.n5047 VSS.n5046 0.121642
R4881 VSS.n2265 VSS.n2261 0.120292
R4882 VSS.n2267 VSS.n2265 0.120292
R4883 VSS.n2269 VSS.n2267 0.120292
R4884 VSS.n2274 VSS.n2269 0.120292
R4885 VSS.n2276 VSS.n2274 0.120292
R4886 VSS.n2278 VSS.n2276 0.120292
R4887 VSS.n2280 VSS.n2278 0.120292
R4888 VSS.n2285 VSS.n2280 0.120292
R4889 VSS.n2286 VSS.n2285 0.120292
R4890 VSS.n2293 VSS.n2289 0.120292
R4891 VSS.n2295 VSS.n2293 0.120292
R4892 VSS.n2297 VSS.n2295 0.120292
R4893 VSS.n2302 VSS.n2297 0.120292
R4894 VSS.n2304 VSS.n2302 0.120292
R4895 VSS.n2306 VSS.n2304 0.120292
R4896 VSS.n2308 VSS.n2306 0.120292
R4897 VSS.n2313 VSS.n2308 0.120292
R4898 VSS.n2314 VSS.n2313 0.120292
R4899 VSS.n2321 VSS.n2317 0.120292
R4900 VSS.n2323 VSS.n2321 0.120292
R4901 VSS.n2325 VSS.n2323 0.120292
R4902 VSS.n2330 VSS.n2325 0.120292
R4903 VSS.n2332 VSS.n2330 0.120292
R4904 VSS.n2334 VSS.n2332 0.120292
R4905 VSS.n2336 VSS.n2334 0.120292
R4906 VSS.n2341 VSS.n2336 0.120292
R4907 VSS.n2342 VSS.n2341 0.120292
R4908 VSS.n2347 VSS.n2346 0.120292
R4909 VSS.n2244 VSS.n2243 0.120292
R4910 VSS.n2135 VSS.n2134 0.120292
R4911 VSS.n2141 VSS.n2140 0.120292
R4912 VSS.n2145 VSS.n2121 0.120292
R4913 VSS.n2147 VSS.n2145 0.120292
R4914 VSS.n2150 VSS.n2147 0.120292
R4915 VSS.n2152 VSS.n2150 0.120292
R4916 VSS.n2153 VSS.n2152 0.120292
R4917 VSS.n2157 VSS.n2118 0.120292
R4918 VSS.n2159 VSS.n2157 0.120292
R4919 VSS.n2162 VSS.n2159 0.120292
R4920 VSS.n2164 VSS.n2162 0.120292
R4921 VSS.n2165 VSS.n2164 0.120292
R4922 VSS.n6268 VSS.n6267 0.120292
R4923 VSS.n6274 VSS.n6273 0.120292
R4924 VSS.n6280 VSS.n6278 0.120292
R4925 VSS.n6283 VSS.n6280 0.120292
R4926 VSS.n6285 VSS.n6283 0.120292
R4927 VSS.n6286 VSS.n6285 0.120292
R4928 VSS.n6292 VSS.n6290 0.120292
R4929 VSS.n6295 VSS.n6292 0.120292
R4930 VSS.n6297 VSS.n6295 0.120292
R4931 VSS.n6298 VSS.n6297 0.120292
R4932 VSS.n5074 VSS.n5073 0.119998
R4933 VSS.n2365 VSS.n2364 0.119058
R4934 VSS.n2360 VSS.n1864 0.119058
R4935 VSS.n5817 VSS.n5816 0.118209
R4936 VSS.n2709 VSS.n2708 0.112194
R4937 VSS.n2699 VSS.n2502 0.112194
R4938 VSS.n4407 VSS.n4360 0.109769
R4939 VSS.n4302 VSS.n3892 0.109769
R4940 VSS.n4286 VSS.n4273 0.109769
R4941 VSS.n4267 VSS.n4260 0.109769
R4942 VSS.n7094 VSS.n7081 0.109769
R4943 VSS.n7649 VSS.n7644 0.109764
R4944 VSS.n7681 VSS.n7676 0.109764
R4945 VSS.n7713 VSS.n7708 0.109764
R4946 VSS.n5705 VSS.n5700 0.109764
R4947 VSS.n5737 VSS.n5732 0.109764
R4948 VSS.n5769 VSS.n5764 0.109764
R4949 VSS.n2628 VSS.n2625 0.109764
R4950 VSS.n2570 VSS.n2552 0.109764
R4951 VSS.n4630 VSS.n4355 0.109764
R4952 VSS.n4619 VSS.n4365 0.109764
R4953 VSS.n4319 VSS.n4284 0.109764
R4954 VSS.n5156 VSS.n5151 0.109764
R4955 VSS.n5143 VSS.n2421 0.109764
R4956 VSS.n4690 VSS.n4689 0.109764
R4957 VSS.n4740 VSS.n4735 0.109764
R4958 VSS.n4726 VSS.n4100 0.109764
R4959 VSS.n5205 VSS.n2402 0.109764
R4960 VSS.n4085 VSS.n4084 0.109764
R4961 VSS.n3977 VSS.n3942 0.109764
R4962 VSS.n3969 VSS.n2383 0.109764
R4963 VSS.n2597 VSS.n2527 0.109764
R4964 VSS.n767 VSS.n313 0.109764
R4965 VSS.n659 VSS.n319 0.109764
R4966 VSS.n7045 VSS.n7041 0.109764
R4967 VSS.n7062 VSS.n7061 0.109764
R4968 VSS.n7072 VSS.n751 0.109764
R4969 VSS.n7456 VSS.n7452 0.109764
R4970 VSS.n7374 VSS.n7373 0.109764
R4971 VSS.n7618 VSS.n64 0.109764
R4972 VSS.n7171 VSS.n7166 0.109764
R4973 VSS.n7157 VSS.n722 0.109764
R4974 VSS.n6895 VSS.n717 0.109764
R4975 VSS.n6920 VSS.n45 0.109764
R4976 VSS.n6864 VSS.n6855 0.109764
R4977 VSS.n6964 VSS.n26 0.109764
R4978 VSS.n4604 VSS.n4370 0.109764
R4979 VSS.n528 VSS.n527 0.109764
R4980 VSS.n5255 VSS.n3905 0.108274
R4981 VSS.n665 VSS.n627 0.108274
R4982 VSS.n7177 VSS.n7103 0.108274
R4983 VSS.n842 VSS.n812 0.108274
R4984 VSS.n6991 VSS.n917 0.108269
R4985 VSS.n879 VSS.n871 0.108269
R4986 VSS.n4059 VSS.n3991 0.108269
R4987 VSS.n4824 VSS.n4197 0.108269
R4988 VSS.n4648 VSS.n4647 0.108269
R4989 VSS.n4312 VSS.n3889 0.108269
R4990 VSS.n5276 VSS.n3887 0.108269
R4991 VSS.n4340 VSS.n4336 0.108269
R4992 VSS.n4846 VSS.n4116 0.108269
R4993 VSS.n5149 VSS.n4126 0.108269
R4994 VSS.n5133 VSS.n5127 0.108269
R4995 VSS.n5211 VSS.n4101 0.108269
R4996 VSS.n5195 VSS.n5189 0.108269
R4997 VSS.n4664 VSS.n4663 0.108269
R4998 VSS.n4046 VSS.n4009 0.108269
R4999 VSS.n3975 VSS.n3945 0.108269
R5000 VSS.n3959 VSS.n3953 0.108269
R5001 VSS.n5264 VSS.n5263 0.108269
R5002 VSS.n649 VSS.n643 0.108269
R5003 VSS.n648 VSS.n315 0.108269
R5004 VSS.n635 VSS.n631 0.108269
R5005 VSS.n7076 VSS.n754 0.108269
R5006 VSS.n7051 VSS.n785 0.108269
R5007 VSS.n6668 VSS.n788 0.108269
R5008 VSS.n825 VSS.n790 0.108269
R5009 VSS.n7075 VSS.n7074 0.108269
R5010 VSS.n7198 VSS.n752 0.108269
R5011 VSS.n7408 VSS.n700 0.108269
R5012 VSS.n7379 VSS.n7375 0.108269
R5013 VSS.n7621 VSS.n7620 0.108269
R5014 VSS.n6926 VSS.n6896 0.108269
R5015 VSS.n6910 VSS.n6904 0.108269
R5016 VSS.n7186 VSS.n7185 0.108269
R5017 VSS.n7017 VSS.n851 0.108269
R5018 VSS.n6970 VSS.n6856 0.108269
R5019 VSS.n6954 VSS.n6948 0.108269
R5020 VSS.n836 VSS.n794 0.108269
R5021 VSS.n7638 VSS.n70 0.108269
R5022 VSS.n7670 VSS.n51 0.108269
R5023 VSS.n7702 VSS.n32 0.108269
R5024 VSS.n6890 VSS.n6860 0.108269
R5025 VSS.n6870 VSS.n914 0.108269
R5026 VSS.n907 VSS.n876 0.108269
R5027 VSS.n7252 VSS.n713 0.108269
R5028 VSS.n7147 VSS.n7141 0.108269
R5029 VSS.n7364 VSS.n91 0.108269
R5030 VSS.n5694 VSS.n2427 0.108269
R5031 VSS.n5726 VSS.n2408 0.108269
R5032 VSS.n5758 VSS.n2389 0.108269
R5033 VSS.n4098 VSS.n3938 0.108269
R5034 VSS.n4075 VSS.n4074 0.108269
R5035 VSS.n4002 VSS.n3993 0.108269
R5036 VSS.n4715 VSS.n4105 0.108269
R5037 VSS.n4709 VSS.n4698 0.108269
R5038 VSS.n4133 VSS.n4122 0.108269
R5039 VSS.n4456 VSS.n4357 0.108269
R5040 VSS.n4411 VSS.n4367 0.108269
R5041 VSS.n4375 VSS.n4199 0.108269
R5042 VSS.n4609 VSS.n4204 0.108269
R5043 VSS.n5267 VSS.n3896 0.108269
R5044 VSS.n4351 VSS.n4281 0.108269
R5045 VSS.n4342 VSS.n4292 0.108269
R5046 VSS.n4659 VSS.n4258 0.108269
R5047 VSS.n4621 VSS.n4363 0.108269
R5048 VSS.n4960 VSS.n4956 0.108269
R5049 VSS.n4966 VSS.n4194 0.108269
R5050 VSS.n4813 VSS.n4193 0.108269
R5051 VSS.n4838 VSS.n4748 0.108269
R5052 VSS.n4930 VSS.n4746 0.108269
R5053 VSS.n4916 VSS.n4843 0.108269
R5054 VSS.n4915 VSS.n4119 0.108269
R5055 VSS.n5162 VSS.n4117 0.108269
R5056 VSS.n5122 VSS.n4128 0.108269
R5057 VSS.n4837 VSS.n4805 0.108269
R5058 VSS.n4831 VSS.n4827 0.108269
R5059 VSS.n4808 VSS.n4745 0.108269
R5060 VSS.n4680 VSS.n4225 0.108269
R5061 VSS.n4248 VSS.n4236 0.108269
R5062 VSS.n4676 VSS.n4673 0.108269
R5063 VSS.n4744 VSS.n4743 0.108269
R5064 VSS.n4697 VSS.n4693 0.108269
R5065 VSS.n4732 VSS.n4702 0.108269
R5066 VSS.n4710 VSS.n4704 0.108269
R5067 VSS.n5184 VSS.n4103 0.108269
R5068 VSS.n4250 VSS.n4241 0.108269
R5069 VSS.n4266 VSS.n4244 0.108269
R5070 VSS.n4670 VSS.n4239 0.108269
R5071 VSS.n4024 VSS.n4011 0.108269
R5072 VSS.n4014 VSS.n3910 0.108269
R5073 VSS.n4040 VSS.n4036 0.108269
R5074 VSS.n4023 VSS.n3996 0.108269
R5075 VSS.n4053 VSS.n4049 0.108269
R5076 VSS.n4065 VSS.n4062 0.108269
R5077 VSS.n4001 VSS.n3988 0.108269
R5078 VSS.n4092 VSS.n4088 0.108269
R5079 VSS.n4073 VSS.n3943 0.108269
R5080 VSS.n3947 VSS.n3937 0.108269
R5081 VSS.n4298 VSS.n3900 0.108269
R5082 VSS.n4033 VSS.n3908 0.108269
R5083 VSS.n5775 VSS.n2384 0.108269
R5084 VSS.n3958 VSS.n2386 0.108269
R5085 VSS.n5743 VSS.n2403 0.108269
R5086 VSS.n5194 VSS.n2405 0.108269
R5087 VSS.n5711 VSS.n2422 0.108269
R5088 VSS.n5132 VSS.n2424 0.108269
R5089 VSS.n5611 VSS.n5610 0.108269
R5090 VSS.n2587 VSS.n2548 0.108269
R5091 VSS.n2533 VSS.n2528 0.108269
R5092 VSS.n2581 VSS.n2577 0.108269
R5093 VSS.n2558 VSS.n2553 0.108269
R5094 VSS.n2544 VSS.n2530 0.108269
R5095 VSS.n2608 VSS.n2523 0.108269
R5096 VSS.n2615 VSS.n2611 0.108269
R5097 VSS.n5622 VSS.n5621 0.108269
R5098 VSS.n436 VSS.n425 0.108269
R5099 VSS.n7462 VSS.n310 0.108269
R5100 VSS.n667 VSS.n666 0.108269
R5101 VSS.n678 VSS.n677 0.108269
R5102 VSS.n778 VSS.n777 0.108269
R5103 VSS.n7189 VSS.n7085 0.108269
R5104 VSS.n638 VSS.n629 0.108269
R5105 VSS.n692 VSS.n342 0.108269
R5106 VSS.n7418 VSS.n340 0.108269
R5107 VSS.n7262 VSS.n697 0.108269
R5108 VSS.n7353 VSS.n7258 0.108269
R5109 VSS.n7360 VSS.n702 0.108269
R5110 VSS.n7607 VSS.n7606 0.108269
R5111 VSS.n691 VSS.n417 0.108269
R5112 VSS.n685 VSS.n681 0.108269
R5113 VSS.n420 VSS.n339 0.108269
R5114 VSS.n7126 VSS.n7124 0.108269
R5115 VSS.n7175 VSS.n7174 0.108269
R5116 VSS.n7123 VSS.n7119 0.108269
R5117 VSS.n7136 VSS.n7134 0.108269
R5118 VSS.n7163 VSS.n7132 0.108269
R5119 VSS.n7246 VSS.n7242 0.108269
R5120 VSS.n7146 VSS.n718 0.108269
R5121 VSS.n6898 VSS.n712 0.108269
R5122 VSS.n7096 VSS.n7089 0.108269
R5123 VSS.n7116 VSS.n7106 0.108269
R5124 VSS.n889 VSS.n848 0.108269
R5125 VSS.n843 VSS.n809 0.108269
R5126 VSS.n7027 VSS.n807 0.108269
R5127 VSS.n891 VSS.n884 0.108269
R5128 VSS.n901 VSS.n853 0.108269
R5129 VSS.n909 VSS.n874 0.108269
R5130 VSS.n7001 VSS.n872 0.108269
R5131 VSS.n6884 VSS.n919 0.108269
R5132 VSS.n6871 VSS.n6865 0.108269
R5133 VSS.n6943 VSS.n6858 0.108269
R5134 VSS.n826 VSS.n820 0.108269
R5135 VSS.n815 VSS.n806 0.108269
R5136 VSS.n7719 VSS.n27 0.108269
R5137 VSS.n6953 VSS.n29 0.108269
R5138 VSS.n7687 VSS.n46 0.108269
R5139 VSS.n6909 VSS.n48 0.108269
R5140 VSS.n7655 VSS.n65 0.108269
R5141 VSS.n83 VSS.n67 0.108269
R5142 VSS.n4451 VSS.n4450 0.105167
R5143 VSS.n5277 VSS.n2862 0.105167
R5144 VSS.n4320 VSS.n4308 0.105167
R5145 VSS.n4631 VSS.n4280 0.105167
R5146 VSS.n2596 VSS.n2537 0.105167
R5147 VSS.n2616 VSS.n2521 0.105167
R5148 VSS.n6669 VSS.n6663 0.105167
R5149 VSS.n7060 VSS.n783 0.105167
R5150 VSS.n768 VSS.n763 0.105167
R5151 VSS.n2726 VSS.n309 0.105167
R5152 VSS.n7636 VSS.n72 0.105167
R5153 VSS.n7637 VSS.n7636 0.105167
R5154 VSS.n7668 VSS.n53 0.105167
R5155 VSS.n55 VSS.n53 0.105167
R5156 VSS.n7669 VSS.n7668 0.105167
R5157 VSS.n7700 VSS.n34 0.105167
R5158 VSS.n36 VSS.n34 0.105167
R5159 VSS.n7701 VSS.n7700 0.105167
R5160 VSS.n7732 VSS.n15 0.105167
R5161 VSS.n17 VSS.n15 0.105167
R5162 VSS.n7733 VSS.n7732 0.105167
R5163 VSS.n5692 VSS.n2429 0.105167
R5164 VSS.n5693 VSS.n5692 0.105167
R5165 VSS.n5724 VSS.n2410 0.105167
R5166 VSS.n2412 VSS.n2410 0.105167
R5167 VSS.n5725 VSS.n5724 0.105167
R5168 VSS.n5756 VSS.n2391 0.105167
R5169 VSS.n2393 VSS.n2391 0.105167
R5170 VSS.n5757 VSS.n5756 0.105167
R5171 VSS.n5788 VSS.n2372 0.105167
R5172 VSS.n2374 VSS.n2372 0.105167
R5173 VSS.n5789 VSS.n5788 0.105167
R5174 VSS.n4457 VSS 0.105167
R5175 VSS.n3884 VSS 0.105167
R5176 VSS.n4313 VSS 0.105167
R5177 VSS.n4352 VSS 0.105167
R5178 VSS.n4435 VSS 0.105167
R5179 VSS.n5789 VSS 0.105167
R5180 VSS.n5757 VSS 0.105167
R5181 VSS.n5725 VSS 0.105167
R5182 VSS.n5693 VSS 0.105167
R5183 VSS VSS.n2491 0.105167
R5184 VSS VSS.n5623 0.105167
R5185 VSS.n2589 VSS.n2547 0.105167
R5186 VSS.n2589 VSS.n2588 0.105167
R5187 VSS.n2623 VSS.n2515 0.105167
R5188 VSS.n2624 VSS.n2623 0.105167
R5189 VSS.n2624 VSS.n2514 0.105167
R5190 VSS VSS.n2515 0.105167
R5191 VSS.n2557 VSS 0.105167
R5192 VSS.n2588 VSS 0.105167
R5193 VSS.n2547 VSS.n2546 0.105167
R5194 VSS VSS.n2609 0.105167
R5195 VSS.n5609 VSS 0.105167
R5196 VSS VSS.n2738 0.105167
R5197 VSS.n7463 VSS 0.105167
R5198 VSS.n6679 VSS 0.105167
R5199 VSS.n7052 VSS 0.105167
R5200 VSS.n776 VSS 0.105167
R5201 VSS.n7733 VSS 0.105167
R5202 VSS.n7701 VSS 0.105167
R5203 VSS.n7669 VSS 0.105167
R5204 VSS.n7637 VSS 0.105167
R5205 VSS.n151 VSS 0.105167
R5206 VSS.n6697 VSS.n6695 0.104667
R5207 VSS.n3869 VSS.n3868 0.104667
R5208 VSS.n4514 VSS.n4399 0.104667
R5209 VSS VSS.n4508 0.104667
R5210 VSS.n4569 VSS.n4568 0.104667
R5211 VSS.n4550 VSS 0.104667
R5212 VSS.n5019 VSS.n4187 0.104667
R5213 VSS VSS.n5013 0.104667
R5214 VSS.n5041 VSS.n5039 0.104667
R5215 VSS.n5658 VSS.n5657 0.104667
R5216 VSS.n2470 VSS 0.104667
R5217 VSS.n5087 VSS 0.104667
R5218 VSS VSS.n4877 0.104667
R5219 VSS.n3805 VSS.n2872 0.104667
R5220 VSS VSS.n3770 0.104667
R5221 VSS.n3708 VSS.n2881 0.104667
R5222 VSS VSS.n3672 0.104667
R5223 VSS.n3610 VSS.n2890 0.104667
R5224 VSS VSS.n3574 0.104667
R5225 VSS.n3513 VSS.n2901 0.104667
R5226 VSS VSS.n3477 0.104667
R5227 VSS.n3416 VSS.n2913 0.104667
R5228 VSS VSS.n3380 0.104667
R5229 VSS.n3319 VSS.n3318 0.104667
R5230 VSS.n5456 VSS.n5386 0.104667
R5231 VSS.n2575 VSS.n2574 0.104667
R5232 VSS VSS.n591 0.104667
R5233 VSS VSS.n7531 0.104667
R5234 VSS VSS.n493 0.104667
R5235 VSS.n382 VSS 0.104667
R5236 VSS.n224 VSS 0.104667
R5237 VSS VSS.n7570 0.104667
R5238 VSS VSS.n7318 0.104667
R5239 VSS.n6419 VSS.n1157 0.104667
R5240 VSS VSS.n6398 0.104667
R5241 VSS.n1296 VSS 0.104667
R5242 VSS VSS.n6836 0.104667
R5243 VSS.n6141 VSS.n6140 0.104667
R5244 VSS.n6177 VSS 0.104667
R5245 VSS.n1140 VSS.n1139 0.104146
R5246 VSS.n7750 VSS.n7749 0.103865
R5247 VSS.n4434 VSS.n4433 0.103365
R5248 VSS.n4513 VSS.n4512 0.103365
R5249 VSS.n4571 VSS.n4570 0.103365
R5250 VSS.n5018 VSS.n5017 0.103365
R5251 VSS.n4772 VSS.n4771 0.103365
R5252 VSS.n4857 VSS.n4856 0.103365
R5253 VSS.n5089 VSS.n5088 0.103365
R5254 VSS.n5660 VSS.n5659 0.103365
R5255 VSS.n3804 VSS.n3803 0.103365
R5256 VSS.n3707 VSS.n3706 0.103365
R5257 VSS.n3609 VSS.n3608 0.103365
R5258 VSS.n3512 VSS.n3511 0.103365
R5259 VSS.n3415 VSS.n3414 0.103365
R5260 VSS.n5352 VSS.n2817 0.103365
R5261 VSS.n5455 VSS.n5454 0.103365
R5262 VSS.n2741 VSS.n2740 0.103365
R5263 VSS.n384 VSS.n366 0.103365
R5264 VSS.n384 VSS.n383 0.103365
R5265 VSS.n6571 VSS.n6570 0.103365
R5266 VSS.n6504 VSS.n6503 0.103365
R5267 VSS.n6418 VSS.n6417 0.103365
R5268 VSS.n1293 VSS.n1260 0.103365
R5269 VSS.n6839 VSS.n940 0.103365
R5270 VSS.n6174 VSS.n6142 0.103365
R5271 VSS.n6094 VSS 0.103162
R5272 VSS.n1202 VSS 0.103162
R5273 VSS.n1337 VSS 0.103162
R5274 VSS.n1856 VSS 0.103162
R5275 VSS.n6352 VSS 0.103162
R5276 VSS.n1325 VSS 0.103002
R5277 VSS.n1355 VSS 0.103002
R5278 VSS.n1212 VSS 0.102841
R5279 VSS.n3769 VSS.n2873 0.102547
R5280 VSS.n3671 VSS.n2882 0.102547
R5281 VSS.n3573 VSS.n2891 0.102547
R5282 VSS.n3476 VSS.n2902 0.102547
R5283 VSS.n3379 VSS.n2914 0.102547
R5284 VSS.n2818 VSS.n2815 0.102547
R5285 VSS.n5421 VSS.n5387 0.102547
R5286 VSS.n1090 VSS.n1060 0.102547
R5287 VSS.n1124 VSS.n1107 0.102547
R5288 VSS.n1144 VSS.n1141 0.102547
R5289 VSS.n6397 VSS.n1158 0.102547
R5290 VSS.n1295 VSS.n1294 0.102547
R5291 VSS.n6835 VSS.n941 0.102547
R5292 VSS.n6176 VSS.n6175 0.102547
R5293 VSS.n5354 VSS 0.0999792
R5294 VSS VSS.n6551 0.0999792
R5295 VSS.n2346 VSS 0.0994583
R5296 VSS.n4770 VSS 0.0989375
R5297 VSS.n2134 VSS 0.0981562
R5298 VSS.n2140 VSS 0.0981562
R5299 VSS.n6267 VSS 0.0981562
R5300 VSS.n6273 VSS 0.0981562
R5301 VSS.n2219 VSS.n2113 0.0974697
R5302 VSS.n6278 VSS 0.0968542
R5303 VSS.n6290 VSS 0.0968542
R5304 VSS.n2230 VSS.n2229 0.0963763
R5305 VSS.n3806 VSS 0.095417
R5306 VSS.n3709 VSS 0.095417
R5307 VSS.n2493 VSS.n2492 0.0949964
R5308 VSS.n364 VSS.n363 0.0947708
R5309 VSS.n5626 VSS.n2507 0.0895625
R5310 VSS.n977 VSS.n976 0.0885208
R5311 VSS VSS.n6470 0.0874792
R5312 VSS.n3320 VSS 0.0871183
R5313 VSS VSS.n5422 0.0869583
R5314 VSS.n5457 VSS 0.0855622
R5315 VSS.n4335 VSS.n4294 0.0843334
R5316 VSS.n4277 VSS.n4274 0.0843334
R5317 VSS.n4954 VSS.n4205 0.0843334
R5318 VSS.n4474 VSS.n4403 0.0843334
R5319 VSS.n4794 VSS.n4790 0.0843334
R5320 VSS.n4825 VSS.n4212 0.0843334
R5321 VSS.n4671 VSS.n3920 0.0843334
R5322 VSS.n3913 VSS.n3911 0.0843334
R5323 VSS.n4034 VSS.n2855 0.0843334
R5324 VSS.n4047 VSS.n2851 0.0843334
R5325 VSS.n4060 VSS.n2847 0.0843334
R5326 VSS.n4086 VSS.n2842 0.0843334
R5327 VSS.n5265 VSS.n2859 0.0843334
R5328 VSS.n7200 VSS.n748 0.0843334
R5329 VSS.n636 VSS.n329 0.0843334
R5330 VSS.n7481 VSS.n305 0.0843334
R5331 VSS.n516 VSS.n512 0.0843334
R5332 VSS.n407 VSS.n402 0.0843334
R5333 VSS.n679 VSS.n332 0.0843334
R5334 VSS.n7117 VSS.n739 0.0843334
R5335 VSS.n7164 VSS.n734 0.0843334
R5336 VSS.n7187 VSS.n743 0.0843334
R5337 VSS.n7029 VSS.n804 0.0843334
R5338 VSS.n7015 VSS.n854 0.0843334
R5339 VSS.n7003 VSS.n869 0.0843334
R5340 VSS.n6989 VSS.n920 0.0843334
R5341 VSS.n6972 VSS.n934 0.0843334
R5342 VSS.n4593 VSS.n4589 0.0843334
R5343 VSS.n4980 VSS.n4192 0.0843334
R5344 VSS.n4901 VSS.n4897 0.0843334
R5345 VSS.n5114 VSS.n5107 0.0843334
R5346 VSS.n4932 VSS.n4217 0.0843334
R5347 VSS.n5164 VSS.n4113 0.0843334
R5348 VSS.n5180 VSS.n4106 0.0843334
R5349 VSS.n4691 VSS.n3925 0.0843334
R5350 VSS.n4733 VSS.n3930 0.0843334
R5351 VSS.n5213 VSS.n3934 0.0843334
R5352 VSS.n5332 VSS.n2834 0.0843334
R5353 VSS.n5777 VSS.n2380 0.0843334
R5354 VSS.n5745 VSS.n2399 0.0843334
R5355 VSS.n5713 VSS.n2418 0.0843334
R5356 VSS.n5678 VSS.n2436 0.0843334
R5357 VSS.n617 VSS.n612 0.0843334
R5358 VSS.n7450 VSS.n320 0.0843334
R5359 VSS.n7350 VSS.n7349 0.0843334
R5360 VSS.n7594 VSS.n7591 0.0843334
R5361 VSS.n7420 VSS.n337 0.0843334
R5362 VSS.n7406 VSS.n703 0.0843334
R5363 VSS.n7381 VSS.n709 0.0843334
R5364 VSS.n7240 VSS.n723 0.0843334
R5365 VSS.n6939 VSS.n6928 0.0843334
R5366 VSS.n7039 VSS.n795 0.0843334
R5367 VSS.n7721 VSS.n23 0.0843334
R5368 VSS.n7689 VSS.n42 0.0843334
R5369 VSS.n7657 VSS.n61 0.0843334
R5370 VSS.n187 VSS.n77 0.0843334
R5371 VSS.n5679 VSS.n2435 0.0842037
R5372 VSS.n78 VSS.n76 0.0842037
R5373 VSS.n4325 VSS.n4304 0.0842037
R5374 VSS.n4636 VSS.n4275 0.0842037
R5375 VSS.n4209 VSS.n4207 0.0842037
R5376 VSS.n4972 VSS.n4968 0.0842037
R5377 VSS.n4592 VSS.n4590 0.0842037
R5378 VSS.n4464 VSS.n4413 0.0842037
R5379 VSS.n5113 VSS.n5108 0.0842037
R5380 VSS.n4900 VSS.n4898 0.0842037
R5381 VSS.n4793 VSS.n4791 0.0842037
R5382 VSS.n5173 VSS.n4107 0.0842037
R5383 VSS.n4114 VSS.n4112 0.0842037
R5384 VSS.n4936 VSS.n4215 0.0842037
R5385 VSS.n4946 VSS.n4945 0.0842037
R5386 VSS.n5222 VSS.n3933 0.0842037
R5387 VSS.n5230 VSS.n3928 0.0842037
R5388 VSS.n5238 VSS.n3923 0.0842037
R5389 VSS.n5246 VSS.n3918 0.0842037
R5390 VSS.n3915 VSS.n3912 0.0842037
R5391 VSS.n5325 VSS.n2835 0.0842037
R5392 VSS.n5319 VSS.n5318 0.0842037
R5393 VSS.n5310 VSS.n5309 0.0842037
R5394 VSS.n5301 VSS.n5300 0.0842037
R5395 VSS.n5292 VSS.n5291 0.0842037
R5396 VSS.n5283 VSS.n5282 0.0842037
R5397 VSS.n2381 VSS.n2379 0.0842037
R5398 VSS.n2400 VSS.n2398 0.0842037
R5399 VSS.n2419 VSS.n2417 0.0842037
R5400 VSS.n749 VSS.n747 0.0842037
R5401 VSS.n324 VSS.n322 0.0842037
R5402 VSS.n7442 VSS.n327 0.0842037
R5403 VSS.n7471 VSS.n307 0.0842037
R5404 VSS.n616 VSS.n613 0.0842037
R5405 VSS.n515 VSS.n513 0.0842037
R5406 VSS.n7595 VSS.n7593 0.0842037
R5407 VSS.n7348 VSS.n7346 0.0842037
R5408 VSS.n406 VSS.n403 0.0842037
R5409 VSS.n7390 VSS.n708 0.0842037
R5410 VSS.n7399 VSS.n705 0.0842037
R5411 VSS.n7424 VSS.n335 0.0842037
R5412 VSS.n7434 VSS.n7433 0.0842037
R5413 VSS.n6932 VSS.n6929 0.0842037
R5414 VSS.n7233 VSS.n725 0.0842037
R5415 VSS.n7227 VSS.n7226 0.0842037
R5416 VSS.n7218 VSS.n7217 0.0842037
R5417 VSS.n7209 VSS.n7208 0.0842037
R5418 VSS.n6981 VSS.n933 0.0842037
R5419 VSS.n930 VSS.n922 0.0842037
R5420 VSS.n7007 VSS.n867 0.0842037
R5421 VSS.n864 VSS.n856 0.0842037
R5422 VSS.n7033 VSS.n802 0.0842037
R5423 VSS.n6674 VSS.n797 0.0842037
R5424 VSS.n24 VSS.n22 0.0842037
R5425 VSS.n43 VSS.n41 0.0842037
R5426 VSS.n62 VSS.n60 0.0842037
R5427 VSS.n4854 VSS.n4853 0.0838333
R5428 VSS.n3611 VSS 0.0834875
R5429 VSS.n6139 VSS 0.0826231
R5430 VSS.n7752 VSS 0.0826231
R5431 VSS.n3417 VSS 0.0824502
R5432 VSS.n6420 VSS 0.0821044
R5433 VSS.n2764 VSS.n2762 0.0819275
R5434 VSS.n1106 VSS.n1105 0.08175
R5435 VSS.n4515 VSS 0.0810055
R5436 VSS.n4567 VSS 0.0810055
R5437 VSS.n5020 VSS 0.0810055
R5438 VSS.n5042 VSS 0.0810055
R5439 VSS.n4333 VSS.n4305 0.0808942
R5440 VSS.n4644 VSS.n4276 0.0808942
R5441 VSS.n4952 VSS.n4208 0.0808942
R5442 VSS.n4978 VSS.n4977 0.0808942
R5443 VSS.n4601 VSS.n4600 0.0808942
R5444 VSS.n4472 VSS.n4471 0.0808942
R5445 VSS.n5119 VSS.n5111 0.0808942
R5446 VSS.n4909 VSS.n4908 0.0808942
R5447 VSS.n4802 VSS.n4801 0.0808942
R5448 VSS.n5181 VSS.n4109 0.0808942
R5449 VSS.n5166 VSS.n4111 0.0808942
R5450 VSS.n4224 VSS.n4223 0.0808942
R5451 VSS.n4943 VSS.n4942 0.0808942
R5452 VSS.n5216 VSS.n5215 0.0808942
R5453 VSS.n5228 VSS.n5227 0.0808942
R5454 VSS.n5236 VSS.n5235 0.0808942
R5455 VSS.n5244 VSS.n5243 0.0808942
R5456 VSS.n5252 VSS.n3914 0.0808942
R5457 VSS.n5333 VSS.n2837 0.0808942
R5458 VSS.n5322 VSS.n5321 0.0808942
R5459 VSS.n5313 VSS.n5312 0.0808942
R5460 VSS.n5304 VSS.n5303 0.0808942
R5461 VSS.n5295 VSS.n5294 0.0808942
R5462 VSS.n5286 VSS.n5285 0.0808942
R5463 VSS.n5779 VSS.n2378 0.0808942
R5464 VSS.n5747 VSS.n2397 0.0808942
R5465 VSS.n5715 VSS.n2416 0.0808942
R5466 VSS.n5681 VSS.n2433 0.0808942
R5467 VSS.n7202 VSS.n746 0.0808942
R5468 VSS.n7448 VSS.n323 0.0808942
R5469 VSS.n7440 VSS.n7439 0.0808942
R5470 VSS.n7479 VSS.n7478 0.0808942
R5471 VSS.n624 VSS.n623 0.0808942
R5472 VSS.n524 VSS.n523 0.0808942
R5473 VSS.n7603 VSS.n7602 0.0808942
R5474 VSS.n7342 VSS.n7338 0.0808942
R5475 VSS.n414 VSS.n413 0.0808942
R5476 VSS.n7384 VSS.n7383 0.0808942
R5477 VSS.n7404 VSS.n7403 0.0808942
R5478 VSS.n7396 VSS.n338 0.0808942
R5479 VSS.n7431 VSS.n7430 0.0808942
R5480 VSS.n6940 VSS.n6931 0.0808942
R5481 VSS.n7238 VSS.n7237 0.0808942
R5482 VSS.n7230 VSS.n7229 0.0808942
R5483 VSS.n7221 VSS.n7220 0.0808942
R5484 VSS.n7212 VSS.n7211 0.0808942
R5485 VSS.n6975 VSS.n6974 0.0808942
R5486 VSS.n6987 VSS.n923 0.0808942
R5487 VSS.n925 VSS.n870 0.0808942
R5488 VSS.n7013 VSS.n857 0.0808942
R5489 VSS.n859 VSS.n805 0.0808942
R5490 VSS.n7037 VSS.n7036 0.0808942
R5491 VSS.n7723 VSS.n21 0.0808942
R5492 VSS.n7691 VSS.n40 0.0808942
R5493 VSS.n7659 VSS.n59 0.0808942
R5494 VSS.n7623 VSS.n74 0.0808942
R5495 VSS.n6699 VSS 0.0794216
R5496 VSS VSS.n3865 0.0794216
R5497 VSS VSS.n3767 0.0794216
R5498 VSS VSS.n3669 0.0794216
R5499 VSS VSS.n3571 0.0794216
R5500 VSS VSS.n3474 0.0794216
R5501 VSS VSS.n3377 0.0794216
R5502 VSS.n5355 VSS 0.0794216
R5503 VSS VSS.n5420 0.0794216
R5504 VSS VSS.n6635 0.0794216
R5505 VSS VSS.n6550 0.0794216
R5506 VSS VSS.n6469 0.0794216
R5507 VSS VSS.n6395 0.0794216
R5508 VSS.n1298 VSS 0.0794216
R5509 VSS VSS.n6833 0.0794216
R5510 VSS.n6179 VSS 0.0794216
R5511 VSS.n1258 VSS.n1257 0.0791458
R5512 VSS.n3514 VSS 0.0789924
R5513 VSS.n5656 VSS 0.0785817
R5514 VSS.n2757 VSS.n2756 0.07852
R5515 VSS.n1140 VSS 0.076399
R5516 VSS VSS.n2382 0.0761666
R5517 VSS VSS.n2401 0.0761666
R5518 VSS VSS.n2420 0.0761666
R5519 VSS VSS.n2437 0.0761666
R5520 VSS VSS.n796 0.0761666
R5521 VSS VSS.n25 0.0761666
R5522 VSS VSS.n44 0.0761666
R5523 VSS VSS.n63 0.0761666
R5524 VSS.n7622 VSS 0.0761666
R5525 VSS.n3305 VSS.n2908 0.0757941
R5526 VSS.n6802 VSS.n6801 0.0757941
R5527 VSS.n4341 VSS.n4335 0.0746667
R5528 VSS.n4620 VSS.n4274 0.0746667
R5529 VSS.n4955 VSS.n4954 0.0746667
R5530 VSS.n4475 VSS.n4474 0.0746667
R5531 VSS.n4790 VSS.n4789 0.0746667
R5532 VSS.n4826 VSS.n4825 0.0746667
R5533 VSS.n4672 VSS.n4671 0.0746667
R5534 VSS.n4660 VSS.n3911 0.0746667
R5535 VSS.n4035 VSS.n4034 0.0746667
R5536 VSS.n4048 VSS.n4047 0.0746667
R5537 VSS.n4061 VSS.n4060 0.0746667
R5538 VSS.n4087 VSS.n4086 0.0746667
R5539 VSS.n5266 VSS.n5265 0.0746667
R5540 VSS.n7200 VSS.n7199 0.0746667
R5541 VSS.n637 VSS.n636 0.0746667
R5542 VSS.n7482 VSS.n7481 0.0746667
R5543 VSS.n512 VSS.n511 0.0746667
R5544 VSS.n402 VSS.n401 0.0746667
R5545 VSS.n680 VSS.n679 0.0746667
R5546 VSS.n7118 VSS.n7117 0.0746667
R5547 VSS.n7165 VSS.n7164 0.0746667
R5548 VSS.n7188 VSS.n7187 0.0746667
R5549 VSS.n7029 VSS.n7028 0.0746667
R5550 VSS.n7016 VSS.n7015 0.0746667
R5551 VSS.n7003 VSS.n7002 0.0746667
R5552 VSS.n6990 VSS.n6989 0.0746667
R5553 VSS.n6972 VSS.n6971 0.0746667
R5554 VSS.n4589 VSS.n4588 0.0739167
R5555 VSS VSS.n4603 0.0739167
R5556 VSS.n4303 VSS 0.0739167
R5557 VSS VSS.n4646 0.0739167
R5558 VSS VSS.n4206 0.0739167
R5559 VSS.n4981 VSS.n4980 0.0739167
R5560 VSS.n4967 VSS 0.0739167
R5561 VSS.n4412 VSS 0.0739167
R5562 VSS.n4897 VSS.n4896 0.0739167
R5563 VSS VSS.n4911 0.0739167
R5564 VSS.n5107 VSS.n5106 0.0739167
R5565 VSS VSS.n5121 0.0739167
R5566 VSS VSS.n4804 0.0739167
R5567 VSS.n4932 VSS.n4931 0.0739167
R5568 VSS.n4934 VSS 0.0739167
R5569 VSS.n5164 VSS.n5163 0.0739167
R5570 VSS VSS.n4115 0.0739167
R5571 VSS.n5150 VSS.n4106 0.0739167
R5572 VSS VSS.n5183 0.0739167
R5573 VSS VSS.n4249 0.0739167
R5574 VSS VSS.n4019 0.0739167
R5575 VSS.n4692 VSS.n4691 0.0739167
R5576 VSS VSS.n3998 0.0739167
R5577 VSS.n4734 VSS.n4733 0.0739167
R5578 VSS VSS.n4069 0.0739167
R5579 VSS.n5213 VSS.n5212 0.0739167
R5580 VSS.n4099 VSS 0.0739167
R5581 VSS VSS.n5254 0.0739167
R5582 VSS VSS.n3675 0.0739167
R5583 VSS VSS.n3577 0.0739167
R5584 VSS VSS.n3480 0.0739167
R5585 VSS VSS.n3383 0.0739167
R5586 VSS.n3976 VSS.n2834 0.0739167
R5587 VSS VSS.n5335 0.0739167
R5588 VSS VSS.n3788 0.0739167
R5589 VSS.n5777 VSS.n5776 0.0739167
R5590 VSS.n5745 VSS.n5744 0.0739167
R5591 VSS.n5713 VSS.n5712 0.0739167
R5592 VSS.n5678 VSS.n5677 0.0739167
R5593 VSS.n612 VSS.n611 0.0739167
R5594 VSS VSS.n626 0.0739167
R5595 VSS VSS.n750 0.0739167
R5596 VSS.n7451 VSS.n7450 0.0739167
R5597 VSS VSS.n321 0.0739167
R5598 VSS VSS.n7095 0.0739167
R5599 VSS VSS.n306 0.0739167
R5600 VSS VSS.n526 0.0739167
R5601 VSS.n7350 VSS.n7337 0.0739167
R5602 VSS VSS.n7352 0.0739167
R5603 VSS.n7591 VSS.n7590 0.0739167
R5604 VSS VSS.n7605 0.0739167
R5605 VSS VSS.n416 0.0739167
R5606 VSS.n7420 VSS.n7419 0.0739167
R5607 VSS.n7422 VSS 0.0739167
R5608 VSS.n7407 VSS.n7406 0.0739167
R5609 VSS VSS.n704 0.0739167
R5610 VSS.n7381 VSS.n7380 0.0739167
R5611 VSS.n7253 VSS 0.0739167
R5612 VSS VSS.n7176 0.0739167
R5613 VSS VSS.n890 0.0739167
R5614 VSS VSS.n908 0.0739167
R5615 VSS.n7241 VSS.n7240 0.0739167
R5616 VSS VSS.n724 0.0739167
R5617 VSS.n6928 VSS.n6927 0.0739167
R5618 VSS VSS.n6942 0.0739167
R5619 VSS VSS.n811 0.0739167
R5620 VSS.n7031 VSS 0.0739167
R5621 VSS VSS.n855 0.0739167
R5622 VSS.n7005 VSS 0.0739167
R5623 VSS VSS.n921 0.0739167
R5624 VSS.n6854 VSS 0.0739167
R5625 VSS.n7040 VSS.n7039 0.0739167
R5626 VSS.n7721 VSS.n7720 0.0739167
R5627 VSS.n7689 VSS.n7688 0.0739167
R5628 VSS.n7657 VSS.n7656 0.0739167
R5629 VSS.n188 VSS.n187 0.0739167
R5630 VSS.n364 VSS 0.0734889
R5631 VSS.n6642 VSS.n6641 0.072375
R5632 VSS.n977 VSS 0.0712123
R5633 VSS.n6636 VSS.n1089 0.0702917
R5634 VSS.n4854 VSS 0.0697521
R5635 VSS.n1106 VSS 0.0689647
R5636 VSS VSS.n6636 0.0687292
R5637 VSS.n1258 VSS 0.0681003
R5638 VSS.n552 VSS.n551 0.0676875
R5639 VSS.n6659 VSS.n6658 0.066646
R5640 VSS.n6642 VSS 0.0658527
R5641 VSS.n6372 VSS.n6366 0.0652425
R5642 VSS.n6122 VSS.n6100 0.065125
R5643 VSS.n155 VSS.n153 0.0650833
R5644 VSS.n251 VSS.n93 0.0650833
R5645 VSS.n7279 VSS.n7278 0.0650833
R5646 VSS.n217 VSS.n216 0.0650833
R5647 VSS.n6366 VSS.n6365 0.0647725
R5648 VSS.n493 VSS.n491 0.0645625
R5649 VSS.n1323 VSS.n1322 0.0635975
R5650 VSS.n6661 VSS 0.063
R5651 VSS.n4418 VSS 0.063
R5652 VSS.n4416 VSS 0.063
R5653 VSS.n4503 VSS 0.063
R5654 VSS.n4533 VSS 0.063
R5655 VSS.n5008 VSS 0.063
R5656 VSS.n4752 VSS 0.063
R5657 VSS.n2453 VSS 0.063
R5658 VSS.n3869 VSS 0.063
R5659 VSS.n2893 VSS 0.063
R5660 VSS.n2904 VSS 0.063
R5661 VSS.n2916 VSS 0.063
R5662 VSS.n2814 VSS 0.063
R5663 VSS.n5389 VSS 0.063
R5664 VSS.n5805 VSS 0.063
R5665 VSS.n2507 VSS 0.063
R5666 VSS.n5624 VSS 0.063
R5667 VSS.n2573 VSS 0.063
R5668 VSS.n2565 VSS 0.063
R5669 VSS.n2575 VSS 0.063
R5670 VSS.n5607 VSS 0.063
R5671 VSS.n2722 VSS 0.063
R5672 VSS.n2739 VSS 0.063
R5673 VSS.n6695 VSS 0.063
R5674 VSS.n1089 VSS 0.063
R5675 VSS.n1123 VSS 0.063
R5676 VSS.n1143 VSS 0.063
R5677 VSS.n1174 VSS 0.063
R5678 VSS.n1233 VSS 0.063
R5679 VSS.n957 VSS 0.063
R5680 VSS.n7748 VSS 0.063
R5681 VSS.n6103 VSS 0.063
R5682 VSS.n153 VSS 0.063
R5683 VSS.n5607 VSS.n5606 0.0609167
R5684 VSS VSS.n1138 0.0607775
R5685 VSS.n2261 VSS 0.0603958
R5686 VSS.n2289 VSS 0.0603958
R5687 VSS.n2317 VSS 0.0603958
R5688 VSS VSS.n2246 0.0603958
R5689 VSS VSS.n2245 0.0603958
R5690 VSS VSS.n2244 0.0603958
R5691 VSS.n2355 VSS 0.0603958
R5692 VSS VSS.n2135 0.0603958
R5693 VSS.n2136 VSS 0.0603958
R5694 VSS.n2141 VSS 0.0603958
R5695 VSS VSS.n2121 0.0603958
R5696 VSS.n2153 VSS 0.0603958
R5697 VSS VSS.n2118 0.0603958
R5698 VSS.n2165 VSS 0.0603958
R5699 VSS.n2168 VSS 0.0603958
R5700 VSS VSS.n6268 0.0603958
R5701 VSS.n6269 VSS 0.0603958
R5702 VSS VSS.n6274 0.0603958
R5703 VSS.n6275 VSS 0.0603958
R5704 VSS VSS.n6286 0.0603958
R5705 VSS.n6287 VSS 0.0603958
R5706 VSS.n6298 VSS 0.0603958
R5707 VSS.n6301 VSS 0.0603958
R5708 VSS.n6829 VSS.n958 0.0603075
R5709 VSS.n6182 VSS.n6100 0.0603075
R5710 VSS.n5825 VSS.n5824 0.0600725
R5711 VSS.n1217 VSS.n1216 0.0598752
R5712 VSS.n455 VSS.n454 0.0593542
R5713 VSS VSS.n6698 0.0593235
R5714 VSS.n3866 VSS 0.0593235
R5715 VSS.n4431 VSS 0.0593235
R5716 VSS.n4506 VSS 0.0593235
R5717 VSS.n4551 VSS 0.0593235
R5718 VSS.n5011 VSS 0.0593235
R5719 VSS.n4770 VSS 0.0593235
R5720 VSS.n4155 VSS 0.0593235
R5721 VSS.n2471 VSS 0.0593235
R5722 VSS.n5086 VSS 0.0593235
R5723 VSS.n4875 VSS 0.0593235
R5724 VSS.n3768 VSS 0.0593235
R5725 VSS.n3670 VSS 0.0593235
R5726 VSS.n3572 VSS 0.0593235
R5727 VSS.n3475 VSS 0.0593235
R5728 VSS.n3378 VSS 0.0593235
R5729 VSS VSS.n5354 0.0593235
R5730 VSS.n5422 VSS 0.0593235
R5731 VSS.n5626 VSS 0.0593235
R5732 VSS.n5606 VSS 0.0593235
R5733 VSS.n2743 VSS 0.0593235
R5734 VSS.n551 VSS 0.0593235
R5735 VSS.n454 VSS 0.0593235
R5736 VSS.n589 VSS 0.0593235
R5737 VSS.n7529 VSS 0.0593235
R5738 VSS.n7539 VSS 0.0593235
R5739 VSS.n491 VSS 0.0593235
R5740 VSS.n261 VSS 0.0593235
R5741 VSS.n7278 VSS 0.0593235
R5742 VSS.n251 VSS 0.0593235
R5743 VSS.n216 VSS 0.0593235
R5744 VSS.n225 VSS 0.0593235
R5745 VSS.n7568 VSS 0.0593235
R5746 VSS.n7316 VSS 0.0593235
R5747 VSS.n6636 VSS 0.0593235
R5748 VSS.n6551 VSS 0.0593235
R5749 VSS.n6470 VSS 0.0593235
R5750 VSS.n6396 VSS 0.0593235
R5751 VSS VSS.n1297 0.0593235
R5752 VSS.n6834 VSS 0.0593235
R5753 VSS VSS.n6178 0.0593235
R5754 VSS.n155 VSS 0.0593235
R5755 VSS.n1349 VSS.n1348 0.0584275
R5756 VSS.n591 VSS.n589 0.0583125
R5757 VSS.n975 VSS.n958 0.05737
R5758 VSS.n1098 VSS.n1097 0.057271
R5759 VSS.n3806 VSS.n3805 0.0572708
R5760 VSS.n3709 VSS.n3708 0.0572708
R5761 VSS.n5786 VSS.n5785 0.0564896
R5762 VSS.n5754 VSS.n5753 0.0564896
R5763 VSS.n5722 VSS.n5721 0.0564896
R5764 VSS.n2592 VSS.n2591 0.0564896
R5765 VSS.n2621 VSS.n2620 0.0564896
R5766 VSS.n7730 VSS.n7729 0.0564896
R5767 VSS.n7698 VSS.n7697 0.0564896
R5768 VSS.n7666 VSS.n7665 0.0564896
R5769 VSS.n82 VSS.n80 0.0560583
R5770 VSS.n6908 VSS.n6906 0.0560583
R5771 VSS.n6952 VSS.n6950 0.0560583
R5772 VSS.n5131 VSS.n5129 0.0560583
R5773 VSS.n5193 VSS.n5191 0.0560583
R5774 VSS.n3957 VSS.n3955 0.0560583
R5775 VSS.n4265 VSS.n4263 0.0560583
R5776 VSS.n4455 VSS.n4453 0.0560583
R5777 VSS.n4410 VSS.n4408 0.0560583
R5778 VSS.n4374 VSS.n4372 0.0560583
R5779 VSS.n4297 VSS.n4295 0.0560583
R5780 VSS.n4311 VSS.n4309 0.0560583
R5781 VSS.n4350 VSS.n4282 0.0560583
R5782 VSS.n4651 VSS.n4650 0.0560583
R5783 VSS.n4817 VSS.n4816 0.0560583
R5784 VSS.n4841 VSS.n4840 0.0560583
R5785 VSS.n4914 VSS.n4912 0.0560583
R5786 VSS.n5125 VSS.n5124 0.0560583
R5787 VSS.n4247 VSS.n4235 0.0560583
R5788 VSS.n4229 VSS.n4226 0.0560583
R5789 VSS.n4713 VSS.n4712 0.0560583
R5790 VSS.n5187 VSS.n5186 0.0560583
R5791 VSS.n4018 VSS.n4017 0.0560583
R5792 VSS.n4022 VSS.n4020 0.0560583
R5793 VSS.n4000 VSS.n3987 0.0560583
R5794 VSS.n4072 VSS.n4070 0.0560583
R5795 VSS.n3951 VSS.n3950 0.0560583
R5796 VSS.n5618 VSS.n2509 0.0560583
R5797 VSS.n2561 VSS.n2560 0.0560583
R5798 VSS.n2607 VSS.n2524 0.0560583
R5799 VSS.n435 VSS.n433 0.0560583
R5800 VSS.n7099 VSS.n7098 0.0560583
R5801 VSS.n7461 VSS.n311 0.0560583
R5802 VSS.n670 VSS.n669 0.0560583
R5803 VSS.n829 VSS.n828 0.0560583
R5804 VSS.n7050 VSS.n786 0.0560583
R5805 VSS.n781 VSS.n780 0.0560583
R5806 VSS.n7079 VSS.n7078 0.0560583
R5807 VSS.n652 VSS.n651 0.0560583
R5808 VSS.n695 VSS.n694 0.0560583
R5809 VSS.n7354 VSS.n7257 0.0560583
R5810 VSS.n7610 VSS.n7609 0.0560583
R5811 VSS.n7111 VSS.n7108 0.0560583
R5812 VSS.n7139 VSS.n7138 0.0560583
R5813 VSS.n7145 VSS.n7143 0.0560583
R5814 VSS.n6902 VSS.n6901 0.0560583
R5815 VSS.n846 VSS.n845 0.0560583
R5816 VSS.n894 VSS.n893 0.0560583
R5817 VSS.n912 VSS.n911 0.0560583
R5818 VSS.n6874 VSS.n6873 0.0560583
R5819 VSS.n6946 VSS.n6945 0.0560583
R5820 VSS.n1349 VSS.n1104 0.0558425
R5821 VSS VSS.n1341 0.055725
R5822 VSS.n1323 VSS.n1226 0.0553725
R5823 VSS.n4849 VSS.n4848 0.0551877
R5824 VSS.n7647 VSS.n7646 0.0545568
R5825 VSS.n7679 VSS.n7678 0.0545568
R5826 VSS.n7711 VSS.n7710 0.0545568
R5827 VSS.n6994 VSS.n6993 0.0545568
R5828 VSS.n882 VSS.n881 0.0545568
R5829 VSS.n5703 VSS.n5702 0.0545568
R5830 VSS.n5735 VSS.n5734 0.0545568
R5831 VSS.n5767 VSS.n5766 0.0545568
R5832 VSS.n4058 VSS.n3992 0.0545568
R5833 VSS.n4823 VSS.n4821 0.0545568
R5834 VSS.n4406 VSS.n4404 0.0545568
R5835 VSS.n4607 VSS.n4606 0.0545568
R5836 VSS.n4612 VSS.n4611 0.0545568
R5837 VSS.n4618 VSS.n4366 0.0545568
R5838 VSS.n5275 VSS.n3888 0.0545568
R5839 VSS.n4301 VSS.n4299 0.0545568
R5840 VSS.n5269 VSS.n5268 0.0545568
R5841 VSS.n4290 VSS.n4289 0.0545568
R5842 VSS.n4344 VSS.n4343 0.0545568
R5843 VSS.n4318 VSS.n4316 0.0545568
R5844 VSS.n4339 VSS.n4271 0.0545568
R5845 VSS.n4270 VSS.n4269 0.0545568
R5846 VSS.n4658 VSS.n4259 0.0545568
R5847 VSS.n4623 VSS.n4622 0.0545568
R5848 VSS.n4629 VSS.n4356 0.0545568
R5849 VSS.n4958 VSS.n4957 0.0545568
R5850 VSS.n4965 VSS.n4195 0.0545568
R5851 VSS.n4923 VSS.n4922 0.0545568
R5852 VSS.n4929 VSS.n4747 0.0545568
R5853 VSS.n4919 VSS.n4918 0.0545568
R5854 VSS.n5154 VSS.n5153 0.0545568
R5855 VSS.n5161 VSS.n4118 0.0545568
R5856 VSS.n4132 VSS.n4130 0.0545568
R5857 VSS.n5148 VSS.n4127 0.0545568
R5858 VSS.n5136 VSS.n5135 0.0545568
R5859 VSS.n5141 VSS.n5140 0.0545568
R5860 VSS.n4836 VSS.n4806 0.0545568
R5861 VSS.n4829 VSS.n4828 0.0545568
R5862 VSS.n4811 VSS.n4810 0.0545568
R5863 VSS.n4686 VSS.n4232 0.0545568
R5864 VSS.n4674 VSS.n4234 0.0545568
R5865 VSS.n4683 VSS.n4682 0.0545568
R5866 VSS.n4738 VSS.n4737 0.0545568
R5867 VSS.n4695 VSS.n4694 0.0545568
R5868 VSS.n4708 VSS.n4706 0.0545568
R5869 VSS.n4724 VSS.n4723 0.0545568
R5870 VSS.n4731 VSS.n4703 0.0545568
R5871 VSS.n4719 VSS.n4718 0.0545568
R5872 VSS.n5210 VSS.n4102 0.0545568
R5873 VSS.n5198 VSS.n5197 0.0545568
R5874 VSS.n5203 VSS.n5202 0.0545568
R5875 VSS.n4253 VSS.n4252 0.0545568
R5876 VSS.n4662 VSS.n4661 0.0545568
R5877 VSS.n4669 VSS.n4240 0.0545568
R5878 VSS.n4045 VSS.n4010 0.0545568
R5879 VSS.n4038 VSS.n4037 0.0545568
R5880 VSS.n4027 VSS.n4026 0.0545568
R5881 VSS.n4051 VSS.n4050 0.0545568
R5882 VSS.n4005 VSS.n4004 0.0545568
R5883 VSS.n4081 VSS.n3984 0.0545568
R5884 VSS.n4063 VSS.n3986 0.0545568
R5885 VSS.n4078 VSS.n4077 0.0545568
R5886 VSS.n3980 VSS.n3979 0.0545568
R5887 VSS.n4090 VSS.n4089 0.0545568
R5888 VSS.n4097 VSS.n3939 0.0545568
R5889 VSS.n3974 VSS.n3946 0.0545568
R5890 VSS.n3962 VSS.n3961 0.0545568
R5891 VSS.n3967 VSS.n3966 0.0545568
R5892 VSS.n5258 VSS.n5257 0.0545568
R5893 VSS.n3903 VSS.n3898 0.0545568
R5894 VSS.n4032 VSS.n3909 0.0545568
R5895 VSS.n5774 VSS.n2385 0.0545568
R5896 VSS.n5761 VSS.n5760 0.0545568
R5897 VSS.n5742 VSS.n2404 0.0545568
R5898 VSS.n5729 VSS.n5728 0.0545568
R5899 VSS.n5710 VSS.n2423 0.0545568
R5900 VSS.n5697 VSS.n5696 0.0545568
R5901 VSS.n2626 VSS.n2512 0.0545568
R5902 VSS.n2536 VSS.n2535 0.0545568
R5903 VSS.n2600 VSS.n2599 0.0545568
R5904 VSS.n2569 VSS.n2567 0.0545568
R5905 VSS.n2579 VSS.n2578 0.0545568
R5906 VSS.n2586 VSS.n2549 0.0545568
R5907 VSS.n2543 VSS.n2532 0.0545568
R5908 VSS.n2614 VSS.n2511 0.0545568
R5909 VSS.n5614 VSS.n5613 0.0545568
R5910 VSS.n647 VSS.n645 0.0545568
R5911 VSS.n634 VSS.n532 0.0545568
R5912 VSS.n531 VSS.n432 0.0545568
R5913 VSS.n674 VSS.n430 0.0545568
R5914 VSS.n664 VSS.n628 0.0545568
R5915 VSS.n657 VSS.n656 0.0545568
R5916 VSS.n6667 VSS.n6665 0.0545568
R5917 VSS.n824 VSS.n822 0.0545568
R5918 VSS.n7043 VSS.n7042 0.0545568
R5919 VSS.n760 VSS.n756 0.0545568
R5920 VSS.n7070 VSS.n7069 0.0545568
R5921 VSS.n7065 VSS.n7064 0.0545568
R5922 VSS.n7197 VSS.n753 0.0545568
R5923 VSS.n7093 VSS.n7091 0.0545568
R5924 VSS.n7191 VSS.n7190 0.0545568
R5925 VSS.n7454 VSS.n7453 0.0545568
R5926 VSS.n766 VSS.n764 0.0545568
R5927 VSS.n641 VSS.n640 0.0545568
R5928 VSS.n7411 VSS.n7410 0.0545568
R5929 VSS.n7417 VSS.n341 0.0545568
R5930 VSS.n7261 VSS.n7259 0.0545568
R5931 VSS.n7370 VSS.n7254 0.0545568
R5932 VSS.n7358 VSS.n7256 0.0545568
R5933 VSS.n7367 VSS.n7366 0.0545568
R5934 VSS.n7378 VSS.n89 0.0545568
R5935 VSS.n88 VSS.n84 0.0545568
R5936 VSS.n7616 VSS.n7615 0.0545568
R5937 VSS.n690 VSS.n418 0.0545568
R5938 VSS.n683 VSS.n682 0.0545568
R5939 VSS.n423 VSS.n422 0.0545568
R5940 VSS.n7169 VSS.n7168 0.0545568
R5941 VSS.n7121 VSS.n7120 0.0545568
R5942 VSS.n7129 VSS.n7128 0.0545568
R5943 VSS.n7155 VSS.n7154 0.0545568
R5944 VSS.n7162 VSS.n7133 0.0545568
R5945 VSS.n7150 VSS.n7149 0.0545568
R5946 VSS.n6894 VSS.n6892 0.0545568
R5947 VSS.n7244 VSS.n7243 0.0545568
R5948 VSS.n7251 VSS.n714 0.0545568
R5949 VSS.n6925 VSS.n6897 0.0545568
R5950 VSS.n6913 VSS.n6912 0.0545568
R5951 VSS.n6918 VSS.n6917 0.0545568
R5952 VSS.n7180 VSS.n7179 0.0545568
R5953 VSS.n7101 VSS.n7087 0.0545568
R5954 VSS.n7115 VSS.n7107 0.0545568
R5955 VSS.n7020 VSS.n7019 0.0545568
R5956 VSS.n7026 VSS.n808 0.0545568
R5957 VSS.n888 VSS.n886 0.0545568
R5958 VSS.n899 VSS.n898 0.0545568
R5959 VSS.n906 VSS.n877 0.0545568
R5960 VSS.n7000 VSS.n873 0.0545568
R5961 VSS.n6869 VSS.n6867 0.0545568
R5962 VSS.n6877 VSS.n6876 0.0545568
R5963 VSS.n6882 VSS.n6881 0.0545568
R5964 VSS.n6889 VSS.n6861 0.0545568
R5965 VSS.n6969 VSS.n6857 0.0545568
R5966 VSS.n6957 VSS.n6956 0.0545568
R5967 VSS.n6962 VSS.n6961 0.0545568
R5968 VSS.n841 VSS.n813 0.0545568
R5969 VSS.n834 VSS.n833 0.0545568
R5970 VSS.n818 VSS.n817 0.0545568
R5971 VSS.n7718 VSS.n28 0.0545568
R5972 VSS.n7705 VSS.n7704 0.0545568
R5973 VSS.n7686 VSS.n47 0.0545568
R5974 VSS.n7673 VSS.n7672 0.0545568
R5975 VSS.n7654 VSS.n66 0.0545568
R5976 VSS.n7641 VSS.n7640 0.0545568
R5977 VSS.n1359 VSS 0.0542143
R5978 VSS.n1 VSS 0.0539905
R5979 VSS.n1195 VSS 0.0539905
R5980 VSS.n1185 VSS 0.0539905
R5981 VSS.n1180 VSS 0.0539905
R5982 VSS.n1189 VSS 0.0537667
R5983 VSS.n1329 VSS 0.0537667
R5984 VSS.n6356 VSS 0.0537667
R5985 VSS.n6648 VSS.n1038 0.0537275
R5986 VSS.n7622 VSS.n79 0.0530835
R5987 VSS.n7658 VSS.n63 0.0530835
R5988 VSS.n7690 VSS.n44 0.0530835
R5989 VSS.n7722 VSS.n25 0.0530835
R5990 VSS.n7038 VSS.n796 0.0530835
R5991 VSS.n5680 VSS.n2437 0.0530835
R5992 VSS.n5714 VSS.n2420 0.0530835
R5993 VSS.n5746 VSS.n2401 0.0530835
R5994 VSS.n5778 VSS.n2382 0.0530835
R5995 VSS.n2382 VSS 0.0530835
R5996 VSS.n2401 VSS 0.0530835
R5997 VSS.n2420 VSS 0.0530835
R5998 VSS.n2437 VSS 0.0530835
R5999 VSS VSS.n796 0.0530835
R6000 VSS.n25 VSS 0.0530835
R6001 VSS.n44 VSS 0.0530835
R6002 VSS.n63 VSS 0.0530835
R6003 VSS VSS.n7622 0.0530835
R6004 VSS VSS.n4592 0.0530834
R6005 VSS VSS.n4325 0.0530834
R6006 VSS VSS.n4636 0.0530834
R6007 VSS VSS.n4209 0.0530834
R6008 VSS VSS.n4972 0.0530834
R6009 VSS VSS.n4464 0.0530834
R6010 VSS VSS.n4900 0.0530834
R6011 VSS VSS.n5113 0.0530834
R6012 VSS VSS.n4793 0.0530834
R6013 VSS.n4936 VSS 0.0530834
R6014 VSS VSS.n4112 0.0530834
R6015 VSS VSS.n5173 0.0530834
R6016 VSS.n4946 VSS 0.0530834
R6017 VSS.n5246 VSS 0.0530834
R6018 VSS.n5238 VSS 0.0530834
R6019 VSS.n5230 VSS 0.0530834
R6020 VSS.n5222 VSS 0.0530834
R6021 VSS VSS.n3915 0.0530834
R6022 VSS.n5291 VSS 0.0530834
R6023 VSS.n5300 VSS 0.0530834
R6024 VSS.n5309 VSS 0.0530834
R6025 VSS.n5318 VSS 0.0530834
R6026 VSS VSS.n5325 0.0530834
R6027 VSS.n5282 VSS 0.0530834
R6028 VSS VSS.n2379 0.0530834
R6029 VSS VSS.n2398 0.0530834
R6030 VSS VSS.n2417 0.0530834
R6031 VSS VSS.n2435 0.0530834
R6032 VSS VSS.n616 0.0530834
R6033 VSS VSS.n747 0.0530834
R6034 VSS VSS.n324 0.0530834
R6035 VSS.n7442 VSS 0.0530834
R6036 VSS VSS.n7471 0.0530834
R6037 VSS VSS.n515 0.0530834
R6038 VSS.n7346 VSS 0.0530834
R6039 VSS VSS.n7593 0.0530834
R6040 VSS VSS.n406 0.0530834
R6041 VSS.n7424 VSS 0.0530834
R6042 VSS VSS.n7399 0.0530834
R6043 VSS.n7390 VSS 0.0530834
R6044 VSS.n7434 VSS 0.0530834
R6045 VSS.n7217 VSS 0.0530834
R6046 VSS.n7226 VSS 0.0530834
R6047 VSS VSS.n7233 0.0530834
R6048 VSS VSS.n6932 0.0530834
R6049 VSS.n7208 VSS 0.0530834
R6050 VSS.n7033 VSS 0.0530834
R6051 VSS VSS.n864 0.0530834
R6052 VSS.n7007 VSS 0.0530834
R6053 VSS VSS.n930 0.0530834
R6054 VSS.n6981 VSS 0.0530834
R6055 VSS.n6674 VSS 0.0530834
R6056 VSS VSS.n22 0.0530834
R6057 VSS VSS.n41 0.0530834
R6058 VSS VSS.n60 0.0530834
R6059 VSS VSS.n76 0.0530834
R6060 VSS.n6973 VSS.n6854 0.0530834
R6061 VSS.n6988 VSS.n921 0.0530834
R6062 VSS.n7005 VSS.n7004 0.0530834
R6063 VSS.n7014 VSS.n855 0.0530834
R6064 VSS.n7031 VSS.n7030 0.0530834
R6065 VSS.n811 VSS.n742 0.0530834
R6066 VSS.n6942 VSS.n6941 0.0530834
R6067 VSS.n7239 VSS.n724 0.0530834
R6068 VSS.n908 VSS.n733 0.0530834
R6069 VSS.n890 VSS.n738 0.0530834
R6070 VSS.n7176 VSS.n333 0.0530834
R6071 VSS.n7382 VSS.n7253 0.0530834
R6072 VSS.n7405 VSS.n704 0.0530834
R6073 VSS.n7422 VSS.n7421 0.0530834
R6074 VSS.n416 VSS.n415 0.0530834
R6075 VSS.n7605 VSS.n7604 0.0530834
R6076 VSS.n7352 VSS.n7351 0.0530834
R6077 VSS.n3788 VSS.n2858 0.0530834
R6078 VSS.n5335 VSS.n5334 0.0530834
R6079 VSS.n3383 VSS.n2841 0.0530834
R6080 VSS.n3480 VSS.n2846 0.0530834
R6081 VSS.n3577 VSS.n2850 0.0530834
R6082 VSS.n3675 VSS.n2854 0.0530834
R6083 VSS.n5254 VSS.n5253 0.0530834
R6084 VSS.n5214 VSS.n4099 0.0530834
R6085 VSS.n4069 VSS.n3931 0.0530834
R6086 VSS.n3998 VSS.n3926 0.0530834
R6087 VSS.n4019 VSS.n3921 0.0530834
R6088 VSS.n4249 VSS.n4213 0.0530834
R6089 VSS.n5183 VSS.n5182 0.0530834
R6090 VSS.n5165 VSS.n4115 0.0530834
R6091 VSS.n4934 VSS.n4933 0.0530834
R6092 VSS.n4804 VSS.n4803 0.0530834
R6093 VSS.n5121 VSS.n5120 0.0530834
R6094 VSS.n4911 VSS.n4910 0.0530834
R6095 VSS.n4473 VSS.n4412 0.0530834
R6096 VSS.n4979 VSS.n4967 0.0530834
R6097 VSS.n4603 VSS.n4602 0.0530834
R6098 VSS.n4603 VSS 0.0530834
R6099 VSS.n4646 VSS.n4645 0.0530834
R6100 VSS.n4334 VSS.n4303 0.0530834
R6101 VSS VSS.n4303 0.0530834
R6102 VSS.n4646 VSS 0.0530834
R6103 VSS.n4953 VSS.n4206 0.0530834
R6104 VSS VSS.n4206 0.0530834
R6105 VSS VSS.n4967 0.0530834
R6106 VSS VSS.n4412 0.0530834
R6107 VSS.n4911 VSS 0.0530834
R6108 VSS.n5121 VSS 0.0530834
R6109 VSS.n4804 VSS 0.0530834
R6110 VSS VSS.n4934 0.0530834
R6111 VSS.n4115 VSS 0.0530834
R6112 VSS.n5183 VSS 0.0530834
R6113 VSS.n4249 VSS 0.0530834
R6114 VSS.n4019 VSS 0.0530834
R6115 VSS.n3998 VSS 0.0530834
R6116 VSS.n4069 VSS 0.0530834
R6117 VSS.n4099 VSS 0.0530834
R6118 VSS.n5254 VSS 0.0530834
R6119 VSS.n3675 VSS 0.0530834
R6120 VSS.n3577 VSS 0.0530834
R6121 VSS.n3480 VSS 0.0530834
R6122 VSS.n3383 VSS 0.0530834
R6123 VSS.n5335 VSS 0.0530834
R6124 VSS.n3788 VSS 0.0530834
R6125 VSS.n7480 VSS.n306 0.0530834
R6126 VSS.n626 VSS.n625 0.0530834
R6127 VSS.n626 VSS 0.0530834
R6128 VSS.n7449 VSS.n321 0.0530834
R6129 VSS.n7201 VSS.n750 0.0530834
R6130 VSS.n750 VSS 0.0530834
R6131 VSS VSS.n321 0.0530834
R6132 VSS.n7095 VSS.n330 0.0530834
R6133 VSS.n7095 VSS 0.0530834
R6134 VSS VSS.n306 0.0530834
R6135 VSS.n526 VSS.n525 0.0530834
R6136 VSS.n526 VSS 0.0530834
R6137 VSS.n7352 VSS 0.0530834
R6138 VSS.n7605 VSS 0.0530834
R6139 VSS.n416 VSS 0.0530834
R6140 VSS VSS.n7422 0.0530834
R6141 VSS VSS.n704 0.0530834
R6142 VSS.n7253 VSS 0.0530834
R6143 VSS.n7176 VSS 0.0530834
R6144 VSS.n890 VSS 0.0530834
R6145 VSS.n908 VSS 0.0530834
R6146 VSS VSS.n724 0.0530834
R6147 VSS.n6942 VSS 0.0530834
R6148 VSS.n811 VSS 0.0530834
R6149 VSS VSS.n7031 0.0530834
R6150 VSS VSS.n855 0.0530834
R6151 VSS VSS.n7005 0.0530834
R6152 VSS VSS.n921 0.0530834
R6153 VSS.n6854 VSS 0.0530834
R6154 VSS.n256 VSS 0.0526476
R6155 VSS.n440 VSS 0.0526476
R6156 VSS.n7272 VSS 0.0526476
R6157 VSS.n162 VSS 0.0526476
R6158 VSS.n211 VSS 0.0526476
R6159 VSS.n4595 VSS 0.0525833
R6160 VSS VSS.n4331 0.0525833
R6161 VSS VSS.n4642 0.0525833
R6162 VSS VSS.n4950 0.0525833
R6163 VSS.n4974 VSS 0.0525833
R6164 VSS.n4466 VSS 0.0525833
R6165 VSS.n4903 VSS 0.0525833
R6166 VSS VSS.n5117 0.0525833
R6167 VSS.n4796 VSS 0.0525833
R6168 VSS VSS.n4216 0.0525833
R6169 VSS.n5168 VSS 0.0525833
R6170 VSS VSS.n5179 0.0525833
R6171 VSS.n4938 VSS 0.0525833
R6172 VSS VSS.n3919 0.0525833
R6173 VSS VSS.n3924 0.0525833
R6174 VSS VSS.n3929 0.0525833
R6175 VSS VSS.n5221 0.0525833
R6176 VSS VSS.n5250 0.0525833
R6177 VSS VSS.n2853 0.0525833
R6178 VSS VSS.n2849 0.0525833
R6179 VSS VSS.n2845 0.0525833
R6180 VSS VSS.n2843 0.0525833
R6181 VSS VSS.n5331 0.0525833
R6182 VSS VSS.n2857 0.0525833
R6183 VSS.n5781 VSS 0.0525833
R6184 VSS.n5749 VSS 0.0525833
R6185 VSS.n5717 VSS 0.0525833
R6186 VSS.n5683 VSS 0.0525833
R6187 VSS.n618 VSS 0.0525833
R6188 VSS.n7205 VSS 0.0525833
R6189 VSS VSS.n7446 0.0525833
R6190 VSS VSS.n328 0.0525833
R6191 VSS.n7473 VSS 0.0525833
R6192 VSS.n518 VSS 0.0525833
R6193 VSS VSS.n7344 0.0525833
R6194 VSS.n7597 VSS 0.0525833
R6195 VSS.n408 VSS 0.0525833
R6196 VSS VSS.n336 0.0525833
R6197 VSS.n7400 VSS 0.0525833
R6198 VSS VSS.n7389 0.0525833
R6199 VSS.n7426 VSS 0.0525833
R6200 VSS VSS.n737 0.0525833
R6201 VSS VSS.n735 0.0525833
R6202 VSS.n7234 VSS 0.0525833
R6203 VSS VSS.n6938 0.0525833
R6204 VSS VSS.n741 0.0525833
R6205 VSS VSS.n803 0.0525833
R6206 VSS VSS.n7011 0.0525833
R6207 VSS VSS.n868 0.0525833
R6208 VSS VSS.n6985 0.0525833
R6209 VSS VSS.n6980 0.0525833
R6210 VSS VSS.n6673 0.0525833
R6211 VSS.n7725 VSS 0.0525833
R6212 VSS.n7693 VSS 0.0525833
R6213 VSS.n7661 VSS 0.0525833
R6214 VSS.n7627 VSS 0.0525833
R6215 VSS.n7187 VSS.n742 0.0525626
R6216 VSS.n679 VSS.n333 0.0525626
R6217 VSS.n415 VSS.n402 0.0525626
R6218 VSS.n5265 VSS.n2858 0.0525626
R6219 VSS.n5253 VSS.n3911 0.0525626
R6220 VSS.n4825 VSS.n4213 0.0525626
R6221 VSS.n4803 VSS.n4790 0.0525626
R6222 VSS.n4474 VSS.n4473 0.0525626
R6223 VSS.n4335 VSS.n4334 0.0525626
R6224 VSS.n4645 VSS.n4274 0.0525626
R6225 VSS.n4954 VSS.n4953 0.0525626
R6226 VSS.n4671 VSS.n3921 0.0525626
R6227 VSS.n4034 VSS.n2854 0.0525626
R6228 VSS.n4047 VSS.n2850 0.0525626
R6229 VSS.n4060 VSS.n2846 0.0525626
R6230 VSS.n4086 VSS.n2841 0.0525626
R6231 VSS.n7201 VSS.n7200 0.0525626
R6232 VSS.n636 VSS.n330 0.0525626
R6233 VSS.n7481 VSS.n7480 0.0525626
R6234 VSS.n525 VSS.n512 0.0525626
R6235 VSS.n7117 VSS.n738 0.0525626
R6236 VSS.n7164 VSS.n733 0.0525626
R6237 VSS.n7030 VSS.n7029 0.0525626
R6238 VSS.n7015 VSS.n7014 0.0525626
R6239 VSS.n7004 VSS.n7003 0.0525626
R6240 VSS.n6989 VSS.n6988 0.0525626
R6241 VSS.n6973 VSS.n6972 0.0525626
R6242 VSS.n187 VSS.n79 0.0525625
R6243 VSS.n7658 VSS.n7657 0.0525625
R6244 VSS.n7690 VSS.n7689 0.0525625
R6245 VSS.n7722 VSS.n7721 0.0525625
R6246 VSS.n7039 VSS.n7038 0.0525625
R6247 VSS.n6941 VSS.n6928 0.0525625
R6248 VSS.n7240 VSS.n7239 0.0525625
R6249 VSS.n7382 VSS.n7381 0.0525625
R6250 VSS.n7406 VSS.n7405 0.0525625
R6251 VSS.n7421 VSS.n7420 0.0525625
R6252 VSS.n7604 VSS.n7591 0.0525625
R6253 VSS.n7351 VSS.n7350 0.0525625
R6254 VSS.n5680 VSS.n5678 0.0525625
R6255 VSS.n5714 VSS.n5713 0.0525625
R6256 VSS.n5746 VSS.n5745 0.0525625
R6257 VSS.n5778 VSS.n5777 0.0525625
R6258 VSS.n5334 VSS.n2834 0.0525625
R6259 VSS.n5214 VSS.n5213 0.0525625
R6260 VSS.n4733 VSS.n3931 0.0525625
R6261 VSS.n4691 VSS.n3926 0.0525625
R6262 VSS.n5182 VSS.n4106 0.0525625
R6263 VSS.n5165 VSS.n5164 0.0525625
R6264 VSS.n4933 VSS.n4932 0.0525625
R6265 VSS.n5120 VSS.n5107 0.0525625
R6266 VSS.n4910 VSS.n4897 0.0525625
R6267 VSS.n4980 VSS.n4979 0.0525625
R6268 VSS.n4602 VSS.n4589 0.0525625
R6269 VSS.n625 VSS.n612 0.0525625
R6270 VSS.n7450 VSS.n7449 0.0525625
R6271 VSS.n7544 VSS 0.0524238
R6272 VSS.n538 VSS 0.0524238
R6273 VSS.n358 VSS 0.0524238
R6274 VSS.n5422 VSS.n5389 0.0520625
R6275 VSS.n225 VSS.n224 0.0515417
R6276 VSS.n7570 VSS.n7568 0.0515417
R6277 VSS.n7318 VSS.n7316 0.0515417
R6278 VSS.n6470 VSS.n1143 0.0515417
R6279 VSS.n5599 VSS.n5595 0.0513775
R6280 VSS.n6631 VSS.n1038 0.0513775
R6281 VSS.n6092 VSS.n6091 0.05126
R6282 VSS.n2660 VSS.n2658 0.05126
R6283 VSS.n571 VSS.n114 0.05126
R6284 VSS.n471 VSS.n118 0.05126
R6285 VSS.n7296 VSS.n258 0.05126
R6286 VSS.n283 VSS.n281 0.05126
R6287 VSS.n125 VSS.n123 0.05126
R6288 VSS.n241 VSS.n239 0.05126
R6289 VSS.n7550 VSS.n127 0.05126
R6290 VSS.n7509 VSS.n287 0.05126
R6291 VSS.n7549 VSS.n7547 0.05126
R6292 VSS.n7550 VSS.n291 0.05126
R6293 VSS.n6358 VSS.n6354 0.05126
R6294 VSS.n1854 VSS.n1182 0.05126
R6295 VSS.n1361 VSS.n1357 0.05126
R6296 VSS.n1335 VSS.n1187 0.05126
R6297 VSS.n1331 VSS.n1327 0.05126
R6298 VSS.n1210 VSS.n1191 0.05126
R6299 VSS.n1206 VSS.n1204 0.05126
R6300 VSS.n7757 VSS.n7756 0.051025
R6301 VSS.n6624 VSS.n6623 0.050555
R6302 VSS.n966 VSS.n965 0.0505002
R6303 VSS.n5087 VSS.n5086 0.0499792
R6304 VSS.n5626 VSS.n5624 0.0494583
R6305 VSS.n2197 VSS.n2196 0.0489848
R6306 VSS.n2199 VSS.n2198 0.0489848
R6307 VSS.n7531 VSS.n7529 0.0489375
R6308 VSS.n5806 VSS 0.0487365
R6309 VSS.n1057 VSS.n1056 0.047735
R6310 VSS.n2705 VSS 0.0475
R6311 VSS.n2679 VSS 0.0475
R6312 VSS.n2632 VSS 0.0475
R6313 VSS.n2665 VSS 0.0475
R6314 VSS.n2643 VSS 0.0475
R6315 VSS.n2656 VSS 0.0475
R6316 VSS.n1650 VSS 0.0475
R6317 VSS.n1533 VSS 0.0475
R6318 VSS.n1495 VSS 0.0475
R6319 VSS.n1398 VSS 0.0475
R6320 VSS.n1612 VSS 0.0475
R6321 VSS.n1547 VSS 0.0475
R6322 VSS.n1478 VSS 0.0475
R6323 VSS.n1371 VSS 0.0475
R6324 VSS.n1863 VSS 0.0475
R6325 VSS.n0 VSS 0.0475
R6326 VSS.n6351 VSS.n6350 0.047265
R6327 VSS.n1252 VSS.n1251 0.0469125
R6328 VSS.n7539 VSS.n7537 0.0468542
R6329 VSS.n480 VSS.n479 0.046795
R6330 VSS.n5413 VSS.n5411 0.0464425
R6331 VSS.n4877 VSS.n4875 0.0463333
R6332 VSS.n6578 VSS.n6577 0.046325
R6333 VSS.n6466 VSS.n6461 0.046325
R6334 VSS.n583 VSS.n579 0.0452675
R6335 VSS.n3672 VSS.n3670 0.0447708
R6336 VSS.n984 VSS.n983 0.04468
R6337 VSS.n479 VSS 0.0445116
R6338 VSS.n579 VSS 0.0444436
R6339 VSS.n7517 VSS 0.0443757
R6340 VSS.n7304 VSS 0.0443757
R6341 VSS.n279 VSS 0.0443757
R6342 VSS.n7556 VSS 0.0443757
R6343 VSS.n237 VSS 0.0443757
R6344 VSS.n352 VSS.n351 0.0442502
R6345 VSS.n6090 VSS 0.0439131
R6346 VSS.n1205 VSS 0.0439131
R6347 VSS.n1188 VSS 0.0439131
R6348 VSS.n1328 VSS 0.0439131
R6349 VSS.n1184 VSS 0.0439131
R6350 VSS.n1358 VSS 0.0439131
R6351 VSS.n1179 VSS 0.0439131
R6352 VSS.n124 VSS 0.0439131
R6353 VSS.n286 VSS 0.0439131
R6354 VSS.n2691 VSS 0.0439131
R6355 VSS.n2631 VSS 0.0439131
R6356 VSS.n2642 VSS 0.0439131
R6357 VSS.n2653 VSS 0.0439131
R6358 VSS.n2659 VSS 0.0439131
R6359 VSS.n2663 VSS 0.0439131
R6360 VSS.n2677 VSS 0.0439131
R6361 VSS.n113 VSS 0.0439131
R6362 VSS.n117 VSS 0.0439131
R6363 VSS.n242 VSS 0.0439131
R6364 VSS.n282 VSS 0.0439131
R6365 VSS.n128 VSS 0.0439131
R6366 VSS.n240 VSS 0.0439131
R6367 VSS.n1649 VSS 0.0439131
R6368 VSS.n1531 VSS 0.0439131
R6369 VSS.n1410 VSS 0.0439131
R6370 VSS.n1844 VSS 0.0439131
R6371 VSS.n292 VSS 0.0439131
R6372 VSS.n7548 VSS 0.0439131
R6373 VSS.n1625 VSS 0.0439131
R6374 VSS.n1560 VSS 0.0439131
R6375 VSS.n1491 VSS 0.0439131
R6376 VSS.n1386 VSS 0.0439131
R6377 VSS.n6355 VSS 0.0439131
R6378 VSS.n3868 VSS.n3866 0.0437292
R6379 VSS.n3770 VSS.n3768 0.0437292
R6380 VSS.n2700 VSS 0.0437243
R6381 VSS.n7305 VSS.n7304 0.0436225
R6382 VSS.n279 VSS.n272 0.0436225
R6383 VSS.n7557 VSS.n7556 0.0436225
R6384 VSS.n237 VSS.n230 0.0436225
R6385 VSS.n5361 VSS.n5360 0.043505
R6386 VSS.n6547 VSS.n6546 0.043505
R6387 VSS.n7523 VSS.n7517 0.043035
R6388 VSS.n3564 VSS.n3562 0.042095
R6389 VSS.n6826 VSS.n6822 0.0415075
R6390 VSS.n6189 VSS.n6188 0.0415075
R6391 VSS.n6511 VSS.n6510 0.04139
R6392 VSS.n6703 VSS.n6702 0.0405675
R6393 VSS.n6091 VSS.n6089 0.0402038
R6394 VSS.n241 VSS.n163 0.0400873
R6395 VSS.n4770 VSS.n4752 0.0400833
R6396 VSS.n3531 VSS.n3530 0.0396275
R6397 VSS.n5354 VSS.n2814 0.0390417
R6398 VSS.n6551 VSS.n1123 0.0390417
R6399 VSS.n2435 VSS.n2434 0.0389306
R6400 VSS.n76 VSS.n75 0.0389306
R6401 VSS.n2662 VSS.n2655 0.0383507
R6402 VSS.n160 VSS.n159 0.038335
R6403 VSS.n162 VSS.n160 0.038221
R6404 VSS.n4325 VSS.n4324 0.0381806
R6405 VSS.n4636 VSS.n4635 0.0381806
R6406 VSS.n4639 VSS.n4209 0.0381806
R6407 VSS.n4972 VSS.n4971 0.0381806
R6408 VSS.n4592 VSS.n4591 0.0381806
R6409 VSS.n4464 VSS.n4463 0.0381806
R6410 VSS.n5113 VSS.n5112 0.0381806
R6411 VSS.n4900 VSS.n4899 0.0381806
R6412 VSS.n4793 VSS.n4792 0.0381806
R6413 VSS.n4219 VSS.n4112 0.0381806
R6414 VSS.n5173 VSS.n5172 0.0381806
R6415 VSS.n4937 VSS.n4936 0.0381806
R6416 VSS.n4947 VSS.n4946 0.0381806
R6417 VSS.n5223 VSS.n5222 0.0381806
R6418 VSS.n5231 VSS.n5230 0.0381806
R6419 VSS.n5239 VSS.n5238 0.0381806
R6420 VSS.n5247 VSS.n5246 0.0381806
R6421 VSS.n4328 VSS.n3915 0.0381806
R6422 VSS.n5325 VSS.n5324 0.0381806
R6423 VSS.n5318 VSS.n5317 0.0381806
R6424 VSS.n5309 VSS.n5308 0.0381806
R6425 VSS.n5300 VSS.n5299 0.0381806
R6426 VSS.n5291 VSS.n5290 0.0381806
R6427 VSS.n5282 VSS.n5281 0.0381806
R6428 VSS.n5328 VSS.n2379 0.0381806
R6429 VSS.n5218 VSS.n2398 0.0381806
R6430 VSS.n5176 VSS.n2417 0.0381806
R6431 VSS.n7056 VSS.n747 0.0381806
R6432 VSS.n772 VSS.n324 0.0381806
R6433 VSS.n7443 VSS.n7442 0.0381806
R6434 VSS.n7471 VSS.n7470 0.0381806
R6435 VSS.n616 VSS.n615 0.0381806
R6436 VSS.n515 VSS.n514 0.0381806
R6437 VSS.n7593 VSS.n7592 0.0381806
R6438 VSS.n7346 VSS.n7345 0.0381806
R6439 VSS.n406 VSS.n405 0.0381806
R6440 VSS.n7399 VSS.n7398 0.0381806
R6441 VSS.n7391 VSS.n7390 0.0381806
R6442 VSS.n7425 VSS.n7424 0.0381806
R6443 VSS.n7435 VSS.n7434 0.0381806
R6444 VSS.n6932 VSS.n728 0.0381806
R6445 VSS.n7233 VSS.n7232 0.0381806
R6446 VSS.n7226 VSS.n7225 0.0381806
R6447 VSS.n7217 VSS.n7216 0.0381806
R6448 VSS.n7208 VSS.n7207 0.0381806
R6449 VSS.n6982 VSS.n6981 0.0381806
R6450 VSS.n930 VSS.n929 0.0381806
R6451 VSS.n7008 VSS.n7007 0.0381806
R6452 VSS.n864 VSS.n863 0.0381806
R6453 VSS.n7034 VSS.n7033 0.0381806
R6454 VSS.n6675 VSS.n6674 0.0381806
R6455 VSS.n6977 VSS.n22 0.0381806
R6456 VSS.n6935 VSS.n41 0.0381806
R6457 VSS.n7386 VSS.n60 0.0381806
R6458 VSS.n1319 VSS.n1318 0.0381
R6459 VSS.n3370 VSS.n3368 0.0379825
R6460 VSS.n6435 VSS.n6434 0.037395
R6461 VSS.n3434 VSS.n3433 0.0370425
R6462 VSS.n6126 VSS.n6121 0.0370425
R6463 VSS.n6060 VSS.n6059 0.0370425
R6464 VSS.n6359 VSS.n1178 0.0368605
R6465 VSS.n6392 VSS.n6391 0.03669
R6466 VSS.n3628 VSS.n3627 0.0365725
R6467 VSS.n3467 VSS.n3465 0.0361025
R6468 VSS.n3885 VSS.n2861 0.0356744
R6469 VSS.n4314 VSS.n4307 0.0356744
R6470 VSS.n4353 VSS.n4279 0.0356744
R6471 VSS.n2556 VSS.n2538 0.0356744
R6472 VSS.n2522 VSS.n2520 0.0356744
R6473 VSS.n6678 VSS.n6662 0.0356744
R6474 VSS.n7053 VSS.n784 0.0356744
R6475 VSS.n775 VSS.n762 0.0356744
R6476 VSS.n5474 VSS.n5473 0.0351625
R6477 VSS.n5278 VSS.n2861 0.035093
R6478 VSS.n4321 VSS.n4307 0.035093
R6479 VSS.n4632 VSS.n4279 0.035093
R6480 VSS.n2595 VSS.n2538 0.035093
R6481 VSS.n2617 VSS.n2520 0.035093
R6482 VSS.n6670 VSS.n6662 0.035093
R6483 VSS.n7059 VSS.n784 0.035093
R6484 VSS.n769 VSS.n762 0.035093
R6485 VSS.n1132 VSS.n1131 0.0348752
R6486 VSS VSS.n2168 0.0343542
R6487 VSS VSS.n6301 0.0343542
R6488 VSS.n4452 VSS.n4414 0.0341111
R6489 VSS.n2861 VSS.n2860 0.0341111
R6490 VSS.n4307 VSS.n4306 0.0341111
R6491 VSS.n4329 VSS.n4305 0.0341111
R6492 VSS.n4279 VSS.n4278 0.0341111
R6493 VSS.n4640 VSS.n4276 0.0341111
R6494 VSS.n4211 VSS.n4208 0.0341111
R6495 VSS.n4977 VSS.n4976 0.0341111
R6496 VSS.n4600 VSS.n4599 0.0341111
R6497 VSS.n4471 VSS.n4470 0.0341111
R6498 VSS.n5116 VSS.n5111 0.0341111
R6499 VSS.n4908 VSS.n4907 0.0341111
R6500 VSS.n4801 VSS.n4800 0.0341111
R6501 VSS.n5178 VSS.n4109 0.0341111
R6502 VSS.n4111 VSS.n4110 0.0341111
R6503 VSS.n4223 VSS.n4222 0.0341111
R6504 VSS.n4942 VSS.n4941 0.0341111
R6505 VSS.n5220 VSS.n5216 0.0341111
R6506 VSS.n5227 VSS.n5226 0.0341111
R6507 VSS.n5235 VSS.n5234 0.0341111
R6508 VSS.n5243 VSS.n5242 0.0341111
R6509 VSS.n3917 VSS.n3914 0.0341111
R6510 VSS.n5330 VSS.n2837 0.0341111
R6511 VSS.n5322 VSS.n2838 0.0341111
R6512 VSS.n5313 VSS.n2844 0.0341111
R6513 VSS.n5304 VSS.n2848 0.0341111
R6514 VSS.n5295 VSS.n2852 0.0341111
R6515 VSS.n5286 VSS.n2856 0.0341111
R6516 VSS.n2378 VSS.n2377 0.0341111
R6517 VSS.n2397 VSS.n2396 0.0341111
R6518 VSS.n2416 VSS.n2415 0.0341111
R6519 VSS.n2433 VSS.n2432 0.0341111
R6520 VSS.n2539 VSS.n2538 0.0341111
R6521 VSS.n2520 VSS.n2519 0.0341111
R6522 VSS.n6676 VSS.n6662 0.0341111
R6523 VSS.n7055 VSS.n784 0.0341111
R6524 VSS.n746 VSS.n744 0.0341111
R6525 VSS.n773 VSS.n762 0.0341111
R6526 VSS.n7444 VSS.n323 0.0341111
R6527 VSS.n7439 VSS.n7438 0.0341111
R6528 VSS.n7465 VSS.n308 0.0341111
R6529 VSS.n7478 VSS.n7477 0.0341111
R6530 VSS.n623 VSS.n622 0.0341111
R6531 VSS.n523 VSS.n522 0.0341111
R6532 VSS.n7342 VSS.n7341 0.0341111
R6533 VSS.n413 VSS.n412 0.0341111
R6534 VSS.n7388 VSS.n7384 0.0341111
R6535 VSS.n7403 VSS.n7402 0.0341111
R6536 VSS.n7396 VSS.n7393 0.0341111
R6537 VSS.n7430 VSS.n7429 0.0341111
R6538 VSS.n6937 VSS.n6931 0.0341111
R6539 VSS.n7237 VSS.n7236 0.0341111
R6540 VSS.n7230 VSS.n730 0.0341111
R6541 VSS.n7221 VSS.n736 0.0341111
R6542 VSS.n7212 VSS.n740 0.0341111
R6543 VSS.n6979 VSS.n6975 0.0341111
R6544 VSS.n932 VSS.n923 0.0341111
R6545 VSS.n925 VSS.n924 0.0341111
R6546 VSS.n866 VSS.n857 0.0341111
R6547 VSS.n859 VSS.n858 0.0341111
R6548 VSS.n7036 VSS.n7035 0.0341111
R6549 VSS.n21 VSS.n20 0.0341111
R6550 VSS.n40 VSS.n39 0.0341111
R6551 VSS.n59 VSS.n58 0.0341111
R6552 VSS.n3337 VSS.n3336 0.034105
R6553 VSS.n4462 VSS.n4414 0.0335556
R6554 VSS.n5280 VSS.n2861 0.0335556
R6555 VSS.n4323 VSS.n4307 0.0335556
R6556 VSS.n4326 VSS.n4305 0.0335556
R6557 VSS.n4634 VSS.n4279 0.0335556
R6558 VSS.n4637 VSS.n4276 0.0335556
R6559 VSS.n4949 VSS.n4208 0.0335556
R6560 VSS.n4977 VSS.n4970 0.0335556
R6561 VSS.n4600 VSS.n4597 0.0335556
R6562 VSS.n4471 VSS.n4468 0.0335556
R6563 VSS.n5111 VSS.n5110 0.0335556
R6564 VSS.n4908 VSS.n4905 0.0335556
R6565 VSS.n4801 VSS.n4798 0.0335556
R6566 VSS.n5175 VSS.n4109 0.0335556
R6567 VSS.n5171 VSS.n4111 0.0335556
R6568 VSS.n4223 VSS.n4218 0.0335556
R6569 VSS.n4942 VSS.n4214 0.0335556
R6570 VSS.n5217 VSS.n5216 0.0335556
R6571 VSS.n5227 VSS.n3932 0.0335556
R6572 VSS.n5235 VSS.n3927 0.0335556
R6573 VSS.n5243 VSS.n3922 0.0335556
R6574 VSS.n5249 VSS.n3914 0.0335556
R6575 VSS.n5327 VSS.n2837 0.0335556
R6576 VSS.n5323 VSS.n5322 0.0335556
R6577 VSS.n5316 VSS.n5313 0.0335556
R6578 VSS.n5307 VSS.n5304 0.0335556
R6579 VSS.n5298 VSS.n5295 0.0335556
R6580 VSS.n5289 VSS.n5286 0.0335556
R6581 VSS.n5784 VSS.n2378 0.0335556
R6582 VSS.n5752 VSS.n2397 0.0335556
R6583 VSS.n5720 VSS.n2416 0.0335556
R6584 VSS.n5685 VSS.n2433 0.0335556
R6585 VSS.n2593 VSS.n2538 0.0335556
R6586 VSS.n2619 VSS.n2520 0.0335556
R6587 VSS.n6672 VSS.n6662 0.0335556
R6588 VSS.n7057 VSS.n784 0.0335556
R6589 VSS.n7206 VSS.n746 0.0335556
R6590 VSS.n771 VSS.n762 0.0335556
R6591 VSS.n325 VSS.n323 0.0335556
R6592 VSS.n7439 VSS.n331 0.0335556
R6593 VSS.n7469 VSS.n308 0.0335556
R6594 VSS.n623 VSS.n620 0.0335556
R6595 VSS.n523 VSS.n520 0.0335556
R6596 VSS.n7602 VSS.n7601 0.0335556
R6597 VSS.n7343 VSS.n7342 0.0335556
R6598 VSS.n413 VSS.n410 0.0335556
R6599 VSS.n7385 VSS.n7384 0.0335556
R6600 VSS.n7403 VSS.n707 0.0335556
R6601 VSS.n7397 VSS.n7396 0.0335556
R6602 VSS.n7430 VSS.n334 0.0335556
R6603 VSS.n6934 VSS.n6931 0.0335556
R6604 VSS.n7237 VSS.n727 0.0335556
R6605 VSS.n7231 VSS.n7230 0.0335556
R6606 VSS.n7224 VSS.n7221 0.0335556
R6607 VSS.n7215 VSS.n7212 0.0335556
R6608 VSS.n6976 VSS.n6975 0.0335556
R6609 VSS.n6984 VSS.n923 0.0335556
R6610 VSS.n928 VSS.n925 0.0335556
R6611 VSS.n7010 VSS.n857 0.0335556
R6612 VSS.n862 VSS.n859 0.0335556
R6613 VSS.n7036 VSS.n799 0.0335556
R6614 VSS.n7728 VSS.n21 0.0335556
R6615 VSS.n7696 VSS.n40 0.0335556
R6616 VSS.n7664 VSS.n59 0.0335556
R6617 VSS.n7629 VSS.n74 0.0335556
R6618 VSS.n2245 VSS 0.0330521
R6619 VSS VSS.n2355 0.0330521
R6620 VSS VSS.n2182 0.0330521
R6621 VSS VSS.n6306 0.0330521
R6622 VSS.n3572 VSS.n2893 0.0327917
R6623 VSS.n3858 VSS.n3854 0.032695
R6624 VSS.n3760 VSS.n3757 0.032695
R6625 VSS.n3662 VSS.n3659 0.03246
R6626 VSS.n3320 VSS.n3319 0.0322708
R6627 VSS.n6351 VSS.n6343 0.031755
R6628 VSS.n4596 VSS 0.03175
R6629 VSS VSS.n4593 0.03175
R6630 VSS VSS.n4594 0.03175
R6631 VSS.n4594 VSS 0.03175
R6632 VSS.n4327 VSS 0.03175
R6633 VSS VSS.n4294 0.03175
R6634 VSS.n4332 VSS 0.03175
R6635 VSS.n4332 VSS 0.03175
R6636 VSS.n4638 VSS 0.03175
R6637 VSS VSS.n4277 0.03175
R6638 VSS.n4643 VSS 0.03175
R6639 VSS.n4643 VSS 0.03175
R6640 VSS.n4948 VSS 0.03175
R6641 VSS VSS.n4205 0.03175
R6642 VSS.n4951 VSS 0.03175
R6643 VSS.n4951 VSS 0.03175
R6644 VSS VSS.n4192 0.03175
R6645 VSS VSS.n4973 0.03175
R6646 VSS.n4973 VSS 0.03175
R6647 VSS.n4975 VSS 0.03175
R6648 VSS.n4467 VSS 0.03175
R6649 VSS VSS.n4403 0.03175
R6650 VSS VSS.n4465 0.03175
R6651 VSS.n4465 VSS 0.03175
R6652 VSS.n4904 VSS 0.03175
R6653 VSS VSS.n4901 0.03175
R6654 VSS VSS.n4902 0.03175
R6655 VSS.n4902 VSS 0.03175
R6656 VSS VSS.n5114 0.03175
R6657 VSS.n5118 VSS 0.03175
R6658 VSS.n5118 VSS 0.03175
R6659 VSS.n5115 VSS 0.03175
R6660 VSS.n4797 VSS 0.03175
R6661 VSS VSS.n4794 0.03175
R6662 VSS VSS.n4795 0.03175
R6663 VSS.n4795 VSS 0.03175
R6664 VSS.n4221 VSS 0.03175
R6665 VSS VSS.n4217 0.03175
R6666 VSS VSS.n4935 0.03175
R6667 VSS.n4935 VSS 0.03175
R6668 VSS.n5170 VSS 0.03175
R6669 VSS VSS.n4113 0.03175
R6670 VSS VSS.n5167 0.03175
R6671 VSS.n5167 VSS 0.03175
R6672 VSS.n5180 VSS 0.03175
R6673 VSS VSS.n4108 0.03175
R6674 VSS.n4108 VSS 0.03175
R6675 VSS.n5177 VSS 0.03175
R6676 VSS.n4939 VSS 0.03175
R6677 VSS.n4212 VSS 0.03175
R6678 VSS.n4944 VSS 0.03175
R6679 VSS.n4944 VSS 0.03175
R6680 VSS.n5241 VSS 0.03175
R6681 VSS VSS.n3920 0.03175
R6682 VSS VSS.n5245 0.03175
R6683 VSS.n5245 VSS 0.03175
R6684 VSS.n5232 VSS 0.03175
R6685 VSS VSS.n3925 0.03175
R6686 VSS VSS.n5237 0.03175
R6687 VSS.n5237 VSS 0.03175
R6688 VSS.n5224 VSS 0.03175
R6689 VSS VSS.n3930 0.03175
R6690 VSS VSS.n5229 0.03175
R6691 VSS.n5229 VSS 0.03175
R6692 VSS VSS.n3934 0.03175
R6693 VSS VSS.n3935 0.03175
R6694 VSS VSS.n3935 0.03175
R6695 VSS.n5219 VSS 0.03175
R6696 VSS.n5248 VSS 0.03175
R6697 VSS VSS.n3913 0.03175
R6698 VSS.n5251 VSS 0.03175
R6699 VSS.n5251 VSS 0.03175
R6700 VSS.n5297 VSS 0.03175
R6701 VSS VSS.n2855 0.03175
R6702 VSS.n5293 VSS 0.03175
R6703 VSS.n5293 VSS 0.03175
R6704 VSS.n5306 VSS 0.03175
R6705 VSS VSS.n2851 0.03175
R6706 VSS.n5302 VSS 0.03175
R6707 VSS.n5302 VSS 0.03175
R6708 VSS.n5315 VSS 0.03175
R6709 VSS VSS.n2847 0.03175
R6710 VSS.n5311 VSS 0.03175
R6711 VSS.n5311 VSS 0.03175
R6712 VSS.n2839 VSS 0.03175
R6713 VSS VSS.n2842 0.03175
R6714 VSS.n5320 VSS 0.03175
R6715 VSS.n5320 VSS 0.03175
R6716 VSS.n5332 VSS 0.03175
R6717 VSS VSS.n2836 0.03175
R6718 VSS.n2836 VSS 0.03175
R6719 VSS.n5329 VSS 0.03175
R6720 VSS.n5288 VSS 0.03175
R6721 VSS VSS.n2859 0.03175
R6722 VSS.n5284 VSS 0.03175
R6723 VSS.n5284 VSS 0.03175
R6724 VSS.n5783 VSS 0.03175
R6725 VSS VSS.n2380 0.03175
R6726 VSS VSS.n5780 0.03175
R6727 VSS.n5780 VSS 0.03175
R6728 VSS.n5751 VSS 0.03175
R6729 VSS VSS.n2399 0.03175
R6730 VSS VSS.n5748 0.03175
R6731 VSS.n5748 VSS 0.03175
R6732 VSS.n5719 VSS 0.03175
R6733 VSS VSS.n2418 0.03175
R6734 VSS VSS.n5716 0.03175
R6735 VSS.n5716 VSS 0.03175
R6736 VSS.n5684 VSS 0.03175
R6737 VSS VSS.n2436 0.03175
R6738 VSS VSS.n5682 0.03175
R6739 VSS.n5682 VSS 0.03175
R6740 VSS.n619 VSS 0.03175
R6741 VSS VSS.n617 0.03175
R6742 VSS VSS.n614 0.03175
R6743 VSS.n614 VSS 0.03175
R6744 VSS.n745 VSS 0.03175
R6745 VSS VSS.n748 0.03175
R6746 VSS VSS.n7203 0.03175
R6747 VSS.n7203 VSS 0.03175
R6748 VSS.n326 VSS 0.03175
R6749 VSS VSS.n320 0.03175
R6750 VSS.n7447 VSS 0.03175
R6751 VSS.n7447 VSS 0.03175
R6752 VSS.n7437 VSS 0.03175
R6753 VSS VSS.n329 0.03175
R6754 VSS VSS.n7441 0.03175
R6755 VSS.n7441 VSS 0.03175
R6756 VSS.n7476 VSS 0.03175
R6757 VSS VSS.n305 0.03175
R6758 VSS VSS.n7472 0.03175
R6759 VSS.n7472 VSS 0.03175
R6760 VSS.n519 VSS 0.03175
R6761 VSS VSS.n516 0.03175
R6762 VSS VSS.n517 0.03175
R6763 VSS.n517 VSS 0.03175
R6764 VSS.n7339 VSS 0.03175
R6765 VSS.n7349 VSS 0.03175
R6766 VSS.n7347 VSS 0.03175
R6767 VSS.n7347 VSS 0.03175
R6768 VSS VSS.n7594 0.03175
R6769 VSS VSS.n7596 0.03175
R6770 VSS.n7596 VSS 0.03175
R6771 VSS.n7599 VSS 0.03175
R6772 VSS.n409 VSS 0.03175
R6773 VSS VSS.n407 0.03175
R6774 VSS VSS.n404 0.03175
R6775 VSS.n404 VSS 0.03175
R6776 VSS.n7394 VSS 0.03175
R6777 VSS VSS.n337 0.03175
R6778 VSS VSS.n7423 0.03175
R6779 VSS.n7423 VSS 0.03175
R6780 VSS.n7392 VSS 0.03175
R6781 VSS VSS.n703 0.03175
R6782 VSS VSS.n706 0.03175
R6783 VSS.n706 VSS 0.03175
R6784 VSS VSS.n709 0.03175
R6785 VSS VSS.n710 0.03175
R6786 VSS VSS.n710 0.03175
R6787 VSS.n7387 VSS 0.03175
R6788 VSS.n7427 VSS 0.03175
R6789 VSS.n332 VSS 0.03175
R6790 VSS.n7432 VSS 0.03175
R6791 VSS.n7432 VSS 0.03175
R6792 VSS.n7223 VSS 0.03175
R6793 VSS VSS.n739 0.03175
R6794 VSS.n7219 VSS 0.03175
R6795 VSS.n7219 VSS 0.03175
R6796 VSS.n731 VSS 0.03175
R6797 VSS VSS.n734 0.03175
R6798 VSS.n7228 VSS 0.03175
R6799 VSS.n7228 VSS 0.03175
R6800 VSS.n729 VSS 0.03175
R6801 VSS VSS.n723 0.03175
R6802 VSS VSS.n726 0.03175
R6803 VSS.n726 VSS 0.03175
R6804 VSS.n6939 VSS 0.03175
R6805 VSS VSS.n6930 0.03175
R6806 VSS.n6930 VSS 0.03175
R6807 VSS.n6936 VSS 0.03175
R6808 VSS.n7214 VSS 0.03175
R6809 VSS VSS.n743 0.03175
R6810 VSS.n7210 VSS 0.03175
R6811 VSS.n7210 VSS 0.03175
R6812 VSS.n861 VSS 0.03175
R6813 VSS VSS.n804 0.03175
R6814 VSS VSS.n7032 0.03175
R6815 VSS.n7032 VSS 0.03175
R6816 VSS.n7009 VSS 0.03175
R6817 VSS VSS.n854 0.03175
R6818 VSS.n7012 VSS 0.03175
R6819 VSS.n7012 VSS 0.03175
R6820 VSS.n927 VSS 0.03175
R6821 VSS VSS.n869 0.03175
R6822 VSS VSS.n7006 0.03175
R6823 VSS.n7006 VSS 0.03175
R6824 VSS.n6983 VSS 0.03175
R6825 VSS VSS.n920 0.03175
R6826 VSS.n6986 VSS 0.03175
R6827 VSS.n6986 VSS 0.03175
R6828 VSS VSS.n934 0.03175
R6829 VSS VSS.n935 0.03175
R6830 VSS VSS.n935 0.03175
R6831 VSS.n6978 VSS 0.03175
R6832 VSS.n800 VSS 0.03175
R6833 VSS VSS.n795 0.03175
R6834 VSS VSS.n798 0.03175
R6835 VSS.n798 VSS 0.03175
R6836 VSS.n7727 VSS 0.03175
R6837 VSS VSS.n23 0.03175
R6838 VSS VSS.n7724 0.03175
R6839 VSS.n7724 VSS 0.03175
R6840 VSS.n7695 VSS 0.03175
R6841 VSS VSS.n42 0.03175
R6842 VSS VSS.n7692 0.03175
R6843 VSS.n7692 VSS 0.03175
R6844 VSS.n7663 VSS 0.03175
R6845 VSS VSS.n61 0.03175
R6846 VSS VSS.n7660 0.03175
R6847 VSS.n7660 VSS 0.03175
R6848 VSS.n7628 VSS 0.03175
R6849 VSS VSS.n77 0.03175
R6850 VSS VSS.n7624 0.03175
R6851 VSS.n7624 VSS 0.03175
R6852 VSS.n4334 VSS.n4304 0.0316203
R6853 VSS.n4334 VSS.n4333 0.0316203
R6854 VSS.n4645 VSS.n4275 0.0316203
R6855 VSS.n4645 VSS.n4644 0.0316203
R6856 VSS.n4953 VSS.n4207 0.0316203
R6857 VSS.n4953 VSS.n4952 0.0316203
R6858 VSS.n4979 VSS.n4968 0.0316203
R6859 VSS.n4979 VSS.n4978 0.0316203
R6860 VSS.n4602 VSS.n4590 0.0316203
R6861 VSS.n4602 VSS.n4601 0.0316203
R6862 VSS.n4473 VSS.n4413 0.0316203
R6863 VSS.n4473 VSS.n4472 0.0316203
R6864 VSS.n5120 VSS.n5108 0.0316203
R6865 VSS.n5120 VSS.n5119 0.0316203
R6866 VSS.n4910 VSS.n4898 0.0316203
R6867 VSS.n4910 VSS.n4909 0.0316203
R6868 VSS.n4803 VSS.n4791 0.0316203
R6869 VSS.n4803 VSS.n4802 0.0316203
R6870 VSS.n5182 VSS.n4107 0.0316203
R6871 VSS.n5182 VSS.n5181 0.0316203
R6872 VSS.n5165 VSS.n4114 0.0316203
R6873 VSS.n5166 VSS.n5165 0.0316203
R6874 VSS.n4933 VSS.n4215 0.0316203
R6875 VSS.n4933 VSS.n4224 0.0316203
R6876 VSS.n4945 VSS.n4213 0.0316203
R6877 VSS.n4943 VSS.n4213 0.0316203
R6878 VSS.n5214 VSS.n3933 0.0316203
R6879 VSS.n5215 VSS.n5214 0.0316203
R6880 VSS.n3931 VSS.n3928 0.0316203
R6881 VSS.n5228 VSS.n3931 0.0316203
R6882 VSS.n3926 VSS.n3923 0.0316203
R6883 VSS.n5236 VSS.n3926 0.0316203
R6884 VSS.n3921 VSS.n3918 0.0316203
R6885 VSS.n5244 VSS.n3921 0.0316203
R6886 VSS.n5253 VSS.n3912 0.0316203
R6887 VSS.n5253 VSS.n5252 0.0316203
R6888 VSS.n5334 VSS.n2835 0.0316203
R6889 VSS.n5334 VSS.n5333 0.0316203
R6890 VSS.n5319 VSS.n2841 0.0316203
R6891 VSS.n5321 VSS.n2841 0.0316203
R6892 VSS.n5310 VSS.n2846 0.0316203
R6893 VSS.n5312 VSS.n2846 0.0316203
R6894 VSS.n5301 VSS.n2850 0.0316203
R6895 VSS.n5303 VSS.n2850 0.0316203
R6896 VSS.n5292 VSS.n2854 0.0316203
R6897 VSS.n5294 VSS.n2854 0.0316203
R6898 VSS.n5283 VSS.n2858 0.0316203
R6899 VSS.n5285 VSS.n2858 0.0316203
R6900 VSS.n5778 VSS.n2381 0.0316203
R6901 VSS.n5779 VSS.n5778 0.0316203
R6902 VSS.n5746 VSS.n2400 0.0316203
R6903 VSS.n5747 VSS.n5746 0.0316203
R6904 VSS.n5714 VSS.n2419 0.0316203
R6905 VSS.n5715 VSS.n5714 0.0316203
R6906 VSS.n5680 VSS.n5679 0.0316203
R6907 VSS.n5681 VSS.n5680 0.0316203
R6908 VSS.n7201 VSS.n749 0.0316203
R6909 VSS.n7202 VSS.n7201 0.0316203
R6910 VSS.n7449 VSS.n322 0.0316203
R6911 VSS.n7449 VSS.n7448 0.0316203
R6912 VSS.n330 VSS.n327 0.0316203
R6913 VSS.n7440 VSS.n330 0.0316203
R6914 VSS.n7480 VSS.n307 0.0316203
R6915 VSS.n7480 VSS.n7479 0.0316203
R6916 VSS.n625 VSS.n613 0.0316203
R6917 VSS.n625 VSS.n624 0.0316203
R6918 VSS.n525 VSS.n513 0.0316203
R6919 VSS.n525 VSS.n524 0.0316203
R6920 VSS.n7604 VSS.n7603 0.0316203
R6921 VSS.n415 VSS.n403 0.0316203
R6922 VSS.n415 VSS.n414 0.0316203
R6923 VSS.n7382 VSS.n708 0.0316203
R6924 VSS.n7383 VSS.n7382 0.0316203
R6925 VSS.n7405 VSS.n705 0.0316203
R6926 VSS.n7405 VSS.n7404 0.0316203
R6927 VSS.n7421 VSS.n335 0.0316203
R6928 VSS.n7421 VSS.n338 0.0316203
R6929 VSS.n7433 VSS.n333 0.0316203
R6930 VSS.n7431 VSS.n333 0.0316203
R6931 VSS.n6941 VSS.n6929 0.0316203
R6932 VSS.n6941 VSS.n6940 0.0316203
R6933 VSS.n7239 VSS.n725 0.0316203
R6934 VSS.n7239 VSS.n7238 0.0316203
R6935 VSS.n7227 VSS.n733 0.0316203
R6936 VSS.n7229 VSS.n733 0.0316203
R6937 VSS.n7218 VSS.n738 0.0316203
R6938 VSS.n7220 VSS.n738 0.0316203
R6939 VSS.n7209 VSS.n742 0.0316203
R6940 VSS.n7211 VSS.n742 0.0316203
R6941 VSS.n6973 VSS.n933 0.0316203
R6942 VSS.n6974 VSS.n6973 0.0316203
R6943 VSS.n6988 VSS.n922 0.0316203
R6944 VSS.n6988 VSS.n6987 0.0316203
R6945 VSS.n7004 VSS.n867 0.0316203
R6946 VSS.n7004 VSS.n870 0.0316203
R6947 VSS.n7014 VSS.n856 0.0316203
R6948 VSS.n7014 VSS.n7013 0.0316203
R6949 VSS.n7030 VSS.n802 0.0316203
R6950 VSS.n7030 VSS.n805 0.0316203
R6951 VSS.n7038 VSS.n797 0.0316203
R6952 VSS.n7038 VSS.n7037 0.0316203
R6953 VSS.n7722 VSS.n24 0.0316203
R6954 VSS.n7723 VSS.n7722 0.0316203
R6955 VSS.n7690 VSS.n43 0.0316203
R6956 VSS.n7691 VSS.n7690 0.0316203
R6957 VSS.n7658 VSS.n62 0.0316203
R6958 VSS.n7659 VSS.n7658 0.0316203
R6959 VSS.n79 VSS.n78 0.0316203
R6960 VSS.n359 VSS.n358 0.0314025
R6961 VSS.n2471 VSS.n2453 0.0307083
R6962 VSS.n6834 VSS.n957 0.0307083
R6963 VSS.n6178 VSS.n6103 0.0307083
R6964 VSS.n1206 VSS.n1196 0.0303642
R6965 VSS.n537 VSS.n287 0.0303642
R6966 VSS.n439 VSS.n114 0.0303642
R6967 VSS.n7271 VSS.n283 0.0303642
R6968 VSS.n357 VSS.n118 0.0303642
R6969 VSS.n258 VSS.n257 0.0303642
R6970 VSS.n210 VSS.n125 0.0303642
R6971 VSS.n7549 VSS.n7545 0.0303642
R6972 VSS.n6358 VSS.n6357 0.0303642
R6973 VSS.n1182 VSS.n1181 0.0303642
R6974 VSS.n1361 VSS.n1360 0.0303642
R6975 VSS.n1187 VSS.n1186 0.0303642
R6976 VSS.n1331 VSS.n1330 0.0303642
R6977 VSS.n1191 VSS.n1190 0.0303642
R6978 VSS.n6359 VSS.n1194 0.0303642
R6979 VSS.n2441 VSS.n2440 0.0286252
R6980 VSS.n3477 VSS.n3475 0.028625
R6981 VSS.n3823 VSS.n3822 0.0283475
R6982 VSS.n3726 VSS.n3725 0.0283475
R6983 VSS.n2286 VSS 0.0278438
R6984 VSS.n2314 VSS 0.0278438
R6985 VSS.n2342 VSS 0.0278438
R6986 VSS.n5785 VSS.n2375 0.0278438
R6987 VSS.n5753 VSS.n2394 0.0278438
R6988 VSS.n5721 VSS.n2413 0.0278438
R6989 VSS.n5687 VSS.n5686 0.0278438
R6990 VSS.n2592 VSS.n2540 0.0278438
R6991 VSS.n2620 VSS.n2518 0.0278438
R6992 VSS.n7729 VSS.n18 0.0278438
R6993 VSS.n7697 VSS.n37 0.0278438
R6994 VSS.n7665 VSS.n56 0.0278438
R6995 VSS.n7631 VSS.n7630 0.0278438
R6996 VSS.n5457 VSS.n5456 0.0275833
R6997 VSS.n3524 VSS.n3523 0.0270627
R6998 VSS.n6698 VSS.n6661 0.0265417
R6999 VSS.n2743 VSS.n2722 0.0265417
R7000 VSS.n6398 VSS.n6396 0.0260208
R7001 VSS.n1458 VSS.n1384 0.02588
R7002 VSS.n1585 VSS.n1562 0.02588
R7003 VSS.n1733 VSS.n1611 0.02588
R7004 VSS.n7550 VSS.n112 0.02588
R7005 VSS.n7550 VSS.n284 0.02588
R7006 VSS.n7550 VSS.n116 0.02588
R7007 VSS.n7550 VSS.n120 0.02588
R7008 VSS.n1705 VSS.n1634 0.02588
R7009 VSS.n7552 VSS.n7550 0.02588
R7010 VSS.n7550 VSS.n122 0.02588
R7011 VSS.n1732 VSS.n1730 0.02588
R7012 VSS.n1733 VSS.n1629 0.02588
R7013 VSS.n1776 VSS.n1532 0.02588
R7014 VSS.n1776 VSS.n1546 0.02588
R7015 VSS.n1605 VSS.n1577 0.02588
R7016 VSS.n1775 VSS.n1773 0.02588
R7017 VSS.n1776 VSS.n1564 0.02588
R7018 VSS.n1776 VSS.n1568 0.02588
R7019 VSS.n1845 VSS.n1477 0.02588
R7020 VSS.n1853 VSS.n1362 0.02588
R7021 VSS.n1470 VSS.n1397 0.02588
R7022 VSS.n1845 VSS.n1843 0.02588
R7023 VSS.n1526 VSS.n1506 0.02588
R7024 VSS.n1758 VSS.n1544 0.02588
R7025 VSS.n1747 VSS.n1573 0.02588
R7026 VSS.n1715 VSS.n1647 0.02588
R7027 VSS.n1685 VSS.n1639 0.02588
R7028 VSS.n1733 VSS.n1645 0.02588
R7029 VSS.n1733 VSS.n1641 0.02588
R7030 VSS.n1695 VSS.n1637 0.02588
R7031 VSS.n1733 VSS.n1630 0.02588
R7032 VSS.n1733 VSS.n1632 0.02588
R7033 VSS.n1735 VSS.n1570 0.02588
R7034 VSS.n1776 VSS.n1578 0.02588
R7035 VSS.n1776 VSS.n1574 0.02588
R7036 VSS.n1817 VSS.n1511 0.02588
R7037 VSS.n1830 VSS.n1508 0.02588
R7038 VSS.n1845 VSS.n1524 0.02588
R7039 VSS.n1845 VSS.n1512 0.02588
R7040 VSS.n1853 VSS.n1394 0.02588
R7041 VSS.n1420 VSS.n1364 0.02588
R7042 VSS.n1853 VSS.n1366 0.02588
R7043 VSS.n1427 VSS.n1393 0.02588
R7044 VSS.n1811 VSS.n1515 0.02588
R7045 VSS.n1797 VSS.n1523 0.02588
R7046 VSS.n1845 VSS.n1516 0.02588
R7047 VSS.n1845 VSS.n1520 0.02588
R7048 VSS.n1853 VSS.n1390 0.02588
R7049 VSS.n1449 VSS.n1368 0.02588
R7050 VSS.n1853 VSS.n1370 0.02588
R7051 VSS.n1439 VSS.n1389 0.02588
R7052 VSS.n1779 VSS.n1518 0.02588
R7053 VSS.n1787 VSS.n1493 0.02588
R7054 VSS.n1596 VSS.n1566 0.02588
R7055 VSS.n1664 VSS.n1644 0.02588
R7056 VSS.n1675 VSS.n1627 0.02588
R7057 VSS.n7550 VSS.n293 0.02588
R7058 VSS.n1733 VSS.n1624 0.02588
R7059 VSS.n1776 VSS.n1559 0.02588
R7060 VSS.n1845 VSS.n1490 0.02588
R7061 VSS.n1853 VSS.n1385 0.02588
R7062 VSS.n1413 VSS.n1409 0.02588
R7063 VSS.n1853 VSS.n1852 0.02588
R7064 VSS.n542 VSS.n538 0.0252925
R7065 VSS.n256 VSS.n255 0.0245875
R7066 VSS.n7273 VSS.n7272 0.0245875
R7067 VSS.n212 VSS.n211 0.0245875
R7068 VSS.n2696 VSS 0.024
R7069 VSS.n2705 VSS 0.024
R7070 VSS.n2656 VSS 0.024
R7071 VSS.n2654 VSS 0.024
R7072 VSS VSS.n289 0.024
R7073 VSS.n2347 VSS 0.0239375
R7074 VSS.n6275 VSS 0.0239375
R7075 VSS.n6287 VSS 0.0239375
R7076 VSS.n6314 VSS.n6313 0.0233646
R7077 VSS.n444 VSS.n440 0.023295
R7078 VSS.n4432 VSS.n4431 0.0228958
R7079 VSS.n4508 VSS.n4506 0.0228958
R7080 VSS.n4551 VSS.n4550 0.0228958
R7081 VSS.n5013 VSS.n5011 0.0228958
R7082 VSS.n2243 VSS 0.0226354
R7083 VSS.n2136 VSS 0.0226354
R7084 VSS.n6269 VSS 0.0226354
R7085 VSS.n1383 VSS 0.0224565
R7086 VSS.n1382 VSS 0.0224565
R7087 VSS.n1561 VSS 0.0224565
R7088 VSS.n1558 VSS 0.0224565
R7089 VSS.n1643 VSS 0.0224565
R7090 VSS.n1628 VSS 0.0224565
R7091 VSS.n1636 VSS 0.0224565
R7092 VSS.n1631 VSS 0.0224565
R7093 VSS.n294 VSS 0.0224565
R7094 VSS.n285 VSS 0.0224565
R7095 VSS.n115 VSS 0.0224565
R7096 VSS.n259 VSS 0.0224565
R7097 VSS.n119 VSS 0.0224565
R7098 VSS.n1646 VSS 0.0224565
R7099 VSS.n1640 VSS 0.0224565
R7100 VSS.n1633 VSS 0.0224565
R7101 VSS.n1635 VSS 0.0224565
R7102 VSS.n121 VSS 0.0224565
R7103 VSS.n126 VSS 0.0224565
R7104 VSS.n1731 VSS 0.0224565
R7105 VSS.n1648 VSS 0.0224565
R7106 VSS.n1565 VSS 0.0224565
R7107 VSS.n1563 VSS 0.0224565
R7108 VSS.n1543 VSS 0.0224565
R7109 VSS.n1545 VSS 0.0224565
R7110 VSS.n1576 VSS 0.0224565
R7111 VSS.n1579 VSS 0.0224565
R7112 VSS.n1774 VSS 0.0224565
R7113 VSS.n1567 VSS 0.0224565
R7114 VSS.n1514 VSS 0.0224565
R7115 VSS.n1521 VSS 0.0224565
R7116 VSS.n1517 VSS 0.0224565
R7117 VSS.n1494 VSS 0.0224565
R7118 VSS.n1396 VSS 0.0224565
R7119 VSS.n1395 VSS 0.0224565
R7120 VSS.n1408 VSS 0.0224565
R7121 VSS.n1411 VSS 0.0224565
R7122 VSS.n1505 VSS 0.0224565
R7123 VSS.n1525 VSS 0.0224565
R7124 VSS.n1572 VSS 0.0224565
R7125 VSS.n1571 VSS 0.0224565
R7126 VSS.n1638 VSS 0.0224565
R7127 VSS.n1642 VSS 0.0224565
R7128 VSS.n1569 VSS 0.0224565
R7129 VSS.n1575 VSS 0.0224565
R7130 VSS.n1510 VSS 0.0224565
R7131 VSS.n1509 VSS 0.0224565
R7132 VSS.n1507 VSS 0.0224565
R7133 VSS.n1513 VSS 0.0224565
R7134 VSS.n1363 VSS 0.0224565
R7135 VSS.n1365 VSS 0.0224565
R7136 VSS.n1392 VSS 0.0224565
R7137 VSS.n1391 VSS 0.0224565
R7138 VSS.n1522 VSS 0.0224565
R7139 VSS.n1519 VSS 0.0224565
R7140 VSS.n1367 VSS 0.0224565
R7141 VSS.n1369 VSS 0.0224565
R7142 VSS.n1388 VSS 0.0224565
R7143 VSS.n1387 VSS 0.0224565
R7144 VSS.n1492 VSS 0.0224565
R7145 VSS.n1489 VSS 0.0224565
R7146 VSS.n1626 VSS 0.0224565
R7147 VSS.n1623 VSS 0.0224565
R7148 VSS.n2661 VSS.n2656 0.0220983
R7149 VSS.n162 VSS 0.0216803
R7150 VSS.n4397 VSS.n4396 0.0213335
R7151 VSS.n4379 VSS.n4378 0.0213335
R7152 VSS.n4185 VSS.n4184 0.0213335
R7153 VSS.n5037 VSS.n5036 0.0213335
R7154 VSS VSS.n83 0.0213333
R7155 VSS VSS.n6909 0.0213333
R7156 VSS VSS.n6953 0.0213333
R7157 VSS.n6160 VSS 0.0213333
R7158 VSS.n6841 VSS.n6840 0.0213333
R7159 VSS.n1292 VSS.n1291 0.0213333
R7160 VSS.n6416 VSS.n6415 0.0213333
R7161 VSS.n6502 VSS.n6501 0.0213333
R7162 VSS.n6991 VSS.n6990 0.0213333
R7163 VSS.n7002 VSS.n871 0.0213333
R7164 VSS.n7590 VSS.n7589 0.0213333
R7165 VSS.n7319 VSS.n7294 0.0213333
R7166 VSS.n7576 VSS.n7575 0.0213333
R7167 VSS.n189 VSS.n188 0.0213333
R7168 VSS.n7571 VSS.n107 0.0213333
R7169 VSS.n218 VSS.n201 0.0213333
R7170 VSS.n222 VSS.n184 0.0213333
R7171 VSS.n381 VSS.n380 0.0213333
R7172 VSS.n2246 VSS 0.0213333
R7173 VSS VSS.n5132 0.0213333
R7174 VSS VSS.n5194 0.0213333
R7175 VSS VSS.n3958 0.0213333
R7176 VSS VSS.n5439 0.0213333
R7177 VSS.n5351 VSS.n5349 0.0213333
R7178 VSS.n3413 VSS.n3411 0.0213333
R7179 VSS.n3510 VSS.n3508 0.0213333
R7180 VSS.n3607 VSS.n3605 0.0213333
R7181 VSS.n4061 VSS.n4059 0.0213333
R7182 VSS.n4769 VSS.n4768 0.0213333
R7183 VSS.n5014 VSS.n5006 0.0213333
R7184 VSS.n4775 VSS.n4774 0.0213333
R7185 VSS.n4789 VSS.n4788 0.0213333
R7186 VSS.n4826 VSS.n4824 0.0213333
R7187 VSS VSS.n4266 0.0213333
R7188 VSS.n4487 VSS.n4486 0.0213333
R7189 VSS VSS.n4456 0.0213333
R7190 VSS VSS.n4407 0.0213333
R7191 VSS VSS.n4411 0.0213333
R7192 VSS.n4548 VSS.n4547 0.0213333
R7193 VSS.n4992 VSS.n4991 0.0213333
R7194 VSS.n4982 VSS.n4981 0.0213333
R7195 VSS.n4509 VSS.n4501 0.0213333
R7196 VSS.n4574 VSS.n4573 0.0213333
R7197 VSS.n4588 VSS.n4587 0.0213333
R7198 VSS VSS.n4375 0.0213333
R7199 VSS.n4604 VSS 0.0213333
R7200 VSS.n4955 VSS.n4204 0.0213333
R7201 VSS.n4620 VSS.n4619 0.0213333
R7202 VSS VSS.n4298 0.0213333
R7203 VSS VSS.n3883 0.0213333
R7204 VSS VSS.n4302 0.0213333
R7205 VSS.n5267 VSS.n5266 0.0213333
R7206 VSS VSS.n4312 0.0213333
R7207 VSS VSS.n4351 0.0213333
R7208 VSS.n4342 VSS.n4341 0.0213333
R7209 VSS.n4341 VSS.n4340 0.0213333
R7210 VSS.n4267 VSS 0.0213333
R7211 VSS.n4660 VSS.n4659 0.0213333
R7212 VSS.n4647 VSS 0.0213333
R7213 VSS VSS.n4273 0.0213333
R7214 VSS.n4621 VSS.n4620 0.0213333
R7215 VSS.n4956 VSS.n4955 0.0213333
R7216 VSS VSS.n4193 0.0213333
R7217 VSS VSS.n4966 0.0213333
R7218 VSS.n4476 VSS.n4475 0.0213333
R7219 VSS.n4436 VSS 0.0213333
R7220 VSS.n5106 VSS.n5105 0.0213333
R7221 VSS.n4878 VSS.n4871 0.0213333
R7222 VSS.n5092 VSS.n5091 0.0213333
R7223 VSS.n5677 VSS.n5676 0.0213333
R7224 VSS.n4151 VSS.n4150 0.0213333
R7225 VSS.n5663 VSS.n5662 0.0213333
R7226 VSS.n2468 VSS.n2467 0.0213333
R7227 VSS.n4882 VSS.n4881 0.0213333
R7228 VSS.n4896 VSS.n4895 0.0213333
R7229 VSS.n5163 VSS.n4116 0.0213333
R7230 VSS.n4838 VSS 0.0213333
R7231 VSS.n4916 VSS 0.0213333
R7232 VSS VSS.n4915 0.0213333
R7233 VSS.n5151 VSS.n5150 0.0213333
R7234 VSS.n5163 VSS.n5162 0.0213333
R7235 VSS.n5150 VSS.n5149 0.0213333
R7236 VSS.n5133 VSS 0.0213333
R7237 VSS.n5712 VSS.n2421 0.0213333
R7238 VSS.n5122 VSS 0.0213333
R7239 VSS VSS.n4133 0.0213333
R7240 VSS VSS.n4837 0.0213333
R7241 VSS.n4827 VSS.n4826 0.0213333
R7242 VSS.n4931 VSS.n4745 0.0213333
R7243 VSS.n4931 VSS.n4930 0.0213333
R7244 VSS VSS.n4248 0.0213333
R7245 VSS.n4692 VSS.n4690 0.0213333
R7246 VSS VSS.n4225 0.0213333
R7247 VSS VSS.n4744 0.0213333
R7248 VSS.n4735 VSS.n4734 0.0213333
R7249 VSS.n4693 VSS.n4692 0.0213333
R7250 VSS VSS.n4709 0.0213333
R7251 VSS.n4710 VSS 0.0213333
R7252 VSS.n5212 VSS.n4100 0.0213333
R7253 VSS.n4734 VSS.n4732 0.0213333
R7254 VSS.n5212 VSS.n5211 0.0213333
R7255 VSS.n5195 VSS 0.0213333
R7256 VSS.n5744 VSS.n2402 0.0213333
R7257 VSS.n5184 VSS 0.0213333
R7258 VSS VSS.n4105 0.0213333
R7259 VSS.n4250 VSS 0.0213333
R7260 VSS.n4663 VSS.n4660 0.0213333
R7261 VSS.n4672 VSS.n4670 0.0213333
R7262 VSS.n4673 VSS.n4672 0.0213333
R7263 VSS.n4048 VSS.n4046 0.0213333
R7264 VSS VSS.n3910 0.0213333
R7265 VSS.n4024 VSS 0.0213333
R7266 VSS VSS.n4023 0.0213333
R7267 VSS.n4049 VSS.n4048 0.0213333
R7268 VSS.n4002 VSS 0.0213333
R7269 VSS VSS.n4001 0.0213333
R7270 VSS.n4087 VSS.n4085 0.0213333
R7271 VSS.n4062 VSS.n4061 0.0213333
R7272 VSS.n4074 VSS 0.0213333
R7273 VSS VSS.n4073 0.0213333
R7274 VSS.n3977 VSS.n3976 0.0213333
R7275 VSS.n4088 VSS.n4087 0.0213333
R7276 VSS.n3976 VSS.n3975 0.0213333
R7277 VSS.n3959 VSS 0.0213333
R7278 VSS.n5776 VSS.n2383 0.0213333
R7279 VSS VSS.n3937 0.0213333
R7280 VSS VSS.n4098 0.0213333
R7281 VSS.n5255 VSS 0.0213333
R7282 VSS.n5266 VSS.n5264 0.0213333
R7283 VSS.n4035 VSS.n4033 0.0213333
R7284 VSS.n4036 VSS.n4035 0.0213333
R7285 VSS.n3705 VSS.n3703 0.0213333
R7286 VSS VSS.n3787 0.0213333
R7287 VSS.n3776 VSS.n3771 0.0213333
R7288 VSS.n3690 VSS 0.0213333
R7289 VSS VSS.n3689 0.0213333
R7290 VSS.n3678 VSS.n3673 0.0213333
R7291 VSS.n3592 VSS 0.0213333
R7292 VSS VSS.n3591 0.0213333
R7293 VSS.n3580 VSS.n3575 0.0213333
R7294 VSS.n3495 VSS 0.0213333
R7295 VSS VSS.n3494 0.0213333
R7296 VSS.n3483 VSS.n3478 0.0213333
R7297 VSS.n3398 VSS 0.0213333
R7298 VSS VSS.n3397 0.0213333
R7299 VSS.n3386 VSS.n3381 0.0213333
R7300 VSS.n5353 VSS.n2816 0.0213333
R7301 VSS.n5440 VSS 0.0213333
R7302 VSS.n5453 VSS.n5451 0.0213333
R7303 VSS VSS.n2833 0.0213333
R7304 VSS.n5336 VSS 0.0213333
R7305 VSS.n3789 VSS 0.0213333
R7306 VSS.n3802 VSS.n3800 0.0213333
R7307 VSS.n3611 VSS.n3610 0.0213333
R7308 VSS.n5429 VSS.n5423 0.0213333
R7309 VSS.n5790 VSS 0.0213333
R7310 VSS.n5776 VSS.n5775 0.0213333
R7311 VSS.n5758 VSS 0.0213333
R7312 VSS.n5744 VSS.n5743 0.0213333
R7313 VSS.n5726 VSS 0.0213333
R7314 VSS.n5712 VSS.n5711 0.0213333
R7315 VSS.n5694 VSS 0.0213333
R7316 VSS VSS.n2490 0.0213333
R7317 VSS VSS.n5622 0.0213333
R7318 VSS.n2533 VSS 0.0213333
R7319 VSS.n2558 VSS 0.0213333
R7320 VSS VSS.n2587 0.0213333
R7321 VSS VSS.n2608 0.0213333
R7322 VSS.n5610 VSS 0.0213333
R7323 VSS.n494 VSS.n469 0.0213333
R7324 VSS.n387 VSS.n386 0.0213333
R7325 VSS.n401 VSS.n400 0.0213333
R7326 VSS VSS.n436 0.0213333
R7327 VSS VSS.n2737 0.0213333
R7328 VSS.n7536 VSS.n7492 0.0213333
R7329 VSS.n7096 VSS 0.0213333
R7330 VSS VSS.n7462 0.0213333
R7331 VSS.n499 VSS.n498 0.0213333
R7332 VSS.n7532 VSS.n7506 0.0213333
R7333 VSS.n597 VSS.n596 0.0213333
R7334 VSS.n611 VSS.n610 0.0213333
R7335 VSS.n637 VSS.n635 0.0213333
R7336 VSS.n527 VSS 0.0213333
R7337 VSS.n680 VSS.n678 0.0213333
R7338 VSS.n666 VSS 0.0213333
R7339 VSS VSS.n665 0.0213333
R7340 VSS.n7451 VSS.n319 0.0213333
R7341 VSS.n826 VSS 0.0213333
R7342 VSS.n6680 VSS 0.0213333
R7343 VSS VSS.n825 0.0213333
R7344 VSS.n7041 VSS.n7040 0.0213333
R7345 VSS VSS.n7051 0.0213333
R7346 VSS.n777 VSS 0.0213333
R7347 VSS.n7199 VSS.n751 0.0213333
R7348 VSS.n7199 VSS.n7198 0.0213333
R7349 VSS VSS.n7094 0.0213333
R7350 VSS.n7189 VSS.n7188 0.0213333
R7351 VSS.n7076 VSS 0.0213333
R7352 VSS VSS.n7075 0.0213333
R7353 VSS.n7452 VSS.n7451 0.0213333
R7354 VSS.n638 VSS.n637 0.0213333
R7355 VSS.n649 VSS 0.0213333
R7356 VSS VSS.n648 0.0213333
R7357 VSS.n7483 VSS.n7482 0.0213333
R7358 VSS.n511 VSS.n510 0.0213333
R7359 VSS.n592 VSS.n567 0.0213333
R7360 VSS.n7323 VSS.n7322 0.0213333
R7361 VSS.n7337 VSS.n7336 0.0213333
R7362 VSS.n7408 VSS.n7407 0.0213333
R7363 VSS.n692 VSS 0.0213333
R7364 VSS VSS.n7262 0.0213333
R7365 VSS.n7353 VSS 0.0213333
R7366 VSS.n7380 VSS.n7374 0.0213333
R7367 VSS.n7407 VSS.n702 0.0213333
R7368 VSS.n7380 VSS.n7379 0.0213333
R7369 VSS VSS.n7621 0.0213333
R7370 VSS.n7656 VSS.n64 0.0213333
R7371 VSS.n7606 VSS 0.0213333
R7372 VSS VSS.n91 0.0213333
R7373 VSS VSS.n691 0.0213333
R7374 VSS.n681 VSS.n680 0.0213333
R7375 VSS.n7419 VSS.n339 0.0213333
R7376 VSS.n7419 VSS.n7418 0.0213333
R7377 VSS VSS.n7175 0.0213333
R7378 VSS.n7166 VSS.n7165 0.0213333
R7379 VSS.n7126 VSS 0.0213333
R7380 VSS.n7136 VSS 0.0213333
R7381 VSS.n7241 VSS.n722 0.0213333
R7382 VSS.n7165 VSS.n7163 0.0213333
R7383 VSS.n7147 VSS 0.0213333
R7384 VSS VSS.n7146 0.0213333
R7385 VSS.n6927 VSS.n6895 0.0213333
R7386 VSS.n7242 VSS.n7241 0.0213333
R7387 VSS.n6927 VSS.n6926 0.0213333
R7388 VSS.n6910 VSS 0.0213333
R7389 VSS.n7688 VSS.n45 0.0213333
R7390 VSS VSS.n712 0.0213333
R7391 VSS VSS.n7252 0.0213333
R7392 VSS.n7177 VSS 0.0213333
R7393 VSS.n7188 VSS.n7186 0.0213333
R7394 VSS.n7118 VSS.n7116 0.0213333
R7395 VSS.n7119 VSS.n7118 0.0213333
R7396 VSS.n7017 VSS.n7016 0.0213333
R7397 VSS.n843 VSS 0.0213333
R7398 VSS VSS.n889 0.0213333
R7399 VSS.n891 VSS 0.0213333
R7400 VSS.n7016 VSS.n853 0.0213333
R7401 VSS VSS.n907 0.0213333
R7402 VSS.n909 VSS 0.0213333
R7403 VSS.n7002 VSS.n7001 0.0213333
R7404 VSS VSS.n6870 0.0213333
R7405 VSS.n6871 VSS 0.0213333
R7406 VSS.n6971 VSS.n6855 0.0213333
R7407 VSS.n6990 VSS.n919 0.0213333
R7408 VSS.n6971 VSS.n6970 0.0213333
R7409 VSS.n6954 VSS 0.0213333
R7410 VSS.n7720 VSS.n26 0.0213333
R7411 VSS.n6943 VSS 0.0213333
R7412 VSS VSS.n6890 0.0213333
R7413 VSS VSS.n842 0.0213333
R7414 VSS.n7040 VSS.n794 0.0213333
R7415 VSS.n7028 VSS.n806 0.0213333
R7416 VSS.n7028 VSS.n7027 0.0213333
R7417 VSS.n6569 VSS.n6568 0.0213333
R7418 VSS.n1075 VSS 0.0213333
R7419 VSS.n6638 VSS.n1087 0.0213333
R7420 VSS.n6555 VSS 0.0213333
R7421 VSS.n1109 VSS 0.0213333
R7422 VSS.n6553 VSS.n1121 0.0213333
R7423 VSS.n6488 VSS 0.0213333
R7424 VSS VSS.n6487 0.0213333
R7425 VSS.n6476 VSS.n6472 0.0213333
R7426 VSS.n6402 VSS 0.0213333
R7427 VSS.n1160 VSS 0.0213333
R7428 VSS.n6400 VSS.n1172 0.0213333
R7429 VSS.n1278 VSS 0.0213333
R7430 VSS VSS.n1277 0.0213333
R7431 VSS.n1266 VSS.n1262 0.0213333
R7432 VSS.n6838 VSS.n955 0.0213333
R7433 VSS VSS.n6159 0.0213333
R7434 VSS.n6149 VSS.n6143 0.0213333
R7435 VSS VSS.n937 0.0213333
R7436 VSS VSS.n6853 0.0213333
R7437 VSS VSS.n1074 0.0213333
R7438 VSS.n6640 VSS.n1059 0.0213333
R7439 VSS.n6173 VSS.n6172 0.0213333
R7440 VSS.n7734 VSS 0.0213333
R7441 VSS.n7720 VSS.n7719 0.0213333
R7442 VSS.n7702 VSS 0.0213333
R7443 VSS.n7688 VSS.n7687 0.0213333
R7444 VSS.n7670 VSS 0.0213333
R7445 VSS.n7656 VSS.n7655 0.0213333
R7446 VSS.n7638 VSS 0.0213333
R7447 VSS VSS.n150 0.0213333
R7448 VSS.n1 VSS.n0 0.0211485
R7449 VSS VSS.n1 0.0211485
R7450 VSS.n5806 VSS.n5805 0.0208125
R7451 VSS.n7544 VSS.n7543 0.0205925
R7452 VSS.n3380 VSS.n3378 0.0202917
R7453 VSS.n6097 VSS.n6096 0.02024
R7454 VSS.n6098 VSS.n6097 0.02024
R7455 VSS.n576 VSS.n575 0.02024
R7456 VSS.n577 VSS.n576 0.02024
R7457 VSS.n476 VSS.n475 0.02024
R7458 VSS.n477 VSS.n476 0.02024
R7459 VSS.n7301 VSS.n7300 0.02024
R7460 VSS.n7302 VSS.n7301 0.02024
R7461 VSS.n276 VSS.n275 0.02024
R7462 VSS.n277 VSS.n276 0.02024
R7463 VSS.n7553 VSS.n111 0.02024
R7464 VSS.n7554 VSS.n7553 0.02024
R7465 VSS.n234 VSS.n233 0.02024
R7466 VSS.n235 VSS.n234 0.02024
R7467 VSS.n7514 VSS.n7513 0.02024
R7468 VSS.n7515 VSS.n7514 0.02024
R7469 VSS.n1860 VSS.n1859 0.02024
R7470 VSS.n1859 VSS.n1858 0.02024
R7471 VSS.n1352 VSS.n1351 0.02024
R7472 VSS.n1353 VSS.n1352 0.02024
R7473 VSS.n1333 VSS.n1332 0.02024
R7474 VSS.n1338 VSS.n1332 0.02024
R7475 VSS.n6361 VSS.n1177 0.02024
R7476 VSS.n6362 VSS.n6361 0.02024
R7477 VSS.n1208 VSS.n1207 0.02024
R7478 VSS.n1213 VSS.n1207 0.02024
R7479 VSS.n1199 VSS.n1198 0.02024
R7480 VSS.n1200 VSS.n1199 0.02024
R7481 VSS.n2708 VSS 0.0198529
R7482 VSS.n2699 VSS 0.0198529
R7483 VSS.n2664 VSS.t94 0.01977
R7484 VSS.t94 VSS.n2662 0.01977
R7485 VSS.n2678 VSS.t43 0.01977
R7486 VSS.t43 VSS.n2676 0.01977
R7487 VSS.n2692 VSS.t42 0.01977
R7488 VSS.t42 VSS.n2690 0.01977
R7489 VSS.n7550 VSS.t11 0.01977
R7490 VSS.n1722 VSS.t11 0.01977
R7491 VSS.n1722 VSS.t39 0.01977
R7492 VSS.n1722 VSS.t29 0.01977
R7493 VSS.n1837 VSS.t6 0.01977
R7494 VSS.t17 VSS.n1845 0.01977
R7495 VSS.n1846 VSS.t17 0.01977
R7496 VSS.n1837 VSS.t33 0.01977
R7497 VSS.t13 VSS.n1733 0.01977
R7498 VSS.n1764 VSS.t13 0.01977
R7499 VSS.n1764 VSS.t21 0.01977
R7500 VSS.n1722 VSS.t26 0.01977
R7501 VSS.n1764 VSS.t15 0.01977
R7502 VSS.n1722 VSS.t23 0.01977
R7503 VSS.n1764 VSS.t7 0.01977
R7504 VSS.n1764 VSS.t36 0.01977
R7505 VSS.n1837 VSS.t1 0.01977
R7506 VSS.n1837 VSS.t27 0.01977
R7507 VSS.n1846 VSS.t37 0.01977
R7508 VSS.n1846 VSS.t25 0.01977
R7509 VSS.n1837 VSS.t35 0.01977
R7510 VSS.n1846 VSS.t38 0.01977
R7511 VSS.n1846 VSS.t20 0.01977
R7512 VSS.n1846 VSS.t9 0.01977
R7513 VSS.n1837 VSS.t14 0.01977
R7514 VSS.t28 VSS.n1776 0.01977
R7515 VSS.n1837 VSS.t28 0.01977
R7516 VSS.n1764 VSS.t3 0.01977
R7517 VSS.n1764 VSS.t31 0.01977
R7518 VSS.n1722 VSS.t0 0.01977
R7519 VSS.n1722 VSS.t8 0.01977
R7520 VSS.n1722 VSS.t19 0.01977
R7521 VSS.n1764 VSS.t10 0.01977
R7522 VSS.n1837 VSS.t2 0.01977
R7523 VSS.n1846 VSS.t34 0.01977
R7524 VSS.n6359 VSS.t24 0.01977
R7525 VSS.t12 VSS.n1853 0.01977
R7526 VSS.n6359 VSS.t12 0.01977
R7527 VSS.n6359 VSS.t4 0.01977
R7528 VSS.n6359 VSS.t30 0.01977
R7529 VSS.n6359 VSS.t16 0.01977
R7530 VSS.n6359 VSS.t32 0.01977
R7531 VSS.n6359 VSS.t18 0.01977
R7532 VSS.n1846 VSS.t22 0.01977
R7533 VSS.n6359 VSS.t5 0.01977
R7534 VSS.n2698 VSS.n2696 0.0195238
R7535 VSS.n2693 VSS 0.0195238
R7536 VSS VSS.n2704 0.0195238
R7537 VSS.n2707 VSS.n2705 0.0195238
R7538 VSS.n2636 VSS 0.0195238
R7539 VSS.n2647 VSS 0.0195238
R7540 VSS VSS.n2671 0.0195238
R7541 VSS VSS.n2685 0.0195238
R7542 VSS VSS.n161 0.0195238
R7543 VSS.n1654 VSS 0.0195238
R7544 VSS.n1537 VSS 0.0195238
R7545 VSS.n1401 VSS 0.0195238
R7546 VSS.n1498 VSS 0.0195238
R7547 VSS.n290 VSS 0.0195238
R7548 VSS VSS.n1619 0.0195238
R7549 VSS VSS.n1554 0.0195238
R7550 VSS VSS.n1485 0.0195238
R7551 VSS VSS.n1378 0.0195238
R7552 VSS.n1297 VSS.n1296 0.01925
R7553 VSS.n6141 VSS.n6139 0.0187292
R7554 VSS.n7752 VSS.n7751 0.0187292
R7555 VSS.n3417 VSS.n3416 0.0182083
R7556 VSS.n83 VSS.n82 0.0178611
R7557 VSS.n6909 VSS.n6908 0.0178611
R7558 VSS.n6953 VSS.n6952 0.0178611
R7559 VSS.n6161 VSS.n6160 0.0178611
R7560 VSS.n7294 VSS.n7293 0.0178611
R7561 VSS.n107 VSS.n106 0.0178611
R7562 VSS.n184 VSS.n183 0.0178611
R7563 VSS.n380 VSS.n379 0.0178611
R7564 VSS.n5132 VSS.n5131 0.0178611
R7565 VSS.n5194 VSS.n5193 0.0178611
R7566 VSS.n3958 VSS.n3957 0.0178611
R7567 VSS.n5439 VSS.n5438 0.0178611
R7568 VSS.n4768 VSS.n4767 0.0178611
R7569 VSS.n5006 VSS.n5005 0.0178611
R7570 VSS.n4266 VSS.n4265 0.0178611
R7571 VSS.n4456 VSS.n4455 0.0178611
R7572 VSS.n4411 VSS.n4410 0.0178611
R7573 VSS.n4547 VSS.n4546 0.0178611
R7574 VSS.n4501 VSS.n4500 0.0178611
R7575 VSS.n4375 VSS.n4374 0.0178611
R7576 VSS.n4298 VSS.n4297 0.0178611
R7577 VSS.n3883 VSS.n3882 0.0178611
R7578 VSS.n4312 VSS.n4311 0.0178611
R7579 VSS.n4351 VSS.n4350 0.0178611
R7580 VSS.n4650 VSS.n4647 0.0178611
R7581 VSS.n4816 VSS.n4193 0.0178611
R7582 VSS.n4437 VSS.n4436 0.0178611
R7583 VSS.n4871 VSS.n4870 0.0178611
R7584 VSS.n4150 VSS.n4149 0.0178611
R7585 VSS.n2467 VSS.n2466 0.0178611
R7586 VSS.n4840 VSS.n4838 0.0178611
R7587 VSS.n4915 VSS.n4914 0.0178611
R7588 VSS.n5124 VSS.n5122 0.0178611
R7589 VSS.n4248 VSS.n4247 0.0178611
R7590 VSS.n4744 VSS.n4226 0.0178611
R7591 VSS.n4712 VSS.n4710 0.0178611
R7592 VSS.n5186 VSS.n5184 0.0178611
R7593 VSS.n4017 VSS.n3910 0.0178611
R7594 VSS.n4023 VSS.n4022 0.0178611
R7595 VSS.n4001 VSS.n4000 0.0178611
R7596 VSS.n4073 VSS.n4072 0.0178611
R7597 VSS.n3950 VSS.n3937 0.0178611
R7598 VSS.n3787 VSS.n3786 0.0178611
R7599 VSS.n3689 VSS.n3688 0.0178611
R7600 VSS.n3591 VSS.n3590 0.0178611
R7601 VSS.n3494 VSS.n3493 0.0178611
R7602 VSS.n3397 VSS.n3396 0.0178611
R7603 VSS.n2833 VSS.n2832 0.0178611
R7604 VSS.n5622 VSS.n2509 0.0178611
R7605 VSS.n2560 VSS.n2558 0.0178611
R7606 VSS.n2608 VSS.n2607 0.0178611
R7607 VSS.n469 VSS.n468 0.0178611
R7608 VSS.n436 VSS.n435 0.0178611
R7609 VSS.n2737 VSS.n2736 0.0178611
R7610 VSS.n7098 VSS.n7096 0.0178611
R7611 VSS.n7462 VSS.n7461 0.0178611
R7612 VSS.n7506 VSS.n7505 0.0178611
R7613 VSS.n669 VSS.n666 0.0178611
R7614 VSS.n828 VSS.n826 0.0178611
R7615 VSS.n6681 VSS.n6680 0.0178611
R7616 VSS.n7051 VSS.n7050 0.0178611
R7617 VSS.n780 VSS.n777 0.0178611
R7618 VSS.n7078 VSS.n7076 0.0178611
R7619 VSS.n651 VSS.n649 0.0178611
R7620 VSS.n567 VSS.n566 0.0178611
R7621 VSS.n694 VSS.n692 0.0178611
R7622 VSS.n7354 VSS.n7353 0.0178611
R7623 VSS.n7609 VSS.n7606 0.0178611
R7624 VSS.n7175 VSS.n7108 0.0178611
R7625 VSS.n7138 VSS.n7136 0.0178611
R7626 VSS.n7146 VSS.n7145 0.0178611
R7627 VSS.n6901 VSS.n712 0.0178611
R7628 VSS.n845 VSS.n843 0.0178611
R7629 VSS.n893 VSS.n891 0.0178611
R7630 VSS.n911 VSS.n909 0.0178611
R7631 VSS.n6873 VSS.n6871 0.0178611
R7632 VSS.n6945 VSS.n6943 0.0178611
R7633 VSS.n1076 VSS.n1075 0.0178611
R7634 VSS.n1110 VSS.n1109 0.0178611
R7635 VSS.n6487 VSS.n6486 0.0178611
R7636 VSS.n1161 VSS.n1160 0.0178611
R7637 VSS.n1277 VSS.n1276 0.0178611
R7638 VSS.n943 VSS.n937 0.0178611
R7639 VSS.n6423 VSS.n6422 0.0176877
R7640 VSS.n4461 VSS.n4451 0.0175455
R7641 VSS.n4461 VSS 0.0175455
R7642 VSS VSS.n4459 0.0175455
R7643 VSS.n4459 VSS 0.0175455
R7644 VSS.n5279 VSS.n2862 0.0175455
R7645 VSS.n5279 VSS 0.0175455
R7646 VSS VSS.n3886 0.0175455
R7647 VSS.n3886 VSS 0.0175455
R7648 VSS.n4322 VSS.n4308 0.0175455
R7649 VSS.n4322 VSS 0.0175455
R7650 VSS VSS.n4315 0.0175455
R7651 VSS.n4315 VSS 0.0175455
R7652 VSS.n4633 VSS.n4280 0.0175455
R7653 VSS.n4633 VSS 0.0175455
R7654 VSS VSS.n4354 0.0175455
R7655 VSS.n4354 VSS 0.0175455
R7656 VSS VSS.n4487 0.0175455
R7657 VSS.n4510 VSS 0.0175455
R7658 VSS.n4573 VSS 0.0175455
R7659 VSS.n4377 VSS 0.0175455
R7660 VSS VSS.n4992 0.0175455
R7661 VSS.n5015 VSS 0.0175455
R7662 VSS.n4774 VSS 0.0175455
R7663 VSS.n4750 VSS 0.0175455
R7664 VSS.n5662 VSS 0.0175455
R7665 VSS.n2439 VSS 0.0175455
R7666 VSS.n5091 VSS.n4135 0.0175455
R7667 VSS.n5091 VSS 0.0175455
R7668 VSS.n4136 VSS 0.0175455
R7669 VSS.n4881 VSS 0.0175455
R7670 VSS.n4879 VSS 0.0175455
R7671 VSS.n3802 VSS 0.0175455
R7672 VSS VSS.n3771 0.0175455
R7673 VSS.n3771 VSS 0.0175455
R7674 VSS.n3705 VSS 0.0175455
R7675 VSS VSS.n3673 0.0175455
R7676 VSS.n3673 VSS 0.0175455
R7677 VSS.n3607 VSS 0.0175455
R7678 VSS VSS.n3575 0.0175455
R7679 VSS.n3575 VSS 0.0175455
R7680 VSS.n3510 VSS 0.0175455
R7681 VSS VSS.n3478 0.0175455
R7682 VSS.n3478 VSS 0.0175455
R7683 VSS.n3413 VSS 0.0175455
R7684 VSS VSS.n3381 0.0175455
R7685 VSS.n3381 VSS 0.0175455
R7686 VSS.n5351 VSS 0.0175455
R7687 VSS.n5353 VSS 0.0175455
R7688 VSS VSS.n5353 0.0175455
R7689 VSS.n5453 VSS 0.0175455
R7690 VSS VSS.n5423 0.0175455
R7691 VSS.n5423 VSS 0.0175455
R7692 VSS.n5787 VSS.n2374 0.0175455
R7693 VSS.n5787 VSS 0.0175455
R7694 VSS VSS.n2376 0.0175455
R7695 VSS.n2376 VSS 0.0175455
R7696 VSS.n5755 VSS.n2393 0.0175455
R7697 VSS.n5755 VSS 0.0175455
R7698 VSS VSS.n2395 0.0175455
R7699 VSS.n2395 VSS 0.0175455
R7700 VSS.n5723 VSS.n2412 0.0175455
R7701 VSS.n5723 VSS 0.0175455
R7702 VSS VSS.n2414 0.0175455
R7703 VSS.n2414 VSS 0.0175455
R7704 VSS.n5691 VSS.n2430 0.0175455
R7705 VSS.n5691 VSS 0.0175455
R7706 VSS VSS.n5689 0.0175455
R7707 VSS.n5689 VSS 0.0175455
R7708 VSS.n2492 VSS 0.0175455
R7709 VSS.n2517 VSS.n2514 0.0175455
R7710 VSS.n2517 VSS 0.0175455
R7711 VSS.n2622 VSS 0.0175455
R7712 VSS.n2622 VSS 0.0175455
R7713 VSS.n2594 VSS.n2537 0.0175455
R7714 VSS.n2594 VSS 0.0175455
R7715 VSS.n2555 VSS 0.0175455
R7716 VSS.n2555 VSS 0.0175455
R7717 VSS.n2546 VSS.n2545 0.0175455
R7718 VSS.n2545 VSS 0.0175455
R7719 VSS.n2590 VSS 0.0175455
R7720 VSS.n2590 VSS 0.0175455
R7721 VSS.n2618 VSS.n2521 0.0175455
R7722 VSS.n2618 VSS 0.0175455
R7723 VSS VSS.n2610 0.0175455
R7724 VSS.n2610 VSS 0.0175455
R7725 VSS.n7468 VSS.n309 0.0175455
R7726 VSS.n7468 VSS 0.0175455
R7727 VSS VSS.n7466 0.0175455
R7728 VSS.n7466 VSS 0.0175455
R7729 VSS.n6671 VSS.n6663 0.0175455
R7730 VSS.n6671 VSS 0.0175455
R7731 VSS.n6677 VSS 0.0175455
R7732 VSS.n6677 VSS 0.0175455
R7733 VSS.n7058 VSS.n783 0.0175455
R7734 VSS.n7058 VSS 0.0175455
R7735 VSS.n7054 VSS 0.0175455
R7736 VSS.n7054 VSS 0.0175455
R7737 VSS.n770 VSS.n763 0.0175455
R7738 VSS.n770 VSS 0.0175455
R7739 VSS.n774 VSS 0.0175455
R7740 VSS.n774 VSS 0.0175455
R7741 VSS.n596 VSS.n552 0.0175455
R7742 VSS.n596 VSS 0.0175455
R7743 VSS.n593 VSS 0.0175455
R7744 VSS.n7537 VSS.n7536 0.0175455
R7745 VSS.n7536 VSS 0.0175455
R7746 VSS.n7533 VSS 0.0175455
R7747 VSS.n498 VSS.n455 0.0175455
R7748 VSS.n498 VSS 0.0175455
R7749 VSS.n495 VSS 0.0175455
R7750 VSS.n386 VSS 0.0175455
R7751 VSS.n344 VSS 0.0175455
R7752 VSS.n218 VSS.n217 0.0175455
R7753 VSS.n218 VSS 0.0175455
R7754 VSS.n221 VSS 0.0175455
R7755 VSS.n7575 VSS.n93 0.0175455
R7756 VSS.n7575 VSS 0.0175455
R7757 VSS.n7572 VSS 0.0175455
R7758 VSS.n7322 VSS.n7279 0.0175455
R7759 VSS.n7322 VSS 0.0175455
R7760 VSS.n7320 VSS 0.0175455
R7761 VSS.n6641 VSS.n6640 0.0175455
R7762 VSS.n6640 VSS 0.0175455
R7763 VSS.n6638 VSS 0.0175455
R7764 VSS.n6638 VSS 0.0175455
R7765 VSS.n6569 VSS 0.0175455
R7766 VSS VSS.n6553 0.0175455
R7767 VSS.n6553 VSS 0.0175455
R7768 VSS.n6502 VSS 0.0175455
R7769 VSS VSS.n6472 0.0175455
R7770 VSS.n6472 VSS 0.0175455
R7771 VSS.n6416 VSS 0.0175455
R7772 VSS VSS.n6400 0.0175455
R7773 VSS.n6400 VSS 0.0175455
R7774 VSS.n1292 VSS 0.0175455
R7775 VSS VSS.n1262 0.0175455
R7776 VSS.n1262 VSS 0.0175455
R7777 VSS.n6840 VSS 0.0175455
R7778 VSS.n6838 VSS 0.0175455
R7779 VSS.n6838 VSS 0.0175455
R7780 VSS VSS.n6143 0.0175455
R7781 VSS.n6173 VSS 0.0175455
R7782 VSS.n6173 VSS 0.0175455
R7783 VSS.n7731 VSS.n17 0.0175455
R7784 VSS.n7731 VSS 0.0175455
R7785 VSS VSS.n19 0.0175455
R7786 VSS.n19 VSS 0.0175455
R7787 VSS.n7699 VSS.n36 0.0175455
R7788 VSS.n7699 VSS 0.0175455
R7789 VSS VSS.n38 0.0175455
R7790 VSS.n38 VSS 0.0175455
R7791 VSS.n7667 VSS.n55 0.0175455
R7792 VSS.n7667 VSS 0.0175455
R7793 VSS VSS.n57 0.0175455
R7794 VSS.n57 VSS 0.0175455
R7795 VSS.n7635 VSS.n73 0.0175455
R7796 VSS.n7635 VSS 0.0175455
R7797 VSS VSS.n7633 0.0175455
R7798 VSS.n7633 VSS 0.0175455
R7799 VSS.n143 VSS.n142 0.0173919
R7800 VSS.n7647 VSS.n7644 0.0173919
R7801 VSS.n7679 VSS.n7676 0.0173919
R7802 VSS.n7711 VSS.n7708 0.0173919
R7803 VSS.n6842 VSS.n6841 0.0173919
R7804 VSS.n1291 VSS.n1290 0.0173919
R7805 VSS.n6415 VSS.n6414 0.0173919
R7806 VSS.n6501 VSS.n6500 0.0173919
R7807 VSS.n6993 VSS.n6991 0.0173919
R7808 VSS.n881 VSS.n871 0.0173919
R7809 VSS.n7589 VSS.n7588 0.0173919
R7810 VSS.n7284 VSS.n7283 0.0173919
R7811 VSS.n7577 VSS.n7576 0.0173919
R7812 VSS.n190 VSS.n189 0.0173919
R7813 VSS.n97 VSS.n96 0.0173919
R7814 VSS.n201 VSS.n200 0.0173919
R7815 VSS.n2483 VSS.n2482 0.0173919
R7816 VSS.n5703 VSS.n5700 0.0173919
R7817 VSS.n5735 VSS.n5732 0.0173919
R7818 VSS.n5767 VSS.n5764 0.0173919
R7819 VSS.n5349 VSS.n5348 0.0173919
R7820 VSS.n3411 VSS.n3410 0.0173919
R7821 VSS.n3508 VSS.n3507 0.0173919
R7822 VSS.n3605 VSS.n3604 0.0173919
R7823 VSS.n4059 VSS.n4058 0.0173919
R7824 VSS.n4776 VSS.n4775 0.0173919
R7825 VSS.n4788 VSS.n4787 0.0173919
R7826 VSS.n4998 VSS.n4997 0.0173919
R7827 VSS.n4824 VSS.n4823 0.0173919
R7828 VSS.n4486 VSS.n4485 0.0173919
R7829 VSS.n4449 VSS.n4448 0.0173919
R7830 VSS.n4407 VSS.n4406 0.0173919
R7831 VSS.n4991 VSS.n4990 0.0173919
R7832 VSS.n4983 VSS.n4982 0.0173919
R7833 VSS.n4539 VSS.n4538 0.0173919
R7834 VSS.n4575 VSS.n4574 0.0173919
R7835 VSS.n4491 VSS.n4490 0.0173919
R7836 VSS.n4587 VSS.n4586 0.0173919
R7837 VSS.n4606 VSS.n4604 0.0173919
R7838 VSS.n4611 VSS.n4204 0.0173919
R7839 VSS.n4619 VSS.n4618 0.0173919
R7840 VSS.n5276 VSS.n5275 0.0173919
R7841 VSS.n4302 VSS.n4301 0.0173919
R7842 VSS.n5268 VSS.n5267 0.0173919
R7843 VSS.n4289 VSS.n4273 0.0173919
R7844 VSS.n4343 VSS.n4342 0.0173919
R7845 VSS.n4319 VSS.n4318 0.0173919
R7846 VSS.n4340 VSS.n4339 0.0173919
R7847 VSS.n4269 VSS.n4267 0.0173919
R7848 VSS.n4659 VSS.n4658 0.0173919
R7849 VSS.n4622 VSS.n4621 0.0173919
R7850 VSS.n4630 VSS.n4629 0.0173919
R7851 VSS.n4958 VSS.n4956 0.0173919
R7852 VSS.n4966 VSS.n4965 0.0173919
R7853 VSS.n4477 VSS.n4476 0.0173919
R7854 VSS.n5105 VSS.n5104 0.0173919
R7855 VSS.n4861 VSS.n4860 0.0173919
R7856 VSS.n5093 VSS.n5092 0.0173919
R7857 VSS.n5676 VSS.n5675 0.0173919
R7858 VSS.n4140 VSS.n4139 0.0173919
R7859 VSS.n5664 VSS.n5663 0.0173919
R7860 VSS.n4883 VSS.n4882 0.0173919
R7861 VSS.n4758 VSS.n4757 0.0173919
R7862 VSS.n4895 VSS.n4894 0.0173919
R7863 VSS.n4922 VSS.n4116 0.0173919
R7864 VSS.n4930 VSS.n4929 0.0173919
R7865 VSS.n4918 VSS.n4916 0.0173919
R7866 VSS.n5154 VSS.n5151 0.0173919
R7867 VSS.n5162 VSS.n5161 0.0173919
R7868 VSS.n4133 VSS.n4132 0.0173919
R7869 VSS.n5149 VSS.n5148 0.0173919
R7870 VSS.n5135 VSS.n5133 0.0173919
R7871 VSS.n5141 VSS.n2421 0.0173919
R7872 VSS.n4837 VSS.n4836 0.0173919
R7873 VSS.n4829 VSS.n4827 0.0173919
R7874 VSS.n4810 VSS.n4745 0.0173919
R7875 VSS.n4690 VSS.n4232 0.0173919
R7876 VSS.n4674 VSS.n4673 0.0173919
R7877 VSS.n4682 VSS.n4225 0.0173919
R7878 VSS.n4738 VSS.n4735 0.0173919
R7879 VSS.n4695 VSS.n4693 0.0173919
R7880 VSS.n4709 VSS.n4708 0.0173919
R7881 VSS.n4724 VSS.n4100 0.0173919
R7882 VSS.n4732 VSS.n4731 0.0173919
R7883 VSS.n4718 VSS.n4105 0.0173919
R7884 VSS.n5211 VSS.n5210 0.0173919
R7885 VSS.n5197 VSS.n5195 0.0173919
R7886 VSS.n5203 VSS.n2402 0.0173919
R7887 VSS.n4252 VSS.n4250 0.0173919
R7888 VSS.n4663 VSS.n4662 0.0173919
R7889 VSS.n4670 VSS.n4669 0.0173919
R7890 VSS.n4046 VSS.n4045 0.0173919
R7891 VSS.n4038 VSS.n4036 0.0173919
R7892 VSS.n4026 VSS.n4024 0.0173919
R7893 VSS.n4051 VSS.n4049 0.0173919
R7894 VSS.n4004 VSS.n4002 0.0173919
R7895 VSS.n4085 VSS.n3984 0.0173919
R7896 VSS.n4063 VSS.n4062 0.0173919
R7897 VSS.n4077 VSS.n4074 0.0173919
R7898 VSS.n3979 VSS.n3977 0.0173919
R7899 VSS.n4090 VSS.n4088 0.0173919
R7900 VSS.n4098 VSS.n4097 0.0173919
R7901 VSS.n3975 VSS.n3974 0.0173919
R7902 VSS.n3961 VSS.n3959 0.0173919
R7903 VSS.n3967 VSS.n2383 0.0173919
R7904 VSS.n5257 VSS.n5255 0.0173919
R7905 VSS.n5264 VSS.n3898 0.0173919
R7906 VSS.n4033 VSS.n4032 0.0173919
R7907 VSS.n3703 VSS.n3702 0.0173919
R7908 VSS.n3777 VSS.n3776 0.0173919
R7909 VSS.n3691 VSS.n3690 0.0173919
R7910 VSS.n3679 VSS.n3678 0.0173919
R7911 VSS.n3593 VSS.n3592 0.0173919
R7912 VSS.n3581 VSS.n3580 0.0173919
R7913 VSS.n3496 VSS.n3495 0.0173919
R7914 VSS.n3484 VSS.n3483 0.0173919
R7915 VSS.n3399 VSS.n3398 0.0173919
R7916 VSS.n3387 VSS.n3386 0.0173919
R7917 VSS.n5337 VSS.n5336 0.0173919
R7918 VSS.n2825 VSS.n2816 0.0173919
R7919 VSS.n5441 VSS.n5440 0.0173919
R7920 VSS.n5451 VSS.n5450 0.0173919
R7921 VSS.n3790 VSS.n3789 0.0173919
R7922 VSS.n3800 VSS.n3799 0.0173919
R7923 VSS.n3872 VSS.n3871 0.0173919
R7924 VSS.n5803 VSS.n5802 0.0173919
R7925 VSS.n5430 VSS.n5429 0.0173919
R7926 VSS.n5791 VSS.n5790 0.0173919
R7927 VSS.n5775 VSS.n5774 0.0173919
R7928 VSS.n5760 VSS.n5758 0.0173919
R7929 VSS.n5743 VSS.n5742 0.0173919
R7930 VSS.n5728 VSS.n5726 0.0173919
R7931 VSS.n5711 VSS.n5710 0.0173919
R7932 VSS.n5696 VSS.n5694 0.0173919
R7933 VSS.n2457 VSS.n2456 0.0173919
R7934 VSS.n2490 VSS.n2489 0.0173919
R7935 VSS.n2626 VSS.n2625 0.0173919
R7936 VSS.n2535 VSS.n2533 0.0173919
R7937 VSS.n2599 VSS.n2597 0.0173919
R7938 VSS.n2570 VSS.n2569 0.0173919
R7939 VSS.n2579 VSS.n2577 0.0173919
R7940 VSS.n2587 VSS.n2586 0.0173919
R7941 VSS.n2544 VSS.n2543 0.0173919
R7942 VSS.n2615 VSS.n2614 0.0173919
R7943 VSS.n5613 VSS.n5610 0.0173919
R7944 VSS.n388 VSS.n387 0.0173919
R7945 VSS.n400 VSS.n399 0.0173919
R7946 VSS.n461 VSS.n460 0.0173919
R7947 VSS.n7492 VSS.n7491 0.0173919
R7948 VSS.n648 VSS.n647 0.0173919
R7949 VSS.n500 VSS.n499 0.0173919
R7950 VSS.n560 VSS.n559 0.0173919
R7951 VSS.n598 VSS.n597 0.0173919
R7952 VSS.n7496 VSS.n7495 0.0173919
R7953 VSS.n610 VSS.n609 0.0173919
R7954 VSS.n635 VSS.n634 0.0173919
R7955 VSS.n527 VSS.n432 0.0173919
R7956 VSS.n678 VSS.n430 0.0173919
R7957 VSS.n665 VSS.n664 0.0173919
R7958 VSS.n657 VSS.n319 0.0173919
R7959 VSS.n6668 VSS.n6667 0.0173919
R7960 VSS.n825 VSS.n824 0.0173919
R7961 VSS.n7043 VSS.n7041 0.0173919
R7962 VSS.n7075 VSS.n756 0.0173919
R7963 VSS.n7070 VSS.n751 0.0173919
R7964 VSS.n7064 VSS.n7061 0.0173919
R7965 VSS.n7198 VSS.n7197 0.0173919
R7966 VSS.n7094 VSS.n7093 0.0173919
R7967 VSS.n7190 VSS.n7189 0.0173919
R7968 VSS.n7454 VSS.n7452 0.0173919
R7969 VSS.n767 VSS.n766 0.0173919
R7970 VSS.n640 VSS.n638 0.0173919
R7971 VSS.n7484 VSS.n7483 0.0173919
R7972 VSS.n2728 VSS.n2727 0.0173919
R7973 VSS.n510 VSS.n509 0.0173919
R7974 VSS.n7324 VSS.n7323 0.0173919
R7975 VSS.n370 VSS.n369 0.0173919
R7976 VSS.n7336 VSS.n7335 0.0173919
R7977 VSS.n7410 VSS.n7408 0.0173919
R7978 VSS.n7418 VSS.n7417 0.0173919
R7979 VSS.n7262 VSS.n7261 0.0173919
R7980 VSS.n7374 VSS.n7254 0.0173919
R7981 VSS.n7358 VSS.n702 0.0173919
R7982 VSS.n7366 VSS.n91 0.0173919
R7983 VSS.n7379 VSS.n7378 0.0173919
R7984 VSS.n7621 VSS.n84 0.0173919
R7985 VSS.n7616 VSS.n64 0.0173919
R7986 VSS.n691 VSS.n690 0.0173919
R7987 VSS.n683 VSS.n681 0.0173919
R7988 VSS.n422 VSS.n339 0.0173919
R7989 VSS.n7169 VSS.n7166 0.0173919
R7990 VSS.n7121 VSS.n7119 0.0173919
R7991 VSS.n7128 VSS.n7126 0.0173919
R7992 VSS.n7155 VSS.n722 0.0173919
R7993 VSS.n7163 VSS.n7162 0.0173919
R7994 VSS.n7149 VSS.n7147 0.0173919
R7995 VSS.n6895 VSS.n6894 0.0173919
R7996 VSS.n7244 VSS.n7242 0.0173919
R7997 VSS.n7252 VSS.n7251 0.0173919
R7998 VSS.n6926 VSS.n6925 0.0173919
R7999 VSS.n6912 VSS.n6910 0.0173919
R8000 VSS.n6918 VSS.n45 0.0173919
R8001 VSS.n7179 VSS.n7177 0.0173919
R8002 VSS.n7186 VSS.n7087 0.0173919
R8003 VSS.n7116 VSS.n7115 0.0173919
R8004 VSS.n7019 VSS.n7017 0.0173919
R8005 VSS.n7027 VSS.n7026 0.0173919
R8006 VSS.n889 VSS.n888 0.0173919
R8007 VSS.n899 VSS.n853 0.0173919
R8008 VSS.n907 VSS.n906 0.0173919
R8009 VSS.n7001 VSS.n7000 0.0173919
R8010 VSS.n6870 VSS.n6869 0.0173919
R8011 VSS.n6876 VSS.n6855 0.0173919
R8012 VSS.n6882 VSS.n919 0.0173919
R8013 VSS.n6890 VSS.n6889 0.0173919
R8014 VSS.n6970 VSS.n6969 0.0173919
R8015 VSS.n6956 VSS.n6954 0.0173919
R8016 VSS.n6962 VSS.n26 0.0173919
R8017 VSS.n842 VSS.n841 0.0173919
R8018 VSS.n834 VSS.n794 0.0173919
R8019 VSS.n817 VSS.n806 0.0173919
R8020 VSS.n6568 VSS.n6567 0.0173919
R8021 VSS.n1087 VSS.n1086 0.0173919
R8022 VSS.n6556 VSS.n6555 0.0173919
R8023 VSS.n1121 VSS.n1120 0.0173919
R8024 VSS.n6489 VSS.n6488 0.0173919
R8025 VSS.n6477 VSS.n6476 0.0173919
R8026 VSS.n6403 VSS.n6402 0.0173919
R8027 VSS.n1172 VSS.n1171 0.0173919
R8028 VSS.n1279 VSS.n1278 0.0173919
R8029 VSS.n1267 VSS.n1266 0.0173919
R8030 VSS.n6853 VSS.n6852 0.0173919
R8031 VSS.n955 VSS.n954 0.0173919
R8032 VSS.n6159 VSS.n6158 0.0173919
R8033 VSS.n6150 VSS.n6149 0.0173919
R8034 VSS.n1074 VSS.n1073 0.0173919
R8035 VSS.n1065 VSS.n1059 0.0173919
R8036 VSS.n6693 VSS.n6692 0.0173919
R8037 VSS.n7747 VSS.n7746 0.0173919
R8038 VSS.n6172 VSS.n6171 0.0173919
R8039 VSS.n7735 VSS.n7734 0.0173919
R8040 VSS.n7719 VSS.n7718 0.0173919
R8041 VSS.n7704 VSS.n7702 0.0173919
R8042 VSS.n7687 VSS.n7686 0.0173919
R8043 VSS.n7672 VSS.n7670 0.0173919
R8044 VSS.n7655 VSS.n7654 0.0173919
R8045 VSS.n7640 VSS.n7638 0.0173919
R8046 VSS.n174 VSS.n173 0.0173919
R8047 VSS.n150 VSS.n149 0.0173919
R8048 VSS.n6095 VSS 0.017343
R8049 VSS.n6099 VSS 0.017343
R8050 VSS.n1197 VSS 0.017343
R8051 VSS VSS.n1201 0.017343
R8052 VSS VSS.n1209 0.017343
R8053 VSS.n1214 VSS 0.017343
R8054 VSS.n1176 VSS 0.017343
R8055 VSS.n6363 VSS 0.017343
R8056 VSS VSS.n1334 0.017343
R8057 VSS VSS.n1339 0.017343
R8058 VSS.n1339 VSS 0.017343
R8059 VSS.n1350 VSS 0.017343
R8060 VSS VSS.n1354 0.017343
R8061 VSS VSS.n1861 0.017343
R8062 VSS.n1857 VSS 0.017343
R8063 VSS.n6100 VSS.n6099 0.0171826
R8064 VSS.n1201 VSS.n958 0.0171826
R8065 VSS.n6366 VSS.n6363 0.0171826
R8066 VSS.n1354 VSS.n1349 0.0171826
R8067 VSS.n1857 VSS.n1038 0.0171826
R8068 VSS.n6420 VSS.n6419 0.0171667
R8069 VSS.n1323 VSS.n1214 0.0170222
R8070 VSS VSS.n7757 0.0168222
R8071 VSS.n3427 VSS.n3426 0.016646
R8072 VSS.n1764 VSS.n1743 0.0163425
R8073 VSS.n1837 VSS.n1826 0.0163425
R8074 VSS.n1846 VSS.n1466 0.0163425
R8075 VSS.n1837 VSS.n1786 0.0163425
R8076 VSS.n1764 VSS.n1601 0.0163425
R8077 VSS.n1765 VSS.n1764 0.0163425
R8078 VSS.n1722 VSS.n1671 0.0163425
R8079 VSS.n6359 VSS.n1862 0.0163425
R8080 VSS.n6359 VSS.n1183 0.0163425
R8081 VSS.n6359 VSS.n1342 0.0163425
R8082 VSS.n6360 VSS.n6359 0.0163425
R8083 VSS.n6359 VSS.n1324 0.0163425
R8084 VSS.n6359 VSS.n1192 0.0163425
R8085 VSS.n6359 VSS.n1193 0.0163425
R8086 VSS.n6129 VSS.n6128 0.0161252
R8087 VSS.n4 VSS.n3 0.0161252
R8088 VSS.n4509 VSS 0.016125
R8089 VSS VSS.n4548 0.016125
R8090 VSS.n5014 VSS 0.016125
R8091 VSS VSS.n4769 0.016125
R8092 VSS VSS.n2468 0.016125
R8093 VSS VSS.n4151 0.016125
R8094 VSS.n4878 VSS 0.016125
R8095 VSS.n592 VSS 0.016125
R8096 VSS.n7532 VSS 0.016125
R8097 VSS.n494 VSS 0.016125
R8098 VSS VSS.n381 0.016125
R8099 VSS VSS.n222 0.016125
R8100 VSS.n7571 VSS 0.016125
R8101 VSS.n7319 VSS 0.016125
R8102 VSS.n1462 VSS.n1381 0.0157702
R8103 VSS.n1587 VSS.n1557 0.0157702
R8104 VSS.n1707 VSS.n1637 0.0157702
R8105 VSS.n1728 VSS.n1647 0.0157702
R8106 VSS.n1775 VSS.n1580 0.0157702
R8107 VSS.n1771 VSS.n1566 0.0157702
R8108 VSS.n1472 VSS.n1364 0.0157702
R8109 VSS.n1528 VSS.n1511 0.0157702
R8110 VSS.n1757 VSS.n1573 0.0157702
R8111 VSS.n1749 VSS.n1570 0.0157702
R8112 VSS.n1714 VSS.n1634 0.0157702
R8113 VSS.n1687 VSS.n1644 0.0157702
R8114 VSS.n1694 VSS.n1639 0.0157702
R8115 VSS.n1737 VSS.n1577 0.0157702
R8116 VSS.n1819 VSS.n1508 0.0157702
R8117 VSS.n1832 VSS.n1515 0.0157702
R8118 VSS.n1422 VSS.n1393 0.0157702
R8119 VSS.n1429 VSS.n1368 0.0157702
R8120 VSS.n1810 VSS.n1523 0.0157702
R8121 VSS.n1799 VSS.n1518 0.0157702
R8122 VSS.n1451 VSS.n1389 0.0157702
R8123 VSS.n1441 VSS.n1384 0.0157702
R8124 VSS.n1778 VSS.n1493 0.0157702
R8125 VSS.n1789 VSS.n1488 0.0157702
R8126 VSS.n1595 VSS.n1562 0.0157702
R8127 VSS.n1663 VSS.n1627 0.0157702
R8128 VSS.n1677 VSS.n1622 0.0157702
R8129 VSS.n1412 VSS.n1397 0.0157702
R8130 VSS.n1297 VSS.n1233 0.0156042
R8131 VSS.n1764 VSS.n1591 0.0155925
R8132 VSS.n1722 VSS.n1701 0.0155925
R8133 VSS.n1722 VSS.n1711 0.0155925
R8134 VSS.n1722 VSS.n1721 0.0155925
R8135 VSS.n1723 VSS.n1722 0.0155925
R8136 VSS.n1764 VSS.n1610 0.0155925
R8137 VSS.n1837 VSS.n1816 0.0155925
R8138 VSS.n1846 VSS.n1476 0.0155925
R8139 VSS.n1847 VSS.n1846 0.0155925
R8140 VSS.n1838 VSS.n1837 0.0155925
R8141 VSS.n1764 VSS.n1753 0.0155925
R8142 VSS.n1764 VSS.n1763 0.0155925
R8143 VSS.n1722 VSS.n1691 0.0155925
R8144 VSS.n1837 VSS.n1836 0.0155925
R8145 VSS.n1846 VSS.n1436 0.0155925
R8146 VSS.n1846 VSS.n1426 0.0155925
R8147 VSS.n1837 VSS.n1806 0.0155925
R8148 VSS.n1846 VSS.n1446 0.0155925
R8149 VSS.n1846 VSS.n1456 0.0155925
R8150 VSS.n1837 VSS.n1796 0.0155925
R8151 VSS.n1722 VSS.n1681 0.0155925
R8152 VSS.n7545 VSS.n7544 0.0151004
R8153 VSS.n538 VSS.n537 0.0151004
R8154 VSS.n358 VSS.n357 0.0151004
R8155 VSS.n6321 VSS.n6320 0.0150187
R8156 VSS VSS.n6351 0.0149369
R8157 VSS.n257 VSS.n256 0.0148765
R8158 VSS.n440 VSS.n439 0.0148765
R8159 VSS.n7272 VSS.n7271 0.0148765
R8160 VSS.n211 VSS.n210 0.0148765
R8161 VSS.n479 VSS.n472 0.0146
R8162 VSS.n3378 VSS.n2916 0.0145625
R8163 VSS.n7757 VSS 0.0144825
R8164 VSS.n579 VSS.n572 0.0143762
R8165 VSS.n7556 VSS.n109 0.0141524
R8166 VSS.n7517 VSS.n7510 0.0141524
R8167 VSS.n2708 VSS.n2707 0.0141524
R8168 VSS.n7304 VSS.n7297 0.0141524
R8169 VSS.n280 VSS.n279 0.0141524
R8170 VSS.n238 VSS.n237 0.0141524
R8171 VSS.n160 VSS 0.01413
R8172 VSS.n1190 VSS.n1189 0.0137575
R8173 VSS.n1330 VSS.n1329 0.0137575
R8174 VSS.n6357 VSS.n6356 0.0137575
R8175 VSS.n6308 VSS.n6307 0.0136341
R8176 VSS.n1196 VSS.n1195 0.0135337
R8177 VSS.n1186 VSS.n1185 0.0135337
R8178 VSS.n1181 VSS.n1180 0.0135337
R8179 VSS.n3621 VSS.n3620 0.013521
R8180 VSS.n4515 VSS.n4514 0.0135208
R8181 VSS.n4569 VSS.n4567 0.0135208
R8182 VSS.n5020 VSS.n5019 0.0135208
R8183 VSS.n5042 VSS.n5041 0.0135208
R8184 VSS.n4516 VSS.n4515 0.0133116
R8185 VSS.n4567 VSS.n4566 0.0133116
R8186 VSS.n5021 VSS.n5020 0.0133116
R8187 VSS.n5043 VSS.n5042 0.0133116
R8188 VSS.n5656 VSS.n5655 0.0133116
R8189 VSS.n1360 VSS.n1359 0.0133099
R8190 VSS.n3807 VSS.n3806 0.0132939
R8191 VSS.n3710 VSS.n3709 0.0132939
R8192 VSS.n3612 VSS.n3611 0.0132939
R8193 VSS.n3515 VSS.n3514 0.0132939
R8194 VSS.n3418 VSS.n3417 0.0132939
R8195 VSS.n3321 VSS.n3320 0.0132939
R8196 VSS.n5458 VSS.n5457 0.0132939
R8197 VSS.n5807 VSS.n5806 0.0132939
R8198 VSS.n6421 VSS.n6420 0.0132939
R8199 VSS.n6139 VSS.n6138 0.0132939
R8200 VSS.n7753 VSS.n7752 0.0132939
R8201 VSS.n6506 VSS.n6505 0.013121
R8202 VSS.n6094 VSS.n6093 0.0128095
R8203 VSS.n1203 VSS.n1202 0.0128095
R8204 VSS.n1337 VSS.n1336 0.0128095
R8205 VSS.n1856 VSS.n1855 0.0128095
R8206 VSS.n6353 VSS.n6352 0.0128095
R8207 VSS.n1326 VSS.n1325 0.0125857
R8208 VSS.n1356 VSS.n1355 0.0125857
R8209 VSS.n6089 VSS.n1194 0.0124386
R8210 VSS.n1212 VSS.n1211 0.0123619
R8211 VSS.n1463 VSS 0.01225
R8212 VSS VSS.n1461 0.01225
R8213 VSS.n1461 VSS 0.01225
R8214 VSS.n1588 VSS 0.01225
R8215 VSS VSS.n1584 0.01225
R8216 VSS.n1584 VSS 0.01225
R8217 VSS VSS.n1662 0.01225
R8218 VSS.n1668 VSS 0.01225
R8219 VSS.n1668 VSS 0.01225
R8220 VSS VSS.n1693 0.01225
R8221 VSS.n1698 VSS 0.01225
R8222 VSS.n1698 VSS 0.01225
R8223 VSS VSS.n1713 0.01225
R8224 VSS.n1718 VSS 0.01225
R8225 VSS.n1718 VSS 0.01225
R8226 VSS.n1708 VSS 0.01225
R8227 VSS VSS.n1704 0.01225
R8228 VSS.n1704 VSS 0.01225
R8229 VSS VSS.n1661 0.01225
R8230 VSS VSS.n1727 0.01225
R8231 VSS.n1727 VSS 0.01225
R8232 VSS.n1598 VSS 0.01225
R8233 VSS VSS.n1594 0.01225
R8234 VSS.n1594 VSS 0.01225
R8235 VSS.n1760 VSS 0.01225
R8236 VSS VSS.n1756 0.01225
R8237 VSS.n1756 VSS 0.01225
R8238 VSS.n1607 VSS 0.01225
R8239 VSS VSS.n1604 0.01225
R8240 VSS.n1604 VSS 0.01225
R8241 VSS VSS.n1581 0.01225
R8242 VSS VSS.n1770 0.01225
R8243 VSS.n1770 VSS 0.01225
R8244 VSS.n1813 VSS 0.01225
R8245 VSS VSS.n1809 0.01225
R8246 VSS.n1809 VSS 0.01225
R8247 VSS VSS.n1777 0.01225
R8248 VSS.n1782 VSS 0.01225
R8249 VSS.n1782 VSS 0.01225
R8250 VSS.n1473 VSS 0.01225
R8251 VSS VSS.n1469 0.01225
R8252 VSS.n1469 VSS 0.01225
R8253 VSS.n1416 VSS 0.01225
R8254 VSS.n1850 VSS 0.01225
R8255 VSS VSS.n1850 0.01225
R8256 VSS.n1529 VSS 0.01225
R8257 VSS.n1841 VSS 0.01225
R8258 VSS VSS.n1841 0.01225
R8259 VSS.n1750 VSS 0.01225
R8260 VSS VSS.n1746 0.01225
R8261 VSS.n1746 VSS 0.01225
R8262 VSS.n1688 VSS 0.01225
R8263 VSS VSS.n1684 0.01225
R8264 VSS.n1684 VSS 0.01225
R8265 VSS VSS.n1734 0.01225
R8266 VSS.n1739 VSS 0.01225
R8267 VSS.n1739 VSS 0.01225
R8268 VSS.n1820 VSS 0.01225
R8269 VSS.n1823 VSS 0.01225
R8270 VSS.n1823 VSS 0.01225
R8271 VSS.n1833 VSS 0.01225
R8272 VSS VSS.n1829 0.01225
R8273 VSS.n1829 VSS 0.01225
R8274 VSS.n1423 VSS 0.01225
R8275 VSS VSS.n1419 0.01225
R8276 VSS.n1419 VSS 0.01225
R8277 VSS.n1430 VSS 0.01225
R8278 VSS.n1433 VSS 0.01225
R8279 VSS.n1433 VSS 0.01225
R8280 VSS.n1803 VSS 0.01225
R8281 VSS.n1801 VSS 0.01225
R8282 VSS.n1801 VSS 0.01225
R8283 VSS VSS.n1448 0.01225
R8284 VSS.n1453 VSS 0.01225
R8285 VSS.n1453 VSS 0.01225
R8286 VSS VSS.n1438 0.01225
R8287 VSS.n1443 VSS 0.01225
R8288 VSS.n1443 VSS 0.01225
R8289 VSS.n1790 VSS 0.01225
R8290 VSS.n1793 VSS 0.01225
R8291 VSS.n1793 VSS 0.01225
R8292 VSS.n1678 VSS 0.01225
R8293 VSS VSS.n1674 0.01225
R8294 VSS.n1674 VSS 0.01225
R8295 VSS.n4431 VSS.n4418 0.0119583
R8296 VSS.n4506 VSS.n4503 0.0119583
R8297 VSS.n4551 VSS.n4533 0.0119583
R8298 VSS.n5011 VSS.n5008 0.0119583
R8299 VSS.n2194 VSS.n2183 0.0114881
R8300 VSS.n353 VSS.n352 0.0114223
R8301 VSS.n4850 VSS.n4849 0.0114072
R8302 VSS.n4398 VSS.n4397 0.0114072
R8303 VSS.n4380 VSS.n4379 0.0114072
R8304 VSS.n4186 VSS.n4185 0.0114072
R8305 VSS.n5038 VSS.n5037 0.0114072
R8306 VSS.n2442 VSS.n2441 0.0114072
R8307 VSS.n3622 VSS.n3621 0.0113921
R8308 VSS.n3525 VSS.n3524 0.0113921
R8309 VSS.n3428 VSS.n3427 0.0113921
R8310 VSS.n3331 VSS.n3330 0.0113921
R8311 VSS.n5468 VSS.n5467 0.0113921
R8312 VSS.n5820 VSS.n5817 0.0113921
R8313 VSS.n6658 VSS.n6657 0.0113921
R8314 VSS.n1099 VSS.n1098 0.0113921
R8315 VSS.n1133 VSS.n1132 0.0113921
R8316 VSS.n6425 VSS.n6423 0.0113921
R8317 VSS.n1218 VSS.n1217 0.0113921
R8318 VSS.n967 VSS.n966 0.0113921
R8319 VSS.n6130 VSS.n6129 0.0113921
R8320 VSS.n5 VSS.n4 0.0113921
R8321 VSS.n6644 VSS.n6642 0.0112192
R8322 VSS.n1862 VSS 0.0105121
R8323 VSS VSS.n1183 0.0105121
R8324 VSS.n1342 VSS 0.0105121
R8325 VSS.n6360 VSS 0.0105121
R8326 VSS.n1324 VSS 0.0105121
R8327 VSS VSS.n1192 0.0105121
R8328 VSS VSS.n1193 0.0105121
R8329 VSS VSS.n1462 0.0105121
R8330 VSS VSS.n1587 0.0105121
R8331 VSS VSS.n1663 0.0105121
R8332 VSS VSS.n1694 0.0105121
R8333 VSS VSS.n1707 0.0105121
R8334 VSS VSS.n1728 0.0105121
R8335 VSS VSS.n1595 0.0105121
R8336 VSS VSS.n1757 0.0105121
R8337 VSS VSS.n1580 0.0105121
R8338 VSS VSS.n1771 0.0105121
R8339 VSS VSS.n1810 0.0105121
R8340 VSS VSS.n1778 0.0105121
R8341 VSS VSS.n1472 0.0105121
R8342 VSS VSS.n1412 0.0105121
R8343 VSS VSS.n1528 0.0105121
R8344 VSS VSS.n1749 0.0105121
R8345 VSS VSS.n1714 0.0105121
R8346 VSS VSS.n1687 0.0105121
R8347 VSS VSS.n1737 0.0105121
R8348 VSS VSS.n1819 0.0105121
R8349 VSS VSS.n1832 0.0105121
R8350 VSS VSS.n1422 0.0105121
R8351 VSS VSS.n1429 0.0105121
R8352 VSS VSS.n1799 0.0105121
R8353 VSS VSS.n1451 0.0105121
R8354 VSS VSS.n1441 0.0105121
R8355 VSS VSS.n1789 0.0105121
R8356 VSS VSS.n1677 0.0105121
R8357 VSS.n1465 VSS.n1464 0.01037
R8358 VSS.n1590 VSS.n1589 0.01037
R8359 VSS.n1710 VSS.n1702 0.01037
R8360 VSS.n1710 VSS.n1709 0.01037
R8361 VSS.n1725 VSS.n1724 0.01037
R8362 VSS.n1609 VSS.n1608 0.01037
R8363 VSS.n1767 VSS.n1766 0.01037
R8364 VSS.n1475 VSS.n1474 0.01037
R8365 VSS.n1839 VSS.n1530 0.01037
R8366 VSS.n1840 VSS.n1839 0.01037
R8367 VSS.n1762 VSS.n1761 0.01037
R8368 VSS.n1752 VSS.n1751 0.01037
R8369 VSS.n1720 VSS.n1719 0.01037
R8370 VSS.n1690 VSS.n1689 0.01037
R8371 VSS.n1700 VSS.n1699 0.01037
R8372 VSS.n1742 VSS.n1740 0.01037
R8373 VSS.n1742 VSS.n1741 0.01037
R8374 VSS.n1825 VSS.n1824 0.01037
R8375 VSS.n1835 VSS.n1827 0.01037
R8376 VSS.n1835 VSS.n1834 0.01037
R8377 VSS.n1425 VSS.n1424 0.01037
R8378 VSS.n1435 VSS.n1434 0.01037
R8379 VSS.n1815 VSS.n1814 0.01037
R8380 VSS.n1805 VSS.n1804 0.01037
R8381 VSS.n1455 VSS.n1454 0.01037
R8382 VSS.n1445 VSS.n1444 0.01037
R8383 VSS.n1785 VSS.n1783 0.01037
R8384 VSS.n1785 VSS.n1784 0.01037
R8385 VSS.n1795 VSS.n1794 0.01037
R8386 VSS.n1600 VSS.n1599 0.01037
R8387 VSS.n1670 VSS.n1669 0.01037
R8388 VSS.n1680 VSS.n1679 0.01037
R8389 VSS.n1849 VSS.n1848 0.01037
R8390 VSS.n365 VSS.n362 0.0100354
R8391 VSS VSS.n1459 0.0100119
R8392 VSS VSS.n1460 0.0100119
R8393 VSS VSS.n1586 0.0100119
R8394 VSS VSS.n1582 0.0100119
R8395 VSS VSS.n1665 0.0100119
R8396 VSS VSS.n1667 0.0100119
R8397 VSS VSS.n1696 0.0100119
R8398 VSS VSS.n1697 0.0100119
R8399 VSS VSS.n7511 0.0100119
R8400 VSS VSS.n573 0.0100119
R8401 VSS VSS.n473 0.0100119
R8402 VSS VSS.n7298 0.0100119
R8403 VSS VSS.n273 0.0100119
R8404 VSS VSS.n1716 0.0100119
R8405 VSS VSS.n1717 0.0100119
R8406 VSS VSS.n1706 0.0100119
R8407 VSS VSS.n1703 0.0100119
R8408 VSS.n7551 VSS 0.0100119
R8409 VSS VSS.n231 0.0100119
R8410 VSS.n1729 VSS 0.0100119
R8411 VSS VSS.n1726 0.0100119
R8412 VSS VSS.n1597 0.0100119
R8413 VSS VSS.n1592 0.0100119
R8414 VSS VSS.n1759 0.0100119
R8415 VSS VSS.n1754 0.0100119
R8416 VSS VSS.n1606 0.0100119
R8417 VSS VSS.n1602 0.0100119
R8418 VSS.n1772 VSS 0.0100119
R8419 VSS VSS.n1768 0.0100119
R8420 VSS VSS.n1812 0.0100119
R8421 VSS VSS.n1807 0.0100119
R8422 VSS VSS.n1780 0.0100119
R8423 VSS VSS.n1781 0.0100119
R8424 VSS VSS.n1471 0.0100119
R8425 VSS VSS.n1467 0.0100119
R8426 VSS VSS.n1414 0.0100119
R8427 VSS.n1851 VSS 0.0100119
R8428 VSS VSS.n1527 0.0100119
R8429 VSS.n1842 VSS 0.0100119
R8430 VSS VSS.n1748 0.0100119
R8431 VSS VSS.n1744 0.0100119
R8432 VSS VSS.n1686 0.0100119
R8433 VSS VSS.n1682 0.0100119
R8434 VSS VSS.n1736 0.0100119
R8435 VSS VSS.n1738 0.0100119
R8436 VSS VSS.n1818 0.0100119
R8437 VSS VSS.n1822 0.0100119
R8438 VSS VSS.n1831 0.0100119
R8439 VSS VSS.n1828 0.0100119
R8440 VSS VSS.n1421 0.0100119
R8441 VSS VSS.n1417 0.0100119
R8442 VSS VSS.n1428 0.0100119
R8443 VSS VSS.n1432 0.0100119
R8444 VSS VSS.n1798 0.0100119
R8445 VSS VSS.n1800 0.0100119
R8446 VSS VSS.n1450 0.0100119
R8447 VSS VSS.n1452 0.0100119
R8448 VSS VSS.n1440 0.0100119
R8449 VSS VSS.n1442 0.0100119
R8450 VSS VSS.n1788 0.0100119
R8451 VSS VSS.n1792 0.0100119
R8452 VSS VSS.n1676 0.0100119
R8453 VSS VSS.n1672 0.0100119
R8454 VSS.n2669 VSS.n2668 0.00946062
R8455 VSS.n2683 VSS.n2682 0.00946062
R8456 VSS.n1617 VSS.n1616 0.00946062
R8457 VSS.n1552 VSS.n1551 0.00946062
R8458 VSS.n1483 VSS.n1482 0.00946062
R8459 VSS.n1376 VSS.n1375 0.00946062
R8460 VSS.n2649 VSS.n2645 0.00946026
R8461 VSS.n2638 VSS.n2635 0.00946026
R8462 VSS.n1656 VSS.n1652 0.00946026
R8463 VSS.n1539 VSS.n1535 0.00946026
R8464 VSS.n1404 VSS.n1403 0.00946026
R8465 VSS.n1501 VSS.n1500 0.00946026
R8466 VSS.n2699 VSS.n2698 0.00922857
R8467 VSS.n1259 VSS.n1258 0.00897165
R8468 VSS.n2703 VSS.n2702 0.00896
R8469 VSS.n2638 VSS.n2637 0.00896
R8470 VSS.n2649 VSS.n2648 0.00896
R8471 VSS.n2670 VSS.n2669 0.00896
R8472 VSS.n2684 VSS.n2683 0.00896
R8473 VSS.n2695 VSS.n2694 0.00896
R8474 VSS.n1656 VSS.n1655 0.00896
R8475 VSS.n1539 VSS.n1538 0.00896
R8476 VSS.n1501 VSS.n1499 0.00896
R8477 VSS.n291 VSS.n288 0.00896
R8478 VSS.n1618 VSS.n1617 0.00896
R8479 VSS.n1553 VSS.n1552 0.00896
R8480 VSS.n1484 VSS.n1483 0.00896
R8481 VSS.n1377 VSS.n1376 0.00896
R8482 VSS.n1404 VSS.n1402 0.00896
R8483 VSS.n6396 VSS.n1174 0.00883333
R8484 VSS.n6698 VSS.n6697 0.0083125
R8485 VSS.n2743 VSS.n2742 0.0083125
R8486 VSS.n6572 VSS.n1106 0.00810719
R8487 VSS.n979 VSS.n978 0.0079343
R8488 VSS.n3514 VSS.n3513 0.00779167
R8489 VSS.n7512 VSS 0.0076315
R8490 VSS.n7516 VSS 0.0076315
R8491 VSS VSS.n7516 0.0076315
R8492 VSS.n574 VSS 0.0076315
R8493 VSS.n578 VSS 0.0076315
R8494 VSS VSS.n578 0.0076315
R8495 VSS.n474 VSS 0.0076315
R8496 VSS.n478 VSS 0.0076315
R8497 VSS VSS.n478 0.0076315
R8498 VSS.n7299 VSS 0.0076315
R8499 VSS.n7303 VSS 0.0076315
R8500 VSS VSS.n7303 0.0076315
R8501 VSS.n274 VSS 0.0076315
R8502 VSS.n278 VSS 0.0076315
R8503 VSS VSS.n278 0.0076315
R8504 VSS.n110 VSS 0.0076315
R8505 VSS.n7555 VSS 0.0076315
R8506 VSS VSS.n7555 0.0076315
R8507 VSS.n232 VSS 0.0076315
R8508 VSS.n236 VSS 0.0076315
R8509 VSS VSS.n236 0.0076315
R8510 VSS.n4855 VSS.n4854 0.00742521
R8511 VSS.n5634 VSS.n2502 0.007315
R8512 VSS.n2764 VSS.n2709 0.007315
R8513 VSS.n5467 VSS.n5466 0.00727101
R8514 VSS.n4855 VSS.n4852 0.00638643
R8515 VSS.n5658 VSS.n5656 0.00622917
R8516 VSS.n3475 VSS.n2904 0.00622917
R8517 VSS.n2633 VSS.n2632 0.00610795
R8518 VSS.n2633 VSS 0.00610795
R8519 VSS.n2640 VSS 0.00610795
R8520 VSS.n2640 VSS 0.00610795
R8521 VSS.n2651 VSS.n2643 0.00610795
R8522 VSS.n2651 VSS 0.00610795
R8523 VSS.n2646 VSS 0.00610795
R8524 VSS VSS.n2646 0.00610795
R8525 VSS.n2666 VSS.n2665 0.00610795
R8526 VSS.n2666 VSS 0.00610795
R8527 VSS.n2673 VSS 0.00610795
R8528 VSS.n2673 VSS 0.00610795
R8529 VSS.n2680 VSS.n2679 0.00610795
R8530 VSS.n2680 VSS 0.00610795
R8531 VSS.n2687 VSS 0.00610795
R8532 VSS.n2687 VSS 0.00610795
R8533 VSS.n1658 VSS.n1650 0.00610795
R8534 VSS.n1658 VSS 0.00610795
R8535 VSS.n1653 VSS 0.00610795
R8536 VSS VSS.n1653 0.00610795
R8537 VSS.n1541 VSS.n1533 0.00610795
R8538 VSS.n1541 VSS 0.00610795
R8539 VSS.n1536 VSS 0.00610795
R8540 VSS VSS.n1536 0.00610795
R8541 VSS.n1406 VSS.n1398 0.00610795
R8542 VSS.n1406 VSS 0.00610795
R8543 VSS.n1400 VSS 0.00610795
R8544 VSS VSS.n1400 0.00610795
R8545 VSS.n1503 VSS.n1495 0.00610795
R8546 VSS.n1503 VSS 0.00610795
R8547 VSS.n1497 VSS 0.00610795
R8548 VSS VSS.n1497 0.00610795
R8549 VSS.n1613 VSS.n1612 0.00610795
R8550 VSS.n1613 VSS 0.00610795
R8551 VSS.n1620 VSS 0.00610795
R8552 VSS.n1620 VSS 0.00610795
R8553 VSS.n1548 VSS.n1547 0.00610795
R8554 VSS.n1548 VSS 0.00610795
R8555 VSS.n1555 VSS 0.00610795
R8556 VSS.n1555 VSS 0.00610795
R8557 VSS.n1479 VSS.n1478 0.00610795
R8558 VSS.n1479 VSS 0.00610795
R8559 VSS.n1486 VSS 0.00610795
R8560 VSS.n1486 VSS 0.00610795
R8561 VSS.n1372 VSS.n1371 0.00610795
R8562 VSS.n1372 VSS 0.00610795
R8563 VSS.n1379 VSS 0.00610795
R8564 VSS.n1379 VSS 0.00610795
R8565 VSS.n5820 VSS.n5819 0.00585961
R8566 VSS.n978 VSS.n977 0.00585961
R8567 VSS.n6573 VSS.n6572 0.00568672
R8568 VSS VSS.n1212 0.00563311
R8569 VSS.n2369 VSS.n2368 0.00557629
R8570 VSS.n2364 VSS.n2363 0.00557629
R8571 VSS.n1325 VSS 0.0054727
R8572 VSS.n1355 VSS 0.0054727
R8573 VSS VSS.n6094 0.00531229
R8574 VSS.n1202 VSS 0.00531229
R8575 VSS VSS.n1337 0.00531229
R8576 VSS VSS.n1856 0.00531229
R8577 VSS.n6352 VSS 0.00531229
R8578 VSS.n2708 VSS.n2701 0.00526062
R8579 VSS.n1743 VSS.n1742 0.00523021
R8580 VSS.n1826 VSS.n1825 0.00523021
R8581 VSS.n1466 VSS.n1465 0.00523021
R8582 VSS.n1786 VSS.n1785 0.00523021
R8583 VSS.n1601 VSS.n1600 0.00523021
R8584 VSS.n1766 VSS.n1765 0.00523021
R8585 VSS.n1671 VSS.n1670 0.00523021
R8586 VSS.n1862 VSS.n1859 0.00523021
R8587 VSS.n1352 VSS.n1183 0.00523021
R8588 VSS.n1342 VSS.n1332 0.00523021
R8589 VSS.n6361 VSS.n6360 0.00523021
R8590 VSS.n1324 VSS.n1207 0.00523021
R8591 VSS.n1199 VSS.n1192 0.00523021
R8592 VSS.n6097 VSS.n1193 0.00523021
R8593 VSS.n1591 VSS.n1590 0.00523013
R8594 VSS.n1701 VSS.n1700 0.00523013
R8595 VSS.n1711 VSS.n1710 0.00523013
R8596 VSS.n1721 VSS.n1720 0.00523013
R8597 VSS.n1724 VSS.n1723 0.00523013
R8598 VSS.n1610 VSS.n1609 0.00523013
R8599 VSS.n1816 VSS.n1815 0.00523013
R8600 VSS.n1476 VSS.n1475 0.00523013
R8601 VSS.n1848 VSS.n1847 0.00523013
R8602 VSS.n1839 VSS.n1838 0.00523013
R8603 VSS.n1753 VSS.n1752 0.00523013
R8604 VSS.n1763 VSS.n1762 0.00523013
R8605 VSS.n1691 VSS.n1690 0.00523013
R8606 VSS.n1836 VSS.n1835 0.00523013
R8607 VSS.n1436 VSS.n1435 0.00523013
R8608 VSS.n1426 VSS.n1425 0.00523013
R8609 VSS.n1806 VSS.n1805 0.00523013
R8610 VSS.n1446 VSS.n1445 0.00523013
R8611 VSS.n1456 VSS.n1455 0.00523013
R8612 VSS.n1796 VSS.n1795 0.00523013
R8613 VSS.n1681 VSS.n1680 0.00523013
R8614 VSS.n6332 VSS.n6331 0.0052
R8615 VSS.n6331 VSS.n1864 0.0050825
R8616 VSS.n1259 VSS.n1256 0.00482227
R8617 VSS.n2701 VSS.n2700 0.00476029
R8618 VSS.n6091 VSS.n6090 0.00476028
R8619 VSS.n2692 VSS.n2631 0.00476028
R8620 VSS.n2678 VSS.n2642 0.00476028
R8621 VSS.n2664 VSS.n2653 0.00476028
R8622 VSS.n2660 VSS.n2659 0.00476028
R8623 VSS.n2664 VSS.n2663 0.00476028
R8624 VSS.n2678 VSS.n2677 0.00476028
R8625 VSS.n2692 VSS.n2691 0.00476028
R8626 VSS.n114 VSS.n113 0.00476028
R8627 VSS.n118 VSS.n117 0.00476028
R8628 VSS.n258 VSS.n242 0.00476028
R8629 VSS.n283 VSS.n282 0.00476028
R8630 VSS.n125 VSS.n124 0.00476028
R8631 VSS.n241 VSS.n240 0.00476028
R8632 VSS.n7550 VSS.n128 0.00476028
R8633 VSS.n1733 VSS.n1649 0.00476028
R8634 VSS.n1776 VSS.n1531 0.00476028
R8635 VSS.n1845 VSS.n1844 0.00476028
R8636 VSS.n287 VSS.n286 0.00476028
R8637 VSS.n7549 VSS.n7548 0.00476028
R8638 VSS.n7550 VSS.n292 0.00476028
R8639 VSS.n1733 VSS.n1625 0.00476028
R8640 VSS.n1776 VSS.n1560 0.00476028
R8641 VSS.n1845 VSS.n1491 0.00476028
R8642 VSS.n1853 VSS.n1386 0.00476028
R8643 VSS.n6358 VSS.n6355 0.00476028
R8644 VSS.n1182 VSS.n1179 0.00476028
R8645 VSS.n1361 VSS.n1358 0.00476028
R8646 VSS.n1187 VSS.n1184 0.00476028
R8647 VSS.n1331 VSS.n1328 0.00476028
R8648 VSS.n1191 VSS.n1188 0.00476028
R8649 VSS.n1206 VSS.n1205 0.00476028
R8650 VSS.n1853 VSS.n1410 0.00476028
R8651 VSS.n2675 VSS.n2664 0.00473
R8652 VSS.n2689 VSS.n2678 0.00473
R8653 VSS.n2676 VSS.n2675 0.00473
R8654 VSS.n2701 VSS.n2692 0.00473
R8655 VSS.n2690 VSS.n2689 0.00473
R8656 VSS.n576 VSS.n112 0.00473
R8657 VSS.n476 VSS.n284 0.00473
R8658 VSS.n276 VSS.n116 0.00473
R8659 VSS.n7301 VSS.n120 0.00473
R8660 VSS.n7550 VSS.n283 0.00473
R8661 VSS.n7550 VSS.n258 0.00473
R8662 VSS.n7553 VSS.n7552 0.00473
R8663 VSS.n234 VSS.n122 0.00473
R8664 VSS.n7550 VSS.n241 0.00473
R8665 VSS.n1776 VSS.n1775 0.00473
R8666 VSS.n1845 VSS.n1506 0.00473
R8667 VSS.n1776 VSS.n1544 0.00473
R8668 VSS.n1733 VSS.n1732 0.00473
R8669 VSS.n1733 VSS.n1647 0.00473
R8670 VSS.n7550 VSS.n125 0.00473
R8671 VSS.n1722 VSS.n1647 0.00473
R8672 VSS.n1733 VSS.n1639 0.00473
R8673 VSS.n7550 VSS.n118 0.00473
R8674 VSS.n1733 VSS.n1637 0.00473
R8675 VSS.n1764 VSS.n1577 0.00473
R8676 VSS.n1733 VSS.n1634 0.00473
R8677 VSS.n1776 VSS.n1570 0.00473
R8678 VSS.n1776 VSS.n1573 0.00473
R8679 VSS.n1845 VSS.n1508 0.00473
R8680 VSS.n1845 VSS.n1515 0.00473
R8681 VSS.n1846 VSS.n1393 0.00473
R8682 VSS.n1776 VSS.n1577 0.00473
R8683 VSS.n1837 VSS.n1515 0.00473
R8684 VSS.n1845 VSS.n1523 0.00473
R8685 VSS.n1845 VSS.n1493 0.00473
R8686 VSS.n1845 VSS.n1518 0.00473
R8687 VSS.n1776 VSS.n1566 0.00473
R8688 VSS.n1776 VSS.n1562 0.00473
R8689 VSS.n1733 VSS.n1627 0.00473
R8690 VSS.n1733 VSS.n1644 0.00473
R8691 VSS.n7550 VSS.n114 0.00473
R8692 VSS.n7550 VSS.n287 0.00473
R8693 VSS.n7514 VSS.n293 0.00473
R8694 VSS.n7550 VSS.n7549 0.00473
R8695 VSS.n1733 VSS.n1622 0.00473
R8696 VSS.n1776 VSS.n1557 0.00473
R8697 VSS.n1845 VSS.n1488 0.00473
R8698 VSS.n1853 VSS.n1381 0.00473
R8699 VSS.n6359 VSS.n6358 0.00473
R8700 VSS.n1853 VSS.n1384 0.00473
R8701 VSS.n6359 VSS.n1182 0.00473
R8702 VSS.n1853 VSS.n1389 0.00473
R8703 VSS.n6359 VSS.n1361 0.00473
R8704 VSS.n1853 VSS.n1368 0.00473
R8705 VSS.n6359 VSS.n1187 0.00473
R8706 VSS.n1853 VSS.n1393 0.00473
R8707 VSS.n6359 VSS.n1331 0.00473
R8708 VSS.n1853 VSS.n1364 0.00473
R8709 VSS.n6359 VSS.n1191 0.00473
R8710 VSS.n1853 VSS.n1397 0.00473
R8711 VSS.n6359 VSS.n1206 0.00473
R8712 VSS.n1845 VSS.n1511 0.00473
R8713 VSS.n1853 VSS.n1409 0.00473
R8714 VSS.n2705 VSS.n2702 0.00426062
R8715 VSS.n2696 VSS.n2695 0.00426062
R8716 VSS.n289 VSS.n288 0.00426062
R8717 VSS.n2471 VSS.n2470 0.00414583
R8718 VSS.n6836 VSS.n6834 0.00414583
R8719 VSS.n6178 VSS.n6177 0.00414583
R8720 VSS.n2655 VSS.n2654 0.00390244
R8721 VSS.n365 VSS.n364 0.00379404
R8722 VSS.n3817 VSS.n3816 0.00378492
R8723 VSS.n3720 VSS.n3719 0.00378492
R8724 VSS.n2362 VSS.n2361 0.00335545
R8725 VSS.n2367 VSS.n2366 0.00335545
R8726 VSS.n2366 VSS.n2365 0.00334133
R8727 VSS.n2361 VSS.n2360 0.00334133
R8728 VSS.n1863 VSS.n1178 0.00327702
R8729 VSS.n2661 VSS.n2660 0.00306417
R8730 VSS.n6330 VSS.n6326 0.00298917
R8731 VSS.n2224 VSS.n2223 0.00296757
R8732 VSS.n2223 VSS.n2222 0.00296757
R8733 VSS.n2662 VSS.n2661 0.00295776
R8734 VSS.n6351 VSS.n1863 0.00290614
R8735 VSS.n2675 VSS.n2652 0.00288062
R8736 VSS.n2675 VSS.n2674 0.00288062
R8737 VSS.n2689 VSS.n2641 0.00288031
R8738 VSS.n2689 VSS.n2688 0.00288031
R8739 VSS.n1732 VSS.n1659 0.00288031
R8740 VSS.n1544 VSS.n1542 0.00288031
R8741 VSS.n1409 VSS.n1407 0.00288031
R8742 VSS.n1506 VSS.n1504 0.00288031
R8743 VSS.n1622 VSS.n1621 0.00288031
R8744 VSS.n1557 VSS.n1556 0.00288031
R8745 VSS.n1488 VSS.n1487 0.00288031
R8746 VSS.n1381 VSS.n1380 0.00288031
R8747 VSS.n1384 VSS.n1383 0.00288014
R8748 VSS.n1562 VSS.n1561 0.00288014
R8749 VSS.n1733 VSS.n1628 0.00288014
R8750 VSS.n7550 VSS.n285 0.00288014
R8751 VSS.n7550 VSS.n115 0.00288014
R8752 VSS.n7550 VSS.n119 0.00288014
R8753 VSS.n7550 VSS.n259 0.00288014
R8754 VSS.n1634 VSS.n1633 0.00288014
R8755 VSS.n7550 VSS.n121 0.00288014
R8756 VSS.n7550 VSS.n126 0.00288014
R8757 VSS.n1732 VSS.n1731 0.00288014
R8758 VSS.n1733 VSS.n1648 0.00288014
R8759 VSS.n1776 VSS.n1545 0.00288014
R8760 VSS.n1776 VSS.n1563 0.00288014
R8761 VSS.n1577 VSS.n1576 0.00288014
R8762 VSS.n1775 VSS.n1774 0.00288014
R8763 VSS.n1776 VSS.n1567 0.00288014
R8764 VSS.n1776 VSS.n1579 0.00288014
R8765 VSS.n1845 VSS.n1494 0.00288014
R8766 VSS.n1853 VSS.n1395 0.00288014
R8767 VSS.n1397 VSS.n1396 0.00288014
R8768 VSS.n1845 VSS.n1525 0.00288014
R8769 VSS.n1506 VSS.n1505 0.00288014
R8770 VSS.n1544 VSS.n1543 0.00288014
R8771 VSS.n1573 VSS.n1572 0.00288014
R8772 VSS.n1647 VSS.n1646 0.00288014
R8773 VSS.n1639 VSS.n1638 0.00288014
R8774 VSS.n1733 VSS.n1642 0.00288014
R8775 VSS.n1733 VSS.n1640 0.00288014
R8776 VSS.n1637 VSS.n1636 0.00288014
R8777 VSS.n1733 VSS.n1631 0.00288014
R8778 VSS.n1733 VSS.n1635 0.00288014
R8779 VSS.n1570 VSS.n1569 0.00288014
R8780 VSS.n1776 VSS.n1575 0.00288014
R8781 VSS.n1776 VSS.n1571 0.00288014
R8782 VSS.n1511 VSS.n1510 0.00288014
R8783 VSS.n1508 VSS.n1507 0.00288014
R8784 VSS.n1845 VSS.n1513 0.00288014
R8785 VSS.n1845 VSS.n1509 0.00288014
R8786 VSS.n1853 VSS.n1365 0.00288014
R8787 VSS.n1364 VSS.n1363 0.00288014
R8788 VSS.n1853 VSS.n1391 0.00288014
R8789 VSS.n1393 VSS.n1392 0.00288014
R8790 VSS.n1515 VSS.n1514 0.00288014
R8791 VSS.n1523 VSS.n1522 0.00288014
R8792 VSS.n1845 VSS.n1519 0.00288014
R8793 VSS.n1845 VSS.n1521 0.00288014
R8794 VSS.n1853 VSS.n1369 0.00288014
R8795 VSS.n1368 VSS.n1367 0.00288014
R8796 VSS.n1853 VSS.n1387 0.00288014
R8797 VSS.n1389 VSS.n1388 0.00288014
R8798 VSS.n1518 VSS.n1517 0.00288014
R8799 VSS.n1493 VSS.n1492 0.00288014
R8800 VSS.n1566 VSS.n1565 0.00288014
R8801 VSS.n1644 VSS.n1643 0.00288014
R8802 VSS.n1627 VSS.n1626 0.00288014
R8803 VSS.n7550 VSS.n294 0.00288014
R8804 VSS.n1733 VSS.n1623 0.00288014
R8805 VSS.n1776 VSS.n1558 0.00288014
R8806 VSS.n1845 VSS.n1489 0.00288014
R8807 VSS.n1853 VSS.n1382 0.00288014
R8808 VSS.n1409 VSS.n1408 0.00288014
R8809 VSS.n1853 VSS.n1411 0.00288014
R8810 VSS.n3281 VSS.n3280 0.00258771
R8811 VSS.n6020 VSS.n1949 0.00258771
R8812 VSS.n1991 VSS.n1971 0.00258771
R8813 VSS.n1908 VSS.n1907 0.00258771
R8814 VSS.n3330 VSS.n3329 0.00258351
R8815 VSS.n6645 VSS.n6644 0.00257469
R8816 VSS.n2359 VSS.n2358 0.00253147
R8817 VSS.n2234 VSS.n2233 0.00253147
R8818 VSS.n2234 VSS.n2110 0.00250667
R8819 VSS.n2359 VSS.n2239 0.00250667
R8820 VSS.n4880 VSS.n4879 0.00239617
R8821 VSS.n7321 VSS.n7320 0.00239617
R8822 VSS.n2639 VSS.n2638 0.00238
R8823 VSS.n2650 VSS.n2649 0.00238
R8824 VSS.n2669 VSS.n2667 0.00238
R8825 VSS.n2683 VSS.n2681 0.00238
R8826 VSS.n1657 VSS.n1656 0.00238
R8827 VSS.n1540 VSS.n1539 0.00238
R8828 VSS.n1405 VSS.n1404 0.00238
R8829 VSS.n1502 VSS.n1501 0.00238
R8830 VSS.n1617 VSS.n1614 0.00238
R8831 VSS.n1552 VSS.n1549 0.00238
R8832 VSS.n1483 VSS.n1480 0.00238
R8833 VSS.n1376 VSS.n1373 0.00238
R8834 VSS.n4511 VSS.n4487 0.00225009
R8835 VSS.n4573 VSS.n4572 0.00225009
R8836 VSS.n5016 VSS.n4992 0.00225009
R8837 VSS.n4774 VSS.n4773 0.00225009
R8838 VSS.n5662 VSS.n5661 0.00225009
R8839 VSS.n5091 VSS.n5090 0.00225009
R8840 VSS.n596 VSS.n595 0.00225009
R8841 VSS.n7536 VSS.n7535 0.00225009
R8842 VSS.n498 VSS.n497 0.00225009
R8843 VSS.n386 VSS.n385 0.00225009
R8844 VSS.n220 VSS.n218 0.00225009
R8845 VSS.n7575 VSS.n7574 0.00225009
R8846 VSS.n7517 VSS 0.00213006
R8847 VSS.n7304 VSS 0.00213006
R8848 VSS.n279 VSS 0.00213006
R8849 VSS.n7556 VSS 0.00213006
R8850 VSS.n237 VSS 0.00213006
R8851 VSS.n163 VSS.n162 0.00206853
R8852 VSS.n3574 VSS.n3572 0.0020625
R8853 VSS.n579 VSS 0.00206214
R8854 VSS.n6330 VSS.n6329 0.00201061
R8855 VSS.n7287 VSS.n7285 0.00200697
R8856 VSS.n7292 VSS.n7291 0.00200697
R8857 VSS.n7580 VSS.n7578 0.00200697
R8858 VSS.n100 VSS.n98 0.00200697
R8859 VSS.n105 VSS.n104 0.00200697
R8860 VSS.n199 VSS.n198 0.00200697
R8861 VSS.n4786 VSS.n4785 0.00200697
R8862 VSS.n4454 VSS.n4359 0.00200697
R8863 VSS.n4484 VSS.n4483 0.00200697
R8864 VSS.n4405 VSS.n4361 0.00200697
R8865 VSS.n4409 VSS.n4369 0.00200697
R8866 VSS.n4986 VSS.n4984 0.00200697
R8867 VSS.n4578 VSS.n4576 0.00200697
R8868 VSS.n4494 VSS.n4492 0.00200697
R8869 VSS.n4499 VSS.n4498 0.00200697
R8870 VSS.n4613 VSS.n4610 0.00200697
R8871 VSS.n3881 VSS.n3880 0.00200697
R8872 VSS.n5274 VSS.n5273 0.00200697
R8873 VSS.n4300 VSS.n3893 0.00200697
R8874 VSS.n5270 VSS.n3897 0.00200697
R8875 VSS.n4349 VSS.n4348 0.00200697
R8876 VSS.n4288 VSS.n4287 0.00200697
R8877 VSS.n4345 VSS.n4293 0.00200697
R8878 VSS.n4338 VSS.n4337 0.00200697
R8879 VSS.n4268 VSS.n4262 0.00200697
R8880 VSS.n4657 VSS.n4656 0.00200697
R8881 VSS.n4624 VSS.n4364 0.00200697
R8882 VSS.n4959 VSS.n4203 0.00200697
R8883 VSS.n4373 VSS.n4200 0.00200697
R8884 VSS.n4964 VSS.n4963 0.00200697
R8885 VSS.n4480 VSS.n4478 0.00200697
R8886 VSS.n4864 VSS.n4862 0.00200697
R8887 VSS.n4869 VSS.n4868 0.00200697
R8888 VSS.n5096 VSS.n5094 0.00200697
R8889 VSS.n4143 VSS.n4141 0.00200697
R8890 VSS.n4148 VSS.n4147 0.00200697
R8891 VSS.n5667 VSS.n5665 0.00200697
R8892 VSS.n4886 VSS.n4884 0.00200697
R8893 VSS.n4761 VSS.n4759 0.00200697
R8894 VSS.n4766 VSS.n4765 0.00200697
R8895 VSS.n4928 VSS.n4927 0.00200697
R8896 VSS.n4839 VSS.n4749 0.00200697
R8897 VSS.n4917 VSS.n4844 0.00200697
R8898 VSS.n5160 VSS.n5159 0.00200697
R8899 VSS.n4913 VSS.n4120 0.00200697
R8900 VSS.n5147 VSS.n5146 0.00200697
R8901 VSS.n5134 VSS.n5128 0.00200697
R8902 VSS.n4835 VSS.n4834 0.00200697
R8903 VSS.n4830 VSS.n4820 0.00200697
R8904 VSS.n4815 VSS.n4814 0.00200697
R8905 VSS.n4675 VSS.n4238 0.00200697
R8906 VSS.n4246 VSS.n4237 0.00200697
R8907 VSS.n4696 VSS.n4231 0.00200697
R8908 VSS.n4228 VSS.n4227 0.00200697
R8909 VSS.n4730 VSS.n4729 0.00200697
R8910 VSS.n4711 VSS.n4705 0.00200697
R8911 VSS.n5209 VSS.n5208 0.00200697
R8912 VSS.n5196 VSS.n5190 0.00200697
R8913 VSS.n4251 VSS.n4242 0.00200697
R8914 VSS.n4257 VSS.n4256 0.00200697
R8915 VSS.n4264 VSS.n4245 0.00200697
R8916 VSS.n4039 VSS.n4030 0.00200697
R8917 VSS.n4016 VSS.n4015 0.00200697
R8918 VSS.n4025 VSS.n4012 0.00200697
R8919 VSS.n4052 VSS.n4008 0.00200697
R8920 VSS.n4021 VSS.n3997 0.00200697
R8921 VSS.n4003 VSS.n3994 0.00200697
R8922 VSS.n4064 VSS.n3990 0.00200697
R8923 VSS.n3999 VSS.n3989 0.00200697
R8924 VSS.n4091 VSS.n3983 0.00200697
R8925 VSS.n4071 VSS.n3944 0.00200697
R8926 VSS.n3973 VSS.n3972 0.00200697
R8927 VSS.n3960 VSS.n3954 0.00200697
R8928 VSS.n5256 VSS.n3906 0.00200697
R8929 VSS.n3904 VSS.n3899 0.00200697
R8930 VSS.n4296 VSS.n3901 0.00200697
R8931 VSS.n3780 VSS.n3778 0.00200697
R8932 VSS.n3785 VSS.n3784 0.00200697
R8933 VSS.n3694 VSS.n3692 0.00200697
R8934 VSS.n3682 VSS.n3680 0.00200697
R8935 VSS.n3687 VSS.n3686 0.00200697
R8936 VSS.n3596 VSS.n3594 0.00200697
R8937 VSS.n3584 VSS.n3582 0.00200697
R8938 VSS.n3589 VSS.n3588 0.00200697
R8939 VSS.n3499 VSS.n3497 0.00200697
R8940 VSS.n3487 VSS.n3485 0.00200697
R8941 VSS.n3492 VSS.n3491 0.00200697
R8942 VSS.n3402 VSS.n3400 0.00200697
R8943 VSS.n3390 VSS.n3388 0.00200697
R8944 VSS.n3395 VSS.n3394 0.00200697
R8945 VSS.n5340 VSS.n5338 0.00200697
R8946 VSS.n2828 VSS.n2826 0.00200697
R8947 VSS.n5443 VSS.n5442 0.00200697
R8948 VSS.n3792 VSS.n3791 0.00200697
R8949 VSS.n3798 VSS.n3797 0.00200697
R8950 VSS.n5433 VSS.n5431 0.00200697
R8951 VSS.n5437 VSS.n5436 0.00200697
R8952 VSS.n5773 VSS.n5772 0.00200697
R8953 VSS.n3956 VSS.n2387 0.00200697
R8954 VSS.n5741 VSS.n5740 0.00200697
R8955 VSS.n5192 VSS.n2406 0.00200697
R8956 VSS.n5709 VSS.n5708 0.00200697
R8957 VSS.n5130 VSS.n2425 0.00200697
R8958 VSS.n2460 VSS.n2458 0.00200697
R8959 VSS.n2465 VSS.n2464 0.00200697
R8960 VSS.n2534 VSS.n2529 0.00200697
R8961 VSS.n2580 VSS.n2563 0.00200697
R8962 VSS.n2559 VSS.n2554 0.00200697
R8963 VSS.n2542 VSS.n2531 0.00200697
R8964 VSS.n2613 VSS.n2612 0.00200697
R8965 VSS.n5620 VSS.n5619 0.00200697
R8966 VSS.n398 VSS.n397 0.00200697
R8967 VSS.n2735 VSS.n2734 0.00200697
R8968 VSS.n7460 VSS.n7459 0.00200697
R8969 VSS.n646 VSS.n316 0.00200697
R8970 VSS.n502 VSS.n501 0.00200697
R8971 VSS.n601 VSS.n599 0.00200697
R8972 VSS.n7499 VSS.n7497 0.00200697
R8973 VSS.n7504 VSS.n7503 0.00200697
R8974 VSS.n633 VSS.n632 0.00200697
R8975 VSS.n676 VSS.n675 0.00200697
R8976 VSS.n663 VSS.n662 0.00200697
R8977 VSS.n6666 VSS.n789 0.00200697
R8978 VSS.n823 VSS.n791 0.00200697
R8979 VSS.n779 VSS.n761 0.00200697
R8980 VSS.n759 VSS.n757 0.00200697
R8981 VSS.n7196 VSS.n7195 0.00200697
R8982 VSS.n7092 VSS.n7082 0.00200697
R8983 VSS.n7192 VSS.n7086 0.00200697
R8984 VSS.n639 VSS.n630 0.00200697
R8985 VSS.n7487 VSS.n7485 0.00200697
R8986 VSS.n508 VSS.n507 0.00200697
R8987 VSS.n7327 VSS.n7325 0.00200697
R8988 VSS.n373 VSS.n371 0.00200697
R8989 VSS.n378 VSS.n377 0.00200697
R8990 VSS.n7416 VSS.n7415 0.00200697
R8991 VSS.n693 VSS.n343 0.00200697
R8992 VSS.n7260 VSS.n698 0.00200697
R8993 VSS.n7359 VSS.n7357 0.00200697
R8994 VSS.n7356 VSS.n7355 0.00200697
R8995 VSS.n7377 VSS.n7376 0.00200697
R8996 VSS.n87 VSS.n85 0.00200697
R8997 VSS.n689 VSS.n688 0.00200697
R8998 VSS.n684 VSS.n429 0.00200697
R8999 VSS.n434 VSS.n426 0.00200697
R9000 VSS.n7122 VSS.n7113 0.00200697
R9001 VSS.n7110 VSS.n7109 0.00200697
R9002 VSS.n7161 VSS.n7160 0.00200697
R9003 VSS.n7137 VSS.n7135 0.00200697
R9004 VSS.n7245 VSS.n721 0.00200697
R9005 VSS.n7144 VSS.n719 0.00200697
R9006 VSS.n6924 VSS.n6923 0.00200697
R9007 VSS.n6911 VSS.n6905 0.00200697
R9008 VSS.n7178 VSS.n7104 0.00200697
R9009 VSS.n7102 VSS.n7088 0.00200697
R9010 VSS.n7097 VSS.n7090 0.00200697
R9011 VSS.n7025 VSS.n7024 0.00200697
R9012 VSS.n844 VSS.n810 0.00200697
R9013 VSS.n887 VSS.n849 0.00200697
R9014 VSS.n900 VSS.n897 0.00200697
R9015 VSS.n892 VSS.n885 0.00200697
R9016 VSS.n905 VSS.n904 0.00200697
R9017 VSS.n6999 VSS.n6998 0.00200697
R9018 VSS.n910 VSS.n875 0.00200697
R9019 VSS.n6868 VSS.n915 0.00200697
R9020 VSS.n6883 VSS.n6880 0.00200697
R9021 VSS.n6872 VSS.n6866 0.00200697
R9022 VSS.n6968 VSS.n6967 0.00200697
R9023 VSS.n6955 VSS.n6949 0.00200697
R9024 VSS.n840 VSS.n839 0.00200697
R9025 VSS.n835 VSS.n832 0.00200697
R9026 VSS.n827 VSS.n821 0.00200697
R9027 VSS.n1085 VSS.n1084 0.00200697
R9028 VSS.n1079 VSS.n1077 0.00200697
R9029 VSS.n6559 VSS.n6557 0.00200697
R9030 VSS.n1119 VSS.n1118 0.00200697
R9031 VSS.n1113 VSS.n1111 0.00200697
R9032 VSS.n6492 VSS.n6490 0.00200697
R9033 VSS.n6480 VSS.n6478 0.00200697
R9034 VSS.n6485 VSS.n6484 0.00200697
R9035 VSS.n6406 VSS.n6404 0.00200697
R9036 VSS.n1170 VSS.n1169 0.00200697
R9037 VSS.n1164 VSS.n1162 0.00200697
R9038 VSS.n1282 VSS.n1280 0.00200697
R9039 VSS.n1270 VSS.n1268 0.00200697
R9040 VSS.n1275 VSS.n1274 0.00200697
R9041 VSS.n6851 VSS.n6850 0.00200697
R9042 VSS.n953 VSS.n952 0.00200697
R9043 VSS.n6157 VSS.n6156 0.00200697
R9044 VSS.n6153 VSS.n6151 0.00200697
R9045 VSS.n1072 VSS.n1071 0.00200697
R9046 VSS.n1068 VSS.n1066 0.00200697
R9047 VSS.n6170 VSS.n6169 0.00200697
R9048 VSS.n6164 VSS.n6162 0.00200697
R9049 VSS.n7717 VSS.n7716 0.00200697
R9050 VSS.n6951 VSS.n30 0.00200697
R9051 VSS.n7685 VSS.n7684 0.00200697
R9052 VSS.n6907 VSS.n49 0.00200697
R9053 VSS.n7653 VSS.n7652 0.00200697
R9054 VSS.n81 VSS.n68 0.00200697
R9055 VSS.n177 VSS.n175 0.00200697
R9056 VSS.n182 VSS.n181 0.00200697
R9057 VSS.n145 VSS.n144 0.00200683
R9058 VSS.n7649 VSS.n7648 0.00200683
R9059 VSS.n7681 VSS.n7680 0.00200683
R9060 VSS.n7713 VSS.n7712 0.00200683
R9061 VSS.n2485 VSS.n2484 0.00200683
R9062 VSS.n5705 VSS.n5704 0.00200683
R9063 VSS.n5737 VSS.n5736 0.00200683
R9064 VSS.n5769 VSS.n5768 0.00200683
R9065 VSS.n4778 VSS.n4777 0.00200683
R9066 VSS.n5000 VSS.n4999 0.00200683
R9067 VSS.n4447 VSS.n4446 0.00200683
R9068 VSS.n4989 VSS.n4988 0.00200683
R9069 VSS.n4541 VSS.n4540 0.00200683
R9070 VSS.n4605 VSS.n4370 0.00200683
R9071 VSS.n4617 VSS.n4365 0.00200683
R9072 VSS.n4317 VSS.n4284 0.00200683
R9073 VSS.n4628 VSS.n4355 0.00200683
R9074 VSS.n5156 VSS.n5155 0.00200683
R9075 VSS.n5143 VSS.n5142 0.00200683
R9076 VSS.n4689 VSS.n4688 0.00200683
R9077 VSS.n4740 VSS.n4739 0.00200683
R9078 VSS.n4726 VSS.n4725 0.00200683
R9079 VSS.n5205 VSS.n5204 0.00200683
R9080 VSS.n4084 VSS.n4083 0.00200683
R9081 VSS.n3978 VSS.n3942 0.00200683
R9082 VSS.n3969 VSS.n3968 0.00200683
R9083 VSS.n5449 VSS.n5448 0.00200683
R9084 VSS.n5801 VSS.n5800 0.00200683
R9085 VSS.n2628 VSS.n2627 0.00200683
R9086 VSS.n2598 VSS.n2527 0.00200683
R9087 VSS.n2568 VSS.n2552 0.00200683
R9088 VSS.n390 VSS.n389 0.00200683
R9089 VSS.n463 VSS.n462 0.00200683
R9090 VSS.n7490 VSS.n7489 0.00200683
R9091 VSS.n562 VSS.n561 0.00200683
R9092 VSS.n529 VSS.n528 0.00200683
R9093 VSS.n659 VSS.n658 0.00200683
R9094 VSS.n7045 VSS.n7044 0.00200683
R9095 VSS.n7072 VSS.n7071 0.00200683
R9096 VSS.n7063 VSS.n7062 0.00200683
R9097 VSS.n7456 VSS.n7455 0.00200683
R9098 VSS.n765 VSS.n313 0.00200683
R9099 VSS.n2730 VSS.n2729 0.00200683
R9100 VSS.n7373 VSS.n7372 0.00200683
R9101 VSS.n7618 VSS.n7617 0.00200683
R9102 VSS.n7171 VSS.n7170 0.00200683
R9103 VSS.n7157 VSS.n7156 0.00200683
R9104 VSS.n6893 VSS.n717 0.00200683
R9105 VSS.n6920 VSS.n6919 0.00200683
R9106 VSS.n6875 VSS.n6864 0.00200683
R9107 VSS.n6964 VSS.n6963 0.00200683
R9108 VSS.n6691 VSS.n6690 0.00200683
R9109 VSS.n7745 VSS.n7744 0.00200683
R9110 VSS.n5004 VSS.n5003 0.00200677
R9111 VSS.n4545 VSS.n4544 0.00200677
R9112 VSS.n467 VSS.n466 0.00200677
R9113 VSS.n6683 VSS.n6682 0.00200674
R9114 VSS.n2201 VSS.n2200 0.002
R9115 VSS.n6089 VSS.n1 0.00199514
R9116 VSS.n479 VSS 0.00199422
R9117 VSS.n4510 VSS.n4509 0.00192045
R9118 VSS.n4548 VSS.n4377 0.00192045
R9119 VSS.n5015 VSS.n5014 0.00192045
R9120 VSS.n4769 VSS.n4750 0.00192045
R9121 VSS.n2468 VSS.n2439 0.00192045
R9122 VSS.n4151 VSS.n4136 0.00192045
R9123 VSS.n4879 VSS.n4878 0.00192045
R9124 VSS.n593 VSS.n592 0.00192045
R9125 VSS.n7533 VSS.n7532 0.00192045
R9126 VSS.n495 VSS.n494 0.00192045
R9127 VSS.n381 VSS.n344 0.00192045
R9128 VSS.n222 VSS.n221 0.00192045
R9129 VSS.n7572 VSS.n7571 0.00192045
R9130 VSS.n7320 VSS.n7319 0.00192045
R9131 VSS.n2256 VSS.n2255 0.00178939
R9132 VSS.n4330 VSS.n4327 0.00175017
R9133 VSS.n4641 VSS.n4638 0.00175017
R9134 VSS.n4950 VSS.n4210 0.00175017
R9135 VSS.n5179 VSS.n5174 0.00175017
R9136 VSS.n4220 VSS.n4216 0.00175017
R9137 VSS.n4940 VSS.n4938 0.00175017
R9138 VSS.n5221 VSS.n3936 0.00175017
R9139 VSS.n5240 VSS.n3919 0.00175017
R9140 VSS.n5250 VSS.n3916 0.00175017
R9141 VSS.n5331 VSS.n5326 0.00175017
R9142 VSS.n2843 VSS.n2840 0.00175017
R9143 VSS.n5314 VSS.n2845 0.00175017
R9144 VSS.n5305 VSS.n2849 0.00175017
R9145 VSS.n5296 VSS.n2853 0.00175017
R9146 VSS.n5287 VSS.n2857 0.00175017
R9147 VSS.n2623 VSS.n2516 0.00175017
R9148 VSS.n2591 VSS.n2541 0.00175017
R9149 VSS.n7204 VSS.n745 0.00175017
R9150 VSS.n7445 VSS.n326 0.00175017
R9151 VSS.n7436 VSS.n328 0.00175017
R9152 VSS.n7389 VSS.n711 0.00175017
R9153 VSS.n7395 VSS.n336 0.00175017
R9154 VSS.n7428 VSS.n7426 0.00175017
R9155 VSS.n6938 VSS.n6933 0.00175017
R9156 VSS.n735 VSS.n732 0.00175017
R9157 VSS.n7222 VSS.n737 0.00175017
R9158 VSS.n7213 VSS.n741 0.00175017
R9159 VSS.n6980 VSS.n936 0.00175017
R9160 VSS.n6985 VSS.n931 0.00175017
R9161 VSS.n926 VSS.n868 0.00175017
R9162 VSS.n7011 VSS.n865 0.00175017
R9163 VSS.n860 VSS.n803 0.00175017
R9164 VSS.n6673 VSS.n801 0.00175017
R9165 VSS.n1873 VSS.n1872 0.00173379
R9166 VSS.n1872 VSS.n1871 0.00173379
R9167 VSS.n6325 VSS.n6324 0.00152605
R9168 VSS.n6331 VSS.n6325 0.00151551
R9169 VSS.n2367 VSS.n2234 0.00150431
R9170 VSS.n2362 VSS.n2359 0.00150431
R9171 VSS.n2211 VSS.n2210 0.0015
R9172 VSS.n2230 VSS.n2220 0.0015
R9173 VSS.n5261 VSS.n3905 0.00149521
R9174 VSS.n661 VSS.n627 0.00149521
R9175 VSS.n7183 VSS.n7103 0.00149521
R9176 VSS.n838 VSS.n812 0.00149521
R9177 VSS.n7289 VSS.n7288 0.00149516
R9178 VSS.n7585 VSS.n7581 0.00149516
R9179 VSS.n102 VSS.n101 0.00149516
R9180 VSS.n197 VSS.n193 0.00149516
R9181 VSS.n4783 VSS.n4782 0.00149516
R9182 VSS.n4987 VSS.n4191 0.00149516
R9183 VSS.n4496 VSS.n4495 0.00149516
R9184 VSS.n4583 VSS.n4579 0.00149516
R9185 VSS.n4614 VSS.n4609 0.00149516
R9186 VSS.n3879 VSS.n2864 0.00149516
R9187 VSS.n5272 VSS.n3887 0.00149516
R9188 VSS.n5271 VSS.n3896 0.00149516
R9189 VSS.n5272 VSS.n3889 0.00149516
R9190 VSS.n4346 VSS.n4292 0.00149516
R9191 VSS.n4336 VSS.n4261 0.00149516
R9192 VSS.n4655 VSS.n4258 0.00149516
R9193 VSS.n4648 VSS.n4261 0.00149516
R9194 VSS.n4625 VSS.n4363 0.00149516
R9195 VSS.n4961 VSS.n4960 0.00149516
R9196 VSS.n4962 VSS.n4197 0.00149516
R9197 VSS.n4482 VSS.n4402 0.00149516
R9198 VSS.n4445 VSS.n4415 0.00149516
R9199 VSS.n4866 VSS.n4865 0.00149516
R9200 VSS.n5101 VSS.n5097 0.00149516
R9201 VSS.n4145 VSS.n4144 0.00149516
R9202 VSS.n5672 VSS.n5668 0.00149516
R9203 VSS.n4763 VSS.n4762 0.00149516
R9204 VSS.n4891 VSS.n4887 0.00149516
R9205 VSS.n4926 VSS.n4746 0.00149516
R9206 VSS.n4925 VSS.n4846 0.00149516
R9207 VSS.n5158 VSS.n4117 0.00149516
R9208 VSS.n5145 VSS.n4126 0.00149516
R9209 VSS.n4832 VSS.n4831 0.00149516
R9210 VSS.n4833 VSS.n4808 0.00149516
R9211 VSS.n4677 VSS.n4676 0.00149516
R9212 VSS.n4742 VSS.n4697 0.00149516
R9213 VSS.n4728 VSS.n4702 0.00149516
R9214 VSS.n4728 VSS.n4704 0.00149516
R9215 VSS.n5207 VSS.n4101 0.00149516
R9216 VSS.n5207 VSS.n4103 0.00149516
R9217 VSS.n4665 VSS.n4664 0.00149516
R9218 VSS.n4665 VSS.n4244 0.00149516
R9219 VSS.n4666 VSS.n4239 0.00149516
R9220 VSS.n4041 VSS.n4040 0.00149516
R9221 VSS.n4042 VSS.n4009 0.00149516
R9222 VSS.n4054 VSS.n4053 0.00149516
R9223 VSS.n4055 VSS.n3991 0.00149516
R9224 VSS.n4066 VSS.n4065 0.00149516
R9225 VSS.n4066 VSS.n3988 0.00149516
R9226 VSS.n4093 VSS.n4092 0.00149516
R9227 VSS.n4093 VSS.n3943 0.00149516
R9228 VSS.n3971 VSS.n3945 0.00149516
R9229 VSS.n3971 VSS.n3947 0.00149516
R9230 VSS.n5263 VSS.n5262 0.00149516
R9231 VSS.n5262 VSS.n3900 0.00149516
R9232 VSS.n5261 VSS.n3908 0.00149516
R9233 VSS.n3782 VSS.n3781 0.00149516
R9234 VSS.n3699 VSS.n3695 0.00149516
R9235 VSS.n3684 VSS.n3683 0.00149516
R9236 VSS.n3601 VSS.n3597 0.00149516
R9237 VSS.n3586 VSS.n3585 0.00149516
R9238 VSS.n3504 VSS.n3500 0.00149516
R9239 VSS.n3489 VSS.n3488 0.00149516
R9240 VSS.n3407 VSS.n3403 0.00149516
R9241 VSS.n3392 VSS.n3391 0.00149516
R9242 VSS.n5345 VSS.n5341 0.00149516
R9243 VSS.n2829 VSS.n2824 0.00149516
R9244 VSS.n2829 VSS.n2820 0.00149516
R9245 VSS.n3795 VSS.n3794 0.00149516
R9246 VSS.n3879 VSS.n3875 0.00149516
R9247 VSS.n5435 VSS.n5434 0.00149516
R9248 VSS.n5435 VSS.n5427 0.00149516
R9249 VSS.n5771 VSS.n2384 0.00149516
R9250 VSS.n5771 VSS.n2386 0.00149516
R9251 VSS.n5739 VSS.n2403 0.00149516
R9252 VSS.n5739 VSS.n2405 0.00149516
R9253 VSS.n5707 VSS.n2422 0.00149516
R9254 VSS.n5707 VSS.n2424 0.00149516
R9255 VSS.n2462 VSS.n2461 0.00149516
R9256 VSS.n2582 VSS.n2581 0.00149516
R9257 VSS.n2582 VSS.n2553 0.00149516
R9258 VSS.n2603 VSS.n2530 0.00149516
R9259 VSS.n2604 VSS.n2523 0.00149516
R9260 VSS.n2611 VSS.n2510 0.00149516
R9261 VSS.n5621 VSS.n2510 0.00149516
R9262 VSS.n395 VSS.n394 0.00149516
R9263 VSS.n7501 VSS.n7500 0.00149516
R9264 VSS.n606 VSS.n602 0.00149516
R9265 VSS.n631 VSS.n533 0.00149516
R9266 VSS.n677 VSS.n431 0.00149516
R9267 VSS.n7047 VSS.n788 0.00149516
R9268 VSS.n7047 VSS.n785 0.00149516
R9269 VSS.n7194 VSS.n752 0.00149516
R9270 VSS.n7193 VSS.n7085 0.00149516
R9271 VSS.n7194 VSS.n754 0.00149516
R9272 VSS.n661 VSS.n629 0.00149516
R9273 VSS.n660 VSS.n643 0.00149516
R9274 VSS.n7488 VSS.n304 0.00149516
R9275 VSS.n505 VSS.n503 0.00149516
R9276 VSS.n375 VSS.n374 0.00149516
R9277 VSS.n7332 VSS.n7328 0.00149516
R9278 VSS.n7414 VSS.n340 0.00149516
R9279 VSS.n7413 VSS.n700 0.00149516
R9280 VSS.n7361 VSS.n7360 0.00149516
R9281 VSS.n7375 VSS.n86 0.00149516
R9282 VSS.n686 VSS.n685 0.00149516
R9283 VSS.n687 VSS.n420 0.00149516
R9284 VSS.n7173 VSS.n7123 0.00149516
R9285 VSS.n7159 VSS.n7132 0.00149516
R9286 VSS.n7247 VSS.n7246 0.00149516
R9287 VSS.n7247 VSS.n718 0.00149516
R9288 VSS.n6922 VSS.n6896 0.00149516
R9289 VSS.n6922 VSS.n6898 0.00149516
R9290 VSS.n7185 VSS.n7184 0.00149516
R9291 VSS.n7184 VSS.n7089 0.00149516
R9292 VSS.n7183 VSS.n7106 0.00149516
R9293 VSS.n7023 VSS.n807 0.00149516
R9294 VSS.n7022 VSS.n851 0.00149516
R9295 VSS.n902 VSS.n901 0.00149516
R9296 VSS.n903 VSS.n879 0.00149516
R9297 VSS.n6997 VSS.n872 0.00149516
R9298 VSS.n6996 VSS.n917 0.00149516
R9299 VSS.n6885 VSS.n6884 0.00149516
R9300 VSS.n6885 VSS.n6865 0.00149516
R9301 VSS.n6966 VSS.n6856 0.00149516
R9302 VSS.n6966 VSS.n6858 0.00149516
R9303 VSS.n837 VSS.n836 0.00149516
R9304 VSS.n837 VSS.n820 0.00149516
R9305 VSS.n838 VSS.n815 0.00149516
R9306 VSS.n1082 VSS.n1081 0.00149516
R9307 VSS.n6564 VSS.n6560 0.00149516
R9308 VSS.n1116 VSS.n1115 0.00149516
R9309 VSS.n6497 VSS.n6493 0.00149516
R9310 VSS.n6482 VSS.n6481 0.00149516
R9311 VSS.n6411 VSS.n6407 0.00149516
R9312 VSS.n1167 VSS.n1166 0.00149516
R9313 VSS.n1287 VSS.n1283 0.00149516
R9314 VSS.n1272 VSS.n1271 0.00149516
R9315 VSS.n6849 VSS.n6845 0.00149516
R9316 VSS.n950 VSS.n949 0.00149516
R9317 VSS.n6154 VSS.n6148 0.00149516
R9318 VSS.n1069 VSS.n1064 0.00149516
R9319 VSS.n6167 VSS.n6166 0.00149516
R9320 VSS.n6167 VSS.n6145 0.00149516
R9321 VSS.n7715 VSS.n27 0.00149516
R9322 VSS.n7715 VSS.n29 0.00149516
R9323 VSS.n7683 VSS.n46 0.00149516
R9324 VSS.n7683 VSS.n48 0.00149516
R9325 VSS.n7651 VSS.n65 0.00149516
R9326 VSS.n7651 VSS.n67 0.00149516
R9327 VSS.n179 VSS.n178 0.00149516
R9328 VSS.n7289 VSS.n7281 0.00149516
R9329 VSS.n7585 VSS.n92 0.00149516
R9330 VSS.n102 VSS.n94 0.00149516
R9331 VSS.n197 VSS.n186 0.00149516
R9332 VSS.n4626 VSS.n4357 0.00149516
R9333 VSS.n4482 VSS.n4401 0.00149516
R9334 VSS.n4615 VSS.n4367 0.00149516
R9335 VSS.n4583 VSS.n4376 0.00149516
R9336 VSS.n4496 VSS.n4488 0.00149516
R9337 VSS.n4347 VSS.n4281 0.00149516
R9338 VSS.n4961 VSS.n4199 0.00149516
R9339 VSS.n4962 VSS.n4194 0.00149516
R9340 VSS.n4866 VSS.n4858 0.00149516
R9341 VSS.n5101 VSS.n4134 0.00149516
R9342 VSS.n4145 VSS.n4137 0.00149516
R9343 VSS.n5672 VSS.n2438 0.00149516
R9344 VSS.n4891 VSS.n4847 0.00149516
R9345 VSS.n4763 VSS.n4755 0.00149516
R9346 VSS.n4926 VSS.n4748 0.00149516
R9347 VSS.n4925 VSS.n4843 0.00149516
R9348 VSS.n5158 VSS.n4119 0.00149516
R9349 VSS.n5157 VSS.n4122 0.00149516
R9350 VSS.n5144 VSS.n5127 0.00149516
R9351 VSS.n5145 VSS.n4128 0.00149516
R9352 VSS.n4833 VSS.n4805 0.00149516
R9353 VSS.n4832 VSS.n4813 0.00149516
R9354 VSS.n4677 VSS.n4236 0.00149516
R9355 VSS.n4680 VSS.n4233 0.00149516
R9356 VSS.n4743 VSS.n4742 0.00149516
R9357 VSS.n4741 VSS.n4698 0.00149516
R9358 VSS.n4727 VSS.n4715 0.00149516
R9359 VSS.n5206 VSS.n5189 0.00149516
R9360 VSS.n4666 VSS.n4241 0.00149516
R9361 VSS.n4041 VSS.n4014 0.00149516
R9362 VSS.n4042 VSS.n4011 0.00149516
R9363 VSS.n4054 VSS.n3996 0.00149516
R9364 VSS.n4055 VSS.n3993 0.00149516
R9365 VSS.n4075 VSS.n3985 0.00149516
R9366 VSS.n4094 VSS.n3938 0.00149516
R9367 VSS.n3970 VSS.n3953 0.00149516
R9368 VSS.n3782 VSS.n3774 0.00149516
R9369 VSS.n3699 VSS.n3674 0.00149516
R9370 VSS.n3684 VSS.n3676 0.00149516
R9371 VSS.n3601 VSS.n3576 0.00149516
R9372 VSS.n3586 VSS.n3578 0.00149516
R9373 VSS.n3504 VSS.n3479 0.00149516
R9374 VSS.n3489 VSS.n3481 0.00149516
R9375 VSS.n3407 VSS.n3382 0.00149516
R9376 VSS.n3392 VSS.n3384 0.00149516
R9377 VSS.n5345 VSS.n2819 0.00149516
R9378 VSS.n5447 VSS.n5424 0.00149516
R9379 VSS.n5799 VSS.n2371 0.00149516
R9380 VSS.n5770 VSS.n2389 0.00149516
R9381 VSS.n5738 VSS.n2408 0.00149516
R9382 VSS.n5706 VSS.n2427 0.00149516
R9383 VSS.n2462 VSS.n2454 0.00149516
R9384 VSS.n2486 VSS.n2476 0.00149516
R9385 VSS.n2603 VSS.n2528 0.00149516
R9386 VSS.n2583 VSS.n2548 0.00149516
R9387 VSS.n5611 VSS.n2629 0.00149516
R9388 VSS.n2732 VSS.n2723 0.00149516
R9389 VSS.n7458 VSS.n310 0.00149516
R9390 VSS.n7457 VSS.n315 0.00149516
R9391 VSS.n505 VSS.n437 0.00149516
R9392 VSS.n606 VSS.n535 0.00149516
R9393 VSS.n7501 VSS.n7493 0.00149516
R9394 VSS.n667 VSS.n533 0.00149516
R9395 VSS.n7046 VSS.n790 0.00149516
R9396 VSS.n778 VSS.n758 0.00149516
R9397 VSS.n7074 VSS.n7073 0.00149516
R9398 VSS.n563 VSS.n553 0.00149516
R9399 VSS.n7332 VSS.n7263 0.00149516
R9400 VSS.n375 VSS.n367 0.00149516
R9401 VSS.n7414 VSS.n342 0.00149516
R9402 VSS.n7413 VSS.n697 0.00149516
R9403 VSS.n7361 VSS.n7258 0.00149516
R9404 VSS.n7364 VSS.n7255 0.00149516
R9405 VSS.n7620 VSS.n7619 0.00149516
R9406 VSS.n7607 VSS.n86 0.00149516
R9407 VSS.n687 VSS.n417 0.00149516
R9408 VSS.n686 VSS.n425 0.00149516
R9409 VSS.n7174 VSS.n7173 0.00149516
R9410 VSS.n7172 VSS.n7124 0.00149516
R9411 VSS.n7159 VSS.n7134 0.00149516
R9412 VSS.n7158 VSS.n7141 0.00149516
R9413 VSS.n7248 VSS.n713 0.00149516
R9414 VSS.n6921 VSS.n6904 0.00149516
R9415 VSS.n7023 VSS.n809 0.00149516
R9416 VSS.n7022 VSS.n848 0.00149516
R9417 VSS.n902 VSS.n884 0.00149516
R9418 VSS.n903 VSS.n876 0.00149516
R9419 VSS.n6997 VSS.n874 0.00149516
R9420 VSS.n6996 VSS.n914 0.00149516
R9421 VSS.n6886 VSS.n6860 0.00149516
R9422 VSS.n6965 VSS.n6948 0.00149516
R9423 VSS.n1082 VSS.n1061 0.00149516
R9424 VSS.n6564 VSS.n6554 0.00149516
R9425 VSS.n1116 VSS.n1108 0.00149516
R9426 VSS.n6497 VSS.n6473 0.00149516
R9427 VSS.n6482 VSS.n6474 0.00149516
R9428 VSS.n6411 VSS.n6401 0.00149516
R9429 VSS.n1167 VSS.n1159 0.00149516
R9430 VSS.n1287 VSS.n1263 0.00149516
R9431 VSS.n1272 VSS.n1264 0.00149516
R9432 VSS.n6849 VSS.n939 0.00149516
R9433 VSS.n950 VSS.n942 0.00149516
R9434 VSS.n7743 VSS.n14 0.00149516
R9435 VSS.n7714 VSS.n32 0.00149516
R9436 VSS.n7682 VSS.n51 0.00149516
R9437 VSS.n7650 VSS.n70 0.00149516
R9438 VSS.n179 VSS.n171 0.00149516
R9439 VSS.n146 VSS.n136 0.00149516
R9440 VSS.n6309 VSS.n6308 0.00146193
R9441 VSS.n5631 VSS.n5630 0.00125069
R9442 VSS.n5598 VSS.n5597 0.00125069
R9443 VSS.n2571 VSS.n2565 0.0012504
R9444 VSS.n2113 VSS.n2112 0.00118497
R9445 VSS.n2112 VSS.n2111 0.00118497
R9446 VSS.n6134 VSS.n6133 0.00114286
R9447 VSS.n974 VSS.n970 0.00114286
R9448 VSS.n1225 VSS.n1221 0.00114286
R9449 VSS.n6431 VSS.n6429 0.00114286
R9450 VSS.n1136 VSS.n1130 0.00114286
R9451 VSS.n1103 VSS.n1096 0.00114286
R9452 VSS.n6654 VSS.n6652 0.00114286
R9453 VSS.n4162 VSS.n4158 0.00114286
R9454 VSS.n548 VSS.n546 0.00114286
R9455 VSS.n450 VSS.n448 0.00114286
R9456 VSS.n6629 VSS.n6628 0.00114286
R9457 VSS.n12 VSS.n8 0.00114286
R9458 VSS.n3568 VSS.n3567 0.00114281
R9459 VSS.n3471 VSS.n3470 0.00114281
R9460 VSS.n3374 VSS.n3373 0.00114281
R9461 VSS.n5358 VSS.n2812 0.00114281
R9462 VSS.n5417 VSS.n5416 0.00114281
R9463 VSS.n6341 VSS.n6337 0.00114266
R9464 VSS.n2752 VSS.n298 0.00114214
R9465 VSS.n5643 VSS.n5642 0.00114214
R9466 VSS.n247 VSS.n243 0.00114214
R9467 VSS.n7268 VSS.n7264 0.00114214
R9468 VSS.n208 VSS.n204 0.00114214
R9469 VSS.n133 VSS.n129 0.00114214
R9470 VSS.n3760 VSS.n3758 0.00114214
R9471 VSS.n3662 VSS.n3660 0.00114214
R9472 VSS.n3858 VSS.n3856 0.00114214
R9473 VSS.n2499 VSS.n2496 0.00106587
R9474 VSS.n7522 VSS.n7521 0.00106587
R9475 VSS.n360 VSS.n347 0.00106587
R9476 VSS.n484 VSS.n481 0.00106587
R9477 VSS.n7309 VSS.n7306 0.00106587
R9478 VSS.n7561 VSS.n7558 0.00106587
R9479 VSS.n1231 VSS.n1230 0.00106587
R9480 VSS.n6371 VSS.n6370 0.00106587
R9481 VSS.n1347 VSS.n1346 0.00106587
R9482 VSS.n2762 VSS.n2719 0.00106586
R9483 VSS.n359 VSS.n350 0.00106586
R9484 VSS.n7311 VSS.n7310 0.00106586
R9485 VSS.n7563 VSS.n7562 0.00106586
R9486 VSS.n6350 VSS.n6349 0.00106582
R9487 VSS.n2747 VSS.n2746 0.00106068
R9488 VSS.n4428 VSS.n4427 0.00106068
R9489 VSS.n6349 VSS.n6348 0.00106068
R9490 VSS.n2719 VSS.n2718 0.00106064
R9491 VSS.n350 VSS.n349 0.00106064
R9492 VSS.n7312 VSS.n7311 0.00106064
R9493 VSS.n7564 VSS.n7563 0.00106064
R9494 VSS.n7523 VSS.n7522 0.00106063
R9495 VSS.n347 VSS.n346 0.00106063
R9496 VSS.n481 VSS.n480 0.00106063
R9497 VSS.n7306 VSS.n7305 0.00106063
R9498 VSS.n7558 VSS.n7557 0.00106063
R9499 VSS.n1348 VSS.n1347 0.00106063
R9500 VSS.n1341 VSS.n1340 0.00106063
R9501 VSS.n6372 VSS.n6371 0.00106063
R9502 VSS.n1322 VSS.n1231 0.00106063
R9503 VSS.n6348 VSS.n6347 0.00104326
R9504 VSS.n4428 VSS.n4426 0.00104326
R9505 VSS.n2751 VSS.n2747 0.00104326
R9506 VSS.n2500 VSS.n2495 0.00104326
R9507 VSS.n3862 VSS.n3861 0.00104325
R9508 VSS.n3764 VSS.n3763 0.00104325
R9509 VSS.n3666 VSS.n3665 0.00104325
R9510 VSS.n5464 VSS.n5460 0.00104325
R9511 VSS.n3327 VSS.n3323 0.00104325
R9512 VSS.n3424 VSS.n3420 0.00104325
R9513 VSS.n3521 VSS.n3517 0.00104325
R9514 VSS.n3618 VSS.n3614 0.00104325
R9515 VSS.n3716 VSS.n3712 0.00104325
R9516 VSS.n3813 VSS.n3809 0.00104325
R9517 VSS.n5813 VSS.n5809 0.00104325
R9518 VSS.n7524 VSS.n7508 0.00104317
R9519 VSS.n6186 VSS.n6182 0.00104317
R9520 VSS.n6547 VSS.n1126 0.00104317
R9521 VSS.n6466 VSS.n1146 0.00104317
R9522 VSS.n6392 VSS.n6373 0.00104317
R9523 VSS.n1321 VSS.n1319 0.00104317
R9524 VSS.n6343 VSS.n6342 0.00104317
R9525 VSS.n5413 VSS.n5412 0.00104317
R9526 VSS.n3564 VSS.n3563 0.00104317
R9527 VSS.n3467 VSS.n3466 0.00104317
R9528 VSS.n3370 VSS.n3369 0.00104317
R9529 VSS.n5360 VSS.n5359 0.00104317
R9530 VSS.n2255 VSS.n2254 0.00103939
R9531 VSS.n2255 VSS.n2252 0.00103403
R9532 VSS.n4173 VSS.n4169 0.00103325
R9533 VSS.n4180 VSS.n4176 0.00103325
R9534 VSS.n4385 VSS.n4381 0.00103325
R9535 VSS.n4392 VSS.n4388 0.00103325
R9536 VSS.n2447 VSS.n2443 0.00103325
R9537 VSS.n584 VSS.n570 0.00103325
R9538 VSS.n4166 VSS.n4165 0.00103325
R9539 VSS.n2474 VSS.n2451 0.00103325
R9540 VSS.n5082 VSS.n4152 0.00103325
R9541 VSS.n4164 VSS.n4163 0.00103325
R9542 VSS.n4168 VSS.n4167 0.00103325
R9543 VSS.n4175 VSS.n4174 0.00103325
R9544 VSS.n4554 VSS.n4531 0.00103325
R9545 VSS.n4387 VSS.n4386 0.00103325
R9546 VSS.n585 VSS.n584 0.00103325
R9547 VSS.n271 VSS.n270 0.00103325
R9548 VSS.n229 VSS.n169 0.00103325
R9549 VSS.n229 VSS.n228 0.00103325
R9550 VSS.n6828 VSS.n6827 0.00103325
R9551 VSS.n2500 VSS.n2499 0.00103324
R9552 VSS.n2751 VSS.n2750 0.00103324
R9553 VSS.n4426 VSS.n4425 0.00103324
R9554 VSS.n6347 VSS.n6346 0.00103324
R9555 VSS.n5464 VSS.n5463 0.00103323
R9556 VSS.n3327 VSS.n3326 0.00103323
R9557 VSS.n3424 VSS.n3423 0.00103323
R9558 VSS.n3521 VSS.n3520 0.00103323
R9559 VSS.n3618 VSS.n3617 0.00103323
R9560 VSS.n3716 VSS.n3715 0.00103323
R9561 VSS.n3813 VSS.n3812 0.00103323
R9562 VSS.n5813 VSS.n5812 0.00103323
R9563 VSS.n300 VSS.n299 0.00103323
R9564 VSS.n249 VSS.n248 0.00103323
R9565 VSS.n7270 VSS.n7269 0.00103323
R9566 VSS.n135 VSS.n134 0.00103323
R9567 VSS.n3765 VSS.n3764 0.00103323
R9568 VSS.n3667 VSS.n3666 0.00103323
R9569 VSS.n3863 VSS.n3862 0.00103323
R9570 VSS.n4419 VSS.n4395 0.00103319
R9571 VSS.n4522 VSS.n4520 0.00103319
R9572 VSS.n4530 VSS.n4527 0.00103319
R9573 VSS.n4562 VSS.n4561 0.00103319
R9574 VSS.n4555 VSS.n4183 0.00103319
R9575 VSS.n5027 VSS.n5025 0.00103319
R9576 VSS.n5035 VSS.n5032 0.00103319
R9577 VSS.n5049 VSS.n5047 0.00103319
R9578 VSS.n5057 VSS.n5054 0.00103319
R9579 VSS.n5065 VSS.n5063 0.00103319
R9580 VSS.n5076 VSS.n5074 0.00103319
R9581 VSS.n5077 VSS.n2450 0.00103319
R9582 VSS.n5651 VSS.n5650 0.00103319
R9583 VSS.n5650 VSS.n5648 0.00103319
R9584 VSS.n5652 VSS.n2450 0.00103319
R9585 VSS.n5081 VSS.n5076 0.00103319
R9586 VSS.n5069 VSS.n5065 0.00103319
R9587 VSS.n5062 VSS.n5057 0.00103319
R9588 VSS.n5053 VSS.n5049 0.00103319
R9589 VSS.n5046 VSS.n5035 0.00103319
R9590 VSS.n5031 VSS.n5027 0.00103319
R9591 VSS.n5024 VSS.n4183 0.00103319
R9592 VSS.n4561 VSS.n4559 0.00103319
R9593 VSS.n4563 VSS.n4530 0.00103319
R9594 VSS.n4526 VSS.n4522 0.00103319
R9595 VSS.n4519 VSS.n4395 0.00103319
R9596 VSS.n583 VSS.n582 0.00103319
R9597 VSS.n582 VSS.n580 0.00103319
R9598 VSS.n272 VSS.n267 0.00103319
R9599 VSS.n267 VSS.n265 0.00103319
R9600 VSS.n230 VSS.n166 0.00103319
R9601 VSS.n166 VSS.n164 0.00103319
R9602 VSS.n6830 VSS.n6829 0.00103319
R9603 VSS.n7524 VSS.n7523 0.00103317
R9604 VSS.n1348 VSS.n1126 0.00103317
R9605 VSS.n1341 VSS.n1146 0.00103317
R9606 VSS.n6373 VSS.n6372 0.00103317
R9607 VSS.n1322 VSS.n1321 0.00103317
R9608 VSS.n6188 VSS.n6186 0.00103317
R9609 VSS.n7521 VSS.n7518 0.0010331
R9610 VSS.n4162 VSS.n4161 0.0010331
R9611 VSS.n546 VSS.n545 0.0010331
R9612 VSS.n448 VSS.n447 0.0010331
R9613 VSS.n1346 VSS.n1343 0.0010331
R9614 VSS.n6465 VSS.n6464 0.0010331
R9615 VSS.n6370 VSS.n6367 0.0010331
R9616 VSS.n1230 VSS.n1227 0.0010331
R9617 VSS.n6135 VSS.n6134 0.0010331
R9618 VSS.n974 VSS.n973 0.0010331
R9619 VSS.n1225 VSS.n1224 0.0010331
R9620 VSS.n6429 VSS.n6428 0.0010331
R9621 VSS.n1130 VSS.n1129 0.0010331
R9622 VSS.n1103 VSS.n1102 0.0010331
R9623 VSS.n6628 VSS.n6627 0.0010331
R9624 VSS.n6652 VSS.n6651 0.0010331
R9625 VSS.n12 VSS.n11 0.0010331
R9626 VSS.n3569 VSS.n3568 0.00103308
R9627 VSS.n3472 VSS.n3471 0.00103308
R9628 VSS.n3375 VSS.n3374 0.00103308
R9629 VSS.n5358 VSS.n5357 0.00103308
R9630 VSS.n5418 VSS.n5417 0.00103308
R9631 VSS.n6341 VSS.n6340 0.00103305
R9632 VSS.n5644 VSS.n5643 0.00103293
R9633 VSS.n7543 VSS.n298 0.00103293
R9634 VSS.n255 VSS.n247 0.00103293
R9635 VSS.n7273 VSS.n7268 0.00103293
R9636 VSS.n212 VSS.n208 0.00103293
R9637 VSS.n159 VSS.n133 0.00103293
R9638 VSS.n3856 VSS.n3855 0.00103293
R9639 VSS.n3758 VSS.n2870 0.00103293
R9640 VSS.n3660 VSS.n2879 0.00103293
R9641 VSS.n2367 VSS.n2107 0.00102396
R9642 VSS.n2362 VSS.n2236 0.00102396
R9643 VSS.n5472 VSS.n5471 0.00102352
R9644 VSS.n3335 VSS.n3334 0.00102352
R9645 VSS.n3432 VSS.n3431 0.00102352
R9646 VSS.n3529 VSS.n3528 0.00102352
R9647 VSS.n3626 VSS.n3625 0.00102352
R9648 VSS.n3724 VSS.n3723 0.00102352
R9649 VSS.n3821 VSS.n3820 0.00102352
R9650 VSS.n5823 VSS.n5822 0.00102352
R9651 VSS.n2755 VSS.n2754 0.00102352
R9652 VSS.n5072 VSS.n5071 0.00102352
R9653 VSS.n4421 VSS.n4420 0.00102352
R9654 VSS.n541 VSS.n540 0.00102352
R9655 VSS.n443 VSS.n442 0.00102352
R9656 VSS.n6125 VSS.n6124 0.00102352
R9657 VSS.n982 VSS.n981 0.00102352
R9658 VSS.n1254 VSS.n1253 0.00102352
R9659 VSS.n6509 VSS.n6508 0.00102352
R9660 VSS.n6576 VSS.n6575 0.00102352
R9661 VSS.n6633 VSS.n6632 0.00102352
R9662 VSS.n6647 VSS.n1058 0.00102352
R9663 VSS.n6701 VSS.n1037 0.00102352
R9664 VSS.n7755 VSS.n13 0.00102352
R9665 VSS.n2761 VSS.n2760 0.00102351
R9666 VSS.n486 VSS.n485 0.0010235
R9667 VSS.n6127 VSS.n6126 0.0010235
R9668 VSS.n6434 VSS.n6432 0.0010235
R9669 VSS.n6510 VSS.n1137 0.0010235
R9670 VSS.n6631 VSS.n6630 0.0010235
R9671 VSS.n2194 VSS.n2193 0.00101844
R9672 VSS.n3809 VSS.n2871 0.00101835
R9673 VSS.n3712 VSS.n2880 0.00101835
R9674 VSS.n3614 VSS.n2889 0.00101835
R9675 VSS.n3517 VSS.n2900 0.00101835
R9676 VSS.n3420 VSS.n2912 0.00101835
R9677 VSS.n3323 VSS.n3317 0.00101835
R9678 VSS.n5460 VSS.n5385 0.00101835
R9679 VSS.n5809 VSS.n2370 0.00101835
R9680 VSS.n4158 VSS.n4153 0.00101832
R9681 VSS.n548 VSS.n547 0.00101832
R9682 VSS.n450 VSS.n449 0.00101832
R9683 VSS.n6133 VSS.n6127 0.00101832
R9684 VSS.n970 VSS.n964 0.00101832
R9685 VSS.n1221 VSS.n1215 0.00101832
R9686 VSS.n6432 VSS.n6431 0.00101832
R9687 VSS.n1137 VSS.n1136 0.00101832
R9688 VSS.n1096 VSS.n1093 0.00101832
R9689 VSS.n6654 VSS.n6653 0.00101832
R9690 VSS.n6630 VSS.n6629 0.00101832
R9691 VSS.n8 VSS.n2 0.00101832
R9692 VSS.n487 VSS.n486 0.00101831
R9693 VSS.n2762 VSS.n2761 0.0010183
R9694 VSS.n2756 VSS.n2755 0.0010183
R9695 VSS.n5071 VSS.n5070 0.0010183
R9696 VSS.n540 VSS.n539 0.0010183
R9697 VSS.n442 VSS.n441 0.0010183
R9698 VSS.n6126 VSS.n6125 0.0010183
R9699 VSS.n983 VSS.n982 0.0010183
R9700 VSS.n1253 VSS.n1252 0.0010183
R9701 VSS.n6434 VSS.n6433 0.0010183
R9702 VSS.n6510 VSS.n6509 0.0010183
R9703 VSS.n6577 VSS.n6576 0.0010183
R9704 VSS.n1058 VSS.n1057 0.0010183
R9705 VSS.n6632 VSS.n6631 0.0010183
R9706 VSS.n6350 VSS.n1037 0.0010183
R9707 VSS.n6059 VSS.n13 0.0010183
R9708 VSS.n3822 VSS.n3821 0.0010183
R9709 VSS.n3725 VSS.n3724 0.0010183
R9710 VSS.n3627 VSS.n3626 0.0010183
R9711 VSS.n3530 VSS.n3529 0.0010183
R9712 VSS.n3433 VSS.n3432 0.0010183
R9713 VSS.n3336 VSS.n3335 0.0010183
R9714 VSS.n5473 VSS.n5472 0.0010183
R9715 VSS.n5824 VSS.n5823 0.0010183
R9716 VSS.n2771 VSS.n2766 0.00101562
R9717 VSS.n6620 VSS.n6618 0.00101562
R9718 VSS.n1050 VSS.n1045 0.00101562
R9719 VSS.n6525 VSS.n6523 0.00101562
R9720 VSS.n6543 VSS.n6541 0.00101562
R9721 VSS.n6193 VSS.n6088 0.00101562
R9722 VSS.n6115 VSS.n6110 0.00101562
R9723 VSS.n6819 VSS.n6817 0.00101562
R9724 VSS.n1315 VSS.n1313 0.00101562
R9725 VSS.n6388 VSS.n6386 0.00101562
R9726 VSS.n1870 VSS.n1865 0.00101218
R9727 VSS.n5060 VSS.n5058 0.0010119
R9728 VSS.n6331 VSS.n6330 0.00100876
R9729 VSS.n2869 VSS.n2868 0.00100763
R9730 VSS.n2910 VSS.n2909 0.00100763
R9731 VSS.n2105 VSS.n2104 0.00100763
R9732 VSS.n5392 VSS.n5391 0.00100763
R9733 VSS.n5383 VSS.n5382 0.00100763
R9734 VSS.n2808 VSS.n2807 0.00100763
R9735 VSS.n3315 VSS.n3314 0.00100763
R9736 VSS.n2919 VSS.n2918 0.00100763
R9737 VSS.n2907 VSS.n2906 0.00100763
R9738 VSS.n2898 VSS.n2897 0.00100763
R9739 VSS.n2896 VSS.n2895 0.00100763
R9740 VSS.n2887 VSS.n2886 0.00100763
R9741 VSS.n2885 VSS.n2884 0.00100763
R9742 VSS.n2878 VSS.n2877 0.00100763
R9743 VSS.n2876 VSS.n2875 0.00100763
R9744 VSS.n998 VSS.n997 0.00100763
R9745 VSS.n6592 VSS.n6591 0.00100763
R9746 VSS.n6620 VSS.n6619 0.00100763
R9747 VSS.n1050 VSS.n1049 0.00100763
R9748 VSS.n3851 VSS.n3850 0.00100763
R9749 VSS.n6525 VSS.n6524 0.00100763
R9750 VSS.n6543 VSS.n6542 0.00100763
R9751 VSS.n6074 VSS.n6073 0.00100763
R9752 VSS.n6193 VSS.n6192 0.00100763
R9753 VSS.n6115 VSS.n6114 0.00100763
R9754 VSS.n6819 VSS.n6818 0.00100763
R9755 VSS.n1315 VSS.n1314 0.00100763
R9756 VSS.n1245 VSS.n1244 0.00100763
R9757 VSS.n6388 VSS.n6387 0.00100763
R9758 VSS.n6442 VSS.n6441 0.00100763
R9759 VSS.n6458 VSS.n6457 0.00100763
R9760 VSS.n5583 VSS.n5579 0.00100763
R9761 VSS.n6320 VSS.n6319 0.00100757
R9762 VSS.n4172 VSS.n4170 0.00100756
R9763 VSS.n4179 VSS.n4177 0.00100756
R9764 VSS.n4384 VSS.n4382 0.00100756
R9765 VSS.n4391 VSS.n4389 0.00100756
R9766 VSS.n2446 VSS.n2444 0.00100756
R9767 VSS.n2772 VSS.n2771 0.00100756
R9768 VSS.n7287 VSS.n7286 0.001007
R9769 VSS.n7291 VSS.n7290 0.001007
R9770 VSS.n7580 VSS.n7579 0.001007
R9771 VSS.n100 VSS.n99 0.001007
R9772 VSS.n104 VSS.n103 0.001007
R9773 VSS.n198 VSS.n185 0.001007
R9774 VSS.n4785 VSS.n4784 0.001007
R9775 VSS.n4453 VSS.n4359 0.001007
R9776 VSS.n4404 VSS.n4361 0.001007
R9777 VSS.n4408 VSS.n4369 0.001007
R9778 VSS.n4986 VSS.n4985 0.001007
R9779 VSS.n4578 VSS.n4577 0.001007
R9780 VSS.n4494 VSS.n4493 0.001007
R9781 VSS.n4498 VSS.n4497 0.001007
R9782 VSS.n4613 VSS.n4612 0.001007
R9783 VSS.n3880 VSS.n2863 0.001007
R9784 VSS.n5273 VSS.n3888 0.001007
R9785 VSS.n4299 VSS.n3893 0.001007
R9786 VSS.n5270 VSS.n5269 0.001007
R9787 VSS.n4348 VSS.n4282 0.001007
R9788 VSS.n4290 VSS.n4287 0.001007
R9789 VSS.n4345 VSS.n4344 0.001007
R9790 VSS.n4337 VSS.n4271 0.001007
R9791 VSS.n4270 VSS.n4262 0.001007
R9792 VSS.n4656 VSS.n4259 0.001007
R9793 VSS.n4624 VSS.n4623 0.001007
R9794 VSS.n4957 VSS.n4203 0.001007
R9795 VSS.n4372 VSS.n4200 0.001007
R9796 VSS.n4963 VSS.n4195 0.001007
R9797 VSS.n4480 VSS.n4479 0.001007
R9798 VSS.n4483 VSS.n4400 0.001007
R9799 VSS.n4864 VSS.n4863 0.001007
R9800 VSS.n4868 VSS.n4867 0.001007
R9801 VSS.n5096 VSS.n5095 0.001007
R9802 VSS.n4143 VSS.n4142 0.001007
R9803 VSS.n4147 VSS.n4146 0.001007
R9804 VSS.n5667 VSS.n5666 0.001007
R9805 VSS.n4886 VSS.n4885 0.001007
R9806 VSS.n4761 VSS.n4760 0.001007
R9807 VSS.n4765 VSS.n4764 0.001007
R9808 VSS.n4927 VSS.n4747 0.001007
R9809 VSS.n4841 VSS.n4749 0.001007
R9810 VSS.n4919 VSS.n4844 0.001007
R9811 VSS.n5159 VSS.n4118 0.001007
R9812 VSS.n4912 VSS.n4120 0.001007
R9813 VSS.n5146 VSS.n4127 0.001007
R9814 VSS.n5136 VSS.n5128 0.001007
R9815 VSS.n4834 VSS.n4806 0.001007
R9816 VSS.n4828 VSS.n4820 0.001007
R9817 VSS.n4817 VSS.n4814 0.001007
R9818 VSS.n4238 VSS.n4234 0.001007
R9819 VSS.n4237 VSS.n4235 0.001007
R9820 VSS.n4694 VSS.n4231 0.001007
R9821 VSS.n4229 VSS.n4228 0.001007
R9822 VSS.n4729 VSS.n4703 0.001007
R9823 VSS.n4713 VSS.n4705 0.001007
R9824 VSS.n5208 VSS.n4102 0.001007
R9825 VSS.n5198 VSS.n5190 0.001007
R9826 VSS.n4253 VSS.n4242 0.001007
R9827 VSS.n4661 VSS.n4256 0.001007
R9828 VSS.n4263 VSS.n4245 0.001007
R9829 VSS.n4037 VSS.n4030 0.001007
R9830 VSS.n4018 VSS.n4015 0.001007
R9831 VSS.n4027 VSS.n4012 0.001007
R9832 VSS.n4050 VSS.n4008 0.001007
R9833 VSS.n4020 VSS.n3997 0.001007
R9834 VSS.n4005 VSS.n3994 0.001007
R9835 VSS.n3990 VSS.n3986 0.001007
R9836 VSS.n3989 VSS.n3987 0.001007
R9837 VSS.n4089 VSS.n3983 0.001007
R9838 VSS.n4070 VSS.n3944 0.001007
R9839 VSS.n3972 VSS.n3946 0.001007
R9840 VSS.n3962 VSS.n3954 0.001007
R9841 VSS.n5258 VSS.n3906 0.001007
R9842 VSS.n3904 VSS.n3903 0.001007
R9843 VSS.n4295 VSS.n3901 0.001007
R9844 VSS.n3780 VSS.n3779 0.001007
R9845 VSS.n3784 VSS.n3783 0.001007
R9846 VSS.n3694 VSS.n3693 0.001007
R9847 VSS.n3682 VSS.n3681 0.001007
R9848 VSS.n3686 VSS.n3685 0.001007
R9849 VSS.n3596 VSS.n3595 0.001007
R9850 VSS.n3584 VSS.n3583 0.001007
R9851 VSS.n3588 VSS.n3587 0.001007
R9852 VSS.n3499 VSS.n3498 0.001007
R9853 VSS.n3487 VSS.n3486 0.001007
R9854 VSS.n3491 VSS.n3490 0.001007
R9855 VSS.n3402 VSS.n3401 0.001007
R9856 VSS.n3390 VSS.n3389 0.001007
R9857 VSS.n3394 VSS.n3393 0.001007
R9858 VSS.n5340 VSS.n5339 0.001007
R9859 VSS.n2828 VSS.n2827 0.001007
R9860 VSS.n5443 VSS.n5425 0.001007
R9861 VSS.n3792 VSS.n3773 0.001007
R9862 VSS.n3797 VSS.n3796 0.001007
R9863 VSS.n5433 VSS.n5432 0.001007
R9864 VSS.n5436 VSS.n5426 0.001007
R9865 VSS.n5772 VSS.n2385 0.001007
R9866 VSS.n3955 VSS.n2387 0.001007
R9867 VSS.n5740 VSS.n2404 0.001007
R9868 VSS.n5191 VSS.n2406 0.001007
R9869 VSS.n5708 VSS.n2423 0.001007
R9870 VSS.n5129 VSS.n2425 0.001007
R9871 VSS.n2460 VSS.n2459 0.001007
R9872 VSS.n2464 VSS.n2463 0.001007
R9873 VSS.n2578 VSS.n2563 0.001007
R9874 VSS.n2561 VSS.n2554 0.001007
R9875 VSS.n2532 VSS.n2531 0.001007
R9876 VSS.n2536 VSS.n2529 0.001007
R9877 VSS.n2612 VSS.n2511 0.001007
R9878 VSS.n5619 VSS.n5618 0.001007
R9879 VSS.n397 VSS.n396 0.001007
R9880 VSS.n2734 VSS.n2733 0.001007
R9881 VSS.n7459 VSS.n311 0.001007
R9882 VSS.n645 VSS.n316 0.001007
R9883 VSS.n601 VSS.n600 0.001007
R9884 VSS.n7499 VSS.n7498 0.001007
R9885 VSS.n7503 VSS.n7502 0.001007
R9886 VSS.n632 VSS.n532 0.001007
R9887 VSS.n675 VSS.n674 0.001007
R9888 VSS.n6665 VSS.n789 0.001007
R9889 VSS.n822 VSS.n791 0.001007
R9890 VSS.n781 VSS.n761 0.001007
R9891 VSS.n760 VSS.n759 0.001007
R9892 VSS.n7195 VSS.n753 0.001007
R9893 VSS.n7091 VSS.n7082 0.001007
R9894 VSS.n7192 VSS.n7191 0.001007
R9895 VSS.n641 VSS.n630 0.001007
R9896 VSS.n662 VSS.n628 0.001007
R9897 VSS.n7487 VSS.n7486 0.001007
R9898 VSS.n507 VSS.n506 0.001007
R9899 VSS.n502 VSS.n438 0.001007
R9900 VSS.n7327 VSS.n7326 0.001007
R9901 VSS.n373 VSS.n372 0.001007
R9902 VSS.n377 VSS.n376 0.001007
R9903 VSS.n7415 VSS.n341 0.001007
R9904 VSS.n695 VSS.n343 0.001007
R9905 VSS.n7259 VSS.n698 0.001007
R9906 VSS.n7357 VSS.n7256 0.001007
R9907 VSS.n7356 VSS.n7257 0.001007
R9908 VSS.n7376 VSS.n89 0.001007
R9909 VSS.n88 VSS.n87 0.001007
R9910 VSS.n688 VSS.n418 0.001007
R9911 VSS.n682 VSS.n429 0.001007
R9912 VSS.n433 VSS.n426 0.001007
R9913 VSS.n7120 VSS.n7113 0.001007
R9914 VSS.n7111 VSS.n7110 0.001007
R9915 VSS.n7160 VSS.n7133 0.001007
R9916 VSS.n7139 VSS.n7135 0.001007
R9917 VSS.n7243 VSS.n721 0.001007
R9918 VSS.n7143 VSS.n719 0.001007
R9919 VSS.n6923 VSS.n6897 0.001007
R9920 VSS.n6913 VSS.n6905 0.001007
R9921 VSS.n7180 VSS.n7104 0.001007
R9922 VSS.n7102 VSS.n7101 0.001007
R9923 VSS.n7099 VSS.n7090 0.001007
R9924 VSS.n7024 VSS.n808 0.001007
R9925 VSS.n846 VSS.n810 0.001007
R9926 VSS.n886 VSS.n849 0.001007
R9927 VSS.n898 VSS.n897 0.001007
R9928 VSS.n894 VSS.n885 0.001007
R9929 VSS.n904 VSS.n877 0.001007
R9930 VSS.n6998 VSS.n873 0.001007
R9931 VSS.n912 VSS.n875 0.001007
R9932 VSS.n6867 VSS.n915 0.001007
R9933 VSS.n6881 VSS.n6880 0.001007
R9934 VSS.n6874 VSS.n6866 0.001007
R9935 VSS.n6967 VSS.n6857 0.001007
R9936 VSS.n6957 VSS.n6949 0.001007
R9937 VSS.n839 VSS.n813 0.001007
R9938 VSS.n833 VSS.n832 0.001007
R9939 VSS.n829 VSS.n821 0.001007
R9940 VSS.n1084 VSS.n1083 0.001007
R9941 VSS.n1079 VSS.n1078 0.001007
R9942 VSS.n6559 VSS.n6558 0.001007
R9943 VSS.n1118 VSS.n1117 0.001007
R9944 VSS.n1113 VSS.n1112 0.001007
R9945 VSS.n6492 VSS.n6491 0.001007
R9946 VSS.n6480 VSS.n6479 0.001007
R9947 VSS.n6484 VSS.n6483 0.001007
R9948 VSS.n6406 VSS.n6405 0.001007
R9949 VSS.n1169 VSS.n1168 0.001007
R9950 VSS.n1164 VSS.n1163 0.001007
R9951 VSS.n1282 VSS.n1281 0.001007
R9952 VSS.n1270 VSS.n1269 0.001007
R9953 VSS.n1274 VSS.n1273 0.001007
R9954 VSS.n6850 VSS.n938 0.001007
R9955 VSS.n952 VSS.n951 0.001007
R9956 VSS.n6156 VSS.n6155 0.001007
R9957 VSS.n6153 VSS.n6152 0.001007
R9958 VSS.n1071 VSS.n1070 0.001007
R9959 VSS.n1068 VSS.n1067 0.001007
R9960 VSS.n6169 VSS.n6168 0.001007
R9961 VSS.n6164 VSS.n6163 0.001007
R9962 VSS.n7716 VSS.n28 0.001007
R9963 VSS.n6950 VSS.n30 0.001007
R9964 VSS.n7684 VSS.n47 0.001007
R9965 VSS.n6906 VSS.n49 0.001007
R9966 VSS.n7652 VSS.n66 0.001007
R9967 VSS.n80 VSS.n68 0.001007
R9968 VSS.n177 VSS.n176 0.001007
R9969 VSS.n181 VSS.n180 0.001007
R9970 VSS.n141 VSS.n140 0.001007
R9971 VSS.n7646 VSS.n7643 0.001007
R9972 VSS.n7678 VSS.n7675 0.001007
R9973 VSS.n7710 VSS.n7707 0.001007
R9974 VSS.n7587 VSS.n7586 0.001007
R9975 VSS.n192 VSS.n191 0.001007
R9976 VSS.n2481 VSS.n2480 0.001007
R9977 VSS.n5702 VSS.n5699 0.001007
R9978 VSS.n5734 VSS.n5731 0.001007
R9979 VSS.n5766 VSS.n5763 0.001007
R9980 VSS.n4994 VSS.n4993 0.001007
R9981 VSS.n4780 VSS.n4779 0.001007
R9982 VSS.n4996 VSS.n4995 0.001007
R9983 VSS.n4444 VSS.n4443 0.001007
R9984 VSS.n4535 VSS.n4534 0.001007
R9985 VSS.n4189 VSS.n4188 0.001007
R9986 VSS.n4537 VSS.n4536 0.001007
R9987 VSS.n4585 VSS.n4584 0.001007
R9988 VSS.n4607 VSS.n4371 0.001007
R9989 VSS.n4616 VSS.n4366 0.001007
R9990 VSS.n4310 VSS.n3890 0.001007
R9991 VSS.n4316 VSS.n4283 0.001007
R9992 VSS.n4649 VSS.n4272 0.001007
R9993 VSS.n4627 VSS.n4356 0.001007
R9994 VSS.n4822 VSS.n4196 0.001007
R9995 VSS.n4439 VSS.n4438 0.001007
R9996 VSS.n5103 VSS.n5102 0.001007
R9997 VSS.n5674 VSS.n5673 0.001007
R9998 VSS.n4893 VSS.n4892 0.001007
R9999 VSS.n4921 VSS.n4845 0.001007
R10000 VSS.n5153 VSS.n4125 0.001007
R10001 VSS.n4131 VSS.n4123 0.001007
R10002 VSS.n5140 VSS.n5139 0.001007
R10003 VSS.n5123 VSS.n4129 0.001007
R10004 VSS.n4809 VSS.n4807 0.001007
R10005 VSS.n4687 VSS.n4686 0.001007
R10006 VSS.n4681 VSS.n4679 0.001007
R10007 VSS.n4737 VSS.n4701 0.001007
R10008 VSS.n4707 VSS.n4699 0.001007
R10009 VSS.n4723 VSS.n4721 0.001007
R10010 VSS.n4717 VSS.n4716 0.001007
R10011 VSS.n5202 VSS.n5201 0.001007
R10012 VSS.n5185 VSS.n4104 0.001007
R10013 VSS.n4668 VSS.n4667 0.001007
R10014 VSS.n4044 VSS.n4043 0.001007
R10015 VSS.n4057 VSS.n4056 0.001007
R10016 VSS.n4082 VSS.n4081 0.001007
R10017 VSS.n4076 VSS.n4068 0.001007
R10018 VSS.n3980 VSS.n3941 0.001007
R10019 VSS.n4096 VSS.n4095 0.001007
R10020 VSS.n3966 VSS.n3965 0.001007
R10021 VSS.n3949 VSS.n3948 0.001007
R10022 VSS.n4031 VSS.n3907 0.001007
R10023 VSS.n3701 VSS.n3700 0.001007
R10024 VSS.n3603 VSS.n3602 0.001007
R10025 VSS.n3506 VSS.n3505 0.001007
R10026 VSS.n3409 VSS.n3408 0.001007
R10027 VSS.n5347 VSS.n5346 0.001007
R10028 VSS.n5446 VSS.n5445 0.001007
R10029 VSS.n2831 VSS.n2830 0.001007
R10030 VSS.n3874 VSS.n3873 0.001007
R10031 VSS.n5798 VSS.n5797 0.001007
R10032 VSS.n5793 VSS.n5792 0.001007
R10033 VSS.n5759 VSS.n2390 0.001007
R10034 VSS.n5727 VSS.n2409 0.001007
R10035 VSS.n5695 VSS.n2428 0.001007
R10036 VSS.n2488 VSS.n2487 0.001007
R10037 VSS.n2513 VSS.n2512 0.001007
R10038 VSS.n2600 VSS.n2526 0.001007
R10039 VSS.n2567 VSS.n2551 0.001007
R10040 VSS.n2585 VSS.n2584 0.001007
R10041 VSS.n2606 VSS.n2605 0.001007
R10042 VSS.n5612 VSS.n2630 0.001007
R10043 VSS.n457 VSS.n456 0.001007
R10044 VSS.n392 VSS.n391 0.001007
R10045 VSS.n459 VSS.n458 0.001007
R10046 VSS.n558 VSS.n557 0.001007
R10047 VSS.n608 VSS.n607 0.001007
R10048 VSS.n531 VSS.n530 0.001007
R10049 VSS.n668 VSS.n534 0.001007
R10050 VSS.n656 VSS.n654 0.001007
R10051 VSS.n6685 VSS.n6684 0.001007
R10052 VSS.n7042 VSS.n793 0.001007
R10053 VSS.n7049 VSS.n7048 0.001007
R10054 VSS.n7069 VSS.n7068 0.001007
R10055 VSS.n7065 VSS.n782 0.001007
R10056 VSS.n7077 VSS.n755 0.001007
R10057 VSS.n7453 VSS.n318 0.001007
R10058 VSS.n764 VSS.n312 0.001007
R10059 VSS.n650 VSS.n644 0.001007
R10060 VSS.n302 VSS.n301 0.001007
R10061 VSS.n2725 VSS.n2724 0.001007
R10062 VSS.n565 VSS.n564 0.001007
R10063 VSS.n7334 VSS.n7333 0.001007
R10064 VSS.n7409 VSS.n699 0.001007
R10065 VSS.n7371 VSS.n7370 0.001007
R10066 VSS.n7365 VSS.n7363 0.001007
R10067 VSS.n7615 VSS.n7614 0.001007
R10068 VSS.n7608 VSS.n90 0.001007
R10069 VSS.n421 VSS.n419 0.001007
R10070 VSS.n7168 VSS.n7131 0.001007
R10071 VSS.n7127 VSS.n7125 0.001007
R10072 VSS.n7154 VSS.n7152 0.001007
R10073 VSS.n7148 VSS.n7142 0.001007
R10074 VSS.n6892 VSS.n716 0.001007
R10075 VSS.n7250 VSS.n7249 0.001007
R10076 VSS.n6917 VSS.n6916 0.001007
R10077 VSS.n6900 VSS.n6899 0.001007
R10078 VSS.n7114 VSS.n7105 0.001007
R10079 VSS.n7018 VSS.n850 0.001007
R10080 VSS.n880 VSS.n878 0.001007
R10081 VSS.n6992 VSS.n916 0.001007
R10082 VSS.n6877 VSS.n6863 0.001007
R10083 VSS.n6888 VSS.n6887 0.001007
R10084 VSS.n6961 VSS.n6960 0.001007
R10085 VSS.n6944 VSS.n6859 0.001007
R10086 VSS.n816 VSS.n814 0.001007
R10087 VSS.n6566 VSS.n6565 0.001007
R10088 VSS.n6499 VSS.n6498 0.001007
R10089 VSS.n6413 VSS.n6412 0.001007
R10090 VSS.n1289 VSS.n1288 0.001007
R10091 VSS.n6844 VSS.n6843 0.001007
R10092 VSS.n945 VSS.n944 0.001007
R10093 VSS.n6687 VSS.n6686 0.001007
R10094 VSS.n7742 VSS.n7741 0.001007
R10095 VSS.n7737 VSS.n7736 0.001007
R10096 VSS.n7703 VSS.n33 0.001007
R10097 VSS.n7671 VSS.n52 0.001007
R10098 VSS.n7639 VSS.n71 0.001007
R10099 VSS.n148 VSS.n147 0.001007
R10100 VSS.n4309 VSS.n3891 0.00100685
R10101 VSS.n4652 VSS.n4651 0.00100685
R10102 VSS.n4442 VSS.n4440 0.00100685
R10103 VSS.n5126 VSS.n5125 0.00100685
R10104 VSS.n5188 VSS.n5187 0.00100685
R10105 VSS.n3952 VSS.n3951 0.00100685
R10106 VSS.n2823 VSS.n2821 0.00100685
R10107 VSS.n3878 VSS.n3876 0.00100685
R10108 VSS.n2525 VSS.n2524 0.00100685
R10109 VSS.n671 VSS.n670 0.00100685
R10110 VSS.n787 VSS.n786 0.00100685
R10111 VSS.n7080 VSS.n7079 0.00100685
R10112 VSS.n653 VSS.n652 0.00100685
R10113 VSS.n556 VSS.n554 0.00100685
R10114 VSS.n7611 VSS.n7610 0.00100685
R10115 VSS.n6903 VSS.n6902 0.00100685
R10116 VSS.n6947 VSS.n6946 0.00100685
R10117 VSS.n948 VSS.n946 0.00100685
R10118 VSS.n6848 VSS.n6847 0.00100685
R10119 VSS.n1286 VSS.n1285 0.00100685
R10120 VSS.n6410 VSS.n6409 0.00100685
R10121 VSS.n6496 VSS.n6495 0.00100685
R10122 VSS.n6995 VSS.n6994 0.00100685
R10123 VSS.n883 VSS.n882 0.00100685
R10124 VSS.n7584 VSS.n7583 0.00100685
R10125 VSS.n196 VSS.n195 0.00100685
R10126 VSS.n5344 VSS.n5343 0.00100685
R10127 VSS.n3406 VSS.n3405 0.00100685
R10128 VSS.n3503 VSS.n3502 0.00100685
R10129 VSS.n3600 VSS.n3599 0.00100685
R10130 VSS.n3995 VSS.n3992 0.00100685
R10131 VSS.n4821 VSS.n4198 0.00100685
R10132 VSS.n4582 VSS.n4580 0.00100685
R10133 VSS.n5100 VSS.n5099 0.00100685
R10134 VSS.n5671 VSS.n5670 0.00100685
R10135 VSS.n4890 VSS.n4888 0.00100685
R10136 VSS.n4924 VSS.n4923 0.00100685
R10137 VSS.n4130 VSS.n4124 0.00100685
R10138 VSS.n4812 VSS.n4811 0.00100685
R10139 VSS.n4684 VSS.n4683 0.00100685
R10140 VSS.n4706 VSS.n4700 0.00100685
R10141 VSS.n4720 VSS.n4719 0.00100685
R10142 VSS.n4243 VSS.n4240 0.00100685
R10143 VSS.n4013 VSS.n4010 0.00100685
R10144 VSS.n4079 VSS.n4078 0.00100685
R10145 VSS.n3940 VSS.n3939 0.00100685
R10146 VSS.n5260 VSS.n3909 0.00100685
R10147 VSS.n3698 VSS.n3697 0.00100685
R10148 VSS.n5796 VSS.n5794 0.00100685
R10149 VSS.n5762 VSS.n5761 0.00100685
R10150 VSS.n5730 VSS.n5729 0.00100685
R10151 VSS.n5698 VSS.n5697 0.00100685
R10152 VSS.n2479 VSS.n2477 0.00100685
R10153 VSS.n2550 VSS.n2549 0.00100685
R10154 VSS.n5615 VSS.n5614 0.00100685
R10155 VSS.n605 VSS.n603 0.00100685
R10156 VSS.n7331 VSS.n7329 0.00100685
R10157 VSS.n7412 VSS.n7411 0.00100685
R10158 VSS.n7368 VSS.n7367 0.00100685
R10159 VSS.n424 VSS.n423 0.00100685
R10160 VSS.n7130 VSS.n7129 0.00100685
R10161 VSS.n7151 VSS.n7150 0.00100685
R10162 VSS.n715 VSS.n714 0.00100685
R10163 VSS.n7182 VSS.n7107 0.00100685
R10164 VSS.n7021 VSS.n7020 0.00100685
R10165 VSS.n6862 VSS.n6861 0.00100685
R10166 VSS.n819 VSS.n818 0.00100685
R10167 VSS.n6563 VSS.n6562 0.00100685
R10168 VSS.n7740 VSS.n7738 0.00100685
R10169 VSS.n7706 VSS.n7705 0.00100685
R10170 VSS.n7674 VSS.n7673 0.00100685
R10171 VSS.n7642 VSS.n7641 0.00100685
R10172 VSS.n139 VSS.n137 0.00100685
R10173 VSS.n3811 VSS.n3810 0.00100593
R10174 VSS.n3714 VSS.n3713 0.00100593
R10175 VSS.n3616 VSS.n3615 0.00100593
R10176 VSS.n3519 VSS.n3518 0.00100593
R10177 VSS.n3422 VSS.n3421 0.00100593
R10178 VSS.n3325 VSS.n3324 0.00100593
R10179 VSS.n5462 VSS.n5461 0.00100593
R10180 VSS.n5811 VSS.n5810 0.00100593
R10181 VSS.n6650 VSS.n6649 0.00100593
R10182 VSS.n1101 VSS.n1100 0.00100593
R10183 VSS.n1128 VSS.n1127 0.00100593
R10184 VSS.n6427 VSS.n6426 0.00100593
R10185 VSS.n1223 VSS.n1222 0.00100593
R10186 VSS.n972 VSS.n971 0.00100593
R10187 VSS.n6137 VSS.n6136 0.00100593
R10188 VSS.n10 VSS.n9 0.00100593
R10189 VSS.n2498 VSS.n2497 0.00100588
R10190 VSS.n1100 VSS.n1099 0.00100584
R10191 VSS.n6426 VSS.n6425 0.00100584
R10192 VSS.n5591 VSS.n5589 0.00100509
R10193 VSS.n5591 VSS.n5590 0.00100509
R10194 VSS.n988 VSS.n963 0.00100509
R10195 VSS.n999 VSS.n988 0.00100509
R10196 VSS.n6582 VSS.n1092 0.00100509
R10197 VSS.n6593 VSS.n6582 0.00100509
R10198 VSS.n6611 VSS.n6606 0.00100509
R10199 VSS.n6612 VSS.n6611 0.00100509
R10200 VSS.n1052 VSS.n1039 0.00100509
R10201 VSS.n1052 VSS.n1051 0.00100509
R10202 VSS.n1036 VSS.n1030 0.00100509
R10203 VSS.n1036 VSS.n1035 0.00100509
R10204 VSS.n3843 VSS.n2867 0.00100509
R10205 VSS.n3849 VSS.n3843 0.00100509
R10206 VSS.n3827 VSS.n2869 0.00100509
R10207 VSS.n3833 VSS.n3827 0.00100509
R10208 VSS.n3438 VSS.n2910 0.00100509
R10209 VSS.n3444 VSS.n3438 0.00100509
R10210 VSS.n5829 VSS.n2105 0.00100509
R10211 VSS.n5835 VSS.n5829 0.00100509
R10212 VSS.n5400 VSS.n5392 0.00100509
R10213 VSS.n5406 VSS.n5400 0.00100509
R10214 VSS.n5478 VSS.n5383 0.00100509
R10215 VSS.n5484 VSS.n5478 0.00100509
R10216 VSS.n5372 VSS.n2808 0.00100509
R10217 VSS.n5372 VSS.n5371 0.00100509
R10218 VSS.n3341 VSS.n3315 0.00100509
R10219 VSS.n3347 VSS.n3341 0.00100509
R10220 VSS.n3357 VSS.n2919 0.00100509
R10221 VSS.n3363 VSS.n3357 0.00100509
R10222 VSS.n3454 VSS.n2907 0.00100509
R10223 VSS.n3460 VSS.n3454 0.00100509
R10224 VSS.n3535 VSS.n2898 0.00100509
R10225 VSS.n3541 VSS.n3535 0.00100509
R10226 VSS.n3551 VSS.n2896 0.00100509
R10227 VSS.n3557 VSS.n3551 0.00100509
R10228 VSS.n3632 VSS.n2887 0.00100509
R10229 VSS.n3638 VSS.n3632 0.00100509
R10230 VSS.n3648 VSS.n2885 0.00100509
R10231 VSS.n3654 VSS.n3648 0.00100509
R10232 VSS.n3730 VSS.n2878 0.00100509
R10233 VSS.n3736 VSS.n3730 0.00100509
R10234 VSS.n3746 VSS.n2876 0.00100509
R10235 VSS.n3752 VSS.n3746 0.00100509
R10236 VSS.n6516 VSS.n6515 0.00100509
R10237 VSS.n6534 VSS.n6533 0.00100509
R10238 VSS.n6064 VSS.n6058 0.00100509
R10239 VSS.n6075 VSS.n6064 0.00100509
R10240 VSS.n6194 VSS.n6081 0.00100509
R10241 VSS.n6117 VSS.n6104 0.00100509
R10242 VSS.n6117 VSS.n6116 0.00100509
R10243 VSS.n6815 VSS.n6809 0.00100509
R10244 VSS.n1311 VSS.n1305 0.00100509
R10245 VSS.n1247 VSS.n1235 0.00100509
R10246 VSS.n1247 VSS.n1246 0.00100509
R10247 VSS.n6379 VSS.n6374 0.00100509
R10248 VSS.n6385 VSS.n6379 0.00100509
R10249 VSS.n6439 VSS.n1155 0.00100509
R10250 VSS.n6440 VSS.n6439 0.00100509
R10251 VSS.n6450 VSS.n1148 0.00100509
R10252 VSS.n6456 VSS.n6450 0.00100509
R10253 VSS.n5584 VSS.n5578 0.00100509
R10254 VSS.n5584 VSS.n5583 0.00100509
R10255 VSS.n5592 VSS.n2772 0.00100509
R10256 VSS.n1154 VSS.n1153 0.00100509
R10257 VSS.n6541 VSS.n6540 0.00100509
R10258 VSS.n6523 VSS.n6522 0.00100509
R10259 VSS.n6618 VSS.n6617 0.00100509
R10260 VSS.n361 VSS.n345 0.00100462
R10261 VSS.n5821 VSS.n5815 0.00100462
R10262 VSS.n354 VSS.n353 0.00100462
R10263 VSS.n5574 VSS.n5573 0.00100381
R10264 VSS.n993 VSS.n989 0.00100381
R10265 VSS.n6587 VSS.n6583 0.00100381
R10266 VSS.n6617 VSS.n6613 0.00100381
R10267 VSS.n1044 VSS.n1040 0.00100381
R10268 VSS.n6712 VSS.n6711 0.00100381
R10269 VSS.n3848 VSS.n3844 0.00100381
R10270 VSS.n3832 VSS.n3828 0.00100381
R10271 VSS.n3443 VSS.n3439 0.00100381
R10272 VSS.n5834 VSS.n5830 0.00100381
R10273 VSS.n5405 VSS.n5401 0.00100381
R10274 VSS.n5483 VSS.n5479 0.00100381
R10275 VSS.n5370 VSS.n5366 0.00100381
R10276 VSS.n3346 VSS.n3342 0.00100381
R10277 VSS.n3362 VSS.n3358 0.00100381
R10278 VSS.n3459 VSS.n3455 0.00100381
R10279 VSS.n3540 VSS.n3536 0.00100381
R10280 VSS.n3556 VSS.n3552 0.00100381
R10281 VSS.n3637 VSS.n3633 0.00100381
R10282 VSS.n3653 VSS.n3649 0.00100381
R10283 VSS.n3735 VSS.n3731 0.00100381
R10284 VSS.n3751 VSS.n3747 0.00100381
R10285 VSS.n6522 VSS.n6518 0.00100381
R10286 VSS.n6540 VSS.n6536 0.00100381
R10287 VSS.n6069 VSS.n6065 0.00100381
R10288 VSS.n6086 VSS.n6082 0.00100381
R10289 VSS.n6109 VSS.n6105 0.00100381
R10290 VSS.n6814 VSS.n6810 0.00100381
R10291 VSS.n1310 VSS.n1306 0.00100381
R10292 VSS.n1240 VSS.n1236 0.00100381
R10293 VSS.n6384 VSS.n6380 0.00100381
R10294 VSS.n1153 VSS.n1149 0.00100381
R10295 VSS.n6455 VSS.n6451 0.00100381
R10296 VSS.n5572 VSS.n5563 0.00100381
R10297 VSS.n3818 VSS.n3817 0.0010038
R10298 VSS.n3721 VSS.n3720 0.0010038
R10299 VSS.n3623 VSS.n3622 0.0010038
R10300 VSS.n3526 VSS.n3525 0.0010038
R10301 VSS.n3429 VSS.n3428 0.0010038
R10302 VSS.n3332 VSS.n3331 0.0010038
R10303 VSS.n5469 VSS.n5468 0.0010038
R10304 VSS.n6657 VSS.n6656 0.0010038
R10305 VSS.n1134 VSS.n1133 0.0010038
R10306 VSS.n6425 VSS.n6424 0.0010038
R10307 VSS.n1219 VSS.n1218 0.0010038
R10308 VSS.n968 VSS.n967 0.0010038
R10309 VSS.n6131 VSS.n6130 0.0010038
R10310 VSS.n6 VSS.n5 0.0010038
R10311 VSS.n3819 VSS.n3818 0.00100371
R10312 VSS.n3722 VSS.n3721 0.00100371
R10313 VSS.n3624 VSS.n3623 0.00100371
R10314 VSS.n3527 VSS.n3526 0.00100371
R10315 VSS.n3430 VSS.n3429 0.00100371
R10316 VSS.n3333 VSS.n3332 0.00100371
R10317 VSS.n5470 VSS.n5469 0.00100371
R10318 VSS.n6656 VSS.n6655 0.00100371
R10319 VSS.n1095 VSS.n1094 0.00100371
R10320 VSS.n1135 VSS.n1134 0.00100371
R10321 VSS.n1220 VSS.n1219 0.00100371
R10322 VSS.n969 VSS.n968 0.00100371
R10323 VSS.n6132 VSS.n6131 0.00100371
R10324 VSS.n7 VSS.n6 0.00100371
R10325 VSS.n6713 VSS.n6712 0.00100369
R10326 VSS.n5573 VSS.n5572 0.00100369
R10327 VSS.n2238 VSS.n2237 0.00100208
R10328 VSS.n2109 VSS.n2108 0.00100208
R10329 VSS.n6328 VSS.n6327 0.00100208
R10330 VSS.n5597 VSS.n5596 0.00100206
R10331 VSS.n6345 VSS.n6344 0.00100116
R10332 VSS.n3860 VSS.n3859 0.00100116
R10333 VSS.n4424 VSS.n4423 0.00100116
R10334 VSS.n4524 VSS.n4523 0.00100116
R10335 VSS.n4557 VSS.n4556 0.00100116
R10336 VSS.n5029 VSS.n5028 0.00100116
R10337 VSS.n5051 VSS.n5050 0.00100116
R10338 VSS.n4160 VSS.n4159 0.00100116
R10339 VSS.n5646 VSS.n5645 0.00100116
R10340 VSS.n5079 VSS.n5078 0.00100116
R10341 VSS.n5067 VSS.n5066 0.00100116
R10342 VSS.n3762 VSS.n3761 0.00100116
R10343 VSS.n3664 VSS.n3663 0.00100116
R10344 VSS.n3566 VSS.n3565 0.00100116
R10345 VSS.n3469 VSS.n3468 0.00100116
R10346 VSS.n3372 VSS.n3371 0.00100116
R10347 VSS.n2811 VSS.n2810 0.00100116
R10348 VSS.n5415 VSS.n5414 0.00100116
R10349 VSS.n6336 VSS.n6335 0.00100116
R10350 VSS.n2759 VSS.n2758 0.00100116
R10351 VSS.n2749 VSS.n2748 0.00100116
R10352 VSS.n544 VSS.n543 0.00100116
R10353 VSS.n446 VSS.n445 0.00100116
R10354 VSS.n569 VSS.n568 0.00100116
R10355 VSS.n7520 VSS.n7519 0.00100116
R10356 VSS.n296 VSS.n295 0.00100116
R10357 VSS.n483 VSS.n482 0.00100116
R10358 VSS.n269 VSS.n268 0.00100116
R10359 VSS.n7266 VSS.n7265 0.00100116
R10360 VSS.n245 VSS.n244 0.00100116
R10361 VSS.n206 VSS.n205 0.00100116
R10362 VSS.n168 VSS.n167 0.00100116
R10363 VSS.n7560 VSS.n7559 0.00100116
R10364 VSS.n7308 VSS.n7307 0.00100116
R10365 VSS.n6626 VSS.n6625 0.00100116
R10366 VSS.n1345 VSS.n1344 0.00100116
R10367 VSS.n6463 VSS.n6462 0.00100116
R10368 VSS.n6369 VSS.n6368 0.00100116
R10369 VSS.n1229 VSS.n1228 0.00100116
R10370 VSS.n6824 VSS.n6823 0.00100116
R10371 VSS.n6184 VSS.n6183 0.00100116
R10372 VSS.n131 VSS.n130 0.00100116
R10373 VSS.n2652 VSS.n2651 0.00100062
R10374 VSS.n2674 VSS.n2673 0.00100062
R10375 VSS.n4625 VSS.n4360 0.00100058
R10376 VSS.n5271 VSS.n3892 0.00100058
R10377 VSS.n4346 VSS.n4286 0.00100058
R10378 VSS.n4655 VSS.n4260 0.00100058
R10379 VSS.n3795 VSS.n3772 0.00100058
R10380 VSS.n7193 VSS.n7081 0.00100058
R10381 VSS.n6154 VSS.n6146 0.00100058
R10382 VSS.n1069 VSS.n1062 0.00100058
R10383 VSS.n2107 VSS.n2106 0.0010004
R10384 VSS.n2236 VSS.n2235 0.0010004
R10385 VSS.n298 VSS.n297 0.00100034
R10386 VSS.n247 VSS.n246 0.00100034
R10387 VSS.n7268 VSS.n7267 0.00100034
R10388 VSS.n208 VSS.n207 0.00100034
R10389 VSS.n133 VSS.n132 0.00100034
R10390 VSS.n2700 VSS.n2699 0.00100033
R10391 VSS.n2641 VSS.n2640 0.00100031
R10392 VSS.n2688 VSS.n2687 0.00100031
R10393 VSS.n1659 VSS.n1658 0.00100031
R10394 VSS.n1542 VSS.n1541 0.00100031
R10395 VSS.n1407 VSS.n1406 0.00100031
R10396 VSS.n1504 VSS.n1503 0.00100031
R10397 VSS.n1621 VSS.n1620 0.00100031
R10398 VSS.n1556 VSS.n1555 0.00100031
R10399 VSS.n1487 VSS.n1486 0.00100031
R10400 VSS.n1380 VSS.n1379 0.00100031
R10401 VSS.n6343 VSS.n6341 0.00100024
R10402 VSS.n6689 VSS.n6683 0.00100023
R10403 VSS.n3568 VSS.n3564 0.00100022
R10404 VSS.n3471 VSS.n3467 0.00100022
R10405 VSS.n3374 VSS.n3370 0.00100022
R10406 VSS.n5360 VSS.n5358 0.00100022
R10407 VSS.n5417 VSS.n5413 0.00100022
R10408 VSS.n5073 VSS.n4162 0.00100021
R10409 VSS.n546 VSS.n542 0.00100021
R10410 VSS.n448 VSS.n444 0.00100021
R10411 VSS.n6182 VSS.n6101 0.00100021
R10412 VSS.n975 VSS.n974 0.00100021
R10413 VSS.n1226 VSS.n1225 0.00100021
R10414 VSS.n1104 VSS.n1103 0.00100021
R10415 VSS.n6652 VSS.n6648 0.00100021
R10416 VSS.n6466 VSS.n6465 0.00100021
R10417 VSS.n7756 VSS.n12 0.00100021
R10418 VSS.n5003 VSS.n5002 0.0010002
R10419 VSS.n4544 VSS.n4543 0.0010002
R10420 VSS.n466 VSS.n465 0.0010002
R10421 VSS.n4331 VSS.n4330 0.00100017
R10422 VSS.n4642 VSS.n4641 0.00100017
R10423 VSS.n4948 VSS.n4210 0.00100017
R10424 VSS.n5170 VSS.n5169 0.00100017
R10425 VSS.n5177 VSS.n5174 0.00100017
R10426 VSS.n5169 VSS.n5168 0.00100017
R10427 VSS.n4221 VSS.n4220 0.00100017
R10428 VSS.n4940 VSS.n4939 0.00100017
R10429 VSS.n5233 VSS.n5232 0.00100017
R10430 VSS.n5225 VSS.n5224 0.00100017
R10431 VSS.n5219 VSS.n3936 0.00100017
R10432 VSS.n5225 VSS.n3929 0.00100017
R10433 VSS.n5233 VSS.n3924 0.00100017
R10434 VSS.n5241 VSS.n5240 0.00100017
R10435 VSS.n5248 VSS.n3916 0.00100017
R10436 VSS.n5329 VSS.n5326 0.00100017
R10437 VSS.n2840 VSS.n2839 0.00100017
R10438 VSS.n5315 VSS.n5314 0.00100017
R10439 VSS.n5306 VSS.n5305 0.00100017
R10440 VSS.n5297 VSS.n5296 0.00100017
R10441 VSS.n5288 VSS.n5287 0.00100017
R10442 VSS.n5453 VSS.n5452 0.00100017
R10443 VSS.n5788 VSS.n2373 0.00100017
R10444 VSS.n5786 VSS.n2373 0.00100017
R10445 VSS.n5783 VSS.n5782 0.00100017
R10446 VSS.n5782 VSS.n5781 0.00100017
R10447 VSS.n5756 VSS.n2392 0.00100017
R10448 VSS.n5754 VSS.n2392 0.00100017
R10449 VSS.n5751 VSS.n5750 0.00100017
R10450 VSS.n5750 VSS.n5749 0.00100017
R10451 VSS.n5724 VSS.n2411 0.00100017
R10452 VSS.n5722 VSS.n2411 0.00100017
R10453 VSS.n5719 VSS.n5718 0.00100017
R10454 VSS.n5718 VSS.n5717 0.00100017
R10455 VSS.n2621 VSS.n2516 0.00100017
R10456 VSS.n2589 VSS.n2541 0.00100017
R10457 VSS.n7205 VSS.n7204 0.00100017
R10458 VSS.n7446 VSS.n7445 0.00100017
R10459 VSS.n7437 VSS.n7436 0.00100017
R10460 VSS.n7476 VSS.n7475 0.00100017
R10461 VSS.n7600 VSS.n7599 0.00100017
R10462 VSS.n7340 VSS.n7339 0.00100017
R10463 VSS.n7401 VSS.n7392 0.00100017
R10464 VSS.n7387 VSS.n711 0.00100017
R10465 VSS.n7401 VSS.n7400 0.00100017
R10466 VSS.n7395 VSS.n7394 0.00100017
R10467 VSS.n7428 VSS.n7427 0.00100017
R10468 VSS.n7235 VSS.n729 0.00100017
R10469 VSS.n6936 VSS.n6933 0.00100017
R10470 VSS.n7235 VSS.n7234 0.00100017
R10471 VSS.n732 VSS.n731 0.00100017
R10472 VSS.n7223 VSS.n7222 0.00100017
R10473 VSS.n7214 VSS.n7213 0.00100017
R10474 VSS.n6978 VSS.n936 0.00100017
R10475 VSS.n6983 VSS.n931 0.00100017
R10476 VSS.n927 VSS.n926 0.00100017
R10477 VSS.n7009 VSS.n865 0.00100017
R10478 VSS.n861 VSS.n860 0.00100017
R10479 VSS.n801 VSS.n800 0.00100017
R10480 VSS.n7732 VSS.n16 0.00100017
R10481 VSS.n7730 VSS.n16 0.00100017
R10482 VSS.n7727 VSS.n7726 0.00100017
R10483 VSS.n7726 VSS.n7725 0.00100017
R10484 VSS.n7700 VSS.n35 0.00100017
R10485 VSS.n7698 VSS.n35 0.00100017
R10486 VSS.n7695 VSS.n7694 0.00100017
R10487 VSS.n7694 VSS.n7693 0.00100017
R10488 VSS.n7668 VSS.n54 0.00100017
R10489 VSS.n7666 VSS.n54 0.00100017
R10490 VSS.n7663 VSS.n7662 0.00100017
R10491 VSS.n7662 VSS.n7661 0.00100017
R10492 VSS.n7627 VSS.n7626 0.00100017
R10493 VSS.n3802 VSS.n3801 0.00100017
R10494 VSS.n3705 VSS.n3704 0.00100017
R10495 VSS.n3607 VSS.n3606 0.00100017
R10496 VSS.n3510 VSS.n3509 0.00100017
R10497 VSS.n3413 VSS.n3412 0.00100017
R10498 VSS.n5351 VSS.n5350 0.00100017
R10499 VSS.n5606 VSS.n5605 0.00100017
R10500 VSS.n7539 VSS.n7538 0.00100017
R10501 VSS.n7278 VSS.n7277 0.00100017
R10502 VSS.n155 VSS.n154 0.00100017
R10503 VSS.n4330 VSS.n4329 0.00100017
R10504 VSS.n4641 VSS.n4640 0.00100017
R10505 VSS.n4211 VSS.n4210 0.00100017
R10506 VSS.n4970 VSS.n4969 0.00100017
R10507 VSS.n4599 VSS.n4598 0.00100017
R10508 VSS.n4470 VSS.n4469 0.00100017
R10509 VSS.n5110 VSS.n5109 0.00100017
R10510 VSS.n4907 VSS.n4906 0.00100017
R10511 VSS.n4800 VSS.n4799 0.00100017
R10512 VSS.n5175 VSS.n5174 0.00100017
R10513 VSS.n4220 VSS.n4218 0.00100017
R10514 VSS.n4941 VSS.n4940 0.00100017
R10515 VSS.n5217 VSS.n3936 0.00100017
R10516 VSS.n5240 VSS.n3922 0.00100017
R10517 VSS.n3917 VSS.n3916 0.00100017
R10518 VSS.n5327 VSS.n5326 0.00100017
R10519 VSS.n5323 VSS.n2840 0.00100017
R10520 VSS.n5314 VSS.n2844 0.00100017
R10521 VSS.n5305 VSS.n2848 0.00100017
R10522 VSS.n5296 VSS.n2852 0.00100017
R10523 VSS.n5287 VSS.n2856 0.00100017
R10524 VSS.n2517 VSS.n2516 0.00100017
R10525 VSS.n2545 VSS.n2541 0.00100017
R10526 VSS.n7204 VSS.n744 0.00100017
R10527 VSS.n7445 VSS.n7444 0.00100017
R10528 VSS.n7436 VSS.n331 0.00100017
R10529 VSS.n7475 VSS.n7474 0.00100017
R10530 VSS.n622 VSS.n621 0.00100017
R10531 VSS.n522 VSS.n521 0.00100017
R10532 VSS.n7601 VSS.n7600 0.00100017
R10533 VSS.n7341 VSS.n7340 0.00100017
R10534 VSS.n412 VSS.n411 0.00100017
R10535 VSS.n7385 VSS.n711 0.00100017
R10536 VSS.n7397 VSS.n7395 0.00100017
R10537 VSS.n7429 VSS.n7428 0.00100017
R10538 VSS.n6934 VSS.n6933 0.00100017
R10539 VSS.n7231 VSS.n732 0.00100017
R10540 VSS.n7222 VSS.n736 0.00100017
R10541 VSS.n7213 VSS.n740 0.00100017
R10542 VSS.n6976 VSS.n936 0.00100017
R10543 VSS.n932 VSS.n931 0.00100017
R10544 VSS.n926 VSS.n924 0.00100017
R10545 VSS.n866 VSS.n865 0.00100017
R10546 VSS.n860 VSS.n858 0.00100017
R10547 VSS.n7035 VSS.n801 0.00100017
R10548 VSS.n7585 VSS.n7584 0.00100016
R10549 VSS.n197 VSS.n196 0.00100016
R10550 VSS.n4583 VSS.n4582 0.00100016
R10551 VSS.n4962 VSS.n4198 0.00100016
R10552 VSS.n5101 VSS.n5100 0.00100016
R10553 VSS.n5672 VSS.n5671 0.00100016
R10554 VSS.n4891 VSS.n4890 0.00100016
R10555 VSS.n4925 VSS.n4924 0.00100016
R10556 VSS.n5157 VSS.n4124 0.00100016
R10557 VSS.n4833 VSS.n4812 0.00100016
R10558 VSS.n4684 VSS.n4233 0.00100016
R10559 VSS.n4741 VSS.n4700 0.00100016
R10560 VSS.n4727 VSS.n4720 0.00100016
R10561 VSS.n4666 VSS.n4243 0.00100016
R10562 VSS.n4042 VSS.n4013 0.00100016
R10563 VSS.n4055 VSS.n3995 0.00100016
R10564 VSS.n4079 VSS.n3985 0.00100016
R10565 VSS.n4094 VSS.n3940 0.00100016
R10566 VSS.n5261 VSS.n5260 0.00100016
R10567 VSS.n3699 VSS.n3698 0.00100016
R10568 VSS.n3601 VSS.n3600 0.00100016
R10569 VSS.n3504 VSS.n3503 0.00100016
R10570 VSS.n3407 VSS.n3406 0.00100016
R10571 VSS.n5345 VSS.n5344 0.00100016
R10572 VSS.n5799 VSS.n5796 0.00100016
R10573 VSS.n5770 VSS.n5762 0.00100016
R10574 VSS.n5738 VSS.n5730 0.00100016
R10575 VSS.n5706 VSS.n5698 0.00100016
R10576 VSS.n2486 VSS.n2479 0.00100016
R10577 VSS.n2583 VSS.n2550 0.00100016
R10578 VSS.n5615 VSS.n2629 0.00100016
R10579 VSS.n606 VSS.n605 0.00100016
R10580 VSS.n7332 VSS.n7331 0.00100016
R10581 VSS.n7413 VSS.n7412 0.00100016
R10582 VSS.n7368 VSS.n7255 0.00100016
R10583 VSS.n687 VSS.n424 0.00100016
R10584 VSS.n7172 VSS.n7130 0.00100016
R10585 VSS.n7158 VSS.n7151 0.00100016
R10586 VSS.n7248 VSS.n715 0.00100016
R10587 VSS.n7183 VSS.n7182 0.00100016
R10588 VSS.n7022 VSS.n7021 0.00100016
R10589 VSS.n903 VSS.n883 0.00100016
R10590 VSS.n6996 VSS.n6995 0.00100016
R10591 VSS.n6886 VSS.n6862 0.00100016
R10592 VSS.n838 VSS.n819 0.00100016
R10593 VSS.n6564 VSS.n6563 0.00100016
R10594 VSS.n6497 VSS.n6496 0.00100016
R10595 VSS.n6411 VSS.n6410 0.00100016
R10596 VSS.n1287 VSS.n1286 0.00100016
R10597 VSS.n6849 VSS.n6848 0.00100016
R10598 VSS.n7743 VSS.n7740 0.00100016
R10599 VSS.n7714 VSS.n7706 0.00100016
R10600 VSS.n7682 VSS.n7674 0.00100016
R10601 VSS.n7650 VSS.n7642 0.00100016
R10602 VSS.n146 VSS.n139 0.00100016
R10603 VSS.n5272 VSS.n3891 0.00100015
R10604 VSS.n4652 VSS.n4261 0.00100015
R10605 VSS.n4445 VSS.n4442 0.00100015
R10606 VSS.n5145 VSS.n5126 0.00100015
R10607 VSS.n5207 VSS.n5188 0.00100015
R10608 VSS.n3971 VSS.n3952 0.00100015
R10609 VSS.n2829 VSS.n2823 0.00100015
R10610 VSS.n3879 VSS.n3878 0.00100015
R10611 VSS.n2604 VSS.n2525 0.00100015
R10612 VSS.n671 VSS.n533 0.00100015
R10613 VSS.n7047 VSS.n787 0.00100015
R10614 VSS.n7194 VSS.n7080 0.00100015
R10615 VSS.n660 VSS.n653 0.00100015
R10616 VSS.n563 VSS.n556 0.00100015
R10617 VSS.n7611 VSS.n86 0.00100015
R10618 VSS.n6922 VSS.n6903 0.00100015
R10619 VSS.n6966 VSS.n6947 0.00100015
R10620 VSS.n950 VSS.n948 0.00100015
R10621 VSS.n146 VSS.n145 0.00100015
R10622 VSS.n7650 VSS.n7649 0.00100015
R10623 VSS.n7682 VSS.n7681 0.00100015
R10624 VSS.n7714 VSS.n7713 0.00100015
R10625 VSS.n2486 VSS.n2485 0.00100015
R10626 VSS.n5706 VSS.n5705 0.00100015
R10627 VSS.n5738 VSS.n5737 0.00100015
R10628 VSS.n5770 VSS.n5769 0.00100015
R10629 VSS.n4783 VSS.n4778 0.00100015
R10630 VSS.n5002 VSS.n5000 0.00100015
R10631 VSS.n4446 VSS.n4445 0.00100015
R10632 VSS.n4988 VSS.n4987 0.00100015
R10633 VSS.n4543 VSS.n4541 0.00100015
R10634 VSS.n4614 VSS.n4370 0.00100015
R10635 VSS.n4615 VSS.n4365 0.00100015
R10636 VSS.n4347 VSS.n4284 0.00100015
R10637 VSS.n4626 VSS.n4355 0.00100015
R10638 VSS.n5157 VSS.n5156 0.00100015
R10639 VSS.n5144 VSS.n5143 0.00100015
R10640 VSS.n4689 VSS.n4233 0.00100015
R10641 VSS.n4741 VSS.n4740 0.00100015
R10642 VSS.n4727 VSS.n4726 0.00100015
R10643 VSS.n5206 VSS.n5205 0.00100015
R10644 VSS.n4084 VSS.n3985 0.00100015
R10645 VSS.n4094 VSS.n3942 0.00100015
R10646 VSS.n3970 VSS.n3969 0.00100015
R10647 VSS.n5448 VSS.n5447 0.00100015
R10648 VSS.n5800 VSS.n5799 0.00100015
R10649 VSS.n2629 VSS.n2628 0.00100015
R10650 VSS.n2604 VSS.n2527 0.00100015
R10651 VSS.n2583 VSS.n2552 0.00100015
R10652 VSS.n395 VSS.n390 0.00100015
R10653 VSS.n465 VSS.n463 0.00100015
R10654 VSS.n7489 VSS.n7488 0.00100015
R10655 VSS.n563 VSS.n562 0.00100015
R10656 VSS.n528 VSS.n431 0.00100015
R10657 VSS.n660 VSS.n659 0.00100015
R10658 VSS.n7046 VSS.n7045 0.00100015
R10659 VSS.n7073 VSS.n7072 0.00100015
R10660 VSS.n7062 VSS.n758 0.00100015
R10661 VSS.n7457 VSS.n7456 0.00100015
R10662 VSS.n7458 VSS.n313 0.00100015
R10663 VSS.n2732 VSS.n2730 0.00100015
R10664 VSS.n7373 VSS.n7255 0.00100015
R10665 VSS.n7619 VSS.n7618 0.00100015
R10666 VSS.n7172 VSS.n7171 0.00100015
R10667 VSS.n7158 VSS.n7157 0.00100015
R10668 VSS.n7248 VSS.n717 0.00100015
R10669 VSS.n6921 VSS.n6920 0.00100015
R10670 VSS.n6886 VSS.n6864 0.00100015
R10671 VSS.n6965 VSS.n6964 0.00100015
R10672 VSS.n6690 VSS.n6689 0.00100015
R10673 VSS.n7744 VSS.n7743 0.00100015
R10674 VSS.n3870 VSS.n3869 0.00100011
R10675 VSS.n2576 VSS.n2575 0.00100011
R10676 VSS.n6695 VSS.n6694 0.00100011
R10677 VSS.n4880 VSS.n4857 0.00100011
R10678 VSS.n7321 VSS.n7280 0.00100011
R10679 VSS.n7525 VSS.n7524 0.0010001
R10680 VSS.n6186 VSS.n6185 0.0010001
R10681 VSS.n1126 VSS.n1125 0.0010001
R10682 VSS.n1146 VSS.n1145 0.0010001
R10683 VSS.n6373 VSS.n1175 0.0010001
R10684 VSS.n1321 VSS.n1320 0.0010001
R10685 VSS.n4512 VSS.n4511 0.00100009
R10686 VSS.n4511 VSS.n4510 0.00100009
R10687 VSS.n4572 VSS.n4571 0.00100009
R10688 VSS.n4572 VSS.n4377 0.00100009
R10689 VSS.n5017 VSS.n5016 0.00100009
R10690 VSS.n5016 VSS.n5015 0.00100009
R10691 VSS.n4773 VSS.n4772 0.00100009
R10692 VSS.n4773 VSS.n4750 0.00100009
R10693 VSS.n5661 VSS.n5660 0.00100009
R10694 VSS.n5661 VSS.n2439 0.00100009
R10695 VSS.n5090 VSS.n5089 0.00100009
R10696 VSS.n5090 VSS.n4136 0.00100009
R10697 VSS.n5805 VSS.n5804 0.00100009
R10698 VSS.n595 VSS.n594 0.00100009
R10699 VSS.n595 VSS.n593 0.00100009
R10700 VSS.n7535 VSS.n7534 0.00100009
R10701 VSS.n7535 VSS.n7533 0.00100009
R10702 VSS.n497 VSS.n496 0.00100009
R10703 VSS.n497 VSS.n495 0.00100009
R10704 VSS.n385 VSS.n384 0.00100009
R10705 VSS.n385 VSS.n344 0.00100009
R10706 VSS.n220 VSS.n219 0.00100009
R10707 VSS.n221 VSS.n220 0.00100009
R10708 VSS.n7574 VSS.n7573 0.00100009
R10709 VSS.n7574 VSS.n7572 0.00100009
R10710 VSS.n6638 VSS.n6637 0.00100009
R10711 VSS.n6553 VSS.n6552 0.00100009
R10712 VSS.n6472 VSS.n6471 0.00100009
R10713 VSS.n6400 VSS.n6399 0.00100009
R10714 VSS.n1262 VSS.n1261 0.00100009
R10715 VSS.n6838 VSS.n6837 0.00100009
R10716 VSS.n7749 VSS.n7748 0.00100009
R10717 VSS.n6173 VSS.n6144 0.00100009
R10718 VSS.n5650 VSS.n5649 0.00100008
R10719 VSS.n2450 VSS.n2449 0.00100008
R10720 VSS.n5076 VSS.n5075 0.00100008
R10721 VSS.n5065 VSS.n5064 0.00100008
R10722 VSS.n5057 VSS.n5056 0.00100008
R10723 VSS.n5049 VSS.n5048 0.00100008
R10724 VSS.n5035 VSS.n5034 0.00100008
R10725 VSS.n5027 VSS.n5026 0.00100008
R10726 VSS.n4183 VSS.n4182 0.00100008
R10727 VSS.n4561 VSS.n4560 0.00100008
R10728 VSS.n4530 VSS.n4529 0.00100008
R10729 VSS.n4522 VSS.n4521 0.00100008
R10730 VSS.n4395 VSS.n4394 0.00100008
R10731 VSS.n582 VSS.n581 0.00100008
R10732 VSS.n267 VSS.n266 0.00100008
R10733 VSS.n166 VSS.n165 0.00100008
R10734 VSS.n6831 VSS.n6830 0.00100008
R10735 VSS.n4155 VSS.n4154 0.00100007
R10736 VSS.n4881 VSS.n4880 0.00100007
R10737 VSS.n7322 VSS.n7321 0.00100007
R10738 VSS.n454 VSS.n453 0.00100007
R10739 VSS.n204 VSS.n203 0.00100006
R10740 VSS.n3814 VSS.n3813 0.00100006
R10741 VSS.n3717 VSS.n3716 0.00100006
R10742 VSS.n3619 VSS.n3618 0.00100006
R10743 VSS.n3522 VSS.n3521 0.00100006
R10744 VSS.n3425 VSS.n3424 0.00100006
R10745 VSS.n3328 VSS.n3327 0.00100006
R10746 VSS.n5465 VSS.n5464 0.00100006
R10747 VSS.n5814 VSS.n5813 0.00100006
R10748 VSS.n3862 VSS.n3858 0.00100006
R10749 VSS.n3764 VSS.n3760 0.00100006
R10750 VSS.n3666 VSS.n3662 0.00100006
R10751 VSS.n216 VSS.n202 0.00100006
R10752 VSS.n251 VSS.n250 0.00100006
R10753 VSS.n551 VSS.n536 0.00100006
R10754 VSS.n2753 VSS.n2751 0.00100006
R10755 VSS.n4426 VSS.n4422 0.00100006
R10756 VSS.n5642 VSS.n2500 0.00100006
R10757 VSS.n2368 VSS.n2367 0.00100006
R10758 VSS.n2363 VSS.n2362 0.00100006
R10759 VSS.n584 VSS.n583 0.00100005
R10760 VSS.n272 VSS.n271 0.00100005
R10761 VSS.n230 VSS.n229 0.00100005
R10762 VSS.n6829 VSS.n6828 0.00100005
R10763 VSS.n6319 VSS.n6309 0.00100002
R10764 VSS.n2195 VSS.n2194 0.00100002
R10765 VSS.n6320 VSS.n1878 0.00100001
R10766 VSS.n4391 VSS.n4390 0.001
R10767 VSS.n4384 VSS.n4383 0.001
R10768 VSS.n4179 VSS.n4178 0.001
R10769 VSS.n4172 VSS.n4171 0.001
R10770 VSS.n2446 VSS.n2445 0.001
R10771 VSS.n963 VSS.n962 0.001
R10772 VSS.n1092 VSS.n1091 0.001
R10773 VSS.n2867 VSS.n2866 0.001
R10774 VSS.n6523 VSS.n6517 0.001
R10775 VSS.n6541 VSS.n6535 0.001
R10776 VSS.n6058 VSS.n6057 0.001
R10777 VSS.n6088 VSS.n6087 0.001
R10778 VSS.n6817 VSS.n6816 0.001
R10779 VSS.n1313 VSS.n1312 0.001
R10780 VSS.n1235 VSS.n1234 0.001
R10781 VSS.n1155 VSS.n1154 0.001
R10782 VSS.n1148 VSS.n1147 0.001
R10783 VSS.n5060 VSS.n5059 0.001
R10784 VSS.n146 VSS.n141 0.001
R10785 VSS.n7650 VSS.n7643 0.001
R10786 VSS.n7682 VSS.n7675 0.001
R10787 VSS.n7714 VSS.n7707 0.001
R10788 VSS.n7586 VSS.n7585 0.001
R10789 VSS.n197 VSS.n192 0.001
R10790 VSS.n2486 VSS.n2481 0.001
R10791 VSS.n5706 VSS.n5699 0.001
R10792 VSS.n5738 VSS.n5731 0.001
R10793 VSS.n5770 VSS.n5763 0.001
R10794 VSS.n5002 VSS.n4994 0.001
R10795 VSS.n4783 VSS.n4780 0.001
R10796 VSS.n5002 VSS.n4996 0.001
R10797 VSS.n4445 VSS.n4444 0.001
R10798 VSS.n4543 VSS.n4535 0.001
R10799 VSS.n4987 VSS.n4189 0.001
R10800 VSS.n4543 VSS.n4537 0.001
R10801 VSS.n4584 VSS.n4583 0.001
R10802 VSS.n4614 VSS.n4371 0.001
R10803 VSS.n4616 VSS.n4615 0.001
R10804 VSS.n5272 VSS.n3890 0.001
R10805 VSS.n4347 VSS.n4283 0.001
R10806 VSS.n4272 VSS.n4261 0.001
R10807 VSS.n4627 VSS.n4626 0.001
R10808 VSS.n4962 VSS.n4196 0.001
R10809 VSS.n4445 VSS.n4439 0.001
R10810 VSS.n5102 VSS.n5101 0.001
R10811 VSS.n5673 VSS.n5672 0.001
R10812 VSS.n4892 VSS.n4891 0.001
R10813 VSS.n4925 VSS.n4845 0.001
R10814 VSS.n5157 VSS.n4125 0.001
R10815 VSS.n5157 VSS.n4123 0.001
R10816 VSS.n5144 VSS.n5139 0.001
R10817 VSS.n5145 VSS.n4129 0.001
R10818 VSS.n4833 VSS.n4807 0.001
R10819 VSS.n4687 VSS.n4233 0.001
R10820 VSS.n4679 VSS.n4233 0.001
R10821 VSS.n4741 VSS.n4701 0.001
R10822 VSS.n4741 VSS.n4699 0.001
R10823 VSS.n4727 VSS.n4721 0.001
R10824 VSS.n4727 VSS.n4716 0.001
R10825 VSS.n5206 VSS.n5201 0.001
R10826 VSS.n5207 VSS.n4104 0.001
R10827 VSS.n4667 VSS.n4666 0.001
R10828 VSS.n4043 VSS.n4042 0.001
R10829 VSS.n4056 VSS.n4055 0.001
R10830 VSS.n4082 VSS.n3985 0.001
R10831 VSS.n4068 VSS.n3985 0.001
R10832 VSS.n4094 VSS.n3941 0.001
R10833 VSS.n4095 VSS.n4094 0.001
R10834 VSS.n3970 VSS.n3965 0.001
R10835 VSS.n3971 VSS.n3948 0.001
R10836 VSS.n5261 VSS.n3907 0.001
R10837 VSS.n3700 VSS.n3699 0.001
R10838 VSS.n3602 VSS.n3601 0.001
R10839 VSS.n3505 VSS.n3504 0.001
R10840 VSS.n3408 VSS.n3407 0.001
R10841 VSS.n5346 VSS.n5345 0.001
R10842 VSS.n5447 VSS.n5446 0.001
R10843 VSS.n2830 VSS.n2829 0.001
R10844 VSS.n3879 VSS.n3874 0.001
R10845 VSS.n5799 VSS.n5798 0.001
R10846 VSS.n5799 VSS.n5793 0.001
R10847 VSS.n5770 VSS.n2390 0.001
R10848 VSS.n5738 VSS.n2409 0.001
R10849 VSS.n5706 VSS.n2428 0.001
R10850 VSS.n2487 VSS.n2486 0.001
R10851 VSS.n2629 VSS.n2513 0.001
R10852 VSS.n2604 VSS.n2526 0.001
R10853 VSS.n2583 VSS.n2551 0.001
R10854 VSS.n2584 VSS.n2583 0.001
R10855 VSS.n2605 VSS.n2604 0.001
R10856 VSS.n2630 VSS.n2629 0.001
R10857 VSS.n465 VSS.n457 0.001
R10858 VSS.n395 VSS.n392 0.001
R10859 VSS.n465 VSS.n459 0.001
R10860 VSS.n7488 VSS.n302 0.001
R10861 VSS.n563 VSS.n558 0.001
R10862 VSS.n607 VSS.n606 0.001
R10863 VSS.n530 VSS.n431 0.001
R10864 VSS.n534 VSS.n533 0.001
R10865 VSS.n660 VSS.n654 0.001
R10866 VSS.n6689 VSS.n6685 0.001
R10867 VSS.n7046 VSS.n793 0.001
R10868 VSS.n7048 VSS.n7047 0.001
R10869 VSS.n7073 VSS.n7068 0.001
R10870 VSS.n782 VSS.n758 0.001
R10871 VSS.n7194 VSS.n755 0.001
R10872 VSS.n7457 VSS.n318 0.001
R10873 VSS.n7458 VSS.n312 0.001
R10874 VSS.n660 VSS.n644 0.001
R10875 VSS.n2732 VSS.n2725 0.001
R10876 VSS.n564 VSS.n563 0.001
R10877 VSS.n7333 VSS.n7332 0.001
R10878 VSS.n7413 VSS.n699 0.001
R10879 VSS.n7371 VSS.n7255 0.001
R10880 VSS.n7363 VSS.n7255 0.001
R10881 VSS.n7619 VSS.n7614 0.001
R10882 VSS.n90 VSS.n86 0.001
R10883 VSS.n687 VSS.n419 0.001
R10884 VSS.n7172 VSS.n7131 0.001
R10885 VSS.n7172 VSS.n7125 0.001
R10886 VSS.n7158 VSS.n7152 0.001
R10887 VSS.n7158 VSS.n7142 0.001
R10888 VSS.n7248 VSS.n716 0.001
R10889 VSS.n7249 VSS.n7248 0.001
R10890 VSS.n6921 VSS.n6916 0.001
R10891 VSS.n6922 VSS.n6899 0.001
R10892 VSS.n7183 VSS.n7105 0.001
R10893 VSS.n7022 VSS.n850 0.001
R10894 VSS.n903 VSS.n878 0.001
R10895 VSS.n6996 VSS.n916 0.001
R10896 VSS.n6886 VSS.n6863 0.001
R10897 VSS.n6887 VSS.n6886 0.001
R10898 VSS.n6965 VSS.n6960 0.001
R10899 VSS.n6966 VSS.n6859 0.001
R10900 VSS.n838 VSS.n814 0.001
R10901 VSS.n6565 VSS.n6564 0.001
R10902 VSS.n6498 VSS.n6497 0.001
R10903 VSS.n6412 VSS.n6411 0.001
R10904 VSS.n1288 VSS.n1287 0.001
R10905 VSS.n6849 VSS.n6844 0.001
R10906 VSS.n950 VSS.n945 0.001
R10907 VSS.n6689 VSS.n6687 0.001
R10908 VSS.n7743 VSS.n7742 0.001
R10909 VSS.n7743 VSS.n7737 0.001
R10910 VSS.n7714 VSS.n33 0.001
R10911 VSS.n7682 VSS.n52 0.001
R10912 VSS.n7650 VSS.n71 0.001
R10913 VSS.n147 VSS.n146 0.001
R10914 VSS.n355 VSS.n354 0.001
R10915 VSS.n5564 VSS.n2772 0.001
R10916 VSS.n2492 VSS.n2475 0.001
R10917 VSS.n5585 VSS.n5584 0.001
R10918 VSS.n7289 VSS.n7287 0.001
R10919 VSS.n7291 VSS.n7289 0.001
R10920 VSS.n7585 VSS.n7580 0.001
R10921 VSS.n102 VSS.n100 0.001
R10922 VSS.n104 VSS.n102 0.001
R10923 VSS.n198 VSS.n197 0.001
R10924 VSS.n4785 VSS.n4783 0.001
R10925 VSS.n4483 VSS.n4482 0.001
R10926 VSS.n4626 VSS.n4359 0.001
R10927 VSS.n4615 VSS.n4369 0.001
R10928 VSS.n4987 VSS.n4986 0.001
R10929 VSS.n4583 VSS.n4578 0.001
R10930 VSS.n4496 VSS.n4494 0.001
R10931 VSS.n4498 VSS.n4496 0.001
R10932 VSS.n4614 VSS.n4613 0.001
R10933 VSS.n3880 VSS.n3879 0.001
R10934 VSS.n5273 VSS.n5272 0.001
R10935 VSS.n5271 VSS.n5270 0.001
R10936 VSS.n5271 VSS.n3893 0.001
R10937 VSS.n4348 VSS.n4347 0.001
R10938 VSS.n4346 VSS.n4345 0.001
R10939 VSS.n4346 VSS.n4287 0.001
R10940 VSS.n4337 VSS.n4261 0.001
R10941 VSS.n4656 VSS.n4655 0.001
R10942 VSS.n4655 VSS.n4262 0.001
R10943 VSS.n4625 VSS.n4624 0.001
R10944 VSS.n4625 VSS.n4361 0.001
R10945 VSS.n4961 VSS.n4203 0.001
R10946 VSS.n4961 VSS.n4200 0.001
R10947 VSS.n4963 VSS.n4962 0.001
R10948 VSS.n4482 VSS.n4480 0.001
R10949 VSS.n4866 VSS.n4864 0.001
R10950 VSS.n4868 VSS.n4866 0.001
R10951 VSS.n5101 VSS.n5096 0.001
R10952 VSS.n4145 VSS.n4143 0.001
R10953 VSS.n4147 VSS.n4145 0.001
R10954 VSS.n5672 VSS.n5667 0.001
R10955 VSS.n4891 VSS.n4886 0.001
R10956 VSS.n4763 VSS.n4761 0.001
R10957 VSS.n4765 VSS.n4763 0.001
R10958 VSS.n4927 VSS.n4926 0.001
R10959 VSS.n4926 VSS.n4749 0.001
R10960 VSS.n4925 VSS.n4844 0.001
R10961 VSS.n5159 VSS.n5158 0.001
R10962 VSS.n5158 VSS.n4120 0.001
R10963 VSS.n5146 VSS.n5145 0.001
R10964 VSS.n5144 VSS.n5128 0.001
R10965 VSS.n4834 VSS.n4833 0.001
R10966 VSS.n4832 VSS.n4820 0.001
R10967 VSS.n4832 VSS.n4814 0.001
R10968 VSS.n4677 VSS.n4238 0.001
R10969 VSS.n4677 VSS.n4237 0.001
R10970 VSS.n4742 VSS.n4231 0.001
R10971 VSS.n4742 VSS.n4228 0.001
R10972 VSS.n4729 VSS.n4728 0.001
R10973 VSS.n4728 VSS.n4705 0.001
R10974 VSS.n5208 VSS.n5207 0.001
R10975 VSS.n5206 VSS.n5190 0.001
R10976 VSS.n4666 VSS.n4242 0.001
R10977 VSS.n4665 VSS.n4256 0.001
R10978 VSS.n4665 VSS.n4245 0.001
R10979 VSS.n4041 VSS.n4030 0.001
R10980 VSS.n4041 VSS.n4015 0.001
R10981 VSS.n4042 VSS.n4012 0.001
R10982 VSS.n4054 VSS.n4008 0.001
R10983 VSS.n4054 VSS.n3997 0.001
R10984 VSS.n4055 VSS.n3994 0.001
R10985 VSS.n4066 VSS.n3990 0.001
R10986 VSS.n4066 VSS.n3989 0.001
R10987 VSS.n4093 VSS.n3983 0.001
R10988 VSS.n4093 VSS.n3944 0.001
R10989 VSS.n3972 VSS.n3971 0.001
R10990 VSS.n3970 VSS.n3954 0.001
R10991 VSS.n5261 VSS.n3906 0.001
R10992 VSS.n5262 VSS.n3904 0.001
R10993 VSS.n5262 VSS.n3901 0.001
R10994 VSS.n3782 VSS.n3780 0.001
R10995 VSS.n3784 VSS.n3782 0.001
R10996 VSS.n3699 VSS.n3694 0.001
R10997 VSS.n3684 VSS.n3682 0.001
R10998 VSS.n3686 VSS.n3684 0.001
R10999 VSS.n3601 VSS.n3596 0.001
R11000 VSS.n3586 VSS.n3584 0.001
R11001 VSS.n3588 VSS.n3586 0.001
R11002 VSS.n3504 VSS.n3499 0.001
R11003 VSS.n3489 VSS.n3487 0.001
R11004 VSS.n3491 VSS.n3489 0.001
R11005 VSS.n3407 VSS.n3402 0.001
R11006 VSS.n3392 VSS.n3390 0.001
R11007 VSS.n3394 VSS.n3392 0.001
R11008 VSS.n5345 VSS.n5340 0.001
R11009 VSS.n2829 VSS.n2828 0.001
R11010 VSS.n5447 VSS.n5443 0.001
R11011 VSS.n3797 VSS.n3795 0.001
R11012 VSS.n3795 VSS.n3792 0.001
R11013 VSS.n5435 VSS.n5433 0.001
R11014 VSS.n5436 VSS.n5435 0.001
R11015 VSS.n5772 VSS.n5771 0.001
R11016 VSS.n5771 VSS.n2387 0.001
R11017 VSS.n5740 VSS.n5739 0.001
R11018 VSS.n5739 VSS.n2406 0.001
R11019 VSS.n5708 VSS.n5707 0.001
R11020 VSS.n5707 VSS.n2425 0.001
R11021 VSS.n2462 VSS.n2460 0.001
R11022 VSS.n2464 VSS.n2462 0.001
R11023 VSS.n2603 VSS.n2529 0.001
R11024 VSS.n2582 VSS.n2563 0.001
R11025 VSS.n2582 VSS.n2554 0.001
R11026 VSS.n2603 VSS.n2531 0.001
R11027 VSS.n2612 VSS.n2510 0.001
R11028 VSS.n5619 VSS.n2510 0.001
R11029 VSS.n397 VSS.n395 0.001
R11030 VSS.n2734 VSS.n2732 0.001
R11031 VSS.n7459 VSS.n7458 0.001
R11032 VSS.n505 VSS.n502 0.001
R11033 VSS.n606 VSS.n601 0.001
R11034 VSS.n7501 VSS.n7499 0.001
R11035 VSS.n7503 VSS.n7501 0.001
R11036 VSS.n632 VSS.n533 0.001
R11037 VSS.n675 VSS.n431 0.001
R11038 VSS.n662 VSS.n661 0.001
R11039 VSS.n7047 VSS.n789 0.001
R11040 VSS.n7046 VSS.n791 0.001
R11041 VSS.n761 VSS.n758 0.001
R11042 VSS.n7073 VSS.n759 0.001
R11043 VSS.n7195 VSS.n7194 0.001
R11044 VSS.n7193 VSS.n7192 0.001
R11045 VSS.n7193 VSS.n7082 0.001
R11046 VSS.n7457 VSS.n316 0.001
R11047 VSS.n661 VSS.n630 0.001
R11048 VSS.n7488 VSS.n7487 0.001
R11049 VSS.n507 VSS.n505 0.001
R11050 VSS.n7332 VSS.n7327 0.001
R11051 VSS.n375 VSS.n373 0.001
R11052 VSS.n377 VSS.n375 0.001
R11053 VSS.n7415 VSS.n7414 0.001
R11054 VSS.n7414 VSS.n343 0.001
R11055 VSS.n7413 VSS.n698 0.001
R11056 VSS.n7361 VSS.n7357 0.001
R11057 VSS.n7361 VSS.n7356 0.001
R11058 VSS.n7376 VSS.n86 0.001
R11059 VSS.n7619 VSS.n87 0.001
R11060 VSS.n688 VSS.n687 0.001
R11061 VSS.n686 VSS.n429 0.001
R11062 VSS.n686 VSS.n426 0.001
R11063 VSS.n7173 VSS.n7113 0.001
R11064 VSS.n7173 VSS.n7110 0.001
R11065 VSS.n7160 VSS.n7159 0.001
R11066 VSS.n7159 VSS.n7135 0.001
R11067 VSS.n7247 VSS.n721 0.001
R11068 VSS.n7247 VSS.n719 0.001
R11069 VSS.n6923 VSS.n6922 0.001
R11070 VSS.n6921 VSS.n6905 0.001
R11071 VSS.n7183 VSS.n7104 0.001
R11072 VSS.n7184 VSS.n7102 0.001
R11073 VSS.n7184 VSS.n7090 0.001
R11074 VSS.n7024 VSS.n7023 0.001
R11075 VSS.n7023 VSS.n810 0.001
R11076 VSS.n7022 VSS.n849 0.001
R11077 VSS.n902 VSS.n897 0.001
R11078 VSS.n902 VSS.n885 0.001
R11079 VSS.n904 VSS.n903 0.001
R11080 VSS.n6998 VSS.n6997 0.001
R11081 VSS.n6997 VSS.n875 0.001
R11082 VSS.n6996 VSS.n915 0.001
R11083 VSS.n6885 VSS.n6880 0.001
R11084 VSS.n6885 VSS.n6866 0.001
R11085 VSS.n6967 VSS.n6966 0.001
R11086 VSS.n6965 VSS.n6949 0.001
R11087 VSS.n839 VSS.n838 0.001
R11088 VSS.n837 VSS.n832 0.001
R11089 VSS.n837 VSS.n821 0.001
R11090 VSS.n1084 VSS.n1082 0.001
R11091 VSS.n1082 VSS.n1079 0.001
R11092 VSS.n6564 VSS.n6559 0.001
R11093 VSS.n1118 VSS.n1116 0.001
R11094 VSS.n1116 VSS.n1113 0.001
R11095 VSS.n6497 VSS.n6492 0.001
R11096 VSS.n6482 VSS.n6480 0.001
R11097 VSS.n6484 VSS.n6482 0.001
R11098 VSS.n6411 VSS.n6406 0.001
R11099 VSS.n1169 VSS.n1167 0.001
R11100 VSS.n1167 VSS.n1164 0.001
R11101 VSS.n1287 VSS.n1282 0.001
R11102 VSS.n1272 VSS.n1270 0.001
R11103 VSS.n1274 VSS.n1272 0.001
R11104 VSS.n6850 VSS.n6849 0.001
R11105 VSS.n952 VSS.n950 0.001
R11106 VSS.n6154 VSS.n6153 0.001
R11107 VSS.n6156 VSS.n6154 0.001
R11108 VSS.n1069 VSS.n1068 0.001
R11109 VSS.n1071 VSS.n1069 0.001
R11110 VSS.n6169 VSS.n6167 0.001
R11111 VSS.n6167 VSS.n6164 0.001
R11112 VSS.n7716 VSS.n7715 0.001
R11113 VSS.n7715 VSS.n30 0.001
R11114 VSS.n7684 VSS.n7683 0.001
R11115 VSS.n7683 VSS.n49 0.001
R11116 VSS.n7652 VSS.n7651 0.001
R11117 VSS.n7651 VSS.n68 0.001
R11118 VSS.n179 VSS.n177 0.001
R11119 VSS.n181 VSS.n179 0.001
R11120 VSS.n2771 VSS.n2770 0.001
R11121 VSS.n5592 VSS.n5591 0.001
R11122 VSS.n988 VSS.n987 0.001
R11123 VSS.n6582 VSS.n6581 0.001
R11124 VSS.n6611 VSS.n6610 0.001
R11125 VSS.n1053 VSS.n1052 0.001
R11126 VSS.n1035 VSS.n1034 0.001
R11127 VSS.n3843 VSS.n3842 0.001
R11128 VSS.n3827 VSS.n3826 0.001
R11129 VSS.n3438 VSS.n3437 0.001
R11130 VSS.n5829 VSS.n5828 0.001
R11131 VSS.n5400 VSS.n5399 0.001
R11132 VSS.n5478 VSS.n5477 0.001
R11133 VSS.n5373 VSS.n5372 0.001
R11134 VSS.n3341 VSS.n3340 0.001
R11135 VSS.n3357 VSS.n3356 0.001
R11136 VSS.n3454 VSS.n3453 0.001
R11137 VSS.n3535 VSS.n3534 0.001
R11138 VSS.n3551 VSS.n3550 0.001
R11139 VSS.n3632 VSS.n3631 0.001
R11140 VSS.n3648 VSS.n3647 0.001
R11141 VSS.n3730 VSS.n3729 0.001
R11142 VSS.n3746 VSS.n3745 0.001
R11143 VSS.n6515 VSS.n6514 0.001
R11144 VSS.n6533 VSS.n6532 0.001
R11145 VSS.n6064 VSS.n6063 0.001
R11146 VSS.n6081 VSS.n6080 0.001
R11147 VSS.n6118 VSS.n6117 0.001
R11148 VSS.n6809 VSS.n6808 0.001
R11149 VSS.n1305 VSS.n1304 0.001
R11150 VSS.n1248 VSS.n1247 0.001
R11151 VSS.n6379 VSS.n6378 0.001
R11152 VSS.n6439 VSS.n6438 0.001
R11153 VSS.n6450 VSS.n6449 0.001
R11154 VSS.n5169 VSS.n4110 0.001
R11155 VSS.n5226 VSS.n5225 0.001
R11156 VSS.n5234 VSS.n5233 0.001
R11157 VSS.n2376 VSS.n2373 0.001
R11158 VSS.n5782 VSS.n2377 0.001
R11159 VSS.n2395 VSS.n2392 0.001
R11160 VSS.n5750 VSS.n2396 0.001
R11161 VSS.n2414 VSS.n2411 0.001
R11162 VSS.n5718 VSS.n2415 0.001
R11163 VSS.n5689 VSS.n5688 0.001
R11164 VSS.n2432 VSS.n2431 0.001
R11165 VSS.n7402 VSS.n7401 0.001
R11166 VSS.n7236 VSS.n7235 0.001
R11167 VSS.n19 VSS.n16 0.001
R11168 VSS.n7726 VSS.n20 0.001
R11169 VSS.n38 VSS.n35 0.001
R11170 VSS.n7694 VSS.n39 0.001
R11171 VSS.n57 VSS.n54 0.001
R11172 VSS.n7662 VSS.n58 0.001
R11173 VSS.n7633 VSS.n7632 0.001
R11174 VSS.n7626 VSS.n7625 0.001
R11175 VSS.n5636 VSS.n5635 0.000990196
R11176 VSS.n2713 VSS.n2712 0.000990196
R11177 VSS.n5604 VSS.n5603 0.000990196
R11178 VSS.n5602 VSS.n5601 0.000990196
R11179 VSS VSS.n1323 0.000820819
R11180 VSS.n2220 VSS.n2219 0.000801468
R11181 VSS.n3803 VSS.n2873 0.000760417
R11182 VSS.n3706 VSS.n2882 0.000760417
R11183 VSS.n3608 VSS.n2891 0.000760417
R11184 VSS.n3511 VSS.n2902 0.000760417
R11185 VSS.n3414 VSS.n2914 0.000760417
R11186 VSS.n5352 VSS.n2818 0.000760417
R11187 VSS.n5454 VSS.n5387 0.000760417
R11188 VSS.n6639 VSS.n1060 0.000760417
R11189 VSS.n6570 VSS.n1107 0.000760417
R11190 VSS.n6503 VSS.n1141 0.000760417
R11191 VSS.n6417 VSS.n1158 0.000760417
R11192 VSS.n1294 VSS.n1293 0.000760417
R11193 VSS.n6839 VSS.n941 0.000760417
R11194 VSS.n6175 VSS.n6174 0.000760417
R11195 VSS.n2219 VSS.n2211 0.00073829
R11196 VSS.n2219 VSS.n2218 0.00073829
R11197 VSS.n2218 VSS.n2217 0.00073829
R11198 VSS.n6735 VSS.n6734 0.000712971
R11199 VSS.n6717 VSS.n6716 0.000712971
R11200 VSS.n2952 VSS.n2945 0.000712971
R11201 VSS.n2951 VSS.n2946 0.000712971
R11202 VSS.n3047 VSS.n3046 0.000712971
R11203 VSS.n3045 VSS.n3012 0.000712971
R11204 VSS.n3040 VSS.n3030 0.000712971
R11205 VSS.n3039 VSS.n3031 0.000712971
R11206 VSS.n3068 VSS.n3067 0.000712971
R11207 VSS.n3065 VSS.n3064 0.000712971
R11208 VSS.n3063 VSS.n2991 0.000712971
R11209 VSS.n3062 VSS.n2992 0.000712971
R11210 VSS.n3060 VSS.n2997 0.000712971
R11211 VSS.n3059 VSS.n2998 0.000712971
R11212 VSS.n3057 VSS.n3003 0.000712971
R11213 VSS.n3056 VSS.n3004 0.000712971
R11214 VSS.n3054 VSS.n3009 0.000712971
R11215 VSS.n3053 VSS.n3010 0.000712971
R11216 VSS.n3076 VSS.n3069 0.000712971
R11217 VSS.n3075 VSS.n3070 0.000712971
R11218 VSS.n3043 VSS.n3018 0.000712971
R11219 VSS.n3042 VSS.n3019 0.000712971
R11220 VSS.n3037 VSS.n3034 0.000712971
R11221 VSS.n3036 VSS.n3035 0.000712971
R11222 VSS.n3276 VSS.n3275 0.000712971
R11223 VSS.n3278 VSS.n3277 0.000712971
R11224 VSS.n3072 VSS.n3071 0.000712971
R11225 VSS.n3273 VSS.n3272 0.000712971
R11226 VSS.n5526 VSS.n2092 0.000712971
R11227 VSS.n5525 VSS.n2092 0.000712971
R11228 VSS.n5854 VSS.n2097 0.000712971
R11229 VSS.n5838 VSS.n5837 0.000712971
R11230 VSS.n3306 VSS.n3305 0.000712971
R11231 VSS.n5937 VSS.n5934 0.000712971
R11232 VSS.n5936 VSS.n5935 0.000712971
R11233 VSS.n6034 VSS.n6033 0.000712971
R11234 VSS.n6036 VSS.n6035 0.000712971
R11235 VSS.n6040 VSS.n1948 0.000712971
R11236 VSS.n6042 VSS.n6041 0.000712971
R11237 VSS.n6046 VSS.n1945 0.000712971
R11238 VSS.n6048 VSS.n6047 0.000712971
R11239 VSS.n6052 VSS.n1943 0.000712971
R11240 VSS.n6054 VSS.n6053 0.000712971
R11241 VSS.n6801 VSS.n6800 0.000712971
R11242 VSS.n5948 VSS.n5916 0.000712971
R11243 VSS.n5949 VSS.n5915 0.000712971
R11244 VSS.n5909 VSS.n5908 0.000712971
R11245 VSS.n5906 VSS.n5905 0.000712971
R11246 VSS.n5898 VSS.n5897 0.000712971
R11247 VSS.n5896 VSS.n5895 0.000712971
R11248 VSS.n5901 VSS.n5900 0.000712971
R11249 VSS.n5903 VSS.n5902 0.000712971
R11250 VSS.n5911 VSS.n2008 0.000712971
R11251 VSS.n5913 VSS.n5912 0.000712971
R11252 VSS.n5946 VSS.n5925 0.000712971
R11253 VSS.n5945 VSS.n5926 0.000712971
R11254 VSS.n5942 VSS.n5928 0.000712971
R11255 VSS.n5941 VSS.n5929 0.000712971
R11256 VSS.n5939 VSS.n5932 0.000712971
R11257 VSS.n5938 VSS.n5933 0.000712971
R11258 VSS.n5873 VSS.n2074 0.000712971
R11259 VSS.n5871 VSS.n2079 0.000712971
R11260 VSS.n5866 VSS.n2088 0.000712971
R11261 VSS.n5868 VSS.n2081 0.000712971
R11262 VSS.n5872 VSS.n2078 0.000712971
R11263 VSS.n5874 VSS.n2077 0.000712971
R11264 VSS.n5558 VSS.n2075 0.000712971
R11265 VSS.n5560 VSS.n5559 0.000712971
R11266 VSS.n6743 VSS.n1023 0.000712971
R11267 VSS.n6742 VSS.n1023 0.000712971
R11268 VSS.n5891 VSS.n2073 0.000712971
R11269 VSS.n5890 VSS.n5889 0.000712971
R11270 VSS.n5894 VSS.n2014 0.000712971
R11271 VSS.n5893 VSS.n2015 0.000712971
R11272 VSS.n6246 VSS.n6245 0.000712971
R11273 VSS.n6244 VSS.n1897 0.000712971
R11274 VSS.n2777 VSS.n2776 0.000712971
R11275 VSS.n2778 VSS.n2773 0.000712971
R11276 VSS.n5867 VSS.n2087 0.000712971
R11277 VSS.n5865 VSS.n2090 0.000712971
R11278 VSS.n2089 VSS.n1895 0.000712971
R11279 VSS.n6253 VSS.n1896 0.000712971
R11280 VSS.n6250 VSS.n6249 0.000712971
R11281 VSS.n6248 VSS.n6247 0.000712971
R11282 VSS.n5888 VSS.n5886 0.000712971
R11283 VSS.n5885 VSS.n5884 0.000712971
R11284 VSS.n5878 VSS.n5877 0.000712971
R11285 VSS.n5562 VSS.n5561 0.000712971
R11286 VSS.n5633 VSS.n5631 0.000684314
R11287 VSS.n5640 VSS.n5638 0.000684314
R11288 VSS.n5629 VSS.n2505 0.000684314
R11289 VSS.n2715 VSS.n2710 0.000684314
R11290 VSS.n5600 VSS.n2765 0.000684314
R11291 VSS.n6505 VSS.n1140 0.000672891
R11292 VSS.n6100 VSS 0.00066041
R11293 VSS VSS.n958 0.00066041
R11294 VSS.n6366 VSS 0.00066041
R11295 VSS VSS.n1349 0.00066041
R11296 VSS VSS.n1038 0.00066041
R11297 VSS.n6241 VSS.n1900 0.000606486
R11298 VSS.n6242 VSS.n1899 0.000606486
R11299 VSS.n6747 VSS.n1020 0.000606486
R11300 VSS.n6746 VSS.n6745 0.000606486
R11301 VSS.n3116 VSS.n3115 0.000606486
R11302 VSS.n3114 VSS.n3113 0.000606486
R11303 VSS.n3106 VSS.n2980 0.000606486
R11304 VSS.n3105 VSS.n3104 0.000606486
R11305 VSS.n3097 VSS.n2983 0.000606486
R11306 VSS.n3096 VSS.n3095 0.000606486
R11307 VSS.n3088 VSS.n2986 0.000606486
R11308 VSS.n3087 VSS.n3086 0.000606486
R11309 VSS.n3080 VSS.n2989 0.000606486
R11310 VSS.n3079 VSS.n3078 0.000606486
R11311 VSS.n3073 VSS.n2961 0.000606486
R11312 VSS.n3256 VSS.n3255 0.000606486
R11313 VSS.n3253 VSS.n2964 0.000606486
R11314 VSS.n3251 VSS.n2965 0.000606486
R11315 VSS.n3249 VSS.n2968 0.000606486
R11316 VSS.n3247 VSS.n2969 0.000606486
R11317 VSS.n3245 VSS.n2972 0.000606486
R11318 VSS.n3243 VSS.n2973 0.000606486
R11319 VSS.n3241 VSS.n2976 0.000606486
R11320 VSS.n3239 VSS.n2977 0.000606486
R11321 VSS.n3236 VSS.n3235 0.000606486
R11322 VSS.n3023 VSS.n3022 0.000606486
R11323 VSS.n5550 VSS.n5549 0.000606486
R11324 VSS.n5548 VSS.n5547 0.000606486
R11325 VSS.n3024 VSS.n2785 0.000606486
R11326 VSS.n5504 VSS.n5503 0.000606486
R11327 VSS.n5502 VSS.n5501 0.000606486
R11328 VSS.n5499 VSS.n2790 0.000606486
R11329 VSS.n5508 VSS.n5506 0.000606486
R11330 VSS.n5556 VSS.n5555 0.000606486
R11331 VSS.n5557 VSS.n2076 0.000606486
R11332 VSS.n5507 VSS.n2080 0.000606486
R11333 VSS.n3283 VSS.n3282 0.000606486
R11334 VSS.n3269 VSS.n2955 0.000606486
R11335 VSS.n3270 VSS.n2954 0.000606486
R11336 VSS.n2958 VSS.n2957 0.000606486
R11337 VSS.n3163 VSS.n3162 0.000606486
R11338 VSS.n3266 VSS.n3265 0.000606486
R11339 VSS.n3267 VSS.n3263 0.000606486
R11340 VSS.n3259 VSS.n3258 0.000606486
R11341 VSS.n3260 VSS.n2956 0.000606486
R11342 VSS.n3083 VSS.n2963 0.000606486
R11343 VSS.n3084 VSS.n3082 0.000606486
R11344 VSS.n2995 VSS.n2993 0.000606486
R11345 VSS.n2994 VSS.n2990 0.000606486
R11346 VSS.n3286 VSS.n3285 0.000606486
R11347 VSS.n3290 VSS.n3289 0.000606486
R11348 VSS.n3173 VSS.n3172 0.000606486
R11349 VSS.n3151 VSS.n3150 0.000606486
R11350 VSS.n3179 VSS.n3145 0.000606486
R11351 VSS.n3177 VSS.n3176 0.000606486
R11352 VSS.n3160 VSS.n3159 0.000606486
R11353 VSS.n3158 VSS.n3157 0.000606486
R11354 VSS.n3093 VSS.n3090 0.000606486
R11355 VSS.n3092 VSS.n2967 0.000606486
R11356 VSS.n3000 VSS.n2987 0.000606486
R11357 VSS.n3001 VSS.n2999 0.000606486
R11358 VSS.n3170 VSS.n3149 0.000606486
R11359 VSS.n3169 VSS.n2939 0.000606486
R11360 VSS.n3165 VSS.n3153 0.000606486
R11361 VSS.n3167 VSS.n3166 0.000606486
R11362 VSS.n3190 VSS.n3189 0.000606486
R11363 VSS.n3155 VSS.n3154 0.000606486
R11364 VSS.n3201 VSS.n3200 0.000606486
R11365 VSS.n3194 VSS.n3193 0.000606486
R11366 VSS.n3101 VSS.n2971 0.000606486
R11367 VSS.n3102 VSS.n3099 0.000606486
R11368 VSS.n3007 VSS.n3005 0.000606486
R11369 VSS.n3006 VSS.n2984 0.000606486
R11370 VSS.n3184 VSS.n3181 0.000606486
R11371 VSS.n3183 VSS.n2936 0.000606486
R11372 VSS.n3187 VSS.n3139 0.000606486
R11373 VSS.n3186 VSS.n3144 0.000606486
R11374 VSS.n3141 VSS.n3140 0.000606486
R11375 VSS.n3143 VSS.n3142 0.000606486
R11376 VSS.n3211 VSS.n3210 0.000606486
R11377 VSS.n3147 VSS.n3146 0.000606486
R11378 VSS.n3226 VSS.n3225 0.000606486
R11379 VSS.n3215 VSS.n3214 0.000606486
R11380 VSS.n3049 VSS.n2981 0.000606486
R11381 VSS.n3051 VSS.n3048 0.000606486
R11382 VSS.n3208 VSS.n3133 0.000606486
R11383 VSS.n3207 VSS.n2933 0.000606486
R11384 VSS.n3203 VSS.n3135 0.000606486
R11385 VSS.n3205 VSS.n3204 0.000606486
R11386 VSS.n3196 VSS.n3195 0.000606486
R11387 VSS.n3198 VSS.n3197 0.000606486
R11388 VSS.n3111 VSS.n3108 0.000606486
R11389 VSS.n3110 VSS.n2975 0.000606486
R11390 VSS.n3232 VSS.n3231 0.000606486
R11391 VSS.n3137 VSS.n3136 0.000606486
R11392 VSS.n3127 VSS.n3126 0.000606486
R11393 VSS.n3128 VSS.n3125 0.000606486
R11394 VSS.n3015 VSS.n3014 0.000606486
R11395 VSS.n3016 VSS.n3013 0.000606486
R11396 VSS.n3217 VSS.n2931 0.000606486
R11397 VSS.n3309 VSS.n3308 0.000606486
R11398 VSS.n3229 VSS.n3131 0.000606486
R11399 VSS.n3228 VSS.n3132 0.000606486
R11400 VSS.n3234 VSS.n3123 0.000606486
R11401 VSS.n3233 VSS.n3124 0.000606486
R11402 VSS.n3119 VSS.n3118 0.000606486
R11403 VSS.n3122 VSS.n3121 0.000606486
R11404 VSS.n3221 VSS.n3220 0.000606486
R11405 VSS.n3223 VSS.n3219 0.000606486
R11406 VSS.n5531 VSS.n2798 0.000606486
R11407 VSS.n5533 VSS.n2797 0.000606486
R11408 VSS.n3026 VSS.n2786 0.000606486
R11409 VSS.n3028 VSS.n3020 0.000606486
R11410 VSS.n2922 VSS.n2921 0.000606486
R11411 VSS.n2924 VSS.n2923 0.000606486
R11412 VSS.n5536 VSS.n2794 0.000606486
R11413 VSS.n5535 VSS.n2795 0.000606486
R11414 VSS.n5541 VSS.n2791 0.000606486
R11415 VSS.n5539 VSS.n2792 0.000606486
R11416 VSS.n5545 VSS.n2787 0.000606486
R11417 VSS.n5544 VSS.n5543 0.000606486
R11418 VSS.n5520 VSS.n5519 0.000606486
R11419 VSS.n5493 VSS.n2793 0.000606486
R11420 VSS.n5524 VSS.n2091 0.000606486
R11421 VSS.n5523 VSS.n5522 0.000606486
R11422 VSS.n5553 VSS.n5552 0.000606486
R11423 VSS.n3032 VSS.n2783 0.000606486
R11424 VSS.n5487 VSS.n2799 0.000606486
R11425 VSS.n5486 VSS.n2800 0.000606486
R11426 VSS.n5497 VSS.n5494 0.000606486
R11427 VSS.n5496 VSS.n5495 0.000606486
R11428 VSS.n5516 VSS.n5515 0.000606486
R11429 VSS.n5518 VSS.n5517 0.000606486
R11430 VSS.n5510 VSS.n5509 0.000606486
R11431 VSS.n5512 VSS.n5511 0.000606486
R11432 VSS.n5527 VSS.n5490 0.000606486
R11433 VSS.n5528 VSS.n5489 0.000606486
R11434 VSS.n6235 VSS.n6234 0.000606486
R11435 VSS.n2069 VSS.n2025 0.000606486
R11436 VSS.n2067 VSS.n2026 0.000606486
R11437 VSS.n2065 VSS.n2036 0.000606486
R11438 VSS.n2063 VSS.n2037 0.000606486
R11439 VSS.n2061 VSS.n2060 0.000606486
R11440 VSS.n5956 VSS.n5955 0.000606486
R11441 VSS.n5919 VSS.n2006 0.000606486
R11442 VSS.n5987 VSS.n1952 0.000606486
R11443 VSS.n5988 VSS.n1959 0.000606486
R11444 VSS.n5986 VSS.n1958 0.000606486
R11445 VSS.n5985 VSS.n5984 0.000606486
R11446 VSS.n5920 VSS.n1963 0.000606486
R11447 VSS.n1968 VSS.n1967 0.000606486
R11448 VSS.n5969 VSS.n5968 0.000606486
R11449 VSS.n5967 VSS.n5966 0.000606486
R11450 VSS.n5963 VSS.n5962 0.000606486
R11451 VSS.n2046 VSS.n2045 0.000606486
R11452 VSS.n2052 VSS.n2044 0.000606486
R11453 VSS.n2051 VSS.n2050 0.000606486
R11454 VSS.n6233 VSS.n1903 0.000606486
R11455 VSS.n6006 VSS.n6005 0.000606486
R11456 VSS.n6010 VSS.n6009 0.000606486
R11457 VSS.n6012 VSS.n6011 0.000606486
R11458 VSS.n1947 VSS.n1946 0.000606486
R11459 VSS.n1990 VSS.n1989 0.000606486
R11460 VSS.n1977 VSS.n1918 0.000606486
R11461 VSS.n2055 VSS.n2054 0.000606486
R11462 VSS.n2058 VSS.n2042 0.000606486
R11463 VSS.n2057 VSS.n2043 0.000606486
R11464 VSS.n2041 VSS.n2039 0.000606486
R11465 VSS.n2040 VSS.n2009 0.000606486
R11466 VSS.n1980 VSS.n1979 0.000606486
R11467 VSS.n1987 VSS.n1986 0.000606486
R11468 VSS.n6221 VSS.n1920 0.000606486
R11469 VSS.n6223 VSS.n1919 0.000606486
R11470 VSS.n6217 VSS.n1924 0.000606486
R11471 VSS.n6219 VSS.n1923 0.000606486
R11472 VSS.n5960 VSS.n5959 0.000606486
R11473 VSS.n5958 VSS.n2004 0.000606486
R11474 VSS.n5951 VSS.n2007 0.000606486
R11475 VSS.n5953 VSS.n5952 0.000606486
R11476 VSS.n1996 VSS.n1993 0.000606486
R11477 VSS.n1999 VSS.n1969 0.000606486
R11478 VSS.n1998 VSS.n1970 0.000606486
R11479 VSS.n2003 VSS.n2002 0.000606486
R11480 VSS.n2001 VSS.n1922 0.000606486
R11481 VSS.n6788 VSS.n6787 0.000606486
R11482 VSS.n1973 VSS.n1972 0.000606486
R11483 VSS.n6794 VSS.n6793 0.000606486
R11484 VSS.n6792 VSS.n6791 0.000606486
R11485 VSS.n5922 VSS.n1964 0.000606486
R11486 VSS.n5923 VSS.n5917 0.000606486
R11487 VSS.n6785 VSS.n1003 0.000606486
R11488 VSS.n5973 VSS.n5972 0.000606486
R11489 VSS.n5971 VSS.n1004 0.000606486
R11490 VSS.n5977 VSS.n5976 0.000606486
R11491 VSS.n5975 VSS.n1926 0.000606486
R11492 VSS.n5982 VSS.n1965 0.000606486
R11493 VSS.n5981 VSS.n5980 0.000606486
R11494 VSS.n6213 VSS.n1928 0.000606486
R11495 VSS.n6215 VSS.n1927 0.000606486
R11496 VSS.n6209 VSS.n1931 0.000606486
R11497 VSS.n6210 VSS.n1930 0.000606486
R11498 VSS.n5991 VSS.n5990 0.000606486
R11499 VSS.n5943 VSS.n1960 0.000606486
R11500 VSS.n6797 VSS.n6796 0.000606486
R11501 VSS.n6000 VSS.n1929 0.000606486
R11502 VSS.n5999 VSS.n5998 0.000606486
R11503 VSS.n6003 VSS.n1956 0.000606486
R11504 VSS.n6002 VSS.n5997 0.000606486
R11505 VSS.n5994 VSS.n5993 0.000606486
R11506 VSS.n5996 VSS.n5995 0.000606486
R11507 VSS.n1938 VSS.n1937 0.000606486
R11508 VSS.n1936 VSS.n1935 0.000606486
R11509 VSS.n1944 VSS.n1939 0.000606486
R11510 VSS.n6202 VSS.n1941 0.000606486
R11511 VSS.n6207 VSS.n1933 0.000606486
R11512 VSS.n6205 VSS.n1934 0.000606486
R11513 VSS.n6018 VSS.n6014 0.000606486
R11514 VSS.n6017 VSS.n6016 0.000606486
R11515 VSS.n6024 VSS.n6023 0.000606486
R11516 VSS.n6022 VSS.n1954 0.000606486
R11517 VSS.n6029 VSS.n1950 0.000606486
R11518 VSS.n6027 VSS.n6026 0.000606486
R11519 VSS.n5930 VSS.n1951 0.000606486
R11520 VSS.n6031 VSS.n6030 0.000606486
R11521 VSS.n6039 VSS.n6038 0.000606486
R11522 VSS.n6045 VSS.n6044 0.000606486
R11523 VSS.n6051 VSS.n6050 0.000606486
R11524 VSS.n6201 VSS.n1942 0.000606486
R11525 VSS.n6798 VSS.n961 0.000606486
R11526 VSS.n6784 VSS.n1005 0.000606486
R11527 VSS.n1995 VSS.n1008 0.000606486
R11528 VSS.n6772 VSS.n6771 0.000606486
R11529 VSS.n1975 VSS.n1012 0.000606486
R11530 VSS.n1984 VSS.n1983 0.000606486
R11531 VSS.n1982 VSS.n1981 0.000606486
R11532 VSS.n1906 VSS.n1021 0.000606486
R11533 VSS.n6227 VSS.n1915 0.000606486
R11534 VSS.n6225 VSS.n1916 0.000606486
R11535 VSS.n1911 VSS.n1910 0.000606486
R11536 VSS.n1913 VSS.n1912 0.000606486
R11537 VSS.n6231 VSS.n1904 0.000606486
R11538 VSS.n6229 VSS.n1905 0.000606486
R11539 VSS.n2033 VSS.n2032 0.000606486
R11540 VSS.n2034 VSS.n2031 0.000606486
R11541 VSS.n2029 VSS.n2011 0.000606486
R11542 VSS.n2030 VSS.n2028 0.000606486
R11543 VSS.n6762 VSS.n6761 0.000606486
R11544 VSS.n6765 VSS.n6764 0.000606486
R11545 VSS.n6738 VSS.n6737 0.000606486
R11546 VSS.n6740 VSS.n6736 0.000606486
R11547 VSS.n6757 VSS.n6756 0.000606486
R11548 VSS.n6759 VSS.n6758 0.000606486
R11549 VSS.n6604 VSS.n6603 0.000606486
R11550 VSS.n6598 VSS.n6597 0.000606486
R11551 VSS.n6752 VSS.n6751 0.000606486
R11552 VSS.n6754 VSS.n6753 0.000606486
R11553 VSS.n6749 VSS.n6748 0.000606486
R11554 VSS.n6237 VSS.n6236 0.000606486
R11555 VSS.n2023 VSS.n2022 0.000606486
R11556 VSS.n6240 VSS.n6239 0.000606486
R11557 VSS.n2021 VSS.n2019 0.000606486
R11558 VSS.n2020 VSS.n2013 0.000606486
R11559 VSS.n2072 VSS.n2016 0.000606486
R11560 VSS.n2071 VSS.n2017 0.000606486
R11561 VSS.n2085 VSS.n2082 0.000606486
R11562 VSS.n2084 VSS.n2083 0.000606486
R11563 VSS.n5883 VSS.n5882 0.000606486
R11564 VSS.n5881 VSS.n5880 0.000606486
R11565 VSS.n2196 VSS.n2195 0.000594191
R11566 VSS.n2200 VSS.n2197 0.000593164
R11567 VSS.n6312 VSS.n6311 0.000578781
R11568 VSS.n6311 VSS.n6310 0.000578781
R11569 VSS.n2189 VSS.n2188 0.000578781
R11570 VSS.n2188 VSS.n2187 0.000578781
R11571 VSS.n2193 VSS.n2190 0.000560257
R11572 VSS.n2193 VSS.n2192 0.000560257
R11573 VSS.n2192 VSS.n2191 0.000560257
R11574 VSS.n6303 VSS.n1027 0.000539391
R11575 VSS.n6304 VSS.n6303 0.000539391
R11576 VSS.n6259 VSS.n6258 0.000539391
R11577 VSS.n6258 VSS.n6257 0.000539391
R11578 VSS.n6255 VSS.n1894 0.000539391
R11579 VSS.n6256 VSS.n6255 0.000539391
R11580 VSS.n1026 VSS.n1025 0.000539391
R11581 VSS.n1025 VSS.n1024 0.000539391
R11582 VSS.n6720 VSS.n6719 0.000539391
R11583 VSS.n6719 VSS.n6718 0.000539391
R11584 VSS.n6723 VSS.n6722 0.000539391
R11585 VSS.n6722 VSS.n6721 0.000539391
R11586 VSS.n6732 VSS.n6731 0.000539391
R11587 VSS.n6733 VSS.n6732 0.000539391
R11588 VSS.n6730 VSS.n6729 0.000539391
R11589 VSS.n6729 VSS.n6728 0.000539391
R11590 VSS.n6726 VSS.n6725 0.000539391
R11591 VSS.n6725 VSS.n6724 0.000539391
R11592 VSS.n2095 VSS.n2094 0.000539391
R11593 VSS.n2126 VSS.n2125 0.000539391
R11594 VSS.n2125 VSS.n2124 0.000539391
R11595 VSS.n2129 VSS.n2128 0.000539391
R11596 VSS.n2128 VSS.n2127 0.000539391
R11597 VSS.n2094 VSS.n2093 0.000539391
R11598 VSS.n5859 VSS.n5858 0.000539391
R11599 VSS.t88 VSS.n5859 0.000539391
R11600 VSS.n5857 VSS.n5856 0.000539391
R11601 VSS.n5856 VSS.n5855 0.000539391
R11602 VSS.n5852 VSS.n2096 0.000539391
R11603 VSS.n5853 VSS.n5852 0.000539391
R11604 VSS.n5850 VSS.n5849 0.000539391
R11605 VSS.n5851 VSS.n5850 0.000539391
R11606 VSS.n5848 VSS.n5847 0.000539391
R11607 VSS.n5847 VSS.n5846 0.000539391
R11608 VSS.n5844 VSS.n5843 0.000539391
R11609 VSS.n5843 VSS.n5842 0.000539391
R11610 VSS.n5841 VSS.n5840 0.000539391
R11611 VSS.n5840 VSS.n5839 0.000539391
R11612 VSS.n2100 VSS.n2099 0.000539391
R11613 VSS.n2099 VSS.n2098 0.000539391
R11614 VSS.n2179 VSS.n2178 0.000539391
R11615 VSS.n2180 VSS.n2179 0.000539391
R11616 VSS.n2116 VSS.n2115 0.000539391
R11617 VSS.n2115 VSS.n2114 0.000539391
R11618 VSS.n2207 VSS.n2206 0.000539391
R11619 VSS.n2206 VSS.n2205 0.000539391
R11620 VSS.n2204 VSS.n2203 0.000539391
R11621 VSS.n2203 VSS.n2202 0.000539391
R11622 VSS.n1881 VSS.n1880 0.000539391
R11623 VSS.n1880 VSS.n1879 0.000539391
R11624 VSS.n1884 VSS.n1883 0.000539391
R11625 VSS.n1883 VSS.n1882 0.000539391
R11626 VSS.n1869 VSS.n1868 0.000539391
R11627 VSS.n1868 VSS.n1867 0.000539391
R11628 VSS.n2257 VSS.n2256 0.000539391
R11629 VSS.n2254 VSS.n2253 0.000539391
R11630 VSS.n6262 VSS.n6261 0.000539391
R11631 VSS.n6261 VSS.n6260 0.000539391
R11632 VSS.n2251 VSS.n2250 0.000539391
R11633 VSS.n2250 VSS.n2249 0.000539391
R11634 VSS.n5861 VSS.n1893 0.000539391
R11635 VSS.n5862 VSS.n5861 0.000539391
R11636 VSS.n7543 VSS.n300 0.000533349
R11637 VSS.n2754 VSS.n2753 0.000533349
R11638 VSS.n7543 VSS.n7542 0.000533349
R11639 VSS.n2757 VSS.n2720 0.000533349
R11640 VSS.n2760 VSS.n2757 0.000533349
R11641 VSS.n5642 VSS.n2501 0.000533349
R11642 VSS.n4422 VSS.n4421 0.000533349
R11643 VSS.n4519 VSS.n4392 0.000533349
R11644 VSS.n4519 VSS.n4518 0.000533349
R11645 VSS.n4563 VSS.n4385 0.000533349
R11646 VSS.n4564 VSS.n4563 0.000533349
R11647 VSS.n5024 VSS.n4180 0.000533349
R11648 VSS.n5024 VSS.n5023 0.000533349
R11649 VSS.n5046 VSS.n4173 0.000533349
R11650 VSS.n5046 VSS.n5045 0.000533349
R11651 VSS.n5062 VSS.n5061 0.000533349
R11652 VSS.n5062 VSS.n4166 0.000533349
R11653 VSS.n5073 VSS.n5072 0.000533349
R11654 VSS.n5652 VSS.n2447 0.000533349
R11655 VSS.n5653 VSS.n5652 0.000533349
R11656 VSS.n5648 VSS.n5647 0.000533349
R11657 VSS.n5648 VSS.n2474 0.000533349
R11658 VSS.n5081 VSS.n5080 0.000533349
R11659 VSS.n5082 VSS.n5081 0.000533349
R11660 VSS.n5069 VSS.n5068 0.000533349
R11661 VSS.n5069 VSS.n4164 0.000533349
R11662 VSS.n5053 VSS.n5052 0.000533349
R11663 VSS.n5053 VSS.n4168 0.000533349
R11664 VSS.n5031 VSS.n5030 0.000533349
R11665 VSS.n5031 VSS.n4175 0.000533349
R11666 VSS.n4559 VSS.n4558 0.000533349
R11667 VSS.n4559 VSS.n4554 0.000533349
R11668 VSS.n4526 VSS.n4525 0.000533349
R11669 VSS.n4526 VSS.n4387 0.000533349
R11670 VSS.n7508 VSS.n7507 0.000533349
R11671 VSS.n542 VSS.n541 0.000533349
R11672 VSS.n444 VSS.n443 0.000533349
R11673 VSS.n359 VSS.n356 0.000533349
R11674 VSS.n485 VSS.n470 0.000533349
R11675 VSS.n360 VSS.n359 0.000533349
R11676 VSS.n485 VSS.n484 0.000533349
R11677 VSS.n255 VSS.n249 0.000533349
R11678 VSS.n7310 VSS.n7295 0.000533349
R11679 VSS.n255 VSS.n254 0.000533349
R11680 VSS.n7310 VSS.n7309 0.000533349
R11681 VSS.n7273 VSS.n7270 0.000533349
R11682 VSS.n7274 VSS.n7273 0.000533349
R11683 VSS.n265 VSS.n264 0.000533349
R11684 VSS.n212 VSS.n209 0.000533349
R11685 VSS.n7562 VSS.n108 0.000533349
R11686 VSS.n7562 VSS.n7561 0.000533349
R11687 VSS.n213 VSS.n212 0.000533349
R11688 VSS.n159 VSS.n135 0.000533349
R11689 VSS.n159 VSS.n158 0.000533349
R11690 VSS.n6188 VSS.n6187 0.000533349
R11691 VSS.n6182 VSS.n6181 0.000533349
R11692 VSS.n1319 VSS.n1300 0.000533349
R11693 VSS.n6393 VSS.n6392 0.000533349
R11694 VSS.n6467 VSS.n6466 0.000533349
R11695 VSS.n6548 VSS.n6547 0.000533349
R11696 VSS.n6702 VSS.n6701 0.000533349
R11697 VSS.n6124 VSS.n6122 0.000533349
R11698 VSS.n981 VSS.n975 0.000533349
R11699 VSS.n1254 VSS.n1226 0.000533349
R11700 VSS.n6365 VSS.n6364 0.000533349
R11701 VSS.n6508 VSS.n1138 0.000533349
R11702 VSS.n6575 VSS.n1104 0.000533349
R11703 VSS.n6648 VSS.n6647 0.000533349
R11704 VSS.n6633 VSS.n6624 0.000533349
R11705 VSS.n6826 VSS.n6825 0.000533349
R11706 VSS.n6827 VSS.n6826 0.000533349
R11707 VSS.n7756 VSS.n7755 0.000533349
R11708 VSS.n6334 VSS.n6333 0.000533349
R11709 VSS.n6343 VSS.n6334 0.000533349
R11710 VSS.n5390 VSS.n5384 0.000533349
R11711 VSS.n5413 VSS.n5390 0.000533349
R11712 VSS.n3858 VSS.n3857 0.000533349
R11713 VSS.n5471 VSS.n5465 0.000533349
R11714 VSS.n3334 VSS.n3328 0.000533349
R11715 VSS.n3431 VSS.n3425 0.000533349
R11716 VSS.n3528 VSS.n3522 0.000533349
R11717 VSS.n3625 VSS.n3619 0.000533349
R11718 VSS.n3723 VSS.n3717 0.000533349
R11719 VSS.n3820 VSS.n3814 0.000533349
R11720 VSS.n3760 VSS.n3759 0.000533349
R11721 VSS.n3662 VSS.n3661 0.000533349
R11722 VSS.n2894 VSS.n2888 0.000533349
R11723 VSS.n3564 VSS.n2894 0.000533349
R11724 VSS.n2905 VSS.n2899 0.000533349
R11725 VSS.n3467 VSS.n2905 0.000533349
R11726 VSS.n2917 VSS.n2911 0.000533349
R11727 VSS.n3370 VSS.n2917 0.000533349
R11728 VSS.n3316 VSS.n2809 0.000533349
R11729 VSS.n5360 VSS.n2809 0.000533349
R11730 VSS.n5822 VSS.n5814 0.000533349
R11731 VSS.n5600 VSS.n5599 0.000516685
R11732 VSS.n2764 VSS.n2715 0.000516685
R11733 VSS.n2765 VSS.n2764 0.000516685
R11734 VSS.n5641 VSS.n5640 0.000516685
R11735 VSS.n5638 VSS.n5634 0.000516685
R11736 VSS.n5634 VSS.n5629 0.000516685
R11737 VSS.n5634 VSS.n5633 0.000516685
R11738 VSS.n5599 VSS.n5598 0.000516685
R11739 VSS.n2764 VSS.n2763 0.000516685
R11740 VSS.n2200 VSS.n2199 0.000516018
R11741 VSS.n2219 VSS.n2201 0.000516018
R11742 VSS.n6319 VSS.n6314 0.000513139
R11743 VSS.n5595 VSS.n5594 0.000511116
R11744 VSS.n5576 VSS.n5575 0.000511116
R11745 VSS.n5570 VSS.n5569 0.000511116
R11746 VSS.n5568 VSS.n5567 0.000511116
R11747 VSS.n2768 VSS.n2767 0.000511116
R11748 VSS.n3840 VSS.n3839 0.000511116
R11749 VSS.n3838 VSS.n3837 0.000511116
R11750 VSS.n3824 VSS.n3823 0.000511116
R11751 VSS.n3757 VSS.n3756 0.000511116
R11752 VSS.n3743 VSS.n3742 0.000511116
R11753 VSS.n3741 VSS.n3740 0.000511116
R11754 VSS.n3727 VSS.n3726 0.000511116
R11755 VSS.n3659 VSS.n3658 0.000511116
R11756 VSS.n3645 VSS.n3644 0.000511116
R11757 VSS.n3643 VSS.n3642 0.000511116
R11758 VSS.n3629 VSS.n3628 0.000511116
R11759 VSS.n3562 VSS.n3561 0.000511116
R11760 VSS.n3548 VSS.n3547 0.000511116
R11761 VSS.n3546 VSS.n3545 0.000511116
R11762 VSS.n3532 VSS.n3531 0.000511116
R11763 VSS.n3465 VSS.n3464 0.000511116
R11764 VSS.n3451 VSS.n3450 0.000511116
R11765 VSS.n3449 VSS.n3448 0.000511116
R11766 VSS.n3435 VSS.n3434 0.000511116
R11767 VSS.n3368 VSS.n3367 0.000511116
R11768 VSS.n3354 VSS.n3353 0.000511116
R11769 VSS.n3352 VSS.n3351 0.000511116
R11770 VSS.n3338 VSS.n3337 0.000511116
R11771 VSS.n5362 VSS.n5361 0.000511116
R11772 VSS.n5376 VSS.n5375 0.000511116
R11773 VSS.n5378 VSS.n5377 0.000511116
R11774 VSS.n5475 VSS.n5474 0.000511116
R11775 VSS.n5411 VSS.n5410 0.000511116
R11776 VSS.n5397 VSS.n5396 0.000511116
R11777 VSS.n5395 VSS.n5394 0.000511116
R11778 VSS.n5826 VSS.n5825 0.000511116
R11779 VSS.n6707 VSS.n6706 0.000511116
R11780 VSS.n1056 VSS.n1055 0.000511116
R11781 VSS.n1047 VSS.n1046 0.000511116
R11782 VSS.n6061 VSS.n6060 0.000511116
R11783 VSS.n6071 VSS.n6070 0.000511116
R11784 VSS.n6078 VSS.n6077 0.000511116
R11785 VSS.n6190 VSS.n6189 0.000511116
R11786 VSS.n6121 VSS.n6120 0.000511116
R11787 VSS.n6112 VSS.n6111 0.000511116
R11788 VSS.n6806 VSS.n6805 0.000511116
R11789 VSS.n6822 VSS.n6821 0.000511116
R11790 VSS.n985 VSS.n984 0.000511116
R11791 VSS.n995 VSS.n994 0.000511116
R11792 VSS.n1302 VSS.n1301 0.000511116
R11793 VSS.n1318 VSS.n1317 0.000511116
R11794 VSS.n1251 VSS.n1250 0.000511116
R11795 VSS.n1242 VSS.n1241 0.000511116
R11796 VSS.n6376 VSS.n6375 0.000511116
R11797 VSS.n6391 VSS.n6390 0.000511116
R11798 VSS.n6436 VSS.n6435 0.000511116
R11799 VSS.n6445 VSS.n6444 0.000511116
R11800 VSS.n6447 VSS.n6446 0.000511116
R11801 VSS.n6461 VSS.n6460 0.000511116
R11802 VSS.n6512 VSS.n6511 0.000511116
R11803 VSS.n6528 VSS.n6527 0.000511116
R11804 VSS.n6530 VSS.n6529 0.000511116
R11805 VSS.n6546 VSS.n6545 0.000511116
R11806 VSS.n6579 VSS.n6578 0.000511116
R11807 VSS.n6589 VSS.n6588 0.000511116
R11808 VSS.n6608 VSS.n6607 0.000511116
R11809 VSS.n6623 VSS.n6622 0.000511116
R11810 VSS.n6704 VSS.n6703 0.000511116
R11811 VSS.n3854 VSS.n3853 0.000511116
R11812 VSS.n5581 VSS.n5580 0.000511116
R11813 VSS.n3846 VSS.n3845 0.000511116
R11814 VSS.n3830 VSS.n3829 0.000511116
R11815 VSS.n3749 VSS.n3748 0.000511116
R11816 VSS.n3733 VSS.n3732 0.000511116
R11817 VSS.n3651 VSS.n3650 0.000511116
R11818 VSS.n3635 VSS.n3634 0.000511116
R11819 VSS.n3554 VSS.n3553 0.000511116
R11820 VSS.n3538 VSS.n3537 0.000511116
R11821 VSS.n3457 VSS.n3456 0.000511116
R11822 VSS.n3441 VSS.n3440 0.000511116
R11823 VSS.n3360 VSS.n3359 0.000511116
R11824 VSS.n3344 VSS.n3343 0.000511116
R11825 VSS.n5368 VSS.n5367 0.000511116
R11826 VSS.n5481 VSS.n5480 0.000511116
R11827 VSS.n5403 VSS.n5402 0.000511116
R11828 VSS.n5832 VSS.n5831 0.000511116
R11829 VSS.n6067 VSS.n6066 0.000511116
R11830 VSS.n6084 VSS.n6083 0.000511116
R11831 VSS.n6107 VSS.n6106 0.000511116
R11832 VSS.n6812 VSS.n6811 0.000511116
R11833 VSS.n991 VSS.n990 0.000511116
R11834 VSS.n1308 VSS.n1307 0.000511116
R11835 VSS.n1238 VSS.n1237 0.000511116
R11836 VSS.n6382 VSS.n6381 0.000511116
R11837 VSS.n1151 VSS.n1150 0.000511116
R11838 VSS.n6453 VSS.n6452 0.000511116
R11839 VSS.n6520 VSS.n6519 0.000511116
R11840 VSS.n6538 VSS.n6537 0.000511116
R11841 VSS.n6585 VSS.n6584 0.000511116
R11842 VSS.n6615 VSS.n6614 0.000511116
R11843 VSS.n1042 VSS.n1041 0.000511116
R11844 VSS.n1032 VSS.n1031 0.000511116
R11845 VSS.n1878 VSS.n1870 0.000509989
R11846 VSS.n1878 VSS.n1877 0.000507583
R11847 VSS.n6319 VSS.n6318 0.000506803
R11848 VSS.n6318 VSS.n6317 0.000506803
R11849 VSS.n2239 VSS.n2238 0.000505632
R11850 VSS.n2358 VSS.n2357 0.000505632
R11851 VSS.n2110 VSS.n2109 0.000505632
R11852 VSS.n2233 VSS.n2232 0.000505632
R11853 VSS.n6324 VSS.n6323 0.000505632
R11854 VSS.n6329 VSS.n6328 0.000505632
R11855 VSS.n5640 VSS.n5639 0.000505597
R11856 VSS.n5633 VSS.n5632 0.000505597
R11857 VSS.n2715 VSS.n2714 0.000505597
R11858 VSS.n5602 VSS.n5600 0.000505597
R11859 VSS.n2505 VSS.n2504 0.000505597
R11860 VSS.n5638 VSS.n5637 0.000505597
R11861 VSS.n5629 VSS.n5628 0.000505597
R11862 VSS.n5565 VSS.n5564 0.000505094
R11863 VSS.n999 VSS.n993 0.000505094
R11864 VSS.n999 VSS.n998 0.000505094
R11865 VSS.n6593 VSS.n6587 0.000505094
R11866 VSS.n6593 VSS.n6592 0.000505094
R11867 VSS.n6620 VSS.n6612 0.000505094
R11868 VSS.n1051 VSS.n1044 0.000505094
R11869 VSS.n1051 VSS.n1050 0.000505094
R11870 VSS.n6710 VSS.n6709 0.000505094
R11871 VSS.n6711 VSS.n1036 0.000505094
R11872 VSS.n6711 VSS.n6710 0.000505094
R11873 VSS.n3849 VSS.n3848 0.000505094
R11874 VSS.n3851 VSS.n3849 0.000505094
R11875 VSS.n3833 VSS.n3832 0.000505094
R11876 VSS.n3835 VSS.n3833 0.000505094
R11877 VSS.n3835 VSS.n3834 0.000505094
R11878 VSS.n3444 VSS.n3443 0.000505094
R11879 VSS.n3446 VSS.n3444 0.000505094
R11880 VSS.n3446 VSS.n3445 0.000505094
R11881 VSS.n5835 VSS.n5834 0.000505094
R11882 VSS.n5835 VSS.n2103 0.000505094
R11883 VSS.n2103 VSS.n2102 0.000505094
R11884 VSS.n5406 VSS.n5405 0.000505094
R11885 VSS.n5408 VSS.n5406 0.000505094
R11886 VSS.n5408 VSS.n5407 0.000505094
R11887 VSS.n5484 VSS.n5483 0.000505094
R11888 VSS.n5484 VSS.n5381 0.000505094
R11889 VSS.n5381 VSS.n5380 0.000505094
R11890 VSS.n5371 VSS.n5370 0.000505094
R11891 VSS.n5371 VSS.n5365 0.000505094
R11892 VSS.n5365 VSS.n5364 0.000505094
R11893 VSS.n3347 VSS.n3346 0.000505094
R11894 VSS.n3349 VSS.n3347 0.000505094
R11895 VSS.n3349 VSS.n3348 0.000505094
R11896 VSS.n3363 VSS.n3362 0.000505094
R11897 VSS.n3365 VSS.n3363 0.000505094
R11898 VSS.n3365 VSS.n3364 0.000505094
R11899 VSS.n3460 VSS.n3459 0.000505094
R11900 VSS.n3462 VSS.n3460 0.000505094
R11901 VSS.n3462 VSS.n3461 0.000505094
R11902 VSS.n3541 VSS.n3540 0.000505094
R11903 VSS.n3543 VSS.n3541 0.000505094
R11904 VSS.n3543 VSS.n3542 0.000505094
R11905 VSS.n3557 VSS.n3556 0.000505094
R11906 VSS.n3559 VSS.n3557 0.000505094
R11907 VSS.n3559 VSS.n3558 0.000505094
R11908 VSS.n3638 VSS.n3637 0.000505094
R11909 VSS.n3640 VSS.n3638 0.000505094
R11910 VSS.n3640 VSS.n3639 0.000505094
R11911 VSS.n3654 VSS.n3653 0.000505094
R11912 VSS.n3656 VSS.n3654 0.000505094
R11913 VSS.n3656 VSS.n3655 0.000505094
R11914 VSS.n3736 VSS.n3735 0.000505094
R11915 VSS.n3738 VSS.n3736 0.000505094
R11916 VSS.n3738 VSS.n3737 0.000505094
R11917 VSS.n3752 VSS.n3751 0.000505094
R11918 VSS.n3754 VSS.n3752 0.000505094
R11919 VSS.n3754 VSS.n3753 0.000505094
R11920 VSS.n6525 VSS.n6516 0.000505094
R11921 VSS.n6543 VSS.n6534 0.000505094
R11922 VSS.n6075 VSS.n6069 0.000505094
R11923 VSS.n6075 VSS.n6074 0.000505094
R11924 VSS.n6194 VSS.n6086 0.000505094
R11925 VSS.n6194 VSS.n6193 0.000505094
R11926 VSS.n6116 VSS.n6109 0.000505094
R11927 VSS.n6116 VSS.n6115 0.000505094
R11928 VSS.n6815 VSS.n6814 0.000505094
R11929 VSS.n6819 VSS.n6815 0.000505094
R11930 VSS.n1311 VSS.n1310 0.000505094
R11931 VSS.n1315 VSS.n1311 0.000505094
R11932 VSS.n1246 VSS.n1240 0.000505094
R11933 VSS.n1246 VSS.n1245 0.000505094
R11934 VSS.n6385 VSS.n6384 0.000505094
R11935 VSS.n6388 VSS.n6385 0.000505094
R11936 VSS.n6442 VSS.n6440 0.000505094
R11937 VSS.n6456 VSS.n6455 0.000505094
R11938 VSS.n6458 VSS.n6456 0.000505094
R11939 VSS.n5578 VSS.n5574 0.000505094
R11940 VSS.n6346 VSS.n6345 0.00050467
R11941 VSS.n3864 VSS.n3863 0.00050467
R11942 VSS.n5056 VSS.n5055 0.00050467
R11943 VSS.n4425 VSS.n4424 0.00050467
R11944 VSS.n4394 VSS.n4393 0.00050467
R11945 VSS.n4529 VSS.n4528 0.00050467
R11946 VSS.n4182 VSS.n4181 0.00050467
R11947 VSS.n5034 VSS.n5033 0.00050467
R11948 VSS.n4161 VSS.n4160 0.00050467
R11949 VSS.n2449 VSS.n2448 0.00050467
R11950 VSS.n3812 VSS.n3811 0.00050467
R11951 VSS.n3766 VSS.n3765 0.00050467
R11952 VSS.n3715 VSS.n3714 0.00050467
R11953 VSS.n3668 VSS.n3667 0.00050467
R11954 VSS.n3617 VSS.n3616 0.00050467
R11955 VSS.n3570 VSS.n3569 0.00050467
R11956 VSS.n3520 VSS.n3519 0.00050467
R11957 VSS.n3473 VSS.n3472 0.00050467
R11958 VSS.n3423 VSS.n3422 0.00050467
R11959 VSS.n3376 VSS.n3375 0.00050467
R11960 VSS.n3326 VSS.n3325 0.00050467
R11961 VSS.n5357 VSS.n5356 0.00050467
R11962 VSS.n5463 VSS.n5462 0.00050467
R11963 VSS.n5812 VSS.n5811 0.00050467
R11964 VSS.n5419 VSS.n5418 0.00050467
R11965 VSS.n6340 VSS.n6339 0.00050467
R11966 VSS.n2760 VSS.n2759 0.00050467
R11967 VSS.n2750 VSS.n2749 0.00050467
R11968 VSS.n545 VSS.n544 0.00050467
R11969 VSS.n447 VSS.n446 0.00050467
R11970 VSS.n7542 VSS.n7541 0.00050467
R11971 VSS.n2747 VSS.n2745 0.00050467
R11972 VSS.n297 VSS.n296 0.00050467
R11973 VSS.n2718 VSS.n2717 0.00050467
R11974 VSS.n4429 VSS.n4428 0.00050467
R11975 VSS.n4392 VSS.n4391 0.00050467
R11976 VSS.n4518 VSS.n4517 0.00050467
R11977 VSS.n4385 VSS.n4384 0.00050467
R11978 VSS.n4565 VSS.n4564 0.00050467
R11979 VSS.n4180 VSS.n4179 0.00050467
R11980 VSS.n5023 VSS.n5022 0.00050467
R11981 VSS.n4173 VSS.n4172 0.00050467
R11982 VSS.n5045 VSS.n5044 0.00050467
R11983 VSS.n5061 VSS.n5060 0.00050467
R11984 VSS.n4851 VSS.n4166 0.00050467
R11985 VSS.n4158 VSS.n4157 0.00050467
R11986 VSS.n2447 VSS.n2446 0.00050467
R11987 VSS.n5654 VSS.n5653 0.00050467
R11988 VSS.n5647 VSS.n5646 0.00050467
R11989 VSS.n2474 VSS.n2473 0.00050467
R11990 VSS.n5080 VSS.n5079 0.00050467
R11991 VSS.n5083 VSS.n5082 0.00050467
R11992 VSS.n5068 VSS.n5067 0.00050467
R11993 VSS.n4872 VSS.n4164 0.00050467
R11994 VSS.n5052 VSS.n5051 0.00050467
R11995 VSS.n4753 VSS.n4168 0.00050467
R11996 VSS.n5030 VSS.n5029 0.00050467
R11997 VSS.n5009 VSS.n4175 0.00050467
R11998 VSS.n4558 VSS.n4557 0.00050467
R11999 VSS.n4554 VSS.n4553 0.00050467
R12000 VSS.n4525 VSS.n4524 0.00050467
R12001 VSS.n4504 VSS.n4387 0.00050467
R12002 VSS.n2499 VSS.n2498 0.00050467
R12003 VSS.n2495 VSS.n2494 0.00050467
R12004 VSS.n549 VSS.n548 0.00050467
R12005 VSS.n7521 VSS.n7520 0.00050467
R12006 VSS.n7526 VSS.n7525 0.00050467
R12007 VSS.n451 VSS.n450 0.00050467
R12008 VSS.n570 VSS.n569 0.00050467
R12009 VSS.n586 VSS.n585 0.00050467
R12010 VSS.n356 VSS.n355 0.00050467
R12011 VSS.n488 VSS.n487 0.00050467
R12012 VSS.n484 VSS.n483 0.00050467
R12013 VSS.n361 VSS.n360 0.00050467
R12014 VSS.n349 VSS.n348 0.00050467
R12015 VSS.n7267 VSS.n7266 0.00050467
R12016 VSS.n246 VSS.n245 0.00050467
R12017 VSS.n254 VSS.n253 0.00050467
R12018 VSS.n7275 VSS.n7274 0.00050467
R12019 VSS.n270 VSS.n269 0.00050467
R12020 VSS.n264 VSS.n263 0.00050467
R12021 VSS.n207 VSS.n206 0.00050467
R12022 VSS.n214 VSS.n213 0.00050467
R12023 VSS.n7561 VSS.n7560 0.00050467
R12024 VSS.n7565 VSS.n7564 0.00050467
R12025 VSS.n7309 VSS.n7308 0.00050467
R12026 VSS.n7313 VSS.n7312 0.00050467
R12027 VSS.n6651 VSS.n6650 0.00050467
R12028 VSS.n6627 VSS.n6626 0.00050467
R12029 VSS.n1102 VSS.n1101 0.00050467
R12030 VSS.n6549 VSS.n6548 0.00050467
R12031 VSS.n1129 VSS.n1128 0.00050467
R12032 VSS.n6468 VSS.n6467 0.00050467
R12033 VSS.n6428 VSS.n6427 0.00050467
R12034 VSS.n6394 VSS.n6393 0.00050467
R12035 VSS.n1224 VSS.n1223 0.00050467
R12036 VSS.n1300 VSS.n1299 0.00050467
R12037 VSS.n973 VSS.n972 0.00050467
R12038 VSS.n6832 VSS.n6831 0.00050467
R12039 VSS.n6137 VSS.n6135 0.00050467
R12040 VSS.n11 VSS.n10 0.00050467
R12041 VSS.n132 VSS.n131 0.00050467
R12042 VSS.n158 VSS.n157 0.00050467
R12043 VSS.n169 VSS.n168 0.00050467
R12044 VSS.n228 VSS.n227 0.00050467
R12045 VSS.n6181 VSS.n6180 0.00050467
R12046 VSS.n6185 VSS.n6184 0.00050467
R12047 VSS.n6124 VSS.n6123 0.00050467
R12048 VSS.n6133 VSS.n6132 0.00050467
R12049 VSS.n981 VSS.n980 0.00050467
R12050 VSS.n970 VSS.n969 0.00050467
R12051 VSS.n1255 VSS.n1254 0.00050467
R12052 VSS.n1221 VSS.n1220 0.00050467
R12053 VSS.n6364 VSS.n1156 0.00050467
R12054 VSS.n6431 VSS.n6430 0.00050467
R12055 VSS.n6508 VSS.n6507 0.00050467
R12056 VSS.n1136 VSS.n1135 0.00050467
R12057 VSS.n6575 VSS.n6574 0.00050467
R12058 VSS.n1096 VSS.n1095 0.00050467
R12059 VSS.n6647 VSS.n6646 0.00050467
R12060 VSS.n6655 VSS.n6654 0.00050467
R12061 VSS.n6634 VSS.n6633 0.00050467
R12062 VSS.n1346 VSS.n1345 0.00050467
R12063 VSS.n6464 VSS.n6463 0.00050467
R12064 VSS.n6370 VSS.n6369 0.00050467
R12065 VSS.n1230 VSS.n1229 0.00050467
R12066 VSS.n6825 VSS.n6824 0.00050467
R12067 VSS.n6701 VSS.n6700 0.00050467
R12068 VSS.n7755 VSS.n7754 0.00050467
R12069 VSS.n8 VSS.n7 0.00050467
R12070 VSS.n6337 VSS.n6336 0.00050467
R12071 VSS.n5416 VSS.n5415 0.00050467
R12072 VSS.n3861 VSS.n3860 0.00050467
R12073 VSS.n5460 VSS.n5459 0.00050467
R12074 VSS.n5471 VSS.n5470 0.00050467
R12075 VSS.n3323 VSS.n3322 0.00050467
R12076 VSS.n3334 VSS.n3333 0.00050467
R12077 VSS.n3420 VSS.n3419 0.00050467
R12078 VSS.n3431 VSS.n3430 0.00050467
R12079 VSS.n3517 VSS.n3516 0.00050467
R12080 VSS.n3528 VSS.n3527 0.00050467
R12081 VSS.n3614 VSS.n3613 0.00050467
R12082 VSS.n3625 VSS.n3624 0.00050467
R12083 VSS.n3712 VSS.n3711 0.00050467
R12084 VSS.n3723 VSS.n3722 0.00050467
R12085 VSS.n3809 VSS.n3808 0.00050467
R12086 VSS.n3820 VSS.n3819 0.00050467
R12087 VSS.n3763 VSS.n3762 0.00050467
R12088 VSS.n3665 VSS.n3664 0.00050467
R12089 VSS.n3567 VSS.n3566 0.00050467
R12090 VSS.n3470 VSS.n3469 0.00050467
R12091 VSS.n3373 VSS.n3372 0.00050467
R12092 VSS.n2812 VSS.n2811 0.00050467
R12093 VSS.n5809 VSS.n5808 0.00050467
R12094 VSS.n5822 VSS.n5821 0.00050467
R12095 VSS.n4851 VSS.n4850 0.000504623
R12096 VSS.n4852 VSS.n4851 0.000504623
R12097 VSS.n4517 VSS.n4398 0.000504623
R12098 VSS.n4517 VSS.n4516 0.000504623
R12099 VSS.n4565 VSS.n4380 0.000504623
R12100 VSS.n4566 VSS.n4565 0.000504623
R12101 VSS.n5022 VSS.n4186 0.000504623
R12102 VSS.n5022 VSS.n5021 0.000504623
R12103 VSS.n5044 VSS.n5038 0.000504623
R12104 VSS.n5044 VSS.n5043 0.000504623
R12105 VSS.n5654 VSS.n2442 0.000504623
R12106 VSS.n5655 VSS.n5654 0.000504623
R12107 VSS.n3808 VSS.n3807 0.000504623
R12108 VSS.n3711 VSS.n3710 0.000504623
R12109 VSS.n3613 VSS.n3612 0.000504623
R12110 VSS.n3516 VSS.n3515 0.000504623
R12111 VSS.n3419 VSS.n3418 0.000504623
R12112 VSS.n3322 VSS.n3321 0.000504623
R12113 VSS.n5459 VSS.n5458 0.000504623
R12114 VSS.n5808 VSS.n5807 0.000504623
R12115 VSS.n5821 VSS.n5820 0.000504623
R12116 VSS.n362 VSS.n361 0.000504623
R12117 VSS.n6646 VSS.n6645 0.000504623
R12118 VSS.n6574 VSS.n6573 0.000504623
R12119 VSS.n6507 VSS.n6506 0.000504623
R12120 VSS.n6421 VSS.n1156 0.000504623
R12121 VSS.n6427 VSS.n6421 0.000504623
R12122 VSS.n1256 VSS.n1255 0.000504623
R12123 VSS.n980 VSS.n979 0.000504623
R12124 VSS.n6138 VSS.n6137 0.000504623
R12125 VSS.n7754 VSS.n7753 0.000504623
R12126 VSS.n2357 VSS.n2356 0.000504168
R12127 VSS.n2232 VSS.n2231 0.000504168
R12128 VSS.n6323 VSS.n6322 0.000504168
R12129 VSS.n2504 VSS.n2503 0.000504146
R12130 VSS.n5637 VSS.n5636 0.000504146
R12131 VSS.n5628 VSS.n5627 0.000504146
R12132 VSS.n2714 VSS.n2713 0.000504146
R12133 VSS.n5603 VSS.n5602 0.000504146
R12134 VSS.n2712 VSS.n2711 0.000504146
R12135 VSS.n5571 VSS.n5570 0.000503113
R12136 VSS.n5567 VSS.n5566 0.000503113
R12137 VSS.n2769 VSS.n2768 0.000503113
R12138 VSS.n3841 VSS.n3840 0.000503113
R12139 VSS.n3837 VSS.n3836 0.000503113
R12140 VSS.n3825 VSS.n3824 0.000503113
R12141 VSS.n3756 VSS.n3755 0.000503113
R12142 VSS.n3744 VSS.n3743 0.000503113
R12143 VSS.n3740 VSS.n3739 0.000503113
R12144 VSS.n3728 VSS.n3727 0.000503113
R12145 VSS.n3658 VSS.n3657 0.000503113
R12146 VSS.n3646 VSS.n3645 0.000503113
R12147 VSS.n3642 VSS.n3641 0.000503113
R12148 VSS.n3630 VSS.n3629 0.000503113
R12149 VSS.n3561 VSS.n3560 0.000503113
R12150 VSS.n3549 VSS.n3548 0.000503113
R12151 VSS.n3545 VSS.n3544 0.000503113
R12152 VSS.n3533 VSS.n3532 0.000503113
R12153 VSS.n3464 VSS.n3463 0.000503113
R12154 VSS.n3452 VSS.n3451 0.000503113
R12155 VSS.n3448 VSS.n3447 0.000503113
R12156 VSS.n3436 VSS.n3435 0.000503113
R12157 VSS.n3367 VSS.n3366 0.000503113
R12158 VSS.n3355 VSS.n3354 0.000503113
R12159 VSS.n3351 VSS.n3350 0.000503113
R12160 VSS.n3339 VSS.n3338 0.000503113
R12161 VSS.n5363 VSS.n5362 0.000503113
R12162 VSS.n5375 VSS.n5374 0.000503113
R12163 VSS.n5379 VSS.n5378 0.000503113
R12164 VSS.n5476 VSS.n5475 0.000503113
R12165 VSS.n5410 VSS.n5409 0.000503113
R12166 VSS.n5398 VSS.n5397 0.000503113
R12167 VSS.n5394 VSS.n5393 0.000503113
R12168 VSS.n5827 VSS.n5826 0.000503113
R12169 VSS.n6708 VSS.n6707 0.000503113
R12170 VSS.n1055 VSS.n1054 0.000503113
R12171 VSS.n1048 VSS.n1047 0.000503113
R12172 VSS.n6062 VSS.n6061 0.000503113
R12173 VSS.n6072 VSS.n6071 0.000503113
R12174 VSS.n6079 VSS.n6078 0.000503113
R12175 VSS.n6191 VSS.n6190 0.000503113
R12176 VSS.n6120 VSS.n6119 0.000503113
R12177 VSS.n6113 VSS.n6112 0.000503113
R12178 VSS.n6807 VSS.n6806 0.000503113
R12179 VSS.n6821 VSS.n6820 0.000503113
R12180 VSS.n986 VSS.n985 0.000503113
R12181 VSS.n996 VSS.n995 0.000503113
R12182 VSS.n1303 VSS.n1302 0.000503113
R12183 VSS.n1317 VSS.n1316 0.000503113
R12184 VSS.n1250 VSS.n1249 0.000503113
R12185 VSS.n1243 VSS.n1242 0.000503113
R12186 VSS.n6377 VSS.n6376 0.000503113
R12187 VSS.n6390 VSS.n6389 0.000503113
R12188 VSS.n6437 VSS.n6436 0.000503113
R12189 VSS.n6444 VSS.n6443 0.000503113
R12190 VSS.n6448 VSS.n6447 0.000503113
R12191 VSS.n6460 VSS.n6459 0.000503113
R12192 VSS.n6513 VSS.n6512 0.000503113
R12193 VSS.n6527 VSS.n6526 0.000503113
R12194 VSS.n6531 VSS.n6530 0.000503113
R12195 VSS.n6545 VSS.n6544 0.000503113
R12196 VSS.n6580 VSS.n6579 0.000503113
R12197 VSS.n6590 VSS.n6589 0.000503113
R12198 VSS.n6609 VSS.n6608 0.000503113
R12199 VSS.n6622 VSS.n6621 0.000503113
R12200 VSS.n6705 VSS.n6704 0.000503113
R12201 VSS.n3853 VSS.n3852 0.000503113
R12202 VSS.n5594 VSS.n5593 0.000503113
R12203 VSS.n6454 VSS.n6453 0.000503113
R12204 VSS.n1152 VSS.n1151 0.000503113
R12205 VSS.n6383 VSS.n6382 0.000503113
R12206 VSS.n1239 VSS.n1238 0.000503113
R12207 VSS.n1309 VSS.n1308 0.000503113
R12208 VSS.n992 VSS.n991 0.000503113
R12209 VSS.n6813 VSS.n6812 0.000503113
R12210 VSS.n6108 VSS.n6107 0.000503113
R12211 VSS.n6085 VSS.n6084 0.000503113
R12212 VSS.n6068 VSS.n6067 0.000503113
R12213 VSS.n6539 VSS.n6538 0.000503113
R12214 VSS.n6521 VSS.n6520 0.000503113
R12215 VSS.n1033 VSS.n1032 0.000503113
R12216 VSS.n6616 VSS.n6615 0.000503113
R12217 VSS.n6586 VSS.n6585 0.000503113
R12218 VSS.n1043 VSS.n1042 0.000503113
R12219 VSS.n3831 VSS.n3830 0.000503113
R12220 VSS.n3847 VSS.n3846 0.000503113
R12221 VSS.n3750 VSS.n3749 0.000503113
R12222 VSS.n3734 VSS.n3733 0.000503113
R12223 VSS.n3652 VSS.n3651 0.000503113
R12224 VSS.n3636 VSS.n3635 0.000503113
R12225 VSS.n3555 VSS.n3554 0.000503113
R12226 VSS.n3539 VSS.n3538 0.000503113
R12227 VSS.n3458 VSS.n3457 0.000503113
R12228 VSS.n3442 VSS.n3441 0.000503113
R12229 VSS.n3361 VSS.n3360 0.000503113
R12230 VSS.n3345 VSS.n3344 0.000503113
R12231 VSS.n5369 VSS.n5368 0.000503113
R12232 VSS.n5482 VSS.n5481 0.000503113
R12233 VSS.n5404 VSS.n5403 0.000503113
R12234 VSS.n5833 VSS.n5832 0.000503113
R12235 VSS.n5577 VSS.n5576 0.000503113
R12236 VSS.n5582 VSS.n5581 0.000503113
R12237 VSS.n7285 VSS.n7284 0.000502702
R12238 VSS.n98 VSS.n97 0.000502702
R12239 VSS.n4999 VSS.n4998 0.000502702
R12240 VSS.n4448 VSS.n4447 0.000502702
R12241 VSS.n4540 VSS.n4539 0.000502702
R12242 VSS.n4492 VSS.n4491 0.000502702
R12243 VSS.n4618 VSS.n4617 0.000502702
R12244 VSS.n3882 VSS.n3881 0.000502702
R12245 VSS.n4311 VSS.n4310 0.000502702
R12246 VSS.n4318 VSS.n4317 0.000502702
R12247 VSS.n4650 VSS.n4649 0.000502702
R12248 VSS.n4629 VSS.n4628 0.000502702
R12249 VSS.n4959 VSS.n4958 0.000502702
R12250 VSS.n4438 VSS.n4437 0.000502702
R12251 VSS.n4862 VSS.n4861 0.000502702
R12252 VSS.n4141 VSS.n4140 0.000502702
R12253 VSS.n4759 VSS.n4758 0.000502702
R12254 VSS.n4929 VSS.n4928 0.000502702
R12255 VSS.n5161 VSS.n5160 0.000502702
R12256 VSS.n4914 VSS.n4913 0.000502702
R12257 VSS.n4132 VSS.n4131 0.000502702
R12258 VSS.n5142 VSS.n5141 0.000502702
R12259 VSS.n4830 VSS.n4829 0.000502702
R12260 VSS.n4675 VSS.n4674 0.000502702
R12261 VSS.n4247 VSS.n4246 0.000502702
R12262 VSS.n4682 VSS.n4681 0.000502702
R12263 VSS.n4696 VSS.n4695 0.000502702
R12264 VSS.n4227 VSS.n4226 0.000502702
R12265 VSS.n4708 VSS.n4707 0.000502702
R12266 VSS.n4731 VSS.n4730 0.000502702
R12267 VSS.n4712 VSS.n4711 0.000502702
R12268 VSS.n4718 VSS.n4717 0.000502702
R12269 VSS.n5204 VSS.n5203 0.000502702
R12270 VSS.n4265 VSS.n4264 0.000502702
R12271 VSS.n4039 VSS.n4038 0.000502702
R12272 VSS.n4017 VSS.n4016 0.000502702
R12273 VSS.n4026 VSS.n4025 0.000502702
R12274 VSS.n4052 VSS.n4051 0.000502702
R12275 VSS.n4022 VSS.n4021 0.000502702
R12276 VSS.n4004 VSS.n4003 0.000502702
R12277 VSS.n4064 VSS.n4063 0.000502702
R12278 VSS.n4000 VSS.n3999 0.000502702
R12279 VSS.n4077 VSS.n4076 0.000502702
R12280 VSS.n4091 VSS.n4090 0.000502702
R12281 VSS.n4072 VSS.n4071 0.000502702
R12282 VSS.n4097 VSS.n4096 0.000502702
R12283 VSS.n3968 VSS.n3967 0.000502702
R12284 VSS.n4297 VSS.n4296 0.000502702
R12285 VSS.n3778 VSS.n3777 0.000502702
R12286 VSS.n3786 VSS.n3785 0.000502702
R12287 VSS.n3692 VSS.n3691 0.000502702
R12288 VSS.n3680 VSS.n3679 0.000502702
R12289 VSS.n3688 VSS.n3687 0.000502702
R12290 VSS.n3594 VSS.n3593 0.000502702
R12291 VSS.n3582 VSS.n3581 0.000502702
R12292 VSS.n3590 VSS.n3589 0.000502702
R12293 VSS.n3497 VSS.n3496 0.000502702
R12294 VSS.n3485 VSS.n3484 0.000502702
R12295 VSS.n3493 VSS.n3492 0.000502702
R12296 VSS.n3400 VSS.n3399 0.000502702
R12297 VSS.n3388 VSS.n3387 0.000502702
R12298 VSS.n3396 VSS.n3395 0.000502702
R12299 VSS.n5338 VSS.n5337 0.000502702
R12300 VSS.n5450 VSS.n5449 0.000502702
R12301 VSS.n3873 VSS.n3872 0.000502702
R12302 VSS.n5431 VSS.n5430 0.000502702
R12303 VSS.n5438 VSS.n5437 0.000502702
R12304 VSS.n5792 VSS.n5791 0.000502702
R12305 VSS.n5774 VSS.n5773 0.000502702
R12306 VSS.n3957 VSS.n3956 0.000502702
R12307 VSS.n5760 VSS.n5759 0.000502702
R12308 VSS.n5742 VSS.n5741 0.000502702
R12309 VSS.n5193 VSS.n5192 0.000502702
R12310 VSS.n5728 VSS.n5727 0.000502702
R12311 VSS.n5710 VSS.n5709 0.000502702
R12312 VSS.n5131 VSS.n5130 0.000502702
R12313 VSS.n5696 VSS.n5695 0.000502702
R12314 VSS.n2458 VSS.n2457 0.000502702
R12315 VSS.n2466 VSS.n2465 0.000502702
R12316 VSS.n2489 VSS.n2488 0.000502702
R12317 VSS.n2599 VSS.n2598 0.000502702
R12318 VSS.n2580 VSS.n2579 0.000502702
R12319 VSS.n2560 VSS.n2559 0.000502702
R12320 VSS.n2586 VSS.n2585 0.000502702
R12321 VSS.n2543 VSS.n2542 0.000502702
R12322 VSS.n2614 VSS.n2613 0.000502702
R12323 VSS.n5620 VSS.n2509 0.000502702
R12324 VSS.n5613 VSS.n5612 0.000502702
R12325 VSS.n462 VSS.n461 0.000502702
R12326 VSS.n561 VSS.n560 0.000502702
R12327 VSS.n7497 VSS.n7496 0.000502702
R12328 VSS.n658 VSS.n657 0.000502702
R12329 VSS.n7044 VSS.n7043 0.000502702
R12330 VSS.n7050 VSS.n7049 0.000502702
R12331 VSS.n7071 VSS.n7070 0.000502702
R12332 VSS.n7064 VSS.n7063 0.000502702
R12333 VSS.n7078 VSS.n7077 0.000502702
R12334 VSS.n7455 VSS.n7454 0.000502702
R12335 VSS.n766 VSS.n765 0.000502702
R12336 VSS.n651 VSS.n650 0.000502702
R12337 VSS.n2729 VSS.n2728 0.000502702
R12338 VSS.n371 VSS.n370 0.000502702
R12339 VSS.n7417 VSS.n7416 0.000502702
R12340 VSS.n7359 VSS.n7358 0.000502702
R12341 VSS.n7355 VSS.n7354 0.000502702
R12342 VSS.n7366 VSS.n7365 0.000502702
R12343 VSS.n7617 VSS.n7616 0.000502702
R12344 VSS.n684 VSS.n683 0.000502702
R12345 VSS.n7122 VSS.n7121 0.000502702
R12346 VSS.n7109 VSS.n7108 0.000502702
R12347 VSS.n7128 VSS.n7127 0.000502702
R12348 VSS.n7162 VSS.n7161 0.000502702
R12349 VSS.n7138 VSS.n7137 0.000502702
R12350 VSS.n7149 VSS.n7148 0.000502702
R12351 VSS.n7245 VSS.n7244 0.000502702
R12352 VSS.n7145 VSS.n7144 0.000502702
R12353 VSS.n7251 VSS.n7250 0.000502702
R12354 VSS.n6919 VSS.n6918 0.000502702
R12355 VSS.n7098 VSS.n7097 0.000502702
R12356 VSS.n7026 VSS.n7025 0.000502702
R12357 VSS.n845 VSS.n844 0.000502702
R12358 VSS.n888 VSS.n887 0.000502702
R12359 VSS.n900 VSS.n899 0.000502702
R12360 VSS.n893 VSS.n892 0.000502702
R12361 VSS.n906 VSS.n905 0.000502702
R12362 VSS.n7000 VSS.n6999 0.000502702
R12363 VSS.n911 VSS.n910 0.000502702
R12364 VSS.n6869 VSS.n6868 0.000502702
R12365 VSS.n6883 VSS.n6882 0.000502702
R12366 VSS.n6873 VSS.n6872 0.000502702
R12367 VSS.n6889 VSS.n6888 0.000502702
R12368 VSS.n6963 VSS.n6962 0.000502702
R12369 VSS.n828 VSS.n827 0.000502702
R12370 VSS.n1086 VSS.n1085 0.000502702
R12371 VSS.n1077 VSS.n1076 0.000502702
R12372 VSS.n6557 VSS.n6556 0.000502702
R12373 VSS.n1120 VSS.n1119 0.000502702
R12374 VSS.n1111 VSS.n1110 0.000502702
R12375 VSS.n6490 VSS.n6489 0.000502702
R12376 VSS.n6478 VSS.n6477 0.000502702
R12377 VSS.n6486 VSS.n6485 0.000502702
R12378 VSS.n6404 VSS.n6403 0.000502702
R12379 VSS.n1171 VSS.n1170 0.000502702
R12380 VSS.n1162 VSS.n1161 0.000502702
R12381 VSS.n1280 VSS.n1279 0.000502702
R12382 VSS.n1268 VSS.n1267 0.000502702
R12383 VSS.n1276 VSS.n1275 0.000502702
R12384 VSS.n6852 VSS.n6851 0.000502702
R12385 VSS.n6692 VSS.n6691 0.000502702
R12386 VSS.n6171 VSS.n6170 0.000502702
R12387 VSS.n6162 VSS.n6161 0.000502702
R12388 VSS.n7736 VSS.n7735 0.000502702
R12389 VSS.n7718 VSS.n7717 0.000502702
R12390 VSS.n6952 VSS.n6951 0.000502702
R12391 VSS.n7704 VSS.n7703 0.000502702
R12392 VSS.n7686 VSS.n7685 0.000502702
R12393 VSS.n6908 VSS.n6907 0.000502702
R12394 VSS.n7672 VSS.n7671 0.000502702
R12395 VSS.n7654 VSS.n7653 0.000502702
R12396 VSS.n82 VSS.n81 0.000502702
R12397 VSS.n7640 VSS.n7639 0.000502702
R12398 VSS.n175 VSS.n174 0.000502702
R12399 VSS.n183 VSS.n182 0.000502702
R12400 VSS.n149 VSS.n148 0.000502702
R12401 VSS.n144 VSS.n143 0.000502702
R12402 VSS.n7648 VSS.n7647 0.000502702
R12403 VSS.n7680 VSS.n7679 0.000502702
R12404 VSS.n7712 VSS.n7711 0.000502702
R12405 VSS.n2484 VSS.n2483 0.000502702
R12406 VSS.n5704 VSS.n5703 0.000502702
R12407 VSS.n5736 VSS.n5735 0.000502702
R12408 VSS.n5768 VSS.n5767 0.000502702
R12409 VSS.n4777 VSS.n4776 0.000502702
R12410 VSS.n4485 VSS.n4484 0.000502702
R12411 VSS.n4406 VSS.n4405 0.000502702
R12412 VSS.n4990 VSS.n4989 0.000502702
R12413 VSS.n4586 VSS.n4585 0.000502702
R12414 VSS.n4606 VSS.n4605 0.000502702
R12415 VSS.n4301 VSS.n4300 0.000502702
R12416 VSS.n4289 VSS.n4288 0.000502702
R12417 VSS.n4269 VSS.n4268 0.000502702
R12418 VSS.n4894 VSS.n4893 0.000502702
R12419 VSS.n5124 VSS.n5123 0.000502702
R12420 VSS.n4810 VSS.n4809 0.000502702
R12421 VSS.n5186 VSS.n5185 0.000502702
R12422 VSS.n4669 VSS.n4668 0.000502702
R12423 VSS.n3950 VSS.n3949 0.000502702
R12424 VSS.n2832 VSS.n2831 0.000502702
R12425 VSS.n3791 VSS.n3790 0.000502702
R12426 VSS.n5802 VSS.n5801 0.000502702
R12427 VSS.n2627 VSS.n2626 0.000502702
R12428 VSS.n2569 VSS.n2568 0.000502702
R12429 VSS.n2607 VSS.n2606 0.000502702
R12430 VSS.n389 VSS.n388 0.000502702
R12431 VSS.n7491 VSS.n7490 0.000502702
R12432 VSS.n501 VSS.n500 0.000502702
R12433 VSS.n609 VSS.n608 0.000502702
R12434 VSS.n529 VSS.n432 0.000502702
R12435 VSS.n664 VSS.n663 0.000502702
R12436 VSS.n6682 VSS.n6681 0.000502702
R12437 VSS.n7093 VSS.n7092 0.000502702
R12438 VSS.n7335 VSS.n7334 0.000502702
R12439 VSS.n7609 VSS.n7608 0.000502702
R12440 VSS.n422 VSS.n421 0.000502702
R12441 VSS.n6901 VSS.n6900 0.000502702
R12442 VSS.n6945 VSS.n6944 0.000502702
R12443 VSS.n6158 VSS.n6157 0.000502702
R12444 VSS.n944 VSS.n943 0.000502702
R12445 VSS.n1073 VSS.n1072 0.000502702
R12446 VSS.n7746 VSS.n7745 0.000502702
R12447 VSS.n7293 VSS.n7292 0.000502702
R12448 VSS.n7588 VSS.n7587 0.000502702
R12449 VSS.n7578 VSS.n7577 0.000502702
R12450 VSS.n106 VSS.n105 0.000502702
R12451 VSS.n191 VSS.n190 0.000502702
R12452 VSS.n200 VSS.n199 0.000502702
R12453 VSS.n5005 VSS.n5004 0.000502702
R12454 VSS.n4787 VSS.n4786 0.000502702
R12455 VSS.n4455 VSS.n4454 0.000502702
R12456 VSS.n4410 VSS.n4409 0.000502702
R12457 VSS.n4546 VSS.n4545 0.000502702
R12458 VSS.n4984 VSS.n4983 0.000502702
R12459 VSS.n4576 VSS.n4575 0.000502702
R12460 VSS.n4500 VSS.n4499 0.000502702
R12461 VSS.n4611 VSS.n4610 0.000502702
R12462 VSS.n5275 VSS.n5274 0.000502702
R12463 VSS.n5268 VSS.n3897 0.000502702
R12464 VSS.n4350 VSS.n4349 0.000502702
R12465 VSS.n4343 VSS.n4293 0.000502702
R12466 VSS.n4339 VSS.n4338 0.000502702
R12467 VSS.n4658 VSS.n4657 0.000502702
R12468 VSS.n4622 VSS.n4364 0.000502702
R12469 VSS.n4374 VSS.n4373 0.000502702
R12470 VSS.n4823 VSS.n4822 0.000502702
R12471 VSS.n4965 VSS.n4964 0.000502702
R12472 VSS.n4478 VSS.n4477 0.000502702
R12473 VSS.n4870 VSS.n4869 0.000502702
R12474 VSS.n5104 VSS.n5103 0.000502702
R12475 VSS.n5094 VSS.n5093 0.000502702
R12476 VSS.n4149 VSS.n4148 0.000502702
R12477 VSS.n5675 VSS.n5674 0.000502702
R12478 VSS.n5665 VSS.n5664 0.000502702
R12479 VSS.n4884 VSS.n4883 0.000502702
R12480 VSS.n4767 VSS.n4766 0.000502702
R12481 VSS.n4840 VSS.n4839 0.000502702
R12482 VSS.n4922 VSS.n4921 0.000502702
R12483 VSS.n4918 VSS.n4917 0.000502702
R12484 VSS.n5155 VSS.n5154 0.000502702
R12485 VSS.n5148 VSS.n5147 0.000502702
R12486 VSS.n5135 VSS.n5134 0.000502702
R12487 VSS.n4836 VSS.n4835 0.000502702
R12488 VSS.n4816 VSS.n4815 0.000502702
R12489 VSS.n4688 VSS.n4232 0.000502702
R12490 VSS.n4739 VSS.n4738 0.000502702
R12491 VSS.n4725 VSS.n4724 0.000502702
R12492 VSS.n5210 VSS.n5209 0.000502702
R12493 VSS.n5197 VSS.n5196 0.000502702
R12494 VSS.n4252 VSS.n4251 0.000502702
R12495 VSS.n4662 VSS.n4257 0.000502702
R12496 VSS.n4045 VSS.n4044 0.000502702
R12497 VSS.n4058 VSS.n4057 0.000502702
R12498 VSS.n4083 VSS.n3984 0.000502702
R12499 VSS.n3979 VSS.n3978 0.000502702
R12500 VSS.n3974 VSS.n3973 0.000502702
R12501 VSS.n3961 VSS.n3960 0.000502702
R12502 VSS.n5257 VSS.n5256 0.000502702
R12503 VSS.n3899 VSS.n3898 0.000502702
R12504 VSS.n4032 VSS.n4031 0.000502702
R12505 VSS.n3702 VSS.n3701 0.000502702
R12506 VSS.n3604 VSS.n3603 0.000502702
R12507 VSS.n3507 VSS.n3506 0.000502702
R12508 VSS.n3410 VSS.n3409 0.000502702
R12509 VSS.n5348 VSS.n5347 0.000502702
R12510 VSS.n2826 VSS.n2825 0.000502702
R12511 VSS.n5442 VSS.n5441 0.000502702
R12512 VSS.n3799 VSS.n3798 0.000502702
R12513 VSS.n2535 VSS.n2534 0.000502702
R12514 VSS.n468 VSS.n467 0.000502702
R12515 VSS.n399 VSS.n398 0.000502702
R12516 VSS.n2736 VSS.n2735 0.000502702
R12517 VSS.n7461 VSS.n7460 0.000502702
R12518 VSS.n647 VSS.n646 0.000502702
R12519 VSS.n599 VSS.n598 0.000502702
R12520 VSS.n7505 VSS.n7504 0.000502702
R12521 VSS.n634 VSS.n633 0.000502702
R12522 VSS.n676 VSS.n430 0.000502702
R12523 VSS.n669 VSS.n668 0.000502702
R12524 VSS.n6667 VSS.n6666 0.000502702
R12525 VSS.n824 VSS.n823 0.000502702
R12526 VSS.n780 VSS.n779 0.000502702
R12527 VSS.n757 VSS.n756 0.000502702
R12528 VSS.n7197 VSS.n7196 0.000502702
R12529 VSS.n7190 VSS.n7086 0.000502702
R12530 VSS.n640 VSS.n639 0.000502702
R12531 VSS.n7485 VSS.n7484 0.000502702
R12532 VSS.n509 VSS.n508 0.000502702
R12533 VSS.n566 VSS.n565 0.000502702
R12534 VSS.n7325 VSS.n7324 0.000502702
R12535 VSS.n379 VSS.n378 0.000502702
R12536 VSS.n694 VSS.n693 0.000502702
R12537 VSS.n7410 VSS.n7409 0.000502702
R12538 VSS.n7261 VSS.n7260 0.000502702
R12539 VSS.n7372 VSS.n7254 0.000502702
R12540 VSS.n7378 VSS.n7377 0.000502702
R12541 VSS.n85 VSS.n84 0.000502702
R12542 VSS.n690 VSS.n689 0.000502702
R12543 VSS.n435 VSS.n434 0.000502702
R12544 VSS.n7170 VSS.n7169 0.000502702
R12545 VSS.n7156 VSS.n7155 0.000502702
R12546 VSS.n6894 VSS.n6893 0.000502702
R12547 VSS.n6925 VSS.n6924 0.000502702
R12548 VSS.n6912 VSS.n6911 0.000502702
R12549 VSS.n7179 VSS.n7178 0.000502702
R12550 VSS.n7088 VSS.n7087 0.000502702
R12551 VSS.n7115 VSS.n7114 0.000502702
R12552 VSS.n7019 VSS.n7018 0.000502702
R12553 VSS.n881 VSS.n880 0.000502702
R12554 VSS.n6993 VSS.n6992 0.000502702
R12555 VSS.n6876 VSS.n6875 0.000502702
R12556 VSS.n6969 VSS.n6968 0.000502702
R12557 VSS.n6956 VSS.n6955 0.000502702
R12558 VSS.n841 VSS.n840 0.000502702
R12559 VSS.n835 VSS.n834 0.000502702
R12560 VSS.n817 VSS.n816 0.000502702
R12561 VSS.n6567 VSS.n6566 0.000502702
R12562 VSS.n6500 VSS.n6499 0.000502702
R12563 VSS.n6414 VSS.n6413 0.000502702
R12564 VSS.n1290 VSS.n1289 0.000502702
R12565 VSS.n6843 VSS.n6842 0.000502702
R12566 VSS.n954 VSS.n953 0.000502702
R12567 VSS.n6151 VSS.n6150 0.000502702
R12568 VSS.n1066 VSS.n1065 0.000502702
R12569 VSS.n6700 VSS.n6699 0.000502311
R12570 VSS.n3865 VSS.n3864 0.000502311
R12571 VSS.n3767 VSS.n3766 0.000502311
R12572 VSS.n3669 VSS.n3668 0.000502311
R12573 VSS.n2494 VSS.n2493 0.000502311
R12574 VSS.n7276 VSS.n7275 0.000502311
R12575 VSS.n253 VSS.n252 0.000502311
R12576 VSS.n7566 VSS.n7565 0.000502311
R12577 VSS.n7314 VSS.n7313 0.000502311
R12578 VSS.n157 VSS.n156 0.000502311
R12579 VSS.n4430 VSS.n4429 0.000502311
R12580 VSS.n4505 VSS.n4504 0.000502311
R12581 VSS.n4553 VSS.n4552 0.000502311
R12582 VSS.n5010 VSS.n5009 0.000502311
R12583 VSS.n4754 VSS.n4753 0.000502311
R12584 VSS.n4157 VSS.n4156 0.000502311
R12585 VSS.n2473 VSS.n2472 0.000502311
R12586 VSS.n5084 VSS.n5083 0.000502311
R12587 VSS.n4873 VSS.n4872 0.000502311
R12588 VSS.n3571 VSS.n3570 0.000502311
R12589 VSS.n3474 VSS.n3473 0.000502311
R12590 VSS.n3377 VSS.n3376 0.000502311
R12591 VSS.n5356 VSS.n5355 0.000502311
R12592 VSS.n5420 VSS.n5419 0.000502311
R12593 VSS.n6339 VSS.n6338 0.000502311
R12594 VSS.n2717 VSS.n2716 0.000502311
R12595 VSS.n2745 VSS.n2744 0.000502311
R12596 VSS.n550 VSS.n549 0.000502311
R12597 VSS.n452 VSS.n451 0.000502311
R12598 VSS.n587 VSS.n586 0.000502311
R12599 VSS.n7527 VSS.n7526 0.000502311
R12600 VSS.n7541 VSS.n7540 0.000502311
R12601 VSS.n489 VSS.n488 0.000502311
R12602 VSS.n263 VSS.n262 0.000502311
R12603 VSS.n215 VSS.n214 0.000502311
R12604 VSS.n227 VSS.n226 0.000502311
R12605 VSS.n6635 VSS.n6634 0.000502311
R12606 VSS.n6550 VSS.n6549 0.000502311
R12607 VSS.n6469 VSS.n6468 0.000502311
R12608 VSS.n6395 VSS.n6394 0.000502311
R12609 VSS.n1299 VSS.n1298 0.000502311
R12610 VSS.n6833 VSS.n6832 0.000502311
R12611 VSS.n6180 VSS.n6179 0.000502311
R12612 VSS.n5593 VSS.n5592 0.000501541
R12613 VSS.n6455 VSS.n6454 0.000501541
R12614 VSS.n6449 VSS.n6448 0.000501541
R12615 VSS.n1153 VSS.n1152 0.000501541
R12616 VSS.n6438 VSS.n6437 0.000501541
R12617 VSS.n6384 VSS.n6383 0.000501541
R12618 VSS.n6378 VSS.n6377 0.000501541
R12619 VSS.n1240 VSS.n1239 0.000501541
R12620 VSS.n1249 VSS.n1248 0.000501541
R12621 VSS.n1310 VSS.n1309 0.000501541
R12622 VSS.n1304 VSS.n1303 0.000501541
R12623 VSS.n993 VSS.n992 0.000501541
R12624 VSS.n987 VSS.n986 0.000501541
R12625 VSS.n6814 VSS.n6813 0.000501541
R12626 VSS.n6808 VSS.n6807 0.000501541
R12627 VSS.n6109 VSS.n6108 0.000501541
R12628 VSS.n6119 VSS.n6118 0.000501541
R12629 VSS.n6086 VSS.n6085 0.000501541
R12630 VSS.n6080 VSS.n6079 0.000501541
R12631 VSS.n6069 VSS.n6068 0.000501541
R12632 VSS.n6063 VSS.n6062 0.000501541
R12633 VSS.n6540 VSS.n6539 0.000501541
R12634 VSS.n6532 VSS.n6531 0.000501541
R12635 VSS.n6522 VSS.n6521 0.000501541
R12636 VSS.n6514 VSS.n6513 0.000501541
R12637 VSS.n1034 VSS.n1033 0.000501541
R12638 VSS.n6617 VSS.n6616 0.000501541
R12639 VSS.n6610 VSS.n6609 0.000501541
R12640 VSS.n6587 VSS.n6586 0.000501541
R12641 VSS.n6581 VSS.n6580 0.000501541
R12642 VSS.n1044 VSS.n1043 0.000501541
R12643 VSS.n1054 VSS.n1053 0.000501541
R12644 VSS.n3832 VSS.n3831 0.000501541
R12645 VSS.n3826 VSS.n3825 0.000501541
R12646 VSS.n3848 VSS.n3847 0.000501541
R12647 VSS.n3842 VSS.n3841 0.000501541
R12648 VSS.n3751 VSS.n3750 0.000501541
R12649 VSS.n3745 VSS.n3744 0.000501541
R12650 VSS.n3735 VSS.n3734 0.000501541
R12651 VSS.n3729 VSS.n3728 0.000501541
R12652 VSS.n3653 VSS.n3652 0.000501541
R12653 VSS.n3647 VSS.n3646 0.000501541
R12654 VSS.n3637 VSS.n3636 0.000501541
R12655 VSS.n3631 VSS.n3630 0.000501541
R12656 VSS.n3556 VSS.n3555 0.000501541
R12657 VSS.n3550 VSS.n3549 0.000501541
R12658 VSS.n3540 VSS.n3539 0.000501541
R12659 VSS.n3534 VSS.n3533 0.000501541
R12660 VSS.n3459 VSS.n3458 0.000501541
R12661 VSS.n3453 VSS.n3452 0.000501541
R12662 VSS.n3443 VSS.n3442 0.000501541
R12663 VSS.n3437 VSS.n3436 0.000501541
R12664 VSS.n3362 VSS.n3361 0.000501541
R12665 VSS.n3356 VSS.n3355 0.000501541
R12666 VSS.n3346 VSS.n3345 0.000501541
R12667 VSS.n3340 VSS.n3339 0.000501541
R12668 VSS.n5370 VSS.n5369 0.000501541
R12669 VSS.n5374 VSS.n5373 0.000501541
R12670 VSS.n5483 VSS.n5482 0.000501541
R12671 VSS.n5477 VSS.n5476 0.000501541
R12672 VSS.n5405 VSS.n5404 0.000501541
R12673 VSS.n5399 VSS.n5398 0.000501541
R12674 VSS.n5834 VSS.n5833 0.000501541
R12675 VSS.n5828 VSS.n5827 0.000501541
R12676 VSS.n5583 VSS.n5582 0.000501541
R12677 VSS.n5572 VSS.n5571 0.000501541
R12678 VSS.n5578 VSS.n5577 0.000501541
R12679 VSS.n5566 VSS.n5565 0.000501541
R12680 VSS.n2771 VSS.n2769 0.000501541
R12681 VSS.n998 VSS.n996 0.000501541
R12682 VSS.n6592 VSS.n6590 0.000501541
R12683 VSS.n6621 VSS.n6620 0.000501541
R12684 VSS.n1050 VSS.n1048 0.000501541
R12685 VSS.n6709 VSS.n6708 0.000501541
R12686 VSS.n6711 VSS.n6705 0.000501541
R12687 VSS.n3852 VSS.n3851 0.000501541
R12688 VSS.n3836 VSS.n3835 0.000501541
R12689 VSS.n3447 VSS.n3446 0.000501541
R12690 VSS.n5393 VSS.n2103 0.000501541
R12691 VSS.n5409 VSS.n5408 0.000501541
R12692 VSS.n5381 VSS.n5379 0.000501541
R12693 VSS.n5365 VSS.n5363 0.000501541
R12694 VSS.n3350 VSS.n3349 0.000501541
R12695 VSS.n3366 VSS.n3365 0.000501541
R12696 VSS.n3463 VSS.n3462 0.000501541
R12697 VSS.n3544 VSS.n3543 0.000501541
R12698 VSS.n3560 VSS.n3559 0.000501541
R12699 VSS.n3641 VSS.n3640 0.000501541
R12700 VSS.n3657 VSS.n3656 0.000501541
R12701 VSS.n3739 VSS.n3738 0.000501541
R12702 VSS.n3755 VSS.n3754 0.000501541
R12703 VSS.n6526 VSS.n6525 0.000501541
R12704 VSS.n6544 VSS.n6543 0.000501541
R12705 VSS.n6074 VSS.n6072 0.000501541
R12706 VSS.n6193 VSS.n6191 0.000501541
R12707 VSS.n6115 VSS.n6113 0.000501541
R12708 VSS.n6820 VSS.n6819 0.000501541
R12709 VSS.n1316 VSS.n1315 0.000501541
R12710 VSS.n1245 VSS.n1243 0.000501541
R12711 VSS.n6389 VSS.n6388 0.000501541
R12712 VSS.n6443 VSS.n6442 0.000501541
R12713 VSS.n6459 VSS.n6458 0.000501541
R12714 VSS.n6099 VSS.n6098 0.000500621
R12715 VSS.n6096 VSS.n6095 0.000500621
R12716 VSS.n6093 VSS.n6092 0.000500621
R12717 VSS.n1461 VSS.n1457 0.000500621
R12718 VSS.n1463 VSS.n1457 0.000500621
R12719 VSS.n1464 VSS.n1463 0.000500621
R12720 VSS.n1589 VSS.n1584 0.000500621
R12721 VSS.n1589 VSS.n1588 0.000500621
R12722 VSS.n1584 VSS.n1583 0.000500621
R12723 VSS.n2707 VSS.n2706 0.000500621
R12724 VSS.n2704 VSS.n2703 0.000500621
R12725 VSS.n2634 VSS.n2633 0.000500621
R12726 VSS.n2640 VSS.n2634 0.000500621
R12727 VSS.n2640 VSS.n2639 0.000500621
R12728 VSS.n2637 VSS.n2636 0.000500621
R12729 VSS.n2646 VSS.n2644 0.000500621
R12730 VSS.n2651 VSS.n2644 0.000500621
R12731 VSS.n2651 VSS.n2650 0.000500621
R12732 VSS.n2648 VSS.n2647 0.000500621
R12733 VSS.n2658 VSS.n2657 0.000500621
R12734 VSS.n2671 VSS.n2670 0.000500621
R12735 VSS.n2667 VSS.n2666 0.000500621
R12736 VSS.n2673 VSS.n2667 0.000500621
R12737 VSS.n2673 VSS.n2672 0.000500621
R12738 VSS.n2685 VSS.n2684 0.000500621
R12739 VSS.n2681 VSS.n2680 0.000500621
R12740 VSS.n2687 VSS.n2681 0.000500621
R12741 VSS.n2687 VSS.n2686 0.000500621
R12742 VSS.n2694 VSS.n2693 0.000500621
R12743 VSS.n2698 VSS.n2697 0.000500621
R12744 VSS.n572 VSS.n571 0.000500621
R12745 VSS.n578 VSS.n577 0.000500621
R12746 VSS.n575 VSS.n574 0.000500621
R12747 VSS.n472 VSS.n471 0.000500621
R12748 VSS.n478 VSS.n477 0.000500621
R12749 VSS.n475 VSS.n474 0.000500621
R12750 VSS.n7297 VSS.n7296 0.000500621
R12751 VSS.n7303 VSS.n7302 0.000500621
R12752 VSS.n7300 VSS.n7299 0.000500621
R12753 VSS.n278 VSS.n277 0.000500621
R12754 VSS.n275 VSS.n274 0.000500621
R12755 VSS.n281 VSS.n280 0.000500621
R12756 VSS.n1709 VSS.n1704 0.000500621
R12757 VSS.n1709 VSS.n1708 0.000500621
R12758 VSS.n123 VSS.n109 0.000500621
R12759 VSS.n7555 VSS.n7554 0.000500621
R12760 VSS.n111 VSS.n110 0.000500621
R12761 VSS.n236 VSS.n235 0.000500621
R12762 VSS.n233 VSS.n232 0.000500621
R12763 VSS.n239 VSS.n238 0.000500621
R12764 VSS.n161 VSS.n127 0.000500621
R12765 VSS.n1653 VSS.n1651 0.000500621
R12766 VSS.n1658 VSS.n1651 0.000500621
R12767 VSS.n1658 VSS.n1657 0.000500621
R12768 VSS.n1727 VSS.n1725 0.000500621
R12769 VSS.n1725 VSS.n1661 0.000500621
R12770 VSS.n1661 VSS.n1660 0.000500621
R12771 VSS.n1655 VSS.n1654 0.000500621
R12772 VSS.n1536 VSS.n1534 0.000500621
R12773 VSS.n1541 VSS.n1534 0.000500621
R12774 VSS.n1541 VSS.n1540 0.000500621
R12775 VSS.n1538 VSS.n1537 0.000500621
R12776 VSS.n1608 VSS.n1604 0.000500621
R12777 VSS.n1608 VSS.n1607 0.000500621
R12778 VSS.n1604 VSS.n1603 0.000500621
R12779 VSS.n1770 VSS.n1767 0.000500621
R12780 VSS.n1767 VSS.n1581 0.000500621
R12781 VSS.n1770 VSS.n1769 0.000500621
R12782 VSS.n1474 VSS.n1469 0.000500621
R12783 VSS.n1474 VSS.n1473 0.000500621
R12784 VSS.n1469 VSS.n1468 0.000500621
R12785 VSS.n1400 VSS.n1399 0.000500621
R12786 VSS.n1406 VSS.n1399 0.000500621
R12787 VSS.n1406 VSS.n1405 0.000500621
R12788 VSS.n1499 VSS.n1498 0.000500621
R12789 VSS.n1497 VSS.n1496 0.000500621
R12790 VSS.n1503 VSS.n1496 0.000500621
R12791 VSS.n1503 VSS.n1502 0.000500621
R12792 VSS.n1841 VSS.n1840 0.000500621
R12793 VSS.n1530 VSS.n1529 0.000500621
R12794 VSS.n1761 VSS.n1756 0.000500621
R12795 VSS.n1761 VSS.n1760 0.000500621
R12796 VSS.n1756 VSS.n1755 0.000500621
R12797 VSS.n1751 VSS.n1746 0.000500621
R12798 VSS.n1751 VSS.n1750 0.000500621
R12799 VSS.n1746 VSS.n1745 0.000500621
R12800 VSS.n1713 VSS.n1712 0.000500621
R12801 VSS.n1719 VSS.n1713 0.000500621
R12802 VSS.n1719 VSS.n1718 0.000500621
R12803 VSS.n1689 VSS.n1684 0.000500621
R12804 VSS.n1689 VSS.n1688 0.000500621
R12805 VSS.n1684 VSS.n1683 0.000500621
R12806 VSS.n1693 VSS.n1692 0.000500621
R12807 VSS.n1699 VSS.n1693 0.000500621
R12808 VSS.n1699 VSS.n1698 0.000500621
R12809 VSS.n1740 VSS.n1734 0.000500621
R12810 VSS.n1740 VSS.n1739 0.000500621
R12811 VSS.n1823 VSS.n1821 0.000500621
R12812 VSS.n1821 VSS.n1820 0.000500621
R12813 VSS.n1824 VSS.n1823 0.000500621
R12814 VSS.n1834 VSS.n1829 0.000500621
R12815 VSS.n1834 VSS.n1833 0.000500621
R12816 VSS.n1424 VSS.n1419 0.000500621
R12817 VSS.n1424 VSS.n1423 0.000500621
R12818 VSS.n1419 VSS.n1418 0.000500621
R12819 VSS.n1433 VSS.n1431 0.000500621
R12820 VSS.n1431 VSS.n1430 0.000500621
R12821 VSS.n1434 VSS.n1433 0.000500621
R12822 VSS.n1814 VSS.n1809 0.000500621
R12823 VSS.n1814 VSS.n1813 0.000500621
R12824 VSS.n1809 VSS.n1808 0.000500621
R12825 VSS.n1804 VSS.n1803 0.000500621
R12826 VSS.n1803 VSS.n1802 0.000500621
R12827 VSS.n1802 VSS.n1801 0.000500621
R12828 VSS.n1448 VSS.n1447 0.000500621
R12829 VSS.n1454 VSS.n1448 0.000500621
R12830 VSS.n1454 VSS.n1453 0.000500621
R12831 VSS.n1438 VSS.n1437 0.000500621
R12832 VSS.n1444 VSS.n1438 0.000500621
R12833 VSS.n1444 VSS.n1443 0.000500621
R12834 VSS.n1783 VSS.n1777 0.000500621
R12835 VSS.n1783 VSS.n1782 0.000500621
R12836 VSS.n1793 VSS.n1791 0.000500621
R12837 VSS.n1791 VSS.n1790 0.000500621
R12838 VSS.n1794 VSS.n1793 0.000500621
R12839 VSS.n1599 VSS.n1594 0.000500621
R12840 VSS.n1599 VSS.n1598 0.000500621
R12841 VSS.n1594 VSS.n1593 0.000500621
R12842 VSS.n1668 VSS.n1666 0.000500621
R12843 VSS.n1669 VSS.n1662 0.000500621
R12844 VSS.n1669 VSS.n1668 0.000500621
R12845 VSS.n1679 VSS.n1674 0.000500621
R12846 VSS.n1679 VSS.n1678 0.000500621
R12847 VSS.n1674 VSS.n1673 0.000500621
R12848 VSS.n7516 VSS.n7515 0.000500621
R12849 VSS.n7513 VSS.n7512 0.000500621
R12850 VSS.n7510 VSS.n7509 0.000500621
R12851 VSS.n7547 VSS.n7546 0.000500621
R12852 VSS.n291 VSS.n290 0.000500621
R12853 VSS.n1620 VSS.n1615 0.000500621
R12854 VSS.n1614 VSS.n1613 0.000500621
R12855 VSS.n1620 VSS.n1614 0.000500621
R12856 VSS.n1619 VSS.n1618 0.000500621
R12857 VSS.n1555 VSS.n1550 0.000500621
R12858 VSS.n1549 VSS.n1548 0.000500621
R12859 VSS.n1555 VSS.n1549 0.000500621
R12860 VSS.n1554 VSS.n1553 0.000500621
R12861 VSS.n1486 VSS.n1481 0.000500621
R12862 VSS.n1480 VSS.n1479 0.000500621
R12863 VSS.n1486 VSS.n1480 0.000500621
R12864 VSS.n1485 VSS.n1484 0.000500621
R12865 VSS.n1379 VSS.n1374 0.000500621
R12866 VSS.n1373 VSS.n1372 0.000500621
R12867 VSS.n1379 VSS.n1373 0.000500621
R12868 VSS.n1378 VSS.n1377 0.000500621
R12869 VSS.n6354 VSS.n6353 0.000500621
R12870 VSS.n1858 VSS.n1857 0.000500621
R12871 VSS.n1861 VSS.n1860 0.000500621
R12872 VSS.n1855 VSS.n1854 0.000500621
R12873 VSS.n1354 VSS.n1353 0.000500621
R12874 VSS.n1351 VSS.n1350 0.000500621
R12875 VSS.n1357 VSS.n1356 0.000500621
R12876 VSS.n1339 VSS.n1338 0.000500621
R12877 VSS.n1334 VSS.n1333 0.000500621
R12878 VSS.n1336 VSS.n1335 0.000500621
R12879 VSS.n6363 VSS.n6362 0.000500621
R12880 VSS.n1177 VSS.n1176 0.000500621
R12881 VSS.n1327 VSS.n1326 0.000500621
R12882 VSS.n1214 VSS.n1213 0.000500621
R12883 VSS.n1209 VSS.n1208 0.000500621
R12884 VSS.n1211 VSS.n1210 0.000500621
R12885 VSS.n1201 VSS.n1200 0.000500621
R12886 VSS.n1198 VSS.n1197 0.000500621
R12887 VSS.n1204 VSS.n1203 0.000500621
R12888 VSS.n1416 VSS.n1415 0.000500621
R12889 VSS.n1849 VSS.n1416 0.000500621
R12890 VSS.n1850 VSS.n1849 0.000500621
R12891 VSS.n1402 VSS.n1401 0.000500621
R12892 VSS.n1459 VSS.n1458 0.00050031
R12893 VSS.n1586 VSS.n1585 0.00050031
R12894 VSS.n1667 VSS.n1611 0.00050031
R12895 VSS.n573 VSS.n112 0.00050031
R12896 VSS.n473 VSS.n284 0.00050031
R12897 VSS.n273 VSS.n116 0.00050031
R12898 VSS.n7298 VSS.n120 0.00050031
R12899 VSS.n1706 VSS.n1705 0.00050031
R12900 VSS.n7552 VSS.n7551 0.00050031
R12901 VSS.n231 VSS.n122 0.00050031
R12902 VSS.n1730 VSS.n1729 0.00050031
R12903 VSS.n1726 VSS.n1629 0.00050031
R12904 VSS.n1754 VSS.n1532 0.00050031
R12905 VSS.n1592 VSS.n1546 0.00050031
R12906 VSS.n1606 VSS.n1605 0.00050031
R12907 VSS.n1773 VSS.n1772 0.00050031
R12908 VSS.n1768 VSS.n1564 0.00050031
R12909 VSS.n1602 VSS.n1568 0.00050031
R12910 VSS.n1781 VSS.n1477 0.00050031
R12911 VSS.n1467 VSS.n1362 0.00050031
R12912 VSS.n1471 VSS.n1470 0.00050031
R12913 VSS.n1843 VSS.n1842 0.00050031
R12914 VSS.n1527 VSS.n1526 0.00050031
R12915 VSS.n1759 VSS.n1758 0.00050031
R12916 VSS.n1748 VSS.n1747 0.00050031
R12917 VSS.n1716 VSS.n1715 0.00050031
R12918 VSS.n1686 VSS.n1685 0.00050031
R12919 VSS.n1682 VSS.n1645 0.00050031
R12920 VSS.n1717 VSS.n1641 0.00050031
R12921 VSS.n1696 VSS.n1695 0.00050031
R12922 VSS.n1697 VSS.n1630 0.00050031
R12923 VSS.n1703 VSS.n1632 0.00050031
R12924 VSS.n1736 VSS.n1735 0.00050031
R12925 VSS.n1738 VSS.n1578 0.00050031
R12926 VSS.n1744 VSS.n1574 0.00050031
R12927 VSS.n1818 VSS.n1817 0.00050031
R12928 VSS.n1831 VSS.n1830 0.00050031
R12929 VSS.n1828 VSS.n1524 0.00050031
R12930 VSS.n1822 VSS.n1512 0.00050031
R12931 VSS.n1417 VSS.n1394 0.00050031
R12932 VSS.n1421 VSS.n1420 0.00050031
R12933 VSS.n1432 VSS.n1366 0.00050031
R12934 VSS.n1428 VSS.n1427 0.00050031
R12935 VSS.n1812 VSS.n1811 0.00050031
R12936 VSS.n1798 VSS.n1797 0.00050031
R12937 VSS.n1800 VSS.n1516 0.00050031
R12938 VSS.n1807 VSS.n1520 0.00050031
R12939 VSS.n1452 VSS.n1390 0.00050031
R12940 VSS.n1450 VSS.n1449 0.00050031
R12941 VSS.n1442 VSS.n1370 0.00050031
R12942 VSS.n1440 VSS.n1439 0.00050031
R12943 VSS.n1780 VSS.n1779 0.00050031
R12944 VSS.n1788 VSS.n1787 0.00050031
R12945 VSS.n1597 VSS.n1596 0.00050031
R12946 VSS.n1665 VSS.n1664 0.00050031
R12947 VSS.n1676 VSS.n1675 0.00050031
R12948 VSS.n7511 VSS.n293 0.00050031
R12949 VSS.n1672 VSS.n1624 0.00050031
R12950 VSS.n1582 VSS.n1559 0.00050031
R12951 VSS.n1792 VSS.n1490 0.00050031
R12952 VSS.n1460 VSS.n1385 0.00050031
R12953 VSS.n1414 VSS.n1413 0.00050031
R12954 VSS.n1852 VSS.n1851 0.00050031
R12955 VSS.n4461 VSS.n4460 0.000500172
R12956 VSS.n4459 VSS.n4458 0.000500172
R12957 VSS.n5279 VSS.n5278 0.000500172
R12958 VSS.n3886 VSS.n3885 0.000500172
R12959 VSS.n4322 VSS.n4321 0.000500172
R12960 VSS.n4315 VSS.n4314 0.000500172
R12961 VSS.n4327 VSS.n4326 0.000500172
R12962 VSS.n4331 VSS.n4326 0.000500172
R12963 VSS.n4333 VSS.n4294 0.000500172
R12964 VSS.n4333 VSS.n4332 0.000500172
R12965 VSS.n4304 VSS.n4294 0.000500172
R12966 VSS.n4332 VSS.n4304 0.000500172
R12967 VSS.n4633 VSS.n4632 0.000500172
R12968 VSS.n4354 VSS.n4353 0.000500172
R12969 VSS.n4644 VSS.n4277 0.000500172
R12970 VSS.n4644 VSS.n4643 0.000500172
R12971 VSS.n4277 VSS.n4275 0.000500172
R12972 VSS.n4643 VSS.n4275 0.000500172
R12973 VSS.n4638 VSS.n4637 0.000500172
R12974 VSS.n4642 VSS.n4637 0.000500172
R12975 VSS.n4950 VSS.n4949 0.000500172
R12976 VSS.n4949 VSS.n4948 0.000500172
R12977 VSS.n4952 VSS.n4205 0.000500172
R12978 VSS.n4952 VSS.n4951 0.000500172
R12979 VSS.n4207 VSS.n4205 0.000500172
R12980 VSS.n4951 VSS.n4207 0.000500172
R12981 VSS.n4976 VSS.n4974 0.000500172
R12982 VSS.n4976 VSS.n4975 0.000500172
R12983 VSS.n4973 VSS.n4968 0.000500172
R12984 VSS.n4597 VSS.n4595 0.000500172
R12985 VSS.n4597 VSS.n4596 0.000500172
R12986 VSS.n4594 VSS.n4590 0.000500172
R12987 VSS.n4468 VSS.n4466 0.000500172
R12988 VSS.n4468 VSS.n4467 0.000500172
R12989 VSS.n4465 VSS.n4413 0.000500172
R12990 VSS.n4434 VSS.n4416 0.000500172
R12991 VSS.n4433 VSS.n4432 0.000500172
R12992 VSS.n4418 VSS.n4417 0.000500172
R12993 VSS.n4514 VSS.n4513 0.000500172
R12994 VSS.n4508 VSS.n4507 0.000500172
R12995 VSS.n4503 VSS.n4502 0.000500172
R12996 VSS.n4570 VSS.n4569 0.000500172
R12997 VSS.n4550 VSS.n4549 0.000500172
R12998 VSS.n4533 VSS.n4532 0.000500172
R12999 VSS.n5019 VSS.n5018 0.000500172
R13000 VSS.n5013 VSS.n5012 0.000500172
R13001 VSS.n5008 VSS.n5007 0.000500172
R13002 VSS.n5041 VSS.n5040 0.000500172
R13003 VSS.n4771 VSS.n4770 0.000500172
R13004 VSS.n4752 VSS.n4751 0.000500172
R13005 VSS.n4856 VSS.n4855 0.000500172
R13006 VSS.n2453 VSS.n2452 0.000500172
R13007 VSS.n2470 VSS.n2469 0.000500172
R13008 VSS.n5659 VSS.n5658 0.000500172
R13009 VSS.n5086 VSS.n5085 0.000500172
R13010 VSS.n5088 VSS.n5087 0.000500172
R13011 VSS.n4875 VSS.n4874 0.000500172
R13012 VSS.n4877 VSS.n4876 0.000500172
R13013 VSS.n5117 VSS.n5116 0.000500172
R13014 VSS.n5116 VSS.n5115 0.000500172
R13015 VSS.n5119 VSS.n5118 0.000500172
R13016 VSS.n4905 VSS.n4903 0.000500172
R13017 VSS.n4905 VSS.n4904 0.000500172
R13018 VSS.n4902 VSS.n4898 0.000500172
R13019 VSS.n4798 VSS.n4796 0.000500172
R13020 VSS.n4798 VSS.n4797 0.000500172
R13021 VSS.n4795 VSS.n4791 0.000500172
R13022 VSS.n5179 VSS.n5178 0.000500172
R13023 VSS.n5178 VSS.n5177 0.000500172
R13024 VSS.n5180 VSS.n4107 0.000500172
R13025 VSS.n4108 VSS.n4107 0.000500172
R13026 VSS.n5181 VSS.n4108 0.000500172
R13027 VSS.n5181 VSS.n5180 0.000500172
R13028 VSS.n5171 VSS.n5168 0.000500172
R13029 VSS.n5171 VSS.n5170 0.000500172
R13030 VSS.n5167 VSS.n4114 0.000500172
R13031 VSS.n4114 VSS.n4113 0.000500172
R13032 VSS.n5167 VSS.n5166 0.000500172
R13033 VSS.n5166 VSS.n4113 0.000500172
R13034 VSS.n4222 VSS.n4216 0.000500172
R13035 VSS.n4222 VSS.n4221 0.000500172
R13036 VSS.n4224 VSS.n4217 0.000500172
R13037 VSS.n4935 VSS.n4224 0.000500172
R13038 VSS.n4217 VSS.n4215 0.000500172
R13039 VSS.n4935 VSS.n4215 0.000500172
R13040 VSS.n4938 VSS.n4214 0.000500172
R13041 VSS.n4939 VSS.n4214 0.000500172
R13042 VSS.n4944 VSS.n4943 0.000500172
R13043 VSS.n4943 VSS.n4212 0.000500172
R13044 VSS.n4945 VSS.n4212 0.000500172
R13045 VSS.n4945 VSS.n4944 0.000500172
R13046 VSS.n5221 VSS.n5220 0.000500172
R13047 VSS.n5220 VSS.n5219 0.000500172
R13048 VSS.n3934 VSS.n3933 0.000500172
R13049 VSS.n3935 VSS.n3933 0.000500172
R13050 VSS.n5215 VSS.n3935 0.000500172
R13051 VSS.n5215 VSS.n3934 0.000500172
R13052 VSS.n3932 VSS.n3929 0.000500172
R13053 VSS.n5224 VSS.n3932 0.000500172
R13054 VSS.n3930 VSS.n3928 0.000500172
R13055 VSS.n5229 VSS.n3928 0.000500172
R13056 VSS.n5229 VSS.n5228 0.000500172
R13057 VSS.n5228 VSS.n3930 0.000500172
R13058 VSS.n3927 VSS.n3924 0.000500172
R13059 VSS.n5232 VSS.n3927 0.000500172
R13060 VSS.n3925 VSS.n3923 0.000500172
R13061 VSS.n5237 VSS.n3923 0.000500172
R13062 VSS.n5237 VSS.n5236 0.000500172
R13063 VSS.n5236 VSS.n3925 0.000500172
R13064 VSS.n5242 VSS.n3919 0.000500172
R13065 VSS.n5242 VSS.n5241 0.000500172
R13066 VSS.n5244 VSS.n3920 0.000500172
R13067 VSS.n5245 VSS.n5244 0.000500172
R13068 VSS.n3920 VSS.n3918 0.000500172
R13069 VSS.n5245 VSS.n3918 0.000500172
R13070 VSS.n5250 VSS.n5249 0.000500172
R13071 VSS.n5249 VSS.n5248 0.000500172
R13072 VSS.n5252 VSS.n3913 0.000500172
R13073 VSS.n5252 VSS.n5251 0.000500172
R13074 VSS.n3913 VSS.n3912 0.000500172
R13075 VSS.n5251 VSS.n3912 0.000500172
R13076 VSS.n5331 VSS.n5330 0.000500172
R13077 VSS.n5330 VSS.n5329 0.000500172
R13078 VSS.n5332 VSS.n2835 0.000500172
R13079 VSS.n2836 VSS.n2835 0.000500172
R13080 VSS.n5333 VSS.n2836 0.000500172
R13081 VSS.n5333 VSS.n5332 0.000500172
R13082 VSS.n2843 VSS.n2838 0.000500172
R13083 VSS.n2839 VSS.n2838 0.000500172
R13084 VSS.n5321 VSS.n2842 0.000500172
R13085 VSS.n5321 VSS.n5320 0.000500172
R13086 VSS.n5319 VSS.n2842 0.000500172
R13087 VSS.n5320 VSS.n5319 0.000500172
R13088 VSS.n5316 VSS.n2845 0.000500172
R13089 VSS.n5316 VSS.n5315 0.000500172
R13090 VSS.n5312 VSS.n2847 0.000500172
R13091 VSS.n5312 VSS.n5311 0.000500172
R13092 VSS.n5310 VSS.n2847 0.000500172
R13093 VSS.n5311 VSS.n5310 0.000500172
R13094 VSS.n5307 VSS.n2849 0.000500172
R13095 VSS.n5307 VSS.n5306 0.000500172
R13096 VSS.n5303 VSS.n2851 0.000500172
R13097 VSS.n5303 VSS.n5302 0.000500172
R13098 VSS.n5301 VSS.n2851 0.000500172
R13099 VSS.n5302 VSS.n5301 0.000500172
R13100 VSS.n5298 VSS.n2853 0.000500172
R13101 VSS.n5298 VSS.n5297 0.000500172
R13102 VSS.n5294 VSS.n2855 0.000500172
R13103 VSS.n5294 VSS.n5293 0.000500172
R13104 VSS.n5292 VSS.n2855 0.000500172
R13105 VSS.n5293 VSS.n5292 0.000500172
R13106 VSS.n5289 VSS.n2857 0.000500172
R13107 VSS.n5289 VSS.n5288 0.000500172
R13108 VSS.n5285 VSS.n2859 0.000500172
R13109 VSS.n5285 VSS.n5284 0.000500172
R13110 VSS.n5283 VSS.n2859 0.000500172
R13111 VSS.n5284 VSS.n5283 0.000500172
R13112 VSS.n3866 VSS.n2865 0.000500172
R13113 VSS.n3868 VSS.n3867 0.000500172
R13114 VSS.n3816 VSS.n3815 0.000500172
R13115 VSS.n3805 VSS.n3804 0.000500172
R13116 VSS.n3803 VSS.n3771 0.000500172
R13117 VSS.n3803 VSS.n3802 0.000500172
R13118 VSS.n3768 VSS.n2874 0.000500172
R13119 VSS.n3770 VSS.n3769 0.000500172
R13120 VSS.n3719 VSS.n3718 0.000500172
R13121 VSS.n3708 VSS.n3707 0.000500172
R13122 VSS.n3706 VSS.n3673 0.000500172
R13123 VSS.n3706 VSS.n3705 0.000500172
R13124 VSS.n3670 VSS.n2883 0.000500172
R13125 VSS.n3672 VSS.n3671 0.000500172
R13126 VSS.n3610 VSS.n3609 0.000500172
R13127 VSS.n3608 VSS.n3575 0.000500172
R13128 VSS.n3608 VSS.n3607 0.000500172
R13129 VSS.n3574 VSS.n3573 0.000500172
R13130 VSS.n2893 VSS.n2892 0.000500172
R13131 VSS.n3513 VSS.n3512 0.000500172
R13132 VSS.n3511 VSS.n3478 0.000500172
R13133 VSS.n3511 VSS.n3510 0.000500172
R13134 VSS.n3477 VSS.n3476 0.000500172
R13135 VSS.n2904 VSS.n2903 0.000500172
R13136 VSS.n3416 VSS.n3415 0.000500172
R13137 VSS.n3414 VSS.n3381 0.000500172
R13138 VSS.n3414 VSS.n3413 0.000500172
R13139 VSS.n3380 VSS.n3379 0.000500172
R13140 VSS.n2916 VSS.n2915 0.000500172
R13141 VSS.n3319 VSS.n2817 0.000500172
R13142 VSS.n5353 VSS.n5352 0.000500172
R13143 VSS.n5352 VSS.n5351 0.000500172
R13144 VSS.n5354 VSS.n2815 0.000500172
R13145 VSS.n2814 VSS.n2813 0.000500172
R13146 VSS.n5456 VSS.n5455 0.000500172
R13147 VSS.n5819 VSS.n5818 0.000500172
R13148 VSS.n5389 VSS.n5388 0.000500172
R13149 VSS.n5422 VSS.n5421 0.000500172
R13150 VSS.n5454 VSS.n5423 0.000500172
R13151 VSS.n5454 VSS.n5453 0.000500172
R13152 VSS.n2376 VSS.n2375 0.000500172
R13153 VSS.n5787 VSS.n2375 0.000500172
R13154 VSS.n5787 VSS.n5786 0.000500172
R13155 VSS.n5788 VSS.n5787 0.000500172
R13156 VSS.n5784 VSS.n5781 0.000500172
R13157 VSS.n5784 VSS.n5783 0.000500172
R13158 VSS.n2381 VSS.n2380 0.000500172
R13159 VSS.n5780 VSS.n2381 0.000500172
R13160 VSS.n5780 VSS.n5779 0.000500172
R13161 VSS.n5779 VSS.n2380 0.000500172
R13162 VSS.n2395 VSS.n2394 0.000500172
R13163 VSS.n5755 VSS.n2394 0.000500172
R13164 VSS.n5755 VSS.n5754 0.000500172
R13165 VSS.n5756 VSS.n5755 0.000500172
R13166 VSS.n5752 VSS.n5749 0.000500172
R13167 VSS.n5752 VSS.n5751 0.000500172
R13168 VSS.n2400 VSS.n2399 0.000500172
R13169 VSS.n5748 VSS.n2400 0.000500172
R13170 VSS.n5748 VSS.n5747 0.000500172
R13171 VSS.n5747 VSS.n2399 0.000500172
R13172 VSS.n2414 VSS.n2413 0.000500172
R13173 VSS.n5723 VSS.n2413 0.000500172
R13174 VSS.n5723 VSS.n5722 0.000500172
R13175 VSS.n5724 VSS.n5723 0.000500172
R13176 VSS.n5720 VSS.n5717 0.000500172
R13177 VSS.n5720 VSS.n5719 0.000500172
R13178 VSS.n2419 VSS.n2418 0.000500172
R13179 VSS.n5716 VSS.n2419 0.000500172
R13180 VSS.n5716 VSS.n5715 0.000500172
R13181 VSS.n5715 VSS.n2418 0.000500172
R13182 VSS.n5689 VSS.n5687 0.000500172
R13183 VSS.n5691 VSS.n5687 0.000500172
R13184 VSS.n5691 VSS.n5690 0.000500172
R13185 VSS.n5692 VSS.n5691 0.000500172
R13186 VSS.n5685 VSS.n5683 0.000500172
R13187 VSS.n5685 VSS.n5684 0.000500172
R13188 VSS.n5682 VSS.n5681 0.000500172
R13189 VSS.n5626 VSS.n5625 0.000500172
R13190 VSS.n2507 VSS.n2506 0.000500172
R13191 VSS.n5624 VSS.n2508 0.000500172
R13192 VSS.n2518 VSS.n2517 0.000500172
R13193 VSS.n2623 VSS.n2622 0.000500172
R13194 VSS.n2622 VSS.n2621 0.000500172
R13195 VSS.n2622 VSS.n2518 0.000500172
R13196 VSS.n2595 VSS.n2594 0.000500172
R13197 VSS.n2556 VSS.n2555 0.000500172
R13198 VSS.n2574 VSS.n2564 0.000500172
R13199 VSS.n2573 VSS.n2572 0.000500172
R13200 VSS.n2545 VSS.n2540 0.000500172
R13201 VSS.n2591 VSS.n2590 0.000500172
R13202 VSS.n2590 VSS.n2540 0.000500172
R13203 VSS.n2590 VSS.n2589 0.000500172
R13204 VSS.n2618 VSS.n2617 0.000500172
R13205 VSS.n2610 VSS.n2522 0.000500172
R13206 VSS.n5608 VSS.n5607 0.000500172
R13207 VSS.n2742 VSS.n2741 0.000500172
R13208 VSS.n2722 VSS.n2721 0.000500172
R13209 VSS.n2740 VSS.n2739 0.000500172
R13210 VSS.n6671 VSS.n6670 0.000500172
R13211 VSS.n6678 VSS.n6677 0.000500172
R13212 VSS.n7059 VSS.n7058 0.000500172
R13213 VSS.n7054 VSS.n7053 0.000500172
R13214 VSS.n7206 VSS.n745 0.000500172
R13215 VSS.n7206 VSS.n7205 0.000500172
R13216 VSS.n7203 VSS.n749 0.000500172
R13217 VSS.n749 VSS.n748 0.000500172
R13218 VSS.n7202 VSS.n748 0.000500172
R13219 VSS.n7203 VSS.n7202 0.000500172
R13220 VSS.n770 VSS.n769 0.000500172
R13221 VSS.n775 VSS.n774 0.000500172
R13222 VSS.n7447 VSS.n322 0.000500172
R13223 VSS.n322 VSS.n320 0.000500172
R13224 VSS.n7448 VSS.n320 0.000500172
R13225 VSS.n7448 VSS.n7447 0.000500172
R13226 VSS.n326 VSS.n325 0.000500172
R13227 VSS.n7446 VSS.n325 0.000500172
R13228 VSS.n7438 VSS.n328 0.000500172
R13229 VSS.n7438 VSS.n7437 0.000500172
R13230 VSS.n7440 VSS.n329 0.000500172
R13231 VSS.n7441 VSS.n7440 0.000500172
R13232 VSS.n329 VSS.n327 0.000500172
R13233 VSS.n7441 VSS.n327 0.000500172
R13234 VSS.n7468 VSS.n7467 0.000500172
R13235 VSS.n7466 VSS.n7464 0.000500172
R13236 VSS.n7472 VSS.n307 0.000500172
R13237 VSS.n7477 VSS.n7473 0.000500172
R13238 VSS.n7477 VSS.n7476 0.000500172
R13239 VSS.n624 VSS.n614 0.000500172
R13240 VSS.n620 VSS.n618 0.000500172
R13241 VSS.n620 VSS.n619 0.000500172
R13242 VSS.n520 VSS.n518 0.000500172
R13243 VSS.n520 VSS.n519 0.000500172
R13244 VSS.n517 VSS.n513 0.000500172
R13245 VSS.n589 VSS.n588 0.000500172
R13246 VSS.n591 VSS.n590 0.000500172
R13247 VSS.n7529 VSS.n7528 0.000500172
R13248 VSS.n7531 VSS.n7530 0.000500172
R13249 VSS.n491 VSS.n490 0.000500172
R13250 VSS.n493 VSS.n492 0.000500172
R13251 VSS.n366 VSS.n365 0.000500172
R13252 VSS.n261 VSS.n260 0.000500172
R13253 VSS.n383 VSS.n382 0.000500172
R13254 VSS.n225 VSS.n170 0.000500172
R13255 VSS.n224 VSS.n223 0.000500172
R13256 VSS.n7568 VSS.n7567 0.000500172
R13257 VSS.n7570 VSS.n7569 0.000500172
R13258 VSS.n7316 VSS.n7315 0.000500172
R13259 VSS.n7318 VSS.n7317 0.000500172
R13260 VSS.n7598 VSS.n7597 0.000500172
R13261 VSS.n7599 VSS.n7598 0.000500172
R13262 VSS.n7595 VSS.n7594 0.000500172
R13263 VSS.n7596 VSS.n7595 0.000500172
R13264 VSS.n7344 VSS.n7343 0.000500172
R13265 VSS.n7349 VSS.n7338 0.000500172
R13266 VSS.n7349 VSS.n7348 0.000500172
R13267 VSS.n7348 VSS.n7347 0.000500172
R13268 VSS.n410 VSS.n408 0.000500172
R13269 VSS.n410 VSS.n409 0.000500172
R13270 VSS.n414 VSS.n404 0.000500172
R13271 VSS.n7389 VSS.n7388 0.000500172
R13272 VSS.n7388 VSS.n7387 0.000500172
R13273 VSS.n709 VSS.n708 0.000500172
R13274 VSS.n710 VSS.n708 0.000500172
R13275 VSS.n7383 VSS.n710 0.000500172
R13276 VSS.n7383 VSS.n709 0.000500172
R13277 VSS.n7400 VSS.n707 0.000500172
R13278 VSS.n7392 VSS.n707 0.000500172
R13279 VSS.n706 VSS.n705 0.000500172
R13280 VSS.n705 VSS.n703 0.000500172
R13281 VSS.n7404 VSS.n706 0.000500172
R13282 VSS.n7404 VSS.n703 0.000500172
R13283 VSS.n7393 VSS.n336 0.000500172
R13284 VSS.n7394 VSS.n7393 0.000500172
R13285 VSS.n338 VSS.n337 0.000500172
R13286 VSS.n7423 VSS.n338 0.000500172
R13287 VSS.n337 VSS.n335 0.000500172
R13288 VSS.n7423 VSS.n335 0.000500172
R13289 VSS.n7426 VSS.n334 0.000500172
R13290 VSS.n7427 VSS.n334 0.000500172
R13291 VSS.n7432 VSS.n7431 0.000500172
R13292 VSS.n7431 VSS.n332 0.000500172
R13293 VSS.n7433 VSS.n332 0.000500172
R13294 VSS.n7433 VSS.n7432 0.000500172
R13295 VSS.n6938 VSS.n6937 0.000500172
R13296 VSS.n6937 VSS.n6936 0.000500172
R13297 VSS.n6939 VSS.n6929 0.000500172
R13298 VSS.n6930 VSS.n6929 0.000500172
R13299 VSS.n6940 VSS.n6930 0.000500172
R13300 VSS.n6940 VSS.n6939 0.000500172
R13301 VSS.n7234 VSS.n727 0.000500172
R13302 VSS.n729 VSS.n727 0.000500172
R13303 VSS.n725 VSS.n723 0.000500172
R13304 VSS.n726 VSS.n725 0.000500172
R13305 VSS.n7238 VSS.n726 0.000500172
R13306 VSS.n7238 VSS.n723 0.000500172
R13307 VSS.n735 VSS.n730 0.000500172
R13308 VSS.n731 VSS.n730 0.000500172
R13309 VSS.n7229 VSS.n734 0.000500172
R13310 VSS.n7229 VSS.n7228 0.000500172
R13311 VSS.n7227 VSS.n734 0.000500172
R13312 VSS.n7228 VSS.n7227 0.000500172
R13313 VSS.n7224 VSS.n737 0.000500172
R13314 VSS.n7224 VSS.n7223 0.000500172
R13315 VSS.n7220 VSS.n739 0.000500172
R13316 VSS.n7220 VSS.n7219 0.000500172
R13317 VSS.n7218 VSS.n739 0.000500172
R13318 VSS.n7219 VSS.n7218 0.000500172
R13319 VSS.n7215 VSS.n741 0.000500172
R13320 VSS.n7215 VSS.n7214 0.000500172
R13321 VSS.n7211 VSS.n743 0.000500172
R13322 VSS.n7211 VSS.n7210 0.000500172
R13323 VSS.n7209 VSS.n743 0.000500172
R13324 VSS.n7210 VSS.n7209 0.000500172
R13325 VSS.n6980 VSS.n6979 0.000500172
R13326 VSS.n6979 VSS.n6978 0.000500172
R13327 VSS.n6974 VSS.n934 0.000500172
R13328 VSS.n6974 VSS.n935 0.000500172
R13329 VSS.n934 VSS.n933 0.000500172
R13330 VSS.n935 VSS.n933 0.000500172
R13331 VSS.n6985 VSS.n6984 0.000500172
R13332 VSS.n6984 VSS.n6983 0.000500172
R13333 VSS.n6987 VSS.n920 0.000500172
R13334 VSS.n6987 VSS.n6986 0.000500172
R13335 VSS.n922 VSS.n920 0.000500172
R13336 VSS.n6986 VSS.n922 0.000500172
R13337 VSS.n928 VSS.n868 0.000500172
R13338 VSS.n928 VSS.n927 0.000500172
R13339 VSS.n870 VSS.n869 0.000500172
R13340 VSS.n7006 VSS.n870 0.000500172
R13341 VSS.n869 VSS.n867 0.000500172
R13342 VSS.n7006 VSS.n867 0.000500172
R13343 VSS.n7011 VSS.n7010 0.000500172
R13344 VSS.n7010 VSS.n7009 0.000500172
R13345 VSS.n7013 VSS.n854 0.000500172
R13346 VSS.n7013 VSS.n7012 0.000500172
R13347 VSS.n856 VSS.n854 0.000500172
R13348 VSS.n7012 VSS.n856 0.000500172
R13349 VSS.n862 VSS.n803 0.000500172
R13350 VSS.n862 VSS.n861 0.000500172
R13351 VSS.n805 VSS.n804 0.000500172
R13352 VSS.n7032 VSS.n805 0.000500172
R13353 VSS.n804 VSS.n802 0.000500172
R13354 VSS.n7032 VSS.n802 0.000500172
R13355 VSS.n6673 VSS.n799 0.000500172
R13356 VSS.n800 VSS.n799 0.000500172
R13357 VSS.n798 VSS.n797 0.000500172
R13358 VSS.n797 VSS.n795 0.000500172
R13359 VSS.n7037 VSS.n798 0.000500172
R13360 VSS.n7037 VSS.n795 0.000500172
R13361 VSS.n6661 VSS.n6660 0.000500172
R13362 VSS.n6697 VSS.n6696 0.000500172
R13363 VSS.n6644 VSS.n6643 0.000500172
R13364 VSS.n6640 VSS.n6639 0.000500172
R13365 VSS.n6639 VSS.n6638 0.000500172
R13366 VSS.n6636 VSS.n1090 0.000500172
R13367 VSS.n1089 VSS.n1088 0.000500172
R13368 VSS.n6572 VSS.n6571 0.000500172
R13369 VSS.n6570 VSS.n6569 0.000500172
R13370 VSS.n6570 VSS.n6553 0.000500172
R13371 VSS.n6551 VSS.n1124 0.000500172
R13372 VSS.n1123 VSS.n1122 0.000500172
R13373 VSS.n6505 VSS.n6504 0.000500172
R13374 VSS.n6503 VSS.n6502 0.000500172
R13375 VSS.n6503 VSS.n6472 0.000500172
R13376 VSS.n6470 VSS.n1144 0.000500172
R13377 VSS.n1143 VSS.n1142 0.000500172
R13378 VSS.n6419 VSS.n6418 0.000500172
R13379 VSS.n6417 VSS.n6416 0.000500172
R13380 VSS.n6417 VSS.n6400 0.000500172
R13381 VSS.n6398 VSS.n6397 0.000500172
R13382 VSS.n1174 VSS.n1173 0.000500172
R13383 VSS.n1260 VSS.n1259 0.000500172
R13384 VSS.n1293 VSS.n1292 0.000500172
R13385 VSS.n1293 VSS.n1262 0.000500172
R13386 VSS.n1296 VSS.n1295 0.000500172
R13387 VSS.n1233 VSS.n1232 0.000500172
R13388 VSS.n978 VSS.n940 0.000500172
R13389 VSS.n6840 VSS.n6839 0.000500172
R13390 VSS.n6839 VSS.n6838 0.000500172
R13391 VSS.n6836 VSS.n6835 0.000500172
R13392 VSS.n957 VSS.n956 0.000500172
R13393 VSS.n6142 VSS.n6141 0.000500172
R13394 VSS.n7751 VSS.n7750 0.000500172
R13395 VSS.n6103 VSS.n6102 0.000500172
R13396 VSS.n6177 VSS.n6176 0.000500172
R13397 VSS.n6174 VSS.n6143 0.000500172
R13398 VSS.n6174 VSS.n6173 0.000500172
R13399 VSS.n19 VSS.n18 0.000500172
R13400 VSS.n7731 VSS.n18 0.000500172
R13401 VSS.n7731 VSS.n7730 0.000500172
R13402 VSS.n7732 VSS.n7731 0.000500172
R13403 VSS.n7728 VSS.n7725 0.000500172
R13404 VSS.n7728 VSS.n7727 0.000500172
R13405 VSS.n24 VSS.n23 0.000500172
R13406 VSS.n7724 VSS.n24 0.000500172
R13407 VSS.n7724 VSS.n7723 0.000500172
R13408 VSS.n7723 VSS.n23 0.000500172
R13409 VSS.n38 VSS.n37 0.000500172
R13410 VSS.n7699 VSS.n37 0.000500172
R13411 VSS.n7699 VSS.n7698 0.000500172
R13412 VSS.n7700 VSS.n7699 0.000500172
R13413 VSS.n7696 VSS.n7693 0.000500172
R13414 VSS.n7696 VSS.n7695 0.000500172
R13415 VSS.n43 VSS.n42 0.000500172
R13416 VSS.n7692 VSS.n43 0.000500172
R13417 VSS.n7692 VSS.n7691 0.000500172
R13418 VSS.n7691 VSS.n42 0.000500172
R13419 VSS.n57 VSS.n56 0.000500172
R13420 VSS.n7667 VSS.n56 0.000500172
R13421 VSS.n7667 VSS.n7666 0.000500172
R13422 VSS.n7668 VSS.n7667 0.000500172
R13423 VSS.n7664 VSS.n7661 0.000500172
R13424 VSS.n7664 VSS.n7663 0.000500172
R13425 VSS.n62 VSS.n61 0.000500172
R13426 VSS.n7660 VSS.n62 0.000500172
R13427 VSS.n7660 VSS.n7659 0.000500172
R13428 VSS.n7659 VSS.n61 0.000500172
R13429 VSS.n7633 VSS.n7631 0.000500172
R13430 VSS.n7635 VSS.n7631 0.000500172
R13431 VSS.n7635 VSS.n7634 0.000500172
R13432 VSS.n7636 VSS.n7635 0.000500172
R13433 VSS.n7629 VSS.n7627 0.000500172
R13434 VSS.n7629 VSS.n7628 0.000500172
R13435 VSS.n7624 VSS.n7623 0.000500172
R13436 VSS.n7623 VSS.n77 0.000500172
R13437 VSS.n153 VSS.n152 0.000500172
R13438 VSS.n4462 VSS.n4461 0.000500086
R13439 VSS.n4459 VSS.n4452 0.000500086
R13440 VSS.n5280 VSS.n5279 0.000500086
R13441 VSS.n3886 VSS.n2860 0.000500086
R13442 VSS.n4323 VSS.n4322 0.000500086
R13443 VSS.n4315 VSS.n4306 0.000500086
R13444 VSS.n4634 VSS.n4633 0.000500086
R13445 VSS.n4354 VSS.n4278 0.000500086
R13446 VSS.n2555 VSS.n2539 0.000500086
R13447 VSS.n2594 VSS.n2593 0.000500086
R13448 VSS.n2610 VSS.n2519 0.000500086
R13449 VSS.n2619 VSS.n2618 0.000500086
R13450 VSS.n6672 VSS.n6671 0.000500086
R13451 VSS.n6677 VSS.n6676 0.000500086
R13452 VSS.n7058 VSS.n7057 0.000500086
R13453 VSS.n7055 VSS.n7054 0.000500086
R13454 VSS.n771 VSS.n770 0.000500086
R13455 VSS.n774 VSS.n773 0.000500086
R13456 VSS.n7469 VSS.n7468 0.000500086
R13457 VSS.n7466 VSS.n7465 0.000500086
R13458 VDD.n330 VDD 646.457
R13459 VDD.n99 VDD.n98 469.212
R13460 VDD.n23 VDD 459.156
R13461 VDD.n244 VDD 454.192
R13462 VDD.n314 VDD.n310 304.469
R13463 VDD.n265 VDD.n264 301.644
R13464 VDD.n282 VDD.n281 301.644
R13465 VDD.n290 VDD.n289 301.644
R13466 VDD.n44 VDD.n43 301.644
R13467 VDD.n60 VDD.n59 301.644
R13468 VDD.n68 VDD.n67 301.644
R13469 VDD.n249 VDD.n248 292.5
R13470 VDD.n257 VDD.n256 292.5
R13471 VDD.n237 VDD.n236 292.5
R13472 VDD.n229 VDD.n228 292.5
R13473 VDD.n303 VDD.n302 292.5
R13474 VDD.n86 VDD.n85 292.5
R13475 VDD.n5 VDD.n4 292.5
R13476 VDD.n8 VDD.n7 292.5
R13477 VDD.n28 VDD.n27 292.5
R13478 VDD.n36 VDD.n35 292.5
R13479 VDD.n16 VDD.n15 292.5
R13480 VDD.n328 VDD 279.115
R13481 VDD.t36 VDD.t116 274.072
R13482 VDD VDD.t34 258.938
R13483 VDD VDD.t66 258.481
R13484 VDD.t94 VDD.t114 208.496
R13485 VDD VDD.t142 200.089
R13486 VDD.t44 VDD 193.022
R13487 VDD.t54 VDD 193.022
R13488 VDD.t46 VDD 182.952
R13489 VDD.t82 VDD 182.952
R13490 VDD.t87 VDD.t2 179.595
R13491 VDD.t62 VDD 176.238
R13492 VDD.t98 VDD 176.238
R13493 VDD.t89 VDD.t12 172.881
R13494 VDD.n280 VDD.n279 170.916
R13495 VDD.n58 VDD.n57 170.916
R13496 VDD.n266 VDD.n263 166.381
R13497 VDD.n45 VDD.n42 166.381
R13498 VDD.n272 VDD.n271 164.215
R13499 VDD.n50 VDD.n19 164.215
R13500 VDD.n234 VDD.n233 160.918
R13501 VDD.n13 VDD.n12 160.918
R13502 VDD.t22 VDD.t36 159.736
R13503 VDD.t134 VDD.t120 159.736
R13504 VDD.t38 VDD.t46 159.452
R13505 VDD.t58 VDD.t56 159.452
R13506 VDD.t48 VDD.t82 159.452
R13507 VDD.t132 VDD.t78 159.452
R13508 VDD.t2 VDD.t90 159.452
R13509 VDD.n247 VDD.t25 158.06
R13510 VDD.n255 VDD.t31 158.06
R13511 VDD.n26 VDD.t51 158.06
R13512 VDD.n34 VDD.t29 158.06
R13513 VDD.n326 VDD.t9 152.879
R13514 VDD.n0 VDD.t1 151.633
R13515 VDD.n319 VDD.t143 151.633
R13516 VDD.n321 VDD.t97 149.696
R13517 VDD.n92 VDD.t113 149.696
R13518 VDD.t24 VDD.t44 149.382
R13519 VDD.t50 VDD.t54 149.382
R13520 VDD.n331 VDD.n330 147.387
R13521 VDD.t10 VDD.n243 146.025
R13522 VDD.t100 VDD.n22 146.025
R13523 VDD.n274 VDD.t75 145.868
R13524 VDD.n288 VDD.t21 145.868
R13525 VDD.n52 VDD.t107 145.868
R13526 VDD.n66 VDD.t131 145.868
R13527 VDD.t90 VDD.t89 142.668
R13528 VDD.t142 VDD.t96 141.239
R13529 VDD.t70 VDD.t74 140.989
R13530 VDD.t110 VDD.t14 140.989
R13531 VDD.t16 VDD.t20 140.989
R13532 VDD.t102 VDD.t106 140.989
R13533 VDD.t140 VDD.t124 140.989
R13534 VDD.t126 VDD.t130 140.989
R13535 VDD.n329 VDD.t8 136.196
R13536 VDD.t76 VDD 135.954
R13537 VDD.t20 VDD.t10 135.954
R13538 VDD.t108 VDD 135.954
R13539 VDD.t130 VDD.t100 135.954
R13540 VDD.t92 VDD.t87 135.954
R13541 VDD.t88 VDD.t0 132.597
R13542 VDD.t0 VDD.t84 132.597
R13543 VDD.t86 VDD.t92 129.24
R13544 VDD.t122 VDD.n242 127.562
R13545 VDD VDD.t30 120.849
R13546 VDD VDD.t28 120.849
R13547 VDD.n98 VDD.n97 120.481
R13548 VDD.t96 VDD 117.7
R13549 VDD.n328 VDD.n327 116.73
R13550 VDD.n243 VDD.n231 116.73
R13551 VDD.n22 VDD.n10 116.73
R13552 VDD.t118 VDD 112.656
R13553 VDD.t74 VDD.t58 112.457
R13554 VDD.t106 VDD.t132 112.457
R13555 VDD VDD.t64 110.778
R13556 VDD VDD.t68 110.778
R13557 VDD.n313 VDD.n312 108.525
R13558 VDD.t114 VDD.t22 107.612
R13559 VDD.t34 VDD.t115 102.567
R13560 VDD.t18 VDD.t60 102.385
R13561 VDD.t128 VDD.t4 102.385
R13562 VDD.n98 VDD.t84 102.385
R13563 VDD.t72 VDD.t80 100.707
R13564 VDD.t104 VDD.t138 100.707
R13565 VDD.t12 VDD.t85 92.315
R13566 VDD.t14 VDD.t6 83.9228
R13567 VDD.t124 VDD.t40 83.9228
R13568 VDD.t32 VDD.t136 82.2443
R13569 VDD.t26 VDD.t52 82.2443
R13570 VDD.n302 VDD.t37 77.3934
R13571 VDD.n228 VDD.t95 77.3934
R13572 VDD.n236 VDD.t57 77.3934
R13573 VDD.n256 VDD.t47 77.3934
R13574 VDD.n248 VDD.t45 77.3934
R13575 VDD.n264 VDD.t81 77.3934
R13576 VDD.n281 VDD.t61 77.3934
R13577 VDD.n289 VDD.t123 77.3934
R13578 VDD.n310 VDD.t121 77.3934
R13579 VDD.n7 VDD.t93 77.3934
R13580 VDD.n4 VDD.t91 77.3934
R13581 VDD.n85 VDD.t99 77.3934
R13582 VDD.n15 VDD.t79 77.3934
R13583 VDD.n35 VDD.t83 77.3934
R13584 VDD.n27 VDD.t55 77.3934
R13585 VDD.n43 VDD.t139 77.3934
R13586 VDD.n59 VDD.t5 77.3934
R13587 VDD.n67 VDD.t63 77.3934
R13588 VDD.n314 VDD.n313 68.8164
R13589 VDD.t85 VDD.t98 67.1383
R13590 VDD.t120 VDD.t118 63.8943
R13591 VDD.n330 VDD.n329 61.4756
R13592 VDD VDD.t112 60.4245
R13593 VDD.t136 VDD.t72 58.7461
R13594 VDD.t52 VDD.t104 58.7461
R13595 VDD.t115 VDD.t94 57.1686
R13596 VDD.n311 VDD.t117 57.1305
R13597 VDD.n311 VDD.t119 57.1305
R13598 VDD.t6 VDD.t18 57.0676
R13599 VDD.t40 VDD.t128 57.0676
R13600 VDD VDD.t32 50.3539
R13601 VDD VDD.t110 50.3539
R13602 VDD VDD.t26 50.3539
R13603 VDD VDD.t140 50.3539
R13604 VDD.n242 VDD 48.7616
R13605 VDD.n242 VDD 48.6754
R13606 VDD.t116 VDD.t134 42.0359
R13607 VDD.n329 VDD 42.0359
R13608 VDD.n302 VDD.t23 41.0422
R13609 VDD.n228 VDD.t35 41.0422
R13610 VDD.n236 VDD.t59 41.0422
R13611 VDD.n256 VDD.t39 41.0422
R13612 VDD.n248 VDD.t65 41.0422
R13613 VDD.n264 VDD.t137 41.0422
R13614 VDD.n281 VDD.t7 41.0422
R13615 VDD.n289 VDD.t11 41.0422
R13616 VDD.n310 VDD.t135 41.0422
R13617 VDD.n7 VDD.t67 41.0422
R13618 VDD.n4 VDD.t3 41.0422
R13619 VDD.n85 VDD.t13 41.0422
R13620 VDD.n15 VDD.t133 41.0422
R13621 VDD.n35 VDD.t49 41.0422
R13622 VDD.n27 VDD.t69 41.0422
R13623 VDD.n43 VDD.t53 41.0422
R13624 VDD.n59 VDD.t41 41.0422
R13625 VDD.n67 VDD.t101 41.0422
R13626 VDD.t80 VDD.t76 40.2832
R13627 VDD.t56 VDD 40.2832
R13628 VDD.t138 VDD.t108 40.2832
R13629 VDD.t78 VDD 40.2832
R13630 VDD.t60 VDD.t16 38.6047
R13631 VDD.t4 VDD.t126 38.6047
R13632 VDD.n312 VDD.t42 34.8005
R13633 VDD.n312 VDD.t43 34.8005
R13634 VDD.n267 VDD.n262 34.6358
R13635 VDD.n46 VDD.n41 34.6358
R13636 VDD.n254 VDD.n241 34.6358
R13637 VDD.n262 VDD.n240 34.6358
R13638 VDD.n287 VDD.n286 34.6358
R13639 VDD.n295 VDD.n231 34.6358
R13640 VDD.n296 VDD.n295 34.6358
R13641 VDD.n297 VDD.n296 34.6358
R13642 VDD.n301 VDD.n300 34.6358
R13643 VDD.n304 VDD.n301 34.6358
R13644 VDD.n308 VDD.n226 34.6358
R13645 VDD.n309 VDD.n308 34.6358
R13646 VDD.n315 VDD.n224 34.6358
R13647 VDD.n327 VDD.n222 34.6358
R13648 VDD.n91 VDD.n2 34.6358
R13649 VDD.n84 VDD.n83 34.6358
R13650 VDD.n87 VDD.n84 34.6358
R13651 VDD.n79 VDD.n78 34.6358
R13652 VDD.n80 VDD.n79 34.6358
R13653 VDD.n73 VDD.n10 34.6358
R13654 VDD.n74 VDD.n73 34.6358
R13655 VDD.n75 VDD.n74 34.6358
R13656 VDD.n33 VDD.n21 34.6358
R13657 VDD.n41 VDD.n20 34.6358
R13658 VDD.n65 VDD.n64 34.6358
R13659 VDD.t66 VDD.t86 30.2125
R13660 VDD.n273 VDD.n272 28.9887
R13661 VDD.n51 VDD.n50 28.9887
R13662 VDD.n142 VDD.t146 27.8779
R13663 VDD.n151 VDD.t148 27.8779
R13664 VDD.n160 VDD.t147 27.8779
R13665 VDD.n280 VDD.n278 27.4829
R13666 VDD.n58 VDD.n56 27.4829
R13667 VDD.n263 VDD.t33 26.5955
R13668 VDD.n263 VDD.t73 26.5955
R13669 VDD.n271 VDD.t77 26.5955
R13670 VDD.n271 VDD.t71 26.5955
R13671 VDD.n279 VDD.t111 26.5955
R13672 VDD.n279 VDD.t15 26.5955
R13673 VDD.n233 VDD.t19 26.5955
R13674 VDD.n233 VDD.t17 26.5955
R13675 VDD.n42 VDD.t27 26.5955
R13676 VDD.n42 VDD.t105 26.5955
R13677 VDD.n19 VDD.t109 26.5955
R13678 VDD.n19 VDD.t103 26.5955
R13679 VDD.n57 VDD.t141 26.5955
R13680 VDD.n57 VDD.t125 26.5955
R13681 VDD.n12 VDD.t129 26.5955
R13682 VDD.n12 VDD.t127 26.5955
R13683 VDD.n320 VDD.n319 25.977
R13684 VDD.n93 VDD.n0 25.977
R13685 VDD.n321 VDD.n320 24.4711
R13686 VDD.n93 VDD.n92 24.4711
R13687 VDD.n331 VDD.n221 23.7181
R13688 VDD.n246 VDD.n244 23.7181
R13689 VDD.n283 VDD.n280 23.7181
R13690 VDD.n319 VDD.n224 23.7181
R13691 VDD.n321 VDD.n222 23.7181
R13692 VDD.n92 VDD.n91 23.7181
R13693 VDD.n25 VDD.n23 23.7181
R13694 VDD.n61 VDD.n58 23.7181
R13695 VDD.n291 VDD.n290 19.9534
R13696 VDD.n69 VDD.n68 19.9534
R13697 VDD.n327 VDD.n326 18.4476
R13698 VDD.n266 VDD.n265 18.0711
R13699 VDD.n45 VDD.n44 18.0711
R13700 VDD.n283 VDD.n282 17.3181
R13701 VDD.n61 VDD.n60 17.3181
R13702 VDD.n326 VDD.n221 16.1887
R13703 VDD.n272 VDD.n239 15.4358
R13704 VDD.n50 VDD.n18 15.4358
R13705 VDD.n265 VDD.n239 14.6829
R13706 VDD.n44 VDD.n18 14.6829
R13707 VDD.n290 VDD.n231 14.6829
R13708 VDD.n68 VDD.n10 14.6829
R13709 VDD.n243 VDD.t122 13.4281
R13710 VDD.n22 VDD.t62 13.4281
R13711 VDD.n97 VDD.n0 12.8005
R13712 VDD.n250 VDD.n247 10.5417
R13713 VDD.n258 VDD.n255 10.5417
R13714 VDD.n282 VDD.n234 10.5417
R13715 VDD.n29 VDD.n26 10.5417
R13716 VDD.n37 VDD.n34 10.5417
R13717 VDD.n60 VDD.n13 10.5417
R13718 VDD.n198 VDD.n197 10.416
R13719 VDD.t64 VDD.t24 10.0712
R13720 VDD.t68 VDD.t50 10.0712
R13721 VDD.n249 VDD.n241 9.84252
R13722 VDD.n278 VDD.n237 9.84252
R13723 VDD.n300 VDD.n229 9.84252
R13724 VDD.n78 VDD.n8 9.84252
R13725 VDD.n28 VDD.n21 9.84252
R13726 VDD.n56 VDD.n16 9.84252
R13727 VDD.n274 VDD.n273 9.41227
R13728 VDD.n288 VDD.n287 9.41227
R13729 VDD.n52 VDD.n51 9.41227
R13730 VDD.n66 VDD.n65 9.41227
R13731 VDD.n87 VDD.n86 9.35848
R13732 VDD.t112 VDD.t88 8.39273
R13733 VDD.n247 VDD.n246 8.28285
R13734 VDD.n255 VDD.n254 8.28285
R13735 VDD.n26 VDD.n25 8.28285
R13736 VDD.n34 VDD.n33 8.28285
R13737 VDD.n257 VDD.n240 7.20722
R13738 VDD.n303 VDD.n226 7.20722
R13739 VDD.n83 VDD.n5 7.20722
R13740 VDD.n36 VDD.n20 7.20722
R13741 VDD.n286 VDD.n234 6.77697
R13742 VDD.n64 VDD.n13 6.77697
R13743 VDD.n258 VDD.n257 6.72319
R13744 VDD.n304 VDD.n303 6.72319
R13745 VDD.n80 VDD.n5 6.72319
R13746 VDD.n37 VDD.n36 6.72319
R13747 VDD.n314 VDD.n309 5.27109
R13748 VDD.t8 VDD.n328 5.04475
R13749 VDD VDD.t70 5.03584
R13750 VDD VDD.t102 5.03584
R13751 VDD VDD.n244 4.68175
R13752 VDD VDD.n23 4.68175
R13753 VDD.n251 VDD.n250 4.6505
R13754 VDD.n272 VDD.n270 4.6505
R13755 VDD.n276 VDD.n275 4.6505
R13756 VDD.n280 VDD.n235 4.6505
R13757 VDD.n298 VDD.n297 4.6505
R13758 VDD.n319 VDD.n318 4.6505
R13759 VDD.n322 VDD.n321 4.6505
R13760 VDD.n327 VDD.n325 4.6505
R13761 VDD.n246 VDD.n245 4.6505
R13762 VDD.n252 VDD.n241 4.6505
R13763 VDD.n254 VDD.n253 4.6505
R13764 VDD.n259 VDD.n258 4.6505
R13765 VDD.n260 VDD.n240 4.6505
R13766 VDD.n262 VDD.n261 4.6505
R13767 VDD.n268 VDD.n267 4.6505
R13768 VDD.n269 VDD.n239 4.6505
R13769 VDD.n273 VDD.n238 4.6505
R13770 VDD.n278 VDD.n277 4.6505
R13771 VDD.n284 VDD.n283 4.6505
R13772 VDD.n286 VDD.n285 4.6505
R13773 VDD.n287 VDD.n232 4.6505
R13774 VDD.n292 VDD.n291 4.6505
R13775 VDD.n293 VDD.n231 4.6505
R13776 VDD.n295 VDD.n294 4.6505
R13777 VDD.n296 VDD.n230 4.6505
R13778 VDD.n300 VDD.n299 4.6505
R13779 VDD.n301 VDD.n227 4.6505
R13780 VDD.n305 VDD.n304 4.6505
R13781 VDD.n306 VDD.n226 4.6505
R13782 VDD.n308 VDD.n307 4.6505
R13783 VDD.n309 VDD.n225 4.6505
R13784 VDD.n316 VDD.n315 4.6505
R13785 VDD.n317 VDD.n224 4.6505
R13786 VDD.n320 VDD.n223 4.6505
R13787 VDD.n323 VDD.n222 4.6505
R13788 VDD.n324 VDD.n221 4.6505
R13789 VDD.n332 VDD.n331 4.6505
R13790 VDD.n25 VDD.n24 4.6505
R13791 VDD.n30 VDD.n29 4.6505
R13792 VDD.n31 VDD.n21 4.6505
R13793 VDD.n33 VDD.n32 4.6505
R13794 VDD.n38 VDD.n37 4.6505
R13795 VDD.n39 VDD.n20 4.6505
R13796 VDD.n41 VDD.n40 4.6505
R13797 VDD.n47 VDD.n46 4.6505
R13798 VDD.n48 VDD.n18 4.6505
R13799 VDD.n50 VDD.n49 4.6505
R13800 VDD.n51 VDD.n17 4.6505
R13801 VDD.n54 VDD.n53 4.6505
R13802 VDD.n56 VDD.n55 4.6505
R13803 VDD.n58 VDD.n14 4.6505
R13804 VDD.n62 VDD.n61 4.6505
R13805 VDD.n64 VDD.n63 4.6505
R13806 VDD.n65 VDD.n11 4.6505
R13807 VDD.n70 VDD.n69 4.6505
R13808 VDD.n71 VDD.n10 4.6505
R13809 VDD.n73 VDD.n72 4.6505
R13810 VDD.n74 VDD.n9 4.6505
R13811 VDD.n76 VDD.n75 4.6505
R13812 VDD.n78 VDD.n77 4.6505
R13813 VDD.n79 VDD.n6 4.6505
R13814 VDD.n81 VDD.n80 4.6505
R13815 VDD.n83 VDD.n82 4.6505
R13816 VDD.n84 VDD.n3 4.6505
R13817 VDD.n88 VDD.n87 4.6505
R13818 VDD.n89 VDD.n2 4.6505
R13819 VDD.n91 VDD.n90 4.6505
R13820 VDD.n92 VDD.n1 4.6505
R13821 VDD.n94 VDD.n93 4.6505
R13822 VDD.n95 VDD.n0 4.6505
R13823 VDD.n97 VDD.n96 4.6505
R13824 VDD.n86 VDD.n2 4.57193
R13825 VDD.n342 VDD 4.39723
R13826 VDD.n250 VDD.n249 4.0879
R13827 VDD.n275 VDD.n237 4.0879
R13828 VDD.n297 VDD.n229 4.0879
R13829 VDD.n75 VDD.n8 4.0879
R13830 VDD.n29 VDD.n28 4.0879
R13831 VDD.n53 VDD.n16 4.0879
R13832 VDD.n115 VDD 4.05613
R13833 VDD.n137 VDD 2.29217
R13834 VDD.n162 VDD 2.29217
R13835 VDD.n267 VDD.n266 1.88285
R13836 VDD.n46 VDD.n45 1.88285
R13837 VDD.t30 VDD.t38 1.67895
R13838 VDD.t28 VDD.t48 1.67895
R13839 VDD.n140 VDD.n138 1.57342
R13840 VDD.n141 VDD.n140 1.57342
R13841 VDD.n149 VDD.n147 1.57342
R13842 VDD.n150 VDD.n149 1.57342
R13843 VDD.n158 VDD.n156 1.57342
R13844 VDD.n159 VDD.n158 1.57342
R13845 VDD VDD.n354 1.4367
R13846 VDD.n333 VDD 1.34425
R13847 VDD.n139 VDD 0.828181
R13848 VDD.n148 VDD 0.828181
R13849 VDD.n157 VDD 0.828181
R13850 VDD.n139 VDD 0.827501
R13851 VDD.n148 VDD 0.827501
R13852 VDD.n157 VDD 0.827501
R13853 VDD.n194 VDD.n191 0.579775
R13854 VDD.n275 VDD.n274 0.376971
R13855 VDD.n291 VDD.n288 0.376971
R13856 VDD.n315 VDD.n314 0.376971
R13857 VDD.n53 VDD.n52 0.376971
R13858 VDD.n69 VDD.n66 0.376971
R13859 VDD VDD.n143 0.3755
R13860 VDD VDD.n152 0.3755
R13861 VDD.n184 VDD.n183 0.355402
R13862 VDD.n313 VDD.n311 0.322282
R13863 VDD.n134 VDD 0.234474
R13864 VDD.n140 VDD.n139 0.232147
R13865 VDD.n149 VDD.n148 0.232147
R13866 VDD.n158 VDD.n157 0.232147
R13867 VDD.n99 VDD 0.207531
R13868 VDD.n99 VDD 0.129576
R13869 VDD.n252 VDD.n251 0.120292
R13870 VDD.n260 VDD.n259 0.120292
R13871 VDD.n269 VDD.n268 0.120292
R13872 VDD.n270 VDD.n269 0.120292
R13873 VDD.n276 VDD.n238 0.120292
R13874 VDD.n284 VDD.n235 0.120292
R13875 VDD.n285 VDD.n284 0.120292
R13876 VDD.n285 VDD.n232 0.120292
R13877 VDD.n292 VDD.n232 0.120292
R13878 VDD.n298 VDD.n230 0.120292
R13879 VDD.n299 VDD.n298 0.120292
R13880 VDD.n299 VDD.n227 0.120292
R13881 VDD.n305 VDD.n227 0.120292
R13882 VDD.n306 VDD.n305 0.120292
R13883 VDD.n307 VDD.n306 0.120292
R13884 VDD.n307 VDD.n225 0.120292
R13885 VDD.n316 VDD.n225 0.120292
R13886 VDD.n317 VDD.n316 0.120292
R13887 VDD.n318 VDD.n223 0.120292
R13888 VDD.n322 VDD.n223 0.120292
R13889 VDD.n325 VDD.n323 0.120292
R13890 VDD.n31 VDD.n30 0.120292
R13891 VDD.n39 VDD.n38 0.120292
R13892 VDD.n48 VDD.n47 0.120292
R13893 VDD.n49 VDD.n48 0.120292
R13894 VDD.n54 VDD.n17 0.120292
R13895 VDD.n62 VDD.n14 0.120292
R13896 VDD.n63 VDD.n62 0.120292
R13897 VDD.n63 VDD.n11 0.120292
R13898 VDD.n70 VDD.n11 0.120292
R13899 VDD.n76 VDD.n9 0.120292
R13900 VDD.n77 VDD.n76 0.120292
R13901 VDD.n77 VDD.n6 0.120292
R13902 VDD.n81 VDD.n6 0.120292
R13903 VDD.n82 VDD.n81 0.120292
R13904 VDD.n82 VDD.n3 0.120292
R13905 VDD.n88 VDD.n3 0.120292
R13906 VDD.n89 VDD.n88 0.120292
R13907 VDD.n90 VDD.n89 0.120292
R13908 VDD.n95 VDD.n94 0.120292
R13909 VDD.n218 VDD.n217 0.119058
R13910 VDD.n345 VDD.n344 0.119058
R13911 VDD.n143 VDD 0.117487
R13912 VDD.n152 VDD 0.117487
R13913 VDD.n136 VDD 0.117222
R13914 VDD.n163 VDD 0.105191
R13915 VDD.t149 VDD 0.104171
R13916 VDD.n94 VDD 0.0994583
R13917 VDD.n251 VDD 0.0981562
R13918 VDD.n259 VDD 0.0981562
R13919 VDD.n30 VDD 0.0981562
R13920 VDD.n38 VDD 0.0981562
R13921 VDD.n268 VDD 0.0968542
R13922 VDD VDD.n235 0.0968542
R13923 VDD.n47 VDD 0.0968542
R13924 VDD VDD.n14 0.0968542
R13925 VDD.n147 VDD.n146 0.0914585
R13926 VDD.n156 VDD.n155 0.0914585
R13927 VDD.n161 VDD.n160 0.0888625
R13928 VDD.n164 VDD.n163 0.0878059
R13929 VDD.t144 VDD 0.0806706
R13930 VDD.t145 VDD 0.0806706
R13931 VDD.t149 VDD 0.0806706
R13932 VDD.t144 VDD 0.0805539
R13933 VDD.t145 VDD 0.0805539
R13934 VDD.t149 VDD 0.0805539
R13935 VDD.n165 VDD.n164 0.0799118
R13936 VDD.n245 VDD 0.0603958
R13937 VDD VDD.n252 0.0603958
R13938 VDD.n253 VDD 0.0603958
R13939 VDD VDD.n260 0.0603958
R13940 VDD.n261 VDD 0.0603958
R13941 VDD VDD.n238 0.0603958
R13942 VDD VDD.n276 0.0603958
R13943 VDD.n277 VDD 0.0603958
R13944 VDD VDD.n292 0.0603958
R13945 VDD.n293 VDD 0.0603958
R13946 VDD.n294 VDD 0.0603958
R13947 VDD VDD.n230 0.0603958
R13948 VDD.n318 VDD 0.0603958
R13949 VDD.n323 VDD 0.0603958
R13950 VDD VDD.n324 0.0603958
R13951 VDD.n332 VDD 0.0603958
R13952 VDD.n24 VDD 0.0603958
R13953 VDD VDD.n31 0.0603958
R13954 VDD.n32 VDD 0.0603958
R13955 VDD VDD.n39 0.0603958
R13956 VDD.n40 VDD 0.0603958
R13957 VDD VDD.n17 0.0603958
R13958 VDD VDD.n54 0.0603958
R13959 VDD.n55 VDD 0.0603958
R13960 VDD VDD.n70 0.0603958
R13961 VDD.n71 VDD 0.0603958
R13962 VDD.n72 VDD 0.0603958
R13963 VDD VDD.n9 0.0603958
R13964 VDD VDD.n1 0.0603958
R13965 VDD VDD.n95 0.0603958
R13966 VDD.n96 VDD 0.0603958
R13967 VDD.n138 VDD.n137 0.049413
R13968 VDD.n127 VDD 0.0482381
R13969 VDD.n135 VDD.n134 0.0466957
R13970 VDD.n143 VDD.n142 0.0466957
R13971 VDD.n143 VDD.n133 0.0466957
R13972 VDD.n152 VDD.n151 0.0466957
R13973 VDD.n152 VDD.n132 0.0466957
R13974 VDD.n125 VDD 0.0430763
R13975 VDD.n126 VDD 0.0430763
R13976 VDD.n163 VDD.n162 0.0394617
R13977 VDD.n128 VDD.n127 0.0390868
R13978 VDD VDD.n293 0.0382604
R13979 VDD VDD.n71 0.0382604
R13980 VDD.n168 VDD.n167 0.0357941
R13981 VDD.n325 VDD 0.03175
R13982 VDD VDD.n332 0.03175
R13983 VDD.n96 VDD 0.03175
R13984 VDD VDD.n99 0.03175
R13985 VDD.n166 VDD.n131 0.0294373
R13986 VDD.n164 VDD.n161 0.0287781
R13987 VDD.n270 VDD 0.0278438
R13988 VDD.n294 VDD 0.0278438
R13989 VDD VDD.n317 0.0278438
R13990 VDD.n49 VDD 0.0278438
R13991 VDD.n72 VDD 0.0278438
R13992 VDD.n90 VDD 0.0278438
R13993 VDD.n137 VDD.n136 0.0270767
R13994 VDD.n125 VDD.t149 0.024
R13995 VDD.n126 VDD.t145 0.024
R13996 VDD.t145 VDD.n125 0.024
R13997 VDD.n128 VDD.t144 0.024
R13998 VDD.t144 VDD.n126 0.024
R13999 VDD.n261 VDD 0.0239375
R14000 VDD.n277 VDD 0.0239375
R14001 VDD VDD.n322 0.0239375
R14002 VDD.n40 VDD 0.0239375
R14003 VDD.n55 VDD 0.0239375
R14004 VDD.n178 VDD.n177 0.0233549
R14005 VDD.n174 VDD.n171 0.0233549
R14006 VDD.n123 VDD.n122 0.0233549
R14007 VDD.n245 VDD 0.0226354
R14008 VDD.n253 VDD 0.0226354
R14009 VDD.n324 VDD 0.0226354
R14010 VDD.n24 VDD 0.0226354
R14011 VDD.n32 VDD 0.0226354
R14012 VDD.n205 VDD.n203 0.0222634
R14013 VDD.n214 VDD.n213 0.0222634
R14014 VDD.n1 VDD 0.0213333
R14015 VDD.n146 VDD 0.0209545
R14016 VDD.n155 VDD 0.0209545
R14017 VDD.n144 VDD 0.0150455
R14018 VDD.n153 VDD 0.0150455
R14019 VDD.n130 VDD.n129 0.0137706
R14020 VDD.n209 VDD.n207 0.0101288
R14021 VDD.n215 VDD.n212 0.00918401
R14022 VDD.n206 VDD.n202 0.00868304
R14023 VDD.n129 VDD.n128 0.0073069
R14024 VDD.n351 VDD.n218 0.00633075
R14025 VDD.n350 VDD.n345 0.0052
R14026 VDD.n343 VDD.n342 0.0052
R14027 VDD.n344 VDD.n343 0.0050825
R14028 VDD.n138 VDD.n135 0.00321739
R14029 VDD.n142 VDD.n141 0.00321739
R14030 VDD.n147 VDD.n133 0.00321739
R14031 VDD.n151 VDD.n150 0.00321739
R14032 VDD.n156 VDD.n132 0.00321739
R14033 VDD.n160 VDD.n159 0.00321739
R14034 VDD.n341 VDD.n337 0.00298917
R14035 VDD.n220 VDD.n219 0.00298831
R14036 VDD.n146 VDD.n145 0.00239442
R14037 VDD.n155 VDD.n154 0.00239442
R14038 VDD.n341 VDD.n340 0.00201061
R14039 VDD.n336 VDD.n335 0.00152605
R14040 VDD.n343 VDD.n336 0.00151551
R14041 VDD.n190 VDD.n189 0.00125069
R14042 VDD.n105 VDD.n104 0.00125069
R14043 VDD.n216 VDD.n215 0.0011527
R14044 VDD.n182 VDD.n181 0.00109775
R14045 VDD.n350 VDD.n349 0.00102396
R14046 VDD.n217 VDD.n201 0.00101664
R14047 VDD.n209 VDD.n208 0.00101293
R14048 VDD.n352 VDD.n351 0.00101239
R14049 VDD.n211 VDD.n209 0.00101167
R14050 VDD.n351 VDD.n350 0.00101141
R14051 VDD.n350 VDD.n220 0.00100941
R14052 VDD.n343 VDD.n341 0.00100876
R14053 VDD.n339 VDD.n338 0.00100479
R14054 VDD.n215 VDD.n214 0.00100265
R14055 VDD.n347 VDD.n346 0.00100208
R14056 VDD.n189 VDD.n188 0.00100206
R14057 VDD.n349 VDD.n348 0.0010004
R14058 VDD.n145 VDD.n144 0.0010003
R14059 VDD.n154 VDD.n153 0.0010003
R14060 VDD.n201 VDD.n200 0.00100002
R14061 VDD.n183 VDD.n180 0.000990196
R14062 VDD.n169 VDD.n168 0.000990196
R14063 VDD.n101 VDD.n100 0.000990196
R14064 VDD.n197 VDD.n109 0.000990196
R14065 VDD.n211 VDD.n206 0.000709821
R14066 VDD.n177 VDD.n174 0.000684314
R14067 VDD.n171 VDD.n166 0.000684314
R14068 VDD.n124 VDD.n123 0.000684314
R14069 VDD.n119 VDD.n116 0.000684314
R14070 VDD.n187 VDD.n186 0.000684314
R14071 VDD.n217 VDD.n216 0.000517546
R14072 VDD.n217 VDD.n211 0.000517191
R14073 VDD.n177 VDD.n124 0.000516685
R14074 VDD.n166 VDD.n130 0.000516685
R14075 VDD.n195 VDD.n194 0.000516685
R14076 VDD.n194 VDD.n111 0.000516685
R14077 VDD.n191 VDD.n187 0.000516685
R14078 VDD.n116 VDD.n115 0.000516685
R14079 VDD.n191 VDD.n119 0.000516685
R14080 VDD.n191 VDD.n190 0.000516685
R14081 VDD.n115 VDD.n114 0.000516685
R14082 VDD.n106 VDD.n103 0.000516685
R14083 VDD.n194 VDD.n193 0.000516685
R14084 VDD.n106 VDD.n105 0.000516685
R14085 VDD.n107 VDD.n106 0.000516685
R14086 VDD.n211 VDD.n210 0.000512596
R14087 VDD.n348 VDD.n347 0.000505632
R14088 VDD.n335 VDD.n334 0.000505632
R14089 VDD.n340 VDD.n339 0.000505632
R14090 VDD.n353 VDD.n352 0.000505632
R14091 VDD.n177 VDD.n176 0.000505597
R14092 VDD.n171 VDD.n170 0.000505597
R14093 VDD.n179 VDD.n178 0.000505597
R14094 VDD.n174 VDD.n173 0.000505597
R14095 VDD.n166 VDD.n165 0.000505597
R14096 VDD.n116 VDD.n113 0.000505597
R14097 VDD.n187 VDD.n121 0.000505597
R14098 VDD.n186 VDD.n185 0.000505597
R14099 VDD.n119 VDD.n118 0.000505597
R14100 VDD.n193 VDD.n192 0.000505597
R14101 VDD.n196 VDD.n195 0.000505597
R14102 VDD.n111 VDD.n110 0.000505597
R14103 VDD.n103 VDD.n102 0.000505597
R14104 VDD.n108 VDD.n107 0.000505597
R14105 VDD.n334 VDD.n333 0.000504168
R14106 VDD.n354 VDD.n353 0.000504168
R14107 VDD.n176 VDD.n175 0.000504146
R14108 VDD.n170 VDD.n169 0.000504146
R14109 VDD.n180 VDD.n179 0.000504146
R14110 VDD.n173 VDD.n172 0.000504146
R14111 VDD.n183 VDD.n182 0.000504146
R14112 VDD.n113 VDD.n112 0.000504146
R14113 VDD.n185 VDD.n184 0.000504146
R14114 VDD.n121 VDD.n120 0.000504146
R14115 VDD.n118 VDD.n117 0.000504146
R14116 VDD.n197 VDD.n196 0.000504146
R14117 VDD.n102 VDD.n101 0.000504146
R14118 VDD.n109 VDD.n108 0.000504146
R14119 VDD.n206 VDD.n205 0.000503644
R14120 VDD.n200 VDD.n199 0.000502799
R14121 VDD.n199 VDD.n198 0.000502073
R14122 VDD.n205 VDD.n204 0.000502073
R14123 mimtop1.n51 mimtop1.t4 112.793
R14124 mimtop1.n52 mimtop1.t5 112.416
R14125 mimtop1.n47 mimtop1.n46 109.123
R14126 mimtop1.n52 mimtop1.t1 83.3917
R14127 mimtop1.n51 mimtop1.t0 83.0152
R14128 mimtop1.n48 mimtop1.n47 67.1128
R14129 mimtop1.n46 mimtop1.t3 57.1305
R14130 mimtop1.n46 mimtop1.t2 57.1305
R14131 mimtop1.n45 mimtop1.t6 34.8005
R14132 mimtop1.n45 mimtop1.t7 34.8005
R14133 mimtop1.n54 mimtop1.n53 4.73357
R14134 mimtop1.n66 mimtop1.n65 1.26526
R14135 mimtop1.n71 mimtop1.n70 1.14123
R14136 mimtop1.n53 mimtop1.n51 0.602099
R14137 mimtop1.n38 mimtop1.n37 0.345941
R14138 mimtop1.n6 mimtop1 0.104839
R14139 mimtop1.n6 mimtop1 0.104839
R14140 mimtop1.n6 mimtop1 0.104839
R14141 mimtop1.n6 mimtop1 0.104839
R14142 mimtop1.n6 mimtop1 0.104839
R14143 mimtop1.n6 mimtop1 0.104839
R14144 mimtop1.n6 mimtop1 0.104839
R14145 mimtop1.n6 mimtop1 0.104839
R14146 mimtop1.n36 mimtop1 0.104171
R14147 mimtop1.n36 mimtop1 0.104171
R14148 mimtop1.n36 mimtop1 0.104171
R14149 mimtop1.n36 mimtop1 0.104171
R14150 mimtop1.n36 mimtop1 0.104171
R14151 mimtop1.n36 mimtop1 0.104171
R14152 mimtop1.n36 mimtop1 0.104171
R14153 mimtop1.n36 mimtop1 0.104171
R14154 mimtop1.n47 mimtop1.n45 0.10226
R14155 mimtop1.n13 mimtop1 0.0806706
R14156 mimtop1.n20 mimtop1 0.0806706
R14157 mimtop1.n27 mimtop1 0.0806706
R14158 mimtop1.n6 mimtop1 0.0805539
R14159 mimtop1.n13 mimtop1 0.0805539
R14160 mimtop1.n20 mimtop1 0.0805539
R14161 mimtop1.n27 mimtop1 0.0805539
R14162 mimtop1.n36 mimtop1 0.0805539
R14163 mimtop1.n6 mimtop1 0.0796706
R14164 mimtop1.n37 mimtop1.n36 0.045459
R14165 mimtop1.n35 mimtop1 0.0430763
R14166 mimtop1.n26 mimtop1 0.0430763
R14167 mimtop1.n19 mimtop1 0.0430763
R14168 mimtop1.n12 mimtop1 0.0430763
R14169 mimtop1.n11 mimtop1 0.0430763
R14170 mimtop1.n18 mimtop1 0.0430763
R14171 mimtop1.n25 mimtop1 0.0430763
R14172 mimtop1.n34 mimtop1 0.0430763
R14173 mimtop1.n28 mimtop1 0.0430763
R14174 mimtop1.n24 mimtop1 0.0430763
R14175 mimtop1.n17 mimtop1 0.0430763
R14176 mimtop1.n10 mimtop1 0.0430763
R14177 mimtop1.n9 mimtop1 0.0430763
R14178 mimtop1.n16 mimtop1 0.0430763
R14179 mimtop1.n23 mimtop1 0.0430763
R14180 mimtop1.n29 mimtop1 0.0430763
R14181 mimtop1.n33 mimtop1 0.0430763
R14182 mimtop1.n22 mimtop1 0.0430763
R14183 mimtop1.n15 mimtop1 0.0430763
R14184 mimtop1.n8 mimtop1 0.0430763
R14185 mimtop1.n7 mimtop1 0.0430763
R14186 mimtop1.n14 mimtop1 0.0430763
R14187 mimtop1.n21 mimtop1 0.0430763
R14188 mimtop1.n32 mimtop1 0.0430763
R14189 mimtop1.n30 mimtop1 0.0430763
R14190 mimtop1.n1 mimtop1 0.0430763
R14191 mimtop1.n3 mimtop1 0.0430763
R14192 mimtop1.n5 mimtop1 0.0430763
R14193 mimtop1.n31 mimtop1 0.0419101
R14194 mimtop1.n6 mimtop1 0.0417933
R14195 mimtop1.n6 mimtop1 0.0417933
R14196 mimtop1.n6 mimtop1 0.0417933
R14197 mimtop1.n6 mimtop1 0.0417933
R14198 mimtop1.n6 mimtop1 0.0417933
R14199 mimtop1.n6 mimtop1 0.0417933
R14200 mimtop1.n6 mimtop1 0.0417933
R14201 mimtop1.n13 mimtop1 0.0409101
R14202 mimtop1.n13 mimtop1 0.0409101
R14203 mimtop1.n13 mimtop1 0.0409101
R14204 mimtop1.n13 mimtop1 0.0409101
R14205 mimtop1.n13 mimtop1 0.0409101
R14206 mimtop1.n13 mimtop1 0.0409101
R14207 mimtop1.n13 mimtop1 0.0409101
R14208 mimtop1.n20 mimtop1 0.0409101
R14209 mimtop1.n20 mimtop1 0.0409101
R14210 mimtop1.n20 mimtop1 0.0409101
R14211 mimtop1.n20 mimtop1 0.0409101
R14212 mimtop1.n20 mimtop1 0.0409101
R14213 mimtop1.n20 mimtop1 0.0409101
R14214 mimtop1.n20 mimtop1 0.0409101
R14215 mimtop1.n27 mimtop1 0.0409101
R14216 mimtop1.n27 mimtop1 0.0409101
R14217 mimtop1.n27 mimtop1 0.0409101
R14218 mimtop1.n27 mimtop1 0.0409101
R14219 mimtop1.n27 mimtop1 0.0409101
R14220 mimtop1.n27 mimtop1 0.0409101
R14221 mimtop1.n27 mimtop1 0.0409101
R14222 mimtop1.n36 mimtop1 0.0409101
R14223 mimtop1.n36 mimtop1 0.0409101
R14224 mimtop1.n36 mimtop1 0.0409101
R14225 mimtop1.n36 mimtop1 0.0409101
R14226 mimtop1.n36 mimtop1 0.0409101
R14227 mimtop1.n36 mimtop1 0.0409101
R14228 mimtop1.n36 mimtop1 0.0409101
R14229 mimtop1.n4 mimtop1 0.0409101
R14230 mimtop1.n2 mimtop1 0.0409101
R14231 mimtop1.n0 mimtop1 0.0409101
R14232 mimtop1.n37 mimtop1 0.0355945
R14233 mimtop1.n72 mimtop1.n71 0.0326167
R14234 mimtop1.n36 mimtop1.n35 0.024
R14235 mimtop1.n27 mimtop1.n26 0.024
R14236 mimtop1.n20 mimtop1.n19 0.024
R14237 mimtop1.n13 mimtop1.n12 0.024
R14238 mimtop1.n13 mimtop1.n11 0.024
R14239 mimtop1.n20 mimtop1.n18 0.024
R14240 mimtop1.n27 mimtop1.n25 0.024
R14241 mimtop1.n36 mimtop1.n34 0.024
R14242 mimtop1.n36 mimtop1.n28 0.024
R14243 mimtop1.n27 mimtop1.n24 0.024
R14244 mimtop1.n28 mimtop1.n27 0.024
R14245 mimtop1.n20 mimtop1.n17 0.024
R14246 mimtop1.n13 mimtop1.n10 0.024
R14247 mimtop1.n13 mimtop1.n9 0.024
R14248 mimtop1.n20 mimtop1.n16 0.024
R14249 mimtop1.n27 mimtop1.n23 0.024
R14250 mimtop1.n36 mimtop1.n29 0.024
R14251 mimtop1.n36 mimtop1.n33 0.024
R14252 mimtop1.n27 mimtop1.n22 0.024
R14253 mimtop1.n20 mimtop1.n15 0.024
R14254 mimtop1.n13 mimtop1.n8 0.024
R14255 mimtop1.n7 mimtop1.n6 0.024
R14256 mimtop1.n13 mimtop1.n7 0.024
R14257 mimtop1.n14 mimtop1.n13 0.024
R14258 mimtop1.n20 mimtop1.n14 0.024
R14259 mimtop1.n21 mimtop1.n20 0.024
R14260 mimtop1.n27 mimtop1.n21 0.024
R14261 mimtop1.n36 mimtop1.n32 0.024
R14262 mimtop1.n36 mimtop1.n30 0.024
R14263 mimtop1.n27 mimtop1.n1 0.024
R14264 mimtop1.n20 mimtop1.n3 0.024
R14265 mimtop1.n13 mimtop1.n5 0.024
R14266 mimtop1.n13 mimtop1.n4 0.024
R14267 mimtop1.n20 mimtop1.n2 0.024
R14268 mimtop1.n27 mimtop1.n0 0.024
R14269 mimtop1.n36 mimtop1.n31 0.024
R14270 mimtop1.n60 mimtop1.n59 0.0224263
R14271 mimtop1.n57 mimtop1.n56 0.01925
R14272 mimtop1.n63 mimtop1.n62 0.01925
R14273 mimtop1.n72 mimtop1.n41 0.0174148
R14274 mimtop1.n41 mimtop1.n40 0.0150648
R14275 mimtop1.n56 mimtop1.n55 0.0134654
R14276 mimtop1.n66 mimtop1.n44 0.0133252
R14277 mimtop1.n53 mimtop1.n52 0.0125466
R14278 mimtop1.n67 mimtop1.n66 0.0121627
R14279 mimtop1.n50 mimtop1.n49 0.0099718
R14280 mimtop1.n61 mimtop1.n60 0.0099718
R14281 mimtop1.n43 mimtop1.n42 0.00847576
R14282 mimtop1.n69 mimtop1.n68 0.00847576
R14283 mimtop1.n58 mimtop1.n57 0.00496429
R14284 mimtop1.n64 mimtop1.n63 0.00496429
R14285 mimtop1.n65 mimtop1.n61 0.00478082
R14286 mimtop1.n54 mimtop1.n50 0.00478082
R14287 mimtop1.n73 mimtop1.n72 0.00392883
R14288 mimtop1 mimtop1.n74 0.00300672
R14289 mimtop1.n72 mimtop1.n39 0.00275583
R14290 mimtop1.n39 mimtop1.n38 0.00250494
R14291 mimtop1.n74 mimtop1.n73 0.00250494
R14292 mimtop1.n70 mimtop1.n67 0.00175815
R14293 mimtop1.n44 mimtop1.n43 0.00163939
R14294 mimtop1.n70 mimtop1.n69 0.00138099
R14295 mimtop1.n58 mimtop1.n48 0.00100108
R14296 mimtop1.n65 mimtop1.n58 0.000687305
R14297 mimtop1.n58 mimtop1.n54 0.000687305
R14298 mimtop1.n65 mimtop1.n64 0.000687305
R14299 mimtop1.n36 mimtop1.t45 0.000499999
R14300 mimtop1.n27 mimtop1.t37 0.000499999
R14301 mimtop1.n20 mimtop1.t31 0.000499999
R14302 mimtop1.n13 mimtop1.t17 0.000499999
R14303 mimtop1.n6 mimtop1.t8 0.000499999
R14304 mimtop1.n6 mimtop1.t23 0.000499999
R14305 mimtop1.n13 mimtop1.t30 0.000499999
R14306 mimtop1.n20 mimtop1.t44 0.000499999
R14307 mimtop1.n27 mimtop1.t12 0.000499999
R14308 mimtop1.n36 mimtop1.t19 0.000499999
R14309 mimtop1.n36 mimtop1.t28 0.000499999
R14310 mimtop1.n27 mimtop1.t22 0.000499999
R14311 mimtop1.n20 mimtop1.t16 0.000499999
R14312 mimtop1.n13 mimtop1.t41 0.000499999
R14313 mimtop1.n6 mimtop1.t34 0.000499999
R14314 mimtop1.n6 mimtop1.t46 0.000499999
R14315 mimtop1.n13 mimtop1.t13 0.000499999
R14316 mimtop1.n20 mimtop1.t27 0.000499999
R14317 mimtop1.n27 mimtop1.t33 0.000499999
R14318 mimtop1.n36 mimtop1.t40 0.000499999
R14319 mimtop1.n36 mimtop1.t14 0.000499999
R14320 mimtop1.n27 mimtop1.t47 0.000499999
R14321 mimtop1.n20 mimtop1.t39 0.000499999
R14322 mimtop1.n13 mimtop1.t26 0.000499999
R14323 mimtop1.n6 mimtop1.t20 0.000499999
R14324 mimtop1.n6 mimtop1.t29 0.000499999
R14325 mimtop1.n13 mimtop1.t36 0.000499999
R14326 mimtop1.n20 mimtop1.t11 0.000499999
R14327 mimtop1.n27 mimtop1.t18 0.000499999
R14328 mimtop1.n36 mimtop1.t25 0.000499999
R14329 mimtop1.n36 mimtop1.t38 0.000499999
R14330 mimtop1.n27 mimtop1.t32 0.000499999
R14331 mimtop1.n20 mimtop1.t24 0.000499999
R14332 mimtop1.n13 mimtop1.t10 0.000499999
R14333 mimtop1.n6 mimtop1.t43 0.000499999
R14334 mimtop1.n6 mimtop1.t15 0.000499999
R14335 mimtop1.n13 mimtop1.t21 0.000499999
R14336 mimtop1.n20 mimtop1.t35 0.000499999
R14337 mimtop1.n27 mimtop1.t42 0.000499999
R14338 mimtop1.n36 mimtop1.t9 0.000499999
R14339 mimbot1.n10 mimbot1.t45 112.416
R14340 mimbot1.n9 mimbot1.t44 109.835
R14341 mimbot1.n3 mimbot1.n1 108.15
R14342 mimbot1.n9 mimbot1.t1 82.5823
R14343 mimbot1.n2 mimbot1.t43 57.1305
R14344 mimbot1.n2 mimbot1.t42 57.1305
R14345 mimbot1.n11 mimbot1.n10 47.8363
R14346 mimbot1.n11 mimbot1.t0 34.9023
R14347 mimbot1.n1 mimbot1.t47 34.8005
R14348 mimbot1.n1 mimbot1.t46 34.8005
R14349 mimbot1.n12 mimbot1.n11 24.469
R14350 mimbot1.n725 mimbot1.n26 2.24852
R14351 mimbot1.n4 mimbot1.n3 2.1391
R14352 mimbot1.n25 mimbot1.n24 2.04132
R14353 mimbot1.n6 mimbot1.n0 1.7055
R14354 mimbot1.n26 mimbot1.n25 1.7055
R14355 mimbot1.n10 mimbot1.n9 0.606804
R14356 mimbot1.n725 mimbot1 0.530984
R14357 mimbot1.n724 mimbot1 0.0953952
R14358 mimbot1.n724 mimbot1 0.0936132
R14359 mimbot1.n80 mimbot1.n79 0.0659051
R14360 mimbot1.n75 mimbot1.n74 0.0659051
R14361 mimbot1.n103 mimbot1.n102 0.0659051
R14362 mimbot1.n99 mimbot1.n98 0.0659051
R14363 mimbot1.n126 mimbot1.n125 0.0659051
R14364 mimbot1.n122 mimbot1.n121 0.0659051
R14365 mimbot1.n143 mimbot1.n142 0.0659051
R14366 mimbot1.n597 mimbot1.n596 0.0659051
R14367 mimbot1.n605 mimbot1.n604 0.0659051
R14368 mimbot1.n612 mimbot1.n611 0.0659051
R14369 mimbot1.n631 mimbot1.n630 0.0659051
R14370 mimbot1.n644 mimbot1.n643 0.0659051
R14371 mimbot1.n651 mimbot1.n650 0.0659051
R14372 mimbot1.n663 mimbot1.n662 0.0659051
R14373 mimbot1.n679 mimbot1.n678 0.0659051
R14374 mimbot1.n570 mimbot1.n476 0.0659051
R14375 mimbot1.n424 mimbot1.n354 0.0659051
R14376 mimbot1.n702 mimbot1.n268 0.0659051
R14377 mimbot1.n586 mimbot1.n580 0.0659051
R14378 mimbot1.n584 mimbot1.n582 0.0659051
R14379 mimbot1.n518 mimbot1.n468 0.0659051
R14380 mimbot1.n387 mimbot1.n348 0.0659051
R14381 mimbot1.n306 mimbot1.n248 0.0659051
R14382 mimbot1.n228 mimbot1.n38 0.0659051
R14383 mimbot1.n139 mimbot1.n138 0.0659051
R14384 mimbot1.n632 mimbot1.n622 0.05126
R14385 mimbot1.n645 mimbot1.n635 0.05126
R14386 mimbot1.n652 mimbot1.n619 0.05126
R14387 mimbot1.n664 mimbot1.n658 0.05126
R14388 mimbot1.n680 mimbot1.n670 0.05126
R14389 mimbot1.n613 mimbot1.n608 0.05126
R14390 mimbot1.n681 mimbot1.n603 0.05126
R14391 mimbot1.n692 mimbot1.n475 0.05126
R14392 mimbot1.n695 mimbot1.n355 0.05126
R14393 mimbot1.n718 mimbot1.n267 0.05126
R14394 mimbot1.n598 mimbot1.n588 0.05126
R14395 mimbot1.n583 mimbot1.n577 0.05126
R14396 mimbot1.n681 mimbot1.n587 0.05126
R14397 mimbot1.n692 mimbot1.n469 0.05126
R14398 mimbot1.n695 mimbot1.n349 0.05126
R14399 mimbot1.n718 mimbot1.n249 0.05126
R14400 mimbot1.n723 mimbot1.n37 0.05126
R14401 mimbot1.n150 mimbot1.n136 0.05126
R14402 mimbot1.n144 mimbot1.n53 0.05126
R14403 mimbot1.n133 mimbot1.n113 0.05126
R14404 mimbot1.n127 mimbot1.n56 0.05126
R14405 mimbot1.n110 mimbot1.n90 0.05126
R14406 mimbot1.n104 mimbot1.n59 0.05126
R14407 mimbot1.n87 mimbot1.n66 0.05126
R14408 mimbot1.n81 mimbot1.n78 0.05126
R14409 mimbot1.n723 mimbot1.n722 0.05126
R14410 mimbot1.n62 mimbot1 0.0475
R14411 mimbot1.n76 mimbot1 0.0475
R14412 mimbot1.n68 mimbot1 0.0475
R14413 mimbot1.n100 mimbot1 0.0475
R14414 mimbot1.n92 mimbot1 0.0475
R14415 mimbot1.n123 mimbot1 0.0475
R14416 mimbot1.n115 mimbot1 0.0475
R14417 mimbot1.n140 mimbot1 0.0475
R14418 mimbot1.n590 mimbot1 0.0475
R14419 mimbot1.n157 mimbot1 0.0475
R14420 mimbot1.n606 mimbot1 0.0475
R14421 mimbot1.n609 mimbot1 0.0475
R14422 mimbot1.n624 mimbot1 0.0475
R14423 mimbot1.n637 mimbot1 0.0475
R14424 mimbot1.n648 mimbot1 0.0475
R14425 mimbot1.n660 mimbot1 0.0475
R14426 mimbot1.n672 mimbot1 0.0475
R14427 mimbot1.n574 mimbot1 0.0475
R14428 mimbot1.n422 mimbot1 0.0475
R14429 mimbot1.n699 mimbot1 0.0475
R14430 mimbot1.n521 mimbot1 0.0475
R14431 mimbot1.n390 mimbot1 0.0475
R14432 mimbot1.n309 mimbot1 0.0475
R14433 mimbot1.n231 mimbot1 0.0475
R14434 mimbot1.n79 mimbot1 0.0439131
R14435 mimbot1.n75 mimbot1 0.0439131
R14436 mimbot1.n102 mimbot1 0.0439131
R14437 mimbot1.n99 mimbot1 0.0439131
R14438 mimbot1.n125 mimbot1 0.0439131
R14439 mimbot1.n122 mimbot1 0.0439131
R14440 mimbot1.n142 mimbot1 0.0439131
R14441 mimbot1.n597 mimbot1 0.0439131
R14442 mimbot1.n604 mimbot1 0.0439131
R14443 mimbot1.n611 mimbot1 0.0439131
R14444 mimbot1.n631 mimbot1 0.0439131
R14445 mimbot1.n644 mimbot1 0.0439131
R14446 mimbot1.n650 mimbot1 0.0439131
R14447 mimbot1.n662 mimbot1 0.0439131
R14448 mimbot1.n679 mimbot1 0.0439131
R14449 mimbot1.n476 mimbot1 0.0439131
R14450 mimbot1.n354 mimbot1 0.0439131
R14451 mimbot1.n268 mimbot1 0.0439131
R14452 mimbot1.n580 mimbot1 0.0439131
R14453 mimbot1.n582 mimbot1 0.0439131
R14454 mimbot1.n468 mimbot1 0.0439131
R14455 mimbot1.n348 mimbot1 0.0439131
R14456 mimbot1.n248 mimbot1 0.0439131
R14457 mimbot1.n38 mimbot1 0.0439131
R14458 mimbot1.n139 mimbot1 0.0439131
R14459 mimbot1.n608 mimbot1.n607 0.0422331
R14460 mimbot1.n151 mimbot1.n52 0.0383507
R14461 mimbot1.n626 mimbot1.n623 0.0367203
R14462 mimbot1.n639 mimbot1.n636 0.0367203
R14463 mimbot1.n657 mimbot1.n656 0.0367203
R14464 mimbot1.n669 mimbot1.n668 0.0367203
R14465 mimbot1.n674 mimbot1.n671 0.0367203
R14466 mimbot1.n618 mimbot1.n617 0.0367203
R14467 mimbot1.n592 mimbot1.n589 0.0367203
R14468 mimbot1.n149 mimbot1.n148 0.0367203
R14469 mimbot1.n117 mimbot1.n114 0.0367203
R14470 mimbot1.n132 mimbot1.n131 0.0367203
R14471 mimbot1.n94 mimbot1.n91 0.0367203
R14472 mimbot1.n109 mimbot1.n108 0.0367203
R14473 mimbot1.n70 mimbot1.n67 0.0367203
R14474 mimbot1.n86 mimbot1.n85 0.0367203
R14475 mimbot1.n724 mimbot1.n27 0.0365333
R14476 mimbot1.n628 mimbot1.n622 0.03622
R14477 mimbot1.n641 mimbot1.n635 0.03622
R14478 mimbot1.n653 mimbot1.n652 0.03622
R14479 mimbot1.n665 mimbot1.n664 0.03622
R14480 mimbot1.n676 mimbot1.n670 0.03622
R14481 mimbot1.n614 mimbot1.n613 0.03622
R14482 mimbot1.n594 mimbot1.n588 0.03622
R14483 mimbot1.n145 mimbot1.n144 0.03622
R14484 mimbot1.n119 mimbot1.n113 0.03622
R14485 mimbot1.n128 mimbot1.n127 0.03622
R14486 mimbot1.n96 mimbot1.n90 0.03622
R14487 mimbot1.n105 mimbot1.n104 0.03622
R14488 mimbot1.n72 mimbot1.n66 0.03622
R14489 mimbot1.n82 mimbot1.n81 0.03622
R14490 mimbot1.n136 mimbot1.n52 0.0335645
R14491 mimbot1.n406 mimbot1.n371 0.0334526
R14492 mimbot1.n407 mimbot1.n351 0.0334526
R14493 mimbot1.n219 mimbot1.n41 0.0334526
R14494 mimbot1.n217 mimbot1.n216 0.0334526
R14495 mimbot1.n284 mimbot1.n283 0.0334526
R14496 mimbot1.n286 mimbot1.n251 0.0334526
R14497 mimbot1.n274 mimbot1.n273 0.0334526
R14498 mimbot1.n275 mimbot1.n262 0.0334526
R14499 mimbot1.n327 mimbot1.n326 0.0334526
R14500 mimbot1.n328 mimbot1.n254 0.0334526
R14501 mimbot1.n378 mimbot1.n346 0.0334526
R14502 mimbot1.n377 mimbot1.n376 0.0334526
R14503 mimbot1.n397 mimbot1.n396 0.0334526
R14504 mimbot1.n398 mimbot1.n365 0.0334526
R14505 mimbot1.n417 mimbot1.n368 0.0334526
R14506 mimbot1.n416 mimbot1.n415 0.0334526
R14507 mimbot1.n496 mimbot1.n495 0.0334526
R14508 mimbot1.n498 mimbot1.n471 0.0334526
R14509 mimbot1.n686 mimbot1.n685 0.0334526
R14510 mimbot1.n690 mimbot1.n488 0.0334526
R14511 mimbot1.n540 mimbot1.n479 0.0334526
R14512 mimbot1.n539 mimbot1.n538 0.0334526
R14513 mimbot1.n562 mimbot1.n482 0.0334526
R14514 mimbot1.n561 mimbot1.n560 0.0334526
R14515 mimbot1.n550 mimbot1.n549 0.0334526
R14516 mimbot1.n551 mimbot1.n485 0.0334526
R14517 mimbot1.n529 mimbot1.n474 0.0334526
R14518 mimbot1.n527 mimbot1.n526 0.0334526
R14519 mimbot1.n448 mimbot1.n359 0.0334526
R14520 mimbot1.n447 mimbot1.n446 0.0334526
R14521 mimbot1.n437 mimbot1.n363 0.0334526
R14522 mimbot1.n436 mimbot1.n435 0.0334526
R14523 mimbot1.n459 mimbot1.n356 0.0334526
R14524 mimbot1.n457 mimbot1.n456 0.0334526
R14525 mimbot1.n710 mimbot1.n266 0.0334526
R14526 mimbot1.n716 mimbot1.n715 0.0334526
R14527 mimbot1.n239 mimbot1.n50 0.0334526
R14528 mimbot1.n238 mimbot1.n237 0.0334526
R14529 mimbot1.n164 mimbot1.n30 0.0334526
R14530 mimbot1.n163 mimbot1.n162 0.0334526
R14531 mimbot1.n339 mimbot1.n256 0.0334526
R14532 mimbot1.n337 mimbot1.n336 0.0334526
R14533 mimbot1.n175 mimbot1.n47 0.0334526
R14534 mimbot1.n173 mimbot1.n172 0.0334526
R14535 mimbot1.n186 mimbot1.n33 0.0334526
R14536 mimbot1.n184 mimbot1.n183 0.0334526
R14537 mimbot1.n317 mimbot1.n260 0.0334526
R14538 mimbot1.n315 mimbot1.n314 0.0334526
R14539 mimbot1.n208 mimbot1.n44 0.0334526
R14540 mimbot1.n207 mimbot1.n206 0.0334526
R14541 mimbot1.n197 mimbot1.n36 0.0334526
R14542 mimbot1.n196 mimbot1.n195 0.0334526
R14543 mimbot1.n297 mimbot1.n246 0.0334526
R14544 mimbot1.n295 mimbot1.n294 0.0334526
R14545 mimbot1.n509 mimbot1.n466 0.0334526
R14546 mimbot1.n507 mimbot1.n506 0.0334526
R14547 mimbot1.n583 mimbot1.n581 0.03246
R14548 mimbot1.n682 mimbot1.n522 0.0309349
R14549 mimbot1.n693 mimbot1.n391 0.0309349
R14550 mimbot1.n696 mimbot1.n310 0.0309349
R14551 mimbot1.n719 mimbot1.n232 0.0309349
R14552 mimbot1.n720 mimbot1.n719 0.0303642
R14553 mimbot1.n623 mimbot1.n598 0.0303642
R14554 mimbot1.n636 mimbot1.n632 0.0303642
R14555 mimbot1.n658 mimbot1.n657 0.0303642
R14556 mimbot1.n680 mimbot1.n669 0.0303642
R14557 mimbot1.n671 mimbot1.n645 0.0303642
R14558 mimbot1.n619 mimbot1.n618 0.0303642
R14559 mimbot1.n682 mimbot1.n575 0.0303642
R14560 mimbot1.n693 mimbot1.n430 0.0303642
R14561 mimbot1.n700 mimbot1.n696 0.0303642
R14562 mimbot1.n589 mimbot1.n577 0.0303642
R14563 mimbot1.n150 mimbot1.n149 0.0303642
R14564 mimbot1.n114 mimbot1.n53 0.0303642
R14565 mimbot1.n133 mimbot1.n132 0.0303642
R14566 mimbot1.n91 mimbot1.n56 0.0303642
R14567 mimbot1.n110 mimbot1.n109 0.0303642
R14568 mimbot1.n67 mimbot1.n59 0.0303642
R14569 mimbot1.n87 mimbot1.n86 0.0303642
R14570 mimbot1.n23 mimbot1.n22 0.0295323
R14571 mimbot1.n695 mimbot1.n344 0.02588
R14572 mimbot1.n218 mimbot1.n40 0.02588
R14573 mimbot1.n152 mimbot1.n51 0.02588
R14574 mimbot1.n718 mimbot1.n244 0.02588
R14575 mimbot1.n374 mimbot1.n350 0.02588
R14576 mimbot1.n695 mimbot1.n366 0.02588
R14577 mimbot1.n695 mimbot1.n367 0.02588
R14578 mimbot1.n414 mimbot1.n361 0.02588
R14579 mimbot1.n394 mimbot1.n362 0.02588
R14580 mimbot1.n692 mimbot1.n464 0.02588
R14581 mimbot1.n681 mimbot1.n576 0.02588
R14582 mimbot1.n681 mimbot1.n600 0.02588
R14583 mimbot1.n681 mimbot1.n621 0.02588
R14584 mimbot1.n681 mimbot1.n634 0.02588
R14585 mimbot1.n681 mimbot1.n647 0.02588
R14586 mimbot1.n536 mimbot1.n480 0.02588
R14587 mimbot1.n558 mimbot1.n483 0.02588
R14588 mimbot1.n681 mimbot1.n601 0.02588
R14589 mimbot1.n572 mimbot1.n483 0.02588
R14590 mimbot1.n528 mimbot1.n477 0.02588
R14591 mimbot1.n692 mimbot1.n472 0.02588
R14592 mimbot1.n687 mimbot1.n478 0.02588
R14593 mimbot1.n692 mimbot1.n691 0.02588
R14594 mimbot1.n692 mimbot1.n487 0.02588
R14595 mimbot1.n423 mimbot1.n353 0.02588
R14596 mimbot1.n695 mimbot1.n360 0.02588
R14597 mimbot1.n444 mimbot1.n357 0.02588
R14598 mimbot1.n695 mimbot1.n364 0.02588
R14599 mimbot1.n433 mimbot1.n352 0.02588
R14600 mimbot1.n547 mimbot1.n481 0.02588
R14601 mimbot1.n692 mimbot1.n486 0.02588
R14602 mimbot1.n692 mimbot1.n484 0.02588
R14603 mimbot1.n458 mimbot1.n353 0.02588
R14604 mimbot1.n695 mimbot1.n358 0.02588
R14605 mimbot1.n717 mimbot1.n705 0.02588
R14606 mimbot1.n717 mimbot1.n706 0.02588
R14607 mimbot1.n718 mimbot1.n252 0.02588
R14608 mimbot1.n723 mimbot1.n28 0.02588
R14609 mimbot1.n235 mimbot1.n51 0.02588
R14610 mimbot1.n723 mimbot1.n49 0.02588
R14611 mimbot1.n160 mimbot1.n29 0.02588
R14612 mimbot1.n324 mimbot1.n265 0.02588
R14613 mimbot1.n338 mimbot1.n253 0.02588
R14614 mimbot1.n718 mimbot1.n264 0.02588
R14615 mimbot1.n718 mimbot1.n255 0.02588
R14616 mimbot1.n723 mimbot1.n31 0.02588
R14617 mimbot1.n174 mimbot1.n48 0.02588
R14618 mimbot1.n723 mimbot1.n46 0.02588
R14619 mimbot1.n185 mimbot1.n32 0.02588
R14620 mimbot1.n271 mimbot1.n257 0.02588
R14621 mimbot1.n316 mimbot1.n263 0.02588
R14622 mimbot1.n718 mimbot1.n258 0.02588
R14623 mimbot1.n718 mimbot1.n261 0.02588
R14624 mimbot1.n723 mimbot1.n34 0.02588
R14625 mimbot1.n204 mimbot1.n45 0.02588
R14626 mimbot1.n723 mimbot1.n43 0.02588
R14627 mimbot1.n193 mimbot1.n35 0.02588
R14628 mimbot1.n285 mimbot1.n259 0.02588
R14629 mimbot1.n296 mimbot1.n250 0.02588
R14630 mimbot1.n694 mimbot1.n370 0.02588
R14631 mimbot1.n497 mimbot1.n473 0.02588
R14632 mimbot1.n508 mimbot1.n470 0.02588
R14633 mimbot1.n681 mimbot1.n579 0.02588
R14634 mimbot1.n516 mimbot1.n465 0.02588
R14635 mimbot1.n692 mimbot1.n467 0.02588
R14636 mimbot1.n385 mimbot1.n345 0.02588
R14637 mimbot1.n695 mimbot1.n347 0.02588
R14638 mimbot1.n304 mimbot1.n245 0.02588
R14639 mimbot1.n718 mimbot1.n247 0.02588
R14640 mimbot1.n226 mimbot1.n42 0.02588
R14641 mimbot1.n723 mimbot1.n39 0.02588
R14642 mimbot1.n151 mimbot1.n134 0.02588
R14643 mimbot1.n151 mimbot1.n55 0.02588
R14644 mimbot1.n151 mimbot1.n111 0.02588
R14645 mimbot1.n151 mimbot1.n58 0.02588
R14646 mimbot1.n151 mimbot1.n88 0.02588
R14647 mimbot1.n151 mimbot1.n61 0.02588
R14648 mimbot1.n151 mimbot1.n64 0.02588
R14649 mimbot1.n62 mimbot1 0.024
R14650 mimbot1.n606 mimbot1 0.024
R14651 mimbot1 mimbot1.n585 0.024
R14652 mimbot1.n137 mimbot1 0.024
R14653 mimbot1.n6 mimbot1.n5 0.023003
R14654 mimbot1.n371 mimbot1 0.0224565
R14655 mimbot1.n351 mimbot1 0.0224565
R14656 mimbot1.n41 mimbot1 0.0224565
R14657 mimbot1.n216 mimbot1 0.0224565
R14658 mimbot1.n283 mimbot1 0.0224565
R14659 mimbot1.n251 mimbot1 0.0224565
R14660 mimbot1.n273 mimbot1 0.0224565
R14661 mimbot1.n262 mimbot1 0.0224565
R14662 mimbot1.n326 mimbot1 0.0224565
R14663 mimbot1.n254 mimbot1 0.0224565
R14664 mimbot1.n346 mimbot1 0.0224565
R14665 mimbot1.n376 mimbot1 0.0224565
R14666 mimbot1.n396 mimbot1 0.0224565
R14667 mimbot1.n365 mimbot1 0.0224565
R14668 mimbot1.n368 mimbot1 0.0224565
R14669 mimbot1.n415 mimbot1 0.0224565
R14670 mimbot1.n495 mimbot1 0.0224565
R14671 mimbot1.n471 mimbot1 0.0224565
R14672 mimbot1.n685 mimbot1 0.0224565
R14673 mimbot1.n488 mimbot1 0.0224565
R14674 mimbot1.n479 mimbot1 0.0224565
R14675 mimbot1.n538 mimbot1 0.0224565
R14676 mimbot1.n482 mimbot1 0.0224565
R14677 mimbot1.n560 mimbot1 0.0224565
R14678 mimbot1.n549 mimbot1 0.0224565
R14679 mimbot1.n485 mimbot1 0.0224565
R14680 mimbot1.n474 mimbot1 0.0224565
R14681 mimbot1.n526 mimbot1 0.0224565
R14682 mimbot1.n359 mimbot1 0.0224565
R14683 mimbot1.n446 mimbot1 0.0224565
R14684 mimbot1.n363 mimbot1 0.0224565
R14685 mimbot1.n435 mimbot1 0.0224565
R14686 mimbot1.n356 mimbot1 0.0224565
R14687 mimbot1.n456 mimbot1 0.0224565
R14688 mimbot1.n266 mimbot1 0.0224565
R14689 mimbot1.n716 mimbot1 0.0224565
R14690 mimbot1.n50 mimbot1 0.0224565
R14691 mimbot1.n237 mimbot1 0.0224565
R14692 mimbot1.n30 mimbot1 0.0224565
R14693 mimbot1.n162 mimbot1 0.0224565
R14694 mimbot1.n256 mimbot1 0.0224565
R14695 mimbot1.n336 mimbot1 0.0224565
R14696 mimbot1.n47 mimbot1 0.0224565
R14697 mimbot1.n172 mimbot1 0.0224565
R14698 mimbot1.n33 mimbot1 0.0224565
R14699 mimbot1.n183 mimbot1 0.0224565
R14700 mimbot1.n260 mimbot1 0.0224565
R14701 mimbot1.n314 mimbot1 0.0224565
R14702 mimbot1.n44 mimbot1 0.0224565
R14703 mimbot1.n206 mimbot1 0.0224565
R14704 mimbot1.n36 mimbot1 0.0224565
R14705 mimbot1.n195 mimbot1 0.0224565
R14706 mimbot1.n246 mimbot1 0.0224565
R14707 mimbot1.n294 mimbot1 0.0224565
R14708 mimbot1.n466 mimbot1 0.0224565
R14709 mimbot1.n506 mimbot1 0.0224565
R14710 mimbot1.n411 mimbot1.n403 0.0222621
R14711 mimbot1.n279 mimbot1.n269 0.0222621
R14712 mimbot1.n332 mimbot1.n322 0.0222621
R14713 mimbot1.n382 mimbot1.n372 0.0222621
R14714 mimbot1.n402 mimbot1.n392 0.0222621
R14715 mimbot1.n421 mimbot1.n412 0.0222621
R14716 mimbot1.n684 mimbot1.n683 0.0222621
R14717 mimbot1.n544 mimbot1.n534 0.0222621
R14718 mimbot1.n566 mimbot1.n556 0.0222621
R14719 mimbot1.n555 mimbot1.n545 0.0222621
R14720 mimbot1.n533 mimbot1.n532 0.0222621
R14721 mimbot1.n452 mimbot1.n442 0.0222621
R14722 mimbot1.n441 mimbot1.n431 0.0222621
R14723 mimbot1.n463 mimbot1.n462 0.0222621
R14724 mimbot1.n711 mimbot1.n708 0.0222621
R14725 mimbot1.n243 mimbot1.n233 0.0222621
R14726 mimbot1.n168 mimbot1.n158 0.0222621
R14727 mimbot1.n343 mimbot1.n342 0.0222621
R14728 mimbot1.n223 mimbot1.n222 0.0222621
R14729 mimbot1.n190 mimbot1.n189 0.0222621
R14730 mimbot1.n179 mimbot1.n178 0.0222621
R14731 mimbot1.n321 mimbot1.n320 0.0222621
R14732 mimbot1.n212 mimbot1.n202 0.0222621
R14733 mimbot1.n201 mimbot1.n191 0.0222621
R14734 mimbot1.n301 mimbot1.n300 0.0222621
R14735 mimbot1.n290 mimbot1.n289 0.0222621
R14736 mimbot1.n513 mimbot1.n512 0.0222621
R14737 mimbot1.n502 mimbot1.n501 0.0222621
R14738 mimbot1.n63 mimbot1.n62 0.0220558
R14739 mimbot1.n15 mimbot1.n14 0.0218613
R14740 mimbot1.n8 mimbot1.n7 0.0205382
R14741 mimbot1.n19 mimbot1.n18 0.0205382
R14742 mimbot1.n627 mimbot1.n626 0.02024
R14743 mimbot1.n628 mimbot1.n627 0.02024
R14744 mimbot1.n640 mimbot1.n639 0.02024
R14745 mimbot1.n641 mimbot1.n640 0.02024
R14746 mimbot1.n656 mimbot1.n649 0.02024
R14747 mimbot1.n653 mimbot1.n649 0.02024
R14748 mimbot1.n668 mimbot1.n661 0.02024
R14749 mimbot1.n665 mimbot1.n661 0.02024
R14750 mimbot1.n675 mimbot1.n674 0.02024
R14751 mimbot1.n676 mimbot1.n675 0.02024
R14752 mimbot1.n617 mimbot1.n610 0.02024
R14753 mimbot1.n614 mimbot1.n610 0.02024
R14754 mimbot1.n593 mimbot1.n592 0.02024
R14755 mimbot1.n594 mimbot1.n593 0.02024
R14756 mimbot1.n148 mimbot1.n141 0.02024
R14757 mimbot1.n145 mimbot1.n141 0.02024
R14758 mimbot1.n118 mimbot1.n117 0.02024
R14759 mimbot1.n119 mimbot1.n118 0.02024
R14760 mimbot1.n131 mimbot1.n124 0.02024
R14761 mimbot1.n128 mimbot1.n124 0.02024
R14762 mimbot1.n95 mimbot1.n94 0.02024
R14763 mimbot1.n96 mimbot1.n95 0.02024
R14764 mimbot1.n108 mimbot1.n101 0.02024
R14765 mimbot1.n105 mimbot1.n101 0.02024
R14766 mimbot1.n71 mimbot1.n70 0.02024
R14767 mimbot1.n72 mimbot1.n71 0.02024
R14768 mimbot1.n85 mimbot1.n77 0.02024
R14769 mimbot1.n82 mimbot1.n77 0.02024
R14770 mimbot1.n522 mimbot1.n521 0.0200244
R14771 mimbot1.n391 mimbot1.n390 0.0200244
R14772 mimbot1.n310 mimbot1.n309 0.0200244
R14773 mimbot1.n232 mimbot1.n231 0.0200244
R14774 mimbot1.n86 mimbot1.n76 0.0200242
R14775 mimbot1.n68 mimbot1.n67 0.0200242
R14776 mimbot1.n109 mimbot1.n100 0.0200242
R14777 mimbot1.n92 mimbot1.n91 0.0200242
R14778 mimbot1.n132 mimbot1.n123 0.0200242
R14779 mimbot1.n115 mimbot1.n114 0.0200242
R14780 mimbot1.n149 mimbot1.n140 0.0200242
R14781 mimbot1.n590 mimbot1.n589 0.0200242
R14782 mimbot1.n720 mimbot1.n157 0.0200242
R14783 mimbot1.n618 mimbot1.n609 0.0200242
R14784 mimbot1.n624 mimbot1.n623 0.0200242
R14785 mimbot1.n637 mimbot1.n636 0.0200242
R14786 mimbot1.n657 mimbot1.n648 0.0200242
R14787 mimbot1.n669 mimbot1.n660 0.0200242
R14788 mimbot1.n672 mimbot1.n671 0.0200242
R14789 mimbot1.n575 mimbot1.n574 0.0200242
R14790 mimbot1.n430 mimbot1.n422 0.0200242
R14791 mimbot1.n700 mimbot1.n699 0.0200242
R14792 mimbot1.n695 mimbot1.t38 0.01977
R14793 mimbot1.n696 mimbot1.t38 0.01977
R14794 mimbot1.n695 mimbot1.t22 0.01977
R14795 mimbot1.n696 mimbot1.t22 0.01977
R14796 mimbot1.n681 mimbot1.t29 0.01977
R14797 mimbot1.n682 mimbot1.t29 0.01977
R14798 mimbot1.t6 mimbot1.n681 0.01977
R14799 mimbot1.n682 mimbot1.t6 0.01977
R14800 mimbot1.n681 mimbot1.t34 0.01977
R14801 mimbot1.n682 mimbot1.t34 0.01977
R14802 mimbot1.n692 mimbot1.t36 0.01977
R14803 mimbot1.n693 mimbot1.t36 0.01977
R14804 mimbot1.n681 mimbot1.t3 0.01977
R14805 mimbot1.n682 mimbot1.t3 0.01977
R14806 mimbot1.n692 mimbot1.t23 0.01977
R14807 mimbot1.n693 mimbot1.t23 0.01977
R14808 mimbot1.t13 mimbot1.n692 0.01977
R14809 mimbot1.n693 mimbot1.t13 0.01977
R14810 mimbot1.n681 mimbot1.t20 0.01977
R14811 mimbot1.n682 mimbot1.t20 0.01977
R14812 mimbot1.n692 mimbot1.t39 0.01977
R14813 mimbot1.n693 mimbot1.t39 0.01977
R14814 mimbot1.n692 mimbot1.t28 0.01977
R14815 mimbot1.n693 mimbot1.t28 0.01977
R14816 mimbot1.n695 mimbot1.t14 0.01977
R14817 mimbot1.n696 mimbot1.t14 0.01977
R14818 mimbot1.n718 mimbot1.t7 0.01977
R14819 mimbot1.n719 mimbot1.t7 0.01977
R14820 mimbot1.t17 mimbot1.n718 0.01977
R14821 mimbot1.n719 mimbot1.t17 0.01977
R14822 mimbot1.t25 mimbot1.n695 0.01977
R14823 mimbot1.n696 mimbot1.t25 0.01977
R14824 mimbot1.n718 mimbot1.t31 0.01977
R14825 mimbot1.n719 mimbot1.t31 0.01977
R14826 mimbot1.n718 mimbot1.t2 0.01977
R14827 mimbot1.n719 mimbot1.t2 0.01977
R14828 mimbot1.n695 mimbot1.t10 0.01977
R14829 mimbot1.n696 mimbot1.t10 0.01977
R14830 mimbot1.n718 mimbot1.t16 0.01977
R14831 mimbot1.n719 mimbot1.t16 0.01977
R14832 mimbot1.n718 mimbot1.t37 0.01977
R14833 mimbot1.n719 mimbot1.t37 0.01977
R14834 mimbot1.n718 mimbot1.t27 0.01977
R14835 mimbot1.n719 mimbot1.t27 0.01977
R14836 mimbot1.n695 mimbot1.t33 0.01977
R14837 mimbot1.n696 mimbot1.t33 0.01977
R14838 mimbot1.n695 mimbot1.t5 0.01977
R14839 mimbot1.n696 mimbot1.t5 0.01977
R14840 mimbot1.n692 mimbot1.t19 0.01977
R14841 mimbot1.n693 mimbot1.t19 0.01977
R14842 mimbot1.n692 mimbot1.t8 0.01977
R14843 mimbot1.n693 mimbot1.t8 0.01977
R14844 mimbot1.n681 mimbot1.t15 0.01977
R14845 mimbot1.n682 mimbot1.t15 0.01977
R14846 mimbot1.n681 mimbot1.t26 0.01977
R14847 mimbot1.n682 mimbot1.t26 0.01977
R14848 mimbot1.n681 mimbot1.t41 0.01977
R14849 mimbot1.n682 mimbot1.t41 0.01977
R14850 mimbot1.n692 mimbot1.t32 0.01977
R14851 mimbot1.n693 mimbot1.t32 0.01977
R14852 mimbot1.n695 mimbot1.t18 0.01977
R14853 mimbot1.n696 mimbot1.t18 0.01977
R14854 mimbot1.n718 mimbot1.t12 0.01977
R14855 mimbot1.n719 mimbot1.t12 0.01977
R14856 mimbot1.n723 mimbot1.t4 0.01977
R14857 mimbot1.n151 mimbot1.t4 0.01977
R14858 mimbot1.n723 mimbot1.t30 0.01977
R14859 mimbot1.n151 mimbot1.t30 0.01977
R14860 mimbot1.n723 mimbot1.t21 0.01977
R14861 mimbot1.n151 mimbot1.t21 0.01977
R14862 mimbot1.n723 mimbot1.t9 0.01977
R14863 mimbot1.n151 mimbot1.t9 0.01977
R14864 mimbot1.n723 mimbot1.t35 0.01977
R14865 mimbot1.n151 mimbot1.t35 0.01977
R14866 mimbot1.n723 mimbot1.t24 0.01977
R14867 mimbot1.n151 mimbot1.t24 0.01977
R14868 mimbot1.n723 mimbot1.t11 0.01977
R14869 mimbot1.n151 mimbot1.t11 0.01977
R14870 mimbot1.n723 mimbot1.t40 0.01977
R14871 mimbot1.t40 mimbot1.n151 0.01977
R14872 mimbot1.n80 mimbot1 0.0195238
R14873 mimbot1.n74 mimbot1 0.0195238
R14874 mimbot1.n103 mimbot1 0.0195238
R14875 mimbot1.n98 mimbot1 0.0195238
R14876 mimbot1.n126 mimbot1 0.0195238
R14877 mimbot1.n121 mimbot1 0.0195238
R14878 mimbot1.n143 mimbot1 0.0195238
R14879 mimbot1.n596 mimbot1 0.0195238
R14880 mimbot1 mimbot1.n27 0.0195238
R14881 mimbot1 mimbot1.n605 0.0195238
R14882 mimbot1.n612 mimbot1 0.0195238
R14883 mimbot1.n630 mimbot1 0.0195238
R14884 mimbot1.n643 mimbot1 0.0195238
R14885 mimbot1.n651 mimbot1 0.0195238
R14886 mimbot1.n663 mimbot1 0.0195238
R14887 mimbot1.n678 mimbot1 0.0195238
R14888 mimbot1 mimbot1.n570 0.0195238
R14889 mimbot1 mimbot1.n424 0.0195238
R14890 mimbot1 mimbot1.n702 0.0195238
R14891 mimbot1.n586 mimbot1 0.0195238
R14892 mimbot1.n585 mimbot1.n584 0.0195238
R14893 mimbot1 mimbot1.n518 0.0195238
R14894 mimbot1 mimbot1.n387 0.0195238
R14895 mimbot1 mimbot1.n306 0.0195238
R14896 mimbot1 mimbot1.n228 0.0195238
R14897 mimbot1.n138 mimbot1.n137 0.0195238
R14898 mimbot1.n215 mimbot1.n214 0.0188601
R14899 mimbot1.n375 mimbot1.n373 0.0188601
R14900 mimbot1.n413 mimbot1.n369 0.0188601
R14901 mimbot1.n395 mimbot1.n393 0.0188601
R14902 mimbot1.n537 mimbot1.n535 0.0188601
R14903 mimbot1.n559 mimbot1.n557 0.0188601
R14904 mimbot1.n525 mimbot1.n524 0.0188601
R14905 mimbot1.n491 mimbot1.n490 0.0188601
R14906 mimbot1.n445 mimbot1.n443 0.0188601
R14907 mimbot1.n434 mimbot1.n432 0.0188601
R14908 mimbot1.n548 mimbot1.n546 0.0188601
R14909 mimbot1.n455 mimbot1.n454 0.0188601
R14910 mimbot1.n709 mimbot1.n707 0.0188601
R14911 mimbot1.n236 mimbot1.n234 0.0188601
R14912 mimbot1.n161 mimbot1.n159 0.0188601
R14913 mimbot1.n325 mimbot1.n323 0.0188601
R14914 mimbot1.n335 mimbot1.n334 0.0188601
R14915 mimbot1.n171 mimbot1.n170 0.0188601
R14916 mimbot1.n182 mimbot1.n181 0.0188601
R14917 mimbot1.n272 mimbot1.n270 0.0188601
R14918 mimbot1.n313 mimbot1.n312 0.0188601
R14919 mimbot1.n205 mimbot1.n203 0.0188601
R14920 mimbot1.n194 mimbot1.n192 0.0188601
R14921 mimbot1.n282 mimbot1.n281 0.0188601
R14922 mimbot1.n293 mimbot1.n292 0.0188601
R14923 mimbot1.n405 mimbot1.n404 0.0188601
R14924 mimbot1.n494 mimbot1.n493 0.0188601
R14925 mimbot1.n505 mimbot1.n504 0.0188601
R14926 mimbot1.n221 mimbot1.n218 0.01836
R14927 mimbot1.n380 mimbot1.n374 0.01836
R14928 mimbot1.n419 mimbot1.n414 0.01836
R14929 mimbot1.n400 mimbot1.n394 0.01836
R14930 mimbot1.n542 mimbot1.n536 0.01836
R14931 mimbot1.n564 mimbot1.n558 0.01836
R14932 mimbot1.n531 mimbot1.n528 0.01836
R14933 mimbot1.n688 mimbot1.n687 0.01836
R14934 mimbot1.n450 mimbot1.n444 0.01836
R14935 mimbot1.n439 mimbot1.n433 0.01836
R14936 mimbot1.n553 mimbot1.n547 0.01836
R14937 mimbot1.n461 mimbot1.n458 0.01836
R14938 mimbot1.n713 mimbot1.n706 0.01836
R14939 mimbot1.n241 mimbot1.n235 0.01836
R14940 mimbot1.n166 mimbot1.n160 0.01836
R14941 mimbot1.n330 mimbot1.n324 0.01836
R14942 mimbot1.n341 mimbot1.n338 0.01836
R14943 mimbot1.n177 mimbot1.n174 0.01836
R14944 mimbot1.n188 mimbot1.n185 0.01836
R14945 mimbot1.n277 mimbot1.n271 0.01836
R14946 mimbot1.n319 mimbot1.n316 0.01836
R14947 mimbot1.n210 mimbot1.n204 0.01836
R14948 mimbot1.n199 mimbot1.n193 0.01836
R14949 mimbot1.n288 mimbot1.n285 0.01836
R14950 mimbot1.n299 mimbot1.n296 0.01836
R14951 mimbot1.n409 mimbot1.n370 0.01836
R14952 mimbot1.n500 mimbot1.n497 0.01836
R14953 mimbot1.n511 mimbot1.n508 0.01836
R14954 mimbot1.n721 mimbot1.n152 0.01648
R14955 mimbot1.n572 mimbot1.n567 0.01648
R14956 mimbot1.n429 mimbot1.n423 0.01648
R14957 mimbot1.n705 mimbot1.n701 0.01648
R14958 mimbot1.n516 mimbot1.n514 0.01648
R14959 mimbot1.n385 mimbot1.n383 0.01648
R14960 mimbot1.n304 mimbot1.n302 0.01648
R14961 mimbot1.n226 mimbot1.n224 0.01648
R14962 mimbot1.n215 mimbot1.n42 0.0157702
R14963 mimbot1.n696 mimbot1.n279 0.0157702
R14964 mimbot1.n696 mimbot1.n332 0.0157702
R14965 mimbot1.n375 mimbot1.n345 0.0157702
R14966 mimbot1.n693 mimbot1.n382 0.0157702
R14967 mimbot1.n693 mimbot1.n402 0.0157702
R14968 mimbot1.n694 mimbot1.n369 0.0157702
R14969 mimbot1.n395 mimbot1.n361 0.0157702
R14970 mimbot1.n683 mimbot1.n682 0.0157702
R14971 mimbot1.n537 mimbot1.n478 0.0157702
R14972 mimbot1.n682 mimbot1.n544 0.0157702
R14973 mimbot1.n559 mimbot1.n481 0.0157702
R14974 mimbot1.n682 mimbot1.n555 0.0157702
R14975 mimbot1.n682 mimbot1.n566 0.0157702
R14976 mimbot1.n682 mimbot1.n533 0.0157702
R14977 mimbot1.n525 mimbot1.n473 0.0157702
R14978 mimbot1.n490 mimbot1.n477 0.0157702
R14979 mimbot1.n445 mimbot1.n352 0.0157702
R14980 mimbot1.n434 mimbot1.n362 0.0157702
R14981 mimbot1.n693 mimbot1.n441 0.0157702
R14982 mimbot1.n693 mimbot1.n452 0.0157702
R14983 mimbot1.n548 mimbot1.n480 0.0157702
R14984 mimbot1.n693 mimbot1.n463 0.0157702
R14985 mimbot1.n455 mimbot1.n357 0.0157702
R14986 mimbot1.n711 mimbot1.n696 0.0157702
R14987 mimbot1.n707 mimbot1.n265 0.0157702
R14988 mimbot1.n236 mimbot1.n29 0.0157702
R14989 mimbot1.n161 mimbot1.n48 0.0157702
R14990 mimbot1.n719 mimbot1.n168 0.0157702
R14991 mimbot1.n719 mimbot1.n243 0.0157702
R14992 mimbot1.n325 mimbot1.n253 0.0157702
R14993 mimbot1.n696 mimbot1.n343 0.0157702
R14994 mimbot1.n335 mimbot1.n257 0.0157702
R14995 mimbot1.n719 mimbot1.n223 0.0157702
R14996 mimbot1.n171 mimbot1.n32 0.0157702
R14997 mimbot1.n182 mimbot1.n45 0.0157702
R14998 mimbot1.n719 mimbot1.n190 0.0157702
R14999 mimbot1.n719 mimbot1.n179 0.0157702
R15000 mimbot1.n272 mimbot1.n263 0.0157702
R15001 mimbot1.n696 mimbot1.n321 0.0157702
R15002 mimbot1.n313 mimbot1.n259 0.0157702
R15003 mimbot1.n205 mimbot1.n35 0.0157702
R15004 mimbot1.n194 mimbot1.n40 0.0157702
R15005 mimbot1.n719 mimbot1.n201 0.0157702
R15006 mimbot1.n719 mimbot1.n212 0.0157702
R15007 mimbot1.n282 mimbot1.n250 0.0157702
R15008 mimbot1.n293 mimbot1.n245 0.0157702
R15009 mimbot1.n696 mimbot1.n301 0.0157702
R15010 mimbot1.n696 mimbot1.n290 0.0157702
R15011 mimbot1.n405 mimbot1.n350 0.0157702
R15012 mimbot1.n693 mimbot1.n411 0.0157702
R15013 mimbot1.n693 mimbot1.n421 0.0157702
R15014 mimbot1.n494 mimbot1.n470 0.0157702
R15015 mimbot1.n505 mimbot1.n465 0.0157702
R15016 mimbot1.n682 mimbot1.n513 0.0157702
R15017 mimbot1.n682 mimbot1.n502 0.0157702
R15018 mimbot1.n18 mimbot1.n17 0.0143192
R15019 mimbot1 mimbot1.n724 0.0138019
R15020 mimbot1 mimbot1.n725 0.0128348
R15021 mimbot1 mimbot1.n403 0.01225
R15022 mimbot1.n408 mimbot1 0.01225
R15023 mimbot1.n408 mimbot1 0.01225
R15024 mimbot1.n222 mimbot1 0.01225
R15025 mimbot1.n220 mimbot1 0.01225
R15026 mimbot1.n220 mimbot1 0.01225
R15027 mimbot1.n289 mimbot1 0.01225
R15028 mimbot1.n287 mimbot1 0.01225
R15029 mimbot1.n287 mimbot1 0.01225
R15030 mimbot1 mimbot1.n269 0.01225
R15031 mimbot1.n276 mimbot1 0.01225
R15032 mimbot1.n276 mimbot1 0.01225
R15033 mimbot1 mimbot1.n322 0.01225
R15034 mimbot1.n329 mimbot1 0.01225
R15035 mimbot1.n329 mimbot1 0.01225
R15036 mimbot1 mimbot1.n372 0.01225
R15037 mimbot1.n379 mimbot1 0.01225
R15038 mimbot1.n379 mimbot1 0.01225
R15039 mimbot1 mimbot1.n392 0.01225
R15040 mimbot1.n399 mimbot1 0.01225
R15041 mimbot1.n399 mimbot1 0.01225
R15042 mimbot1 mimbot1.n412 0.01225
R15043 mimbot1.n418 mimbot1 0.01225
R15044 mimbot1.n418 mimbot1 0.01225
R15045 mimbot1.n501 mimbot1 0.01225
R15046 mimbot1.n499 mimbot1 0.01225
R15047 mimbot1.n499 mimbot1 0.01225
R15048 mimbot1.n684 mimbot1 0.01225
R15049 mimbot1.n689 mimbot1 0.01225
R15050 mimbot1 mimbot1.n689 0.01225
R15051 mimbot1 mimbot1.n534 0.01225
R15052 mimbot1.n541 mimbot1 0.01225
R15053 mimbot1.n541 mimbot1 0.01225
R15054 mimbot1 mimbot1.n556 0.01225
R15055 mimbot1.n563 mimbot1 0.01225
R15056 mimbot1.n563 mimbot1 0.01225
R15057 mimbot1 mimbot1.n545 0.01225
R15058 mimbot1.n552 mimbot1 0.01225
R15059 mimbot1.n552 mimbot1 0.01225
R15060 mimbot1.n532 mimbot1 0.01225
R15061 mimbot1.n530 mimbot1 0.01225
R15062 mimbot1.n530 mimbot1 0.01225
R15063 mimbot1 mimbot1.n442 0.01225
R15064 mimbot1.n449 mimbot1 0.01225
R15065 mimbot1.n449 mimbot1 0.01225
R15066 mimbot1 mimbot1.n431 0.01225
R15067 mimbot1.n438 mimbot1 0.01225
R15068 mimbot1.n438 mimbot1 0.01225
R15069 mimbot1.n462 mimbot1 0.01225
R15070 mimbot1.n460 mimbot1 0.01225
R15071 mimbot1.n460 mimbot1 0.01225
R15072 mimbot1 mimbot1.n708 0.01225
R15073 mimbot1 mimbot1.n714 0.01225
R15074 mimbot1.n714 mimbot1 0.01225
R15075 mimbot1 mimbot1.n233 0.01225
R15076 mimbot1.n240 mimbot1 0.01225
R15077 mimbot1.n240 mimbot1 0.01225
R15078 mimbot1 mimbot1.n158 0.01225
R15079 mimbot1.n165 mimbot1 0.01225
R15080 mimbot1.n165 mimbot1 0.01225
R15081 mimbot1.n342 mimbot1 0.01225
R15082 mimbot1.n340 mimbot1 0.01225
R15083 mimbot1.n340 mimbot1 0.01225
R15084 mimbot1.n178 mimbot1 0.01225
R15085 mimbot1.n176 mimbot1 0.01225
R15086 mimbot1.n176 mimbot1 0.01225
R15087 mimbot1.n189 mimbot1 0.01225
R15088 mimbot1.n187 mimbot1 0.01225
R15089 mimbot1.n187 mimbot1 0.01225
R15090 mimbot1.n320 mimbot1 0.01225
R15091 mimbot1.n318 mimbot1 0.01225
R15092 mimbot1.n318 mimbot1 0.01225
R15093 mimbot1 mimbot1.n202 0.01225
R15094 mimbot1.n209 mimbot1 0.01225
R15095 mimbot1.n209 mimbot1 0.01225
R15096 mimbot1 mimbot1.n191 0.01225
R15097 mimbot1.n198 mimbot1 0.01225
R15098 mimbot1.n198 mimbot1 0.01225
R15099 mimbot1.n300 mimbot1 0.01225
R15100 mimbot1.n298 mimbot1 0.01225
R15101 mimbot1.n298 mimbot1 0.01225
R15102 mimbot1.n512 mimbot1 0.01225
R15103 mimbot1.n510 mimbot1 0.01225
R15104 mimbot1.n510 mimbot1 0.01225
R15105 mimbot1.n607 mimbot1.n603 0.0116498
R15106 mimbot1.n3 mimbot1.n2 0.0105709
R15107 mimbot1 mimbot1.n405 0.0105121
R15108 mimbot1 mimbot1.n215 0.0105121
R15109 mimbot1 mimbot1.n282 0.0105121
R15110 mimbot1 mimbot1.n272 0.0105121
R15111 mimbot1 mimbot1.n325 0.0105121
R15112 mimbot1 mimbot1.n375 0.0105121
R15113 mimbot1 mimbot1.n395 0.0105121
R15114 mimbot1 mimbot1.n369 0.0105121
R15115 mimbot1 mimbot1.n494 0.0105121
R15116 mimbot1.n490 mimbot1 0.0105121
R15117 mimbot1 mimbot1.n537 0.0105121
R15118 mimbot1 mimbot1.n559 0.0105121
R15119 mimbot1 mimbot1.n548 0.0105121
R15120 mimbot1 mimbot1.n525 0.0105121
R15121 mimbot1 mimbot1.n445 0.0105121
R15122 mimbot1 mimbot1.n434 0.0105121
R15123 mimbot1 mimbot1.n455 0.0105121
R15124 mimbot1 mimbot1.n707 0.0105121
R15125 mimbot1 mimbot1.n236 0.0105121
R15126 mimbot1 mimbot1.n161 0.0105121
R15127 mimbot1 mimbot1.n335 0.0105121
R15128 mimbot1 mimbot1.n171 0.0105121
R15129 mimbot1 mimbot1.n182 0.0105121
R15130 mimbot1 mimbot1.n313 0.0105121
R15131 mimbot1 mimbot1.n205 0.0105121
R15132 mimbot1 mimbot1.n194 0.0105121
R15133 mimbot1 mimbot1.n293 0.0105121
R15134 mimbot1 mimbot1.n505 0.0105121
R15135 mimbot1.n214 mimbot1.n213 0.01037
R15136 mimbot1.n221 mimbot1.n213 0.01037
R15137 mimbot1.n381 mimbot1.n373 0.01037
R15138 mimbot1.n381 mimbot1.n380 0.01037
R15139 mimbot1.n420 mimbot1.n413 0.01037
R15140 mimbot1.n420 mimbot1.n419 0.01037
R15141 mimbot1.n401 mimbot1.n393 0.01037
R15142 mimbot1.n401 mimbot1.n400 0.01037
R15143 mimbot1.n543 mimbot1.n535 0.01037
R15144 mimbot1.n543 mimbot1.n542 0.01037
R15145 mimbot1.n565 mimbot1.n557 0.01037
R15146 mimbot1.n565 mimbot1.n564 0.01037
R15147 mimbot1.n524 mimbot1.n523 0.01037
R15148 mimbot1.n531 mimbot1.n523 0.01037
R15149 mimbot1.n491 mimbot1.n489 0.01037
R15150 mimbot1.n688 mimbot1.n489 0.01037
R15151 mimbot1.n451 mimbot1.n443 0.01037
R15152 mimbot1.n451 mimbot1.n450 0.01037
R15153 mimbot1.n440 mimbot1.n432 0.01037
R15154 mimbot1.n440 mimbot1.n439 0.01037
R15155 mimbot1.n554 mimbot1.n546 0.01037
R15156 mimbot1.n554 mimbot1.n553 0.01037
R15157 mimbot1.n454 mimbot1.n453 0.01037
R15158 mimbot1.n461 mimbot1.n453 0.01037
R15159 mimbot1.n712 mimbot1.n709 0.01037
R15160 mimbot1.n713 mimbot1.n712 0.01037
R15161 mimbot1.n242 mimbot1.n234 0.01037
R15162 mimbot1.n242 mimbot1.n241 0.01037
R15163 mimbot1.n167 mimbot1.n159 0.01037
R15164 mimbot1.n167 mimbot1.n166 0.01037
R15165 mimbot1.n331 mimbot1.n323 0.01037
R15166 mimbot1.n331 mimbot1.n330 0.01037
R15167 mimbot1.n334 mimbot1.n333 0.01037
R15168 mimbot1.n341 mimbot1.n333 0.01037
R15169 mimbot1.n170 mimbot1.n169 0.01037
R15170 mimbot1.n177 mimbot1.n169 0.01037
R15171 mimbot1.n181 mimbot1.n180 0.01037
R15172 mimbot1.n188 mimbot1.n180 0.01037
R15173 mimbot1.n278 mimbot1.n270 0.01037
R15174 mimbot1.n278 mimbot1.n277 0.01037
R15175 mimbot1.n312 mimbot1.n311 0.01037
R15176 mimbot1.n319 mimbot1.n311 0.01037
R15177 mimbot1.n211 mimbot1.n203 0.01037
R15178 mimbot1.n211 mimbot1.n210 0.01037
R15179 mimbot1.n200 mimbot1.n192 0.01037
R15180 mimbot1.n200 mimbot1.n199 0.01037
R15181 mimbot1.n281 mimbot1.n280 0.01037
R15182 mimbot1.n288 mimbot1.n280 0.01037
R15183 mimbot1.n292 mimbot1.n291 0.01037
R15184 mimbot1.n299 mimbot1.n291 0.01037
R15185 mimbot1.n410 mimbot1.n404 0.01037
R15186 mimbot1.n410 mimbot1.n409 0.01037
R15187 mimbot1.n493 mimbot1.n492 0.01037
R15188 mimbot1.n500 mimbot1.n492 0.01037
R15189 mimbot1.n504 mimbot1.n503 0.01037
R15190 mimbot1.n511 mimbot1.n503 0.01037
R15191 mimbot1 mimbot1.n406 0.0100119
R15192 mimbot1 mimbot1.n407 0.0100119
R15193 mimbot1 mimbot1.n219 0.0100119
R15194 mimbot1.n217 mimbot1 0.0100119
R15195 mimbot1.n284 mimbot1 0.0100119
R15196 mimbot1 mimbot1.n286 0.0100119
R15197 mimbot1 mimbot1.n274 0.0100119
R15198 mimbot1 mimbot1.n275 0.0100119
R15199 mimbot1 mimbot1.n327 0.0100119
R15200 mimbot1 mimbot1.n328 0.0100119
R15201 mimbot1 mimbot1.n378 0.0100119
R15202 mimbot1 mimbot1.n377 0.0100119
R15203 mimbot1 mimbot1.n397 0.0100119
R15204 mimbot1 mimbot1.n398 0.0100119
R15205 mimbot1 mimbot1.n417 0.0100119
R15206 mimbot1 mimbot1.n416 0.0100119
R15207 mimbot1.n496 mimbot1 0.0100119
R15208 mimbot1 mimbot1.n498 0.0100119
R15209 mimbot1.n686 mimbot1 0.0100119
R15210 mimbot1.n690 mimbot1 0.0100119
R15211 mimbot1 mimbot1.n540 0.0100119
R15212 mimbot1 mimbot1.n539 0.0100119
R15213 mimbot1 mimbot1.n562 0.0100119
R15214 mimbot1 mimbot1.n561 0.0100119
R15215 mimbot1 mimbot1.n550 0.0100119
R15216 mimbot1 mimbot1.n551 0.0100119
R15217 mimbot1 mimbot1.n529 0.0100119
R15218 mimbot1.n527 mimbot1 0.0100119
R15219 mimbot1 mimbot1.n448 0.0100119
R15220 mimbot1 mimbot1.n447 0.0100119
R15221 mimbot1 mimbot1.n437 0.0100119
R15222 mimbot1 mimbot1.n436 0.0100119
R15223 mimbot1 mimbot1.n459 0.0100119
R15224 mimbot1.n457 mimbot1 0.0100119
R15225 mimbot1 mimbot1.n710 0.0100119
R15226 mimbot1.n715 mimbot1 0.0100119
R15227 mimbot1 mimbot1.n239 0.0100119
R15228 mimbot1 mimbot1.n238 0.0100119
R15229 mimbot1 mimbot1.n164 0.0100119
R15230 mimbot1 mimbot1.n163 0.0100119
R15231 mimbot1 mimbot1.n339 0.0100119
R15232 mimbot1.n337 mimbot1 0.0100119
R15233 mimbot1 mimbot1.n175 0.0100119
R15234 mimbot1.n173 mimbot1 0.0100119
R15235 mimbot1 mimbot1.n186 0.0100119
R15236 mimbot1.n184 mimbot1 0.0100119
R15237 mimbot1 mimbot1.n317 0.0100119
R15238 mimbot1.n315 mimbot1 0.0100119
R15239 mimbot1 mimbot1.n208 0.0100119
R15240 mimbot1 mimbot1.n207 0.0100119
R15241 mimbot1 mimbot1.n197 0.0100119
R15242 mimbot1 mimbot1.n196 0.0100119
R15243 mimbot1 mimbot1.n297 0.0100119
R15244 mimbot1.n295 mimbot1 0.0100119
R15245 mimbot1 mimbot1.n509 0.0100119
R15246 mimbot1.n507 mimbot1 0.0100119
R15247 mimbot1.n16 mimbot1.n15 0.00991089
R15248 mimbot1.n522 mimbot1.n514 0.00946062
R15249 mimbot1.n391 mimbot1.n383 0.00946062
R15250 mimbot1.n310 mimbot1.n302 0.00946062
R15251 mimbot1.n232 mimbot1.n224 0.00946062
R15252 mimbot1.n721 mimbot1.n720 0.00946026
R15253 mimbot1.n575 mimbot1.n567 0.00946026
R15254 mimbot1.n430 mimbot1.n429 0.00946026
R15255 mimbot1.n701 mimbot1.n700 0.00946026
R15256 mimbot1.n567 mimbot1.n475 0.00896
R15257 mimbot1.n429 mimbot1.n355 0.00896
R15258 mimbot1.n701 mimbot1.n267 0.00896
R15259 mimbot1.n587 mimbot1.n581 0.00896
R15260 mimbot1.n514 mimbot1.n469 0.00896
R15261 mimbot1.n383 mimbot1.n349 0.00896
R15262 mimbot1.n302 mimbot1.n249 0.00896
R15263 mimbot1.n224 mimbot1.n37 0.00896
R15264 mimbot1.n722 mimbot1.n721 0.00896
R15265 mimbot1.n21 mimbot1.n20 0.0082163
R15266 mimbot1.n22 mimbot1.n21 0.00815306
R15267 mimbot1.n84 mimbot1.n76 0.00610795
R15268 mimbot1.n84 mimbot1 0.00610795
R15269 mimbot1 mimbot1.n83 0.00610795
R15270 mimbot1.n83 mimbot1 0.00610795
R15271 mimbot1.n69 mimbot1.n68 0.00610795
R15272 mimbot1.n69 mimbot1 0.00610795
R15273 mimbot1.n73 mimbot1 0.00610795
R15274 mimbot1 mimbot1.n73 0.00610795
R15275 mimbot1.n107 mimbot1.n100 0.00610795
R15276 mimbot1.n107 mimbot1 0.00610795
R15277 mimbot1 mimbot1.n106 0.00610795
R15278 mimbot1.n106 mimbot1 0.00610795
R15279 mimbot1.n93 mimbot1.n92 0.00610795
R15280 mimbot1.n93 mimbot1 0.00610795
R15281 mimbot1.n97 mimbot1 0.00610795
R15282 mimbot1 mimbot1.n97 0.00610795
R15283 mimbot1.n130 mimbot1.n123 0.00610795
R15284 mimbot1.n130 mimbot1 0.00610795
R15285 mimbot1 mimbot1.n129 0.00610795
R15286 mimbot1.n129 mimbot1 0.00610795
R15287 mimbot1.n116 mimbot1.n115 0.00610795
R15288 mimbot1.n116 mimbot1 0.00610795
R15289 mimbot1.n120 mimbot1 0.00610795
R15290 mimbot1 mimbot1.n120 0.00610795
R15291 mimbot1.n147 mimbot1.n140 0.00610795
R15292 mimbot1.n147 mimbot1 0.00610795
R15293 mimbot1 mimbot1.n146 0.00610795
R15294 mimbot1.n146 mimbot1 0.00610795
R15295 mimbot1.n591 mimbot1.n590 0.00610795
R15296 mimbot1.n591 mimbot1 0.00610795
R15297 mimbot1.n595 mimbot1 0.00610795
R15298 mimbot1 mimbot1.n595 0.00610795
R15299 mimbot1.n157 mimbot1.n156 0.00610795
R15300 mimbot1.n156 mimbot1 0.00610795
R15301 mimbot1 mimbot1.n155 0.00610795
R15302 mimbot1.n155 mimbot1 0.00610795
R15303 mimbot1.n616 mimbot1.n609 0.00610795
R15304 mimbot1.n616 mimbot1 0.00610795
R15305 mimbot1 mimbot1.n615 0.00610795
R15306 mimbot1.n615 mimbot1 0.00610795
R15307 mimbot1.n625 mimbot1.n624 0.00610795
R15308 mimbot1.n625 mimbot1 0.00610795
R15309 mimbot1.n629 mimbot1 0.00610795
R15310 mimbot1 mimbot1.n629 0.00610795
R15311 mimbot1.n638 mimbot1.n637 0.00610795
R15312 mimbot1.n638 mimbot1 0.00610795
R15313 mimbot1.n642 mimbot1 0.00610795
R15314 mimbot1 mimbot1.n642 0.00610795
R15315 mimbot1.n655 mimbot1.n648 0.00610795
R15316 mimbot1.n655 mimbot1 0.00610795
R15317 mimbot1 mimbot1.n654 0.00610795
R15318 mimbot1.n654 mimbot1 0.00610795
R15319 mimbot1.n667 mimbot1.n660 0.00610795
R15320 mimbot1.n667 mimbot1 0.00610795
R15321 mimbot1 mimbot1.n666 0.00610795
R15322 mimbot1.n666 mimbot1 0.00610795
R15323 mimbot1.n673 mimbot1.n672 0.00610795
R15324 mimbot1.n673 mimbot1 0.00610795
R15325 mimbot1.n677 mimbot1 0.00610795
R15326 mimbot1 mimbot1.n677 0.00610795
R15327 mimbot1.n574 mimbot1.n573 0.00610795
R15328 mimbot1.n573 mimbot1 0.00610795
R15329 mimbot1.n571 mimbot1 0.00610795
R15330 mimbot1.n571 mimbot1 0.00610795
R15331 mimbot1.n427 mimbot1.n422 0.00610795
R15332 mimbot1.n427 mimbot1 0.00610795
R15333 mimbot1 mimbot1.n425 0.00610795
R15334 mimbot1.n425 mimbot1 0.00610795
R15335 mimbot1.n699 mimbot1.n698 0.00610795
R15336 mimbot1 mimbot1.n698 0.00610795
R15337 mimbot1.n704 mimbot1 0.00610795
R15338 mimbot1.n704 mimbot1 0.00610795
R15339 mimbot1.n521 mimbot1.n520 0.00610795
R15340 mimbot1.n520 mimbot1 0.00610795
R15341 mimbot1 mimbot1.n519 0.00610795
R15342 mimbot1.n519 mimbot1 0.00610795
R15343 mimbot1.n390 mimbot1.n389 0.00610795
R15344 mimbot1.n389 mimbot1 0.00610795
R15345 mimbot1 mimbot1.n388 0.00610795
R15346 mimbot1.n388 mimbot1 0.00610795
R15347 mimbot1.n309 mimbot1.n308 0.00610795
R15348 mimbot1.n308 mimbot1 0.00610795
R15349 mimbot1 mimbot1.n307 0.00610795
R15350 mimbot1.n307 mimbot1 0.00610795
R15351 mimbot1.n231 mimbot1.n230 0.00610795
R15352 mimbot1.n230 mimbot1 0.00610795
R15353 mimbot1 mimbot1.n229 0.00610795
R15354 mimbot1.n229 mimbot1 0.00610795
R15355 mimbot1.n13 mimbot1.n8 0.00527099
R15356 mimbot1.n23 mimbot1.n19 0.00527099
R15357 mimbot1.n279 mimbot1.n278 0.00523013
R15358 mimbot1.n332 mimbot1.n331 0.00523013
R15359 mimbot1.n382 mimbot1.n381 0.00523013
R15360 mimbot1.n402 mimbot1.n401 0.00523013
R15361 mimbot1.n683 mimbot1.n489 0.00523013
R15362 mimbot1.n544 mimbot1.n543 0.00523013
R15363 mimbot1.n555 mimbot1.n554 0.00523013
R15364 mimbot1.n566 mimbot1.n565 0.00523013
R15365 mimbot1.n533 mimbot1.n523 0.00523013
R15366 mimbot1.n441 mimbot1.n440 0.00523013
R15367 mimbot1.n452 mimbot1.n451 0.00523013
R15368 mimbot1.n463 mimbot1.n453 0.00523013
R15369 mimbot1.n712 mimbot1.n711 0.00523013
R15370 mimbot1.n168 mimbot1.n167 0.00523013
R15371 mimbot1.n243 mimbot1.n242 0.00523013
R15372 mimbot1.n343 mimbot1.n333 0.00523013
R15373 mimbot1.n223 mimbot1.n213 0.00523013
R15374 mimbot1.n190 mimbot1.n180 0.00523013
R15375 mimbot1.n179 mimbot1.n169 0.00523013
R15376 mimbot1.n321 mimbot1.n311 0.00523013
R15377 mimbot1.n201 mimbot1.n200 0.00523013
R15378 mimbot1.n212 mimbot1.n211 0.00523013
R15379 mimbot1.n301 mimbot1.n291 0.00523013
R15380 mimbot1.n290 mimbot1.n280 0.00523013
R15381 mimbot1.n411 mimbot1.n410 0.00523013
R15382 mimbot1.n421 mimbot1.n420 0.00523013
R15383 mimbot1.n513 mimbot1.n503 0.00523013
R15384 mimbot1.n502 mimbot1.n492 0.00523013
R15385 mimbot1.n724 mimbot1.n723 0.00501124
R15386 mimbot1.n632 mimbot1.n631 0.00476028
R15387 mimbot1.n645 mimbot1.n644 0.00476028
R15388 mimbot1.n650 mimbot1.n619 0.00476028
R15389 mimbot1.n662 mimbot1.n658 0.00476028
R15390 mimbot1.n680 mimbot1.n679 0.00476028
R15391 mimbot1.n611 mimbot1.n608 0.00476028
R15392 mimbot1.n681 mimbot1.n604 0.00476028
R15393 mimbot1.n692 mimbot1.n476 0.00476028
R15394 mimbot1.n695 mimbot1.n354 0.00476028
R15395 mimbot1.n718 mimbot1.n268 0.00476028
R15396 mimbot1.n598 mimbot1.n597 0.00476028
R15397 mimbot1.n582 mimbot1.n577 0.00476028
R15398 mimbot1.n681 mimbot1.n580 0.00476028
R15399 mimbot1.n692 mimbot1.n468 0.00476028
R15400 mimbot1.n695 mimbot1.n348 0.00476028
R15401 mimbot1.n718 mimbot1.n248 0.00476028
R15402 mimbot1.n723 mimbot1.n38 0.00476028
R15403 mimbot1.n150 mimbot1.n139 0.00476028
R15404 mimbot1.n142 mimbot1.n53 0.00476028
R15405 mimbot1.n133 mimbot1.n122 0.00476028
R15406 mimbot1.n125 mimbot1.n56 0.00476028
R15407 mimbot1.n110 mimbot1.n99 0.00476028
R15408 mimbot1.n102 mimbot1.n59 0.00476028
R15409 mimbot1.n87 mimbot1.n75 0.00476028
R15410 mimbot1.n79 mimbot1.n78 0.00476028
R15411 mimbot1.n24 mimbot1.n16 0.0047517
R15412 mimbot1.n410 mimbot1.n344 0.00473
R15413 mimbot1.n280 mimbot1.n244 0.00473
R15414 mimbot1.n695 mimbot1.n352 0.00473
R15415 mimbot1.n696 mimbot1.n253 0.00473
R15416 mimbot1.n695 mimbot1.n361 0.00473
R15417 mimbot1.n696 mimbot1.n263 0.00473
R15418 mimbot1.n401 mimbot1.n366 0.00473
R15419 mimbot1.n420 mimbot1.n367 0.00473
R15420 mimbot1.n492 mimbot1.n464 0.00473
R15421 mimbot1.n627 mimbot1.n576 0.00473
R15422 mimbot1.n649 mimbot1.n600 0.00473
R15423 mimbot1.n640 mimbot1.n621 0.00473
R15424 mimbot1.n675 mimbot1.n634 0.00473
R15425 mimbot1.n661 mimbot1.n647 0.00473
R15426 mimbot1.n681 mimbot1.n680 0.00473
R15427 mimbot1.n682 mimbot1.n478 0.00473
R15428 mimbot1.n681 mimbot1.n619 0.00473
R15429 mimbot1.n682 mimbot1.n481 0.00473
R15430 mimbot1.n610 mimbot1.n601 0.00473
R15431 mimbot1.n681 mimbot1.n608 0.00473
R15432 mimbot1.n682 mimbot1.n483 0.00473
R15433 mimbot1.n523 mimbot1.n472 0.00473
R15434 mimbot1.n692 mimbot1.n477 0.00473
R15435 mimbot1.n693 mimbot1.n361 0.00473
R15436 mimbot1.n681 mimbot1.n645 0.00473
R15437 mimbot1.n682 mimbot1.n477 0.00473
R15438 mimbot1.n691 mimbot1.n489 0.00473
R15439 mimbot1.n543 mimbot1.n487 0.00473
R15440 mimbot1.n692 mimbot1.n478 0.00473
R15441 mimbot1.n693 mimbot1.n362 0.00473
R15442 mimbot1.n451 mimbot1.n360 0.00473
R15443 mimbot1.n440 mimbot1.n364 0.00473
R15444 mimbot1.n692 mimbot1.n480 0.00473
R15445 mimbot1.n693 mimbot1.n352 0.00473
R15446 mimbot1.n681 mimbot1.n658 0.00473
R15447 mimbot1.n682 mimbot1.n480 0.00473
R15448 mimbot1.n554 mimbot1.n486 0.00473
R15449 mimbot1.n565 mimbot1.n484 0.00473
R15450 mimbot1.n692 mimbot1.n481 0.00473
R15451 mimbot1.n693 mimbot1.n357 0.00473
R15452 mimbot1.n692 mimbot1.n483 0.00473
R15453 mimbot1.n693 mimbot1.n353 0.00473
R15454 mimbot1.n453 mimbot1.n358 0.00473
R15455 mimbot1.n695 mimbot1.n353 0.00473
R15456 mimbot1.n717 mimbot1.n696 0.00473
R15457 mimbot1.n712 mimbot1.n252 0.00473
R15458 mimbot1.n718 mimbot1.n717 0.00473
R15459 mimbot1.n719 mimbot1.n51 0.00473
R15460 mimbot1.n242 mimbot1.n28 0.00473
R15461 mimbot1.n167 mimbot1.n49 0.00473
R15462 mimbot1.n718 mimbot1.n265 0.00473
R15463 mimbot1.n719 mimbot1.n29 0.00473
R15464 mimbot1.n695 mimbot1.n357 0.00473
R15465 mimbot1.n696 mimbot1.n265 0.00473
R15466 mimbot1.n333 mimbot1.n264 0.00473
R15467 mimbot1.n331 mimbot1.n255 0.00473
R15468 mimbot1.n718 mimbot1.n253 0.00473
R15469 mimbot1.n719 mimbot1.n48 0.00473
R15470 mimbot1.n169 mimbot1.n31 0.00473
R15471 mimbot1.n180 mimbot1.n46 0.00473
R15472 mimbot1.n718 mimbot1.n257 0.00473
R15473 mimbot1.n719 mimbot1.n32 0.00473
R15474 mimbot1.n695 mimbot1.n362 0.00473
R15475 mimbot1.n696 mimbot1.n257 0.00473
R15476 mimbot1.n311 mimbot1.n258 0.00473
R15477 mimbot1.n278 mimbot1.n261 0.00473
R15478 mimbot1.n718 mimbot1.n263 0.00473
R15479 mimbot1.n719 mimbot1.n45 0.00473
R15480 mimbot1.n718 mimbot1.n250 0.00473
R15481 mimbot1.n719 mimbot1.n40 0.00473
R15482 mimbot1.n211 mimbot1.n34 0.00473
R15483 mimbot1.n200 mimbot1.n43 0.00473
R15484 mimbot1.n718 mimbot1.n259 0.00473
R15485 mimbot1.n719 mimbot1.n35 0.00473
R15486 mimbot1.n695 mimbot1.n694 0.00473
R15487 mimbot1.n696 mimbot1.n259 0.00473
R15488 mimbot1.n695 mimbot1.n350 0.00473
R15489 mimbot1.n696 mimbot1.n250 0.00473
R15490 mimbot1.n692 mimbot1.n470 0.00473
R15491 mimbot1.n693 mimbot1.n350 0.00473
R15492 mimbot1.n692 mimbot1.n473 0.00473
R15493 mimbot1.n694 mimbot1.n693 0.00473
R15494 mimbot1.n681 mimbot1.n632 0.00473
R15495 mimbot1.n682 mimbot1.n473 0.00473
R15496 mimbot1.n681 mimbot1.n598 0.00473
R15497 mimbot1.n682 mimbot1.n470 0.00473
R15498 mimbot1.n593 mimbot1.n579 0.00473
R15499 mimbot1.n681 mimbot1.n577 0.00473
R15500 mimbot1.n682 mimbot1.n465 0.00473
R15501 mimbot1.n503 mimbot1.n467 0.00473
R15502 mimbot1.n692 mimbot1.n465 0.00473
R15503 mimbot1.n693 mimbot1.n345 0.00473
R15504 mimbot1.n381 mimbot1.n347 0.00473
R15505 mimbot1.n695 mimbot1.n345 0.00473
R15506 mimbot1.n696 mimbot1.n245 0.00473
R15507 mimbot1.n291 mimbot1.n247 0.00473
R15508 mimbot1.n718 mimbot1.n245 0.00473
R15509 mimbot1.n719 mimbot1.n42 0.00473
R15510 mimbot1.n213 mimbot1.n39 0.00473
R15511 mimbot1.n723 mimbot1.n42 0.00473
R15512 mimbot1.n151 mimbot1.n150 0.00473
R15513 mimbot1.n141 mimbot1.n134 0.00473
R15514 mimbot1.n723 mimbot1.n40 0.00473
R15515 mimbot1.n151 mimbot1.n53 0.00473
R15516 mimbot1.n118 mimbot1.n55 0.00473
R15517 mimbot1.n723 mimbot1.n35 0.00473
R15518 mimbot1.n151 mimbot1.n133 0.00473
R15519 mimbot1.n124 mimbot1.n111 0.00473
R15520 mimbot1.n723 mimbot1.n45 0.00473
R15521 mimbot1.n151 mimbot1.n56 0.00473
R15522 mimbot1.n95 mimbot1.n58 0.00473
R15523 mimbot1.n723 mimbot1.n32 0.00473
R15524 mimbot1.n151 mimbot1.n110 0.00473
R15525 mimbot1.n101 mimbot1.n88 0.00473
R15526 mimbot1.n723 mimbot1.n48 0.00473
R15527 mimbot1.n151 mimbot1.n59 0.00473
R15528 mimbot1.n71 mimbot1.n61 0.00473
R15529 mimbot1.n723 mimbot1.n29 0.00473
R15530 mimbot1.n151 mimbot1.n87 0.00473
R15531 mimbot1.n77 mimbot1.n64 0.00473
R15532 mimbot1.n723 mimbot1.n51 0.00473
R15533 mimbot1.n585 mimbot1.n581 0.00426062
R15534 mimbot1.n137 mimbot1.n52 0.00390244
R15535 mimbot1.n78 mimbot1.n63 0.00305965
R15536 mimbot1.n151 mimbot1.n63 0.00296185
R15537 mimbot1.n154 mimbot1.n51 0.00288031
R15538 mimbot1.n681 mimbot1.n599 0.00288031
R15539 mimbot1.n681 mimbot1.n620 0.00288031
R15540 mimbot1.n681 mimbot1.n633 0.00288031
R15541 mimbot1.n681 mimbot1.n646 0.00288031
R15542 mimbot1.n681 mimbot1.n659 0.00288031
R15543 mimbot1.n681 mimbot1.n602 0.00288031
R15544 mimbot1.n568 mimbot1.n483 0.00288031
R15545 mimbot1.n426 mimbot1.n353 0.00288031
R15546 mimbot1.n717 mimbot1.n697 0.00288031
R15547 mimbot1.n681 mimbot1.n578 0.00288031
R15548 mimbot1.n517 mimbot1.n465 0.00288031
R15549 mimbot1.n386 mimbot1.n345 0.00288031
R15550 mimbot1.n305 mimbot1.n245 0.00288031
R15551 mimbot1.n227 mimbot1.n42 0.00288031
R15552 mimbot1.n151 mimbot1.n135 0.00288031
R15553 mimbot1.n151 mimbot1.n54 0.00288031
R15554 mimbot1.n151 mimbot1.n112 0.00288031
R15555 mimbot1.n151 mimbot1.n57 0.00288031
R15556 mimbot1.n151 mimbot1.n89 0.00288031
R15557 mimbot1.n151 mimbot1.n60 0.00288031
R15558 mimbot1.n151 mimbot1.n65 0.00288031
R15559 mimbot1.n695 mimbot1.n351 0.00288014
R15560 mimbot1.n216 mimbot1.n40 0.00288014
R15561 mimbot1.n718 mimbot1.n251 0.00288014
R15562 mimbot1.n376 mimbot1.n350 0.00288014
R15563 mimbot1.n695 mimbot1.n365 0.00288014
R15564 mimbot1.n695 mimbot1.n368 0.00288014
R15565 mimbot1.n415 mimbot1.n361 0.00288014
R15566 mimbot1.n396 mimbot1.n362 0.00288014
R15567 mimbot1.n692 mimbot1.n471 0.00288014
R15568 mimbot1.n538 mimbot1.n480 0.00288014
R15569 mimbot1.n560 mimbot1.n483 0.00288014
R15570 mimbot1.n526 mimbot1.n477 0.00288014
R15571 mimbot1.n692 mimbot1.n474 0.00288014
R15572 mimbot1.n685 mimbot1.n478 0.00288014
R15573 mimbot1.n692 mimbot1.n488 0.00288014
R15574 mimbot1.n692 mimbot1.n479 0.00288014
R15575 mimbot1.n695 mimbot1.n359 0.00288014
R15576 mimbot1.n446 mimbot1.n357 0.00288014
R15577 mimbot1.n695 mimbot1.n363 0.00288014
R15578 mimbot1.n435 mimbot1.n352 0.00288014
R15579 mimbot1.n549 mimbot1.n481 0.00288014
R15580 mimbot1.n692 mimbot1.n485 0.00288014
R15581 mimbot1.n692 mimbot1.n482 0.00288014
R15582 mimbot1.n456 mimbot1.n353 0.00288014
R15583 mimbot1.n695 mimbot1.n356 0.00288014
R15584 mimbot1.n717 mimbot1.n716 0.00288014
R15585 mimbot1.n718 mimbot1.n266 0.00288014
R15586 mimbot1.n723 mimbot1.n50 0.00288014
R15587 mimbot1.n237 mimbot1.n51 0.00288014
R15588 mimbot1.n723 mimbot1.n30 0.00288014
R15589 mimbot1.n162 mimbot1.n29 0.00288014
R15590 mimbot1.n326 mimbot1.n265 0.00288014
R15591 mimbot1.n336 mimbot1.n253 0.00288014
R15592 mimbot1.n718 mimbot1.n256 0.00288014
R15593 mimbot1.n718 mimbot1.n254 0.00288014
R15594 mimbot1.n723 mimbot1.n47 0.00288014
R15595 mimbot1.n172 mimbot1.n48 0.00288014
R15596 mimbot1.n723 mimbot1.n33 0.00288014
R15597 mimbot1.n183 mimbot1.n32 0.00288014
R15598 mimbot1.n273 mimbot1.n257 0.00288014
R15599 mimbot1.n314 mimbot1.n263 0.00288014
R15600 mimbot1.n718 mimbot1.n260 0.00288014
R15601 mimbot1.n718 mimbot1.n262 0.00288014
R15602 mimbot1.n723 mimbot1.n44 0.00288014
R15603 mimbot1.n206 mimbot1.n45 0.00288014
R15604 mimbot1.n723 mimbot1.n36 0.00288014
R15605 mimbot1.n195 mimbot1.n35 0.00288014
R15606 mimbot1.n283 mimbot1.n259 0.00288014
R15607 mimbot1.n294 mimbot1.n250 0.00288014
R15608 mimbot1.n694 mimbot1.n371 0.00288014
R15609 mimbot1.n495 mimbot1.n473 0.00288014
R15610 mimbot1.n506 mimbot1.n470 0.00288014
R15611 mimbot1.n692 mimbot1.n466 0.00288014
R15612 mimbot1.n695 mimbot1.n346 0.00288014
R15613 mimbot1.n718 mimbot1.n246 0.00288014
R15614 mimbot1.n723 mimbot1.n41 0.00288014
R15615 mimbot1.n721 mimbot1.n153 0.00238
R15616 mimbot1.n569 mimbot1.n567 0.00238
R15617 mimbot1.n429 mimbot1.n428 0.00238
R15618 mimbot1.n703 mimbot1.n701 0.00238
R15619 mimbot1.n515 mimbot1.n514 0.00238
R15620 mimbot1.n384 mimbot1.n383 0.00238
R15621 mimbot1.n303 mimbot1.n302 0.00238
R15622 mimbot1.n225 mimbot1.n224 0.00238
R15623 mimbot1.n607 mimbot1.n606 0.00231712
R15624 mimbot1.n156 mimbot1.n154 0.00175031
R15625 mimbot1.n625 mimbot1.n599 0.00175031
R15626 mimbot1.n655 mimbot1.n620 0.00175031
R15627 mimbot1.n638 mimbot1.n633 0.00175031
R15628 mimbot1.n673 mimbot1.n646 0.00175031
R15629 mimbot1.n667 mimbot1.n659 0.00175031
R15630 mimbot1.n616 mimbot1.n602 0.00175031
R15631 mimbot1.n573 mimbot1.n568 0.00175031
R15632 mimbot1.n426 mimbot1.n425 0.00175031
R15633 mimbot1.n698 mimbot1.n697 0.00175031
R15634 mimbot1.n591 mimbot1.n578 0.00175031
R15635 mimbot1.n520 mimbot1.n517 0.00175031
R15636 mimbot1.n389 mimbot1.n386 0.00175031
R15637 mimbot1.n308 mimbot1.n305 0.00175031
R15638 mimbot1.n230 mimbot1.n227 0.00175031
R15639 mimbot1.n147 mimbot1.n135 0.00175031
R15640 mimbot1.n116 mimbot1.n54 0.00175031
R15641 mimbot1.n130 mimbot1.n112 0.00175031
R15642 mimbot1.n93 mimbot1.n57 0.00175031
R15643 mimbot1.n107 mimbot1.n89 0.00175031
R15644 mimbot1.n69 mimbot1.n60 0.00175031
R15645 mimbot1.n84 mimbot1.n65 0.00175031
R15646 mimbot1.n13 mimbot1.n12 0.00112135
R15647 mimbot1.n155 mimbot1.n154 0.00100031
R15648 mimbot1.n629 mimbot1.n599 0.00100031
R15649 mimbot1.n654 mimbot1.n620 0.00100031
R15650 mimbot1.n642 mimbot1.n633 0.00100031
R15651 mimbot1.n677 mimbot1.n646 0.00100031
R15652 mimbot1.n666 mimbot1.n659 0.00100031
R15653 mimbot1.n615 mimbot1.n602 0.00100031
R15654 mimbot1.n571 mimbot1.n568 0.00100031
R15655 mimbot1.n427 mimbot1.n426 0.00100031
R15656 mimbot1.n704 mimbot1.n697 0.00100031
R15657 mimbot1.n595 mimbot1.n578 0.00100031
R15658 mimbot1.n519 mimbot1.n517 0.00100031
R15659 mimbot1.n388 mimbot1.n386 0.00100031
R15660 mimbot1.n307 mimbot1.n305 0.00100031
R15661 mimbot1.n229 mimbot1.n227 0.00100031
R15662 mimbot1.n146 mimbot1.n135 0.00100031
R15663 mimbot1.n120 mimbot1.n54 0.00100031
R15664 mimbot1.n129 mimbot1.n112 0.00100031
R15665 mimbot1.n97 mimbot1.n57 0.00100031
R15666 mimbot1.n106 mimbot1.n89 0.00100031
R15667 mimbot1.n73 mimbot1.n60 0.00100031
R15668 mimbot1.n83 mimbot1.n65 0.00100031
R15669 mimbot1.n26 mimbot1.n6 0.000784848
R15670 mimbot1.n5 mimbot1.n4 0.000784848
R15671 mimbot1.n24 mimbot1.n13 0.000687305
R15672 mimbot1.n24 mimbot1.n23 0.000687305
R15673 mimbot1.n222 mimbot1.n214 0.000500621
R15674 mimbot1.n220 mimbot1.n214 0.000500621
R15675 mimbot1.n222 mimbot1.n221 0.000500621
R15676 mimbot1.n221 mimbot1.n220 0.000500621
R15677 mimbot1.n156 mimbot1.n153 0.000500621
R15678 mimbot1.n155 mimbot1.n153 0.000500621
R15679 mimbot1.n156 mimbot1.n152 0.000500621
R15680 mimbot1.n155 mimbot1.n152 0.000500621
R15681 mimbot1.n373 mimbot1.n372 0.000500621
R15682 mimbot1.n379 mimbot1.n373 0.000500621
R15683 mimbot1.n380 mimbot1.n372 0.000500621
R15684 mimbot1.n380 mimbot1.n379 0.000500621
R15685 mimbot1.n413 mimbot1.n412 0.000500621
R15686 mimbot1.n418 mimbot1.n413 0.000500621
R15687 mimbot1.n419 mimbot1.n412 0.000500621
R15688 mimbot1.n419 mimbot1.n418 0.000500621
R15689 mimbot1.n393 mimbot1.n392 0.000500621
R15690 mimbot1.n399 mimbot1.n393 0.000500621
R15691 mimbot1.n400 mimbot1.n392 0.000500621
R15692 mimbot1.n400 mimbot1.n399 0.000500621
R15693 mimbot1.n626 mimbot1.n625 0.000500621
R15694 mimbot1.n630 mimbot1.n622 0.000500621
R15695 mimbot1.n629 mimbot1.n628 0.000500621
R15696 mimbot1.n625 mimbot1.n576 0.000500621
R15697 mimbot1.n629 mimbot1.n576 0.000500621
R15698 mimbot1.n639 mimbot1.n638 0.000500621
R15699 mimbot1.n643 mimbot1.n635 0.000500621
R15700 mimbot1.n642 mimbot1.n641 0.000500621
R15701 mimbot1.n656 mimbot1.n655 0.000500621
R15702 mimbot1.n652 mimbot1.n651 0.000500621
R15703 mimbot1.n654 mimbot1.n653 0.000500621
R15704 mimbot1.n655 mimbot1.n600 0.000500621
R15705 mimbot1.n654 mimbot1.n600 0.000500621
R15706 mimbot1.n638 mimbot1.n621 0.000500621
R15707 mimbot1.n642 mimbot1.n621 0.000500621
R15708 mimbot1.n668 mimbot1.n667 0.000500621
R15709 mimbot1.n664 mimbot1.n663 0.000500621
R15710 mimbot1.n666 mimbot1.n665 0.000500621
R15711 mimbot1.n674 mimbot1.n673 0.000500621
R15712 mimbot1.n678 mimbot1.n670 0.000500621
R15713 mimbot1.n677 mimbot1.n676 0.000500621
R15714 mimbot1.n673 mimbot1.n634 0.000500621
R15715 mimbot1.n677 mimbot1.n634 0.000500621
R15716 mimbot1.n667 mimbot1.n647 0.000500621
R15717 mimbot1.n666 mimbot1.n647 0.000500621
R15718 mimbot1.n535 mimbot1.n534 0.000500621
R15719 mimbot1.n541 mimbot1.n535 0.000500621
R15720 mimbot1.n542 mimbot1.n534 0.000500621
R15721 mimbot1.n542 mimbot1.n541 0.000500621
R15722 mimbot1.n557 mimbot1.n556 0.000500621
R15723 mimbot1.n563 mimbot1.n557 0.000500621
R15724 mimbot1.n564 mimbot1.n556 0.000500621
R15725 mimbot1.n564 mimbot1.n563 0.000500621
R15726 mimbot1.n617 mimbot1.n616 0.000500621
R15727 mimbot1.n613 mimbot1.n612 0.000500621
R15728 mimbot1.n615 mimbot1.n614 0.000500621
R15729 mimbot1.n616 mimbot1.n601 0.000500621
R15730 mimbot1.n615 mimbot1.n601 0.000500621
R15731 mimbot1.n605 mimbot1.n603 0.000500621
R15732 mimbot1.n573 mimbot1.n572 0.000500621
R15733 mimbot1.n573 mimbot1.n569 0.000500621
R15734 mimbot1.n572 mimbot1.n571 0.000500621
R15735 mimbot1.n571 mimbot1.n569 0.000500621
R15736 mimbot1.n532 mimbot1.n524 0.000500621
R15737 mimbot1.n530 mimbot1.n524 0.000500621
R15738 mimbot1.n532 mimbot1.n531 0.000500621
R15739 mimbot1.n531 mimbot1.n530 0.000500621
R15740 mimbot1.n570 mimbot1.n475 0.000500621
R15741 mimbot1.n684 mimbot1.n491 0.000500621
R15742 mimbot1.n689 mimbot1.n491 0.000500621
R15743 mimbot1.n688 mimbot1.n684 0.000500621
R15744 mimbot1.n689 mimbot1.n688 0.000500621
R15745 mimbot1.n425 mimbot1.n423 0.000500621
R15746 mimbot1.n427 mimbot1.n423 0.000500621
R15747 mimbot1.n428 mimbot1.n425 0.000500621
R15748 mimbot1.n428 mimbot1.n427 0.000500621
R15749 mimbot1.n443 mimbot1.n442 0.000500621
R15750 mimbot1.n449 mimbot1.n443 0.000500621
R15751 mimbot1.n450 mimbot1.n442 0.000500621
R15752 mimbot1.n450 mimbot1.n449 0.000500621
R15753 mimbot1.n432 mimbot1.n431 0.000500621
R15754 mimbot1.n438 mimbot1.n432 0.000500621
R15755 mimbot1.n439 mimbot1.n431 0.000500621
R15756 mimbot1.n439 mimbot1.n438 0.000500621
R15757 mimbot1.n546 mimbot1.n545 0.000500621
R15758 mimbot1.n552 mimbot1.n546 0.000500621
R15759 mimbot1.n553 mimbot1.n545 0.000500621
R15760 mimbot1.n553 mimbot1.n552 0.000500621
R15761 mimbot1.n462 mimbot1.n454 0.000500621
R15762 mimbot1.n460 mimbot1.n454 0.000500621
R15763 mimbot1.n462 mimbot1.n461 0.000500621
R15764 mimbot1.n461 mimbot1.n460 0.000500621
R15765 mimbot1.n424 mimbot1.n355 0.000500621
R15766 mimbot1.n705 mimbot1.n698 0.000500621
R15767 mimbot1.n703 mimbot1.n698 0.000500621
R15768 mimbot1.n705 mimbot1.n704 0.000500621
R15769 mimbot1.n704 mimbot1.n703 0.000500621
R15770 mimbot1.n709 mimbot1.n708 0.000500621
R15771 mimbot1.n714 mimbot1.n709 0.000500621
R15772 mimbot1.n713 mimbot1.n708 0.000500621
R15773 mimbot1.n714 mimbot1.n713 0.000500621
R15774 mimbot1.n702 mimbot1.n267 0.000500621
R15775 mimbot1.n234 mimbot1.n233 0.000500621
R15776 mimbot1.n240 mimbot1.n234 0.000500621
R15777 mimbot1.n241 mimbot1.n233 0.000500621
R15778 mimbot1.n241 mimbot1.n240 0.000500621
R15779 mimbot1.n159 mimbot1.n158 0.000500621
R15780 mimbot1.n165 mimbot1.n159 0.000500621
R15781 mimbot1.n166 mimbot1.n158 0.000500621
R15782 mimbot1.n166 mimbot1.n165 0.000500621
R15783 mimbot1.n323 mimbot1.n322 0.000500621
R15784 mimbot1.n329 mimbot1.n323 0.000500621
R15785 mimbot1.n330 mimbot1.n322 0.000500621
R15786 mimbot1.n330 mimbot1.n329 0.000500621
R15787 mimbot1.n342 mimbot1.n334 0.000500621
R15788 mimbot1.n340 mimbot1.n334 0.000500621
R15789 mimbot1.n342 mimbot1.n341 0.000500621
R15790 mimbot1.n341 mimbot1.n340 0.000500621
R15791 mimbot1.n178 mimbot1.n170 0.000500621
R15792 mimbot1.n176 mimbot1.n170 0.000500621
R15793 mimbot1.n178 mimbot1.n177 0.000500621
R15794 mimbot1.n177 mimbot1.n176 0.000500621
R15795 mimbot1.n189 mimbot1.n181 0.000500621
R15796 mimbot1.n187 mimbot1.n181 0.000500621
R15797 mimbot1.n189 mimbot1.n188 0.000500621
R15798 mimbot1.n188 mimbot1.n187 0.000500621
R15799 mimbot1.n270 mimbot1.n269 0.000500621
R15800 mimbot1.n276 mimbot1.n270 0.000500621
R15801 mimbot1.n277 mimbot1.n269 0.000500621
R15802 mimbot1.n277 mimbot1.n276 0.000500621
R15803 mimbot1.n320 mimbot1.n312 0.000500621
R15804 mimbot1.n318 mimbot1.n312 0.000500621
R15805 mimbot1.n320 mimbot1.n319 0.000500621
R15806 mimbot1.n319 mimbot1.n318 0.000500621
R15807 mimbot1.n203 mimbot1.n202 0.000500621
R15808 mimbot1.n209 mimbot1.n203 0.000500621
R15809 mimbot1.n210 mimbot1.n202 0.000500621
R15810 mimbot1.n210 mimbot1.n209 0.000500621
R15811 mimbot1.n192 mimbot1.n191 0.000500621
R15812 mimbot1.n198 mimbot1.n192 0.000500621
R15813 mimbot1.n199 mimbot1.n191 0.000500621
R15814 mimbot1.n199 mimbot1.n198 0.000500621
R15815 mimbot1.n289 mimbot1.n281 0.000500621
R15816 mimbot1.n287 mimbot1.n281 0.000500621
R15817 mimbot1.n289 mimbot1.n288 0.000500621
R15818 mimbot1.n288 mimbot1.n287 0.000500621
R15819 mimbot1.n300 mimbot1.n292 0.000500621
R15820 mimbot1.n298 mimbot1.n292 0.000500621
R15821 mimbot1.n300 mimbot1.n299 0.000500621
R15822 mimbot1.n299 mimbot1.n298 0.000500621
R15823 mimbot1.n404 mimbot1.n403 0.000500621
R15824 mimbot1.n408 mimbot1.n404 0.000500621
R15825 mimbot1.n409 mimbot1.n403 0.000500621
R15826 mimbot1.n409 mimbot1.n408 0.000500621
R15827 mimbot1.n501 mimbot1.n493 0.000500621
R15828 mimbot1.n499 mimbot1.n493 0.000500621
R15829 mimbot1.n501 mimbot1.n500 0.000500621
R15830 mimbot1.n500 mimbot1.n499 0.000500621
R15831 mimbot1.n512 mimbot1.n504 0.000500621
R15832 mimbot1.n510 mimbot1.n504 0.000500621
R15833 mimbot1.n512 mimbot1.n511 0.000500621
R15834 mimbot1.n511 mimbot1.n510 0.000500621
R15835 mimbot1.n592 mimbot1.n591 0.000500621
R15836 mimbot1.n596 mimbot1.n588 0.000500621
R15837 mimbot1.n595 mimbot1.n594 0.000500621
R15838 mimbot1.n584 mimbot1.n583 0.000500621
R15839 mimbot1.n587 mimbot1.n586 0.000500621
R15840 mimbot1.n591 mimbot1.n579 0.000500621
R15841 mimbot1.n595 mimbot1.n579 0.000500621
R15842 mimbot1.n520 mimbot1.n516 0.000500621
R15843 mimbot1.n519 mimbot1.n516 0.000500621
R15844 mimbot1.n520 mimbot1.n515 0.000500621
R15845 mimbot1.n519 mimbot1.n515 0.000500621
R15846 mimbot1.n518 mimbot1.n469 0.000500621
R15847 mimbot1.n389 mimbot1.n385 0.000500621
R15848 mimbot1.n388 mimbot1.n385 0.000500621
R15849 mimbot1.n389 mimbot1.n384 0.000500621
R15850 mimbot1.n388 mimbot1.n384 0.000500621
R15851 mimbot1.n387 mimbot1.n349 0.000500621
R15852 mimbot1.n308 mimbot1.n304 0.000500621
R15853 mimbot1.n307 mimbot1.n304 0.000500621
R15854 mimbot1.n308 mimbot1.n303 0.000500621
R15855 mimbot1.n307 mimbot1.n303 0.000500621
R15856 mimbot1.n306 mimbot1.n249 0.000500621
R15857 mimbot1.n230 mimbot1.n226 0.000500621
R15858 mimbot1.n229 mimbot1.n226 0.000500621
R15859 mimbot1.n230 mimbot1.n225 0.000500621
R15860 mimbot1.n229 mimbot1.n225 0.000500621
R15861 mimbot1.n228 mimbot1.n37 0.000500621
R15862 mimbot1.n138 mimbot1.n136 0.000500621
R15863 mimbot1.n148 mimbot1.n147 0.000500621
R15864 mimbot1.n146 mimbot1.n145 0.000500621
R15865 mimbot1.n144 mimbot1.n143 0.000500621
R15866 mimbot1.n147 mimbot1.n134 0.000500621
R15867 mimbot1.n146 mimbot1.n134 0.000500621
R15868 mimbot1.n117 mimbot1.n116 0.000500621
R15869 mimbot1.n120 mimbot1.n119 0.000500621
R15870 mimbot1.n121 mimbot1.n113 0.000500621
R15871 mimbot1.n116 mimbot1.n55 0.000500621
R15872 mimbot1.n120 mimbot1.n55 0.000500621
R15873 mimbot1.n131 mimbot1.n130 0.000500621
R15874 mimbot1.n129 mimbot1.n128 0.000500621
R15875 mimbot1.n127 mimbot1.n126 0.000500621
R15876 mimbot1.n130 mimbot1.n111 0.000500621
R15877 mimbot1.n129 mimbot1.n111 0.000500621
R15878 mimbot1.n94 mimbot1.n93 0.000500621
R15879 mimbot1.n97 mimbot1.n96 0.000500621
R15880 mimbot1.n98 mimbot1.n90 0.000500621
R15881 mimbot1.n93 mimbot1.n58 0.000500621
R15882 mimbot1.n97 mimbot1.n58 0.000500621
R15883 mimbot1.n108 mimbot1.n107 0.000500621
R15884 mimbot1.n106 mimbot1.n105 0.000500621
R15885 mimbot1.n104 mimbot1.n103 0.000500621
R15886 mimbot1.n107 mimbot1.n88 0.000500621
R15887 mimbot1.n106 mimbot1.n88 0.000500621
R15888 mimbot1.n70 mimbot1.n69 0.000500621
R15889 mimbot1.n73 mimbot1.n72 0.000500621
R15890 mimbot1.n74 mimbot1.n66 0.000500621
R15891 mimbot1.n69 mimbot1.n61 0.000500621
R15892 mimbot1.n73 mimbot1.n61 0.000500621
R15893 mimbot1.n85 mimbot1.n84 0.000500621
R15894 mimbot1.n83 mimbot1.n82 0.000500621
R15895 mimbot1.n81 mimbot1.n80 0.000500621
R15896 mimbot1.n84 mimbot1.n64 0.000500621
R15897 mimbot1.n83 mimbot1.n64 0.000500621
R15898 mimbot1.n722 mimbot1.n27 0.000500621
R15899 mimbot1.n407 mimbot1.n344 0.00050031
R15900 mimbot1.n218 mimbot1.n217 0.00050031
R15901 mimbot1.n286 mimbot1.n244 0.00050031
R15902 mimbot1.n377 mimbot1.n374 0.00050031
R15903 mimbot1.n398 mimbot1.n366 0.00050031
R15904 mimbot1.n417 mimbot1.n367 0.00050031
R15905 mimbot1.n416 mimbot1.n414 0.00050031
R15906 mimbot1.n397 mimbot1.n394 0.00050031
R15907 mimbot1.n498 mimbot1.n464 0.00050031
R15908 mimbot1.n539 mimbot1.n536 0.00050031
R15909 mimbot1.n561 mimbot1.n558 0.00050031
R15910 mimbot1.n528 mimbot1.n527 0.00050031
R15911 mimbot1.n529 mimbot1.n472 0.00050031
R15912 mimbot1.n687 mimbot1.n686 0.00050031
R15913 mimbot1.n691 mimbot1.n690 0.00050031
R15914 mimbot1.n540 mimbot1.n487 0.00050031
R15915 mimbot1.n448 mimbot1.n360 0.00050031
R15916 mimbot1.n447 mimbot1.n444 0.00050031
R15917 mimbot1.n437 mimbot1.n364 0.00050031
R15918 mimbot1.n436 mimbot1.n433 0.00050031
R15919 mimbot1.n550 mimbot1.n547 0.00050031
R15920 mimbot1.n551 mimbot1.n486 0.00050031
R15921 mimbot1.n562 mimbot1.n484 0.00050031
R15922 mimbot1.n458 mimbot1.n457 0.00050031
R15923 mimbot1.n459 mimbot1.n358 0.00050031
R15924 mimbot1.n715 mimbot1.n706 0.00050031
R15925 mimbot1.n710 mimbot1.n252 0.00050031
R15926 mimbot1.n239 mimbot1.n28 0.00050031
R15927 mimbot1.n238 mimbot1.n235 0.00050031
R15928 mimbot1.n164 mimbot1.n49 0.00050031
R15929 mimbot1.n163 mimbot1.n160 0.00050031
R15930 mimbot1.n327 mimbot1.n324 0.00050031
R15931 mimbot1.n338 mimbot1.n337 0.00050031
R15932 mimbot1.n339 mimbot1.n264 0.00050031
R15933 mimbot1.n328 mimbot1.n255 0.00050031
R15934 mimbot1.n175 mimbot1.n31 0.00050031
R15935 mimbot1.n174 mimbot1.n173 0.00050031
R15936 mimbot1.n186 mimbot1.n46 0.00050031
R15937 mimbot1.n185 mimbot1.n184 0.00050031
R15938 mimbot1.n274 mimbot1.n271 0.00050031
R15939 mimbot1.n316 mimbot1.n315 0.00050031
R15940 mimbot1.n317 mimbot1.n258 0.00050031
R15941 mimbot1.n275 mimbot1.n261 0.00050031
R15942 mimbot1.n208 mimbot1.n34 0.00050031
R15943 mimbot1.n207 mimbot1.n204 0.00050031
R15944 mimbot1.n197 mimbot1.n43 0.00050031
R15945 mimbot1.n196 mimbot1.n193 0.00050031
R15946 mimbot1.n285 mimbot1.n284 0.00050031
R15947 mimbot1.n296 mimbot1.n295 0.00050031
R15948 mimbot1.n406 mimbot1.n370 0.00050031
R15949 mimbot1.n497 mimbot1.n496 0.00050031
R15950 mimbot1.n508 mimbot1.n507 0.00050031
R15951 mimbot1.n509 mimbot1.n467 0.00050031
R15952 mimbot1.n378 mimbot1.n347 0.00050031
R15953 mimbot1.n297 mimbot1.n247 0.00050031
R15954 mimbot1.n219 mimbot1.n39 0.00050031
R15955 clk.n1 clk.t3 229.433
R15956 clk.n0 clk.t2 229.04
R15957 clk.n1 clk.t1 158.886
R15958 clk.n0 clk.t0 158.46
R15959 clk.n7 clk 38.8978
R15960 clk.n8 clk.n0 8.7103
R15961 clk.n2 clk.n1 7.39078
R15962 clk.n4 clk.n3 3.46717
R15963 clk clk.n8 3.16209
R15964 clk.n6 clk.n4 3.03598
R15965 clk.n7 clk.n6 2.61367
R15966 clk.n8 clk.n7 2.26586
R15967 clk.n4 clk.n2 1.06717
R15968 clk.n3 clk 1.06717
R15969 clk.n6 clk.n5 0.00666568
C0 a_3724_38568# phi1_n 8.88e-21
C1 mimbot1 a_3227_38050# 0.0119f
C2 sky130_fd_sc_hd__inv_1_0.A sky130_fd_sc_hd__inv_1_1.A 0.0104f
C3 sky130_fd_sc_hd__inv_1_2.A sky130_fd_sc_hd__inv_1_0.A 0.0876f
C4 mimbot1 a_3227_37506# 0.00858f
C5 a_4041_38050# a_4041_37506# 0.0137f
C6 phi1 a_3172_38568# 0.0991f
C7 sky130_fd_sc_hd__inv_1_3.Y a_3227_38050# 0.0536f
C8 VDD a_2944_38050# 0.198f
C9 sky130_fd_sc_hd__inv_1_3.Y a_3227_37506# 0.00861f
C10 a_2201_38050# a_2590_38050# 7.09e-19
C11 VDD a_2944_37506# 0.202f
C12 sky130_fd_sc_hd__nand2_1_0.Y a_2944_38050# 2.42e-19
C13 a_2307_38050# a_2484_38050# 0.16f
C14 phi1_n a_2024_38050# 0.00446f
C15 vcm sky130_fd_sc_hd__inv_1_2.Y 0.216f
C16 phi1_n a_2024_37506# 1.73e-19
C17 a_3724_36936# sky130_fd_sc_hd__inv_1_3.A 0.191f
C18 mimbot1 phi2_n 0.16f
C19 a_2201_37506# a_2590_37506# 7.09e-19
C20 a_2307_37506# a_2484_37506# 0.16f
C21 sky130_fd_sc_hd__nand2_1_1.Y a_2944_37506# 1.85e-19
C22 sky130_fd_sc_hd__dlymetal6s6s_1_3.A a_4147_38050# 6.53e-19
C23 sky130_fd_sc_hd__inv_1_2.Y a_3510_38050# 0.0222f
C24 mimbot1 mimtop1 1.27p
C25 sky130_fd_sc_hd__inv_1_3.Y phi2_n 0.00921f
C26 sky130_fd_sc_hd__inv_1_2.Y a_3510_37506# 0.0264f
C27 sky130_fd_sc_hd__dlymetal6s6s_1_5.A a_4147_37506# 6.53e-19
C28 a_3121_37506# sky130_fd_sc_hd__inv_1_1.A 1.91e-20
C29 mimtop2 a_2590_38050# 0.0398f
C30 VDD sky130_fd_sc_hd__dlymetal6s6s_1_2.A 0.237f
C31 VDD phi1_n 1.05f
C32 mimtop1 sky130_fd_sc_hd__inv_1_3.Y 0.00363f
C33 sky130_fd_sc_hd__nand2_1_0.Y sky130_fd_sc_hd__dlymetal6s6s_1_2.A 6.15e-19
C34 VDD sky130_fd_sc_hd__dlymetal6s6s_1_4.A 0.247f
C35 mimtop2 a_2590_37506# 0.0383f
C36 phi1_n sky130_fd_sc_hd__nand2_1_0.Y 0.00628f
C37 phi1_n sky130_fd_sc_hd__nand2_1_1.Y 2.53e-19
C38 sky130_fd_sc_hd__dlymetal6s6s_1_5.A phi2 7.55e-19
C39 sky130_fd_sc_hd__nand2_1_1.Y sky130_fd_sc_hd__dlymetal6s6s_1_4.A 6.68e-19
C40 phi1_n a_3172_36936# 1.3e-20
C41 vcm mimbot1 0.769p
C42 mimtop1 a_1794_38050# 2.18e-19
C43 mimtop1 a_1798_37826# 2.3e-19
C44 vcm sky130_fd_sc_hd__inv_1_3.Y 0.21f
C45 mimbot1 a_3510_38050# 0.00204f
C46 a_4041_38050# a_4324_38050# 0.0145f
C47 sky130_fd_sc_hd__inv_1_2.Y a_4041_38050# 0.00151f
C48 a_4147_38050# a_4147_37506# 0.0126f
C49 mimbot1 a_3510_37506# 0.00154f
C50 sky130_fd_sc_hd__inv_1_2.Y a_4041_37506# 3.08e-19
C51 sky130_fd_sc_hd__inv_1_3.Y a_3510_38050# 0.063f
C52 a_4041_37506# a_4324_37506# 0.0145f
C53 VDD a_3227_38050# 0.168f
C54 a_2024_38050# phi2_n 1.12e-19
C55 sky130_fd_sc_hd__inv_1_3.Y a_3510_37506# 0.0273f
C56 vcm a_1794_38050# 2.27e-19
C57 sky130_fd_sc_hd__nand2_1_0.Y a_3227_38050# 1.44e-19
C58 a_2484_38050# a_2590_38050# 0.322f
C59 VDD a_3227_37506# 0.173f
C60 phi1_n a_2307_38050# 0.00322f
C61 a_2024_37506# phi2_n 0.00574f
C62 a_3172_38568# phi2 3.43e-21
C63 mimtop1 a_2024_38050# 1.81e-19
C64 a_2484_38050# a_2590_37506# 4.65e-19
C65 vcm a_1798_37826# 2.3e-19
C66 a_2590_38050# a_2484_37506# 4.65e-19
C67 phi1_n a_2307_37506# 8.42e-20
C68 mimtop1 a_2024_37506# 2.14e-21
C69 sky130_fd_sc_hd__nand2_1_1.Y a_3227_37506# 1.19e-19
C70 a_2484_37506# a_2590_37506# 0.322f
C71 a_3227_38050# a_3172_36936# 1.02e-19
C72 a_3227_37506# a_3172_36936# 0.00449f
C73 VDD phi2_n 0.919f
C74 a_3404_37506# sky130_fd_sc_hd__inv_1_1.A 2.97e-20
C75 sky130_fd_sc_hd__nand2_1_0.Y phi2_n 2.59e-20
C76 mimbot1 a_4041_38050# 0.00226f
C77 VDD mimtop1 1.58f
C78 vcm a_2024_38050# 0.0628f
C79 sky130_fd_sc_hd__nand2_1_1.Y phi2_n 0.00587f
C80 mimtop1 sky130_fd_sc_hd__nand2_1_0.Y 0.0311f
C81 vcm a_2024_37506# 0.0611f
C82 sky130_fd_sc_hd__inv_1_3.Y a_4041_38050# 0.0039f
C83 a_3172_36936# phi2_n 0.224f
C84 mimtop1 sky130_fd_sc_hd__nand2_1_1.Y 0.0297f
C85 sky130_fd_sc_hd__inv_1_3.Y a_4041_37506# 0.00678f
C86 mimtop1 a_3172_36936# 2.61e-19
C87 sky130_fd_sc_hd__inv_1_0.A a_2944_38050# 6.92e-21
C88 VDD vcm 46.2f
C89 sky130_fd_sc_hd__inv_1_2.Y a_4324_38050# 6.66e-19
C90 vcm sky130_fd_sc_hd__nand2_1_0.Y 0.179f
C91 a_4324_38050# a_4324_37506# 0.0137f
C92 sky130_fd_sc_hd__inv_1_2.Y a_4324_37506# 1.31e-19
C93 vcm sky130_fd_sc_hd__nand2_1_1.Y 0.171f
C94 a_3724_38568# a_4041_38050# 7.18e-20
C95 a_3864_37506# sky130_fd_sc_hd__inv_1_1.A 0.00215f
C96 VDD a_3510_38050# 0.178f
C97 a_2307_38050# phi2_n 8.17e-20
C98 phi1 sky130_fd_sc_hd__inv_1_2.A 0.00272f
C99 VDD a_3510_37506# 0.181f
C100 sky130_fd_sc_hd__nand2_1_0.Y a_3510_38050# 7.34e-20
C101 a_2590_38050# sky130_fd_sc_hd__dlymetal6s6s_1_2.A 0.153f
C102 phi1_n a_2590_38050# 0.00604f
C103 a_2307_37506# phi2_n 0.00283f
C104 mimtop1 a_2307_38050# 0.0012f
C105 phi1_n a_2590_37506# 1.2e-19
C106 clk sky130_fd_sc_hd__inv_1_4.Y 0.0908f
C107 sky130_fd_sc_hd__inv_1_0.A phi1_n 1.03e-20
C108 a_2590_37506# sky130_fd_sc_hd__dlymetal6s6s_1_4.A 0.153f
C109 sky130_fd_sc_hd__nand2_1_1.Y a_3510_37506# 2.97e-20
C110 a_2944_38050# a_3121_38050# 0.16f
C111 sky130_fd_sc_hd__dlymetal6s6s_1_5.A sky130_fd_sc_hd__inv_1_1.A 0.00211f
C112 a_2944_37506# a_3121_37506# 0.16f
C113 mimbot1 a_4324_38050# 0.00152f
C114 mimbot1 sky130_fd_sc_hd__inv_1_2.Y 0.165f
C115 vcm a_2307_38050# 0.0198f
C116 vcm a_2307_37506# 0.0173f
C117 sky130_fd_sc_hd__inv_1_3.Y a_4324_38050# 0.00181f
C118 sky130_fd_sc_hd__inv_1_2.Y sky130_fd_sc_hd__inv_1_3.Y 0.279f
C119 VDD a_4041_38050# 0.204f
C120 sky130_fd_sc_hd__inv_1_3.Y a_4324_37506# 0.00309f
C121 sky130_fd_sc_hd__dlymetal6s6s_1_2.A a_3121_38050# 0.0146f
C122 VDD a_4041_37506# 0.204f
C123 phi1 mimtop2 0.0558f
C124 phi1_n a_3121_38050# 4.05e-19
C125 sky130_fd_sc_hd__inv_1_0.A a_3227_38050# 1.31e-20
C126 a_3864_38050# a_3724_36936# 1.92e-19
C127 sky130_fd_sc_hd__dlymetal6s6s_1_4.A a_3121_37506# 0.0146f
C128 a_3864_37506# a_3724_36936# 0.00416f
C129 phi1 a_3724_36936# 3.94e-20
C130 a_4430_38050# a_4430_37506# 0.0126f
C131 sky130_fd_sc_hd__inv_1_2.Y a_1798_37826# 1.16e-19
C132 sky130_fd_sc_hd__inv_1_2.A a_4147_38050# 0.0111f
C133 a_4147_37506# sky130_fd_sc_hd__inv_1_1.A 0.00429f
C134 sky130_fd_sc_hd__inv_1_2.Y a_3724_38568# 0.171f
C135 a_3172_38568# sky130_fd_sc_hd__inv_1_2.A 7.06e-21
C136 a_2590_38050# phi2_n 1.28e-19
C137 sky130_fd_sc_hd__inv_1_2.A a_4147_37506# 3.52e-21
C138 a_2590_37506# phi2_n 0.00393f
C139 mimtop1 a_2590_38050# 5.6e-19
C140 mimbot1 sky130_fd_sc_hd__inv_1_3.Y 0.134f
C141 sky130_fd_sc_hd__inv_1_1.A phi2 0.00236f
C142 sky130_fd_sc_hd__dlymetal6s6s_1_3.A a_3724_36936# 3.61e-19
C143 a_3121_38050# a_3227_38050# 0.319f
C144 sky130_fd_sc_hd__dlymetal6s6s_1_5.A a_3724_36936# 0.00883f
C145 sky130_fd_sc_hd__inv_1_2.Y a_2024_38050# 3.29e-20
C146 a_3121_38050# a_3227_37506# 4.65e-19
C147 a_3227_38050# a_3121_37506# 4.65e-19
C148 sky130_fd_sc_hd__inv_1_2.Y a_2024_37506# 0.0647f
C149 a_3121_37506# a_3227_37506# 0.319f
C150 mimbot1 a_1794_38050# 4.99e-20
C151 vcm a_2590_38050# 5.29e-19
C152 mimbot1 a_1798_37826# 4.07e-20
C153 vcm a_2590_37506# 3.01e-20
C154 mimbot1 a_3724_38568# 0.00827f
C155 VDD a_4324_38050# 0.204f
C156 VDD sky130_fd_sc_hd__inv_1_2.Y 0.646f
C157 mimtop2 a_3172_38568# 4.98e-20
C158 VDD a_4324_37506# 0.204f
C159 a_3121_37506# phi2_n 4.05e-19
C160 sky130_fd_sc_hd__inv_1_2.Y sky130_fd_sc_hd__nand2_1_0.Y 6.3e-20
C161 sky130_fd_sc_hd__inv_1_2.Y sky130_fd_sc_hd__nand2_1_1.Y 0.345f
C162 sky130_fd_sc_hd__inv_1_0.A a_3510_38050# 4.96e-19
C163 a_4041_38050# sky130_fd_sc_hd__inv_1_3.A 2.42e-19
C164 mimbot1 a_2024_38050# -1.06e-34
C165 sky130_fd_sc_hd__inv_1_2.Y a_3172_36936# 2.28e-19
C166 mimtop2 phi2 0.0684f
C167 a_4041_37506# sky130_fd_sc_hd__inv_1_3.A 0.00232f
C168 mimbot1 a_2024_37506# 5.1e-36
C169 phi1 a_2944_38050# 5.55e-20
C170 sky130_fd_sc_hd__inv_1_2.A a_4430_38050# 1.97e-19
C171 a_4430_37506# sky130_fd_sc_hd__inv_1_1.A 0.157f
C172 sky130_fd_sc_hd__inv_1_3.Y a_2024_38050# 0.0542f
C173 a_3724_36936# phi2 0.224f
C174 VDD mimbot1 1.7f
C175 a_3121_38050# a_3510_38050# 7.09e-19
C176 mimbot1 sky130_fd_sc_hd__nand2_1_0.Y 0.0025f
C177 a_3227_38050# a_3404_38050# 0.16f
C178 sky130_fd_sc_hd__inv_1_2.Y a_2307_38050# 3.29e-20
C179 mimbot1 sky130_fd_sc_hd__nand2_1_1.Y 9.9e-19
C180 VDD sky130_fd_sc_hd__inv_1_3.Y 0.905f
C181 phi1 sky130_fd_sc_hd__dlymetal6s6s_1_2.A 2e-20
C182 sky130_fd_sc_hd__inv_1_2.Y a_2307_37506# 0.0525f
C183 phi1 phi1_n 0.785f
C184 sky130_fd_sc_hd__inv_1_0.A a_4041_38050# 0.00325f
C185 sky130_fd_sc_hd__inv_1_3.Y sky130_fd_sc_hd__nand2_1_0.Y 0.282f
C186 mimbot1 a_3172_36936# 0.00895f
C187 a_3121_37506# a_3510_37506# 7.09e-19
C188 a_3227_37506# a_3404_37506# 0.16f
C189 sky130_fd_sc_hd__inv_1_3.Y sky130_fd_sc_hd__nand2_1_1.Y 7.86e-19
C190 sky130_fd_sc_hd__inv_1_3.Y a_3172_36936# 0.215f
C191 VDD a_1794_38050# 2.98e-21
C192 phi1_n clk 0.00371f
C193 sky130_fd_sc_hd__nand2_1_0.Y a_1794_38050# 0.00989f
C194 VDD a_1798_37826# 2.25e-20
C195 VDD a_3724_38568# 0.368f
C196 a_2024_38050# a_2024_37506# 0.0126f
C197 a_4324_38050# sky130_fd_sc_hd__inv_1_3.A 1.37e-19
C198 sky130_fd_sc_hd__nand2_1_1.Y a_1798_37826# 0.00984f
C199 mimbot1 a_2307_38050# 0.00381f
C200 a_4324_37506# sky130_fd_sc_hd__inv_1_3.A 8.38e-19
C201 mimbot1 a_2307_37506# 0.00194f
C202 phi1 a_3227_38050# 2.7e-20
C203 sky130_fd_sc_hd__inv_1_3.Y a_2307_38050# 0.0535f
C204 VDD a_2024_38050# 0.25f
C205 VDD a_2024_37506# 0.254f
C206 sky130_fd_sc_hd__nand2_1_0.Y a_2024_38050# 0.284f
C207 a_2024_38050# sky130_fd_sc_hd__nand2_1_1.Y 4.65e-19
C208 sky130_fd_sc_hd__nand2_1_0.Y a_2024_37506# 4.65e-19
C209 a_2944_37506# phi2 1.22e-19
C210 sky130_fd_sc_hd__nand2_1_1.Y a_2024_37506# 0.311f
C211 a_3404_38050# a_3510_38050# 0.322f
C212 sky130_fd_sc_hd__inv_1_2.Y a_2590_38050# 3.29e-20
C213 a_3172_38568# phi1_n 0.225f
C214 a_3510_38050# a_3404_37506# 4.65e-19
C215 a_3404_38050# a_3510_37506# 4.65e-19
C216 sky130_fd_sc_hd__inv_1_2.Y a_2590_37506# 0.0533f
C217 sky130_fd_sc_hd__inv_1_0.A a_4324_38050# 0.0126f
C218 mimbot1 sky130_fd_sc_hd__inv_1_3.A 2.31e-19
C219 phi1 mimtop1 0.0818f
C220 a_3404_37506# a_3510_37506# 0.322f
C221 sky130_fd_sc_hd__inv_1_2.Y sky130_fd_sc_hd__inv_1_0.A 0.0271f
C222 VDD sky130_fd_sc_hd__nand2_1_0.Y 0.384f
C223 VDD sky130_fd_sc_hd__nand2_1_1.Y 0.445f
C224 sky130_fd_sc_hd__inv_1_3.Y sky130_fd_sc_hd__inv_1_3.A 0.221f
C225 VDD a_3172_36936# 0.415f
C226 sky130_fd_sc_hd__nand2_1_0.Y sky130_fd_sc_hd__nand2_1_1.Y 0.0138f
C227 sky130_fd_sc_hd__dlymetal6s6s_1_4.A phi2 4.55e-19
C228 mimtop1 clk 0.175f
C229 a_2201_38050# a_2201_37506# 0.0137f
C230 vcm phi1 0.213f
C231 mimbot1 a_2590_38050# 0.0178f
C232 sky130_fd_sc_hd__inv_1_1.A a_3724_36936# 0.00335f
C233 a_3172_38568# a_3227_38050# 0.00449f
C234 sky130_fd_sc_hd__inv_1_2.Y a_3121_38050# 0.00905f
C235 mimbot1 a_2590_37506# 0.0174f
C236 a_3724_38568# sky130_fd_sc_hd__inv_1_3.A 3.37e-20
C237 sky130_fd_sc_hd__inv_1_2.A a_3724_36936# 3.37e-20
C238 phi1 a_3510_38050# 6.18e-20
C239 a_3172_38568# a_3227_37506# 1.02e-19
C240 sky130_fd_sc_hd__inv_1_2.Y a_3121_37506# 0.0474f
C241 sky130_fd_sc_hd__inv_1_3.Y a_2590_38050# 0.0541f
C242 vcm clk 0.00409f
C243 mimtop2 a_2201_38050# 0.00635f
C244 VDD a_2307_38050# 0.169f
C245 mimtop2 a_2201_37506# 0.00804f
C246 VDD a_2307_37506# 0.173f
C247 sky130_fd_sc_hd__nand2_1_0.Y a_2307_38050# 0.00235f
C248 sky130_fd_sc_hd__inv_1_0.A sky130_fd_sc_hd__inv_1_3.Y 0.0075f
C249 a_3227_37506# phi2 4.88e-20
C250 sky130_fd_sc_hd__nand2_1_1.Y a_2307_37506# 0.00182f
C251 a_3172_38568# phi2_n 1.3e-20
C252 a_3510_38050# sky130_fd_sc_hd__dlymetal6s6s_1_3.A 0.153f
C253 mimtop1 a_3172_38568# 1.48e-20
C254 a_3510_37506# sky130_fd_sc_hd__dlymetal6s6s_1_5.A 0.153f
C255 a_3864_38050# a_4041_38050# 0.16f
C256 mimbot1 a_3121_38050# 0.0137f
C257 phi2_n phi2 0.647f
C258 a_3724_38568# sky130_fd_sc_hd__inv_1_0.A 0.00343f
C259 mimbot1 a_3121_37506# 0.0122f
C260 VDD sky130_fd_sc_hd__inv_1_3.A 0.449f
C261 mimtop1 phi2 0.0506f
C262 sky130_fd_sc_hd__inv_1_3.Y a_3121_38050# 0.0595f
C263 a_3864_37506# a_4041_37506# 0.16f
C264 sky130_fd_sc_hd__inv_1_3.Y a_3121_37506# 0.00644f
C265 a_2201_38050# a_2484_38050# 0.0145f
C266 vcm a_3172_38568# 0.00117f
C267 a_2307_38050# a_2307_37506# 0.0126f
C268 a_2201_37506# a_2484_37506# 0.0145f
C269 sky130_fd_sc_hd__dlymetal6s6s_1_3.A a_4041_38050# 0.0146f
C270 sky130_fd_sc_hd__inv_1_2.Y a_3404_38050# 0.0267f
C271 vcm phi2 0.0265f
C272 sky130_fd_sc_hd__inv_1_2.Y a_3404_37506# 0.0413f
C273 sky130_fd_sc_hd__dlymetal6s6s_1_5.A a_4041_37506# 0.0146f
C274 a_2944_37506# sky130_fd_sc_hd__inv_1_1.A 6.92e-21
C275 mimtop2 a_2484_38050# 0.0392f
C276 VDD a_2590_38050# 0.173f
C277 sky130_fd_sc_hd__nand2_1_0.Y a_2590_38050# 5.61e-19
C278 VDD a_2590_37506# 0.179f
C279 mimtop2 a_2484_37506# 0.0419f
C280 VDD sky130_fd_sc_hd__inv_1_0.A 0.443f
C281 a_3510_37506# phi2 6.99e-20
C282 sky130_fd_sc_hd__nand2_1_1.Y a_2590_37506# 4.28e-19
C283 phi1_n sky130_fd_sc_hd__inv_1_4.Y 9.78e-20
C284 mimbot1 a_3404_38050# 0.0067f
C285 a_4041_38050# a_4147_38050# 0.319f
C286 sky130_fd_sc_hd__inv_1_2.Y a_3864_38050# 0.00426f
C287 mimbot1 a_3404_37506# 0.00549f
C288 a_4041_38050# a_4147_37506# 4.65e-19
C289 a_4147_38050# a_4041_37506# 4.65e-19
C290 sky130_fd_sc_hd__inv_1_2.Y a_3864_37506# 0.00146f
C291 sky130_fd_sc_hd__inv_1_3.Y a_3404_38050# 0.0607f
C292 phi1 sky130_fd_sc_hd__inv_1_2.Y 0.252f
C293 a_4041_37506# a_4147_37506# 0.319f
C294 VDD a_3121_38050# 0.195f
C295 sky130_fd_sc_hd__inv_1_3.Y a_3404_37506# 0.021f
C296 sky130_fd_sc_hd__nand2_1_0.Y a_3121_38050# 2.37e-19
C297 VDD a_3121_37506# 0.202f
C298 phi1_n a_2201_38050# 0.005f
C299 a_2484_38050# a_2484_37506# 0.0137f
C300 phi1_n a_2201_37506# 2.36e-19
C301 sky130_fd_sc_hd__inv_1_2.Y clk 2.81e-19
C302 sky130_fd_sc_hd__nand2_1_1.Y a_3121_37506# 2.65e-19
C303 a_3121_38050# a_3172_36936# 1.21e-19
C304 sky130_fd_sc_hd__inv_1_2.Y sky130_fd_sc_hd__dlymetal6s6s_1_3.A 0.00594f
C305 a_3121_37506# a_3172_36936# 0.00736f
C306 sky130_fd_sc_hd__inv_1_2.Y sky130_fd_sc_hd__dlymetal6s6s_1_5.A 0.003f
C307 a_3227_37506# sky130_fd_sc_hd__inv_1_1.A 1.31e-20
C308 mimtop2 sky130_fd_sc_hd__dlymetal6s6s_1_2.A 6.84e-19
C309 mimtop2 phi1_n 0.069f
C310 mimbot1 a_3864_38050# 0.00163f
C311 mimtop2 sky130_fd_sc_hd__dlymetal6s6s_1_4.A 4.9e-19
C312 phi1 mimbot1 0.0894f
C313 sky130_fd_sc_hd__inv_1_3.Y a_3864_38050# 0.00768f
C314 sky130_fd_sc_hd__inv_1_3.Y a_3864_37506# 0.0141f
C315 phi1 sky130_fd_sc_hd__inv_1_3.Y 1.81e-19
C316 sky130_fd_sc_hd__inv_1_1.A phi2_n 6.18e-21
C317 a_2484_38050# a_2944_38050# 7.12e-19
C318 mimtop1 sky130_fd_sc_hd__inv_1_4.Y 0.0294f
C319 mimbot1 clk 0.00965f
C320 a_2484_37506# a_2944_37506# 7.12e-19
C321 a_4041_38050# a_4430_38050# 7.09e-19
C322 a_4147_38050# a_4324_38050# 0.16f
C323 mimbot1 sky130_fd_sc_hd__dlymetal6s6s_1_3.A 0.00195f
C324 sky130_fd_sc_hd__inv_1_2.Y a_4147_38050# 0.00169f
C325 clk sky130_fd_sc_hd__inv_1_3.Y 0.0518f
C326 a_3172_38568# sky130_fd_sc_hd__inv_1_2.Y 0.207f
C327 sky130_fd_sc_hd__inv_1_2.Y a_4147_37506# 3.38e-19
C328 sky130_fd_sc_hd__inv_1_3.Y sky130_fd_sc_hd__dlymetal6s6s_1_3.A 0.0176f
C329 a_3724_38568# a_3864_38050# 0.00416f
C330 a_4041_37506# a_4430_37506# 7.09e-19
C331 a_4147_37506# a_4324_37506# 0.16f
C332 VDD a_3404_38050# 0.194f
C333 a_2201_38050# phi2_n 2.48e-19
C334 a_3724_38568# a_3864_37506# 1.92e-19
C335 sky130_fd_sc_hd__inv_1_3.Y sky130_fd_sc_hd__dlymetal6s6s_1_5.A 0.0282f
C336 vcm sky130_fd_sc_hd__inv_1_4.Y 0.00464f
C337 phi1 a_3724_38568# 0.221f
C338 VDD a_3404_37506# 0.202f
C339 a_2484_38050# sky130_fd_sc_hd__dlymetal6s6s_1_2.A 0.0135f
C340 sky130_fd_sc_hd__nand2_1_0.Y a_3404_38050# 1.52e-19
C341 a_2201_37506# phi2_n 0.00468f
C342 phi1_n a_2484_38050# 0.00489f
C343 sky130_fd_sc_hd__inv_1_2.Y phi2 2.22e-20
C344 mimtop1 a_2201_38050# 6.37e-19
C345 a_2590_38050# a_2590_37506# 0.0126f
C346 phi1_n a_2484_37506# 2.17e-19
C347 mimtop1 a_2201_37506# 3.04e-20
C348 sky130_fd_sc_hd__nand2_1_1.Y a_3404_37506# 1.74e-19
C349 a_3404_38050# a_3172_36936# 1.86e-19
C350 a_2484_37506# sky130_fd_sc_hd__dlymetal6s6s_1_4.A 0.0135f
C351 a_3404_37506# a_3172_36936# 0.00358f
C352 a_2944_38050# a_2944_37506# 0.0126f
C353 mimtop2 phi2_n 0.0664f
C354 a_3724_38568# sky130_fd_sc_hd__dlymetal6s6s_1_3.A 0.00883f
C355 a_3510_37506# sky130_fd_sc_hd__inv_1_1.A 3.81e-19
C356 mimbot1 a_4147_38050# 0.0029f
C357 a_3724_38568# sky130_fd_sc_hd__dlymetal6s6s_1_5.A 3.61e-19
C358 mimbot1 a_3172_38568# 0.028f
C359 mimtop1 mimtop2 0.0211f
C360 vcm a_2201_38050# 0.037f
C361 vcm a_2201_37506# 0.0366f
C362 sky130_fd_sc_hd__inv_1_3.Y a_4147_38050# 0.00255f
C363 a_3724_36936# phi2_n 8.34e-21
C364 a_3172_38568# sky130_fd_sc_hd__inv_1_3.Y 6.64e-20
C365 VDD a_3864_38050# 0.205f
C366 sky130_fd_sc_hd__inv_1_3.Y a_4147_37506# 0.00493f
C367 VDD a_3864_37506# 0.205f
C368 sky130_fd_sc_hd__dlymetal6s6s_1_2.A a_2944_38050# 0.35f
C369 phi1_n a_2944_38050# 6.38e-19
C370 VDD phi1 0.54f
C371 mimbot1 phi2 0.126f
C372 a_2944_38050# sky130_fd_sc_hd__dlymetal6s6s_1_4.A 4.65e-19
C373 sky130_fd_sc_hd__dlymetal6s6s_1_2.A a_2944_37506# 4.65e-19
C374 phi1_n a_2944_37506# 7.06e-20
C375 sky130_fd_sc_hd__inv_1_0.A a_3121_38050# 1.91e-20
C376 sky130_fd_sc_hd__dlymetal6s6s_1_4.A a_2944_37506# 0.35f
C377 vcm mimtop2 0.108p
C378 sky130_fd_sc_hd__inv_1_3.Y phi2 0.248f
C379 a_4324_38050# a_4430_38050# 0.322f
C380 sky130_fd_sc_hd__inv_1_2.Y a_4430_38050# 7.49e-19
C381 phi1 a_3172_36936# 1.79e-21
C382 a_4430_38050# a_4324_37506# 4.65e-19
C383 a_4324_38050# a_4430_37506# 4.65e-19
C384 VDD clk 0.337f
C385 sky130_fd_sc_hd__inv_1_2.Y a_4430_37506# 1.72e-19
C386 sky130_fd_sc_hd__inv_1_2.A a_4041_38050# 0.00231f
C387 a_4324_37506# a_4430_37506# 0.322f
C388 a_4041_37506# sky130_fd_sc_hd__inv_1_1.A 0.00325f
C389 clk sky130_fd_sc_hd__nand2_1_0.Y 0.126f
C390 a_3172_38568# a_3724_38568# 6.05e-19
C391 VDD sky130_fd_sc_hd__dlymetal6s6s_1_3.A 0.245f
C392 a_2484_38050# phi2_n 2.56e-19
C393 sky130_fd_sc_hd__inv_1_2.A a_4041_37506# 2.42e-19
C394 clk sky130_fd_sc_hd__nand2_1_1.Y 0.00909f
C395 VDD sky130_fd_sc_hd__dlymetal6s6s_1_5.A 0.245f
C396 phi1_n sky130_fd_sc_hd__dlymetal6s6s_1_2.A 0.00235f
C397 a_2484_37506# phi2_n 0.00678f
C398 mimtop1 a_2484_38050# 5.19e-19
C399 sky130_fd_sc_hd__dlymetal6s6s_1_2.A sky130_fd_sc_hd__dlymetal6s6s_1_4.A 0.0137f
C400 phi1_n sky130_fd_sc_hd__dlymetal6s6s_1_4.A 3.28e-19
C401 a_3724_38568# phi2 4.02e-20
C402 a_3121_38050# a_3121_37506# 0.0137f
C403 mimbot1 a_4430_38050# 3.99e-19
C404 vcm a_2484_38050# 0.00609f
C405 vcm a_2484_37506# 0.00547f
C406 sky130_fd_sc_hd__inv_1_3.Y a_4430_38050# 0.00134f
C407 VDD a_4147_38050# 0.17f
C408 a_2944_38050# phi2_n 7.18e-20
C409 VDD a_3172_38568# 0.417f
C410 sky130_fd_sc_hd__inv_1_3.Y a_4430_37506# 0.00242f
C411 sky130_fd_sc_hd__dlymetal6s6s_1_2.A a_3227_38050# 6.53e-19
C412 VDD a_4147_37506# 0.17f
C413 phi1_n a_3227_38050# 0.0012f
C414 a_2944_37506# phi2_n 5.64e-19
C415 sky130_fd_sc_hd__inv_1_0.A a_3404_38050# 1.2e-19
C416 sky130_fd_sc_hd__dlymetal6s6s_1_4.A a_3227_37506# 6.53e-19
C417 VDD phi2 0.611f
C418 a_3172_38568# a_3172_36936# 0.00101f
C419 sky130_fd_sc_hd__inv_1_2.Y sky130_fd_sc_hd__inv_1_4.Y 0.0521f
C420 a_4041_37506# a_3724_36936# 7.18e-20
C421 sky130_fd_sc_hd__inv_1_2.Y sky130_fd_sc_hd__inv_1_1.A 8.25e-20
C422 sky130_fd_sc_hd__inv_1_2.A a_4324_38050# 8.38e-19
C423 a_4324_37506# sky130_fd_sc_hd__inv_1_1.A 0.0126f
C424 sky130_fd_sc_hd__inv_1_2.Y sky130_fd_sc_hd__inv_1_2.A 0.22f
C425 sky130_fd_sc_hd__dlymetal6s6s_1_2.A phi2_n 3.23e-19
C426 phi1_n phi2_n 0.00349f
C427 sky130_fd_sc_hd__inv_1_2.A a_4324_37506# 1.37e-19
C428 a_3172_36936# phi2 0.103f
C429 sky130_fd_sc_hd__dlymetal6s6s_1_4.A phi2_n 0.00187f
C430 mimtop1 phi1_n 0.0657f
C431 a_3121_38050# a_3404_38050# 0.0145f
C432 sky130_fd_sc_hd__inv_1_2.Y a_2201_38050# 1.32e-20
C433 a_3227_38050# a_3227_37506# 0.0126f
C434 sky130_fd_sc_hd__inv_1_2.Y a_2201_37506# 0.0467f
C435 sky130_fd_sc_hd__inv_1_0.A a_3864_38050# 0.00215f
C436 a_3121_37506# a_3404_37506# 0.0145f
C437 mimbot1 sky130_fd_sc_hd__inv_1_4.Y 0.00182f
C438 phi1 sky130_fd_sc_hd__inv_1_0.A 0.00225f
C439 vcm phi1_n 0.24f
C440 mimbot1 sky130_fd_sc_hd__inv_1_2.A 0.00628f
C441 VDD a_4430_38050# 0.178f
C442 mimtop2 sky130_fd_sc_hd__inv_1_2.Y 0.08f
C443 sky130_fd_sc_hd__inv_1_3.Y sky130_fd_sc_hd__inv_1_1.A 0.0364f
C444 VDD a_4430_37506# 0.178f
C445 a_3227_37506# phi2_n 0.0012f
C446 sky130_fd_sc_hd__inv_1_0.A sky130_fd_sc_hd__dlymetal6s6s_1_3.A 0.00211f
C447 a_4147_38050# sky130_fd_sc_hd__inv_1_3.A 3.52e-21
C448 mimbot1 a_2201_38050# 0.00172f
C449 a_4147_37506# sky130_fd_sc_hd__inv_1_3.A 0.0111f
C450 mimbot1 a_2201_37506# 8.06e-19
C451 sky130_fd_sc_hd__inv_1_3.Y a_2201_38050# 0.0599f
C452 sky130_fd_sc_hd__inv_1_3.A phi2 0.00305f
C453 mimtop1 phi2_n 0.08f
C454 a_3724_38568# sky130_fd_sc_hd__inv_1_2.A 0.19f
C455 mimbot1 mimtop2 1.61f
C456 sky130_fd_sc_hd__inv_1_2.Y a_2484_38050# 1.32e-20
C457 mimtop2 sky130_fd_sc_hd__inv_1_3.Y 0.0818f
C458 a_3404_38050# a_3404_37506# 0.0137f
C459 sky130_fd_sc_hd__inv_1_2.Y a_2484_37506# 0.0447f
C460 sky130_fd_sc_hd__inv_1_0.A a_4147_38050# 0.00429f
C461 mimbot1 a_3724_36936# 7.45e-19
C462 a_3172_38568# sky130_fd_sc_hd__inv_1_0.A 1.89e-19
C463 vcm phi2_n 0.031f
C464 sky130_fd_sc_hd__inv_1_3.Y a_3724_36936# 0.174f
C465 vcm mimtop1 0.11p
C466 VDD sky130_fd_sc_hd__inv_1_4.Y 0.303f
C467 sky130_fd_sc_hd__nand2_1_0.Y sky130_fd_sc_hd__inv_1_4.Y 7.79e-19
C468 VDD sky130_fd_sc_hd__inv_1_1.A 0.441f
C469 a_2024_38050# a_2201_38050# 0.16f
C470 VDD sky130_fd_sc_hd__inv_1_2.A 0.414f
C471 sky130_fd_sc_hd__inv_1_4.Y sky130_fd_sc_hd__nand2_1_1.Y 0.0702f
C472 a_2024_37506# a_2201_37506# 0.16f
C473 mimbot1 a_2484_38050# 0.002f
C474 a_3404_38050# a_3864_38050# 7.12e-19
C475 a_4430_37506# sky130_fd_sc_hd__inv_1_3.A 2.14e-19
C476 sky130_fd_sc_hd__inv_1_1.A a_3172_36936# 1.58e-20
C477 a_3172_38568# a_3121_38050# 0.00736f
C478 sky130_fd_sc_hd__inv_1_2.Y a_2944_38050# 0.00629f
C479 mimbot1 a_2484_37506# 0.00109f
C480 phi1 a_3404_38050# 2.92e-21
C481 a_3724_38568# a_3724_36936# 0.00102f
C482 a_3172_38568# a_3121_37506# 1.21e-19
C483 sky130_fd_sc_hd__inv_1_2.Y a_2944_37506# 0.0631f
C484 sky130_fd_sc_hd__inv_1_3.Y a_2484_38050# 0.0584f
C485 a_3404_37506# a_3864_37506# 7.12e-19
C486 VDD a_2201_38050# 0.195f
C487 sky130_fd_sc_hd__nand2_1_0.Y a_2201_38050# 0.0195f
C488 VDD a_2201_37506# 0.203f
C489 sky130_fd_sc_hd__nand2_1_1.Y a_2201_37506# 0.019f
C490 a_3404_38050# sky130_fd_sc_hd__dlymetal6s6s_1_3.A 0.0135f
C491 sky130_fd_sc_hd__inv_1_2.Y sky130_fd_sc_hd__dlymetal6s6s_1_2.A 0.00223f
C492 sky130_fd_sc_hd__inv_1_2.Y phi1_n 0.0113f
C493 a_3510_38050# a_3510_37506# 0.0126f
C494 VDD mimtop2 1.66f
C495 sky130_fd_sc_hd__inv_1_2.Y sky130_fd_sc_hd__dlymetal6s6s_1_4.A 0.0667f
C496 sky130_fd_sc_hd__inv_1_0.A a_4430_38050# 0.157f
C497 a_3404_37506# sky130_fd_sc_hd__dlymetal6s6s_1_5.A 0.0135f
C498 mimtop2 sky130_fd_sc_hd__nand2_1_0.Y 6.91e-19
C499 mimbot1 a_2944_38050# 0.0295f
C500 mimtop2 sky130_fd_sc_hd__nand2_1_1.Y 5.76e-19
C501 mimbot1 a_2944_37506# 0.0244f
C502 a_3864_38050# a_3864_37506# 0.0126f
C503 VDD a_3724_36936# 0.367f
C504 mimtop2 a_3172_36936# 4.27e-20
C505 sky130_fd_sc_hd__inv_1_3.Y a_2944_38050# 0.0576f
C506 sky130_fd_sc_hd__inv_1_3.Y a_2944_37506# 0.00384f
C507 a_2201_38050# a_2307_38050# 0.319f
C508 a_2201_38050# a_2307_37506# 4.65e-19
C509 a_2307_38050# a_2201_37506# 4.65e-19
C510 a_3172_36936# a_3724_36936# 6.05e-19
C511 a_2201_37506# a_2307_37506# 0.319f
C512 mimbot1 sky130_fd_sc_hd__dlymetal6s6s_1_2.A 0.0575f
C513 sky130_fd_sc_hd__dlymetal6s6s_1_3.A a_3864_38050# 0.35f
C514 mimbot1 phi1_n 0.147f
C515 sky130_fd_sc_hd__inv_1_1.A sky130_fd_sc_hd__inv_1_3.A 0.0988f
C516 a_3172_38568# a_3404_38050# 0.00358f
C517 sky130_fd_sc_hd__inv_1_2.Y a_3227_38050# 0.0138f
C518 mimbot1 sky130_fd_sc_hd__dlymetal6s6s_1_4.A 0.0578f
C519 sky130_fd_sc_hd__dlymetal6s6s_1_3.A a_3864_37506# 4.65e-19
C520 a_3864_38050# sky130_fd_sc_hd__dlymetal6s6s_1_5.A 4.65e-19
C521 sky130_fd_sc_hd__inv_1_2.A sky130_fd_sc_hd__inv_1_3.A 4.25e-19
C522 phi1 sky130_fd_sc_hd__dlymetal6s6s_1_3.A 7.55e-19
C523 sky130_fd_sc_hd__inv_1_2.Y a_3227_37506# 0.0548f
C524 a_3172_38568# a_3404_37506# 1.86e-19
C525 sky130_fd_sc_hd__inv_1_3.Y sky130_fd_sc_hd__dlymetal6s6s_1_2.A 0.0884f
C526 phi1_n sky130_fd_sc_hd__inv_1_3.Y 0.0056f
C527 sky130_fd_sc_hd__dlymetal6s6s_1_5.A a_3864_37506# 0.35f
C528 VDD a_2484_38050# 0.194f
C529 mimtop2 a_2307_38050# 0.0175f
C530 sky130_fd_sc_hd__inv_1_3.Y sky130_fd_sc_hd__dlymetal6s6s_1_4.A 0.00188f
C531 mimtop2 a_2307_37506# 0.0188f
C532 sky130_fd_sc_hd__nand2_1_0.Y a_2484_38050# 0.00112f
C533 VDD a_2484_37506# 0.201f
C534 a_3404_37506# phi2 4.84e-21
C535 sky130_fd_sc_hd__nand2_1_1.Y a_2484_37506# 0.00117f
C536 sky130_fd_sc_hd__inv_1_2.Y phi2_n 1.74e-19
C537 sky130_fd_sc_hd__dlymetal6s6s_1_3.A sky130_fd_sc_hd__dlymetal6s6s_1_5.A 0.0137f
C538 mimtop1 sky130_fd_sc_hd__inv_1_2.Y 0.00212f
C539 phi2 VSS 1.47f
C540 phi2_n VSS 0.811f
C541 sky130_fd_sc_hd__inv_1_3.A VSS 0.532f
C542 a_3724_36936# VSS 0.501f
C543 a_3172_36936# VSS 0.548f
C544 sky130_fd_sc_hd__inv_1_1.A VSS 0.589f
C545 a_1798_37826# VSS 0.00195f
C546 a_4430_37506# VSS 0.241f
C547 a_4324_37506# VSS 0.228f
C548 a_4147_37506# VSS 0.217f
C549 a_4041_37506# VSS 0.22f
C550 a_3864_37506# VSS 0.248f
C551 sky130_fd_sc_hd__dlymetal6s6s_1_5.A VSS 0.258f
C552 a_3510_37506# VSS 0.222f
C553 a_3404_37506# VSS 0.202f
C554 a_3227_37506# VSS 0.201f
C555 a_3121_37506# VSS 0.202f
C556 a_2944_37506# VSS 0.231f
C557 sky130_fd_sc_hd__dlymetal6s6s_1_4.A VSS 0.24f
C558 a_2590_37506# VSS 0.209f
C559 a_2484_37506# VSS 0.201f
C560 a_2307_37506# VSS 0.202f
C561 a_2201_37506# VSS 0.203f
C562 a_2024_37506# VSS 0.229f
C563 sky130_fd_sc_hd__nand2_1_1.Y VSS 0.325f
C564 sky130_fd_sc_hd__inv_1_4.Y VSS 0.337f
C565 a_1794_38050# VSS 0.00199f
C566 a_4430_38050# VSS 0.241f
C567 a_4324_38050# VSS 0.228f
C568 a_4147_38050# VSS 0.217f
C569 a_4041_38050# VSS 0.22f
C570 a_3864_38050# VSS 0.248f
C571 sky130_fd_sc_hd__dlymetal6s6s_1_3.A VSS 0.258f
C572 a_3510_38050# VSS 0.225f
C573 a_3404_38050# VSS 0.212f
C574 a_3227_38050# VSS 0.213f
C575 a_3121_38050# VSS 0.213f
C576 a_2944_38050# VSS 0.245f
C577 sky130_fd_sc_hd__dlymetal6s6s_1_2.A VSS 0.256f
C578 a_2590_38050# VSS 0.222f
C579 a_2484_38050# VSS 0.212f
C580 a_2307_38050# VSS 0.215f
C581 a_2201_38050# VSS 0.214f
C582 a_2024_38050# VSS 0.291f
C583 sky130_fd_sc_hd__nand2_1_0.Y VSS 0.468f
C584 sky130_fd_sc_hd__inv_1_3.Y VSS 1.15f
C585 clk VSS 0.729f
C586 phi1_n VSS 1.08f
C587 sky130_fd_sc_hd__inv_1_0.A VSS 0.588f
C588 sky130_fd_sc_hd__inv_1_2.A VSS 0.497f
C589 a_3724_38568# VSS 0.501f
C590 sky130_fd_sc_hd__inv_1_2.Y VSS 1.53f
C591 a_3172_38568# VSS 0.546f
C592 mimtop2 VSS 1.31p
C593 mimtop1 VSS 0.104p
C594 mimbot1 VSS 0.956p
C595 phi1 VSS 1.81f
C596 vcm VSS 23.8p
C597 VDD VSS 1.18p
C598 mimbot1.n0 VSS 0.0407f
C599 mimbot1.t47 VSS 0.00487f
C600 mimbot1.t46 VSS 0.00487f
C601 mimbot1.n1 VSS 0.0329f
C602 mimbot1.t43 VSS 0.00487f
C603 mimbot1.t42 VSS 0.00487f
C604 mimbot1.n2 VSS 0.00974f
C605 mimbot1.n3 VSS 0.231f
C606 mimbot1.n4 VSS 0.801f
C607 mimbot1.n5 VSS 0.0222f
C608 mimbot1.n6 VSS 0.0222f
C609 mimbot1.n7 VSS 0.0108f
C610 mimbot1.n8 VSS 0.00572f
C611 mimbot1.t45 VSS 0.0192f
C612 mimbot1.t44 VSS 0.0188f
C613 mimbot1.t1 VSS 0.0248f
C614 mimbot1.n9 VSS 0.0914f
C615 mimbot1.n10 VSS 0.0734f
C616 mimbot1.t0 VSS 0.00491f
C617 mimbot1.n11 VSS 0.0425f
C618 mimbot1.n12 VSS 0.066f
C619 mimbot1.n13 VSS 0.0312f
C620 mimbot1.n14 VSS 0.00948f
C621 mimbot1.n15 VSS 0.00663f
C622 mimbot1.n16 VSS 0.00642f
C623 mimbot1.n18 VSS 0.0108f
C624 mimbot1.n19 VSS 0.00572f
C625 mimbot1.n20 VSS 0.0066f
C626 mimbot1.n21 VSS 0.00642f
C627 mimbot1.n22 VSS 0.0136f
C628 mimbot1.n23 VSS 0.0274f
C629 mimbot1.n24 VSS 0.594f
C630 mimbot1.n25 VSS 0.612f
C631 mimbot1.n26 VSS 0.702f
C632 mimbot1.n27 VSS 0.0868f
C633 mimbot1.n28 VSS 0.265f
C634 mimbot1.t11 VSS 16.9f
C635 mimbot1.n29 VSS 5.28f
C636 mimbot1.n30 VSS 0.764f
C637 mimbot1.n31 VSS 0.265f
C638 mimbot1.t35 VSS 16.9f
C639 mimbot1.n32 VSS 5.28f
C640 mimbot1.n33 VSS 0.764f
C641 mimbot1.n34 VSS 0.265f
C642 mimbot1.t21 VSS 16.9f
C643 mimbot1.n35 VSS 5.28f
C644 mimbot1.n36 VSS 0.764f
C645 mimbot1.n37 VSS 0.132f
C646 mimbot1.n38 VSS 0.393f
C647 mimbot1.n39 VSS 0.265f
C648 mimbot1.t30 VSS 16.9f
C649 mimbot1.n40 VSS 5.28f
C650 mimbot1.n41 VSS 0.764f
C651 mimbot1.n42 VSS 5.28f
C652 mimbot1.t4 VSS 16.9f
C653 mimbot1.n43 VSS 0.265f
C654 mimbot1.n44 VSS 0.764f
C655 mimbot1.n45 VSS 5.28f
C656 mimbot1.t9 VSS 16.9f
C657 mimbot1.n46 VSS 0.265f
C658 mimbot1.n47 VSS 0.764f
C659 mimbot1.n48 VSS 5.28f
C660 mimbot1.t24 VSS 16.9f
C661 mimbot1.n49 VSS 0.265f
C662 mimbot1.n50 VSS 0.764f
C663 mimbot1.n51 VSS 4.27f
C664 mimbot1.n52 VSS 0.362f
C665 mimbot1.n53 VSS 2.64f
C666 mimbot1.n54 VSS 0.139f
C667 mimbot1.n55 VSS 0.265f
C668 mimbot1.n56 VSS 2.64f
C669 mimbot1.n57 VSS 0.139f
C670 mimbot1.n58 VSS 0.265f
C671 mimbot1.n59 VSS 2.64f
C672 mimbot1.n60 VSS 0.139f
C673 mimbot1.n61 VSS 0.265f
C674 mimbot1.n62 VSS 0.855f
C675 mimbot1.n63 VSS 0.0458f
C676 mimbot1.n64 VSS 0.265f
C677 mimbot1.n65 VSS 0.139f
C678 mimbot1.n66 VSS 0.193f
C679 mimbot1.n67 VSS 0.354f
C680 mimbot1.n68 VSS 0.264f
C681 mimbot1.n69 VSS 0.311f
C682 mimbot1.n70 VSS 0.127f
C683 mimbot1.n71 VSS 0.126f
C684 mimbot1.n72 VSS 0.124f
C685 mimbot1.n73 VSS 0.646f
C686 mimbot1.n74 VSS 0.134f
C687 mimbot1.n75 VSS 0.393f
C688 mimbot1.n76 VSS 0.264f
C689 mimbot1.n77 VSS 0.126f
C690 mimbot1.n78 VSS 2.74f
C691 mimbot1.n79 VSS 0.393f
C692 mimbot1.n80 VSS 0.134f
C693 mimbot1.n81 VSS 0.193f
C694 mimbot1.n82 VSS 0.124f
C695 mimbot1.n83 VSS 0.646f
C696 mimbot1.n84 VSS 0.311f
C697 mimbot1.n85 VSS 0.127f
C698 mimbot1.n86 VSS 0.354f
C699 mimbot1.n87 VSS 2.64f
C700 mimbot1.n88 VSS 0.265f
C701 mimbot1.n89 VSS 0.139f
C702 mimbot1.n90 VSS 0.193f
C703 mimbot1.n91 VSS 0.354f
C704 mimbot1.n92 VSS 0.264f
C705 mimbot1.n93 VSS 0.311f
C706 mimbot1.n94 VSS 0.127f
C707 mimbot1.n95 VSS 0.126f
C708 mimbot1.n96 VSS 0.124f
C709 mimbot1.n97 VSS 0.646f
C710 mimbot1.n98 VSS 0.134f
C711 mimbot1.n99 VSS 0.393f
C712 mimbot1.n100 VSS 0.264f
C713 mimbot1.n101 VSS 0.126f
C714 mimbot1.n102 VSS 0.393f
C715 mimbot1.n103 VSS 0.134f
C716 mimbot1.n104 VSS 0.193f
C717 mimbot1.n105 VSS 0.124f
C718 mimbot1.n106 VSS 0.646f
C719 mimbot1.n107 VSS 0.311f
C720 mimbot1.n108 VSS 0.127f
C721 mimbot1.n109 VSS 0.354f
C722 mimbot1.n110 VSS 2.64f
C723 mimbot1.n111 VSS 0.265f
C724 mimbot1.n112 VSS 0.139f
C725 mimbot1.n113 VSS 0.193f
C726 mimbot1.n114 VSS 0.354f
C727 mimbot1.n115 VSS 0.264f
C728 mimbot1.n116 VSS 0.311f
C729 mimbot1.n117 VSS 0.127f
C730 mimbot1.n118 VSS 0.126f
C731 mimbot1.n119 VSS 0.124f
C732 mimbot1.n120 VSS 0.646f
C733 mimbot1.n121 VSS 0.134f
C734 mimbot1.n122 VSS 0.393f
C735 mimbot1.n123 VSS 0.264f
C736 mimbot1.n124 VSS 0.126f
C737 mimbot1.n125 VSS 0.393f
C738 mimbot1.n126 VSS 0.134f
C739 mimbot1.n127 VSS 0.193f
C740 mimbot1.n128 VSS 0.124f
C741 mimbot1.n129 VSS 0.646f
C742 mimbot1.n130 VSS 0.311f
C743 mimbot1.n131 VSS 0.127f
C744 mimbot1.n132 VSS 0.354f
C745 mimbot1.n133 VSS 2.64f
C746 mimbot1.n134 VSS 0.265f
C747 mimbot1.n135 VSS 0.139f
C748 mimbot1.n136 VSS 0.188f
C749 mimbot1.n137 VSS 0.233f
C750 mimbot1.n138 VSS 0.134f
C751 mimbot1.n139 VSS 0.393f
C752 mimbot1.n140 VSS 0.264f
C753 mimbot1.n141 VSS 0.126f
C754 mimbot1.n142 VSS 0.393f
C755 mimbot1.n143 VSS 0.134f
C756 mimbot1.n144 VSS 0.193f
C757 mimbot1.n145 VSS 0.124f
C758 mimbot1.n146 VSS 0.646f
C759 mimbot1.n147 VSS 0.311f
C760 mimbot1.n148 VSS 0.127f
C761 mimbot1.n149 VSS 0.354f
C762 mimbot1.n150 VSS 2.64f
C763 mimbot1.n151 VSS 85.8f
C764 mimbot1.t40 VSS 16.9f
C765 mimbot1.n152 VSS 0.37f
C766 mimbot1.n153 VSS 0.193f
C767 mimbot1.n154 VSS 0.139f
C768 mimbot1.n155 VSS 0.646f
C769 mimbot1.n156 VSS 0.311f
C770 mimbot1.n157 VSS 0.264f
C771 mimbot1.t7 VSS 16.9f
C772 mimbot1.n158 VSS 0.218f
C773 mimbot1.n159 VSS 0.258f
C774 mimbot1.n160 VSS 0.386f
C775 mimbot1.n161 VSS 0.702f
C776 mimbot1.n162 VSS 0.764f
C777 mimbot1.n163 VSS 0.27f
C778 mimbot1.n164 VSS 0.27f
C779 mimbot1.n165 VSS 0.148f
C780 mimbot1.n166 VSS 0.248f
C781 mimbot1.n167 VSS 0.28f
C782 mimbot1.n168 VSS 0.644f
C783 mimbot1.t2 VSS 16.9f
C784 mimbot1.n169 VSS 0.28f
C785 mimbot1.n170 VSS 0.258f
C786 mimbot1.n171 VSS 0.702f
C787 mimbot1.n172 VSS 0.764f
C788 mimbot1.n173 VSS 0.27f
C789 mimbot1.n174 VSS 0.386f
C790 mimbot1.n175 VSS 0.27f
C791 mimbot1.n176 VSS 0.148f
C792 mimbot1.n177 VSS 0.248f
C793 mimbot1.n178 VSS 0.218f
C794 mimbot1.n179 VSS 0.644f
C795 mimbot1.n180 VSS 0.28f
C796 mimbot1.n181 VSS 0.258f
C797 mimbot1.n182 VSS 0.702f
C798 mimbot1.n183 VSS 0.764f
C799 mimbot1.n184 VSS 0.27f
C800 mimbot1.n185 VSS 0.386f
C801 mimbot1.n186 VSS 0.27f
C802 mimbot1.n187 VSS 0.148f
C803 mimbot1.n188 VSS 0.248f
C804 mimbot1.n189 VSS 0.218f
C805 mimbot1.n190 VSS 0.644f
C806 mimbot1.t16 VSS 16.9f
C807 mimbot1.t37 VSS 16.9f
C808 mimbot1.n191 VSS 0.218f
C809 mimbot1.n192 VSS 0.258f
C810 mimbot1.n193 VSS 0.386f
C811 mimbot1.n194 VSS 0.702f
C812 mimbot1.n195 VSS 0.764f
C813 mimbot1.n196 VSS 0.27f
C814 mimbot1.n197 VSS 0.27f
C815 mimbot1.n198 VSS 0.148f
C816 mimbot1.n199 VSS 0.248f
C817 mimbot1.n200 VSS 0.28f
C818 mimbot1.n201 VSS 0.644f
C819 mimbot1.n202 VSS 0.218f
C820 mimbot1.n203 VSS 0.258f
C821 mimbot1.n204 VSS 0.386f
C822 mimbot1.n205 VSS 0.702f
C823 mimbot1.n206 VSS 0.764f
C824 mimbot1.n207 VSS 0.27f
C825 mimbot1.n208 VSS 0.27f
C826 mimbot1.n209 VSS 0.148f
C827 mimbot1.n210 VSS 0.248f
C828 mimbot1.n211 VSS 0.28f
C829 mimbot1.n212 VSS 0.644f
C830 mimbot1.t27 VSS 16.9f
C831 mimbot1.n213 VSS 0.28f
C832 mimbot1.n214 VSS 0.258f
C833 mimbot1.n215 VSS 0.702f
C834 mimbot1.n216 VSS 0.764f
C835 mimbot1.n217 VSS 0.27f
C836 mimbot1.n218 VSS 0.386f
C837 mimbot1.n219 VSS 0.27f
C838 mimbot1.n220 VSS 0.148f
C839 mimbot1.n221 VSS 0.248f
C840 mimbot1.n222 VSS 0.218f
C841 mimbot1.n223 VSS 0.644f
C842 mimbot1.t12 VSS 16.9f
C843 mimbot1.n224 VSS 0.205f
C844 mimbot1.n225 VSS 0.193f
C845 mimbot1.n226 VSS 0.37f
C846 mimbot1.n227 VSS 0.139f
C847 mimbot1.n228 VSS 0.134f
C848 mimbot1.n229 VSS 0.646f
C849 mimbot1.n230 VSS 0.311f
C850 mimbot1.n231 VSS 0.264f
C851 mimbot1.n232 VSS 0.284f
C852 mimbot1.t31 VSS 16.9f
C853 mimbot1.n233 VSS 0.218f
C854 mimbot1.n234 VSS 0.258f
C855 mimbot1.n235 VSS 0.386f
C856 mimbot1.n236 VSS 0.702f
C857 mimbot1.n237 VSS 0.764f
C858 mimbot1.n238 VSS 0.27f
C859 mimbot1.n239 VSS 0.27f
C860 mimbot1.n240 VSS 0.148f
C861 mimbot1.n241 VSS 0.248f
C862 mimbot1.n242 VSS 0.28f
C863 mimbot1.n243 VSS 0.644f
C864 mimbot1.n244 VSS 0.265f
C865 mimbot1.n245 VSS 5.28f
C866 mimbot1.n246 VSS 0.764f
C867 mimbot1.n247 VSS 0.265f
C868 mimbot1.n248 VSS 0.393f
C869 mimbot1.n249 VSS 0.132f
C870 mimbot1.n250 VSS 5.28f
C871 mimbot1.n251 VSS 0.764f
C872 mimbot1.n252 VSS 0.265f
C873 mimbot1.n253 VSS 5.28f
C874 mimbot1.n254 VSS 0.764f
C875 mimbot1.n255 VSS 0.265f
C876 mimbot1.n256 VSS 0.764f
C877 mimbot1.n257 VSS 5.28f
C878 mimbot1.n258 VSS 0.265f
C879 mimbot1.n259 VSS 5.28f
C880 mimbot1.n260 VSS 0.764f
C881 mimbot1.n261 VSS 0.265f
C882 mimbot1.n262 VSS 0.764f
C883 mimbot1.n263 VSS 5.28f
C884 mimbot1.n264 VSS 0.265f
C885 mimbot1.n265 VSS 5.28f
C886 mimbot1.n266 VSS 0.764f
C887 mimbot1.n267 VSS 0.132f
C888 mimbot1.n268 VSS 0.393f
C889 mimbot1.n269 VSS 0.218f
C890 mimbot1.n270 VSS 0.258f
C891 mimbot1.n271 VSS 0.386f
C892 mimbot1.n272 VSS 0.702f
C893 mimbot1.n273 VSS 0.764f
C894 mimbot1.n274 VSS 0.27f
C895 mimbot1.n275 VSS 0.27f
C896 mimbot1.n276 VSS 0.148f
C897 mimbot1.n277 VSS 0.248f
C898 mimbot1.n278 VSS 0.28f
C899 mimbot1.n279 VSS 0.644f
C900 mimbot1.t5 VSS 16.9f
C901 mimbot1.n280 VSS 0.28f
C902 mimbot1.n281 VSS 0.258f
C903 mimbot1.n282 VSS 0.702f
C904 mimbot1.n283 VSS 0.764f
C905 mimbot1.n284 VSS 0.27f
C906 mimbot1.n285 VSS 0.386f
C907 mimbot1.n286 VSS 0.27f
C908 mimbot1.n287 VSS 0.148f
C909 mimbot1.n288 VSS 0.248f
C910 mimbot1.n289 VSS 0.218f
C911 mimbot1.n290 VSS 0.644f
C912 mimbot1.n291 VSS 0.28f
C913 mimbot1.n292 VSS 0.258f
C914 mimbot1.n293 VSS 0.702f
C915 mimbot1.n294 VSS 0.764f
C916 mimbot1.n295 VSS 0.27f
C917 mimbot1.n296 VSS 0.386f
C918 mimbot1.n297 VSS 0.27f
C919 mimbot1.n298 VSS 0.148f
C920 mimbot1.n299 VSS 0.248f
C921 mimbot1.n300 VSS 0.218f
C922 mimbot1.n301 VSS 0.644f
C923 mimbot1.t18 VSS 16.9f
C924 mimbot1.n302 VSS 0.205f
C925 mimbot1.n303 VSS 0.193f
C926 mimbot1.n304 VSS 0.37f
C927 mimbot1.n305 VSS 0.139f
C928 mimbot1.n306 VSS 0.134f
C929 mimbot1.n307 VSS 0.646f
C930 mimbot1.n308 VSS 0.311f
C931 mimbot1.n309 VSS 0.264f
C932 mimbot1.n310 VSS 0.284f
C933 mimbot1.t33 VSS 16.9f
C934 mimbot1.n311 VSS 0.28f
C935 mimbot1.n312 VSS 0.258f
C936 mimbot1.n313 VSS 0.702f
C937 mimbot1.n314 VSS 0.764f
C938 mimbot1.n315 VSS 0.27f
C939 mimbot1.n316 VSS 0.386f
C940 mimbot1.n317 VSS 0.27f
C941 mimbot1.n318 VSS 0.148f
C942 mimbot1.n319 VSS 0.248f
C943 mimbot1.n320 VSS 0.218f
C944 mimbot1.n321 VSS 0.644f
C945 mimbot1.t22 VSS 16.9f
C946 mimbot1.n322 VSS 0.218f
C947 mimbot1.n323 VSS 0.258f
C948 mimbot1.n324 VSS 0.386f
C949 mimbot1.n325 VSS 0.702f
C950 mimbot1.n326 VSS 0.764f
C951 mimbot1.n327 VSS 0.27f
C952 mimbot1.n328 VSS 0.27f
C953 mimbot1.n329 VSS 0.148f
C954 mimbot1.n330 VSS 0.248f
C955 mimbot1.n331 VSS 0.28f
C956 mimbot1.n332 VSS 0.644f
C957 mimbot1.t10 VSS 16.9f
C958 mimbot1.n333 VSS 0.28f
C959 mimbot1.n334 VSS 0.258f
C960 mimbot1.n335 VSS 0.702f
C961 mimbot1.n336 VSS 0.764f
C962 mimbot1.n337 VSS 0.27f
C963 mimbot1.n338 VSS 0.386f
C964 mimbot1.n339 VSS 0.27f
C965 mimbot1.n340 VSS 0.148f
C966 mimbot1.n341 VSS 0.248f
C967 mimbot1.n342 VSS 0.218f
C968 mimbot1.n343 VSS 0.644f
C969 mimbot1.t38 VSS 16.9f
C970 mimbot1.t14 VSS 16.9f
C971 mimbot1.n344 VSS 0.265f
C972 mimbot1.n345 VSS 5.28f
C973 mimbot1.n346 VSS 0.764f
C974 mimbot1.n347 VSS 0.265f
C975 mimbot1.n348 VSS 0.393f
C976 mimbot1.n349 VSS 0.132f
C977 mimbot1.n350 VSS 5.28f
C978 mimbot1.n351 VSS 0.764f
C979 mimbot1.n352 VSS 5.28f
C980 mimbot1.n353 VSS 4.27f
C981 mimbot1.n354 VSS 0.393f
C982 mimbot1.n355 VSS 0.132f
C983 mimbot1.n356 VSS 0.764f
C984 mimbot1.n357 VSS 5.28f
C985 mimbot1.n358 VSS 0.265f
C986 mimbot1.n359 VSS 0.764f
C987 mimbot1.n360 VSS 0.265f
C988 mimbot1.n361 VSS 5.28f
C989 mimbot1.n362 VSS 5.28f
C990 mimbot1.n363 VSS 0.764f
C991 mimbot1.n364 VSS 0.265f
C992 mimbot1.n365 VSS 0.764f
C993 mimbot1.n366 VSS 0.265f
C994 mimbot1.n367 VSS 0.265f
C995 mimbot1.n368 VSS 0.764f
C996 mimbot1.n369 VSS 0.702f
C997 mimbot1.n370 VSS 0.386f
C998 mimbot1.n371 VSS 0.764f
C999 mimbot1.n372 VSS 0.218f
C1000 mimbot1.n373 VSS 0.258f
C1001 mimbot1.n374 VSS 0.386f
C1002 mimbot1.n375 VSS 0.702f
C1003 mimbot1.n376 VSS 0.764f
C1004 mimbot1.n377 VSS 0.27f
C1005 mimbot1.n378 VSS 0.27f
C1006 mimbot1.n379 VSS 0.148f
C1007 mimbot1.n380 VSS 0.248f
C1008 mimbot1.n381 VSS 0.28f
C1009 mimbot1.n382 VSS 0.644f
C1010 mimbot1.n383 VSS 0.205f
C1011 mimbot1.n384 VSS 0.193f
C1012 mimbot1.n385 VSS 0.37f
C1013 mimbot1.n386 VSS 0.139f
C1014 mimbot1.n387 VSS 0.134f
C1015 mimbot1.n388 VSS 0.646f
C1016 mimbot1.n389 VSS 0.311f
C1017 mimbot1.n390 VSS 0.264f
C1018 mimbot1.n391 VSS 0.284f
C1019 mimbot1.t32 VSS 16.9f
C1020 mimbot1.n392 VSS 0.218f
C1021 mimbot1.n393 VSS 0.258f
C1022 mimbot1.n394 VSS 0.386f
C1023 mimbot1.n395 VSS 0.702f
C1024 mimbot1.n396 VSS 0.764f
C1025 mimbot1.n397 VSS 0.27f
C1026 mimbot1.n398 VSS 0.27f
C1027 mimbot1.n399 VSS 0.148f
C1028 mimbot1.n400 VSS 0.248f
C1029 mimbot1.n401 VSS 0.28f
C1030 mimbot1.n402 VSS 0.644f
C1031 mimbot1.n403 VSS 0.218f
C1032 mimbot1.n404 VSS 0.258f
C1033 mimbot1.n405 VSS 0.702f
C1034 mimbot1.n406 VSS 0.27f
C1035 mimbot1.n407 VSS 0.27f
C1036 mimbot1.n408 VSS 0.148f
C1037 mimbot1.n409 VSS 0.248f
C1038 mimbot1.n410 VSS 0.28f
C1039 mimbot1.n411 VSS 0.644f
C1040 mimbot1.n412 VSS 0.218f
C1041 mimbot1.n413 VSS 0.258f
C1042 mimbot1.n414 VSS 0.386f
C1043 mimbot1.n415 VSS 0.764f
C1044 mimbot1.n416 VSS 0.27f
C1045 mimbot1.n417 VSS 0.27f
C1046 mimbot1.n418 VSS 0.148f
C1047 mimbot1.n419 VSS 0.248f
C1048 mimbot1.n420 VSS 0.28f
C1049 mimbot1.n421 VSS 0.644f
C1050 mimbot1.t8 VSS 16.9f
C1051 mimbot1.t19 VSS 16.9f
C1052 mimbot1.t36 VSS 16.9f
C1053 mimbot1.n422 VSS 0.264f
C1054 mimbot1.n423 VSS 0.37f
C1055 mimbot1.n424 VSS 0.134f
C1056 mimbot1.n425 VSS 0.311f
C1057 mimbot1.n426 VSS 0.139f
C1058 mimbot1.n427 VSS 0.646f
C1059 mimbot1.n428 VSS 0.193f
C1060 mimbot1.n429 VSS 0.205f
C1061 mimbot1.n430 VSS 0.288f
C1062 mimbot1.t23 VSS 16.9f
C1063 mimbot1.n431 VSS 0.218f
C1064 mimbot1.n432 VSS 0.258f
C1065 mimbot1.n433 VSS 0.386f
C1066 mimbot1.n434 VSS 0.702f
C1067 mimbot1.n435 VSS 0.764f
C1068 mimbot1.n436 VSS 0.27f
C1069 mimbot1.n437 VSS 0.27f
C1070 mimbot1.n438 VSS 0.148f
C1071 mimbot1.n439 VSS 0.248f
C1072 mimbot1.n440 VSS 0.28f
C1073 mimbot1.n441 VSS 0.644f
C1074 mimbot1.n442 VSS 0.218f
C1075 mimbot1.n443 VSS 0.258f
C1076 mimbot1.n444 VSS 0.386f
C1077 mimbot1.n445 VSS 0.702f
C1078 mimbot1.n446 VSS 0.764f
C1079 mimbot1.n447 VSS 0.27f
C1080 mimbot1.n448 VSS 0.27f
C1081 mimbot1.n449 VSS 0.148f
C1082 mimbot1.n450 VSS 0.248f
C1083 mimbot1.n451 VSS 0.28f
C1084 mimbot1.n452 VSS 0.644f
C1085 mimbot1.n453 VSS 0.28f
C1086 mimbot1.n454 VSS 0.258f
C1087 mimbot1.n455 VSS 0.702f
C1088 mimbot1.n456 VSS 0.764f
C1089 mimbot1.n457 VSS 0.27f
C1090 mimbot1.n458 VSS 0.386f
C1091 mimbot1.n459 VSS 0.27f
C1092 mimbot1.n460 VSS 0.148f
C1093 mimbot1.n461 VSS 0.248f
C1094 mimbot1.n462 VSS 0.218f
C1095 mimbot1.n463 VSS 0.644f
C1096 mimbot1.t28 VSS 16.9f
C1097 mimbot1.t39 VSS 16.9f
C1098 mimbot1.n464 VSS 0.265f
C1099 mimbot1.n465 VSS 5.28f
C1100 mimbot1.n466 VSS 0.764f
C1101 mimbot1.n467 VSS 0.265f
C1102 mimbot1.n468 VSS 0.393f
C1103 mimbot1.n469 VSS 0.132f
C1104 mimbot1.n470 VSS 5.28f
C1105 mimbot1.n471 VSS 0.764f
C1106 mimbot1.n472 VSS 0.265f
C1107 mimbot1.n473 VSS 5.28f
C1108 mimbot1.n474 VSS 0.764f
C1109 mimbot1.n475 VSS 0.132f
C1110 mimbot1.n476 VSS 0.393f
C1111 mimbot1.n477 VSS 5.28f
C1112 mimbot1.n478 VSS 5.28f
C1113 mimbot1.n479 VSS 0.764f
C1114 mimbot1.n480 VSS 5.28f
C1115 mimbot1.n481 VSS 5.28f
C1116 mimbot1.n482 VSS 0.764f
C1117 mimbot1.n483 VSS 4.27f
C1118 mimbot1.n484 VSS 0.265f
C1119 mimbot1.n485 VSS 0.764f
C1120 mimbot1.n486 VSS 0.265f
C1121 mimbot1.n487 VSS 0.265f
C1122 mimbot1.n488 VSS 0.764f
C1123 mimbot1.n489 VSS 0.28f
C1124 mimbot1.n490 VSS 0.702f
C1125 mimbot1.n491 VSS 0.258f
C1126 mimbot1.t26 VSS 16.9f
C1127 mimbot1.n492 VSS 0.28f
C1128 mimbot1.n493 VSS 0.258f
C1129 mimbot1.n494 VSS 0.702f
C1130 mimbot1.n495 VSS 0.764f
C1131 mimbot1.n496 VSS 0.27f
C1132 mimbot1.n497 VSS 0.386f
C1133 mimbot1.n498 VSS 0.27f
C1134 mimbot1.n499 VSS 0.148f
C1135 mimbot1.n500 VSS 0.248f
C1136 mimbot1.n501 VSS 0.218f
C1137 mimbot1.n502 VSS 0.644f
C1138 mimbot1.n503 VSS 0.28f
C1139 mimbot1.n504 VSS 0.258f
C1140 mimbot1.n505 VSS 0.702f
C1141 mimbot1.n506 VSS 0.764f
C1142 mimbot1.n507 VSS 0.27f
C1143 mimbot1.n508 VSS 0.386f
C1144 mimbot1.n509 VSS 0.27f
C1145 mimbot1.n510 VSS 0.148f
C1146 mimbot1.n511 VSS 0.248f
C1147 mimbot1.n512 VSS 0.218f
C1148 mimbot1.n513 VSS 0.644f
C1149 mimbot1.t41 VSS 16.9f
C1150 mimbot1.n514 VSS 0.205f
C1151 mimbot1.n515 VSS 0.193f
C1152 mimbot1.n516 VSS 0.37f
C1153 mimbot1.n517 VSS 0.139f
C1154 mimbot1.n518 VSS 0.134f
C1155 mimbot1.n519 VSS 0.646f
C1156 mimbot1.n520 VSS 0.311f
C1157 mimbot1.n521 VSS 0.264f
C1158 mimbot1.n522 VSS 0.284f
C1159 mimbot1.t15 VSS 16.9f
C1160 mimbot1.n523 VSS 0.28f
C1161 mimbot1.n524 VSS 0.258f
C1162 mimbot1.n525 VSS 0.702f
C1163 mimbot1.n526 VSS 0.764f
C1164 mimbot1.n527 VSS 0.27f
C1165 mimbot1.n528 VSS 0.386f
C1166 mimbot1.n529 VSS 0.27f
C1167 mimbot1.n530 VSS 0.148f
C1168 mimbot1.n531 VSS 0.248f
C1169 mimbot1.n532 VSS 0.218f
C1170 mimbot1.n533 VSS 0.644f
C1171 mimbot1.t3 VSS 16.9f
C1172 mimbot1.t29 VSS 16.9f
C1173 mimbot1.n534 VSS 0.218f
C1174 mimbot1.n535 VSS 0.258f
C1175 mimbot1.n536 VSS 0.386f
C1176 mimbot1.n537 VSS 0.702f
C1177 mimbot1.n538 VSS 0.764f
C1178 mimbot1.n539 VSS 0.27f
C1179 mimbot1.n540 VSS 0.27f
C1180 mimbot1.n541 VSS 0.148f
C1181 mimbot1.n542 VSS 0.248f
C1182 mimbot1.n543 VSS 0.28f
C1183 mimbot1.n544 VSS 0.644f
C1184 mimbot1.n545 VSS 0.218f
C1185 mimbot1.n546 VSS 0.258f
C1186 mimbot1.n547 VSS 0.386f
C1187 mimbot1.n548 VSS 0.702f
C1188 mimbot1.n549 VSS 0.764f
C1189 mimbot1.n550 VSS 0.27f
C1190 mimbot1.n551 VSS 0.27f
C1191 mimbot1.n552 VSS 0.148f
C1192 mimbot1.n553 VSS 0.248f
C1193 mimbot1.n554 VSS 0.28f
C1194 mimbot1.n555 VSS 0.644f
C1195 mimbot1.t20 VSS 16.9f
C1196 mimbot1.n556 VSS 0.218f
C1197 mimbot1.n557 VSS 0.258f
C1198 mimbot1.n558 VSS 0.386f
C1199 mimbot1.n559 VSS 0.702f
C1200 mimbot1.n560 VSS 0.764f
C1201 mimbot1.n561 VSS 0.27f
C1202 mimbot1.n562 VSS 0.27f
C1203 mimbot1.n563 VSS 0.148f
C1204 mimbot1.n564 VSS 0.248f
C1205 mimbot1.n565 VSS 0.28f
C1206 mimbot1.n566 VSS 0.644f
C1207 mimbot1.n567 VSS 0.205f
C1208 mimbot1.n568 VSS 0.139f
C1209 mimbot1.n569 VSS 0.193f
C1210 mimbot1.n570 VSS 0.134f
C1211 mimbot1.n571 VSS 0.646f
C1212 mimbot1.n572 VSS 0.37f
C1213 mimbot1.n573 VSS 0.311f
C1214 mimbot1.n574 VSS 0.264f
C1215 mimbot1.n575 VSS 0.288f
C1216 mimbot1.t34 VSS 16.9f
C1217 mimbot1.n576 VSS 0.265f
C1218 mimbot1.n577 VSS 2.64f
C1219 mimbot1.n578 VSS 0.139f
C1220 mimbot1.n579 VSS 0.265f
C1221 mimbot1.n580 VSS 0.393f
C1222 mimbot1.n581 VSS 0.0987f
C1223 mimbot1.n582 VSS 0.393f
C1224 mimbot1.n583 VSS 0.185f
C1225 mimbot1.n584 VSS 0.134f
C1226 mimbot1.n585 VSS 0.238f
C1227 mimbot1.n586 VSS 0.134f
C1228 mimbot1.n587 VSS 0.132f
C1229 mimbot1.n588 VSS 0.193f
C1230 mimbot1.n589 VSS 0.354f
C1231 mimbot1.n590 VSS 0.264f
C1232 mimbot1.n591 VSS 0.311f
C1233 mimbot1.n592 VSS 0.127f
C1234 mimbot1.n593 VSS 0.126f
C1235 mimbot1.n594 VSS 0.124f
C1236 mimbot1.n595 VSS 0.646f
C1237 mimbot1.n596 VSS 0.134f
C1238 mimbot1.n597 VSS 0.393f
C1239 mimbot1.n598 VSS 2.64f
C1240 mimbot1.n599 VSS 0.139f
C1241 mimbot1.n600 VSS 0.265f
C1242 mimbot1.n601 VSS 0.265f
C1243 mimbot1.n602 VSS 0.139f
C1244 mimbot1.n603 VSS 0.157f
C1245 mimbot1.n604 VSS 0.393f
C1246 mimbot1.n605 VSS 0.134f
C1247 mimbot1.n606 VSS 0.316f
C1248 mimbot1.n607 VSS 0.324f
C1249 mimbot1.n608 VSS 2.74f
C1250 mimbot1.n609 VSS 0.264f
C1251 mimbot1.n610 VSS 0.126f
C1252 mimbot1.n611 VSS 0.393f
C1253 mimbot1.n612 VSS 0.134f
C1254 mimbot1.n613 VSS 0.193f
C1255 mimbot1.n614 VSS 0.124f
C1256 mimbot1.n615 VSS 0.646f
C1257 mimbot1.n616 VSS 0.311f
C1258 mimbot1.n617 VSS 0.127f
C1259 mimbot1.n618 VSS 0.354f
C1260 mimbot1.n619 VSS 2.64f
C1261 mimbot1.n620 VSS 0.139f
C1262 mimbot1.n621 VSS 0.265f
C1263 mimbot1.n622 VSS 0.193f
C1264 mimbot1.n623 VSS 0.354f
C1265 mimbot1.n624 VSS 0.264f
C1266 mimbot1.n625 VSS 0.311f
C1267 mimbot1.n626 VSS 0.127f
C1268 mimbot1.n627 VSS 0.126f
C1269 mimbot1.n628 VSS 0.124f
C1270 mimbot1.n629 VSS 0.646f
C1271 mimbot1.n630 VSS 0.134f
C1272 mimbot1.n631 VSS 0.393f
C1273 mimbot1.n632 VSS 2.64f
C1274 mimbot1.n633 VSS 0.139f
C1275 mimbot1.n634 VSS 0.265f
C1276 mimbot1.n635 VSS 0.193f
C1277 mimbot1.n636 VSS 0.354f
C1278 mimbot1.n637 VSS 0.264f
C1279 mimbot1.n638 VSS 0.311f
C1280 mimbot1.n639 VSS 0.127f
C1281 mimbot1.n640 VSS 0.126f
C1282 mimbot1.n641 VSS 0.124f
C1283 mimbot1.n642 VSS 0.646f
C1284 mimbot1.n643 VSS 0.134f
C1285 mimbot1.n644 VSS 0.393f
C1286 mimbot1.n645 VSS 2.64f
C1287 mimbot1.n646 VSS 0.139f
C1288 mimbot1.n647 VSS 0.265f
C1289 mimbot1.n648 VSS 0.264f
C1290 mimbot1.n649 VSS 0.126f
C1291 mimbot1.n650 VSS 0.393f
C1292 mimbot1.n651 VSS 0.134f
C1293 mimbot1.n652 VSS 0.193f
C1294 mimbot1.n653 VSS 0.124f
C1295 mimbot1.n654 VSS 0.646f
C1296 mimbot1.n655 VSS 0.311f
C1297 mimbot1.n656 VSS 0.127f
C1298 mimbot1.n657 VSS 0.354f
C1299 mimbot1.n658 VSS 2.64f
C1300 mimbot1.n659 VSS 0.139f
C1301 mimbot1.n660 VSS 0.264f
C1302 mimbot1.n661 VSS 0.126f
C1303 mimbot1.n662 VSS 0.393f
C1304 mimbot1.n663 VSS 0.134f
C1305 mimbot1.n664 VSS 0.193f
C1306 mimbot1.n665 VSS 0.124f
C1307 mimbot1.n666 VSS 0.646f
C1308 mimbot1.n667 VSS 0.311f
C1309 mimbot1.n668 VSS 0.127f
C1310 mimbot1.n669 VSS 0.354f
C1311 mimbot1.n670 VSS 0.193f
C1312 mimbot1.n671 VSS 0.354f
C1313 mimbot1.n672 VSS 0.264f
C1314 mimbot1.n673 VSS 0.311f
C1315 mimbot1.n674 VSS 0.127f
C1316 mimbot1.n675 VSS 0.126f
C1317 mimbot1.n676 VSS 0.124f
C1318 mimbot1.n677 VSS 0.646f
C1319 mimbot1.n678 VSS 0.134f
C1320 mimbot1.n679 VSS 0.393f
C1321 mimbot1.n680 VSS 2.64f
C1322 mimbot1.n681 VSS 84.6f
C1323 mimbot1.t6 VSS 16.9f
C1324 mimbot1.n682 VSS 92.7f
C1325 mimbot1.n683 VSS 0.644f
C1326 mimbot1.n684 VSS 0.218f
C1327 mimbot1.n685 VSS 0.764f
C1328 mimbot1.n686 VSS 0.27f
C1329 mimbot1.n687 VSS 0.386f
C1330 mimbot1.n688 VSS 0.248f
C1331 mimbot1.n689 VSS 0.148f
C1332 mimbot1.n690 VSS 0.27f
C1333 mimbot1.n691 VSS 0.265f
C1334 mimbot1.n692 VSS 84.6f
C1335 mimbot1.t13 VSS 16.9f
C1336 mimbot1.n693 VSS 92.7f
C1337 mimbot1.n694 VSS 5.28f
C1338 mimbot1.n695 VSS 84.6f
C1339 mimbot1.t25 VSS 16.9f
C1340 mimbot1.n696 VSS 92.7f
C1341 mimbot1.n697 VSS 0.139f
C1342 mimbot1.n698 VSS 0.311f
C1343 mimbot1.n699 VSS 0.264f
C1344 mimbot1.n700 VSS 0.288f
C1345 mimbot1.n701 VSS 0.205f
C1346 mimbot1.n702 VSS 0.134f
C1347 mimbot1.n703 VSS 0.193f
C1348 mimbot1.n704 VSS 0.646f
C1349 mimbot1.n705 VSS 0.37f
C1350 mimbot1.n706 VSS 0.386f
C1351 mimbot1.n707 VSS 0.702f
C1352 mimbot1.n708 VSS 0.218f
C1353 mimbot1.n709 VSS 0.258f
C1354 mimbot1.n710 VSS 0.27f
C1355 mimbot1.n711 VSS 0.644f
C1356 mimbot1.n712 VSS 0.28f
C1357 mimbot1.n713 VSS 0.248f
C1358 mimbot1.n714 VSS 0.148f
C1359 mimbot1.n715 VSS 0.27f
C1360 mimbot1.n716 VSS 0.764f
C1361 mimbot1.n717 VSS 4.27f
C1362 mimbot1.n718 VSS 84.6f
C1363 mimbot1.t17 VSS 16.9f
C1364 mimbot1.n719 VSS 92.7f
C1365 mimbot1.n720 VSS 0.288f
C1366 mimbot1.n721 VSS 0.205f
C1367 mimbot1.n722 VSS 0.132f
C1368 mimbot1.n723 VSS 84.6f
C1369 mimbot1.n724 VSS 0.672f
C1370 mimbot1.n725 VSS 3.19f
C1371 mimtop1.t28 VSS 15.7f
C1372 mimtop1.t42 VSS 15.7f
C1373 mimtop1.n0 VSS 8.84f
C1374 mimtop1.t32 VSS 15.7f
C1375 mimtop1.n1 VSS 8.84f
C1376 mimtop1.t18 VSS 15.7f
C1377 mimtop1.t35 VSS 15.7f
C1378 mimtop1.n2 VSS 8.84f
C1379 mimtop1.t24 VSS 15.7f
C1380 mimtop1.n3 VSS 8.84f
C1381 mimtop1.t11 VSS 15.7f
C1382 mimtop1.t21 VSS 15.7f
C1383 mimtop1.n4 VSS 8.84f
C1384 mimtop1.t10 VSS 15.7f
C1385 mimtop1.n5 VSS 8.84f
C1386 mimtop1.t36 VSS 15.7f
C1387 mimtop1.t8 VSS 15.7f
C1388 mimtop1.t46 VSS 15.7f
C1389 mimtop1.t20 VSS 15.7f
C1390 mimtop1.t15 VSS 15.7f
C1391 mimtop1.t43 VSS 15.7f
C1392 mimtop1.t29 VSS 15.7f
C1393 mimtop1.t34 VSS 15.7f
C1394 mimtop1.t23 VSS 15.7f
C1395 mimtop1.n6 VSS 98.1f
C1396 mimtop1.n7 VSS 8.84f
C1397 mimtop1.t26 VSS 15.7f
C1398 mimtop1.n8 VSS 8.84f
C1399 mimtop1.t13 VSS 15.7f
C1400 mimtop1.n9 VSS 8.84f
C1401 mimtop1.t41 VSS 15.7f
C1402 mimtop1.n10 VSS 8.84f
C1403 mimtop1.t30 VSS 15.7f
C1404 mimtop1.n11 VSS 8.84f
C1405 mimtop1.n12 VSS 8.84f
C1406 mimtop1.t17 VSS 15.7f
C1407 mimtop1.n13 VSS 70.7f
C1408 mimtop1.n14 VSS 8.84f
C1409 mimtop1.t39 VSS 15.7f
C1410 mimtop1.n15 VSS 8.84f
C1411 mimtop1.t27 VSS 15.7f
C1412 mimtop1.n16 VSS 8.84f
C1413 mimtop1.t16 VSS 15.7f
C1414 mimtop1.n17 VSS 8.84f
C1415 mimtop1.t44 VSS 15.7f
C1416 mimtop1.n18 VSS 8.84f
C1417 mimtop1.n19 VSS 8.84f
C1418 mimtop1.t31 VSS 15.7f
C1419 mimtop1.n20 VSS 70.7f
C1420 mimtop1.n21 VSS 8.84f
C1421 mimtop1.t47 VSS 15.7f
C1422 mimtop1.n22 VSS 8.84f
C1423 mimtop1.t33 VSS 15.7f
C1424 mimtop1.n23 VSS 8.84f
C1425 mimtop1.t22 VSS 15.7f
C1426 mimtop1.n24 VSS 8.84f
C1427 mimtop1.t12 VSS 15.7f
C1428 mimtop1.n25 VSS 8.84f
C1429 mimtop1.n26 VSS 8.84f
C1430 mimtop1.t37 VSS 15.7f
C1431 mimtop1.n27 VSS 70.7f
C1432 mimtop1.n28 VSS 8.84f
C1433 mimtop1.n29 VSS 8.84f
C1434 mimtop1.t40 VSS 15.7f
C1435 mimtop1.t38 VSS 15.7f
C1436 mimtop1.n30 VSS 8.84f
C1437 mimtop1.n31 VSS 8.82f
C1438 mimtop1.t9 VSS 15.7f
C1439 mimtop1.t25 VSS 15.7f
C1440 mimtop1.n32 VSS 8.84f
C1441 mimtop1.n33 VSS 8.84f
C1442 mimtop1.t14 VSS 15.7f
C1443 mimtop1.t19 VSS 15.7f
C1444 mimtop1.n34 VSS 8.84f
C1445 mimtop1.n35 VSS 8.84f
C1446 mimtop1.t45 VSS 15.7f
C1447 mimtop1.n36 VSS 97.9f
C1448 mimtop1.n37 VSS 1.8f
C1449 mimtop1.n38 VSS 1.55f
C1450 mimtop1.n39 VSS 0.00537f
C1451 mimtop1.n40 VSS 0.00473f
C1452 mimtop1.n41 VSS 7.24e-19
C1453 mimtop1.n42 VSS 0.00393f
C1454 mimtop1.n43 VSS 0.0035f
C1455 mimtop1.n44 VSS 0.0102f
C1456 mimtop1.t6 VSS 0.00192f
C1457 mimtop1.t7 VSS 0.00192f
C1458 mimtop1.n45 VSS 0.00384f
C1459 mimtop1.t3 VSS 0.00192f
C1460 mimtop1.t2 VSS 0.00192f
C1461 mimtop1.n46 VSS 0.0128f
C1462 mimtop1.n47 VSS 0.0113f
C1463 mimtop1.n48 VSS 0.042f
C1464 mimtop1.n49 VSS 0.00269f
C1465 mimtop1.n50 VSS 0.00251f
C1466 mimtop1.t4 VSS 0.00758f
C1467 mimtop1.t0 VSS 0.00947f
C1468 mimtop1.n51 VSS 0.0341f
C1469 mimtop1.t5 VSS 0.00755f
C1470 mimtop1.t1 VSS 0.00951f
C1471 mimtop1.n52 VSS 0.0177f
C1472 mimtop1.n53 VSS 0.137f
C1473 mimtop1.n54 VSS 0.0983f
C1474 mimtop1.n56 VSS 0.00454f
C1475 mimtop1.n57 VSS 0.00241f
C1476 mimtop1.n58 VSS 0.0271f
C1477 mimtop1.n59 VSS 0.00409f
C1478 mimtop1.n60 VSS 0.00269f
C1479 mimtop1.n61 VSS 0.00251f
C1480 mimtop1.n62 VSS 0.00454f
C1481 mimtop1.n63 VSS 0.00241f
C1482 mimtop1.n64 VSS 0.0201f
C1483 mimtop1.n65 VSS 0.159f
C1484 mimtop1.n66 VSS 0.0952f
C1485 mimtop1.n67 VSS 0.00918f
C1486 mimtop1.n68 VSS 0.00415f
C1487 mimtop1.n69 VSS 0.00351f
C1488 mimtop1.n71 VSS 0.00495f
C1489 mimtop1.n72 VSS 0.0304f
C1490 mimtop1.n73 VSS 0.0267f
C1491 mimtop1.n74 VSS 0.0067f
C1492 VDD.t84 VSS 0.0101f
C1493 VDD.t1 VSS 0.00281f
C1494 VDD.n0 VSS 0.00378f
C1495 VDD.n1 VSS 7.61e-19
C1496 VDD.t113 VSS 0.00281f
C1497 VDD.n2 VSS 9.53e-19
C1498 VDD.n3 VSS 0.00226f
C1499 VDD.t3 VSS 0.00122f
C1500 VDD.t91 VSS 3.55e-19
C1501 VDD.n4 VSS 0.0013f
C1502 VDD.n5 VSS 0.00167f
C1503 VDD.n6 VSS 0.00226f
C1504 VDD.t67 VSS 0.00122f
C1505 VDD.t93 VSS 3.55e-19
C1506 VDD.n7 VSS 0.0013f
C1507 VDD.n8 VSS 0.00155f
C1508 VDD.n9 VSS 0.00169f
C1509 VDD.n10 VSS 0.00404f
C1510 VDD.n11 VSS 0.00226f
C1511 VDD.t129 VSS 6.91e-19
C1512 VDD.t127 VSS 6.91e-19
C1513 VDD.n12 VSS 0.00158f
C1514 VDD.n13 VSS 0.0027f
C1515 VDD.n14 VSS 0.00204f
C1516 VDD.t133 VSS 0.00122f
C1517 VDD.t79 VSS 3.55e-19
C1518 VDD.n15 VSS 0.0013f
C1519 VDD.n16 VSS 0.00155f
C1520 VDD.n17 VSS 0.00169f
C1521 VDD.n18 VSS 3.48e-19
C1522 VDD.t109 VSS 6.91e-19
C1523 VDD.t103 VSS 6.91e-19
C1524 VDD.n19 VSS 0.00164f
C1525 VDD.n20 VSS 8.01e-19
C1526 VDD.n21 VSS 7.46e-19
C1527 VDD.t0 VSS 0.0114f
C1528 VDD.t88 VSS 0.00608f
C1529 VDD.t112 VSS 0.00297f
C1530 VDD.t98 VSS 0.0105f
C1531 VDD.t85 VSS 0.00688f
C1532 VDD.t12 VSS 0.0114f
C1533 VDD.t89 VSS 0.0136f
C1534 VDD.t90 VSS 0.013f
C1535 VDD.t2 VSS 0.0146f
C1536 VDD.t87 VSS 0.0136f
C1537 VDD.t92 VSS 0.0114f
C1538 VDD.t86 VSS 0.00683f
C1539 VDD.t66 VSS 0.0125f
C1540 VDD.t62 VSS 0.00818f
C1541 VDD.n22 VSS 0.00838f
C1542 VDD.t100 VSS 0.0122f
C1543 VDD.t130 VSS 0.0119f
C1544 VDD.t126 VSS 0.00775f
C1545 VDD.t4 VSS 0.00608f
C1546 VDD.t128 VSS 0.00688f
C1547 VDD.t40 VSS 0.00608f
C1548 VDD.t124 VSS 0.0097f
C1549 VDD.t140 VSS 0.00825f
C1550 VDD.t78 VSS 0.00862f
C1551 VDD.t132 VSS 0.0117f
C1552 VDD.t106 VSS 0.0109f
C1553 VDD.t102 VSS 0.0063f
C1554 VDD.t108 VSS 0.0076f
C1555 VDD.t138 VSS 0.00608f
C1556 VDD.t104 VSS 0.00688f
C1557 VDD.t52 VSS 0.00608f
C1558 VDD.t26 VSS 0.00572f
C1559 VDD.t82 VSS 0.0148f
C1560 VDD.t48 VSS 0.00695f
C1561 VDD.t28 VSS 0.00529f
C1562 VDD.t54 VSS 0.0148f
C1563 VDD.t50 VSS 0.00688f
C1564 VDD.t68 VSS 0.00521f
C1565 VDD.n23 VSS 0.013f
C1566 VDD.n24 VSS 7.74e-19
C1567 VDD.n25 VSS 3.7e-19
C1568 VDD.t51 VSS 0.0028f
C1569 VDD.n26 VSS 0.00289f
C1570 VDD.t69 VSS 0.00122f
C1571 VDD.t55 VSS 3.55e-19
C1572 VDD.n27 VSS 0.0013f
C1573 VDD.n28 VSS 0.00155f
C1574 VDD.n29 VSS 7e-19
C1575 VDD.n30 VSS 0.00205f
C1576 VDD.n31 VSS 0.00169f
C1577 VDD.n32 VSS 7.74e-19
C1578 VDD.n33 VSS 4.96e-19
C1579 VDD.t29 VSS 0.0028f
C1580 VDD.n34 VSS 0.00289f
C1581 VDD.t49 VSS 0.00122f
C1582 VDD.t83 VSS 3.55e-19
C1583 VDD.n35 VSS 0.0013f
C1584 VDD.n36 VSS 0.00167f
C1585 VDD.n37 VSS 5.22e-19
C1586 VDD.n38 VSS 0.00205f
C1587 VDD.n39 VSS 0.00169f
C1588 VDD.n40 VSS 7.86e-19
C1589 VDD.n41 VSS 8e-19
C1590 VDD.t27 VSS 6.91e-19
C1591 VDD.t105 VSS 6.91e-19
C1592 VDD.n42 VSS 0.00158f
C1593 VDD.t53 VSS 0.00122f
C1594 VDD.t139 VSS 3.55e-19
C1595 VDD.n43 VSS 0.00134f
C1596 VDD.n44 VSS 0.00202f
C1597 VDD.n45 VSS 0.002f
C1598 VDD.n46 VSS 4.22e-19
C1599 VDD.n47 VSS 0.00204f
C1600 VDD.n48 VSS 0.00226f
C1601 VDD.n49 VSS 0.00139f
C1602 VDD.n50 VSS 0.00353f
C1603 VDD.n51 VSS 4.44e-19
C1604 VDD.t107 VSS 0.00283f
C1605 VDD.n52 VSS 0.00441f
C1606 VDD.n53 VSS 5.83e-19
C1607 VDD.n54 VSS 0.00169f
C1608 VDD.n55 VSS 7.86e-19
C1609 VDD.n56 VSS 6.64e-19
C1610 VDD.t141 VSS 6.91e-19
C1611 VDD.t125 VSS 6.91e-19
C1612 VDD.n57 VSS 0.00163f
C1613 VDD.n58 VSS 0.00273f
C1614 VDD.t41 VSS 0.00122f
C1615 VDD.t5 VSS 3.55e-19
C1616 VDD.n59 VSS 0.00134f
C1617 VDD.n60 VSS 0.00196f
C1618 VDD.n61 VSS 4.74e-19
C1619 VDD.n62 VSS 0.00226f
C1620 VDD.n63 VSS 0.00226f
C1621 VDD.n64 VSS 4.78e-19
C1622 VDD.n65 VSS 5.09e-19
C1623 VDD.t131 VSS 0.00283f
C1624 VDD.n66 VSS 0.00441f
C1625 VDD.t101 VSS 0.00122f
C1626 VDD.t63 VSS 3.55e-19
C1627 VDD.n67 VSS 0.00134f
C1628 VDD.n68 VSS 0.00204f
C1629 VDD.n69 VSS 2.35e-19
C1630 VDD.n70 VSS 0.00169f
C1631 VDD.n71 VSS 9.21e-19
C1632 VDD.n72 VSS 8.23e-19
C1633 VDD.n73 VSS 8e-19
C1634 VDD.n74 VSS 8e-19
C1635 VDD.n75 VSS 9.79e-19
C1636 VDD.n76 VSS 0.00226f
C1637 VDD.n77 VSS 0.00226f
C1638 VDD.n78 VSS 7.46e-19
C1639 VDD.n79 VSS 8e-19
C1640 VDD.n80 VSS 8.01e-19
C1641 VDD.n81 VSS 0.00226f
C1642 VDD.n82 VSS 0.00226f
C1643 VDD.n83 VSS 8.01e-19
C1644 VDD.n84 VSS 8e-19
C1645 VDD.t13 VSS 0.00122f
C1646 VDD.t99 VSS 3.55e-19
C1647 VDD.n85 VSS 0.0013f
C1648 VDD.n86 VSS 0.00158f
C1649 VDD.n87 VSS 7.4e-19
C1650 VDD.n88 VSS 0.00226f
C1651 VDD.n89 VSS 0.00226f
C1652 VDD.n90 VSS 0.00139f
C1653 VDD.n91 VSS 6.74e-19
C1654 VDD.n92 VSS 0.00416f
C1655 VDD.n93 VSS 5.83e-19
C1656 VDD.n94 VSS 0.00206f
C1657 VDD.n95 VSS 0.00169f
C1658 VDD.n96 VSS 8.6e-19
C1659 VDD.n97 VSS 0.00387f
C1660 VDD.n98 VSS 0.0313f
C1661 VDD.n99 VSS 0.0354f
C1662 VDD.n100 VSS 0.00408f
C1663 VDD.n101 VSS 0.00411f
C1664 VDD.n102 VSS 0.00408f
C1665 VDD.n103 VSS 0.00408f
C1666 VDD.n104 VSS 0.00416f
C1667 VDD.n105 VSS 0.015f
C1668 VDD.n106 VSS 3.72f
C1669 VDD.n107 VSS 0.00408f
C1670 VDD.n108 VSS 0.00408f
C1671 VDD.n109 VSS 0.00408f
C1672 VDD.n110 VSS 0.00408f
C1673 VDD.n111 VSS 0.00408f
C1674 VDD.n112 VSS 0.00408f
C1675 VDD.n113 VSS 0.00408f
C1676 VDD.n114 VSS 0.00408f
C1677 VDD.n115 VSS 1.77f
C1678 VDD.n116 VSS 0.00408f
C1679 VDD.n117 VSS 0.00411f
C1680 VDD.n118 VSS 0.00408f
C1681 VDD.n119 VSS 0.00408f
C1682 VDD.n120 VSS 0.00408f
C1683 VDD.n121 VSS 0.00408f
C1684 VDD.n122 VSS 0.00408f
C1685 VDD.n123 VSS 0.00408f
C1686 VDD.n124 VSS 0.00418f
C1687 VDD.t144 VSS 4.73f
C1688 VDD.t145 VSS 4.73f
C1689 VDD.t149 VSS 5.39f
C1690 VDD.n125 VSS 1.71f
C1691 VDD.n126 VSS 1.71f
C1692 VDD.n127 VSS 0.038f
C1693 VDD.n128 VSS 0.759f
C1694 VDD.n129 VSS 0.0316f
C1695 VDD.n130 VSS 0.00238f
C1696 VDD.n131 VSS 0.0511f
C1697 VDD.n132 VSS 0.484f
C1698 VDD.n133 VSS 0.484f
C1699 VDD.n134 VSS 0.103f
C1700 VDD.n135 VSS 0.484f
C1701 VDD.n136 VSS 0.0512f
C1702 VDD.n137 VSS 0.0116f
C1703 VDD.n138 VSS -0.0813f
C1704 VDD.n139 VSS 0.00133f
C1705 VDD.n140 VSS -0.0588f
C1706 VDD.n141 VSS -0.0728f
C1707 VDD.t146 VSS 1.5f
C1708 VDD.n142 VSS 0.484f
C1709 VDD.n143 VSS 0.205f
C1710 VDD.n144 VSS 0.0304f
C1711 VDD.n145 VSS 0.0497f
C1712 VDD.n146 VSS 0.0507f
C1713 VDD.n147 VSS -0.0728f
C1714 VDD.n148 VSS 0.00133f
C1715 VDD.n149 VSS -0.0588f
C1716 VDD.n150 VSS -0.0728f
C1717 VDD.t148 VSS 1.5f
C1718 VDD.n151 VSS 0.484f
C1719 VDD.n152 VSS 0.205f
C1720 VDD.n153 VSS 0.0304f
C1721 VDD.n154 VSS 0.0497f
C1722 VDD.n155 VSS 0.0507f
C1723 VDD.n156 VSS -0.0728f
C1724 VDD.n157 VSS 0.00133f
C1725 VDD.n158 VSS -0.0588f
C1726 VDD.n159 VSS -0.0813f
C1727 VDD.t147 VSS 1.5f
C1728 VDD.n160 VSS 0.487f
C1729 VDD.n161 VSS 0.0584f
C1730 VDD.n162 VSS 0.0114f
C1731 VDD.n163 VSS 0.0427f
C1732 VDD.n164 VSS 0.0151f
C1733 VDD.n165 VSS 0.00532f
C1734 VDD.n166 VSS 0.00515f
C1735 VDD.n167 VSS 0.0051f
C1736 VDD.n168 VSS 0.00238f
C1737 VDD.n169 VSS 0.00408f
C1738 VDD.n170 VSS 0.00408f
C1739 VDD.n171 VSS 0.00408f
C1740 VDD.n172 VSS 0.00408f
C1741 VDD.n173 VSS 0.00408f
C1742 VDD.n174 VSS 0.00408f
C1743 VDD.n175 VSS 0.00408f
C1744 VDD.n176 VSS 0.00408f
C1745 VDD.n177 VSS 0.00408f
C1746 VDD.n178 VSS 0.00408f
C1747 VDD.n179 VSS 0.00408f
C1748 VDD.n180 VSS 0.00408f
C1749 VDD.n181 VSS 0.00449f
C1750 VDD.n182 VSS 0.0147f
C1751 VDD.n183 VSS 0.0236f
C1752 VDD.n184 VSS 0.0236f
C1753 VDD.n185 VSS 0.00473f
C1754 VDD.n186 VSS 0.00473f
C1755 VDD.n187 VSS 0.00408f
C1756 VDD.n188 VSS 0.00408f
C1757 VDD.n189 VSS 0.00416f
C1758 VDD.n190 VSS 0.015f
C1759 VDD.n191 VSS 0.258f
C1760 VDD.n192 VSS 0.00408f
C1761 VDD.n193 VSS 0.00408f
C1762 VDD.n194 VSS 0.258f
C1763 VDD.n195 VSS 0.00473f
C1764 VDD.n196 VSS 0.00473f
C1765 VDD.n197 VSS 0.693f
C1766 VDD.n198 VSS 0.698f
C1767 VDD.n199 VSS 0.00693f
C1768 VDD.n200 VSS 0.00693f
C1769 VDD.n202 VSS 0.00358f
C1770 VDD.n203 VSS 0.00358f
C1771 VDD.n204 VSS 0.00815f
C1772 VDD.n205 VSS 0.00115f
C1773 VDD.n206 VSS 0.00115f
C1774 VDD.n207 VSS 0.00244f
C1775 VDD.n208 VSS 3.72f
C1776 VDD.n210 VSS 0.00246f
C1777 VDD.n211 VSS 0.00117f
C1778 VDD.n212 VSS 0.00247f
C1779 VDD.n213 VSS 0.00355f
C1780 VDD.n214 VSS 0.01f
C1781 VDD.n215 VSS 0.00108f
C1782 VDD.n216 VSS 0.0081f
C1783 VDD.n217 VSS 0.0571f
C1784 VDD.n218 VSS 0.0536f
C1785 VDD.n219 VSS 0.00803f
C1786 VDD.n220 VSS 6.49e-19
C1787 VDD.n221 VSS 4.61e-19
C1788 VDD.n222 VSS 6.74e-19
C1789 VDD.n223 VSS 0.00226f
C1790 VDD.n224 VSS 6.74e-19
C1791 VDD.t143 VSS 0.00281f
C1792 VDD.n225 VSS 0.00226f
C1793 VDD.n226 VSS 8.01e-19
C1794 VDD.n227 VSS 0.00226f
C1795 VDD.t35 VSS 0.00122f
C1796 VDD.t95 VSS 3.55e-19
C1797 VDD.n228 VSS 0.0013f
C1798 VDD.n229 VSS 0.00155f
C1799 VDD.n230 VSS 0.00169f
C1800 VDD.n231 VSS 0.00404f
C1801 VDD.n232 VSS 0.00226f
C1802 VDD.t19 VSS 6.91e-19
C1803 VDD.t17 VSS 6.91e-19
C1804 VDD.n233 VSS 0.00158f
C1805 VDD.n234 VSS 0.0027f
C1806 VDD.n235 VSS 0.00204f
C1807 VDD.t59 VSS 0.00122f
C1808 VDD.t57 VSS 3.55e-19
C1809 VDD.n236 VSS 0.0013f
C1810 VDD.n237 VSS 0.00155f
C1811 VDD.n238 VSS 0.00169f
C1812 VDD.n239 VSS 3.48e-19
C1813 VDD.n240 VSS 8.01e-19
C1814 VDD.n241 VSS 7.46e-19
C1815 VDD.t96 VSS 0.0111f
C1816 VDD.t142 VSS 0.0147f
C1817 VDD.t118 VSS 0.00759f
C1818 VDD.t120 VSS 0.00961f
C1819 VDD.t134 VSS 0.00867f
C1820 VDD.t116 VSS 0.0136f
C1821 VDD.t36 VSS 0.0186f
C1822 VDD.t22 VSS 0.0115f
C1823 VDD.t114 VSS 0.0136f
C1824 VDD.t94 VSS 0.0114f
C1825 VDD.t115 VSS 0.00687f
C1826 VDD.t34 VSS 0.0155f
C1827 VDD.n242 VSS 0.0097f
C1828 VDD.t122 VSS 0.00608f
C1829 VDD.n243 VSS 0.00838f
C1830 VDD.t10 VSS 0.0122f
C1831 VDD.t20 VSS 0.0119f
C1832 VDD.t16 VSS 0.00775f
C1833 VDD.t60 VSS 0.00608f
C1834 VDD.t18 VSS 0.00688f
C1835 VDD.t6 VSS 0.00608f
C1836 VDD.t14 VSS 0.0097f
C1837 VDD.t110 VSS 0.00825f
C1838 VDD.t56 VSS 0.00862f
C1839 VDD.t58 VSS 0.0117f
C1840 VDD.t74 VSS 0.0109f
C1841 VDD.t70 VSS 0.0063f
C1842 VDD.t76 VSS 0.0076f
C1843 VDD.t80 VSS 0.00608f
C1844 VDD.t72 VSS 0.00688f
C1845 VDD.t136 VSS 0.00608f
C1846 VDD.t32 VSS 0.00572f
C1847 VDD.t46 VSS 0.0148f
C1848 VDD.t38 VSS 0.00695f
C1849 VDD.t30 VSS 0.00529f
C1850 VDD.t44 VSS 0.0148f
C1851 VDD.t24 VSS 0.00688f
C1852 VDD.t64 VSS 0.00521f
C1853 VDD.n244 VSS 0.0131f
C1854 VDD.n245 VSS 7.74e-19
C1855 VDD.n246 VSS 3.7e-19
C1856 VDD.t25 VSS 0.0028f
C1857 VDD.n247 VSS 0.00289f
C1858 VDD.t65 VSS 0.00122f
C1859 VDD.t45 VSS 3.55e-19
C1860 VDD.n248 VSS 0.0013f
C1861 VDD.n249 VSS 0.00155f
C1862 VDD.n250 VSS 7e-19
C1863 VDD.n251 VSS 0.00205f
C1864 VDD.n252 VSS 0.00169f
C1865 VDD.n253 VSS 7.74e-19
C1866 VDD.n254 VSS 4.96e-19
C1867 VDD.t31 VSS 0.0028f
C1868 VDD.n255 VSS 0.00289f
C1869 VDD.t39 VSS 0.00122f
C1870 VDD.t47 VSS 3.55e-19
C1871 VDD.n256 VSS 0.0013f
C1872 VDD.n257 VSS 0.00167f
C1873 VDD.n258 VSS 5.22e-19
C1874 VDD.n259 VSS 0.00205f
C1875 VDD.n260 VSS 0.00169f
C1876 VDD.n261 VSS 7.86e-19
C1877 VDD.n262 VSS 8e-19
C1878 VDD.t33 VSS 6.91e-19
C1879 VDD.t73 VSS 6.91e-19
C1880 VDD.n263 VSS 0.00158f
C1881 VDD.t137 VSS 0.00122f
C1882 VDD.t81 VSS 3.55e-19
C1883 VDD.n264 VSS 0.00134f
C1884 VDD.n265 VSS 0.00202f
C1885 VDD.n266 VSS 0.002f
C1886 VDD.n267 VSS 4.22e-19
C1887 VDD.n268 VSS 0.00204f
C1888 VDD.n269 VSS 0.00226f
C1889 VDD.n270 VSS 0.00139f
C1890 VDD.t77 VSS 6.91e-19
C1891 VDD.t71 VSS 6.91e-19
C1892 VDD.n271 VSS 0.00164f
C1893 VDD.n272 VSS 0.00353f
C1894 VDD.n273 VSS 4.44e-19
C1895 VDD.t75 VSS 0.00283f
C1896 VDD.n274 VSS 0.00441f
C1897 VDD.n275 VSS 5.83e-19
C1898 VDD.n276 VSS 0.00169f
C1899 VDD.n277 VSS 7.86e-19
C1900 VDD.n278 VSS 6.64e-19
C1901 VDD.t111 VSS 6.91e-19
C1902 VDD.t15 VSS 6.91e-19
C1903 VDD.n279 VSS 0.00163f
C1904 VDD.n280 VSS 0.00273f
C1905 VDD.t7 VSS 0.00122f
C1906 VDD.t61 VSS 3.55e-19
C1907 VDD.n281 VSS 0.00134f
C1908 VDD.n282 VSS 0.00196f
C1909 VDD.n283 VSS 4.74e-19
C1910 VDD.n284 VSS 0.00226f
C1911 VDD.n285 VSS 0.00226f
C1912 VDD.n286 VSS 4.78e-19
C1913 VDD.n287 VSS 5.09e-19
C1914 VDD.t21 VSS 0.00283f
C1915 VDD.n288 VSS 0.00441f
C1916 VDD.t11 VSS 0.00122f
C1917 VDD.t123 VSS 3.55e-19
C1918 VDD.n289 VSS 0.00134f
C1919 VDD.n290 VSS 0.00204f
C1920 VDD.n291 VSS 2.35e-19
C1921 VDD.n292 VSS 0.00169f
C1922 VDD.n293 VSS 9.21e-19
C1923 VDD.n294 VSS 8.23e-19
C1924 VDD.n295 VSS 8e-19
C1925 VDD.n296 VSS 8e-19
C1926 VDD.n297 VSS 9.79e-19
C1927 VDD.n298 VSS 0.00226f
C1928 VDD.n299 VSS 0.00226f
C1929 VDD.n300 VSS 7.46e-19
C1930 VDD.n301 VSS 8e-19
C1931 VDD.t23 VSS 0.00122f
C1932 VDD.t37 VSS 3.55e-19
C1933 VDD.n302 VSS 0.0013f
C1934 VDD.n303 VSS 0.00167f
C1935 VDD.n304 VSS 8.01e-19
C1936 VDD.n305 VSS 0.00226f
C1937 VDD.n306 VSS 0.00226f
C1938 VDD.n307 VSS 0.00226f
C1939 VDD.n308 VSS 8e-19
C1940 VDD.n309 VSS 4.61e-19
C1941 VDD.t135 VSS 0.00122f
C1942 VDD.t121 VSS 3.55e-19
C1943 VDD.n310 VSS 0.00135f
C1944 VDD.t117 VSS 3.71e-19
C1945 VDD.t119 VSS 3.71e-19
C1946 VDD.n311 VSS 7.42e-19
C1947 VDD.t42 VSS 3.71e-19
C1948 VDD.t43 VSS 3.71e-19
C1949 VDD.n312 VSS 0.00246f
C1950 VDD.n313 VSS 0.00208f
C1951 VDD.n314 VSS 0.00312f
C1952 VDD.n315 VSS 4.04e-19
C1953 VDD.n316 VSS 0.00226f
C1954 VDD.n317 VSS 0.00139f
C1955 VDD.n318 VSS 0.00169f
C1956 VDD.n319 VSS 0.00391f
C1957 VDD.n320 VSS 5.83e-19
C1958 VDD.t97 VSS 0.00281f
C1959 VDD.n321 VSS 0.00416f
C1960 VDD.n322 VSS 0.00135f
C1961 VDD.n323 VSS 0.00169f
C1962 VDD.n324 VSS 7.74e-19
C1963 VDD.n325 VSS 0.00142f
C1964 VDD.t9 VSS 0.00272f
C1965 VDD.n326 VSS 0.00279f
C1966 VDD.n327 VSS 0.00409f
C1967 VDD.n328 VSS 0.0137f
C1968 VDD.t8 VSS 0.00607f
C1969 VDD.n329 VSS 0.0117f
C1970 VDD.n330 VSS 0.00548f
C1971 VDD.n331 VSS 0.00728f
C1972 VDD.n332 VSS 8.6e-19
C1973 VDD.n333 VSS 0.0141f
C1974 VDD.n334 VSS 0.0028f
C1975 VDD.n335 VSS 0.00209f
C1976 VDD.n336 VSS 6.74e-19
C1977 VDD.n337 VSS 0.00804f
C1978 VDD.n338 VSS 0.00279f
C1979 VDD.n339 VSS 0.0028f
C1980 VDD.n340 VSS 0.00253f
C1981 VDD.n341 VSS 6.6e-19
C1982 VDD.n342 VSS 1.92f
C1983 VDD.n343 VSS 0.00405f
C1984 VDD.n344 VSS 0.0536f
C1985 VDD.n345 VSS 0.0537f
C1986 VDD.n346 VSS 0.00279f
C1987 VDD.n347 VSS 0.0028f
C1988 VDD.n348 VSS 0.00187f
C1989 VDD.n349 VSS 6.42e-19
C1990 VDD.n350 VSS 0.00405f
C1991 VDD.n352 VSS 0.0028f
C1992 VDD.n353 VSS 0.0028f
C1993 VDD.n354 VSS 0.015f
C1994 vcm.n0 VSS 2.37f
C1995 vcm.n1 VSS 0.243f
C1996 vcm.n2 VSS 2.37f
C1997 vcm.n3 VSS 0.243f
C1998 vcm.n4 VSS 2.37f
C1999 vcm.n5 VSS 0.243f
C2000 vcm.n6 VSS 2.37f
C2001 vcm.n7 VSS 0.243f
C2002 vcm.t58 VSS 7.38f
C2003 vcm.n8 VSS 0.504f
C2004 vcm.n9 VSS 2.38f
C2005 vcm.n10 VSS 0.251f
C2006 vcm.n11 VSS 0.0571f
C2007 vcm.n12 VSS -0.399f
C2008 vcm.n13 VSS 0.0142f
C2009 vcm.n14 VSS 0.504f
C2010 vcm.n15 VSS 2.38f
C2011 vcm.n16 VSS 0.251f
C2012 vcm.n17 VSS 0.0571f
C2013 vcm.n18 VSS -0.399f
C2014 vcm.n19 VSS 0.405f
C2015 vcm.n20 VSS -0.0315f
C2016 vcm.n21 VSS -0.342f
C2017 vcm.n22 VSS -0.288f
C2018 vcm.n23 VSS 0.428f
C2019 vcm.n24 VSS -0.0316f
C2020 vcm.n25 VSS -0.365f
C2021 vcm.n26 VSS -0.288f
C2022 vcm.n27 VSS -0.358f
C2023 vcm.n28 VSS 2.37f
C2024 vcm.n29 VSS 1.01f
C2025 vcm.n30 VSS 0.242f
C2026 vcm.n31 VSS 0.157f
C2027 vcm.n32 VSS -0.358f
C2028 vcm.n33 VSS 0.0139f
C2029 vcm.n34 VSS 0.405f
C2030 vcm.n35 VSS -0.0313f
C2031 vcm.n36 VSS 2.37f
C2032 vcm.n37 VSS 0.243f
C2033 vcm.n38 VSS -0.358f
C2034 vcm.t21 VSS 7.38f
C2035 vcm.n39 VSS 2.37f
C2036 vcm.n40 VSS 1.01f
C2037 vcm.n41 VSS 0.242f
C2038 vcm.n42 VSS 0.157f
C2039 vcm.n43 VSS -0.358f
C2040 vcm.n44 VSS 0.428f
C2041 vcm.n45 VSS -0.0316f
C2042 vcm.n46 VSS -0.365f
C2043 vcm.n47 VSS -0.288f
C2044 vcm.n48 VSS -0.342f
C2045 vcm.n49 VSS -0.288f
C2046 vcm.n50 VSS -0.358f
C2047 vcm.t52 VSS 7.39f
C2048 vcm.n51 VSS 2.37f
C2049 vcm.n52 VSS 1.01f
C2050 vcm.n53 VSS 0.242f
C2051 vcm.n54 VSS 0.157f
C2052 vcm.n55 VSS -0.358f
C2053 vcm.n56 VSS 0.0142f
C2054 vcm.n57 VSS 0.428f
C2055 vcm.n58 VSS -0.0316f
C2056 vcm.n59 VSS -0.365f
C2057 vcm.n60 VSS -0.288f
C2058 vcm.n61 VSS -0.358f
C2059 vcm.t41 VSS 7.39f
C2060 vcm.n62 VSS 2.37f
C2061 vcm.n63 VSS 1.01f
C2062 vcm.n64 VSS 0.242f
C2063 vcm.n65 VSS 0.157f
C2064 vcm.n66 VSS -0.358f
C2065 vcm.n67 VSS 0.0139f
C2066 vcm.n68 VSS 0.405f
C2067 vcm.n69 VSS -0.0313f
C2068 vcm.n70 VSS 2.37f
C2069 vcm.n71 VSS 0.243f
C2070 vcm.n72 VSS 2.37f
C2071 vcm.n73 VSS 0.243f
C2072 vcm.n74 VSS -0.358f
C2073 vcm.t15 VSS 7.39f
C2074 vcm.n75 VSS 2.37f
C2075 vcm.n76 VSS 1.01f
C2076 vcm.n77 VSS 0.242f
C2077 vcm.n78 VSS 0.157f
C2078 vcm.n79 VSS -0.358f
C2079 vcm.n80 VSS 0.405f
C2080 vcm.n81 VSS -0.0315f
C2081 vcm.n82 VSS -0.342f
C2082 vcm.n83 VSS -0.288f
C2083 vcm.n84 VSS -0.358f
C2084 vcm.t8 VSS 7.39f
C2085 vcm.n85 VSS 2.37f
C2086 vcm.n86 VSS 1.01f
C2087 vcm.n87 VSS 0.242f
C2088 vcm.n88 VSS 0.157f
C2089 vcm.n89 VSS -0.358f
C2090 vcm.n90 VSS 0.428f
C2091 vcm.n91 VSS -0.0316f
C2092 vcm.n92 VSS -0.365f
C2093 vcm.n93 VSS -0.288f
C2094 vcm.n94 VSS -0.342f
C2095 vcm.n95 VSS -0.288f
C2096 vcm.n96 VSS -0.358f
C2097 vcm.t53 VSS 7.39f
C2098 vcm.n97 VSS 2.37f
C2099 vcm.n98 VSS 1.01f
C2100 vcm.n99 VSS 0.242f
C2101 vcm.n100 VSS 0.157f
C2102 vcm.n101 VSS -0.358f
C2103 vcm.n102 VSS 0.0142f
C2104 vcm.n103 VSS 2.37f
C2105 vcm.n104 VSS 0.243f
C2106 vcm.n105 VSS -0.358f
C2107 vcm.t16 VSS 7.39f
C2108 vcm.n106 VSS 2.37f
C2109 vcm.n107 VSS 1.01f
C2110 vcm.n108 VSS 0.242f
C2111 vcm.n109 VSS 0.157f
C2112 vcm.n110 VSS -0.358f
C2113 vcm.n111 VSS 0.405f
C2114 vcm.n112 VSS -0.0315f
C2115 vcm.n113 VSS -0.342f
C2116 vcm.n114 VSS -0.288f
C2117 vcm.n115 VSS 0.428f
C2118 vcm.n116 VSS -0.0316f
C2119 vcm.n117 VSS -0.365f
C2120 vcm.n118 VSS -0.288f
C2121 vcm.n119 VSS 0.332f
C2122 vcm.t44 VSS 7.39f
C2123 vcm.n120 VSS 2.39f
C2124 vcm.n121 VSS -0.38f
C2125 vcm.n122 VSS 0.156f
C2126 vcm.n123 VSS 0.146f
C2127 vcm.n124 VSS 0.0527f
C2128 vcm.n125 VSS 0.0394f
C2129 vcm.n126 VSS 0.0394f
C2130 vcm.n128 VSS 1.02f
C2131 vcm.n130 VSS 0.0527f
C2132 vcm.n131 VSS 0.0394f
C2133 vcm.n132 VSS 0.0394f
C2134 vcm.n133 VSS 0.0527f
C2135 vcm.n134 VSS 0.0394f
C2136 vcm.n135 VSS 0.0394f
C2137 vcm.n136 VSS 0.0527f
C2138 vcm.n137 VSS 0.0394f
C2139 vcm.n138 VSS 0.0394f
C2140 vcm.n139 VSS 0.0527f
C2141 vcm.n140 VSS 0.0394f
C2142 vcm.n141 VSS 0.0394f
C2143 vcm.n143 VSS 1.1f
C2144 vcm.n144 VSS 0.146f
C2145 vcm.n146 VSS 0.243f
C2146 vcm.n147 VSS 0.0587f
C2147 vcm.n148 VSS 2.37f
C2148 vcm.t73 VSS 7.38f
C2149 vcm.n149 VSS 2.38f
C2150 vcm.n150 VSS 2.38f
C2151 vcm.t70 VSS 7.38f
C2152 vcm.n151 VSS 2.38f
C2153 vcm.t68 VSS 7.38f
C2154 vcm.n152 VSS 0.504f
C2155 vcm.n153 VSS 2.38f
C2156 vcm.n154 VSS 0.251f
C2157 vcm.n155 VSS 0.0571f
C2158 vcm.n156 VSS -0.399f
C2159 vcm.n157 VSS 0.0145f
C2160 vcm.n158 VSS -0.288f
C2161 vcm.n159 VSS -0.358f
C2162 vcm.n160 VSS 2.37f
C2163 vcm.n161 VSS 1.01f
C2164 vcm.n162 VSS 0.159f
C2165 vcm.n163 VSS 0.242f
C2166 vcm.n164 VSS 0.242f
C2167 vcm.n165 VSS -0.358f
C2168 vcm.n166 VSS 0.0145f
C2169 vcm.n167 VSS -0.288f
C2170 vcm.n168 VSS -0.358f
C2171 vcm.n169 VSS 2.37f
C2172 vcm.n170 VSS 1.01f
C2173 vcm.n171 VSS 0.159f
C2174 vcm.n172 VSS 0.242f
C2175 vcm.n173 VSS 0.242f
C2176 vcm.n174 VSS -0.358f
C2177 vcm.n175 VSS 0.0145f
C2178 vcm.n176 VSS -0.288f
C2179 vcm.n177 VSS -0.358f
C2180 vcm.t74 VSS 7.38f
C2181 vcm.n178 VSS 2.37f
C2182 vcm.n179 VSS 1.01f
C2183 vcm.n180 VSS 0.159f
C2184 vcm.n181 VSS 0.242f
C2185 vcm.n182 VSS 0.242f
C2186 vcm.n183 VSS -0.358f
C2187 vcm.n184 VSS 0.0145f
C2188 vcm.n185 VSS -0.288f
C2189 vcm.n186 VSS -0.358f
C2190 vcm.n187 VSS 2.37f
C2191 vcm.n188 VSS 1.01f
C2192 vcm.n189 VSS 0.159f
C2193 vcm.n190 VSS 0.242f
C2194 vcm.n191 VSS 0.242f
C2195 vcm.n192 VSS -0.358f
C2196 vcm.n193 VSS 0.0145f
C2197 vcm.n194 VSS -0.288f
C2198 vcm.n195 VSS -0.399f
C2199 vcm.t77 VSS 7.39f
C2200 vcm.n196 VSS 2.39f
C2201 vcm.n197 VSS 0.324f
C2202 vcm.n198 VSS 0.193f
C2203 vcm.n199 VSS 0.211f
C2204 vcm.n200 VSS 0.0445f
C2205 vcm.n201 VSS 0.0445f
C2206 vcm.n203 VSS 1f
C2207 vcm.n204 VSS 1f
C2208 vcm.n205 VSS 0.146f
C2209 vcm.n207 VSS 2.38f
C2210 vcm.n208 VSS 2.37f
C2211 vcm.t61 VSS 7.38f
C2212 vcm.n209 VSS 2.38f
C2213 vcm.n210 VSS 2.38f
C2214 vcm.n211 VSS 0.504f
C2215 vcm.n212 VSS 2.38f
C2216 vcm.n213 VSS 0.251f
C2217 vcm.n214 VSS 0.0571f
C2218 vcm.n215 VSS -0.399f
C2219 vcm.n216 VSS 0.405f
C2220 vcm.n217 VSS -0.0315f
C2221 vcm.n218 VSS -0.342f
C2222 vcm.n219 VSS -0.288f
C2223 vcm.n220 VSS -0.358f
C2224 vcm.t36 VSS 7.38f
C2225 vcm.n221 VSS 2.37f
C2226 vcm.n222 VSS 1.01f
C2227 vcm.n223 VSS 0.159f
C2228 vcm.n224 VSS 0.242f
C2229 vcm.n225 VSS 0.242f
C2230 vcm.n226 VSS -0.358f
C2231 vcm.n227 VSS 0.405f
C2232 vcm.n228 VSS -0.0315f
C2233 vcm.n229 VSS -0.342f
C2234 vcm.n230 VSS -0.288f
C2235 vcm.n231 VSS -0.358f
C2236 vcm.t86 VSS 7.38f
C2237 vcm.n232 VSS 2.37f
C2238 vcm.n233 VSS 1.01f
C2239 vcm.n234 VSS 0.159f
C2240 vcm.n235 VSS 0.242f
C2241 vcm.n236 VSS 0.242f
C2242 vcm.n237 VSS -0.358f
C2243 vcm.n238 VSS 0.428f
C2244 vcm.n239 VSS -0.0316f
C2245 vcm.n240 VSS -0.365f
C2246 vcm.n241 VSS -0.288f
C2247 vcm.n242 VSS -0.358f
C2248 vcm.n243 VSS 2.37f
C2249 vcm.n244 VSS 1.01f
C2250 vcm.n245 VSS 0.159f
C2251 vcm.n246 VSS 0.242f
C2252 vcm.n247 VSS 0.242f
C2253 vcm.n248 VSS -0.358f
C2254 vcm.n249 VSS 0.405f
C2255 vcm.n250 VSS -0.0315f
C2256 vcm.n251 VSS -0.342f
C2257 vcm.n252 VSS -0.288f
C2258 vcm.n253 VSS -0.358f
C2259 vcm.t13 VSS 7.39f
C2260 vcm.n254 VSS 2.37f
C2261 vcm.n255 VSS 1.01f
C2262 vcm.n256 VSS 0.149f
C2263 vcm.n257 VSS 0.244f
C2264 vcm.n258 VSS 0.249f
C2265 vcm.n259 VSS -0.358f
C2266 vcm.n260 VSS 0.405f
C2267 vcm.n261 VSS -0.0297f
C2268 vcm.n262 VSS -0.341f
C2269 vcm.n263 VSS -0.288f
C2270 vcm.n264 VSS 0.243f
C2271 vcm.n265 VSS 0.0587f
C2272 vcm.n266 VSS -0.399f
C2273 vcm.t67 VSS 7.38f
C2274 vcm.n267 VSS 2.39f
C2275 vcm.n268 VSS 0.324f
C2276 vcm.n269 VSS 0.193f
C2277 vcm.n270 VSS 0.211f
C2278 vcm.n271 VSS 0.0445f
C2279 vcm.n272 VSS 0.0445f
C2280 vcm.n274 VSS 1.01f
C2281 vcm.n275 VSS 1.01f
C2282 vcm.n276 VSS 0.146f
C2283 vcm.n278 VSS 0.0527f
C2284 vcm.n279 VSS 0.0394f
C2285 vcm.n280 VSS 0.0394f
C2286 vcm.n281 VSS 0.243f
C2287 vcm.n282 VSS 0.0589f
C2288 vcm.n283 VSS 2.38f
C2289 vcm.t84 VSS 7.39f
C2290 vcm.n284 VSS 2.37f
C2291 vcm.t49 VSS 7.39f
C2292 vcm.n285 VSS 2.37f
C2293 vcm.t79 VSS 7.39f
C2294 vcm.n286 VSS 2.37f
C2295 vcm.t23 VSS 7.38f
C2296 vcm.n287 VSS 0.504f
C2297 vcm.n288 VSS 2.38f
C2298 vcm.n289 VSS 0.251f
C2299 vcm.n290 VSS 0.0571f
C2300 vcm.n291 VSS -0.399f
C2301 vcm.n292 VSS 0.428f
C2302 vcm.n293 VSS -0.0316f
C2303 vcm.n294 VSS -0.365f
C2304 vcm.n295 VSS -0.288f
C2305 vcm.n296 VSS -0.358f
C2306 vcm.n297 VSS 2.37f
C2307 vcm.n298 VSS 1.01f
C2308 vcm.n299 VSS 0.159f
C2309 vcm.n300 VSS 0.242f
C2310 vcm.n301 VSS 0.242f
C2311 vcm.n302 VSS -0.358f
C2312 vcm.n303 VSS 0.405f
C2313 vcm.n304 VSS -0.0315f
C2314 vcm.n305 VSS -0.342f
C2315 vcm.n306 VSS -0.288f
C2316 vcm.n307 VSS -0.358f
C2317 vcm.n308 VSS 2.37f
C2318 vcm.n309 VSS 1.01f
C2319 vcm.n310 VSS 0.159f
C2320 vcm.n311 VSS 0.242f
C2321 vcm.n312 VSS 0.242f
C2322 vcm.n313 VSS -0.358f
C2323 vcm.n314 VSS 0.405f
C2324 vcm.n315 VSS -0.0315f
C2325 vcm.n316 VSS -0.342f
C2326 vcm.n317 VSS -0.288f
C2327 vcm.n318 VSS -0.358f
C2328 vcm.n319 VSS 2.37f
C2329 vcm.n320 VSS 1.01f
C2330 vcm.n321 VSS 0.149f
C2331 vcm.n322 VSS 0.244f
C2332 vcm.n323 VSS 0.249f
C2333 vcm.n324 VSS -0.358f
C2334 vcm.n325 VSS 0.404f
C2335 vcm.n326 VSS -0.0298f
C2336 vcm.n327 VSS -0.341f
C2337 vcm.n328 VSS -0.288f
C2338 vcm.n329 VSS -0.358f
C2339 vcm.n330 VSS 2.37f
C2340 vcm.n331 VSS 1.01f
C2341 vcm.n332 VSS 0.159f
C2342 vcm.n333 VSS 0.242f
C2343 vcm.n334 VSS 0.242f
C2344 vcm.n335 VSS -0.358f
C2345 vcm.n336 VSS 0.404f
C2346 vcm.n337 VSS -0.0297f
C2347 vcm.n338 VSS -0.341f
C2348 vcm.n339 VSS -0.288f
C2349 vcm.n340 VSS -0.399f
C2350 vcm.t57 VSS 7.38f
C2351 vcm.n341 VSS 2.39f
C2352 vcm.n342 VSS 0.324f
C2353 vcm.n343 VSS 0.193f
C2354 vcm.n344 VSS 0.211f
C2355 vcm.n345 VSS 0.0445f
C2356 vcm.n346 VSS 0.0445f
C2357 vcm.n348 VSS 0.996f
C2358 vcm.n349 VSS 0.996f
C2359 vcm.t37 VSS 7.39f
C2360 vcm.n350 VSS 0.404f
C2361 vcm.n351 VSS -0.0298f
C2362 vcm.n352 VSS -0.341f
C2363 vcm.n353 VSS 0.404f
C2364 vcm.n354 VSS -0.0297f
C2365 vcm.n355 VSS -0.341f
C2366 vcm.n356 VSS 2.37f
C2367 vcm.n357 VSS 2.38f
C2368 vcm.t35 VSS 7.39f
C2369 vcm.n358 VSS 2.37f
C2370 vcm.n359 VSS 2.37f
C2371 vcm.n360 VSS 0.504f
C2372 vcm.n361 VSS 2.38f
C2373 vcm.n362 VSS 0.251f
C2374 vcm.n363 VSS 0.0571f
C2375 vcm.n364 VSS -0.399f
C2376 vcm.n365 VSS 0.405f
C2377 vcm.n366 VSS -0.0315f
C2378 vcm.n367 VSS -0.342f
C2379 vcm.n368 VSS 0.405f
C2380 vcm.n369 VSS -0.0315f
C2381 vcm.n370 VSS -0.342f
C2382 vcm.n371 VSS -0.288f
C2383 vcm.n372 VSS -0.358f
C2384 vcm.t54 VSS 7.38f
C2385 vcm.n373 VSS 2.37f
C2386 vcm.n374 VSS 1.01f
C2387 vcm.n375 VSS 0.159f
C2388 vcm.n376 VSS 0.242f
C2389 vcm.n377 VSS 0.242f
C2390 vcm.n378 VSS -0.358f
C2391 vcm.n379 VSS 0.404f
C2392 vcm.n380 VSS -0.0298f
C2393 vcm.n381 VSS -0.341f
C2394 vcm.n382 VSS 0.428f
C2395 vcm.n383 VSS -0.0316f
C2396 vcm.n384 VSS -0.365f
C2397 vcm.n385 VSS -0.288f
C2398 vcm.n386 VSS -0.358f
C2399 vcm.t45 VSS 7.39f
C2400 vcm.n387 VSS 2.37f
C2401 vcm.n388 VSS 1.01f
C2402 vcm.n389 VSS 0.149f
C2403 vcm.n390 VSS 0.244f
C2404 vcm.n391 VSS 0.249f
C2405 vcm.n392 VSS -0.358f
C2406 vcm.n393 VSS 0.404f
C2407 vcm.n394 VSS -0.0297f
C2408 vcm.n395 VSS -0.341f
C2409 vcm.n396 VSS 0.404f
C2410 vcm.n397 VSS -0.0297f
C2411 vcm.n398 VSS -0.341f
C2412 vcm.n399 VSS -0.288f
C2413 vcm.n400 VSS -0.358f
C2414 vcm.n401 VSS 2.37f
C2415 vcm.n402 VSS 1.01f
C2416 vcm.n403 VSS 0.159f
C2417 vcm.n404 VSS 0.242f
C2418 vcm.n405 VSS 0.242f
C2419 vcm.n406 VSS -0.358f
C2420 vcm.n407 VSS 0.404f
C2421 vcm.n408 VSS -0.0297f
C2422 vcm.n409 VSS -0.341f
C2423 vcm.n410 VSS 0.404f
C2424 vcm.n411 VSS -0.0297f
C2425 vcm.n412 VSS -0.341f
C2426 vcm.n413 VSS -0.288f
C2427 vcm.n414 VSS -0.358f
C2428 vcm.t46 VSS 7.38f
C2429 vcm.n415 VSS 2.37f
C2430 vcm.n416 VSS 1.01f
C2431 vcm.n417 VSS 0.159f
C2432 vcm.n418 VSS 0.242f
C2433 vcm.n419 VSS 0.242f
C2434 vcm.n420 VSS -0.358f
C2435 vcm.n421 VSS -0.288f
C2436 vcm.n422 VSS -0.399f
C2437 vcm.n423 VSS 2.39f
C2438 vcm.n424 VSS 0.326f
C2439 vcm.n425 VSS 0.243f
C2440 vcm.n426 VSS 0.0583f
C2441 vcm.n427 VSS 0.192f
C2442 vcm.n428 VSS 0.211f
C2443 vcm.n429 VSS 0.0445f
C2444 vcm.n430 VSS 0.0445f
C2445 vcm.n432 VSS 0.0527f
C2446 vcm.n433 VSS 0.0394f
C2447 vcm.n434 VSS 0.0394f
C2448 vcm.n436 VSS 0.146f
C2449 vcm.n438 VSS 0.959f
C2450 vcm.n439 VSS 0.959f
C2451 vcm.n440 VSS 0.146f
C2452 vcm.n442 VSS 0.0527f
C2453 vcm.n443 VSS 0.0394f
C2454 vcm.n444 VSS 0.0394f
C2455 vcm.n445 VSS 2.38f
C2456 vcm.t31 VSS 7.39f
C2457 vcm.n446 VSS 2.37f
C2458 vcm.n447 VSS 2.38f
C2459 vcm.t28 VSS 7.39f
C2460 vcm.n448 VSS 2.37f
C2461 vcm.n449 VSS 0.504f
C2462 vcm.n450 VSS 2.37f
C2463 vcm.n451 VSS 0.251f
C2464 vcm.n452 VSS 0.0571f
C2465 vcm.n453 VSS -0.399f
C2466 vcm.n454 VSS -0.288f
C2467 vcm.n455 VSS -0.358f
C2468 vcm.t38 VSS 7.39f
C2469 vcm.n456 VSS 2.37f
C2470 vcm.n457 VSS 1.01f
C2471 vcm.n458 VSS 0.149f
C2472 vcm.n459 VSS 0.244f
C2473 vcm.n460 VSS 0.249f
C2474 vcm.n461 VSS -0.358f
C2475 vcm.n462 VSS -0.288f
C2476 vcm.n463 VSS -0.358f
C2477 vcm.n464 VSS 2.37f
C2478 vcm.n465 VSS 1.01f
C2479 vcm.n466 VSS 0.159f
C2480 vcm.n467 VSS 0.242f
C2481 vcm.n468 VSS 0.242f
C2482 vcm.n469 VSS -0.358f
C2483 vcm.n470 VSS -0.288f
C2484 vcm.n471 VSS -0.358f
C2485 vcm.t22 VSS 7.38f
C2486 vcm.n472 VSS 2.37f
C2487 vcm.n473 VSS 1.01f
C2488 vcm.n474 VSS 0.159f
C2489 vcm.n475 VSS 0.242f
C2490 vcm.n476 VSS 0.242f
C2491 vcm.n477 VSS -0.358f
C2492 vcm.n478 VSS -0.288f
C2493 vcm.n479 VSS -0.358f
C2494 vcm.n480 VSS 2.37f
C2495 vcm.n481 VSS 1.01f
C2496 vcm.n482 VSS 0.159f
C2497 vcm.n483 VSS 0.242f
C2498 vcm.n484 VSS 0.242f
C2499 vcm.n485 VSS -0.358f
C2500 vcm.n486 VSS -0.288f
C2501 vcm.n487 VSS 0.332f
C2502 vcm.t24 VSS 7.38f
C2503 vcm.n488 VSS 2.39f
C2504 vcm.n489 VSS -0.38f
C2505 vcm.n490 VSS 0.156f
C2506 vcm.n491 VSS 0.177f
C2507 vcm.n492 VSS 0.194f
C2508 vcm.n493 VSS 0.211f
C2509 vcm.n494 VSS 0.0445f
C2510 vcm.n495 VSS 0.0445f
C2511 vcm.n497 VSS 1.03f
C2512 vcm.n498 VSS 1.03f
C2513 vcm.n499 VSS 0.243f
C2514 vcm.n500 VSS 0.329f
C2515 vcm.t60 VSS 7.38f
C2516 vcm.n501 VSS 2.39f
C2517 vcm.n502 VSS 2.38f
C2518 vcm.t66 VSS 7.39f
C2519 vcm.n503 VSS 2.37f
C2520 vcm.t59 VSS 7.38f
C2521 vcm.n504 VSS 2.38f
C2522 vcm.n505 VSS 2.38f
C2523 vcm.n506 VSS 0.504f
C2524 vcm.n507 VSS 2.38f
C2525 vcm.n508 VSS 0.251f
C2526 vcm.n509 VSS 0.0571f
C2527 vcm.n510 VSS -0.399f
C2528 vcm.n511 VSS 0.404f
C2529 vcm.n512 VSS -0.0297f
C2530 vcm.n513 VSS -0.341f
C2531 vcm.n514 VSS -0.288f
C2532 vcm.n515 VSS -0.358f
C2533 vcm.t72 VSS 7.38f
C2534 vcm.n516 VSS 2.37f
C2535 vcm.n517 VSS 1.01f
C2536 vcm.n518 VSS 0.159f
C2537 vcm.n519 VSS 0.242f
C2538 vcm.n520 VSS 0.242f
C2539 vcm.n521 VSS -0.358f
C2540 vcm.n522 VSS 0.404f
C2541 vcm.n523 VSS -0.0298f
C2542 vcm.n524 VSS -0.341f
C2543 vcm.n525 VSS -0.288f
C2544 vcm.n526 VSS -0.358f
C2545 vcm.t65 VSS 7.38f
C2546 vcm.n527 VSS 2.37f
C2547 vcm.n528 VSS 1.01f
C2548 vcm.n529 VSS 0.159f
C2549 vcm.n530 VSS 0.242f
C2550 vcm.n531 VSS 0.242f
C2551 vcm.n532 VSS -0.358f
C2552 vcm.n533 VSS 0.404f
C2553 vcm.n534 VSS -0.0298f
C2554 vcm.n535 VSS -0.341f
C2555 vcm.n536 VSS -0.288f
C2556 vcm.n537 VSS -0.358f
C2557 vcm.n538 VSS 2.37f
C2558 vcm.n539 VSS 1.01f
C2559 vcm.n540 VSS 0.159f
C2560 vcm.n541 VSS 0.242f
C2561 vcm.n542 VSS 0.242f
C2562 vcm.n543 VSS -0.358f
C2563 vcm.n544 VSS 0.404f
C2564 vcm.n545 VSS -0.0298f
C2565 vcm.n546 VSS -0.341f
C2566 vcm.n547 VSS -0.288f
C2567 vcm.n548 VSS -0.358f
C2568 vcm.n549 VSS 2.37f
C2569 vcm.n550 VSS 1.01f
C2570 vcm.n551 VSS 0.159f
C2571 vcm.n552 VSS 0.242f
C2572 vcm.n553 VSS 0.242f
C2573 vcm.n554 VSS -0.358f
C2574 vcm.n555 VSS 0.404f
C2575 vcm.n556 VSS -0.0297f
C2576 vcm.n557 VSS -0.341f
C2577 vcm.n558 VSS -0.288f
C2578 vcm.n559 VSS -0.399f
C2579 vcm.n560 VSS 0.0568f
C2580 vcm.n561 VSS 0.19f
C2581 vcm.n562 VSS 0.211f
C2582 vcm.n563 VSS 0.0445f
C2583 vcm.n564 VSS 0.0445f
C2584 vcm.n566 VSS 0.0527f
C2585 vcm.n567 VSS 0.0394f
C2586 vcm.n568 VSS 0.0394f
C2587 vcm.n570 VSS 0.146f
C2588 vcm.n572 VSS 0.952f
C2589 vcm.n573 VSS 0.952f
C2590 vcm.n574 VSS 0.146f
C2591 vcm.n576 VSS 0.0527f
C2592 vcm.n577 VSS 0.0394f
C2593 vcm.n578 VSS 0.0394f
C2594 vcm.t48 VSS 7.39f
C2595 vcm.n579 VSS 0.404f
C2596 vcm.n580 VSS -0.0298f
C2597 vcm.n581 VSS -0.341f
C2598 vcm.n582 VSS 0.404f
C2599 vcm.n583 VSS -0.0297f
C2600 vcm.n584 VSS -0.341f
C2601 vcm.n585 VSS 2.37f
C2602 vcm.n586 VSS 2.38f
C2603 vcm.t47 VSS 7.39f
C2604 vcm.n587 VSS 0.404f
C2605 vcm.n588 VSS -0.0298f
C2606 vcm.n589 VSS -0.341f
C2607 vcm.n590 VSS 0.404f
C2608 vcm.n591 VSS -0.0297f
C2609 vcm.n592 VSS -0.341f
C2610 vcm.n593 VSS 2.37f
C2611 vcm.n594 VSS 2.38f
C2612 vcm.t62 VSS 7.39f
C2613 vcm.n595 VSS 0.504f
C2614 vcm.n596 VSS 2.37f
C2615 vcm.n597 VSS 0.251f
C2616 vcm.n598 VSS 0.0571f
C2617 vcm.n599 VSS -0.399f
C2618 vcm.n600 VSS 0.404f
C2619 vcm.n601 VSS -0.0297f
C2620 vcm.n602 VSS -0.341f
C2621 vcm.n603 VSS 0.404f
C2622 vcm.n604 VSS -0.0298f
C2623 vcm.n605 VSS -0.341f
C2624 vcm.n606 VSS -0.288f
C2625 vcm.n607 VSS -0.358f
C2626 vcm.n608 VSS 2.37f
C2627 vcm.n609 VSS 1.01f
C2628 vcm.n610 VSS 0.159f
C2629 vcm.n611 VSS 0.242f
C2630 vcm.n612 VSS 0.242f
C2631 vcm.n613 VSS -0.358f
C2632 vcm.n614 VSS 0.404f
C2633 vcm.n615 VSS -0.0297f
C2634 vcm.n616 VSS -0.341f
C2635 vcm.n617 VSS 0.404f
C2636 vcm.n618 VSS -0.0297f
C2637 vcm.n619 VSS -0.341f
C2638 vcm.n620 VSS -0.288f
C2639 vcm.n621 VSS -0.358f
C2640 vcm.t55 VSS 7.38f
C2641 vcm.n622 VSS 2.37f
C2642 vcm.n623 VSS 1.01f
C2643 vcm.n624 VSS 0.159f
C2644 vcm.n625 VSS 0.242f
C2645 vcm.n626 VSS 0.242f
C2646 vcm.n627 VSS -0.358f
C2647 vcm.n628 VSS -0.288f
C2648 vcm.n629 VSS -0.358f
C2649 vcm.n630 VSS 2.37f
C2650 vcm.n631 VSS 1.01f
C2651 vcm.n632 VSS 0.159f
C2652 vcm.n633 VSS 0.242f
C2653 vcm.n634 VSS 0.242f
C2654 vcm.n635 VSS -0.358f
C2655 vcm.n636 VSS 0.404f
C2656 vcm.n637 VSS -0.0297f
C2657 vcm.n638 VSS -0.341f
C2658 vcm.n639 VSS 0.404f
C2659 vcm.n640 VSS -0.0297f
C2660 vcm.n641 VSS -0.341f
C2661 vcm.n642 VSS -0.288f
C2662 vcm.n643 VSS -0.358f
C2663 vcm.t56 VSS 7.38f
C2664 vcm.n644 VSS 2.37f
C2665 vcm.n645 VSS 1.01f
C2666 vcm.n646 VSS 0.159f
C2667 vcm.n647 VSS 0.242f
C2668 vcm.n648 VSS 0.242f
C2669 vcm.n649 VSS -0.358f
C2670 vcm.n650 VSS -0.288f
C2671 vcm.n651 VSS -0.38f
C2672 vcm.n652 VSS 2.37f
C2673 vcm.n653 VSS 0.504f
C2674 vcm.n654 VSS 0.193f
C2675 vcm.n655 VSS 0.175f
C2676 vcm.n656 VSS 0.185f
C2677 vcm.n657 VSS 0.211f
C2678 vcm.n658 VSS 0.0445f
C2679 vcm.n659 VSS 0.0445f
C2680 vcm.n661 VSS 1.04f
C2681 vcm.n662 VSS 1.04f
C2682 vcm.n663 VSS 0.156f
C2683 vcm.n664 VSS 2.38f
C2684 vcm.t43 VSS 7.39f
C2685 vcm.n665 VSS 0.0142f
C2686 vcm.n666 VSS 2.37f
C2687 vcm.n667 VSS 2.38f
C2688 vcm.t40 VSS 7.39f
C2689 vcm.n668 VSS 0.0142f
C2690 vcm.n669 VSS 2.37f
C2691 vcm.n670 VSS 0.504f
C2692 vcm.n671 VSS 2.38f
C2693 vcm.n672 VSS 0.251f
C2694 vcm.n673 VSS 0.0571f
C2695 vcm.n674 VSS -0.399f
C2696 vcm.n675 VSS 0.13f
C2697 vcm.n676 VSS 1.73f
C2698 vcm.n677 VSS 0.189f
C2699 vcm.n678 VSS -0.135f
C2700 vcm.n679 VSS -0.288f
C2701 vcm.n680 VSS -0.358f
C2702 vcm.t51 VSS 7.38f
C2703 vcm.n681 VSS 2.37f
C2704 vcm.n682 VSS 1.01f
C2705 vcm.n683 VSS 0.159f
C2706 vcm.n684 VSS 0.242f
C2707 vcm.n685 VSS 0.242f
C2708 vcm.n686 VSS -0.358f
C2709 vcm.n687 VSS -0.288f
C2710 vcm.n688 VSS -0.358f
C2711 vcm.n689 VSS 2.37f
C2712 vcm.n690 VSS 1.01f
C2713 vcm.n691 VSS 0.159f
C2714 vcm.n692 VSS 0.242f
C2715 vcm.n693 VSS 0.242f
C2716 vcm.n694 VSS -0.358f
C2717 vcm.n695 VSS 0.0139f
C2718 vcm.n696 VSS -0.288f
C2719 vcm.n697 VSS -0.358f
C2720 vcm.t30 VSS 7.38f
C2721 vcm.n698 VSS 2.37f
C2722 vcm.n699 VSS 1.01f
C2723 vcm.n700 VSS 0.159f
C2724 vcm.n701 VSS 0.242f
C2725 vcm.n702 VSS 0.242f
C2726 vcm.n703 VSS -0.358f
C2727 vcm.n704 VSS -0.288f
C2728 vcm.n705 VSS -0.358f
C2729 vcm.n706 VSS 2.37f
C2730 vcm.n707 VSS 1.01f
C2731 vcm.n708 VSS 0.159f
C2732 vcm.n709 VSS 0.242f
C2733 vcm.n710 VSS 0.242f
C2734 vcm.n711 VSS -0.358f
C2735 vcm.n712 VSS 0.0139f
C2736 vcm.n713 VSS -0.288f
C2737 vcm.n714 VSS -0.38f
C2738 vcm.t33 VSS 7.38f
C2739 vcm.n715 VSS 2.39f
C2740 vcm.n716 VSS 0.331f
C2741 vcm.n717 VSS 0.178f
C2742 vcm.n718 VSS 0.195f
C2743 vcm.n719 VSS 0.211f
C2744 vcm.n720 VSS 0.0445f
C2745 vcm.n721 VSS 0.0445f
C2746 vcm.n723 VSS 0.0527f
C2747 vcm.n724 VSS 0.0394f
C2748 vcm.n725 VSS 0.0394f
C2749 vcm.n727 VSS 0.146f
C2750 vcm.n729 VSS 1.71f
C2751 vcm.n730 VSS 4.37f
C2752 vcm.n731 VSS 2.58f
C2753 vcm.n732 VSS 0.146f
C2754 vcm.n734 VSS 0.0527f
C2755 vcm.n735 VSS 0.0394f
C2756 vcm.n736 VSS 0.0394f
C2757 vcm.n737 VSS 0.506f
C2758 vcm.t76 VSS 7.38f
C2759 vcm.n738 VSS 2.37f
C2760 vcm.n739 VSS 2.38f
C2761 vcm.t82 VSS 7.39f
C2762 vcm.n740 VSS 0.0145f
C2763 vcm.n741 VSS 2.37f
C2764 vcm.t75 VSS 7.39f
C2765 vcm.n742 VSS 0.0145f
C2766 vcm.n743 VSS 2.37f
C2767 vcm.n744 VSS 2.38f
C2768 vcm.t85 VSS 7.39f
C2769 vcm.n745 VSS 0.504f
C2770 vcm.n746 VSS 2.37f
C2771 vcm.n747 VSS 0.251f
C2772 vcm.n748 VSS 0.0571f
C2773 vcm.n749 VSS -0.399f
C2774 vcm.n750 VSS 0.197f
C2775 vcm.n751 VSS 0.0782f
C2776 vcm.t4 VSS 0.00751f
C2777 vcm.t0 VSS 0.00797f
C2778 vcm.n752 VSS 0.0334f
C2779 vcm.t1 VSS 0.00797f
C2780 vcm.n753 VSS 0.0278f
C2781 vcm.t5 VSS 0.00186f
C2782 vcm.n754 VSS 0.0138f
C2783 vcm.t7 VSS 0.00749f
C2784 vcm.t2 VSS 0.00796f
C2785 vcm.n755 VSS 0.0331f
C2786 vcm.t3 VSS 0.00796f
C2787 vcm.n756 VSS 0.0273f
C2788 vcm.t6 VSS 0.00184f
C2789 vcm.n757 VSS 0.0131f
C2790 vcm.n758 VSS 0.0464f
C2791 vcm.n759 VSS 3.39f
C2792 vcm.n760 VSS 0.0769f
C2793 vcm.n761 VSS 1.28f
C2794 vcm.n762 VSS -0.475f
C2795 vcm.n763 VSS 0.0144f
C2796 vcm.n764 VSS 0.0452f
C2797 vcm.n765 VSS -0.178f
C2798 vcm.n766 VSS -0.288f
C2799 vcm.n767 VSS -0.358f
C2800 vcm.n768 VSS 2.37f
C2801 vcm.n769 VSS 1.01f
C2802 vcm.n770 VSS 0.159f
C2803 vcm.n771 VSS 0.242f
C2804 vcm.n772 VSS 0.242f
C2805 vcm.n773 VSS -0.358f
C2806 vcm.n774 VSS 0.0145f
C2807 vcm.n775 VSS -0.288f
C2808 vcm.n776 VSS -0.358f
C2809 vcm.t80 VSS 7.38f
C2810 vcm.n777 VSS 2.37f
C2811 vcm.n778 VSS 1.01f
C2812 vcm.n779 VSS 0.159f
C2813 vcm.n780 VSS 0.242f
C2814 vcm.n781 VSS 0.242f
C2815 vcm.n782 VSS -0.358f
C2816 vcm.n783 VSS -0.288f
C2817 vcm.n784 VSS -0.358f
C2818 vcm.n785 VSS 2.37f
C2819 vcm.n786 VSS 1.01f
C2820 vcm.n787 VSS 0.159f
C2821 vcm.n788 VSS 0.242f
C2822 vcm.n789 VSS 0.242f
C2823 vcm.n790 VSS -0.358f
C2824 vcm.n791 VSS -0.288f
C2825 vcm.n792 VSS -0.358f
C2826 vcm.n793 VSS 2.37f
C2827 vcm.n794 VSS 1.01f
C2828 vcm.n795 VSS 0.149f
C2829 vcm.n796 VSS 0.244f
C2830 vcm.n797 VSS 0.249f
C2831 vcm.n798 VSS -0.358f
C2832 vcm.n799 VSS 0.0145f
C2833 vcm.n800 VSS -0.288f
C2834 vcm.n801 VSS -0.38f
C2835 vcm.n802 VSS 0.193f
C2836 vcm.n803 VSS 0.174f
C2837 vcm.n804 VSS 0.185f
C2838 vcm.n805 VSS 0.211f
C2839 vcm.n806 VSS 0.0445f
C2840 vcm.n807 VSS 0.0445f
C2841 vcm.n809 VSS 1.07f
C2842 vcm.n810 VSS 1.07f
C2843 vcm.n811 VSS 0.243f
C2844 vcm.n812 VSS 0.33f
C2845 vcm.t64 VSS 7.38f
C2846 vcm.n813 VSS 2.39f
C2847 vcm.n814 VSS 2.38f
C2848 vcm.t71 VSS 7.39f
C2849 vcm.n815 VSS 2.37f
C2850 vcm.t63 VSS 7.39f
C2851 vcm.n816 VSS 2.37f
C2852 vcm.t69 VSS 7.39f
C2853 vcm.n817 VSS 0.405f
C2854 vcm.n818 VSS -0.0315f
C2855 vcm.n819 VSS -0.342f
C2856 vcm.n820 VSS 0.428f
C2857 vcm.n821 VSS -0.0316f
C2858 vcm.n822 VSS -0.365f
C2859 vcm.n823 VSS 2.37f
C2860 vcm.n824 VSS 0.504f
C2861 vcm.n825 VSS 2.38f
C2862 vcm.n826 VSS 0.251f
C2863 vcm.n827 VSS 0.0571f
C2864 vcm.n828 VSS -0.399f
C2865 vcm.n829 VSS 0.404f
C2866 vcm.n830 VSS -0.0297f
C2867 vcm.n831 VSS -0.341f
C2868 vcm.n832 VSS 0.404f
C2869 vcm.n833 VSS -0.0297f
C2870 vcm.n834 VSS -0.341f
C2871 vcm.n835 VSS -0.288f
C2872 vcm.n836 VSS -0.358f
C2873 vcm.t78 VSS 7.38f
C2874 vcm.n837 VSS 2.37f
C2875 vcm.n838 VSS 1.01f
C2876 vcm.n839 VSS 0.159f
C2877 vcm.n840 VSS 0.242f
C2878 vcm.n841 VSS 0.242f
C2879 vcm.n842 VSS -0.358f
C2880 vcm.n843 VSS -0.288f
C2881 vcm.n844 VSS -0.358f
C2882 vcm.n845 VSS 2.37f
C2883 vcm.n846 VSS 1.01f
C2884 vcm.n847 VSS 0.159f
C2885 vcm.n848 VSS 0.242f
C2886 vcm.n849 VSS 0.242f
C2887 vcm.n850 VSS -0.358f
C2888 vcm.n851 VSS 0.404f
C2889 vcm.n852 VSS -0.0297f
C2890 vcm.n853 VSS -0.341f
C2891 vcm.n854 VSS 0.405f
C2892 vcm.n855 VSS -0.0315f
C2893 vcm.n856 VSS -0.342f
C2894 vcm.n857 VSS -0.288f
C2895 vcm.n858 VSS -0.358f
C2896 vcm.n859 VSS 2.37f
C2897 vcm.n860 VSS 1.01f
C2898 vcm.n861 VSS 0.149f
C2899 vcm.n862 VSS 0.244f
C2900 vcm.n863 VSS 0.249f
C2901 vcm.n864 VSS -0.358f
C2902 vcm.n865 VSS 0.404f
C2903 vcm.n866 VSS -0.0297f
C2904 vcm.n867 VSS -0.341f
C2905 vcm.n868 VSS 0.405f
C2906 vcm.n869 VSS -0.0298f
C2907 vcm.n870 VSS -0.341f
C2908 vcm.n871 VSS -0.288f
C2909 vcm.n872 VSS -0.358f
C2910 vcm.n873 VSS 2.37f
C2911 vcm.n874 VSS 1.01f
C2912 vcm.n875 VSS 0.159f
C2913 vcm.n876 VSS 0.242f
C2914 vcm.n877 VSS 0.242f
C2915 vcm.n878 VSS -0.358f
C2916 vcm.n879 VSS 0.428f
C2917 vcm.n880 VSS -0.0316f
C2918 vcm.n881 VSS -0.365f
C2919 vcm.n882 VSS 0.405f
C2920 vcm.n883 VSS -0.0315f
C2921 vcm.n884 VSS -0.342f
C2922 vcm.n885 VSS -0.288f
C2923 vcm.n886 VSS -0.399f
C2924 vcm.n887 VSS 0.0564f
C2925 vcm.n888 VSS 0.19f
C2926 vcm.n889 VSS 0.211f
C2927 vcm.n890 VSS 0.0445f
C2928 vcm.n891 VSS 0.0445f
C2929 vcm.n893 VSS 0.0527f
C2930 vcm.n894 VSS 0.0394f
C2931 vcm.n895 VSS 0.0394f
C2932 vcm.n897 VSS 0.146f
C2933 vcm.n899 VSS 0.985f
C2934 vcm.n900 VSS 0.985f
C2935 vcm.n901 VSS 0.146f
C2936 vcm.n903 VSS 0.0527f
C2937 vcm.n904 VSS 0.0394f
C2938 vcm.n905 VSS 0.0394f
C2939 vcm.n906 VSS 0.332f
C2940 vcm.t12 VSS 7.38f
C2941 vcm.n907 VSS 2.39f
C2942 vcm.n908 VSS 2.38f
C2943 vcm.t19 VSS 7.39f
C2944 vcm.n909 VSS 2.37f
C2945 vcm.t11 VSS 7.39f
C2946 vcm.n910 VSS 2.37f
C2947 vcm.t17 VSS 7.39f
C2948 vcm.n911 VSS 2.37f
C2949 vcm.t25 VSS 7.38f
C2950 vcm.n912 VSS 0.504f
C2951 vcm.n913 VSS 2.38f
C2952 vcm.n914 VSS 0.251f
C2953 vcm.n915 VSS 0.0571f
C2954 vcm.n916 VSS -0.399f
C2955 vcm.n917 VSS -0.288f
C2956 vcm.n918 VSS -0.358f
C2957 vcm.n919 VSS 2.37f
C2958 vcm.n920 VSS 1.01f
C2959 vcm.n921 VSS 0.159f
C2960 vcm.n922 VSS 0.242f
C2961 vcm.n923 VSS 0.242f
C2962 vcm.n924 VSS -0.358f
C2963 vcm.n925 VSS -0.288f
C2964 vcm.n926 VSS -0.358f
C2965 vcm.n927 VSS 2.37f
C2966 vcm.n928 VSS 1.01f
C2967 vcm.n929 VSS 0.149f
C2968 vcm.n930 VSS 0.244f
C2969 vcm.n931 VSS 0.249f
C2970 vcm.n932 VSS -0.358f
C2971 vcm.n933 VSS -0.288f
C2972 vcm.n934 VSS -0.358f
C2973 vcm.n935 VSS 2.37f
C2974 vcm.n936 VSS 1.01f
C2975 vcm.n937 VSS 0.159f
C2976 vcm.n938 VSS 0.242f
C2977 vcm.n939 VSS 0.242f
C2978 vcm.n940 VSS -0.358f
C2979 vcm.n941 VSS -0.288f
C2980 vcm.n942 VSS -0.358f
C2981 vcm.n943 VSS 2.37f
C2982 vcm.n944 VSS 1.01f
C2983 vcm.n945 VSS 0.159f
C2984 vcm.n946 VSS 0.242f
C2985 vcm.n947 VSS 0.242f
C2986 vcm.n948 VSS -0.358f
C2987 vcm.n949 VSS -0.288f
C2988 vcm.n950 VSS -0.38f
C2989 vcm.n951 VSS 0.156f
C2990 vcm.n952 VSS 0.177f
C2991 vcm.n953 VSS 0.194f
C2992 vcm.n954 VSS 0.211f
C2993 vcm.n955 VSS 0.0445f
C2994 vcm.n956 VSS 0.0445f
C2995 vcm.n958 VSS 1.01f
C2996 vcm.n959 VSS 1.01f
C2997 vcm.n960 VSS 0.146f
C2998 vcm.n962 VSS 0.332f
C2999 vcm.t83 VSS 7.38f
C3000 vcm.n963 VSS 2.39f
C3001 vcm.n964 VSS 2.38f
C3002 vcm.t9 VSS 7.39f
C3003 vcm.n965 VSS 2.37f
C3004 vcm.t81 VSS 7.39f
C3005 vcm.n966 VSS 0.404f
C3006 vcm.n967 VSS -0.0297f
C3007 vcm.n968 VSS -0.341f
C3008 vcm.n969 VSS 2.37f
C3009 vcm.n970 VSS 2.38f
C3010 vcm.t14 VSS 7.39f
C3011 vcm.n971 VSS 0.504f
C3012 vcm.n972 VSS 2.37f
C3013 vcm.n973 VSS 0.251f
C3014 vcm.n974 VSS 0.0571f
C3015 vcm.n975 VSS -0.399f
C3016 vcm.n976 VSS 0.404f
C3017 vcm.n977 VSS -0.0298f
C3018 vcm.n978 VSS -0.341f
C3019 vcm.n979 VSS -0.288f
C3020 vcm.n980 VSS -0.358f
C3021 vcm.n981 VSS 2.37f
C3022 vcm.n982 VSS 1.01f
C3023 vcm.n983 VSS 0.149f
C3024 vcm.n984 VSS 0.244f
C3025 vcm.n985 VSS 0.249f
C3026 vcm.n986 VSS -0.358f
C3027 vcm.n987 VSS 0.404f
C3028 vcm.n988 VSS -0.0297f
C3029 vcm.n989 VSS -0.341f
C3030 vcm.n990 VSS -0.288f
C3031 vcm.n991 VSS -0.358f
C3032 vcm.t87 VSS 7.38f
C3033 vcm.n992 VSS 2.37f
C3034 vcm.n993 VSS 1.01f
C3035 vcm.n994 VSS 0.159f
C3036 vcm.n995 VSS 0.242f
C3037 vcm.n996 VSS 0.242f
C3038 vcm.n997 VSS -0.358f
C3039 vcm.n998 VSS -0.288f
C3040 vcm.n999 VSS -0.358f
C3041 vcm.n1000 VSS 2.37f
C3042 vcm.n1001 VSS 1.01f
C3043 vcm.n1002 VSS 0.159f
C3044 vcm.n1003 VSS 0.242f
C3045 vcm.n1004 VSS 0.242f
C3046 vcm.n1005 VSS -0.358f
C3047 vcm.n1006 VSS 0.404f
C3048 vcm.n1007 VSS -0.0297f
C3049 vcm.n1008 VSS -0.341f
C3050 vcm.n1009 VSS -0.288f
C3051 vcm.n1010 VSS -0.358f
C3052 vcm.n1011 VSS 2.37f
C3053 vcm.n1012 VSS 1.01f
C3054 vcm.n1013 VSS 0.159f
C3055 vcm.n1014 VSS 0.242f
C3056 vcm.n1015 VSS 0.242f
C3057 vcm.n1016 VSS -0.358f
C3058 vcm.n1017 VSS 0.405f
C3059 vcm.n1018 VSS -0.0315f
C3060 vcm.n1019 VSS -0.342f
C3061 vcm.n1020 VSS -0.288f
C3062 vcm.n1021 VSS -0.38f
C3063 vcm.n1022 VSS 0.156f
C3064 vcm.n1023 VSS 0.177f
C3065 vcm.n1024 VSS 0.194f
C3066 vcm.n1025 VSS 0.211f
C3067 vcm.n1026 VSS 0.0445f
C3068 vcm.n1027 VSS 0.0445f
C3069 vcm.n1029 VSS 0.995f
C3070 vcm.t32 VSS 7.39f
C3071 vcm.n1030 VSS 0.177f
C3072 vcm.n1031 VSS 0.193f
C3073 vcm.n1032 VSS 0.428f
C3074 vcm.n1033 VSS -0.0316f
C3075 vcm.n1034 VSS -0.365f
C3076 vcm.n1035 VSS 2.37f
C3077 vcm.n1036 VSS 2.38f
C3078 vcm.t29 VSS 7.38f
C3079 vcm.n1037 VSS 2.38f
C3080 vcm.t39 VSS 7.39f
C3081 vcm.n1038 VSS 0.404f
C3082 vcm.n1039 VSS -0.0297f
C3083 vcm.n1040 VSS -0.341f
C3084 vcm.n1041 VSS 2.37f
C3085 vcm.n1042 VSS 0.504f
C3086 vcm.n1043 VSS 2.38f
C3087 vcm.n1044 VSS 0.251f
C3088 vcm.n1045 VSS 0.0571f
C3089 vcm.n1046 VSS -0.399f
C3090 vcm.n1047 VSS 0.405f
C3091 vcm.n1048 VSS -0.0315f
C3092 vcm.n1049 VSS -0.342f
C3093 vcm.n1050 VSS -0.288f
C3094 vcm.n1051 VSS -0.358f
C3095 vcm.t50 VSS 7.38f
C3096 vcm.n1052 VSS 2.37f
C3097 vcm.n1053 VSS 1.01f
C3098 vcm.n1054 VSS 0.159f
C3099 vcm.n1055 VSS 0.242f
C3100 vcm.n1056 VSS 0.242f
C3101 vcm.n1057 VSS -0.358f
C3102 vcm.n1058 VSS -0.288f
C3103 vcm.n1059 VSS -0.358f
C3104 vcm.n1060 VSS 2.37f
C3105 vcm.n1061 VSS 1.01f
C3106 vcm.n1062 VSS 0.159f
C3107 vcm.n1063 VSS 0.242f
C3108 vcm.n1064 VSS 0.242f
C3109 vcm.n1065 VSS -0.358f
C3110 vcm.n1066 VSS 0.404f
C3111 vcm.n1067 VSS -0.0298f
C3112 vcm.n1068 VSS -0.341f
C3113 vcm.n1069 VSS -0.288f
C3114 vcm.n1070 VSS -0.358f
C3115 vcm.n1071 VSS 2.37f
C3116 vcm.n1072 VSS 1.01f
C3117 vcm.n1073 VSS 0.159f
C3118 vcm.n1074 VSS 0.242f
C3119 vcm.n1075 VSS 0.242f
C3120 vcm.n1076 VSS -0.358f
C3121 vcm.n1077 VSS 0.404f
C3122 vcm.n1078 VSS -0.0297f
C3123 vcm.n1079 VSS -0.341f
C3124 vcm.n1080 VSS -0.288f
C3125 vcm.n1081 VSS -0.358f
C3126 vcm.t42 VSS 7.38f
C3127 vcm.n1082 VSS 2.37f
C3128 vcm.n1083 VSS 1.01f
C3129 vcm.n1084 VSS 0.159f
C3130 vcm.n1085 VSS 0.242f
C3131 vcm.n1086 VSS 0.242f
C3132 vcm.n1087 VSS -0.358f
C3133 vcm.n1088 VSS -0.288f
C3134 vcm.n1089 VSS -0.38f
C3135 vcm.n1090 VSS 2.37f
C3136 vcm.n1091 VSS 0.503f
C3137 vcm.n1092 VSS 0.185f
C3138 vcm.n1093 VSS 0.211f
C3139 vcm.n1094 VSS 0.0445f
C3140 vcm.n1095 VSS 0.0445f
C3141 vcm.n1096 VSS 0.995f
C3142 vcm.n1097 VSS 0.146f
C3143 vcm.n1099 VSS 0.0527f
C3144 vcm.n1100 VSS 0.0394f
C3145 vcm.n1101 VSS 0.0394f
C3146 vcm.n1103 VSS 1.01f
C3147 vcm.n1104 VSS 1.01f
C3148 vcm.n1105 VSS 0.146f
C3149 vcm.n1107 VSS 0.0527f
C3150 vcm.n1108 VSS 0.0394f
C3151 vcm.n1109 VSS 0.0394f
C3152 vcm.n1110 VSS 2.38f
C3153 vcm.n1111 VSS 2.38f
C3154 vcm.t18 VSS 7.39f
C3155 vcm.n1112 VSS 2.37f
C3156 vcm.t26 VSS 7.38f
C3157 vcm.n1113 VSS 2.38f
C3158 vcm.t34 VSS 7.39f
C3159 vcm.n1114 VSS 0.504f
C3160 vcm.n1115 VSS 2.37f
C3161 vcm.n1116 VSS 0.251f
C3162 vcm.n1117 VSS 0.0571f
C3163 vcm.n1118 VSS -0.399f
C3164 vcm.n1119 VSS 0.428f
C3165 vcm.n1120 VSS -0.0316f
C3166 vcm.n1121 VSS -0.365f
C3167 vcm.n1122 VSS -0.288f
C3168 vcm.n1123 VSS -0.358f
C3169 vcm.n1124 VSS 2.37f
C3170 vcm.n1125 VSS 1.01f
C3171 vcm.n1126 VSS 0.159f
C3172 vcm.n1127 VSS 0.242f
C3173 vcm.n1128 VSS 0.242f
C3174 vcm.n1129 VSS -0.358f
C3175 vcm.n1130 VSS 0.404f
C3176 vcm.n1131 VSS -0.0298f
C3177 vcm.n1132 VSS -0.341f
C3178 vcm.n1133 VSS -0.288f
C3179 vcm.n1134 VSS -0.358f
C3180 vcm.n1135 VSS 2.37f
C3181 vcm.n1136 VSS 1.01f
C3182 vcm.n1137 VSS 0.159f
C3183 vcm.n1138 VSS 0.242f
C3184 vcm.n1139 VSS 0.242f
C3185 vcm.n1140 VSS -0.358f
C3186 vcm.n1141 VSS 0.404f
C3187 vcm.n1142 VSS -0.0298f
C3188 vcm.n1143 VSS -0.341f
C3189 vcm.n1144 VSS -0.288f
C3190 vcm.n1145 VSS -0.358f
C3191 vcm.n1146 VSS 2.37f
C3192 vcm.n1147 VSS 1.01f
C3193 vcm.n1148 VSS 0.159f
C3194 vcm.n1149 VSS 0.242f
C3195 vcm.n1150 VSS 0.242f
C3196 vcm.n1151 VSS -0.358f
C3197 vcm.n1152 VSS 0.404f
C3198 vcm.n1153 VSS -0.0298f
C3199 vcm.n1154 VSS -0.341f
C3200 vcm.n1155 VSS -0.288f
C3201 vcm.n1156 VSS -0.358f
C3202 vcm.t27 VSS 7.38f
C3203 vcm.n1157 VSS 2.37f
C3204 vcm.n1158 VSS 1.01f
C3205 vcm.n1159 VSS 0.159f
C3206 vcm.n1160 VSS 0.242f
C3207 vcm.n1161 VSS 0.242f
C3208 vcm.n1162 VSS -0.358f
C3209 vcm.n1163 VSS 0.405f
C3210 vcm.n1164 VSS -0.0315f
C3211 vcm.n1165 VSS -0.342f
C3212 vcm.n1166 VSS -0.288f
C3213 vcm.n1167 VSS 0.177f
C3214 vcm.n1168 VSS 0.193f
C3215 vcm.n1169 VSS -0.38f
C3216 vcm.t20 VSS 7.38f
C3217 vcm.n1170 VSS 2.37f
C3218 vcm.n1171 VSS 0.503f
C3219 vcm.n1172 VSS 0.185f
C3220 vcm.n1173 VSS 0.211f
C3221 vcm.n1174 VSS 0.0445f
C3222 vcm.n1175 VSS 0.0445f
C3223 vcm.n1177 VSS 1.01f
C3224 vcm.n1178 VSS 1.01f
C3225 vcm.n1179 VSS 0.146f
C3226 vcm.n1181 VSS 0.332f
C3227 vcm.t10 VSS 7.39f
C3228 vcm.n1182 VSS 2.39f
C3229 vcm.n1183 VSS -0.38f
C3230 vcm.n1184 VSS 0.156f
C3231 vcm.n1185 VSS 0.177f
C3232 vcm.n1186 VSS 0.194f
C3233 vcm.n1187 VSS 0.211f
C3234 vcm.n1188 VSS 0.0445f
C3235 vcm.n1189 VSS 0.0445f
C3236 vcm.n1191 VSS 1f
C3237 vcm.n1192 VSS 1f
C3238 vcm.n1193 VSS 0.0445f
C3239 vcm.n1194 VSS 0.0445f
C3240 vcm.n1195 VSS 0.211f
C3241 vcm.n1196 VSS 0.194f
C3242 vcm.n1197 VSS 0.177f
.ends

