magic
tech sky130A
magscale 1 2
timestamp 1698671014
<< error_p >>
rect -77 -89 -19 -83
rect -77 -123 -65 -89
rect -77 -129 -19 -123
<< nwell >>
rect -161 -79 161 91
<< pmoshvt >>
rect -63 -42 -33 42
rect 33 -42 63 42
<< pdiff >>
rect -125 30 -63 42
rect -125 -30 -113 30
rect -79 -30 -63 30
rect -125 -42 -63 -30
rect -33 30 33 42
rect -33 -30 -17 30
rect 17 -30 33 30
rect -33 -42 33 -30
rect 63 30 125 42
rect 63 -30 79 30
rect 113 -30 125 30
rect 63 -42 125 -30
<< pdiffc >>
rect -113 -30 -79 30
rect -17 -30 17 30
rect 79 -30 113 30
<< poly >>
rect -63 42 -33 68
rect 33 42 63 68
rect -63 -57 -33 -42
rect 33 -57 63 -42
rect -63 -73 63 -57
rect -81 -87 63 -73
rect -81 -89 -15 -87
rect -81 -123 -65 -89
rect -31 -123 -15 -89
rect -81 -139 -15 -123
<< polycont >>
rect -65 -123 -31 -89
<< locali >>
rect -113 30 -79 46
rect -113 -46 -79 -30
rect -17 30 17 84
rect -17 -46 17 -30
rect 79 30 113 46
rect 79 -46 113 -30
rect -81 -123 -65 -89
rect -31 -123 -15 -89
<< viali >>
rect -113 -30 -79 30
rect 79 -30 113 30
rect -65 -123 -31 -89
<< metal1 >>
rect -119 30 119 42
rect -119 -30 -113 30
rect -79 -30 79 30
rect 113 -30 119 30
rect -119 -42 119 -30
rect -77 -89 -19 -83
rect -77 -123 -65 -89
rect -31 -123 -19 -89
rect -77 -129 -19 -123
<< properties >>
string FIXED_BBOX -210 -208 210 208
string gencell sky130_fd_pr__pfet_01v8_hvt
string library sky130
string parameters w 0.42 l 0.15 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
