magic
tech sky130A
magscale 1 2
timestamp 1706706162
<< nwell >>
rect 116 1874 1020 1994
rect 460 678 494 680
rect 552 678 586 680
rect 644 678 678 680
rect 392 606 1020 678
<< psubdiff >>
rect 154 1310 982 1326
rect 154 1308 644 1310
rect 154 1306 554 1308
rect 154 1304 274 1306
rect 154 1270 186 1304
rect 220 1272 274 1304
rect 308 1302 458 1306
rect 308 1272 368 1302
rect 220 1270 368 1272
rect 154 1268 368 1270
rect 402 1272 458 1302
rect 492 1274 554 1306
rect 588 1276 644 1308
rect 678 1308 982 1310
rect 678 1276 740 1308
rect 588 1274 740 1276
rect 774 1306 982 1308
rect 774 1274 832 1306
rect 492 1272 832 1274
rect 866 1304 982 1306
rect 866 1272 920 1304
rect 402 1270 920 1272
rect 954 1270 982 1304
rect 402 1268 982 1270
rect 154 1246 982 1268
<< nsubdiff >>
rect 154 1940 982 1950
rect 154 1938 556 1940
rect 154 1904 184 1938
rect 218 1936 462 1938
rect 218 1904 276 1936
rect 154 1902 276 1904
rect 310 1902 366 1936
rect 400 1904 462 1936
rect 496 1906 556 1938
rect 590 1938 826 1940
rect 590 1906 646 1938
rect 496 1904 646 1906
rect 680 1904 736 1938
rect 770 1906 826 1938
rect 860 1938 982 1940
rect 860 1906 918 1938
rect 770 1904 918 1906
rect 952 1904 982 1938
rect 400 1902 982 1904
rect 154 1896 982 1902
rect 430 646 460 680
rect 494 646 552 680
rect 586 646 644 680
rect 678 678 982 680
rect 678 646 734 678
rect 430 644 734 646
rect 768 644 826 678
rect 860 644 918 678
rect 952 644 982 678
<< psubdiffcont >>
rect 186 1270 220 1304
rect 274 1272 308 1306
rect 368 1268 402 1302
rect 458 1272 492 1306
rect 554 1274 588 1308
rect 644 1276 678 1310
rect 740 1274 774 1308
rect 832 1272 866 1306
rect 920 1270 954 1304
<< nsubdiffcont >>
rect 184 1904 218 1938
rect 276 1902 310 1936
rect 366 1902 400 1936
rect 462 1904 496 1938
rect 556 1906 590 1940
rect 646 1904 680 1938
rect 736 1904 770 1938
rect 826 1906 860 1940
rect 918 1904 952 1938
rect 460 646 494 680
rect 552 646 586 680
rect 644 646 678 680
rect 734 644 768 678
rect 826 644 860 678
rect 918 644 952 678
<< locali >>
rect 154 1940 982 1950
rect 154 1938 556 1940
rect 154 1904 184 1938
rect 218 1936 462 1938
rect 218 1904 276 1936
rect 154 1902 276 1904
rect 310 1902 366 1936
rect 400 1904 462 1936
rect 496 1906 556 1938
rect 590 1938 826 1940
rect 590 1906 646 1938
rect 496 1904 646 1906
rect 680 1904 736 1938
rect 770 1906 826 1938
rect 860 1938 982 1940
rect 860 1906 918 1938
rect 770 1904 918 1906
rect 952 1904 982 1938
rect 400 1902 982 1904
rect 154 1894 982 1902
rect 608 1552 790 1592
rect 154 1310 982 1326
rect 154 1308 644 1310
rect 154 1306 554 1308
rect 154 1304 274 1306
rect 154 1270 186 1304
rect 220 1272 274 1304
rect 308 1302 458 1306
rect 308 1272 368 1302
rect 220 1270 368 1272
rect 154 1268 368 1270
rect 402 1272 458 1302
rect 492 1274 554 1306
rect 588 1276 644 1308
rect 678 1308 982 1310
rect 678 1276 740 1308
rect 588 1274 740 1276
rect 774 1306 982 1308
rect 774 1274 832 1306
rect 492 1272 832 1274
rect 866 1304 982 1306
rect 866 1272 920 1304
rect 402 1270 920 1272
rect 954 1270 982 1304
rect 402 1268 982 1270
rect 154 1246 982 1268
rect 598 978 806 1018
rect 430 646 460 680
rect 494 646 552 680
rect 586 646 644 680
rect 678 678 982 680
rect 678 646 734 678
rect 430 644 734 646
rect 768 644 826 678
rect 860 644 918 678
rect 952 644 982 678
<< viali >>
rect 276 1696 310 1730
rect 184 1552 218 1586
rect 360 1560 394 1594
rect 508 1558 542 1592
rect 876 1556 910 1590
rect 496 980 530 1014
rect 872 980 906 1014
<< metal1 >>
rect 974 1832 1278 1946
rect 258 1740 328 1756
rect 258 1730 552 1740
rect 258 1696 276 1730
rect 310 1696 552 1730
rect 258 1690 552 1696
rect 258 1682 328 1690
rect 66 1586 238 1602
rect 66 1552 184 1586
rect 218 1552 238 1586
rect 66 1536 238 1552
rect 342 1598 408 1606
rect 500 1598 552 1690
rect 342 1546 348 1598
rect 400 1546 408 1598
rect 494 1592 558 1598
rect 494 1558 508 1592
rect 542 1558 558 1592
rect 494 1546 558 1558
rect 854 1592 932 1602
rect 342 1542 408 1546
rect 854 1540 868 1592
rect 920 1540 932 1592
rect 854 1536 932 1540
rect 106 1190 442 1382
rect 458 1272 492 1306
rect 554 1274 588 1308
rect 644 1276 678 1310
rect 740 1274 774 1308
rect 832 1272 866 1306
rect 854 1026 922 1030
rect 144 1024 542 1026
rect 144 972 352 1024
rect 404 1014 542 1024
rect 404 980 496 1014
rect 530 980 542 1014
rect 404 972 542 980
rect 144 968 542 972
rect 854 974 860 1026
rect 914 974 922 1026
rect 854 968 922 974
rect 144 966 432 968
rect 1076 742 1278 1832
rect 460 646 494 680
rect 552 646 586 680
rect 644 646 678 680
rect 734 644 768 678
rect 972 644 1278 742
<< via1 >>
rect 348 1594 400 1598
rect 348 1560 360 1594
rect 360 1560 394 1594
rect 394 1560 400 1594
rect 348 1546 400 1560
rect 868 1590 920 1592
rect 868 1556 876 1590
rect 876 1556 910 1590
rect 910 1556 920 1590
rect 868 1540 920 1556
rect 352 972 404 1024
rect 860 1014 914 1026
rect 860 980 872 1014
rect 872 980 906 1014
rect 906 980 914 1014
rect 860 974 914 980
<< metal2 >>
rect 342 1598 408 1606
rect 342 1546 348 1598
rect 400 1566 408 1598
rect 854 1592 928 1602
rect 400 1546 414 1566
rect 342 1024 414 1546
rect 342 972 352 1024
rect 404 972 414 1024
rect 342 968 414 972
rect 854 1540 868 1592
rect 920 1540 928 1592
rect 854 1026 928 1540
rect 854 974 860 1026
rect 914 974 928 1026
rect 854 968 928 974
use sky130_fd_sc_hd__inv_1  x1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 430 0 1 1334
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x2
timestamp 1701704242
transform 1 0 706 0 1 1334
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x3
timestamp 1701704242
transform -1 0 982 0 -1 1238
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x4
timestamp 1701704242
transform -1 0 706 0 -1 1238
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  x5 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 430 0 1 1334
box -38 -48 314 592
<< labels >>
flabel metal1 144 966 352 1026 0 FreeSans 320 0 0 0 ring_osil
port 1 nsew
flabel metal1 1076 644 1278 1946 0 FreeSans 320 0 0 0 vdd
port 2 nsew
flabel space 106 1190 459 1382 0 FreeSans 320 0 0 0 gnd
port 4 nsew
flabel metal1 66 1536 184 1602 0 FreeSans 320 0 0 0 en
port 0 nsew
<< end >>
