** sch_path: /foss/designs/hgu_goss/hgu/xschem/hgu_top_block.sch
.subckt hgu_top_block VDD VSS
+ result[0],result[1],result[2],result[3],result[4],result[5],result[6],result[7] EXT_CLK vip vin sel_bit[0],sel_bit[1]
+ sample_delay_cap_ctrl_code[0],sample_delay_cap_ctrl_code[1],sample_delay_cap_ctrl_code[2],sample_delay_cap_ctrl_code[3],sample_delay_cap_ctrl_code[4],sample_delay_cap_ctrl_code[5],sample_delay_cap_ctrl_code[6],sample_delay_cap_ctrl_code[7],sample_delay_cap_ctrl_code[8],sample_delay_cap_ctrl_code[9],sample_delay_cap_ctrl_code[10],sample_delay_cap_ctrl_code[11],sample_delay_cap_ctrl_code[12],sample_delay_cap_ctrl_code[13],sample_delay_cap_ctrl_code[14],sample_delay_cap_ctrl_code[15]
+ async_resetb_delay_cap_ctrl_code[0],async_resetb_delay_cap_ctrl_code[1],async_resetb_delay_cap_ctrl_code[2],async_resetb_delay_cap_ctrl_code[3]
+ async_setb_delay_cap_ctrl_code[0],async_setb_delay_cap_ctrl_code[1],async_setb_delay_cap_ctrl_code[2],async_setb_delay_cap_ctrl_code[3] async_delay_offset sample_delay_offset
+ retimer_delay_code[0],retimer_delay_code[1],retimer_delay_code[2],retimer_delay_code[3] retimer_delay_offset
*.ipin VDD
*.ipin VSS
*.opin result[0],result[1],result[2],result[3],result[4],result[5],result[6],result[7]
*.ipin EXT_CLK
*.ipin vip
*.ipin vin
*.ipin sel_bit[0],sel_bit[1]
*.ipin
*+ sample_delay_cap_ctrl_code[0],sample_delay_cap_ctrl_code[1],sample_delay_cap_ctrl_code[2],sample_delay_cap_ctrl_code[3],sample_delay_cap_ctrl_code[4],sample_delay_cap_ctrl_code[5],sample_delay_cap_ctrl_code[6],sample_delay_cap_ctrl_code[7],sample_delay_cap_ctrl_code[8],sample_delay_cap_ctrl_code[9],sample_delay_cap_ctrl_code[10],sample_delay_cap_ctrl_code[11],sample_delay_cap_ctrl_code[12],sample_delay_cap_ctrl_code[13],sample_delay_cap_ctrl_code[14],sample_delay_cap_ctrl_code[15]
*.ipin
*+ async_resetb_delay_cap_ctrl_code[0],async_resetb_delay_cap_ctrl_code[1],async_resetb_delay_cap_ctrl_code[2],async_resetb_delay_cap_ctrl_code[3]
*.ipin
*+ async_setb_delay_cap_ctrl_code[0],async_setb_delay_cap_ctrl_code[1],async_setb_delay_cap_ctrl_code[2],async_setb_delay_cap_ctrl_code[3]
*.ipin async_delay_offset
*.ipin sample_delay_offset
*.ipin retimer_delay_code[0],retimer_delay_code[1],retimer_delay_code[2],retimer_delay_code[3]
*.ipin retimer_delay_offset
x1 sar_clk result[0] result[1] result[2] result[3] result[4] result[5] result[6] result[7]
+ sample_clk sel_bit[0] sel_bit[1] sample_clk_b VDD VSS EXT_CLK COMP_RESULT result_sw[1] result_sw[2]
+ result_sw[3] result_sw[4] result_sw[5] result_sw[6] result_sw[7] READY result_sw_b[1] result_sw_b[2]
+ result_sw_b[3] result_sw_b[4] result_sw_b[5] result_sw_b[6] result_sw_b[7] result2_sw[1] result2_sw[2]
+ result2_sw[3] result2_sw[4] result2_sw[5] result2_sw[6] result2_sw[7] result2_sw_b[1] result2_sw_b[2]
+ result2_sw_b[3] result2_sw_b[4] result2_sw_b[5] result2_sw_b[6] result2_sw_b[7] sample_delay_cap_ctrl_code[0]
+ sample_delay_cap_ctrl_code[1] sample_delay_cap_ctrl_code[2] sample_delay_cap_ctrl_code[3] sample_delay_cap_ctrl_code[4]
+ sample_delay_cap_ctrl_code[5] sample_delay_cap_ctrl_code[6] sample_delay_cap_ctrl_code[7] sample_delay_cap_ctrl_code[8]
+ sample_delay_cap_ctrl_code[9] sample_delay_cap_ctrl_code[10] sample_delay_cap_ctrl_code[11] sample_delay_cap_ctrl_code[12]
+ sample_delay_cap_ctrl_code[13] sample_delay_cap_ctrl_code[14] sample_delay_cap_ctrl_code[15] async_resetb_delay_cap_ctrl_code[0]
+ async_resetb_delay_cap_ctrl_code[1] async_resetb_delay_cap_ctrl_code[2] async_resetb_delay_cap_ctrl_code[3]
+ async_setb_delay_cap_ctrl_code[0] async_setb_delay_cap_ctrl_code[1] async_setb_delay_cap_ctrl_code[2]
+ async_setb_delay_cap_ctrl_code[3] async_delay_offset sample_delay_offset retimer_delay_offset retimer_delay_code[0]
+ retimer_delay_code[1] retimer_delay_code[2] retimer_delay_code[3] hgu_sarlogic
x2 READY tah_vn COMP_RESULT net11 tah_vp sar_clk VDD VSS hgu_comp
x3 sw5 swd4 sw3 result_sw[2] swd2 sw2 swd6 swd5 result_sw[1] sw4 sw6 result2_sw[2] result2_sw[1]
+ swd3 VSS VREF tah_vp tah_vp tah_vp tah_vp tah_vp tah_vp tah_vp tah_vp tah_vp tah_vp tah_vp tah_vp tah_vp
+ tah_vp VDD hgu_cdac_half
x4 net4 net8 net2 result_sw_b[2] net10 net1 net6 net7 result_sw_b[1] net3 net5 result2_sw_b[2]
+ result2_sw_b[1] net9 VSS VREF tah_vn tah_vn tah_vn tah_vn tah_vn tah_vn tah_vn tah_vn tah_vn tah_vn tah_vn tah_vn
+ tah_vn tah_vn VDD hgu_cdac_half
x21 sample_clk VDD VSS sample_clk_b tah_vp vip vin tah_vn hgu_tah_flat
x6 result2_sw[3] result2_sw[6] result2_sw[4] result2_sw[5] result2_sw[7] sw2 sw5 sw3 sw4 sw6 VDD VSS
+ hgu_cdac_sw_buffer
x7 result_sw[3] result_sw[6] result_sw[4] result_sw[5] result_sw[7] swd2 swd5 swd3 swd4 swd6 VDD VSS
+ hgu_cdac_sw_buffer
x8 result2_sw_b[3] result2_sw_b[6] result2_sw_b[4] result2_sw_b[5] result2_sw_b[7] net1 net4 net2
+ net3 net5 VDD VSS hgu_cdac_sw_buffer
x9 result_sw_b[3] result_sw_b[6] result_sw_b[4] result_sw_b[5] result_sw_b[7] net10 net7 net9 net8
+ net6 VDD VSS hgu_cdac_sw_buffer
V1 VREF GND 0.9
.save i(v1)
**.ends

* expanding   symbol:  ../xschem/hgu_sarlogic.sym # of pins=21
** sym_path: /foss/designs/hgu_goss/hgu/xschem/hgu_sarlogic.sym
** sch_path: /foss/designs/hgu_goss/hgu/xschem/hgu_sarlogic.sch
.subckt hgu_sarlogic sar_clk sar_result[0] sar_result[1] sar_result[2] sar_result[3] sar_result[4]
+ sar_result[5] sar_result[6] sar_result[7] sample_clk sel_bit[0] sel_bit[1] sample_clk_b VDD VSS EXT_CLK
+ COMP_RESULT vdd_sw[1] vdd_sw[2] vdd_sw[3] vdd_sw[4] vdd_sw[5] vdd_sw[6] vdd_sw[7] READY vdd_sw_b[1] vdd_sw_b[2]
+ vdd_sw_b[3] vdd_sw_b[4] vdd_sw_b[5] vdd_sw_b[6] vdd_sw_b[7] vss_sw[1] vss_sw[2] vss_sw[3] vss_sw[4] vss_sw[5]
+ vss_sw[6] vss_sw[7] vss_sw_b[1] vss_sw_b[2] vss_sw_b[3] vss_sw_b[4] vss_sw_b[5] vss_sw_b[6] vss_sw_b[7]
+ sample_delay_cap_ctrl_code[0] sample_delay_cap_ctrl_code[1] sample_delay_cap_ctrl_code[2] sample_delay_cap_ctrl_code[3]
+ sample_delay_cap_ctrl_code[4] sample_delay_cap_ctrl_code[5] sample_delay_cap_ctrl_code[6] sample_delay_cap_ctrl_code[7]
+ sample_delay_cap_ctrl_code[8] sample_delay_cap_ctrl_code[9] sample_delay_cap_ctrl_code[10] sample_delay_cap_ctrl_code[11]
+ sample_delay_cap_ctrl_code[12] sample_delay_cap_ctrl_code[13] sample_delay_cap_ctrl_code[14] sample_delay_cap_ctrl_code[15]
+ async_resetb_delay_cap_ctrl_code[0] async_resetb_delay_cap_ctrl_code[1] async_resetb_delay_cap_ctrl_code[2]
+ async_resetb_delay_cap_ctrl_code[3] async_setb_delay_cap_ctrl_code[0] async_setb_delay_cap_ctrl_code[1]
+ async_setb_delay_cap_ctrl_code[2] async_setb_delay_cap_ctrl_code[3] async_delay_offset sample_delay_offset retimer_eob_delay_offset
+ retimer_delay_code[0] retimer_delay_code[1] retimer_delay_code[2] retimer_delay_code[3]
*.ipin VDD
*.ipin VSS
*.ipin COMP_RESULT
*.ipin READY
*.ipin EXT_CLK
*.opin sar_clk
*.opin
*+ sar_result[0],sar_result[1],sar_result[2],sar_result[3],sar_result[4],sar_result[5],sar_result[6],sar_result[7]
*.opin sample_clk
*.ipin sel_bit[0],sel_bit[1]
*.ipin
*+ sample_delay_cap_ctrl_code[0],sample_delay_cap_ctrl_code[1],sample_delay_cap_ctrl_code[2],sample_delay_cap_ctrl_code[3],sample_delay_cap_ctrl_code[4],sample_delay_cap_ctrl_code[5],sample_delay_cap_ctrl_code[6],sample_delay_cap_ctrl_code[7],sample_delay_cap_ctrl_code[8],sample_delay_cap_ctrl_code[9],sample_delay_cap_ctrl_code[10],sample_delay_cap_ctrl_code[11],sample_delay_cap_ctrl_code[12],sample_delay_cap_ctrl_code[13],sample_delay_cap_ctrl_code[14],sample_delay_cap_ctrl_code[15]
*.opin sample_clk_b
*.opin vdd_sw[1],vdd_sw[2],vdd_sw[3],vdd_sw[4],vdd_sw[5],vdd_sw[6],vdd_sw[7]
*.opin vdd_sw_b[1],vdd_sw_b[2],vdd_sw_b[3],vdd_sw_b[4],vdd_sw_b[5],vdd_sw_b[6],vdd_sw_b[7]
*.opin vss_sw[1],vss_sw[2],vss_sw[3],vss_sw[4],vss_sw[5],vss_sw[6],vss_sw[7]
*.opin vss_sw_b[1],vss_sw_b[2],vss_sw_b[3],vss_sw_b[4],vss_sw_b[5],vss_sw_b[6],vss_sw_b[7]
*.ipin
*+ async_resetb_delay_cap_ctrl_code[0],async_resetb_delay_cap_ctrl_code[1],async_resetb_delay_cap_ctrl_code[2],async_resetb_delay_cap_ctrl_code[3]
*.ipin
*+ async_setb_delay_cap_ctrl_code[0],async_setb_delay_cap_ctrl_code[1],async_setb_delay_cap_ctrl_code[2],async_setb_delay_cap_ctrl_code[3]
*.ipin async_delay_offset
*.ipin sample_delay_offset
*.ipin retimer_delay_code[0],retimer_delay_code[1],retimer_delay_code[2],retimer_delay_code[3]
*.ipin retimer_eob_delay_offset
x1 sar_clk VDD VSS sample_clk EOB READY async_delay_offset async_resetb_delay_cap_ctrl_code[0]
+ async_resetb_delay_cap_ctrl_code[1] async_resetb_delay_cap_ctrl_code[2] async_resetb_delay_cap_ctrl_code[3]
+ async_setb_delay_cap_ctrl_code[0] async_setb_delay_cap_ctrl_code[1] async_setb_delay_cap_ctrl_code[2]
+ async_setb_delay_cap_ctrl_code[3] hgu_clk_async
x2 sample_clk_b VDD VSS EXT_CLK VSS VSS sample_clk sample_delay_cap_ctrl_code[0]
+ sample_delay_cap_ctrl_code[1] sample_delay_cap_ctrl_code[2] sample_delay_cap_ctrl_code[3] sample_delay_cap_ctrl_code[4]
+ sample_delay_cap_ctrl_code[5] sample_delay_cap_ctrl_code[6] sample_delay_cap_ctrl_code[7] sample_delay_cap_ctrl_code[8]
+ sample_delay_cap_ctrl_code[9] sample_delay_cap_ctrl_code[10] sample_delay_cap_ctrl_code[11] sample_delay_cap_ctrl_code[12]
+ sample_delay_cap_ctrl_code[13] sample_delay_cap_ctrl_code[14] sample_delay_cap_ctrl_code[15] sample_delay_offset hgu_clk_sample
x3 sel_bit[0] sel_bit[1] EOB sar_clk sar_result_temp[0] sar_result_temp[1] sar_result_temp[2]
+ sar_result_temp[3] sar_result_temp[4] sar_result_temp[5] sar_result_temp[6] sar_result_temp[7] COMP_RESULT check[0]
+ check[1] check[2] check[3] check[4] check[5] check[6] sample_clk_b VDD VSS hgu_sarlogic_8bit_logic
x4 VDD VSS vdd_sw[1] vdd_sw[2] vdd_sw[3] vdd_sw[4] vdd_sw[5] vdd_sw[6] vdd_sw[7] vdd_sw_b[1]
+ vdd_sw_b[2] vdd_sw_b[3] vdd_sw_b[4] vdd_sw_b[5] vdd_sw_b[6] vdd_sw_b[7] sar_result_temp[1] sar_result_temp[2]
+ sar_result_temp[3] sar_result_temp[4] sar_result_temp[5] sar_result_temp[6] sar_result_temp[7] vss_sw[1] vss_sw[2]
+ vss_sw[3] vss_sw[4] vss_sw[5] vss_sw[6] vss_sw[7] check[0] check[1] check[2] check[3] check[4] check[5]
+ check[6] vss_sw_b[1] vss_sw_b[2] vss_sw_b[3] vss_sw_b[4] vss_sw_b[5] vss_sw_b[6] vss_sw_b[7] sar_clk
+ sample_clk_b hgu_sarlogic_sw_ctrl
x5 VDD VSS sar_result_temp[0] sar_result_temp[1] sar_result_temp[2] sar_result_temp[3]
+ sar_result_temp[4] sar_result_temp[5] sar_result_temp[6] sar_result_temp[7] EOB retimer_delay_code[0]
+ retimer_delay_code[1] retimer_delay_code[2] retimer_delay_code[3] retimer_eob_delay_offset sar_result[0] sar_result[1]
+ sar_result[2] sar_result[3] sar_result[4] sar_result[5] sar_result[6] sar_result[7] hgu_sarlogic_retimer
.ends


* expanding   symbol:  ../xschem/hgu_comp.sym # of pins=8
** sym_path: /foss/designs/hgu_goss/hgu/xschem/hgu_comp.sym
** sch_path: /foss/designs/hgu_goss/hgu/xschem/hgu_comp.sch
.subckt hgu_comp ready cdac_vn comp_outp comp_outn cdac_vp clk VDD VSS
*.ipin cdac_vn
*.ipin cdac_vp
*.ipin VSS
*.ipin VDD
*.ipin clk
*.opin ready
*.opin comp_outp
*.opin comp_outn
XM1 net1 clk VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=4 nf=4 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4 Y X Q VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM5 X Y P VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM6 X Y VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM7 Y X VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM8 X clk VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM9 P clk VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM10 Y clk VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM11 Q clk VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM16 RS_n RS_p VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.84 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM17 RS_p RS_n VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.84 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM19 RS_p Y_inv VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.84 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM23 RS_n X_inv VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.84 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 P cdac_vp net1 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=8 nf=8 ad='int((nf+1)/2) * W / nf * 0.29' as='int((nf+2)/2) * W / nf * 0.29'
+ pd='2*int((nf+1)/2) * (W / nf + 0.29)' ps='2*int((nf+2)/2) * (W / nf + 0.29)' nrd='0.29 / W ' nrs='0.29 / W '
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 Q cdac_vn net1 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=8 nf=8 ad='int((nf+1)/2) * W / nf * 0.29' as='int((nf+2)/2) * W / nf * 0.29'
+ pd='2*int((nf+1)/2) * (W / nf + 0.29)' ps='2*int((nf+2)/2) * (W / nf + 0.29)' nrd='0.29 / W ' nrs='0.29 / W '
+ sa=0 sb=0 sd=0 mult=1 m=1
XM12 X_inv X VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.84 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM13 X_inv X VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM14 X_drive X_inv VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=2.52 nf=3 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM15 X_drive X_inv VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1.38 nf=3 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM18 Y_inv Y VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.84 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM20 Y_inv Y VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM21 Y_drive Y_inv VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=2.52 nf=3 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM22 Y_drive Y_inv VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1.38 nf=3 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM24 net2 Y_drive X_drive VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.84 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM25 net2 X_drive Y_drive VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.84 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM26 net2 Y_drive net3 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.84 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM27 net3 X_drive VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.84 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM28 ready net2 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.84 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM29 ready net2 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM30 net4 RS_p VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.84 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM31 net4 RS_p VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM32 comp_outp net4 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=2.52 nf=3 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM33 comp_outp net4 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1.38 nf=3 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM34 net5 RS_n VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.84 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM35 net5 RS_n VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM36 comp_outn net5 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=2.52 nf=3 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM37 comp_outn net5 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1.38 nf=3 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  ../xschem/hgu_cdac_half.sym # of pins=31
** sym_path: /foss/designs/hgu_goss/hgu/xschem/hgu_cdac_half.sym
** sch_path: /foss/designs/hgu_goss/hgu/xschem/hgu_cdac_half.sch
.subckt hgu_cdac_half d<5> db<4> d<3> db<1> db<2> d<2> db<6> db<5> db<0> d<4> d<6> d<1> d<0> db<3>
+ VSS VREF tb<0> tb<1> tb<2> tb<4> tb<5> tb<6> t<0> tb<3> t<1> t<2> t<3> t<4> t<5> t<6> VDD
*.iopin d<6>
*.iopin d<5>
*.iopin d<4>
*.iopin d<3>
*.iopin d<2>
*.iopin d<1>
*.iopin d<0>
*.iopin db<6>
*.iopin db<5>
*.iopin db<4>
*.iopin db<3>
*.iopin db<2>
*.iopin db<1>
*.iopin db<0>
*.ipin VSS
*.ipin VREF
*.iopin t<6>
*.iopin t<5>
*.iopin t<4>
*.iopin t<3>
*.iopin t<2>
*.iopin t<1>
*.iopin t<0>
*.iopin tb<6>
*.iopin tb<5>
*.iopin tb<4>
*.iopin tb<3>
*.iopin tb<2>
*.iopin tb<1>
*.iopin tb<0>
*.ipin VDD
x1 sw5 sw1 sw0 sw2 sw6 sw4 sw3 t<6> t<5> t<4> t<3> t<2> t<1> t<0> VSS t<0> hgu_cdac_8bit_array
x2 VREF d<4> d<1> d<2> d<3> d<5> d<6> d<0> sw2 sw3 sw4 sw5 sw0 sw1 sw6 VSS VDD hgu_cdac_drv
x3 swd5 swd1 swd0 swd2 swd6 swd4 swd3 tb<6> tb<5> tb<4> tb<3> tb<2> tb<1> tb<0> VSS tb<0>
+ hgu_cdac_8bit_array
x4 VREF db<4> db<1> db<2> db<3> db<5> db<6> db<0> swd2 swd3 swd4 swd5 swd0 swd1 swd6 VSS VDD
+ hgu_cdac_drv
.ends


* expanding   symbol:  ../xschem/hgu_cdac_sw_buffer.sym # of pins=12
** sym_path: /foss/designs/hgu_goss/hgu/xschem/hgu_cdac_sw_buffer.sym
** sch_path: /foss/designs/hgu_goss/hgu/xschem/hgu_cdac_sw_buffer.sch
.subckt hgu_cdac_sw_buffer sar_val<3> sar_val<6> sar_val<4> sar_val<5> sar_val<7> sw<2> sw<5> sw<3>
+ sw<4> sw<6> VDD VSS
*.ipin sar_val<7>
*.opin sw<6>
*.opin sw<5>
*.opin sw<4>
*.opin sw<3>
*.opin sw<2>
*.ipin sar_val<6>
*.ipin sar_val<5>
*.ipin sar_val<4>
*.ipin sar_val<3>
*.ipin VDD
*.ipin VSS
x9 sar_val<7> VSS VSS VDD VDD net1 sky130_fd_sc_hd__buf_1
x10 net1 VSS VSS VDD VDD net2 sky130_fd_sc_hd__buf_4
x11 net2 VSS VSS VDD VDD sw<6> sky130_fd_sc_hd__buf_16
x1 net3 VSS VSS VDD VDD sw<5> sky130_fd_sc_hd__buf_4
x2 net4 VSS VSS VDD VDD sw<4> sky130_fd_sc_hd__buf_4
x3 sar_val<6> VSS VSS VDD VDD net3 sky130_fd_sc_hd__buf_1
x4 sar_val<5> VSS VSS VDD VDD net4 sky130_fd_sc_hd__buf_1
x5 sar_val<4> VSS VSS VDD VDD sw<3> sky130_fd_sc_hd__buf_1
x6 sar_val<3> VSS VSS VDD VDD sw<2> sky130_fd_sc_hd__buf_1
x7 VSS VSS VSS VDD VDD net5 sky130_fd_sc_hd__buf_1
x8 VSS VSS VSS VDD VDD net6 sky130_fd_sc_hd__buf_1
x12 VSS VSS VSS VDD VDD net7 sky130_fd_sc_hd__buf_1
.ends


* expanding   symbol:  ../xschem/hgu_clk_async.sym # of pins=9
** sym_path: /foss/designs/hgu_goss/hgu/xschem/hgu_clk_async.sym
** sch_path: /foss/designs/hgu_goss/hgu/xschem/hgu_clk_async.sch
.subckt hgu_clk_async ASYNC_CLK_SAR VDD VSS sample_clk EOB READY delay_offset
+ async_resetb_delay_ctrl_code[0] async_resetb_delay_ctrl_code[1] async_resetb_delay_ctrl_code[2] async_resetb_delay_ctrl_code[3]
+ async_setb_delay_ctrl_code[0] async_setb_delay_ctrl_code[1] async_setb_delay_ctrl_code[2] async_setb_delay_ctrl_code[3]
*.ipin VDD
*.opin ASYNC_CLK_SAR
*.ipin VSS
*.ipin sample_clk
*.ipin EOB
*.ipin READY
*.ipin
*+ async_resetb_delay_ctrl_code[0],async_resetb_delay_ctrl_code[1],async_resetb_delay_ctrl_code[2],async_resetb_delay_ctrl_code[3]
*.ipin
*+ async_setb_delay_ctrl_code[0],async_setb_delay_ctrl_code[1],async_setb_delay_ctrl_code[2],async_setb_delay_ctrl_code[3]
*.ipin delay_offset
x3 net1 VSS sample_clk VSS VSS vDD VDD net4 sky130_fd_sc_hd__mux2_1
x8 net4 VSS EOB VSS VSS vDD VDD ASYNC_CLK_SAR sky130_fd_sc_hd__mux2_1
x27 sample_clk VDD net5 net6 VSS VSS vDD VDD net1 net7 sky130_fd_sc_hd__dfbbp_1
x9 net2 VSS VSS vDD VDD net6 sky130_fd_sc_hd__inv_1
x10 net3 VSS VSS vDD VDD net5 sky130_fd_sc_hd__inv_1
x2 VDD READY net2 VSS async_setb_delay_ctrl_code[0] async_setb_delay_ctrl_code[1]
+ async_setb_delay_ctrl_code[2] async_setb_delay_ctrl_code[3] delay_offset hgu_delay_no_code
x4 VDD ASYNC_CLK_SAR net3 VSS async_resetb_delay_ctrl_code[0] async_resetb_delay_ctrl_code[1]
+ async_resetb_delay_ctrl_code[2] async_resetb_delay_ctrl_code[3] delay_offset hgu_delay_no_code
C3 net3 VSS 5f m=1
C1 net2 VSS 5f m=1
C2 net4 VSS 5f m=1
C4 net1 VSS 5f m=1
.ends


* expanding   symbol:  ../xschem/hgu_clk_sample.sym # of pins=12
** sym_path: /foss/designs/hgu_goss/hgu/xschem/hgu_clk_sample.sym
** sch_path: /foss/designs/hgu_goss/hgu/xschem/hgu_clk_sample.sch
.subckt hgu_clk_sample SAMPLE_CLK_b VDD VSS CLK RESET SET SAMPLE_CLK CAP_CTRL_CODE0[0]
+ CAP_CTRL_CODE0[1] CAP_CTRL_CODE0[2] CAP_CTRL_CODE0[3] CAP_CTRL_CODE1[0] CAP_CTRL_CODE1[1] CAP_CTRL_CODE1[2]
+ CAP_CTRL_CODE1[3] CAP_CTRL_CODE2[0] CAP_CTRL_CODE2[1] CAP_CTRL_CODE2[2] CAP_CTRL_CODE2[3] CAP_CTRL_CODE3[0]
+ CAP_CTRL_CODE3[1] CAP_CTRL_CODE3[2] CAP_CTRL_CODE3[3] sample_delay_offset
*.ipin VDD
*.ipin VSS
*.ipin SET
*.ipin RESET
*.ipin CLK
*.opin SAMPLE_CLK
*.opin SAMPLE_CLK_b
*.ipin CAP_CTRL_CODE1[0],CAP_CTRL_CODE1[1],CAP_CTRL_CODE1[2],CAP_CTRL_CODE1[3]
*.ipin CAP_CTRL_CODE2[0],CAP_CTRL_CODE2[1],CAP_CTRL_CODE2[2],CAP_CTRL_CODE2[3]
*.ipin CAP_CTRL_CODE3[0],CAP_CTRL_CODE3[1],CAP_CTRL_CODE3[2],CAP_CTRL_CODE3[3]
*.ipin CAP_CTRL_CODE0[0],CAP_CTRL_CODE0[1],CAP_CTRL_CODE0[2],CAP_CTRL_CODE0[3]
*.ipin sample_delay_offset
x1 VDD VSS CLK net2 RESET SET hgu_clk_div
x2 net8 net2 VDD VSS CAP_CTRL_CODE0[0] CAP_CTRL_CODE0[1] CAP_CTRL_CODE0[2] CAP_CTRL_CODE0[3]
+ CAP_CTRL_CODE1[0] CAP_CTRL_CODE1[1] CAP_CTRL_CODE1[2] CAP_CTRL_CODE1[3] CAP_CTRL_CODE2[0] CAP_CTRL_CODE2[1]
+ CAP_CTRL_CODE2[2] CAP_CTRL_CODE2[3] CAP_CTRL_CODE3[0] CAP_CTRL_CODE3[1] CAP_CTRL_CODE3[2] CAP_CTRL_CODE3[3]
+ sample_delay_offset hgu_delay
x7 net8 VSS VSS vDD VDD net1 sky130_fd_sc_hd__inv_1
C1 net1 VSS 5f m=1
C2 net2 VSS 5f m=1
C3 net8 VSS 5f m=1
x3 net2 net1 VSS VSS vDD VDD net4 sky130_fd_sc_hd__nand2_1
XM7 net7 net3 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM8 net7 net3 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1.26 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM9 net5 net4 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM10 net5 net4 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM11 net6 net5 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM12 net6 net5 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1.26 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM13 net4 VSS net3 VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1.9 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM14 net4 VDD net3 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM18 SAMPLE_CLK_b net7 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1.26 nf=3 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM17 SAMPLE_CLK_b net7 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=3.78 nf=3 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM15 SAMPLE_CLK net6 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1.26 nf=3 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM16 SAMPLE_CLK net6 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=3.78 nf=3 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  ../xschem/hgu_sarlogic_8bit_logic.sym # of pins=9
** sym_path: /foss/designs/hgu_goss/hgu/xschem/hgu_sarlogic_8bit_logic.sym
** sch_path: /foss/designs/hgu_goss/hgu/xschem/hgu_sarlogic_8bit_logic.sch
.subckt hgu_sarlogic_8bit_logic sel_bit[0] sel_bit[1] EOB clk_sar D[0] D[1] D[2] D[3] D[4] D[5] D[6]
+ D[7] comparator_out check[0] check[1] check[2] check[3] check[4] check[5] check[6] reset VDD VSS
*.ipin clk_sar
*.ipin VDD
*.ipin VSS
*.ipin comparator_out
*.ipin reset
*.opin EOB
*.opin D[0],D[1],D[2],D[3],D[4],D[5],D[6],D[7]
*.opin check[0],check[1],check[2],check[3],check[4],check[5],check[6]
*.ipin sel_bit[0],sel_bit[1]
x20 clk_sar_buff EOB VDD resetb VSS VSS VDD VDD net1 net4 sky130_fd_sc_hd__dfbbp_1
x27 clk_sar_buff net1 resetb VDD VSS VSS VDD VDD check[6] net5 sky130_fd_sc_hd__dfbbp_1
x30 clk_sar_buff check[6] resetb VDD VSS VSS VDD VDD check[5] net6 sky130_fd_sc_hd__dfbbp_1
x33 clk_sar_buff check[5] resetb VDD VSS VSS VDD VDD check[4] net7 sky130_fd_sc_hd__dfbbp_1
x36 clk_sar_buff check[4] resetb VDD VSS VSS VDD VDD check[3] net8 sky130_fd_sc_hd__dfbbp_1
x39 clk_sar_buff check[3] resetb VDD VSS VSS VDD VDD check[2] net9 sky130_fd_sc_hd__dfbbp_1
x42 clk_sar_buff check[2] resetb VDD VSS VSS VDD VDD check[1] net10 sky130_fd_sc_hd__dfbbp_1
x45 clk_sar_buff check[1] resetb VDD VSS VSS VDD VDD check[0] net11 sky130_fd_sc_hd__dfbbp_1
x48 clk_sar_buff check[0] resetb VDD VSS VSS VDD VDD net3 net12 sky130_fd_sc_hd__dfbbp_1
x51 D[6] comparator_out_buff resetb net4 VSS VSS VDD VDD D[7] net13 sky130_fd_sc_hd__dfbbp_1
x54 D[5] comparator_out_buff resetb net5 VSS VSS VDD VDD D[6] net14 sky130_fd_sc_hd__dfbbp_1
x57 D[4] comparator_out_buff resetb net6 VSS VSS VDD VDD D[5] net15 sky130_fd_sc_hd__dfbbp_1
x60 D[3] comparator_out_buff resetb net7 VSS VSS VDD VDD D[4] net16 sky130_fd_sc_hd__dfbbp_1
x63 D[2] comparator_out_buff resetb net8 VSS VSS VDD VDD D[3] net17 sky130_fd_sc_hd__dfbbp_1
x66 D[1] comparator_out_buff resetb net9 VSS VSS VDD VDD D[2] net18 sky130_fd_sc_hd__dfbbp_1
x69 D[0] comparator_out_buff resetb net10 VSS VSS VDD VDD D[1] net19 sky130_fd_sc_hd__dfbbp_1
x72 net2 comparator_out_buff resetb net11 VSS VSS VDD VDD D[0] net20 sky130_fd_sc_hd__dfbbp_1
x75 VSS VSS resetb net21 VSS VSS VDD VDD net2 net22 sky130_fd_sc_hd__dfbbp_1
x77 EOB VSS VSS VDD VDD net21 sky130_fd_sc_hd__inv_1
x78 check[2] check[1] check[0] net3 sel_bit[0] sel_bit[1] VSS VSS VDD VDD EOB
+ sky130_fd_sc_hd__mux4_4
C2[17] resetb VSS 5f m=1
C2[16] resetb VSS 5f m=1
C2[15] resetb VSS 5f m=1
C2[14] resetb VSS 5f m=1
C2[13] resetb VSS 5f m=1
C2[12] resetb VSS 5f m=1
C2[11] resetb VSS 5f m=1
C2[10] resetb VSS 5f m=1
C2[9] resetb VSS 5f m=1
C2[8] resetb VSS 5f m=1
C2[7] resetb VSS 5f m=1
C2[6] resetb VSS 5f m=1
C2[5] resetb VSS 5f m=1
C2[4] resetb VSS 5f m=1
C2[3] resetb VSS 5f m=1
C2[2] resetb VSS 5f m=1
C2[1] resetb VSS 5f m=1
C2[0] resetb VSS 5f m=1
C2 net1 VSS 5f m=1
C3 check[6] VSS 5f m=1
C4 check[5] VSS 5f m=1
C5 check[4] VSS 5f m=1
C6 check[3] VSS 5f m=1
C7 check[2] VSS 5f m=1
C8 check[1] VSS 5f m=1
C9 check[0] VSS 5f m=1
C10 net3 VSS 5f m=1
C11 EOB VSS 5f m=1
C12 D[6] VSS 5f m=1
C13 D[5] VSS 5f m=1
C14 D[4] VSS 5f m=1
C15 D[3] VSS 5f m=1
C16 D[2] VSS 5f m=1
C17 D[1] VSS 5f m=1
C18 D[0] VSS 5f m=1
C19 net2 VSS 5f m=1
C20 D[7] VSS 5f m=1
C21 D[6] VSS 5f m=1
C22 D[5] VSS 5f m=1
C23 D[4] VSS 5f m=1
C24 D[3] VSS 5f m=1
C25 D[2] VSS 5f m=1
C26 D[1] VSS 5f m=1
C27 D[0] VSS 5f m=1
C28 net5 VSS 5f m=1
C29 net6 VSS 5f m=1
C30 net7 VSS 5f m=1
C31 net8 VSS 5f m=1
C32 net9 VSS 5f m=1
C33 net10 VSS 5f m=1
C34 net11 VSS 5f m=1
C35 net21 VSS 5f m=1
C36 clk_sar_buff VSS 5f m=1
x1 reset VSS VSS VDD VDD net23 sky130_fd_sc_hd__buf_1
x2 clk_sar VSS VSS VDD VDD net24 sky130_fd_sc_hd__buf_1
x3 net23 VSS VSS VDD VDD net25 sky130_fd_sc_hd__buf_4
x4 net25 VSS VSS VDD VDD resetb sky130_fd_sc_hd__buf_16
x5 net24 VSS VSS VDD VDD clk_sar_buff sky130_fd_sc_hd__buf_4
x6 comparator_out VSS VSS VDD VDD net26 sky130_fd_sc_hd__buf_1
x7 net26 VSS VSS VDD VDD comparator_out_buff sky130_fd_sc_hd__buf_4
C1[17] comparator_out_buff VSS 5f m=1
C1[16] comparator_out_buff VSS 5f m=1
C1[15] comparator_out_buff VSS 5f m=1
C1[14] comparator_out_buff VSS 5f m=1
C1[13] comparator_out_buff VSS 5f m=1
C1[12] comparator_out_buff VSS 5f m=1
C1[11] comparator_out_buff VSS 5f m=1
C1[10] comparator_out_buff VSS 5f m=1
C1[9] comparator_out_buff VSS 5f m=1
C1[8] comparator_out_buff VSS 5f m=1
C1[7] comparator_out_buff VSS 5f m=1
C1[6] comparator_out_buff VSS 5f m=1
C1[5] comparator_out_buff VSS 5f m=1
C1[4] comparator_out_buff VSS 5f m=1
C1[3] comparator_out_buff VSS 5f m=1
C1[2] comparator_out_buff VSS 5f m=1
C1[1] comparator_out_buff VSS 5f m=1
C1[0] comparator_out_buff VSS 5f m=1
.ends


* expanding   symbol:  ../xschem/hgu_sarlogic_sw_ctrl.sym # of pins=10
** sym_path: /foss/designs/hgu_goss/hgu/xschem/hgu_sarlogic_sw_ctrl.sym
** sch_path: /foss/designs/hgu_goss/hgu/xschem/hgu_sarlogic_sw_ctrl.sch
.subckt hgu_sarlogic_sw_ctrl VDD VSS vdd_sw[1] vdd_sw[2] vdd_sw[3] vdd_sw[4] vdd_sw[5] vdd_sw[6]
+ vdd_sw[7] vdd_sw_b[1] vdd_sw_b[2] vdd_sw_b[3] vdd_sw_b[4] vdd_sw_b[5] vdd_sw_b[6] vdd_sw_b[7] D[1] D[2] D[3]
+ D[4] D[5] D[6] D[7] vss_sw[1] vss_sw[2] vss_sw[3] vss_sw[4] vss_sw[5] vss_sw[6] vss_sw[7] check[0]
+ check[1] check[2] check[3] check[4] check[5] check[6] vss_sw_b[1] vss_sw_b[2] vss_sw_b[3] vss_sw_b[4]
+ vss_sw_b[5] vss_sw_b[6] vss_sw_b[7] READY reset
*.opin vdd_sw[1],vdd_sw[2],vdd_sw[3],vdd_sw[4],vdd_sw[5],vdd_sw[6],vdd_sw[7]
*.opin vdd_sw_b[1],vdd_sw_b[2],vdd_sw_b[3],vdd_sw_b[4],vdd_sw_b[5],vdd_sw_b[6],vdd_sw_b[7]
*.opin vss_sw[1],vss_sw[2],vss_sw[3],vss_sw[4],vss_sw[5],vss_sw[6],vss_sw[7]
*.opin vss_sw_b[1],vss_sw_b[2],vss_sw_b[3],vss_sw_b[4],vss_sw_b[5],vss_sw_b[6],vss_sw_b[7]
*.ipin VDD
*.ipin VSS
*.ipin READY
*.ipin D[1],D[2],D[3],D[4],D[5],D[6],D[7]
*.ipin check[0],check[1],check[2],check[3],check[4],check[5],check[6]
*.ipin reset
x4 net1 D[7] VDD resetb VSS VSS VDD VDD vdd_sw[7] vdd_sw_b[7] sky130_fd_sc_hd__dfbbn_1
x5 net2 D[7] resetb VDD VSS VSS VDD VDD vss_sw[7] vss_sw_b[7] sky130_fd_sc_hd__dfbbn_1
x19 net3 D[6] VDD resetb VSS VSS VDD VDD vdd_sw[6] vdd_sw_b[6] sky130_fd_sc_hd__dfbbn_1
x21 net4 D[6] resetb VDD VSS VSS VDD VDD vss_sw[6] vss_sw_b[6] sky130_fd_sc_hd__dfbbn_1
x23 net5 D[5] VDD resetb VSS VSS VDD VDD vdd_sw[5] vdd_sw_b[5] sky130_fd_sc_hd__dfbbn_1
x24 net6 D[5] resetb VDD VSS VSS VDD VDD vss_sw[5] vss_sw_b[5] sky130_fd_sc_hd__dfbbn_1
x25 net7 D[4] VDD resetb VSS VSS VDD VDD vdd_sw[4] vdd_sw_b[4] sky130_fd_sc_hd__dfbbn_1
x26 net8 D[4] resetb VDD VSS VSS VDD VDD vss_sw[4] vss_sw_b[4] sky130_fd_sc_hd__dfbbn_1
x28 net9 D[3] VDD resetb VSS VSS VDD VDD vdd_sw[3] vdd_sw_b[3] sky130_fd_sc_hd__dfbbn_1
x29 net10 D[3] resetb VDD VSS VSS VDD VDD vss_sw[3] vss_sw_b[3] sky130_fd_sc_hd__dfbbn_1
x31 net11 D[2] VDD resetb VSS VSS VDD VDD vdd_sw[2] vdd_sw_b[2] sky130_fd_sc_hd__dfbbn_1
x32 net12 D[2] resetb VDD VSS VSS VDD VDD vss_sw[2] vss_sw_b[2] sky130_fd_sc_hd__dfbbn_1
x34 net13 D[1] VDD resetb VSS VSS VDD VDD vdd_sw[1] vdd_sw_b[1] sky130_fd_sc_hd__dfbbn_1
x35 net14 D[1] resetb VDD VSS VSS VDD VDD vss_sw[1] vss_sw_b[1] sky130_fd_sc_hd__dfbbn_1
x6 VSS READY_buff check[6] VSS VSS VDD VDD net1 sky130_fd_sc_hd__mux2_1
x7 VSS READY_buff check[6] VSS VSS VDD VDD net2 sky130_fd_sc_hd__mux2_1
x8 VSS READY_buff check[5] VSS VSS VDD VDD net3 sky130_fd_sc_hd__mux2_1
x9 VSS READY_buff check[5] VSS VSS VDD VDD net4 sky130_fd_sc_hd__mux2_1
x10 VSS READY_buff check[4] VSS VSS VDD VDD net5 sky130_fd_sc_hd__mux2_1
x11 VSS READY_buff check[4] VSS VSS VDD VDD net6 sky130_fd_sc_hd__mux2_1
x12 VSS READY_buff check[3] VSS VSS VDD VDD net7 sky130_fd_sc_hd__mux2_1
x13 VSS READY_buff check[3] VSS VSS VDD VDD net8 sky130_fd_sc_hd__mux2_1
x14 VSS READY_buff check[2] VSS VSS VDD VDD net9 sky130_fd_sc_hd__mux2_1
x15 VSS READY_buff check[2] VSS VSS VDD VDD net10 sky130_fd_sc_hd__mux2_1
x16 VSS READY_buff check[1] VSS VSS VDD VDD net11 sky130_fd_sc_hd__mux2_1
x17 VSS READY_buff check[1] VSS VSS VDD VDD net12 sky130_fd_sc_hd__mux2_1
x18 VSS READY_buff check[0] VSS VSS VDD VDD net13 sky130_fd_sc_hd__mux2_1
x20 VSS READY_buff check[0] VSS VSS VDD VDD net14 sky130_fd_sc_hd__mux2_1
x1 reset VSS VSS VDD VDD net15 sky130_fd_sc_hd__buf_1
x3 net15 VSS VSS VDD VDD net16 sky130_fd_sc_hd__buf_4
x2 net16 VSS VSS VDD VDD resetb sky130_fd_sc_hd__buf_16
x22 READY VSS VSS VDD VDD net17 sky130_fd_sc_hd__buf_1
x27 net17 VSS VSS VDD VDD net18 sky130_fd_sc_hd__buf_4
x30 net18 VSS VSS VDD VDD READY_buff sky130_fd_sc_hd__buf_16
.ends


* expanding   symbol:  /foss/designs/hgu_goss/hgu/xschem/hgu_sarlogic_retimer.sym # of pins=7
** sym_path: /foss/designs/hgu_goss/hgu/xschem/hgu_sarlogic_retimer.sym
** sch_path: /foss/designs/hgu_goss/hgu/xschem/hgu_sarlogic_retimer.sch
.subckt hgu_sarlogic_retimer VDD VSS sar_logic[0] sar_logic[1] sar_logic[2] sar_logic[3]
+ sar_logic[4] sar_logic[5] sar_logic[6] sar_logic[7] eob delay_code[0] delay_code[1] delay_code[2] delay_code[3]
+ delay_offset sar_retimer[0] sar_retimer[1] sar_retimer[2] sar_retimer[3] sar_retimer[4] sar_retimer[5]
+ sar_retimer[6] sar_retimer[7]
*.ipin
*+ sar_logic[0],sar_logic[1],sar_logic[2],sar_logic[3],sar_logic[4],sar_logic[5],sar_logic[6],sar_logic[7]
*.opin
*+ sar_retimer[0],sar_retimer[1],sar_retimer[2],sar_retimer[3],sar_retimer[4],sar_retimer[5],sar_retimer[6],sar_retimer[7]
*.ipin eob
*.ipin VDD
*.ipin VSS
*.ipin delay_code[0],delay_code[1],delay_code[2],delay_code[3]
*.ipin delay_offset
x1[0] eob_delay sar_logic[0] VDD VDD VSS VSS VDD VDD sar_retimer[0] net2[7] sky130_fd_sc_hd__dfbbp_1
x1[1] eob_delay sar_logic[1] VDD VDD VSS VSS VDD VDD sar_retimer[1] net2[6] sky130_fd_sc_hd__dfbbp_1
x1[2] eob_delay sar_logic[2] VDD VDD VSS VSS VDD VDD sar_retimer[2] net2[5] sky130_fd_sc_hd__dfbbp_1
x1[3] eob_delay sar_logic[3] VDD VDD VSS VSS VDD VDD sar_retimer[3] net2[4] sky130_fd_sc_hd__dfbbp_1
x1[4] eob_delay sar_logic[4] VDD VDD VSS VSS VDD VDD sar_retimer[4] net2[3] sky130_fd_sc_hd__dfbbp_1
x1[5] eob_delay sar_logic[5] VDD VDD VSS VSS VDD VDD sar_retimer[5] net2[2] sky130_fd_sc_hd__dfbbp_1
x1[6] eob_delay sar_logic[6] VDD VDD VSS VSS VDD VDD sar_retimer[6] net2[1] sky130_fd_sc_hd__dfbbp_1
x1[7] eob_delay sar_logic[7] VDD VDD VSS VSS VDD VDD sar_retimer[7] net2[0] sky130_fd_sc_hd__dfbbp_1
x2 VDD eob net1 VSS delay_code[0] delay_code[1] delay_code[2] delay_code[3] delay_offset
+ hgu_delay_no_code
x3 net1 VSS VSS VDD VDD eob_delay sky130_fd_sc_hd__buf_2
.ends


* expanding   symbol:  ../xschem/hgu_cdac_8bit_array.sym # of pins=16
** sym_path: /foss/designs/hgu_goss/hgu/xschem/hgu_cdac_8bit_array.sym
** sch_path: /foss/designs/hgu_goss/hgu/xschem/hgu_cdac_8bit_array.sch
.subckt hgu_cdac_8bit_array drv<31:0> drv<1:0> drv<0> drv<3:0> drv<63:0> drv<15:0> drv<7:0>
+ tah<63:0> tah<31:0> tah<15:0> tah<7:0> tah<3:0> tah<1:0> tah<0> SUB tu
*.iopin drv<0>
*.iopin drv<1:0>
*.iopin drv<3:0>
*.iopin drv<7:0>
*.iopin drv<15:0>
*.iopin drv<31:0>
*.iopin drv<63:0>
*.iopin tah<0>
*.iopin tah<1:0>
*.iopin tah<3:0>
*.iopin tah<7:0>
*.iopin tah<15:0>
*.iopin tah<31:0>
*.iopin tah<63:0>
*.iopin SUB
*.iopin tu

.ends


* expanding   symbol:  ../xschem/hgu_cdac_drv.sym # of pins=17
** sym_path: /foss/designs/hgu_goss/hgu/xschem/hgu_cdac_drv.sym
** sch_path: /foss/designs/hgu_goss/hgu/xschem/hgu_cdac_drv.sch
.subckt hgu_cdac_drv VREF SAR<4> SAR<1> SAR<2> SAR<3> SAR<5> SAR<6> SAR<0> C<3:0> C<7:0> C<15:0>
+ C<31:0> C<0> C<1:0> C<63:0> VSS VDD
*.ipin VREF
*.ipin VSS
*.ipin SAR<6>
*.ipin SAR<5>
*.ipin SAR<4>
*.ipin SAR<3>
*.ipin SAR<2>
*.ipin SAR<1>
*.ipin SAR<0>
*.opin C<63:0>
*.opin C<31:0>
*.opin C<15:0>
*.opin C<7:0>
*.opin C<3:0>
*.opin C<1:0>
*.opin C<0>
*.ipin VDD
x7[63] VDD SAR<6> C<63:0> VSS VREF hgu_inverter
x7[62] VDD SAR<6> C<63:0> VSS VREF hgu_inverter
x7[61] VDD SAR<6> C<63:0> VSS VREF hgu_inverter
x7[60] VDD SAR<6> C<63:0> VSS VREF hgu_inverter
x7[59] VDD SAR<6> C<63:0> VSS VREF hgu_inverter
x7[58] VDD SAR<6> C<63:0> VSS VREF hgu_inverter
x7[57] VDD SAR<6> C<63:0> VSS VREF hgu_inverter
x7[56] VDD SAR<6> C<63:0> VSS VREF hgu_inverter
x7[55] VDD SAR<6> C<63:0> VSS VREF hgu_inverter
x7[54] VDD SAR<6> C<63:0> VSS VREF hgu_inverter
x7[53] VDD SAR<6> C<63:0> VSS VREF hgu_inverter
x7[52] VDD SAR<6> C<63:0> VSS VREF hgu_inverter
x7[51] VDD SAR<6> C<63:0> VSS VREF hgu_inverter
x7[50] VDD SAR<6> C<63:0> VSS VREF hgu_inverter
x7[49] VDD SAR<6> C<63:0> VSS VREF hgu_inverter
x7[48] VDD SAR<6> C<63:0> VSS VREF hgu_inverter
x7[47] VDD SAR<6> C<63:0> VSS VREF hgu_inverter
x7[46] VDD SAR<6> C<63:0> VSS VREF hgu_inverter
x7[45] VDD SAR<6> C<63:0> VSS VREF hgu_inverter
x7[44] VDD SAR<6> C<63:0> VSS VREF hgu_inverter
x7[43] VDD SAR<6> C<63:0> VSS VREF hgu_inverter
x7[42] VDD SAR<6> C<63:0> VSS VREF hgu_inverter
x7[41] VDD SAR<6> C<63:0> VSS VREF hgu_inverter
x7[40] VDD SAR<6> C<63:0> VSS VREF hgu_inverter
x7[39] VDD SAR<6> C<63:0> VSS VREF hgu_inverter
x7[38] VDD SAR<6> C<63:0> VSS VREF hgu_inverter
x7[37] VDD SAR<6> C<63:0> VSS VREF hgu_inverter
x7[36] VDD SAR<6> C<63:0> VSS VREF hgu_inverter
x7[35] VDD SAR<6> C<63:0> VSS VREF hgu_inverter
x7[34] VDD SAR<6> C<63:0> VSS VREF hgu_inverter
x7[33] VDD SAR<6> C<63:0> VSS VREF hgu_inverter
x7[32] VDD SAR<6> C<63:0> VSS VREF hgu_inverter
x7[31] VDD SAR<6> C<63:0> VSS VREF hgu_inverter
x7[30] VDD SAR<6> C<63:0> VSS VREF hgu_inverter
x7[29] VDD SAR<6> C<63:0> VSS VREF hgu_inverter
x7[28] VDD SAR<6> C<63:0> VSS VREF hgu_inverter
x7[27] VDD SAR<6> C<63:0> VSS VREF hgu_inverter
x7[26] VDD SAR<6> C<63:0> VSS VREF hgu_inverter
x7[25] VDD SAR<6> C<63:0> VSS VREF hgu_inverter
x7[24] VDD SAR<6> C<63:0> VSS VREF hgu_inverter
x7[23] VDD SAR<6> C<63:0> VSS VREF hgu_inverter
x7[22] VDD SAR<6> C<63:0> VSS VREF hgu_inverter
x7[21] VDD SAR<6> C<63:0> VSS VREF hgu_inverter
x7[20] VDD SAR<6> C<63:0> VSS VREF hgu_inverter
x7[19] VDD SAR<6> C<63:0> VSS VREF hgu_inverter
x7[18] VDD SAR<6> C<63:0> VSS VREF hgu_inverter
x7[17] VDD SAR<6> C<63:0> VSS VREF hgu_inverter
x7[16] VDD SAR<6> C<63:0> VSS VREF hgu_inverter
x7[15] VDD SAR<6> C<63:0> VSS VREF hgu_inverter
x7[14] VDD SAR<6> C<63:0> VSS VREF hgu_inverter
x7[13] VDD SAR<6> C<63:0> VSS VREF hgu_inverter
x7[12] VDD SAR<6> C<63:0> VSS VREF hgu_inverter
x7[11] VDD SAR<6> C<63:0> VSS VREF hgu_inverter
x7[10] VDD SAR<6> C<63:0> VSS VREF hgu_inverter
x7[9] VDD SAR<6> C<63:0> VSS VREF hgu_inverter
x7[8] VDD SAR<6> C<63:0> VSS VREF hgu_inverter
x7[7] VDD SAR<6> C<63:0> VSS VREF hgu_inverter
x7[6] VDD SAR<6> C<63:0> VSS VREF hgu_inverter
x7[5] VDD SAR<6> C<63:0> VSS VREF hgu_inverter
x7[4] VDD SAR<6> C<63:0> VSS VREF hgu_inverter
x7[3] VDD SAR<6> C<63:0> VSS VREF hgu_inverter
x7[2] VDD SAR<6> C<63:0> VSS VREF hgu_inverter
x7[1] VDD SAR<6> C<63:0> VSS VREF hgu_inverter
x7[0] VDD SAR<6> C<63:0> VSS VREF hgu_inverter
x1 VDD SAR<0> C<0> VSS VREF hgu_inverter
x2[1] VDD SAR<1> C<1:0> VSS VREF hgu_inverter
x2[0] VDD SAR<1> C<1:0> VSS VREF hgu_inverter
x3[3] VDD SAR<2> C<3:0> VSS VREF hgu_inverter
x3[2] VDD SAR<2> C<3:0> VSS VREF hgu_inverter
x3[1] VDD SAR<2> C<3:0> VSS VREF hgu_inverter
x3[0] VDD SAR<2> C<3:0> VSS VREF hgu_inverter
x4[7] VDD SAR<3> C<7:0> VSS VREF hgu_inverter
x4[6] VDD SAR<3> C<7:0> VSS VREF hgu_inverter
x4[5] VDD SAR<3> C<7:0> VSS VREF hgu_inverter
x4[4] VDD SAR<3> C<7:0> VSS VREF hgu_inverter
x4[3] VDD SAR<3> C<7:0> VSS VREF hgu_inverter
x4[2] VDD SAR<3> C<7:0> VSS VREF hgu_inverter
x4[1] VDD SAR<3> C<7:0> VSS VREF hgu_inverter
x4[0] VDD SAR<3> C<7:0> VSS VREF hgu_inverter
x5[15] VDD SAR<4> C<15:0> VSS VREF hgu_inverter
x5[14] VDD SAR<4> C<15:0> VSS VREF hgu_inverter
x5[13] VDD SAR<4> C<15:0> VSS VREF hgu_inverter
x5[12] VDD SAR<4> C<15:0> VSS VREF hgu_inverter
x5[11] VDD SAR<4> C<15:0> VSS VREF hgu_inverter
x5[10] VDD SAR<4> C<15:0> VSS VREF hgu_inverter
x5[9] VDD SAR<4> C<15:0> VSS VREF hgu_inverter
x5[8] VDD SAR<4> C<15:0> VSS VREF hgu_inverter
x5[7] VDD SAR<4> C<15:0> VSS VREF hgu_inverter
x5[6] VDD SAR<4> C<15:0> VSS VREF hgu_inverter
x5[5] VDD SAR<4> C<15:0> VSS VREF hgu_inverter
x5[4] VDD SAR<4> C<15:0> VSS VREF hgu_inverter
x5[3] VDD SAR<4> C<15:0> VSS VREF hgu_inverter
x5[2] VDD SAR<4> C<15:0> VSS VREF hgu_inverter
x5[1] VDD SAR<4> C<15:0> VSS VREF hgu_inverter
x5[0] VDD SAR<4> C<15:0> VSS VREF hgu_inverter
x6[31] VDD SAR<5> C<31:0> VSS VREF hgu_inverter
x6[30] VDD SAR<5> C<31:0> VSS VREF hgu_inverter
x6[29] VDD SAR<5> C<31:0> VSS VREF hgu_inverter
x6[28] VDD SAR<5> C<31:0> VSS VREF hgu_inverter
x6[27] VDD SAR<5> C<31:0> VSS VREF hgu_inverter
x6[26] VDD SAR<5> C<31:0> VSS VREF hgu_inverter
x6[25] VDD SAR<5> C<31:0> VSS VREF hgu_inverter
x6[24] VDD SAR<5> C<31:0> VSS VREF hgu_inverter
x6[23] VDD SAR<5> C<31:0> VSS VREF hgu_inverter
x6[22] VDD SAR<5> C<31:0> VSS VREF hgu_inverter
x6[21] VDD SAR<5> C<31:0> VSS VREF hgu_inverter
x6[20] VDD SAR<5> C<31:0> VSS VREF hgu_inverter
x6[19] VDD SAR<5> C<31:0> VSS VREF hgu_inverter
x6[18] VDD SAR<5> C<31:0> VSS VREF hgu_inverter
x6[17] VDD SAR<5> C<31:0> VSS VREF hgu_inverter
x6[16] VDD SAR<5> C<31:0> VSS VREF hgu_inverter
x6[15] VDD SAR<5> C<31:0> VSS VREF hgu_inverter
x6[14] VDD SAR<5> C<31:0> VSS VREF hgu_inverter
x6[13] VDD SAR<5> C<31:0> VSS VREF hgu_inverter
x6[12] VDD SAR<5> C<31:0> VSS VREF hgu_inverter
x6[11] VDD SAR<5> C<31:0> VSS VREF hgu_inverter
x6[10] VDD SAR<5> C<31:0> VSS VREF hgu_inverter
x6[9] VDD SAR<5> C<31:0> VSS VREF hgu_inverter
x6[8] VDD SAR<5> C<31:0> VSS VREF hgu_inverter
x6[7] VDD SAR<5> C<31:0> VSS VREF hgu_inverter
x6[6] VDD SAR<5> C<31:0> VSS VREF hgu_inverter
x6[5] VDD SAR<5> C<31:0> VSS VREF hgu_inverter
x6[4] VDD SAR<5> C<31:0> VSS VREF hgu_inverter
x6[3] VDD SAR<5> C<31:0> VSS VREF hgu_inverter
x6[2] VDD SAR<5> C<31:0> VSS VREF hgu_inverter
x6[1] VDD SAR<5> C<31:0> VSS VREF hgu_inverter
x6[0] VDD SAR<5> C<31:0> VSS VREF hgu_inverter
.ends


* expanding   symbol:  ../xschem/hgu_delay_no_code.sym # of pins=6
** sym_path: /foss/designs/hgu_goss/hgu/xschem/hgu_delay_no_code.sym
** sch_path: /foss/designs/hgu_goss/hgu/xschem/hgu_delay_no_code.sch
.subckt hgu_delay_no_code VDD IN OUT VSS code[0] code[1] code[2] code[3] code_offset
*.ipin IN
*.ipin VDD
*.ipin VSS
*.opin OUT
*.ipin code[0],code[1],code[2],code[3]
*.ipin code_offset
XM13 OUT Uc net2 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM15 net2 Uc VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM46 OUT Uc net1 VDD sky130_fd_pr__pfet_01v8_hvt L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM47 net1 Uc VDD VDD sky130_fd_pr__pfet_01v8_hvt L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
x2 code[0] VSS Uc net5 hgu_sw_cap
x3[1] code[1] VSS Uc net6[1] hgu_sw_cap
x3[0] code[1] VSS Uc net6[0] hgu_sw_cap
x4[3] code[2] VSS Uc net7[3] hgu_sw_cap
x4[2] code[2] VSS Uc net7[2] hgu_sw_cap
x4[1] code[2] VSS Uc net7[1] hgu_sw_cap
x4[0] code[2] VSS Uc net7[0] hgu_sw_cap
x5[7] net3 Uc VDD net9[7] hgu_sw_cap_pmos
x5[6] net3 Uc VDD net9[6] hgu_sw_cap_pmos
x5[5] net3 Uc VDD net9[5] hgu_sw_cap_pmos
x5[4] net3 Uc VDD net9[4] hgu_sw_cap_pmos
x5[3] net3 Uc VDD net9[3] hgu_sw_cap_pmos
x5[2] net3 Uc VDD net9[2] hgu_sw_cap_pmos
x5[1] net3 Uc VDD net9[1] hgu_sw_cap_pmos
x5[0] net3 Uc VDD net9[0] hgu_sw_cap_pmos
x10 code[3] VSS VSS VDD VDD net3 sky130_fd_sc_hd__inv_1
x7 code_offset VSS Uc net8 hgu_sw_cap
x6 net4 Uc VDD net10 hgu_sw_cap_pmos
x11 code_offset VSS VSS VDD VDD net4 sky130_fd_sc_hd__inv_1
x8 VDD IN Uc hgu_pfet_hvt_stack_in_delay
x9 IN Uc VSS hgu_nfet_hvt_stack_in_delay
XM48 VSS OUT net1 VDD sky130_fd_pr__pfet_01v8_hvt L=0.15 W=0.84 nf=2 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM1 VDD OUT net2 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.84 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  ../xschem/hgu_clk_div.sym # of pins=6
** sym_path: /foss/designs/hgu_goss/hgu/xschem/hgu_clk_div.sym
** sch_path: /foss/designs/hgu_goss/hgu/xschem/hgu_clk_div.sch
.subckt hgu_clk_div VDD VSS CLK DIV_CLK RESET SET
*.opin DIV_CLK
*.ipin SET
*.ipin RESET
*.ipin CLK
*.ipin VDD
*.ipin VSS
x2 CLK D_loop net1 net2 VSS VSS vDD VDD DIV_CLK D_loop sky130_fd_sc_hd__dfbbp_1
x3 SET VSS VSS vDD VDD net2 sky130_fd_sc_hd__inv_1
x4 RESET VSS VSS vDD VDD net1 sky130_fd_sc_hd__inv_1
.ends


* expanding   symbol:  ../xschem/hgu_delay.sym # of pins=9
** sym_path: /foss/designs/hgu_goss/hgu/xschem/hgu_delay.sym
** sch_path: /foss/designs/hgu_goss/hgu/xschem/hgu_delay.sch
.subckt hgu_delay OUT IN VDD VSS SAMPLE_CODE0[0] SAMPLE_CODE0[1] SAMPLE_CODE0[2] SAMPLE_CODE0[3]
+ SAMPLE_CODE1[0] SAMPLE_CODE1[1] SAMPLE_CODE1[2] SAMPLE_CODE1[3] SAMPLE_CODE2[0] SAMPLE_CODE2[1] SAMPLE_CODE2[2]
+ SAMPLE_CODE2[3] SAMPLE_CODE3[0] SAMPLE_CODE3[1] SAMPLE_CODE3[2] SAMPLE_CODE3[3] sample_delay_offset
*.ipin IN
*.ipin VDD
*.ipin VSS
*.opin OUT
*.ipin SAMPLE_CODE1[0],SAMPLE_CODE1[1],SAMPLE_CODE1[2],SAMPLE_CODE1[3]
*.ipin SAMPLE_CODE2[0],SAMPLE_CODE2[1],SAMPLE_CODE2[2],SAMPLE_CODE2[3]
*.ipin SAMPLE_CODE3[0],SAMPLE_CODE3[1],SAMPLE_CODE3[2],SAMPLE_CODE3[3]
*.ipin SAMPLE_CODE0[0],SAMPLE_CODE0[1],SAMPLE_CODE0[2],SAMPLE_CODE0[3]
*.ipin sample_delay_offset
x4 VDD IN net1 VSS SAMPLE_CODE0[0] SAMPLE_CODE0[1] SAMPLE_CODE0[2] SAMPLE_CODE0[3]
+ sample_delay_offset hgu_delay_no_code
x1 VDD net1 net2 VSS SAMPLE_CODE1[0] SAMPLE_CODE1[1] SAMPLE_CODE1[2] SAMPLE_CODE1[3]
+ sample_delay_offset hgu_delay_no_code
x2 VDD net2 net3 VSS SAMPLE_CODE2[0] SAMPLE_CODE2[1] SAMPLE_CODE2[2] SAMPLE_CODE2[3]
+ sample_delay_offset hgu_delay_no_code
x3 VDD net3 OUT VSS SAMPLE_CODE3[0] SAMPLE_CODE3[1] SAMPLE_CODE3[2] SAMPLE_CODE3[3]
+ sample_delay_offset hgu_delay_no_code
.ends


* expanding   symbol:  ../xschem/hgu_cdac_unit.sym # of pins=3
** sym_path: /foss/designs/hgu_goss/hgu/xschem/hgu_cdac_unit.sym
** sch_path: /foss/designs/hgu_goss/hgu/xschem/hgu_cdac_unit.sch
*.subckt hgu_cdac_unit CTOP CBOT SUB  csize=1
*.iopin CTOP
*.iopin CBOT
*.iopin SUB
* x1 CTOP CBOT SUB hgu_cdac_unit
*.ends


* expanding   symbol:  ../xschem/hgu_inverter.sym # of pins=5
** sym_path: /foss/designs/hgu_goss/hgu/xschem/hgu_inverter.sym
** sch_path: /foss/designs/hgu_goss/hgu/xschem/hgu_inverter.sch
.subckt hgu_inverter VDD IN OUT VSS VREF
*.ipin IN
*.ipin VREF
*.ipin VSS
*.opin OUT
*.ipin VDD
XM2 OUT IN VREF VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.84 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 OUT IN VSS VSS sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  /foss/designs/hgu_goss/hgu/xschem/hgu_sw_cap.sym # of pins=4
** sym_path: /foss/designs/hgu_goss/hgu/xschem/hgu_sw_cap.sym
** sch_path: /foss/designs/hgu_goss/hgu/xschem/hgu_sw_cap.sch
.subckt hgu_sw_cap SW VSS DELAY_SIGNAL floating
*.ipin SW
*.ipin VSS
*.iopin DELAY_SIGNAL
*.iopin floating
XM14 DELAY_SIGNAL SW floating VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
*x2 floating VSS VSS hgu_cdac_unit
.ends


* expanding   symbol:  /foss/designs/hgu_goss/hgu/xschem/hgu_sw_cap_pmos.sym # of pins=4
** sym_path: /foss/designs/hgu_goss/hgu/xschem/hgu_sw_cap_pmos.sym
** sch_path: /foss/designs/hgu_goss/hgu/xschem/hgu_sw_cap_pmos.sch
.subckt hgu_sw_cap_pmos SW DELAY_SIGNAL VDD floating
*.ipin SW
*.ipin VDD
*.iopin DELAY_SIGNAL
*.iopin floating
XM16 floating SW DELAY_SIGNAL VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
*x1 VDD floating VDD hgu_cdac_unit
.ends


* expanding   symbol:
*+  /foss/designs/hgu_goss/hgu/xschem/../../../hgu_goss/hgu/xschem/hgu_pfet_hvt_stack_in_delay.sym # of pins=3
** sym_path:
*+ /foss/designs/hgu_goss/hgu/xschem/../../../hgu_goss/hgu/xschem/hgu_pfet_hvt_stack_in_delay.sym
** sch_path:
*+ /foss/designs/hgu_goss/hgu/xschem/../../../hgu_goss/hgu/xschem/hgu_pfet_hvt_stack_in_delay.sch
.subckt hgu_pfet_hvt_stack_in_delay VDD input_stack output_stack
*.ipin VDD
*.ipin input_stack
*.iopin output_stack
XM1 output_stack input_stack net1 VDD sky130_fd_pr__pfet_01v8_hvt L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 net1 input_stack net2 VDD sky130_fd_pr__pfet_01v8_hvt L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 net2 input_stack net3 VDD sky130_fd_pr__pfet_01v8_hvt L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 net3 input_stack net4 VDD sky130_fd_pr__pfet_01v8_hvt L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 net4 input_stack net5 VDD sky130_fd_pr__pfet_01v8_hvt L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM6 net5 input_stack VDD VDD sky130_fd_pr__pfet_01v8_hvt L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:
*+  /foss/designs/hgu_goss/hgu/xschem/../../../hgu_goss/hgu/xschem/hgu_nfet_hvt_stack_in_delay.sym # of pins=3
** sym_path:
*+ /foss/designs/hgu_goss/hgu/xschem/../../../hgu_goss/hgu/xschem/hgu_nfet_hvt_stack_in_delay.sym
** sch_path:
*+ /foss/designs/hgu_goss/hgu/xschem/../../../hgu_goss/hgu/xschem/hgu_nfet_hvt_stack_in_delay.sch
.subckt hgu_nfet_hvt_stack_in_delay input_stack output_stack VSS
*.ipin VSS
*.ipin input_stack
*.iopin output_stack
XM1 output_stack input_stack net1 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 net1 input_stack net2 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 net2 input_stack net3 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 net3 input_stack net4 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 net4 input_stack net5 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM6 net5 input_stack net6 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM7 net6 input_stack net7 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM8 net7 input_stack net8 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM9 net8 input_stack net9 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM10 net9 input_stack net10 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM11 net10 input_stack net11 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM12 net11 input_stack net12 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM13 net12 input_stack net13 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM14 net13 input_stack net14 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM15 net14 input_stack net15 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM16 net15 input_stack VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.end
