magic
tech sky130A
magscale 1 2
timestamp 1697348449
<< error_p >>
rect -29 401 29 407
rect -29 367 -17 401
rect -29 361 29 367
rect -29 -367 29 -361
rect -29 -401 -17 -367
rect -29 -407 29 -401
<< nwell >>
rect -211 -539 211 539
<< pmos >>
rect -15 -320 15 320
<< pdiff >>
rect -73 308 -15 320
rect -73 -308 -61 308
rect -27 -308 -15 308
rect -73 -320 -15 -308
rect 15 308 73 320
rect 15 -308 27 308
rect 61 -308 73 308
rect 15 -320 73 -308
<< pdiffc >>
rect -61 -308 -27 308
rect 27 -308 61 308
<< nsubdiff >>
rect -175 469 -79 503
rect 79 469 175 503
rect -175 407 -141 469
rect 141 407 175 469
rect -175 -469 -141 -407
rect 141 -469 175 -407
rect -175 -503 -79 -469
rect 79 -503 175 -469
<< nsubdiffcont >>
rect -79 469 79 503
rect -175 -407 -141 407
rect 141 -407 175 407
rect -79 -503 79 -469
<< poly >>
rect -33 401 33 417
rect -33 367 -17 401
rect 17 367 33 401
rect -33 351 33 367
rect -15 320 15 351
rect -15 -351 15 -320
rect -33 -367 33 -351
rect -33 -401 -17 -367
rect 17 -401 33 -367
rect -33 -417 33 -401
<< polycont >>
rect -17 367 17 401
rect -17 -401 17 -367
<< locali >>
rect -175 469 -79 503
rect 79 469 175 503
rect -175 407 -141 469
rect 141 407 175 469
rect -33 367 -17 401
rect 17 367 33 401
rect -61 308 -27 324
rect -61 -324 -27 -308
rect 27 308 61 324
rect 27 -324 61 -308
rect -33 -401 -17 -367
rect 17 -401 33 -367
rect -175 -469 -141 -407
rect 141 -469 175 -407
rect -175 -503 -79 -469
rect 79 -503 175 -469
<< viali >>
rect -17 367 17 401
rect -61 -308 -27 308
rect 27 -308 61 308
rect -17 -401 17 -367
<< metal1 >>
rect -29 401 29 407
rect -29 367 -17 401
rect 17 367 29 401
rect -29 361 29 367
rect -67 308 -21 320
rect -67 -308 -61 308
rect -27 -308 -21 308
rect -67 -320 -21 -308
rect 21 308 67 320
rect 21 -308 27 308
rect 61 -308 67 308
rect 21 -320 67 -308
rect -29 -367 29 -361
rect -29 -401 -17 -367
rect 17 -401 29 -367
rect -29 -407 29 -401
<< properties >>
string FIXED_BBOX -158 -486 158 486
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 3.2 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
