* NGSPICE file created from hgu_sarlogic.ext - technology: sky130A

.subckt hgu_clk_async x3.S eob x2.IN x4.x7.SW x8.X x4.code[2] x4.code[1] x2.x10.A
+ x2.code[1] x2.code[2] x4.x2.SW x4.x10.A x2.x2.SW vss vdd
X0 x4.x5[7].floating x4.x10.Y x4.x9.output_stack vdd sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X1 x2.x9.output_stack x2.code[2] x2.x4[3].floating vss sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X2 x4.x3[1].floating x4.code[1] x4.x9.output_stack vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X3 x10.Y x10.A vss vss sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X4 a_1373_1841# eob vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_2200_1841# x3.S vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 x4.x9.output_stack x4.x10.Y x4.x5[7].floating vdd sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X7 x9.Y x9.A vss vss sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X8 a_n6207_n1487# x2.IN a_n6295_n1487# vss sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X9 a_n6207_n797# x2.IN a_n6295_n935# vss sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X10 a_n6182_1940# x8.X a_n6270_2078# vdd sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X11 vss x8.X a_n6207_n277# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X12 vss a_1771_1775# x3.X vss sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X13 a_n397_1077# x4.x9.output_stack vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X14 x4.x9.output_stack x4.code[2] x4.x4[3].floating vss sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X15 a_n6135_413# x8.X a_n6207_413# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X16 vdd x9.Y a_1363_798# vdd sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X17 a_1307_1909# x3.X a_944_1775# vss sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X18 a_818_1106# a_618_824# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X19 a_618_824# x10.Y vss vss sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X20 vss vdd a_2077_824# vss sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X21 a_n397_736# x4.x9.output_stack x10.A vss sky130_fd_pr__nfet_01v8 ad=0.0651 pd=0.73 as=0.122 ps=1.42 w=0.42 l=0.15
X22 a_2134_1909# x3.A0 a_1771_1775# vss sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X23 a_1159_798# x3.S vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X24 a_1403_1582# vss a_944_1775# vdd sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X25 a_n397_n2289# x9.A vss vdd sky130_fd_pr__pfet_01v8_hvt ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X26 a_2230_1582# vss a_1771_1775# vdd sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X27 a_1094_1190# a_305_798# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0819 ps=0.81 w=0.42 l=0.15
X28 a_1296_1190# a_1159_798# a_860_798# vdd sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X29 vss x9.Y a_724_824# vss sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.12 ps=1.08 w=0.42 l=0.15
X30 vdd x4.x7.SW x4.x6.SW vdd sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X31 a_618_824# x10.Y vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.154 ps=1.34 w=0.64 l=0.15
X32 a_n6207_n1# x8.X a_n6295_n1# vss sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X33 a_1363_798# a_1631_1008# a_1577_1106# vdd sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X34 x2.x4[3].floating x2.code[2] x2.x9.output_stack vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X35 a_n6207_689# x8.X a_n6295_551# vss sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X36 vss a_944_1775# x8.X vss sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X37 a_n397_n1948# x2.x9.output_stack x9.A vss sky130_fd_pr__nfet_01v8 ad=0.0651 pd=0.73 as=0.122 ps=1.42 w=0.42 l=0.15
X38 a_n6182_1664# x8.X a_n6270_1526# vdd sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X39 a_210_798# a_305_798# vss vss sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X40 a_n6182_n3152# x2.IN a_n6270_n3014# vdd sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X41 a_944_1775# vss a_1086_1909# vss sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X42 a_n397_1077# x10.A vss vdd sky130_fd_pr__pfet_01v8_hvt ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X43 a_n6135_n1073# x2.IN a_n6207_n1073# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X44 vdd x9.Y a_305_798# vdd sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.123 ps=1.17 w=0.42 l=0.15
X45 x2.x4[3].floating x2.code[2] x2.x9.output_stack vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X46 a_n6207_n277# x8.X a_n6295_n277# vss sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X47 vss a_305_798# x27.Q_N vss sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X48 a_n6135_n1349# x2.IN a_n6207_n1349# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X49 x10.Y x10.A vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X50 vss x9.A a_n397_n2289# vdd sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0651 ps=0.73 w=0.42 l=0.15
X51 a_n6207_n1073# x2.IN a_n6295_n1211# vss sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X52 x2.x9.output_stack x4.x7.SW x2.x7.floating vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X53 x4.x10.Y x4.x10.A vss vss sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X54 a_210_798# a_305_798# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X55 x4.x4[3].floating x4.code[2] x4.x9.output_stack vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X56 x2.x9.output_stack x2.IN a_n6270_n2738# vdd sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X57 vdd a_1373_1841# a_1403_1582# vdd sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X58 vdd a_305_798# x27.Q_N vdd sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X59 a_n6207_n1349# x2.IN a_n6295_n1487# vss sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X60 a_724_824# a_860_798# a_305_798# vss sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0864 ps=0.91 w=0.64 l=0.15
X61 x4.x9.output_stack x4.x10.Y x4.x5[7].floating vdd sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X62 a_n397_n2289# x2.x9.output_stack vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X63 a_n6135_n139# x8.X a_n6207_n139# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X64 a_2077_824# a_1159_798# a_1631_1008# vss sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X65 a_n397_736# x4.x9.output_stack vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X66 a_1159_798# x3.S vss vss sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X67 a_860_798# a_1159_798# a_1094_824# vss sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.066 ps=0.745 w=0.36 l=0.15
X68 vss x9.Y a_1499_824# vss sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.101 ps=0.99 w=0.42 l=0.15
X69 vss a_210_798# x3.A0 vss sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X70 x2.x9.output_stack x2.IN a_n6207_n1763# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X71 x4.x9.output_stack x8.X a_n6207_689# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X72 a_1913_1909# x3.S vss vss sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X73 a_n6207_275# x8.X a_n6295_275# vss sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X74 a_2077_824# a_1158_1098# a_1631_1008# vdd sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X75 a_n6207_n1763# x2.IN a_n6295_n1763# vss sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X76 vss a_1159_798# a_1158_1098# vss sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X77 a_305_798# a_618_824# a_724_824# vss sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X78 a_n397_n1948# x2.x9.output_stack vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X79 vss a_1363_798# a_1298_824# vss sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0935 ps=0.965 w=0.64 l=0.15
X80 x4.x9.output_stack x8.X a_n6270_1526# vdd sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X81 a_1086_1909# eob vss vss sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X82 x4.x5[7].floating x4.x10.Y x4.x9.output_stack vdd sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X83 x2.x9.output_stack x2.x6.SW x2.x6.floating vdd sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X84 a_n6207_n139# x8.X a_n6295_n277# vss sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X85 x9.Y x9.A vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X86 vss x4.x7.SW x4.x6.SW vss sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X87 x4.x9.output_stack x4.x10.Y x4.x5[7].floating vdd sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X88 a_n6135_n1073# x2.IN a_n6207_n935# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X89 vdd x2.IN a_n6270_n3290# vdd sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X90 x2.x2.floating x2.x2.SW x2.x9.output_stack vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.124 ps=1.43 w=0.42 l=0.15
X91 vdd a_1771_1775# x3.X vdd sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X92 a_1094_824# a_305_798# vss vss sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0588 ps=0.7 w=0.42 l=0.15
X93 a_305_798# a_860_798# a_818_1106# vdd sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0882 ps=1.05 w=0.84 l=0.15
X94 x4.x9.output_stack x4.x6.SW x4.x6.floating vdd sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X95 a_n6135_n139# x8.X a_n6207_n1# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X96 vdd a_1363_798# a_1296_1190# vdd sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X97 vss x4.x7.SW x2.x6.SW vss sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X98 x2.x9.output_stack x2.x10.Y x2.x5[7].floating vdd sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X99 a_n397_1077# x4.x9.output_stack x10.A vdd sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.122 ps=1.42 w=0.42 l=0.15
X100 x4.x4[3].floating x4.code[2] x4.x9.output_stack vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X101 a_n397_n1948# x9.A vdd vss sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X102 a_n6135_137# x8.X a_n6207_275# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X103 a_n6182_1940# x8.X a_n6270_1802# vdd sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X104 vdd a_2200_1841# a_2230_1582# vdd sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X105 a_1875_1190# a_1363_798# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X106 x2.x9.output_stack x2.x10.Y x2.x5[7].floating vdd sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X107 a_n6135_n1625# x2.IN a_n6207_n1625# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X108 a_n6207_137# x8.X a_n6295_n1# vss sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X109 a_1577_1106# a_618_824# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X110 vdd a_944_1775# x8.X vdd sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X111 x4.x9.output_stack x4.x7.SW x4.x7.floating vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X112 x4.x9.output_stack x4.code[1] x4.x3[1].floating vss sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X113 x2.x10.Y x2.x10.A vss vss sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X114 a_1298_824# a_1158_1098# a_860_798# vss sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.0711 ps=0.755 w=0.36 l=0.15
X115 a_n6182_n2876# x2.IN a_n6270_n3014# vdd sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X116 a_n6207_n935# x2.IN a_n6295_n935# vss sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X117 a_1771_1775# x3.A0 a_1913_1582# vdd sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X118 a_n6207_n1625# x2.IN a_n6295_n1763# vss sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X119 vdd x8.X a_n6270_2078# vdd sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X120 x2.x9.output_stack x2.x10.Y x2.x5[7].floating vdd sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X121 a_1913_1582# x3.S vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X122 a_1499_824# a_1631_1008# a_1363_798# vss sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0864 ps=0.91 w=0.64 l=0.15
X123 vdd x9.A a_n397_n1948# vss sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0651 ps=0.73 w=0.42 l=0.15
X124 x4.x5[7].floating x4.x10.Y x4.x9.output_stack vdd sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X125 x2.x9.output_stack x2.x10.Y x2.x5[7].floating vdd sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X126 x4.x9.output_stack x4.x10.Y x4.x5[7].floating vdd sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X127 a_944_1775# x3.X a_1086_1582# vdd sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X128 a_n6207_551# x8.X a_n6295_551# vss sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X129 a_1086_1582# eob vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X130 a_1363_798# a_618_824# a_1499_824# vss sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X131 a_1631_1008# a_1159_798# a_1875_1190# vdd sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X132 a_n6135_137# x8.X a_n6207_137# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X133 a_n6182_1664# x8.X a_n6270_1802# vdd sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X134 a_n6135_n1349# x2.IN a_n6207_n1211# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X135 a_1631_1008# a_1158_1098# a_1875_824# vss sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0671 ps=0.75 w=0.36 l=0.15
X136 a_1875_824# a_1363_798# vss vss sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.084 ps=0.82 w=0.42 l=0.15
X137 vdd x10.A a_n397_736# vss sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0651 ps=0.73 w=0.42 l=0.15
X138 a_n6207_n1211# x2.IN a_n6295_n1211# vss sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X139 vdd a_1159_798# a_1158_1098# vdd sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X140 a_1373_1841# eob vss vss sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X141 a_2200_1841# x3.S vss vss sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X142 a_n397_736# x10.A vdd vss sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X143 a_n397_n2289# x2.x9.output_stack x9.A vdd sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.122 ps=1.42 w=0.42 l=0.15
X144 x4.x5[7].floating x4.x10.Y x4.x9.output_stack vdd sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X145 x4.x9.output_stack x4.code[2] x4.x4[3].floating vss sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X146 a_n6182_n2876# x2.IN a_n6270_n2738# vdd sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X147 x2.x9.output_stack x2.code[1] x2.x3[1].floating vss sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X148 a_860_798# a_1158_1098# a_1094_1190# vdd sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0924 ps=0.86 w=0.42 l=0.15
X149 vdd x4.x7.SW x2.x6.SW vdd sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X150 x2.x5[7].floating x2.x10.Y x2.x9.output_stack vdd sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X151 a_n6135_413# x8.X a_n6207_551# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X152 vss a_1373_1841# a_1307_1909# vss sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X153 a_1771_1775# vss a_1913_1909# vss sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X154 vss a_2200_1841# a_2134_1909# vss sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X155 x2.x5[7].floating x2.x10.Y x2.x9.output_stack vdd sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X156 x2.x5[7].floating x2.x10.Y x2.x9.output_stack vdd sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X157 a_n6207_413# x8.X a_n6295_275# vss sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X158 x2.x10.Y x2.x10.A vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X159 vss x2.IN a_n6207_n797# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X160 vdd a_210_798# x3.A0 vdd sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X161 vdd vdd a_2077_824# vdd sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0662 ps=0.735 w=0.42 l=0.15
X162 x2.x5[7].floating x2.x10.Y x2.x9.output_stack vdd sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X163 x4.x2.floating x4.x2.SW x4.x9.output_stack vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.124 ps=1.43 w=0.42 l=0.15
X164 x4.x10.Y x4.x10.A vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X165 a_n6182_n3152# x2.IN a_n6270_n3290# vdd sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X166 vss x10.A a_n397_1077# vdd sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0651 ps=0.73 w=0.42 l=0.15
X167 x2.x9.output_stack x2.code[2] x2.x4[3].floating vss sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X168 x2.x3[1].floating x2.code[1] x2.x9.output_stack vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X169 a_n6135_n1625# x2.IN a_n6207_n1487# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
.ends

.subckt hgu_clk_sample set reset x2.x4.x7.SW x2.x4.code[2] x2.x4.code[1] x2.x1.code[2]
+ x2.x1.code[1] x2.x1.x2.SW x2.x2.code[2] x2.x2.code[1] x2.x3.code[2] x2.x3.code[1]
+ x2.x3.x2.SW x2.x1.x10.A x2.x3.x10.A sample_clk_b sample_clk clk x2.x2.x10.A x2.x4.x2.SW
+ x2.x4.x10.A x2.x2.x2.SW vdd vss
X0 a_11371_5456# x2.x1.IN a_11283_5456# vss sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X1 vss a_3106_6090# a_3041_6494# vss sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X2 x2.x4.x2.floating x2.x4.x2.SW x2.x4.x9.output_stack vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.124 ps=1.43 w=0.42 l=0.15
X3 a_4687_7397# x3.A a_4599_7535# vdd sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X4 x2.x1.x5[7].floating x2.x1.x10.Y x2.x1.x9.output_stack vdd sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X5 x7.A x2.x3.x9.output_stack a_4047_2819# vdd sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.0651 ps=0.73 w=0.42 l=0.15
X6 a_2325_6090# x1.x3.Y vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X7 a_10112_1680# x2.x3.IN a_10024_1818# vdd sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X8 x2.x4.x9.output_stack x2.x4.x10.Y x2.x4.x5[7].floating vdd sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X9 a_10472_6534# x2.x4.x9.output_stack x2.x1.IN vdd sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.122 ps=1.42 w=0.42 l=0.15
X10 a_3340_6116# a_2932_6494# a_3106_6090# vdd sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X11 a_10065_3897# x2.x3.IN a_9977_3897# vss sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X12 a_2325_6090# a_2151_6116# a_2465_6482# vss sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X13 a_11396_7121# x2.x1.IN a_11308_6983# vdd sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X14 x2.x1.x10.Y x2.x1.x10.A vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X15 x2.x4.x10.Y x2.x4.x10.A vss vss sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X16 a_2151_6116# a_1870_6122# a_2058_6116# vdd sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X17 a_4734_5594# x3.A a_4662_5594# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X18 x2.x2.x5[7].floating x2.x2.x10.Y x2.x2.x9.output_stack vdd sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X19 vss a_2678_2626# sample_clk vss sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X20 a_16846_3483# x2.x2.IN a_16774_3483# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X21 x2.x2.x6.SW x2.x4.x7.SW vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X22 vdd a_3106_6090# a_3813_6132# vdd sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X23 vdd x7.Y x3.Y vdd sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X24 x2.x3.x9.output_stack x2.x3.code[2] x2.x3.x4[3].floating vss sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X25 vdd a_2678_2626# sample_clk vdd sky130_fd_pr__pfet_01v8 ad=0.391 pd=3.14 as=0.208 ps=1.59 w=1.26 l=0.15
X26 a_17181_6534# x2.x1.x9.output_stack x2.x2.IN vdd sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.122 ps=1.42 w=0.42 l=0.15
X27 x3.A a_3813_6132# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X28 x2.x2.x7.floating x2.x4.x7.SW x2.x2.x9.output_stack vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X29 x2.x1.x9.output_stack x2.x1.x6.SW x2.x1.x6.floating vdd sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X30 a_10472_6193# x2.x1.IN vdd vss sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X31 vdd x2.x3.x10.A x2.x3.x10.Y vdd sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X32 vdd a_2678_2006# sample_clk_b vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.391 ps=3.14 w=1.26 l=0.15
X33 a_4662_5180# x3.A a_4574_5180# vss sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X34 vss x2.x1.IN a_11371_5180# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X35 a_16846_3759# x2.x2.IN a_16774_3759# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X36 a_4047_3022# x7.A vdd vss sky130_fd_pr__nfet_01v8 ad=0.0651 pd=0.73 as=0.0693 ps=0.75 w=0.42 l=0.15
X37 a_11371_5870# x2.x1.IN a_11283_5732# vss sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X38 x2.x1.x9.output_stack x2.x1.x10.Y x2.x1.x5[7].floating vdd sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X39 a_16774_4173# x2.x2.IN vss vss sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X40 x2.x3.x5[7].floating x2.x3.x10.Y x2.x3.x9.output_stack vdd sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X41 x2.x4.x9.output_stack x2.x4.code[2] x2.x4.x4[3].floating vss sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X42 a_4662_5456# x3.A a_4574_5456# vss sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X43 a_11443_5318# x2.x1.IN a_11371_5456# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X44 x2.x1.x5[7].floating x2.x1.x10.Y x2.x1.x9.output_stack vdd sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X45 a_16774_3345# x2.x2.IN a_16686_3345# vss sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X46 x2.x3.x9.output_stack x2.x3.x10.Y x2.x3.x5[7].floating vdd sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X47 x2.x4.x5[7].floating x2.x4.x10.Y x2.x4.x9.output_stack vdd sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X48 a_17181_6534# x2.x2.IN vss vdd sky130_fd_pr__pfet_01v8_hvt ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X49 x2.x1.x9.output_stack x2.x4.x7.SW x2.x1.x7.floating vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X50 vdd a_3056_2150# a_2678_2006# vdd sky130_fd_pr__pfet_01v8 ad=0.365 pd=3.1 as=0.365 ps=3.1 w=1.26 l=0.15
X51 x2.x3.x5[7].floating x2.x3.x10.Y x2.x3.x9.output_stack vdd sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X52 x2.x1.x9.output_stack x2.x1.x10.Y x2.x1.x5[7].floating vdd sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X53 x1.x4.Y reset vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X54 a_10137_3759# x2.x3.IN a_10065_3897# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X55 vss a_2678_2006# sample_clk_b vss sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X56 x2.x2.x9.output_stack x2.x2.x10.Y x2.x2.x5[7].floating vdd sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X57 x2.x1.x5[7].floating x2.x1.x10.Y x2.x1.x9.output_stack vdd sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X58 a_11371_6146# x2.x1.IN a_11283_6008# vss sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X59 a_4687_7121# x3.A a_4599_6983# vdd sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X60 x2.x2.x4[3].floating x2.x2.code[2] x2.x2.x9.output_stack vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X61 vdd x2.x4.x7.SW x2.x1.x6.SW vdd sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X62 a_11371_5318# x2.x1.IN a_11283_5180# vss sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X63 a_10112_2232# x2.x3.IN a_10024_2094# vdd sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X64 a_4047_2819# x7.A vss vdd sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.0693 ps=0.75 w=0.42 l=0.15
X65 x2.x2.x9.output_stack x2.x2.code[2] x2.x2.x4[3].floating vss sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X66 a_2058_6116# x1.x2.D vss vss sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X67 a_10065_3483# x2.x3.IN a_9977_3345# vss sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X68 vss clk a_1704_6122# vss sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X69 a_10472_6193# x2.x4.x9.output_stack vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X70 x2.x1.x9.output_stack x2.x1.code[1] x2.x1.x3[1].floating vss sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X71 x2.x2.x6.floating x2.x2.x6.SW x2.x2.x9.output_stack vdd sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X72 vss x3.A a_4662_5180# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X73 a_4662_5870# x3.A a_4574_5732# vss sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X74 a_11443_5870# x2.x1.IN a_11371_5870# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X75 a_10065_3759# x2.x3.IN a_9977_3621# vss sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X76 x2.x2.x4[3].floating x2.x2.code[2] x2.x2.x9.output_stack vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X77 vdd a_3056_2936# a_2678_2626# vdd sky130_fd_pr__pfet_01v8 ad=0.365 pd=3.1 as=0.365 ps=3.1 w=1.26 l=0.15
X78 vss a_2325_6090# a_2259_6494# vss sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X79 a_3106_6090# x1.x3.Y vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X80 x2.x4.x9.output_stack x2.x4.x10.Y x2.x4.x5[7].floating vdd sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X81 a_16846_4035# x2.x2.IN a_16774_4173# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X82 x2.x4.x5[7].floating x2.x4.x10.Y x2.x4.x9.output_stack vdd sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X83 a_17181_6193# x2.x1.x9.output_stack vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X84 a_4734_5318# x3.A a_4662_5456# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X85 x2.x3.x6.SW x2.x4.x7.SW vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X86 x2.x3.x9.output_stack x2.x3.x10.Y x2.x3.x5[7].floating vdd sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X87 sample_clk a_2678_2626# vss vss sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X88 vdd a_3106_6090# a_3018_6116# vdd sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X89 x2.x4.x9.output_stack x2.x4.x7.SW x2.x4.x7.floating vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X90 a_16846_3207# x2.x2.IN a_16774_3345# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X91 vss x2.x2.x9.output_stack a_10756_3022# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X92 sample_clk a_2678_2626# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X93 vss x7.A x7.Y vss sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X94 a_3106_6090# a_2932_6494# a_3222_6482# vss sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X95 vdd x2.x1.IN a_10472_6193# vss sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0651 ps=0.73 w=0.42 l=0.15
X96 a_11371_5732# x2.x1.IN a_11283_5732# vss sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X97 x2.x3.x9.output_stack x2.x3.x10.Y x2.x3.x5[7].floating vdd sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X98 vdd x7.A a_4047_3022# vss sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X99 a_11396_7397# x2.x1.IN a_11308_7259# vdd sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X100 a_3222_6482# x1.x3.Y vss vss sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X101 x1.x2.D a_3106_6090# vss vss sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X102 a_4662_6146# x3.A a_4574_6008# vss sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X103 x2.x1.x9.output_stack x2.x1.IN a_11371_6146# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X104 vdd a_2619_6316# a_2569_6116# vdd sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X105 x2.x3.x4[3].floating x2.x3.code[2] x2.x3.x9.output_stack vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X106 vdd x2.x4.x7.SW x2.x4.x6.SW vdd sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X107 a_4662_5318# x3.A a_4574_5180# vss sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X108 a_16774_4035# x2.x2.IN a_16686_3897# vss sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X109 a_11443_5318# x2.x1.IN a_11371_5318# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X110 a_10472_6534# x2.x1.IN vss vdd sky130_fd_pr__pfet_01v8_hvt ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X111 x2.x4.x3[1].floating x2.x4.code[1] x2.x4.x9.output_stack vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X112 a_10137_3483# x2.x3.IN a_10065_3483# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X113 x2.x2.x9.output_stack x2.x2.code[1] x2.x2.x3[1].floating vss sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X114 a_16774_3207# x2.x2.IN x2.x2.x9.output_stack vss sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X115 x2.x1.x5[7].floating x2.x1.x10.Y x2.x1.x9.output_stack vdd sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X116 vdd x2.x2.IN a_17181_6193# vss sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0651 ps=0.73 w=0.42 l=0.15
X117 a_16821_1956# x2.x2.IN a_16733_2094# vdd sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X118 vdd x2.x2.x9.output_stack a_10756_2819# vdd sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X119 a_2465_6482# a_2619_6316# a_2325_6090# vss sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X120 x2.x4.x9.output_stack x2.x4.code[1] x2.x4.x3[1].floating vss sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X121 x2.x2.x5[7].floating x2.x2.x10.Y x2.x2.x9.output_stack vdd sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X122 x2.x1.x9.output_stack x2.x1.code[2] x2.x1.x4[3].floating vss sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X123 x2.x2.x9.output_stack x2.x2.x2.SW x2.x2.x2.floating vss sky130_fd_pr__nfet_01v8 ad=0.124 pd=1.43 as=0.122 ps=1.42 w=0.42 l=0.15
X124 x2.x1.x4[3].floating x2.x1.code[2] x2.x1.x9.output_stack vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X125 a_4734_5870# x3.A a_4662_5870# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X126 a_10137_3759# x2.x3.IN a_10065_3759# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X127 a_2235_6116# a_1704_6122# a_2151_6116# vdd sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X128 a_3553_3025# x3.A x3.Y vss sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X129 a_11371_6008# x2.x1.IN a_11283_6008# vss sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X130 a_10065_4173# x2.x3.IN vss vss sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X131 vss x7.A a_4047_2819# vdd sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X132 vdd a_2619_6316# a_3340_6116# vdd sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X133 a_10065_3345# x2.x3.IN a_9977_3345# vss sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X134 vss x3.Y a_3056_2936# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X135 a_1870_6122# a_1704_6122# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X136 x2.x1.x9.output_stack x2.x1.IN a_11308_6983# vdd sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X137 a_4662_5732# x3.A a_4574_5732# vss sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X138 a_11443_5594# x2.x1.IN a_11371_5732# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X139 a_4687_7397# x3.A a_4599_7259# vdd sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X140 x2.x4.x9.output_stack x3.A a_4662_6146# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X141 x1.x3.Y set vss vss sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X142 a_16774_3621# x2.x2.IN a_16686_3621# vss sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X143 vss x2.x2.x10.A x2.x2.x10.Y vss sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X144 x2.x4.x9.output_stack x2.x4.x6.SW x2.x4.x6.floating vdd sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X145 a_16846_4035# x2.x2.IN a_16774_4035# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X146 a_4734_5318# x3.A a_4662_5318# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X147 vss a_2678_2626# sample_clk vss sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X148 a_16821_1680# x2.x2.IN vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X149 x2.x3.x9.output_stack x2.x3.code[1] x2.x3.x3[1].floating vss sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X150 a_16846_3207# x2.x2.IN a_16774_3207# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X151 x2.x3.IN x2.x2.x9.output_stack a_10756_3022# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0651 ps=0.73 w=0.42 l=0.15
X152 a_2058_6116# x1.x2.D vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X153 vdd a_2678_2626# sample_clk vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.391 ps=3.14 w=1.26 l=0.15
X154 vss a_3056_2936# a_2678_2626# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X155 x2.x4.x9.output_stack x2.x4.code[2] x2.x4.x4[3].floating vss sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X156 x2.x3.x9.output_stack x2.x3.x2.SW x2.x3.x2.floating vss sky130_fd_pr__nfet_01v8 ad=0.124 pd=1.43 as=0.122 ps=1.42 w=0.42 l=0.15
X157 x2.x4.x10.Y x2.x4.x10.A vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X158 a_3018_6116# a_1870_6122# a_2932_6494# vdd sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X159 x2.x4.x4[3].floating x2.x4.code[2] x2.x4.x9.output_stack vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X160 a_16821_1956# x2.x2.IN a_16733_1818# vdd sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X161 a_11396_7121# x2.x1.IN a_11308_7259# vdd sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X162 a_2932_6494# a_1870_6122# a_2837_6438# vss sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X163 x2.x3.x5[7].floating x2.x3.x10.Y x2.x3.x9.output_stack vdd sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X164 a_4662_6008# x3.A a_4574_6008# vss sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X165 a_11443_5870# x2.x1.IN a_11371_6008# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X166 vdd a_2325_6090# a_2235_6116# vdd sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X167 x2.x1.x9.output_stack x2.x1.x10.Y x2.x1.x5[7].floating vdd sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X168 a_10137_4035# x2.x3.IN a_10065_4173# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X169 x2.x3.x7.floating x2.x4.x7.SW x2.x3.x9.output_stack vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X170 vss x2.x1.IN a_10472_6534# vdd sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0651 ps=0.73 w=0.42 l=0.15
X171 a_10137_3207# x2.x3.IN a_10065_3345# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X172 x2.x1.x10.Y x2.x1.x10.A vss vss sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X173 a_3041_6494# a_1704_6122# a_2932_6494# vss sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X174 x2.x4.x9.output_stack x3.A a_4599_6983# vdd sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X175 x2.x1.x2.floating x2.x1.x2.SW x2.x1.x9.output_stack vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.124 ps=1.43 w=0.42 l=0.15
X176 a_4734_5594# x3.A a_4662_5732# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X177 x2.x2.x9.output_stack x2.x2.code[2] x2.x2.x4[3].floating vss sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X178 a_16846_3483# x2.x2.IN a_16774_3621# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X179 x2.x2.x9.output_stack x2.x2.x10.Y x2.x2.x5[7].floating vdd sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X180 x2.x3.IN x2.x2.x9.output_stack a_10756_2819# vdd sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.0651 ps=0.73 w=0.42 l=0.15
X181 a_10756_3022# x2.x3.IN vdd vss sky130_fd_pr__nfet_01v8 ad=0.0651 pd=0.73 as=0.0693 ps=0.75 w=0.42 l=0.15
X182 a_2151_6116# a_1704_6122# a_2058_6116# vss sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X183 vss x2.x2.IN a_17181_6534# vdd sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0651 ps=0.73 w=0.42 l=0.15
X184 vdd x1.x4.Y a_2619_6316# vdd sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X185 a_10065_4035# x2.x3.IN a_9977_3897# vss sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X186 x2.x3.x6.floating x2.x3.x6.SW x2.x3.x9.output_stack vdd sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X187 a_10065_3207# x2.x3.IN x2.x3.x9.output_stack vss sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X188 vdd x7.A x7.Y vdd sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X189 vdd x2.x1.IN a_11308_7535# vdd sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X190 vss x1.x4.Y a_2619_6316# vss sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X191 x2.x4.x9.output_stack x2.x4.x10.Y x2.x4.x5[7].floating vdd sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X192 a_10112_1956# x2.x3.IN a_10024_2094# vdd sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X193 vdd a_2678_2006# sample_clk_b vdd sky130_fd_pr__pfet_01v8 ad=0.391 pd=3.14 as=0.208 ps=1.59 w=1.26 l=0.15
X194 a_2790_6116# a_2325_6090# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X195 x2.x4.x5[7].floating x2.x4.x10.Y x2.x4.x9.output_stack vdd sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X196 x2.x2.x6.SW x2.x4.x7.SW vss vss sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X197 a_4687_7121# x3.A a_4599_7259# vdd sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X198 vss x2.x3.x9.output_stack a_4047_3022# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X199 x2.x2.x5[7].floating x2.x2.x10.Y x2.x2.x9.output_stack vdd sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X200 x3.A a_3813_6132# vss vss sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X201 a_4734_5870# x3.A a_4662_6008# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X202 vss x2.x3.x10.A x2.x3.x10.Y vss sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X203 x2.x3.x9.output_stack x2.x3.code[2] x2.x3.x4[3].floating vss sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X204 a_16821_2232# x2.x2.IN x2.x2.x9.output_stack vdd sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X205 a_2837_6438# a_2325_6090# vss vss sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X206 x1.x4.Y reset vss vss sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X207 a_2465_6482# x1.x3.Y vss vss sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X208 x1.x2.D a_3106_6090# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X209 x2.x3.x4[3].floating x2.x3.code[2] x2.x3.x9.output_stack vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X210 vss x7.Y a_3553_3025# vss sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X211 vss x2.x4.x7.SW x2.x1.x6.SW vss sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X212 x2.x1.x9.output_stack x2.x1.x10.Y x2.x1.x5[7].floating vdd sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X213 a_10756_2819# x2.x3.IN vss vdd sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.0693 ps=0.75 w=0.42 l=0.15
X214 a_2569_6116# a_2151_6116# a_2325_6090# vdd sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X215 x2.x1.x9.output_stack x2.x1.code[2] x2.x1.x4[3].floating vss sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X216 a_16821_1680# x2.x2.IN a_16733_1818# vdd sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X217 vss a_2678_2006# sample_clk_b vss sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X218 x2.x2.x9.output_stack x2.x2.x10.Y x2.x2.x5[7].floating vdd sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X219 a_16774_3897# x2.x2.IN a_16686_3897# vss sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X220 x3.Y x3.A vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X221 x2.x2.x3[1].floating x2.x2.code[1] x2.x2.x9.output_stack vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X222 vss a_3106_6090# a_3813_6132# vss sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X223 x2.x4.x5[7].floating x2.x4.x10.Y x2.x4.x9.output_stack vdd sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X224 x2.x3.x9.output_stack x2.x3.x10.Y x2.x3.x5[7].floating vdd sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X225 a_10065_3621# x2.x3.IN a_9977_3621# vss sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X226 vdd x2.x3.x9.output_stack a_4047_2819# vdd sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X227 x2.x3.x5[7].floating x2.x3.x10.Y x2.x3.x9.output_stack vdd sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X228 vdd x3.Y a_3056_2936# vdd sky130_fd_pr__pfet_01v8 ad=0.406 pd=3.38 as=0.406 ps=3.38 w=1.4 l=0.15
X229 a_10472_6193# x2.x4.x9.output_stack x2.x1.IN vss sky130_fd_pr__nfet_01v8 ad=0.0651 pd=0.73 as=0.122 ps=1.42 w=0.42 l=0.15
X230 x2.x1.x4[3].floating x2.x1.code[2] x2.x1.x9.output_stack vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X231 a_11371_5594# x2.x1.IN a_11283_5456# vss sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X232 a_10137_4035# x2.x3.IN a_10065_4035# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X233 a_10137_3207# x2.x3.IN a_10065_3207# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X234 a_10112_1680# x2.x3.IN vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X235 vdd x3.A a_4599_7535# vdd sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X236 x2.x2.x9.output_stack x2.x2.x10.Y x2.x2.x5[7].floating vdd sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X237 a_10472_6534# x2.x4.x9.output_stack vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X238 a_1870_6122# a_1704_6122# vss vss sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X239 a_17181_6193# x2.x1.x9.output_stack x2.x2.IN vss sky130_fd_pr__nfet_01v8 ad=0.0651 pd=0.73 as=0.122 ps=1.42 w=0.42 l=0.15
X240 a_10112_1956# x2.x3.IN a_10024_1818# vdd sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X241 vdd x2.x3.IN a_10756_3022# vss sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X242 a_2259_6494# a_1870_6122# a_2151_6116# vss sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X243 vdd clk a_1704_6122# vdd sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X244 a_11396_7397# x2.x1.IN a_11308_7535# vdd sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X245 a_17181_6534# x2.x1.x9.output_stack vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X246 vss x2.x4.x7.SW x2.x4.x6.SW vss sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X247 x2.x4.x9.output_stack x2.x4.x10.Y x2.x4.x5[7].floating vdd sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X248 sample_clk_b a_2678_2006# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X249 x2.x3.x6.SW x2.x4.x7.SW vss vss sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X250 x2.x1.x3[1].floating x2.x1.code[1] x2.x1.x9.output_stack vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X251 vdd x2.x2.x10.A x2.x2.x10.Y vdd sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X252 a_17181_6193# x2.x2.IN vdd vss sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X253 a_16846_3759# x2.x2.IN a_16774_3897# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X254 x3.Y vdd a_3056_2150# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X255 x2.x3.x3[1].floating x2.x3.code[1] x2.x3.x9.output_stack vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X256 a_3222_6482# a_2619_6316# a_3106_6090# vss sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X257 x7.A x2.x3.x9.output_stack a_4047_3022# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0651 ps=0.73 w=0.42 l=0.15
X258 a_10137_3483# x2.x3.IN a_10065_3621# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X259 a_16821_2232# x2.x2.IN a_16733_2094# vdd sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X260 x2.x4.x4[3].floating x2.x4.code[2] x2.x4.x9.output_stack vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X261 a_4662_5594# x3.A a_4574_5456# vss sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X262 a_11443_5594# x2.x1.IN a_11371_5594# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X263 x3.Y vss a_3056_2150# vdd sky130_fd_pr__pfet_01v8 ad=0.551 pd=4.38 as=0.551 ps=4.38 w=1.9 l=0.15
X264 a_16774_3483# x2.x2.IN a_16686_3345# vss sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X265 vss a_3056_2150# a_2678_2006# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X266 x1.x3.Y set vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X267 a_2932_6494# a_1704_6122# a_2790_6116# vdd sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X268 vss x2.x3.IN a_10756_2819# vdd sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X269 a_11371_5180# x2.x1.IN a_11283_5180# vss sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X270 a_16774_3759# x2.x2.IN a_16686_3621# vss sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X271 sample_clk_b a_2678_2006# vss vss sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X272 a_10112_2232# x2.x3.IN x2.x3.x9.output_stack vdd sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X273 x2.x2.x5[7].floating x2.x2.x10.Y x2.x2.x9.output_stack vdd sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
.ends

.subckt hgu_sarlogic_8bit_logic sel_bit[0] sel_bit[1] x1.A eob x6.A D[7] D[6] x30.D
+ D[5] x48.D x33.D x45.D x36.D x42.D x39.D D[2] D[3] D[1] D[4] D[0] x2.A VSS VDD
X0 VDD a_10680_2340# D[3] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X1 VDD a_8289_4086# x45.D VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X2 VDD D[0] a_8236_3239# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3 VDD a_2389_5648# eob VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.135 ps=1.27 w=1 l=0.15
X4 a_12030_3213# a_11856_3239# a_12146_3239# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X5 VDD a_1338_5674# x5.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6 a_4971_4801# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X7 a_2147_5083# a_1682_4775# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X8 a_1822_4801# x4.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X9 a_11330_2340# a_11628_2640# a_11564_2732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0924 ps=0.86 w=0.42 l=0.15
X10 VSS a_12030_3213# a_12737_3239# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X11 a_4213_3239# a_4367_3213# a_4073_3213# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X12 a_8591_4801# x33.D VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X13 a_9710_4296# a_9238_4086# a_9954_4478# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X14 VSS x30.Q_N a_7185_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.101 ps=0.99 w=0.42 l=0.15
X15 VDD a_11250_4775# a_11160_5167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X16 VSS a_5992_4086# x45.Q_N VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X17 a_3599_2340# a_3912_2366# a_4018_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X18 x72.Q_N a_7246_3213# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X19 VSS x27.Q_N a_4018_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.12 ps=1.08 w=0.42 l=0.15
X20 a_4854_3213# x77.Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X21 a_7072_3239# a_5844_3239# a_6930_3521# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X22 a_9442_4086# a_8697_4112# a_9578_4112# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X23 VSS x4.X a_9151_3213# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X24 VDD a_7246_3213# a_7158_3605# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X25 VDD a_5897_4086# x48.D VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X26 a_11089_4112# x4.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.154 ps=1.34 w=0.64 l=0.15
X27 a_4793_2366# a_4925_2550# a_4657_2340# VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0864 ps=0.91 w=0.64 l=0.15
X28 VDD x75.Q a_5844_3239# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X29 a_6978_4801# a_6466_4775# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X30 a_4388_2732# a_3599_2340# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0819 ps=0.81 w=0.42 l=0.15
X31 a_2788_5674# x42.D VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.107 ps=1 w=0.42 l=0.15
X32 a_10794_3239# a_10628_3239# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X33 VSS D[0] a_8236_3239# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X34 VDD x4.X a_4368_4775# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X35 a_9465_4801# a_8403_4801# a_9370_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X36 VSS a_1511_4112# x4.X VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X37 a_12048_4394# a_11089_4112# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X38 a_9101_3521# a_8683_3605# a_8857_3213# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X39 a_7247_4775# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X40 VDD a_6846_4086# a_6845_4386# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X41 VSS x20.Q_N a_1626_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.12 ps=1.08 w=0.42 l=0.15
X42 D[2] a_12737_3239# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X43 a_11250_4775# a_11076_5167# a_11390_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X44 a_4680_3239# a_3452_3239# a_4538_3521# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X45 a_2479_2648# a_1520_2366# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X46 VDD a_4854_3213# a_4766_3605# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X47 a_11184_4801# a_10795_4801# a_11076_5167# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X48 a_2784_5996# x42.D VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=0.995 as=0.154 ps=1.34 w=0.64 l=0.15
X49 a_4593_4112# a_4453_4386# a_4155_4086# VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.0711 ps=0.755 w=0.36 l=0.15
X50 a_1996_2732# a_1207_2340# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0819 ps=0.81 w=0.42 l=0.15
X51 a_7181_3239# a_5844_3239# a_7072_3239# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X52 a_6198_3239# x7.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X53 x4.X a_1511_4112# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X54 a_2265_2340# a_1520_2366# a_2401_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X55 a_12031_4775# a_11857_4801# a_12147_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X56 VSS x75.Q a_5844_3239# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X57 VDD VDD a_1976_4775# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X58 VSS a_7050_4086# a_6985_4112# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0935 ps=0.965 w=0.64 l=0.15
X59 a_1762_2340# a_2060_2640# a_1996_2732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0924 ps=0.86 w=0.42 l=0.15
X60 VDD x45.D a_2969_6040# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.138 ps=1.16 w=0.64 l=0.15
X61 a_2883_5674# a_2853_5648# a_2788_5674# VSS sky130_fd_pr__nfet_01v8 ad=0.072 pd=0.76 as=0.066 ps=0.745 w=0.36 l=0.15
X62 a_7562_4478# a_7050_4086# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X63 a_10775_2340# a_11088_2366# a_11194_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X64 a_6504_2648# a_6304_2366# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X65 a_4214_4801# a_4368_4775# a_4074_4775# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X66 VSS x36.Q_N a_11194_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.12 ps=1.08 w=0.42 l=0.15
X67 a_10794_3239# a_10628_3239# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X68 a_1511_4112# x4.A VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X69 a_4855_4775# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X70 a_7073_4801# a_5845_4801# a_6931_5083# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X71 VDD a_4454_4086# a_4453_4386# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X72 VDD a_7247_4775# a_7159_5167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X73 x4.A a_897_4112# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X74 VDD a_1338_5674# x5.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X75 x30.Q_N a_7247_4775# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X76 x4.X a_1511_4112# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X77 a_12345_2732# a_11833_2340# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X78 VSS x48.D a_5372_4112# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X79 a_8803_4112# a_8939_4086# a_8384_4086# VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0864 ps=0.91 w=0.64 l=0.15
X80 VSS x4.X a_9152_4775# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X81 a_3806_3239# VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X82 VDD x20.Q_N a_1207_2340# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.123 ps=1.17 w=0.42 l=0.15
X83 VSS x45.D a_2993_5674# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0786 ps=0.805 w=0.42 l=0.15
X84 VSS VDD a_8803_4112# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.12 ps=1.08 w=0.42 l=0.15
X85 VSS a_10776_4086# x39.Q_N VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X86 a_6291_3605# a_5844_3239# a_6198_3239# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X87 x75.Q_N a_4854_3213# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X88 VSS x5.X a_8237_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X89 VSS a_6465_3213# a_6399_3239# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X90 a_1822_4801# a_1976_4775# a_1682_4775# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X91 VDD a_10775_2340# x63.Q_N VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X92 a_9102_5083# a_8684_5167# a_8858_4775# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X93 a_11856_3239# a_10628_3239# a_11714_3521# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X94 a_4681_4801# a_3453_4801# a_4539_5083# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X95 VDD a_4855_4775# a_4767_5167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X96 a_9953_2366# a_9441_2340# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.084 ps=0.82 w=0.42 l=0.15
X97 x39.D a_12738_4801# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X98 a_11769_4112# a_11629_4386# a_11331_4086# VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.0711 ps=0.755 w=0.36 l=0.15
X99 a_1112_2340# a_1207_2340# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X100 x7.X a_929_3238# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X101 a_2579_4801# x4.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X102 a_4155_4086# a_4453_4386# a_4389_4478# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0924 ps=0.86 w=0.42 l=0.15
X103 a_7480_3521# a_7072_3239# a_7246_3213# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X104 VSS VDD a_9578_4112# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.101 ps=0.99 w=0.42 l=0.15
X105 a_5992_4086# a_6305_4112# a_6411_4112# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X106 VDD x7.X a_12547_2366# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0662 ps=0.735 w=0.42 l=0.15
X107 a_6199_4801# x30.D VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X108 a_7182_4801# a_5845_4801# a_7073_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X109 VSS VDD a_6411_4112# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.12 ps=1.08 w=0.42 l=0.15
X110 VDD x4.X a_6759_3213# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X111 x33.Q_N a_9639_4775# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X112 VSS x27.Q_N a_4793_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.101 ps=0.99 w=0.42 l=0.15
X113 a_3899_3605# a_3452_3239# a_3806_3239# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X114 VSS x5.X a_5845_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X115 D[1] a_10345_3239# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X116 a_6710_5083# a_6292_5167# a_6466_4775# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X117 a_11195_4112# a_11331_4086# a_10776_4086# VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0864 ps=0.91 w=0.64 l=0.15
X118 a_6375_3605# a_5844_3239# a_6291_3605# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X119 a_2969_6040# a_2853_5648# a_2883_5674# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.16 as=0.0567 ps=0.69 w=0.42 l=0.15
X120 a_8288_2340# a_8383_2340# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X121 a_10795_4801# a_10629_4801# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X122 a_7050_4086# a_6305_4112# a_7186_4112# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X123 a_11965_3239# a_10628_3239# a_11856_3239# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X124 a_12102_4296# a_11629_4386# a_12346_4112# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0671 ps=0.75 w=0.36 l=0.15
X125 VSS a_2463_4775# a_3170_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X126 a_11970_4112# a_12102_4296# a_11834_4086# VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0864 ps=0.91 w=0.64 l=0.15
X127 VDD a_3505_4086# x48.Q VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X128 a_8590_3239# x7.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X129 VDD VSS a_3452_3239# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X130 x4.X a_1511_4112# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X131 a_4113_4394# a_3913_4112# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X132 VSS a_11834_4086# a_11769_4112# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0935 ps=0.965 w=0.64 l=0.15
X133 a_3807_4801# x27.D VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X134 a_4790_4801# a_3453_4801# a_4681_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X135 VSS x20.Q_N a_2401_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.101 ps=0.99 w=0.42 l=0.15
X136 VDD a_929_3238# x7.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X137 a_1511_4112# x4.A VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X138 a_11564_2366# a_10775_2340# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0588 ps=0.7 w=0.42 l=0.15
X139 a_7763_2366# a_6844_2640# a_7317_2550# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X140 a_11714_3521# a_11249_3213# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X141 a_11857_4801# a_10629_4801# a_11715_5083# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X142 x4.A a_897_4112# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X143 a_6292_5167# a_5845_4801# a_6199_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X144 VDD a_1207_2340# x51.Q_N VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X145 a_3983_3605# a_3452_3239# a_3899_3605# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X146 a_2389_5648# a_3258_5648# a_2883_5674# VSS sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X147 a_5896_2340# a_5991_2340# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X148 VSS a_6466_4775# a_6400_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X149 a_4658_4086# a_3913_4112# a_4794_4112# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X150 VDD a_2463_4775# a_3170_4801# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X151 a_7481_5083# a_7073_4801# a_7247_4775# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X152 a_9237_2340# D[3] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X153 VDD x1.A a_621_4112# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X154 a_9173_4112# a_8384_4086# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0588 ps=0.7 w=0.42 l=0.15
X155 VDD x7.X a_2979_2366# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0662 ps=0.735 w=0.42 l=0.15
X156 VDD a_11833_2340# a_11766_2732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X157 VSS VSS a_3452_3239# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X158 VDD a_9442_4086# a_9375_4478# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X159 VDD x30.Q_N a_7049_2340# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X160 a_4317_3521# a_3899_3605# a_4073_3213# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X161 a_6376_5167# a_5845_4801# a_6292_5167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X162 a_3900_5167# a_3453_4801# a_3807_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X163 VSS a_8383_2340# x60.Q_N VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X164 a_11249_3213# x39.Q_N VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X165 x7.X a_929_3238# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X166 a_1227_4801# a_1061_4801# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X167 a_4074_4775# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X168 a_8997_3239# x42.Q_N VSS VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X169 a_8591_4801# x33.D VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X170 a_11289_4394# a_11089_4112# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X171 a_1511_4112# x4.A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X172 x4.X a_1511_4112# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X173 x75.Q a_5561_3239# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X174 a_11966_4801# a_10629_4801# a_11857_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X175 a_9376_2366# a_9236_2640# a_8938_2340# VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.0711 ps=0.755 w=0.36 l=0.15
X176 eob a_2389_5648# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X177 a_6781_4112# a_5992_4086# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0588 ps=0.7 w=0.42 l=0.15
X178 x77.Y eob VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X179 x5.X a_1338_5674# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X180 a_9237_2340# D[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X181 a_11715_5083# a_11250_4775# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X182 x27.Q_N a_4855_4775# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X183 a_3984_5167# a_3453_4801# a_3900_5167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X184 a_8791_3239# a_8402_3239# a_8683_3605# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X185 a_11089_4112# x4.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X186 a_5991_2340# a_6546_2340# a_6504_2648# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0882 ps=1.05 w=0.84 l=0.15
X187 a_11075_3605# a_10794_3239# a_10982_3239# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X188 VDD x48.D a_5372_4112# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0662 ps=0.735 w=0.42 l=0.15
X189 VDD a_11629_2340# a_11628_2640# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X190 a_9638_3213# a_9464_3239# a_9754_3239# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X191 a_5088_3521# a_4680_3239# a_4854_3213# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X192 x4.X a_1511_4112# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X193 VDD VDD a_9442_4086# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X194 a_6984_2366# a_6844_2640# a_6546_2340# VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.0711 ps=0.755 w=0.36 l=0.15
X195 VDD x4.X a_4367_3213# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X196 VDD a_929_3238# x7.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X197 a_7318_4296# a_6846_4086# a_7562_4478# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X198 VSS a_9441_2340# a_9376_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0935 ps=0.965 w=0.64 l=0.15
X199 a_4318_5083# a_3900_5167# a_4074_4775# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X200 x36.D a_10346_4801# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X201 VDD a_1511_4112# x4.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X202 a_12548_4112# a_11629_4386# a_12102_4296# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X203 a_12101_2550# a_11629_2340# a_12345_2732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X204 VSS x5.X a_3453_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X205 a_11250_4775# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X206 a_4453_2340# D[5] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X207 a_3373_5674# a_3258_5648# a_2389_5648# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.6 as=0.0729 ps=0.81 w=0.54 l=0.15
X208 VSS x4.X a_6759_3213# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X209 VSS x1.A a_621_4112# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X210 a_1762_2340# a_2061_2340# a_1996_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.066 ps=0.745 w=0.36 l=0.15
X211 a_9550_3605# a_8402_3239# a_9464_3239# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X212 a_8998_4801# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X213 x4.X a_1511_4112# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X214 a_7049_2340# a_7317_2550# a_7263_2648# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X215 a_6198_3239# x7.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X216 VSS x7.X a_7763_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X217 a_2398_4801# a_1061_4801# a_2289_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X218 VSS a_11629_2340# a_11628_2640# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X219 VDD a_6759_3213# a_7480_3521# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X220 a_3877_5674# a_2853_5648# a_3373_5674# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.072 ps=0.76 w=0.36 l=0.15
X221 a_9656_4394# a_8697_4112# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X222 a_7185_2366# a_7317_2550# a_7049_2340# VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0864 ps=0.91 w=0.64 l=0.15
X223 a_10155_2366# a_9237_2340# a_9709_2550# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X224 a_1926_5083# a_1508_5167# a_1682_4775# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X225 a_9370_4801# a_8858_4775# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X226 VDD VDD a_11834_4086# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X227 a_3504_2340# a_3599_2340# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X228 a_11076_5167# a_10795_4801# a_10983_4801# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X229 a_8792_4801# a_8403_4801# a_8684_5167# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X230 a_5089_5083# a_4681_4801# a_4855_4775# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X231 x4.X a_1511_4112# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X232 VDD a_2061_2340# a_2060_2640# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X233 a_3671_5674# x48.Q VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0819 ps=0.81 w=0.42 l=0.15
X234 a_4453_2340# D[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X235 a_4657_2340# a_4925_2550# a_4871_2648# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X236 a_3806_3239# VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X237 x5.X a_1338_5674# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X238 a_9639_4775# a_9465_4801# a_9755_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X239 VDD a_12030_3213# a_12737_3239# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X240 a_4970_3239# a_4367_3213# a_4854_3213# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X241 a_8857_3213# a_8683_3605# a_8997_3239# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X242 a_3600_4086# a_4155_4086# a_4113_4394# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0882 ps=1.05 w=0.84 l=0.15
X243 a_8383_2340# a_8696_2366# a_8802_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X244 VDD a_6465_3213# a_6375_3605# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X245 VSS x48.D a_3877_5674# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.066 ps=0.745 w=0.42 l=0.15
X246 VSS a_2463_4775# a_2398_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X247 VSS a_8289_4086# x45.D VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X248 x5.A a_1062_5674# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X249 VDD x48.D a_3876_6040# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.0974 ps=0.97 w=0.64 l=0.15
X250 a_11390_4801# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X251 VSS a_5991_2340# x57.Q_N VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X252 a_4590_2732# a_4453_2340# a_4154_2340# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X253 VDD a_8288_2340# D[4] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X254 VSS x7.X a_10155_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X255 a_9953_2732# a_9441_2340# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X256 a_8289_4086# a_8384_4086# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X257 a_2697_5083# a_2289_4801# a_2463_4775# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X258 a_9551_5167# a_8403_4801# a_9465_4801# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X259 a_9441_2340# a_8696_2366# a_9577_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X260 a_6199_4801# x30.D VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X261 a_11630_4086# x5.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X262 VSS x4.X a_6760_4775# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X263 a_5170_4112# a_4658_4086# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.084 ps=0.82 w=0.42 l=0.15
X264 a_10680_2340# a_10775_2340# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X265 VSS sel_bit[1] a_3258_5648# VSS sky130_fd_pr__nfet_01v8 ad=0.0819 pd=0.81 as=0.113 ps=1.38 w=0.42 l=0.15
X266 a_9173_4478# a_8384_4086# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0819 ps=0.81 w=0.42 l=0.15
X267 VDD sel_bit[1] a_3258_5648# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X268 x30.D a_5562_4801# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X269 VDD a_6760_4775# a_7481_5083# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X270 a_4389_4112# a_3600_4086# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0588 ps=0.7 w=0.42 l=0.15
X271 a_5372_4112# a_4454_4086# a_4926_4296# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X272 a_9375_4478# a_9238_4086# a_8939_4086# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X273 VSS a_2061_2340# a_2060_2640# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X274 a_6465_3213# a_6291_3605# a_6605_3239# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X275 VSS a_5897_4086# x48.D VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X276 a_6399_3239# a_6010_3239# a_6291_3605# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X277 VSS a_3599_2340# x54.Q_N VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X278 eob a_2389_5648# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.335 ps=2.67 w=1 l=0.15
X279 VDD x5.X a_1061_4801# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X280 VDD a_5896_2340# D[5] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X281 VDD x27.Q_N a_3599_2340# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.123 ps=1.17 w=0.42 l=0.15
X282 a_11389_3239# a_11543_3213# a_11249_3213# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X283 VDD a_4658_4086# a_4591_4478# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X284 VDD a_9237_2340# a_9236_2640# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X285 a_5897_4086# a_5992_4086# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X286 a_8289_4086# a_8384_4086# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X287 a_6304_2366# x4.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X288 a_3807_4801# x27.D VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X289 a_12146_3239# x39.Q_N VSS VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X290 VSS a_12031_4775# a_12738_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X291 a_6781_4478# a_5992_4086# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0819 ps=0.81 w=0.42 l=0.15
X292 VSS a_1112_2340# D[7] VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X293 a_12146_3239# a_11543_3213# a_12030_3213# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X294 a_6983_4478# a_6846_4086# a_6547_4086# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X295 VDD VDD a_8384_4086# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.123 ps=1.17 w=0.42 l=0.15
X296 a_9238_4086# x5.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X297 a_12047_2648# a_11088_2366# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X298 a_6546_2340# a_6844_2640# a_6780_2732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0924 ps=0.86 w=0.42 l=0.15
X299 a_1520_2366# x4.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.154 ps=1.34 w=0.64 l=0.15
X300 a_4585_3239# a_4073_3213# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X301 VDD a_6466_4775# a_6376_5167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X302 VSS a_7049_2340# a_6984_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0935 ps=0.965 w=0.64 l=0.15
X303 a_11564_2732# a_10775_2340# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0819 ps=0.81 w=0.42 l=0.15
X304 x4.X a_1511_4112# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X305 a_11766_2732# a_11629_2340# a_11330_2340# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X306 a_11833_2340# a_11088_2366# a_11969_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X307 a_4971_4801# a_4368_4775# a_4855_4775# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X308 a_4155_4086# a_4454_4086# a_4389_4112# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.066 ps=0.745 w=0.36 l=0.15
X309 a_10156_4112# a_9237_4386# a_9710_4296# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X310 a_7072_3239# a_6010_3239# a_6977_3239# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X311 a_4007_3239# a_3618_3239# a_3899_3605# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X312 a_8858_4775# a_8684_5167# a_8998_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X313 x4.X a_1511_4112# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X314 VDD x4.X a_11544_4775# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X315 a_6305_4112# x4.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.154 ps=1.34 w=0.64 l=0.15
X316 a_4018_2366# a_4154_2340# a_3599_2340# VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0864 ps=0.91 w=0.64 l=0.15
X317 a_5897_4086# a_5992_4086# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X318 VDD a_12031_4775# a_12738_4801# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X319 a_3912_2366# x4.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X320 a_7158_3605# a_6010_3239# a_7072_3239# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X321 a_12346_4112# a_11834_4086# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.084 ps=0.82 w=0.42 l=0.15
X322 a_9578_4112# a_9710_4296# a_9442_4086# VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0864 ps=0.91 w=0.64 l=0.15
X323 a_12548_4112# a_11630_4086# a_12102_4296# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X324 VDD a_8384_4086# x42.Q_N VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X325 VSS a_9237_2340# a_9236_2640# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X326 a_4925_2550# a_4452_2640# a_5169_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0671 ps=0.75 w=0.36 l=0.15
X327 VDD VDD a_5992_4086# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.123 ps=1.17 w=0.42 l=0.15
X328 x4.A a_897_4112# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X329 VSS a_4657_2340# a_4592_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0935 ps=0.965 w=0.64 l=0.15
X330 x5.A a_1062_5674# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X331 x4.X a_1511_4112# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X332 a_2579_4801# a_1976_4775# a_2463_4775# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X333 VDD x36.Q_N a_10775_2340# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.123 ps=1.17 w=0.42 l=0.15
X334 a_4680_3239# a_3618_3239# a_4585_3239# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X335 a_6466_4775# a_6292_5167# a_6606_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X336 VDD x4.A a_1511_4112# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X337 a_3913_4112# x4.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.154 ps=1.34 w=0.64 l=0.15
X338 a_1626_2366# a_1762_2340# a_1207_2340# VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0864 ps=0.91 w=0.64 l=0.15
X339 VSS a_9638_3213# a_10345_3239# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X340 VDD a_9151_3213# a_9101_3521# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X341 a_1112_2340# a_1207_2340# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X342 a_11390_4801# a_11544_4775# a_11250_4775# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X343 VSS a_6846_4086# a_6845_4386# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X344 a_4766_3605# a_3618_3239# a_4680_3239# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X345 VDD a_11630_4086# a_11629_4386# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X346 x75.Q_N a_4854_3213# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X347 a_2533_2550# a_2060_2640# a_2777_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0671 ps=0.75 w=0.36 l=0.15
X348 a_2401_2366# a_2533_2550# a_2265_2340# VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0864 ps=0.91 w=0.64 l=0.15
X349 a_12147_4801# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X350 VSS x39.D a_12548_4112# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X351 a_12147_4801# a_11544_4775# a_12031_4775# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X352 a_10982_3239# x7.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X353 a_4586_4801# a_4074_4775# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X354 a_2198_2732# a_2061_2340# a_1762_2340# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X355 a_8857_3213# x42.Q_N VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X356 a_8403_4801# a_8237_4801# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X357 a_4008_4801# a_3619_4801# a_3900_5167# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X358 a_7073_4801# a_6011_4801# a_6978_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X359 x66.Q_N a_12030_3213# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X360 VDD a_6759_3213# a_6709_3521# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X361 a_7159_5167# a_6011_4801# a_7073_4801# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X362 a_4454_4086# x5.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X363 VSS a_4454_4086# a_4453_4386# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X364 a_8897_4394# a_8697_4112# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X365 a_12030_3213# x39.Q_N VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X366 D[1] a_10345_3239# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X367 VDD x5.A a_1338_5674# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X368 a_3373_5674# a_2853_5648# a_3648_5972# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.164 ps=1.33 w=0.42 l=0.15
X369 a_11331_4086# a_11629_4386# a_11565_4478# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0924 ps=0.86 w=0.42 l=0.15
X370 a_11856_3239# a_10794_3239# a_11761_3239# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X371 a_8697_4112# x4.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X372 a_8683_3605# a_8402_3239# a_8590_3239# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X373 D[0] a_7953_3239# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X374 a_6011_4801# a_5845_4801# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X375 VSS x36.Q_N a_11969_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.101 ps=0.99 w=0.42 l=0.15
X376 a_4681_4801# a_3619_4801# a_4586_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X377 VDD a_9152_4775# a_9102_5083# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X378 VSS a_3505_4086# x48.Q VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X379 a_4767_5167# a_3619_4801# a_4681_4801# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X380 x4.X a_1511_4112# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X381 VSS VDD a_1976_4775# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X382 a_5170_4478# a_4658_4086# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X383 a_4112_2648# a_3912_2366# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X384 VDD a_3504_2340# D[6] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X385 VSS a_9639_4775# a_10346_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X386 a_2463_4775# x4.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X387 a_3505_4086# a_3600_4086# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X388 a_4389_4478# a_3600_4086# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0819 ps=0.81 w=0.42 l=0.15
X389 VDD x7.X a_7763_2366# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0662 ps=0.735 w=0.42 l=0.15
X390 VSS a_929_3238# x7.X VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X391 VSS a_2389_5648# eob VSS sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X392 VDD a_1976_4775# a_2697_5083# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X393 x4.A a_897_4112# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X394 x27.Q_N a_4855_4775# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X395 a_6411_4112# a_6547_4086# a_5992_4086# VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0864 ps=0.91 w=0.64 l=0.15
X396 VDD x4.A a_1511_4112# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X397 a_8858_4775# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X398 a_10983_4801# x36.D VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X399 VDD a_6760_4775# a_6710_5083# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X400 a_7318_4296# a_6845_4386# a_7562_4112# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0671 ps=0.75 w=0.36 l=0.15
X401 VDD a_9639_4775# a_10346_4801# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X402 a_12031_4775# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X403 a_1720_2648# a_1520_2366# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X404 VSS a_4073_3213# a_4007_3239# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X405 a_3505_4086# a_3600_4086# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X406 VSS a_9638_3213# a_9573_3239# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X407 a_2289_4801# a_1061_4801# a_2147_5083# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X408 a_6845_2340# D[4] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X409 VDD a_2463_4775# a_2375_5167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X410 a_7561_2366# a_7049_2340# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.084 ps=0.82 w=0.42 l=0.15
X411 a_7763_2366# a_6845_2340# a_7317_2550# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X412 x36.D a_10346_4801# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X413 VDD a_1511_4112# x4.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X414 VDD a_9441_2340# a_9374_2732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X415 VSS VDD a_7186_4112# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.101 ps=0.99 w=0.42 l=0.15
X416 a_8684_5167# a_8403_4801# a_8591_4801# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X417 a_11857_4801# a_10795_4801# a_11762_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X418 VDD x7.X a_10155_2366# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0662 ps=0.735 w=0.42 l=0.15
X419 a_8938_2340# a_9237_2340# a_9172_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.066 ps=0.745 w=0.36 l=0.15
X420 a_6930_3521# a_6465_3213# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X421 VDD a_897_4112# x4.A VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X422 a_3600_4086# a_3913_4112# a_4019_4112# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X423 a_1511_4112# x4.A VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X424 VSS VDD a_4019_4112# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.12 ps=1.08 w=0.42 l=0.15
X425 a_12346_4478# a_11834_4086# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X426 a_11288_2648# a_11088_2366# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X427 x75.Q a_5561_3239# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X428 x77.Y eob VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X429 VDD a_9238_4086# a_9237_4386# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X430 a_11493_3521# a_11075_3605# a_11249_3213# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X431 a_3373_5674# sel_bit[1] a_2389_5648# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X432 VDD a_3600_4086# x48.Q_N VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X433 a_9710_4296# a_9237_4386# a_9954_4112# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0671 ps=0.75 w=0.36 l=0.15
X434 a_6845_2340# D[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X435 x4.X a_1511_4112# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X436 a_6546_2340# a_6845_2340# a_6780_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.066 ps=0.745 w=0.36 l=0.15
X437 VSS a_12030_3213# a_11965_3239# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X438 a_11075_3605# a_10628_3239# a_10982_3239# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X439 x69.Q_N a_9638_3213# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X440 a_1415_4801# eob VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X441 VSS a_11249_3213# a_11183_3239# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X442 VDD x5.X a_10629_4801# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X443 x36.Q_N a_12031_4775# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X444 VSS a_929_3238# x7.X VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X445 a_5371_2366# a_4452_2640# a_4925_2550# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X446 VSS a_4074_4775# a_4008_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X447 a_2993_5674# sel_bit[0] a_2883_5674# VSS sky130_fd_pr__nfet_01v8 ad=0.0786 pd=0.805 as=0.072 ps=0.76 w=0.36 l=0.15
X448 VDD x39.D a_12548_4112# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0662 ps=0.735 w=0.42 l=0.15
X449 VSS a_10680_2340# D[3] VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X450 VDD x4.A a_1511_4112# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X451 VSS a_1511_4112# x4.X VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X452 a_12264_3521# a_11856_3239# a_12030_3213# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X453 VSS a_9639_4775# a_9574_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X454 VSS a_2389_5648# eob VSS sky130_fd_pr__nfet_01v8 ad=0.107 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X455 VSS a_1338_5674# x5.X VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X456 a_6931_5083# a_6466_4775# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X457 a_10776_4086# a_11089_4112# a_11195_4112# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X458 VDD x4.X a_11543_3213# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X459 a_3619_4801# a_3453_4801# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X460 VSS VDD a_11195_4112# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.12 ps=1.08 w=0.42 l=0.15
X461 a_2289_4801# a_1227_4801# a_2194_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X462 x33.D a_7954_4801# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X463 a_11494_5083# a_11076_5167# a_11250_4775# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X464 VDD x27.Q_N a_4657_2340# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X465 a_2979_2366# a_2060_2640# a_2533_2550# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X466 a_11159_3605# a_10628_3239# a_11075_3605# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X467 x30.D a_5562_4801# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X468 VDD a_7050_4086# a_6983_4478# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X469 a_9754_3239# x42.Q_N VSS VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X470 a_1508_5167# a_1061_4801# a_1415_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X471 a_9754_3239# a_9151_3213# a_9638_3213# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X472 VSS a_1682_4775# a_1616_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X473 a_9655_2648# a_8696_2366# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X474 VDD a_1511_4112# x4.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X475 a_8384_4086# a_8939_4086# a_8897_4394# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0882 ps=1.05 w=0.84 l=0.15
X476 x7.A a_653_3238# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X477 a_6605_3239# x45.Q_N VSS VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X478 a_7764_4112# a_6845_4386# a_7318_4296# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X479 a_3899_3605# a_3618_3239# a_3806_3239# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X480 a_8938_2340# a_9236_2640# a_9172_2732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0924 ps=0.86 w=0.42 l=0.15
X481 a_12547_2366# a_11628_2640# a_12101_2550# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X482 a_9954_4112# a_9442_4086# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.084 ps=0.82 w=0.42 l=0.15
X483 x20.Q_N a_2463_4775# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X484 a_11076_5167# a_10629_4801# a_10983_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X485 VSS a_12031_4775# a_11966_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X486 VDD a_1511_4112# x4.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X487 VDD x20.Q_N a_2265_2340# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X488 a_1592_5167# a_1061_4801# a_1508_5167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X489 a_8696_2366# x4.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.154 ps=1.34 w=0.64 l=0.15
X490 a_10680_2340# a_10775_2340# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X491 a_5169_2366# a_4657_2340# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.084 ps=0.82 w=0.42 l=0.15
X492 a_3599_2340# a_4154_2340# a_4112_2648# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0882 ps=1.05 w=0.84 l=0.15
X493 a_12265_5083# a_11857_4801# a_12031_4775# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X494 a_10982_3239# x7.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X495 a_7246_3213# a_7072_3239# a_7362_3239# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X496 VDD x3.A a_897_4112# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X497 VDD VDD a_7050_4086# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X498 VDD x7.A a_929_3238# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X499 a_4592_2366# a_4452_2640# a_4154_2340# VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.0711 ps=0.755 w=0.36 l=0.15
X500 a_8402_3239# a_8236_3239# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X501 a_4538_3521# a_4073_3213# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X502 a_4926_4296# a_4454_4086# a_5170_4478# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X503 a_10776_4086# a_11331_4086# a_11289_4394# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0882 ps=1.05 w=0.84 l=0.15
X504 VDD x36.Q_N a_11833_2340# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X505 a_9709_2550# a_9237_2340# a_9953_2732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X506 a_2061_2340# D[6] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X507 VSS x5.X a_1061_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X508 a_2777_2366# a_2265_2340# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.084 ps=0.82 w=0.42 l=0.15
X509 a_1207_2340# a_1762_2340# a_1720_2648# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0882 ps=1.05 w=0.84 l=0.15
X510 a_9755_4801# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X511 a_2979_2366# a_2061_2340# a_2533_2550# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X512 VSS x4.X a_4367_3213# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X513 VSS a_1338_5674# x5.X VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X514 a_9755_4801# a_9152_4775# a_9639_4775# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X515 a_6606_4801# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X516 a_11565_4112# a_10776_4086# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0588 ps=0.7 w=0.42 l=0.15
X517 a_8802_2366# a_8938_2340# a_8383_2340# VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0864 ps=0.91 w=0.64 l=0.15
X518 a_11088_2366# x4.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.154 ps=1.34 w=0.64 l=0.15
X519 VSS x7.X a_5371_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X520 VDD a_4657_2340# a_4590_2732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X521 a_6010_3239# a_5844_3239# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X522 VDD a_4367_3213# a_5088_3521# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X523 a_7264_4394# a_6305_4112# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X524 a_8402_3239# a_8236_3239# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X525 VSS x33.Q_N a_8802_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.12 ps=1.08 w=0.42 l=0.15
X526 a_9638_3213# x42.Q_N VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X527 VDD a_1511_4112# x4.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X528 VSS a_10775_2340# x63.Q_N VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X529 x4.X a_1511_4112# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X530 a_11834_4086# a_12102_4296# a_12048_4394# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X531 a_3648_5972# x48.Q VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.164 pd=1.33 as=0.0864 ps=0.91 w=0.64 l=0.15
X532 a_6400_4801# a_6011_4801# a_6292_5167# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X533 a_10983_4801# x36.D VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X534 a_6846_4086# x5.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X535 a_11768_2366# a_11628_2640# a_11330_2340# VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.0711 ps=0.755 w=0.36 l=0.15
X536 a_2061_2340# D[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X537 a_4539_5083# a_4074_4775# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X538 a_2265_2340# a_2533_2550# a_2479_2648# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X539 a_6605_3239# a_6759_3213# a_6465_3213# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X540 a_7247_4775# a_7073_4801# a_7363_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X541 a_12102_4296# a_11630_4086# a_12346_4478# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X542 a_11761_3239# a_11249_3213# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X543 VSS x33.Q_N a_9577_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.101 ps=0.99 w=0.42 l=0.15
X544 VDD a_9638_3213# a_10345_3239# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X545 VDD a_1511_4112# x4.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X546 a_4872_4394# a_3913_4112# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X547 VSS a_8384_4086# x42.Q_N VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X548 a_11331_4086# a_11630_4086# a_11565_4112# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.066 ps=0.745 w=0.36 l=0.15
X549 VDD a_8383_2340# x60.Q_N VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X550 a_5991_2340# a_6304_2366# a_6410_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X551 a_6010_3239# a_5844_3239# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X552 VDD a_4073_3213# a_3983_3605# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X553 VSS x30.Q_N a_6410_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.12 ps=1.08 w=0.42 l=0.15
X554 a_9464_3239# a_8236_3239# a_9322_3521# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X555 VDD a_9638_3213# a_9550_3605# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X556 VDD a_897_4112# x4.A VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X557 VSS x4.X a_11543_3213# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X558 a_11194_2366# a_11330_2340# a_10775_2340# VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0864 ps=0.91 w=0.64 l=0.15
X559 a_7561_2732# a_7049_2340# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X560 a_9377_4112# a_9237_4386# a_8939_4086# VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.0711 ps=0.755 w=0.36 l=0.15
X561 VSS x4.A a_1511_4112# VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X562 a_7049_2340# a_6304_2366# a_7185_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X563 VSS x4.X a_4368_4775# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X564 a_9238_4086# x5.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X565 a_12101_2550# a_11628_2640# a_12345_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0671 ps=0.75 w=0.36 l=0.15
X566 x5.X a_1338_5674# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X567 eob a_2389_5648# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.175 ps=1.35 w=1 l=0.15
X568 VDD a_11543_3213# a_12264_3521# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X569 x27.D a_3170_4801# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X570 VDD a_4368_4775# a_5089_5083# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X571 VDD a_1511_4112# x4.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X572 a_11969_2366# a_12101_2550# a_11833_2340# VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0864 ps=0.91 w=0.64 l=0.15
X573 VSS a_11833_2340# a_11768_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0935 ps=0.965 w=0.64 l=0.15
X574 a_4073_3213# a_3899_3605# a_4213_3239# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X575 a_9639_4775# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X576 VSS a_7246_3213# a_7953_3239# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X577 VSS a_1207_2340# x51.Q_N VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X578 a_8403_4801# a_8237_4801# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X579 a_6985_4112# a_6845_4386# a_6547_4086# VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.0711 ps=0.755 w=0.36 l=0.15
X580 a_9573_3239# a_8236_3239# a_9464_3239# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X581 a_11942_3605# a_10794_3239# a_11856_3239# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X582 a_4854_3213# a_4680_3239# a_4970_3239# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X583 a_4657_2340# a_3912_2366# a_4793_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X584 x66.Q_N a_12030_3213# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X585 a_1415_4801# eob VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X586 VSS a_9442_4086# a_9377_4112# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0935 ps=0.965 w=0.64 l=0.15
X587 VDD a_12030_3213# a_11942_3605# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X588 a_4591_4478# a_4454_4086# a_4155_4086# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X589 a_4154_2340# a_4452_2640# a_4388_2732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0924 ps=0.86 w=0.42 l=0.15
X590 VDD D[1] a_10628_3239# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X591 a_9954_4478# a_9442_4086# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X592 VDD a_10681_4086# x42.D VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X593 a_8896_2648# a_8696_2366# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X594 VDD a_11249_3213# a_11159_3605# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X595 VDD a_4074_4775# a_3984_5167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X596 a_11762_4801# a_11250_4775# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X597 a_9322_3521# a_8857_3213# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X598 a_9172_2366# a_8383_2340# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0588 ps=0.7 w=0.42 l=0.15
X599 a_9465_4801# a_8237_4801# a_9323_5083# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X600 VSS a_4854_3213# a_5561_3239# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X601 VDD a_9639_4775# a_9551_5167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X602 a_6011_4801# a_5845_4801# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X603 VDD x4.X a_9152_4775# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X604 VSS x45.D a_7764_4112# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X605 D[0] a_7953_3239# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X606 VSS x4.X a_11544_4775# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X607 VSS a_11630_4086# a_11629_4386# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X608 a_1520_2366# x4.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X609 VDD x2.A a_1062_5674# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X610 a_7186_4112# a_7318_4296# a_7050_4086# VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0864 ps=0.91 w=0.64 l=0.15
X611 a_10156_4112# a_9238_4086# a_9710_4296# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X612 VDD a_11544_4775# a_12265_5083# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X613 a_3618_3239# a_3452_3239# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X614 VDD a_5992_4086# x45.Q_N VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X615 a_8683_3605# a_8236_3239# a_8590_3239# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X616 VDD VDD a_3600_4086# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.123 ps=1.17 w=0.42 l=0.15
X617 a_11249_3213# a_11075_3605# a_11389_3239# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X618 x72.Q_N a_7246_3213# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X619 VSS a_8857_3213# a_8791_3239# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X620 VDD a_1682_4775# a_1592_5167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X621 x3.A a_621_4112# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X622 a_6780_2366# a_5991_2340# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0588 ps=0.7 w=0.42 l=0.15
X623 VSS a_2265_2340# a_2200_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0935 ps=0.965 w=0.64 l=0.15
X624 VSS x6.A a_653_3238# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X625 a_4074_4775# a_3900_5167# a_4214_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X626 VSS D[1] a_10628_3239# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X627 VSS x4.A a_1511_4112# VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X628 a_4454_4086# x5.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X629 VSS a_7247_4775# a_7954_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X630 a_6547_4086# a_6845_4386# a_6781_4478# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0924 ps=0.86 w=0.42 l=0.15
X631 a_10681_4086# a_10776_4086# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X632 a_11943_5167# a_10795_4801# a_11857_4801# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X633 a_11088_2366# x4.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X634 a_9872_3521# a_9464_3239# a_9638_3213# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X635 x5.X a_1338_5674# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X636 a_3876_6040# sel_bit[0] a_3373_5674# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0974 pd=0.97 as=0.0567 ps=0.69 w=0.42 l=0.15
X637 a_11565_4478# a_10776_4086# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0819 ps=0.81 w=0.42 l=0.15
X638 VDD a_1511_4112# x4.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X639 a_4794_4112# a_4926_4296# a_4658_4086# VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0864 ps=0.91 w=0.64 l=0.15
X640 a_4855_4775# a_4681_4801# a_4971_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X641 a_9574_4801# a_8237_4801# a_9465_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X642 a_8384_4086# a_8697_4112# a_8803_4112# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X643 a_11767_4478# a_11630_4086# a_11331_4086# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X644 VDD a_12031_4775# a_11943_5167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X645 x36.Q_N a_12031_4775# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X646 D[2] a_12737_3239# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X647 a_9323_5083# a_8858_4775# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X648 VSS x42.D a_10156_4112# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X649 VDD a_5991_2340# x57.Q_N VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X650 a_8767_3605# a_8236_3239# a_8683_3605# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X651 a_3618_3239# a_3452_3239# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X652 a_2194_4801# a_1682_4775# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X653 a_1682_4775# a_1508_5167# a_1822_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X654 VDD a_7247_4775# a_7954_4801# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X655 VSS a_1511_4112# x4.X VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X656 a_5169_2732# a_4657_2340# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X657 a_6465_3213# x45.Q_N VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X658 VSS a_4855_4775# a_5562_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X659 a_10681_4086# a_10776_4086# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X660 a_1616_4801# a_1227_4801# a_1508_5167# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X661 VDD a_4367_3213# a_4317_3521# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X662 VSS a_897_4112# x4.A VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X663 x7.A a_653_3238# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X664 a_6505_4394# a_6305_4112# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X665 a_9709_2550# a_9236_2640# a_9953_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0671 ps=0.75 w=0.36 l=0.15
X666 a_2463_4775# a_2289_4801# a_2579_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X667 x33.D a_7954_4801# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X668 VDD VDD a_10776_4086# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.123 ps=1.17 w=0.42 l=0.15
X669 a_1511_4112# x4.A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X670 VSS a_3600_4086# x48.Q_N VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X671 VDD a_3599_2340# x54.Q_N VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X672 a_1207_2340# a_1520_2366# a_1626_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X673 a_8684_5167# a_8237_4801# a_8591_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X674 VSS a_8858_4775# a_8792_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X675 VDD a_4855_4775# a_5562_4801# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X676 a_6305_4112# x4.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X677 a_3373_5674# sel_bit[0] a_3671_5674# VSS sky130_fd_pr__nfet_01v8 ad=0.072 pd=0.76 as=0.0671 ps=0.75 w=0.36 l=0.15
X678 a_2777_2732# a_2265_2340# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X679 a_6291_3605# a_6010_3239# a_6198_3239# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X680 a_2883_5674# sel_bit[0] a_2784_5996# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.105 ps=0.995 w=0.42 l=0.15
X681 a_9873_5083# a_9465_4801# a_9639_4775# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X682 VSS x5.X a_10629_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X683 a_11629_2340# D[2] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X684 VSS x2.A a_1062_5674# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X685 a_2375_5167# a_1227_4801# a_2289_4801# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X686 VDD a_1112_2340# D[7] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X687 x69.Q_N a_9638_3213# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X688 VDD a_10776_4086# x39.Q_N VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X689 a_11834_4086# a_11089_4112# a_11970_4112# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X690 VDD x7.X a_5371_2366# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0662 ps=0.735 w=0.42 l=0.15
X691 x20.Q_N a_2463_4775# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X692 VDD x5.X a_8237_4801# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X693 x3.A a_621_4112# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X694 VDD x33.Q_N a_9441_2340# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X695 a_8768_5167# a_8237_4801# a_8684_5167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X696 a_6709_3521# a_6291_3605# a_6465_3213# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X697 a_4019_4112# a_4155_4086# a_3600_4086# VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0864 ps=0.91 w=0.64 l=0.15
X698 x7.X a_929_3238# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X699 VSS x4.A a_1511_4112# VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X700 a_7317_2550# a_6845_2340# a_7561_2732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X701 a_6466_4775# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X702 a_3913_4112# x4.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X703 a_3619_4801# a_3453_4801# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X704 VSS a_8288_2340# D[4] VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X705 VDD a_11543_3213# a_11493_3521# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X706 a_4926_4296# a_4453_4386# a_5170_4112# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0671 ps=0.75 w=0.36 l=0.15
X707 VSS a_9238_4086# a_9237_4386# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X708 a_4789_3239# a_3452_3239# a_4680_3239# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X709 VDD a_4368_4775# a_4318_5083# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X710 VSS a_11250_4775# a_11184_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X711 VSS a_4658_4086# a_4593_4112# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0935 ps=0.965 w=0.64 l=0.15
X712 a_11629_2340# D[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X713 VSS a_7246_3213# a_7181_3239# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X714 VDD x5.X a_5845_4801# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X715 x30.Q_N a_7247_4775# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X716 VDD a_7049_2340# a_6982_2732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X717 a_5371_2366# a_4453_2340# a_4925_2550# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X718 a_4388_2366# a_3599_2340# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0588 ps=0.7 w=0.42 l=0.15
X719 VSS a_1511_4112# x4.X VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X720 VSS VDD a_4794_4112# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.101 ps=0.99 w=0.42 l=0.15
X721 a_8383_2340# a_8938_2340# a_8896_2648# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0882 ps=1.05 w=0.84 l=0.15
X722 a_10795_4801# a_10629_4801# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X723 VDD x45.D a_7764_4112# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0662 ps=0.735 w=0.42 l=0.15
X724 a_9442_4086# a_9710_4296# a_9656_4394# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X725 a_6292_5167# a_6011_4801# a_6199_4801# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X726 VSS a_5896_2340# D[5] VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X727 eob a_2389_5648# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.218 ps=1.97 w=0.65 l=0.15
X728 VDD a_1976_4775# a_1926_5083# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X729 a_11160_5167# a_10629_4801# a_11076_5167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X730 a_1511_4112# x4.A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X731 a_8288_2340# a_8383_2340# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X732 VSS a_4854_3213# a_4789_3239# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X733 VSS a_1511_4112# x4.X VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X734 a_1996_2366# a_1207_2340# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0588 ps=0.7 w=0.42 l=0.15
X735 x39.D a_12738_4801# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X736 a_4073_3213# x77.Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X737 a_8997_3239# a_9151_3213# a_8857_3213# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X738 a_3900_5167# a_3619_4801# a_3807_4801# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X739 VDD a_11544_4775# a_11494_5083# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X740 a_4154_2340# a_4453_2340# a_4388_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.066 ps=0.745 w=0.36 l=0.15
X741 VSS x3.A a_897_4112# VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X742 VDD a_6845_2340# a_6844_2640# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X743 VSS x7.A a_929_3238# VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X744 x33.Q_N a_9639_4775# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X745 a_9441_2340# a_9709_2550# a_9655_2648# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X746 VDD a_11834_4086# a_11767_4478# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X747 a_5896_2340# a_5991_2340# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X748 VDD a_9151_3213# a_9872_3521# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X749 a_10775_2340# a_11330_2340# a_11288_2648# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0882 ps=1.05 w=0.84 l=0.15
X750 a_12345_2366# a_11833_2340# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.084 ps=0.82 w=0.42 l=0.15
X751 VDD x42.D a_10156_4112# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0662 ps=0.735 w=0.42 l=0.15
X752 a_9577_2366# a_9709_2550# a_9441_2340# VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0864 ps=0.91 w=0.64 l=0.15
X753 a_12547_2366# a_11629_2340# a_12101_2550# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X754 x7.X a_929_3238# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X755 VSS a_7247_4775# a_7182_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X756 a_9172_2732# a_8383_2340# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0819 ps=0.81 w=0.42 l=0.15
X757 VSS VDD a_11970_4112# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.101 ps=0.99 w=0.42 l=0.15
X758 a_9374_2732# a_9237_2340# a_8938_2340# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X759 VDD x4.X a_9151_3213# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X760 a_1227_4801# a_1061_4801# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X761 x4.X a_1511_4112# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X762 VDD a_4453_2340# a_4452_2640# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X763 a_2389_5648# sel_bit[1] a_2883_5674# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0729 pd=0.81 as=0.14 ps=1.6 w=0.54 l=0.15
X764 VDD a_2389_5648# eob VDD sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X765 x27.D a_3170_4801# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X766 VSS a_6845_2340# a_6844_2640# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X767 a_7362_3239# x45.Q_N VSS VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X768 a_7263_2648# a_6304_2366# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X769 a_7362_3239# a_6759_3213# a_7246_3213# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X770 VSS a_1511_4112# x4.X VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X771 a_5992_4086# a_6547_4086# a_6505_4394# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0882 ps=1.05 w=0.84 l=0.15
X772 VDD a_8857_3213# a_8767_3605# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X773 a_4213_3239# x77.Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X774 VSS a_4855_4775# a_4790_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X775 a_6780_2732# a_5991_2340# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0819 ps=0.81 w=0.42 l=0.15
X776 a_5372_4112# a_4453_4386# a_4926_4296# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X777 VDD x33.Q_N a_8383_2340# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.123 ps=1.17 w=0.42 l=0.15
X778 a_11833_2340# a_12101_2550# a_12047_2648# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X779 a_6982_2732# a_6845_2340# a_6546_2340# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X780 a_4925_2550# a_4453_2340# a_5169_2732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X781 a_11330_2340# a_11629_2340# a_11564_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.066 ps=0.745 w=0.36 l=0.15
X782 VSS x7.X a_12547_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X783 VDD x4.X a_6760_4775# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X784 a_8998_4801# a_9152_4775# a_8858_4775# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X785 a_10155_2366# a_9236_2640# a_9709_2550# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X786 a_7562_4112# a_7050_4086# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.084 ps=0.82 w=0.42 l=0.15
X787 VDD a_9152_4775# a_9873_5083# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X788 VSS a_1511_4112# x4.X VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X789 a_7764_4112# a_6846_4086# a_7318_4296# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X790 VSS a_4453_2340# a_4452_2640# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X791 a_6304_2366# x4.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.154 ps=1.34 w=0.64 l=0.15
X792 a_9369_3239# a_8857_3213# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X793 a_4970_3239# x77.Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X794 a_4871_2648# a_3912_2366# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X795 VSS x5.A a_1338_5674# VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X796 VSS a_897_4112# x4.A VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X797 a_8939_4086# a_9238_4086# a_9173_4112# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.066 ps=0.745 w=0.36 l=0.15
X798 a_8590_3239# x7.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X799 VDD a_7246_3213# a_7953_3239# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X800 VDD x30.Q_N a_5991_2340# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.123 ps=1.17 w=0.42 l=0.15
X801 a_2533_2550# a_2061_2340# a_2777_2732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X802 a_1682_4775# x4.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X803 VDD x5.X a_3453_4801# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X804 VDD VDD a_4658_4086# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X805 a_7050_4086# a_7318_4296# a_7264_4394# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X806 VDD x6.A a_653_3238# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X807 x4.X a_1511_4112# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X808 a_2200_2366# a_2060_2640# a_1762_2340# VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.0711 ps=0.755 w=0.36 l=0.15
X809 a_2853_5648# sel_bit[0] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X810 a_2853_5648# sel_bit[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X811 a_8696_2366# x4.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X812 a_6606_4801# a_6760_4775# a_6466_4775# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X813 VSS a_1511_4112# x4.X VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X814 VSS a_3504_2340# D[6] VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X815 a_11630_4086# x5.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X816 a_3912_2366# x4.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.154 ps=1.34 w=0.64 l=0.15
X817 a_6977_3239# a_6465_3213# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X818 a_6846_4086# x5.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X819 a_11389_3239# x39.Q_N VSS VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X820 VDD a_8858_4775# a_8768_5167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X821 a_7363_4801# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X822 a_8939_4086# a_9237_4386# a_9173_4478# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0924 ps=0.86 w=0.42 l=0.15
X823 a_7363_4801# a_6760_4775# a_7247_4775# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X824 a_6547_4086# a_6846_4086# a_6781_4112# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.066 ps=0.745 w=0.36 l=0.15
X825 a_9464_3239# a_8402_3239# a_9369_3239# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X826 VDD a_4854_3213# a_5561_3239# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X827 a_4214_4801# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X828 x4.X a_1511_4112# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X829 a_4658_4086# a_4926_4296# a_4872_4394# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X830 a_8697_4112# x4.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.154 ps=1.34 w=0.64 l=0.15
X831 VSS x7.X a_2979_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X832 VDD a_2265_2340# a_2198_2732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X833 a_1508_5167# a_1227_4801# a_1415_4801# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X834 a_6410_2366# a_6546_2340# a_5991_2340# VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0864 ps=0.91 w=0.64 l=0.15
X835 VSS a_10681_4086# x42.D VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X836 a_7317_2550# a_6844_2640# a_7561_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0671 ps=0.75 w=0.36 l=0.15
X837 a_3504_2340# a_3599_2340# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X838 a_11183_3239# a_10794_3239# a_11075_3605# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X839 a_7246_3213# x45.Q_N VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
.ends

.subckt hgu_sarlogic_sw_ctrl x35.Q x32.Q x29.Q x26.Q x24.Q x21.Q x5.Q x31.Q x28.Q
+ x25.Q x23.Q x19.Q VDD_SW[7] D[2] D[3] D[4] D[5] D[6] x5.D x20.S x17.S x15.S x13.S
+ x11.S x9.S x7.S x34.Q_N x31.Q_N x28.Q_N x25.Q_N x23.Q_N x19.Q_N VDD_SW_b[7] x35.Q_N
+ x32.Q_N x29.Q_N x26.Q_N x24.Q_N x21.Q_N x5.Q_N D[1] x34.Q x22.A x1.A VSS VDD
X0 a_3420_212# x9.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 VSS VDD a_10509_601# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X2 a_11539_1642# VSS a_11325_1642# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.193 ps=1.34 w=0.42 l=0.15
X3 VSS VDD a_7769_n62# VSS sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.109 ps=1.03 w=0.42 l=0.15
X4 VDD a_15293_601# a_16024_909# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X5 VSS a_5812_212# a_5813_n88# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6 a_5927_n62# a_5812_212# a_5504_106# VSS sky130_fd_pr__nfet_01v8 ad=0.116 pd=1.09 as=0.0486 ps=0.63 w=0.36 l=0.15
X7 a_5323_2457# x30.A VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 VDD x3.X a_939_2457# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_5271_n62# x2.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X10 a_13300_993# a_11987_627# a_13216_993# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0787 pd=0.795 as=0.0567 ps=0.69 w=0.42 l=0.15
X11 VDD VDD a_10509_601# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.17 ps=1.81 w=0.64 l=0.15
X12 VDD x16.X a_11987_627# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X13 a_14887_1642# x9.A1 a_14428_1467# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X14 a_7896_106# a_8205_n88# a_8140_n62# VSS sky130_fd_pr__nfet_01v8 ad=0.0486 pd=0.63 as=0.066 ps=0.745 w=0.36 l=0.15
X15 VSS a_9742_n88# x29.Q_N VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X16 VSS a_14857_1289# a_14791_1315# VSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X17 VDD a_1415_895# a_2136_627# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X18 VDD a_8591_895# a_8516_993# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0956 pd=0.875 as=0.0787 ps=0.795 w=0.42 l=0.15
X19 x7.X a_1757_1642# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.113 ps=1.04 w=0.65 l=0.15
X20 a_1501_122# a_1029_n88# a_1745_304# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X21 a_8933_1642# x9.A1 a_8861_1642# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X22 a_8933_1315# a_8679_1642# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.145 ps=1.11 w=0.42 l=0.15
X23 a_9154_1315# x9.A1 a_8933_1642# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X24 VSS D[6] a_4338_n62# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X25 VDD x17.S a_13461_1642# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.118 ps=1.4 w=0.42 l=0.15
X26 a_10983_895# a_10824_993# a_11123_627# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.109 ps=1.03 w=0.64 l=0.15
X27 VSS x17.S a_13461_1642# VSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.109 ps=1.36 w=0.42 l=0.15
X28 VDD D[2] a_13906_n62# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X29 a_16298_n62# a_15381_n88# a_15853_122# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0675 ps=0.735 w=0.36 l=0.15
X30 a_15518_304# a_15381_n88# a_15072_106# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X31 x19.Q_N a_3807_895# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X32 a_8731_627# a_8117_601# a_8591_895# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X33 a_10041_993# a_9595_627# a_9949_627# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0651 ps=0.73 w=0.42 l=0.15
X34 a_5462_220# a_5271_n62# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X35 VSS x16.X a_11987_627# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X36 x9.A1 a_5323_2457# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X37 a_15608_993# a_14545_627# a_15464_909# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X38 a_9949_627# D[3] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X39 VDD a_76_1467# x6.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X40 VDD a_15293_601# a_15243_909# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X41 a_8545_n62# a_8677_122# a_8409_n88# VSS sky130_fd_pr__nfet_01v8 ad=0.0974 pd=0.97 as=0.0864 ps=0.91 w=0.64 l=0.15
X42 a_11325_1642# x9.A1 a_11253_1642# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X43 VDD a_12134_n88# x32.Q_N VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X44 a_15585_n88# a_15853_122# a_15799_220# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X45 a_11325_1315# a_11071_1642# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.145 ps=1.11 w=0.42 l=0.15
X46 VDD a_13193_n88# a_13126_304# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X47 VDD x30.A a_5323_2457# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X48 a_10532_n62# a_9742_n88# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0703 ps=0.755 w=0.42 l=0.15
X49 a_1028_212# x7.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X50 a_5319_1642# x9.A1 a_4860_1467# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X51 a_10801_n88# a_10055_n62# a_10937_n62# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X52 a_8921_304# a_8409_n88# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X53 VSS a_3420_212# a_3421_n88# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X54 VSS a_5289_1289# a_5223_1315# VSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X55 a_3807_895# x2.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.132 pd=1.22 as=0.0956 ps=0.875 w=0.42 l=0.15
X56 a_15380_212# x20.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X57 VSS a_7823_601# a_7757_627# VSS sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0671 ps=0.75 w=0.42 l=0.15
X58 a_2773_627# D[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X59 a_12433_993# a_12153_627# a_12341_627# VSS sky130_fd_pr__nfet_01v8 ad=0.0675 pd=0.735 as=0.066 ps=0.745 w=0.36 l=0.15
X60 VDD x11.S a_6753_1642# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.0767 ps=0.785 w=0.42 l=0.15
X61 VSS VDD a_8545_n62# VSS sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0974 ps=0.97 w=0.42 l=0.15
X62 a_12134_n88# a_12680_106# a_12638_220# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.132 pd=1.22 as=0.0882 ps=1.05 w=0.84 l=0.15
X63 VSS x11.S a_6760_1315# VSS sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.0693 ps=0.75 w=0.42 l=0.15
X64 VSS a_305_2457# x3.X VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X65 VDD a_12607_601# a_12517_993# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X66 a_6753_1642# VSS a_6539_1642# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.193 ps=1.34 w=0.42 l=0.15
X67 a_7757_627# a_7203_627# a_7649_993# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0675 ps=0.735 w=0.36 l=0.15
X68 x25.Q a_9312_627# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X69 VSS VDD a_8117_601# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X70 VSS x3.X a_939_2457# VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X71 a_2927_1642# x9.A1 a_2468_1467# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X72 a_4862_90# a_4958_n88# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X73 VDD a_13375_895# a_14096_627# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X74 VSS x5.D a_1946_n62# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X75 a_487_n62# x2.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X76 x30.A a_4689_2457# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X77 VDD a_5323_2457# x9.A1 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X78 x9.A1 a_5323_2457# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X79 VSS a_2897_1289# a_2831_1315# VSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X80 VDD x13.S a_8679_1642# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.118 ps=1.4 w=0.42 l=0.15
X81 VDD VDD a_1233_n88# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X82 VDD a_7681_1289# a_7711_1642# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X83 VSS x13.S a_8679_1642# VSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.109 ps=1.36 w=0.42 l=0.15
X84 VDD x20.S a_16323_1642# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.0767 ps=0.785 w=0.42 l=0.15
X85 VSS VDD a_941_601# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X86 VSS x20.S a_16330_1315# VSS sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.0693 ps=0.75 w=0.42 l=0.15
X87 a_6730_n62# a_5813_n88# a_6285_122# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0675 ps=0.735 w=0.36 l=0.15
X88 a_10596_212# x15.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X89 a_5950_304# a_5813_n88# a_5504_106# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X90 a_15143_627# a_15293_601# a_14999_601# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X91 a_3732_993# a_2419_627# a_3648_993# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0787 pd=0.795 as=0.0567 ps=0.69 w=0.42 l=0.15
X92 a_13126_304# a_12989_n88# a_12680_106# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X93 VSS a_939_2457# x2.X VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X94 a_16323_1642# VSS a_16109_1642# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.193 ps=1.34 w=0.42 l=0.15
X95 VDD VDD a_941_601# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.17 ps=1.81 w=0.64 l=0.15
X96 a_3070_220# a_2879_n62# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X97 VDD x1.A a_29_2457# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X98 a_13216_993# a_12153_627# a_13072_909# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X99 a_7557_627# D[4] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X100 VSS a_14428_1467# x18.X VSS sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X101 a_14945_n62# a_15072_106# a_14526_n88# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.03 as=0.0864 ps=0.91 w=0.64 l=0.15
X102 x9.A1 a_5323_2457# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X103 VSS a_8591_895# a_8539_627# VSS sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.066 ps=0.745 w=0.42 l=0.15
X104 VDD a_6199_895# a_6124_993# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0956 pd=0.875 as=0.0787 ps=0.795 w=0.42 l=0.15
X105 VSS a_7350_n88# x26.Q_N VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X106 x34.Q_N a_15767_895# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X107 VSS a_8409_n88# a_8319_n62# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.116 ps=1.09 w=0.64 l=0.15
X108 a_13193_n88# a_13461_122# a_13407_220# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X109 VDD x30.A a_5323_2457# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X110 VSS a_939_2457# x2.X VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X111 a_678_220# a_487_n62# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X112 a_1415_895# x2.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.132 pd=1.22 as=0.0956 ps=0.875 w=0.42 l=0.15
X113 VDD VDD a_8117_601# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.17 ps=1.81 w=0.64 l=0.15
X114 a_9644_1467# VSS a_9786_1642# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X115 a_12937_304# a_12134_n88# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0787 pd=0.795 as=0.0956 ps=0.875 w=0.42 l=0.15
X116 a_4862_90# a_4958_n88# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X117 a_12988_212# x17.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X118 VSS a_10983_895# a_11704_627# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X119 VSS a_5431_601# a_5365_627# VSS sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0671 ps=0.75 w=0.42 l=0.15
X120 a_15495_n62# a_15380_212# a_15072_106# VSS sky130_fd_pr__nfet_01v8 ad=0.116 pd=1.09 as=0.0486 ps=0.63 w=0.36 l=0.15
X121 VSS a_15380_212# a_15381_n88# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X122 VDD D[3] a_11514_n62# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X123 a_10041_993# a_9761_627# a_9949_627# VSS sky130_fd_pr__nfet_01v8 ad=0.0675 pd=0.735 as=0.066 ps=0.745 w=0.36 l=0.15
X124 VSS VDD a_6153_n62# VSS sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0974 ps=0.97 w=0.42 l=0.15
X125 VDD a_9644_1467# x14.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X126 a_9786_1642# x15.S VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X127 VDD a_14857_1289# a_14887_1642# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X128 x2.X a_939_2457# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X129 a_9786_1315# x15.S VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X130 x17.X a_13715_1642# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.158 ps=1.39 w=1 l=0.15
X131 VDD a_10215_601# a_10125_993# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X132 a_7769_n62# a_7896_106# a_7350_n88# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.03 as=0.0864 ps=0.91 w=0.64 l=0.15
X133 a_939_2457# x3.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X134 VDD a_5725_601# a_5675_909# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X135 a_5365_627# a_4811_627# a_5257_993# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0675 ps=0.735 w=0.36 l=0.15
X136 x23.Q a_6920_627# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X137 a_8140_n62# a_7350_n88# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0703 ps=0.755 w=0.42 l=0.15
X138 a_14733_627# D[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X139 VDD a_5323_2457# x9.A1 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X140 a_6153_n62# a_6285_122# a_6017_n88# VSS sky130_fd_pr__nfet_01v8 ad=0.0974 pd=0.97 as=0.0864 ps=0.91 w=0.64 l=0.15
X141 VSS x3.A a_305_2457# VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X142 a_2470_90# a_2566_n88# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X143 a_8409_n88# a_7663_n62# a_8545_n62# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X144 VSS D[2] a_13906_n62# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X145 a_11069_122# a_10597_n88# a_11313_304# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X146 a_76_1467# x9.A1 a_218_1315# VSS sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X147 a_15799_220# a_14839_n62# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X148 x9.A1 a_5323_2457# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X149 VDD a_3333_601# a_4064_909# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X150 a_10931_627# a_9761_627# a_10824_993# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0486 ps=0.63 w=0.36 l=0.15
X151 a_6529_304# a_6017_n88# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X152 VSS a_1028_212# a_1029_n88# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X153 a_7615_1315# VSS a_7252_1467# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X154 a_1340_993# a_27_627# a_1256_993# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0787 pd=0.795 as=0.0567 ps=0.69 w=0.42 l=0.15
X155 VDD a_5323_2457# x9.A1 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X156 a_1978_1315# x9.A1 a_1757_1642# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X157 a_12036_1467# VSS a_12178_1642# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X158 a_5165_627# D[5] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X159 x2.X a_939_2457# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X160 VSS a_939_2457# x2.X VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X161 x19.Q a_4528_627# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X162 VSS a_6199_895# a_6147_627# VSS sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.066 ps=0.745 w=0.42 l=0.15
X163 a_9742_n88# a_10288_106# a_10246_220# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.132 pd=1.22 as=0.0882 ps=1.05 w=0.84 l=0.15
X164 a_15030_220# a_14839_n62# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X165 VSS a_4958_n88# x24.Q_N VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X166 VSS x1.A a_29_2457# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X167 VDD VDD a_14526_n88# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0956 pd=0.875 as=0.132 ps=1.22 w=0.42 l=0.15
X168 VSS a_6017_n88# a_5927_n62# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.116 ps=1.09 w=0.64 l=0.15
X169 a_8335_627# a_7823_601# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.116 pd=1.09 as=0.166 ps=1.8 w=0.64 l=0.15
X170 a_8921_n62# a_8409_n88# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0882 ps=0.84 w=0.42 l=0.15
X171 x9.A1 a_5323_2457# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X172 a_13715_1642# x9.A1 a_13643_1642# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X173 VSS a_2468_1467# x8.X VSS sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X174 a_13715_1315# a_13461_1642# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.145 ps=1.11 w=0.42 l=0.15
X175 a_8848_909# a_8432_993# a_8591_895# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.132 ps=1.22 w=0.84 l=0.15
X176 a_10545_304# a_9742_n88# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0787 pd=0.795 as=0.0956 ps=0.875 w=0.42 l=0.15
X177 a_2470_90# a_2566_n88# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X178 VDD x30.A a_5323_2457# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X179 VSS a_939_2457# x2.X VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X180 VDD a_941_601# a_891_909# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X181 a_581_627# a_27_627# a_473_993# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0675 ps=0.735 w=0.36 l=0.15
X182 a_4338_n62# a_3421_n88# a_3893_122# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0675 ps=0.735 w=0.36 l=0.15
X183 x9.A1 a_5323_2457# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X184 a_5575_627# a_5725_601# a_5431_601# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X185 a_13103_n62# a_12988_212# a_12680_106# VSS sky130_fd_pr__nfet_01v8 ad=0.116 pd=1.09 as=0.0486 ps=0.63 w=0.36 l=0.15
X186 a_3558_304# a_3421_n88# a_3112_106# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X187 VDD a_10596_212# a_10597_n88# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X188 a_15072_106# a_15381_n88# a_15316_n62# VSS sky130_fd_pr__nfet_01v8 ad=0.0486 pd=0.63 as=0.066 ps=0.745 w=0.36 l=0.15
X189 x3.X a_305_2457# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X190 a_3648_993# a_2585_627# a_3504_909# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X191 a_8677_122# a_8204_212# a_8921_n62# VSS sky130_fd_pr__nfet_01v8 ad=0.0675 pd=0.735 as=0.0671 ps=0.75 w=0.36 l=0.15
X192 a_5504_106# a_5812_212# a_5761_304# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0787 ps=0.795 w=0.42 l=0.15
X193 VSS a_12036_1467# x16.X VSS sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X194 a_5377_n62# a_5504_106# a_4958_n88# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.03 as=0.0864 ps=0.91 w=0.64 l=0.15
X195 a_12341_627# D[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X196 a_939_2457# x3.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X197 VDD a_3333_601# a_3283_909# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X198 a_7350_n88# a_7663_n62# a_7769_n62# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X199 a_5675_909# a_5257_993# a_5431_601# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X200 a_7967_627# x2.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0974 pd=0.97 as=0.0882 ps=0.84 w=0.42 l=0.15
X201 VDD a_5323_2457# x9.A1 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X202 VDD a_2897_1289# a_2927_1642# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X203 a_10801_n88# a_11069_122# a_11015_220# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X204 VDD a_5323_2457# x9.A1 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X205 a_9761_627# a_9595_627# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X206 a_13407_220# a_12447_n62# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X207 a_381_627# x5.D VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X208 VSS a_647_601# a_581_627# VSS sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0671 ps=0.75 w=0.42 l=0.15
X209 VSS a_8591_895# a_9312_627# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X210 VDD x15.S a_11539_1642# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.0767 ps=0.785 w=0.42 l=0.15
X211 a_14430_90# a_14526_n88# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X212 a_8204_212# x13.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X213 VDD D[4] a_9122_n62# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X214 VSS x15.S a_11546_1315# VSS sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.0693 ps=0.75 w=0.42 l=0.15
X215 VSS VDD a_14945_n62# VSS sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.109 ps=1.03 w=0.42 l=0.15
X216 VSS a_174_n88# x5.Q_N VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X217 VSS a_3039_601# a_2973_627# VSS sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0671 ps=0.75 w=0.42 l=0.15
X218 x13.X a_8933_1642# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.113 ps=1.04 w=0.65 l=0.15
X219 VSS a_12988_212# a_12989_n88# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X220 VDD a_5323_2457# x9.A1 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X221 VSS a_305_2457# x3.X VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X222 VDD_SW[7] a_2136_627# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X223 x23.Q_N a_6199_895# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X224 VDD VDD a_4958_n88# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0956 pd=0.875 as=0.132 ps=1.22 w=0.42 l=0.15
X225 a_8677_122# a_8205_n88# a_8921_304# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X226 VSS a_939_2457# x2.X VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X227 a_16037_1642# a_15855_1642# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X228 a_14857_1289# x20.S VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X229 x34.Q a_16488_627# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X230 x30.A a_4689_2457# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X231 a_791_627# a_941_601# a_647_601# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X232 x2.X a_939_2457# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X233 a_14857_1289# x20.S VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X234 a_4149_1642# VSS a_4149_1315# VSS sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X235 x20.X a_16109_1642# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.158 ps=1.39 w=1 l=0.15
X236 a_7823_601# x2.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X237 a_9761_627# a_9595_627# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X238 a_6456_909# a_6040_993# a_6199_895# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.132 ps=1.22 w=0.84 l=0.15
X239 VSS D[3] a_11514_n62# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X240 x9.A1 a_5323_2457# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X241 a_8731_627# x2.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.03 as=0.0703 ps=0.755 w=0.42 l=0.15
X242 a_891_909# a_473_993# a_647_601# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X243 a_3183_627# a_3333_601# a_3039_601# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X244 a_10824_993# a_9595_627# a_10727_627# VSS sky130_fd_pr__nfet_01v8 ad=0.0486 pd=0.63 as=0.116 ps=1.09 w=0.36 l=0.15
X245 VSS a_939_2457# x2.X VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X246 a_1166_304# a_1029_n88# a_720_106# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X247 a_10983_895# x2.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.132 pd=1.22 as=0.0956 ps=0.875 w=0.42 l=0.15
X248 a_5431_601# a_5257_993# a_5575_627# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.0974 ps=0.97 w=0.64 l=0.15
X249 a_14430_90# a_14526_n88# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X250 VDD a_9646_90# x29.Q VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X251 a_1256_993# a_193_627# a_1112_909# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X252 a_6285_122# a_5812_212# a_6529_n62# VSS sky130_fd_pr__nfet_01v8 ad=0.0675 pd=0.735 as=0.0671 ps=0.75 w=0.36 l=0.15
X253 VSS a_4862_90# x24.Q VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X254 a_3112_106# a_3420_212# a_3369_304# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0787 ps=0.795 w=0.42 l=0.15
X255 VSS x27.A a_4689_2457# VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X256 a_12465_1289# x17.S VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X257 a_2985_n62# a_3112_106# a_2566_n88# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.03 as=0.0864 ps=0.91 w=0.64 l=0.15
X258 VDD x7.S a_1971_1642# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.0767 ps=0.785 w=0.42 l=0.15
X259 a_7252_1467# x9.A1 a_7394_1315# VSS sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X260 a_12465_1289# x17.S VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X261 a_5896_909# a_5431_601# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X262 a_15907_627# a_15293_601# a_15767_895# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X263 a_1757_1642# VSS a_1757_1315# VSS sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X264 VSS x7.S a_1978_1315# VSS sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.0693 ps=0.75 w=0.42 l=0.15
X265 a_3283_909# a_2865_993# a_3039_601# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X266 a_5575_627# x2.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0974 pd=0.97 as=0.0882 ps=0.84 w=0.42 l=0.15
X267 a_1233_n88# a_1501_122# a_1447_220# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X268 a_939_2457# x3.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X269 a_6529_n62# a_6017_n88# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0882 ps=0.84 w=0.42 l=0.15
X270 a_8153_304# a_7350_n88# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0787 pd=0.795 as=0.0956 ps=0.875 w=0.42 l=0.15
X271 VSS a_939_2457# x2.X VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X272 a_8539_627# a_7369_627# a_8432_993# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0486 ps=0.63 w=0.36 l=0.15
X273 a_12038_90# a_12134_n88# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X274 a_7733_993# a_7369_627# a_7649_993# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X275 a_5812_212# x11.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X276 VSS VDD a_5377_n62# VSS sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.109 ps=1.03 w=0.42 l=0.15
X277 VDD a_12901_601# a_13632_909# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X278 VDD a_8204_212# a_8205_n88# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X279 a_593_n62# a_720_106# a_174_n88# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.03 as=0.0864 ps=0.91 w=0.64 l=0.15
X280 a_2831_1315# VSS a_2468_1467# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X281 VDD x22.A a_4413_2457# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X282 a_3535_n62# a_3420_212# a_3112_106# VSS sky130_fd_pr__nfet_01v8 ad=0.116 pd=1.09 as=0.0486 ps=0.63 w=0.36 l=0.15
X283 x2.X a_939_2457# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X284 a_16097_304# a_15585_n88# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X285 VSS a_14999_601# a_14933_627# VSS sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0671 ps=0.75 w=0.42 l=0.15
X286 a_5504_106# a_5813_n88# a_5748_n62# VSS sky130_fd_pr__nfet_01v8 ad=0.0486 pd=0.63 as=0.066 ps=0.745 w=0.36 l=0.15
X287 x19.Q_N a_3807_895# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X288 a_16330_1315# x9.A1 a_16109_1642# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X289 a_7663_n62# x2.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.17 pd=1.81 as=0.154 ps=1.34 w=0.64 l=0.15
X290 VSS a_15767_895# a_15715_627# VSS sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.066 ps=0.745 w=0.42 l=0.15
X291 VDD a_5323_2457# x9.A1 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X292 a_5323_2457# x30.A VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X293 VDD VDD a_8409_n88# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X294 VSS a_15585_n88# a_15495_n62# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.116 ps=1.09 w=0.64 l=0.15
X295 VSS a_76_1467# x6.X VSS sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X296 a_4958_n88# a_5271_n62# a_5377_n62# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X297 x31.Q a_14096_627# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X298 a_5431_601# x2.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X299 a_4064_909# a_3648_993# a_3807_895# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.132 ps=1.22 w=0.84 l=0.15
X300 a_3839_220# a_2879_n62# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X301 x2.X a_939_2457# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X302 a_4077_1642# a_3895_1642# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X303 a_7369_627# a_7203_627# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X304 a_14428_1467# x9.A1 a_14570_1315# VSS sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X305 a_2897_1289# x9.S VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X306 VDD x14.X a_9595_627# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X307 VDD VDD a_174_n88# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0956 pd=0.875 as=0.132 ps=1.22 w=0.42 l=0.15
X308 VDD a_5323_2457# x9.A1 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X309 x9.A1 a_5323_2457# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X310 a_2897_1289# x9.S VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X311 a_791_627# x2.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0974 pd=0.97 as=0.0882 ps=0.84 w=0.42 l=0.15
X312 a_13906_n62# a_12989_n88# a_13461_122# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0675 ps=0.735 w=0.36 l=0.15
X313 x9.X a_4149_1642# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.158 ps=1.39 w=1 l=0.15
X314 a_10908_993# a_9595_627# a_10824_993# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0787 pd=0.795 as=0.0567 ps=0.69 w=0.42 l=0.15
X315 a_12038_90# a_12134_n88# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X316 VDD a_7254_90# x26.Q VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X317 a_2879_n62# x2.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X318 a_720_106# a_1028_212# a_977_304# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0787 ps=0.795 w=0.42 l=0.15
X319 VSS a_2470_90# x21.Q VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X320 VDD_SW_b[7] a_1415_895# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X321 a_6339_627# a_5725_601# a_6199_895# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X322 a_3504_909# a_3039_601# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X323 VDD VDD a_2566_n88# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0956 pd=0.875 as=0.132 ps=1.22 w=0.42 l=0.15
X324 a_3183_627# x2.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0974 pd=0.97 as=0.0882 ps=0.84 w=0.42 l=0.15
X325 a_15072_106# a_15380_212# a_15329_304# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0787 ps=0.795 w=0.42 l=0.15
X326 VSS D[4] a_9122_n62# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X327 VSS a_939_2457# x2.X VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X328 a_12495_1642# x9.A1 a_12036_1467# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X329 a_1685_1642# a_1503_1642# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X330 VSS a_12465_1289# a_12399_1315# VSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X331 a_6147_627# a_4977_627# a_6040_993# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0486 ps=0.63 w=0.36 l=0.15
X332 a_15243_909# a_14825_993# a_14999_601# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X333 a_218_1642# x7.S VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X334 a_647_601# a_473_993# a_791_627# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.0974 ps=0.97 w=0.64 l=0.15
X335 a_5341_993# a_4977_627# a_5257_993# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X336 a_7369_627# a_7203_627# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X337 a_8432_993# a_7203_627# a_8335_627# VSS sky130_fd_pr__nfet_01v8 ad=0.0486 pd=0.63 as=0.116 ps=1.09 w=0.36 l=0.15
X338 VDD a_10509_601# a_11240_909# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X339 a_218_1315# x7.S VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X340 VSS x14.X a_9595_627# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X341 a_13929_1642# VSS a_13715_1642# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.193 ps=1.34 w=0.42 l=0.15
X342 a_1143_n62# a_1028_212# a_720_106# VSS sky130_fd_pr__nfet_01v8 ad=0.116 pd=1.09 as=0.0486 ps=0.63 w=0.36 l=0.15
X343 a_174_n88# a_487_n62# a_593_n62# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X344 a_6339_627# x2.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.03 as=0.0703 ps=0.755 w=0.42 l=0.15
X345 a_3112_106# a_3421_n88# a_3356_n62# VSS sky130_fd_pr__nfet_01v8 ad=0.0486 pd=0.63 as=0.066 ps=0.745 w=0.36 l=0.15
X346 a_647_601# x2.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X347 a_3039_601# a_2865_993# a_3183_627# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.0974 ps=0.97 w=0.64 l=0.15
X348 VDD a_9742_n88# x29.Q_N VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X349 VSS x22.A a_4413_2457# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X350 a_16298_n62# a_15380_212# a_15853_122# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.0567 ps=0.69 w=0.42 l=0.15
X351 a_5271_n62# x2.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.17 pd=1.81 as=0.154 ps=1.34 w=0.64 l=0.15
X352 VSS a_13193_n88# a_13103_n62# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.116 ps=1.09 w=0.64 l=0.15
X353 VDD VDD a_6017_n88# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X354 VDD x20.S a_15855_1642# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.118 ps=1.4 w=0.42 l=0.15
X355 a_4860_1467# x9.A1 a_5002_1315# VSS sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X356 VSS x20.S a_15855_1642# VSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.109 ps=1.36 w=0.42 l=0.15
X357 a_15511_627# a_14999_601# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.116 pd=1.09 as=0.166 ps=1.8 w=0.64 l=0.15
X358 a_5323_2457# x30.A VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X359 a_15316_n62# a_14526_n88# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0703 ps=0.755 w=0.42 l=0.15
X360 a_2566_n88# a_2879_n62# a_2985_n62# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X361 VSS VDD a_593_n62# VSS sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.109 ps=1.03 w=0.42 l=0.15
X362 x34.Q_N a_15767_895# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X363 VDD a_10983_895# a_11704_627# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X364 a_4370_1315# x9.A1 a_4149_1642# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X365 a_8591_895# a_8432_993# a_8731_627# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.109 ps=1.03 w=0.64 l=0.15
X366 a_3039_601# x2.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X367 x3.X a_305_2457# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X368 VDD a_10801_n88# a_10734_304# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X369 a_1447_220# a_487_n62# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X370 a_16024_909# a_15608_993# a_15767_895# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.132 ps=1.22 w=0.84 l=0.15
X371 a_6539_1642# VSS a_6539_1315# VSS sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X372 VDD x12.X a_7203_627# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X373 VSS VDD a_2985_n62# VSS sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.109 ps=1.03 w=0.42 l=0.15
X374 x2.X a_939_2457# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X375 VDD a_4689_2457# x30.A VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X376 VSS x3.X a_939_2457# VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X377 a_11514_n62# a_10597_n88# a_11069_122# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0675 ps=0.735 w=0.36 l=0.15
X378 a_7649_993# a_7203_627# a_7557_627# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0651 ps=0.73 w=0.42 l=0.15
X379 a_2468_1467# x9.A1 a_2610_1315# VSS sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X380 a_10824_993# a_9761_627# a_10680_909# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X381 VSS a_9644_1467# x14.X VSS sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X382 a_1112_909# a_647_601# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X383 a_14839_n62# x2.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X384 VSS a_13375_895# a_13323_627# VSS sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.066 ps=0.745 w=0.42 l=0.15
X385 x31.Q_N a_13375_895# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X386 x2.X a_939_2457# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X387 x17.X a_13715_1642# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.113 ps=1.04 w=0.65 l=0.15
X388 a_16109_1642# VSS a_16109_1315# VSS sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X389 a_12680_106# a_12988_212# a_12937_304# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0787 ps=0.795 w=0.42 l=0.15
X390 VSS a_14430_90# x35.Q VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X391 a_15853_122# a_15380_212# a_16097_n62# VSS sky130_fd_pr__nfet_01v8 ad=0.0675 pd=0.735 as=0.0671 ps=0.75 w=0.36 l=0.15
X392 VSS VDD a_5725_601# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X393 a_15464_909# a_14999_601# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X394 a_15143_627# x2.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0974 pd=0.97 as=0.0882 ps=0.84 w=0.42 l=0.15
X395 a_6040_993# a_4811_627# a_5943_627# VSS sky130_fd_pr__nfet_01v8 ad=0.0486 pd=0.63 as=0.116 ps=1.09 w=0.36 l=0.15
X396 a_16097_n62# a_15585_n88# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0882 ps=0.84 w=0.42 l=0.15
X397 VSS x12.X a_7203_627# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X398 a_8516_993# a_7203_627# a_8432_993# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0787 pd=0.795 as=0.0567 ps=0.69 w=0.42 l=0.15
X399 VDD VDD a_5725_601# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.17 ps=1.81 w=0.64 l=0.15
X400 a_10596_212# x15.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X401 a_11546_1315# x9.A1 a_11325_1642# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X402 VDD a_5289_1289# a_5319_1642# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X403 a_5323_2457# x30.A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X404 VSS VDD a_3761_n62# VSS sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0974 ps=0.97 w=0.42 l=0.15
X405 VSS a_4689_2457# x30.A VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X406 a_193_627# a_27_627# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X407 a_2973_627# a_2419_627# a_2865_993# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0675 ps=0.735 w=0.36 l=0.15
X408 x19.Q a_4528_627# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X409 a_12553_n62# a_12680_106# a_12134_n88# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.03 as=0.0864 ps=0.91 w=0.64 l=0.15
X410 a_557_993# a_193_627# a_473_993# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X411 a_3947_627# a_3333_601# a_3807_895# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X412 a_14999_601# a_14825_993# a_15143_627# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.0974 ps=0.97 w=0.64 l=0.15
X413 a_14526_n88# a_14839_n62# a_14945_n62# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X414 a_3761_n62# a_3893_122# a_3625_n88# VSS sky130_fd_pr__nfet_01v8 ad=0.0974 pd=0.97 as=0.0864 ps=0.91 w=0.64 l=0.15
X415 a_6199_895# a_6040_993# a_6339_627# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.109 ps=1.03 w=0.64 l=0.15
X416 VDD x9.S a_3895_1642# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.118 ps=1.4 w=0.42 l=0.15
X417 a_14791_1315# VSS a_14428_1467# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X418 a_4149_1642# x9.A1 a_4077_1642# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X419 VSS x9.S a_3895_1642# VSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.109 ps=1.36 w=0.42 l=0.15
X420 a_6467_1642# a_6285_1642# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X421 VDD a_941_601# a_1672_909# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X422 a_7649_993# a_7369_627# a_7557_627# VSS sky130_fd_pr__nfet_01v8 ad=0.0675 pd=0.735 as=0.066 ps=0.745 w=0.36 l=0.15
X423 a_6017_n88# a_5271_n62# a_6153_n62# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X424 a_4149_1315# a_3895_1642# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.145 ps=1.11 w=0.42 l=0.15
X425 a_14999_601# x2.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X426 a_5257_993# a_4811_627# a_5165_627# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0651 ps=0.73 w=0.42 l=0.15
X427 VSS a_78_90# x5.Q VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X428 a_487_n62# x2.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.17 pd=1.81 as=0.154 ps=1.34 w=0.64 l=0.15
X429 VDD a_7823_601# a_7733_993# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X430 x11.X a_6539_1642# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.158 ps=1.39 w=1 l=0.15
X431 a_7252_1467# VSS a_7394_1642# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X432 a_2773_627# D[6] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X433 a_4137_304# a_3625_n88# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X434 a_193_627# a_27_627# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X435 VDD a_8591_895# a_9312_627# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X436 a_6730_n62# a_5812_212# a_6285_122# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.0567 ps=0.69 w=0.42 l=0.15
X437 a_720_106# a_1029_n88# a_964_n62# VSS sky130_fd_pr__nfet_01v8 ad=0.0486 pd=0.63 as=0.066 ps=0.745 w=0.36 l=0.15
X438 VSS a_3807_895# a_3755_627# VSS sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.066 ps=0.745 w=0.42 l=0.15
X439 a_12447_n62# x2.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X440 VDD a_7350_n88# x26.Q_N VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X441 VSS a_2566_n88# x21.Q_N VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X442 x9.A1 a_5323_2457# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X443 VDD VDD a_12134_n88# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0956 pd=0.875 as=0.132 ps=1.22 w=0.42 l=0.15
X444 VSS a_3625_n88# a_3535_n62# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.116 ps=1.09 w=0.64 l=0.15
X445 a_15853_122# a_15381_n88# a_16097_304# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X446 VDD a_8409_n88# a_8342_304# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X447 VDD a_7252_1467# x12.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X448 a_7394_1642# x13.S VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X449 VDD a_12465_1289# a_12495_1642# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X450 a_5943_627# a_5431_601# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.116 pd=1.09 as=0.166 ps=1.8 w=0.64 l=0.15
X451 a_13119_627# a_12607_601# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.116 pd=1.09 as=0.166 ps=1.8 w=0.64 l=0.15
X452 a_1757_1642# x9.A1 a_1685_1642# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X453 a_7394_1315# x13.S VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X454 a_5748_n62# a_4958_n88# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0703 ps=0.755 w=0.42 l=0.15
X455 x2.X a_939_2457# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X456 VSS VDD a_3333_601# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X457 VDD a_15767_895# a_15692_993# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0956 pd=0.875 as=0.0787 ps=0.795 w=0.42 l=0.15
X458 a_13072_909# a_12607_601# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X459 a_1757_1315# a_1503_1642# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.145 ps=1.11 w=0.42 l=0.15
X460 a_15715_627# a_14545_627# a_15608_993# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0486 ps=0.63 w=0.36 l=0.15
X461 a_9122_n62# a_8205_n88# a_8677_122# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0675 ps=0.735 w=0.36 l=0.15
X462 a_6124_993# a_4811_627# a_6040_993# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0787 pd=0.795 as=0.0567 ps=0.69 w=0.42 l=0.15
X463 VSS x3.X a_939_2457# VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X464 VDD VDD a_3333_601# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.17 ps=1.81 w=0.64 l=0.15
X465 a_10711_n62# a_10596_212# a_10288_106# VSS sky130_fd_pr__nfet_01v8 ad=0.116 pd=1.09 as=0.0486 ps=0.63 w=0.36 l=0.15
X466 a_7350_n88# a_7896_106# a_7854_220# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.132 pd=1.22 as=0.0882 ps=1.05 w=0.84 l=0.15
X467 a_1946_n62# a_1029_n88# a_1501_122# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0675 ps=0.735 w=0.36 l=0.15
X468 a_15907_627# x2.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.03 as=0.0703 ps=0.755 w=0.42 l=0.15
X469 VDD a_4860_1467# x10.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X470 a_5002_1642# x11.S VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X471 a_5002_1315# x11.S VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X472 a_5223_1315# VSS a_4860_1467# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X473 a_9147_1642# VSS a_8933_1642# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.193 ps=1.34 w=0.42 l=0.15
X474 VDD_SW[7] a_2136_627# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X475 VSS VDD a_15721_n62# VSS sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0974 ps=0.97 w=0.42 l=0.15
X476 a_10161_n62# a_10288_106# a_9742_n88# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.03 as=0.0864 ps=0.91 w=0.64 l=0.15
X477 x28.Q_N a_10983_895# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X478 a_12638_220# a_12447_n62# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X479 VSS a_12038_90# x32.Q VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X480 VDD a_305_2457# x3.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X481 a_473_993# a_27_627# a_381_627# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0651 ps=0.73 w=0.42 l=0.15
X482 a_3807_895# a_3648_993# a_3947_627# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.109 ps=1.03 w=0.64 l=0.15
X483 a_14933_627# a_14379_627# a_14825_993# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0675 ps=0.735 w=0.36 l=0.15
X484 VDD x3.X a_939_2457# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X485 a_6760_1315# x9.A1 a_6539_1642# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X486 VSS a_6199_895# a_6920_627# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X487 a_15329_304# a_14526_n88# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0787 pd=0.795 as=0.0956 ps=0.875 w=0.42 l=0.15
X488 a_11015_220# a_10055_n62# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X489 x34.Q a_16488_627# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X490 a_15721_n62# a_15853_122# a_15585_n88# VSS sky130_fd_pr__nfet_01v8 ad=0.0974 pd=0.97 as=0.0864 ps=0.91 w=0.64 l=0.15
X491 a_5257_993# a_4977_627# a_5165_627# VSS sky130_fd_pr__nfet_01v8 ad=0.0675 pd=0.735 as=0.066 ps=0.745 w=0.36 l=0.15
X492 VDD D[5] a_6730_n62# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X493 x9.A1 a_5323_2457# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X494 x20.X a_16109_1642# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.113 ps=1.04 w=0.65 l=0.15
X495 VSS VDD a_12553_n62# VSS sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.109 ps=1.03 w=0.42 l=0.15
X496 a_14909_993# a_14545_627# a_14825_993# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X497 a_535_1642# x9.A1 a_76_1467# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X498 VDD a_5431_601# a_5341_993# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X499 a_964_n62# a_174_n88# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0703 ps=0.755 w=0.42 l=0.15
X500 VSS a_505_1289# a_439_1315# VSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X501 VSS a_10596_212# a_10597_n88# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X502 a_12680_106# a_12989_n88# a_12924_n62# VSS sky130_fd_pr__nfet_01v8 ad=0.0486 pd=0.63 as=0.066 ps=0.745 w=0.36 l=0.15
X503 a_4338_n62# a_3420_212# a_3893_122# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.0567 ps=0.69 w=0.42 l=0.15
X504 VDD a_939_2457# x2.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X505 a_10055_n62# x2.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X506 VDD a_4958_n88# x24.Q_N VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X507 VDD VDD a_9742_n88# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0956 pd=0.875 as=0.132 ps=1.22 w=0.42 l=0.15
X508 a_8409_n88# a_8677_122# a_8623_220# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X509 VDD a_6017_n88# a_5950_304# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X510 VSS a_1233_n88# a_1143_n62# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.116 ps=1.09 w=0.64 l=0.15
X511 a_3551_627# a_3039_601# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.116 pd=1.09 as=0.166 ps=1.8 w=0.64 l=0.15
X512 a_14733_627# D[1] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X513 x9.A1 a_5323_2457# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X514 VSS x30.A a_5323_2457# VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X515 a_3356_n62# a_2566_n88# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0703 ps=0.755 w=0.42 l=0.15
X516 VSS a_14526_n88# x35.Q_N VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X517 VDD a_13375_895# a_13300_993# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0956 pd=0.875 as=0.0787 ps=0.795 w=0.42 l=0.15
X518 a_13323_627# a_12153_627# a_13216_993# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0486 ps=0.63 w=0.36 l=0.15
X519 VDD x7.S a_1503_1642# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.118 ps=1.4 w=0.42 l=0.15
X520 a_12399_1315# VSS a_12036_1467# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X521 VSS x7.S a_1503_1642# VSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.109 ps=1.36 w=0.42 l=0.15
X522 a_8204_212# x13.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X523 VSS VDD a_15293_601# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X524 VDD a_939_2457# x2.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X525 a_13515_627# x2.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.03 as=0.0703 ps=0.755 w=0.42 l=0.15
X526 a_13936_1315# x9.A1 a_13715_1642# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X527 VDD VDD a_15293_601# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.17 ps=1.81 w=0.64 l=0.15
X528 a_9949_627# D[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X529 VSS VDD a_13329_n62# VSS sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0974 ps=0.97 w=0.42 l=0.15
X530 a_7681_1289# x13.S VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X531 VSS a_1415_895# a_1363_627# VSS sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.066 ps=0.745 w=0.42 l=0.15
X532 a_10246_220# a_10055_n62# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X533 a_3893_122# a_3420_212# a_4137_n62# VSS sky130_fd_pr__nfet_01v8 ad=0.0675 pd=0.735 as=0.0671 ps=0.75 w=0.36 l=0.15
X534 a_13515_627# a_12901_601# a_13375_895# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X535 a_7681_1289# x13.S VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X536 a_6285_122# a_5813_n88# a_6529_304# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X537 a_15767_895# a_15608_993# a_15907_627# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.109 ps=1.03 w=0.64 l=0.15
X538 x30.A a_4689_2457# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X539 VSS a_5323_2457# x9.A1 VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X540 a_5761_304# a_4958_n88# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0787 pd=0.795 as=0.0956 ps=0.875 w=0.42 l=0.15
X541 x31.Q a_14096_627# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X542 a_12541_627# a_11987_627# a_12433_993# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0675 ps=0.735 w=0.36 l=0.15
X543 VSS a_3807_895# a_4528_627# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X544 VDD a_12901_601# a_12851_909# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X545 VDD x3.A a_305_2457# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X546 a_76_1467# VSS a_218_1642# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X547 a_13329_n62# a_13461_122# a_13193_n88# VSS sky130_fd_pr__nfet_01v8 ad=0.0974 pd=0.97 as=0.0864 ps=0.91 w=0.64 l=0.15
X548 a_15585_n88# a_14839_n62# a_15721_n62# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X549 a_4137_n62# a_3625_n88# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0882 ps=0.84 w=0.42 l=0.15
X550 a_3420_212# x9.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X551 VDD a_174_n88# x5.Q_N VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X552 a_12517_993# a_12153_627# a_12433_993# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X553 a_6539_1642# x9.A1 a_6467_1642# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X554 a_8591_895# x2.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.132 pd=1.22 as=0.0956 ps=0.875 w=0.42 l=0.15
X555 a_6539_1315# a_6285_1642# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.145 ps=1.11 w=0.42 l=0.15
X556 VDD a_5812_212# a_5813_n88# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X557 a_14825_993# a_14379_627# a_14733_627# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0651 ps=0.73 w=0.42 l=0.15
X558 x9.A1 a_5323_2457# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X559 a_13705_304# a_13193_n88# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X560 x25.Q_N a_8591_895# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X561 x9.X a_4149_1642# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.113 ps=1.04 w=0.65 l=0.15
X562 a_10288_106# a_10597_n88# a_10532_n62# VSS sky130_fd_pr__nfet_01v8 ad=0.0486 pd=0.63 as=0.066 ps=0.745 w=0.36 l=0.15
X563 a_6017_n88# a_6285_122# a_6231_220# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X564 a_8623_220# a_7663_n62# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X565 VSS a_12607_601# a_12541_627# VSS sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0671 ps=0.75 w=0.42 l=0.15
X566 a_12341_627# D[2] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X567 VDD a_939_2457# x2.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X568 a_11253_1642# a_11071_1642# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X569 a_16109_1642# x9.A1 a_16037_1642# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X570 a_473_993# a_193_627# a_381_627# VSS sky130_fd_pr__nfet_01v8 ad=0.0675 pd=0.735 as=0.066 ps=0.745 w=0.36 l=0.15
X571 VDD_SW_b[7] a_1415_895# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X572 a_9646_90# a_9742_n88# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X573 x28.Q a_11704_627# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X574 VSS a_12134_n88# x32.Q_N VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X575 a_10073_1289# x15.S VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X576 a_16109_1315# a_15855_1642# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.145 ps=1.11 w=0.42 l=0.15
X577 x9.A1 a_5323_2457# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X578 VSS x30.A a_5323_2457# VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X579 a_10073_1289# x15.S VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X580 x15.X a_11325_1642# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.158 ps=1.39 w=1 l=0.15
X581 VDD a_647_601# a_557_993# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X582 a_1672_909# a_1256_993# a_1415_895# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.132 ps=1.22 w=0.84 l=0.15
X583 a_4977_627# a_4811_627# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X584 a_5812_212# x11.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X585 VSS a_8204_212# a_8205_n88# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X586 a_8319_n62# a_8204_212# a_7896_106# VSS sky130_fd_pr__nfet_01v8 ad=0.116 pd=1.09 as=0.0486 ps=0.63 w=0.36 l=0.15
X587 a_11123_627# x2.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.03 as=0.0703 ps=0.755 w=0.42 l=0.15
X588 VDD a_939_2457# x2.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X589 x2.X a_939_2457# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X590 VDD a_3039_601# a_2949_993# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X591 VDD a_4862_90# x24.Q VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X592 a_7557_627# D[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X593 x9.A1 a_5323_2457# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X594 a_12751_627# a_12901_601# a_12607_601# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X595 a_939_2457# x3.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X596 VSS a_5323_2457# x9.A1 VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X597 a_10734_304# a_10597_n88# a_10288_106# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X598 a_11123_627# a_10509_601# a_10983_895# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X599 VSS D[5] a_6730_n62# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X600 a_3893_122# a_3421_n88# a_4137_304# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X601 a_13375_895# a_13216_993# a_13515_627# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.109 ps=1.03 w=0.64 l=0.15
X602 a_1159_627# a_647_601# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.116 pd=1.09 as=0.166 ps=1.8 w=0.64 l=0.15
X603 VDD a_3807_895# a_3732_993# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0956 pd=0.875 as=0.0787 ps=0.795 w=0.42 l=0.15
X604 VDD a_10509_601# a_10459_909# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X605 a_10937_n62# a_11069_122# a_10801_n88# VSS sky130_fd_pr__nfet_01v8 ad=0.0974 pd=0.97 as=0.0864 ps=0.91 w=0.64 l=0.15
X606 a_3755_627# a_2585_627# a_3648_993# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0486 ps=0.63 w=0.36 l=0.15
X607 a_12851_909# a_12433_993# a_12607_601# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X608 a_13193_n88# a_12447_n62# a_13329_n62# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X609 a_4977_627# a_4811_627# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X610 a_6199_895# x2.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.132 pd=1.22 as=0.0956 ps=0.875 w=0.42 l=0.15
X611 a_10125_993# a_9761_627# a_10041_993# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X612 a_1028_212# x7.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X613 VDD a_3420_212# a_3421_n88# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X614 VSS a_5323_2457# x9.A1 VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X615 a_9646_90# a_9742_n88# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X616 VSS a_15767_895# a_16488_627# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X617 VDD D[1] a_16298_n62# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X618 a_3947_627# x2.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.03 as=0.0703 ps=0.755 w=0.42 l=0.15
X619 a_15380_212# x20.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X620 a_11313_304# a_10801_n88# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X621 x2.X a_939_2457# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X622 a_12036_1467# x9.A1 a_12178_1315# VSS sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X623 a_2879_n62# x2.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.17 pd=1.81 as=0.154 ps=1.34 w=0.64 l=0.15
X624 a_977_304# a_174_n88# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0787 pd=0.795 as=0.0956 ps=0.875 w=0.42 l=0.15
X625 x7.X a_1757_1642# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.158 ps=1.39 w=1 l=0.15
X626 VDD x17.S a_13929_1642# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.0767 ps=0.785 w=0.42 l=0.15
X627 VSS a_10215_601# a_10149_627# VSS sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0671 ps=0.75 w=0.42 l=0.15
X628 VSS VDD a_10937_n62# VSS sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0974 ps=0.97 w=0.42 l=0.15
X629 VDD a_305_2457# x3.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X630 VSS x17.S a_13936_1315# VSS sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.0693 ps=0.75 w=0.42 l=0.15
X631 a_7254_90# a_7350_n88# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X632 a_12924_n62# a_12134_n88# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0703 ps=0.755 w=0.42 l=0.15
X633 x31.Q_N a_13375_895# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X634 VDD a_8117_601# a_8848_909# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X635 VDD VDD a_3625_n88# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X636 VDD a_939_2457# x2.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X637 a_3369_304# a_2566_n88# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0787 pd=0.795 as=0.0956 ps=0.875 w=0.42 l=0.15
X638 a_10149_627# a_9595_627# a_10041_993# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0675 ps=0.735 w=0.36 l=0.15
X639 a_10103_1642# x9.A1 a_9644_1467# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X640 a_2585_627# a_2419_627# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X641 VSS a_1415_895# a_2136_627# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X642 VSS x30.A a_5323_2457# VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X643 VSS a_10073_1289# a_10007_1315# VSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X644 VDD x10.X a_4811_627# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X645 a_2949_993# a_2585_627# a_2865_993# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X646 a_14825_993# a_14545_627# a_14733_627# VSS sky130_fd_pr__nfet_01v8 ad=0.0675 pd=0.735 as=0.066 ps=0.745 w=0.36 l=0.15
X647 a_505_1289# x7.S VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X648 a_505_1289# x7.S VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X649 a_13632_909# a_13216_993# a_13375_895# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.132 ps=1.22 w=0.84 l=0.15
X650 x9.A1 a_5323_2457# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X651 x3.X a_305_2457# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X652 VDD a_2470_90# x21.Q VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X653 a_5165_627# D[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X654 VDD a_14999_601# a_14909_993# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X655 a_14526_n88# a_15072_106# a_15030_220# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.132 pd=1.22 as=0.0882 ps=1.05 w=0.84 l=0.15
X656 x3.A a_29_2457# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X657 VDD a_939_2457# x2.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X658 a_939_2457# x3.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X659 a_13906_n62# a_12988_212# a_13461_122# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.0567 ps=0.69 w=0.42 l=0.15
X660 VDD x27.A a_4689_2457# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X661 VSS a_5323_2457# x9.A1 VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X662 a_10288_106# a_10596_212# a_10545_304# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0787 ps=0.795 w=0.42 l=0.15
X663 VSS a_10983_895# a_10931_627# VSS sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.066 ps=0.745 w=0.42 l=0.15
X664 a_13461_122# a_12988_212# a_13705_n62# VSS sky130_fd_pr__nfet_01v8 ad=0.0675 pd=0.735 as=0.0671 ps=0.75 w=0.36 l=0.15
X665 VSS a_5323_2457# x9.A1 VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X666 VDD a_1415_895# a_1340_993# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0956 pd=0.875 as=0.0787 ps=0.795 w=0.42 l=0.15
X667 a_1363_627# a_193_627# a_1256_993# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0486 ps=0.63 w=0.36 l=0.15
X668 a_2585_627# a_2419_627# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X669 a_12751_627# x2.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0974 pd=0.97 as=0.0882 ps=0.84 w=0.42 l=0.15
X670 a_3648_993# a_2419_627# a_3551_627# VSS sky130_fd_pr__nfet_01v8 ad=0.0486 pd=0.63 as=0.116 ps=1.09 w=0.36 l=0.15
X671 a_13705_n62# a_13193_n88# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0882 ps=0.84 w=0.42 l=0.15
X672 VDD a_939_2457# x2.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X673 VSS x10.X a_4811_627# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X674 a_7254_90# a_7350_n88# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X675 VSS a_5323_2457# x9.A1 VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X676 a_1555_627# x2.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.03 as=0.0703 ps=0.755 w=0.42 l=0.15
X677 a_12988_212# x17.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X678 a_8342_304# a_8205_n88# a_7896_106# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X679 a_8432_993# a_7369_627# a_8288_909# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X680 VDD a_15380_212# a_15381_n88# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X681 x11.X a_6539_1642# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.113 ps=1.04 w=0.65 l=0.15
X682 a_8933_1642# VSS a_8933_1315# VSS sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X683 a_439_1315# VSS a_76_1467# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X684 VDD a_8117_601# a_8067_909# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X685 VDD x13.S a_9147_1642# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.0767 ps=0.785 w=0.42 l=0.15
X686 x25.Q a_9312_627# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X687 VSS VDD a_1369_n62# VSS sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0974 ps=0.97 w=0.42 l=0.15
X688 a_10359_627# a_10509_601# a_10215_601# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X689 x30.A a_4689_2457# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X690 VSS x13.S a_9154_1315# VSS sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.0693 ps=0.75 w=0.42 l=0.15
X691 a_1555_627# a_941_601# a_1415_895# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X692 a_12607_601# a_12433_993# a_12751_627# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.0974 ps=0.97 w=0.64 l=0.15
X693 a_5323_2457# x30.A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X694 x2.X a_939_2457# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X695 a_13643_1642# a_13461_1642# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X696 a_14839_n62# x2.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.17 pd=1.81 as=0.154 ps=1.34 w=0.64 l=0.15
X697 VSS a_7252_1467# x12.X VSS sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X698 VDD VDD a_15585_n88# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X699 a_381_627# x5.D VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X700 a_1369_n62# a_1501_122# a_1233_n88# VSS sky130_fd_pr__nfet_01v8 ad=0.0974 pd=0.97 as=0.0864 ps=0.91 w=0.64 l=0.15
X701 a_12134_n88# a_12447_n62# a_12553_n62# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X702 a_10007_1315# VSS a_9644_1467# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X703 VDD x8.X a_2419_627# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X704 a_10459_909# a_10041_993# a_10215_601# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X705 a_3625_n88# a_2879_n62# a_3761_n62# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X706 a_14428_1467# VSS a_14570_1642# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X707 a_12607_601# x2.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X708 a_2865_993# a_2419_627# a_2773_627# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0651 ps=0.73 w=0.42 l=0.15
X709 VDD a_1028_212# a_1029_n88# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X710 VSS a_13375_895# a_14096_627# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X711 a_14545_627# a_14379_627# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X712 a_11240_909# a_10824_993# a_10983_895# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.132 ps=1.22 w=0.84 l=0.15
X713 VDD a_14428_1467# x18.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X714 a_14570_1642# x20.S VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X715 a_1745_304# a_1233_n88# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X716 x9.A1 a_5323_2457# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X717 a_14570_1315# x20.S VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X718 VDD a_6199_895# a_6920_627# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X719 a_11514_n62# a_10596_212# a_11069_122# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.0567 ps=0.69 w=0.42 l=0.15
X720 VSS a_4860_1467# x10.X VSS sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X721 VDD a_14430_90# x35.Q VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X722 a_939_2457# x3.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X723 a_13461_122# a_12989_n88# a_13705_304# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X724 x3.A a_29_2457# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X725 a_11325_1642# VSS a_11325_1315# VSS sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X726 a_10727_627# a_10215_601# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.116 pd=1.09 as=0.166 ps=1.8 w=0.64 l=0.15
X727 a_10680_909# a_10215_601# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X728 x28.Q_N a_10983_895# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X729 VDD a_939_2457# x2.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X730 VDD a_5725_601# a_6456_909# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X731 VSS D[1] a_16298_n62# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X732 a_11313_n62# a_10801_n88# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0882 ps=0.84 w=0.42 l=0.15
X733 VSS x8.X a_2419_627# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X734 x2.X a_939_2457# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X735 a_15608_993# a_14379_627# a_15511_627# VSS sky130_fd_pr__nfet_01v8 ad=0.0486 pd=0.63 as=0.116 ps=1.09 w=0.36 l=0.15
X736 a_14545_627# a_14379_627# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X737 a_6040_993# a_4977_627# a_5896_909# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X738 VSS a_5323_2457# x9.A1 VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X739 a_4958_n88# a_5504_106# a_5462_220# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.132 pd=1.22 as=0.0882 ps=1.05 w=0.84 l=0.15
X740 x23.Q a_6920_627# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X741 a_10215_601# a_10041_993# a_10359_627# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.0974 ps=0.97 w=0.64 l=0.15
X742 a_4860_1467# VSS a_5002_1642# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X743 a_1415_895# a_1256_993# a_1555_627# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.109 ps=1.03 w=0.64 l=0.15
X744 a_11069_122# a_10596_212# a_11313_n62# VSS sky130_fd_pr__nfet_01v8 ad=0.0675 pd=0.735 as=0.0671 ps=0.75 w=0.36 l=0.15
X745 a_8861_1642# a_8679_1642# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X746 VDD x15.S a_11071_1642# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.118 ps=1.4 w=0.42 l=0.15
X747 a_5323_2457# x30.A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X748 x2.X a_939_2457# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X749 a_9742_n88# a_10055_n62# a_10161_n62# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X750 VDD a_10073_1289# a_10103_1642# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X751 VSS x15.S a_11071_1642# VSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.109 ps=1.36 w=0.42 l=0.15
X752 a_1233_n88# a_487_n62# a_1369_n62# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X753 a_10359_627# x2.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0974 pd=0.97 as=0.0882 ps=0.84 w=0.42 l=0.15
X754 x3.X a_305_2457# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X755 a_1256_993# a_27_627# a_1159_627# VSS sky130_fd_pr__nfet_01v8 ad=0.0486 pd=0.63 as=0.116 ps=1.09 w=0.36 l=0.15
X756 a_10215_601# x2.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X757 VSS a_5323_2457# x9.A1 VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X758 VDD a_78_90# x5.Q VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X759 x27.A a_4413_2457# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X760 a_15767_895# x2.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.132 pd=1.22 as=0.0956 ps=0.875 w=0.42 l=0.15
X761 a_12153_627# a_11987_627# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X762 a_7967_627# a_8117_601# a_7823_601# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X763 VDD D[6] a_4338_n62# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X764 VDD x18.X a_14379_627# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X765 VDD x3.X a_939_2457# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X766 VSS VDD a_10161_n62# VSS sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.109 ps=1.03 w=0.42 l=0.15
X767 a_78_90# a_174_n88# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X768 a_2468_1467# VSS a_2610_1642# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X769 VDD a_12988_212# a_12989_n88# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X770 VSS a_9646_90# x29.Q VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X771 a_7896_106# a_8204_212# a_8153_304# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0787 ps=0.795 w=0.42 l=0.15
X772 VDD a_3807_895# a_4528_627# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X773 VDD a_2566_n88# x21.Q_N VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X774 VDD a_3625_n88# a_3558_304# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X775 VDD a_2468_1467# x8.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X776 a_2610_1642# x9.S VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X777 a_8067_909# a_7649_993# a_7823_601# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X778 x2.X a_939_2457# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X779 a_2610_1315# x9.S VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X780 VDD a_10983_895# a_10908_993# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0956 pd=0.875 as=0.0787 ps=0.795 w=0.42 l=0.15
X781 a_12447_n62# x2.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.17 pd=1.81 as=0.154 ps=1.34 w=0.64 l=0.15
X782 VDD VDD a_13193_n88# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X783 a_174_n88# a_720_106# a_678_220# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.132 pd=1.22 as=0.0882 ps=1.05 w=0.84 l=0.15
X784 VSS VDD a_12901_601# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X785 a_2865_993# a_2585_627# a_2773_627# VSS sky130_fd_pr__nfet_01v8 ad=0.0675 pd=0.735 as=0.066 ps=0.745 w=0.36 l=0.15
X786 a_12153_627# a_11987_627# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X787 a_7663_n62# x2.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X788 a_9122_n62# a_8204_212# a_8677_122# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.0567 ps=0.69 w=0.42 l=0.15
X789 a_15692_993# a_14379_627# a_15608_993# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0787 pd=0.795 as=0.0567 ps=0.69 w=0.42 l=0.15
X790 VSS x18.X a_14379_627# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X791 VDD x9.S a_4363_1642# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.0767 ps=0.785 w=0.42 l=0.15
X792 VDD VDD a_12901_601# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.17 ps=1.81 w=0.64 l=0.15
X793 VDD a_12036_1467# x16.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X794 a_12178_1642# x17.S VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X795 a_9644_1467# x9.A1 a_9786_1315# VSS sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X796 VSS x9.S a_4370_1315# VSS sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.0693 ps=0.75 w=0.42 l=0.15
X797 a_12178_1315# x17.S VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X798 a_2566_n88# a_3112_106# a_3070_220# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.132 pd=1.22 as=0.0882 ps=1.05 w=0.84 l=0.15
X799 x25.Q_N a_8591_895# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X800 VDD a_4689_2457# x30.A VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X801 VDD VDD a_7350_n88# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0956 pd=0.875 as=0.132 ps=1.22 w=0.42 l=0.15
X802 a_1946_n62# a_1028_212# a_1501_122# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.0567 ps=0.69 w=0.42 l=0.15
X803 a_4363_1642# VSS a_4149_1642# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.193 ps=1.34 w=0.42 l=0.15
X804 VDD a_12038_90# x32.Q VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X805 a_1501_122# a_1028_212# a_1745_n62# VSS sky130_fd_pr__nfet_01v8 ad=0.0675 pd=0.735 as=0.0671 ps=0.75 w=0.36 l=0.15
X806 a_78_90# a_174_n88# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X807 VDD x6.X a_27_627# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X808 x28.Q a_11704_627# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X809 x2.X a_939_2457# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X810 a_7711_1642# x9.A1 a_7252_1467# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X811 a_1745_n62# a_1233_n88# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0882 ps=0.84 w=0.42 l=0.15
X812 VSS a_4689_2457# x30.A VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X813 x15.X a_11325_1642# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.113 ps=1.04 w=0.65 l=0.15
X814 VSS a_7681_1289# a_7615_1315# VSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X815 a_13375_895# x2.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.132 pd=1.22 as=0.0956 ps=0.875 w=0.42 l=0.15
X816 VDD x5.D a_1946_n62# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X817 VDD a_505_1289# a_535_1642# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X818 x13.X a_8933_1642# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.158 ps=1.39 w=1 l=0.15
X819 a_13216_993# a_11987_627# a_13119_627# VSS sky130_fd_pr__nfet_01v8 ad=0.0486 pd=0.63 as=0.116 ps=1.09 w=0.36 l=0.15
X820 a_7823_601# a_7649_993# a_7967_627# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.0974 ps=0.97 w=0.64 l=0.15
X821 x27.A a_4413_2457# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X822 a_1971_1642# VSS a_1757_1642# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.193 ps=1.34 w=0.42 l=0.15
X823 x23.Q_N a_6199_895# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X824 VSS a_7254_90# x26.Q VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X825 a_12433_993# a_11987_627# a_12341_627# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0651 ps=0.73 w=0.42 l=0.15
X826 a_7854_220# a_7663_n62# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X827 VDD x11.S a_6285_1642# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.118 ps=1.4 w=0.42 l=0.15
X828 a_3625_n88# a_3893_122# a_3839_220# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X829 VSS x11.S a_6285_1642# VSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.109 ps=1.36 w=0.42 l=0.15
X830 VDD a_1233_n88# a_1166_304# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X831 a_8288_909# a_7823_601# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X832 a_13715_1642# VSS a_13715_1315# VSS sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X833 VDD a_14526_n88# x35.Q_N VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X834 VDD a_15767_895# a_16488_627# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X835 a_10055_n62# x2.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.17 pd=1.81 as=0.154 ps=1.34 w=0.64 l=0.15
X836 VSS x6.X a_27_627# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X837 VSS a_10801_n88# a_10711_n62# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.116 ps=1.09 w=0.64 l=0.15
X838 VDD a_15585_n88# a_15518_304# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X839 VDD VDD a_10801_n88# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X840 a_6231_220# a_5271_n62# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X841 a_5289_1289# x11.S VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X842 x2.X a_939_2457# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X843 a_5289_1289# x11.S VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
.ends

.subckt hgu_sarlogic_retimer eob x2.code[2] x2.code[1] x2.x10.A x1[1].D x1[2].D x1[5].D
+ x1[4].D x1[1].Q x1[0].Q x1[3].Q x1[2].Q x1[5].Q x1[4].Q x1[7].Q x1[6].Q x1[6].D
+ x1[7].D x1[3].D x1[0].D x2.x7.SW x2.x2.SW VSS VDD
X0 a_14018_6401# a_13844_6793# a_14158_6427# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X1 x1[3].Q a_17898_6427# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X2 a_16654_5787# a_16236_5787# a_16410_5761# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X3 a_16410_7041# a_16236_7067# a_16550_7433# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X4 VSS a_17191_5121# a_17126_5147# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X5 a_13751_5147# x1[6].D VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X6 a_16922_6109# a_16410_5761# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X7 VSS a_16410_5121# a_16344_5147# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X8 VSS eob a_12385_8002# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X9 a_14530_7389# a_14018_7041# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X10 x1[2].Q a_15506_6427# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X11 a_14483_5787# a_14018_5761# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X12 a_16410_5761# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X13 a_18195_9356# x2.x9.output_stack VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X14 x3.X a_18499_9105# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X15 VDD a_16704_7267# a_16654_7067# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X16 VDD a_17191_7041# a_17898_7083# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X17 x2.x3[1].floating x2.code[1] x2.x9.output_stack VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X18 VSS x3.X a_13397_7073# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X19 x1[0].Q_N a_14799_7041# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X20 VDD VDD a_14312_6401# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X21 a_16236_5787# a_15955_5793# a_16143_5787# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X22 VDD x3.X a_13397_5147# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X23 a_14262_7067# a_13844_7067# a_14018_7041# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X24 a_16143_6427# x1[3].D VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X25 a_14734_7445# a_13397_7073# a_14625_7445# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X26 a_14915_6153# a_14312_5987# a_14799_5761# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X27 a_13928_5513# a_13397_5147# a_13844_5513# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X28 VSS a_14018_7041# a_13952_7445# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X29 a_16236_7067# a_15789_7073# a_16143_7067# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X30 VSS a_14799_5761# a_14734_6165# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X31 a_13844_5787# a_13563_5793# a_13751_5787# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X32 VDD VDD a_16704_7267# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X33 VDD a_17191_5761# a_17898_5803# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X34 a_14018_7041# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X35 a_13751_6427# x1[2].D VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X36 a_16654_6709# a_16236_6793# a_16410_6401# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X37 VDD a_17191_6401# a_17103_6793# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X38 VSS x3.X a_13397_5147# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X39 a_14018_7041# a_13844_7067# a_14158_7433# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X40 a_15033_7067# a_14625_7445# a_14799_7041# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X41 VDD a_16410_6401# a_16320_6793# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X42 VDD x3.X a_15789_5793# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X43 a_16410_5761# a_16236_5787# a_16550_6153# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X44 a_16875_5429# a_16410_5121# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X45 a_13844_7067# a_13397_7073# a_13751_7067# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X46 VSS VDD a_16704_7267# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X47 x1[1].Q a_17898_7083# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X48 a_14483_6709# a_14018_6401# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X49 a_17103_5787# a_15955_5793# a_17017_6165# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X50 VDD a_16704_7267# a_17425_7067# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X51 a_14530_6109# a_14018_5761# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X52 a_17307_6153# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X53 VSS a_14018_5121# a_13952_5147# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X54 a_16550_6427# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X55 VDD a_14799_7041# a_15506_7083# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X56 a_15955_7073# a_15789_7073# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X57 a_16922_5147# a_16410_5121# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X58 VDD a_14312_5121# a_14262_5429# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X59 x1[0].Q a_15506_7083# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X60 a_17191_6401# a_17017_6427# a_17307_6427# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X61 a_14711_5787# a_13563_5793# a_14625_6165# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X62 x2.x9.output_stack x2.x10.Y x2.x5[7].floating VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X63 a_12385_8278# eob a_12297_8278# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X64 a_14915_6153# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X65 VSS VDD a_16704_5121# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X66 VDD VDD a_14312_5121# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X67 VSS VDD a_14312_6401# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X68 VSS a_17191_6401# a_17898_6427# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X69 a_16143_5147# x1[7].D VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X70 a_17017_6165# a_15789_5793# a_16875_5787# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X71 a_18195_9015# x2.x9.output_stack VSS VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X72 a_16320_6793# a_15789_6427# a_16236_6793# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X73 VDD a_14799_5761# a_15506_5803# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X74 x1[7].Q_N a_17191_5121# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X75 VDD a_17191_5121# a_17103_5513# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X76 a_14915_5147# a_14312_5121# a_14799_5121# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X77 a_13751_5147# x1[6].D VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X78 a_17191_7041# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X79 VDD a_14018_6401# a_13928_6793# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X80 x1[2].Q_N a_14799_6401# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X81 VDD x3.X a_13397_5793# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X82 a_14018_5761# a_13844_5787# a_14158_6153# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X83 VDD a_16410_5121# a_16320_5513# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X84 a_16550_6427# a_16704_6401# a_16410_6401# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X85 x2.x10.Y x2.x10.A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X86 a_14158_6427# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X87 a_16410_5121# a_16236_5513# a_16550_5147# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X88 VDD a_14312_5121# a_15033_5429# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X89 a_17017_7445# a_15955_7073# a_16922_7389# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X90 a_16344_5147# a_15955_5147# a_16236_5513# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X91 a_18195_9356# x2.x9.output_stack x3.A VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.122 ps=1.42 w=0.42 l=0.15
X92 a_14625_7445# a_13397_7073# a_14483_7067# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X93 VDD a_14799_7041# a_14711_7067# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X94 a_14530_5147# a_14018_5121# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X95 a_12385_8692# eob a_12297_8554# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X96 a_15955_7073# a_15789_7073# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X97 a_17191_7041# a_17017_7445# a_17307_7433# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X98 a_14799_6401# a_14625_6427# a_14915_6427# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X99 x1[6].Q_N a_14799_5121# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X100 a_13952_5147# a_13563_5147# a_13844_5513# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X101 x1[1].Q_N a_17191_7041# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X102 VSS a_14799_6401# a_15506_6427# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X103 a_14799_5761# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X104 x1[3].Q a_17898_6427# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X105 VSS x3.X a_15789_5793# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X106 a_16143_5787# x1[5].D VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X107 a_15955_5147# a_15789_5147# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X108 a_17425_5787# a_17017_6165# a_17191_5761# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X109 x2.x9.output_stack x2.x10.Y x2.x5[7].floating VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X110 x2.x9.output_stack x2.code[2] x2.x4[3].floating VSS sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X111 a_14625_5147# a_13563_5147# a_14530_5147# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X112 a_12385_8968# eob a_12297_8830# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X113 a_12457_8140# eob a_12385_8278# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X114 a_17126_7445# a_15789_7073# a_17017_7445# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X115 a_13563_6427# a_13397_6427# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X116 a_13751_5787# x1[4].D VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X117 VSS a_17191_5761# a_17126_6165# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X118 a_16320_5513# a_15789_5147# a_16236_5513# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X119 x2.x9.output_stack x2.x7.SW x2.x7.floating VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X120 a_18195_9015# x3.A VDD VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X121 x1[2].Q a_15506_6427# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X122 VDD a_14018_5121# a_13928_5513# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X123 a_16410_6401# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X124 VSS a_16410_5761# a_16344_6165# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X125 a_15955_5147# a_15789_5147# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X126 x3.X a_18499_9105# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X127 a_16550_7433# a_16704_7267# a_16410_7041# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X128 VDD a_16704_5987# a_16654_5787# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X129 x2.x9.output_stack x2.x10.Y x2.x5[7].floating VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X130 a_13563_6427# a_13397_6427# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X131 x1[4].Q_N a_14799_5761# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X132 x1[7].Q a_17898_5147# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X133 a_14018_5121# a_13844_5513# a_14158_5147# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X134 a_16236_6793# a_15955_6427# a_16143_6427# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X135 a_16875_7067# a_16410_7041# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X136 a_14262_5787# a_13844_5787# a_14018_5761# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X137 a_13928_7067# a_13397_7073# a_13844_7067# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X138 x1[6].Q a_15506_5147# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X139 a_17191_5761# a_17017_6165# a_17307_6153# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X140 VDD x2.x7.SW x2.x6.SW VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X141 a_14799_7041# a_14625_7445# a_14915_7433# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X142 VDD eob a_12322_10357# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X143 a_13844_6793# a_13563_6427# a_13751_6427# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X144 a_17425_6709# a_17017_6427# a_17191_6401# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X145 VDD VDD a_16704_5987# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X146 x1[5].Q_N a_17191_5761# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X147 VDD a_14312_7267# a_14262_7067# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X148 VSS x3.X a_13397_5793# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X149 a_14018_5761# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X150 x2.x9.output_stack x2.code[1] x2.x3[1].floating VSS sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X151 a_14734_6427# a_13397_6427# a_14625_6427# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X152 a_15033_5787# a_14625_6165# a_14799_5761# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X153 a_12457_8692# eob a_12385_8692# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X154 a_16236_6793# a_15789_6427# a_16143_6427# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X155 x1[5].Q a_17898_5803# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X156 a_12410_9943# eob a_12322_9805# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X157 VDD a_16704_6401# a_16654_6709# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X158 a_17103_6793# a_15955_6427# a_17017_6427# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X159 a_14734_6165# a_13397_5793# a_14625_6165# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X160 VDD a_16704_5987# a_17425_5787# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X161 a_16550_7433# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X162 VSS a_14799_6401# a_14734_6427# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X163 VSS a_14018_5761# a_13952_6165# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X164 a_16236_5787# a_15789_5793# a_16143_5787# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X165 a_16410_5121# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X166 a_13844_6793# a_13397_6427# a_13751_6427# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X167 VDD a_17191_6401# a_17898_6427# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X168 a_15955_5793# a_15789_5793# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X169 a_16550_6153# a_16704_5987# a_16410_5761# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X170 a_16654_5429# a_16236_5513# a_16410_5121# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X171 x2.x9.output_stack eob a_12385_8968# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X172 a_14711_6793# a_13563_6427# a_14625_6427# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X173 x1[4].Q a_15506_5803# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X174 VDD VDD a_14312_7267# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X175 a_13844_5787# a_13397_5793# a_13751_5787# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X176 VSS VDD a_16704_5987# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X177 a_14262_6709# a_13844_6793# a_14018_6401# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X178 a_16236_5513# a_15955_5147# a_16143_5147# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X179 a_16143_7067# x1[1].D VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X180 VSS a_17191_7041# a_17898_7083# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X181 a_14483_5429# a_14018_5121# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X182 VSS VDD a_14312_7267# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X183 a_16550_5147# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X184 a_12385_8554# eob a_12297_8554# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X185 a_17307_6427# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X186 a_17307_6427# a_16704_6401# a_17191_6401# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X187 a_14799_5761# a_14625_6165# a_14915_6153# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X188 a_13844_5513# a_13563_5147# a_13751_5147# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X189 a_13751_7067# x1[0].D VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X190 VDD a_14312_7267# a_15033_7067# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X191 VDD a_17191_7041# a_17103_7067# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X192 a_15033_6709# a_14625_6427# a_14799_6401# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X193 a_17017_6427# a_15789_6427# a_16875_6709# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X194 a_13563_7073# a_13397_7073# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X195 a_17191_5121# a_17017_5147# a_17307_5147# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X196 a_17191_5761# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X197 VDD a_16410_7041# a_16320_7067# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X198 a_14915_6427# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X199 VSS a_17191_5121# a_17898_5147# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X200 VDD a_16704_6401# a_17425_6709# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X201 a_17103_5513# a_15955_5147# a_17017_5147# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X202 VSS VDD a_14312_5121# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X203 x2.x5[7].floating x2.x10.Y x2.x9.output_stack VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X204 VDD x3.A a_18499_9105# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X205 VDD x3.A a_18195_9015# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0651 ps=0.73 w=0.42 l=0.15
X206 a_14158_7433# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X207 VSS x3.A a_18499_9105# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X208 VDD a_14799_6401# a_15506_6427# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X209 x2.x5[7].floating x2.x10.Y x2.x9.output_stack VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X210 x1[3].Q_N a_17191_6401# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X211 a_14625_6165# a_13397_5793# a_14483_5787# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X212 x1[6].Q_N a_14799_5121# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X213 a_14711_5513# a_13563_5147# a_14625_5147# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X214 a_12410_9943# eob a_12322_10081# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X215 a_16344_7445# a_15955_7073# a_16236_7067# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X216 VDD a_14799_5761# a_14711_5787# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X217 a_16550_5147# a_16704_5121# a_16410_5121# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X218 a_18195_9356# x3.A VSS VDD sky130_fd_pr__pfet_01v8_hvt ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X219 a_17017_6427# a_15955_6427# a_16922_6427# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X220 VSS a_14799_7041# a_15506_7083# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X221 a_14799_6401# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X222 a_14158_6427# a_14312_6401# a_14018_6401# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X223 a_14158_5147# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X224 a_12410_10219# eob a_12322_10357# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X225 a_13952_7445# a_13563_7073# a_13844_7067# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X226 a_16320_7067# a_15789_7073# a_16236_7067# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X227 a_17307_7433# a_16704_7267# a_17191_7041# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X228 a_17017_6165# a_15955_5793# a_16922_6109# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X229 a_17017_5147# a_15789_5147# a_16875_5429# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X230 VDD x3.X a_15789_6427# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X231 x2.x5[7].floating x2.x10.Y x2.x9.output_stack VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X232 a_14625_7445# a_13563_7073# a_14530_7389# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X233 VDD a_14018_7041# a_13928_7067# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X234 a_15955_5793# a_15789_5793# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X235 a_14799_5121# a_14625_5147# a_14915_5147# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X236 VDD a_18499_9105# x3.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X237 a_12457_8416# eob a_12385_8554# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X238 a_17126_6427# a_15789_6427# a_17017_6427# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X239 VSS a_14799_5121# a_15506_5147# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X240 a_13563_7073# a_13397_7073# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X241 a_16143_6427# x1[3].D VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X242 x1[7].Q a_17898_5147# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X243 x2.x9.output_stack eob a_12322_9805# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X244 x1[0].Q_N a_14799_7041# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X245 VSS x3.X a_15789_6427# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X246 a_17126_6165# a_15789_5793# a_17017_6165# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X247 a_13563_5147# a_13397_5147# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X248 a_16875_5787# a_16410_5761# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X249 x1[6].Q a_15506_5147# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X250 a_12385_8140# eob a_12297_8002# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X251 a_13751_6427# x1[2].D VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X252 VSS a_17191_6401# a_17126_6427# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X253 a_13928_5787# a_13397_5793# a_13844_5787# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X254 VSS a_16410_6401# a_16344_6427# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X255 x1[1].Q_N a_17191_7041# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X256 a_13563_5147# a_13397_5147# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X257 a_14018_6401# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X258 VDD VDD a_16704_6401# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X259 a_14799_5121# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X260 a_12385_8416# eob a_12297_8278# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X261 a_14158_7433# a_14312_7267# a_14018_7041# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X262 a_16654_7067# a_16236_7067# a_16410_7041# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X263 VDD a_14312_5987# a_14262_5787# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X264 a_17307_6153# a_16704_5987# a_17191_5761# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X265 VDD x3.X a_13397_6427# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X266 a_14483_7067# a_14018_7041# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X267 x1[1].Q a_17898_7083# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X268 x2.x9.output_stack x2.x10.Y x2.x5[7].floating VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X269 VSS a_14799_7041# a_14734_7445# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X270 a_16410_7041# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X271 a_17425_5429# a_17017_5147# a_17191_5121# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X272 x1[0].Q a_15506_7083# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X273 VSS x3.X a_13397_6427# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X274 a_16875_6709# a_16410_6401# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X275 x1[4].Q_N a_14799_5761# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X276 VDD VDD a_14312_5987# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X277 a_14734_5147# a_13397_5147# a_14625_5147# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X278 x2.x10.Y x2.x10.A VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X279 a_16236_7067# a_15955_7073# a_16143_7067# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X280 a_16236_5513# a_15789_5147# a_16143_5147# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X281 a_16143_5787# x1[5].D VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X282 x2.x2.floating x2.x2.SW x2.x9.output_stack VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.124 ps=1.43 w=0.42 l=0.15
X283 a_16550_6153# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X284 VDD a_16704_5121# a_16654_5429# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X285 VSS a_14799_5121# a_14734_5147# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X286 a_13844_7067# a_13563_7073# a_13751_7067# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X287 a_17307_7433# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X288 VSS a_14018_6401# a_13952_6427# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X289 VSS x3.A a_18195_9356# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0651 ps=0.73 w=0.42 l=0.15
X290 VDD a_14312_6401# a_14262_6709# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X291 a_13751_5787# x1[4].D VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X292 VDD a_14312_5987# a_15033_5787# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X293 VDD a_17191_5121# a_17898_5147# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X294 a_13844_5513# a_13397_5147# a_13751_5147# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X295 VDD a_17191_5761# a_17103_5787# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X296 a_17191_6401# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X297 a_16922_6427# a_16410_6401# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X298 VDD VDD a_16704_5121# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X299 a_14018_5121# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X300 a_14915_7433# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X301 VDD x3.X a_15789_7073# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X302 VSS VDD a_16704_6401# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X303 a_13563_5793# a_13397_5793# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X304 a_14158_6153# a_14312_5987# a_14018_5761# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X305 VDD a_16410_5761# a_16320_5787# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X306 a_14262_5429# a_13844_5513# a_14018_5121# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X307 a_12410_10219# eob a_12322_10081# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X308 x2.x9.output_stack x2.x6.SW x2.x6.floating VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X309 x2.x4[3].floating x2.code[2] x2.x9.output_stack VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X310 a_12385_8830# eob a_12297_8830# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X311 a_12457_8140# eob a_12385_8140# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X312 VSS a_17191_5761# a_17898_5803# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X313 a_17103_7067# a_15955_7073# a_17017_7445# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X314 VSS VDD a_14312_5987# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X315 a_17307_5147# a_16704_5121# a_17191_5121# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X316 a_17307_5147# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X317 x1[5].Q a_17898_5803# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X318 a_12457_8416# eob a_12385_8416# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X319 x1[3].Q_N a_17191_6401# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X320 a_15033_5429# a_14625_5147# a_14799_5121# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X321 a_14711_7067# a_13563_7073# a_14625_7445# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X322 a_14915_6427# a_14312_6401# a_14799_6401# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X323 x1[4].Q a_15506_5803# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X324 a_14625_6427# a_13397_6427# a_14483_6709# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X325 VDD a_14799_6401# a_14711_6793# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X326 a_14915_5147# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X327 VDD a_16704_5121# a_17425_5429# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X328 a_12385_8002# eob a_12297_8002# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X329 a_16410_6401# a_16236_6793# a_16550_6427# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X330 a_14158_6153# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X331 a_17017_7445# a_15789_7073# a_16875_7067# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X332 VDD a_14312_6401# a_15033_6709# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X333 a_16344_6427# a_15955_6427# a_16236_6793# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X334 a_16320_5787# a_15789_5793# a_16236_5787# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X335 VDD a_14799_5121# a_15506_5147# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X336 x1[7].Q_N a_17191_5121# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X337 VSS x2.x7.SW x2.x6.SW VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X338 x2.x9.output_stack x2.code[2] x2.x4[3].floating VSS sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X339 a_16922_7389# a_16410_7041# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X340 a_14530_6427# a_14018_6401# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X341 VDD a_14018_5761# a_13928_5787# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X342 a_17191_5121# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X343 VSS a_18499_9105# x3.X VSS sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X344 VDD x3.X a_13397_7073# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X345 a_16344_6165# a_15955_5793# a_16236_5787# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X346 x2.x5[7].floating x2.x10.Y x2.x9.output_stack VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X347 a_13952_6427# a_13563_6427# a_13844_6793# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X348 x1[2].Q_N a_14799_6401# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X349 VSS a_14799_5761# a_15506_5803# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X350 a_17017_5147# a_15955_5147# a_16922_5147# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X351 a_16143_7067# x1[1].D VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X352 a_15955_6427# a_15789_6427# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X353 a_14158_5147# a_14312_5121# a_14018_5121# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X354 x2.x4[3].floating x2.code[2] x2.x9.output_stack VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X355 VSS x3.X a_15789_7073# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X356 a_14625_6427# a_13563_6427# a_14530_6427# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X357 a_13952_6165# a_13563_5793# a_13844_5787# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X358 VDD x3.X a_15789_5147# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X359 a_12457_8692# eob a_12385_8830# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X360 a_13751_7067# x1[0].D VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X361 a_14915_7433# a_14312_7267# a_14799_7041# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X362 VSS a_17191_7041# a_17126_7445# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X363 a_13928_6793# a_13397_6427# a_13844_6793# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X364 a_14625_6165# a_13563_5793# a_14530_6109# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X365 a_14625_5147# a_13397_5147# a_14483_5429# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X366 VSS a_16410_7041# a_16344_7445# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X367 a_15955_6427# a_15789_6427# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X368 a_17126_5147# a_15789_5147# a_17017_5147# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X369 VDD a_14799_5121# a_14711_5513# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X370 a_14799_7041# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X371 x1[5].Q_N a_17191_5761# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X372 a_18195_9015# x2.x9.output_stack x3.A VSS sky130_fd_pr__nfet_01v8 ad=0.0651 pd=0.73 as=0.122 ps=1.42 w=0.42 l=0.15
X373 a_17425_7067# a_17017_7445# a_17191_7041# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X374 a_13563_5793# a_13397_5793# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X375 a_16143_5147# x1[7].D VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X376 VSS x3.X a_15789_5147# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt hgu_sarlogic ready ext_clk sample_clk sample_clk_b sar_clk VSS VDD sel_bit[0]
+ sel_bit[1] sar_result[1] sar_result[2] sar_result[3] sar_result[5] sar_result[4]
+ sar_result[6] sar_result[7] sar_result[0] sample_delay_cap_ctrl_code[2] sample_delay_cap_ctrl_code[1]
+ sample_delay_cap_ctrl_code[0] sample_delay_cap_ctrl_code[6] sample_delay_cap_ctrl_code[5]
+ sample_delay_cap_ctrl_code[4] sample_delay_offset sample_delay_cap_ctrl_code[3]
+ sample_delay_cap_ctrl_code[7] sample_delay_cap_ctrl_code[11] sample_delay_cap_ctrl_code[15]
+ async_setb_delay_cap_ctrl_code[2] async_setb_delay_cap_ctrl_code[1] async_setb_delay_cap_ctrl_code[0]
+ async_resetb_delay_cap_ctrl_code[0] async_resetb_delay_cap_ctrl_code[1] async_resetb_delay_cap_ctrl_code[2]
+ async_setb_delay_cap_ctrl_code[3] async_resetb_delay_cap_ctrl_code[3] async_delay_offset
+ retimer_eob_delay_offset retimer_delay_code[3] retimer_delay_code[2] retimer_delay_code[1]
+ retimer_delay_code[0] comp_result vss_sw[7] vss_sw[6] vss_sw[5] vss_sw[4] vss_sw[3]
+ vss_sw[2] vss_sw[1] vdd_sw[7] vdd_sw[6] vdd_sw[5] vdd_sw[4] vdd_sw[3] vdd_sw[2]
+ vdd_sw[1] vss_sw_b[7] vss_sw_b[6] vss_sw_b[5] vss_sw_b[4] vss_sw_b[3] vss_sw_b[2]
+ vss_sw_b[1] vdd_sw_b[1] vdd_sw_b[2] vdd_sw_b[3] vdd_sw_b[4] vdd_sw_b[5] vdd_sw_b[6]
+ vdd_sw_b[7] sample_delay_cap_ctrl_code[9] sample_delay_cap_ctrl_code[8] sample_delay_cap_ctrl_code[14]
+ sample_delay_cap_ctrl_code[13] sample_delay_cap_ctrl_code[12] sample_delay_cap_ctrl_code[10]
Xx1 sample_clk x5/eob ready async_delay_offset sar_clk async_resetb_delay_cap_ctrl_code[2]
+ async_resetb_delay_cap_ctrl_code[1] async_setb_delay_cap_ctrl_code[3] async_setb_delay_cap_ctrl_code[1]
+ async_setb_delay_cap_ctrl_code[2] async_resetb_delay_cap_ctrl_code[0] async_resetb_delay_cap_ctrl_code[3]
+ async_setb_delay_cap_ctrl_code[0] VSS VDD hgu_clk_async
Xx2 VSS VSS sample_delay_offset sample_delay_cap_ctrl_code[2] sample_delay_cap_ctrl_code[1]
+ sample_delay_cap_ctrl_code[6] sample_delay_cap_ctrl_code[5] sample_delay_cap_ctrl_code[4]
+ sample_delay_cap_ctrl_code[10] sample_delay_cap_ctrl_code[9] sample_delay_cap_ctrl_code[14]
+ sample_delay_cap_ctrl_code[13] sample_delay_cap_ctrl_code[12] sample_delay_cap_ctrl_code[7]
+ sample_delay_cap_ctrl_code[15] sample_clk_b sample_clk ext_clk sample_delay_cap_ctrl_code[11]
+ sample_delay_cap_ctrl_code[0] sample_delay_cap_ctrl_code[3] sample_delay_cap_ctrl_code[8]
+ VDD VSS hgu_clk_sample
Xx3 sel_bit[0] sel_bit[1] sample_clk_b x5/eob comp_result x4/x5.D x4/D[6] x4/x7.S
+ x4/D[5] x4/x20.S x4/x9.S x4/x17.S x4/x11.S x4/x15.S x4/x13.S x4/D[2] x4/D[3] x4/D[1]
+ x4/D[4] x3/D[0] sar_clk VSS VDD hgu_sarlogic_8bit_logic
Xx4 vss_sw[1] vss_sw[2] vss_sw[3] vss_sw[4] vss_sw[5] vss_sw[6] vss_sw[7] vdd_sw[2]
+ vdd_sw[3] vdd_sw[4] vdd_sw[5] vdd_sw[6] vdd_sw[7] x4/D[2] x4/D[3] x4/D[4] x4/D[5]
+ x4/D[6] x4/x5.D x4/x20.S x4/x17.S x4/x15.S x4/x13.S x4/x11.S x4/x9.S x4/x7.S vdd_sw_b[1]
+ vdd_sw_b[2] vdd_sw_b[3] vdd_sw_b[4] vdd_sw_b[5] vdd_sw_b[6] vdd_sw_b[7] vss_sw_b[1]
+ vss_sw_b[2] vss_sw_b[3] vss_sw_b[4] vss_sw_b[5] vss_sw_b[6] vss_sw_b[7] x4/D[1]
+ vdd_sw[1] sar_clk sample_clk_b VSS VDD hgu_sarlogic_sw_ctrl
Xx5 x5/eob retimer_delay_code[2] retimer_delay_code[1] retimer_delay_code[3] x4/D[1]
+ x4/D[2] x4/D[5] x4/D[4] sar_result[1] sar_result[0] sar_result[3] sar_result[2]
+ sar_result[5] sar_result[4] sar_result[7] sar_result[6] x4/D[6] x4/x5.D x4/D[3]
+ x3/D[0] retimer_eob_delay_offset retimer_delay_code[0] VSS VDD hgu_sarlogic_retimer
.ends

