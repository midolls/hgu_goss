magic
tech sky130A
magscale 1 2
timestamp 1697393286
<< pwell >>
rect 1926 3419 1947 3468
<< metal1 >>
rect 750 4461 3032 4468
rect 750 4412 838 4461
rect 750 4360 757 4412
rect 809 4409 838 4412
rect 890 4409 902 4461
rect 954 4409 966 4461
rect 1018 4409 1030 4461
rect 1082 4409 1094 4461
rect 1146 4409 1158 4461
rect 1210 4409 1222 4461
rect 1274 4409 1286 4461
rect 1338 4409 1350 4461
rect 1402 4409 1414 4461
rect 1466 4409 1478 4461
rect 1530 4409 1542 4461
rect 1594 4409 1606 4461
rect 1658 4409 1670 4461
rect 1722 4409 1734 4461
rect 1786 4409 1996 4461
rect 2048 4409 2060 4461
rect 2112 4409 2124 4461
rect 2176 4409 2188 4461
rect 2240 4409 2252 4461
rect 2304 4409 2316 4461
rect 2368 4409 2380 4461
rect 2432 4409 2444 4461
rect 2496 4409 2508 4461
rect 2560 4409 2572 4461
rect 2624 4409 2636 4461
rect 2688 4409 2700 4461
rect 2752 4409 2764 4461
rect 2816 4409 2828 4461
rect 2880 4409 2892 4461
rect 2944 4412 3032 4461
rect 2944 4409 2973 4412
rect 809 4402 2973 4409
rect 809 4360 822 4402
rect 750 4348 822 4360
rect 750 4296 757 4348
rect 809 4296 822 4348
rect 750 4284 822 4296
rect 750 4232 757 4284
rect 809 4232 822 4284
rect 750 4220 822 4232
rect 750 4168 757 4220
rect 809 4168 822 4220
rect 750 4156 822 4168
rect 750 4104 757 4156
rect 809 4104 822 4156
rect 750 4092 822 4104
rect 750 4040 757 4092
rect 809 4040 822 4092
rect 750 4028 822 4040
rect 750 3976 757 4028
rect 809 3976 822 4028
rect 750 3964 822 3976
rect 750 3912 757 3964
rect 809 3912 822 3964
rect 750 3900 822 3912
rect 750 3848 757 3900
rect 809 3848 822 3900
rect 750 3836 822 3848
rect 750 3784 757 3836
rect 809 3784 822 3836
rect 750 3772 822 3784
rect 750 3720 757 3772
rect 809 3720 822 3772
rect 750 3708 822 3720
rect 750 3656 757 3708
rect 809 3656 822 3708
rect 750 3644 822 3656
rect 750 3592 757 3644
rect 809 3592 822 3644
rect 750 3580 822 3592
rect 750 3528 757 3580
rect 809 3528 822 3580
rect 750 3516 822 3528
rect 750 3464 757 3516
rect 809 3464 822 3516
rect 750 3452 822 3464
rect 750 3400 757 3452
rect 809 3400 822 3452
rect 750 3198 822 3400
rect 750 3146 757 3198
rect 809 3146 822 3198
rect 750 3134 822 3146
rect 750 3082 757 3134
rect 809 3082 822 3134
rect 750 3070 822 3082
rect 750 3018 757 3070
rect 809 3018 822 3070
rect 750 3006 822 3018
rect 750 2954 757 3006
rect 809 2954 822 3006
rect 750 2942 822 2954
rect 750 2890 757 2942
rect 809 2890 822 2942
rect 750 2878 822 2890
rect 750 2826 757 2878
rect 809 2826 822 2878
rect 750 2814 822 2826
rect 750 2762 757 2814
rect 809 2762 822 2814
rect 750 2750 822 2762
rect 750 2698 757 2750
rect 809 2698 822 2750
rect 750 2686 822 2698
rect 750 2634 757 2686
rect 809 2634 822 2686
rect 750 2622 822 2634
rect 750 2570 757 2622
rect 809 2570 822 2622
rect 750 2558 822 2570
rect 750 2506 757 2558
rect 809 2506 822 2558
rect 750 2494 822 2506
rect 750 2442 757 2494
rect 809 2442 822 2494
rect 750 2430 822 2442
rect 750 2378 757 2430
rect 809 2378 822 2430
rect 750 2366 822 2378
rect 750 2314 757 2366
rect 809 2314 822 2366
rect 750 2302 822 2314
rect 750 2250 757 2302
rect 809 2250 822 2302
rect 750 2238 822 2250
rect 750 2186 757 2238
rect 809 2196 822 2238
rect 850 3331 878 4374
rect 906 3359 934 4402
rect 962 3331 990 4374
rect 1018 3359 1046 4402
rect 1074 3331 1102 4374
rect 1130 3359 1158 4402
rect 1186 3331 1214 4374
rect 1242 3359 1270 4402
rect 1298 3331 1326 4374
rect 1354 3359 1382 4402
rect 1410 3331 1438 4374
rect 1466 3359 1494 4402
rect 1522 3331 1550 4374
rect 1578 3359 1606 4402
rect 1634 3331 1662 4374
rect 1690 3359 1718 4402
rect 1746 3331 1774 4374
rect 1802 3359 1830 4402
rect 1858 4367 1924 4374
rect 1858 4315 1865 4367
rect 1917 4315 1924 4367
rect 1858 4303 1924 4315
rect 1858 4251 1865 4303
rect 1917 4251 1924 4303
rect 1858 4239 1924 4251
rect 1858 4187 1865 4239
rect 1917 4187 1924 4239
rect 1858 4175 1924 4187
rect 1858 4123 1865 4175
rect 1917 4123 1924 4175
rect 1858 4111 1924 4123
rect 1858 4059 1865 4111
rect 1917 4059 1924 4111
rect 1858 4047 1924 4059
rect 1858 3995 1865 4047
rect 1917 3995 1924 4047
rect 1858 3983 1924 3995
rect 1858 3931 1865 3983
rect 1917 3931 1924 3983
rect 1858 3919 1924 3931
rect 1858 3867 1865 3919
rect 1917 3867 1924 3919
rect 1858 3855 1924 3867
rect 1858 3803 1865 3855
rect 1917 3803 1924 3855
rect 1858 3791 1924 3803
rect 1858 3739 1865 3791
rect 1917 3739 1924 3791
rect 1858 3727 1924 3739
rect 1858 3675 1865 3727
rect 1917 3675 1924 3727
rect 1858 3663 1924 3675
rect 1858 3611 1865 3663
rect 1917 3611 1924 3663
rect 1858 3599 1924 3611
rect 1858 3547 1865 3599
rect 1917 3547 1924 3599
rect 1858 3535 1924 3547
rect 1858 3483 1865 3535
rect 1917 3483 1924 3535
rect 1858 3471 1924 3483
rect 1858 3419 1865 3471
rect 1917 3419 1924 3471
rect 1858 3407 1924 3419
rect 1858 3355 1865 3407
rect 1917 3355 1924 3407
rect 1952 3359 1980 4402
rect 1858 3331 1924 3355
rect 2008 3331 2036 4374
rect 2064 3359 2092 4402
rect 2120 3331 2148 4374
rect 2176 3359 2204 4402
rect 2232 3331 2260 4374
rect 2288 3359 2316 4402
rect 2344 3331 2372 4374
rect 2400 3359 2428 4402
rect 2456 3331 2484 4374
rect 2512 3359 2540 4402
rect 2568 3331 2596 4374
rect 2624 3359 2652 4402
rect 2680 3331 2708 4374
rect 2736 3359 2764 4402
rect 2792 3331 2820 4374
rect 2848 3359 2876 4402
rect 2904 3331 2932 4374
rect 850 3325 2932 3331
rect 850 3273 902 3325
rect 954 3273 966 3325
rect 1018 3273 1030 3325
rect 1082 3273 1094 3325
rect 1146 3273 1158 3325
rect 1210 3273 1222 3325
rect 1274 3273 1286 3325
rect 1338 3273 1350 3325
rect 1402 3273 1414 3325
rect 1466 3273 1478 3325
rect 1530 3273 1542 3325
rect 1594 3273 1606 3325
rect 1658 3273 1670 3325
rect 1722 3273 1734 3325
rect 1786 3273 1798 3325
rect 1850 3273 1932 3325
rect 1984 3273 1996 3325
rect 2048 3273 2060 3325
rect 2112 3273 2124 3325
rect 2176 3273 2188 3325
rect 2240 3273 2252 3325
rect 2304 3273 2316 3325
rect 2368 3273 2380 3325
rect 2432 3273 2444 3325
rect 2496 3273 2508 3325
rect 2560 3273 2572 3325
rect 2624 3273 2636 3325
rect 2688 3273 2700 3325
rect 2752 3273 2764 3325
rect 2816 3273 2828 3325
rect 2880 3273 2932 3325
rect 850 3267 2932 3273
rect 850 2224 878 3267
rect 906 2196 934 3239
rect 962 2224 990 3267
rect 1018 2196 1046 3239
rect 1074 2224 1102 3267
rect 1130 2196 1158 3239
rect 1186 2224 1214 3267
rect 1242 2196 1270 3239
rect 1298 2224 1326 3267
rect 1354 2196 1382 3239
rect 1410 2224 1438 3267
rect 1466 2196 1494 3239
rect 1522 2224 1550 3267
rect 1578 2196 1606 3239
rect 1634 2224 1662 3267
rect 1690 2196 1718 3239
rect 1746 2224 1774 3267
rect 1858 3243 1924 3267
rect 1802 2196 1830 3239
rect 1858 3191 1865 3243
rect 1917 3191 1924 3243
rect 1858 3179 1924 3191
rect 1858 3127 1865 3179
rect 1917 3127 1924 3179
rect 1858 3115 1924 3127
rect 1858 3063 1865 3115
rect 1917 3063 1924 3115
rect 1858 3051 1924 3063
rect 1858 2999 1865 3051
rect 1917 2999 1924 3051
rect 1858 2987 1924 2999
rect 1858 2935 1865 2987
rect 1917 2935 1924 2987
rect 1858 2923 1924 2935
rect 1858 2871 1865 2923
rect 1917 2871 1924 2923
rect 1858 2859 1924 2871
rect 1858 2807 1865 2859
rect 1917 2807 1924 2859
rect 1858 2795 1924 2807
rect 1858 2743 1865 2795
rect 1917 2743 1924 2795
rect 1858 2731 1924 2743
rect 1858 2679 1865 2731
rect 1917 2679 1924 2731
rect 1858 2667 1924 2679
rect 1858 2615 1865 2667
rect 1917 2615 1924 2667
rect 1858 2603 1924 2615
rect 1858 2551 1865 2603
rect 1917 2551 1924 2603
rect 1858 2539 1924 2551
rect 1858 2487 1865 2539
rect 1917 2487 1924 2539
rect 1858 2475 1924 2487
rect 1858 2423 1865 2475
rect 1917 2423 1924 2475
rect 1858 2411 1924 2423
rect 1858 2359 1865 2411
rect 1917 2359 1924 2411
rect 1858 2347 1924 2359
rect 1858 2295 1865 2347
rect 1917 2295 1924 2347
rect 1858 2283 1924 2295
rect 1858 2231 1865 2283
rect 1917 2231 1924 2283
rect 1858 2224 1924 2231
rect 1952 2196 1980 3239
rect 2008 2224 2036 3267
rect 2064 2196 2092 3239
rect 2120 2224 2148 3267
rect 2176 2196 2204 3239
rect 2232 2224 2260 3267
rect 2288 2196 2316 3239
rect 2344 2224 2372 3267
rect 2400 2196 2428 3239
rect 2456 2224 2484 3267
rect 2512 2196 2540 3239
rect 2568 2224 2596 3267
rect 2624 2196 2652 3239
rect 2680 2224 2708 3267
rect 2736 2196 2764 3239
rect 2792 2224 2820 3267
rect 2848 2196 2876 3239
rect 2904 2224 2932 3267
rect 2960 4360 2973 4402
rect 3025 4360 3032 4412
rect 2960 4348 3032 4360
rect 2960 4296 2973 4348
rect 3025 4296 3032 4348
rect 2960 4284 3032 4296
rect 2960 4232 2973 4284
rect 3025 4232 3032 4284
rect 2960 4220 3032 4232
rect 2960 4168 2973 4220
rect 3025 4168 3032 4220
rect 2960 4156 3032 4168
rect 2960 4104 2973 4156
rect 3025 4104 3032 4156
rect 2960 4092 3032 4104
rect 2960 4040 2973 4092
rect 3025 4040 3032 4092
rect 2960 4028 3032 4040
rect 2960 3976 2973 4028
rect 3025 3976 3032 4028
rect 2960 3964 3032 3976
rect 2960 3912 2973 3964
rect 3025 3912 3032 3964
rect 2960 3900 3032 3912
rect 2960 3848 2973 3900
rect 3025 3848 3032 3900
rect 2960 3836 3032 3848
rect 2960 3784 2973 3836
rect 3025 3784 3032 3836
rect 2960 3772 3032 3784
rect 2960 3720 2973 3772
rect 3025 3720 3032 3772
rect 2960 3708 3032 3720
rect 2960 3656 2973 3708
rect 3025 3656 3032 3708
rect 2960 3644 3032 3656
rect 2960 3592 2973 3644
rect 3025 3592 3032 3644
rect 2960 3580 3032 3592
rect 2960 3528 2973 3580
rect 3025 3528 3032 3580
rect 2960 3516 3032 3528
rect 2960 3464 2973 3516
rect 3025 3464 3032 3516
rect 2960 3452 3032 3464
rect 2960 3400 2973 3452
rect 3025 3400 3032 3452
rect 2960 3198 3032 3400
rect 2960 3146 2973 3198
rect 3025 3146 3032 3198
rect 2960 3134 3032 3146
rect 2960 3082 2973 3134
rect 3025 3082 3032 3134
rect 2960 3070 3032 3082
rect 2960 3018 2973 3070
rect 3025 3018 3032 3070
rect 2960 3006 3032 3018
rect 2960 2954 2973 3006
rect 3025 2954 3032 3006
rect 2960 2942 3032 2954
rect 2960 2890 2973 2942
rect 3025 2890 3032 2942
rect 2960 2878 3032 2890
rect 2960 2826 2973 2878
rect 3025 2826 3032 2878
rect 2960 2814 3032 2826
rect 2960 2762 2973 2814
rect 3025 2762 3032 2814
rect 2960 2750 3032 2762
rect 2960 2698 2973 2750
rect 3025 2698 3032 2750
rect 2960 2686 3032 2698
rect 2960 2634 2973 2686
rect 3025 2634 3032 2686
rect 2960 2622 3032 2634
rect 2960 2570 2973 2622
rect 3025 2570 3032 2622
rect 2960 2558 3032 2570
rect 2960 2506 2973 2558
rect 3025 2506 3032 2558
rect 2960 2494 3032 2506
rect 2960 2442 2973 2494
rect 3025 2442 3032 2494
rect 2960 2430 3032 2442
rect 2960 2378 2973 2430
rect 3025 2378 3032 2430
rect 2960 2366 3032 2378
rect 2960 2314 2973 2366
rect 3025 2314 3032 2366
rect 2960 2302 3032 2314
rect 2960 2250 2973 2302
rect 3025 2250 3032 2302
rect 2960 2238 3032 2250
rect 2960 2196 2973 2238
rect 809 2189 2973 2196
rect 809 2186 838 2189
rect 750 2137 838 2186
rect 890 2137 902 2189
rect 954 2137 966 2189
rect 1018 2137 1030 2189
rect 1082 2137 1094 2189
rect 1146 2137 1158 2189
rect 1210 2137 1222 2189
rect 1274 2137 1286 2189
rect 1338 2137 1350 2189
rect 1402 2137 1414 2189
rect 1466 2137 1478 2189
rect 1530 2137 1542 2189
rect 1594 2137 1606 2189
rect 1658 2137 1670 2189
rect 1722 2137 1734 2189
rect 1786 2137 1996 2189
rect 2048 2137 2060 2189
rect 2112 2137 2124 2189
rect 2176 2137 2188 2189
rect 2240 2137 2252 2189
rect 2304 2137 2316 2189
rect 2368 2137 2380 2189
rect 2432 2137 2444 2189
rect 2496 2137 2508 2189
rect 2560 2137 2572 2189
rect 2624 2137 2636 2189
rect 2688 2137 2700 2189
rect 2752 2137 2764 2189
rect 2816 2137 2828 2189
rect 2880 2137 2892 2189
rect 2944 2186 2973 2189
rect 3025 2186 3032 2238
rect 2944 2137 3032 2186
rect 750 2130 3032 2137
<< via1 >>
rect 757 4360 809 4412
rect 838 4409 890 4461
rect 902 4409 954 4461
rect 966 4409 1018 4461
rect 1030 4409 1082 4461
rect 1094 4409 1146 4461
rect 1158 4409 1210 4461
rect 1222 4409 1274 4461
rect 1286 4409 1338 4461
rect 1350 4409 1402 4461
rect 1414 4409 1466 4461
rect 1478 4409 1530 4461
rect 1542 4409 1594 4461
rect 1606 4409 1658 4461
rect 1670 4409 1722 4461
rect 1734 4409 1786 4461
rect 1996 4409 2048 4461
rect 2060 4409 2112 4461
rect 2124 4409 2176 4461
rect 2188 4409 2240 4461
rect 2252 4409 2304 4461
rect 2316 4409 2368 4461
rect 2380 4409 2432 4461
rect 2444 4409 2496 4461
rect 2508 4409 2560 4461
rect 2572 4409 2624 4461
rect 2636 4409 2688 4461
rect 2700 4409 2752 4461
rect 2764 4409 2816 4461
rect 2828 4409 2880 4461
rect 2892 4409 2944 4461
rect 757 4296 809 4348
rect 757 4232 809 4284
rect 757 4168 809 4220
rect 757 4104 809 4156
rect 757 4040 809 4092
rect 757 3976 809 4028
rect 757 3912 809 3964
rect 757 3848 809 3900
rect 757 3784 809 3836
rect 757 3720 809 3772
rect 757 3656 809 3708
rect 757 3592 809 3644
rect 757 3528 809 3580
rect 757 3464 809 3516
rect 757 3400 809 3452
rect 757 3146 809 3198
rect 757 3082 809 3134
rect 757 3018 809 3070
rect 757 2954 809 3006
rect 757 2890 809 2942
rect 757 2826 809 2878
rect 757 2762 809 2814
rect 757 2698 809 2750
rect 757 2634 809 2686
rect 757 2570 809 2622
rect 757 2506 809 2558
rect 757 2442 809 2494
rect 757 2378 809 2430
rect 757 2314 809 2366
rect 757 2250 809 2302
rect 757 2186 809 2238
rect 1865 4315 1917 4367
rect 1865 4251 1917 4303
rect 1865 4187 1917 4239
rect 1865 4123 1917 4175
rect 1865 4059 1917 4111
rect 1865 3995 1917 4047
rect 1865 3931 1917 3983
rect 1865 3867 1917 3919
rect 1865 3803 1917 3855
rect 1865 3739 1917 3791
rect 1865 3675 1917 3727
rect 1865 3611 1917 3663
rect 1865 3547 1917 3599
rect 1865 3483 1917 3535
rect 1865 3419 1917 3471
rect 1865 3355 1917 3407
rect 902 3273 954 3325
rect 966 3273 1018 3325
rect 1030 3273 1082 3325
rect 1094 3273 1146 3325
rect 1158 3273 1210 3325
rect 1222 3273 1274 3325
rect 1286 3273 1338 3325
rect 1350 3273 1402 3325
rect 1414 3273 1466 3325
rect 1478 3273 1530 3325
rect 1542 3273 1594 3325
rect 1606 3273 1658 3325
rect 1670 3273 1722 3325
rect 1734 3273 1786 3325
rect 1798 3273 1850 3325
rect 1932 3273 1984 3325
rect 1996 3273 2048 3325
rect 2060 3273 2112 3325
rect 2124 3273 2176 3325
rect 2188 3273 2240 3325
rect 2252 3273 2304 3325
rect 2316 3273 2368 3325
rect 2380 3273 2432 3325
rect 2444 3273 2496 3325
rect 2508 3273 2560 3325
rect 2572 3273 2624 3325
rect 2636 3273 2688 3325
rect 2700 3273 2752 3325
rect 2764 3273 2816 3325
rect 2828 3273 2880 3325
rect 1865 3191 1917 3243
rect 1865 3127 1917 3179
rect 1865 3063 1917 3115
rect 1865 2999 1917 3051
rect 1865 2935 1917 2987
rect 1865 2871 1917 2923
rect 1865 2807 1917 2859
rect 1865 2743 1917 2795
rect 1865 2679 1917 2731
rect 1865 2615 1917 2667
rect 1865 2551 1917 2603
rect 1865 2487 1917 2539
rect 1865 2423 1917 2475
rect 1865 2359 1917 2411
rect 1865 2295 1917 2347
rect 1865 2231 1917 2283
rect 2973 4360 3025 4412
rect 2973 4296 3025 4348
rect 2973 4232 3025 4284
rect 2973 4168 3025 4220
rect 2973 4104 3025 4156
rect 2973 4040 3025 4092
rect 2973 3976 3025 4028
rect 2973 3912 3025 3964
rect 2973 3848 3025 3900
rect 2973 3784 3025 3836
rect 2973 3720 3025 3772
rect 2973 3656 3025 3708
rect 2973 3592 3025 3644
rect 2973 3528 3025 3580
rect 2973 3464 3025 3516
rect 2973 3400 3025 3452
rect 2973 3146 3025 3198
rect 2973 3082 3025 3134
rect 2973 3018 3025 3070
rect 2973 2954 3025 3006
rect 2973 2890 3025 2942
rect 2973 2826 3025 2878
rect 2973 2762 3025 2814
rect 2973 2698 3025 2750
rect 2973 2634 3025 2686
rect 2973 2570 3025 2622
rect 2973 2506 3025 2558
rect 2973 2442 3025 2494
rect 2973 2378 3025 2430
rect 2973 2314 3025 2366
rect 2973 2250 3025 2302
rect 838 2137 890 2189
rect 902 2137 954 2189
rect 966 2137 1018 2189
rect 1030 2137 1082 2189
rect 1094 2137 1146 2189
rect 1158 2137 1210 2189
rect 1222 2137 1274 2189
rect 1286 2137 1338 2189
rect 1350 2137 1402 2189
rect 1414 2137 1466 2189
rect 1478 2137 1530 2189
rect 1542 2137 1594 2189
rect 1606 2137 1658 2189
rect 1670 2137 1722 2189
rect 1734 2137 1786 2189
rect 1996 2137 2048 2189
rect 2060 2137 2112 2189
rect 2124 2137 2176 2189
rect 2188 2137 2240 2189
rect 2252 2137 2304 2189
rect 2316 2137 2368 2189
rect 2380 2137 2432 2189
rect 2444 2137 2496 2189
rect 2508 2137 2560 2189
rect 2572 2137 2624 2189
rect 2636 2137 2688 2189
rect 2700 2137 2752 2189
rect 2764 2137 2816 2189
rect 2828 2137 2880 2189
rect 2892 2137 2944 2189
rect 2973 2186 3025 2238
<< metal2 >>
rect 750 4461 1836 4468
rect 750 4412 838 4461
rect 750 4360 757 4412
rect 809 4409 838 4412
rect 890 4409 902 4461
rect 954 4409 966 4461
rect 1018 4409 1030 4461
rect 1082 4409 1094 4461
rect 1146 4409 1158 4461
rect 1210 4409 1222 4461
rect 1274 4409 1286 4461
rect 1338 4409 1350 4461
rect 1402 4409 1414 4461
rect 1466 4409 1478 4461
rect 1530 4409 1542 4461
rect 1594 4409 1606 4461
rect 1658 4409 1670 4461
rect 1722 4409 1734 4461
rect 1786 4409 1836 4461
rect 809 4402 1836 4409
rect 809 4360 816 4402
rect 1864 4374 1918 4468
rect 1946 4461 3032 4468
rect 1946 4409 1996 4461
rect 2048 4409 2060 4461
rect 2112 4409 2124 4461
rect 2176 4409 2188 4461
rect 2240 4409 2252 4461
rect 2304 4409 2316 4461
rect 2368 4409 2380 4461
rect 2432 4409 2444 4461
rect 2496 4409 2508 4461
rect 2560 4409 2572 4461
rect 2624 4409 2636 4461
rect 2688 4409 2700 4461
rect 2752 4409 2764 4461
rect 2816 4409 2828 4461
rect 2880 4409 2892 4461
rect 2944 4412 3032 4461
rect 2944 4409 2973 4412
rect 1946 4402 2973 4409
rect 750 4348 816 4360
rect 750 4296 757 4348
rect 809 4318 816 4348
rect 844 4367 2938 4374
rect 844 4346 1865 4367
rect 809 4296 1835 4318
rect 750 4290 1835 4296
rect 1863 4315 1865 4346
rect 1917 4346 2938 4367
rect 2966 4360 2973 4402
rect 3025 4360 3032 4412
rect 2966 4348 3032 4360
rect 1917 4315 1919 4346
rect 2966 4318 2973 4348
rect 1863 4303 1919 4315
rect 750 4284 816 4290
rect 750 4232 757 4284
rect 809 4232 816 4284
rect 1863 4262 1865 4303
rect 844 4251 1865 4262
rect 1917 4262 1919 4303
rect 1947 4296 2973 4318
rect 3025 4296 3032 4348
rect 1947 4290 3032 4296
rect 2966 4284 3032 4290
rect 1917 4251 2938 4262
rect 844 4239 2938 4251
rect 844 4234 1865 4239
rect 750 4220 816 4232
rect 750 4168 757 4220
rect 809 4206 816 4220
rect 809 4178 1835 4206
rect 1863 4187 1865 4234
rect 1917 4234 2938 4239
rect 1917 4187 1919 4234
rect 2966 4232 2973 4284
rect 3025 4232 3032 4284
rect 2966 4220 3032 4232
rect 2966 4206 2973 4220
rect 809 4168 816 4178
rect 750 4156 816 4168
rect 750 4104 757 4156
rect 809 4104 816 4156
rect 1863 4175 1919 4187
rect 1947 4178 2973 4206
rect 1863 4150 1865 4175
rect 844 4123 1865 4150
rect 1917 4150 1919 4175
rect 2966 4168 2973 4178
rect 3025 4168 3032 4220
rect 2966 4156 3032 4168
rect 1917 4123 2938 4150
rect 844 4122 2938 4123
rect 750 4094 816 4104
rect 1863 4111 1919 4122
rect 750 4092 1835 4094
rect 750 4040 757 4092
rect 809 4066 1835 4092
rect 809 4040 816 4066
rect 750 4028 816 4040
rect 1863 4059 1865 4111
rect 1917 4059 1919 4111
rect 2966 4104 2973 4156
rect 3025 4104 3032 4156
rect 2966 4094 3032 4104
rect 1947 4092 3032 4094
rect 1947 4066 2973 4092
rect 1863 4047 1919 4059
rect 1863 4038 1865 4047
rect 750 3976 757 4028
rect 809 3982 816 4028
rect 844 4010 1865 4038
rect 1863 3995 1865 4010
rect 1917 4038 1919 4047
rect 2966 4040 2973 4066
rect 3025 4040 3032 4092
rect 1917 4010 2938 4038
rect 2966 4028 3032 4040
rect 1917 3995 1919 4010
rect 1863 3983 1919 3995
rect 809 3976 1835 3982
rect 750 3964 1835 3976
rect 750 3912 757 3964
rect 809 3954 1835 3964
rect 809 3912 816 3954
rect 1863 3931 1865 3983
rect 1917 3931 1919 3983
rect 2966 3982 2973 4028
rect 1947 3976 2973 3982
rect 3025 3976 3032 4028
rect 1947 3964 3032 3976
rect 1947 3954 2973 3964
rect 1863 3926 1919 3931
rect 750 3900 816 3912
rect 750 3848 757 3900
rect 809 3870 816 3900
rect 844 3919 2938 3926
rect 844 3898 1865 3919
rect 809 3848 1835 3870
rect 750 3842 1835 3848
rect 1863 3867 1865 3898
rect 1917 3898 2938 3919
rect 2966 3912 2973 3954
rect 3025 3912 3032 3964
rect 2966 3900 3032 3912
rect 1917 3867 1919 3898
rect 2966 3870 2973 3900
rect 1863 3855 1919 3867
rect 750 3836 816 3842
rect 750 3784 757 3836
rect 809 3784 816 3836
rect 1863 3814 1865 3855
rect 844 3803 1865 3814
rect 1917 3814 1919 3855
rect 1947 3848 2973 3870
rect 3025 3848 3032 3900
rect 1947 3842 3032 3848
rect 2966 3836 3032 3842
rect 1917 3803 2938 3814
rect 844 3791 2938 3803
rect 844 3786 1865 3791
rect 750 3772 816 3784
rect 750 3720 757 3772
rect 809 3758 816 3772
rect 809 3730 1835 3758
rect 1863 3739 1865 3786
rect 1917 3786 2938 3791
rect 1917 3739 1919 3786
rect 2966 3784 2973 3836
rect 3025 3784 3032 3836
rect 2966 3772 3032 3784
rect 2966 3758 2973 3772
rect 809 3720 816 3730
rect 750 3708 816 3720
rect 750 3656 757 3708
rect 809 3656 816 3708
rect 1863 3727 1919 3739
rect 1947 3730 2973 3758
rect 1863 3702 1865 3727
rect 844 3675 1865 3702
rect 1917 3702 1919 3727
rect 2966 3720 2973 3730
rect 3025 3720 3032 3772
rect 2966 3708 3032 3720
rect 1917 3675 2938 3702
rect 844 3674 2938 3675
rect 750 3646 816 3656
rect 1863 3663 1919 3674
rect 750 3644 1835 3646
rect 750 3592 757 3644
rect 809 3618 1835 3644
rect 809 3592 816 3618
rect 750 3580 816 3592
rect 1863 3611 1865 3663
rect 1917 3611 1919 3663
rect 2966 3656 2973 3708
rect 3025 3656 3032 3708
rect 2966 3646 3032 3656
rect 1947 3644 3032 3646
rect 1947 3618 2973 3644
rect 1863 3599 1919 3611
rect 1863 3590 1865 3599
rect 750 3528 757 3580
rect 809 3534 816 3580
rect 844 3562 1865 3590
rect 1863 3547 1865 3562
rect 1917 3590 1919 3599
rect 2966 3592 2973 3618
rect 3025 3592 3032 3644
rect 1917 3562 2938 3590
rect 2966 3580 3032 3592
rect 1917 3547 1919 3562
rect 1863 3535 1919 3547
rect 809 3528 1835 3534
rect 750 3516 1835 3528
rect 750 3464 757 3516
rect 809 3506 1835 3516
rect 809 3464 816 3506
rect 1863 3483 1865 3535
rect 1917 3483 1919 3535
rect 2966 3534 2973 3580
rect 1947 3528 2973 3534
rect 3025 3528 3032 3580
rect 1947 3516 3032 3528
rect 1947 3506 2973 3516
rect 1863 3478 1919 3483
rect 750 3452 816 3464
rect 750 3400 757 3452
rect 809 3422 816 3452
rect 844 3471 2938 3478
rect 844 3450 1865 3471
rect 809 3400 1835 3422
rect 750 3355 1835 3400
rect 1863 3419 1865 3450
rect 1917 3450 2938 3471
rect 2966 3464 2973 3506
rect 3025 3464 3032 3516
rect 2966 3452 3032 3464
rect 1917 3419 1919 3450
rect 2966 3422 2973 3452
rect 1863 3407 1919 3419
rect 1863 3355 1865 3407
rect 1917 3355 1919 3407
rect 1947 3400 2973 3422
rect 3025 3400 3032 3452
rect 1947 3355 3032 3400
rect 750 3354 816 3355
rect 1863 3327 1919 3355
rect 2966 3354 3032 3355
rect 824 3326 2958 3327
rect 750 3325 3032 3326
rect 750 3273 902 3325
rect 954 3273 966 3325
rect 1018 3273 1030 3325
rect 1082 3273 1094 3325
rect 1146 3273 1158 3325
rect 1210 3273 1222 3325
rect 1274 3273 1286 3325
rect 1338 3273 1350 3325
rect 1402 3273 1414 3325
rect 1466 3273 1478 3325
rect 1530 3273 1542 3325
rect 1594 3273 1606 3325
rect 1658 3273 1670 3325
rect 1722 3273 1734 3325
rect 1786 3273 1798 3325
rect 1850 3273 1932 3325
rect 1984 3273 1996 3325
rect 2048 3273 2060 3325
rect 2112 3273 2124 3325
rect 2176 3273 2188 3325
rect 2240 3273 2252 3325
rect 2304 3273 2316 3325
rect 2368 3273 2380 3325
rect 2432 3273 2444 3325
rect 2496 3273 2508 3325
rect 2560 3273 2572 3325
rect 2624 3273 2636 3325
rect 2688 3273 2700 3325
rect 2752 3273 2764 3325
rect 2816 3273 2828 3325
rect 2880 3273 3032 3325
rect 750 3272 3032 3273
rect 824 3271 2958 3272
rect 750 3243 816 3244
rect 1863 3243 1919 3271
rect 2966 3243 3032 3244
rect 750 3198 1835 3243
rect 750 3146 757 3198
rect 809 3176 1835 3198
rect 1863 3191 1865 3243
rect 1917 3191 1919 3243
rect 1863 3179 1919 3191
rect 809 3146 816 3176
rect 1863 3148 1865 3179
rect 750 3134 816 3146
rect 750 3082 757 3134
rect 809 3092 816 3134
rect 844 3127 1865 3148
rect 1917 3148 1919 3179
rect 1947 3198 3032 3243
rect 1947 3176 2973 3198
rect 1917 3127 2938 3148
rect 844 3120 2938 3127
rect 2966 3146 2973 3176
rect 3025 3146 3032 3198
rect 2966 3134 3032 3146
rect 1863 3115 1919 3120
rect 809 3082 1835 3092
rect 750 3070 1835 3082
rect 750 3018 757 3070
rect 809 3064 1835 3070
rect 809 3018 816 3064
rect 1863 3063 1865 3115
rect 1917 3063 1919 3115
rect 2966 3092 2973 3134
rect 1947 3082 2973 3092
rect 3025 3082 3032 3134
rect 1947 3070 3032 3082
rect 1947 3064 2973 3070
rect 1863 3051 1919 3063
rect 1863 3036 1865 3051
rect 750 3006 816 3018
rect 844 3008 1865 3036
rect 750 2954 757 3006
rect 809 2980 816 3006
rect 1863 2999 1865 3008
rect 1917 3036 1919 3051
rect 1917 3008 2938 3036
rect 2966 3018 2973 3064
rect 3025 3018 3032 3070
rect 1917 2999 1919 3008
rect 1863 2987 1919 2999
rect 809 2954 1835 2980
rect 750 2952 1835 2954
rect 750 2942 816 2952
rect 750 2890 757 2942
rect 809 2890 816 2942
rect 1863 2935 1865 2987
rect 1917 2935 1919 2987
rect 2966 3006 3032 3018
rect 2966 2980 2973 3006
rect 1947 2954 2973 2980
rect 3025 2954 3032 3006
rect 1947 2952 3032 2954
rect 1863 2924 1919 2935
rect 2966 2942 3032 2952
rect 844 2923 2938 2924
rect 844 2896 1865 2923
rect 750 2878 816 2890
rect 750 2826 757 2878
rect 809 2868 816 2878
rect 1863 2871 1865 2896
rect 1917 2896 2938 2923
rect 1917 2871 1919 2896
rect 809 2840 1835 2868
rect 1863 2859 1919 2871
rect 2966 2890 2973 2942
rect 3025 2890 3032 2942
rect 2966 2878 3032 2890
rect 2966 2868 2973 2878
rect 809 2826 816 2840
rect 750 2814 816 2826
rect 750 2762 757 2814
rect 809 2762 816 2814
rect 1863 2812 1865 2859
rect 844 2807 1865 2812
rect 1917 2812 1919 2859
rect 1947 2840 2973 2868
rect 2966 2826 2973 2840
rect 3025 2826 3032 2878
rect 2966 2814 3032 2826
rect 1917 2807 2938 2812
rect 844 2795 2938 2807
rect 844 2784 1865 2795
rect 750 2756 816 2762
rect 750 2750 1835 2756
rect 750 2698 757 2750
rect 809 2728 1835 2750
rect 1863 2743 1865 2784
rect 1917 2784 2938 2795
rect 1917 2743 1919 2784
rect 2966 2762 2973 2814
rect 3025 2762 3032 2814
rect 2966 2756 3032 2762
rect 1863 2731 1919 2743
rect 809 2698 816 2728
rect 1863 2700 1865 2731
rect 750 2686 816 2698
rect 750 2634 757 2686
rect 809 2644 816 2686
rect 844 2679 1865 2700
rect 1917 2700 1919 2731
rect 1947 2750 3032 2756
rect 1947 2728 2973 2750
rect 1917 2679 2938 2700
rect 844 2672 2938 2679
rect 2966 2698 2973 2728
rect 3025 2698 3032 2750
rect 2966 2686 3032 2698
rect 1863 2667 1919 2672
rect 809 2634 1835 2644
rect 750 2622 1835 2634
rect 750 2570 757 2622
rect 809 2616 1835 2622
rect 809 2570 816 2616
rect 1863 2615 1865 2667
rect 1917 2615 1919 2667
rect 2966 2644 2973 2686
rect 1947 2634 2973 2644
rect 3025 2634 3032 2686
rect 1947 2622 3032 2634
rect 1947 2616 2973 2622
rect 1863 2603 1919 2615
rect 1863 2588 1865 2603
rect 750 2558 816 2570
rect 844 2560 1865 2588
rect 750 2506 757 2558
rect 809 2532 816 2558
rect 1863 2551 1865 2560
rect 1917 2588 1919 2603
rect 1917 2560 2938 2588
rect 2966 2570 2973 2616
rect 3025 2570 3032 2622
rect 1917 2551 1919 2560
rect 1863 2539 1919 2551
rect 809 2506 1835 2532
rect 750 2504 1835 2506
rect 750 2494 816 2504
rect 750 2442 757 2494
rect 809 2442 816 2494
rect 1863 2487 1865 2539
rect 1917 2487 1919 2539
rect 2966 2558 3032 2570
rect 2966 2532 2973 2558
rect 1947 2506 2973 2532
rect 3025 2506 3032 2558
rect 1947 2504 3032 2506
rect 1863 2476 1919 2487
rect 2966 2494 3032 2504
rect 844 2475 2938 2476
rect 844 2448 1865 2475
rect 750 2430 816 2442
rect 750 2378 757 2430
rect 809 2420 816 2430
rect 1863 2423 1865 2448
rect 1917 2448 2938 2475
rect 1917 2423 1919 2448
rect 809 2392 1835 2420
rect 1863 2411 1919 2423
rect 2966 2442 2973 2494
rect 3025 2442 3032 2494
rect 2966 2430 3032 2442
rect 2966 2420 2973 2430
rect 809 2378 816 2392
rect 750 2366 816 2378
rect 750 2314 757 2366
rect 809 2314 816 2366
rect 1863 2364 1865 2411
rect 844 2359 1865 2364
rect 1917 2364 1919 2411
rect 1947 2392 2973 2420
rect 2966 2378 2973 2392
rect 3025 2378 3032 2430
rect 2966 2366 3032 2378
rect 1917 2359 2938 2364
rect 844 2347 2938 2359
rect 844 2336 1865 2347
rect 750 2308 816 2314
rect 750 2302 1835 2308
rect 750 2250 757 2302
rect 809 2280 1835 2302
rect 1863 2295 1865 2336
rect 1917 2336 2938 2347
rect 1917 2295 1919 2336
rect 2966 2314 2973 2366
rect 3025 2314 3032 2366
rect 2966 2308 3032 2314
rect 1863 2283 1919 2295
rect 809 2250 816 2280
rect 1863 2252 1865 2283
rect 750 2238 816 2250
rect 750 2186 757 2238
rect 809 2196 816 2238
rect 844 2231 1865 2252
rect 1917 2252 1919 2283
rect 1947 2302 3032 2308
rect 1947 2280 2973 2302
rect 1917 2231 2938 2252
rect 844 2224 2938 2231
rect 2966 2250 2973 2280
rect 3025 2250 3032 2302
rect 2966 2238 3032 2250
rect 809 2189 1836 2196
rect 809 2186 838 2189
rect 750 2137 838 2186
rect 890 2137 902 2189
rect 954 2137 966 2189
rect 1018 2137 1030 2189
rect 1082 2137 1094 2189
rect 1146 2137 1158 2189
rect 1210 2137 1222 2189
rect 1274 2137 1286 2189
rect 1338 2137 1350 2189
rect 1402 2137 1414 2189
rect 1466 2137 1478 2189
rect 1530 2137 1542 2189
rect 1594 2137 1606 2189
rect 1658 2137 1670 2189
rect 1722 2137 1734 2189
rect 1786 2137 1836 2189
rect 750 2130 1836 2137
rect 1864 2130 1918 2224
rect 2966 2196 2973 2238
rect 1946 2189 2973 2196
rect 1946 2137 1996 2189
rect 2048 2137 2060 2189
rect 2112 2137 2124 2189
rect 2176 2137 2188 2189
rect 2240 2137 2252 2189
rect 2304 2137 2316 2189
rect 2368 2137 2380 2189
rect 2432 2137 2444 2189
rect 2496 2137 2508 2189
rect 2560 2137 2572 2189
rect 2624 2137 2636 2189
rect 2688 2137 2700 2189
rect 2752 2137 2764 2189
rect 2816 2137 2828 2189
rect 2880 2137 2892 2189
rect 2944 2186 2973 2189
rect 3025 2186 3032 2238
rect 2944 2137 3032 2186
rect 1946 2130 3032 2137
<< labels >>
flabel metal2 1769 4292 1799 4314 0 FreeSans 200 0 0 0 sky130_fd_pr__cap_vpp_11p5x11p7_m1m2_noshield_0.C0
flabel metal2 1871 4192 1913 4228 0 FreeSans 200 0 0 0 sky130_fd_pr__cap_vpp_11p5x11p7_m1m2_noshield_0.C1
flabel pwell 1926 3419 1947 3468 0 FreeSans 1600 0 0 0 sky130_fd_pr__cap_vpp_11p5x11p7_m1m2_noshield_0.SUB
<< end >>
